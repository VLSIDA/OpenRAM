**************************************************
* OpenRAM generated memory.
* Words: 1024
* Data bits: 128
* Banks: 2
* Column mux: 2:1
**************************************************

* ptx M{0} {1} n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p

* ptx M{0} {1} p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p

.SUBCKT pnand2_1 A B Z vdd gnd
Mpnand2_pmos1 vdd A Z vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand2_pmos2 Z B vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand2_nmos1 Z B net1 gnd n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand2_nmos2 net1 A gnd gnd n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
.ENDS pnand2_1

.SUBCKT pnand3_1 A B C Z vdd gnd
Mpnand3_pmos1 vdd A Z vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand3_pmos2 Z B vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand3_pmos3 Z C vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand3_nmos1 Z C net1 gnd n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand3_nmos2 net1 B net2 gnd n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand3_nmos3 net2 A gnd gnd n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
.ENDS pnand3_1

* ptx M{0} {1} n m=1 w=1.2u l=0.6u pd=3.6u ps=3.6u as=1.8p ad=1.8p

* ptx M{0} {1} p m=1 w=3.6u l=0.6u pd=8.4u ps=8.4u as=5.4p ad=5.4p

.SUBCKT pnor2_1 A B Z vdd gnd
Mpnor2_pmos1 vdd A net1 vdd p m=1 w=3.6u l=0.6u pd=8.4u ps=8.4u as=5.4p ad=5.4p
Mpnor2_pmos2 net1 B Z vdd p m=1 w=3.6u l=0.6u pd=8.4u ps=8.4u as=5.4p ad=5.4p
Mpnor2_nmos1 Z A gnd gnd n m=1 w=1.2u l=0.6u pd=3.6u ps=3.6u as=1.8p ad=1.8p
Mpnor2_nmos2 Z B gnd gnd n m=1 w=1.2u l=0.6u pd=3.6u ps=3.6u as=1.8p ad=1.8p
.ENDS pnor2_1

.SUBCKT pinv_1 A Z vdd gnd
Mpinv_pmos Z A vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpinv_nmos Z A gnd gnd n m=1 w=1.2u l=0.6u pd=3.6u ps=3.6u as=1.8p ad=1.8p
.ENDS pinv_1

* ptx M{0} {1} n m=2 w=1.2u l=0.6u pd=3.6u ps=3.6u as=1.8p ad=1.8p

* ptx M{0} {1} p m=2 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p

.SUBCKT pinv_2 A Z vdd gnd
Mpinv_pmos Z A vdd vdd p m=2 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpinv_nmos Z A gnd gnd n m=2 w=1.2u l=0.6u pd=3.6u ps=3.6u as=1.8p ad=1.8p
.ENDS pinv_2

* ptx M{0} {1} n m=3 w=1.65u l=0.6u pd=4.5u ps=4.5u as=2.475p ad=2.475p

* ptx M{0} {1} p m=3 w=3.15u l=0.6u pd=7.5u ps=7.5u as=4.725p ad=4.725p

.SUBCKT pinv_3 A Z vdd gnd
Mpinv_pmos Z A vdd vdd p m=3 w=3.15u l=0.6u pd=7.5u ps=7.5u as=4.725p ad=4.725p
Mpinv_nmos Z A gnd gnd n m=3 w=1.65u l=0.6u pd=4.5u ps=4.5u as=2.475p ad=2.475p
.ENDS pinv_3

* ptx M{0} {1} n m=5 w=1.95u l=0.6u pd=5.1u ps=5.1u as=2.925p ad=2.925p

* ptx M{0} {1} p m=5 w=3.9u l=0.6u pd=9.0u ps=9.0u as=5.85p ad=5.85p

.SUBCKT pinv_4 A Z vdd gnd
Mpinv_pmos Z A vdd vdd p m=5 w=3.9u l=0.6u pd=9.0u ps=9.0u as=5.85p ad=5.85p
Mpinv_nmos Z A gnd gnd n m=5 w=1.95u l=0.6u pd=5.1u ps=5.1u as=2.925p ad=2.925p
.ENDS pinv_4

* ptx M{0} {1} n m=10 w=1.95u l=0.6u pd=5.1u ps=5.1u as=2.925p ad=2.925p

* ptx M{0} {1} p m=10 w=3.9u l=0.6u pd=9.0u ps=9.0u as=5.85p ad=5.85p

.SUBCKT pinv_5 A Z vdd gnd
Mpinv_pmos Z A vdd vdd p m=10 w=3.9u l=0.6u pd=9.0u ps=9.0u as=5.85p ad=5.85p
Mpinv_nmos Z A gnd gnd n m=10 w=1.95u l=0.6u pd=5.1u ps=5.1u as=2.925p ad=2.925p
.ENDS pinv_5
*master-slave flip-flop with both output and inverted ouput

.subckt ms_flop din dout dout_bar clk vdd gnd
xmaster din mout mout_bar clk clk_bar vdd gnd dlatch
xslave mout_bar dout_bar dout clk_bar clk_nn vdd gnd dlatch
.ends flop

.subckt dlatch din dout dout_bar clk clk_bar vdd gnd
*clk inverter
mPff1 clk_bar clk vdd vdd p W=1.8u L=0.6u m=1
mNff1 clk_bar clk gnd gnd n W=0.9u L=0.6u m=1

*transmission gate 1
mtmP1 din clk int1 vdd p W=1.8u L=0.6u m=1
mtmN1 din clk_bar int1 gnd n W=0.9u L=0.6u m=1

*foward inverter
mPff3 dout_bar int1 vdd vdd p W=1.8u L=0.6u m=1
mNff3 dout_bar int1 gnd gnd n W=0.9u L=0.6u m=1

*backward inverter
mPff4 dout dout_bar vdd vdd p W=1.8u L=0.6u m=1
mNf4 dout dout_bar gnd gnd n W=0.9u L=0.6u m=1

*transmission gate 2
mtmP2 int1 clk_bar dout vdd p W=1.8u L=0.6u m=1
mtmN2 int1 clk dout gnd n W=0.9u L=0.6u m=1
.ends dlatch


.SUBCKT msf_control din[0] din[1] din[2] dout[0] dout_bar[0] dout[1] dout_bar[1] dout[2] dout_bar[2] clk vdd gnd
XXdff0 din[0] dout[0] dout_bar[0] clk vdd gnd ms_flop
XXdff1 din[1] dout[1] dout_bar[1] clk vdd gnd ms_flop
XXdff2 din[2] dout[2] dout_bar[2] clk vdd gnd ms_flop
.ENDS msf_control

*********************** "cell_6t" ******************************
.SUBCKT replica_cell_6t bl br wl vdd gnd
M_1 gnd net_2 vdd vdd p W='0.9u' L=1.2u
M_2 net_2 gnd vdd vdd p W='0.9u' L=1.2u
M_3 br wl net_2 gnd n W='1.2u' L=0.6u
M_4 bl wl gnd gnd n W='1.2u' L=0.6u
M_5 net_2 gnd gnd gnd n W='2.4u' L=0.6u
M_6 gnd net_2 gnd gnd n W='2.4u' L=0.6u
.ENDS	$ replica_cell_6t

*********************** "cell_6t" ******************************
.SUBCKT cell_6t bl br wl vdd gnd
M_1 net_1 net_2 vdd vdd p W='0.9u' L=1.2u
M_2 net_2 net_1 vdd vdd p W='0.9u' L=1.2u
M_3 br wl net_2 gnd n W='1.2u' L=0.6u
M_4 bl wl net_1 gnd n W='1.2u' L=0.6u
M_5 net_2 net_1 gnd gnd n W='2.4u' L=0.6u
M_6 net_1 net_2 gnd gnd n W='2.4u' L=0.6u
.ENDS	$ cell_6t

.SUBCKT bitline_load bl[0] br[0] wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] vdd gnd
Xbit_r0_c0 bl[0] br[0] wl[0] vdd gnd cell_6t
Xbit_r1_c0 bl[0] br[0] wl[1] vdd gnd cell_6t
Xbit_r2_c0 bl[0] br[0] wl[2] vdd gnd cell_6t
Xbit_r3_c0 bl[0] br[0] wl[3] vdd gnd cell_6t
Xbit_r4_c0 bl[0] br[0] wl[4] vdd gnd cell_6t
Xbit_r5_c0 bl[0] br[0] wl[5] vdd gnd cell_6t
Xbit_r6_c0 bl[0] br[0] wl[6] vdd gnd cell_6t
Xbit_r7_c0 bl[0] br[0] wl[7] vdd gnd cell_6t
Xbit_r8_c0 bl[0] br[0] wl[8] vdd gnd cell_6t
Xbit_r9_c0 bl[0] br[0] wl[9] vdd gnd cell_6t
Xbit_r10_c0 bl[0] br[0] wl[10] vdd gnd cell_6t
Xbit_r11_c0 bl[0] br[0] wl[11] vdd gnd cell_6t
Xbit_r12_c0 bl[0] br[0] wl[12] vdd gnd cell_6t
Xbit_r13_c0 bl[0] br[0] wl[13] vdd gnd cell_6t
Xbit_r14_c0 bl[0] br[0] wl[14] vdd gnd cell_6t
Xbit_r15_c0 bl[0] br[0] wl[15] vdd gnd cell_6t
Xbit_r16_c0 bl[0] br[0] wl[16] vdd gnd cell_6t
Xbit_r17_c0 bl[0] br[0] wl[17] vdd gnd cell_6t
Xbit_r18_c0 bl[0] br[0] wl[18] vdd gnd cell_6t
Xbit_r19_c0 bl[0] br[0] wl[19] vdd gnd cell_6t
Xbit_r20_c0 bl[0] br[0] wl[20] vdd gnd cell_6t
Xbit_r21_c0 bl[0] br[0] wl[21] vdd gnd cell_6t
Xbit_r22_c0 bl[0] br[0] wl[22] vdd gnd cell_6t
Xbit_r23_c0 bl[0] br[0] wl[23] vdd gnd cell_6t
Xbit_r24_c0 bl[0] br[0] wl[24] vdd gnd cell_6t
Xbit_r25_c0 bl[0] br[0] wl[25] vdd gnd cell_6t
Xbit_r26_c0 bl[0] br[0] wl[26] vdd gnd cell_6t
Xbit_r27_c0 bl[0] br[0] wl[27] vdd gnd cell_6t
Xbit_r28_c0 bl[0] br[0] wl[28] vdd gnd cell_6t
Xbit_r29_c0 bl[0] br[0] wl[29] vdd gnd cell_6t
Xbit_r30_c0 bl[0] br[0] wl[30] vdd gnd cell_6t
Xbit_r31_c0 bl[0] br[0] wl[31] vdd gnd cell_6t
Xbit_r32_c0 bl[0] br[0] wl[32] vdd gnd cell_6t
Xbit_r33_c0 bl[0] br[0] wl[33] vdd gnd cell_6t
Xbit_r34_c0 bl[0] br[0] wl[34] vdd gnd cell_6t
Xbit_r35_c0 bl[0] br[0] wl[35] vdd gnd cell_6t
Xbit_r36_c0 bl[0] br[0] wl[36] vdd gnd cell_6t
Xbit_r37_c0 bl[0] br[0] wl[37] vdd gnd cell_6t
Xbit_r38_c0 bl[0] br[0] wl[38] vdd gnd cell_6t
Xbit_r39_c0 bl[0] br[0] wl[39] vdd gnd cell_6t
Xbit_r40_c0 bl[0] br[0] wl[40] vdd gnd cell_6t
Xbit_r41_c0 bl[0] br[0] wl[41] vdd gnd cell_6t
Xbit_r42_c0 bl[0] br[0] wl[42] vdd gnd cell_6t
Xbit_r43_c0 bl[0] br[0] wl[43] vdd gnd cell_6t
Xbit_r44_c0 bl[0] br[0] wl[44] vdd gnd cell_6t
Xbit_r45_c0 bl[0] br[0] wl[45] vdd gnd cell_6t
Xbit_r46_c0 bl[0] br[0] wl[46] vdd gnd cell_6t
Xbit_r47_c0 bl[0] br[0] wl[47] vdd gnd cell_6t
Xbit_r48_c0 bl[0] br[0] wl[48] vdd gnd cell_6t
Xbit_r49_c0 bl[0] br[0] wl[49] vdd gnd cell_6t
Xbit_r50_c0 bl[0] br[0] wl[50] vdd gnd cell_6t
Xbit_r51_c0 bl[0] br[0] wl[51] vdd gnd cell_6t
.ENDS bitline_load

.SUBCKT pinv_6 A Z vdd gnd
Mpinv_pmos Z A vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpinv_nmos Z A gnd gnd n m=1 w=1.2u l=0.6u pd=3.6u ps=3.6u as=1.8p ad=1.8p
.ENDS pinv_6

.SUBCKT delay_chain in out vdd gnd
Xdinv0 in s1 vdd gnd pinv_6
Xdinv1 s1 s2n1 vdd gnd pinv_6
Xdinv2 s1 s2n2 vdd gnd pinv_6
Xdinv3 s1 s2 vdd gnd pinv_6
Xdinv4 s2 s3n1 vdd gnd pinv_6
Xdinv5 s2 s3n2 vdd gnd pinv_6
Xdinv6 s2 s3 vdd gnd pinv_6
Xdinv7 s3 s4n1 vdd gnd pinv_6
Xdinv8 s3 s4n2 vdd gnd pinv_6
Xdinv9 s3 s4 vdd gnd pinv_6
Xdinv10 s4 s5n1 vdd gnd pinv_6
Xdinv11 s4 s5n2 vdd gnd pinv_6
Xdinv12 s4 out vdd gnd pinv_6
.ENDS delay_chain

.SUBCKT pinv_7 A Z vdd gnd
Mpinv_pmos Z A vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpinv_nmos Z A gnd gnd n m=1 w=1.2u l=0.6u pd=3.6u ps=3.6u as=1.8p ad=1.8p
.ENDS pinv_7

* ptx M{0} {1} p m=1 w=1.2u l=0.6u pd=3.6u ps=3.6u as=1.8p ad=1.8p

.SUBCKT replica_bitline en out vdd gnd
Xrbl_inv bl[0] out vdd gnd pinv_7
Mrbl_access_tx vdd delayed_en bl[0] vdd p m=1 w=1.2u l=0.6u pd=3.6u ps=3.6u as=1.8p ad=1.8p
Xdelay_chain en delayed_en vdd gnd delay_chain
Xbitcell bl[0] br[0] delayed_en vdd gnd replica_cell_6t
Xload bl[0] br[0] gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd vdd gnd bitline_load
.ENDS replica_bitline

.SUBCKT control_logic csb web oeb clk s_en w_en tri_en tri_en_bar clk_bar clk_buf vdd gnd
Xmsf_control oeb csb web oe_bar oe cs_bar cs we_bar we clk_buf vdd gnd msf_control
Xinv_clk1_bar clk clk1_bar vdd gnd pinv_2
Xinv_clk2 clk1_bar clk2 vdd gnd pinv_3
Xinv_clk_bar clk2 clk_bar vdd gnd pinv_4
Xinv_clk_buf clk_bar clk_buf vdd gnd pinv_5
Xnand3_rblk_bar clk_bar oe cs rblk_bar vdd gnd pnand3_1
Xinv_rblk rblk_bar rblk vdd gnd pinv_1
Xnor2_tri_en clk_buf oe_bar tri_en vdd gnd pnor2_1
Xnand2_tri_en clk_bar oe tri_en_bar vdd gnd pnand2_1
Xinv_s_en pre_s_en_bar s_en vdd gnd pinv_1
Xinv_pre_s_en_bar pre_s_en pre_s_en_bar vdd gnd pinv_1
Xnand3_w_en_bar clk_bar cs we w_en_bar vdd gnd pnand3_1
Xinv_pre_w_en w_en_bar pre_w_en vdd gnd pinv_1
Xinv_pre_w_en_bar pre_w_en pre_w_en_bar vdd gnd pinv_1
Xinv_w_en2 pre_w_en_bar w_en vdd gnd pinv_1
Xreplica_bitline rblk pre_s_en vdd gnd replica_bitline
.ENDS control_logic

.SUBCKT bitcell_array bl[0] br[0] bl[1] br[1] bl[2] br[2] bl[3] br[3] bl[4] br[4] bl[5] br[5] bl[6] br[6] bl[7] br[7] bl[8] br[8] bl[9] br[9] bl[10] br[10] bl[11] br[11] bl[12] br[12] bl[13] br[13] bl[14] br[14] bl[15] br[15] bl[16] br[16] bl[17] br[17] bl[18] br[18] bl[19] br[19] bl[20] br[20] bl[21] br[21] bl[22] br[22] bl[23] br[23] bl[24] br[24] bl[25] br[25] bl[26] br[26] bl[27] br[27] bl[28] br[28] bl[29] br[29] bl[30] br[30] bl[31] br[31] bl[32] br[32] bl[33] br[33] bl[34] br[34] bl[35] br[35] bl[36] br[36] bl[37] br[37] bl[38] br[38] bl[39] br[39] bl[40] br[40] bl[41] br[41] bl[42] br[42] bl[43] br[43] bl[44] br[44] bl[45] br[45] bl[46] br[46] bl[47] br[47] bl[48] br[48] bl[49] br[49] bl[50] br[50] bl[51] br[51] bl[52] br[52] bl[53] br[53] bl[54] br[54] bl[55] br[55] bl[56] br[56] bl[57] br[57] bl[58] br[58] bl[59] br[59] bl[60] br[60] bl[61] br[61] bl[62] br[62] bl[63] br[63] bl[64] br[64] bl[65] br[65] bl[66] br[66] bl[67] br[67] bl[68] br[68] bl[69] br[69] bl[70] br[70] bl[71] br[71] bl[72] br[72] bl[73] br[73] bl[74] br[74] bl[75] br[75] bl[76] br[76] bl[77] br[77] bl[78] br[78] bl[79] br[79] bl[80] br[80] bl[81] br[81] bl[82] br[82] bl[83] br[83] bl[84] br[84] bl[85] br[85] bl[86] br[86] bl[87] br[87] bl[88] br[88] bl[89] br[89] bl[90] br[90] bl[91] br[91] bl[92] br[92] bl[93] br[93] bl[94] br[94] bl[95] br[95] bl[96] br[96] bl[97] br[97] bl[98] br[98] bl[99] br[99] bl[100] br[100] bl[101] br[101] bl[102] br[102] bl[103] br[103] bl[104] br[104] bl[105] br[105] bl[106] br[106] bl[107] br[107] bl[108] br[108] bl[109] br[109] bl[110] br[110] bl[111] br[111] bl[112] br[112] bl[113] br[113] bl[114] br[114] bl[115] br[115] bl[116] br[116] bl[117] br[117] bl[118] br[118] bl[119] br[119] bl[120] br[120] bl[121] br[121] bl[122] br[122] bl[123] br[123] bl[124] br[124] bl[125] br[125] bl[126] br[126] bl[127] br[127] bl[128] br[128] bl[129] br[129] bl[130] br[130] bl[131] br[131] bl[132] br[132] bl[133] br[133] bl[134] br[134] bl[135] br[135] bl[136] br[136] bl[137] br[137] bl[138] br[138] bl[139] br[139] bl[140] br[140] bl[141] br[141] bl[142] br[142] bl[143] br[143] bl[144] br[144] bl[145] br[145] bl[146] br[146] bl[147] br[147] bl[148] br[148] bl[149] br[149] bl[150] br[150] bl[151] br[151] bl[152] br[152] bl[153] br[153] bl[154] br[154] bl[155] br[155] bl[156] br[156] bl[157] br[157] bl[158] br[158] bl[159] br[159] bl[160] br[160] bl[161] br[161] bl[162] br[162] bl[163] br[163] bl[164] br[164] bl[165] br[165] bl[166] br[166] bl[167] br[167] bl[168] br[168] bl[169] br[169] bl[170] br[170] bl[171] br[171] bl[172] br[172] bl[173] br[173] bl[174] br[174] bl[175] br[175] bl[176] br[176] bl[177] br[177] bl[178] br[178] bl[179] br[179] bl[180] br[180] bl[181] br[181] bl[182] br[182] bl[183] br[183] bl[184] br[184] bl[185] br[185] bl[186] br[186] bl[187] br[187] bl[188] br[188] bl[189] br[189] bl[190] br[190] bl[191] br[191] bl[192] br[192] bl[193] br[193] bl[194] br[194] bl[195] br[195] bl[196] br[196] bl[197] br[197] bl[198] br[198] bl[199] br[199] bl[200] br[200] bl[201] br[201] bl[202] br[202] bl[203] br[203] bl[204] br[204] bl[205] br[205] bl[206] br[206] bl[207] br[207] bl[208] br[208] bl[209] br[209] bl[210] br[210] bl[211] br[211] bl[212] br[212] bl[213] br[213] bl[214] br[214] bl[215] br[215] bl[216] br[216] bl[217] br[217] bl[218] br[218] bl[219] br[219] bl[220] br[220] bl[221] br[221] bl[222] br[222] bl[223] br[223] bl[224] br[224] bl[225] br[225] bl[226] br[226] bl[227] br[227] bl[228] br[228] bl[229] br[229] bl[230] br[230] bl[231] br[231] bl[232] br[232] bl[233] br[233] bl[234] br[234] bl[235] br[235] bl[236] br[236] bl[237] br[237] bl[238] br[238] bl[239] br[239] bl[240] br[240] bl[241] br[241] bl[242] br[242] bl[243] br[243] bl[244] br[244] bl[245] br[245] bl[246] br[246] bl[247] br[247] bl[248] br[248] bl[249] br[249] bl[250] br[250] bl[251] br[251] bl[252] br[252] bl[253] br[253] bl[254] br[254] bl[255] br[255] wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] wl[128] wl[129] wl[130] wl[131] wl[132] wl[133] wl[134] wl[135] wl[136] wl[137] wl[138] wl[139] wl[140] wl[141] wl[142] wl[143] wl[144] wl[145] wl[146] wl[147] wl[148] wl[149] wl[150] wl[151] wl[152] wl[153] wl[154] wl[155] wl[156] wl[157] wl[158] wl[159] wl[160] wl[161] wl[162] wl[163] wl[164] wl[165] wl[166] wl[167] wl[168] wl[169] wl[170] wl[171] wl[172] wl[173] wl[174] wl[175] wl[176] wl[177] wl[178] wl[179] wl[180] wl[181] wl[182] wl[183] wl[184] wl[185] wl[186] wl[187] wl[188] wl[189] wl[190] wl[191] wl[192] wl[193] wl[194] wl[195] wl[196] wl[197] wl[198] wl[199] wl[200] wl[201] wl[202] wl[203] wl[204] wl[205] wl[206] wl[207] wl[208] wl[209] wl[210] wl[211] wl[212] wl[213] wl[214] wl[215] wl[216] wl[217] wl[218] wl[219] wl[220] wl[221] wl[222] wl[223] wl[224] wl[225] wl[226] wl[227] wl[228] wl[229] wl[230] wl[231] wl[232] wl[233] wl[234] wl[235] wl[236] wl[237] wl[238] wl[239] wl[240] wl[241] wl[242] wl[243] wl[244] wl[245] wl[246] wl[247] wl[248] wl[249] wl[250] wl[251] wl[252] wl[253] wl[254] wl[255] vdd gnd
Xbit_r0_c0 bl[0] br[0] wl[0] vdd gnd cell_6t
Xbit_r1_c0 bl[0] br[0] wl[1] vdd gnd cell_6t
Xbit_r2_c0 bl[0] br[0] wl[2] vdd gnd cell_6t
Xbit_r3_c0 bl[0] br[0] wl[3] vdd gnd cell_6t
Xbit_r4_c0 bl[0] br[0] wl[4] vdd gnd cell_6t
Xbit_r5_c0 bl[0] br[0] wl[5] vdd gnd cell_6t
Xbit_r6_c0 bl[0] br[0] wl[6] vdd gnd cell_6t
Xbit_r7_c0 bl[0] br[0] wl[7] vdd gnd cell_6t
Xbit_r8_c0 bl[0] br[0] wl[8] vdd gnd cell_6t
Xbit_r9_c0 bl[0] br[0] wl[9] vdd gnd cell_6t
Xbit_r10_c0 bl[0] br[0] wl[10] vdd gnd cell_6t
Xbit_r11_c0 bl[0] br[0] wl[11] vdd gnd cell_6t
Xbit_r12_c0 bl[0] br[0] wl[12] vdd gnd cell_6t
Xbit_r13_c0 bl[0] br[0] wl[13] vdd gnd cell_6t
Xbit_r14_c0 bl[0] br[0] wl[14] vdd gnd cell_6t
Xbit_r15_c0 bl[0] br[0] wl[15] vdd gnd cell_6t
Xbit_r16_c0 bl[0] br[0] wl[16] vdd gnd cell_6t
Xbit_r17_c0 bl[0] br[0] wl[17] vdd gnd cell_6t
Xbit_r18_c0 bl[0] br[0] wl[18] vdd gnd cell_6t
Xbit_r19_c0 bl[0] br[0] wl[19] vdd gnd cell_6t
Xbit_r20_c0 bl[0] br[0] wl[20] vdd gnd cell_6t
Xbit_r21_c0 bl[0] br[0] wl[21] vdd gnd cell_6t
Xbit_r22_c0 bl[0] br[0] wl[22] vdd gnd cell_6t
Xbit_r23_c0 bl[0] br[0] wl[23] vdd gnd cell_6t
Xbit_r24_c0 bl[0] br[0] wl[24] vdd gnd cell_6t
Xbit_r25_c0 bl[0] br[0] wl[25] vdd gnd cell_6t
Xbit_r26_c0 bl[0] br[0] wl[26] vdd gnd cell_6t
Xbit_r27_c0 bl[0] br[0] wl[27] vdd gnd cell_6t
Xbit_r28_c0 bl[0] br[0] wl[28] vdd gnd cell_6t
Xbit_r29_c0 bl[0] br[0] wl[29] vdd gnd cell_6t
Xbit_r30_c0 bl[0] br[0] wl[30] vdd gnd cell_6t
Xbit_r31_c0 bl[0] br[0] wl[31] vdd gnd cell_6t
Xbit_r32_c0 bl[0] br[0] wl[32] vdd gnd cell_6t
Xbit_r33_c0 bl[0] br[0] wl[33] vdd gnd cell_6t
Xbit_r34_c0 bl[0] br[0] wl[34] vdd gnd cell_6t
Xbit_r35_c0 bl[0] br[0] wl[35] vdd gnd cell_6t
Xbit_r36_c0 bl[0] br[0] wl[36] vdd gnd cell_6t
Xbit_r37_c0 bl[0] br[0] wl[37] vdd gnd cell_6t
Xbit_r38_c0 bl[0] br[0] wl[38] vdd gnd cell_6t
Xbit_r39_c0 bl[0] br[0] wl[39] vdd gnd cell_6t
Xbit_r40_c0 bl[0] br[0] wl[40] vdd gnd cell_6t
Xbit_r41_c0 bl[0] br[0] wl[41] vdd gnd cell_6t
Xbit_r42_c0 bl[0] br[0] wl[42] vdd gnd cell_6t
Xbit_r43_c0 bl[0] br[0] wl[43] vdd gnd cell_6t
Xbit_r44_c0 bl[0] br[0] wl[44] vdd gnd cell_6t
Xbit_r45_c0 bl[0] br[0] wl[45] vdd gnd cell_6t
Xbit_r46_c0 bl[0] br[0] wl[46] vdd gnd cell_6t
Xbit_r47_c0 bl[0] br[0] wl[47] vdd gnd cell_6t
Xbit_r48_c0 bl[0] br[0] wl[48] vdd gnd cell_6t
Xbit_r49_c0 bl[0] br[0] wl[49] vdd gnd cell_6t
Xbit_r50_c0 bl[0] br[0] wl[50] vdd gnd cell_6t
Xbit_r51_c0 bl[0] br[0] wl[51] vdd gnd cell_6t
Xbit_r52_c0 bl[0] br[0] wl[52] vdd gnd cell_6t
Xbit_r53_c0 bl[0] br[0] wl[53] vdd gnd cell_6t
Xbit_r54_c0 bl[0] br[0] wl[54] vdd gnd cell_6t
Xbit_r55_c0 bl[0] br[0] wl[55] vdd gnd cell_6t
Xbit_r56_c0 bl[0] br[0] wl[56] vdd gnd cell_6t
Xbit_r57_c0 bl[0] br[0] wl[57] vdd gnd cell_6t
Xbit_r58_c0 bl[0] br[0] wl[58] vdd gnd cell_6t
Xbit_r59_c0 bl[0] br[0] wl[59] vdd gnd cell_6t
Xbit_r60_c0 bl[0] br[0] wl[60] vdd gnd cell_6t
Xbit_r61_c0 bl[0] br[0] wl[61] vdd gnd cell_6t
Xbit_r62_c0 bl[0] br[0] wl[62] vdd gnd cell_6t
Xbit_r63_c0 bl[0] br[0] wl[63] vdd gnd cell_6t
Xbit_r64_c0 bl[0] br[0] wl[64] vdd gnd cell_6t
Xbit_r65_c0 bl[0] br[0] wl[65] vdd gnd cell_6t
Xbit_r66_c0 bl[0] br[0] wl[66] vdd gnd cell_6t
Xbit_r67_c0 bl[0] br[0] wl[67] vdd gnd cell_6t
Xbit_r68_c0 bl[0] br[0] wl[68] vdd gnd cell_6t
Xbit_r69_c0 bl[0] br[0] wl[69] vdd gnd cell_6t
Xbit_r70_c0 bl[0] br[0] wl[70] vdd gnd cell_6t
Xbit_r71_c0 bl[0] br[0] wl[71] vdd gnd cell_6t
Xbit_r72_c0 bl[0] br[0] wl[72] vdd gnd cell_6t
Xbit_r73_c0 bl[0] br[0] wl[73] vdd gnd cell_6t
Xbit_r74_c0 bl[0] br[0] wl[74] vdd gnd cell_6t
Xbit_r75_c0 bl[0] br[0] wl[75] vdd gnd cell_6t
Xbit_r76_c0 bl[0] br[0] wl[76] vdd gnd cell_6t
Xbit_r77_c0 bl[0] br[0] wl[77] vdd gnd cell_6t
Xbit_r78_c0 bl[0] br[0] wl[78] vdd gnd cell_6t
Xbit_r79_c0 bl[0] br[0] wl[79] vdd gnd cell_6t
Xbit_r80_c0 bl[0] br[0] wl[80] vdd gnd cell_6t
Xbit_r81_c0 bl[0] br[0] wl[81] vdd gnd cell_6t
Xbit_r82_c0 bl[0] br[0] wl[82] vdd gnd cell_6t
Xbit_r83_c0 bl[0] br[0] wl[83] vdd gnd cell_6t
Xbit_r84_c0 bl[0] br[0] wl[84] vdd gnd cell_6t
Xbit_r85_c0 bl[0] br[0] wl[85] vdd gnd cell_6t
Xbit_r86_c0 bl[0] br[0] wl[86] vdd gnd cell_6t
Xbit_r87_c0 bl[0] br[0] wl[87] vdd gnd cell_6t
Xbit_r88_c0 bl[0] br[0] wl[88] vdd gnd cell_6t
Xbit_r89_c0 bl[0] br[0] wl[89] vdd gnd cell_6t
Xbit_r90_c0 bl[0] br[0] wl[90] vdd gnd cell_6t
Xbit_r91_c0 bl[0] br[0] wl[91] vdd gnd cell_6t
Xbit_r92_c0 bl[0] br[0] wl[92] vdd gnd cell_6t
Xbit_r93_c0 bl[0] br[0] wl[93] vdd gnd cell_6t
Xbit_r94_c0 bl[0] br[0] wl[94] vdd gnd cell_6t
Xbit_r95_c0 bl[0] br[0] wl[95] vdd gnd cell_6t
Xbit_r96_c0 bl[0] br[0] wl[96] vdd gnd cell_6t
Xbit_r97_c0 bl[0] br[0] wl[97] vdd gnd cell_6t
Xbit_r98_c0 bl[0] br[0] wl[98] vdd gnd cell_6t
Xbit_r99_c0 bl[0] br[0] wl[99] vdd gnd cell_6t
Xbit_r100_c0 bl[0] br[0] wl[100] vdd gnd cell_6t
Xbit_r101_c0 bl[0] br[0] wl[101] vdd gnd cell_6t
Xbit_r102_c0 bl[0] br[0] wl[102] vdd gnd cell_6t
Xbit_r103_c0 bl[0] br[0] wl[103] vdd gnd cell_6t
Xbit_r104_c0 bl[0] br[0] wl[104] vdd gnd cell_6t
Xbit_r105_c0 bl[0] br[0] wl[105] vdd gnd cell_6t
Xbit_r106_c0 bl[0] br[0] wl[106] vdd gnd cell_6t
Xbit_r107_c0 bl[0] br[0] wl[107] vdd gnd cell_6t
Xbit_r108_c0 bl[0] br[0] wl[108] vdd gnd cell_6t
Xbit_r109_c0 bl[0] br[0] wl[109] vdd gnd cell_6t
Xbit_r110_c0 bl[0] br[0] wl[110] vdd gnd cell_6t
Xbit_r111_c0 bl[0] br[0] wl[111] vdd gnd cell_6t
Xbit_r112_c0 bl[0] br[0] wl[112] vdd gnd cell_6t
Xbit_r113_c0 bl[0] br[0] wl[113] vdd gnd cell_6t
Xbit_r114_c0 bl[0] br[0] wl[114] vdd gnd cell_6t
Xbit_r115_c0 bl[0] br[0] wl[115] vdd gnd cell_6t
Xbit_r116_c0 bl[0] br[0] wl[116] vdd gnd cell_6t
Xbit_r117_c0 bl[0] br[0] wl[117] vdd gnd cell_6t
Xbit_r118_c0 bl[0] br[0] wl[118] vdd gnd cell_6t
Xbit_r119_c0 bl[0] br[0] wl[119] vdd gnd cell_6t
Xbit_r120_c0 bl[0] br[0] wl[120] vdd gnd cell_6t
Xbit_r121_c0 bl[0] br[0] wl[121] vdd gnd cell_6t
Xbit_r122_c0 bl[0] br[0] wl[122] vdd gnd cell_6t
Xbit_r123_c0 bl[0] br[0] wl[123] vdd gnd cell_6t
Xbit_r124_c0 bl[0] br[0] wl[124] vdd gnd cell_6t
Xbit_r125_c0 bl[0] br[0] wl[125] vdd gnd cell_6t
Xbit_r126_c0 bl[0] br[0] wl[126] vdd gnd cell_6t
Xbit_r127_c0 bl[0] br[0] wl[127] vdd gnd cell_6t
Xbit_r128_c0 bl[0] br[0] wl[128] vdd gnd cell_6t
Xbit_r129_c0 bl[0] br[0] wl[129] vdd gnd cell_6t
Xbit_r130_c0 bl[0] br[0] wl[130] vdd gnd cell_6t
Xbit_r131_c0 bl[0] br[0] wl[131] vdd gnd cell_6t
Xbit_r132_c0 bl[0] br[0] wl[132] vdd gnd cell_6t
Xbit_r133_c0 bl[0] br[0] wl[133] vdd gnd cell_6t
Xbit_r134_c0 bl[0] br[0] wl[134] vdd gnd cell_6t
Xbit_r135_c0 bl[0] br[0] wl[135] vdd gnd cell_6t
Xbit_r136_c0 bl[0] br[0] wl[136] vdd gnd cell_6t
Xbit_r137_c0 bl[0] br[0] wl[137] vdd gnd cell_6t
Xbit_r138_c0 bl[0] br[0] wl[138] vdd gnd cell_6t
Xbit_r139_c0 bl[0] br[0] wl[139] vdd gnd cell_6t
Xbit_r140_c0 bl[0] br[0] wl[140] vdd gnd cell_6t
Xbit_r141_c0 bl[0] br[0] wl[141] vdd gnd cell_6t
Xbit_r142_c0 bl[0] br[0] wl[142] vdd gnd cell_6t
Xbit_r143_c0 bl[0] br[0] wl[143] vdd gnd cell_6t
Xbit_r144_c0 bl[0] br[0] wl[144] vdd gnd cell_6t
Xbit_r145_c0 bl[0] br[0] wl[145] vdd gnd cell_6t
Xbit_r146_c0 bl[0] br[0] wl[146] vdd gnd cell_6t
Xbit_r147_c0 bl[0] br[0] wl[147] vdd gnd cell_6t
Xbit_r148_c0 bl[0] br[0] wl[148] vdd gnd cell_6t
Xbit_r149_c0 bl[0] br[0] wl[149] vdd gnd cell_6t
Xbit_r150_c0 bl[0] br[0] wl[150] vdd gnd cell_6t
Xbit_r151_c0 bl[0] br[0] wl[151] vdd gnd cell_6t
Xbit_r152_c0 bl[0] br[0] wl[152] vdd gnd cell_6t
Xbit_r153_c0 bl[0] br[0] wl[153] vdd gnd cell_6t
Xbit_r154_c0 bl[0] br[0] wl[154] vdd gnd cell_6t
Xbit_r155_c0 bl[0] br[0] wl[155] vdd gnd cell_6t
Xbit_r156_c0 bl[0] br[0] wl[156] vdd gnd cell_6t
Xbit_r157_c0 bl[0] br[0] wl[157] vdd gnd cell_6t
Xbit_r158_c0 bl[0] br[0] wl[158] vdd gnd cell_6t
Xbit_r159_c0 bl[0] br[0] wl[159] vdd gnd cell_6t
Xbit_r160_c0 bl[0] br[0] wl[160] vdd gnd cell_6t
Xbit_r161_c0 bl[0] br[0] wl[161] vdd gnd cell_6t
Xbit_r162_c0 bl[0] br[0] wl[162] vdd gnd cell_6t
Xbit_r163_c0 bl[0] br[0] wl[163] vdd gnd cell_6t
Xbit_r164_c0 bl[0] br[0] wl[164] vdd gnd cell_6t
Xbit_r165_c0 bl[0] br[0] wl[165] vdd gnd cell_6t
Xbit_r166_c0 bl[0] br[0] wl[166] vdd gnd cell_6t
Xbit_r167_c0 bl[0] br[0] wl[167] vdd gnd cell_6t
Xbit_r168_c0 bl[0] br[0] wl[168] vdd gnd cell_6t
Xbit_r169_c0 bl[0] br[0] wl[169] vdd gnd cell_6t
Xbit_r170_c0 bl[0] br[0] wl[170] vdd gnd cell_6t
Xbit_r171_c0 bl[0] br[0] wl[171] vdd gnd cell_6t
Xbit_r172_c0 bl[0] br[0] wl[172] vdd gnd cell_6t
Xbit_r173_c0 bl[0] br[0] wl[173] vdd gnd cell_6t
Xbit_r174_c0 bl[0] br[0] wl[174] vdd gnd cell_6t
Xbit_r175_c0 bl[0] br[0] wl[175] vdd gnd cell_6t
Xbit_r176_c0 bl[0] br[0] wl[176] vdd gnd cell_6t
Xbit_r177_c0 bl[0] br[0] wl[177] vdd gnd cell_6t
Xbit_r178_c0 bl[0] br[0] wl[178] vdd gnd cell_6t
Xbit_r179_c0 bl[0] br[0] wl[179] vdd gnd cell_6t
Xbit_r180_c0 bl[0] br[0] wl[180] vdd gnd cell_6t
Xbit_r181_c0 bl[0] br[0] wl[181] vdd gnd cell_6t
Xbit_r182_c0 bl[0] br[0] wl[182] vdd gnd cell_6t
Xbit_r183_c0 bl[0] br[0] wl[183] vdd gnd cell_6t
Xbit_r184_c0 bl[0] br[0] wl[184] vdd gnd cell_6t
Xbit_r185_c0 bl[0] br[0] wl[185] vdd gnd cell_6t
Xbit_r186_c0 bl[0] br[0] wl[186] vdd gnd cell_6t
Xbit_r187_c0 bl[0] br[0] wl[187] vdd gnd cell_6t
Xbit_r188_c0 bl[0] br[0] wl[188] vdd gnd cell_6t
Xbit_r189_c0 bl[0] br[0] wl[189] vdd gnd cell_6t
Xbit_r190_c0 bl[0] br[0] wl[190] vdd gnd cell_6t
Xbit_r191_c0 bl[0] br[0] wl[191] vdd gnd cell_6t
Xbit_r192_c0 bl[0] br[0] wl[192] vdd gnd cell_6t
Xbit_r193_c0 bl[0] br[0] wl[193] vdd gnd cell_6t
Xbit_r194_c0 bl[0] br[0] wl[194] vdd gnd cell_6t
Xbit_r195_c0 bl[0] br[0] wl[195] vdd gnd cell_6t
Xbit_r196_c0 bl[0] br[0] wl[196] vdd gnd cell_6t
Xbit_r197_c0 bl[0] br[0] wl[197] vdd gnd cell_6t
Xbit_r198_c0 bl[0] br[0] wl[198] vdd gnd cell_6t
Xbit_r199_c0 bl[0] br[0] wl[199] vdd gnd cell_6t
Xbit_r200_c0 bl[0] br[0] wl[200] vdd gnd cell_6t
Xbit_r201_c0 bl[0] br[0] wl[201] vdd gnd cell_6t
Xbit_r202_c0 bl[0] br[0] wl[202] vdd gnd cell_6t
Xbit_r203_c0 bl[0] br[0] wl[203] vdd gnd cell_6t
Xbit_r204_c0 bl[0] br[0] wl[204] vdd gnd cell_6t
Xbit_r205_c0 bl[0] br[0] wl[205] vdd gnd cell_6t
Xbit_r206_c0 bl[0] br[0] wl[206] vdd gnd cell_6t
Xbit_r207_c0 bl[0] br[0] wl[207] vdd gnd cell_6t
Xbit_r208_c0 bl[0] br[0] wl[208] vdd gnd cell_6t
Xbit_r209_c0 bl[0] br[0] wl[209] vdd gnd cell_6t
Xbit_r210_c0 bl[0] br[0] wl[210] vdd gnd cell_6t
Xbit_r211_c0 bl[0] br[0] wl[211] vdd gnd cell_6t
Xbit_r212_c0 bl[0] br[0] wl[212] vdd gnd cell_6t
Xbit_r213_c0 bl[0] br[0] wl[213] vdd gnd cell_6t
Xbit_r214_c0 bl[0] br[0] wl[214] vdd gnd cell_6t
Xbit_r215_c0 bl[0] br[0] wl[215] vdd gnd cell_6t
Xbit_r216_c0 bl[0] br[0] wl[216] vdd gnd cell_6t
Xbit_r217_c0 bl[0] br[0] wl[217] vdd gnd cell_6t
Xbit_r218_c0 bl[0] br[0] wl[218] vdd gnd cell_6t
Xbit_r219_c0 bl[0] br[0] wl[219] vdd gnd cell_6t
Xbit_r220_c0 bl[0] br[0] wl[220] vdd gnd cell_6t
Xbit_r221_c0 bl[0] br[0] wl[221] vdd gnd cell_6t
Xbit_r222_c0 bl[0] br[0] wl[222] vdd gnd cell_6t
Xbit_r223_c0 bl[0] br[0] wl[223] vdd gnd cell_6t
Xbit_r224_c0 bl[0] br[0] wl[224] vdd gnd cell_6t
Xbit_r225_c0 bl[0] br[0] wl[225] vdd gnd cell_6t
Xbit_r226_c0 bl[0] br[0] wl[226] vdd gnd cell_6t
Xbit_r227_c0 bl[0] br[0] wl[227] vdd gnd cell_6t
Xbit_r228_c0 bl[0] br[0] wl[228] vdd gnd cell_6t
Xbit_r229_c0 bl[0] br[0] wl[229] vdd gnd cell_6t
Xbit_r230_c0 bl[0] br[0] wl[230] vdd gnd cell_6t
Xbit_r231_c0 bl[0] br[0] wl[231] vdd gnd cell_6t
Xbit_r232_c0 bl[0] br[0] wl[232] vdd gnd cell_6t
Xbit_r233_c0 bl[0] br[0] wl[233] vdd gnd cell_6t
Xbit_r234_c0 bl[0] br[0] wl[234] vdd gnd cell_6t
Xbit_r235_c0 bl[0] br[0] wl[235] vdd gnd cell_6t
Xbit_r236_c0 bl[0] br[0] wl[236] vdd gnd cell_6t
Xbit_r237_c0 bl[0] br[0] wl[237] vdd gnd cell_6t
Xbit_r238_c0 bl[0] br[0] wl[238] vdd gnd cell_6t
Xbit_r239_c0 bl[0] br[0] wl[239] vdd gnd cell_6t
Xbit_r240_c0 bl[0] br[0] wl[240] vdd gnd cell_6t
Xbit_r241_c0 bl[0] br[0] wl[241] vdd gnd cell_6t
Xbit_r242_c0 bl[0] br[0] wl[242] vdd gnd cell_6t
Xbit_r243_c0 bl[0] br[0] wl[243] vdd gnd cell_6t
Xbit_r244_c0 bl[0] br[0] wl[244] vdd gnd cell_6t
Xbit_r245_c0 bl[0] br[0] wl[245] vdd gnd cell_6t
Xbit_r246_c0 bl[0] br[0] wl[246] vdd gnd cell_6t
Xbit_r247_c0 bl[0] br[0] wl[247] vdd gnd cell_6t
Xbit_r248_c0 bl[0] br[0] wl[248] vdd gnd cell_6t
Xbit_r249_c0 bl[0] br[0] wl[249] vdd gnd cell_6t
Xbit_r250_c0 bl[0] br[0] wl[250] vdd gnd cell_6t
Xbit_r251_c0 bl[0] br[0] wl[251] vdd gnd cell_6t
Xbit_r252_c0 bl[0] br[0] wl[252] vdd gnd cell_6t
Xbit_r253_c0 bl[0] br[0] wl[253] vdd gnd cell_6t
Xbit_r254_c0 bl[0] br[0] wl[254] vdd gnd cell_6t
Xbit_r255_c0 bl[0] br[0] wl[255] vdd gnd cell_6t
Xbit_r0_c1 bl[1] br[1] wl[0] vdd gnd cell_6t
Xbit_r1_c1 bl[1] br[1] wl[1] vdd gnd cell_6t
Xbit_r2_c1 bl[1] br[1] wl[2] vdd gnd cell_6t
Xbit_r3_c1 bl[1] br[1] wl[3] vdd gnd cell_6t
Xbit_r4_c1 bl[1] br[1] wl[4] vdd gnd cell_6t
Xbit_r5_c1 bl[1] br[1] wl[5] vdd gnd cell_6t
Xbit_r6_c1 bl[1] br[1] wl[6] vdd gnd cell_6t
Xbit_r7_c1 bl[1] br[1] wl[7] vdd gnd cell_6t
Xbit_r8_c1 bl[1] br[1] wl[8] vdd gnd cell_6t
Xbit_r9_c1 bl[1] br[1] wl[9] vdd gnd cell_6t
Xbit_r10_c1 bl[1] br[1] wl[10] vdd gnd cell_6t
Xbit_r11_c1 bl[1] br[1] wl[11] vdd gnd cell_6t
Xbit_r12_c1 bl[1] br[1] wl[12] vdd gnd cell_6t
Xbit_r13_c1 bl[1] br[1] wl[13] vdd gnd cell_6t
Xbit_r14_c1 bl[1] br[1] wl[14] vdd gnd cell_6t
Xbit_r15_c1 bl[1] br[1] wl[15] vdd gnd cell_6t
Xbit_r16_c1 bl[1] br[1] wl[16] vdd gnd cell_6t
Xbit_r17_c1 bl[1] br[1] wl[17] vdd gnd cell_6t
Xbit_r18_c1 bl[1] br[1] wl[18] vdd gnd cell_6t
Xbit_r19_c1 bl[1] br[1] wl[19] vdd gnd cell_6t
Xbit_r20_c1 bl[1] br[1] wl[20] vdd gnd cell_6t
Xbit_r21_c1 bl[1] br[1] wl[21] vdd gnd cell_6t
Xbit_r22_c1 bl[1] br[1] wl[22] vdd gnd cell_6t
Xbit_r23_c1 bl[1] br[1] wl[23] vdd gnd cell_6t
Xbit_r24_c1 bl[1] br[1] wl[24] vdd gnd cell_6t
Xbit_r25_c1 bl[1] br[1] wl[25] vdd gnd cell_6t
Xbit_r26_c1 bl[1] br[1] wl[26] vdd gnd cell_6t
Xbit_r27_c1 bl[1] br[1] wl[27] vdd gnd cell_6t
Xbit_r28_c1 bl[1] br[1] wl[28] vdd gnd cell_6t
Xbit_r29_c1 bl[1] br[1] wl[29] vdd gnd cell_6t
Xbit_r30_c1 bl[1] br[1] wl[30] vdd gnd cell_6t
Xbit_r31_c1 bl[1] br[1] wl[31] vdd gnd cell_6t
Xbit_r32_c1 bl[1] br[1] wl[32] vdd gnd cell_6t
Xbit_r33_c1 bl[1] br[1] wl[33] vdd gnd cell_6t
Xbit_r34_c1 bl[1] br[1] wl[34] vdd gnd cell_6t
Xbit_r35_c1 bl[1] br[1] wl[35] vdd gnd cell_6t
Xbit_r36_c1 bl[1] br[1] wl[36] vdd gnd cell_6t
Xbit_r37_c1 bl[1] br[1] wl[37] vdd gnd cell_6t
Xbit_r38_c1 bl[1] br[1] wl[38] vdd gnd cell_6t
Xbit_r39_c1 bl[1] br[1] wl[39] vdd gnd cell_6t
Xbit_r40_c1 bl[1] br[1] wl[40] vdd gnd cell_6t
Xbit_r41_c1 bl[1] br[1] wl[41] vdd gnd cell_6t
Xbit_r42_c1 bl[1] br[1] wl[42] vdd gnd cell_6t
Xbit_r43_c1 bl[1] br[1] wl[43] vdd gnd cell_6t
Xbit_r44_c1 bl[1] br[1] wl[44] vdd gnd cell_6t
Xbit_r45_c1 bl[1] br[1] wl[45] vdd gnd cell_6t
Xbit_r46_c1 bl[1] br[1] wl[46] vdd gnd cell_6t
Xbit_r47_c1 bl[1] br[1] wl[47] vdd gnd cell_6t
Xbit_r48_c1 bl[1] br[1] wl[48] vdd gnd cell_6t
Xbit_r49_c1 bl[1] br[1] wl[49] vdd gnd cell_6t
Xbit_r50_c1 bl[1] br[1] wl[50] vdd gnd cell_6t
Xbit_r51_c1 bl[1] br[1] wl[51] vdd gnd cell_6t
Xbit_r52_c1 bl[1] br[1] wl[52] vdd gnd cell_6t
Xbit_r53_c1 bl[1] br[1] wl[53] vdd gnd cell_6t
Xbit_r54_c1 bl[1] br[1] wl[54] vdd gnd cell_6t
Xbit_r55_c1 bl[1] br[1] wl[55] vdd gnd cell_6t
Xbit_r56_c1 bl[1] br[1] wl[56] vdd gnd cell_6t
Xbit_r57_c1 bl[1] br[1] wl[57] vdd gnd cell_6t
Xbit_r58_c1 bl[1] br[1] wl[58] vdd gnd cell_6t
Xbit_r59_c1 bl[1] br[1] wl[59] vdd gnd cell_6t
Xbit_r60_c1 bl[1] br[1] wl[60] vdd gnd cell_6t
Xbit_r61_c1 bl[1] br[1] wl[61] vdd gnd cell_6t
Xbit_r62_c1 bl[1] br[1] wl[62] vdd gnd cell_6t
Xbit_r63_c1 bl[1] br[1] wl[63] vdd gnd cell_6t
Xbit_r64_c1 bl[1] br[1] wl[64] vdd gnd cell_6t
Xbit_r65_c1 bl[1] br[1] wl[65] vdd gnd cell_6t
Xbit_r66_c1 bl[1] br[1] wl[66] vdd gnd cell_6t
Xbit_r67_c1 bl[1] br[1] wl[67] vdd gnd cell_6t
Xbit_r68_c1 bl[1] br[1] wl[68] vdd gnd cell_6t
Xbit_r69_c1 bl[1] br[1] wl[69] vdd gnd cell_6t
Xbit_r70_c1 bl[1] br[1] wl[70] vdd gnd cell_6t
Xbit_r71_c1 bl[1] br[1] wl[71] vdd gnd cell_6t
Xbit_r72_c1 bl[1] br[1] wl[72] vdd gnd cell_6t
Xbit_r73_c1 bl[1] br[1] wl[73] vdd gnd cell_6t
Xbit_r74_c1 bl[1] br[1] wl[74] vdd gnd cell_6t
Xbit_r75_c1 bl[1] br[1] wl[75] vdd gnd cell_6t
Xbit_r76_c1 bl[1] br[1] wl[76] vdd gnd cell_6t
Xbit_r77_c1 bl[1] br[1] wl[77] vdd gnd cell_6t
Xbit_r78_c1 bl[1] br[1] wl[78] vdd gnd cell_6t
Xbit_r79_c1 bl[1] br[1] wl[79] vdd gnd cell_6t
Xbit_r80_c1 bl[1] br[1] wl[80] vdd gnd cell_6t
Xbit_r81_c1 bl[1] br[1] wl[81] vdd gnd cell_6t
Xbit_r82_c1 bl[1] br[1] wl[82] vdd gnd cell_6t
Xbit_r83_c1 bl[1] br[1] wl[83] vdd gnd cell_6t
Xbit_r84_c1 bl[1] br[1] wl[84] vdd gnd cell_6t
Xbit_r85_c1 bl[1] br[1] wl[85] vdd gnd cell_6t
Xbit_r86_c1 bl[1] br[1] wl[86] vdd gnd cell_6t
Xbit_r87_c1 bl[1] br[1] wl[87] vdd gnd cell_6t
Xbit_r88_c1 bl[1] br[1] wl[88] vdd gnd cell_6t
Xbit_r89_c1 bl[1] br[1] wl[89] vdd gnd cell_6t
Xbit_r90_c1 bl[1] br[1] wl[90] vdd gnd cell_6t
Xbit_r91_c1 bl[1] br[1] wl[91] vdd gnd cell_6t
Xbit_r92_c1 bl[1] br[1] wl[92] vdd gnd cell_6t
Xbit_r93_c1 bl[1] br[1] wl[93] vdd gnd cell_6t
Xbit_r94_c1 bl[1] br[1] wl[94] vdd gnd cell_6t
Xbit_r95_c1 bl[1] br[1] wl[95] vdd gnd cell_6t
Xbit_r96_c1 bl[1] br[1] wl[96] vdd gnd cell_6t
Xbit_r97_c1 bl[1] br[1] wl[97] vdd gnd cell_6t
Xbit_r98_c1 bl[1] br[1] wl[98] vdd gnd cell_6t
Xbit_r99_c1 bl[1] br[1] wl[99] vdd gnd cell_6t
Xbit_r100_c1 bl[1] br[1] wl[100] vdd gnd cell_6t
Xbit_r101_c1 bl[1] br[1] wl[101] vdd gnd cell_6t
Xbit_r102_c1 bl[1] br[1] wl[102] vdd gnd cell_6t
Xbit_r103_c1 bl[1] br[1] wl[103] vdd gnd cell_6t
Xbit_r104_c1 bl[1] br[1] wl[104] vdd gnd cell_6t
Xbit_r105_c1 bl[1] br[1] wl[105] vdd gnd cell_6t
Xbit_r106_c1 bl[1] br[1] wl[106] vdd gnd cell_6t
Xbit_r107_c1 bl[1] br[1] wl[107] vdd gnd cell_6t
Xbit_r108_c1 bl[1] br[1] wl[108] vdd gnd cell_6t
Xbit_r109_c1 bl[1] br[1] wl[109] vdd gnd cell_6t
Xbit_r110_c1 bl[1] br[1] wl[110] vdd gnd cell_6t
Xbit_r111_c1 bl[1] br[1] wl[111] vdd gnd cell_6t
Xbit_r112_c1 bl[1] br[1] wl[112] vdd gnd cell_6t
Xbit_r113_c1 bl[1] br[1] wl[113] vdd gnd cell_6t
Xbit_r114_c1 bl[1] br[1] wl[114] vdd gnd cell_6t
Xbit_r115_c1 bl[1] br[1] wl[115] vdd gnd cell_6t
Xbit_r116_c1 bl[1] br[1] wl[116] vdd gnd cell_6t
Xbit_r117_c1 bl[1] br[1] wl[117] vdd gnd cell_6t
Xbit_r118_c1 bl[1] br[1] wl[118] vdd gnd cell_6t
Xbit_r119_c1 bl[1] br[1] wl[119] vdd gnd cell_6t
Xbit_r120_c1 bl[1] br[1] wl[120] vdd gnd cell_6t
Xbit_r121_c1 bl[1] br[1] wl[121] vdd gnd cell_6t
Xbit_r122_c1 bl[1] br[1] wl[122] vdd gnd cell_6t
Xbit_r123_c1 bl[1] br[1] wl[123] vdd gnd cell_6t
Xbit_r124_c1 bl[1] br[1] wl[124] vdd gnd cell_6t
Xbit_r125_c1 bl[1] br[1] wl[125] vdd gnd cell_6t
Xbit_r126_c1 bl[1] br[1] wl[126] vdd gnd cell_6t
Xbit_r127_c1 bl[1] br[1] wl[127] vdd gnd cell_6t
Xbit_r128_c1 bl[1] br[1] wl[128] vdd gnd cell_6t
Xbit_r129_c1 bl[1] br[1] wl[129] vdd gnd cell_6t
Xbit_r130_c1 bl[1] br[1] wl[130] vdd gnd cell_6t
Xbit_r131_c1 bl[1] br[1] wl[131] vdd gnd cell_6t
Xbit_r132_c1 bl[1] br[1] wl[132] vdd gnd cell_6t
Xbit_r133_c1 bl[1] br[1] wl[133] vdd gnd cell_6t
Xbit_r134_c1 bl[1] br[1] wl[134] vdd gnd cell_6t
Xbit_r135_c1 bl[1] br[1] wl[135] vdd gnd cell_6t
Xbit_r136_c1 bl[1] br[1] wl[136] vdd gnd cell_6t
Xbit_r137_c1 bl[1] br[1] wl[137] vdd gnd cell_6t
Xbit_r138_c1 bl[1] br[1] wl[138] vdd gnd cell_6t
Xbit_r139_c1 bl[1] br[1] wl[139] vdd gnd cell_6t
Xbit_r140_c1 bl[1] br[1] wl[140] vdd gnd cell_6t
Xbit_r141_c1 bl[1] br[1] wl[141] vdd gnd cell_6t
Xbit_r142_c1 bl[1] br[1] wl[142] vdd gnd cell_6t
Xbit_r143_c1 bl[1] br[1] wl[143] vdd gnd cell_6t
Xbit_r144_c1 bl[1] br[1] wl[144] vdd gnd cell_6t
Xbit_r145_c1 bl[1] br[1] wl[145] vdd gnd cell_6t
Xbit_r146_c1 bl[1] br[1] wl[146] vdd gnd cell_6t
Xbit_r147_c1 bl[1] br[1] wl[147] vdd gnd cell_6t
Xbit_r148_c1 bl[1] br[1] wl[148] vdd gnd cell_6t
Xbit_r149_c1 bl[1] br[1] wl[149] vdd gnd cell_6t
Xbit_r150_c1 bl[1] br[1] wl[150] vdd gnd cell_6t
Xbit_r151_c1 bl[1] br[1] wl[151] vdd gnd cell_6t
Xbit_r152_c1 bl[1] br[1] wl[152] vdd gnd cell_6t
Xbit_r153_c1 bl[1] br[1] wl[153] vdd gnd cell_6t
Xbit_r154_c1 bl[1] br[1] wl[154] vdd gnd cell_6t
Xbit_r155_c1 bl[1] br[1] wl[155] vdd gnd cell_6t
Xbit_r156_c1 bl[1] br[1] wl[156] vdd gnd cell_6t
Xbit_r157_c1 bl[1] br[1] wl[157] vdd gnd cell_6t
Xbit_r158_c1 bl[1] br[1] wl[158] vdd gnd cell_6t
Xbit_r159_c1 bl[1] br[1] wl[159] vdd gnd cell_6t
Xbit_r160_c1 bl[1] br[1] wl[160] vdd gnd cell_6t
Xbit_r161_c1 bl[1] br[1] wl[161] vdd gnd cell_6t
Xbit_r162_c1 bl[1] br[1] wl[162] vdd gnd cell_6t
Xbit_r163_c1 bl[1] br[1] wl[163] vdd gnd cell_6t
Xbit_r164_c1 bl[1] br[1] wl[164] vdd gnd cell_6t
Xbit_r165_c1 bl[1] br[1] wl[165] vdd gnd cell_6t
Xbit_r166_c1 bl[1] br[1] wl[166] vdd gnd cell_6t
Xbit_r167_c1 bl[1] br[1] wl[167] vdd gnd cell_6t
Xbit_r168_c1 bl[1] br[1] wl[168] vdd gnd cell_6t
Xbit_r169_c1 bl[1] br[1] wl[169] vdd gnd cell_6t
Xbit_r170_c1 bl[1] br[1] wl[170] vdd gnd cell_6t
Xbit_r171_c1 bl[1] br[1] wl[171] vdd gnd cell_6t
Xbit_r172_c1 bl[1] br[1] wl[172] vdd gnd cell_6t
Xbit_r173_c1 bl[1] br[1] wl[173] vdd gnd cell_6t
Xbit_r174_c1 bl[1] br[1] wl[174] vdd gnd cell_6t
Xbit_r175_c1 bl[1] br[1] wl[175] vdd gnd cell_6t
Xbit_r176_c1 bl[1] br[1] wl[176] vdd gnd cell_6t
Xbit_r177_c1 bl[1] br[1] wl[177] vdd gnd cell_6t
Xbit_r178_c1 bl[1] br[1] wl[178] vdd gnd cell_6t
Xbit_r179_c1 bl[1] br[1] wl[179] vdd gnd cell_6t
Xbit_r180_c1 bl[1] br[1] wl[180] vdd gnd cell_6t
Xbit_r181_c1 bl[1] br[1] wl[181] vdd gnd cell_6t
Xbit_r182_c1 bl[1] br[1] wl[182] vdd gnd cell_6t
Xbit_r183_c1 bl[1] br[1] wl[183] vdd gnd cell_6t
Xbit_r184_c1 bl[1] br[1] wl[184] vdd gnd cell_6t
Xbit_r185_c1 bl[1] br[1] wl[185] vdd gnd cell_6t
Xbit_r186_c1 bl[1] br[1] wl[186] vdd gnd cell_6t
Xbit_r187_c1 bl[1] br[1] wl[187] vdd gnd cell_6t
Xbit_r188_c1 bl[1] br[1] wl[188] vdd gnd cell_6t
Xbit_r189_c1 bl[1] br[1] wl[189] vdd gnd cell_6t
Xbit_r190_c1 bl[1] br[1] wl[190] vdd gnd cell_6t
Xbit_r191_c1 bl[1] br[1] wl[191] vdd gnd cell_6t
Xbit_r192_c1 bl[1] br[1] wl[192] vdd gnd cell_6t
Xbit_r193_c1 bl[1] br[1] wl[193] vdd gnd cell_6t
Xbit_r194_c1 bl[1] br[1] wl[194] vdd gnd cell_6t
Xbit_r195_c1 bl[1] br[1] wl[195] vdd gnd cell_6t
Xbit_r196_c1 bl[1] br[1] wl[196] vdd gnd cell_6t
Xbit_r197_c1 bl[1] br[1] wl[197] vdd gnd cell_6t
Xbit_r198_c1 bl[1] br[1] wl[198] vdd gnd cell_6t
Xbit_r199_c1 bl[1] br[1] wl[199] vdd gnd cell_6t
Xbit_r200_c1 bl[1] br[1] wl[200] vdd gnd cell_6t
Xbit_r201_c1 bl[1] br[1] wl[201] vdd gnd cell_6t
Xbit_r202_c1 bl[1] br[1] wl[202] vdd gnd cell_6t
Xbit_r203_c1 bl[1] br[1] wl[203] vdd gnd cell_6t
Xbit_r204_c1 bl[1] br[1] wl[204] vdd gnd cell_6t
Xbit_r205_c1 bl[1] br[1] wl[205] vdd gnd cell_6t
Xbit_r206_c1 bl[1] br[1] wl[206] vdd gnd cell_6t
Xbit_r207_c1 bl[1] br[1] wl[207] vdd gnd cell_6t
Xbit_r208_c1 bl[1] br[1] wl[208] vdd gnd cell_6t
Xbit_r209_c1 bl[1] br[1] wl[209] vdd gnd cell_6t
Xbit_r210_c1 bl[1] br[1] wl[210] vdd gnd cell_6t
Xbit_r211_c1 bl[1] br[1] wl[211] vdd gnd cell_6t
Xbit_r212_c1 bl[1] br[1] wl[212] vdd gnd cell_6t
Xbit_r213_c1 bl[1] br[1] wl[213] vdd gnd cell_6t
Xbit_r214_c1 bl[1] br[1] wl[214] vdd gnd cell_6t
Xbit_r215_c1 bl[1] br[1] wl[215] vdd gnd cell_6t
Xbit_r216_c1 bl[1] br[1] wl[216] vdd gnd cell_6t
Xbit_r217_c1 bl[1] br[1] wl[217] vdd gnd cell_6t
Xbit_r218_c1 bl[1] br[1] wl[218] vdd gnd cell_6t
Xbit_r219_c1 bl[1] br[1] wl[219] vdd gnd cell_6t
Xbit_r220_c1 bl[1] br[1] wl[220] vdd gnd cell_6t
Xbit_r221_c1 bl[1] br[1] wl[221] vdd gnd cell_6t
Xbit_r222_c1 bl[1] br[1] wl[222] vdd gnd cell_6t
Xbit_r223_c1 bl[1] br[1] wl[223] vdd gnd cell_6t
Xbit_r224_c1 bl[1] br[1] wl[224] vdd gnd cell_6t
Xbit_r225_c1 bl[1] br[1] wl[225] vdd gnd cell_6t
Xbit_r226_c1 bl[1] br[1] wl[226] vdd gnd cell_6t
Xbit_r227_c1 bl[1] br[1] wl[227] vdd gnd cell_6t
Xbit_r228_c1 bl[1] br[1] wl[228] vdd gnd cell_6t
Xbit_r229_c1 bl[1] br[1] wl[229] vdd gnd cell_6t
Xbit_r230_c1 bl[1] br[1] wl[230] vdd gnd cell_6t
Xbit_r231_c1 bl[1] br[1] wl[231] vdd gnd cell_6t
Xbit_r232_c1 bl[1] br[1] wl[232] vdd gnd cell_6t
Xbit_r233_c1 bl[1] br[1] wl[233] vdd gnd cell_6t
Xbit_r234_c1 bl[1] br[1] wl[234] vdd gnd cell_6t
Xbit_r235_c1 bl[1] br[1] wl[235] vdd gnd cell_6t
Xbit_r236_c1 bl[1] br[1] wl[236] vdd gnd cell_6t
Xbit_r237_c1 bl[1] br[1] wl[237] vdd gnd cell_6t
Xbit_r238_c1 bl[1] br[1] wl[238] vdd gnd cell_6t
Xbit_r239_c1 bl[1] br[1] wl[239] vdd gnd cell_6t
Xbit_r240_c1 bl[1] br[1] wl[240] vdd gnd cell_6t
Xbit_r241_c1 bl[1] br[1] wl[241] vdd gnd cell_6t
Xbit_r242_c1 bl[1] br[1] wl[242] vdd gnd cell_6t
Xbit_r243_c1 bl[1] br[1] wl[243] vdd gnd cell_6t
Xbit_r244_c1 bl[1] br[1] wl[244] vdd gnd cell_6t
Xbit_r245_c1 bl[1] br[1] wl[245] vdd gnd cell_6t
Xbit_r246_c1 bl[1] br[1] wl[246] vdd gnd cell_6t
Xbit_r247_c1 bl[1] br[1] wl[247] vdd gnd cell_6t
Xbit_r248_c1 bl[1] br[1] wl[248] vdd gnd cell_6t
Xbit_r249_c1 bl[1] br[1] wl[249] vdd gnd cell_6t
Xbit_r250_c1 bl[1] br[1] wl[250] vdd gnd cell_6t
Xbit_r251_c1 bl[1] br[1] wl[251] vdd gnd cell_6t
Xbit_r252_c1 bl[1] br[1] wl[252] vdd gnd cell_6t
Xbit_r253_c1 bl[1] br[1] wl[253] vdd gnd cell_6t
Xbit_r254_c1 bl[1] br[1] wl[254] vdd gnd cell_6t
Xbit_r255_c1 bl[1] br[1] wl[255] vdd gnd cell_6t
Xbit_r0_c2 bl[2] br[2] wl[0] vdd gnd cell_6t
Xbit_r1_c2 bl[2] br[2] wl[1] vdd gnd cell_6t
Xbit_r2_c2 bl[2] br[2] wl[2] vdd gnd cell_6t
Xbit_r3_c2 bl[2] br[2] wl[3] vdd gnd cell_6t
Xbit_r4_c2 bl[2] br[2] wl[4] vdd gnd cell_6t
Xbit_r5_c2 bl[2] br[2] wl[5] vdd gnd cell_6t
Xbit_r6_c2 bl[2] br[2] wl[6] vdd gnd cell_6t
Xbit_r7_c2 bl[2] br[2] wl[7] vdd gnd cell_6t
Xbit_r8_c2 bl[2] br[2] wl[8] vdd gnd cell_6t
Xbit_r9_c2 bl[2] br[2] wl[9] vdd gnd cell_6t
Xbit_r10_c2 bl[2] br[2] wl[10] vdd gnd cell_6t
Xbit_r11_c2 bl[2] br[2] wl[11] vdd gnd cell_6t
Xbit_r12_c2 bl[2] br[2] wl[12] vdd gnd cell_6t
Xbit_r13_c2 bl[2] br[2] wl[13] vdd gnd cell_6t
Xbit_r14_c2 bl[2] br[2] wl[14] vdd gnd cell_6t
Xbit_r15_c2 bl[2] br[2] wl[15] vdd gnd cell_6t
Xbit_r16_c2 bl[2] br[2] wl[16] vdd gnd cell_6t
Xbit_r17_c2 bl[2] br[2] wl[17] vdd gnd cell_6t
Xbit_r18_c2 bl[2] br[2] wl[18] vdd gnd cell_6t
Xbit_r19_c2 bl[2] br[2] wl[19] vdd gnd cell_6t
Xbit_r20_c2 bl[2] br[2] wl[20] vdd gnd cell_6t
Xbit_r21_c2 bl[2] br[2] wl[21] vdd gnd cell_6t
Xbit_r22_c2 bl[2] br[2] wl[22] vdd gnd cell_6t
Xbit_r23_c2 bl[2] br[2] wl[23] vdd gnd cell_6t
Xbit_r24_c2 bl[2] br[2] wl[24] vdd gnd cell_6t
Xbit_r25_c2 bl[2] br[2] wl[25] vdd gnd cell_6t
Xbit_r26_c2 bl[2] br[2] wl[26] vdd gnd cell_6t
Xbit_r27_c2 bl[2] br[2] wl[27] vdd gnd cell_6t
Xbit_r28_c2 bl[2] br[2] wl[28] vdd gnd cell_6t
Xbit_r29_c2 bl[2] br[2] wl[29] vdd gnd cell_6t
Xbit_r30_c2 bl[2] br[2] wl[30] vdd gnd cell_6t
Xbit_r31_c2 bl[2] br[2] wl[31] vdd gnd cell_6t
Xbit_r32_c2 bl[2] br[2] wl[32] vdd gnd cell_6t
Xbit_r33_c2 bl[2] br[2] wl[33] vdd gnd cell_6t
Xbit_r34_c2 bl[2] br[2] wl[34] vdd gnd cell_6t
Xbit_r35_c2 bl[2] br[2] wl[35] vdd gnd cell_6t
Xbit_r36_c2 bl[2] br[2] wl[36] vdd gnd cell_6t
Xbit_r37_c2 bl[2] br[2] wl[37] vdd gnd cell_6t
Xbit_r38_c2 bl[2] br[2] wl[38] vdd gnd cell_6t
Xbit_r39_c2 bl[2] br[2] wl[39] vdd gnd cell_6t
Xbit_r40_c2 bl[2] br[2] wl[40] vdd gnd cell_6t
Xbit_r41_c2 bl[2] br[2] wl[41] vdd gnd cell_6t
Xbit_r42_c2 bl[2] br[2] wl[42] vdd gnd cell_6t
Xbit_r43_c2 bl[2] br[2] wl[43] vdd gnd cell_6t
Xbit_r44_c2 bl[2] br[2] wl[44] vdd gnd cell_6t
Xbit_r45_c2 bl[2] br[2] wl[45] vdd gnd cell_6t
Xbit_r46_c2 bl[2] br[2] wl[46] vdd gnd cell_6t
Xbit_r47_c2 bl[2] br[2] wl[47] vdd gnd cell_6t
Xbit_r48_c2 bl[2] br[2] wl[48] vdd gnd cell_6t
Xbit_r49_c2 bl[2] br[2] wl[49] vdd gnd cell_6t
Xbit_r50_c2 bl[2] br[2] wl[50] vdd gnd cell_6t
Xbit_r51_c2 bl[2] br[2] wl[51] vdd gnd cell_6t
Xbit_r52_c2 bl[2] br[2] wl[52] vdd gnd cell_6t
Xbit_r53_c2 bl[2] br[2] wl[53] vdd gnd cell_6t
Xbit_r54_c2 bl[2] br[2] wl[54] vdd gnd cell_6t
Xbit_r55_c2 bl[2] br[2] wl[55] vdd gnd cell_6t
Xbit_r56_c2 bl[2] br[2] wl[56] vdd gnd cell_6t
Xbit_r57_c2 bl[2] br[2] wl[57] vdd gnd cell_6t
Xbit_r58_c2 bl[2] br[2] wl[58] vdd gnd cell_6t
Xbit_r59_c2 bl[2] br[2] wl[59] vdd gnd cell_6t
Xbit_r60_c2 bl[2] br[2] wl[60] vdd gnd cell_6t
Xbit_r61_c2 bl[2] br[2] wl[61] vdd gnd cell_6t
Xbit_r62_c2 bl[2] br[2] wl[62] vdd gnd cell_6t
Xbit_r63_c2 bl[2] br[2] wl[63] vdd gnd cell_6t
Xbit_r64_c2 bl[2] br[2] wl[64] vdd gnd cell_6t
Xbit_r65_c2 bl[2] br[2] wl[65] vdd gnd cell_6t
Xbit_r66_c2 bl[2] br[2] wl[66] vdd gnd cell_6t
Xbit_r67_c2 bl[2] br[2] wl[67] vdd gnd cell_6t
Xbit_r68_c2 bl[2] br[2] wl[68] vdd gnd cell_6t
Xbit_r69_c2 bl[2] br[2] wl[69] vdd gnd cell_6t
Xbit_r70_c2 bl[2] br[2] wl[70] vdd gnd cell_6t
Xbit_r71_c2 bl[2] br[2] wl[71] vdd gnd cell_6t
Xbit_r72_c2 bl[2] br[2] wl[72] vdd gnd cell_6t
Xbit_r73_c2 bl[2] br[2] wl[73] vdd gnd cell_6t
Xbit_r74_c2 bl[2] br[2] wl[74] vdd gnd cell_6t
Xbit_r75_c2 bl[2] br[2] wl[75] vdd gnd cell_6t
Xbit_r76_c2 bl[2] br[2] wl[76] vdd gnd cell_6t
Xbit_r77_c2 bl[2] br[2] wl[77] vdd gnd cell_6t
Xbit_r78_c2 bl[2] br[2] wl[78] vdd gnd cell_6t
Xbit_r79_c2 bl[2] br[2] wl[79] vdd gnd cell_6t
Xbit_r80_c2 bl[2] br[2] wl[80] vdd gnd cell_6t
Xbit_r81_c2 bl[2] br[2] wl[81] vdd gnd cell_6t
Xbit_r82_c2 bl[2] br[2] wl[82] vdd gnd cell_6t
Xbit_r83_c2 bl[2] br[2] wl[83] vdd gnd cell_6t
Xbit_r84_c2 bl[2] br[2] wl[84] vdd gnd cell_6t
Xbit_r85_c2 bl[2] br[2] wl[85] vdd gnd cell_6t
Xbit_r86_c2 bl[2] br[2] wl[86] vdd gnd cell_6t
Xbit_r87_c2 bl[2] br[2] wl[87] vdd gnd cell_6t
Xbit_r88_c2 bl[2] br[2] wl[88] vdd gnd cell_6t
Xbit_r89_c2 bl[2] br[2] wl[89] vdd gnd cell_6t
Xbit_r90_c2 bl[2] br[2] wl[90] vdd gnd cell_6t
Xbit_r91_c2 bl[2] br[2] wl[91] vdd gnd cell_6t
Xbit_r92_c2 bl[2] br[2] wl[92] vdd gnd cell_6t
Xbit_r93_c2 bl[2] br[2] wl[93] vdd gnd cell_6t
Xbit_r94_c2 bl[2] br[2] wl[94] vdd gnd cell_6t
Xbit_r95_c2 bl[2] br[2] wl[95] vdd gnd cell_6t
Xbit_r96_c2 bl[2] br[2] wl[96] vdd gnd cell_6t
Xbit_r97_c2 bl[2] br[2] wl[97] vdd gnd cell_6t
Xbit_r98_c2 bl[2] br[2] wl[98] vdd gnd cell_6t
Xbit_r99_c2 bl[2] br[2] wl[99] vdd gnd cell_6t
Xbit_r100_c2 bl[2] br[2] wl[100] vdd gnd cell_6t
Xbit_r101_c2 bl[2] br[2] wl[101] vdd gnd cell_6t
Xbit_r102_c2 bl[2] br[2] wl[102] vdd gnd cell_6t
Xbit_r103_c2 bl[2] br[2] wl[103] vdd gnd cell_6t
Xbit_r104_c2 bl[2] br[2] wl[104] vdd gnd cell_6t
Xbit_r105_c2 bl[2] br[2] wl[105] vdd gnd cell_6t
Xbit_r106_c2 bl[2] br[2] wl[106] vdd gnd cell_6t
Xbit_r107_c2 bl[2] br[2] wl[107] vdd gnd cell_6t
Xbit_r108_c2 bl[2] br[2] wl[108] vdd gnd cell_6t
Xbit_r109_c2 bl[2] br[2] wl[109] vdd gnd cell_6t
Xbit_r110_c2 bl[2] br[2] wl[110] vdd gnd cell_6t
Xbit_r111_c2 bl[2] br[2] wl[111] vdd gnd cell_6t
Xbit_r112_c2 bl[2] br[2] wl[112] vdd gnd cell_6t
Xbit_r113_c2 bl[2] br[2] wl[113] vdd gnd cell_6t
Xbit_r114_c2 bl[2] br[2] wl[114] vdd gnd cell_6t
Xbit_r115_c2 bl[2] br[2] wl[115] vdd gnd cell_6t
Xbit_r116_c2 bl[2] br[2] wl[116] vdd gnd cell_6t
Xbit_r117_c2 bl[2] br[2] wl[117] vdd gnd cell_6t
Xbit_r118_c2 bl[2] br[2] wl[118] vdd gnd cell_6t
Xbit_r119_c2 bl[2] br[2] wl[119] vdd gnd cell_6t
Xbit_r120_c2 bl[2] br[2] wl[120] vdd gnd cell_6t
Xbit_r121_c2 bl[2] br[2] wl[121] vdd gnd cell_6t
Xbit_r122_c2 bl[2] br[2] wl[122] vdd gnd cell_6t
Xbit_r123_c2 bl[2] br[2] wl[123] vdd gnd cell_6t
Xbit_r124_c2 bl[2] br[2] wl[124] vdd gnd cell_6t
Xbit_r125_c2 bl[2] br[2] wl[125] vdd gnd cell_6t
Xbit_r126_c2 bl[2] br[2] wl[126] vdd gnd cell_6t
Xbit_r127_c2 bl[2] br[2] wl[127] vdd gnd cell_6t
Xbit_r128_c2 bl[2] br[2] wl[128] vdd gnd cell_6t
Xbit_r129_c2 bl[2] br[2] wl[129] vdd gnd cell_6t
Xbit_r130_c2 bl[2] br[2] wl[130] vdd gnd cell_6t
Xbit_r131_c2 bl[2] br[2] wl[131] vdd gnd cell_6t
Xbit_r132_c2 bl[2] br[2] wl[132] vdd gnd cell_6t
Xbit_r133_c2 bl[2] br[2] wl[133] vdd gnd cell_6t
Xbit_r134_c2 bl[2] br[2] wl[134] vdd gnd cell_6t
Xbit_r135_c2 bl[2] br[2] wl[135] vdd gnd cell_6t
Xbit_r136_c2 bl[2] br[2] wl[136] vdd gnd cell_6t
Xbit_r137_c2 bl[2] br[2] wl[137] vdd gnd cell_6t
Xbit_r138_c2 bl[2] br[2] wl[138] vdd gnd cell_6t
Xbit_r139_c2 bl[2] br[2] wl[139] vdd gnd cell_6t
Xbit_r140_c2 bl[2] br[2] wl[140] vdd gnd cell_6t
Xbit_r141_c2 bl[2] br[2] wl[141] vdd gnd cell_6t
Xbit_r142_c2 bl[2] br[2] wl[142] vdd gnd cell_6t
Xbit_r143_c2 bl[2] br[2] wl[143] vdd gnd cell_6t
Xbit_r144_c2 bl[2] br[2] wl[144] vdd gnd cell_6t
Xbit_r145_c2 bl[2] br[2] wl[145] vdd gnd cell_6t
Xbit_r146_c2 bl[2] br[2] wl[146] vdd gnd cell_6t
Xbit_r147_c2 bl[2] br[2] wl[147] vdd gnd cell_6t
Xbit_r148_c2 bl[2] br[2] wl[148] vdd gnd cell_6t
Xbit_r149_c2 bl[2] br[2] wl[149] vdd gnd cell_6t
Xbit_r150_c2 bl[2] br[2] wl[150] vdd gnd cell_6t
Xbit_r151_c2 bl[2] br[2] wl[151] vdd gnd cell_6t
Xbit_r152_c2 bl[2] br[2] wl[152] vdd gnd cell_6t
Xbit_r153_c2 bl[2] br[2] wl[153] vdd gnd cell_6t
Xbit_r154_c2 bl[2] br[2] wl[154] vdd gnd cell_6t
Xbit_r155_c2 bl[2] br[2] wl[155] vdd gnd cell_6t
Xbit_r156_c2 bl[2] br[2] wl[156] vdd gnd cell_6t
Xbit_r157_c2 bl[2] br[2] wl[157] vdd gnd cell_6t
Xbit_r158_c2 bl[2] br[2] wl[158] vdd gnd cell_6t
Xbit_r159_c2 bl[2] br[2] wl[159] vdd gnd cell_6t
Xbit_r160_c2 bl[2] br[2] wl[160] vdd gnd cell_6t
Xbit_r161_c2 bl[2] br[2] wl[161] vdd gnd cell_6t
Xbit_r162_c2 bl[2] br[2] wl[162] vdd gnd cell_6t
Xbit_r163_c2 bl[2] br[2] wl[163] vdd gnd cell_6t
Xbit_r164_c2 bl[2] br[2] wl[164] vdd gnd cell_6t
Xbit_r165_c2 bl[2] br[2] wl[165] vdd gnd cell_6t
Xbit_r166_c2 bl[2] br[2] wl[166] vdd gnd cell_6t
Xbit_r167_c2 bl[2] br[2] wl[167] vdd gnd cell_6t
Xbit_r168_c2 bl[2] br[2] wl[168] vdd gnd cell_6t
Xbit_r169_c2 bl[2] br[2] wl[169] vdd gnd cell_6t
Xbit_r170_c2 bl[2] br[2] wl[170] vdd gnd cell_6t
Xbit_r171_c2 bl[2] br[2] wl[171] vdd gnd cell_6t
Xbit_r172_c2 bl[2] br[2] wl[172] vdd gnd cell_6t
Xbit_r173_c2 bl[2] br[2] wl[173] vdd gnd cell_6t
Xbit_r174_c2 bl[2] br[2] wl[174] vdd gnd cell_6t
Xbit_r175_c2 bl[2] br[2] wl[175] vdd gnd cell_6t
Xbit_r176_c2 bl[2] br[2] wl[176] vdd gnd cell_6t
Xbit_r177_c2 bl[2] br[2] wl[177] vdd gnd cell_6t
Xbit_r178_c2 bl[2] br[2] wl[178] vdd gnd cell_6t
Xbit_r179_c2 bl[2] br[2] wl[179] vdd gnd cell_6t
Xbit_r180_c2 bl[2] br[2] wl[180] vdd gnd cell_6t
Xbit_r181_c2 bl[2] br[2] wl[181] vdd gnd cell_6t
Xbit_r182_c2 bl[2] br[2] wl[182] vdd gnd cell_6t
Xbit_r183_c2 bl[2] br[2] wl[183] vdd gnd cell_6t
Xbit_r184_c2 bl[2] br[2] wl[184] vdd gnd cell_6t
Xbit_r185_c2 bl[2] br[2] wl[185] vdd gnd cell_6t
Xbit_r186_c2 bl[2] br[2] wl[186] vdd gnd cell_6t
Xbit_r187_c2 bl[2] br[2] wl[187] vdd gnd cell_6t
Xbit_r188_c2 bl[2] br[2] wl[188] vdd gnd cell_6t
Xbit_r189_c2 bl[2] br[2] wl[189] vdd gnd cell_6t
Xbit_r190_c2 bl[2] br[2] wl[190] vdd gnd cell_6t
Xbit_r191_c2 bl[2] br[2] wl[191] vdd gnd cell_6t
Xbit_r192_c2 bl[2] br[2] wl[192] vdd gnd cell_6t
Xbit_r193_c2 bl[2] br[2] wl[193] vdd gnd cell_6t
Xbit_r194_c2 bl[2] br[2] wl[194] vdd gnd cell_6t
Xbit_r195_c2 bl[2] br[2] wl[195] vdd gnd cell_6t
Xbit_r196_c2 bl[2] br[2] wl[196] vdd gnd cell_6t
Xbit_r197_c2 bl[2] br[2] wl[197] vdd gnd cell_6t
Xbit_r198_c2 bl[2] br[2] wl[198] vdd gnd cell_6t
Xbit_r199_c2 bl[2] br[2] wl[199] vdd gnd cell_6t
Xbit_r200_c2 bl[2] br[2] wl[200] vdd gnd cell_6t
Xbit_r201_c2 bl[2] br[2] wl[201] vdd gnd cell_6t
Xbit_r202_c2 bl[2] br[2] wl[202] vdd gnd cell_6t
Xbit_r203_c2 bl[2] br[2] wl[203] vdd gnd cell_6t
Xbit_r204_c2 bl[2] br[2] wl[204] vdd gnd cell_6t
Xbit_r205_c2 bl[2] br[2] wl[205] vdd gnd cell_6t
Xbit_r206_c2 bl[2] br[2] wl[206] vdd gnd cell_6t
Xbit_r207_c2 bl[2] br[2] wl[207] vdd gnd cell_6t
Xbit_r208_c2 bl[2] br[2] wl[208] vdd gnd cell_6t
Xbit_r209_c2 bl[2] br[2] wl[209] vdd gnd cell_6t
Xbit_r210_c2 bl[2] br[2] wl[210] vdd gnd cell_6t
Xbit_r211_c2 bl[2] br[2] wl[211] vdd gnd cell_6t
Xbit_r212_c2 bl[2] br[2] wl[212] vdd gnd cell_6t
Xbit_r213_c2 bl[2] br[2] wl[213] vdd gnd cell_6t
Xbit_r214_c2 bl[2] br[2] wl[214] vdd gnd cell_6t
Xbit_r215_c2 bl[2] br[2] wl[215] vdd gnd cell_6t
Xbit_r216_c2 bl[2] br[2] wl[216] vdd gnd cell_6t
Xbit_r217_c2 bl[2] br[2] wl[217] vdd gnd cell_6t
Xbit_r218_c2 bl[2] br[2] wl[218] vdd gnd cell_6t
Xbit_r219_c2 bl[2] br[2] wl[219] vdd gnd cell_6t
Xbit_r220_c2 bl[2] br[2] wl[220] vdd gnd cell_6t
Xbit_r221_c2 bl[2] br[2] wl[221] vdd gnd cell_6t
Xbit_r222_c2 bl[2] br[2] wl[222] vdd gnd cell_6t
Xbit_r223_c2 bl[2] br[2] wl[223] vdd gnd cell_6t
Xbit_r224_c2 bl[2] br[2] wl[224] vdd gnd cell_6t
Xbit_r225_c2 bl[2] br[2] wl[225] vdd gnd cell_6t
Xbit_r226_c2 bl[2] br[2] wl[226] vdd gnd cell_6t
Xbit_r227_c2 bl[2] br[2] wl[227] vdd gnd cell_6t
Xbit_r228_c2 bl[2] br[2] wl[228] vdd gnd cell_6t
Xbit_r229_c2 bl[2] br[2] wl[229] vdd gnd cell_6t
Xbit_r230_c2 bl[2] br[2] wl[230] vdd gnd cell_6t
Xbit_r231_c2 bl[2] br[2] wl[231] vdd gnd cell_6t
Xbit_r232_c2 bl[2] br[2] wl[232] vdd gnd cell_6t
Xbit_r233_c2 bl[2] br[2] wl[233] vdd gnd cell_6t
Xbit_r234_c2 bl[2] br[2] wl[234] vdd gnd cell_6t
Xbit_r235_c2 bl[2] br[2] wl[235] vdd gnd cell_6t
Xbit_r236_c2 bl[2] br[2] wl[236] vdd gnd cell_6t
Xbit_r237_c2 bl[2] br[2] wl[237] vdd gnd cell_6t
Xbit_r238_c2 bl[2] br[2] wl[238] vdd gnd cell_6t
Xbit_r239_c2 bl[2] br[2] wl[239] vdd gnd cell_6t
Xbit_r240_c2 bl[2] br[2] wl[240] vdd gnd cell_6t
Xbit_r241_c2 bl[2] br[2] wl[241] vdd gnd cell_6t
Xbit_r242_c2 bl[2] br[2] wl[242] vdd gnd cell_6t
Xbit_r243_c2 bl[2] br[2] wl[243] vdd gnd cell_6t
Xbit_r244_c2 bl[2] br[2] wl[244] vdd gnd cell_6t
Xbit_r245_c2 bl[2] br[2] wl[245] vdd gnd cell_6t
Xbit_r246_c2 bl[2] br[2] wl[246] vdd gnd cell_6t
Xbit_r247_c2 bl[2] br[2] wl[247] vdd gnd cell_6t
Xbit_r248_c2 bl[2] br[2] wl[248] vdd gnd cell_6t
Xbit_r249_c2 bl[2] br[2] wl[249] vdd gnd cell_6t
Xbit_r250_c2 bl[2] br[2] wl[250] vdd gnd cell_6t
Xbit_r251_c2 bl[2] br[2] wl[251] vdd gnd cell_6t
Xbit_r252_c2 bl[2] br[2] wl[252] vdd gnd cell_6t
Xbit_r253_c2 bl[2] br[2] wl[253] vdd gnd cell_6t
Xbit_r254_c2 bl[2] br[2] wl[254] vdd gnd cell_6t
Xbit_r255_c2 bl[2] br[2] wl[255] vdd gnd cell_6t
Xbit_r0_c3 bl[3] br[3] wl[0] vdd gnd cell_6t
Xbit_r1_c3 bl[3] br[3] wl[1] vdd gnd cell_6t
Xbit_r2_c3 bl[3] br[3] wl[2] vdd gnd cell_6t
Xbit_r3_c3 bl[3] br[3] wl[3] vdd gnd cell_6t
Xbit_r4_c3 bl[3] br[3] wl[4] vdd gnd cell_6t
Xbit_r5_c3 bl[3] br[3] wl[5] vdd gnd cell_6t
Xbit_r6_c3 bl[3] br[3] wl[6] vdd gnd cell_6t
Xbit_r7_c3 bl[3] br[3] wl[7] vdd gnd cell_6t
Xbit_r8_c3 bl[3] br[3] wl[8] vdd gnd cell_6t
Xbit_r9_c3 bl[3] br[3] wl[9] vdd gnd cell_6t
Xbit_r10_c3 bl[3] br[3] wl[10] vdd gnd cell_6t
Xbit_r11_c3 bl[3] br[3] wl[11] vdd gnd cell_6t
Xbit_r12_c3 bl[3] br[3] wl[12] vdd gnd cell_6t
Xbit_r13_c3 bl[3] br[3] wl[13] vdd gnd cell_6t
Xbit_r14_c3 bl[3] br[3] wl[14] vdd gnd cell_6t
Xbit_r15_c3 bl[3] br[3] wl[15] vdd gnd cell_6t
Xbit_r16_c3 bl[3] br[3] wl[16] vdd gnd cell_6t
Xbit_r17_c3 bl[3] br[3] wl[17] vdd gnd cell_6t
Xbit_r18_c3 bl[3] br[3] wl[18] vdd gnd cell_6t
Xbit_r19_c3 bl[3] br[3] wl[19] vdd gnd cell_6t
Xbit_r20_c3 bl[3] br[3] wl[20] vdd gnd cell_6t
Xbit_r21_c3 bl[3] br[3] wl[21] vdd gnd cell_6t
Xbit_r22_c3 bl[3] br[3] wl[22] vdd gnd cell_6t
Xbit_r23_c3 bl[3] br[3] wl[23] vdd gnd cell_6t
Xbit_r24_c3 bl[3] br[3] wl[24] vdd gnd cell_6t
Xbit_r25_c3 bl[3] br[3] wl[25] vdd gnd cell_6t
Xbit_r26_c3 bl[3] br[3] wl[26] vdd gnd cell_6t
Xbit_r27_c3 bl[3] br[3] wl[27] vdd gnd cell_6t
Xbit_r28_c3 bl[3] br[3] wl[28] vdd gnd cell_6t
Xbit_r29_c3 bl[3] br[3] wl[29] vdd gnd cell_6t
Xbit_r30_c3 bl[3] br[3] wl[30] vdd gnd cell_6t
Xbit_r31_c3 bl[3] br[3] wl[31] vdd gnd cell_6t
Xbit_r32_c3 bl[3] br[3] wl[32] vdd gnd cell_6t
Xbit_r33_c3 bl[3] br[3] wl[33] vdd gnd cell_6t
Xbit_r34_c3 bl[3] br[3] wl[34] vdd gnd cell_6t
Xbit_r35_c3 bl[3] br[3] wl[35] vdd gnd cell_6t
Xbit_r36_c3 bl[3] br[3] wl[36] vdd gnd cell_6t
Xbit_r37_c3 bl[3] br[3] wl[37] vdd gnd cell_6t
Xbit_r38_c3 bl[3] br[3] wl[38] vdd gnd cell_6t
Xbit_r39_c3 bl[3] br[3] wl[39] vdd gnd cell_6t
Xbit_r40_c3 bl[3] br[3] wl[40] vdd gnd cell_6t
Xbit_r41_c3 bl[3] br[3] wl[41] vdd gnd cell_6t
Xbit_r42_c3 bl[3] br[3] wl[42] vdd gnd cell_6t
Xbit_r43_c3 bl[3] br[3] wl[43] vdd gnd cell_6t
Xbit_r44_c3 bl[3] br[3] wl[44] vdd gnd cell_6t
Xbit_r45_c3 bl[3] br[3] wl[45] vdd gnd cell_6t
Xbit_r46_c3 bl[3] br[3] wl[46] vdd gnd cell_6t
Xbit_r47_c3 bl[3] br[3] wl[47] vdd gnd cell_6t
Xbit_r48_c3 bl[3] br[3] wl[48] vdd gnd cell_6t
Xbit_r49_c3 bl[3] br[3] wl[49] vdd gnd cell_6t
Xbit_r50_c3 bl[3] br[3] wl[50] vdd gnd cell_6t
Xbit_r51_c3 bl[3] br[3] wl[51] vdd gnd cell_6t
Xbit_r52_c3 bl[3] br[3] wl[52] vdd gnd cell_6t
Xbit_r53_c3 bl[3] br[3] wl[53] vdd gnd cell_6t
Xbit_r54_c3 bl[3] br[3] wl[54] vdd gnd cell_6t
Xbit_r55_c3 bl[3] br[3] wl[55] vdd gnd cell_6t
Xbit_r56_c3 bl[3] br[3] wl[56] vdd gnd cell_6t
Xbit_r57_c3 bl[3] br[3] wl[57] vdd gnd cell_6t
Xbit_r58_c3 bl[3] br[3] wl[58] vdd gnd cell_6t
Xbit_r59_c3 bl[3] br[3] wl[59] vdd gnd cell_6t
Xbit_r60_c3 bl[3] br[3] wl[60] vdd gnd cell_6t
Xbit_r61_c3 bl[3] br[3] wl[61] vdd gnd cell_6t
Xbit_r62_c3 bl[3] br[3] wl[62] vdd gnd cell_6t
Xbit_r63_c3 bl[3] br[3] wl[63] vdd gnd cell_6t
Xbit_r64_c3 bl[3] br[3] wl[64] vdd gnd cell_6t
Xbit_r65_c3 bl[3] br[3] wl[65] vdd gnd cell_6t
Xbit_r66_c3 bl[3] br[3] wl[66] vdd gnd cell_6t
Xbit_r67_c3 bl[3] br[3] wl[67] vdd gnd cell_6t
Xbit_r68_c3 bl[3] br[3] wl[68] vdd gnd cell_6t
Xbit_r69_c3 bl[3] br[3] wl[69] vdd gnd cell_6t
Xbit_r70_c3 bl[3] br[3] wl[70] vdd gnd cell_6t
Xbit_r71_c3 bl[3] br[3] wl[71] vdd gnd cell_6t
Xbit_r72_c3 bl[3] br[3] wl[72] vdd gnd cell_6t
Xbit_r73_c3 bl[3] br[3] wl[73] vdd gnd cell_6t
Xbit_r74_c3 bl[3] br[3] wl[74] vdd gnd cell_6t
Xbit_r75_c3 bl[3] br[3] wl[75] vdd gnd cell_6t
Xbit_r76_c3 bl[3] br[3] wl[76] vdd gnd cell_6t
Xbit_r77_c3 bl[3] br[3] wl[77] vdd gnd cell_6t
Xbit_r78_c3 bl[3] br[3] wl[78] vdd gnd cell_6t
Xbit_r79_c3 bl[3] br[3] wl[79] vdd gnd cell_6t
Xbit_r80_c3 bl[3] br[3] wl[80] vdd gnd cell_6t
Xbit_r81_c3 bl[3] br[3] wl[81] vdd gnd cell_6t
Xbit_r82_c3 bl[3] br[3] wl[82] vdd gnd cell_6t
Xbit_r83_c3 bl[3] br[3] wl[83] vdd gnd cell_6t
Xbit_r84_c3 bl[3] br[3] wl[84] vdd gnd cell_6t
Xbit_r85_c3 bl[3] br[3] wl[85] vdd gnd cell_6t
Xbit_r86_c3 bl[3] br[3] wl[86] vdd gnd cell_6t
Xbit_r87_c3 bl[3] br[3] wl[87] vdd gnd cell_6t
Xbit_r88_c3 bl[3] br[3] wl[88] vdd gnd cell_6t
Xbit_r89_c3 bl[3] br[3] wl[89] vdd gnd cell_6t
Xbit_r90_c3 bl[3] br[3] wl[90] vdd gnd cell_6t
Xbit_r91_c3 bl[3] br[3] wl[91] vdd gnd cell_6t
Xbit_r92_c3 bl[3] br[3] wl[92] vdd gnd cell_6t
Xbit_r93_c3 bl[3] br[3] wl[93] vdd gnd cell_6t
Xbit_r94_c3 bl[3] br[3] wl[94] vdd gnd cell_6t
Xbit_r95_c3 bl[3] br[3] wl[95] vdd gnd cell_6t
Xbit_r96_c3 bl[3] br[3] wl[96] vdd gnd cell_6t
Xbit_r97_c3 bl[3] br[3] wl[97] vdd gnd cell_6t
Xbit_r98_c3 bl[3] br[3] wl[98] vdd gnd cell_6t
Xbit_r99_c3 bl[3] br[3] wl[99] vdd gnd cell_6t
Xbit_r100_c3 bl[3] br[3] wl[100] vdd gnd cell_6t
Xbit_r101_c3 bl[3] br[3] wl[101] vdd gnd cell_6t
Xbit_r102_c3 bl[3] br[3] wl[102] vdd gnd cell_6t
Xbit_r103_c3 bl[3] br[3] wl[103] vdd gnd cell_6t
Xbit_r104_c3 bl[3] br[3] wl[104] vdd gnd cell_6t
Xbit_r105_c3 bl[3] br[3] wl[105] vdd gnd cell_6t
Xbit_r106_c3 bl[3] br[3] wl[106] vdd gnd cell_6t
Xbit_r107_c3 bl[3] br[3] wl[107] vdd gnd cell_6t
Xbit_r108_c3 bl[3] br[3] wl[108] vdd gnd cell_6t
Xbit_r109_c3 bl[3] br[3] wl[109] vdd gnd cell_6t
Xbit_r110_c3 bl[3] br[3] wl[110] vdd gnd cell_6t
Xbit_r111_c3 bl[3] br[3] wl[111] vdd gnd cell_6t
Xbit_r112_c3 bl[3] br[3] wl[112] vdd gnd cell_6t
Xbit_r113_c3 bl[3] br[3] wl[113] vdd gnd cell_6t
Xbit_r114_c3 bl[3] br[3] wl[114] vdd gnd cell_6t
Xbit_r115_c3 bl[3] br[3] wl[115] vdd gnd cell_6t
Xbit_r116_c3 bl[3] br[3] wl[116] vdd gnd cell_6t
Xbit_r117_c3 bl[3] br[3] wl[117] vdd gnd cell_6t
Xbit_r118_c3 bl[3] br[3] wl[118] vdd gnd cell_6t
Xbit_r119_c3 bl[3] br[3] wl[119] vdd gnd cell_6t
Xbit_r120_c3 bl[3] br[3] wl[120] vdd gnd cell_6t
Xbit_r121_c3 bl[3] br[3] wl[121] vdd gnd cell_6t
Xbit_r122_c3 bl[3] br[3] wl[122] vdd gnd cell_6t
Xbit_r123_c3 bl[3] br[3] wl[123] vdd gnd cell_6t
Xbit_r124_c3 bl[3] br[3] wl[124] vdd gnd cell_6t
Xbit_r125_c3 bl[3] br[3] wl[125] vdd gnd cell_6t
Xbit_r126_c3 bl[3] br[3] wl[126] vdd gnd cell_6t
Xbit_r127_c3 bl[3] br[3] wl[127] vdd gnd cell_6t
Xbit_r128_c3 bl[3] br[3] wl[128] vdd gnd cell_6t
Xbit_r129_c3 bl[3] br[3] wl[129] vdd gnd cell_6t
Xbit_r130_c3 bl[3] br[3] wl[130] vdd gnd cell_6t
Xbit_r131_c3 bl[3] br[3] wl[131] vdd gnd cell_6t
Xbit_r132_c3 bl[3] br[3] wl[132] vdd gnd cell_6t
Xbit_r133_c3 bl[3] br[3] wl[133] vdd gnd cell_6t
Xbit_r134_c3 bl[3] br[3] wl[134] vdd gnd cell_6t
Xbit_r135_c3 bl[3] br[3] wl[135] vdd gnd cell_6t
Xbit_r136_c3 bl[3] br[3] wl[136] vdd gnd cell_6t
Xbit_r137_c3 bl[3] br[3] wl[137] vdd gnd cell_6t
Xbit_r138_c3 bl[3] br[3] wl[138] vdd gnd cell_6t
Xbit_r139_c3 bl[3] br[3] wl[139] vdd gnd cell_6t
Xbit_r140_c3 bl[3] br[3] wl[140] vdd gnd cell_6t
Xbit_r141_c3 bl[3] br[3] wl[141] vdd gnd cell_6t
Xbit_r142_c3 bl[3] br[3] wl[142] vdd gnd cell_6t
Xbit_r143_c3 bl[3] br[3] wl[143] vdd gnd cell_6t
Xbit_r144_c3 bl[3] br[3] wl[144] vdd gnd cell_6t
Xbit_r145_c3 bl[3] br[3] wl[145] vdd gnd cell_6t
Xbit_r146_c3 bl[3] br[3] wl[146] vdd gnd cell_6t
Xbit_r147_c3 bl[3] br[3] wl[147] vdd gnd cell_6t
Xbit_r148_c3 bl[3] br[3] wl[148] vdd gnd cell_6t
Xbit_r149_c3 bl[3] br[3] wl[149] vdd gnd cell_6t
Xbit_r150_c3 bl[3] br[3] wl[150] vdd gnd cell_6t
Xbit_r151_c3 bl[3] br[3] wl[151] vdd gnd cell_6t
Xbit_r152_c3 bl[3] br[3] wl[152] vdd gnd cell_6t
Xbit_r153_c3 bl[3] br[3] wl[153] vdd gnd cell_6t
Xbit_r154_c3 bl[3] br[3] wl[154] vdd gnd cell_6t
Xbit_r155_c3 bl[3] br[3] wl[155] vdd gnd cell_6t
Xbit_r156_c3 bl[3] br[3] wl[156] vdd gnd cell_6t
Xbit_r157_c3 bl[3] br[3] wl[157] vdd gnd cell_6t
Xbit_r158_c3 bl[3] br[3] wl[158] vdd gnd cell_6t
Xbit_r159_c3 bl[3] br[3] wl[159] vdd gnd cell_6t
Xbit_r160_c3 bl[3] br[3] wl[160] vdd gnd cell_6t
Xbit_r161_c3 bl[3] br[3] wl[161] vdd gnd cell_6t
Xbit_r162_c3 bl[3] br[3] wl[162] vdd gnd cell_6t
Xbit_r163_c3 bl[3] br[3] wl[163] vdd gnd cell_6t
Xbit_r164_c3 bl[3] br[3] wl[164] vdd gnd cell_6t
Xbit_r165_c3 bl[3] br[3] wl[165] vdd gnd cell_6t
Xbit_r166_c3 bl[3] br[3] wl[166] vdd gnd cell_6t
Xbit_r167_c3 bl[3] br[3] wl[167] vdd gnd cell_6t
Xbit_r168_c3 bl[3] br[3] wl[168] vdd gnd cell_6t
Xbit_r169_c3 bl[3] br[3] wl[169] vdd gnd cell_6t
Xbit_r170_c3 bl[3] br[3] wl[170] vdd gnd cell_6t
Xbit_r171_c3 bl[3] br[3] wl[171] vdd gnd cell_6t
Xbit_r172_c3 bl[3] br[3] wl[172] vdd gnd cell_6t
Xbit_r173_c3 bl[3] br[3] wl[173] vdd gnd cell_6t
Xbit_r174_c3 bl[3] br[3] wl[174] vdd gnd cell_6t
Xbit_r175_c3 bl[3] br[3] wl[175] vdd gnd cell_6t
Xbit_r176_c3 bl[3] br[3] wl[176] vdd gnd cell_6t
Xbit_r177_c3 bl[3] br[3] wl[177] vdd gnd cell_6t
Xbit_r178_c3 bl[3] br[3] wl[178] vdd gnd cell_6t
Xbit_r179_c3 bl[3] br[3] wl[179] vdd gnd cell_6t
Xbit_r180_c3 bl[3] br[3] wl[180] vdd gnd cell_6t
Xbit_r181_c3 bl[3] br[3] wl[181] vdd gnd cell_6t
Xbit_r182_c3 bl[3] br[3] wl[182] vdd gnd cell_6t
Xbit_r183_c3 bl[3] br[3] wl[183] vdd gnd cell_6t
Xbit_r184_c3 bl[3] br[3] wl[184] vdd gnd cell_6t
Xbit_r185_c3 bl[3] br[3] wl[185] vdd gnd cell_6t
Xbit_r186_c3 bl[3] br[3] wl[186] vdd gnd cell_6t
Xbit_r187_c3 bl[3] br[3] wl[187] vdd gnd cell_6t
Xbit_r188_c3 bl[3] br[3] wl[188] vdd gnd cell_6t
Xbit_r189_c3 bl[3] br[3] wl[189] vdd gnd cell_6t
Xbit_r190_c3 bl[3] br[3] wl[190] vdd gnd cell_6t
Xbit_r191_c3 bl[3] br[3] wl[191] vdd gnd cell_6t
Xbit_r192_c3 bl[3] br[3] wl[192] vdd gnd cell_6t
Xbit_r193_c3 bl[3] br[3] wl[193] vdd gnd cell_6t
Xbit_r194_c3 bl[3] br[3] wl[194] vdd gnd cell_6t
Xbit_r195_c3 bl[3] br[3] wl[195] vdd gnd cell_6t
Xbit_r196_c3 bl[3] br[3] wl[196] vdd gnd cell_6t
Xbit_r197_c3 bl[3] br[3] wl[197] vdd gnd cell_6t
Xbit_r198_c3 bl[3] br[3] wl[198] vdd gnd cell_6t
Xbit_r199_c3 bl[3] br[3] wl[199] vdd gnd cell_6t
Xbit_r200_c3 bl[3] br[3] wl[200] vdd gnd cell_6t
Xbit_r201_c3 bl[3] br[3] wl[201] vdd gnd cell_6t
Xbit_r202_c3 bl[3] br[3] wl[202] vdd gnd cell_6t
Xbit_r203_c3 bl[3] br[3] wl[203] vdd gnd cell_6t
Xbit_r204_c3 bl[3] br[3] wl[204] vdd gnd cell_6t
Xbit_r205_c3 bl[3] br[3] wl[205] vdd gnd cell_6t
Xbit_r206_c3 bl[3] br[3] wl[206] vdd gnd cell_6t
Xbit_r207_c3 bl[3] br[3] wl[207] vdd gnd cell_6t
Xbit_r208_c3 bl[3] br[3] wl[208] vdd gnd cell_6t
Xbit_r209_c3 bl[3] br[3] wl[209] vdd gnd cell_6t
Xbit_r210_c3 bl[3] br[3] wl[210] vdd gnd cell_6t
Xbit_r211_c3 bl[3] br[3] wl[211] vdd gnd cell_6t
Xbit_r212_c3 bl[3] br[3] wl[212] vdd gnd cell_6t
Xbit_r213_c3 bl[3] br[3] wl[213] vdd gnd cell_6t
Xbit_r214_c3 bl[3] br[3] wl[214] vdd gnd cell_6t
Xbit_r215_c3 bl[3] br[3] wl[215] vdd gnd cell_6t
Xbit_r216_c3 bl[3] br[3] wl[216] vdd gnd cell_6t
Xbit_r217_c3 bl[3] br[3] wl[217] vdd gnd cell_6t
Xbit_r218_c3 bl[3] br[3] wl[218] vdd gnd cell_6t
Xbit_r219_c3 bl[3] br[3] wl[219] vdd gnd cell_6t
Xbit_r220_c3 bl[3] br[3] wl[220] vdd gnd cell_6t
Xbit_r221_c3 bl[3] br[3] wl[221] vdd gnd cell_6t
Xbit_r222_c3 bl[3] br[3] wl[222] vdd gnd cell_6t
Xbit_r223_c3 bl[3] br[3] wl[223] vdd gnd cell_6t
Xbit_r224_c3 bl[3] br[3] wl[224] vdd gnd cell_6t
Xbit_r225_c3 bl[3] br[3] wl[225] vdd gnd cell_6t
Xbit_r226_c3 bl[3] br[3] wl[226] vdd gnd cell_6t
Xbit_r227_c3 bl[3] br[3] wl[227] vdd gnd cell_6t
Xbit_r228_c3 bl[3] br[3] wl[228] vdd gnd cell_6t
Xbit_r229_c3 bl[3] br[3] wl[229] vdd gnd cell_6t
Xbit_r230_c3 bl[3] br[3] wl[230] vdd gnd cell_6t
Xbit_r231_c3 bl[3] br[3] wl[231] vdd gnd cell_6t
Xbit_r232_c3 bl[3] br[3] wl[232] vdd gnd cell_6t
Xbit_r233_c3 bl[3] br[3] wl[233] vdd gnd cell_6t
Xbit_r234_c3 bl[3] br[3] wl[234] vdd gnd cell_6t
Xbit_r235_c3 bl[3] br[3] wl[235] vdd gnd cell_6t
Xbit_r236_c3 bl[3] br[3] wl[236] vdd gnd cell_6t
Xbit_r237_c3 bl[3] br[3] wl[237] vdd gnd cell_6t
Xbit_r238_c3 bl[3] br[3] wl[238] vdd gnd cell_6t
Xbit_r239_c3 bl[3] br[3] wl[239] vdd gnd cell_6t
Xbit_r240_c3 bl[3] br[3] wl[240] vdd gnd cell_6t
Xbit_r241_c3 bl[3] br[3] wl[241] vdd gnd cell_6t
Xbit_r242_c3 bl[3] br[3] wl[242] vdd gnd cell_6t
Xbit_r243_c3 bl[3] br[3] wl[243] vdd gnd cell_6t
Xbit_r244_c3 bl[3] br[3] wl[244] vdd gnd cell_6t
Xbit_r245_c3 bl[3] br[3] wl[245] vdd gnd cell_6t
Xbit_r246_c3 bl[3] br[3] wl[246] vdd gnd cell_6t
Xbit_r247_c3 bl[3] br[3] wl[247] vdd gnd cell_6t
Xbit_r248_c3 bl[3] br[3] wl[248] vdd gnd cell_6t
Xbit_r249_c3 bl[3] br[3] wl[249] vdd gnd cell_6t
Xbit_r250_c3 bl[3] br[3] wl[250] vdd gnd cell_6t
Xbit_r251_c3 bl[3] br[3] wl[251] vdd gnd cell_6t
Xbit_r252_c3 bl[3] br[3] wl[252] vdd gnd cell_6t
Xbit_r253_c3 bl[3] br[3] wl[253] vdd gnd cell_6t
Xbit_r254_c3 bl[3] br[3] wl[254] vdd gnd cell_6t
Xbit_r255_c3 bl[3] br[3] wl[255] vdd gnd cell_6t
Xbit_r0_c4 bl[4] br[4] wl[0] vdd gnd cell_6t
Xbit_r1_c4 bl[4] br[4] wl[1] vdd gnd cell_6t
Xbit_r2_c4 bl[4] br[4] wl[2] vdd gnd cell_6t
Xbit_r3_c4 bl[4] br[4] wl[3] vdd gnd cell_6t
Xbit_r4_c4 bl[4] br[4] wl[4] vdd gnd cell_6t
Xbit_r5_c4 bl[4] br[4] wl[5] vdd gnd cell_6t
Xbit_r6_c4 bl[4] br[4] wl[6] vdd gnd cell_6t
Xbit_r7_c4 bl[4] br[4] wl[7] vdd gnd cell_6t
Xbit_r8_c4 bl[4] br[4] wl[8] vdd gnd cell_6t
Xbit_r9_c4 bl[4] br[4] wl[9] vdd gnd cell_6t
Xbit_r10_c4 bl[4] br[4] wl[10] vdd gnd cell_6t
Xbit_r11_c4 bl[4] br[4] wl[11] vdd gnd cell_6t
Xbit_r12_c4 bl[4] br[4] wl[12] vdd gnd cell_6t
Xbit_r13_c4 bl[4] br[4] wl[13] vdd gnd cell_6t
Xbit_r14_c4 bl[4] br[4] wl[14] vdd gnd cell_6t
Xbit_r15_c4 bl[4] br[4] wl[15] vdd gnd cell_6t
Xbit_r16_c4 bl[4] br[4] wl[16] vdd gnd cell_6t
Xbit_r17_c4 bl[4] br[4] wl[17] vdd gnd cell_6t
Xbit_r18_c4 bl[4] br[4] wl[18] vdd gnd cell_6t
Xbit_r19_c4 bl[4] br[4] wl[19] vdd gnd cell_6t
Xbit_r20_c4 bl[4] br[4] wl[20] vdd gnd cell_6t
Xbit_r21_c4 bl[4] br[4] wl[21] vdd gnd cell_6t
Xbit_r22_c4 bl[4] br[4] wl[22] vdd gnd cell_6t
Xbit_r23_c4 bl[4] br[4] wl[23] vdd gnd cell_6t
Xbit_r24_c4 bl[4] br[4] wl[24] vdd gnd cell_6t
Xbit_r25_c4 bl[4] br[4] wl[25] vdd gnd cell_6t
Xbit_r26_c4 bl[4] br[4] wl[26] vdd gnd cell_6t
Xbit_r27_c4 bl[4] br[4] wl[27] vdd gnd cell_6t
Xbit_r28_c4 bl[4] br[4] wl[28] vdd gnd cell_6t
Xbit_r29_c4 bl[4] br[4] wl[29] vdd gnd cell_6t
Xbit_r30_c4 bl[4] br[4] wl[30] vdd gnd cell_6t
Xbit_r31_c4 bl[4] br[4] wl[31] vdd gnd cell_6t
Xbit_r32_c4 bl[4] br[4] wl[32] vdd gnd cell_6t
Xbit_r33_c4 bl[4] br[4] wl[33] vdd gnd cell_6t
Xbit_r34_c4 bl[4] br[4] wl[34] vdd gnd cell_6t
Xbit_r35_c4 bl[4] br[4] wl[35] vdd gnd cell_6t
Xbit_r36_c4 bl[4] br[4] wl[36] vdd gnd cell_6t
Xbit_r37_c4 bl[4] br[4] wl[37] vdd gnd cell_6t
Xbit_r38_c4 bl[4] br[4] wl[38] vdd gnd cell_6t
Xbit_r39_c4 bl[4] br[4] wl[39] vdd gnd cell_6t
Xbit_r40_c4 bl[4] br[4] wl[40] vdd gnd cell_6t
Xbit_r41_c4 bl[4] br[4] wl[41] vdd gnd cell_6t
Xbit_r42_c4 bl[4] br[4] wl[42] vdd gnd cell_6t
Xbit_r43_c4 bl[4] br[4] wl[43] vdd gnd cell_6t
Xbit_r44_c4 bl[4] br[4] wl[44] vdd gnd cell_6t
Xbit_r45_c4 bl[4] br[4] wl[45] vdd gnd cell_6t
Xbit_r46_c4 bl[4] br[4] wl[46] vdd gnd cell_6t
Xbit_r47_c4 bl[4] br[4] wl[47] vdd gnd cell_6t
Xbit_r48_c4 bl[4] br[4] wl[48] vdd gnd cell_6t
Xbit_r49_c4 bl[4] br[4] wl[49] vdd gnd cell_6t
Xbit_r50_c4 bl[4] br[4] wl[50] vdd gnd cell_6t
Xbit_r51_c4 bl[4] br[4] wl[51] vdd gnd cell_6t
Xbit_r52_c4 bl[4] br[4] wl[52] vdd gnd cell_6t
Xbit_r53_c4 bl[4] br[4] wl[53] vdd gnd cell_6t
Xbit_r54_c4 bl[4] br[4] wl[54] vdd gnd cell_6t
Xbit_r55_c4 bl[4] br[4] wl[55] vdd gnd cell_6t
Xbit_r56_c4 bl[4] br[4] wl[56] vdd gnd cell_6t
Xbit_r57_c4 bl[4] br[4] wl[57] vdd gnd cell_6t
Xbit_r58_c4 bl[4] br[4] wl[58] vdd gnd cell_6t
Xbit_r59_c4 bl[4] br[4] wl[59] vdd gnd cell_6t
Xbit_r60_c4 bl[4] br[4] wl[60] vdd gnd cell_6t
Xbit_r61_c4 bl[4] br[4] wl[61] vdd gnd cell_6t
Xbit_r62_c4 bl[4] br[4] wl[62] vdd gnd cell_6t
Xbit_r63_c4 bl[4] br[4] wl[63] vdd gnd cell_6t
Xbit_r64_c4 bl[4] br[4] wl[64] vdd gnd cell_6t
Xbit_r65_c4 bl[4] br[4] wl[65] vdd gnd cell_6t
Xbit_r66_c4 bl[4] br[4] wl[66] vdd gnd cell_6t
Xbit_r67_c4 bl[4] br[4] wl[67] vdd gnd cell_6t
Xbit_r68_c4 bl[4] br[4] wl[68] vdd gnd cell_6t
Xbit_r69_c4 bl[4] br[4] wl[69] vdd gnd cell_6t
Xbit_r70_c4 bl[4] br[4] wl[70] vdd gnd cell_6t
Xbit_r71_c4 bl[4] br[4] wl[71] vdd gnd cell_6t
Xbit_r72_c4 bl[4] br[4] wl[72] vdd gnd cell_6t
Xbit_r73_c4 bl[4] br[4] wl[73] vdd gnd cell_6t
Xbit_r74_c4 bl[4] br[4] wl[74] vdd gnd cell_6t
Xbit_r75_c4 bl[4] br[4] wl[75] vdd gnd cell_6t
Xbit_r76_c4 bl[4] br[4] wl[76] vdd gnd cell_6t
Xbit_r77_c4 bl[4] br[4] wl[77] vdd gnd cell_6t
Xbit_r78_c4 bl[4] br[4] wl[78] vdd gnd cell_6t
Xbit_r79_c4 bl[4] br[4] wl[79] vdd gnd cell_6t
Xbit_r80_c4 bl[4] br[4] wl[80] vdd gnd cell_6t
Xbit_r81_c4 bl[4] br[4] wl[81] vdd gnd cell_6t
Xbit_r82_c4 bl[4] br[4] wl[82] vdd gnd cell_6t
Xbit_r83_c4 bl[4] br[4] wl[83] vdd gnd cell_6t
Xbit_r84_c4 bl[4] br[4] wl[84] vdd gnd cell_6t
Xbit_r85_c4 bl[4] br[4] wl[85] vdd gnd cell_6t
Xbit_r86_c4 bl[4] br[4] wl[86] vdd gnd cell_6t
Xbit_r87_c4 bl[4] br[4] wl[87] vdd gnd cell_6t
Xbit_r88_c4 bl[4] br[4] wl[88] vdd gnd cell_6t
Xbit_r89_c4 bl[4] br[4] wl[89] vdd gnd cell_6t
Xbit_r90_c4 bl[4] br[4] wl[90] vdd gnd cell_6t
Xbit_r91_c4 bl[4] br[4] wl[91] vdd gnd cell_6t
Xbit_r92_c4 bl[4] br[4] wl[92] vdd gnd cell_6t
Xbit_r93_c4 bl[4] br[4] wl[93] vdd gnd cell_6t
Xbit_r94_c4 bl[4] br[4] wl[94] vdd gnd cell_6t
Xbit_r95_c4 bl[4] br[4] wl[95] vdd gnd cell_6t
Xbit_r96_c4 bl[4] br[4] wl[96] vdd gnd cell_6t
Xbit_r97_c4 bl[4] br[4] wl[97] vdd gnd cell_6t
Xbit_r98_c4 bl[4] br[4] wl[98] vdd gnd cell_6t
Xbit_r99_c4 bl[4] br[4] wl[99] vdd gnd cell_6t
Xbit_r100_c4 bl[4] br[4] wl[100] vdd gnd cell_6t
Xbit_r101_c4 bl[4] br[4] wl[101] vdd gnd cell_6t
Xbit_r102_c4 bl[4] br[4] wl[102] vdd gnd cell_6t
Xbit_r103_c4 bl[4] br[4] wl[103] vdd gnd cell_6t
Xbit_r104_c4 bl[4] br[4] wl[104] vdd gnd cell_6t
Xbit_r105_c4 bl[4] br[4] wl[105] vdd gnd cell_6t
Xbit_r106_c4 bl[4] br[4] wl[106] vdd gnd cell_6t
Xbit_r107_c4 bl[4] br[4] wl[107] vdd gnd cell_6t
Xbit_r108_c4 bl[4] br[4] wl[108] vdd gnd cell_6t
Xbit_r109_c4 bl[4] br[4] wl[109] vdd gnd cell_6t
Xbit_r110_c4 bl[4] br[4] wl[110] vdd gnd cell_6t
Xbit_r111_c4 bl[4] br[4] wl[111] vdd gnd cell_6t
Xbit_r112_c4 bl[4] br[4] wl[112] vdd gnd cell_6t
Xbit_r113_c4 bl[4] br[4] wl[113] vdd gnd cell_6t
Xbit_r114_c4 bl[4] br[4] wl[114] vdd gnd cell_6t
Xbit_r115_c4 bl[4] br[4] wl[115] vdd gnd cell_6t
Xbit_r116_c4 bl[4] br[4] wl[116] vdd gnd cell_6t
Xbit_r117_c4 bl[4] br[4] wl[117] vdd gnd cell_6t
Xbit_r118_c4 bl[4] br[4] wl[118] vdd gnd cell_6t
Xbit_r119_c4 bl[4] br[4] wl[119] vdd gnd cell_6t
Xbit_r120_c4 bl[4] br[4] wl[120] vdd gnd cell_6t
Xbit_r121_c4 bl[4] br[4] wl[121] vdd gnd cell_6t
Xbit_r122_c4 bl[4] br[4] wl[122] vdd gnd cell_6t
Xbit_r123_c4 bl[4] br[4] wl[123] vdd gnd cell_6t
Xbit_r124_c4 bl[4] br[4] wl[124] vdd gnd cell_6t
Xbit_r125_c4 bl[4] br[4] wl[125] vdd gnd cell_6t
Xbit_r126_c4 bl[4] br[4] wl[126] vdd gnd cell_6t
Xbit_r127_c4 bl[4] br[4] wl[127] vdd gnd cell_6t
Xbit_r128_c4 bl[4] br[4] wl[128] vdd gnd cell_6t
Xbit_r129_c4 bl[4] br[4] wl[129] vdd gnd cell_6t
Xbit_r130_c4 bl[4] br[4] wl[130] vdd gnd cell_6t
Xbit_r131_c4 bl[4] br[4] wl[131] vdd gnd cell_6t
Xbit_r132_c4 bl[4] br[4] wl[132] vdd gnd cell_6t
Xbit_r133_c4 bl[4] br[4] wl[133] vdd gnd cell_6t
Xbit_r134_c4 bl[4] br[4] wl[134] vdd gnd cell_6t
Xbit_r135_c4 bl[4] br[4] wl[135] vdd gnd cell_6t
Xbit_r136_c4 bl[4] br[4] wl[136] vdd gnd cell_6t
Xbit_r137_c4 bl[4] br[4] wl[137] vdd gnd cell_6t
Xbit_r138_c4 bl[4] br[4] wl[138] vdd gnd cell_6t
Xbit_r139_c4 bl[4] br[4] wl[139] vdd gnd cell_6t
Xbit_r140_c4 bl[4] br[4] wl[140] vdd gnd cell_6t
Xbit_r141_c4 bl[4] br[4] wl[141] vdd gnd cell_6t
Xbit_r142_c4 bl[4] br[4] wl[142] vdd gnd cell_6t
Xbit_r143_c4 bl[4] br[4] wl[143] vdd gnd cell_6t
Xbit_r144_c4 bl[4] br[4] wl[144] vdd gnd cell_6t
Xbit_r145_c4 bl[4] br[4] wl[145] vdd gnd cell_6t
Xbit_r146_c4 bl[4] br[4] wl[146] vdd gnd cell_6t
Xbit_r147_c4 bl[4] br[4] wl[147] vdd gnd cell_6t
Xbit_r148_c4 bl[4] br[4] wl[148] vdd gnd cell_6t
Xbit_r149_c4 bl[4] br[4] wl[149] vdd gnd cell_6t
Xbit_r150_c4 bl[4] br[4] wl[150] vdd gnd cell_6t
Xbit_r151_c4 bl[4] br[4] wl[151] vdd gnd cell_6t
Xbit_r152_c4 bl[4] br[4] wl[152] vdd gnd cell_6t
Xbit_r153_c4 bl[4] br[4] wl[153] vdd gnd cell_6t
Xbit_r154_c4 bl[4] br[4] wl[154] vdd gnd cell_6t
Xbit_r155_c4 bl[4] br[4] wl[155] vdd gnd cell_6t
Xbit_r156_c4 bl[4] br[4] wl[156] vdd gnd cell_6t
Xbit_r157_c4 bl[4] br[4] wl[157] vdd gnd cell_6t
Xbit_r158_c4 bl[4] br[4] wl[158] vdd gnd cell_6t
Xbit_r159_c4 bl[4] br[4] wl[159] vdd gnd cell_6t
Xbit_r160_c4 bl[4] br[4] wl[160] vdd gnd cell_6t
Xbit_r161_c4 bl[4] br[4] wl[161] vdd gnd cell_6t
Xbit_r162_c4 bl[4] br[4] wl[162] vdd gnd cell_6t
Xbit_r163_c4 bl[4] br[4] wl[163] vdd gnd cell_6t
Xbit_r164_c4 bl[4] br[4] wl[164] vdd gnd cell_6t
Xbit_r165_c4 bl[4] br[4] wl[165] vdd gnd cell_6t
Xbit_r166_c4 bl[4] br[4] wl[166] vdd gnd cell_6t
Xbit_r167_c4 bl[4] br[4] wl[167] vdd gnd cell_6t
Xbit_r168_c4 bl[4] br[4] wl[168] vdd gnd cell_6t
Xbit_r169_c4 bl[4] br[4] wl[169] vdd gnd cell_6t
Xbit_r170_c4 bl[4] br[4] wl[170] vdd gnd cell_6t
Xbit_r171_c4 bl[4] br[4] wl[171] vdd gnd cell_6t
Xbit_r172_c4 bl[4] br[4] wl[172] vdd gnd cell_6t
Xbit_r173_c4 bl[4] br[4] wl[173] vdd gnd cell_6t
Xbit_r174_c4 bl[4] br[4] wl[174] vdd gnd cell_6t
Xbit_r175_c4 bl[4] br[4] wl[175] vdd gnd cell_6t
Xbit_r176_c4 bl[4] br[4] wl[176] vdd gnd cell_6t
Xbit_r177_c4 bl[4] br[4] wl[177] vdd gnd cell_6t
Xbit_r178_c4 bl[4] br[4] wl[178] vdd gnd cell_6t
Xbit_r179_c4 bl[4] br[4] wl[179] vdd gnd cell_6t
Xbit_r180_c4 bl[4] br[4] wl[180] vdd gnd cell_6t
Xbit_r181_c4 bl[4] br[4] wl[181] vdd gnd cell_6t
Xbit_r182_c4 bl[4] br[4] wl[182] vdd gnd cell_6t
Xbit_r183_c4 bl[4] br[4] wl[183] vdd gnd cell_6t
Xbit_r184_c4 bl[4] br[4] wl[184] vdd gnd cell_6t
Xbit_r185_c4 bl[4] br[4] wl[185] vdd gnd cell_6t
Xbit_r186_c4 bl[4] br[4] wl[186] vdd gnd cell_6t
Xbit_r187_c4 bl[4] br[4] wl[187] vdd gnd cell_6t
Xbit_r188_c4 bl[4] br[4] wl[188] vdd gnd cell_6t
Xbit_r189_c4 bl[4] br[4] wl[189] vdd gnd cell_6t
Xbit_r190_c4 bl[4] br[4] wl[190] vdd gnd cell_6t
Xbit_r191_c4 bl[4] br[4] wl[191] vdd gnd cell_6t
Xbit_r192_c4 bl[4] br[4] wl[192] vdd gnd cell_6t
Xbit_r193_c4 bl[4] br[4] wl[193] vdd gnd cell_6t
Xbit_r194_c4 bl[4] br[4] wl[194] vdd gnd cell_6t
Xbit_r195_c4 bl[4] br[4] wl[195] vdd gnd cell_6t
Xbit_r196_c4 bl[4] br[4] wl[196] vdd gnd cell_6t
Xbit_r197_c4 bl[4] br[4] wl[197] vdd gnd cell_6t
Xbit_r198_c4 bl[4] br[4] wl[198] vdd gnd cell_6t
Xbit_r199_c4 bl[4] br[4] wl[199] vdd gnd cell_6t
Xbit_r200_c4 bl[4] br[4] wl[200] vdd gnd cell_6t
Xbit_r201_c4 bl[4] br[4] wl[201] vdd gnd cell_6t
Xbit_r202_c4 bl[4] br[4] wl[202] vdd gnd cell_6t
Xbit_r203_c4 bl[4] br[4] wl[203] vdd gnd cell_6t
Xbit_r204_c4 bl[4] br[4] wl[204] vdd gnd cell_6t
Xbit_r205_c4 bl[4] br[4] wl[205] vdd gnd cell_6t
Xbit_r206_c4 bl[4] br[4] wl[206] vdd gnd cell_6t
Xbit_r207_c4 bl[4] br[4] wl[207] vdd gnd cell_6t
Xbit_r208_c4 bl[4] br[4] wl[208] vdd gnd cell_6t
Xbit_r209_c4 bl[4] br[4] wl[209] vdd gnd cell_6t
Xbit_r210_c4 bl[4] br[4] wl[210] vdd gnd cell_6t
Xbit_r211_c4 bl[4] br[4] wl[211] vdd gnd cell_6t
Xbit_r212_c4 bl[4] br[4] wl[212] vdd gnd cell_6t
Xbit_r213_c4 bl[4] br[4] wl[213] vdd gnd cell_6t
Xbit_r214_c4 bl[4] br[4] wl[214] vdd gnd cell_6t
Xbit_r215_c4 bl[4] br[4] wl[215] vdd gnd cell_6t
Xbit_r216_c4 bl[4] br[4] wl[216] vdd gnd cell_6t
Xbit_r217_c4 bl[4] br[4] wl[217] vdd gnd cell_6t
Xbit_r218_c4 bl[4] br[4] wl[218] vdd gnd cell_6t
Xbit_r219_c4 bl[4] br[4] wl[219] vdd gnd cell_6t
Xbit_r220_c4 bl[4] br[4] wl[220] vdd gnd cell_6t
Xbit_r221_c4 bl[4] br[4] wl[221] vdd gnd cell_6t
Xbit_r222_c4 bl[4] br[4] wl[222] vdd gnd cell_6t
Xbit_r223_c4 bl[4] br[4] wl[223] vdd gnd cell_6t
Xbit_r224_c4 bl[4] br[4] wl[224] vdd gnd cell_6t
Xbit_r225_c4 bl[4] br[4] wl[225] vdd gnd cell_6t
Xbit_r226_c4 bl[4] br[4] wl[226] vdd gnd cell_6t
Xbit_r227_c4 bl[4] br[4] wl[227] vdd gnd cell_6t
Xbit_r228_c4 bl[4] br[4] wl[228] vdd gnd cell_6t
Xbit_r229_c4 bl[4] br[4] wl[229] vdd gnd cell_6t
Xbit_r230_c4 bl[4] br[4] wl[230] vdd gnd cell_6t
Xbit_r231_c4 bl[4] br[4] wl[231] vdd gnd cell_6t
Xbit_r232_c4 bl[4] br[4] wl[232] vdd gnd cell_6t
Xbit_r233_c4 bl[4] br[4] wl[233] vdd gnd cell_6t
Xbit_r234_c4 bl[4] br[4] wl[234] vdd gnd cell_6t
Xbit_r235_c4 bl[4] br[4] wl[235] vdd gnd cell_6t
Xbit_r236_c4 bl[4] br[4] wl[236] vdd gnd cell_6t
Xbit_r237_c4 bl[4] br[4] wl[237] vdd gnd cell_6t
Xbit_r238_c4 bl[4] br[4] wl[238] vdd gnd cell_6t
Xbit_r239_c4 bl[4] br[4] wl[239] vdd gnd cell_6t
Xbit_r240_c4 bl[4] br[4] wl[240] vdd gnd cell_6t
Xbit_r241_c4 bl[4] br[4] wl[241] vdd gnd cell_6t
Xbit_r242_c4 bl[4] br[4] wl[242] vdd gnd cell_6t
Xbit_r243_c4 bl[4] br[4] wl[243] vdd gnd cell_6t
Xbit_r244_c4 bl[4] br[4] wl[244] vdd gnd cell_6t
Xbit_r245_c4 bl[4] br[4] wl[245] vdd gnd cell_6t
Xbit_r246_c4 bl[4] br[4] wl[246] vdd gnd cell_6t
Xbit_r247_c4 bl[4] br[4] wl[247] vdd gnd cell_6t
Xbit_r248_c4 bl[4] br[4] wl[248] vdd gnd cell_6t
Xbit_r249_c4 bl[4] br[4] wl[249] vdd gnd cell_6t
Xbit_r250_c4 bl[4] br[4] wl[250] vdd gnd cell_6t
Xbit_r251_c4 bl[4] br[4] wl[251] vdd gnd cell_6t
Xbit_r252_c4 bl[4] br[4] wl[252] vdd gnd cell_6t
Xbit_r253_c4 bl[4] br[4] wl[253] vdd gnd cell_6t
Xbit_r254_c4 bl[4] br[4] wl[254] vdd gnd cell_6t
Xbit_r255_c4 bl[4] br[4] wl[255] vdd gnd cell_6t
Xbit_r0_c5 bl[5] br[5] wl[0] vdd gnd cell_6t
Xbit_r1_c5 bl[5] br[5] wl[1] vdd gnd cell_6t
Xbit_r2_c5 bl[5] br[5] wl[2] vdd gnd cell_6t
Xbit_r3_c5 bl[5] br[5] wl[3] vdd gnd cell_6t
Xbit_r4_c5 bl[5] br[5] wl[4] vdd gnd cell_6t
Xbit_r5_c5 bl[5] br[5] wl[5] vdd gnd cell_6t
Xbit_r6_c5 bl[5] br[5] wl[6] vdd gnd cell_6t
Xbit_r7_c5 bl[5] br[5] wl[7] vdd gnd cell_6t
Xbit_r8_c5 bl[5] br[5] wl[8] vdd gnd cell_6t
Xbit_r9_c5 bl[5] br[5] wl[9] vdd gnd cell_6t
Xbit_r10_c5 bl[5] br[5] wl[10] vdd gnd cell_6t
Xbit_r11_c5 bl[5] br[5] wl[11] vdd gnd cell_6t
Xbit_r12_c5 bl[5] br[5] wl[12] vdd gnd cell_6t
Xbit_r13_c5 bl[5] br[5] wl[13] vdd gnd cell_6t
Xbit_r14_c5 bl[5] br[5] wl[14] vdd gnd cell_6t
Xbit_r15_c5 bl[5] br[5] wl[15] vdd gnd cell_6t
Xbit_r16_c5 bl[5] br[5] wl[16] vdd gnd cell_6t
Xbit_r17_c5 bl[5] br[5] wl[17] vdd gnd cell_6t
Xbit_r18_c5 bl[5] br[5] wl[18] vdd gnd cell_6t
Xbit_r19_c5 bl[5] br[5] wl[19] vdd gnd cell_6t
Xbit_r20_c5 bl[5] br[5] wl[20] vdd gnd cell_6t
Xbit_r21_c5 bl[5] br[5] wl[21] vdd gnd cell_6t
Xbit_r22_c5 bl[5] br[5] wl[22] vdd gnd cell_6t
Xbit_r23_c5 bl[5] br[5] wl[23] vdd gnd cell_6t
Xbit_r24_c5 bl[5] br[5] wl[24] vdd gnd cell_6t
Xbit_r25_c5 bl[5] br[5] wl[25] vdd gnd cell_6t
Xbit_r26_c5 bl[5] br[5] wl[26] vdd gnd cell_6t
Xbit_r27_c5 bl[5] br[5] wl[27] vdd gnd cell_6t
Xbit_r28_c5 bl[5] br[5] wl[28] vdd gnd cell_6t
Xbit_r29_c5 bl[5] br[5] wl[29] vdd gnd cell_6t
Xbit_r30_c5 bl[5] br[5] wl[30] vdd gnd cell_6t
Xbit_r31_c5 bl[5] br[5] wl[31] vdd gnd cell_6t
Xbit_r32_c5 bl[5] br[5] wl[32] vdd gnd cell_6t
Xbit_r33_c5 bl[5] br[5] wl[33] vdd gnd cell_6t
Xbit_r34_c5 bl[5] br[5] wl[34] vdd gnd cell_6t
Xbit_r35_c5 bl[5] br[5] wl[35] vdd gnd cell_6t
Xbit_r36_c5 bl[5] br[5] wl[36] vdd gnd cell_6t
Xbit_r37_c5 bl[5] br[5] wl[37] vdd gnd cell_6t
Xbit_r38_c5 bl[5] br[5] wl[38] vdd gnd cell_6t
Xbit_r39_c5 bl[5] br[5] wl[39] vdd gnd cell_6t
Xbit_r40_c5 bl[5] br[5] wl[40] vdd gnd cell_6t
Xbit_r41_c5 bl[5] br[5] wl[41] vdd gnd cell_6t
Xbit_r42_c5 bl[5] br[5] wl[42] vdd gnd cell_6t
Xbit_r43_c5 bl[5] br[5] wl[43] vdd gnd cell_6t
Xbit_r44_c5 bl[5] br[5] wl[44] vdd gnd cell_6t
Xbit_r45_c5 bl[5] br[5] wl[45] vdd gnd cell_6t
Xbit_r46_c5 bl[5] br[5] wl[46] vdd gnd cell_6t
Xbit_r47_c5 bl[5] br[5] wl[47] vdd gnd cell_6t
Xbit_r48_c5 bl[5] br[5] wl[48] vdd gnd cell_6t
Xbit_r49_c5 bl[5] br[5] wl[49] vdd gnd cell_6t
Xbit_r50_c5 bl[5] br[5] wl[50] vdd gnd cell_6t
Xbit_r51_c5 bl[5] br[5] wl[51] vdd gnd cell_6t
Xbit_r52_c5 bl[5] br[5] wl[52] vdd gnd cell_6t
Xbit_r53_c5 bl[5] br[5] wl[53] vdd gnd cell_6t
Xbit_r54_c5 bl[5] br[5] wl[54] vdd gnd cell_6t
Xbit_r55_c5 bl[5] br[5] wl[55] vdd gnd cell_6t
Xbit_r56_c5 bl[5] br[5] wl[56] vdd gnd cell_6t
Xbit_r57_c5 bl[5] br[5] wl[57] vdd gnd cell_6t
Xbit_r58_c5 bl[5] br[5] wl[58] vdd gnd cell_6t
Xbit_r59_c5 bl[5] br[5] wl[59] vdd gnd cell_6t
Xbit_r60_c5 bl[5] br[5] wl[60] vdd gnd cell_6t
Xbit_r61_c5 bl[5] br[5] wl[61] vdd gnd cell_6t
Xbit_r62_c5 bl[5] br[5] wl[62] vdd gnd cell_6t
Xbit_r63_c5 bl[5] br[5] wl[63] vdd gnd cell_6t
Xbit_r64_c5 bl[5] br[5] wl[64] vdd gnd cell_6t
Xbit_r65_c5 bl[5] br[5] wl[65] vdd gnd cell_6t
Xbit_r66_c5 bl[5] br[5] wl[66] vdd gnd cell_6t
Xbit_r67_c5 bl[5] br[5] wl[67] vdd gnd cell_6t
Xbit_r68_c5 bl[5] br[5] wl[68] vdd gnd cell_6t
Xbit_r69_c5 bl[5] br[5] wl[69] vdd gnd cell_6t
Xbit_r70_c5 bl[5] br[5] wl[70] vdd gnd cell_6t
Xbit_r71_c5 bl[5] br[5] wl[71] vdd gnd cell_6t
Xbit_r72_c5 bl[5] br[5] wl[72] vdd gnd cell_6t
Xbit_r73_c5 bl[5] br[5] wl[73] vdd gnd cell_6t
Xbit_r74_c5 bl[5] br[5] wl[74] vdd gnd cell_6t
Xbit_r75_c5 bl[5] br[5] wl[75] vdd gnd cell_6t
Xbit_r76_c5 bl[5] br[5] wl[76] vdd gnd cell_6t
Xbit_r77_c5 bl[5] br[5] wl[77] vdd gnd cell_6t
Xbit_r78_c5 bl[5] br[5] wl[78] vdd gnd cell_6t
Xbit_r79_c5 bl[5] br[5] wl[79] vdd gnd cell_6t
Xbit_r80_c5 bl[5] br[5] wl[80] vdd gnd cell_6t
Xbit_r81_c5 bl[5] br[5] wl[81] vdd gnd cell_6t
Xbit_r82_c5 bl[5] br[5] wl[82] vdd gnd cell_6t
Xbit_r83_c5 bl[5] br[5] wl[83] vdd gnd cell_6t
Xbit_r84_c5 bl[5] br[5] wl[84] vdd gnd cell_6t
Xbit_r85_c5 bl[5] br[5] wl[85] vdd gnd cell_6t
Xbit_r86_c5 bl[5] br[5] wl[86] vdd gnd cell_6t
Xbit_r87_c5 bl[5] br[5] wl[87] vdd gnd cell_6t
Xbit_r88_c5 bl[5] br[5] wl[88] vdd gnd cell_6t
Xbit_r89_c5 bl[5] br[5] wl[89] vdd gnd cell_6t
Xbit_r90_c5 bl[5] br[5] wl[90] vdd gnd cell_6t
Xbit_r91_c5 bl[5] br[5] wl[91] vdd gnd cell_6t
Xbit_r92_c5 bl[5] br[5] wl[92] vdd gnd cell_6t
Xbit_r93_c5 bl[5] br[5] wl[93] vdd gnd cell_6t
Xbit_r94_c5 bl[5] br[5] wl[94] vdd gnd cell_6t
Xbit_r95_c5 bl[5] br[5] wl[95] vdd gnd cell_6t
Xbit_r96_c5 bl[5] br[5] wl[96] vdd gnd cell_6t
Xbit_r97_c5 bl[5] br[5] wl[97] vdd gnd cell_6t
Xbit_r98_c5 bl[5] br[5] wl[98] vdd gnd cell_6t
Xbit_r99_c5 bl[5] br[5] wl[99] vdd gnd cell_6t
Xbit_r100_c5 bl[5] br[5] wl[100] vdd gnd cell_6t
Xbit_r101_c5 bl[5] br[5] wl[101] vdd gnd cell_6t
Xbit_r102_c5 bl[5] br[5] wl[102] vdd gnd cell_6t
Xbit_r103_c5 bl[5] br[5] wl[103] vdd gnd cell_6t
Xbit_r104_c5 bl[5] br[5] wl[104] vdd gnd cell_6t
Xbit_r105_c5 bl[5] br[5] wl[105] vdd gnd cell_6t
Xbit_r106_c5 bl[5] br[5] wl[106] vdd gnd cell_6t
Xbit_r107_c5 bl[5] br[5] wl[107] vdd gnd cell_6t
Xbit_r108_c5 bl[5] br[5] wl[108] vdd gnd cell_6t
Xbit_r109_c5 bl[5] br[5] wl[109] vdd gnd cell_6t
Xbit_r110_c5 bl[5] br[5] wl[110] vdd gnd cell_6t
Xbit_r111_c5 bl[5] br[5] wl[111] vdd gnd cell_6t
Xbit_r112_c5 bl[5] br[5] wl[112] vdd gnd cell_6t
Xbit_r113_c5 bl[5] br[5] wl[113] vdd gnd cell_6t
Xbit_r114_c5 bl[5] br[5] wl[114] vdd gnd cell_6t
Xbit_r115_c5 bl[5] br[5] wl[115] vdd gnd cell_6t
Xbit_r116_c5 bl[5] br[5] wl[116] vdd gnd cell_6t
Xbit_r117_c5 bl[5] br[5] wl[117] vdd gnd cell_6t
Xbit_r118_c5 bl[5] br[5] wl[118] vdd gnd cell_6t
Xbit_r119_c5 bl[5] br[5] wl[119] vdd gnd cell_6t
Xbit_r120_c5 bl[5] br[5] wl[120] vdd gnd cell_6t
Xbit_r121_c5 bl[5] br[5] wl[121] vdd gnd cell_6t
Xbit_r122_c5 bl[5] br[5] wl[122] vdd gnd cell_6t
Xbit_r123_c5 bl[5] br[5] wl[123] vdd gnd cell_6t
Xbit_r124_c5 bl[5] br[5] wl[124] vdd gnd cell_6t
Xbit_r125_c5 bl[5] br[5] wl[125] vdd gnd cell_6t
Xbit_r126_c5 bl[5] br[5] wl[126] vdd gnd cell_6t
Xbit_r127_c5 bl[5] br[5] wl[127] vdd gnd cell_6t
Xbit_r128_c5 bl[5] br[5] wl[128] vdd gnd cell_6t
Xbit_r129_c5 bl[5] br[5] wl[129] vdd gnd cell_6t
Xbit_r130_c5 bl[5] br[5] wl[130] vdd gnd cell_6t
Xbit_r131_c5 bl[5] br[5] wl[131] vdd gnd cell_6t
Xbit_r132_c5 bl[5] br[5] wl[132] vdd gnd cell_6t
Xbit_r133_c5 bl[5] br[5] wl[133] vdd gnd cell_6t
Xbit_r134_c5 bl[5] br[5] wl[134] vdd gnd cell_6t
Xbit_r135_c5 bl[5] br[5] wl[135] vdd gnd cell_6t
Xbit_r136_c5 bl[5] br[5] wl[136] vdd gnd cell_6t
Xbit_r137_c5 bl[5] br[5] wl[137] vdd gnd cell_6t
Xbit_r138_c5 bl[5] br[5] wl[138] vdd gnd cell_6t
Xbit_r139_c5 bl[5] br[5] wl[139] vdd gnd cell_6t
Xbit_r140_c5 bl[5] br[5] wl[140] vdd gnd cell_6t
Xbit_r141_c5 bl[5] br[5] wl[141] vdd gnd cell_6t
Xbit_r142_c5 bl[5] br[5] wl[142] vdd gnd cell_6t
Xbit_r143_c5 bl[5] br[5] wl[143] vdd gnd cell_6t
Xbit_r144_c5 bl[5] br[5] wl[144] vdd gnd cell_6t
Xbit_r145_c5 bl[5] br[5] wl[145] vdd gnd cell_6t
Xbit_r146_c5 bl[5] br[5] wl[146] vdd gnd cell_6t
Xbit_r147_c5 bl[5] br[5] wl[147] vdd gnd cell_6t
Xbit_r148_c5 bl[5] br[5] wl[148] vdd gnd cell_6t
Xbit_r149_c5 bl[5] br[5] wl[149] vdd gnd cell_6t
Xbit_r150_c5 bl[5] br[5] wl[150] vdd gnd cell_6t
Xbit_r151_c5 bl[5] br[5] wl[151] vdd gnd cell_6t
Xbit_r152_c5 bl[5] br[5] wl[152] vdd gnd cell_6t
Xbit_r153_c5 bl[5] br[5] wl[153] vdd gnd cell_6t
Xbit_r154_c5 bl[5] br[5] wl[154] vdd gnd cell_6t
Xbit_r155_c5 bl[5] br[5] wl[155] vdd gnd cell_6t
Xbit_r156_c5 bl[5] br[5] wl[156] vdd gnd cell_6t
Xbit_r157_c5 bl[5] br[5] wl[157] vdd gnd cell_6t
Xbit_r158_c5 bl[5] br[5] wl[158] vdd gnd cell_6t
Xbit_r159_c5 bl[5] br[5] wl[159] vdd gnd cell_6t
Xbit_r160_c5 bl[5] br[5] wl[160] vdd gnd cell_6t
Xbit_r161_c5 bl[5] br[5] wl[161] vdd gnd cell_6t
Xbit_r162_c5 bl[5] br[5] wl[162] vdd gnd cell_6t
Xbit_r163_c5 bl[5] br[5] wl[163] vdd gnd cell_6t
Xbit_r164_c5 bl[5] br[5] wl[164] vdd gnd cell_6t
Xbit_r165_c5 bl[5] br[5] wl[165] vdd gnd cell_6t
Xbit_r166_c5 bl[5] br[5] wl[166] vdd gnd cell_6t
Xbit_r167_c5 bl[5] br[5] wl[167] vdd gnd cell_6t
Xbit_r168_c5 bl[5] br[5] wl[168] vdd gnd cell_6t
Xbit_r169_c5 bl[5] br[5] wl[169] vdd gnd cell_6t
Xbit_r170_c5 bl[5] br[5] wl[170] vdd gnd cell_6t
Xbit_r171_c5 bl[5] br[5] wl[171] vdd gnd cell_6t
Xbit_r172_c5 bl[5] br[5] wl[172] vdd gnd cell_6t
Xbit_r173_c5 bl[5] br[5] wl[173] vdd gnd cell_6t
Xbit_r174_c5 bl[5] br[5] wl[174] vdd gnd cell_6t
Xbit_r175_c5 bl[5] br[5] wl[175] vdd gnd cell_6t
Xbit_r176_c5 bl[5] br[5] wl[176] vdd gnd cell_6t
Xbit_r177_c5 bl[5] br[5] wl[177] vdd gnd cell_6t
Xbit_r178_c5 bl[5] br[5] wl[178] vdd gnd cell_6t
Xbit_r179_c5 bl[5] br[5] wl[179] vdd gnd cell_6t
Xbit_r180_c5 bl[5] br[5] wl[180] vdd gnd cell_6t
Xbit_r181_c5 bl[5] br[5] wl[181] vdd gnd cell_6t
Xbit_r182_c5 bl[5] br[5] wl[182] vdd gnd cell_6t
Xbit_r183_c5 bl[5] br[5] wl[183] vdd gnd cell_6t
Xbit_r184_c5 bl[5] br[5] wl[184] vdd gnd cell_6t
Xbit_r185_c5 bl[5] br[5] wl[185] vdd gnd cell_6t
Xbit_r186_c5 bl[5] br[5] wl[186] vdd gnd cell_6t
Xbit_r187_c5 bl[5] br[5] wl[187] vdd gnd cell_6t
Xbit_r188_c5 bl[5] br[5] wl[188] vdd gnd cell_6t
Xbit_r189_c5 bl[5] br[5] wl[189] vdd gnd cell_6t
Xbit_r190_c5 bl[5] br[5] wl[190] vdd gnd cell_6t
Xbit_r191_c5 bl[5] br[5] wl[191] vdd gnd cell_6t
Xbit_r192_c5 bl[5] br[5] wl[192] vdd gnd cell_6t
Xbit_r193_c5 bl[5] br[5] wl[193] vdd gnd cell_6t
Xbit_r194_c5 bl[5] br[5] wl[194] vdd gnd cell_6t
Xbit_r195_c5 bl[5] br[5] wl[195] vdd gnd cell_6t
Xbit_r196_c5 bl[5] br[5] wl[196] vdd gnd cell_6t
Xbit_r197_c5 bl[5] br[5] wl[197] vdd gnd cell_6t
Xbit_r198_c5 bl[5] br[5] wl[198] vdd gnd cell_6t
Xbit_r199_c5 bl[5] br[5] wl[199] vdd gnd cell_6t
Xbit_r200_c5 bl[5] br[5] wl[200] vdd gnd cell_6t
Xbit_r201_c5 bl[5] br[5] wl[201] vdd gnd cell_6t
Xbit_r202_c5 bl[5] br[5] wl[202] vdd gnd cell_6t
Xbit_r203_c5 bl[5] br[5] wl[203] vdd gnd cell_6t
Xbit_r204_c5 bl[5] br[5] wl[204] vdd gnd cell_6t
Xbit_r205_c5 bl[5] br[5] wl[205] vdd gnd cell_6t
Xbit_r206_c5 bl[5] br[5] wl[206] vdd gnd cell_6t
Xbit_r207_c5 bl[5] br[5] wl[207] vdd gnd cell_6t
Xbit_r208_c5 bl[5] br[5] wl[208] vdd gnd cell_6t
Xbit_r209_c5 bl[5] br[5] wl[209] vdd gnd cell_6t
Xbit_r210_c5 bl[5] br[5] wl[210] vdd gnd cell_6t
Xbit_r211_c5 bl[5] br[5] wl[211] vdd gnd cell_6t
Xbit_r212_c5 bl[5] br[5] wl[212] vdd gnd cell_6t
Xbit_r213_c5 bl[5] br[5] wl[213] vdd gnd cell_6t
Xbit_r214_c5 bl[5] br[5] wl[214] vdd gnd cell_6t
Xbit_r215_c5 bl[5] br[5] wl[215] vdd gnd cell_6t
Xbit_r216_c5 bl[5] br[5] wl[216] vdd gnd cell_6t
Xbit_r217_c5 bl[5] br[5] wl[217] vdd gnd cell_6t
Xbit_r218_c5 bl[5] br[5] wl[218] vdd gnd cell_6t
Xbit_r219_c5 bl[5] br[5] wl[219] vdd gnd cell_6t
Xbit_r220_c5 bl[5] br[5] wl[220] vdd gnd cell_6t
Xbit_r221_c5 bl[5] br[5] wl[221] vdd gnd cell_6t
Xbit_r222_c5 bl[5] br[5] wl[222] vdd gnd cell_6t
Xbit_r223_c5 bl[5] br[5] wl[223] vdd gnd cell_6t
Xbit_r224_c5 bl[5] br[5] wl[224] vdd gnd cell_6t
Xbit_r225_c5 bl[5] br[5] wl[225] vdd gnd cell_6t
Xbit_r226_c5 bl[5] br[5] wl[226] vdd gnd cell_6t
Xbit_r227_c5 bl[5] br[5] wl[227] vdd gnd cell_6t
Xbit_r228_c5 bl[5] br[5] wl[228] vdd gnd cell_6t
Xbit_r229_c5 bl[5] br[5] wl[229] vdd gnd cell_6t
Xbit_r230_c5 bl[5] br[5] wl[230] vdd gnd cell_6t
Xbit_r231_c5 bl[5] br[5] wl[231] vdd gnd cell_6t
Xbit_r232_c5 bl[5] br[5] wl[232] vdd gnd cell_6t
Xbit_r233_c5 bl[5] br[5] wl[233] vdd gnd cell_6t
Xbit_r234_c5 bl[5] br[5] wl[234] vdd gnd cell_6t
Xbit_r235_c5 bl[5] br[5] wl[235] vdd gnd cell_6t
Xbit_r236_c5 bl[5] br[5] wl[236] vdd gnd cell_6t
Xbit_r237_c5 bl[5] br[5] wl[237] vdd gnd cell_6t
Xbit_r238_c5 bl[5] br[5] wl[238] vdd gnd cell_6t
Xbit_r239_c5 bl[5] br[5] wl[239] vdd gnd cell_6t
Xbit_r240_c5 bl[5] br[5] wl[240] vdd gnd cell_6t
Xbit_r241_c5 bl[5] br[5] wl[241] vdd gnd cell_6t
Xbit_r242_c5 bl[5] br[5] wl[242] vdd gnd cell_6t
Xbit_r243_c5 bl[5] br[5] wl[243] vdd gnd cell_6t
Xbit_r244_c5 bl[5] br[5] wl[244] vdd gnd cell_6t
Xbit_r245_c5 bl[5] br[5] wl[245] vdd gnd cell_6t
Xbit_r246_c5 bl[5] br[5] wl[246] vdd gnd cell_6t
Xbit_r247_c5 bl[5] br[5] wl[247] vdd gnd cell_6t
Xbit_r248_c5 bl[5] br[5] wl[248] vdd gnd cell_6t
Xbit_r249_c5 bl[5] br[5] wl[249] vdd gnd cell_6t
Xbit_r250_c5 bl[5] br[5] wl[250] vdd gnd cell_6t
Xbit_r251_c5 bl[5] br[5] wl[251] vdd gnd cell_6t
Xbit_r252_c5 bl[5] br[5] wl[252] vdd gnd cell_6t
Xbit_r253_c5 bl[5] br[5] wl[253] vdd gnd cell_6t
Xbit_r254_c5 bl[5] br[5] wl[254] vdd gnd cell_6t
Xbit_r255_c5 bl[5] br[5] wl[255] vdd gnd cell_6t
Xbit_r0_c6 bl[6] br[6] wl[0] vdd gnd cell_6t
Xbit_r1_c6 bl[6] br[6] wl[1] vdd gnd cell_6t
Xbit_r2_c6 bl[6] br[6] wl[2] vdd gnd cell_6t
Xbit_r3_c6 bl[6] br[6] wl[3] vdd gnd cell_6t
Xbit_r4_c6 bl[6] br[6] wl[4] vdd gnd cell_6t
Xbit_r5_c6 bl[6] br[6] wl[5] vdd gnd cell_6t
Xbit_r6_c6 bl[6] br[6] wl[6] vdd gnd cell_6t
Xbit_r7_c6 bl[6] br[6] wl[7] vdd gnd cell_6t
Xbit_r8_c6 bl[6] br[6] wl[8] vdd gnd cell_6t
Xbit_r9_c6 bl[6] br[6] wl[9] vdd gnd cell_6t
Xbit_r10_c6 bl[6] br[6] wl[10] vdd gnd cell_6t
Xbit_r11_c6 bl[6] br[6] wl[11] vdd gnd cell_6t
Xbit_r12_c6 bl[6] br[6] wl[12] vdd gnd cell_6t
Xbit_r13_c6 bl[6] br[6] wl[13] vdd gnd cell_6t
Xbit_r14_c6 bl[6] br[6] wl[14] vdd gnd cell_6t
Xbit_r15_c6 bl[6] br[6] wl[15] vdd gnd cell_6t
Xbit_r16_c6 bl[6] br[6] wl[16] vdd gnd cell_6t
Xbit_r17_c6 bl[6] br[6] wl[17] vdd gnd cell_6t
Xbit_r18_c6 bl[6] br[6] wl[18] vdd gnd cell_6t
Xbit_r19_c6 bl[6] br[6] wl[19] vdd gnd cell_6t
Xbit_r20_c6 bl[6] br[6] wl[20] vdd gnd cell_6t
Xbit_r21_c6 bl[6] br[6] wl[21] vdd gnd cell_6t
Xbit_r22_c6 bl[6] br[6] wl[22] vdd gnd cell_6t
Xbit_r23_c6 bl[6] br[6] wl[23] vdd gnd cell_6t
Xbit_r24_c6 bl[6] br[6] wl[24] vdd gnd cell_6t
Xbit_r25_c6 bl[6] br[6] wl[25] vdd gnd cell_6t
Xbit_r26_c6 bl[6] br[6] wl[26] vdd gnd cell_6t
Xbit_r27_c6 bl[6] br[6] wl[27] vdd gnd cell_6t
Xbit_r28_c6 bl[6] br[6] wl[28] vdd gnd cell_6t
Xbit_r29_c6 bl[6] br[6] wl[29] vdd gnd cell_6t
Xbit_r30_c6 bl[6] br[6] wl[30] vdd gnd cell_6t
Xbit_r31_c6 bl[6] br[6] wl[31] vdd gnd cell_6t
Xbit_r32_c6 bl[6] br[6] wl[32] vdd gnd cell_6t
Xbit_r33_c6 bl[6] br[6] wl[33] vdd gnd cell_6t
Xbit_r34_c6 bl[6] br[6] wl[34] vdd gnd cell_6t
Xbit_r35_c6 bl[6] br[6] wl[35] vdd gnd cell_6t
Xbit_r36_c6 bl[6] br[6] wl[36] vdd gnd cell_6t
Xbit_r37_c6 bl[6] br[6] wl[37] vdd gnd cell_6t
Xbit_r38_c6 bl[6] br[6] wl[38] vdd gnd cell_6t
Xbit_r39_c6 bl[6] br[6] wl[39] vdd gnd cell_6t
Xbit_r40_c6 bl[6] br[6] wl[40] vdd gnd cell_6t
Xbit_r41_c6 bl[6] br[6] wl[41] vdd gnd cell_6t
Xbit_r42_c6 bl[6] br[6] wl[42] vdd gnd cell_6t
Xbit_r43_c6 bl[6] br[6] wl[43] vdd gnd cell_6t
Xbit_r44_c6 bl[6] br[6] wl[44] vdd gnd cell_6t
Xbit_r45_c6 bl[6] br[6] wl[45] vdd gnd cell_6t
Xbit_r46_c6 bl[6] br[6] wl[46] vdd gnd cell_6t
Xbit_r47_c6 bl[6] br[6] wl[47] vdd gnd cell_6t
Xbit_r48_c6 bl[6] br[6] wl[48] vdd gnd cell_6t
Xbit_r49_c6 bl[6] br[6] wl[49] vdd gnd cell_6t
Xbit_r50_c6 bl[6] br[6] wl[50] vdd gnd cell_6t
Xbit_r51_c6 bl[6] br[6] wl[51] vdd gnd cell_6t
Xbit_r52_c6 bl[6] br[6] wl[52] vdd gnd cell_6t
Xbit_r53_c6 bl[6] br[6] wl[53] vdd gnd cell_6t
Xbit_r54_c6 bl[6] br[6] wl[54] vdd gnd cell_6t
Xbit_r55_c6 bl[6] br[6] wl[55] vdd gnd cell_6t
Xbit_r56_c6 bl[6] br[6] wl[56] vdd gnd cell_6t
Xbit_r57_c6 bl[6] br[6] wl[57] vdd gnd cell_6t
Xbit_r58_c6 bl[6] br[6] wl[58] vdd gnd cell_6t
Xbit_r59_c6 bl[6] br[6] wl[59] vdd gnd cell_6t
Xbit_r60_c6 bl[6] br[6] wl[60] vdd gnd cell_6t
Xbit_r61_c6 bl[6] br[6] wl[61] vdd gnd cell_6t
Xbit_r62_c6 bl[6] br[6] wl[62] vdd gnd cell_6t
Xbit_r63_c6 bl[6] br[6] wl[63] vdd gnd cell_6t
Xbit_r64_c6 bl[6] br[6] wl[64] vdd gnd cell_6t
Xbit_r65_c6 bl[6] br[6] wl[65] vdd gnd cell_6t
Xbit_r66_c6 bl[6] br[6] wl[66] vdd gnd cell_6t
Xbit_r67_c6 bl[6] br[6] wl[67] vdd gnd cell_6t
Xbit_r68_c6 bl[6] br[6] wl[68] vdd gnd cell_6t
Xbit_r69_c6 bl[6] br[6] wl[69] vdd gnd cell_6t
Xbit_r70_c6 bl[6] br[6] wl[70] vdd gnd cell_6t
Xbit_r71_c6 bl[6] br[6] wl[71] vdd gnd cell_6t
Xbit_r72_c6 bl[6] br[6] wl[72] vdd gnd cell_6t
Xbit_r73_c6 bl[6] br[6] wl[73] vdd gnd cell_6t
Xbit_r74_c6 bl[6] br[6] wl[74] vdd gnd cell_6t
Xbit_r75_c6 bl[6] br[6] wl[75] vdd gnd cell_6t
Xbit_r76_c6 bl[6] br[6] wl[76] vdd gnd cell_6t
Xbit_r77_c6 bl[6] br[6] wl[77] vdd gnd cell_6t
Xbit_r78_c6 bl[6] br[6] wl[78] vdd gnd cell_6t
Xbit_r79_c6 bl[6] br[6] wl[79] vdd gnd cell_6t
Xbit_r80_c6 bl[6] br[6] wl[80] vdd gnd cell_6t
Xbit_r81_c6 bl[6] br[6] wl[81] vdd gnd cell_6t
Xbit_r82_c6 bl[6] br[6] wl[82] vdd gnd cell_6t
Xbit_r83_c6 bl[6] br[6] wl[83] vdd gnd cell_6t
Xbit_r84_c6 bl[6] br[6] wl[84] vdd gnd cell_6t
Xbit_r85_c6 bl[6] br[6] wl[85] vdd gnd cell_6t
Xbit_r86_c6 bl[6] br[6] wl[86] vdd gnd cell_6t
Xbit_r87_c6 bl[6] br[6] wl[87] vdd gnd cell_6t
Xbit_r88_c6 bl[6] br[6] wl[88] vdd gnd cell_6t
Xbit_r89_c6 bl[6] br[6] wl[89] vdd gnd cell_6t
Xbit_r90_c6 bl[6] br[6] wl[90] vdd gnd cell_6t
Xbit_r91_c6 bl[6] br[6] wl[91] vdd gnd cell_6t
Xbit_r92_c6 bl[6] br[6] wl[92] vdd gnd cell_6t
Xbit_r93_c6 bl[6] br[6] wl[93] vdd gnd cell_6t
Xbit_r94_c6 bl[6] br[6] wl[94] vdd gnd cell_6t
Xbit_r95_c6 bl[6] br[6] wl[95] vdd gnd cell_6t
Xbit_r96_c6 bl[6] br[6] wl[96] vdd gnd cell_6t
Xbit_r97_c6 bl[6] br[6] wl[97] vdd gnd cell_6t
Xbit_r98_c6 bl[6] br[6] wl[98] vdd gnd cell_6t
Xbit_r99_c6 bl[6] br[6] wl[99] vdd gnd cell_6t
Xbit_r100_c6 bl[6] br[6] wl[100] vdd gnd cell_6t
Xbit_r101_c6 bl[6] br[6] wl[101] vdd gnd cell_6t
Xbit_r102_c6 bl[6] br[6] wl[102] vdd gnd cell_6t
Xbit_r103_c6 bl[6] br[6] wl[103] vdd gnd cell_6t
Xbit_r104_c6 bl[6] br[6] wl[104] vdd gnd cell_6t
Xbit_r105_c6 bl[6] br[6] wl[105] vdd gnd cell_6t
Xbit_r106_c6 bl[6] br[6] wl[106] vdd gnd cell_6t
Xbit_r107_c6 bl[6] br[6] wl[107] vdd gnd cell_6t
Xbit_r108_c6 bl[6] br[6] wl[108] vdd gnd cell_6t
Xbit_r109_c6 bl[6] br[6] wl[109] vdd gnd cell_6t
Xbit_r110_c6 bl[6] br[6] wl[110] vdd gnd cell_6t
Xbit_r111_c6 bl[6] br[6] wl[111] vdd gnd cell_6t
Xbit_r112_c6 bl[6] br[6] wl[112] vdd gnd cell_6t
Xbit_r113_c6 bl[6] br[6] wl[113] vdd gnd cell_6t
Xbit_r114_c6 bl[6] br[6] wl[114] vdd gnd cell_6t
Xbit_r115_c6 bl[6] br[6] wl[115] vdd gnd cell_6t
Xbit_r116_c6 bl[6] br[6] wl[116] vdd gnd cell_6t
Xbit_r117_c6 bl[6] br[6] wl[117] vdd gnd cell_6t
Xbit_r118_c6 bl[6] br[6] wl[118] vdd gnd cell_6t
Xbit_r119_c6 bl[6] br[6] wl[119] vdd gnd cell_6t
Xbit_r120_c6 bl[6] br[6] wl[120] vdd gnd cell_6t
Xbit_r121_c6 bl[6] br[6] wl[121] vdd gnd cell_6t
Xbit_r122_c6 bl[6] br[6] wl[122] vdd gnd cell_6t
Xbit_r123_c6 bl[6] br[6] wl[123] vdd gnd cell_6t
Xbit_r124_c6 bl[6] br[6] wl[124] vdd gnd cell_6t
Xbit_r125_c6 bl[6] br[6] wl[125] vdd gnd cell_6t
Xbit_r126_c6 bl[6] br[6] wl[126] vdd gnd cell_6t
Xbit_r127_c6 bl[6] br[6] wl[127] vdd gnd cell_6t
Xbit_r128_c6 bl[6] br[6] wl[128] vdd gnd cell_6t
Xbit_r129_c6 bl[6] br[6] wl[129] vdd gnd cell_6t
Xbit_r130_c6 bl[6] br[6] wl[130] vdd gnd cell_6t
Xbit_r131_c6 bl[6] br[6] wl[131] vdd gnd cell_6t
Xbit_r132_c6 bl[6] br[6] wl[132] vdd gnd cell_6t
Xbit_r133_c6 bl[6] br[6] wl[133] vdd gnd cell_6t
Xbit_r134_c6 bl[6] br[6] wl[134] vdd gnd cell_6t
Xbit_r135_c6 bl[6] br[6] wl[135] vdd gnd cell_6t
Xbit_r136_c6 bl[6] br[6] wl[136] vdd gnd cell_6t
Xbit_r137_c6 bl[6] br[6] wl[137] vdd gnd cell_6t
Xbit_r138_c6 bl[6] br[6] wl[138] vdd gnd cell_6t
Xbit_r139_c6 bl[6] br[6] wl[139] vdd gnd cell_6t
Xbit_r140_c6 bl[6] br[6] wl[140] vdd gnd cell_6t
Xbit_r141_c6 bl[6] br[6] wl[141] vdd gnd cell_6t
Xbit_r142_c6 bl[6] br[6] wl[142] vdd gnd cell_6t
Xbit_r143_c6 bl[6] br[6] wl[143] vdd gnd cell_6t
Xbit_r144_c6 bl[6] br[6] wl[144] vdd gnd cell_6t
Xbit_r145_c6 bl[6] br[6] wl[145] vdd gnd cell_6t
Xbit_r146_c6 bl[6] br[6] wl[146] vdd gnd cell_6t
Xbit_r147_c6 bl[6] br[6] wl[147] vdd gnd cell_6t
Xbit_r148_c6 bl[6] br[6] wl[148] vdd gnd cell_6t
Xbit_r149_c6 bl[6] br[6] wl[149] vdd gnd cell_6t
Xbit_r150_c6 bl[6] br[6] wl[150] vdd gnd cell_6t
Xbit_r151_c6 bl[6] br[6] wl[151] vdd gnd cell_6t
Xbit_r152_c6 bl[6] br[6] wl[152] vdd gnd cell_6t
Xbit_r153_c6 bl[6] br[6] wl[153] vdd gnd cell_6t
Xbit_r154_c6 bl[6] br[6] wl[154] vdd gnd cell_6t
Xbit_r155_c6 bl[6] br[6] wl[155] vdd gnd cell_6t
Xbit_r156_c6 bl[6] br[6] wl[156] vdd gnd cell_6t
Xbit_r157_c6 bl[6] br[6] wl[157] vdd gnd cell_6t
Xbit_r158_c6 bl[6] br[6] wl[158] vdd gnd cell_6t
Xbit_r159_c6 bl[6] br[6] wl[159] vdd gnd cell_6t
Xbit_r160_c6 bl[6] br[6] wl[160] vdd gnd cell_6t
Xbit_r161_c6 bl[6] br[6] wl[161] vdd gnd cell_6t
Xbit_r162_c6 bl[6] br[6] wl[162] vdd gnd cell_6t
Xbit_r163_c6 bl[6] br[6] wl[163] vdd gnd cell_6t
Xbit_r164_c6 bl[6] br[6] wl[164] vdd gnd cell_6t
Xbit_r165_c6 bl[6] br[6] wl[165] vdd gnd cell_6t
Xbit_r166_c6 bl[6] br[6] wl[166] vdd gnd cell_6t
Xbit_r167_c6 bl[6] br[6] wl[167] vdd gnd cell_6t
Xbit_r168_c6 bl[6] br[6] wl[168] vdd gnd cell_6t
Xbit_r169_c6 bl[6] br[6] wl[169] vdd gnd cell_6t
Xbit_r170_c6 bl[6] br[6] wl[170] vdd gnd cell_6t
Xbit_r171_c6 bl[6] br[6] wl[171] vdd gnd cell_6t
Xbit_r172_c6 bl[6] br[6] wl[172] vdd gnd cell_6t
Xbit_r173_c6 bl[6] br[6] wl[173] vdd gnd cell_6t
Xbit_r174_c6 bl[6] br[6] wl[174] vdd gnd cell_6t
Xbit_r175_c6 bl[6] br[6] wl[175] vdd gnd cell_6t
Xbit_r176_c6 bl[6] br[6] wl[176] vdd gnd cell_6t
Xbit_r177_c6 bl[6] br[6] wl[177] vdd gnd cell_6t
Xbit_r178_c6 bl[6] br[6] wl[178] vdd gnd cell_6t
Xbit_r179_c6 bl[6] br[6] wl[179] vdd gnd cell_6t
Xbit_r180_c6 bl[6] br[6] wl[180] vdd gnd cell_6t
Xbit_r181_c6 bl[6] br[6] wl[181] vdd gnd cell_6t
Xbit_r182_c6 bl[6] br[6] wl[182] vdd gnd cell_6t
Xbit_r183_c6 bl[6] br[6] wl[183] vdd gnd cell_6t
Xbit_r184_c6 bl[6] br[6] wl[184] vdd gnd cell_6t
Xbit_r185_c6 bl[6] br[6] wl[185] vdd gnd cell_6t
Xbit_r186_c6 bl[6] br[6] wl[186] vdd gnd cell_6t
Xbit_r187_c6 bl[6] br[6] wl[187] vdd gnd cell_6t
Xbit_r188_c6 bl[6] br[6] wl[188] vdd gnd cell_6t
Xbit_r189_c6 bl[6] br[6] wl[189] vdd gnd cell_6t
Xbit_r190_c6 bl[6] br[6] wl[190] vdd gnd cell_6t
Xbit_r191_c6 bl[6] br[6] wl[191] vdd gnd cell_6t
Xbit_r192_c6 bl[6] br[6] wl[192] vdd gnd cell_6t
Xbit_r193_c6 bl[6] br[6] wl[193] vdd gnd cell_6t
Xbit_r194_c6 bl[6] br[6] wl[194] vdd gnd cell_6t
Xbit_r195_c6 bl[6] br[6] wl[195] vdd gnd cell_6t
Xbit_r196_c6 bl[6] br[6] wl[196] vdd gnd cell_6t
Xbit_r197_c6 bl[6] br[6] wl[197] vdd gnd cell_6t
Xbit_r198_c6 bl[6] br[6] wl[198] vdd gnd cell_6t
Xbit_r199_c6 bl[6] br[6] wl[199] vdd gnd cell_6t
Xbit_r200_c6 bl[6] br[6] wl[200] vdd gnd cell_6t
Xbit_r201_c6 bl[6] br[6] wl[201] vdd gnd cell_6t
Xbit_r202_c6 bl[6] br[6] wl[202] vdd gnd cell_6t
Xbit_r203_c6 bl[6] br[6] wl[203] vdd gnd cell_6t
Xbit_r204_c6 bl[6] br[6] wl[204] vdd gnd cell_6t
Xbit_r205_c6 bl[6] br[6] wl[205] vdd gnd cell_6t
Xbit_r206_c6 bl[6] br[6] wl[206] vdd gnd cell_6t
Xbit_r207_c6 bl[6] br[6] wl[207] vdd gnd cell_6t
Xbit_r208_c6 bl[6] br[6] wl[208] vdd gnd cell_6t
Xbit_r209_c6 bl[6] br[6] wl[209] vdd gnd cell_6t
Xbit_r210_c6 bl[6] br[6] wl[210] vdd gnd cell_6t
Xbit_r211_c6 bl[6] br[6] wl[211] vdd gnd cell_6t
Xbit_r212_c6 bl[6] br[6] wl[212] vdd gnd cell_6t
Xbit_r213_c6 bl[6] br[6] wl[213] vdd gnd cell_6t
Xbit_r214_c6 bl[6] br[6] wl[214] vdd gnd cell_6t
Xbit_r215_c6 bl[6] br[6] wl[215] vdd gnd cell_6t
Xbit_r216_c6 bl[6] br[6] wl[216] vdd gnd cell_6t
Xbit_r217_c6 bl[6] br[6] wl[217] vdd gnd cell_6t
Xbit_r218_c6 bl[6] br[6] wl[218] vdd gnd cell_6t
Xbit_r219_c6 bl[6] br[6] wl[219] vdd gnd cell_6t
Xbit_r220_c6 bl[6] br[6] wl[220] vdd gnd cell_6t
Xbit_r221_c6 bl[6] br[6] wl[221] vdd gnd cell_6t
Xbit_r222_c6 bl[6] br[6] wl[222] vdd gnd cell_6t
Xbit_r223_c6 bl[6] br[6] wl[223] vdd gnd cell_6t
Xbit_r224_c6 bl[6] br[6] wl[224] vdd gnd cell_6t
Xbit_r225_c6 bl[6] br[6] wl[225] vdd gnd cell_6t
Xbit_r226_c6 bl[6] br[6] wl[226] vdd gnd cell_6t
Xbit_r227_c6 bl[6] br[6] wl[227] vdd gnd cell_6t
Xbit_r228_c6 bl[6] br[6] wl[228] vdd gnd cell_6t
Xbit_r229_c6 bl[6] br[6] wl[229] vdd gnd cell_6t
Xbit_r230_c6 bl[6] br[6] wl[230] vdd gnd cell_6t
Xbit_r231_c6 bl[6] br[6] wl[231] vdd gnd cell_6t
Xbit_r232_c6 bl[6] br[6] wl[232] vdd gnd cell_6t
Xbit_r233_c6 bl[6] br[6] wl[233] vdd gnd cell_6t
Xbit_r234_c6 bl[6] br[6] wl[234] vdd gnd cell_6t
Xbit_r235_c6 bl[6] br[6] wl[235] vdd gnd cell_6t
Xbit_r236_c6 bl[6] br[6] wl[236] vdd gnd cell_6t
Xbit_r237_c6 bl[6] br[6] wl[237] vdd gnd cell_6t
Xbit_r238_c6 bl[6] br[6] wl[238] vdd gnd cell_6t
Xbit_r239_c6 bl[6] br[6] wl[239] vdd gnd cell_6t
Xbit_r240_c6 bl[6] br[6] wl[240] vdd gnd cell_6t
Xbit_r241_c6 bl[6] br[6] wl[241] vdd gnd cell_6t
Xbit_r242_c6 bl[6] br[6] wl[242] vdd gnd cell_6t
Xbit_r243_c6 bl[6] br[6] wl[243] vdd gnd cell_6t
Xbit_r244_c6 bl[6] br[6] wl[244] vdd gnd cell_6t
Xbit_r245_c6 bl[6] br[6] wl[245] vdd gnd cell_6t
Xbit_r246_c6 bl[6] br[6] wl[246] vdd gnd cell_6t
Xbit_r247_c6 bl[6] br[6] wl[247] vdd gnd cell_6t
Xbit_r248_c6 bl[6] br[6] wl[248] vdd gnd cell_6t
Xbit_r249_c6 bl[6] br[6] wl[249] vdd gnd cell_6t
Xbit_r250_c6 bl[6] br[6] wl[250] vdd gnd cell_6t
Xbit_r251_c6 bl[6] br[6] wl[251] vdd gnd cell_6t
Xbit_r252_c6 bl[6] br[6] wl[252] vdd gnd cell_6t
Xbit_r253_c6 bl[6] br[6] wl[253] vdd gnd cell_6t
Xbit_r254_c6 bl[6] br[6] wl[254] vdd gnd cell_6t
Xbit_r255_c6 bl[6] br[6] wl[255] vdd gnd cell_6t
Xbit_r0_c7 bl[7] br[7] wl[0] vdd gnd cell_6t
Xbit_r1_c7 bl[7] br[7] wl[1] vdd gnd cell_6t
Xbit_r2_c7 bl[7] br[7] wl[2] vdd gnd cell_6t
Xbit_r3_c7 bl[7] br[7] wl[3] vdd gnd cell_6t
Xbit_r4_c7 bl[7] br[7] wl[4] vdd gnd cell_6t
Xbit_r5_c7 bl[7] br[7] wl[5] vdd gnd cell_6t
Xbit_r6_c7 bl[7] br[7] wl[6] vdd gnd cell_6t
Xbit_r7_c7 bl[7] br[7] wl[7] vdd gnd cell_6t
Xbit_r8_c7 bl[7] br[7] wl[8] vdd gnd cell_6t
Xbit_r9_c7 bl[7] br[7] wl[9] vdd gnd cell_6t
Xbit_r10_c7 bl[7] br[7] wl[10] vdd gnd cell_6t
Xbit_r11_c7 bl[7] br[7] wl[11] vdd gnd cell_6t
Xbit_r12_c7 bl[7] br[7] wl[12] vdd gnd cell_6t
Xbit_r13_c7 bl[7] br[7] wl[13] vdd gnd cell_6t
Xbit_r14_c7 bl[7] br[7] wl[14] vdd gnd cell_6t
Xbit_r15_c7 bl[7] br[7] wl[15] vdd gnd cell_6t
Xbit_r16_c7 bl[7] br[7] wl[16] vdd gnd cell_6t
Xbit_r17_c7 bl[7] br[7] wl[17] vdd gnd cell_6t
Xbit_r18_c7 bl[7] br[7] wl[18] vdd gnd cell_6t
Xbit_r19_c7 bl[7] br[7] wl[19] vdd gnd cell_6t
Xbit_r20_c7 bl[7] br[7] wl[20] vdd gnd cell_6t
Xbit_r21_c7 bl[7] br[7] wl[21] vdd gnd cell_6t
Xbit_r22_c7 bl[7] br[7] wl[22] vdd gnd cell_6t
Xbit_r23_c7 bl[7] br[7] wl[23] vdd gnd cell_6t
Xbit_r24_c7 bl[7] br[7] wl[24] vdd gnd cell_6t
Xbit_r25_c7 bl[7] br[7] wl[25] vdd gnd cell_6t
Xbit_r26_c7 bl[7] br[7] wl[26] vdd gnd cell_6t
Xbit_r27_c7 bl[7] br[7] wl[27] vdd gnd cell_6t
Xbit_r28_c7 bl[7] br[7] wl[28] vdd gnd cell_6t
Xbit_r29_c7 bl[7] br[7] wl[29] vdd gnd cell_6t
Xbit_r30_c7 bl[7] br[7] wl[30] vdd gnd cell_6t
Xbit_r31_c7 bl[7] br[7] wl[31] vdd gnd cell_6t
Xbit_r32_c7 bl[7] br[7] wl[32] vdd gnd cell_6t
Xbit_r33_c7 bl[7] br[7] wl[33] vdd gnd cell_6t
Xbit_r34_c7 bl[7] br[7] wl[34] vdd gnd cell_6t
Xbit_r35_c7 bl[7] br[7] wl[35] vdd gnd cell_6t
Xbit_r36_c7 bl[7] br[7] wl[36] vdd gnd cell_6t
Xbit_r37_c7 bl[7] br[7] wl[37] vdd gnd cell_6t
Xbit_r38_c7 bl[7] br[7] wl[38] vdd gnd cell_6t
Xbit_r39_c7 bl[7] br[7] wl[39] vdd gnd cell_6t
Xbit_r40_c7 bl[7] br[7] wl[40] vdd gnd cell_6t
Xbit_r41_c7 bl[7] br[7] wl[41] vdd gnd cell_6t
Xbit_r42_c7 bl[7] br[7] wl[42] vdd gnd cell_6t
Xbit_r43_c7 bl[7] br[7] wl[43] vdd gnd cell_6t
Xbit_r44_c7 bl[7] br[7] wl[44] vdd gnd cell_6t
Xbit_r45_c7 bl[7] br[7] wl[45] vdd gnd cell_6t
Xbit_r46_c7 bl[7] br[7] wl[46] vdd gnd cell_6t
Xbit_r47_c7 bl[7] br[7] wl[47] vdd gnd cell_6t
Xbit_r48_c7 bl[7] br[7] wl[48] vdd gnd cell_6t
Xbit_r49_c7 bl[7] br[7] wl[49] vdd gnd cell_6t
Xbit_r50_c7 bl[7] br[7] wl[50] vdd gnd cell_6t
Xbit_r51_c7 bl[7] br[7] wl[51] vdd gnd cell_6t
Xbit_r52_c7 bl[7] br[7] wl[52] vdd gnd cell_6t
Xbit_r53_c7 bl[7] br[7] wl[53] vdd gnd cell_6t
Xbit_r54_c7 bl[7] br[7] wl[54] vdd gnd cell_6t
Xbit_r55_c7 bl[7] br[7] wl[55] vdd gnd cell_6t
Xbit_r56_c7 bl[7] br[7] wl[56] vdd gnd cell_6t
Xbit_r57_c7 bl[7] br[7] wl[57] vdd gnd cell_6t
Xbit_r58_c7 bl[7] br[7] wl[58] vdd gnd cell_6t
Xbit_r59_c7 bl[7] br[7] wl[59] vdd gnd cell_6t
Xbit_r60_c7 bl[7] br[7] wl[60] vdd gnd cell_6t
Xbit_r61_c7 bl[7] br[7] wl[61] vdd gnd cell_6t
Xbit_r62_c7 bl[7] br[7] wl[62] vdd gnd cell_6t
Xbit_r63_c7 bl[7] br[7] wl[63] vdd gnd cell_6t
Xbit_r64_c7 bl[7] br[7] wl[64] vdd gnd cell_6t
Xbit_r65_c7 bl[7] br[7] wl[65] vdd gnd cell_6t
Xbit_r66_c7 bl[7] br[7] wl[66] vdd gnd cell_6t
Xbit_r67_c7 bl[7] br[7] wl[67] vdd gnd cell_6t
Xbit_r68_c7 bl[7] br[7] wl[68] vdd gnd cell_6t
Xbit_r69_c7 bl[7] br[7] wl[69] vdd gnd cell_6t
Xbit_r70_c7 bl[7] br[7] wl[70] vdd gnd cell_6t
Xbit_r71_c7 bl[7] br[7] wl[71] vdd gnd cell_6t
Xbit_r72_c7 bl[7] br[7] wl[72] vdd gnd cell_6t
Xbit_r73_c7 bl[7] br[7] wl[73] vdd gnd cell_6t
Xbit_r74_c7 bl[7] br[7] wl[74] vdd gnd cell_6t
Xbit_r75_c7 bl[7] br[7] wl[75] vdd gnd cell_6t
Xbit_r76_c7 bl[7] br[7] wl[76] vdd gnd cell_6t
Xbit_r77_c7 bl[7] br[7] wl[77] vdd gnd cell_6t
Xbit_r78_c7 bl[7] br[7] wl[78] vdd gnd cell_6t
Xbit_r79_c7 bl[7] br[7] wl[79] vdd gnd cell_6t
Xbit_r80_c7 bl[7] br[7] wl[80] vdd gnd cell_6t
Xbit_r81_c7 bl[7] br[7] wl[81] vdd gnd cell_6t
Xbit_r82_c7 bl[7] br[7] wl[82] vdd gnd cell_6t
Xbit_r83_c7 bl[7] br[7] wl[83] vdd gnd cell_6t
Xbit_r84_c7 bl[7] br[7] wl[84] vdd gnd cell_6t
Xbit_r85_c7 bl[7] br[7] wl[85] vdd gnd cell_6t
Xbit_r86_c7 bl[7] br[7] wl[86] vdd gnd cell_6t
Xbit_r87_c7 bl[7] br[7] wl[87] vdd gnd cell_6t
Xbit_r88_c7 bl[7] br[7] wl[88] vdd gnd cell_6t
Xbit_r89_c7 bl[7] br[7] wl[89] vdd gnd cell_6t
Xbit_r90_c7 bl[7] br[7] wl[90] vdd gnd cell_6t
Xbit_r91_c7 bl[7] br[7] wl[91] vdd gnd cell_6t
Xbit_r92_c7 bl[7] br[7] wl[92] vdd gnd cell_6t
Xbit_r93_c7 bl[7] br[7] wl[93] vdd gnd cell_6t
Xbit_r94_c7 bl[7] br[7] wl[94] vdd gnd cell_6t
Xbit_r95_c7 bl[7] br[7] wl[95] vdd gnd cell_6t
Xbit_r96_c7 bl[7] br[7] wl[96] vdd gnd cell_6t
Xbit_r97_c7 bl[7] br[7] wl[97] vdd gnd cell_6t
Xbit_r98_c7 bl[7] br[7] wl[98] vdd gnd cell_6t
Xbit_r99_c7 bl[7] br[7] wl[99] vdd gnd cell_6t
Xbit_r100_c7 bl[7] br[7] wl[100] vdd gnd cell_6t
Xbit_r101_c7 bl[7] br[7] wl[101] vdd gnd cell_6t
Xbit_r102_c7 bl[7] br[7] wl[102] vdd gnd cell_6t
Xbit_r103_c7 bl[7] br[7] wl[103] vdd gnd cell_6t
Xbit_r104_c7 bl[7] br[7] wl[104] vdd gnd cell_6t
Xbit_r105_c7 bl[7] br[7] wl[105] vdd gnd cell_6t
Xbit_r106_c7 bl[7] br[7] wl[106] vdd gnd cell_6t
Xbit_r107_c7 bl[7] br[7] wl[107] vdd gnd cell_6t
Xbit_r108_c7 bl[7] br[7] wl[108] vdd gnd cell_6t
Xbit_r109_c7 bl[7] br[7] wl[109] vdd gnd cell_6t
Xbit_r110_c7 bl[7] br[7] wl[110] vdd gnd cell_6t
Xbit_r111_c7 bl[7] br[7] wl[111] vdd gnd cell_6t
Xbit_r112_c7 bl[7] br[7] wl[112] vdd gnd cell_6t
Xbit_r113_c7 bl[7] br[7] wl[113] vdd gnd cell_6t
Xbit_r114_c7 bl[7] br[7] wl[114] vdd gnd cell_6t
Xbit_r115_c7 bl[7] br[7] wl[115] vdd gnd cell_6t
Xbit_r116_c7 bl[7] br[7] wl[116] vdd gnd cell_6t
Xbit_r117_c7 bl[7] br[7] wl[117] vdd gnd cell_6t
Xbit_r118_c7 bl[7] br[7] wl[118] vdd gnd cell_6t
Xbit_r119_c7 bl[7] br[7] wl[119] vdd gnd cell_6t
Xbit_r120_c7 bl[7] br[7] wl[120] vdd gnd cell_6t
Xbit_r121_c7 bl[7] br[7] wl[121] vdd gnd cell_6t
Xbit_r122_c7 bl[7] br[7] wl[122] vdd gnd cell_6t
Xbit_r123_c7 bl[7] br[7] wl[123] vdd gnd cell_6t
Xbit_r124_c7 bl[7] br[7] wl[124] vdd gnd cell_6t
Xbit_r125_c7 bl[7] br[7] wl[125] vdd gnd cell_6t
Xbit_r126_c7 bl[7] br[7] wl[126] vdd gnd cell_6t
Xbit_r127_c7 bl[7] br[7] wl[127] vdd gnd cell_6t
Xbit_r128_c7 bl[7] br[7] wl[128] vdd gnd cell_6t
Xbit_r129_c7 bl[7] br[7] wl[129] vdd gnd cell_6t
Xbit_r130_c7 bl[7] br[7] wl[130] vdd gnd cell_6t
Xbit_r131_c7 bl[7] br[7] wl[131] vdd gnd cell_6t
Xbit_r132_c7 bl[7] br[7] wl[132] vdd gnd cell_6t
Xbit_r133_c7 bl[7] br[7] wl[133] vdd gnd cell_6t
Xbit_r134_c7 bl[7] br[7] wl[134] vdd gnd cell_6t
Xbit_r135_c7 bl[7] br[7] wl[135] vdd gnd cell_6t
Xbit_r136_c7 bl[7] br[7] wl[136] vdd gnd cell_6t
Xbit_r137_c7 bl[7] br[7] wl[137] vdd gnd cell_6t
Xbit_r138_c7 bl[7] br[7] wl[138] vdd gnd cell_6t
Xbit_r139_c7 bl[7] br[7] wl[139] vdd gnd cell_6t
Xbit_r140_c7 bl[7] br[7] wl[140] vdd gnd cell_6t
Xbit_r141_c7 bl[7] br[7] wl[141] vdd gnd cell_6t
Xbit_r142_c7 bl[7] br[7] wl[142] vdd gnd cell_6t
Xbit_r143_c7 bl[7] br[7] wl[143] vdd gnd cell_6t
Xbit_r144_c7 bl[7] br[7] wl[144] vdd gnd cell_6t
Xbit_r145_c7 bl[7] br[7] wl[145] vdd gnd cell_6t
Xbit_r146_c7 bl[7] br[7] wl[146] vdd gnd cell_6t
Xbit_r147_c7 bl[7] br[7] wl[147] vdd gnd cell_6t
Xbit_r148_c7 bl[7] br[7] wl[148] vdd gnd cell_6t
Xbit_r149_c7 bl[7] br[7] wl[149] vdd gnd cell_6t
Xbit_r150_c7 bl[7] br[7] wl[150] vdd gnd cell_6t
Xbit_r151_c7 bl[7] br[7] wl[151] vdd gnd cell_6t
Xbit_r152_c7 bl[7] br[7] wl[152] vdd gnd cell_6t
Xbit_r153_c7 bl[7] br[7] wl[153] vdd gnd cell_6t
Xbit_r154_c7 bl[7] br[7] wl[154] vdd gnd cell_6t
Xbit_r155_c7 bl[7] br[7] wl[155] vdd gnd cell_6t
Xbit_r156_c7 bl[7] br[7] wl[156] vdd gnd cell_6t
Xbit_r157_c7 bl[7] br[7] wl[157] vdd gnd cell_6t
Xbit_r158_c7 bl[7] br[7] wl[158] vdd gnd cell_6t
Xbit_r159_c7 bl[7] br[7] wl[159] vdd gnd cell_6t
Xbit_r160_c7 bl[7] br[7] wl[160] vdd gnd cell_6t
Xbit_r161_c7 bl[7] br[7] wl[161] vdd gnd cell_6t
Xbit_r162_c7 bl[7] br[7] wl[162] vdd gnd cell_6t
Xbit_r163_c7 bl[7] br[7] wl[163] vdd gnd cell_6t
Xbit_r164_c7 bl[7] br[7] wl[164] vdd gnd cell_6t
Xbit_r165_c7 bl[7] br[7] wl[165] vdd gnd cell_6t
Xbit_r166_c7 bl[7] br[7] wl[166] vdd gnd cell_6t
Xbit_r167_c7 bl[7] br[7] wl[167] vdd gnd cell_6t
Xbit_r168_c7 bl[7] br[7] wl[168] vdd gnd cell_6t
Xbit_r169_c7 bl[7] br[7] wl[169] vdd gnd cell_6t
Xbit_r170_c7 bl[7] br[7] wl[170] vdd gnd cell_6t
Xbit_r171_c7 bl[7] br[7] wl[171] vdd gnd cell_6t
Xbit_r172_c7 bl[7] br[7] wl[172] vdd gnd cell_6t
Xbit_r173_c7 bl[7] br[7] wl[173] vdd gnd cell_6t
Xbit_r174_c7 bl[7] br[7] wl[174] vdd gnd cell_6t
Xbit_r175_c7 bl[7] br[7] wl[175] vdd gnd cell_6t
Xbit_r176_c7 bl[7] br[7] wl[176] vdd gnd cell_6t
Xbit_r177_c7 bl[7] br[7] wl[177] vdd gnd cell_6t
Xbit_r178_c7 bl[7] br[7] wl[178] vdd gnd cell_6t
Xbit_r179_c7 bl[7] br[7] wl[179] vdd gnd cell_6t
Xbit_r180_c7 bl[7] br[7] wl[180] vdd gnd cell_6t
Xbit_r181_c7 bl[7] br[7] wl[181] vdd gnd cell_6t
Xbit_r182_c7 bl[7] br[7] wl[182] vdd gnd cell_6t
Xbit_r183_c7 bl[7] br[7] wl[183] vdd gnd cell_6t
Xbit_r184_c7 bl[7] br[7] wl[184] vdd gnd cell_6t
Xbit_r185_c7 bl[7] br[7] wl[185] vdd gnd cell_6t
Xbit_r186_c7 bl[7] br[7] wl[186] vdd gnd cell_6t
Xbit_r187_c7 bl[7] br[7] wl[187] vdd gnd cell_6t
Xbit_r188_c7 bl[7] br[7] wl[188] vdd gnd cell_6t
Xbit_r189_c7 bl[7] br[7] wl[189] vdd gnd cell_6t
Xbit_r190_c7 bl[7] br[7] wl[190] vdd gnd cell_6t
Xbit_r191_c7 bl[7] br[7] wl[191] vdd gnd cell_6t
Xbit_r192_c7 bl[7] br[7] wl[192] vdd gnd cell_6t
Xbit_r193_c7 bl[7] br[7] wl[193] vdd gnd cell_6t
Xbit_r194_c7 bl[7] br[7] wl[194] vdd gnd cell_6t
Xbit_r195_c7 bl[7] br[7] wl[195] vdd gnd cell_6t
Xbit_r196_c7 bl[7] br[7] wl[196] vdd gnd cell_6t
Xbit_r197_c7 bl[7] br[7] wl[197] vdd gnd cell_6t
Xbit_r198_c7 bl[7] br[7] wl[198] vdd gnd cell_6t
Xbit_r199_c7 bl[7] br[7] wl[199] vdd gnd cell_6t
Xbit_r200_c7 bl[7] br[7] wl[200] vdd gnd cell_6t
Xbit_r201_c7 bl[7] br[7] wl[201] vdd gnd cell_6t
Xbit_r202_c7 bl[7] br[7] wl[202] vdd gnd cell_6t
Xbit_r203_c7 bl[7] br[7] wl[203] vdd gnd cell_6t
Xbit_r204_c7 bl[7] br[7] wl[204] vdd gnd cell_6t
Xbit_r205_c7 bl[7] br[7] wl[205] vdd gnd cell_6t
Xbit_r206_c7 bl[7] br[7] wl[206] vdd gnd cell_6t
Xbit_r207_c7 bl[7] br[7] wl[207] vdd gnd cell_6t
Xbit_r208_c7 bl[7] br[7] wl[208] vdd gnd cell_6t
Xbit_r209_c7 bl[7] br[7] wl[209] vdd gnd cell_6t
Xbit_r210_c7 bl[7] br[7] wl[210] vdd gnd cell_6t
Xbit_r211_c7 bl[7] br[7] wl[211] vdd gnd cell_6t
Xbit_r212_c7 bl[7] br[7] wl[212] vdd gnd cell_6t
Xbit_r213_c7 bl[7] br[7] wl[213] vdd gnd cell_6t
Xbit_r214_c7 bl[7] br[7] wl[214] vdd gnd cell_6t
Xbit_r215_c7 bl[7] br[7] wl[215] vdd gnd cell_6t
Xbit_r216_c7 bl[7] br[7] wl[216] vdd gnd cell_6t
Xbit_r217_c7 bl[7] br[7] wl[217] vdd gnd cell_6t
Xbit_r218_c7 bl[7] br[7] wl[218] vdd gnd cell_6t
Xbit_r219_c7 bl[7] br[7] wl[219] vdd gnd cell_6t
Xbit_r220_c7 bl[7] br[7] wl[220] vdd gnd cell_6t
Xbit_r221_c7 bl[7] br[7] wl[221] vdd gnd cell_6t
Xbit_r222_c7 bl[7] br[7] wl[222] vdd gnd cell_6t
Xbit_r223_c7 bl[7] br[7] wl[223] vdd gnd cell_6t
Xbit_r224_c7 bl[7] br[7] wl[224] vdd gnd cell_6t
Xbit_r225_c7 bl[7] br[7] wl[225] vdd gnd cell_6t
Xbit_r226_c7 bl[7] br[7] wl[226] vdd gnd cell_6t
Xbit_r227_c7 bl[7] br[7] wl[227] vdd gnd cell_6t
Xbit_r228_c7 bl[7] br[7] wl[228] vdd gnd cell_6t
Xbit_r229_c7 bl[7] br[7] wl[229] vdd gnd cell_6t
Xbit_r230_c7 bl[7] br[7] wl[230] vdd gnd cell_6t
Xbit_r231_c7 bl[7] br[7] wl[231] vdd gnd cell_6t
Xbit_r232_c7 bl[7] br[7] wl[232] vdd gnd cell_6t
Xbit_r233_c7 bl[7] br[7] wl[233] vdd gnd cell_6t
Xbit_r234_c7 bl[7] br[7] wl[234] vdd gnd cell_6t
Xbit_r235_c7 bl[7] br[7] wl[235] vdd gnd cell_6t
Xbit_r236_c7 bl[7] br[7] wl[236] vdd gnd cell_6t
Xbit_r237_c7 bl[7] br[7] wl[237] vdd gnd cell_6t
Xbit_r238_c7 bl[7] br[7] wl[238] vdd gnd cell_6t
Xbit_r239_c7 bl[7] br[7] wl[239] vdd gnd cell_6t
Xbit_r240_c7 bl[7] br[7] wl[240] vdd gnd cell_6t
Xbit_r241_c7 bl[7] br[7] wl[241] vdd gnd cell_6t
Xbit_r242_c7 bl[7] br[7] wl[242] vdd gnd cell_6t
Xbit_r243_c7 bl[7] br[7] wl[243] vdd gnd cell_6t
Xbit_r244_c7 bl[7] br[7] wl[244] vdd gnd cell_6t
Xbit_r245_c7 bl[7] br[7] wl[245] vdd gnd cell_6t
Xbit_r246_c7 bl[7] br[7] wl[246] vdd gnd cell_6t
Xbit_r247_c7 bl[7] br[7] wl[247] vdd gnd cell_6t
Xbit_r248_c7 bl[7] br[7] wl[248] vdd gnd cell_6t
Xbit_r249_c7 bl[7] br[7] wl[249] vdd gnd cell_6t
Xbit_r250_c7 bl[7] br[7] wl[250] vdd gnd cell_6t
Xbit_r251_c7 bl[7] br[7] wl[251] vdd gnd cell_6t
Xbit_r252_c7 bl[7] br[7] wl[252] vdd gnd cell_6t
Xbit_r253_c7 bl[7] br[7] wl[253] vdd gnd cell_6t
Xbit_r254_c7 bl[7] br[7] wl[254] vdd gnd cell_6t
Xbit_r255_c7 bl[7] br[7] wl[255] vdd gnd cell_6t
Xbit_r0_c8 bl[8] br[8] wl[0] vdd gnd cell_6t
Xbit_r1_c8 bl[8] br[8] wl[1] vdd gnd cell_6t
Xbit_r2_c8 bl[8] br[8] wl[2] vdd gnd cell_6t
Xbit_r3_c8 bl[8] br[8] wl[3] vdd gnd cell_6t
Xbit_r4_c8 bl[8] br[8] wl[4] vdd gnd cell_6t
Xbit_r5_c8 bl[8] br[8] wl[5] vdd gnd cell_6t
Xbit_r6_c8 bl[8] br[8] wl[6] vdd gnd cell_6t
Xbit_r7_c8 bl[8] br[8] wl[7] vdd gnd cell_6t
Xbit_r8_c8 bl[8] br[8] wl[8] vdd gnd cell_6t
Xbit_r9_c8 bl[8] br[8] wl[9] vdd gnd cell_6t
Xbit_r10_c8 bl[8] br[8] wl[10] vdd gnd cell_6t
Xbit_r11_c8 bl[8] br[8] wl[11] vdd gnd cell_6t
Xbit_r12_c8 bl[8] br[8] wl[12] vdd gnd cell_6t
Xbit_r13_c8 bl[8] br[8] wl[13] vdd gnd cell_6t
Xbit_r14_c8 bl[8] br[8] wl[14] vdd gnd cell_6t
Xbit_r15_c8 bl[8] br[8] wl[15] vdd gnd cell_6t
Xbit_r16_c8 bl[8] br[8] wl[16] vdd gnd cell_6t
Xbit_r17_c8 bl[8] br[8] wl[17] vdd gnd cell_6t
Xbit_r18_c8 bl[8] br[8] wl[18] vdd gnd cell_6t
Xbit_r19_c8 bl[8] br[8] wl[19] vdd gnd cell_6t
Xbit_r20_c8 bl[8] br[8] wl[20] vdd gnd cell_6t
Xbit_r21_c8 bl[8] br[8] wl[21] vdd gnd cell_6t
Xbit_r22_c8 bl[8] br[8] wl[22] vdd gnd cell_6t
Xbit_r23_c8 bl[8] br[8] wl[23] vdd gnd cell_6t
Xbit_r24_c8 bl[8] br[8] wl[24] vdd gnd cell_6t
Xbit_r25_c8 bl[8] br[8] wl[25] vdd gnd cell_6t
Xbit_r26_c8 bl[8] br[8] wl[26] vdd gnd cell_6t
Xbit_r27_c8 bl[8] br[8] wl[27] vdd gnd cell_6t
Xbit_r28_c8 bl[8] br[8] wl[28] vdd gnd cell_6t
Xbit_r29_c8 bl[8] br[8] wl[29] vdd gnd cell_6t
Xbit_r30_c8 bl[8] br[8] wl[30] vdd gnd cell_6t
Xbit_r31_c8 bl[8] br[8] wl[31] vdd gnd cell_6t
Xbit_r32_c8 bl[8] br[8] wl[32] vdd gnd cell_6t
Xbit_r33_c8 bl[8] br[8] wl[33] vdd gnd cell_6t
Xbit_r34_c8 bl[8] br[8] wl[34] vdd gnd cell_6t
Xbit_r35_c8 bl[8] br[8] wl[35] vdd gnd cell_6t
Xbit_r36_c8 bl[8] br[8] wl[36] vdd gnd cell_6t
Xbit_r37_c8 bl[8] br[8] wl[37] vdd gnd cell_6t
Xbit_r38_c8 bl[8] br[8] wl[38] vdd gnd cell_6t
Xbit_r39_c8 bl[8] br[8] wl[39] vdd gnd cell_6t
Xbit_r40_c8 bl[8] br[8] wl[40] vdd gnd cell_6t
Xbit_r41_c8 bl[8] br[8] wl[41] vdd gnd cell_6t
Xbit_r42_c8 bl[8] br[8] wl[42] vdd gnd cell_6t
Xbit_r43_c8 bl[8] br[8] wl[43] vdd gnd cell_6t
Xbit_r44_c8 bl[8] br[8] wl[44] vdd gnd cell_6t
Xbit_r45_c8 bl[8] br[8] wl[45] vdd gnd cell_6t
Xbit_r46_c8 bl[8] br[8] wl[46] vdd gnd cell_6t
Xbit_r47_c8 bl[8] br[8] wl[47] vdd gnd cell_6t
Xbit_r48_c8 bl[8] br[8] wl[48] vdd gnd cell_6t
Xbit_r49_c8 bl[8] br[8] wl[49] vdd gnd cell_6t
Xbit_r50_c8 bl[8] br[8] wl[50] vdd gnd cell_6t
Xbit_r51_c8 bl[8] br[8] wl[51] vdd gnd cell_6t
Xbit_r52_c8 bl[8] br[8] wl[52] vdd gnd cell_6t
Xbit_r53_c8 bl[8] br[8] wl[53] vdd gnd cell_6t
Xbit_r54_c8 bl[8] br[8] wl[54] vdd gnd cell_6t
Xbit_r55_c8 bl[8] br[8] wl[55] vdd gnd cell_6t
Xbit_r56_c8 bl[8] br[8] wl[56] vdd gnd cell_6t
Xbit_r57_c8 bl[8] br[8] wl[57] vdd gnd cell_6t
Xbit_r58_c8 bl[8] br[8] wl[58] vdd gnd cell_6t
Xbit_r59_c8 bl[8] br[8] wl[59] vdd gnd cell_6t
Xbit_r60_c8 bl[8] br[8] wl[60] vdd gnd cell_6t
Xbit_r61_c8 bl[8] br[8] wl[61] vdd gnd cell_6t
Xbit_r62_c8 bl[8] br[8] wl[62] vdd gnd cell_6t
Xbit_r63_c8 bl[8] br[8] wl[63] vdd gnd cell_6t
Xbit_r64_c8 bl[8] br[8] wl[64] vdd gnd cell_6t
Xbit_r65_c8 bl[8] br[8] wl[65] vdd gnd cell_6t
Xbit_r66_c8 bl[8] br[8] wl[66] vdd gnd cell_6t
Xbit_r67_c8 bl[8] br[8] wl[67] vdd gnd cell_6t
Xbit_r68_c8 bl[8] br[8] wl[68] vdd gnd cell_6t
Xbit_r69_c8 bl[8] br[8] wl[69] vdd gnd cell_6t
Xbit_r70_c8 bl[8] br[8] wl[70] vdd gnd cell_6t
Xbit_r71_c8 bl[8] br[8] wl[71] vdd gnd cell_6t
Xbit_r72_c8 bl[8] br[8] wl[72] vdd gnd cell_6t
Xbit_r73_c8 bl[8] br[8] wl[73] vdd gnd cell_6t
Xbit_r74_c8 bl[8] br[8] wl[74] vdd gnd cell_6t
Xbit_r75_c8 bl[8] br[8] wl[75] vdd gnd cell_6t
Xbit_r76_c8 bl[8] br[8] wl[76] vdd gnd cell_6t
Xbit_r77_c8 bl[8] br[8] wl[77] vdd gnd cell_6t
Xbit_r78_c8 bl[8] br[8] wl[78] vdd gnd cell_6t
Xbit_r79_c8 bl[8] br[8] wl[79] vdd gnd cell_6t
Xbit_r80_c8 bl[8] br[8] wl[80] vdd gnd cell_6t
Xbit_r81_c8 bl[8] br[8] wl[81] vdd gnd cell_6t
Xbit_r82_c8 bl[8] br[8] wl[82] vdd gnd cell_6t
Xbit_r83_c8 bl[8] br[8] wl[83] vdd gnd cell_6t
Xbit_r84_c8 bl[8] br[8] wl[84] vdd gnd cell_6t
Xbit_r85_c8 bl[8] br[8] wl[85] vdd gnd cell_6t
Xbit_r86_c8 bl[8] br[8] wl[86] vdd gnd cell_6t
Xbit_r87_c8 bl[8] br[8] wl[87] vdd gnd cell_6t
Xbit_r88_c8 bl[8] br[8] wl[88] vdd gnd cell_6t
Xbit_r89_c8 bl[8] br[8] wl[89] vdd gnd cell_6t
Xbit_r90_c8 bl[8] br[8] wl[90] vdd gnd cell_6t
Xbit_r91_c8 bl[8] br[8] wl[91] vdd gnd cell_6t
Xbit_r92_c8 bl[8] br[8] wl[92] vdd gnd cell_6t
Xbit_r93_c8 bl[8] br[8] wl[93] vdd gnd cell_6t
Xbit_r94_c8 bl[8] br[8] wl[94] vdd gnd cell_6t
Xbit_r95_c8 bl[8] br[8] wl[95] vdd gnd cell_6t
Xbit_r96_c8 bl[8] br[8] wl[96] vdd gnd cell_6t
Xbit_r97_c8 bl[8] br[8] wl[97] vdd gnd cell_6t
Xbit_r98_c8 bl[8] br[8] wl[98] vdd gnd cell_6t
Xbit_r99_c8 bl[8] br[8] wl[99] vdd gnd cell_6t
Xbit_r100_c8 bl[8] br[8] wl[100] vdd gnd cell_6t
Xbit_r101_c8 bl[8] br[8] wl[101] vdd gnd cell_6t
Xbit_r102_c8 bl[8] br[8] wl[102] vdd gnd cell_6t
Xbit_r103_c8 bl[8] br[8] wl[103] vdd gnd cell_6t
Xbit_r104_c8 bl[8] br[8] wl[104] vdd gnd cell_6t
Xbit_r105_c8 bl[8] br[8] wl[105] vdd gnd cell_6t
Xbit_r106_c8 bl[8] br[8] wl[106] vdd gnd cell_6t
Xbit_r107_c8 bl[8] br[8] wl[107] vdd gnd cell_6t
Xbit_r108_c8 bl[8] br[8] wl[108] vdd gnd cell_6t
Xbit_r109_c8 bl[8] br[8] wl[109] vdd gnd cell_6t
Xbit_r110_c8 bl[8] br[8] wl[110] vdd gnd cell_6t
Xbit_r111_c8 bl[8] br[8] wl[111] vdd gnd cell_6t
Xbit_r112_c8 bl[8] br[8] wl[112] vdd gnd cell_6t
Xbit_r113_c8 bl[8] br[8] wl[113] vdd gnd cell_6t
Xbit_r114_c8 bl[8] br[8] wl[114] vdd gnd cell_6t
Xbit_r115_c8 bl[8] br[8] wl[115] vdd gnd cell_6t
Xbit_r116_c8 bl[8] br[8] wl[116] vdd gnd cell_6t
Xbit_r117_c8 bl[8] br[8] wl[117] vdd gnd cell_6t
Xbit_r118_c8 bl[8] br[8] wl[118] vdd gnd cell_6t
Xbit_r119_c8 bl[8] br[8] wl[119] vdd gnd cell_6t
Xbit_r120_c8 bl[8] br[8] wl[120] vdd gnd cell_6t
Xbit_r121_c8 bl[8] br[8] wl[121] vdd gnd cell_6t
Xbit_r122_c8 bl[8] br[8] wl[122] vdd gnd cell_6t
Xbit_r123_c8 bl[8] br[8] wl[123] vdd gnd cell_6t
Xbit_r124_c8 bl[8] br[8] wl[124] vdd gnd cell_6t
Xbit_r125_c8 bl[8] br[8] wl[125] vdd gnd cell_6t
Xbit_r126_c8 bl[8] br[8] wl[126] vdd gnd cell_6t
Xbit_r127_c8 bl[8] br[8] wl[127] vdd gnd cell_6t
Xbit_r128_c8 bl[8] br[8] wl[128] vdd gnd cell_6t
Xbit_r129_c8 bl[8] br[8] wl[129] vdd gnd cell_6t
Xbit_r130_c8 bl[8] br[8] wl[130] vdd gnd cell_6t
Xbit_r131_c8 bl[8] br[8] wl[131] vdd gnd cell_6t
Xbit_r132_c8 bl[8] br[8] wl[132] vdd gnd cell_6t
Xbit_r133_c8 bl[8] br[8] wl[133] vdd gnd cell_6t
Xbit_r134_c8 bl[8] br[8] wl[134] vdd gnd cell_6t
Xbit_r135_c8 bl[8] br[8] wl[135] vdd gnd cell_6t
Xbit_r136_c8 bl[8] br[8] wl[136] vdd gnd cell_6t
Xbit_r137_c8 bl[8] br[8] wl[137] vdd gnd cell_6t
Xbit_r138_c8 bl[8] br[8] wl[138] vdd gnd cell_6t
Xbit_r139_c8 bl[8] br[8] wl[139] vdd gnd cell_6t
Xbit_r140_c8 bl[8] br[8] wl[140] vdd gnd cell_6t
Xbit_r141_c8 bl[8] br[8] wl[141] vdd gnd cell_6t
Xbit_r142_c8 bl[8] br[8] wl[142] vdd gnd cell_6t
Xbit_r143_c8 bl[8] br[8] wl[143] vdd gnd cell_6t
Xbit_r144_c8 bl[8] br[8] wl[144] vdd gnd cell_6t
Xbit_r145_c8 bl[8] br[8] wl[145] vdd gnd cell_6t
Xbit_r146_c8 bl[8] br[8] wl[146] vdd gnd cell_6t
Xbit_r147_c8 bl[8] br[8] wl[147] vdd gnd cell_6t
Xbit_r148_c8 bl[8] br[8] wl[148] vdd gnd cell_6t
Xbit_r149_c8 bl[8] br[8] wl[149] vdd gnd cell_6t
Xbit_r150_c8 bl[8] br[8] wl[150] vdd gnd cell_6t
Xbit_r151_c8 bl[8] br[8] wl[151] vdd gnd cell_6t
Xbit_r152_c8 bl[8] br[8] wl[152] vdd gnd cell_6t
Xbit_r153_c8 bl[8] br[8] wl[153] vdd gnd cell_6t
Xbit_r154_c8 bl[8] br[8] wl[154] vdd gnd cell_6t
Xbit_r155_c8 bl[8] br[8] wl[155] vdd gnd cell_6t
Xbit_r156_c8 bl[8] br[8] wl[156] vdd gnd cell_6t
Xbit_r157_c8 bl[8] br[8] wl[157] vdd gnd cell_6t
Xbit_r158_c8 bl[8] br[8] wl[158] vdd gnd cell_6t
Xbit_r159_c8 bl[8] br[8] wl[159] vdd gnd cell_6t
Xbit_r160_c8 bl[8] br[8] wl[160] vdd gnd cell_6t
Xbit_r161_c8 bl[8] br[8] wl[161] vdd gnd cell_6t
Xbit_r162_c8 bl[8] br[8] wl[162] vdd gnd cell_6t
Xbit_r163_c8 bl[8] br[8] wl[163] vdd gnd cell_6t
Xbit_r164_c8 bl[8] br[8] wl[164] vdd gnd cell_6t
Xbit_r165_c8 bl[8] br[8] wl[165] vdd gnd cell_6t
Xbit_r166_c8 bl[8] br[8] wl[166] vdd gnd cell_6t
Xbit_r167_c8 bl[8] br[8] wl[167] vdd gnd cell_6t
Xbit_r168_c8 bl[8] br[8] wl[168] vdd gnd cell_6t
Xbit_r169_c8 bl[8] br[8] wl[169] vdd gnd cell_6t
Xbit_r170_c8 bl[8] br[8] wl[170] vdd gnd cell_6t
Xbit_r171_c8 bl[8] br[8] wl[171] vdd gnd cell_6t
Xbit_r172_c8 bl[8] br[8] wl[172] vdd gnd cell_6t
Xbit_r173_c8 bl[8] br[8] wl[173] vdd gnd cell_6t
Xbit_r174_c8 bl[8] br[8] wl[174] vdd gnd cell_6t
Xbit_r175_c8 bl[8] br[8] wl[175] vdd gnd cell_6t
Xbit_r176_c8 bl[8] br[8] wl[176] vdd gnd cell_6t
Xbit_r177_c8 bl[8] br[8] wl[177] vdd gnd cell_6t
Xbit_r178_c8 bl[8] br[8] wl[178] vdd gnd cell_6t
Xbit_r179_c8 bl[8] br[8] wl[179] vdd gnd cell_6t
Xbit_r180_c8 bl[8] br[8] wl[180] vdd gnd cell_6t
Xbit_r181_c8 bl[8] br[8] wl[181] vdd gnd cell_6t
Xbit_r182_c8 bl[8] br[8] wl[182] vdd gnd cell_6t
Xbit_r183_c8 bl[8] br[8] wl[183] vdd gnd cell_6t
Xbit_r184_c8 bl[8] br[8] wl[184] vdd gnd cell_6t
Xbit_r185_c8 bl[8] br[8] wl[185] vdd gnd cell_6t
Xbit_r186_c8 bl[8] br[8] wl[186] vdd gnd cell_6t
Xbit_r187_c8 bl[8] br[8] wl[187] vdd gnd cell_6t
Xbit_r188_c8 bl[8] br[8] wl[188] vdd gnd cell_6t
Xbit_r189_c8 bl[8] br[8] wl[189] vdd gnd cell_6t
Xbit_r190_c8 bl[8] br[8] wl[190] vdd gnd cell_6t
Xbit_r191_c8 bl[8] br[8] wl[191] vdd gnd cell_6t
Xbit_r192_c8 bl[8] br[8] wl[192] vdd gnd cell_6t
Xbit_r193_c8 bl[8] br[8] wl[193] vdd gnd cell_6t
Xbit_r194_c8 bl[8] br[8] wl[194] vdd gnd cell_6t
Xbit_r195_c8 bl[8] br[8] wl[195] vdd gnd cell_6t
Xbit_r196_c8 bl[8] br[8] wl[196] vdd gnd cell_6t
Xbit_r197_c8 bl[8] br[8] wl[197] vdd gnd cell_6t
Xbit_r198_c8 bl[8] br[8] wl[198] vdd gnd cell_6t
Xbit_r199_c8 bl[8] br[8] wl[199] vdd gnd cell_6t
Xbit_r200_c8 bl[8] br[8] wl[200] vdd gnd cell_6t
Xbit_r201_c8 bl[8] br[8] wl[201] vdd gnd cell_6t
Xbit_r202_c8 bl[8] br[8] wl[202] vdd gnd cell_6t
Xbit_r203_c8 bl[8] br[8] wl[203] vdd gnd cell_6t
Xbit_r204_c8 bl[8] br[8] wl[204] vdd gnd cell_6t
Xbit_r205_c8 bl[8] br[8] wl[205] vdd gnd cell_6t
Xbit_r206_c8 bl[8] br[8] wl[206] vdd gnd cell_6t
Xbit_r207_c8 bl[8] br[8] wl[207] vdd gnd cell_6t
Xbit_r208_c8 bl[8] br[8] wl[208] vdd gnd cell_6t
Xbit_r209_c8 bl[8] br[8] wl[209] vdd gnd cell_6t
Xbit_r210_c8 bl[8] br[8] wl[210] vdd gnd cell_6t
Xbit_r211_c8 bl[8] br[8] wl[211] vdd gnd cell_6t
Xbit_r212_c8 bl[8] br[8] wl[212] vdd gnd cell_6t
Xbit_r213_c8 bl[8] br[8] wl[213] vdd gnd cell_6t
Xbit_r214_c8 bl[8] br[8] wl[214] vdd gnd cell_6t
Xbit_r215_c8 bl[8] br[8] wl[215] vdd gnd cell_6t
Xbit_r216_c8 bl[8] br[8] wl[216] vdd gnd cell_6t
Xbit_r217_c8 bl[8] br[8] wl[217] vdd gnd cell_6t
Xbit_r218_c8 bl[8] br[8] wl[218] vdd gnd cell_6t
Xbit_r219_c8 bl[8] br[8] wl[219] vdd gnd cell_6t
Xbit_r220_c8 bl[8] br[8] wl[220] vdd gnd cell_6t
Xbit_r221_c8 bl[8] br[8] wl[221] vdd gnd cell_6t
Xbit_r222_c8 bl[8] br[8] wl[222] vdd gnd cell_6t
Xbit_r223_c8 bl[8] br[8] wl[223] vdd gnd cell_6t
Xbit_r224_c8 bl[8] br[8] wl[224] vdd gnd cell_6t
Xbit_r225_c8 bl[8] br[8] wl[225] vdd gnd cell_6t
Xbit_r226_c8 bl[8] br[8] wl[226] vdd gnd cell_6t
Xbit_r227_c8 bl[8] br[8] wl[227] vdd gnd cell_6t
Xbit_r228_c8 bl[8] br[8] wl[228] vdd gnd cell_6t
Xbit_r229_c8 bl[8] br[8] wl[229] vdd gnd cell_6t
Xbit_r230_c8 bl[8] br[8] wl[230] vdd gnd cell_6t
Xbit_r231_c8 bl[8] br[8] wl[231] vdd gnd cell_6t
Xbit_r232_c8 bl[8] br[8] wl[232] vdd gnd cell_6t
Xbit_r233_c8 bl[8] br[8] wl[233] vdd gnd cell_6t
Xbit_r234_c8 bl[8] br[8] wl[234] vdd gnd cell_6t
Xbit_r235_c8 bl[8] br[8] wl[235] vdd gnd cell_6t
Xbit_r236_c8 bl[8] br[8] wl[236] vdd gnd cell_6t
Xbit_r237_c8 bl[8] br[8] wl[237] vdd gnd cell_6t
Xbit_r238_c8 bl[8] br[8] wl[238] vdd gnd cell_6t
Xbit_r239_c8 bl[8] br[8] wl[239] vdd gnd cell_6t
Xbit_r240_c8 bl[8] br[8] wl[240] vdd gnd cell_6t
Xbit_r241_c8 bl[8] br[8] wl[241] vdd gnd cell_6t
Xbit_r242_c8 bl[8] br[8] wl[242] vdd gnd cell_6t
Xbit_r243_c8 bl[8] br[8] wl[243] vdd gnd cell_6t
Xbit_r244_c8 bl[8] br[8] wl[244] vdd gnd cell_6t
Xbit_r245_c8 bl[8] br[8] wl[245] vdd gnd cell_6t
Xbit_r246_c8 bl[8] br[8] wl[246] vdd gnd cell_6t
Xbit_r247_c8 bl[8] br[8] wl[247] vdd gnd cell_6t
Xbit_r248_c8 bl[8] br[8] wl[248] vdd gnd cell_6t
Xbit_r249_c8 bl[8] br[8] wl[249] vdd gnd cell_6t
Xbit_r250_c8 bl[8] br[8] wl[250] vdd gnd cell_6t
Xbit_r251_c8 bl[8] br[8] wl[251] vdd gnd cell_6t
Xbit_r252_c8 bl[8] br[8] wl[252] vdd gnd cell_6t
Xbit_r253_c8 bl[8] br[8] wl[253] vdd gnd cell_6t
Xbit_r254_c8 bl[8] br[8] wl[254] vdd gnd cell_6t
Xbit_r255_c8 bl[8] br[8] wl[255] vdd gnd cell_6t
Xbit_r0_c9 bl[9] br[9] wl[0] vdd gnd cell_6t
Xbit_r1_c9 bl[9] br[9] wl[1] vdd gnd cell_6t
Xbit_r2_c9 bl[9] br[9] wl[2] vdd gnd cell_6t
Xbit_r3_c9 bl[9] br[9] wl[3] vdd gnd cell_6t
Xbit_r4_c9 bl[9] br[9] wl[4] vdd gnd cell_6t
Xbit_r5_c9 bl[9] br[9] wl[5] vdd gnd cell_6t
Xbit_r6_c9 bl[9] br[9] wl[6] vdd gnd cell_6t
Xbit_r7_c9 bl[9] br[9] wl[7] vdd gnd cell_6t
Xbit_r8_c9 bl[9] br[9] wl[8] vdd gnd cell_6t
Xbit_r9_c9 bl[9] br[9] wl[9] vdd gnd cell_6t
Xbit_r10_c9 bl[9] br[9] wl[10] vdd gnd cell_6t
Xbit_r11_c9 bl[9] br[9] wl[11] vdd gnd cell_6t
Xbit_r12_c9 bl[9] br[9] wl[12] vdd gnd cell_6t
Xbit_r13_c9 bl[9] br[9] wl[13] vdd gnd cell_6t
Xbit_r14_c9 bl[9] br[9] wl[14] vdd gnd cell_6t
Xbit_r15_c9 bl[9] br[9] wl[15] vdd gnd cell_6t
Xbit_r16_c9 bl[9] br[9] wl[16] vdd gnd cell_6t
Xbit_r17_c9 bl[9] br[9] wl[17] vdd gnd cell_6t
Xbit_r18_c9 bl[9] br[9] wl[18] vdd gnd cell_6t
Xbit_r19_c9 bl[9] br[9] wl[19] vdd gnd cell_6t
Xbit_r20_c9 bl[9] br[9] wl[20] vdd gnd cell_6t
Xbit_r21_c9 bl[9] br[9] wl[21] vdd gnd cell_6t
Xbit_r22_c9 bl[9] br[9] wl[22] vdd gnd cell_6t
Xbit_r23_c9 bl[9] br[9] wl[23] vdd gnd cell_6t
Xbit_r24_c9 bl[9] br[9] wl[24] vdd gnd cell_6t
Xbit_r25_c9 bl[9] br[9] wl[25] vdd gnd cell_6t
Xbit_r26_c9 bl[9] br[9] wl[26] vdd gnd cell_6t
Xbit_r27_c9 bl[9] br[9] wl[27] vdd gnd cell_6t
Xbit_r28_c9 bl[9] br[9] wl[28] vdd gnd cell_6t
Xbit_r29_c9 bl[9] br[9] wl[29] vdd gnd cell_6t
Xbit_r30_c9 bl[9] br[9] wl[30] vdd gnd cell_6t
Xbit_r31_c9 bl[9] br[9] wl[31] vdd gnd cell_6t
Xbit_r32_c9 bl[9] br[9] wl[32] vdd gnd cell_6t
Xbit_r33_c9 bl[9] br[9] wl[33] vdd gnd cell_6t
Xbit_r34_c9 bl[9] br[9] wl[34] vdd gnd cell_6t
Xbit_r35_c9 bl[9] br[9] wl[35] vdd gnd cell_6t
Xbit_r36_c9 bl[9] br[9] wl[36] vdd gnd cell_6t
Xbit_r37_c9 bl[9] br[9] wl[37] vdd gnd cell_6t
Xbit_r38_c9 bl[9] br[9] wl[38] vdd gnd cell_6t
Xbit_r39_c9 bl[9] br[9] wl[39] vdd gnd cell_6t
Xbit_r40_c9 bl[9] br[9] wl[40] vdd gnd cell_6t
Xbit_r41_c9 bl[9] br[9] wl[41] vdd gnd cell_6t
Xbit_r42_c9 bl[9] br[9] wl[42] vdd gnd cell_6t
Xbit_r43_c9 bl[9] br[9] wl[43] vdd gnd cell_6t
Xbit_r44_c9 bl[9] br[9] wl[44] vdd gnd cell_6t
Xbit_r45_c9 bl[9] br[9] wl[45] vdd gnd cell_6t
Xbit_r46_c9 bl[9] br[9] wl[46] vdd gnd cell_6t
Xbit_r47_c9 bl[9] br[9] wl[47] vdd gnd cell_6t
Xbit_r48_c9 bl[9] br[9] wl[48] vdd gnd cell_6t
Xbit_r49_c9 bl[9] br[9] wl[49] vdd gnd cell_6t
Xbit_r50_c9 bl[9] br[9] wl[50] vdd gnd cell_6t
Xbit_r51_c9 bl[9] br[9] wl[51] vdd gnd cell_6t
Xbit_r52_c9 bl[9] br[9] wl[52] vdd gnd cell_6t
Xbit_r53_c9 bl[9] br[9] wl[53] vdd gnd cell_6t
Xbit_r54_c9 bl[9] br[9] wl[54] vdd gnd cell_6t
Xbit_r55_c9 bl[9] br[9] wl[55] vdd gnd cell_6t
Xbit_r56_c9 bl[9] br[9] wl[56] vdd gnd cell_6t
Xbit_r57_c9 bl[9] br[9] wl[57] vdd gnd cell_6t
Xbit_r58_c9 bl[9] br[9] wl[58] vdd gnd cell_6t
Xbit_r59_c9 bl[9] br[9] wl[59] vdd gnd cell_6t
Xbit_r60_c9 bl[9] br[9] wl[60] vdd gnd cell_6t
Xbit_r61_c9 bl[9] br[9] wl[61] vdd gnd cell_6t
Xbit_r62_c9 bl[9] br[9] wl[62] vdd gnd cell_6t
Xbit_r63_c9 bl[9] br[9] wl[63] vdd gnd cell_6t
Xbit_r64_c9 bl[9] br[9] wl[64] vdd gnd cell_6t
Xbit_r65_c9 bl[9] br[9] wl[65] vdd gnd cell_6t
Xbit_r66_c9 bl[9] br[9] wl[66] vdd gnd cell_6t
Xbit_r67_c9 bl[9] br[9] wl[67] vdd gnd cell_6t
Xbit_r68_c9 bl[9] br[9] wl[68] vdd gnd cell_6t
Xbit_r69_c9 bl[9] br[9] wl[69] vdd gnd cell_6t
Xbit_r70_c9 bl[9] br[9] wl[70] vdd gnd cell_6t
Xbit_r71_c9 bl[9] br[9] wl[71] vdd gnd cell_6t
Xbit_r72_c9 bl[9] br[9] wl[72] vdd gnd cell_6t
Xbit_r73_c9 bl[9] br[9] wl[73] vdd gnd cell_6t
Xbit_r74_c9 bl[9] br[9] wl[74] vdd gnd cell_6t
Xbit_r75_c9 bl[9] br[9] wl[75] vdd gnd cell_6t
Xbit_r76_c9 bl[9] br[9] wl[76] vdd gnd cell_6t
Xbit_r77_c9 bl[9] br[9] wl[77] vdd gnd cell_6t
Xbit_r78_c9 bl[9] br[9] wl[78] vdd gnd cell_6t
Xbit_r79_c9 bl[9] br[9] wl[79] vdd gnd cell_6t
Xbit_r80_c9 bl[9] br[9] wl[80] vdd gnd cell_6t
Xbit_r81_c9 bl[9] br[9] wl[81] vdd gnd cell_6t
Xbit_r82_c9 bl[9] br[9] wl[82] vdd gnd cell_6t
Xbit_r83_c9 bl[9] br[9] wl[83] vdd gnd cell_6t
Xbit_r84_c9 bl[9] br[9] wl[84] vdd gnd cell_6t
Xbit_r85_c9 bl[9] br[9] wl[85] vdd gnd cell_6t
Xbit_r86_c9 bl[9] br[9] wl[86] vdd gnd cell_6t
Xbit_r87_c9 bl[9] br[9] wl[87] vdd gnd cell_6t
Xbit_r88_c9 bl[9] br[9] wl[88] vdd gnd cell_6t
Xbit_r89_c9 bl[9] br[9] wl[89] vdd gnd cell_6t
Xbit_r90_c9 bl[9] br[9] wl[90] vdd gnd cell_6t
Xbit_r91_c9 bl[9] br[9] wl[91] vdd gnd cell_6t
Xbit_r92_c9 bl[9] br[9] wl[92] vdd gnd cell_6t
Xbit_r93_c9 bl[9] br[9] wl[93] vdd gnd cell_6t
Xbit_r94_c9 bl[9] br[9] wl[94] vdd gnd cell_6t
Xbit_r95_c9 bl[9] br[9] wl[95] vdd gnd cell_6t
Xbit_r96_c9 bl[9] br[9] wl[96] vdd gnd cell_6t
Xbit_r97_c9 bl[9] br[9] wl[97] vdd gnd cell_6t
Xbit_r98_c9 bl[9] br[9] wl[98] vdd gnd cell_6t
Xbit_r99_c9 bl[9] br[9] wl[99] vdd gnd cell_6t
Xbit_r100_c9 bl[9] br[9] wl[100] vdd gnd cell_6t
Xbit_r101_c9 bl[9] br[9] wl[101] vdd gnd cell_6t
Xbit_r102_c9 bl[9] br[9] wl[102] vdd gnd cell_6t
Xbit_r103_c9 bl[9] br[9] wl[103] vdd gnd cell_6t
Xbit_r104_c9 bl[9] br[9] wl[104] vdd gnd cell_6t
Xbit_r105_c9 bl[9] br[9] wl[105] vdd gnd cell_6t
Xbit_r106_c9 bl[9] br[9] wl[106] vdd gnd cell_6t
Xbit_r107_c9 bl[9] br[9] wl[107] vdd gnd cell_6t
Xbit_r108_c9 bl[9] br[9] wl[108] vdd gnd cell_6t
Xbit_r109_c9 bl[9] br[9] wl[109] vdd gnd cell_6t
Xbit_r110_c9 bl[9] br[9] wl[110] vdd gnd cell_6t
Xbit_r111_c9 bl[9] br[9] wl[111] vdd gnd cell_6t
Xbit_r112_c9 bl[9] br[9] wl[112] vdd gnd cell_6t
Xbit_r113_c9 bl[9] br[9] wl[113] vdd gnd cell_6t
Xbit_r114_c9 bl[9] br[9] wl[114] vdd gnd cell_6t
Xbit_r115_c9 bl[9] br[9] wl[115] vdd gnd cell_6t
Xbit_r116_c9 bl[9] br[9] wl[116] vdd gnd cell_6t
Xbit_r117_c9 bl[9] br[9] wl[117] vdd gnd cell_6t
Xbit_r118_c9 bl[9] br[9] wl[118] vdd gnd cell_6t
Xbit_r119_c9 bl[9] br[9] wl[119] vdd gnd cell_6t
Xbit_r120_c9 bl[9] br[9] wl[120] vdd gnd cell_6t
Xbit_r121_c9 bl[9] br[9] wl[121] vdd gnd cell_6t
Xbit_r122_c9 bl[9] br[9] wl[122] vdd gnd cell_6t
Xbit_r123_c9 bl[9] br[9] wl[123] vdd gnd cell_6t
Xbit_r124_c9 bl[9] br[9] wl[124] vdd gnd cell_6t
Xbit_r125_c9 bl[9] br[9] wl[125] vdd gnd cell_6t
Xbit_r126_c9 bl[9] br[9] wl[126] vdd gnd cell_6t
Xbit_r127_c9 bl[9] br[9] wl[127] vdd gnd cell_6t
Xbit_r128_c9 bl[9] br[9] wl[128] vdd gnd cell_6t
Xbit_r129_c9 bl[9] br[9] wl[129] vdd gnd cell_6t
Xbit_r130_c9 bl[9] br[9] wl[130] vdd gnd cell_6t
Xbit_r131_c9 bl[9] br[9] wl[131] vdd gnd cell_6t
Xbit_r132_c9 bl[9] br[9] wl[132] vdd gnd cell_6t
Xbit_r133_c9 bl[9] br[9] wl[133] vdd gnd cell_6t
Xbit_r134_c9 bl[9] br[9] wl[134] vdd gnd cell_6t
Xbit_r135_c9 bl[9] br[9] wl[135] vdd gnd cell_6t
Xbit_r136_c9 bl[9] br[9] wl[136] vdd gnd cell_6t
Xbit_r137_c9 bl[9] br[9] wl[137] vdd gnd cell_6t
Xbit_r138_c9 bl[9] br[9] wl[138] vdd gnd cell_6t
Xbit_r139_c9 bl[9] br[9] wl[139] vdd gnd cell_6t
Xbit_r140_c9 bl[9] br[9] wl[140] vdd gnd cell_6t
Xbit_r141_c9 bl[9] br[9] wl[141] vdd gnd cell_6t
Xbit_r142_c9 bl[9] br[9] wl[142] vdd gnd cell_6t
Xbit_r143_c9 bl[9] br[9] wl[143] vdd gnd cell_6t
Xbit_r144_c9 bl[9] br[9] wl[144] vdd gnd cell_6t
Xbit_r145_c9 bl[9] br[9] wl[145] vdd gnd cell_6t
Xbit_r146_c9 bl[9] br[9] wl[146] vdd gnd cell_6t
Xbit_r147_c9 bl[9] br[9] wl[147] vdd gnd cell_6t
Xbit_r148_c9 bl[9] br[9] wl[148] vdd gnd cell_6t
Xbit_r149_c9 bl[9] br[9] wl[149] vdd gnd cell_6t
Xbit_r150_c9 bl[9] br[9] wl[150] vdd gnd cell_6t
Xbit_r151_c9 bl[9] br[9] wl[151] vdd gnd cell_6t
Xbit_r152_c9 bl[9] br[9] wl[152] vdd gnd cell_6t
Xbit_r153_c9 bl[9] br[9] wl[153] vdd gnd cell_6t
Xbit_r154_c9 bl[9] br[9] wl[154] vdd gnd cell_6t
Xbit_r155_c9 bl[9] br[9] wl[155] vdd gnd cell_6t
Xbit_r156_c9 bl[9] br[9] wl[156] vdd gnd cell_6t
Xbit_r157_c9 bl[9] br[9] wl[157] vdd gnd cell_6t
Xbit_r158_c9 bl[9] br[9] wl[158] vdd gnd cell_6t
Xbit_r159_c9 bl[9] br[9] wl[159] vdd gnd cell_6t
Xbit_r160_c9 bl[9] br[9] wl[160] vdd gnd cell_6t
Xbit_r161_c9 bl[9] br[9] wl[161] vdd gnd cell_6t
Xbit_r162_c9 bl[9] br[9] wl[162] vdd gnd cell_6t
Xbit_r163_c9 bl[9] br[9] wl[163] vdd gnd cell_6t
Xbit_r164_c9 bl[9] br[9] wl[164] vdd gnd cell_6t
Xbit_r165_c9 bl[9] br[9] wl[165] vdd gnd cell_6t
Xbit_r166_c9 bl[9] br[9] wl[166] vdd gnd cell_6t
Xbit_r167_c9 bl[9] br[9] wl[167] vdd gnd cell_6t
Xbit_r168_c9 bl[9] br[9] wl[168] vdd gnd cell_6t
Xbit_r169_c9 bl[9] br[9] wl[169] vdd gnd cell_6t
Xbit_r170_c9 bl[9] br[9] wl[170] vdd gnd cell_6t
Xbit_r171_c9 bl[9] br[9] wl[171] vdd gnd cell_6t
Xbit_r172_c9 bl[9] br[9] wl[172] vdd gnd cell_6t
Xbit_r173_c9 bl[9] br[9] wl[173] vdd gnd cell_6t
Xbit_r174_c9 bl[9] br[9] wl[174] vdd gnd cell_6t
Xbit_r175_c9 bl[9] br[9] wl[175] vdd gnd cell_6t
Xbit_r176_c9 bl[9] br[9] wl[176] vdd gnd cell_6t
Xbit_r177_c9 bl[9] br[9] wl[177] vdd gnd cell_6t
Xbit_r178_c9 bl[9] br[9] wl[178] vdd gnd cell_6t
Xbit_r179_c9 bl[9] br[9] wl[179] vdd gnd cell_6t
Xbit_r180_c9 bl[9] br[9] wl[180] vdd gnd cell_6t
Xbit_r181_c9 bl[9] br[9] wl[181] vdd gnd cell_6t
Xbit_r182_c9 bl[9] br[9] wl[182] vdd gnd cell_6t
Xbit_r183_c9 bl[9] br[9] wl[183] vdd gnd cell_6t
Xbit_r184_c9 bl[9] br[9] wl[184] vdd gnd cell_6t
Xbit_r185_c9 bl[9] br[9] wl[185] vdd gnd cell_6t
Xbit_r186_c9 bl[9] br[9] wl[186] vdd gnd cell_6t
Xbit_r187_c9 bl[9] br[9] wl[187] vdd gnd cell_6t
Xbit_r188_c9 bl[9] br[9] wl[188] vdd gnd cell_6t
Xbit_r189_c9 bl[9] br[9] wl[189] vdd gnd cell_6t
Xbit_r190_c9 bl[9] br[9] wl[190] vdd gnd cell_6t
Xbit_r191_c9 bl[9] br[9] wl[191] vdd gnd cell_6t
Xbit_r192_c9 bl[9] br[9] wl[192] vdd gnd cell_6t
Xbit_r193_c9 bl[9] br[9] wl[193] vdd gnd cell_6t
Xbit_r194_c9 bl[9] br[9] wl[194] vdd gnd cell_6t
Xbit_r195_c9 bl[9] br[9] wl[195] vdd gnd cell_6t
Xbit_r196_c9 bl[9] br[9] wl[196] vdd gnd cell_6t
Xbit_r197_c9 bl[9] br[9] wl[197] vdd gnd cell_6t
Xbit_r198_c9 bl[9] br[9] wl[198] vdd gnd cell_6t
Xbit_r199_c9 bl[9] br[9] wl[199] vdd gnd cell_6t
Xbit_r200_c9 bl[9] br[9] wl[200] vdd gnd cell_6t
Xbit_r201_c9 bl[9] br[9] wl[201] vdd gnd cell_6t
Xbit_r202_c9 bl[9] br[9] wl[202] vdd gnd cell_6t
Xbit_r203_c9 bl[9] br[9] wl[203] vdd gnd cell_6t
Xbit_r204_c9 bl[9] br[9] wl[204] vdd gnd cell_6t
Xbit_r205_c9 bl[9] br[9] wl[205] vdd gnd cell_6t
Xbit_r206_c9 bl[9] br[9] wl[206] vdd gnd cell_6t
Xbit_r207_c9 bl[9] br[9] wl[207] vdd gnd cell_6t
Xbit_r208_c9 bl[9] br[9] wl[208] vdd gnd cell_6t
Xbit_r209_c9 bl[9] br[9] wl[209] vdd gnd cell_6t
Xbit_r210_c9 bl[9] br[9] wl[210] vdd gnd cell_6t
Xbit_r211_c9 bl[9] br[9] wl[211] vdd gnd cell_6t
Xbit_r212_c9 bl[9] br[9] wl[212] vdd gnd cell_6t
Xbit_r213_c9 bl[9] br[9] wl[213] vdd gnd cell_6t
Xbit_r214_c9 bl[9] br[9] wl[214] vdd gnd cell_6t
Xbit_r215_c9 bl[9] br[9] wl[215] vdd gnd cell_6t
Xbit_r216_c9 bl[9] br[9] wl[216] vdd gnd cell_6t
Xbit_r217_c9 bl[9] br[9] wl[217] vdd gnd cell_6t
Xbit_r218_c9 bl[9] br[9] wl[218] vdd gnd cell_6t
Xbit_r219_c9 bl[9] br[9] wl[219] vdd gnd cell_6t
Xbit_r220_c9 bl[9] br[9] wl[220] vdd gnd cell_6t
Xbit_r221_c9 bl[9] br[9] wl[221] vdd gnd cell_6t
Xbit_r222_c9 bl[9] br[9] wl[222] vdd gnd cell_6t
Xbit_r223_c9 bl[9] br[9] wl[223] vdd gnd cell_6t
Xbit_r224_c9 bl[9] br[9] wl[224] vdd gnd cell_6t
Xbit_r225_c9 bl[9] br[9] wl[225] vdd gnd cell_6t
Xbit_r226_c9 bl[9] br[9] wl[226] vdd gnd cell_6t
Xbit_r227_c9 bl[9] br[9] wl[227] vdd gnd cell_6t
Xbit_r228_c9 bl[9] br[9] wl[228] vdd gnd cell_6t
Xbit_r229_c9 bl[9] br[9] wl[229] vdd gnd cell_6t
Xbit_r230_c9 bl[9] br[9] wl[230] vdd gnd cell_6t
Xbit_r231_c9 bl[9] br[9] wl[231] vdd gnd cell_6t
Xbit_r232_c9 bl[9] br[9] wl[232] vdd gnd cell_6t
Xbit_r233_c9 bl[9] br[9] wl[233] vdd gnd cell_6t
Xbit_r234_c9 bl[9] br[9] wl[234] vdd gnd cell_6t
Xbit_r235_c9 bl[9] br[9] wl[235] vdd gnd cell_6t
Xbit_r236_c9 bl[9] br[9] wl[236] vdd gnd cell_6t
Xbit_r237_c9 bl[9] br[9] wl[237] vdd gnd cell_6t
Xbit_r238_c9 bl[9] br[9] wl[238] vdd gnd cell_6t
Xbit_r239_c9 bl[9] br[9] wl[239] vdd gnd cell_6t
Xbit_r240_c9 bl[9] br[9] wl[240] vdd gnd cell_6t
Xbit_r241_c9 bl[9] br[9] wl[241] vdd gnd cell_6t
Xbit_r242_c9 bl[9] br[9] wl[242] vdd gnd cell_6t
Xbit_r243_c9 bl[9] br[9] wl[243] vdd gnd cell_6t
Xbit_r244_c9 bl[9] br[9] wl[244] vdd gnd cell_6t
Xbit_r245_c9 bl[9] br[9] wl[245] vdd gnd cell_6t
Xbit_r246_c9 bl[9] br[9] wl[246] vdd gnd cell_6t
Xbit_r247_c9 bl[9] br[9] wl[247] vdd gnd cell_6t
Xbit_r248_c9 bl[9] br[9] wl[248] vdd gnd cell_6t
Xbit_r249_c9 bl[9] br[9] wl[249] vdd gnd cell_6t
Xbit_r250_c9 bl[9] br[9] wl[250] vdd gnd cell_6t
Xbit_r251_c9 bl[9] br[9] wl[251] vdd gnd cell_6t
Xbit_r252_c9 bl[9] br[9] wl[252] vdd gnd cell_6t
Xbit_r253_c9 bl[9] br[9] wl[253] vdd gnd cell_6t
Xbit_r254_c9 bl[9] br[9] wl[254] vdd gnd cell_6t
Xbit_r255_c9 bl[9] br[9] wl[255] vdd gnd cell_6t
Xbit_r0_c10 bl[10] br[10] wl[0] vdd gnd cell_6t
Xbit_r1_c10 bl[10] br[10] wl[1] vdd gnd cell_6t
Xbit_r2_c10 bl[10] br[10] wl[2] vdd gnd cell_6t
Xbit_r3_c10 bl[10] br[10] wl[3] vdd gnd cell_6t
Xbit_r4_c10 bl[10] br[10] wl[4] vdd gnd cell_6t
Xbit_r5_c10 bl[10] br[10] wl[5] vdd gnd cell_6t
Xbit_r6_c10 bl[10] br[10] wl[6] vdd gnd cell_6t
Xbit_r7_c10 bl[10] br[10] wl[7] vdd gnd cell_6t
Xbit_r8_c10 bl[10] br[10] wl[8] vdd gnd cell_6t
Xbit_r9_c10 bl[10] br[10] wl[9] vdd gnd cell_6t
Xbit_r10_c10 bl[10] br[10] wl[10] vdd gnd cell_6t
Xbit_r11_c10 bl[10] br[10] wl[11] vdd gnd cell_6t
Xbit_r12_c10 bl[10] br[10] wl[12] vdd gnd cell_6t
Xbit_r13_c10 bl[10] br[10] wl[13] vdd gnd cell_6t
Xbit_r14_c10 bl[10] br[10] wl[14] vdd gnd cell_6t
Xbit_r15_c10 bl[10] br[10] wl[15] vdd gnd cell_6t
Xbit_r16_c10 bl[10] br[10] wl[16] vdd gnd cell_6t
Xbit_r17_c10 bl[10] br[10] wl[17] vdd gnd cell_6t
Xbit_r18_c10 bl[10] br[10] wl[18] vdd gnd cell_6t
Xbit_r19_c10 bl[10] br[10] wl[19] vdd gnd cell_6t
Xbit_r20_c10 bl[10] br[10] wl[20] vdd gnd cell_6t
Xbit_r21_c10 bl[10] br[10] wl[21] vdd gnd cell_6t
Xbit_r22_c10 bl[10] br[10] wl[22] vdd gnd cell_6t
Xbit_r23_c10 bl[10] br[10] wl[23] vdd gnd cell_6t
Xbit_r24_c10 bl[10] br[10] wl[24] vdd gnd cell_6t
Xbit_r25_c10 bl[10] br[10] wl[25] vdd gnd cell_6t
Xbit_r26_c10 bl[10] br[10] wl[26] vdd gnd cell_6t
Xbit_r27_c10 bl[10] br[10] wl[27] vdd gnd cell_6t
Xbit_r28_c10 bl[10] br[10] wl[28] vdd gnd cell_6t
Xbit_r29_c10 bl[10] br[10] wl[29] vdd gnd cell_6t
Xbit_r30_c10 bl[10] br[10] wl[30] vdd gnd cell_6t
Xbit_r31_c10 bl[10] br[10] wl[31] vdd gnd cell_6t
Xbit_r32_c10 bl[10] br[10] wl[32] vdd gnd cell_6t
Xbit_r33_c10 bl[10] br[10] wl[33] vdd gnd cell_6t
Xbit_r34_c10 bl[10] br[10] wl[34] vdd gnd cell_6t
Xbit_r35_c10 bl[10] br[10] wl[35] vdd gnd cell_6t
Xbit_r36_c10 bl[10] br[10] wl[36] vdd gnd cell_6t
Xbit_r37_c10 bl[10] br[10] wl[37] vdd gnd cell_6t
Xbit_r38_c10 bl[10] br[10] wl[38] vdd gnd cell_6t
Xbit_r39_c10 bl[10] br[10] wl[39] vdd gnd cell_6t
Xbit_r40_c10 bl[10] br[10] wl[40] vdd gnd cell_6t
Xbit_r41_c10 bl[10] br[10] wl[41] vdd gnd cell_6t
Xbit_r42_c10 bl[10] br[10] wl[42] vdd gnd cell_6t
Xbit_r43_c10 bl[10] br[10] wl[43] vdd gnd cell_6t
Xbit_r44_c10 bl[10] br[10] wl[44] vdd gnd cell_6t
Xbit_r45_c10 bl[10] br[10] wl[45] vdd gnd cell_6t
Xbit_r46_c10 bl[10] br[10] wl[46] vdd gnd cell_6t
Xbit_r47_c10 bl[10] br[10] wl[47] vdd gnd cell_6t
Xbit_r48_c10 bl[10] br[10] wl[48] vdd gnd cell_6t
Xbit_r49_c10 bl[10] br[10] wl[49] vdd gnd cell_6t
Xbit_r50_c10 bl[10] br[10] wl[50] vdd gnd cell_6t
Xbit_r51_c10 bl[10] br[10] wl[51] vdd gnd cell_6t
Xbit_r52_c10 bl[10] br[10] wl[52] vdd gnd cell_6t
Xbit_r53_c10 bl[10] br[10] wl[53] vdd gnd cell_6t
Xbit_r54_c10 bl[10] br[10] wl[54] vdd gnd cell_6t
Xbit_r55_c10 bl[10] br[10] wl[55] vdd gnd cell_6t
Xbit_r56_c10 bl[10] br[10] wl[56] vdd gnd cell_6t
Xbit_r57_c10 bl[10] br[10] wl[57] vdd gnd cell_6t
Xbit_r58_c10 bl[10] br[10] wl[58] vdd gnd cell_6t
Xbit_r59_c10 bl[10] br[10] wl[59] vdd gnd cell_6t
Xbit_r60_c10 bl[10] br[10] wl[60] vdd gnd cell_6t
Xbit_r61_c10 bl[10] br[10] wl[61] vdd gnd cell_6t
Xbit_r62_c10 bl[10] br[10] wl[62] vdd gnd cell_6t
Xbit_r63_c10 bl[10] br[10] wl[63] vdd gnd cell_6t
Xbit_r64_c10 bl[10] br[10] wl[64] vdd gnd cell_6t
Xbit_r65_c10 bl[10] br[10] wl[65] vdd gnd cell_6t
Xbit_r66_c10 bl[10] br[10] wl[66] vdd gnd cell_6t
Xbit_r67_c10 bl[10] br[10] wl[67] vdd gnd cell_6t
Xbit_r68_c10 bl[10] br[10] wl[68] vdd gnd cell_6t
Xbit_r69_c10 bl[10] br[10] wl[69] vdd gnd cell_6t
Xbit_r70_c10 bl[10] br[10] wl[70] vdd gnd cell_6t
Xbit_r71_c10 bl[10] br[10] wl[71] vdd gnd cell_6t
Xbit_r72_c10 bl[10] br[10] wl[72] vdd gnd cell_6t
Xbit_r73_c10 bl[10] br[10] wl[73] vdd gnd cell_6t
Xbit_r74_c10 bl[10] br[10] wl[74] vdd gnd cell_6t
Xbit_r75_c10 bl[10] br[10] wl[75] vdd gnd cell_6t
Xbit_r76_c10 bl[10] br[10] wl[76] vdd gnd cell_6t
Xbit_r77_c10 bl[10] br[10] wl[77] vdd gnd cell_6t
Xbit_r78_c10 bl[10] br[10] wl[78] vdd gnd cell_6t
Xbit_r79_c10 bl[10] br[10] wl[79] vdd gnd cell_6t
Xbit_r80_c10 bl[10] br[10] wl[80] vdd gnd cell_6t
Xbit_r81_c10 bl[10] br[10] wl[81] vdd gnd cell_6t
Xbit_r82_c10 bl[10] br[10] wl[82] vdd gnd cell_6t
Xbit_r83_c10 bl[10] br[10] wl[83] vdd gnd cell_6t
Xbit_r84_c10 bl[10] br[10] wl[84] vdd gnd cell_6t
Xbit_r85_c10 bl[10] br[10] wl[85] vdd gnd cell_6t
Xbit_r86_c10 bl[10] br[10] wl[86] vdd gnd cell_6t
Xbit_r87_c10 bl[10] br[10] wl[87] vdd gnd cell_6t
Xbit_r88_c10 bl[10] br[10] wl[88] vdd gnd cell_6t
Xbit_r89_c10 bl[10] br[10] wl[89] vdd gnd cell_6t
Xbit_r90_c10 bl[10] br[10] wl[90] vdd gnd cell_6t
Xbit_r91_c10 bl[10] br[10] wl[91] vdd gnd cell_6t
Xbit_r92_c10 bl[10] br[10] wl[92] vdd gnd cell_6t
Xbit_r93_c10 bl[10] br[10] wl[93] vdd gnd cell_6t
Xbit_r94_c10 bl[10] br[10] wl[94] vdd gnd cell_6t
Xbit_r95_c10 bl[10] br[10] wl[95] vdd gnd cell_6t
Xbit_r96_c10 bl[10] br[10] wl[96] vdd gnd cell_6t
Xbit_r97_c10 bl[10] br[10] wl[97] vdd gnd cell_6t
Xbit_r98_c10 bl[10] br[10] wl[98] vdd gnd cell_6t
Xbit_r99_c10 bl[10] br[10] wl[99] vdd gnd cell_6t
Xbit_r100_c10 bl[10] br[10] wl[100] vdd gnd cell_6t
Xbit_r101_c10 bl[10] br[10] wl[101] vdd gnd cell_6t
Xbit_r102_c10 bl[10] br[10] wl[102] vdd gnd cell_6t
Xbit_r103_c10 bl[10] br[10] wl[103] vdd gnd cell_6t
Xbit_r104_c10 bl[10] br[10] wl[104] vdd gnd cell_6t
Xbit_r105_c10 bl[10] br[10] wl[105] vdd gnd cell_6t
Xbit_r106_c10 bl[10] br[10] wl[106] vdd gnd cell_6t
Xbit_r107_c10 bl[10] br[10] wl[107] vdd gnd cell_6t
Xbit_r108_c10 bl[10] br[10] wl[108] vdd gnd cell_6t
Xbit_r109_c10 bl[10] br[10] wl[109] vdd gnd cell_6t
Xbit_r110_c10 bl[10] br[10] wl[110] vdd gnd cell_6t
Xbit_r111_c10 bl[10] br[10] wl[111] vdd gnd cell_6t
Xbit_r112_c10 bl[10] br[10] wl[112] vdd gnd cell_6t
Xbit_r113_c10 bl[10] br[10] wl[113] vdd gnd cell_6t
Xbit_r114_c10 bl[10] br[10] wl[114] vdd gnd cell_6t
Xbit_r115_c10 bl[10] br[10] wl[115] vdd gnd cell_6t
Xbit_r116_c10 bl[10] br[10] wl[116] vdd gnd cell_6t
Xbit_r117_c10 bl[10] br[10] wl[117] vdd gnd cell_6t
Xbit_r118_c10 bl[10] br[10] wl[118] vdd gnd cell_6t
Xbit_r119_c10 bl[10] br[10] wl[119] vdd gnd cell_6t
Xbit_r120_c10 bl[10] br[10] wl[120] vdd gnd cell_6t
Xbit_r121_c10 bl[10] br[10] wl[121] vdd gnd cell_6t
Xbit_r122_c10 bl[10] br[10] wl[122] vdd gnd cell_6t
Xbit_r123_c10 bl[10] br[10] wl[123] vdd gnd cell_6t
Xbit_r124_c10 bl[10] br[10] wl[124] vdd gnd cell_6t
Xbit_r125_c10 bl[10] br[10] wl[125] vdd gnd cell_6t
Xbit_r126_c10 bl[10] br[10] wl[126] vdd gnd cell_6t
Xbit_r127_c10 bl[10] br[10] wl[127] vdd gnd cell_6t
Xbit_r128_c10 bl[10] br[10] wl[128] vdd gnd cell_6t
Xbit_r129_c10 bl[10] br[10] wl[129] vdd gnd cell_6t
Xbit_r130_c10 bl[10] br[10] wl[130] vdd gnd cell_6t
Xbit_r131_c10 bl[10] br[10] wl[131] vdd gnd cell_6t
Xbit_r132_c10 bl[10] br[10] wl[132] vdd gnd cell_6t
Xbit_r133_c10 bl[10] br[10] wl[133] vdd gnd cell_6t
Xbit_r134_c10 bl[10] br[10] wl[134] vdd gnd cell_6t
Xbit_r135_c10 bl[10] br[10] wl[135] vdd gnd cell_6t
Xbit_r136_c10 bl[10] br[10] wl[136] vdd gnd cell_6t
Xbit_r137_c10 bl[10] br[10] wl[137] vdd gnd cell_6t
Xbit_r138_c10 bl[10] br[10] wl[138] vdd gnd cell_6t
Xbit_r139_c10 bl[10] br[10] wl[139] vdd gnd cell_6t
Xbit_r140_c10 bl[10] br[10] wl[140] vdd gnd cell_6t
Xbit_r141_c10 bl[10] br[10] wl[141] vdd gnd cell_6t
Xbit_r142_c10 bl[10] br[10] wl[142] vdd gnd cell_6t
Xbit_r143_c10 bl[10] br[10] wl[143] vdd gnd cell_6t
Xbit_r144_c10 bl[10] br[10] wl[144] vdd gnd cell_6t
Xbit_r145_c10 bl[10] br[10] wl[145] vdd gnd cell_6t
Xbit_r146_c10 bl[10] br[10] wl[146] vdd gnd cell_6t
Xbit_r147_c10 bl[10] br[10] wl[147] vdd gnd cell_6t
Xbit_r148_c10 bl[10] br[10] wl[148] vdd gnd cell_6t
Xbit_r149_c10 bl[10] br[10] wl[149] vdd gnd cell_6t
Xbit_r150_c10 bl[10] br[10] wl[150] vdd gnd cell_6t
Xbit_r151_c10 bl[10] br[10] wl[151] vdd gnd cell_6t
Xbit_r152_c10 bl[10] br[10] wl[152] vdd gnd cell_6t
Xbit_r153_c10 bl[10] br[10] wl[153] vdd gnd cell_6t
Xbit_r154_c10 bl[10] br[10] wl[154] vdd gnd cell_6t
Xbit_r155_c10 bl[10] br[10] wl[155] vdd gnd cell_6t
Xbit_r156_c10 bl[10] br[10] wl[156] vdd gnd cell_6t
Xbit_r157_c10 bl[10] br[10] wl[157] vdd gnd cell_6t
Xbit_r158_c10 bl[10] br[10] wl[158] vdd gnd cell_6t
Xbit_r159_c10 bl[10] br[10] wl[159] vdd gnd cell_6t
Xbit_r160_c10 bl[10] br[10] wl[160] vdd gnd cell_6t
Xbit_r161_c10 bl[10] br[10] wl[161] vdd gnd cell_6t
Xbit_r162_c10 bl[10] br[10] wl[162] vdd gnd cell_6t
Xbit_r163_c10 bl[10] br[10] wl[163] vdd gnd cell_6t
Xbit_r164_c10 bl[10] br[10] wl[164] vdd gnd cell_6t
Xbit_r165_c10 bl[10] br[10] wl[165] vdd gnd cell_6t
Xbit_r166_c10 bl[10] br[10] wl[166] vdd gnd cell_6t
Xbit_r167_c10 bl[10] br[10] wl[167] vdd gnd cell_6t
Xbit_r168_c10 bl[10] br[10] wl[168] vdd gnd cell_6t
Xbit_r169_c10 bl[10] br[10] wl[169] vdd gnd cell_6t
Xbit_r170_c10 bl[10] br[10] wl[170] vdd gnd cell_6t
Xbit_r171_c10 bl[10] br[10] wl[171] vdd gnd cell_6t
Xbit_r172_c10 bl[10] br[10] wl[172] vdd gnd cell_6t
Xbit_r173_c10 bl[10] br[10] wl[173] vdd gnd cell_6t
Xbit_r174_c10 bl[10] br[10] wl[174] vdd gnd cell_6t
Xbit_r175_c10 bl[10] br[10] wl[175] vdd gnd cell_6t
Xbit_r176_c10 bl[10] br[10] wl[176] vdd gnd cell_6t
Xbit_r177_c10 bl[10] br[10] wl[177] vdd gnd cell_6t
Xbit_r178_c10 bl[10] br[10] wl[178] vdd gnd cell_6t
Xbit_r179_c10 bl[10] br[10] wl[179] vdd gnd cell_6t
Xbit_r180_c10 bl[10] br[10] wl[180] vdd gnd cell_6t
Xbit_r181_c10 bl[10] br[10] wl[181] vdd gnd cell_6t
Xbit_r182_c10 bl[10] br[10] wl[182] vdd gnd cell_6t
Xbit_r183_c10 bl[10] br[10] wl[183] vdd gnd cell_6t
Xbit_r184_c10 bl[10] br[10] wl[184] vdd gnd cell_6t
Xbit_r185_c10 bl[10] br[10] wl[185] vdd gnd cell_6t
Xbit_r186_c10 bl[10] br[10] wl[186] vdd gnd cell_6t
Xbit_r187_c10 bl[10] br[10] wl[187] vdd gnd cell_6t
Xbit_r188_c10 bl[10] br[10] wl[188] vdd gnd cell_6t
Xbit_r189_c10 bl[10] br[10] wl[189] vdd gnd cell_6t
Xbit_r190_c10 bl[10] br[10] wl[190] vdd gnd cell_6t
Xbit_r191_c10 bl[10] br[10] wl[191] vdd gnd cell_6t
Xbit_r192_c10 bl[10] br[10] wl[192] vdd gnd cell_6t
Xbit_r193_c10 bl[10] br[10] wl[193] vdd gnd cell_6t
Xbit_r194_c10 bl[10] br[10] wl[194] vdd gnd cell_6t
Xbit_r195_c10 bl[10] br[10] wl[195] vdd gnd cell_6t
Xbit_r196_c10 bl[10] br[10] wl[196] vdd gnd cell_6t
Xbit_r197_c10 bl[10] br[10] wl[197] vdd gnd cell_6t
Xbit_r198_c10 bl[10] br[10] wl[198] vdd gnd cell_6t
Xbit_r199_c10 bl[10] br[10] wl[199] vdd gnd cell_6t
Xbit_r200_c10 bl[10] br[10] wl[200] vdd gnd cell_6t
Xbit_r201_c10 bl[10] br[10] wl[201] vdd gnd cell_6t
Xbit_r202_c10 bl[10] br[10] wl[202] vdd gnd cell_6t
Xbit_r203_c10 bl[10] br[10] wl[203] vdd gnd cell_6t
Xbit_r204_c10 bl[10] br[10] wl[204] vdd gnd cell_6t
Xbit_r205_c10 bl[10] br[10] wl[205] vdd gnd cell_6t
Xbit_r206_c10 bl[10] br[10] wl[206] vdd gnd cell_6t
Xbit_r207_c10 bl[10] br[10] wl[207] vdd gnd cell_6t
Xbit_r208_c10 bl[10] br[10] wl[208] vdd gnd cell_6t
Xbit_r209_c10 bl[10] br[10] wl[209] vdd gnd cell_6t
Xbit_r210_c10 bl[10] br[10] wl[210] vdd gnd cell_6t
Xbit_r211_c10 bl[10] br[10] wl[211] vdd gnd cell_6t
Xbit_r212_c10 bl[10] br[10] wl[212] vdd gnd cell_6t
Xbit_r213_c10 bl[10] br[10] wl[213] vdd gnd cell_6t
Xbit_r214_c10 bl[10] br[10] wl[214] vdd gnd cell_6t
Xbit_r215_c10 bl[10] br[10] wl[215] vdd gnd cell_6t
Xbit_r216_c10 bl[10] br[10] wl[216] vdd gnd cell_6t
Xbit_r217_c10 bl[10] br[10] wl[217] vdd gnd cell_6t
Xbit_r218_c10 bl[10] br[10] wl[218] vdd gnd cell_6t
Xbit_r219_c10 bl[10] br[10] wl[219] vdd gnd cell_6t
Xbit_r220_c10 bl[10] br[10] wl[220] vdd gnd cell_6t
Xbit_r221_c10 bl[10] br[10] wl[221] vdd gnd cell_6t
Xbit_r222_c10 bl[10] br[10] wl[222] vdd gnd cell_6t
Xbit_r223_c10 bl[10] br[10] wl[223] vdd gnd cell_6t
Xbit_r224_c10 bl[10] br[10] wl[224] vdd gnd cell_6t
Xbit_r225_c10 bl[10] br[10] wl[225] vdd gnd cell_6t
Xbit_r226_c10 bl[10] br[10] wl[226] vdd gnd cell_6t
Xbit_r227_c10 bl[10] br[10] wl[227] vdd gnd cell_6t
Xbit_r228_c10 bl[10] br[10] wl[228] vdd gnd cell_6t
Xbit_r229_c10 bl[10] br[10] wl[229] vdd gnd cell_6t
Xbit_r230_c10 bl[10] br[10] wl[230] vdd gnd cell_6t
Xbit_r231_c10 bl[10] br[10] wl[231] vdd gnd cell_6t
Xbit_r232_c10 bl[10] br[10] wl[232] vdd gnd cell_6t
Xbit_r233_c10 bl[10] br[10] wl[233] vdd gnd cell_6t
Xbit_r234_c10 bl[10] br[10] wl[234] vdd gnd cell_6t
Xbit_r235_c10 bl[10] br[10] wl[235] vdd gnd cell_6t
Xbit_r236_c10 bl[10] br[10] wl[236] vdd gnd cell_6t
Xbit_r237_c10 bl[10] br[10] wl[237] vdd gnd cell_6t
Xbit_r238_c10 bl[10] br[10] wl[238] vdd gnd cell_6t
Xbit_r239_c10 bl[10] br[10] wl[239] vdd gnd cell_6t
Xbit_r240_c10 bl[10] br[10] wl[240] vdd gnd cell_6t
Xbit_r241_c10 bl[10] br[10] wl[241] vdd gnd cell_6t
Xbit_r242_c10 bl[10] br[10] wl[242] vdd gnd cell_6t
Xbit_r243_c10 bl[10] br[10] wl[243] vdd gnd cell_6t
Xbit_r244_c10 bl[10] br[10] wl[244] vdd gnd cell_6t
Xbit_r245_c10 bl[10] br[10] wl[245] vdd gnd cell_6t
Xbit_r246_c10 bl[10] br[10] wl[246] vdd gnd cell_6t
Xbit_r247_c10 bl[10] br[10] wl[247] vdd gnd cell_6t
Xbit_r248_c10 bl[10] br[10] wl[248] vdd gnd cell_6t
Xbit_r249_c10 bl[10] br[10] wl[249] vdd gnd cell_6t
Xbit_r250_c10 bl[10] br[10] wl[250] vdd gnd cell_6t
Xbit_r251_c10 bl[10] br[10] wl[251] vdd gnd cell_6t
Xbit_r252_c10 bl[10] br[10] wl[252] vdd gnd cell_6t
Xbit_r253_c10 bl[10] br[10] wl[253] vdd gnd cell_6t
Xbit_r254_c10 bl[10] br[10] wl[254] vdd gnd cell_6t
Xbit_r255_c10 bl[10] br[10] wl[255] vdd gnd cell_6t
Xbit_r0_c11 bl[11] br[11] wl[0] vdd gnd cell_6t
Xbit_r1_c11 bl[11] br[11] wl[1] vdd gnd cell_6t
Xbit_r2_c11 bl[11] br[11] wl[2] vdd gnd cell_6t
Xbit_r3_c11 bl[11] br[11] wl[3] vdd gnd cell_6t
Xbit_r4_c11 bl[11] br[11] wl[4] vdd gnd cell_6t
Xbit_r5_c11 bl[11] br[11] wl[5] vdd gnd cell_6t
Xbit_r6_c11 bl[11] br[11] wl[6] vdd gnd cell_6t
Xbit_r7_c11 bl[11] br[11] wl[7] vdd gnd cell_6t
Xbit_r8_c11 bl[11] br[11] wl[8] vdd gnd cell_6t
Xbit_r9_c11 bl[11] br[11] wl[9] vdd gnd cell_6t
Xbit_r10_c11 bl[11] br[11] wl[10] vdd gnd cell_6t
Xbit_r11_c11 bl[11] br[11] wl[11] vdd gnd cell_6t
Xbit_r12_c11 bl[11] br[11] wl[12] vdd gnd cell_6t
Xbit_r13_c11 bl[11] br[11] wl[13] vdd gnd cell_6t
Xbit_r14_c11 bl[11] br[11] wl[14] vdd gnd cell_6t
Xbit_r15_c11 bl[11] br[11] wl[15] vdd gnd cell_6t
Xbit_r16_c11 bl[11] br[11] wl[16] vdd gnd cell_6t
Xbit_r17_c11 bl[11] br[11] wl[17] vdd gnd cell_6t
Xbit_r18_c11 bl[11] br[11] wl[18] vdd gnd cell_6t
Xbit_r19_c11 bl[11] br[11] wl[19] vdd gnd cell_6t
Xbit_r20_c11 bl[11] br[11] wl[20] vdd gnd cell_6t
Xbit_r21_c11 bl[11] br[11] wl[21] vdd gnd cell_6t
Xbit_r22_c11 bl[11] br[11] wl[22] vdd gnd cell_6t
Xbit_r23_c11 bl[11] br[11] wl[23] vdd gnd cell_6t
Xbit_r24_c11 bl[11] br[11] wl[24] vdd gnd cell_6t
Xbit_r25_c11 bl[11] br[11] wl[25] vdd gnd cell_6t
Xbit_r26_c11 bl[11] br[11] wl[26] vdd gnd cell_6t
Xbit_r27_c11 bl[11] br[11] wl[27] vdd gnd cell_6t
Xbit_r28_c11 bl[11] br[11] wl[28] vdd gnd cell_6t
Xbit_r29_c11 bl[11] br[11] wl[29] vdd gnd cell_6t
Xbit_r30_c11 bl[11] br[11] wl[30] vdd gnd cell_6t
Xbit_r31_c11 bl[11] br[11] wl[31] vdd gnd cell_6t
Xbit_r32_c11 bl[11] br[11] wl[32] vdd gnd cell_6t
Xbit_r33_c11 bl[11] br[11] wl[33] vdd gnd cell_6t
Xbit_r34_c11 bl[11] br[11] wl[34] vdd gnd cell_6t
Xbit_r35_c11 bl[11] br[11] wl[35] vdd gnd cell_6t
Xbit_r36_c11 bl[11] br[11] wl[36] vdd gnd cell_6t
Xbit_r37_c11 bl[11] br[11] wl[37] vdd gnd cell_6t
Xbit_r38_c11 bl[11] br[11] wl[38] vdd gnd cell_6t
Xbit_r39_c11 bl[11] br[11] wl[39] vdd gnd cell_6t
Xbit_r40_c11 bl[11] br[11] wl[40] vdd gnd cell_6t
Xbit_r41_c11 bl[11] br[11] wl[41] vdd gnd cell_6t
Xbit_r42_c11 bl[11] br[11] wl[42] vdd gnd cell_6t
Xbit_r43_c11 bl[11] br[11] wl[43] vdd gnd cell_6t
Xbit_r44_c11 bl[11] br[11] wl[44] vdd gnd cell_6t
Xbit_r45_c11 bl[11] br[11] wl[45] vdd gnd cell_6t
Xbit_r46_c11 bl[11] br[11] wl[46] vdd gnd cell_6t
Xbit_r47_c11 bl[11] br[11] wl[47] vdd gnd cell_6t
Xbit_r48_c11 bl[11] br[11] wl[48] vdd gnd cell_6t
Xbit_r49_c11 bl[11] br[11] wl[49] vdd gnd cell_6t
Xbit_r50_c11 bl[11] br[11] wl[50] vdd gnd cell_6t
Xbit_r51_c11 bl[11] br[11] wl[51] vdd gnd cell_6t
Xbit_r52_c11 bl[11] br[11] wl[52] vdd gnd cell_6t
Xbit_r53_c11 bl[11] br[11] wl[53] vdd gnd cell_6t
Xbit_r54_c11 bl[11] br[11] wl[54] vdd gnd cell_6t
Xbit_r55_c11 bl[11] br[11] wl[55] vdd gnd cell_6t
Xbit_r56_c11 bl[11] br[11] wl[56] vdd gnd cell_6t
Xbit_r57_c11 bl[11] br[11] wl[57] vdd gnd cell_6t
Xbit_r58_c11 bl[11] br[11] wl[58] vdd gnd cell_6t
Xbit_r59_c11 bl[11] br[11] wl[59] vdd gnd cell_6t
Xbit_r60_c11 bl[11] br[11] wl[60] vdd gnd cell_6t
Xbit_r61_c11 bl[11] br[11] wl[61] vdd gnd cell_6t
Xbit_r62_c11 bl[11] br[11] wl[62] vdd gnd cell_6t
Xbit_r63_c11 bl[11] br[11] wl[63] vdd gnd cell_6t
Xbit_r64_c11 bl[11] br[11] wl[64] vdd gnd cell_6t
Xbit_r65_c11 bl[11] br[11] wl[65] vdd gnd cell_6t
Xbit_r66_c11 bl[11] br[11] wl[66] vdd gnd cell_6t
Xbit_r67_c11 bl[11] br[11] wl[67] vdd gnd cell_6t
Xbit_r68_c11 bl[11] br[11] wl[68] vdd gnd cell_6t
Xbit_r69_c11 bl[11] br[11] wl[69] vdd gnd cell_6t
Xbit_r70_c11 bl[11] br[11] wl[70] vdd gnd cell_6t
Xbit_r71_c11 bl[11] br[11] wl[71] vdd gnd cell_6t
Xbit_r72_c11 bl[11] br[11] wl[72] vdd gnd cell_6t
Xbit_r73_c11 bl[11] br[11] wl[73] vdd gnd cell_6t
Xbit_r74_c11 bl[11] br[11] wl[74] vdd gnd cell_6t
Xbit_r75_c11 bl[11] br[11] wl[75] vdd gnd cell_6t
Xbit_r76_c11 bl[11] br[11] wl[76] vdd gnd cell_6t
Xbit_r77_c11 bl[11] br[11] wl[77] vdd gnd cell_6t
Xbit_r78_c11 bl[11] br[11] wl[78] vdd gnd cell_6t
Xbit_r79_c11 bl[11] br[11] wl[79] vdd gnd cell_6t
Xbit_r80_c11 bl[11] br[11] wl[80] vdd gnd cell_6t
Xbit_r81_c11 bl[11] br[11] wl[81] vdd gnd cell_6t
Xbit_r82_c11 bl[11] br[11] wl[82] vdd gnd cell_6t
Xbit_r83_c11 bl[11] br[11] wl[83] vdd gnd cell_6t
Xbit_r84_c11 bl[11] br[11] wl[84] vdd gnd cell_6t
Xbit_r85_c11 bl[11] br[11] wl[85] vdd gnd cell_6t
Xbit_r86_c11 bl[11] br[11] wl[86] vdd gnd cell_6t
Xbit_r87_c11 bl[11] br[11] wl[87] vdd gnd cell_6t
Xbit_r88_c11 bl[11] br[11] wl[88] vdd gnd cell_6t
Xbit_r89_c11 bl[11] br[11] wl[89] vdd gnd cell_6t
Xbit_r90_c11 bl[11] br[11] wl[90] vdd gnd cell_6t
Xbit_r91_c11 bl[11] br[11] wl[91] vdd gnd cell_6t
Xbit_r92_c11 bl[11] br[11] wl[92] vdd gnd cell_6t
Xbit_r93_c11 bl[11] br[11] wl[93] vdd gnd cell_6t
Xbit_r94_c11 bl[11] br[11] wl[94] vdd gnd cell_6t
Xbit_r95_c11 bl[11] br[11] wl[95] vdd gnd cell_6t
Xbit_r96_c11 bl[11] br[11] wl[96] vdd gnd cell_6t
Xbit_r97_c11 bl[11] br[11] wl[97] vdd gnd cell_6t
Xbit_r98_c11 bl[11] br[11] wl[98] vdd gnd cell_6t
Xbit_r99_c11 bl[11] br[11] wl[99] vdd gnd cell_6t
Xbit_r100_c11 bl[11] br[11] wl[100] vdd gnd cell_6t
Xbit_r101_c11 bl[11] br[11] wl[101] vdd gnd cell_6t
Xbit_r102_c11 bl[11] br[11] wl[102] vdd gnd cell_6t
Xbit_r103_c11 bl[11] br[11] wl[103] vdd gnd cell_6t
Xbit_r104_c11 bl[11] br[11] wl[104] vdd gnd cell_6t
Xbit_r105_c11 bl[11] br[11] wl[105] vdd gnd cell_6t
Xbit_r106_c11 bl[11] br[11] wl[106] vdd gnd cell_6t
Xbit_r107_c11 bl[11] br[11] wl[107] vdd gnd cell_6t
Xbit_r108_c11 bl[11] br[11] wl[108] vdd gnd cell_6t
Xbit_r109_c11 bl[11] br[11] wl[109] vdd gnd cell_6t
Xbit_r110_c11 bl[11] br[11] wl[110] vdd gnd cell_6t
Xbit_r111_c11 bl[11] br[11] wl[111] vdd gnd cell_6t
Xbit_r112_c11 bl[11] br[11] wl[112] vdd gnd cell_6t
Xbit_r113_c11 bl[11] br[11] wl[113] vdd gnd cell_6t
Xbit_r114_c11 bl[11] br[11] wl[114] vdd gnd cell_6t
Xbit_r115_c11 bl[11] br[11] wl[115] vdd gnd cell_6t
Xbit_r116_c11 bl[11] br[11] wl[116] vdd gnd cell_6t
Xbit_r117_c11 bl[11] br[11] wl[117] vdd gnd cell_6t
Xbit_r118_c11 bl[11] br[11] wl[118] vdd gnd cell_6t
Xbit_r119_c11 bl[11] br[11] wl[119] vdd gnd cell_6t
Xbit_r120_c11 bl[11] br[11] wl[120] vdd gnd cell_6t
Xbit_r121_c11 bl[11] br[11] wl[121] vdd gnd cell_6t
Xbit_r122_c11 bl[11] br[11] wl[122] vdd gnd cell_6t
Xbit_r123_c11 bl[11] br[11] wl[123] vdd gnd cell_6t
Xbit_r124_c11 bl[11] br[11] wl[124] vdd gnd cell_6t
Xbit_r125_c11 bl[11] br[11] wl[125] vdd gnd cell_6t
Xbit_r126_c11 bl[11] br[11] wl[126] vdd gnd cell_6t
Xbit_r127_c11 bl[11] br[11] wl[127] vdd gnd cell_6t
Xbit_r128_c11 bl[11] br[11] wl[128] vdd gnd cell_6t
Xbit_r129_c11 bl[11] br[11] wl[129] vdd gnd cell_6t
Xbit_r130_c11 bl[11] br[11] wl[130] vdd gnd cell_6t
Xbit_r131_c11 bl[11] br[11] wl[131] vdd gnd cell_6t
Xbit_r132_c11 bl[11] br[11] wl[132] vdd gnd cell_6t
Xbit_r133_c11 bl[11] br[11] wl[133] vdd gnd cell_6t
Xbit_r134_c11 bl[11] br[11] wl[134] vdd gnd cell_6t
Xbit_r135_c11 bl[11] br[11] wl[135] vdd gnd cell_6t
Xbit_r136_c11 bl[11] br[11] wl[136] vdd gnd cell_6t
Xbit_r137_c11 bl[11] br[11] wl[137] vdd gnd cell_6t
Xbit_r138_c11 bl[11] br[11] wl[138] vdd gnd cell_6t
Xbit_r139_c11 bl[11] br[11] wl[139] vdd gnd cell_6t
Xbit_r140_c11 bl[11] br[11] wl[140] vdd gnd cell_6t
Xbit_r141_c11 bl[11] br[11] wl[141] vdd gnd cell_6t
Xbit_r142_c11 bl[11] br[11] wl[142] vdd gnd cell_6t
Xbit_r143_c11 bl[11] br[11] wl[143] vdd gnd cell_6t
Xbit_r144_c11 bl[11] br[11] wl[144] vdd gnd cell_6t
Xbit_r145_c11 bl[11] br[11] wl[145] vdd gnd cell_6t
Xbit_r146_c11 bl[11] br[11] wl[146] vdd gnd cell_6t
Xbit_r147_c11 bl[11] br[11] wl[147] vdd gnd cell_6t
Xbit_r148_c11 bl[11] br[11] wl[148] vdd gnd cell_6t
Xbit_r149_c11 bl[11] br[11] wl[149] vdd gnd cell_6t
Xbit_r150_c11 bl[11] br[11] wl[150] vdd gnd cell_6t
Xbit_r151_c11 bl[11] br[11] wl[151] vdd gnd cell_6t
Xbit_r152_c11 bl[11] br[11] wl[152] vdd gnd cell_6t
Xbit_r153_c11 bl[11] br[11] wl[153] vdd gnd cell_6t
Xbit_r154_c11 bl[11] br[11] wl[154] vdd gnd cell_6t
Xbit_r155_c11 bl[11] br[11] wl[155] vdd gnd cell_6t
Xbit_r156_c11 bl[11] br[11] wl[156] vdd gnd cell_6t
Xbit_r157_c11 bl[11] br[11] wl[157] vdd gnd cell_6t
Xbit_r158_c11 bl[11] br[11] wl[158] vdd gnd cell_6t
Xbit_r159_c11 bl[11] br[11] wl[159] vdd gnd cell_6t
Xbit_r160_c11 bl[11] br[11] wl[160] vdd gnd cell_6t
Xbit_r161_c11 bl[11] br[11] wl[161] vdd gnd cell_6t
Xbit_r162_c11 bl[11] br[11] wl[162] vdd gnd cell_6t
Xbit_r163_c11 bl[11] br[11] wl[163] vdd gnd cell_6t
Xbit_r164_c11 bl[11] br[11] wl[164] vdd gnd cell_6t
Xbit_r165_c11 bl[11] br[11] wl[165] vdd gnd cell_6t
Xbit_r166_c11 bl[11] br[11] wl[166] vdd gnd cell_6t
Xbit_r167_c11 bl[11] br[11] wl[167] vdd gnd cell_6t
Xbit_r168_c11 bl[11] br[11] wl[168] vdd gnd cell_6t
Xbit_r169_c11 bl[11] br[11] wl[169] vdd gnd cell_6t
Xbit_r170_c11 bl[11] br[11] wl[170] vdd gnd cell_6t
Xbit_r171_c11 bl[11] br[11] wl[171] vdd gnd cell_6t
Xbit_r172_c11 bl[11] br[11] wl[172] vdd gnd cell_6t
Xbit_r173_c11 bl[11] br[11] wl[173] vdd gnd cell_6t
Xbit_r174_c11 bl[11] br[11] wl[174] vdd gnd cell_6t
Xbit_r175_c11 bl[11] br[11] wl[175] vdd gnd cell_6t
Xbit_r176_c11 bl[11] br[11] wl[176] vdd gnd cell_6t
Xbit_r177_c11 bl[11] br[11] wl[177] vdd gnd cell_6t
Xbit_r178_c11 bl[11] br[11] wl[178] vdd gnd cell_6t
Xbit_r179_c11 bl[11] br[11] wl[179] vdd gnd cell_6t
Xbit_r180_c11 bl[11] br[11] wl[180] vdd gnd cell_6t
Xbit_r181_c11 bl[11] br[11] wl[181] vdd gnd cell_6t
Xbit_r182_c11 bl[11] br[11] wl[182] vdd gnd cell_6t
Xbit_r183_c11 bl[11] br[11] wl[183] vdd gnd cell_6t
Xbit_r184_c11 bl[11] br[11] wl[184] vdd gnd cell_6t
Xbit_r185_c11 bl[11] br[11] wl[185] vdd gnd cell_6t
Xbit_r186_c11 bl[11] br[11] wl[186] vdd gnd cell_6t
Xbit_r187_c11 bl[11] br[11] wl[187] vdd gnd cell_6t
Xbit_r188_c11 bl[11] br[11] wl[188] vdd gnd cell_6t
Xbit_r189_c11 bl[11] br[11] wl[189] vdd gnd cell_6t
Xbit_r190_c11 bl[11] br[11] wl[190] vdd gnd cell_6t
Xbit_r191_c11 bl[11] br[11] wl[191] vdd gnd cell_6t
Xbit_r192_c11 bl[11] br[11] wl[192] vdd gnd cell_6t
Xbit_r193_c11 bl[11] br[11] wl[193] vdd gnd cell_6t
Xbit_r194_c11 bl[11] br[11] wl[194] vdd gnd cell_6t
Xbit_r195_c11 bl[11] br[11] wl[195] vdd gnd cell_6t
Xbit_r196_c11 bl[11] br[11] wl[196] vdd gnd cell_6t
Xbit_r197_c11 bl[11] br[11] wl[197] vdd gnd cell_6t
Xbit_r198_c11 bl[11] br[11] wl[198] vdd gnd cell_6t
Xbit_r199_c11 bl[11] br[11] wl[199] vdd gnd cell_6t
Xbit_r200_c11 bl[11] br[11] wl[200] vdd gnd cell_6t
Xbit_r201_c11 bl[11] br[11] wl[201] vdd gnd cell_6t
Xbit_r202_c11 bl[11] br[11] wl[202] vdd gnd cell_6t
Xbit_r203_c11 bl[11] br[11] wl[203] vdd gnd cell_6t
Xbit_r204_c11 bl[11] br[11] wl[204] vdd gnd cell_6t
Xbit_r205_c11 bl[11] br[11] wl[205] vdd gnd cell_6t
Xbit_r206_c11 bl[11] br[11] wl[206] vdd gnd cell_6t
Xbit_r207_c11 bl[11] br[11] wl[207] vdd gnd cell_6t
Xbit_r208_c11 bl[11] br[11] wl[208] vdd gnd cell_6t
Xbit_r209_c11 bl[11] br[11] wl[209] vdd gnd cell_6t
Xbit_r210_c11 bl[11] br[11] wl[210] vdd gnd cell_6t
Xbit_r211_c11 bl[11] br[11] wl[211] vdd gnd cell_6t
Xbit_r212_c11 bl[11] br[11] wl[212] vdd gnd cell_6t
Xbit_r213_c11 bl[11] br[11] wl[213] vdd gnd cell_6t
Xbit_r214_c11 bl[11] br[11] wl[214] vdd gnd cell_6t
Xbit_r215_c11 bl[11] br[11] wl[215] vdd gnd cell_6t
Xbit_r216_c11 bl[11] br[11] wl[216] vdd gnd cell_6t
Xbit_r217_c11 bl[11] br[11] wl[217] vdd gnd cell_6t
Xbit_r218_c11 bl[11] br[11] wl[218] vdd gnd cell_6t
Xbit_r219_c11 bl[11] br[11] wl[219] vdd gnd cell_6t
Xbit_r220_c11 bl[11] br[11] wl[220] vdd gnd cell_6t
Xbit_r221_c11 bl[11] br[11] wl[221] vdd gnd cell_6t
Xbit_r222_c11 bl[11] br[11] wl[222] vdd gnd cell_6t
Xbit_r223_c11 bl[11] br[11] wl[223] vdd gnd cell_6t
Xbit_r224_c11 bl[11] br[11] wl[224] vdd gnd cell_6t
Xbit_r225_c11 bl[11] br[11] wl[225] vdd gnd cell_6t
Xbit_r226_c11 bl[11] br[11] wl[226] vdd gnd cell_6t
Xbit_r227_c11 bl[11] br[11] wl[227] vdd gnd cell_6t
Xbit_r228_c11 bl[11] br[11] wl[228] vdd gnd cell_6t
Xbit_r229_c11 bl[11] br[11] wl[229] vdd gnd cell_6t
Xbit_r230_c11 bl[11] br[11] wl[230] vdd gnd cell_6t
Xbit_r231_c11 bl[11] br[11] wl[231] vdd gnd cell_6t
Xbit_r232_c11 bl[11] br[11] wl[232] vdd gnd cell_6t
Xbit_r233_c11 bl[11] br[11] wl[233] vdd gnd cell_6t
Xbit_r234_c11 bl[11] br[11] wl[234] vdd gnd cell_6t
Xbit_r235_c11 bl[11] br[11] wl[235] vdd gnd cell_6t
Xbit_r236_c11 bl[11] br[11] wl[236] vdd gnd cell_6t
Xbit_r237_c11 bl[11] br[11] wl[237] vdd gnd cell_6t
Xbit_r238_c11 bl[11] br[11] wl[238] vdd gnd cell_6t
Xbit_r239_c11 bl[11] br[11] wl[239] vdd gnd cell_6t
Xbit_r240_c11 bl[11] br[11] wl[240] vdd gnd cell_6t
Xbit_r241_c11 bl[11] br[11] wl[241] vdd gnd cell_6t
Xbit_r242_c11 bl[11] br[11] wl[242] vdd gnd cell_6t
Xbit_r243_c11 bl[11] br[11] wl[243] vdd gnd cell_6t
Xbit_r244_c11 bl[11] br[11] wl[244] vdd gnd cell_6t
Xbit_r245_c11 bl[11] br[11] wl[245] vdd gnd cell_6t
Xbit_r246_c11 bl[11] br[11] wl[246] vdd gnd cell_6t
Xbit_r247_c11 bl[11] br[11] wl[247] vdd gnd cell_6t
Xbit_r248_c11 bl[11] br[11] wl[248] vdd gnd cell_6t
Xbit_r249_c11 bl[11] br[11] wl[249] vdd gnd cell_6t
Xbit_r250_c11 bl[11] br[11] wl[250] vdd gnd cell_6t
Xbit_r251_c11 bl[11] br[11] wl[251] vdd gnd cell_6t
Xbit_r252_c11 bl[11] br[11] wl[252] vdd gnd cell_6t
Xbit_r253_c11 bl[11] br[11] wl[253] vdd gnd cell_6t
Xbit_r254_c11 bl[11] br[11] wl[254] vdd gnd cell_6t
Xbit_r255_c11 bl[11] br[11] wl[255] vdd gnd cell_6t
Xbit_r0_c12 bl[12] br[12] wl[0] vdd gnd cell_6t
Xbit_r1_c12 bl[12] br[12] wl[1] vdd gnd cell_6t
Xbit_r2_c12 bl[12] br[12] wl[2] vdd gnd cell_6t
Xbit_r3_c12 bl[12] br[12] wl[3] vdd gnd cell_6t
Xbit_r4_c12 bl[12] br[12] wl[4] vdd gnd cell_6t
Xbit_r5_c12 bl[12] br[12] wl[5] vdd gnd cell_6t
Xbit_r6_c12 bl[12] br[12] wl[6] vdd gnd cell_6t
Xbit_r7_c12 bl[12] br[12] wl[7] vdd gnd cell_6t
Xbit_r8_c12 bl[12] br[12] wl[8] vdd gnd cell_6t
Xbit_r9_c12 bl[12] br[12] wl[9] vdd gnd cell_6t
Xbit_r10_c12 bl[12] br[12] wl[10] vdd gnd cell_6t
Xbit_r11_c12 bl[12] br[12] wl[11] vdd gnd cell_6t
Xbit_r12_c12 bl[12] br[12] wl[12] vdd gnd cell_6t
Xbit_r13_c12 bl[12] br[12] wl[13] vdd gnd cell_6t
Xbit_r14_c12 bl[12] br[12] wl[14] vdd gnd cell_6t
Xbit_r15_c12 bl[12] br[12] wl[15] vdd gnd cell_6t
Xbit_r16_c12 bl[12] br[12] wl[16] vdd gnd cell_6t
Xbit_r17_c12 bl[12] br[12] wl[17] vdd gnd cell_6t
Xbit_r18_c12 bl[12] br[12] wl[18] vdd gnd cell_6t
Xbit_r19_c12 bl[12] br[12] wl[19] vdd gnd cell_6t
Xbit_r20_c12 bl[12] br[12] wl[20] vdd gnd cell_6t
Xbit_r21_c12 bl[12] br[12] wl[21] vdd gnd cell_6t
Xbit_r22_c12 bl[12] br[12] wl[22] vdd gnd cell_6t
Xbit_r23_c12 bl[12] br[12] wl[23] vdd gnd cell_6t
Xbit_r24_c12 bl[12] br[12] wl[24] vdd gnd cell_6t
Xbit_r25_c12 bl[12] br[12] wl[25] vdd gnd cell_6t
Xbit_r26_c12 bl[12] br[12] wl[26] vdd gnd cell_6t
Xbit_r27_c12 bl[12] br[12] wl[27] vdd gnd cell_6t
Xbit_r28_c12 bl[12] br[12] wl[28] vdd gnd cell_6t
Xbit_r29_c12 bl[12] br[12] wl[29] vdd gnd cell_6t
Xbit_r30_c12 bl[12] br[12] wl[30] vdd gnd cell_6t
Xbit_r31_c12 bl[12] br[12] wl[31] vdd gnd cell_6t
Xbit_r32_c12 bl[12] br[12] wl[32] vdd gnd cell_6t
Xbit_r33_c12 bl[12] br[12] wl[33] vdd gnd cell_6t
Xbit_r34_c12 bl[12] br[12] wl[34] vdd gnd cell_6t
Xbit_r35_c12 bl[12] br[12] wl[35] vdd gnd cell_6t
Xbit_r36_c12 bl[12] br[12] wl[36] vdd gnd cell_6t
Xbit_r37_c12 bl[12] br[12] wl[37] vdd gnd cell_6t
Xbit_r38_c12 bl[12] br[12] wl[38] vdd gnd cell_6t
Xbit_r39_c12 bl[12] br[12] wl[39] vdd gnd cell_6t
Xbit_r40_c12 bl[12] br[12] wl[40] vdd gnd cell_6t
Xbit_r41_c12 bl[12] br[12] wl[41] vdd gnd cell_6t
Xbit_r42_c12 bl[12] br[12] wl[42] vdd gnd cell_6t
Xbit_r43_c12 bl[12] br[12] wl[43] vdd gnd cell_6t
Xbit_r44_c12 bl[12] br[12] wl[44] vdd gnd cell_6t
Xbit_r45_c12 bl[12] br[12] wl[45] vdd gnd cell_6t
Xbit_r46_c12 bl[12] br[12] wl[46] vdd gnd cell_6t
Xbit_r47_c12 bl[12] br[12] wl[47] vdd gnd cell_6t
Xbit_r48_c12 bl[12] br[12] wl[48] vdd gnd cell_6t
Xbit_r49_c12 bl[12] br[12] wl[49] vdd gnd cell_6t
Xbit_r50_c12 bl[12] br[12] wl[50] vdd gnd cell_6t
Xbit_r51_c12 bl[12] br[12] wl[51] vdd gnd cell_6t
Xbit_r52_c12 bl[12] br[12] wl[52] vdd gnd cell_6t
Xbit_r53_c12 bl[12] br[12] wl[53] vdd gnd cell_6t
Xbit_r54_c12 bl[12] br[12] wl[54] vdd gnd cell_6t
Xbit_r55_c12 bl[12] br[12] wl[55] vdd gnd cell_6t
Xbit_r56_c12 bl[12] br[12] wl[56] vdd gnd cell_6t
Xbit_r57_c12 bl[12] br[12] wl[57] vdd gnd cell_6t
Xbit_r58_c12 bl[12] br[12] wl[58] vdd gnd cell_6t
Xbit_r59_c12 bl[12] br[12] wl[59] vdd gnd cell_6t
Xbit_r60_c12 bl[12] br[12] wl[60] vdd gnd cell_6t
Xbit_r61_c12 bl[12] br[12] wl[61] vdd gnd cell_6t
Xbit_r62_c12 bl[12] br[12] wl[62] vdd gnd cell_6t
Xbit_r63_c12 bl[12] br[12] wl[63] vdd gnd cell_6t
Xbit_r64_c12 bl[12] br[12] wl[64] vdd gnd cell_6t
Xbit_r65_c12 bl[12] br[12] wl[65] vdd gnd cell_6t
Xbit_r66_c12 bl[12] br[12] wl[66] vdd gnd cell_6t
Xbit_r67_c12 bl[12] br[12] wl[67] vdd gnd cell_6t
Xbit_r68_c12 bl[12] br[12] wl[68] vdd gnd cell_6t
Xbit_r69_c12 bl[12] br[12] wl[69] vdd gnd cell_6t
Xbit_r70_c12 bl[12] br[12] wl[70] vdd gnd cell_6t
Xbit_r71_c12 bl[12] br[12] wl[71] vdd gnd cell_6t
Xbit_r72_c12 bl[12] br[12] wl[72] vdd gnd cell_6t
Xbit_r73_c12 bl[12] br[12] wl[73] vdd gnd cell_6t
Xbit_r74_c12 bl[12] br[12] wl[74] vdd gnd cell_6t
Xbit_r75_c12 bl[12] br[12] wl[75] vdd gnd cell_6t
Xbit_r76_c12 bl[12] br[12] wl[76] vdd gnd cell_6t
Xbit_r77_c12 bl[12] br[12] wl[77] vdd gnd cell_6t
Xbit_r78_c12 bl[12] br[12] wl[78] vdd gnd cell_6t
Xbit_r79_c12 bl[12] br[12] wl[79] vdd gnd cell_6t
Xbit_r80_c12 bl[12] br[12] wl[80] vdd gnd cell_6t
Xbit_r81_c12 bl[12] br[12] wl[81] vdd gnd cell_6t
Xbit_r82_c12 bl[12] br[12] wl[82] vdd gnd cell_6t
Xbit_r83_c12 bl[12] br[12] wl[83] vdd gnd cell_6t
Xbit_r84_c12 bl[12] br[12] wl[84] vdd gnd cell_6t
Xbit_r85_c12 bl[12] br[12] wl[85] vdd gnd cell_6t
Xbit_r86_c12 bl[12] br[12] wl[86] vdd gnd cell_6t
Xbit_r87_c12 bl[12] br[12] wl[87] vdd gnd cell_6t
Xbit_r88_c12 bl[12] br[12] wl[88] vdd gnd cell_6t
Xbit_r89_c12 bl[12] br[12] wl[89] vdd gnd cell_6t
Xbit_r90_c12 bl[12] br[12] wl[90] vdd gnd cell_6t
Xbit_r91_c12 bl[12] br[12] wl[91] vdd gnd cell_6t
Xbit_r92_c12 bl[12] br[12] wl[92] vdd gnd cell_6t
Xbit_r93_c12 bl[12] br[12] wl[93] vdd gnd cell_6t
Xbit_r94_c12 bl[12] br[12] wl[94] vdd gnd cell_6t
Xbit_r95_c12 bl[12] br[12] wl[95] vdd gnd cell_6t
Xbit_r96_c12 bl[12] br[12] wl[96] vdd gnd cell_6t
Xbit_r97_c12 bl[12] br[12] wl[97] vdd gnd cell_6t
Xbit_r98_c12 bl[12] br[12] wl[98] vdd gnd cell_6t
Xbit_r99_c12 bl[12] br[12] wl[99] vdd gnd cell_6t
Xbit_r100_c12 bl[12] br[12] wl[100] vdd gnd cell_6t
Xbit_r101_c12 bl[12] br[12] wl[101] vdd gnd cell_6t
Xbit_r102_c12 bl[12] br[12] wl[102] vdd gnd cell_6t
Xbit_r103_c12 bl[12] br[12] wl[103] vdd gnd cell_6t
Xbit_r104_c12 bl[12] br[12] wl[104] vdd gnd cell_6t
Xbit_r105_c12 bl[12] br[12] wl[105] vdd gnd cell_6t
Xbit_r106_c12 bl[12] br[12] wl[106] vdd gnd cell_6t
Xbit_r107_c12 bl[12] br[12] wl[107] vdd gnd cell_6t
Xbit_r108_c12 bl[12] br[12] wl[108] vdd gnd cell_6t
Xbit_r109_c12 bl[12] br[12] wl[109] vdd gnd cell_6t
Xbit_r110_c12 bl[12] br[12] wl[110] vdd gnd cell_6t
Xbit_r111_c12 bl[12] br[12] wl[111] vdd gnd cell_6t
Xbit_r112_c12 bl[12] br[12] wl[112] vdd gnd cell_6t
Xbit_r113_c12 bl[12] br[12] wl[113] vdd gnd cell_6t
Xbit_r114_c12 bl[12] br[12] wl[114] vdd gnd cell_6t
Xbit_r115_c12 bl[12] br[12] wl[115] vdd gnd cell_6t
Xbit_r116_c12 bl[12] br[12] wl[116] vdd gnd cell_6t
Xbit_r117_c12 bl[12] br[12] wl[117] vdd gnd cell_6t
Xbit_r118_c12 bl[12] br[12] wl[118] vdd gnd cell_6t
Xbit_r119_c12 bl[12] br[12] wl[119] vdd gnd cell_6t
Xbit_r120_c12 bl[12] br[12] wl[120] vdd gnd cell_6t
Xbit_r121_c12 bl[12] br[12] wl[121] vdd gnd cell_6t
Xbit_r122_c12 bl[12] br[12] wl[122] vdd gnd cell_6t
Xbit_r123_c12 bl[12] br[12] wl[123] vdd gnd cell_6t
Xbit_r124_c12 bl[12] br[12] wl[124] vdd gnd cell_6t
Xbit_r125_c12 bl[12] br[12] wl[125] vdd gnd cell_6t
Xbit_r126_c12 bl[12] br[12] wl[126] vdd gnd cell_6t
Xbit_r127_c12 bl[12] br[12] wl[127] vdd gnd cell_6t
Xbit_r128_c12 bl[12] br[12] wl[128] vdd gnd cell_6t
Xbit_r129_c12 bl[12] br[12] wl[129] vdd gnd cell_6t
Xbit_r130_c12 bl[12] br[12] wl[130] vdd gnd cell_6t
Xbit_r131_c12 bl[12] br[12] wl[131] vdd gnd cell_6t
Xbit_r132_c12 bl[12] br[12] wl[132] vdd gnd cell_6t
Xbit_r133_c12 bl[12] br[12] wl[133] vdd gnd cell_6t
Xbit_r134_c12 bl[12] br[12] wl[134] vdd gnd cell_6t
Xbit_r135_c12 bl[12] br[12] wl[135] vdd gnd cell_6t
Xbit_r136_c12 bl[12] br[12] wl[136] vdd gnd cell_6t
Xbit_r137_c12 bl[12] br[12] wl[137] vdd gnd cell_6t
Xbit_r138_c12 bl[12] br[12] wl[138] vdd gnd cell_6t
Xbit_r139_c12 bl[12] br[12] wl[139] vdd gnd cell_6t
Xbit_r140_c12 bl[12] br[12] wl[140] vdd gnd cell_6t
Xbit_r141_c12 bl[12] br[12] wl[141] vdd gnd cell_6t
Xbit_r142_c12 bl[12] br[12] wl[142] vdd gnd cell_6t
Xbit_r143_c12 bl[12] br[12] wl[143] vdd gnd cell_6t
Xbit_r144_c12 bl[12] br[12] wl[144] vdd gnd cell_6t
Xbit_r145_c12 bl[12] br[12] wl[145] vdd gnd cell_6t
Xbit_r146_c12 bl[12] br[12] wl[146] vdd gnd cell_6t
Xbit_r147_c12 bl[12] br[12] wl[147] vdd gnd cell_6t
Xbit_r148_c12 bl[12] br[12] wl[148] vdd gnd cell_6t
Xbit_r149_c12 bl[12] br[12] wl[149] vdd gnd cell_6t
Xbit_r150_c12 bl[12] br[12] wl[150] vdd gnd cell_6t
Xbit_r151_c12 bl[12] br[12] wl[151] vdd gnd cell_6t
Xbit_r152_c12 bl[12] br[12] wl[152] vdd gnd cell_6t
Xbit_r153_c12 bl[12] br[12] wl[153] vdd gnd cell_6t
Xbit_r154_c12 bl[12] br[12] wl[154] vdd gnd cell_6t
Xbit_r155_c12 bl[12] br[12] wl[155] vdd gnd cell_6t
Xbit_r156_c12 bl[12] br[12] wl[156] vdd gnd cell_6t
Xbit_r157_c12 bl[12] br[12] wl[157] vdd gnd cell_6t
Xbit_r158_c12 bl[12] br[12] wl[158] vdd gnd cell_6t
Xbit_r159_c12 bl[12] br[12] wl[159] vdd gnd cell_6t
Xbit_r160_c12 bl[12] br[12] wl[160] vdd gnd cell_6t
Xbit_r161_c12 bl[12] br[12] wl[161] vdd gnd cell_6t
Xbit_r162_c12 bl[12] br[12] wl[162] vdd gnd cell_6t
Xbit_r163_c12 bl[12] br[12] wl[163] vdd gnd cell_6t
Xbit_r164_c12 bl[12] br[12] wl[164] vdd gnd cell_6t
Xbit_r165_c12 bl[12] br[12] wl[165] vdd gnd cell_6t
Xbit_r166_c12 bl[12] br[12] wl[166] vdd gnd cell_6t
Xbit_r167_c12 bl[12] br[12] wl[167] vdd gnd cell_6t
Xbit_r168_c12 bl[12] br[12] wl[168] vdd gnd cell_6t
Xbit_r169_c12 bl[12] br[12] wl[169] vdd gnd cell_6t
Xbit_r170_c12 bl[12] br[12] wl[170] vdd gnd cell_6t
Xbit_r171_c12 bl[12] br[12] wl[171] vdd gnd cell_6t
Xbit_r172_c12 bl[12] br[12] wl[172] vdd gnd cell_6t
Xbit_r173_c12 bl[12] br[12] wl[173] vdd gnd cell_6t
Xbit_r174_c12 bl[12] br[12] wl[174] vdd gnd cell_6t
Xbit_r175_c12 bl[12] br[12] wl[175] vdd gnd cell_6t
Xbit_r176_c12 bl[12] br[12] wl[176] vdd gnd cell_6t
Xbit_r177_c12 bl[12] br[12] wl[177] vdd gnd cell_6t
Xbit_r178_c12 bl[12] br[12] wl[178] vdd gnd cell_6t
Xbit_r179_c12 bl[12] br[12] wl[179] vdd gnd cell_6t
Xbit_r180_c12 bl[12] br[12] wl[180] vdd gnd cell_6t
Xbit_r181_c12 bl[12] br[12] wl[181] vdd gnd cell_6t
Xbit_r182_c12 bl[12] br[12] wl[182] vdd gnd cell_6t
Xbit_r183_c12 bl[12] br[12] wl[183] vdd gnd cell_6t
Xbit_r184_c12 bl[12] br[12] wl[184] vdd gnd cell_6t
Xbit_r185_c12 bl[12] br[12] wl[185] vdd gnd cell_6t
Xbit_r186_c12 bl[12] br[12] wl[186] vdd gnd cell_6t
Xbit_r187_c12 bl[12] br[12] wl[187] vdd gnd cell_6t
Xbit_r188_c12 bl[12] br[12] wl[188] vdd gnd cell_6t
Xbit_r189_c12 bl[12] br[12] wl[189] vdd gnd cell_6t
Xbit_r190_c12 bl[12] br[12] wl[190] vdd gnd cell_6t
Xbit_r191_c12 bl[12] br[12] wl[191] vdd gnd cell_6t
Xbit_r192_c12 bl[12] br[12] wl[192] vdd gnd cell_6t
Xbit_r193_c12 bl[12] br[12] wl[193] vdd gnd cell_6t
Xbit_r194_c12 bl[12] br[12] wl[194] vdd gnd cell_6t
Xbit_r195_c12 bl[12] br[12] wl[195] vdd gnd cell_6t
Xbit_r196_c12 bl[12] br[12] wl[196] vdd gnd cell_6t
Xbit_r197_c12 bl[12] br[12] wl[197] vdd gnd cell_6t
Xbit_r198_c12 bl[12] br[12] wl[198] vdd gnd cell_6t
Xbit_r199_c12 bl[12] br[12] wl[199] vdd gnd cell_6t
Xbit_r200_c12 bl[12] br[12] wl[200] vdd gnd cell_6t
Xbit_r201_c12 bl[12] br[12] wl[201] vdd gnd cell_6t
Xbit_r202_c12 bl[12] br[12] wl[202] vdd gnd cell_6t
Xbit_r203_c12 bl[12] br[12] wl[203] vdd gnd cell_6t
Xbit_r204_c12 bl[12] br[12] wl[204] vdd gnd cell_6t
Xbit_r205_c12 bl[12] br[12] wl[205] vdd gnd cell_6t
Xbit_r206_c12 bl[12] br[12] wl[206] vdd gnd cell_6t
Xbit_r207_c12 bl[12] br[12] wl[207] vdd gnd cell_6t
Xbit_r208_c12 bl[12] br[12] wl[208] vdd gnd cell_6t
Xbit_r209_c12 bl[12] br[12] wl[209] vdd gnd cell_6t
Xbit_r210_c12 bl[12] br[12] wl[210] vdd gnd cell_6t
Xbit_r211_c12 bl[12] br[12] wl[211] vdd gnd cell_6t
Xbit_r212_c12 bl[12] br[12] wl[212] vdd gnd cell_6t
Xbit_r213_c12 bl[12] br[12] wl[213] vdd gnd cell_6t
Xbit_r214_c12 bl[12] br[12] wl[214] vdd gnd cell_6t
Xbit_r215_c12 bl[12] br[12] wl[215] vdd gnd cell_6t
Xbit_r216_c12 bl[12] br[12] wl[216] vdd gnd cell_6t
Xbit_r217_c12 bl[12] br[12] wl[217] vdd gnd cell_6t
Xbit_r218_c12 bl[12] br[12] wl[218] vdd gnd cell_6t
Xbit_r219_c12 bl[12] br[12] wl[219] vdd gnd cell_6t
Xbit_r220_c12 bl[12] br[12] wl[220] vdd gnd cell_6t
Xbit_r221_c12 bl[12] br[12] wl[221] vdd gnd cell_6t
Xbit_r222_c12 bl[12] br[12] wl[222] vdd gnd cell_6t
Xbit_r223_c12 bl[12] br[12] wl[223] vdd gnd cell_6t
Xbit_r224_c12 bl[12] br[12] wl[224] vdd gnd cell_6t
Xbit_r225_c12 bl[12] br[12] wl[225] vdd gnd cell_6t
Xbit_r226_c12 bl[12] br[12] wl[226] vdd gnd cell_6t
Xbit_r227_c12 bl[12] br[12] wl[227] vdd gnd cell_6t
Xbit_r228_c12 bl[12] br[12] wl[228] vdd gnd cell_6t
Xbit_r229_c12 bl[12] br[12] wl[229] vdd gnd cell_6t
Xbit_r230_c12 bl[12] br[12] wl[230] vdd gnd cell_6t
Xbit_r231_c12 bl[12] br[12] wl[231] vdd gnd cell_6t
Xbit_r232_c12 bl[12] br[12] wl[232] vdd gnd cell_6t
Xbit_r233_c12 bl[12] br[12] wl[233] vdd gnd cell_6t
Xbit_r234_c12 bl[12] br[12] wl[234] vdd gnd cell_6t
Xbit_r235_c12 bl[12] br[12] wl[235] vdd gnd cell_6t
Xbit_r236_c12 bl[12] br[12] wl[236] vdd gnd cell_6t
Xbit_r237_c12 bl[12] br[12] wl[237] vdd gnd cell_6t
Xbit_r238_c12 bl[12] br[12] wl[238] vdd gnd cell_6t
Xbit_r239_c12 bl[12] br[12] wl[239] vdd gnd cell_6t
Xbit_r240_c12 bl[12] br[12] wl[240] vdd gnd cell_6t
Xbit_r241_c12 bl[12] br[12] wl[241] vdd gnd cell_6t
Xbit_r242_c12 bl[12] br[12] wl[242] vdd gnd cell_6t
Xbit_r243_c12 bl[12] br[12] wl[243] vdd gnd cell_6t
Xbit_r244_c12 bl[12] br[12] wl[244] vdd gnd cell_6t
Xbit_r245_c12 bl[12] br[12] wl[245] vdd gnd cell_6t
Xbit_r246_c12 bl[12] br[12] wl[246] vdd gnd cell_6t
Xbit_r247_c12 bl[12] br[12] wl[247] vdd gnd cell_6t
Xbit_r248_c12 bl[12] br[12] wl[248] vdd gnd cell_6t
Xbit_r249_c12 bl[12] br[12] wl[249] vdd gnd cell_6t
Xbit_r250_c12 bl[12] br[12] wl[250] vdd gnd cell_6t
Xbit_r251_c12 bl[12] br[12] wl[251] vdd gnd cell_6t
Xbit_r252_c12 bl[12] br[12] wl[252] vdd gnd cell_6t
Xbit_r253_c12 bl[12] br[12] wl[253] vdd gnd cell_6t
Xbit_r254_c12 bl[12] br[12] wl[254] vdd gnd cell_6t
Xbit_r255_c12 bl[12] br[12] wl[255] vdd gnd cell_6t
Xbit_r0_c13 bl[13] br[13] wl[0] vdd gnd cell_6t
Xbit_r1_c13 bl[13] br[13] wl[1] vdd gnd cell_6t
Xbit_r2_c13 bl[13] br[13] wl[2] vdd gnd cell_6t
Xbit_r3_c13 bl[13] br[13] wl[3] vdd gnd cell_6t
Xbit_r4_c13 bl[13] br[13] wl[4] vdd gnd cell_6t
Xbit_r5_c13 bl[13] br[13] wl[5] vdd gnd cell_6t
Xbit_r6_c13 bl[13] br[13] wl[6] vdd gnd cell_6t
Xbit_r7_c13 bl[13] br[13] wl[7] vdd gnd cell_6t
Xbit_r8_c13 bl[13] br[13] wl[8] vdd gnd cell_6t
Xbit_r9_c13 bl[13] br[13] wl[9] vdd gnd cell_6t
Xbit_r10_c13 bl[13] br[13] wl[10] vdd gnd cell_6t
Xbit_r11_c13 bl[13] br[13] wl[11] vdd gnd cell_6t
Xbit_r12_c13 bl[13] br[13] wl[12] vdd gnd cell_6t
Xbit_r13_c13 bl[13] br[13] wl[13] vdd gnd cell_6t
Xbit_r14_c13 bl[13] br[13] wl[14] vdd gnd cell_6t
Xbit_r15_c13 bl[13] br[13] wl[15] vdd gnd cell_6t
Xbit_r16_c13 bl[13] br[13] wl[16] vdd gnd cell_6t
Xbit_r17_c13 bl[13] br[13] wl[17] vdd gnd cell_6t
Xbit_r18_c13 bl[13] br[13] wl[18] vdd gnd cell_6t
Xbit_r19_c13 bl[13] br[13] wl[19] vdd gnd cell_6t
Xbit_r20_c13 bl[13] br[13] wl[20] vdd gnd cell_6t
Xbit_r21_c13 bl[13] br[13] wl[21] vdd gnd cell_6t
Xbit_r22_c13 bl[13] br[13] wl[22] vdd gnd cell_6t
Xbit_r23_c13 bl[13] br[13] wl[23] vdd gnd cell_6t
Xbit_r24_c13 bl[13] br[13] wl[24] vdd gnd cell_6t
Xbit_r25_c13 bl[13] br[13] wl[25] vdd gnd cell_6t
Xbit_r26_c13 bl[13] br[13] wl[26] vdd gnd cell_6t
Xbit_r27_c13 bl[13] br[13] wl[27] vdd gnd cell_6t
Xbit_r28_c13 bl[13] br[13] wl[28] vdd gnd cell_6t
Xbit_r29_c13 bl[13] br[13] wl[29] vdd gnd cell_6t
Xbit_r30_c13 bl[13] br[13] wl[30] vdd gnd cell_6t
Xbit_r31_c13 bl[13] br[13] wl[31] vdd gnd cell_6t
Xbit_r32_c13 bl[13] br[13] wl[32] vdd gnd cell_6t
Xbit_r33_c13 bl[13] br[13] wl[33] vdd gnd cell_6t
Xbit_r34_c13 bl[13] br[13] wl[34] vdd gnd cell_6t
Xbit_r35_c13 bl[13] br[13] wl[35] vdd gnd cell_6t
Xbit_r36_c13 bl[13] br[13] wl[36] vdd gnd cell_6t
Xbit_r37_c13 bl[13] br[13] wl[37] vdd gnd cell_6t
Xbit_r38_c13 bl[13] br[13] wl[38] vdd gnd cell_6t
Xbit_r39_c13 bl[13] br[13] wl[39] vdd gnd cell_6t
Xbit_r40_c13 bl[13] br[13] wl[40] vdd gnd cell_6t
Xbit_r41_c13 bl[13] br[13] wl[41] vdd gnd cell_6t
Xbit_r42_c13 bl[13] br[13] wl[42] vdd gnd cell_6t
Xbit_r43_c13 bl[13] br[13] wl[43] vdd gnd cell_6t
Xbit_r44_c13 bl[13] br[13] wl[44] vdd gnd cell_6t
Xbit_r45_c13 bl[13] br[13] wl[45] vdd gnd cell_6t
Xbit_r46_c13 bl[13] br[13] wl[46] vdd gnd cell_6t
Xbit_r47_c13 bl[13] br[13] wl[47] vdd gnd cell_6t
Xbit_r48_c13 bl[13] br[13] wl[48] vdd gnd cell_6t
Xbit_r49_c13 bl[13] br[13] wl[49] vdd gnd cell_6t
Xbit_r50_c13 bl[13] br[13] wl[50] vdd gnd cell_6t
Xbit_r51_c13 bl[13] br[13] wl[51] vdd gnd cell_6t
Xbit_r52_c13 bl[13] br[13] wl[52] vdd gnd cell_6t
Xbit_r53_c13 bl[13] br[13] wl[53] vdd gnd cell_6t
Xbit_r54_c13 bl[13] br[13] wl[54] vdd gnd cell_6t
Xbit_r55_c13 bl[13] br[13] wl[55] vdd gnd cell_6t
Xbit_r56_c13 bl[13] br[13] wl[56] vdd gnd cell_6t
Xbit_r57_c13 bl[13] br[13] wl[57] vdd gnd cell_6t
Xbit_r58_c13 bl[13] br[13] wl[58] vdd gnd cell_6t
Xbit_r59_c13 bl[13] br[13] wl[59] vdd gnd cell_6t
Xbit_r60_c13 bl[13] br[13] wl[60] vdd gnd cell_6t
Xbit_r61_c13 bl[13] br[13] wl[61] vdd gnd cell_6t
Xbit_r62_c13 bl[13] br[13] wl[62] vdd gnd cell_6t
Xbit_r63_c13 bl[13] br[13] wl[63] vdd gnd cell_6t
Xbit_r64_c13 bl[13] br[13] wl[64] vdd gnd cell_6t
Xbit_r65_c13 bl[13] br[13] wl[65] vdd gnd cell_6t
Xbit_r66_c13 bl[13] br[13] wl[66] vdd gnd cell_6t
Xbit_r67_c13 bl[13] br[13] wl[67] vdd gnd cell_6t
Xbit_r68_c13 bl[13] br[13] wl[68] vdd gnd cell_6t
Xbit_r69_c13 bl[13] br[13] wl[69] vdd gnd cell_6t
Xbit_r70_c13 bl[13] br[13] wl[70] vdd gnd cell_6t
Xbit_r71_c13 bl[13] br[13] wl[71] vdd gnd cell_6t
Xbit_r72_c13 bl[13] br[13] wl[72] vdd gnd cell_6t
Xbit_r73_c13 bl[13] br[13] wl[73] vdd gnd cell_6t
Xbit_r74_c13 bl[13] br[13] wl[74] vdd gnd cell_6t
Xbit_r75_c13 bl[13] br[13] wl[75] vdd gnd cell_6t
Xbit_r76_c13 bl[13] br[13] wl[76] vdd gnd cell_6t
Xbit_r77_c13 bl[13] br[13] wl[77] vdd gnd cell_6t
Xbit_r78_c13 bl[13] br[13] wl[78] vdd gnd cell_6t
Xbit_r79_c13 bl[13] br[13] wl[79] vdd gnd cell_6t
Xbit_r80_c13 bl[13] br[13] wl[80] vdd gnd cell_6t
Xbit_r81_c13 bl[13] br[13] wl[81] vdd gnd cell_6t
Xbit_r82_c13 bl[13] br[13] wl[82] vdd gnd cell_6t
Xbit_r83_c13 bl[13] br[13] wl[83] vdd gnd cell_6t
Xbit_r84_c13 bl[13] br[13] wl[84] vdd gnd cell_6t
Xbit_r85_c13 bl[13] br[13] wl[85] vdd gnd cell_6t
Xbit_r86_c13 bl[13] br[13] wl[86] vdd gnd cell_6t
Xbit_r87_c13 bl[13] br[13] wl[87] vdd gnd cell_6t
Xbit_r88_c13 bl[13] br[13] wl[88] vdd gnd cell_6t
Xbit_r89_c13 bl[13] br[13] wl[89] vdd gnd cell_6t
Xbit_r90_c13 bl[13] br[13] wl[90] vdd gnd cell_6t
Xbit_r91_c13 bl[13] br[13] wl[91] vdd gnd cell_6t
Xbit_r92_c13 bl[13] br[13] wl[92] vdd gnd cell_6t
Xbit_r93_c13 bl[13] br[13] wl[93] vdd gnd cell_6t
Xbit_r94_c13 bl[13] br[13] wl[94] vdd gnd cell_6t
Xbit_r95_c13 bl[13] br[13] wl[95] vdd gnd cell_6t
Xbit_r96_c13 bl[13] br[13] wl[96] vdd gnd cell_6t
Xbit_r97_c13 bl[13] br[13] wl[97] vdd gnd cell_6t
Xbit_r98_c13 bl[13] br[13] wl[98] vdd gnd cell_6t
Xbit_r99_c13 bl[13] br[13] wl[99] vdd gnd cell_6t
Xbit_r100_c13 bl[13] br[13] wl[100] vdd gnd cell_6t
Xbit_r101_c13 bl[13] br[13] wl[101] vdd gnd cell_6t
Xbit_r102_c13 bl[13] br[13] wl[102] vdd gnd cell_6t
Xbit_r103_c13 bl[13] br[13] wl[103] vdd gnd cell_6t
Xbit_r104_c13 bl[13] br[13] wl[104] vdd gnd cell_6t
Xbit_r105_c13 bl[13] br[13] wl[105] vdd gnd cell_6t
Xbit_r106_c13 bl[13] br[13] wl[106] vdd gnd cell_6t
Xbit_r107_c13 bl[13] br[13] wl[107] vdd gnd cell_6t
Xbit_r108_c13 bl[13] br[13] wl[108] vdd gnd cell_6t
Xbit_r109_c13 bl[13] br[13] wl[109] vdd gnd cell_6t
Xbit_r110_c13 bl[13] br[13] wl[110] vdd gnd cell_6t
Xbit_r111_c13 bl[13] br[13] wl[111] vdd gnd cell_6t
Xbit_r112_c13 bl[13] br[13] wl[112] vdd gnd cell_6t
Xbit_r113_c13 bl[13] br[13] wl[113] vdd gnd cell_6t
Xbit_r114_c13 bl[13] br[13] wl[114] vdd gnd cell_6t
Xbit_r115_c13 bl[13] br[13] wl[115] vdd gnd cell_6t
Xbit_r116_c13 bl[13] br[13] wl[116] vdd gnd cell_6t
Xbit_r117_c13 bl[13] br[13] wl[117] vdd gnd cell_6t
Xbit_r118_c13 bl[13] br[13] wl[118] vdd gnd cell_6t
Xbit_r119_c13 bl[13] br[13] wl[119] vdd gnd cell_6t
Xbit_r120_c13 bl[13] br[13] wl[120] vdd gnd cell_6t
Xbit_r121_c13 bl[13] br[13] wl[121] vdd gnd cell_6t
Xbit_r122_c13 bl[13] br[13] wl[122] vdd gnd cell_6t
Xbit_r123_c13 bl[13] br[13] wl[123] vdd gnd cell_6t
Xbit_r124_c13 bl[13] br[13] wl[124] vdd gnd cell_6t
Xbit_r125_c13 bl[13] br[13] wl[125] vdd gnd cell_6t
Xbit_r126_c13 bl[13] br[13] wl[126] vdd gnd cell_6t
Xbit_r127_c13 bl[13] br[13] wl[127] vdd gnd cell_6t
Xbit_r128_c13 bl[13] br[13] wl[128] vdd gnd cell_6t
Xbit_r129_c13 bl[13] br[13] wl[129] vdd gnd cell_6t
Xbit_r130_c13 bl[13] br[13] wl[130] vdd gnd cell_6t
Xbit_r131_c13 bl[13] br[13] wl[131] vdd gnd cell_6t
Xbit_r132_c13 bl[13] br[13] wl[132] vdd gnd cell_6t
Xbit_r133_c13 bl[13] br[13] wl[133] vdd gnd cell_6t
Xbit_r134_c13 bl[13] br[13] wl[134] vdd gnd cell_6t
Xbit_r135_c13 bl[13] br[13] wl[135] vdd gnd cell_6t
Xbit_r136_c13 bl[13] br[13] wl[136] vdd gnd cell_6t
Xbit_r137_c13 bl[13] br[13] wl[137] vdd gnd cell_6t
Xbit_r138_c13 bl[13] br[13] wl[138] vdd gnd cell_6t
Xbit_r139_c13 bl[13] br[13] wl[139] vdd gnd cell_6t
Xbit_r140_c13 bl[13] br[13] wl[140] vdd gnd cell_6t
Xbit_r141_c13 bl[13] br[13] wl[141] vdd gnd cell_6t
Xbit_r142_c13 bl[13] br[13] wl[142] vdd gnd cell_6t
Xbit_r143_c13 bl[13] br[13] wl[143] vdd gnd cell_6t
Xbit_r144_c13 bl[13] br[13] wl[144] vdd gnd cell_6t
Xbit_r145_c13 bl[13] br[13] wl[145] vdd gnd cell_6t
Xbit_r146_c13 bl[13] br[13] wl[146] vdd gnd cell_6t
Xbit_r147_c13 bl[13] br[13] wl[147] vdd gnd cell_6t
Xbit_r148_c13 bl[13] br[13] wl[148] vdd gnd cell_6t
Xbit_r149_c13 bl[13] br[13] wl[149] vdd gnd cell_6t
Xbit_r150_c13 bl[13] br[13] wl[150] vdd gnd cell_6t
Xbit_r151_c13 bl[13] br[13] wl[151] vdd gnd cell_6t
Xbit_r152_c13 bl[13] br[13] wl[152] vdd gnd cell_6t
Xbit_r153_c13 bl[13] br[13] wl[153] vdd gnd cell_6t
Xbit_r154_c13 bl[13] br[13] wl[154] vdd gnd cell_6t
Xbit_r155_c13 bl[13] br[13] wl[155] vdd gnd cell_6t
Xbit_r156_c13 bl[13] br[13] wl[156] vdd gnd cell_6t
Xbit_r157_c13 bl[13] br[13] wl[157] vdd gnd cell_6t
Xbit_r158_c13 bl[13] br[13] wl[158] vdd gnd cell_6t
Xbit_r159_c13 bl[13] br[13] wl[159] vdd gnd cell_6t
Xbit_r160_c13 bl[13] br[13] wl[160] vdd gnd cell_6t
Xbit_r161_c13 bl[13] br[13] wl[161] vdd gnd cell_6t
Xbit_r162_c13 bl[13] br[13] wl[162] vdd gnd cell_6t
Xbit_r163_c13 bl[13] br[13] wl[163] vdd gnd cell_6t
Xbit_r164_c13 bl[13] br[13] wl[164] vdd gnd cell_6t
Xbit_r165_c13 bl[13] br[13] wl[165] vdd gnd cell_6t
Xbit_r166_c13 bl[13] br[13] wl[166] vdd gnd cell_6t
Xbit_r167_c13 bl[13] br[13] wl[167] vdd gnd cell_6t
Xbit_r168_c13 bl[13] br[13] wl[168] vdd gnd cell_6t
Xbit_r169_c13 bl[13] br[13] wl[169] vdd gnd cell_6t
Xbit_r170_c13 bl[13] br[13] wl[170] vdd gnd cell_6t
Xbit_r171_c13 bl[13] br[13] wl[171] vdd gnd cell_6t
Xbit_r172_c13 bl[13] br[13] wl[172] vdd gnd cell_6t
Xbit_r173_c13 bl[13] br[13] wl[173] vdd gnd cell_6t
Xbit_r174_c13 bl[13] br[13] wl[174] vdd gnd cell_6t
Xbit_r175_c13 bl[13] br[13] wl[175] vdd gnd cell_6t
Xbit_r176_c13 bl[13] br[13] wl[176] vdd gnd cell_6t
Xbit_r177_c13 bl[13] br[13] wl[177] vdd gnd cell_6t
Xbit_r178_c13 bl[13] br[13] wl[178] vdd gnd cell_6t
Xbit_r179_c13 bl[13] br[13] wl[179] vdd gnd cell_6t
Xbit_r180_c13 bl[13] br[13] wl[180] vdd gnd cell_6t
Xbit_r181_c13 bl[13] br[13] wl[181] vdd gnd cell_6t
Xbit_r182_c13 bl[13] br[13] wl[182] vdd gnd cell_6t
Xbit_r183_c13 bl[13] br[13] wl[183] vdd gnd cell_6t
Xbit_r184_c13 bl[13] br[13] wl[184] vdd gnd cell_6t
Xbit_r185_c13 bl[13] br[13] wl[185] vdd gnd cell_6t
Xbit_r186_c13 bl[13] br[13] wl[186] vdd gnd cell_6t
Xbit_r187_c13 bl[13] br[13] wl[187] vdd gnd cell_6t
Xbit_r188_c13 bl[13] br[13] wl[188] vdd gnd cell_6t
Xbit_r189_c13 bl[13] br[13] wl[189] vdd gnd cell_6t
Xbit_r190_c13 bl[13] br[13] wl[190] vdd gnd cell_6t
Xbit_r191_c13 bl[13] br[13] wl[191] vdd gnd cell_6t
Xbit_r192_c13 bl[13] br[13] wl[192] vdd gnd cell_6t
Xbit_r193_c13 bl[13] br[13] wl[193] vdd gnd cell_6t
Xbit_r194_c13 bl[13] br[13] wl[194] vdd gnd cell_6t
Xbit_r195_c13 bl[13] br[13] wl[195] vdd gnd cell_6t
Xbit_r196_c13 bl[13] br[13] wl[196] vdd gnd cell_6t
Xbit_r197_c13 bl[13] br[13] wl[197] vdd gnd cell_6t
Xbit_r198_c13 bl[13] br[13] wl[198] vdd gnd cell_6t
Xbit_r199_c13 bl[13] br[13] wl[199] vdd gnd cell_6t
Xbit_r200_c13 bl[13] br[13] wl[200] vdd gnd cell_6t
Xbit_r201_c13 bl[13] br[13] wl[201] vdd gnd cell_6t
Xbit_r202_c13 bl[13] br[13] wl[202] vdd gnd cell_6t
Xbit_r203_c13 bl[13] br[13] wl[203] vdd gnd cell_6t
Xbit_r204_c13 bl[13] br[13] wl[204] vdd gnd cell_6t
Xbit_r205_c13 bl[13] br[13] wl[205] vdd gnd cell_6t
Xbit_r206_c13 bl[13] br[13] wl[206] vdd gnd cell_6t
Xbit_r207_c13 bl[13] br[13] wl[207] vdd gnd cell_6t
Xbit_r208_c13 bl[13] br[13] wl[208] vdd gnd cell_6t
Xbit_r209_c13 bl[13] br[13] wl[209] vdd gnd cell_6t
Xbit_r210_c13 bl[13] br[13] wl[210] vdd gnd cell_6t
Xbit_r211_c13 bl[13] br[13] wl[211] vdd gnd cell_6t
Xbit_r212_c13 bl[13] br[13] wl[212] vdd gnd cell_6t
Xbit_r213_c13 bl[13] br[13] wl[213] vdd gnd cell_6t
Xbit_r214_c13 bl[13] br[13] wl[214] vdd gnd cell_6t
Xbit_r215_c13 bl[13] br[13] wl[215] vdd gnd cell_6t
Xbit_r216_c13 bl[13] br[13] wl[216] vdd gnd cell_6t
Xbit_r217_c13 bl[13] br[13] wl[217] vdd gnd cell_6t
Xbit_r218_c13 bl[13] br[13] wl[218] vdd gnd cell_6t
Xbit_r219_c13 bl[13] br[13] wl[219] vdd gnd cell_6t
Xbit_r220_c13 bl[13] br[13] wl[220] vdd gnd cell_6t
Xbit_r221_c13 bl[13] br[13] wl[221] vdd gnd cell_6t
Xbit_r222_c13 bl[13] br[13] wl[222] vdd gnd cell_6t
Xbit_r223_c13 bl[13] br[13] wl[223] vdd gnd cell_6t
Xbit_r224_c13 bl[13] br[13] wl[224] vdd gnd cell_6t
Xbit_r225_c13 bl[13] br[13] wl[225] vdd gnd cell_6t
Xbit_r226_c13 bl[13] br[13] wl[226] vdd gnd cell_6t
Xbit_r227_c13 bl[13] br[13] wl[227] vdd gnd cell_6t
Xbit_r228_c13 bl[13] br[13] wl[228] vdd gnd cell_6t
Xbit_r229_c13 bl[13] br[13] wl[229] vdd gnd cell_6t
Xbit_r230_c13 bl[13] br[13] wl[230] vdd gnd cell_6t
Xbit_r231_c13 bl[13] br[13] wl[231] vdd gnd cell_6t
Xbit_r232_c13 bl[13] br[13] wl[232] vdd gnd cell_6t
Xbit_r233_c13 bl[13] br[13] wl[233] vdd gnd cell_6t
Xbit_r234_c13 bl[13] br[13] wl[234] vdd gnd cell_6t
Xbit_r235_c13 bl[13] br[13] wl[235] vdd gnd cell_6t
Xbit_r236_c13 bl[13] br[13] wl[236] vdd gnd cell_6t
Xbit_r237_c13 bl[13] br[13] wl[237] vdd gnd cell_6t
Xbit_r238_c13 bl[13] br[13] wl[238] vdd gnd cell_6t
Xbit_r239_c13 bl[13] br[13] wl[239] vdd gnd cell_6t
Xbit_r240_c13 bl[13] br[13] wl[240] vdd gnd cell_6t
Xbit_r241_c13 bl[13] br[13] wl[241] vdd gnd cell_6t
Xbit_r242_c13 bl[13] br[13] wl[242] vdd gnd cell_6t
Xbit_r243_c13 bl[13] br[13] wl[243] vdd gnd cell_6t
Xbit_r244_c13 bl[13] br[13] wl[244] vdd gnd cell_6t
Xbit_r245_c13 bl[13] br[13] wl[245] vdd gnd cell_6t
Xbit_r246_c13 bl[13] br[13] wl[246] vdd gnd cell_6t
Xbit_r247_c13 bl[13] br[13] wl[247] vdd gnd cell_6t
Xbit_r248_c13 bl[13] br[13] wl[248] vdd gnd cell_6t
Xbit_r249_c13 bl[13] br[13] wl[249] vdd gnd cell_6t
Xbit_r250_c13 bl[13] br[13] wl[250] vdd gnd cell_6t
Xbit_r251_c13 bl[13] br[13] wl[251] vdd gnd cell_6t
Xbit_r252_c13 bl[13] br[13] wl[252] vdd gnd cell_6t
Xbit_r253_c13 bl[13] br[13] wl[253] vdd gnd cell_6t
Xbit_r254_c13 bl[13] br[13] wl[254] vdd gnd cell_6t
Xbit_r255_c13 bl[13] br[13] wl[255] vdd gnd cell_6t
Xbit_r0_c14 bl[14] br[14] wl[0] vdd gnd cell_6t
Xbit_r1_c14 bl[14] br[14] wl[1] vdd gnd cell_6t
Xbit_r2_c14 bl[14] br[14] wl[2] vdd gnd cell_6t
Xbit_r3_c14 bl[14] br[14] wl[3] vdd gnd cell_6t
Xbit_r4_c14 bl[14] br[14] wl[4] vdd gnd cell_6t
Xbit_r5_c14 bl[14] br[14] wl[5] vdd gnd cell_6t
Xbit_r6_c14 bl[14] br[14] wl[6] vdd gnd cell_6t
Xbit_r7_c14 bl[14] br[14] wl[7] vdd gnd cell_6t
Xbit_r8_c14 bl[14] br[14] wl[8] vdd gnd cell_6t
Xbit_r9_c14 bl[14] br[14] wl[9] vdd gnd cell_6t
Xbit_r10_c14 bl[14] br[14] wl[10] vdd gnd cell_6t
Xbit_r11_c14 bl[14] br[14] wl[11] vdd gnd cell_6t
Xbit_r12_c14 bl[14] br[14] wl[12] vdd gnd cell_6t
Xbit_r13_c14 bl[14] br[14] wl[13] vdd gnd cell_6t
Xbit_r14_c14 bl[14] br[14] wl[14] vdd gnd cell_6t
Xbit_r15_c14 bl[14] br[14] wl[15] vdd gnd cell_6t
Xbit_r16_c14 bl[14] br[14] wl[16] vdd gnd cell_6t
Xbit_r17_c14 bl[14] br[14] wl[17] vdd gnd cell_6t
Xbit_r18_c14 bl[14] br[14] wl[18] vdd gnd cell_6t
Xbit_r19_c14 bl[14] br[14] wl[19] vdd gnd cell_6t
Xbit_r20_c14 bl[14] br[14] wl[20] vdd gnd cell_6t
Xbit_r21_c14 bl[14] br[14] wl[21] vdd gnd cell_6t
Xbit_r22_c14 bl[14] br[14] wl[22] vdd gnd cell_6t
Xbit_r23_c14 bl[14] br[14] wl[23] vdd gnd cell_6t
Xbit_r24_c14 bl[14] br[14] wl[24] vdd gnd cell_6t
Xbit_r25_c14 bl[14] br[14] wl[25] vdd gnd cell_6t
Xbit_r26_c14 bl[14] br[14] wl[26] vdd gnd cell_6t
Xbit_r27_c14 bl[14] br[14] wl[27] vdd gnd cell_6t
Xbit_r28_c14 bl[14] br[14] wl[28] vdd gnd cell_6t
Xbit_r29_c14 bl[14] br[14] wl[29] vdd gnd cell_6t
Xbit_r30_c14 bl[14] br[14] wl[30] vdd gnd cell_6t
Xbit_r31_c14 bl[14] br[14] wl[31] vdd gnd cell_6t
Xbit_r32_c14 bl[14] br[14] wl[32] vdd gnd cell_6t
Xbit_r33_c14 bl[14] br[14] wl[33] vdd gnd cell_6t
Xbit_r34_c14 bl[14] br[14] wl[34] vdd gnd cell_6t
Xbit_r35_c14 bl[14] br[14] wl[35] vdd gnd cell_6t
Xbit_r36_c14 bl[14] br[14] wl[36] vdd gnd cell_6t
Xbit_r37_c14 bl[14] br[14] wl[37] vdd gnd cell_6t
Xbit_r38_c14 bl[14] br[14] wl[38] vdd gnd cell_6t
Xbit_r39_c14 bl[14] br[14] wl[39] vdd gnd cell_6t
Xbit_r40_c14 bl[14] br[14] wl[40] vdd gnd cell_6t
Xbit_r41_c14 bl[14] br[14] wl[41] vdd gnd cell_6t
Xbit_r42_c14 bl[14] br[14] wl[42] vdd gnd cell_6t
Xbit_r43_c14 bl[14] br[14] wl[43] vdd gnd cell_6t
Xbit_r44_c14 bl[14] br[14] wl[44] vdd gnd cell_6t
Xbit_r45_c14 bl[14] br[14] wl[45] vdd gnd cell_6t
Xbit_r46_c14 bl[14] br[14] wl[46] vdd gnd cell_6t
Xbit_r47_c14 bl[14] br[14] wl[47] vdd gnd cell_6t
Xbit_r48_c14 bl[14] br[14] wl[48] vdd gnd cell_6t
Xbit_r49_c14 bl[14] br[14] wl[49] vdd gnd cell_6t
Xbit_r50_c14 bl[14] br[14] wl[50] vdd gnd cell_6t
Xbit_r51_c14 bl[14] br[14] wl[51] vdd gnd cell_6t
Xbit_r52_c14 bl[14] br[14] wl[52] vdd gnd cell_6t
Xbit_r53_c14 bl[14] br[14] wl[53] vdd gnd cell_6t
Xbit_r54_c14 bl[14] br[14] wl[54] vdd gnd cell_6t
Xbit_r55_c14 bl[14] br[14] wl[55] vdd gnd cell_6t
Xbit_r56_c14 bl[14] br[14] wl[56] vdd gnd cell_6t
Xbit_r57_c14 bl[14] br[14] wl[57] vdd gnd cell_6t
Xbit_r58_c14 bl[14] br[14] wl[58] vdd gnd cell_6t
Xbit_r59_c14 bl[14] br[14] wl[59] vdd gnd cell_6t
Xbit_r60_c14 bl[14] br[14] wl[60] vdd gnd cell_6t
Xbit_r61_c14 bl[14] br[14] wl[61] vdd gnd cell_6t
Xbit_r62_c14 bl[14] br[14] wl[62] vdd gnd cell_6t
Xbit_r63_c14 bl[14] br[14] wl[63] vdd gnd cell_6t
Xbit_r64_c14 bl[14] br[14] wl[64] vdd gnd cell_6t
Xbit_r65_c14 bl[14] br[14] wl[65] vdd gnd cell_6t
Xbit_r66_c14 bl[14] br[14] wl[66] vdd gnd cell_6t
Xbit_r67_c14 bl[14] br[14] wl[67] vdd gnd cell_6t
Xbit_r68_c14 bl[14] br[14] wl[68] vdd gnd cell_6t
Xbit_r69_c14 bl[14] br[14] wl[69] vdd gnd cell_6t
Xbit_r70_c14 bl[14] br[14] wl[70] vdd gnd cell_6t
Xbit_r71_c14 bl[14] br[14] wl[71] vdd gnd cell_6t
Xbit_r72_c14 bl[14] br[14] wl[72] vdd gnd cell_6t
Xbit_r73_c14 bl[14] br[14] wl[73] vdd gnd cell_6t
Xbit_r74_c14 bl[14] br[14] wl[74] vdd gnd cell_6t
Xbit_r75_c14 bl[14] br[14] wl[75] vdd gnd cell_6t
Xbit_r76_c14 bl[14] br[14] wl[76] vdd gnd cell_6t
Xbit_r77_c14 bl[14] br[14] wl[77] vdd gnd cell_6t
Xbit_r78_c14 bl[14] br[14] wl[78] vdd gnd cell_6t
Xbit_r79_c14 bl[14] br[14] wl[79] vdd gnd cell_6t
Xbit_r80_c14 bl[14] br[14] wl[80] vdd gnd cell_6t
Xbit_r81_c14 bl[14] br[14] wl[81] vdd gnd cell_6t
Xbit_r82_c14 bl[14] br[14] wl[82] vdd gnd cell_6t
Xbit_r83_c14 bl[14] br[14] wl[83] vdd gnd cell_6t
Xbit_r84_c14 bl[14] br[14] wl[84] vdd gnd cell_6t
Xbit_r85_c14 bl[14] br[14] wl[85] vdd gnd cell_6t
Xbit_r86_c14 bl[14] br[14] wl[86] vdd gnd cell_6t
Xbit_r87_c14 bl[14] br[14] wl[87] vdd gnd cell_6t
Xbit_r88_c14 bl[14] br[14] wl[88] vdd gnd cell_6t
Xbit_r89_c14 bl[14] br[14] wl[89] vdd gnd cell_6t
Xbit_r90_c14 bl[14] br[14] wl[90] vdd gnd cell_6t
Xbit_r91_c14 bl[14] br[14] wl[91] vdd gnd cell_6t
Xbit_r92_c14 bl[14] br[14] wl[92] vdd gnd cell_6t
Xbit_r93_c14 bl[14] br[14] wl[93] vdd gnd cell_6t
Xbit_r94_c14 bl[14] br[14] wl[94] vdd gnd cell_6t
Xbit_r95_c14 bl[14] br[14] wl[95] vdd gnd cell_6t
Xbit_r96_c14 bl[14] br[14] wl[96] vdd gnd cell_6t
Xbit_r97_c14 bl[14] br[14] wl[97] vdd gnd cell_6t
Xbit_r98_c14 bl[14] br[14] wl[98] vdd gnd cell_6t
Xbit_r99_c14 bl[14] br[14] wl[99] vdd gnd cell_6t
Xbit_r100_c14 bl[14] br[14] wl[100] vdd gnd cell_6t
Xbit_r101_c14 bl[14] br[14] wl[101] vdd gnd cell_6t
Xbit_r102_c14 bl[14] br[14] wl[102] vdd gnd cell_6t
Xbit_r103_c14 bl[14] br[14] wl[103] vdd gnd cell_6t
Xbit_r104_c14 bl[14] br[14] wl[104] vdd gnd cell_6t
Xbit_r105_c14 bl[14] br[14] wl[105] vdd gnd cell_6t
Xbit_r106_c14 bl[14] br[14] wl[106] vdd gnd cell_6t
Xbit_r107_c14 bl[14] br[14] wl[107] vdd gnd cell_6t
Xbit_r108_c14 bl[14] br[14] wl[108] vdd gnd cell_6t
Xbit_r109_c14 bl[14] br[14] wl[109] vdd gnd cell_6t
Xbit_r110_c14 bl[14] br[14] wl[110] vdd gnd cell_6t
Xbit_r111_c14 bl[14] br[14] wl[111] vdd gnd cell_6t
Xbit_r112_c14 bl[14] br[14] wl[112] vdd gnd cell_6t
Xbit_r113_c14 bl[14] br[14] wl[113] vdd gnd cell_6t
Xbit_r114_c14 bl[14] br[14] wl[114] vdd gnd cell_6t
Xbit_r115_c14 bl[14] br[14] wl[115] vdd gnd cell_6t
Xbit_r116_c14 bl[14] br[14] wl[116] vdd gnd cell_6t
Xbit_r117_c14 bl[14] br[14] wl[117] vdd gnd cell_6t
Xbit_r118_c14 bl[14] br[14] wl[118] vdd gnd cell_6t
Xbit_r119_c14 bl[14] br[14] wl[119] vdd gnd cell_6t
Xbit_r120_c14 bl[14] br[14] wl[120] vdd gnd cell_6t
Xbit_r121_c14 bl[14] br[14] wl[121] vdd gnd cell_6t
Xbit_r122_c14 bl[14] br[14] wl[122] vdd gnd cell_6t
Xbit_r123_c14 bl[14] br[14] wl[123] vdd gnd cell_6t
Xbit_r124_c14 bl[14] br[14] wl[124] vdd gnd cell_6t
Xbit_r125_c14 bl[14] br[14] wl[125] vdd gnd cell_6t
Xbit_r126_c14 bl[14] br[14] wl[126] vdd gnd cell_6t
Xbit_r127_c14 bl[14] br[14] wl[127] vdd gnd cell_6t
Xbit_r128_c14 bl[14] br[14] wl[128] vdd gnd cell_6t
Xbit_r129_c14 bl[14] br[14] wl[129] vdd gnd cell_6t
Xbit_r130_c14 bl[14] br[14] wl[130] vdd gnd cell_6t
Xbit_r131_c14 bl[14] br[14] wl[131] vdd gnd cell_6t
Xbit_r132_c14 bl[14] br[14] wl[132] vdd gnd cell_6t
Xbit_r133_c14 bl[14] br[14] wl[133] vdd gnd cell_6t
Xbit_r134_c14 bl[14] br[14] wl[134] vdd gnd cell_6t
Xbit_r135_c14 bl[14] br[14] wl[135] vdd gnd cell_6t
Xbit_r136_c14 bl[14] br[14] wl[136] vdd gnd cell_6t
Xbit_r137_c14 bl[14] br[14] wl[137] vdd gnd cell_6t
Xbit_r138_c14 bl[14] br[14] wl[138] vdd gnd cell_6t
Xbit_r139_c14 bl[14] br[14] wl[139] vdd gnd cell_6t
Xbit_r140_c14 bl[14] br[14] wl[140] vdd gnd cell_6t
Xbit_r141_c14 bl[14] br[14] wl[141] vdd gnd cell_6t
Xbit_r142_c14 bl[14] br[14] wl[142] vdd gnd cell_6t
Xbit_r143_c14 bl[14] br[14] wl[143] vdd gnd cell_6t
Xbit_r144_c14 bl[14] br[14] wl[144] vdd gnd cell_6t
Xbit_r145_c14 bl[14] br[14] wl[145] vdd gnd cell_6t
Xbit_r146_c14 bl[14] br[14] wl[146] vdd gnd cell_6t
Xbit_r147_c14 bl[14] br[14] wl[147] vdd gnd cell_6t
Xbit_r148_c14 bl[14] br[14] wl[148] vdd gnd cell_6t
Xbit_r149_c14 bl[14] br[14] wl[149] vdd gnd cell_6t
Xbit_r150_c14 bl[14] br[14] wl[150] vdd gnd cell_6t
Xbit_r151_c14 bl[14] br[14] wl[151] vdd gnd cell_6t
Xbit_r152_c14 bl[14] br[14] wl[152] vdd gnd cell_6t
Xbit_r153_c14 bl[14] br[14] wl[153] vdd gnd cell_6t
Xbit_r154_c14 bl[14] br[14] wl[154] vdd gnd cell_6t
Xbit_r155_c14 bl[14] br[14] wl[155] vdd gnd cell_6t
Xbit_r156_c14 bl[14] br[14] wl[156] vdd gnd cell_6t
Xbit_r157_c14 bl[14] br[14] wl[157] vdd gnd cell_6t
Xbit_r158_c14 bl[14] br[14] wl[158] vdd gnd cell_6t
Xbit_r159_c14 bl[14] br[14] wl[159] vdd gnd cell_6t
Xbit_r160_c14 bl[14] br[14] wl[160] vdd gnd cell_6t
Xbit_r161_c14 bl[14] br[14] wl[161] vdd gnd cell_6t
Xbit_r162_c14 bl[14] br[14] wl[162] vdd gnd cell_6t
Xbit_r163_c14 bl[14] br[14] wl[163] vdd gnd cell_6t
Xbit_r164_c14 bl[14] br[14] wl[164] vdd gnd cell_6t
Xbit_r165_c14 bl[14] br[14] wl[165] vdd gnd cell_6t
Xbit_r166_c14 bl[14] br[14] wl[166] vdd gnd cell_6t
Xbit_r167_c14 bl[14] br[14] wl[167] vdd gnd cell_6t
Xbit_r168_c14 bl[14] br[14] wl[168] vdd gnd cell_6t
Xbit_r169_c14 bl[14] br[14] wl[169] vdd gnd cell_6t
Xbit_r170_c14 bl[14] br[14] wl[170] vdd gnd cell_6t
Xbit_r171_c14 bl[14] br[14] wl[171] vdd gnd cell_6t
Xbit_r172_c14 bl[14] br[14] wl[172] vdd gnd cell_6t
Xbit_r173_c14 bl[14] br[14] wl[173] vdd gnd cell_6t
Xbit_r174_c14 bl[14] br[14] wl[174] vdd gnd cell_6t
Xbit_r175_c14 bl[14] br[14] wl[175] vdd gnd cell_6t
Xbit_r176_c14 bl[14] br[14] wl[176] vdd gnd cell_6t
Xbit_r177_c14 bl[14] br[14] wl[177] vdd gnd cell_6t
Xbit_r178_c14 bl[14] br[14] wl[178] vdd gnd cell_6t
Xbit_r179_c14 bl[14] br[14] wl[179] vdd gnd cell_6t
Xbit_r180_c14 bl[14] br[14] wl[180] vdd gnd cell_6t
Xbit_r181_c14 bl[14] br[14] wl[181] vdd gnd cell_6t
Xbit_r182_c14 bl[14] br[14] wl[182] vdd gnd cell_6t
Xbit_r183_c14 bl[14] br[14] wl[183] vdd gnd cell_6t
Xbit_r184_c14 bl[14] br[14] wl[184] vdd gnd cell_6t
Xbit_r185_c14 bl[14] br[14] wl[185] vdd gnd cell_6t
Xbit_r186_c14 bl[14] br[14] wl[186] vdd gnd cell_6t
Xbit_r187_c14 bl[14] br[14] wl[187] vdd gnd cell_6t
Xbit_r188_c14 bl[14] br[14] wl[188] vdd gnd cell_6t
Xbit_r189_c14 bl[14] br[14] wl[189] vdd gnd cell_6t
Xbit_r190_c14 bl[14] br[14] wl[190] vdd gnd cell_6t
Xbit_r191_c14 bl[14] br[14] wl[191] vdd gnd cell_6t
Xbit_r192_c14 bl[14] br[14] wl[192] vdd gnd cell_6t
Xbit_r193_c14 bl[14] br[14] wl[193] vdd gnd cell_6t
Xbit_r194_c14 bl[14] br[14] wl[194] vdd gnd cell_6t
Xbit_r195_c14 bl[14] br[14] wl[195] vdd gnd cell_6t
Xbit_r196_c14 bl[14] br[14] wl[196] vdd gnd cell_6t
Xbit_r197_c14 bl[14] br[14] wl[197] vdd gnd cell_6t
Xbit_r198_c14 bl[14] br[14] wl[198] vdd gnd cell_6t
Xbit_r199_c14 bl[14] br[14] wl[199] vdd gnd cell_6t
Xbit_r200_c14 bl[14] br[14] wl[200] vdd gnd cell_6t
Xbit_r201_c14 bl[14] br[14] wl[201] vdd gnd cell_6t
Xbit_r202_c14 bl[14] br[14] wl[202] vdd gnd cell_6t
Xbit_r203_c14 bl[14] br[14] wl[203] vdd gnd cell_6t
Xbit_r204_c14 bl[14] br[14] wl[204] vdd gnd cell_6t
Xbit_r205_c14 bl[14] br[14] wl[205] vdd gnd cell_6t
Xbit_r206_c14 bl[14] br[14] wl[206] vdd gnd cell_6t
Xbit_r207_c14 bl[14] br[14] wl[207] vdd gnd cell_6t
Xbit_r208_c14 bl[14] br[14] wl[208] vdd gnd cell_6t
Xbit_r209_c14 bl[14] br[14] wl[209] vdd gnd cell_6t
Xbit_r210_c14 bl[14] br[14] wl[210] vdd gnd cell_6t
Xbit_r211_c14 bl[14] br[14] wl[211] vdd gnd cell_6t
Xbit_r212_c14 bl[14] br[14] wl[212] vdd gnd cell_6t
Xbit_r213_c14 bl[14] br[14] wl[213] vdd gnd cell_6t
Xbit_r214_c14 bl[14] br[14] wl[214] vdd gnd cell_6t
Xbit_r215_c14 bl[14] br[14] wl[215] vdd gnd cell_6t
Xbit_r216_c14 bl[14] br[14] wl[216] vdd gnd cell_6t
Xbit_r217_c14 bl[14] br[14] wl[217] vdd gnd cell_6t
Xbit_r218_c14 bl[14] br[14] wl[218] vdd gnd cell_6t
Xbit_r219_c14 bl[14] br[14] wl[219] vdd gnd cell_6t
Xbit_r220_c14 bl[14] br[14] wl[220] vdd gnd cell_6t
Xbit_r221_c14 bl[14] br[14] wl[221] vdd gnd cell_6t
Xbit_r222_c14 bl[14] br[14] wl[222] vdd gnd cell_6t
Xbit_r223_c14 bl[14] br[14] wl[223] vdd gnd cell_6t
Xbit_r224_c14 bl[14] br[14] wl[224] vdd gnd cell_6t
Xbit_r225_c14 bl[14] br[14] wl[225] vdd gnd cell_6t
Xbit_r226_c14 bl[14] br[14] wl[226] vdd gnd cell_6t
Xbit_r227_c14 bl[14] br[14] wl[227] vdd gnd cell_6t
Xbit_r228_c14 bl[14] br[14] wl[228] vdd gnd cell_6t
Xbit_r229_c14 bl[14] br[14] wl[229] vdd gnd cell_6t
Xbit_r230_c14 bl[14] br[14] wl[230] vdd gnd cell_6t
Xbit_r231_c14 bl[14] br[14] wl[231] vdd gnd cell_6t
Xbit_r232_c14 bl[14] br[14] wl[232] vdd gnd cell_6t
Xbit_r233_c14 bl[14] br[14] wl[233] vdd gnd cell_6t
Xbit_r234_c14 bl[14] br[14] wl[234] vdd gnd cell_6t
Xbit_r235_c14 bl[14] br[14] wl[235] vdd gnd cell_6t
Xbit_r236_c14 bl[14] br[14] wl[236] vdd gnd cell_6t
Xbit_r237_c14 bl[14] br[14] wl[237] vdd gnd cell_6t
Xbit_r238_c14 bl[14] br[14] wl[238] vdd gnd cell_6t
Xbit_r239_c14 bl[14] br[14] wl[239] vdd gnd cell_6t
Xbit_r240_c14 bl[14] br[14] wl[240] vdd gnd cell_6t
Xbit_r241_c14 bl[14] br[14] wl[241] vdd gnd cell_6t
Xbit_r242_c14 bl[14] br[14] wl[242] vdd gnd cell_6t
Xbit_r243_c14 bl[14] br[14] wl[243] vdd gnd cell_6t
Xbit_r244_c14 bl[14] br[14] wl[244] vdd gnd cell_6t
Xbit_r245_c14 bl[14] br[14] wl[245] vdd gnd cell_6t
Xbit_r246_c14 bl[14] br[14] wl[246] vdd gnd cell_6t
Xbit_r247_c14 bl[14] br[14] wl[247] vdd gnd cell_6t
Xbit_r248_c14 bl[14] br[14] wl[248] vdd gnd cell_6t
Xbit_r249_c14 bl[14] br[14] wl[249] vdd gnd cell_6t
Xbit_r250_c14 bl[14] br[14] wl[250] vdd gnd cell_6t
Xbit_r251_c14 bl[14] br[14] wl[251] vdd gnd cell_6t
Xbit_r252_c14 bl[14] br[14] wl[252] vdd gnd cell_6t
Xbit_r253_c14 bl[14] br[14] wl[253] vdd gnd cell_6t
Xbit_r254_c14 bl[14] br[14] wl[254] vdd gnd cell_6t
Xbit_r255_c14 bl[14] br[14] wl[255] vdd gnd cell_6t
Xbit_r0_c15 bl[15] br[15] wl[0] vdd gnd cell_6t
Xbit_r1_c15 bl[15] br[15] wl[1] vdd gnd cell_6t
Xbit_r2_c15 bl[15] br[15] wl[2] vdd gnd cell_6t
Xbit_r3_c15 bl[15] br[15] wl[3] vdd gnd cell_6t
Xbit_r4_c15 bl[15] br[15] wl[4] vdd gnd cell_6t
Xbit_r5_c15 bl[15] br[15] wl[5] vdd gnd cell_6t
Xbit_r6_c15 bl[15] br[15] wl[6] vdd gnd cell_6t
Xbit_r7_c15 bl[15] br[15] wl[7] vdd gnd cell_6t
Xbit_r8_c15 bl[15] br[15] wl[8] vdd gnd cell_6t
Xbit_r9_c15 bl[15] br[15] wl[9] vdd gnd cell_6t
Xbit_r10_c15 bl[15] br[15] wl[10] vdd gnd cell_6t
Xbit_r11_c15 bl[15] br[15] wl[11] vdd gnd cell_6t
Xbit_r12_c15 bl[15] br[15] wl[12] vdd gnd cell_6t
Xbit_r13_c15 bl[15] br[15] wl[13] vdd gnd cell_6t
Xbit_r14_c15 bl[15] br[15] wl[14] vdd gnd cell_6t
Xbit_r15_c15 bl[15] br[15] wl[15] vdd gnd cell_6t
Xbit_r16_c15 bl[15] br[15] wl[16] vdd gnd cell_6t
Xbit_r17_c15 bl[15] br[15] wl[17] vdd gnd cell_6t
Xbit_r18_c15 bl[15] br[15] wl[18] vdd gnd cell_6t
Xbit_r19_c15 bl[15] br[15] wl[19] vdd gnd cell_6t
Xbit_r20_c15 bl[15] br[15] wl[20] vdd gnd cell_6t
Xbit_r21_c15 bl[15] br[15] wl[21] vdd gnd cell_6t
Xbit_r22_c15 bl[15] br[15] wl[22] vdd gnd cell_6t
Xbit_r23_c15 bl[15] br[15] wl[23] vdd gnd cell_6t
Xbit_r24_c15 bl[15] br[15] wl[24] vdd gnd cell_6t
Xbit_r25_c15 bl[15] br[15] wl[25] vdd gnd cell_6t
Xbit_r26_c15 bl[15] br[15] wl[26] vdd gnd cell_6t
Xbit_r27_c15 bl[15] br[15] wl[27] vdd gnd cell_6t
Xbit_r28_c15 bl[15] br[15] wl[28] vdd gnd cell_6t
Xbit_r29_c15 bl[15] br[15] wl[29] vdd gnd cell_6t
Xbit_r30_c15 bl[15] br[15] wl[30] vdd gnd cell_6t
Xbit_r31_c15 bl[15] br[15] wl[31] vdd gnd cell_6t
Xbit_r32_c15 bl[15] br[15] wl[32] vdd gnd cell_6t
Xbit_r33_c15 bl[15] br[15] wl[33] vdd gnd cell_6t
Xbit_r34_c15 bl[15] br[15] wl[34] vdd gnd cell_6t
Xbit_r35_c15 bl[15] br[15] wl[35] vdd gnd cell_6t
Xbit_r36_c15 bl[15] br[15] wl[36] vdd gnd cell_6t
Xbit_r37_c15 bl[15] br[15] wl[37] vdd gnd cell_6t
Xbit_r38_c15 bl[15] br[15] wl[38] vdd gnd cell_6t
Xbit_r39_c15 bl[15] br[15] wl[39] vdd gnd cell_6t
Xbit_r40_c15 bl[15] br[15] wl[40] vdd gnd cell_6t
Xbit_r41_c15 bl[15] br[15] wl[41] vdd gnd cell_6t
Xbit_r42_c15 bl[15] br[15] wl[42] vdd gnd cell_6t
Xbit_r43_c15 bl[15] br[15] wl[43] vdd gnd cell_6t
Xbit_r44_c15 bl[15] br[15] wl[44] vdd gnd cell_6t
Xbit_r45_c15 bl[15] br[15] wl[45] vdd gnd cell_6t
Xbit_r46_c15 bl[15] br[15] wl[46] vdd gnd cell_6t
Xbit_r47_c15 bl[15] br[15] wl[47] vdd gnd cell_6t
Xbit_r48_c15 bl[15] br[15] wl[48] vdd gnd cell_6t
Xbit_r49_c15 bl[15] br[15] wl[49] vdd gnd cell_6t
Xbit_r50_c15 bl[15] br[15] wl[50] vdd gnd cell_6t
Xbit_r51_c15 bl[15] br[15] wl[51] vdd gnd cell_6t
Xbit_r52_c15 bl[15] br[15] wl[52] vdd gnd cell_6t
Xbit_r53_c15 bl[15] br[15] wl[53] vdd gnd cell_6t
Xbit_r54_c15 bl[15] br[15] wl[54] vdd gnd cell_6t
Xbit_r55_c15 bl[15] br[15] wl[55] vdd gnd cell_6t
Xbit_r56_c15 bl[15] br[15] wl[56] vdd gnd cell_6t
Xbit_r57_c15 bl[15] br[15] wl[57] vdd gnd cell_6t
Xbit_r58_c15 bl[15] br[15] wl[58] vdd gnd cell_6t
Xbit_r59_c15 bl[15] br[15] wl[59] vdd gnd cell_6t
Xbit_r60_c15 bl[15] br[15] wl[60] vdd gnd cell_6t
Xbit_r61_c15 bl[15] br[15] wl[61] vdd gnd cell_6t
Xbit_r62_c15 bl[15] br[15] wl[62] vdd gnd cell_6t
Xbit_r63_c15 bl[15] br[15] wl[63] vdd gnd cell_6t
Xbit_r64_c15 bl[15] br[15] wl[64] vdd gnd cell_6t
Xbit_r65_c15 bl[15] br[15] wl[65] vdd gnd cell_6t
Xbit_r66_c15 bl[15] br[15] wl[66] vdd gnd cell_6t
Xbit_r67_c15 bl[15] br[15] wl[67] vdd gnd cell_6t
Xbit_r68_c15 bl[15] br[15] wl[68] vdd gnd cell_6t
Xbit_r69_c15 bl[15] br[15] wl[69] vdd gnd cell_6t
Xbit_r70_c15 bl[15] br[15] wl[70] vdd gnd cell_6t
Xbit_r71_c15 bl[15] br[15] wl[71] vdd gnd cell_6t
Xbit_r72_c15 bl[15] br[15] wl[72] vdd gnd cell_6t
Xbit_r73_c15 bl[15] br[15] wl[73] vdd gnd cell_6t
Xbit_r74_c15 bl[15] br[15] wl[74] vdd gnd cell_6t
Xbit_r75_c15 bl[15] br[15] wl[75] vdd gnd cell_6t
Xbit_r76_c15 bl[15] br[15] wl[76] vdd gnd cell_6t
Xbit_r77_c15 bl[15] br[15] wl[77] vdd gnd cell_6t
Xbit_r78_c15 bl[15] br[15] wl[78] vdd gnd cell_6t
Xbit_r79_c15 bl[15] br[15] wl[79] vdd gnd cell_6t
Xbit_r80_c15 bl[15] br[15] wl[80] vdd gnd cell_6t
Xbit_r81_c15 bl[15] br[15] wl[81] vdd gnd cell_6t
Xbit_r82_c15 bl[15] br[15] wl[82] vdd gnd cell_6t
Xbit_r83_c15 bl[15] br[15] wl[83] vdd gnd cell_6t
Xbit_r84_c15 bl[15] br[15] wl[84] vdd gnd cell_6t
Xbit_r85_c15 bl[15] br[15] wl[85] vdd gnd cell_6t
Xbit_r86_c15 bl[15] br[15] wl[86] vdd gnd cell_6t
Xbit_r87_c15 bl[15] br[15] wl[87] vdd gnd cell_6t
Xbit_r88_c15 bl[15] br[15] wl[88] vdd gnd cell_6t
Xbit_r89_c15 bl[15] br[15] wl[89] vdd gnd cell_6t
Xbit_r90_c15 bl[15] br[15] wl[90] vdd gnd cell_6t
Xbit_r91_c15 bl[15] br[15] wl[91] vdd gnd cell_6t
Xbit_r92_c15 bl[15] br[15] wl[92] vdd gnd cell_6t
Xbit_r93_c15 bl[15] br[15] wl[93] vdd gnd cell_6t
Xbit_r94_c15 bl[15] br[15] wl[94] vdd gnd cell_6t
Xbit_r95_c15 bl[15] br[15] wl[95] vdd gnd cell_6t
Xbit_r96_c15 bl[15] br[15] wl[96] vdd gnd cell_6t
Xbit_r97_c15 bl[15] br[15] wl[97] vdd gnd cell_6t
Xbit_r98_c15 bl[15] br[15] wl[98] vdd gnd cell_6t
Xbit_r99_c15 bl[15] br[15] wl[99] vdd gnd cell_6t
Xbit_r100_c15 bl[15] br[15] wl[100] vdd gnd cell_6t
Xbit_r101_c15 bl[15] br[15] wl[101] vdd gnd cell_6t
Xbit_r102_c15 bl[15] br[15] wl[102] vdd gnd cell_6t
Xbit_r103_c15 bl[15] br[15] wl[103] vdd gnd cell_6t
Xbit_r104_c15 bl[15] br[15] wl[104] vdd gnd cell_6t
Xbit_r105_c15 bl[15] br[15] wl[105] vdd gnd cell_6t
Xbit_r106_c15 bl[15] br[15] wl[106] vdd gnd cell_6t
Xbit_r107_c15 bl[15] br[15] wl[107] vdd gnd cell_6t
Xbit_r108_c15 bl[15] br[15] wl[108] vdd gnd cell_6t
Xbit_r109_c15 bl[15] br[15] wl[109] vdd gnd cell_6t
Xbit_r110_c15 bl[15] br[15] wl[110] vdd gnd cell_6t
Xbit_r111_c15 bl[15] br[15] wl[111] vdd gnd cell_6t
Xbit_r112_c15 bl[15] br[15] wl[112] vdd gnd cell_6t
Xbit_r113_c15 bl[15] br[15] wl[113] vdd gnd cell_6t
Xbit_r114_c15 bl[15] br[15] wl[114] vdd gnd cell_6t
Xbit_r115_c15 bl[15] br[15] wl[115] vdd gnd cell_6t
Xbit_r116_c15 bl[15] br[15] wl[116] vdd gnd cell_6t
Xbit_r117_c15 bl[15] br[15] wl[117] vdd gnd cell_6t
Xbit_r118_c15 bl[15] br[15] wl[118] vdd gnd cell_6t
Xbit_r119_c15 bl[15] br[15] wl[119] vdd gnd cell_6t
Xbit_r120_c15 bl[15] br[15] wl[120] vdd gnd cell_6t
Xbit_r121_c15 bl[15] br[15] wl[121] vdd gnd cell_6t
Xbit_r122_c15 bl[15] br[15] wl[122] vdd gnd cell_6t
Xbit_r123_c15 bl[15] br[15] wl[123] vdd gnd cell_6t
Xbit_r124_c15 bl[15] br[15] wl[124] vdd gnd cell_6t
Xbit_r125_c15 bl[15] br[15] wl[125] vdd gnd cell_6t
Xbit_r126_c15 bl[15] br[15] wl[126] vdd gnd cell_6t
Xbit_r127_c15 bl[15] br[15] wl[127] vdd gnd cell_6t
Xbit_r128_c15 bl[15] br[15] wl[128] vdd gnd cell_6t
Xbit_r129_c15 bl[15] br[15] wl[129] vdd gnd cell_6t
Xbit_r130_c15 bl[15] br[15] wl[130] vdd gnd cell_6t
Xbit_r131_c15 bl[15] br[15] wl[131] vdd gnd cell_6t
Xbit_r132_c15 bl[15] br[15] wl[132] vdd gnd cell_6t
Xbit_r133_c15 bl[15] br[15] wl[133] vdd gnd cell_6t
Xbit_r134_c15 bl[15] br[15] wl[134] vdd gnd cell_6t
Xbit_r135_c15 bl[15] br[15] wl[135] vdd gnd cell_6t
Xbit_r136_c15 bl[15] br[15] wl[136] vdd gnd cell_6t
Xbit_r137_c15 bl[15] br[15] wl[137] vdd gnd cell_6t
Xbit_r138_c15 bl[15] br[15] wl[138] vdd gnd cell_6t
Xbit_r139_c15 bl[15] br[15] wl[139] vdd gnd cell_6t
Xbit_r140_c15 bl[15] br[15] wl[140] vdd gnd cell_6t
Xbit_r141_c15 bl[15] br[15] wl[141] vdd gnd cell_6t
Xbit_r142_c15 bl[15] br[15] wl[142] vdd gnd cell_6t
Xbit_r143_c15 bl[15] br[15] wl[143] vdd gnd cell_6t
Xbit_r144_c15 bl[15] br[15] wl[144] vdd gnd cell_6t
Xbit_r145_c15 bl[15] br[15] wl[145] vdd gnd cell_6t
Xbit_r146_c15 bl[15] br[15] wl[146] vdd gnd cell_6t
Xbit_r147_c15 bl[15] br[15] wl[147] vdd gnd cell_6t
Xbit_r148_c15 bl[15] br[15] wl[148] vdd gnd cell_6t
Xbit_r149_c15 bl[15] br[15] wl[149] vdd gnd cell_6t
Xbit_r150_c15 bl[15] br[15] wl[150] vdd gnd cell_6t
Xbit_r151_c15 bl[15] br[15] wl[151] vdd gnd cell_6t
Xbit_r152_c15 bl[15] br[15] wl[152] vdd gnd cell_6t
Xbit_r153_c15 bl[15] br[15] wl[153] vdd gnd cell_6t
Xbit_r154_c15 bl[15] br[15] wl[154] vdd gnd cell_6t
Xbit_r155_c15 bl[15] br[15] wl[155] vdd gnd cell_6t
Xbit_r156_c15 bl[15] br[15] wl[156] vdd gnd cell_6t
Xbit_r157_c15 bl[15] br[15] wl[157] vdd gnd cell_6t
Xbit_r158_c15 bl[15] br[15] wl[158] vdd gnd cell_6t
Xbit_r159_c15 bl[15] br[15] wl[159] vdd gnd cell_6t
Xbit_r160_c15 bl[15] br[15] wl[160] vdd gnd cell_6t
Xbit_r161_c15 bl[15] br[15] wl[161] vdd gnd cell_6t
Xbit_r162_c15 bl[15] br[15] wl[162] vdd gnd cell_6t
Xbit_r163_c15 bl[15] br[15] wl[163] vdd gnd cell_6t
Xbit_r164_c15 bl[15] br[15] wl[164] vdd gnd cell_6t
Xbit_r165_c15 bl[15] br[15] wl[165] vdd gnd cell_6t
Xbit_r166_c15 bl[15] br[15] wl[166] vdd gnd cell_6t
Xbit_r167_c15 bl[15] br[15] wl[167] vdd gnd cell_6t
Xbit_r168_c15 bl[15] br[15] wl[168] vdd gnd cell_6t
Xbit_r169_c15 bl[15] br[15] wl[169] vdd gnd cell_6t
Xbit_r170_c15 bl[15] br[15] wl[170] vdd gnd cell_6t
Xbit_r171_c15 bl[15] br[15] wl[171] vdd gnd cell_6t
Xbit_r172_c15 bl[15] br[15] wl[172] vdd gnd cell_6t
Xbit_r173_c15 bl[15] br[15] wl[173] vdd gnd cell_6t
Xbit_r174_c15 bl[15] br[15] wl[174] vdd gnd cell_6t
Xbit_r175_c15 bl[15] br[15] wl[175] vdd gnd cell_6t
Xbit_r176_c15 bl[15] br[15] wl[176] vdd gnd cell_6t
Xbit_r177_c15 bl[15] br[15] wl[177] vdd gnd cell_6t
Xbit_r178_c15 bl[15] br[15] wl[178] vdd gnd cell_6t
Xbit_r179_c15 bl[15] br[15] wl[179] vdd gnd cell_6t
Xbit_r180_c15 bl[15] br[15] wl[180] vdd gnd cell_6t
Xbit_r181_c15 bl[15] br[15] wl[181] vdd gnd cell_6t
Xbit_r182_c15 bl[15] br[15] wl[182] vdd gnd cell_6t
Xbit_r183_c15 bl[15] br[15] wl[183] vdd gnd cell_6t
Xbit_r184_c15 bl[15] br[15] wl[184] vdd gnd cell_6t
Xbit_r185_c15 bl[15] br[15] wl[185] vdd gnd cell_6t
Xbit_r186_c15 bl[15] br[15] wl[186] vdd gnd cell_6t
Xbit_r187_c15 bl[15] br[15] wl[187] vdd gnd cell_6t
Xbit_r188_c15 bl[15] br[15] wl[188] vdd gnd cell_6t
Xbit_r189_c15 bl[15] br[15] wl[189] vdd gnd cell_6t
Xbit_r190_c15 bl[15] br[15] wl[190] vdd gnd cell_6t
Xbit_r191_c15 bl[15] br[15] wl[191] vdd gnd cell_6t
Xbit_r192_c15 bl[15] br[15] wl[192] vdd gnd cell_6t
Xbit_r193_c15 bl[15] br[15] wl[193] vdd gnd cell_6t
Xbit_r194_c15 bl[15] br[15] wl[194] vdd gnd cell_6t
Xbit_r195_c15 bl[15] br[15] wl[195] vdd gnd cell_6t
Xbit_r196_c15 bl[15] br[15] wl[196] vdd gnd cell_6t
Xbit_r197_c15 bl[15] br[15] wl[197] vdd gnd cell_6t
Xbit_r198_c15 bl[15] br[15] wl[198] vdd gnd cell_6t
Xbit_r199_c15 bl[15] br[15] wl[199] vdd gnd cell_6t
Xbit_r200_c15 bl[15] br[15] wl[200] vdd gnd cell_6t
Xbit_r201_c15 bl[15] br[15] wl[201] vdd gnd cell_6t
Xbit_r202_c15 bl[15] br[15] wl[202] vdd gnd cell_6t
Xbit_r203_c15 bl[15] br[15] wl[203] vdd gnd cell_6t
Xbit_r204_c15 bl[15] br[15] wl[204] vdd gnd cell_6t
Xbit_r205_c15 bl[15] br[15] wl[205] vdd gnd cell_6t
Xbit_r206_c15 bl[15] br[15] wl[206] vdd gnd cell_6t
Xbit_r207_c15 bl[15] br[15] wl[207] vdd gnd cell_6t
Xbit_r208_c15 bl[15] br[15] wl[208] vdd gnd cell_6t
Xbit_r209_c15 bl[15] br[15] wl[209] vdd gnd cell_6t
Xbit_r210_c15 bl[15] br[15] wl[210] vdd gnd cell_6t
Xbit_r211_c15 bl[15] br[15] wl[211] vdd gnd cell_6t
Xbit_r212_c15 bl[15] br[15] wl[212] vdd gnd cell_6t
Xbit_r213_c15 bl[15] br[15] wl[213] vdd gnd cell_6t
Xbit_r214_c15 bl[15] br[15] wl[214] vdd gnd cell_6t
Xbit_r215_c15 bl[15] br[15] wl[215] vdd gnd cell_6t
Xbit_r216_c15 bl[15] br[15] wl[216] vdd gnd cell_6t
Xbit_r217_c15 bl[15] br[15] wl[217] vdd gnd cell_6t
Xbit_r218_c15 bl[15] br[15] wl[218] vdd gnd cell_6t
Xbit_r219_c15 bl[15] br[15] wl[219] vdd gnd cell_6t
Xbit_r220_c15 bl[15] br[15] wl[220] vdd gnd cell_6t
Xbit_r221_c15 bl[15] br[15] wl[221] vdd gnd cell_6t
Xbit_r222_c15 bl[15] br[15] wl[222] vdd gnd cell_6t
Xbit_r223_c15 bl[15] br[15] wl[223] vdd gnd cell_6t
Xbit_r224_c15 bl[15] br[15] wl[224] vdd gnd cell_6t
Xbit_r225_c15 bl[15] br[15] wl[225] vdd gnd cell_6t
Xbit_r226_c15 bl[15] br[15] wl[226] vdd gnd cell_6t
Xbit_r227_c15 bl[15] br[15] wl[227] vdd gnd cell_6t
Xbit_r228_c15 bl[15] br[15] wl[228] vdd gnd cell_6t
Xbit_r229_c15 bl[15] br[15] wl[229] vdd gnd cell_6t
Xbit_r230_c15 bl[15] br[15] wl[230] vdd gnd cell_6t
Xbit_r231_c15 bl[15] br[15] wl[231] vdd gnd cell_6t
Xbit_r232_c15 bl[15] br[15] wl[232] vdd gnd cell_6t
Xbit_r233_c15 bl[15] br[15] wl[233] vdd gnd cell_6t
Xbit_r234_c15 bl[15] br[15] wl[234] vdd gnd cell_6t
Xbit_r235_c15 bl[15] br[15] wl[235] vdd gnd cell_6t
Xbit_r236_c15 bl[15] br[15] wl[236] vdd gnd cell_6t
Xbit_r237_c15 bl[15] br[15] wl[237] vdd gnd cell_6t
Xbit_r238_c15 bl[15] br[15] wl[238] vdd gnd cell_6t
Xbit_r239_c15 bl[15] br[15] wl[239] vdd gnd cell_6t
Xbit_r240_c15 bl[15] br[15] wl[240] vdd gnd cell_6t
Xbit_r241_c15 bl[15] br[15] wl[241] vdd gnd cell_6t
Xbit_r242_c15 bl[15] br[15] wl[242] vdd gnd cell_6t
Xbit_r243_c15 bl[15] br[15] wl[243] vdd gnd cell_6t
Xbit_r244_c15 bl[15] br[15] wl[244] vdd gnd cell_6t
Xbit_r245_c15 bl[15] br[15] wl[245] vdd gnd cell_6t
Xbit_r246_c15 bl[15] br[15] wl[246] vdd gnd cell_6t
Xbit_r247_c15 bl[15] br[15] wl[247] vdd gnd cell_6t
Xbit_r248_c15 bl[15] br[15] wl[248] vdd gnd cell_6t
Xbit_r249_c15 bl[15] br[15] wl[249] vdd gnd cell_6t
Xbit_r250_c15 bl[15] br[15] wl[250] vdd gnd cell_6t
Xbit_r251_c15 bl[15] br[15] wl[251] vdd gnd cell_6t
Xbit_r252_c15 bl[15] br[15] wl[252] vdd gnd cell_6t
Xbit_r253_c15 bl[15] br[15] wl[253] vdd gnd cell_6t
Xbit_r254_c15 bl[15] br[15] wl[254] vdd gnd cell_6t
Xbit_r255_c15 bl[15] br[15] wl[255] vdd gnd cell_6t
Xbit_r0_c16 bl[16] br[16] wl[0] vdd gnd cell_6t
Xbit_r1_c16 bl[16] br[16] wl[1] vdd gnd cell_6t
Xbit_r2_c16 bl[16] br[16] wl[2] vdd gnd cell_6t
Xbit_r3_c16 bl[16] br[16] wl[3] vdd gnd cell_6t
Xbit_r4_c16 bl[16] br[16] wl[4] vdd gnd cell_6t
Xbit_r5_c16 bl[16] br[16] wl[5] vdd gnd cell_6t
Xbit_r6_c16 bl[16] br[16] wl[6] vdd gnd cell_6t
Xbit_r7_c16 bl[16] br[16] wl[7] vdd gnd cell_6t
Xbit_r8_c16 bl[16] br[16] wl[8] vdd gnd cell_6t
Xbit_r9_c16 bl[16] br[16] wl[9] vdd gnd cell_6t
Xbit_r10_c16 bl[16] br[16] wl[10] vdd gnd cell_6t
Xbit_r11_c16 bl[16] br[16] wl[11] vdd gnd cell_6t
Xbit_r12_c16 bl[16] br[16] wl[12] vdd gnd cell_6t
Xbit_r13_c16 bl[16] br[16] wl[13] vdd gnd cell_6t
Xbit_r14_c16 bl[16] br[16] wl[14] vdd gnd cell_6t
Xbit_r15_c16 bl[16] br[16] wl[15] vdd gnd cell_6t
Xbit_r16_c16 bl[16] br[16] wl[16] vdd gnd cell_6t
Xbit_r17_c16 bl[16] br[16] wl[17] vdd gnd cell_6t
Xbit_r18_c16 bl[16] br[16] wl[18] vdd gnd cell_6t
Xbit_r19_c16 bl[16] br[16] wl[19] vdd gnd cell_6t
Xbit_r20_c16 bl[16] br[16] wl[20] vdd gnd cell_6t
Xbit_r21_c16 bl[16] br[16] wl[21] vdd gnd cell_6t
Xbit_r22_c16 bl[16] br[16] wl[22] vdd gnd cell_6t
Xbit_r23_c16 bl[16] br[16] wl[23] vdd gnd cell_6t
Xbit_r24_c16 bl[16] br[16] wl[24] vdd gnd cell_6t
Xbit_r25_c16 bl[16] br[16] wl[25] vdd gnd cell_6t
Xbit_r26_c16 bl[16] br[16] wl[26] vdd gnd cell_6t
Xbit_r27_c16 bl[16] br[16] wl[27] vdd gnd cell_6t
Xbit_r28_c16 bl[16] br[16] wl[28] vdd gnd cell_6t
Xbit_r29_c16 bl[16] br[16] wl[29] vdd gnd cell_6t
Xbit_r30_c16 bl[16] br[16] wl[30] vdd gnd cell_6t
Xbit_r31_c16 bl[16] br[16] wl[31] vdd gnd cell_6t
Xbit_r32_c16 bl[16] br[16] wl[32] vdd gnd cell_6t
Xbit_r33_c16 bl[16] br[16] wl[33] vdd gnd cell_6t
Xbit_r34_c16 bl[16] br[16] wl[34] vdd gnd cell_6t
Xbit_r35_c16 bl[16] br[16] wl[35] vdd gnd cell_6t
Xbit_r36_c16 bl[16] br[16] wl[36] vdd gnd cell_6t
Xbit_r37_c16 bl[16] br[16] wl[37] vdd gnd cell_6t
Xbit_r38_c16 bl[16] br[16] wl[38] vdd gnd cell_6t
Xbit_r39_c16 bl[16] br[16] wl[39] vdd gnd cell_6t
Xbit_r40_c16 bl[16] br[16] wl[40] vdd gnd cell_6t
Xbit_r41_c16 bl[16] br[16] wl[41] vdd gnd cell_6t
Xbit_r42_c16 bl[16] br[16] wl[42] vdd gnd cell_6t
Xbit_r43_c16 bl[16] br[16] wl[43] vdd gnd cell_6t
Xbit_r44_c16 bl[16] br[16] wl[44] vdd gnd cell_6t
Xbit_r45_c16 bl[16] br[16] wl[45] vdd gnd cell_6t
Xbit_r46_c16 bl[16] br[16] wl[46] vdd gnd cell_6t
Xbit_r47_c16 bl[16] br[16] wl[47] vdd gnd cell_6t
Xbit_r48_c16 bl[16] br[16] wl[48] vdd gnd cell_6t
Xbit_r49_c16 bl[16] br[16] wl[49] vdd gnd cell_6t
Xbit_r50_c16 bl[16] br[16] wl[50] vdd gnd cell_6t
Xbit_r51_c16 bl[16] br[16] wl[51] vdd gnd cell_6t
Xbit_r52_c16 bl[16] br[16] wl[52] vdd gnd cell_6t
Xbit_r53_c16 bl[16] br[16] wl[53] vdd gnd cell_6t
Xbit_r54_c16 bl[16] br[16] wl[54] vdd gnd cell_6t
Xbit_r55_c16 bl[16] br[16] wl[55] vdd gnd cell_6t
Xbit_r56_c16 bl[16] br[16] wl[56] vdd gnd cell_6t
Xbit_r57_c16 bl[16] br[16] wl[57] vdd gnd cell_6t
Xbit_r58_c16 bl[16] br[16] wl[58] vdd gnd cell_6t
Xbit_r59_c16 bl[16] br[16] wl[59] vdd gnd cell_6t
Xbit_r60_c16 bl[16] br[16] wl[60] vdd gnd cell_6t
Xbit_r61_c16 bl[16] br[16] wl[61] vdd gnd cell_6t
Xbit_r62_c16 bl[16] br[16] wl[62] vdd gnd cell_6t
Xbit_r63_c16 bl[16] br[16] wl[63] vdd gnd cell_6t
Xbit_r64_c16 bl[16] br[16] wl[64] vdd gnd cell_6t
Xbit_r65_c16 bl[16] br[16] wl[65] vdd gnd cell_6t
Xbit_r66_c16 bl[16] br[16] wl[66] vdd gnd cell_6t
Xbit_r67_c16 bl[16] br[16] wl[67] vdd gnd cell_6t
Xbit_r68_c16 bl[16] br[16] wl[68] vdd gnd cell_6t
Xbit_r69_c16 bl[16] br[16] wl[69] vdd gnd cell_6t
Xbit_r70_c16 bl[16] br[16] wl[70] vdd gnd cell_6t
Xbit_r71_c16 bl[16] br[16] wl[71] vdd gnd cell_6t
Xbit_r72_c16 bl[16] br[16] wl[72] vdd gnd cell_6t
Xbit_r73_c16 bl[16] br[16] wl[73] vdd gnd cell_6t
Xbit_r74_c16 bl[16] br[16] wl[74] vdd gnd cell_6t
Xbit_r75_c16 bl[16] br[16] wl[75] vdd gnd cell_6t
Xbit_r76_c16 bl[16] br[16] wl[76] vdd gnd cell_6t
Xbit_r77_c16 bl[16] br[16] wl[77] vdd gnd cell_6t
Xbit_r78_c16 bl[16] br[16] wl[78] vdd gnd cell_6t
Xbit_r79_c16 bl[16] br[16] wl[79] vdd gnd cell_6t
Xbit_r80_c16 bl[16] br[16] wl[80] vdd gnd cell_6t
Xbit_r81_c16 bl[16] br[16] wl[81] vdd gnd cell_6t
Xbit_r82_c16 bl[16] br[16] wl[82] vdd gnd cell_6t
Xbit_r83_c16 bl[16] br[16] wl[83] vdd gnd cell_6t
Xbit_r84_c16 bl[16] br[16] wl[84] vdd gnd cell_6t
Xbit_r85_c16 bl[16] br[16] wl[85] vdd gnd cell_6t
Xbit_r86_c16 bl[16] br[16] wl[86] vdd gnd cell_6t
Xbit_r87_c16 bl[16] br[16] wl[87] vdd gnd cell_6t
Xbit_r88_c16 bl[16] br[16] wl[88] vdd gnd cell_6t
Xbit_r89_c16 bl[16] br[16] wl[89] vdd gnd cell_6t
Xbit_r90_c16 bl[16] br[16] wl[90] vdd gnd cell_6t
Xbit_r91_c16 bl[16] br[16] wl[91] vdd gnd cell_6t
Xbit_r92_c16 bl[16] br[16] wl[92] vdd gnd cell_6t
Xbit_r93_c16 bl[16] br[16] wl[93] vdd gnd cell_6t
Xbit_r94_c16 bl[16] br[16] wl[94] vdd gnd cell_6t
Xbit_r95_c16 bl[16] br[16] wl[95] vdd gnd cell_6t
Xbit_r96_c16 bl[16] br[16] wl[96] vdd gnd cell_6t
Xbit_r97_c16 bl[16] br[16] wl[97] vdd gnd cell_6t
Xbit_r98_c16 bl[16] br[16] wl[98] vdd gnd cell_6t
Xbit_r99_c16 bl[16] br[16] wl[99] vdd gnd cell_6t
Xbit_r100_c16 bl[16] br[16] wl[100] vdd gnd cell_6t
Xbit_r101_c16 bl[16] br[16] wl[101] vdd gnd cell_6t
Xbit_r102_c16 bl[16] br[16] wl[102] vdd gnd cell_6t
Xbit_r103_c16 bl[16] br[16] wl[103] vdd gnd cell_6t
Xbit_r104_c16 bl[16] br[16] wl[104] vdd gnd cell_6t
Xbit_r105_c16 bl[16] br[16] wl[105] vdd gnd cell_6t
Xbit_r106_c16 bl[16] br[16] wl[106] vdd gnd cell_6t
Xbit_r107_c16 bl[16] br[16] wl[107] vdd gnd cell_6t
Xbit_r108_c16 bl[16] br[16] wl[108] vdd gnd cell_6t
Xbit_r109_c16 bl[16] br[16] wl[109] vdd gnd cell_6t
Xbit_r110_c16 bl[16] br[16] wl[110] vdd gnd cell_6t
Xbit_r111_c16 bl[16] br[16] wl[111] vdd gnd cell_6t
Xbit_r112_c16 bl[16] br[16] wl[112] vdd gnd cell_6t
Xbit_r113_c16 bl[16] br[16] wl[113] vdd gnd cell_6t
Xbit_r114_c16 bl[16] br[16] wl[114] vdd gnd cell_6t
Xbit_r115_c16 bl[16] br[16] wl[115] vdd gnd cell_6t
Xbit_r116_c16 bl[16] br[16] wl[116] vdd gnd cell_6t
Xbit_r117_c16 bl[16] br[16] wl[117] vdd gnd cell_6t
Xbit_r118_c16 bl[16] br[16] wl[118] vdd gnd cell_6t
Xbit_r119_c16 bl[16] br[16] wl[119] vdd gnd cell_6t
Xbit_r120_c16 bl[16] br[16] wl[120] vdd gnd cell_6t
Xbit_r121_c16 bl[16] br[16] wl[121] vdd gnd cell_6t
Xbit_r122_c16 bl[16] br[16] wl[122] vdd gnd cell_6t
Xbit_r123_c16 bl[16] br[16] wl[123] vdd gnd cell_6t
Xbit_r124_c16 bl[16] br[16] wl[124] vdd gnd cell_6t
Xbit_r125_c16 bl[16] br[16] wl[125] vdd gnd cell_6t
Xbit_r126_c16 bl[16] br[16] wl[126] vdd gnd cell_6t
Xbit_r127_c16 bl[16] br[16] wl[127] vdd gnd cell_6t
Xbit_r128_c16 bl[16] br[16] wl[128] vdd gnd cell_6t
Xbit_r129_c16 bl[16] br[16] wl[129] vdd gnd cell_6t
Xbit_r130_c16 bl[16] br[16] wl[130] vdd gnd cell_6t
Xbit_r131_c16 bl[16] br[16] wl[131] vdd gnd cell_6t
Xbit_r132_c16 bl[16] br[16] wl[132] vdd gnd cell_6t
Xbit_r133_c16 bl[16] br[16] wl[133] vdd gnd cell_6t
Xbit_r134_c16 bl[16] br[16] wl[134] vdd gnd cell_6t
Xbit_r135_c16 bl[16] br[16] wl[135] vdd gnd cell_6t
Xbit_r136_c16 bl[16] br[16] wl[136] vdd gnd cell_6t
Xbit_r137_c16 bl[16] br[16] wl[137] vdd gnd cell_6t
Xbit_r138_c16 bl[16] br[16] wl[138] vdd gnd cell_6t
Xbit_r139_c16 bl[16] br[16] wl[139] vdd gnd cell_6t
Xbit_r140_c16 bl[16] br[16] wl[140] vdd gnd cell_6t
Xbit_r141_c16 bl[16] br[16] wl[141] vdd gnd cell_6t
Xbit_r142_c16 bl[16] br[16] wl[142] vdd gnd cell_6t
Xbit_r143_c16 bl[16] br[16] wl[143] vdd gnd cell_6t
Xbit_r144_c16 bl[16] br[16] wl[144] vdd gnd cell_6t
Xbit_r145_c16 bl[16] br[16] wl[145] vdd gnd cell_6t
Xbit_r146_c16 bl[16] br[16] wl[146] vdd gnd cell_6t
Xbit_r147_c16 bl[16] br[16] wl[147] vdd gnd cell_6t
Xbit_r148_c16 bl[16] br[16] wl[148] vdd gnd cell_6t
Xbit_r149_c16 bl[16] br[16] wl[149] vdd gnd cell_6t
Xbit_r150_c16 bl[16] br[16] wl[150] vdd gnd cell_6t
Xbit_r151_c16 bl[16] br[16] wl[151] vdd gnd cell_6t
Xbit_r152_c16 bl[16] br[16] wl[152] vdd gnd cell_6t
Xbit_r153_c16 bl[16] br[16] wl[153] vdd gnd cell_6t
Xbit_r154_c16 bl[16] br[16] wl[154] vdd gnd cell_6t
Xbit_r155_c16 bl[16] br[16] wl[155] vdd gnd cell_6t
Xbit_r156_c16 bl[16] br[16] wl[156] vdd gnd cell_6t
Xbit_r157_c16 bl[16] br[16] wl[157] vdd gnd cell_6t
Xbit_r158_c16 bl[16] br[16] wl[158] vdd gnd cell_6t
Xbit_r159_c16 bl[16] br[16] wl[159] vdd gnd cell_6t
Xbit_r160_c16 bl[16] br[16] wl[160] vdd gnd cell_6t
Xbit_r161_c16 bl[16] br[16] wl[161] vdd gnd cell_6t
Xbit_r162_c16 bl[16] br[16] wl[162] vdd gnd cell_6t
Xbit_r163_c16 bl[16] br[16] wl[163] vdd gnd cell_6t
Xbit_r164_c16 bl[16] br[16] wl[164] vdd gnd cell_6t
Xbit_r165_c16 bl[16] br[16] wl[165] vdd gnd cell_6t
Xbit_r166_c16 bl[16] br[16] wl[166] vdd gnd cell_6t
Xbit_r167_c16 bl[16] br[16] wl[167] vdd gnd cell_6t
Xbit_r168_c16 bl[16] br[16] wl[168] vdd gnd cell_6t
Xbit_r169_c16 bl[16] br[16] wl[169] vdd gnd cell_6t
Xbit_r170_c16 bl[16] br[16] wl[170] vdd gnd cell_6t
Xbit_r171_c16 bl[16] br[16] wl[171] vdd gnd cell_6t
Xbit_r172_c16 bl[16] br[16] wl[172] vdd gnd cell_6t
Xbit_r173_c16 bl[16] br[16] wl[173] vdd gnd cell_6t
Xbit_r174_c16 bl[16] br[16] wl[174] vdd gnd cell_6t
Xbit_r175_c16 bl[16] br[16] wl[175] vdd gnd cell_6t
Xbit_r176_c16 bl[16] br[16] wl[176] vdd gnd cell_6t
Xbit_r177_c16 bl[16] br[16] wl[177] vdd gnd cell_6t
Xbit_r178_c16 bl[16] br[16] wl[178] vdd gnd cell_6t
Xbit_r179_c16 bl[16] br[16] wl[179] vdd gnd cell_6t
Xbit_r180_c16 bl[16] br[16] wl[180] vdd gnd cell_6t
Xbit_r181_c16 bl[16] br[16] wl[181] vdd gnd cell_6t
Xbit_r182_c16 bl[16] br[16] wl[182] vdd gnd cell_6t
Xbit_r183_c16 bl[16] br[16] wl[183] vdd gnd cell_6t
Xbit_r184_c16 bl[16] br[16] wl[184] vdd gnd cell_6t
Xbit_r185_c16 bl[16] br[16] wl[185] vdd gnd cell_6t
Xbit_r186_c16 bl[16] br[16] wl[186] vdd gnd cell_6t
Xbit_r187_c16 bl[16] br[16] wl[187] vdd gnd cell_6t
Xbit_r188_c16 bl[16] br[16] wl[188] vdd gnd cell_6t
Xbit_r189_c16 bl[16] br[16] wl[189] vdd gnd cell_6t
Xbit_r190_c16 bl[16] br[16] wl[190] vdd gnd cell_6t
Xbit_r191_c16 bl[16] br[16] wl[191] vdd gnd cell_6t
Xbit_r192_c16 bl[16] br[16] wl[192] vdd gnd cell_6t
Xbit_r193_c16 bl[16] br[16] wl[193] vdd gnd cell_6t
Xbit_r194_c16 bl[16] br[16] wl[194] vdd gnd cell_6t
Xbit_r195_c16 bl[16] br[16] wl[195] vdd gnd cell_6t
Xbit_r196_c16 bl[16] br[16] wl[196] vdd gnd cell_6t
Xbit_r197_c16 bl[16] br[16] wl[197] vdd gnd cell_6t
Xbit_r198_c16 bl[16] br[16] wl[198] vdd gnd cell_6t
Xbit_r199_c16 bl[16] br[16] wl[199] vdd gnd cell_6t
Xbit_r200_c16 bl[16] br[16] wl[200] vdd gnd cell_6t
Xbit_r201_c16 bl[16] br[16] wl[201] vdd gnd cell_6t
Xbit_r202_c16 bl[16] br[16] wl[202] vdd gnd cell_6t
Xbit_r203_c16 bl[16] br[16] wl[203] vdd gnd cell_6t
Xbit_r204_c16 bl[16] br[16] wl[204] vdd gnd cell_6t
Xbit_r205_c16 bl[16] br[16] wl[205] vdd gnd cell_6t
Xbit_r206_c16 bl[16] br[16] wl[206] vdd gnd cell_6t
Xbit_r207_c16 bl[16] br[16] wl[207] vdd gnd cell_6t
Xbit_r208_c16 bl[16] br[16] wl[208] vdd gnd cell_6t
Xbit_r209_c16 bl[16] br[16] wl[209] vdd gnd cell_6t
Xbit_r210_c16 bl[16] br[16] wl[210] vdd gnd cell_6t
Xbit_r211_c16 bl[16] br[16] wl[211] vdd gnd cell_6t
Xbit_r212_c16 bl[16] br[16] wl[212] vdd gnd cell_6t
Xbit_r213_c16 bl[16] br[16] wl[213] vdd gnd cell_6t
Xbit_r214_c16 bl[16] br[16] wl[214] vdd gnd cell_6t
Xbit_r215_c16 bl[16] br[16] wl[215] vdd gnd cell_6t
Xbit_r216_c16 bl[16] br[16] wl[216] vdd gnd cell_6t
Xbit_r217_c16 bl[16] br[16] wl[217] vdd gnd cell_6t
Xbit_r218_c16 bl[16] br[16] wl[218] vdd gnd cell_6t
Xbit_r219_c16 bl[16] br[16] wl[219] vdd gnd cell_6t
Xbit_r220_c16 bl[16] br[16] wl[220] vdd gnd cell_6t
Xbit_r221_c16 bl[16] br[16] wl[221] vdd gnd cell_6t
Xbit_r222_c16 bl[16] br[16] wl[222] vdd gnd cell_6t
Xbit_r223_c16 bl[16] br[16] wl[223] vdd gnd cell_6t
Xbit_r224_c16 bl[16] br[16] wl[224] vdd gnd cell_6t
Xbit_r225_c16 bl[16] br[16] wl[225] vdd gnd cell_6t
Xbit_r226_c16 bl[16] br[16] wl[226] vdd gnd cell_6t
Xbit_r227_c16 bl[16] br[16] wl[227] vdd gnd cell_6t
Xbit_r228_c16 bl[16] br[16] wl[228] vdd gnd cell_6t
Xbit_r229_c16 bl[16] br[16] wl[229] vdd gnd cell_6t
Xbit_r230_c16 bl[16] br[16] wl[230] vdd gnd cell_6t
Xbit_r231_c16 bl[16] br[16] wl[231] vdd gnd cell_6t
Xbit_r232_c16 bl[16] br[16] wl[232] vdd gnd cell_6t
Xbit_r233_c16 bl[16] br[16] wl[233] vdd gnd cell_6t
Xbit_r234_c16 bl[16] br[16] wl[234] vdd gnd cell_6t
Xbit_r235_c16 bl[16] br[16] wl[235] vdd gnd cell_6t
Xbit_r236_c16 bl[16] br[16] wl[236] vdd gnd cell_6t
Xbit_r237_c16 bl[16] br[16] wl[237] vdd gnd cell_6t
Xbit_r238_c16 bl[16] br[16] wl[238] vdd gnd cell_6t
Xbit_r239_c16 bl[16] br[16] wl[239] vdd gnd cell_6t
Xbit_r240_c16 bl[16] br[16] wl[240] vdd gnd cell_6t
Xbit_r241_c16 bl[16] br[16] wl[241] vdd gnd cell_6t
Xbit_r242_c16 bl[16] br[16] wl[242] vdd gnd cell_6t
Xbit_r243_c16 bl[16] br[16] wl[243] vdd gnd cell_6t
Xbit_r244_c16 bl[16] br[16] wl[244] vdd gnd cell_6t
Xbit_r245_c16 bl[16] br[16] wl[245] vdd gnd cell_6t
Xbit_r246_c16 bl[16] br[16] wl[246] vdd gnd cell_6t
Xbit_r247_c16 bl[16] br[16] wl[247] vdd gnd cell_6t
Xbit_r248_c16 bl[16] br[16] wl[248] vdd gnd cell_6t
Xbit_r249_c16 bl[16] br[16] wl[249] vdd gnd cell_6t
Xbit_r250_c16 bl[16] br[16] wl[250] vdd gnd cell_6t
Xbit_r251_c16 bl[16] br[16] wl[251] vdd gnd cell_6t
Xbit_r252_c16 bl[16] br[16] wl[252] vdd gnd cell_6t
Xbit_r253_c16 bl[16] br[16] wl[253] vdd gnd cell_6t
Xbit_r254_c16 bl[16] br[16] wl[254] vdd gnd cell_6t
Xbit_r255_c16 bl[16] br[16] wl[255] vdd gnd cell_6t
Xbit_r0_c17 bl[17] br[17] wl[0] vdd gnd cell_6t
Xbit_r1_c17 bl[17] br[17] wl[1] vdd gnd cell_6t
Xbit_r2_c17 bl[17] br[17] wl[2] vdd gnd cell_6t
Xbit_r3_c17 bl[17] br[17] wl[3] vdd gnd cell_6t
Xbit_r4_c17 bl[17] br[17] wl[4] vdd gnd cell_6t
Xbit_r5_c17 bl[17] br[17] wl[5] vdd gnd cell_6t
Xbit_r6_c17 bl[17] br[17] wl[6] vdd gnd cell_6t
Xbit_r7_c17 bl[17] br[17] wl[7] vdd gnd cell_6t
Xbit_r8_c17 bl[17] br[17] wl[8] vdd gnd cell_6t
Xbit_r9_c17 bl[17] br[17] wl[9] vdd gnd cell_6t
Xbit_r10_c17 bl[17] br[17] wl[10] vdd gnd cell_6t
Xbit_r11_c17 bl[17] br[17] wl[11] vdd gnd cell_6t
Xbit_r12_c17 bl[17] br[17] wl[12] vdd gnd cell_6t
Xbit_r13_c17 bl[17] br[17] wl[13] vdd gnd cell_6t
Xbit_r14_c17 bl[17] br[17] wl[14] vdd gnd cell_6t
Xbit_r15_c17 bl[17] br[17] wl[15] vdd gnd cell_6t
Xbit_r16_c17 bl[17] br[17] wl[16] vdd gnd cell_6t
Xbit_r17_c17 bl[17] br[17] wl[17] vdd gnd cell_6t
Xbit_r18_c17 bl[17] br[17] wl[18] vdd gnd cell_6t
Xbit_r19_c17 bl[17] br[17] wl[19] vdd gnd cell_6t
Xbit_r20_c17 bl[17] br[17] wl[20] vdd gnd cell_6t
Xbit_r21_c17 bl[17] br[17] wl[21] vdd gnd cell_6t
Xbit_r22_c17 bl[17] br[17] wl[22] vdd gnd cell_6t
Xbit_r23_c17 bl[17] br[17] wl[23] vdd gnd cell_6t
Xbit_r24_c17 bl[17] br[17] wl[24] vdd gnd cell_6t
Xbit_r25_c17 bl[17] br[17] wl[25] vdd gnd cell_6t
Xbit_r26_c17 bl[17] br[17] wl[26] vdd gnd cell_6t
Xbit_r27_c17 bl[17] br[17] wl[27] vdd gnd cell_6t
Xbit_r28_c17 bl[17] br[17] wl[28] vdd gnd cell_6t
Xbit_r29_c17 bl[17] br[17] wl[29] vdd gnd cell_6t
Xbit_r30_c17 bl[17] br[17] wl[30] vdd gnd cell_6t
Xbit_r31_c17 bl[17] br[17] wl[31] vdd gnd cell_6t
Xbit_r32_c17 bl[17] br[17] wl[32] vdd gnd cell_6t
Xbit_r33_c17 bl[17] br[17] wl[33] vdd gnd cell_6t
Xbit_r34_c17 bl[17] br[17] wl[34] vdd gnd cell_6t
Xbit_r35_c17 bl[17] br[17] wl[35] vdd gnd cell_6t
Xbit_r36_c17 bl[17] br[17] wl[36] vdd gnd cell_6t
Xbit_r37_c17 bl[17] br[17] wl[37] vdd gnd cell_6t
Xbit_r38_c17 bl[17] br[17] wl[38] vdd gnd cell_6t
Xbit_r39_c17 bl[17] br[17] wl[39] vdd gnd cell_6t
Xbit_r40_c17 bl[17] br[17] wl[40] vdd gnd cell_6t
Xbit_r41_c17 bl[17] br[17] wl[41] vdd gnd cell_6t
Xbit_r42_c17 bl[17] br[17] wl[42] vdd gnd cell_6t
Xbit_r43_c17 bl[17] br[17] wl[43] vdd gnd cell_6t
Xbit_r44_c17 bl[17] br[17] wl[44] vdd gnd cell_6t
Xbit_r45_c17 bl[17] br[17] wl[45] vdd gnd cell_6t
Xbit_r46_c17 bl[17] br[17] wl[46] vdd gnd cell_6t
Xbit_r47_c17 bl[17] br[17] wl[47] vdd gnd cell_6t
Xbit_r48_c17 bl[17] br[17] wl[48] vdd gnd cell_6t
Xbit_r49_c17 bl[17] br[17] wl[49] vdd gnd cell_6t
Xbit_r50_c17 bl[17] br[17] wl[50] vdd gnd cell_6t
Xbit_r51_c17 bl[17] br[17] wl[51] vdd gnd cell_6t
Xbit_r52_c17 bl[17] br[17] wl[52] vdd gnd cell_6t
Xbit_r53_c17 bl[17] br[17] wl[53] vdd gnd cell_6t
Xbit_r54_c17 bl[17] br[17] wl[54] vdd gnd cell_6t
Xbit_r55_c17 bl[17] br[17] wl[55] vdd gnd cell_6t
Xbit_r56_c17 bl[17] br[17] wl[56] vdd gnd cell_6t
Xbit_r57_c17 bl[17] br[17] wl[57] vdd gnd cell_6t
Xbit_r58_c17 bl[17] br[17] wl[58] vdd gnd cell_6t
Xbit_r59_c17 bl[17] br[17] wl[59] vdd gnd cell_6t
Xbit_r60_c17 bl[17] br[17] wl[60] vdd gnd cell_6t
Xbit_r61_c17 bl[17] br[17] wl[61] vdd gnd cell_6t
Xbit_r62_c17 bl[17] br[17] wl[62] vdd gnd cell_6t
Xbit_r63_c17 bl[17] br[17] wl[63] vdd gnd cell_6t
Xbit_r64_c17 bl[17] br[17] wl[64] vdd gnd cell_6t
Xbit_r65_c17 bl[17] br[17] wl[65] vdd gnd cell_6t
Xbit_r66_c17 bl[17] br[17] wl[66] vdd gnd cell_6t
Xbit_r67_c17 bl[17] br[17] wl[67] vdd gnd cell_6t
Xbit_r68_c17 bl[17] br[17] wl[68] vdd gnd cell_6t
Xbit_r69_c17 bl[17] br[17] wl[69] vdd gnd cell_6t
Xbit_r70_c17 bl[17] br[17] wl[70] vdd gnd cell_6t
Xbit_r71_c17 bl[17] br[17] wl[71] vdd gnd cell_6t
Xbit_r72_c17 bl[17] br[17] wl[72] vdd gnd cell_6t
Xbit_r73_c17 bl[17] br[17] wl[73] vdd gnd cell_6t
Xbit_r74_c17 bl[17] br[17] wl[74] vdd gnd cell_6t
Xbit_r75_c17 bl[17] br[17] wl[75] vdd gnd cell_6t
Xbit_r76_c17 bl[17] br[17] wl[76] vdd gnd cell_6t
Xbit_r77_c17 bl[17] br[17] wl[77] vdd gnd cell_6t
Xbit_r78_c17 bl[17] br[17] wl[78] vdd gnd cell_6t
Xbit_r79_c17 bl[17] br[17] wl[79] vdd gnd cell_6t
Xbit_r80_c17 bl[17] br[17] wl[80] vdd gnd cell_6t
Xbit_r81_c17 bl[17] br[17] wl[81] vdd gnd cell_6t
Xbit_r82_c17 bl[17] br[17] wl[82] vdd gnd cell_6t
Xbit_r83_c17 bl[17] br[17] wl[83] vdd gnd cell_6t
Xbit_r84_c17 bl[17] br[17] wl[84] vdd gnd cell_6t
Xbit_r85_c17 bl[17] br[17] wl[85] vdd gnd cell_6t
Xbit_r86_c17 bl[17] br[17] wl[86] vdd gnd cell_6t
Xbit_r87_c17 bl[17] br[17] wl[87] vdd gnd cell_6t
Xbit_r88_c17 bl[17] br[17] wl[88] vdd gnd cell_6t
Xbit_r89_c17 bl[17] br[17] wl[89] vdd gnd cell_6t
Xbit_r90_c17 bl[17] br[17] wl[90] vdd gnd cell_6t
Xbit_r91_c17 bl[17] br[17] wl[91] vdd gnd cell_6t
Xbit_r92_c17 bl[17] br[17] wl[92] vdd gnd cell_6t
Xbit_r93_c17 bl[17] br[17] wl[93] vdd gnd cell_6t
Xbit_r94_c17 bl[17] br[17] wl[94] vdd gnd cell_6t
Xbit_r95_c17 bl[17] br[17] wl[95] vdd gnd cell_6t
Xbit_r96_c17 bl[17] br[17] wl[96] vdd gnd cell_6t
Xbit_r97_c17 bl[17] br[17] wl[97] vdd gnd cell_6t
Xbit_r98_c17 bl[17] br[17] wl[98] vdd gnd cell_6t
Xbit_r99_c17 bl[17] br[17] wl[99] vdd gnd cell_6t
Xbit_r100_c17 bl[17] br[17] wl[100] vdd gnd cell_6t
Xbit_r101_c17 bl[17] br[17] wl[101] vdd gnd cell_6t
Xbit_r102_c17 bl[17] br[17] wl[102] vdd gnd cell_6t
Xbit_r103_c17 bl[17] br[17] wl[103] vdd gnd cell_6t
Xbit_r104_c17 bl[17] br[17] wl[104] vdd gnd cell_6t
Xbit_r105_c17 bl[17] br[17] wl[105] vdd gnd cell_6t
Xbit_r106_c17 bl[17] br[17] wl[106] vdd gnd cell_6t
Xbit_r107_c17 bl[17] br[17] wl[107] vdd gnd cell_6t
Xbit_r108_c17 bl[17] br[17] wl[108] vdd gnd cell_6t
Xbit_r109_c17 bl[17] br[17] wl[109] vdd gnd cell_6t
Xbit_r110_c17 bl[17] br[17] wl[110] vdd gnd cell_6t
Xbit_r111_c17 bl[17] br[17] wl[111] vdd gnd cell_6t
Xbit_r112_c17 bl[17] br[17] wl[112] vdd gnd cell_6t
Xbit_r113_c17 bl[17] br[17] wl[113] vdd gnd cell_6t
Xbit_r114_c17 bl[17] br[17] wl[114] vdd gnd cell_6t
Xbit_r115_c17 bl[17] br[17] wl[115] vdd gnd cell_6t
Xbit_r116_c17 bl[17] br[17] wl[116] vdd gnd cell_6t
Xbit_r117_c17 bl[17] br[17] wl[117] vdd gnd cell_6t
Xbit_r118_c17 bl[17] br[17] wl[118] vdd gnd cell_6t
Xbit_r119_c17 bl[17] br[17] wl[119] vdd gnd cell_6t
Xbit_r120_c17 bl[17] br[17] wl[120] vdd gnd cell_6t
Xbit_r121_c17 bl[17] br[17] wl[121] vdd gnd cell_6t
Xbit_r122_c17 bl[17] br[17] wl[122] vdd gnd cell_6t
Xbit_r123_c17 bl[17] br[17] wl[123] vdd gnd cell_6t
Xbit_r124_c17 bl[17] br[17] wl[124] vdd gnd cell_6t
Xbit_r125_c17 bl[17] br[17] wl[125] vdd gnd cell_6t
Xbit_r126_c17 bl[17] br[17] wl[126] vdd gnd cell_6t
Xbit_r127_c17 bl[17] br[17] wl[127] vdd gnd cell_6t
Xbit_r128_c17 bl[17] br[17] wl[128] vdd gnd cell_6t
Xbit_r129_c17 bl[17] br[17] wl[129] vdd gnd cell_6t
Xbit_r130_c17 bl[17] br[17] wl[130] vdd gnd cell_6t
Xbit_r131_c17 bl[17] br[17] wl[131] vdd gnd cell_6t
Xbit_r132_c17 bl[17] br[17] wl[132] vdd gnd cell_6t
Xbit_r133_c17 bl[17] br[17] wl[133] vdd gnd cell_6t
Xbit_r134_c17 bl[17] br[17] wl[134] vdd gnd cell_6t
Xbit_r135_c17 bl[17] br[17] wl[135] vdd gnd cell_6t
Xbit_r136_c17 bl[17] br[17] wl[136] vdd gnd cell_6t
Xbit_r137_c17 bl[17] br[17] wl[137] vdd gnd cell_6t
Xbit_r138_c17 bl[17] br[17] wl[138] vdd gnd cell_6t
Xbit_r139_c17 bl[17] br[17] wl[139] vdd gnd cell_6t
Xbit_r140_c17 bl[17] br[17] wl[140] vdd gnd cell_6t
Xbit_r141_c17 bl[17] br[17] wl[141] vdd gnd cell_6t
Xbit_r142_c17 bl[17] br[17] wl[142] vdd gnd cell_6t
Xbit_r143_c17 bl[17] br[17] wl[143] vdd gnd cell_6t
Xbit_r144_c17 bl[17] br[17] wl[144] vdd gnd cell_6t
Xbit_r145_c17 bl[17] br[17] wl[145] vdd gnd cell_6t
Xbit_r146_c17 bl[17] br[17] wl[146] vdd gnd cell_6t
Xbit_r147_c17 bl[17] br[17] wl[147] vdd gnd cell_6t
Xbit_r148_c17 bl[17] br[17] wl[148] vdd gnd cell_6t
Xbit_r149_c17 bl[17] br[17] wl[149] vdd gnd cell_6t
Xbit_r150_c17 bl[17] br[17] wl[150] vdd gnd cell_6t
Xbit_r151_c17 bl[17] br[17] wl[151] vdd gnd cell_6t
Xbit_r152_c17 bl[17] br[17] wl[152] vdd gnd cell_6t
Xbit_r153_c17 bl[17] br[17] wl[153] vdd gnd cell_6t
Xbit_r154_c17 bl[17] br[17] wl[154] vdd gnd cell_6t
Xbit_r155_c17 bl[17] br[17] wl[155] vdd gnd cell_6t
Xbit_r156_c17 bl[17] br[17] wl[156] vdd gnd cell_6t
Xbit_r157_c17 bl[17] br[17] wl[157] vdd gnd cell_6t
Xbit_r158_c17 bl[17] br[17] wl[158] vdd gnd cell_6t
Xbit_r159_c17 bl[17] br[17] wl[159] vdd gnd cell_6t
Xbit_r160_c17 bl[17] br[17] wl[160] vdd gnd cell_6t
Xbit_r161_c17 bl[17] br[17] wl[161] vdd gnd cell_6t
Xbit_r162_c17 bl[17] br[17] wl[162] vdd gnd cell_6t
Xbit_r163_c17 bl[17] br[17] wl[163] vdd gnd cell_6t
Xbit_r164_c17 bl[17] br[17] wl[164] vdd gnd cell_6t
Xbit_r165_c17 bl[17] br[17] wl[165] vdd gnd cell_6t
Xbit_r166_c17 bl[17] br[17] wl[166] vdd gnd cell_6t
Xbit_r167_c17 bl[17] br[17] wl[167] vdd gnd cell_6t
Xbit_r168_c17 bl[17] br[17] wl[168] vdd gnd cell_6t
Xbit_r169_c17 bl[17] br[17] wl[169] vdd gnd cell_6t
Xbit_r170_c17 bl[17] br[17] wl[170] vdd gnd cell_6t
Xbit_r171_c17 bl[17] br[17] wl[171] vdd gnd cell_6t
Xbit_r172_c17 bl[17] br[17] wl[172] vdd gnd cell_6t
Xbit_r173_c17 bl[17] br[17] wl[173] vdd gnd cell_6t
Xbit_r174_c17 bl[17] br[17] wl[174] vdd gnd cell_6t
Xbit_r175_c17 bl[17] br[17] wl[175] vdd gnd cell_6t
Xbit_r176_c17 bl[17] br[17] wl[176] vdd gnd cell_6t
Xbit_r177_c17 bl[17] br[17] wl[177] vdd gnd cell_6t
Xbit_r178_c17 bl[17] br[17] wl[178] vdd gnd cell_6t
Xbit_r179_c17 bl[17] br[17] wl[179] vdd gnd cell_6t
Xbit_r180_c17 bl[17] br[17] wl[180] vdd gnd cell_6t
Xbit_r181_c17 bl[17] br[17] wl[181] vdd gnd cell_6t
Xbit_r182_c17 bl[17] br[17] wl[182] vdd gnd cell_6t
Xbit_r183_c17 bl[17] br[17] wl[183] vdd gnd cell_6t
Xbit_r184_c17 bl[17] br[17] wl[184] vdd gnd cell_6t
Xbit_r185_c17 bl[17] br[17] wl[185] vdd gnd cell_6t
Xbit_r186_c17 bl[17] br[17] wl[186] vdd gnd cell_6t
Xbit_r187_c17 bl[17] br[17] wl[187] vdd gnd cell_6t
Xbit_r188_c17 bl[17] br[17] wl[188] vdd gnd cell_6t
Xbit_r189_c17 bl[17] br[17] wl[189] vdd gnd cell_6t
Xbit_r190_c17 bl[17] br[17] wl[190] vdd gnd cell_6t
Xbit_r191_c17 bl[17] br[17] wl[191] vdd gnd cell_6t
Xbit_r192_c17 bl[17] br[17] wl[192] vdd gnd cell_6t
Xbit_r193_c17 bl[17] br[17] wl[193] vdd gnd cell_6t
Xbit_r194_c17 bl[17] br[17] wl[194] vdd gnd cell_6t
Xbit_r195_c17 bl[17] br[17] wl[195] vdd gnd cell_6t
Xbit_r196_c17 bl[17] br[17] wl[196] vdd gnd cell_6t
Xbit_r197_c17 bl[17] br[17] wl[197] vdd gnd cell_6t
Xbit_r198_c17 bl[17] br[17] wl[198] vdd gnd cell_6t
Xbit_r199_c17 bl[17] br[17] wl[199] vdd gnd cell_6t
Xbit_r200_c17 bl[17] br[17] wl[200] vdd gnd cell_6t
Xbit_r201_c17 bl[17] br[17] wl[201] vdd gnd cell_6t
Xbit_r202_c17 bl[17] br[17] wl[202] vdd gnd cell_6t
Xbit_r203_c17 bl[17] br[17] wl[203] vdd gnd cell_6t
Xbit_r204_c17 bl[17] br[17] wl[204] vdd gnd cell_6t
Xbit_r205_c17 bl[17] br[17] wl[205] vdd gnd cell_6t
Xbit_r206_c17 bl[17] br[17] wl[206] vdd gnd cell_6t
Xbit_r207_c17 bl[17] br[17] wl[207] vdd gnd cell_6t
Xbit_r208_c17 bl[17] br[17] wl[208] vdd gnd cell_6t
Xbit_r209_c17 bl[17] br[17] wl[209] vdd gnd cell_6t
Xbit_r210_c17 bl[17] br[17] wl[210] vdd gnd cell_6t
Xbit_r211_c17 bl[17] br[17] wl[211] vdd gnd cell_6t
Xbit_r212_c17 bl[17] br[17] wl[212] vdd gnd cell_6t
Xbit_r213_c17 bl[17] br[17] wl[213] vdd gnd cell_6t
Xbit_r214_c17 bl[17] br[17] wl[214] vdd gnd cell_6t
Xbit_r215_c17 bl[17] br[17] wl[215] vdd gnd cell_6t
Xbit_r216_c17 bl[17] br[17] wl[216] vdd gnd cell_6t
Xbit_r217_c17 bl[17] br[17] wl[217] vdd gnd cell_6t
Xbit_r218_c17 bl[17] br[17] wl[218] vdd gnd cell_6t
Xbit_r219_c17 bl[17] br[17] wl[219] vdd gnd cell_6t
Xbit_r220_c17 bl[17] br[17] wl[220] vdd gnd cell_6t
Xbit_r221_c17 bl[17] br[17] wl[221] vdd gnd cell_6t
Xbit_r222_c17 bl[17] br[17] wl[222] vdd gnd cell_6t
Xbit_r223_c17 bl[17] br[17] wl[223] vdd gnd cell_6t
Xbit_r224_c17 bl[17] br[17] wl[224] vdd gnd cell_6t
Xbit_r225_c17 bl[17] br[17] wl[225] vdd gnd cell_6t
Xbit_r226_c17 bl[17] br[17] wl[226] vdd gnd cell_6t
Xbit_r227_c17 bl[17] br[17] wl[227] vdd gnd cell_6t
Xbit_r228_c17 bl[17] br[17] wl[228] vdd gnd cell_6t
Xbit_r229_c17 bl[17] br[17] wl[229] vdd gnd cell_6t
Xbit_r230_c17 bl[17] br[17] wl[230] vdd gnd cell_6t
Xbit_r231_c17 bl[17] br[17] wl[231] vdd gnd cell_6t
Xbit_r232_c17 bl[17] br[17] wl[232] vdd gnd cell_6t
Xbit_r233_c17 bl[17] br[17] wl[233] vdd gnd cell_6t
Xbit_r234_c17 bl[17] br[17] wl[234] vdd gnd cell_6t
Xbit_r235_c17 bl[17] br[17] wl[235] vdd gnd cell_6t
Xbit_r236_c17 bl[17] br[17] wl[236] vdd gnd cell_6t
Xbit_r237_c17 bl[17] br[17] wl[237] vdd gnd cell_6t
Xbit_r238_c17 bl[17] br[17] wl[238] vdd gnd cell_6t
Xbit_r239_c17 bl[17] br[17] wl[239] vdd gnd cell_6t
Xbit_r240_c17 bl[17] br[17] wl[240] vdd gnd cell_6t
Xbit_r241_c17 bl[17] br[17] wl[241] vdd gnd cell_6t
Xbit_r242_c17 bl[17] br[17] wl[242] vdd gnd cell_6t
Xbit_r243_c17 bl[17] br[17] wl[243] vdd gnd cell_6t
Xbit_r244_c17 bl[17] br[17] wl[244] vdd gnd cell_6t
Xbit_r245_c17 bl[17] br[17] wl[245] vdd gnd cell_6t
Xbit_r246_c17 bl[17] br[17] wl[246] vdd gnd cell_6t
Xbit_r247_c17 bl[17] br[17] wl[247] vdd gnd cell_6t
Xbit_r248_c17 bl[17] br[17] wl[248] vdd gnd cell_6t
Xbit_r249_c17 bl[17] br[17] wl[249] vdd gnd cell_6t
Xbit_r250_c17 bl[17] br[17] wl[250] vdd gnd cell_6t
Xbit_r251_c17 bl[17] br[17] wl[251] vdd gnd cell_6t
Xbit_r252_c17 bl[17] br[17] wl[252] vdd gnd cell_6t
Xbit_r253_c17 bl[17] br[17] wl[253] vdd gnd cell_6t
Xbit_r254_c17 bl[17] br[17] wl[254] vdd gnd cell_6t
Xbit_r255_c17 bl[17] br[17] wl[255] vdd gnd cell_6t
Xbit_r0_c18 bl[18] br[18] wl[0] vdd gnd cell_6t
Xbit_r1_c18 bl[18] br[18] wl[1] vdd gnd cell_6t
Xbit_r2_c18 bl[18] br[18] wl[2] vdd gnd cell_6t
Xbit_r3_c18 bl[18] br[18] wl[3] vdd gnd cell_6t
Xbit_r4_c18 bl[18] br[18] wl[4] vdd gnd cell_6t
Xbit_r5_c18 bl[18] br[18] wl[5] vdd gnd cell_6t
Xbit_r6_c18 bl[18] br[18] wl[6] vdd gnd cell_6t
Xbit_r7_c18 bl[18] br[18] wl[7] vdd gnd cell_6t
Xbit_r8_c18 bl[18] br[18] wl[8] vdd gnd cell_6t
Xbit_r9_c18 bl[18] br[18] wl[9] vdd gnd cell_6t
Xbit_r10_c18 bl[18] br[18] wl[10] vdd gnd cell_6t
Xbit_r11_c18 bl[18] br[18] wl[11] vdd gnd cell_6t
Xbit_r12_c18 bl[18] br[18] wl[12] vdd gnd cell_6t
Xbit_r13_c18 bl[18] br[18] wl[13] vdd gnd cell_6t
Xbit_r14_c18 bl[18] br[18] wl[14] vdd gnd cell_6t
Xbit_r15_c18 bl[18] br[18] wl[15] vdd gnd cell_6t
Xbit_r16_c18 bl[18] br[18] wl[16] vdd gnd cell_6t
Xbit_r17_c18 bl[18] br[18] wl[17] vdd gnd cell_6t
Xbit_r18_c18 bl[18] br[18] wl[18] vdd gnd cell_6t
Xbit_r19_c18 bl[18] br[18] wl[19] vdd gnd cell_6t
Xbit_r20_c18 bl[18] br[18] wl[20] vdd gnd cell_6t
Xbit_r21_c18 bl[18] br[18] wl[21] vdd gnd cell_6t
Xbit_r22_c18 bl[18] br[18] wl[22] vdd gnd cell_6t
Xbit_r23_c18 bl[18] br[18] wl[23] vdd gnd cell_6t
Xbit_r24_c18 bl[18] br[18] wl[24] vdd gnd cell_6t
Xbit_r25_c18 bl[18] br[18] wl[25] vdd gnd cell_6t
Xbit_r26_c18 bl[18] br[18] wl[26] vdd gnd cell_6t
Xbit_r27_c18 bl[18] br[18] wl[27] vdd gnd cell_6t
Xbit_r28_c18 bl[18] br[18] wl[28] vdd gnd cell_6t
Xbit_r29_c18 bl[18] br[18] wl[29] vdd gnd cell_6t
Xbit_r30_c18 bl[18] br[18] wl[30] vdd gnd cell_6t
Xbit_r31_c18 bl[18] br[18] wl[31] vdd gnd cell_6t
Xbit_r32_c18 bl[18] br[18] wl[32] vdd gnd cell_6t
Xbit_r33_c18 bl[18] br[18] wl[33] vdd gnd cell_6t
Xbit_r34_c18 bl[18] br[18] wl[34] vdd gnd cell_6t
Xbit_r35_c18 bl[18] br[18] wl[35] vdd gnd cell_6t
Xbit_r36_c18 bl[18] br[18] wl[36] vdd gnd cell_6t
Xbit_r37_c18 bl[18] br[18] wl[37] vdd gnd cell_6t
Xbit_r38_c18 bl[18] br[18] wl[38] vdd gnd cell_6t
Xbit_r39_c18 bl[18] br[18] wl[39] vdd gnd cell_6t
Xbit_r40_c18 bl[18] br[18] wl[40] vdd gnd cell_6t
Xbit_r41_c18 bl[18] br[18] wl[41] vdd gnd cell_6t
Xbit_r42_c18 bl[18] br[18] wl[42] vdd gnd cell_6t
Xbit_r43_c18 bl[18] br[18] wl[43] vdd gnd cell_6t
Xbit_r44_c18 bl[18] br[18] wl[44] vdd gnd cell_6t
Xbit_r45_c18 bl[18] br[18] wl[45] vdd gnd cell_6t
Xbit_r46_c18 bl[18] br[18] wl[46] vdd gnd cell_6t
Xbit_r47_c18 bl[18] br[18] wl[47] vdd gnd cell_6t
Xbit_r48_c18 bl[18] br[18] wl[48] vdd gnd cell_6t
Xbit_r49_c18 bl[18] br[18] wl[49] vdd gnd cell_6t
Xbit_r50_c18 bl[18] br[18] wl[50] vdd gnd cell_6t
Xbit_r51_c18 bl[18] br[18] wl[51] vdd gnd cell_6t
Xbit_r52_c18 bl[18] br[18] wl[52] vdd gnd cell_6t
Xbit_r53_c18 bl[18] br[18] wl[53] vdd gnd cell_6t
Xbit_r54_c18 bl[18] br[18] wl[54] vdd gnd cell_6t
Xbit_r55_c18 bl[18] br[18] wl[55] vdd gnd cell_6t
Xbit_r56_c18 bl[18] br[18] wl[56] vdd gnd cell_6t
Xbit_r57_c18 bl[18] br[18] wl[57] vdd gnd cell_6t
Xbit_r58_c18 bl[18] br[18] wl[58] vdd gnd cell_6t
Xbit_r59_c18 bl[18] br[18] wl[59] vdd gnd cell_6t
Xbit_r60_c18 bl[18] br[18] wl[60] vdd gnd cell_6t
Xbit_r61_c18 bl[18] br[18] wl[61] vdd gnd cell_6t
Xbit_r62_c18 bl[18] br[18] wl[62] vdd gnd cell_6t
Xbit_r63_c18 bl[18] br[18] wl[63] vdd gnd cell_6t
Xbit_r64_c18 bl[18] br[18] wl[64] vdd gnd cell_6t
Xbit_r65_c18 bl[18] br[18] wl[65] vdd gnd cell_6t
Xbit_r66_c18 bl[18] br[18] wl[66] vdd gnd cell_6t
Xbit_r67_c18 bl[18] br[18] wl[67] vdd gnd cell_6t
Xbit_r68_c18 bl[18] br[18] wl[68] vdd gnd cell_6t
Xbit_r69_c18 bl[18] br[18] wl[69] vdd gnd cell_6t
Xbit_r70_c18 bl[18] br[18] wl[70] vdd gnd cell_6t
Xbit_r71_c18 bl[18] br[18] wl[71] vdd gnd cell_6t
Xbit_r72_c18 bl[18] br[18] wl[72] vdd gnd cell_6t
Xbit_r73_c18 bl[18] br[18] wl[73] vdd gnd cell_6t
Xbit_r74_c18 bl[18] br[18] wl[74] vdd gnd cell_6t
Xbit_r75_c18 bl[18] br[18] wl[75] vdd gnd cell_6t
Xbit_r76_c18 bl[18] br[18] wl[76] vdd gnd cell_6t
Xbit_r77_c18 bl[18] br[18] wl[77] vdd gnd cell_6t
Xbit_r78_c18 bl[18] br[18] wl[78] vdd gnd cell_6t
Xbit_r79_c18 bl[18] br[18] wl[79] vdd gnd cell_6t
Xbit_r80_c18 bl[18] br[18] wl[80] vdd gnd cell_6t
Xbit_r81_c18 bl[18] br[18] wl[81] vdd gnd cell_6t
Xbit_r82_c18 bl[18] br[18] wl[82] vdd gnd cell_6t
Xbit_r83_c18 bl[18] br[18] wl[83] vdd gnd cell_6t
Xbit_r84_c18 bl[18] br[18] wl[84] vdd gnd cell_6t
Xbit_r85_c18 bl[18] br[18] wl[85] vdd gnd cell_6t
Xbit_r86_c18 bl[18] br[18] wl[86] vdd gnd cell_6t
Xbit_r87_c18 bl[18] br[18] wl[87] vdd gnd cell_6t
Xbit_r88_c18 bl[18] br[18] wl[88] vdd gnd cell_6t
Xbit_r89_c18 bl[18] br[18] wl[89] vdd gnd cell_6t
Xbit_r90_c18 bl[18] br[18] wl[90] vdd gnd cell_6t
Xbit_r91_c18 bl[18] br[18] wl[91] vdd gnd cell_6t
Xbit_r92_c18 bl[18] br[18] wl[92] vdd gnd cell_6t
Xbit_r93_c18 bl[18] br[18] wl[93] vdd gnd cell_6t
Xbit_r94_c18 bl[18] br[18] wl[94] vdd gnd cell_6t
Xbit_r95_c18 bl[18] br[18] wl[95] vdd gnd cell_6t
Xbit_r96_c18 bl[18] br[18] wl[96] vdd gnd cell_6t
Xbit_r97_c18 bl[18] br[18] wl[97] vdd gnd cell_6t
Xbit_r98_c18 bl[18] br[18] wl[98] vdd gnd cell_6t
Xbit_r99_c18 bl[18] br[18] wl[99] vdd gnd cell_6t
Xbit_r100_c18 bl[18] br[18] wl[100] vdd gnd cell_6t
Xbit_r101_c18 bl[18] br[18] wl[101] vdd gnd cell_6t
Xbit_r102_c18 bl[18] br[18] wl[102] vdd gnd cell_6t
Xbit_r103_c18 bl[18] br[18] wl[103] vdd gnd cell_6t
Xbit_r104_c18 bl[18] br[18] wl[104] vdd gnd cell_6t
Xbit_r105_c18 bl[18] br[18] wl[105] vdd gnd cell_6t
Xbit_r106_c18 bl[18] br[18] wl[106] vdd gnd cell_6t
Xbit_r107_c18 bl[18] br[18] wl[107] vdd gnd cell_6t
Xbit_r108_c18 bl[18] br[18] wl[108] vdd gnd cell_6t
Xbit_r109_c18 bl[18] br[18] wl[109] vdd gnd cell_6t
Xbit_r110_c18 bl[18] br[18] wl[110] vdd gnd cell_6t
Xbit_r111_c18 bl[18] br[18] wl[111] vdd gnd cell_6t
Xbit_r112_c18 bl[18] br[18] wl[112] vdd gnd cell_6t
Xbit_r113_c18 bl[18] br[18] wl[113] vdd gnd cell_6t
Xbit_r114_c18 bl[18] br[18] wl[114] vdd gnd cell_6t
Xbit_r115_c18 bl[18] br[18] wl[115] vdd gnd cell_6t
Xbit_r116_c18 bl[18] br[18] wl[116] vdd gnd cell_6t
Xbit_r117_c18 bl[18] br[18] wl[117] vdd gnd cell_6t
Xbit_r118_c18 bl[18] br[18] wl[118] vdd gnd cell_6t
Xbit_r119_c18 bl[18] br[18] wl[119] vdd gnd cell_6t
Xbit_r120_c18 bl[18] br[18] wl[120] vdd gnd cell_6t
Xbit_r121_c18 bl[18] br[18] wl[121] vdd gnd cell_6t
Xbit_r122_c18 bl[18] br[18] wl[122] vdd gnd cell_6t
Xbit_r123_c18 bl[18] br[18] wl[123] vdd gnd cell_6t
Xbit_r124_c18 bl[18] br[18] wl[124] vdd gnd cell_6t
Xbit_r125_c18 bl[18] br[18] wl[125] vdd gnd cell_6t
Xbit_r126_c18 bl[18] br[18] wl[126] vdd gnd cell_6t
Xbit_r127_c18 bl[18] br[18] wl[127] vdd gnd cell_6t
Xbit_r128_c18 bl[18] br[18] wl[128] vdd gnd cell_6t
Xbit_r129_c18 bl[18] br[18] wl[129] vdd gnd cell_6t
Xbit_r130_c18 bl[18] br[18] wl[130] vdd gnd cell_6t
Xbit_r131_c18 bl[18] br[18] wl[131] vdd gnd cell_6t
Xbit_r132_c18 bl[18] br[18] wl[132] vdd gnd cell_6t
Xbit_r133_c18 bl[18] br[18] wl[133] vdd gnd cell_6t
Xbit_r134_c18 bl[18] br[18] wl[134] vdd gnd cell_6t
Xbit_r135_c18 bl[18] br[18] wl[135] vdd gnd cell_6t
Xbit_r136_c18 bl[18] br[18] wl[136] vdd gnd cell_6t
Xbit_r137_c18 bl[18] br[18] wl[137] vdd gnd cell_6t
Xbit_r138_c18 bl[18] br[18] wl[138] vdd gnd cell_6t
Xbit_r139_c18 bl[18] br[18] wl[139] vdd gnd cell_6t
Xbit_r140_c18 bl[18] br[18] wl[140] vdd gnd cell_6t
Xbit_r141_c18 bl[18] br[18] wl[141] vdd gnd cell_6t
Xbit_r142_c18 bl[18] br[18] wl[142] vdd gnd cell_6t
Xbit_r143_c18 bl[18] br[18] wl[143] vdd gnd cell_6t
Xbit_r144_c18 bl[18] br[18] wl[144] vdd gnd cell_6t
Xbit_r145_c18 bl[18] br[18] wl[145] vdd gnd cell_6t
Xbit_r146_c18 bl[18] br[18] wl[146] vdd gnd cell_6t
Xbit_r147_c18 bl[18] br[18] wl[147] vdd gnd cell_6t
Xbit_r148_c18 bl[18] br[18] wl[148] vdd gnd cell_6t
Xbit_r149_c18 bl[18] br[18] wl[149] vdd gnd cell_6t
Xbit_r150_c18 bl[18] br[18] wl[150] vdd gnd cell_6t
Xbit_r151_c18 bl[18] br[18] wl[151] vdd gnd cell_6t
Xbit_r152_c18 bl[18] br[18] wl[152] vdd gnd cell_6t
Xbit_r153_c18 bl[18] br[18] wl[153] vdd gnd cell_6t
Xbit_r154_c18 bl[18] br[18] wl[154] vdd gnd cell_6t
Xbit_r155_c18 bl[18] br[18] wl[155] vdd gnd cell_6t
Xbit_r156_c18 bl[18] br[18] wl[156] vdd gnd cell_6t
Xbit_r157_c18 bl[18] br[18] wl[157] vdd gnd cell_6t
Xbit_r158_c18 bl[18] br[18] wl[158] vdd gnd cell_6t
Xbit_r159_c18 bl[18] br[18] wl[159] vdd gnd cell_6t
Xbit_r160_c18 bl[18] br[18] wl[160] vdd gnd cell_6t
Xbit_r161_c18 bl[18] br[18] wl[161] vdd gnd cell_6t
Xbit_r162_c18 bl[18] br[18] wl[162] vdd gnd cell_6t
Xbit_r163_c18 bl[18] br[18] wl[163] vdd gnd cell_6t
Xbit_r164_c18 bl[18] br[18] wl[164] vdd gnd cell_6t
Xbit_r165_c18 bl[18] br[18] wl[165] vdd gnd cell_6t
Xbit_r166_c18 bl[18] br[18] wl[166] vdd gnd cell_6t
Xbit_r167_c18 bl[18] br[18] wl[167] vdd gnd cell_6t
Xbit_r168_c18 bl[18] br[18] wl[168] vdd gnd cell_6t
Xbit_r169_c18 bl[18] br[18] wl[169] vdd gnd cell_6t
Xbit_r170_c18 bl[18] br[18] wl[170] vdd gnd cell_6t
Xbit_r171_c18 bl[18] br[18] wl[171] vdd gnd cell_6t
Xbit_r172_c18 bl[18] br[18] wl[172] vdd gnd cell_6t
Xbit_r173_c18 bl[18] br[18] wl[173] vdd gnd cell_6t
Xbit_r174_c18 bl[18] br[18] wl[174] vdd gnd cell_6t
Xbit_r175_c18 bl[18] br[18] wl[175] vdd gnd cell_6t
Xbit_r176_c18 bl[18] br[18] wl[176] vdd gnd cell_6t
Xbit_r177_c18 bl[18] br[18] wl[177] vdd gnd cell_6t
Xbit_r178_c18 bl[18] br[18] wl[178] vdd gnd cell_6t
Xbit_r179_c18 bl[18] br[18] wl[179] vdd gnd cell_6t
Xbit_r180_c18 bl[18] br[18] wl[180] vdd gnd cell_6t
Xbit_r181_c18 bl[18] br[18] wl[181] vdd gnd cell_6t
Xbit_r182_c18 bl[18] br[18] wl[182] vdd gnd cell_6t
Xbit_r183_c18 bl[18] br[18] wl[183] vdd gnd cell_6t
Xbit_r184_c18 bl[18] br[18] wl[184] vdd gnd cell_6t
Xbit_r185_c18 bl[18] br[18] wl[185] vdd gnd cell_6t
Xbit_r186_c18 bl[18] br[18] wl[186] vdd gnd cell_6t
Xbit_r187_c18 bl[18] br[18] wl[187] vdd gnd cell_6t
Xbit_r188_c18 bl[18] br[18] wl[188] vdd gnd cell_6t
Xbit_r189_c18 bl[18] br[18] wl[189] vdd gnd cell_6t
Xbit_r190_c18 bl[18] br[18] wl[190] vdd gnd cell_6t
Xbit_r191_c18 bl[18] br[18] wl[191] vdd gnd cell_6t
Xbit_r192_c18 bl[18] br[18] wl[192] vdd gnd cell_6t
Xbit_r193_c18 bl[18] br[18] wl[193] vdd gnd cell_6t
Xbit_r194_c18 bl[18] br[18] wl[194] vdd gnd cell_6t
Xbit_r195_c18 bl[18] br[18] wl[195] vdd gnd cell_6t
Xbit_r196_c18 bl[18] br[18] wl[196] vdd gnd cell_6t
Xbit_r197_c18 bl[18] br[18] wl[197] vdd gnd cell_6t
Xbit_r198_c18 bl[18] br[18] wl[198] vdd gnd cell_6t
Xbit_r199_c18 bl[18] br[18] wl[199] vdd gnd cell_6t
Xbit_r200_c18 bl[18] br[18] wl[200] vdd gnd cell_6t
Xbit_r201_c18 bl[18] br[18] wl[201] vdd gnd cell_6t
Xbit_r202_c18 bl[18] br[18] wl[202] vdd gnd cell_6t
Xbit_r203_c18 bl[18] br[18] wl[203] vdd gnd cell_6t
Xbit_r204_c18 bl[18] br[18] wl[204] vdd gnd cell_6t
Xbit_r205_c18 bl[18] br[18] wl[205] vdd gnd cell_6t
Xbit_r206_c18 bl[18] br[18] wl[206] vdd gnd cell_6t
Xbit_r207_c18 bl[18] br[18] wl[207] vdd gnd cell_6t
Xbit_r208_c18 bl[18] br[18] wl[208] vdd gnd cell_6t
Xbit_r209_c18 bl[18] br[18] wl[209] vdd gnd cell_6t
Xbit_r210_c18 bl[18] br[18] wl[210] vdd gnd cell_6t
Xbit_r211_c18 bl[18] br[18] wl[211] vdd gnd cell_6t
Xbit_r212_c18 bl[18] br[18] wl[212] vdd gnd cell_6t
Xbit_r213_c18 bl[18] br[18] wl[213] vdd gnd cell_6t
Xbit_r214_c18 bl[18] br[18] wl[214] vdd gnd cell_6t
Xbit_r215_c18 bl[18] br[18] wl[215] vdd gnd cell_6t
Xbit_r216_c18 bl[18] br[18] wl[216] vdd gnd cell_6t
Xbit_r217_c18 bl[18] br[18] wl[217] vdd gnd cell_6t
Xbit_r218_c18 bl[18] br[18] wl[218] vdd gnd cell_6t
Xbit_r219_c18 bl[18] br[18] wl[219] vdd gnd cell_6t
Xbit_r220_c18 bl[18] br[18] wl[220] vdd gnd cell_6t
Xbit_r221_c18 bl[18] br[18] wl[221] vdd gnd cell_6t
Xbit_r222_c18 bl[18] br[18] wl[222] vdd gnd cell_6t
Xbit_r223_c18 bl[18] br[18] wl[223] vdd gnd cell_6t
Xbit_r224_c18 bl[18] br[18] wl[224] vdd gnd cell_6t
Xbit_r225_c18 bl[18] br[18] wl[225] vdd gnd cell_6t
Xbit_r226_c18 bl[18] br[18] wl[226] vdd gnd cell_6t
Xbit_r227_c18 bl[18] br[18] wl[227] vdd gnd cell_6t
Xbit_r228_c18 bl[18] br[18] wl[228] vdd gnd cell_6t
Xbit_r229_c18 bl[18] br[18] wl[229] vdd gnd cell_6t
Xbit_r230_c18 bl[18] br[18] wl[230] vdd gnd cell_6t
Xbit_r231_c18 bl[18] br[18] wl[231] vdd gnd cell_6t
Xbit_r232_c18 bl[18] br[18] wl[232] vdd gnd cell_6t
Xbit_r233_c18 bl[18] br[18] wl[233] vdd gnd cell_6t
Xbit_r234_c18 bl[18] br[18] wl[234] vdd gnd cell_6t
Xbit_r235_c18 bl[18] br[18] wl[235] vdd gnd cell_6t
Xbit_r236_c18 bl[18] br[18] wl[236] vdd gnd cell_6t
Xbit_r237_c18 bl[18] br[18] wl[237] vdd gnd cell_6t
Xbit_r238_c18 bl[18] br[18] wl[238] vdd gnd cell_6t
Xbit_r239_c18 bl[18] br[18] wl[239] vdd gnd cell_6t
Xbit_r240_c18 bl[18] br[18] wl[240] vdd gnd cell_6t
Xbit_r241_c18 bl[18] br[18] wl[241] vdd gnd cell_6t
Xbit_r242_c18 bl[18] br[18] wl[242] vdd gnd cell_6t
Xbit_r243_c18 bl[18] br[18] wl[243] vdd gnd cell_6t
Xbit_r244_c18 bl[18] br[18] wl[244] vdd gnd cell_6t
Xbit_r245_c18 bl[18] br[18] wl[245] vdd gnd cell_6t
Xbit_r246_c18 bl[18] br[18] wl[246] vdd gnd cell_6t
Xbit_r247_c18 bl[18] br[18] wl[247] vdd gnd cell_6t
Xbit_r248_c18 bl[18] br[18] wl[248] vdd gnd cell_6t
Xbit_r249_c18 bl[18] br[18] wl[249] vdd gnd cell_6t
Xbit_r250_c18 bl[18] br[18] wl[250] vdd gnd cell_6t
Xbit_r251_c18 bl[18] br[18] wl[251] vdd gnd cell_6t
Xbit_r252_c18 bl[18] br[18] wl[252] vdd gnd cell_6t
Xbit_r253_c18 bl[18] br[18] wl[253] vdd gnd cell_6t
Xbit_r254_c18 bl[18] br[18] wl[254] vdd gnd cell_6t
Xbit_r255_c18 bl[18] br[18] wl[255] vdd gnd cell_6t
Xbit_r0_c19 bl[19] br[19] wl[0] vdd gnd cell_6t
Xbit_r1_c19 bl[19] br[19] wl[1] vdd gnd cell_6t
Xbit_r2_c19 bl[19] br[19] wl[2] vdd gnd cell_6t
Xbit_r3_c19 bl[19] br[19] wl[3] vdd gnd cell_6t
Xbit_r4_c19 bl[19] br[19] wl[4] vdd gnd cell_6t
Xbit_r5_c19 bl[19] br[19] wl[5] vdd gnd cell_6t
Xbit_r6_c19 bl[19] br[19] wl[6] vdd gnd cell_6t
Xbit_r7_c19 bl[19] br[19] wl[7] vdd gnd cell_6t
Xbit_r8_c19 bl[19] br[19] wl[8] vdd gnd cell_6t
Xbit_r9_c19 bl[19] br[19] wl[9] vdd gnd cell_6t
Xbit_r10_c19 bl[19] br[19] wl[10] vdd gnd cell_6t
Xbit_r11_c19 bl[19] br[19] wl[11] vdd gnd cell_6t
Xbit_r12_c19 bl[19] br[19] wl[12] vdd gnd cell_6t
Xbit_r13_c19 bl[19] br[19] wl[13] vdd gnd cell_6t
Xbit_r14_c19 bl[19] br[19] wl[14] vdd gnd cell_6t
Xbit_r15_c19 bl[19] br[19] wl[15] vdd gnd cell_6t
Xbit_r16_c19 bl[19] br[19] wl[16] vdd gnd cell_6t
Xbit_r17_c19 bl[19] br[19] wl[17] vdd gnd cell_6t
Xbit_r18_c19 bl[19] br[19] wl[18] vdd gnd cell_6t
Xbit_r19_c19 bl[19] br[19] wl[19] vdd gnd cell_6t
Xbit_r20_c19 bl[19] br[19] wl[20] vdd gnd cell_6t
Xbit_r21_c19 bl[19] br[19] wl[21] vdd gnd cell_6t
Xbit_r22_c19 bl[19] br[19] wl[22] vdd gnd cell_6t
Xbit_r23_c19 bl[19] br[19] wl[23] vdd gnd cell_6t
Xbit_r24_c19 bl[19] br[19] wl[24] vdd gnd cell_6t
Xbit_r25_c19 bl[19] br[19] wl[25] vdd gnd cell_6t
Xbit_r26_c19 bl[19] br[19] wl[26] vdd gnd cell_6t
Xbit_r27_c19 bl[19] br[19] wl[27] vdd gnd cell_6t
Xbit_r28_c19 bl[19] br[19] wl[28] vdd gnd cell_6t
Xbit_r29_c19 bl[19] br[19] wl[29] vdd gnd cell_6t
Xbit_r30_c19 bl[19] br[19] wl[30] vdd gnd cell_6t
Xbit_r31_c19 bl[19] br[19] wl[31] vdd gnd cell_6t
Xbit_r32_c19 bl[19] br[19] wl[32] vdd gnd cell_6t
Xbit_r33_c19 bl[19] br[19] wl[33] vdd gnd cell_6t
Xbit_r34_c19 bl[19] br[19] wl[34] vdd gnd cell_6t
Xbit_r35_c19 bl[19] br[19] wl[35] vdd gnd cell_6t
Xbit_r36_c19 bl[19] br[19] wl[36] vdd gnd cell_6t
Xbit_r37_c19 bl[19] br[19] wl[37] vdd gnd cell_6t
Xbit_r38_c19 bl[19] br[19] wl[38] vdd gnd cell_6t
Xbit_r39_c19 bl[19] br[19] wl[39] vdd gnd cell_6t
Xbit_r40_c19 bl[19] br[19] wl[40] vdd gnd cell_6t
Xbit_r41_c19 bl[19] br[19] wl[41] vdd gnd cell_6t
Xbit_r42_c19 bl[19] br[19] wl[42] vdd gnd cell_6t
Xbit_r43_c19 bl[19] br[19] wl[43] vdd gnd cell_6t
Xbit_r44_c19 bl[19] br[19] wl[44] vdd gnd cell_6t
Xbit_r45_c19 bl[19] br[19] wl[45] vdd gnd cell_6t
Xbit_r46_c19 bl[19] br[19] wl[46] vdd gnd cell_6t
Xbit_r47_c19 bl[19] br[19] wl[47] vdd gnd cell_6t
Xbit_r48_c19 bl[19] br[19] wl[48] vdd gnd cell_6t
Xbit_r49_c19 bl[19] br[19] wl[49] vdd gnd cell_6t
Xbit_r50_c19 bl[19] br[19] wl[50] vdd gnd cell_6t
Xbit_r51_c19 bl[19] br[19] wl[51] vdd gnd cell_6t
Xbit_r52_c19 bl[19] br[19] wl[52] vdd gnd cell_6t
Xbit_r53_c19 bl[19] br[19] wl[53] vdd gnd cell_6t
Xbit_r54_c19 bl[19] br[19] wl[54] vdd gnd cell_6t
Xbit_r55_c19 bl[19] br[19] wl[55] vdd gnd cell_6t
Xbit_r56_c19 bl[19] br[19] wl[56] vdd gnd cell_6t
Xbit_r57_c19 bl[19] br[19] wl[57] vdd gnd cell_6t
Xbit_r58_c19 bl[19] br[19] wl[58] vdd gnd cell_6t
Xbit_r59_c19 bl[19] br[19] wl[59] vdd gnd cell_6t
Xbit_r60_c19 bl[19] br[19] wl[60] vdd gnd cell_6t
Xbit_r61_c19 bl[19] br[19] wl[61] vdd gnd cell_6t
Xbit_r62_c19 bl[19] br[19] wl[62] vdd gnd cell_6t
Xbit_r63_c19 bl[19] br[19] wl[63] vdd gnd cell_6t
Xbit_r64_c19 bl[19] br[19] wl[64] vdd gnd cell_6t
Xbit_r65_c19 bl[19] br[19] wl[65] vdd gnd cell_6t
Xbit_r66_c19 bl[19] br[19] wl[66] vdd gnd cell_6t
Xbit_r67_c19 bl[19] br[19] wl[67] vdd gnd cell_6t
Xbit_r68_c19 bl[19] br[19] wl[68] vdd gnd cell_6t
Xbit_r69_c19 bl[19] br[19] wl[69] vdd gnd cell_6t
Xbit_r70_c19 bl[19] br[19] wl[70] vdd gnd cell_6t
Xbit_r71_c19 bl[19] br[19] wl[71] vdd gnd cell_6t
Xbit_r72_c19 bl[19] br[19] wl[72] vdd gnd cell_6t
Xbit_r73_c19 bl[19] br[19] wl[73] vdd gnd cell_6t
Xbit_r74_c19 bl[19] br[19] wl[74] vdd gnd cell_6t
Xbit_r75_c19 bl[19] br[19] wl[75] vdd gnd cell_6t
Xbit_r76_c19 bl[19] br[19] wl[76] vdd gnd cell_6t
Xbit_r77_c19 bl[19] br[19] wl[77] vdd gnd cell_6t
Xbit_r78_c19 bl[19] br[19] wl[78] vdd gnd cell_6t
Xbit_r79_c19 bl[19] br[19] wl[79] vdd gnd cell_6t
Xbit_r80_c19 bl[19] br[19] wl[80] vdd gnd cell_6t
Xbit_r81_c19 bl[19] br[19] wl[81] vdd gnd cell_6t
Xbit_r82_c19 bl[19] br[19] wl[82] vdd gnd cell_6t
Xbit_r83_c19 bl[19] br[19] wl[83] vdd gnd cell_6t
Xbit_r84_c19 bl[19] br[19] wl[84] vdd gnd cell_6t
Xbit_r85_c19 bl[19] br[19] wl[85] vdd gnd cell_6t
Xbit_r86_c19 bl[19] br[19] wl[86] vdd gnd cell_6t
Xbit_r87_c19 bl[19] br[19] wl[87] vdd gnd cell_6t
Xbit_r88_c19 bl[19] br[19] wl[88] vdd gnd cell_6t
Xbit_r89_c19 bl[19] br[19] wl[89] vdd gnd cell_6t
Xbit_r90_c19 bl[19] br[19] wl[90] vdd gnd cell_6t
Xbit_r91_c19 bl[19] br[19] wl[91] vdd gnd cell_6t
Xbit_r92_c19 bl[19] br[19] wl[92] vdd gnd cell_6t
Xbit_r93_c19 bl[19] br[19] wl[93] vdd gnd cell_6t
Xbit_r94_c19 bl[19] br[19] wl[94] vdd gnd cell_6t
Xbit_r95_c19 bl[19] br[19] wl[95] vdd gnd cell_6t
Xbit_r96_c19 bl[19] br[19] wl[96] vdd gnd cell_6t
Xbit_r97_c19 bl[19] br[19] wl[97] vdd gnd cell_6t
Xbit_r98_c19 bl[19] br[19] wl[98] vdd gnd cell_6t
Xbit_r99_c19 bl[19] br[19] wl[99] vdd gnd cell_6t
Xbit_r100_c19 bl[19] br[19] wl[100] vdd gnd cell_6t
Xbit_r101_c19 bl[19] br[19] wl[101] vdd gnd cell_6t
Xbit_r102_c19 bl[19] br[19] wl[102] vdd gnd cell_6t
Xbit_r103_c19 bl[19] br[19] wl[103] vdd gnd cell_6t
Xbit_r104_c19 bl[19] br[19] wl[104] vdd gnd cell_6t
Xbit_r105_c19 bl[19] br[19] wl[105] vdd gnd cell_6t
Xbit_r106_c19 bl[19] br[19] wl[106] vdd gnd cell_6t
Xbit_r107_c19 bl[19] br[19] wl[107] vdd gnd cell_6t
Xbit_r108_c19 bl[19] br[19] wl[108] vdd gnd cell_6t
Xbit_r109_c19 bl[19] br[19] wl[109] vdd gnd cell_6t
Xbit_r110_c19 bl[19] br[19] wl[110] vdd gnd cell_6t
Xbit_r111_c19 bl[19] br[19] wl[111] vdd gnd cell_6t
Xbit_r112_c19 bl[19] br[19] wl[112] vdd gnd cell_6t
Xbit_r113_c19 bl[19] br[19] wl[113] vdd gnd cell_6t
Xbit_r114_c19 bl[19] br[19] wl[114] vdd gnd cell_6t
Xbit_r115_c19 bl[19] br[19] wl[115] vdd gnd cell_6t
Xbit_r116_c19 bl[19] br[19] wl[116] vdd gnd cell_6t
Xbit_r117_c19 bl[19] br[19] wl[117] vdd gnd cell_6t
Xbit_r118_c19 bl[19] br[19] wl[118] vdd gnd cell_6t
Xbit_r119_c19 bl[19] br[19] wl[119] vdd gnd cell_6t
Xbit_r120_c19 bl[19] br[19] wl[120] vdd gnd cell_6t
Xbit_r121_c19 bl[19] br[19] wl[121] vdd gnd cell_6t
Xbit_r122_c19 bl[19] br[19] wl[122] vdd gnd cell_6t
Xbit_r123_c19 bl[19] br[19] wl[123] vdd gnd cell_6t
Xbit_r124_c19 bl[19] br[19] wl[124] vdd gnd cell_6t
Xbit_r125_c19 bl[19] br[19] wl[125] vdd gnd cell_6t
Xbit_r126_c19 bl[19] br[19] wl[126] vdd gnd cell_6t
Xbit_r127_c19 bl[19] br[19] wl[127] vdd gnd cell_6t
Xbit_r128_c19 bl[19] br[19] wl[128] vdd gnd cell_6t
Xbit_r129_c19 bl[19] br[19] wl[129] vdd gnd cell_6t
Xbit_r130_c19 bl[19] br[19] wl[130] vdd gnd cell_6t
Xbit_r131_c19 bl[19] br[19] wl[131] vdd gnd cell_6t
Xbit_r132_c19 bl[19] br[19] wl[132] vdd gnd cell_6t
Xbit_r133_c19 bl[19] br[19] wl[133] vdd gnd cell_6t
Xbit_r134_c19 bl[19] br[19] wl[134] vdd gnd cell_6t
Xbit_r135_c19 bl[19] br[19] wl[135] vdd gnd cell_6t
Xbit_r136_c19 bl[19] br[19] wl[136] vdd gnd cell_6t
Xbit_r137_c19 bl[19] br[19] wl[137] vdd gnd cell_6t
Xbit_r138_c19 bl[19] br[19] wl[138] vdd gnd cell_6t
Xbit_r139_c19 bl[19] br[19] wl[139] vdd gnd cell_6t
Xbit_r140_c19 bl[19] br[19] wl[140] vdd gnd cell_6t
Xbit_r141_c19 bl[19] br[19] wl[141] vdd gnd cell_6t
Xbit_r142_c19 bl[19] br[19] wl[142] vdd gnd cell_6t
Xbit_r143_c19 bl[19] br[19] wl[143] vdd gnd cell_6t
Xbit_r144_c19 bl[19] br[19] wl[144] vdd gnd cell_6t
Xbit_r145_c19 bl[19] br[19] wl[145] vdd gnd cell_6t
Xbit_r146_c19 bl[19] br[19] wl[146] vdd gnd cell_6t
Xbit_r147_c19 bl[19] br[19] wl[147] vdd gnd cell_6t
Xbit_r148_c19 bl[19] br[19] wl[148] vdd gnd cell_6t
Xbit_r149_c19 bl[19] br[19] wl[149] vdd gnd cell_6t
Xbit_r150_c19 bl[19] br[19] wl[150] vdd gnd cell_6t
Xbit_r151_c19 bl[19] br[19] wl[151] vdd gnd cell_6t
Xbit_r152_c19 bl[19] br[19] wl[152] vdd gnd cell_6t
Xbit_r153_c19 bl[19] br[19] wl[153] vdd gnd cell_6t
Xbit_r154_c19 bl[19] br[19] wl[154] vdd gnd cell_6t
Xbit_r155_c19 bl[19] br[19] wl[155] vdd gnd cell_6t
Xbit_r156_c19 bl[19] br[19] wl[156] vdd gnd cell_6t
Xbit_r157_c19 bl[19] br[19] wl[157] vdd gnd cell_6t
Xbit_r158_c19 bl[19] br[19] wl[158] vdd gnd cell_6t
Xbit_r159_c19 bl[19] br[19] wl[159] vdd gnd cell_6t
Xbit_r160_c19 bl[19] br[19] wl[160] vdd gnd cell_6t
Xbit_r161_c19 bl[19] br[19] wl[161] vdd gnd cell_6t
Xbit_r162_c19 bl[19] br[19] wl[162] vdd gnd cell_6t
Xbit_r163_c19 bl[19] br[19] wl[163] vdd gnd cell_6t
Xbit_r164_c19 bl[19] br[19] wl[164] vdd gnd cell_6t
Xbit_r165_c19 bl[19] br[19] wl[165] vdd gnd cell_6t
Xbit_r166_c19 bl[19] br[19] wl[166] vdd gnd cell_6t
Xbit_r167_c19 bl[19] br[19] wl[167] vdd gnd cell_6t
Xbit_r168_c19 bl[19] br[19] wl[168] vdd gnd cell_6t
Xbit_r169_c19 bl[19] br[19] wl[169] vdd gnd cell_6t
Xbit_r170_c19 bl[19] br[19] wl[170] vdd gnd cell_6t
Xbit_r171_c19 bl[19] br[19] wl[171] vdd gnd cell_6t
Xbit_r172_c19 bl[19] br[19] wl[172] vdd gnd cell_6t
Xbit_r173_c19 bl[19] br[19] wl[173] vdd gnd cell_6t
Xbit_r174_c19 bl[19] br[19] wl[174] vdd gnd cell_6t
Xbit_r175_c19 bl[19] br[19] wl[175] vdd gnd cell_6t
Xbit_r176_c19 bl[19] br[19] wl[176] vdd gnd cell_6t
Xbit_r177_c19 bl[19] br[19] wl[177] vdd gnd cell_6t
Xbit_r178_c19 bl[19] br[19] wl[178] vdd gnd cell_6t
Xbit_r179_c19 bl[19] br[19] wl[179] vdd gnd cell_6t
Xbit_r180_c19 bl[19] br[19] wl[180] vdd gnd cell_6t
Xbit_r181_c19 bl[19] br[19] wl[181] vdd gnd cell_6t
Xbit_r182_c19 bl[19] br[19] wl[182] vdd gnd cell_6t
Xbit_r183_c19 bl[19] br[19] wl[183] vdd gnd cell_6t
Xbit_r184_c19 bl[19] br[19] wl[184] vdd gnd cell_6t
Xbit_r185_c19 bl[19] br[19] wl[185] vdd gnd cell_6t
Xbit_r186_c19 bl[19] br[19] wl[186] vdd gnd cell_6t
Xbit_r187_c19 bl[19] br[19] wl[187] vdd gnd cell_6t
Xbit_r188_c19 bl[19] br[19] wl[188] vdd gnd cell_6t
Xbit_r189_c19 bl[19] br[19] wl[189] vdd gnd cell_6t
Xbit_r190_c19 bl[19] br[19] wl[190] vdd gnd cell_6t
Xbit_r191_c19 bl[19] br[19] wl[191] vdd gnd cell_6t
Xbit_r192_c19 bl[19] br[19] wl[192] vdd gnd cell_6t
Xbit_r193_c19 bl[19] br[19] wl[193] vdd gnd cell_6t
Xbit_r194_c19 bl[19] br[19] wl[194] vdd gnd cell_6t
Xbit_r195_c19 bl[19] br[19] wl[195] vdd gnd cell_6t
Xbit_r196_c19 bl[19] br[19] wl[196] vdd gnd cell_6t
Xbit_r197_c19 bl[19] br[19] wl[197] vdd gnd cell_6t
Xbit_r198_c19 bl[19] br[19] wl[198] vdd gnd cell_6t
Xbit_r199_c19 bl[19] br[19] wl[199] vdd gnd cell_6t
Xbit_r200_c19 bl[19] br[19] wl[200] vdd gnd cell_6t
Xbit_r201_c19 bl[19] br[19] wl[201] vdd gnd cell_6t
Xbit_r202_c19 bl[19] br[19] wl[202] vdd gnd cell_6t
Xbit_r203_c19 bl[19] br[19] wl[203] vdd gnd cell_6t
Xbit_r204_c19 bl[19] br[19] wl[204] vdd gnd cell_6t
Xbit_r205_c19 bl[19] br[19] wl[205] vdd gnd cell_6t
Xbit_r206_c19 bl[19] br[19] wl[206] vdd gnd cell_6t
Xbit_r207_c19 bl[19] br[19] wl[207] vdd gnd cell_6t
Xbit_r208_c19 bl[19] br[19] wl[208] vdd gnd cell_6t
Xbit_r209_c19 bl[19] br[19] wl[209] vdd gnd cell_6t
Xbit_r210_c19 bl[19] br[19] wl[210] vdd gnd cell_6t
Xbit_r211_c19 bl[19] br[19] wl[211] vdd gnd cell_6t
Xbit_r212_c19 bl[19] br[19] wl[212] vdd gnd cell_6t
Xbit_r213_c19 bl[19] br[19] wl[213] vdd gnd cell_6t
Xbit_r214_c19 bl[19] br[19] wl[214] vdd gnd cell_6t
Xbit_r215_c19 bl[19] br[19] wl[215] vdd gnd cell_6t
Xbit_r216_c19 bl[19] br[19] wl[216] vdd gnd cell_6t
Xbit_r217_c19 bl[19] br[19] wl[217] vdd gnd cell_6t
Xbit_r218_c19 bl[19] br[19] wl[218] vdd gnd cell_6t
Xbit_r219_c19 bl[19] br[19] wl[219] vdd gnd cell_6t
Xbit_r220_c19 bl[19] br[19] wl[220] vdd gnd cell_6t
Xbit_r221_c19 bl[19] br[19] wl[221] vdd gnd cell_6t
Xbit_r222_c19 bl[19] br[19] wl[222] vdd gnd cell_6t
Xbit_r223_c19 bl[19] br[19] wl[223] vdd gnd cell_6t
Xbit_r224_c19 bl[19] br[19] wl[224] vdd gnd cell_6t
Xbit_r225_c19 bl[19] br[19] wl[225] vdd gnd cell_6t
Xbit_r226_c19 bl[19] br[19] wl[226] vdd gnd cell_6t
Xbit_r227_c19 bl[19] br[19] wl[227] vdd gnd cell_6t
Xbit_r228_c19 bl[19] br[19] wl[228] vdd gnd cell_6t
Xbit_r229_c19 bl[19] br[19] wl[229] vdd gnd cell_6t
Xbit_r230_c19 bl[19] br[19] wl[230] vdd gnd cell_6t
Xbit_r231_c19 bl[19] br[19] wl[231] vdd gnd cell_6t
Xbit_r232_c19 bl[19] br[19] wl[232] vdd gnd cell_6t
Xbit_r233_c19 bl[19] br[19] wl[233] vdd gnd cell_6t
Xbit_r234_c19 bl[19] br[19] wl[234] vdd gnd cell_6t
Xbit_r235_c19 bl[19] br[19] wl[235] vdd gnd cell_6t
Xbit_r236_c19 bl[19] br[19] wl[236] vdd gnd cell_6t
Xbit_r237_c19 bl[19] br[19] wl[237] vdd gnd cell_6t
Xbit_r238_c19 bl[19] br[19] wl[238] vdd gnd cell_6t
Xbit_r239_c19 bl[19] br[19] wl[239] vdd gnd cell_6t
Xbit_r240_c19 bl[19] br[19] wl[240] vdd gnd cell_6t
Xbit_r241_c19 bl[19] br[19] wl[241] vdd gnd cell_6t
Xbit_r242_c19 bl[19] br[19] wl[242] vdd gnd cell_6t
Xbit_r243_c19 bl[19] br[19] wl[243] vdd gnd cell_6t
Xbit_r244_c19 bl[19] br[19] wl[244] vdd gnd cell_6t
Xbit_r245_c19 bl[19] br[19] wl[245] vdd gnd cell_6t
Xbit_r246_c19 bl[19] br[19] wl[246] vdd gnd cell_6t
Xbit_r247_c19 bl[19] br[19] wl[247] vdd gnd cell_6t
Xbit_r248_c19 bl[19] br[19] wl[248] vdd gnd cell_6t
Xbit_r249_c19 bl[19] br[19] wl[249] vdd gnd cell_6t
Xbit_r250_c19 bl[19] br[19] wl[250] vdd gnd cell_6t
Xbit_r251_c19 bl[19] br[19] wl[251] vdd gnd cell_6t
Xbit_r252_c19 bl[19] br[19] wl[252] vdd gnd cell_6t
Xbit_r253_c19 bl[19] br[19] wl[253] vdd gnd cell_6t
Xbit_r254_c19 bl[19] br[19] wl[254] vdd gnd cell_6t
Xbit_r255_c19 bl[19] br[19] wl[255] vdd gnd cell_6t
Xbit_r0_c20 bl[20] br[20] wl[0] vdd gnd cell_6t
Xbit_r1_c20 bl[20] br[20] wl[1] vdd gnd cell_6t
Xbit_r2_c20 bl[20] br[20] wl[2] vdd gnd cell_6t
Xbit_r3_c20 bl[20] br[20] wl[3] vdd gnd cell_6t
Xbit_r4_c20 bl[20] br[20] wl[4] vdd gnd cell_6t
Xbit_r5_c20 bl[20] br[20] wl[5] vdd gnd cell_6t
Xbit_r6_c20 bl[20] br[20] wl[6] vdd gnd cell_6t
Xbit_r7_c20 bl[20] br[20] wl[7] vdd gnd cell_6t
Xbit_r8_c20 bl[20] br[20] wl[8] vdd gnd cell_6t
Xbit_r9_c20 bl[20] br[20] wl[9] vdd gnd cell_6t
Xbit_r10_c20 bl[20] br[20] wl[10] vdd gnd cell_6t
Xbit_r11_c20 bl[20] br[20] wl[11] vdd gnd cell_6t
Xbit_r12_c20 bl[20] br[20] wl[12] vdd gnd cell_6t
Xbit_r13_c20 bl[20] br[20] wl[13] vdd gnd cell_6t
Xbit_r14_c20 bl[20] br[20] wl[14] vdd gnd cell_6t
Xbit_r15_c20 bl[20] br[20] wl[15] vdd gnd cell_6t
Xbit_r16_c20 bl[20] br[20] wl[16] vdd gnd cell_6t
Xbit_r17_c20 bl[20] br[20] wl[17] vdd gnd cell_6t
Xbit_r18_c20 bl[20] br[20] wl[18] vdd gnd cell_6t
Xbit_r19_c20 bl[20] br[20] wl[19] vdd gnd cell_6t
Xbit_r20_c20 bl[20] br[20] wl[20] vdd gnd cell_6t
Xbit_r21_c20 bl[20] br[20] wl[21] vdd gnd cell_6t
Xbit_r22_c20 bl[20] br[20] wl[22] vdd gnd cell_6t
Xbit_r23_c20 bl[20] br[20] wl[23] vdd gnd cell_6t
Xbit_r24_c20 bl[20] br[20] wl[24] vdd gnd cell_6t
Xbit_r25_c20 bl[20] br[20] wl[25] vdd gnd cell_6t
Xbit_r26_c20 bl[20] br[20] wl[26] vdd gnd cell_6t
Xbit_r27_c20 bl[20] br[20] wl[27] vdd gnd cell_6t
Xbit_r28_c20 bl[20] br[20] wl[28] vdd gnd cell_6t
Xbit_r29_c20 bl[20] br[20] wl[29] vdd gnd cell_6t
Xbit_r30_c20 bl[20] br[20] wl[30] vdd gnd cell_6t
Xbit_r31_c20 bl[20] br[20] wl[31] vdd gnd cell_6t
Xbit_r32_c20 bl[20] br[20] wl[32] vdd gnd cell_6t
Xbit_r33_c20 bl[20] br[20] wl[33] vdd gnd cell_6t
Xbit_r34_c20 bl[20] br[20] wl[34] vdd gnd cell_6t
Xbit_r35_c20 bl[20] br[20] wl[35] vdd gnd cell_6t
Xbit_r36_c20 bl[20] br[20] wl[36] vdd gnd cell_6t
Xbit_r37_c20 bl[20] br[20] wl[37] vdd gnd cell_6t
Xbit_r38_c20 bl[20] br[20] wl[38] vdd gnd cell_6t
Xbit_r39_c20 bl[20] br[20] wl[39] vdd gnd cell_6t
Xbit_r40_c20 bl[20] br[20] wl[40] vdd gnd cell_6t
Xbit_r41_c20 bl[20] br[20] wl[41] vdd gnd cell_6t
Xbit_r42_c20 bl[20] br[20] wl[42] vdd gnd cell_6t
Xbit_r43_c20 bl[20] br[20] wl[43] vdd gnd cell_6t
Xbit_r44_c20 bl[20] br[20] wl[44] vdd gnd cell_6t
Xbit_r45_c20 bl[20] br[20] wl[45] vdd gnd cell_6t
Xbit_r46_c20 bl[20] br[20] wl[46] vdd gnd cell_6t
Xbit_r47_c20 bl[20] br[20] wl[47] vdd gnd cell_6t
Xbit_r48_c20 bl[20] br[20] wl[48] vdd gnd cell_6t
Xbit_r49_c20 bl[20] br[20] wl[49] vdd gnd cell_6t
Xbit_r50_c20 bl[20] br[20] wl[50] vdd gnd cell_6t
Xbit_r51_c20 bl[20] br[20] wl[51] vdd gnd cell_6t
Xbit_r52_c20 bl[20] br[20] wl[52] vdd gnd cell_6t
Xbit_r53_c20 bl[20] br[20] wl[53] vdd gnd cell_6t
Xbit_r54_c20 bl[20] br[20] wl[54] vdd gnd cell_6t
Xbit_r55_c20 bl[20] br[20] wl[55] vdd gnd cell_6t
Xbit_r56_c20 bl[20] br[20] wl[56] vdd gnd cell_6t
Xbit_r57_c20 bl[20] br[20] wl[57] vdd gnd cell_6t
Xbit_r58_c20 bl[20] br[20] wl[58] vdd gnd cell_6t
Xbit_r59_c20 bl[20] br[20] wl[59] vdd gnd cell_6t
Xbit_r60_c20 bl[20] br[20] wl[60] vdd gnd cell_6t
Xbit_r61_c20 bl[20] br[20] wl[61] vdd gnd cell_6t
Xbit_r62_c20 bl[20] br[20] wl[62] vdd gnd cell_6t
Xbit_r63_c20 bl[20] br[20] wl[63] vdd gnd cell_6t
Xbit_r64_c20 bl[20] br[20] wl[64] vdd gnd cell_6t
Xbit_r65_c20 bl[20] br[20] wl[65] vdd gnd cell_6t
Xbit_r66_c20 bl[20] br[20] wl[66] vdd gnd cell_6t
Xbit_r67_c20 bl[20] br[20] wl[67] vdd gnd cell_6t
Xbit_r68_c20 bl[20] br[20] wl[68] vdd gnd cell_6t
Xbit_r69_c20 bl[20] br[20] wl[69] vdd gnd cell_6t
Xbit_r70_c20 bl[20] br[20] wl[70] vdd gnd cell_6t
Xbit_r71_c20 bl[20] br[20] wl[71] vdd gnd cell_6t
Xbit_r72_c20 bl[20] br[20] wl[72] vdd gnd cell_6t
Xbit_r73_c20 bl[20] br[20] wl[73] vdd gnd cell_6t
Xbit_r74_c20 bl[20] br[20] wl[74] vdd gnd cell_6t
Xbit_r75_c20 bl[20] br[20] wl[75] vdd gnd cell_6t
Xbit_r76_c20 bl[20] br[20] wl[76] vdd gnd cell_6t
Xbit_r77_c20 bl[20] br[20] wl[77] vdd gnd cell_6t
Xbit_r78_c20 bl[20] br[20] wl[78] vdd gnd cell_6t
Xbit_r79_c20 bl[20] br[20] wl[79] vdd gnd cell_6t
Xbit_r80_c20 bl[20] br[20] wl[80] vdd gnd cell_6t
Xbit_r81_c20 bl[20] br[20] wl[81] vdd gnd cell_6t
Xbit_r82_c20 bl[20] br[20] wl[82] vdd gnd cell_6t
Xbit_r83_c20 bl[20] br[20] wl[83] vdd gnd cell_6t
Xbit_r84_c20 bl[20] br[20] wl[84] vdd gnd cell_6t
Xbit_r85_c20 bl[20] br[20] wl[85] vdd gnd cell_6t
Xbit_r86_c20 bl[20] br[20] wl[86] vdd gnd cell_6t
Xbit_r87_c20 bl[20] br[20] wl[87] vdd gnd cell_6t
Xbit_r88_c20 bl[20] br[20] wl[88] vdd gnd cell_6t
Xbit_r89_c20 bl[20] br[20] wl[89] vdd gnd cell_6t
Xbit_r90_c20 bl[20] br[20] wl[90] vdd gnd cell_6t
Xbit_r91_c20 bl[20] br[20] wl[91] vdd gnd cell_6t
Xbit_r92_c20 bl[20] br[20] wl[92] vdd gnd cell_6t
Xbit_r93_c20 bl[20] br[20] wl[93] vdd gnd cell_6t
Xbit_r94_c20 bl[20] br[20] wl[94] vdd gnd cell_6t
Xbit_r95_c20 bl[20] br[20] wl[95] vdd gnd cell_6t
Xbit_r96_c20 bl[20] br[20] wl[96] vdd gnd cell_6t
Xbit_r97_c20 bl[20] br[20] wl[97] vdd gnd cell_6t
Xbit_r98_c20 bl[20] br[20] wl[98] vdd gnd cell_6t
Xbit_r99_c20 bl[20] br[20] wl[99] vdd gnd cell_6t
Xbit_r100_c20 bl[20] br[20] wl[100] vdd gnd cell_6t
Xbit_r101_c20 bl[20] br[20] wl[101] vdd gnd cell_6t
Xbit_r102_c20 bl[20] br[20] wl[102] vdd gnd cell_6t
Xbit_r103_c20 bl[20] br[20] wl[103] vdd gnd cell_6t
Xbit_r104_c20 bl[20] br[20] wl[104] vdd gnd cell_6t
Xbit_r105_c20 bl[20] br[20] wl[105] vdd gnd cell_6t
Xbit_r106_c20 bl[20] br[20] wl[106] vdd gnd cell_6t
Xbit_r107_c20 bl[20] br[20] wl[107] vdd gnd cell_6t
Xbit_r108_c20 bl[20] br[20] wl[108] vdd gnd cell_6t
Xbit_r109_c20 bl[20] br[20] wl[109] vdd gnd cell_6t
Xbit_r110_c20 bl[20] br[20] wl[110] vdd gnd cell_6t
Xbit_r111_c20 bl[20] br[20] wl[111] vdd gnd cell_6t
Xbit_r112_c20 bl[20] br[20] wl[112] vdd gnd cell_6t
Xbit_r113_c20 bl[20] br[20] wl[113] vdd gnd cell_6t
Xbit_r114_c20 bl[20] br[20] wl[114] vdd gnd cell_6t
Xbit_r115_c20 bl[20] br[20] wl[115] vdd gnd cell_6t
Xbit_r116_c20 bl[20] br[20] wl[116] vdd gnd cell_6t
Xbit_r117_c20 bl[20] br[20] wl[117] vdd gnd cell_6t
Xbit_r118_c20 bl[20] br[20] wl[118] vdd gnd cell_6t
Xbit_r119_c20 bl[20] br[20] wl[119] vdd gnd cell_6t
Xbit_r120_c20 bl[20] br[20] wl[120] vdd gnd cell_6t
Xbit_r121_c20 bl[20] br[20] wl[121] vdd gnd cell_6t
Xbit_r122_c20 bl[20] br[20] wl[122] vdd gnd cell_6t
Xbit_r123_c20 bl[20] br[20] wl[123] vdd gnd cell_6t
Xbit_r124_c20 bl[20] br[20] wl[124] vdd gnd cell_6t
Xbit_r125_c20 bl[20] br[20] wl[125] vdd gnd cell_6t
Xbit_r126_c20 bl[20] br[20] wl[126] vdd gnd cell_6t
Xbit_r127_c20 bl[20] br[20] wl[127] vdd gnd cell_6t
Xbit_r128_c20 bl[20] br[20] wl[128] vdd gnd cell_6t
Xbit_r129_c20 bl[20] br[20] wl[129] vdd gnd cell_6t
Xbit_r130_c20 bl[20] br[20] wl[130] vdd gnd cell_6t
Xbit_r131_c20 bl[20] br[20] wl[131] vdd gnd cell_6t
Xbit_r132_c20 bl[20] br[20] wl[132] vdd gnd cell_6t
Xbit_r133_c20 bl[20] br[20] wl[133] vdd gnd cell_6t
Xbit_r134_c20 bl[20] br[20] wl[134] vdd gnd cell_6t
Xbit_r135_c20 bl[20] br[20] wl[135] vdd gnd cell_6t
Xbit_r136_c20 bl[20] br[20] wl[136] vdd gnd cell_6t
Xbit_r137_c20 bl[20] br[20] wl[137] vdd gnd cell_6t
Xbit_r138_c20 bl[20] br[20] wl[138] vdd gnd cell_6t
Xbit_r139_c20 bl[20] br[20] wl[139] vdd gnd cell_6t
Xbit_r140_c20 bl[20] br[20] wl[140] vdd gnd cell_6t
Xbit_r141_c20 bl[20] br[20] wl[141] vdd gnd cell_6t
Xbit_r142_c20 bl[20] br[20] wl[142] vdd gnd cell_6t
Xbit_r143_c20 bl[20] br[20] wl[143] vdd gnd cell_6t
Xbit_r144_c20 bl[20] br[20] wl[144] vdd gnd cell_6t
Xbit_r145_c20 bl[20] br[20] wl[145] vdd gnd cell_6t
Xbit_r146_c20 bl[20] br[20] wl[146] vdd gnd cell_6t
Xbit_r147_c20 bl[20] br[20] wl[147] vdd gnd cell_6t
Xbit_r148_c20 bl[20] br[20] wl[148] vdd gnd cell_6t
Xbit_r149_c20 bl[20] br[20] wl[149] vdd gnd cell_6t
Xbit_r150_c20 bl[20] br[20] wl[150] vdd gnd cell_6t
Xbit_r151_c20 bl[20] br[20] wl[151] vdd gnd cell_6t
Xbit_r152_c20 bl[20] br[20] wl[152] vdd gnd cell_6t
Xbit_r153_c20 bl[20] br[20] wl[153] vdd gnd cell_6t
Xbit_r154_c20 bl[20] br[20] wl[154] vdd gnd cell_6t
Xbit_r155_c20 bl[20] br[20] wl[155] vdd gnd cell_6t
Xbit_r156_c20 bl[20] br[20] wl[156] vdd gnd cell_6t
Xbit_r157_c20 bl[20] br[20] wl[157] vdd gnd cell_6t
Xbit_r158_c20 bl[20] br[20] wl[158] vdd gnd cell_6t
Xbit_r159_c20 bl[20] br[20] wl[159] vdd gnd cell_6t
Xbit_r160_c20 bl[20] br[20] wl[160] vdd gnd cell_6t
Xbit_r161_c20 bl[20] br[20] wl[161] vdd gnd cell_6t
Xbit_r162_c20 bl[20] br[20] wl[162] vdd gnd cell_6t
Xbit_r163_c20 bl[20] br[20] wl[163] vdd gnd cell_6t
Xbit_r164_c20 bl[20] br[20] wl[164] vdd gnd cell_6t
Xbit_r165_c20 bl[20] br[20] wl[165] vdd gnd cell_6t
Xbit_r166_c20 bl[20] br[20] wl[166] vdd gnd cell_6t
Xbit_r167_c20 bl[20] br[20] wl[167] vdd gnd cell_6t
Xbit_r168_c20 bl[20] br[20] wl[168] vdd gnd cell_6t
Xbit_r169_c20 bl[20] br[20] wl[169] vdd gnd cell_6t
Xbit_r170_c20 bl[20] br[20] wl[170] vdd gnd cell_6t
Xbit_r171_c20 bl[20] br[20] wl[171] vdd gnd cell_6t
Xbit_r172_c20 bl[20] br[20] wl[172] vdd gnd cell_6t
Xbit_r173_c20 bl[20] br[20] wl[173] vdd gnd cell_6t
Xbit_r174_c20 bl[20] br[20] wl[174] vdd gnd cell_6t
Xbit_r175_c20 bl[20] br[20] wl[175] vdd gnd cell_6t
Xbit_r176_c20 bl[20] br[20] wl[176] vdd gnd cell_6t
Xbit_r177_c20 bl[20] br[20] wl[177] vdd gnd cell_6t
Xbit_r178_c20 bl[20] br[20] wl[178] vdd gnd cell_6t
Xbit_r179_c20 bl[20] br[20] wl[179] vdd gnd cell_6t
Xbit_r180_c20 bl[20] br[20] wl[180] vdd gnd cell_6t
Xbit_r181_c20 bl[20] br[20] wl[181] vdd gnd cell_6t
Xbit_r182_c20 bl[20] br[20] wl[182] vdd gnd cell_6t
Xbit_r183_c20 bl[20] br[20] wl[183] vdd gnd cell_6t
Xbit_r184_c20 bl[20] br[20] wl[184] vdd gnd cell_6t
Xbit_r185_c20 bl[20] br[20] wl[185] vdd gnd cell_6t
Xbit_r186_c20 bl[20] br[20] wl[186] vdd gnd cell_6t
Xbit_r187_c20 bl[20] br[20] wl[187] vdd gnd cell_6t
Xbit_r188_c20 bl[20] br[20] wl[188] vdd gnd cell_6t
Xbit_r189_c20 bl[20] br[20] wl[189] vdd gnd cell_6t
Xbit_r190_c20 bl[20] br[20] wl[190] vdd gnd cell_6t
Xbit_r191_c20 bl[20] br[20] wl[191] vdd gnd cell_6t
Xbit_r192_c20 bl[20] br[20] wl[192] vdd gnd cell_6t
Xbit_r193_c20 bl[20] br[20] wl[193] vdd gnd cell_6t
Xbit_r194_c20 bl[20] br[20] wl[194] vdd gnd cell_6t
Xbit_r195_c20 bl[20] br[20] wl[195] vdd gnd cell_6t
Xbit_r196_c20 bl[20] br[20] wl[196] vdd gnd cell_6t
Xbit_r197_c20 bl[20] br[20] wl[197] vdd gnd cell_6t
Xbit_r198_c20 bl[20] br[20] wl[198] vdd gnd cell_6t
Xbit_r199_c20 bl[20] br[20] wl[199] vdd gnd cell_6t
Xbit_r200_c20 bl[20] br[20] wl[200] vdd gnd cell_6t
Xbit_r201_c20 bl[20] br[20] wl[201] vdd gnd cell_6t
Xbit_r202_c20 bl[20] br[20] wl[202] vdd gnd cell_6t
Xbit_r203_c20 bl[20] br[20] wl[203] vdd gnd cell_6t
Xbit_r204_c20 bl[20] br[20] wl[204] vdd gnd cell_6t
Xbit_r205_c20 bl[20] br[20] wl[205] vdd gnd cell_6t
Xbit_r206_c20 bl[20] br[20] wl[206] vdd gnd cell_6t
Xbit_r207_c20 bl[20] br[20] wl[207] vdd gnd cell_6t
Xbit_r208_c20 bl[20] br[20] wl[208] vdd gnd cell_6t
Xbit_r209_c20 bl[20] br[20] wl[209] vdd gnd cell_6t
Xbit_r210_c20 bl[20] br[20] wl[210] vdd gnd cell_6t
Xbit_r211_c20 bl[20] br[20] wl[211] vdd gnd cell_6t
Xbit_r212_c20 bl[20] br[20] wl[212] vdd gnd cell_6t
Xbit_r213_c20 bl[20] br[20] wl[213] vdd gnd cell_6t
Xbit_r214_c20 bl[20] br[20] wl[214] vdd gnd cell_6t
Xbit_r215_c20 bl[20] br[20] wl[215] vdd gnd cell_6t
Xbit_r216_c20 bl[20] br[20] wl[216] vdd gnd cell_6t
Xbit_r217_c20 bl[20] br[20] wl[217] vdd gnd cell_6t
Xbit_r218_c20 bl[20] br[20] wl[218] vdd gnd cell_6t
Xbit_r219_c20 bl[20] br[20] wl[219] vdd gnd cell_6t
Xbit_r220_c20 bl[20] br[20] wl[220] vdd gnd cell_6t
Xbit_r221_c20 bl[20] br[20] wl[221] vdd gnd cell_6t
Xbit_r222_c20 bl[20] br[20] wl[222] vdd gnd cell_6t
Xbit_r223_c20 bl[20] br[20] wl[223] vdd gnd cell_6t
Xbit_r224_c20 bl[20] br[20] wl[224] vdd gnd cell_6t
Xbit_r225_c20 bl[20] br[20] wl[225] vdd gnd cell_6t
Xbit_r226_c20 bl[20] br[20] wl[226] vdd gnd cell_6t
Xbit_r227_c20 bl[20] br[20] wl[227] vdd gnd cell_6t
Xbit_r228_c20 bl[20] br[20] wl[228] vdd gnd cell_6t
Xbit_r229_c20 bl[20] br[20] wl[229] vdd gnd cell_6t
Xbit_r230_c20 bl[20] br[20] wl[230] vdd gnd cell_6t
Xbit_r231_c20 bl[20] br[20] wl[231] vdd gnd cell_6t
Xbit_r232_c20 bl[20] br[20] wl[232] vdd gnd cell_6t
Xbit_r233_c20 bl[20] br[20] wl[233] vdd gnd cell_6t
Xbit_r234_c20 bl[20] br[20] wl[234] vdd gnd cell_6t
Xbit_r235_c20 bl[20] br[20] wl[235] vdd gnd cell_6t
Xbit_r236_c20 bl[20] br[20] wl[236] vdd gnd cell_6t
Xbit_r237_c20 bl[20] br[20] wl[237] vdd gnd cell_6t
Xbit_r238_c20 bl[20] br[20] wl[238] vdd gnd cell_6t
Xbit_r239_c20 bl[20] br[20] wl[239] vdd gnd cell_6t
Xbit_r240_c20 bl[20] br[20] wl[240] vdd gnd cell_6t
Xbit_r241_c20 bl[20] br[20] wl[241] vdd gnd cell_6t
Xbit_r242_c20 bl[20] br[20] wl[242] vdd gnd cell_6t
Xbit_r243_c20 bl[20] br[20] wl[243] vdd gnd cell_6t
Xbit_r244_c20 bl[20] br[20] wl[244] vdd gnd cell_6t
Xbit_r245_c20 bl[20] br[20] wl[245] vdd gnd cell_6t
Xbit_r246_c20 bl[20] br[20] wl[246] vdd gnd cell_6t
Xbit_r247_c20 bl[20] br[20] wl[247] vdd gnd cell_6t
Xbit_r248_c20 bl[20] br[20] wl[248] vdd gnd cell_6t
Xbit_r249_c20 bl[20] br[20] wl[249] vdd gnd cell_6t
Xbit_r250_c20 bl[20] br[20] wl[250] vdd gnd cell_6t
Xbit_r251_c20 bl[20] br[20] wl[251] vdd gnd cell_6t
Xbit_r252_c20 bl[20] br[20] wl[252] vdd gnd cell_6t
Xbit_r253_c20 bl[20] br[20] wl[253] vdd gnd cell_6t
Xbit_r254_c20 bl[20] br[20] wl[254] vdd gnd cell_6t
Xbit_r255_c20 bl[20] br[20] wl[255] vdd gnd cell_6t
Xbit_r0_c21 bl[21] br[21] wl[0] vdd gnd cell_6t
Xbit_r1_c21 bl[21] br[21] wl[1] vdd gnd cell_6t
Xbit_r2_c21 bl[21] br[21] wl[2] vdd gnd cell_6t
Xbit_r3_c21 bl[21] br[21] wl[3] vdd gnd cell_6t
Xbit_r4_c21 bl[21] br[21] wl[4] vdd gnd cell_6t
Xbit_r5_c21 bl[21] br[21] wl[5] vdd gnd cell_6t
Xbit_r6_c21 bl[21] br[21] wl[6] vdd gnd cell_6t
Xbit_r7_c21 bl[21] br[21] wl[7] vdd gnd cell_6t
Xbit_r8_c21 bl[21] br[21] wl[8] vdd gnd cell_6t
Xbit_r9_c21 bl[21] br[21] wl[9] vdd gnd cell_6t
Xbit_r10_c21 bl[21] br[21] wl[10] vdd gnd cell_6t
Xbit_r11_c21 bl[21] br[21] wl[11] vdd gnd cell_6t
Xbit_r12_c21 bl[21] br[21] wl[12] vdd gnd cell_6t
Xbit_r13_c21 bl[21] br[21] wl[13] vdd gnd cell_6t
Xbit_r14_c21 bl[21] br[21] wl[14] vdd gnd cell_6t
Xbit_r15_c21 bl[21] br[21] wl[15] vdd gnd cell_6t
Xbit_r16_c21 bl[21] br[21] wl[16] vdd gnd cell_6t
Xbit_r17_c21 bl[21] br[21] wl[17] vdd gnd cell_6t
Xbit_r18_c21 bl[21] br[21] wl[18] vdd gnd cell_6t
Xbit_r19_c21 bl[21] br[21] wl[19] vdd gnd cell_6t
Xbit_r20_c21 bl[21] br[21] wl[20] vdd gnd cell_6t
Xbit_r21_c21 bl[21] br[21] wl[21] vdd gnd cell_6t
Xbit_r22_c21 bl[21] br[21] wl[22] vdd gnd cell_6t
Xbit_r23_c21 bl[21] br[21] wl[23] vdd gnd cell_6t
Xbit_r24_c21 bl[21] br[21] wl[24] vdd gnd cell_6t
Xbit_r25_c21 bl[21] br[21] wl[25] vdd gnd cell_6t
Xbit_r26_c21 bl[21] br[21] wl[26] vdd gnd cell_6t
Xbit_r27_c21 bl[21] br[21] wl[27] vdd gnd cell_6t
Xbit_r28_c21 bl[21] br[21] wl[28] vdd gnd cell_6t
Xbit_r29_c21 bl[21] br[21] wl[29] vdd gnd cell_6t
Xbit_r30_c21 bl[21] br[21] wl[30] vdd gnd cell_6t
Xbit_r31_c21 bl[21] br[21] wl[31] vdd gnd cell_6t
Xbit_r32_c21 bl[21] br[21] wl[32] vdd gnd cell_6t
Xbit_r33_c21 bl[21] br[21] wl[33] vdd gnd cell_6t
Xbit_r34_c21 bl[21] br[21] wl[34] vdd gnd cell_6t
Xbit_r35_c21 bl[21] br[21] wl[35] vdd gnd cell_6t
Xbit_r36_c21 bl[21] br[21] wl[36] vdd gnd cell_6t
Xbit_r37_c21 bl[21] br[21] wl[37] vdd gnd cell_6t
Xbit_r38_c21 bl[21] br[21] wl[38] vdd gnd cell_6t
Xbit_r39_c21 bl[21] br[21] wl[39] vdd gnd cell_6t
Xbit_r40_c21 bl[21] br[21] wl[40] vdd gnd cell_6t
Xbit_r41_c21 bl[21] br[21] wl[41] vdd gnd cell_6t
Xbit_r42_c21 bl[21] br[21] wl[42] vdd gnd cell_6t
Xbit_r43_c21 bl[21] br[21] wl[43] vdd gnd cell_6t
Xbit_r44_c21 bl[21] br[21] wl[44] vdd gnd cell_6t
Xbit_r45_c21 bl[21] br[21] wl[45] vdd gnd cell_6t
Xbit_r46_c21 bl[21] br[21] wl[46] vdd gnd cell_6t
Xbit_r47_c21 bl[21] br[21] wl[47] vdd gnd cell_6t
Xbit_r48_c21 bl[21] br[21] wl[48] vdd gnd cell_6t
Xbit_r49_c21 bl[21] br[21] wl[49] vdd gnd cell_6t
Xbit_r50_c21 bl[21] br[21] wl[50] vdd gnd cell_6t
Xbit_r51_c21 bl[21] br[21] wl[51] vdd gnd cell_6t
Xbit_r52_c21 bl[21] br[21] wl[52] vdd gnd cell_6t
Xbit_r53_c21 bl[21] br[21] wl[53] vdd gnd cell_6t
Xbit_r54_c21 bl[21] br[21] wl[54] vdd gnd cell_6t
Xbit_r55_c21 bl[21] br[21] wl[55] vdd gnd cell_6t
Xbit_r56_c21 bl[21] br[21] wl[56] vdd gnd cell_6t
Xbit_r57_c21 bl[21] br[21] wl[57] vdd gnd cell_6t
Xbit_r58_c21 bl[21] br[21] wl[58] vdd gnd cell_6t
Xbit_r59_c21 bl[21] br[21] wl[59] vdd gnd cell_6t
Xbit_r60_c21 bl[21] br[21] wl[60] vdd gnd cell_6t
Xbit_r61_c21 bl[21] br[21] wl[61] vdd gnd cell_6t
Xbit_r62_c21 bl[21] br[21] wl[62] vdd gnd cell_6t
Xbit_r63_c21 bl[21] br[21] wl[63] vdd gnd cell_6t
Xbit_r64_c21 bl[21] br[21] wl[64] vdd gnd cell_6t
Xbit_r65_c21 bl[21] br[21] wl[65] vdd gnd cell_6t
Xbit_r66_c21 bl[21] br[21] wl[66] vdd gnd cell_6t
Xbit_r67_c21 bl[21] br[21] wl[67] vdd gnd cell_6t
Xbit_r68_c21 bl[21] br[21] wl[68] vdd gnd cell_6t
Xbit_r69_c21 bl[21] br[21] wl[69] vdd gnd cell_6t
Xbit_r70_c21 bl[21] br[21] wl[70] vdd gnd cell_6t
Xbit_r71_c21 bl[21] br[21] wl[71] vdd gnd cell_6t
Xbit_r72_c21 bl[21] br[21] wl[72] vdd gnd cell_6t
Xbit_r73_c21 bl[21] br[21] wl[73] vdd gnd cell_6t
Xbit_r74_c21 bl[21] br[21] wl[74] vdd gnd cell_6t
Xbit_r75_c21 bl[21] br[21] wl[75] vdd gnd cell_6t
Xbit_r76_c21 bl[21] br[21] wl[76] vdd gnd cell_6t
Xbit_r77_c21 bl[21] br[21] wl[77] vdd gnd cell_6t
Xbit_r78_c21 bl[21] br[21] wl[78] vdd gnd cell_6t
Xbit_r79_c21 bl[21] br[21] wl[79] vdd gnd cell_6t
Xbit_r80_c21 bl[21] br[21] wl[80] vdd gnd cell_6t
Xbit_r81_c21 bl[21] br[21] wl[81] vdd gnd cell_6t
Xbit_r82_c21 bl[21] br[21] wl[82] vdd gnd cell_6t
Xbit_r83_c21 bl[21] br[21] wl[83] vdd gnd cell_6t
Xbit_r84_c21 bl[21] br[21] wl[84] vdd gnd cell_6t
Xbit_r85_c21 bl[21] br[21] wl[85] vdd gnd cell_6t
Xbit_r86_c21 bl[21] br[21] wl[86] vdd gnd cell_6t
Xbit_r87_c21 bl[21] br[21] wl[87] vdd gnd cell_6t
Xbit_r88_c21 bl[21] br[21] wl[88] vdd gnd cell_6t
Xbit_r89_c21 bl[21] br[21] wl[89] vdd gnd cell_6t
Xbit_r90_c21 bl[21] br[21] wl[90] vdd gnd cell_6t
Xbit_r91_c21 bl[21] br[21] wl[91] vdd gnd cell_6t
Xbit_r92_c21 bl[21] br[21] wl[92] vdd gnd cell_6t
Xbit_r93_c21 bl[21] br[21] wl[93] vdd gnd cell_6t
Xbit_r94_c21 bl[21] br[21] wl[94] vdd gnd cell_6t
Xbit_r95_c21 bl[21] br[21] wl[95] vdd gnd cell_6t
Xbit_r96_c21 bl[21] br[21] wl[96] vdd gnd cell_6t
Xbit_r97_c21 bl[21] br[21] wl[97] vdd gnd cell_6t
Xbit_r98_c21 bl[21] br[21] wl[98] vdd gnd cell_6t
Xbit_r99_c21 bl[21] br[21] wl[99] vdd gnd cell_6t
Xbit_r100_c21 bl[21] br[21] wl[100] vdd gnd cell_6t
Xbit_r101_c21 bl[21] br[21] wl[101] vdd gnd cell_6t
Xbit_r102_c21 bl[21] br[21] wl[102] vdd gnd cell_6t
Xbit_r103_c21 bl[21] br[21] wl[103] vdd gnd cell_6t
Xbit_r104_c21 bl[21] br[21] wl[104] vdd gnd cell_6t
Xbit_r105_c21 bl[21] br[21] wl[105] vdd gnd cell_6t
Xbit_r106_c21 bl[21] br[21] wl[106] vdd gnd cell_6t
Xbit_r107_c21 bl[21] br[21] wl[107] vdd gnd cell_6t
Xbit_r108_c21 bl[21] br[21] wl[108] vdd gnd cell_6t
Xbit_r109_c21 bl[21] br[21] wl[109] vdd gnd cell_6t
Xbit_r110_c21 bl[21] br[21] wl[110] vdd gnd cell_6t
Xbit_r111_c21 bl[21] br[21] wl[111] vdd gnd cell_6t
Xbit_r112_c21 bl[21] br[21] wl[112] vdd gnd cell_6t
Xbit_r113_c21 bl[21] br[21] wl[113] vdd gnd cell_6t
Xbit_r114_c21 bl[21] br[21] wl[114] vdd gnd cell_6t
Xbit_r115_c21 bl[21] br[21] wl[115] vdd gnd cell_6t
Xbit_r116_c21 bl[21] br[21] wl[116] vdd gnd cell_6t
Xbit_r117_c21 bl[21] br[21] wl[117] vdd gnd cell_6t
Xbit_r118_c21 bl[21] br[21] wl[118] vdd gnd cell_6t
Xbit_r119_c21 bl[21] br[21] wl[119] vdd gnd cell_6t
Xbit_r120_c21 bl[21] br[21] wl[120] vdd gnd cell_6t
Xbit_r121_c21 bl[21] br[21] wl[121] vdd gnd cell_6t
Xbit_r122_c21 bl[21] br[21] wl[122] vdd gnd cell_6t
Xbit_r123_c21 bl[21] br[21] wl[123] vdd gnd cell_6t
Xbit_r124_c21 bl[21] br[21] wl[124] vdd gnd cell_6t
Xbit_r125_c21 bl[21] br[21] wl[125] vdd gnd cell_6t
Xbit_r126_c21 bl[21] br[21] wl[126] vdd gnd cell_6t
Xbit_r127_c21 bl[21] br[21] wl[127] vdd gnd cell_6t
Xbit_r128_c21 bl[21] br[21] wl[128] vdd gnd cell_6t
Xbit_r129_c21 bl[21] br[21] wl[129] vdd gnd cell_6t
Xbit_r130_c21 bl[21] br[21] wl[130] vdd gnd cell_6t
Xbit_r131_c21 bl[21] br[21] wl[131] vdd gnd cell_6t
Xbit_r132_c21 bl[21] br[21] wl[132] vdd gnd cell_6t
Xbit_r133_c21 bl[21] br[21] wl[133] vdd gnd cell_6t
Xbit_r134_c21 bl[21] br[21] wl[134] vdd gnd cell_6t
Xbit_r135_c21 bl[21] br[21] wl[135] vdd gnd cell_6t
Xbit_r136_c21 bl[21] br[21] wl[136] vdd gnd cell_6t
Xbit_r137_c21 bl[21] br[21] wl[137] vdd gnd cell_6t
Xbit_r138_c21 bl[21] br[21] wl[138] vdd gnd cell_6t
Xbit_r139_c21 bl[21] br[21] wl[139] vdd gnd cell_6t
Xbit_r140_c21 bl[21] br[21] wl[140] vdd gnd cell_6t
Xbit_r141_c21 bl[21] br[21] wl[141] vdd gnd cell_6t
Xbit_r142_c21 bl[21] br[21] wl[142] vdd gnd cell_6t
Xbit_r143_c21 bl[21] br[21] wl[143] vdd gnd cell_6t
Xbit_r144_c21 bl[21] br[21] wl[144] vdd gnd cell_6t
Xbit_r145_c21 bl[21] br[21] wl[145] vdd gnd cell_6t
Xbit_r146_c21 bl[21] br[21] wl[146] vdd gnd cell_6t
Xbit_r147_c21 bl[21] br[21] wl[147] vdd gnd cell_6t
Xbit_r148_c21 bl[21] br[21] wl[148] vdd gnd cell_6t
Xbit_r149_c21 bl[21] br[21] wl[149] vdd gnd cell_6t
Xbit_r150_c21 bl[21] br[21] wl[150] vdd gnd cell_6t
Xbit_r151_c21 bl[21] br[21] wl[151] vdd gnd cell_6t
Xbit_r152_c21 bl[21] br[21] wl[152] vdd gnd cell_6t
Xbit_r153_c21 bl[21] br[21] wl[153] vdd gnd cell_6t
Xbit_r154_c21 bl[21] br[21] wl[154] vdd gnd cell_6t
Xbit_r155_c21 bl[21] br[21] wl[155] vdd gnd cell_6t
Xbit_r156_c21 bl[21] br[21] wl[156] vdd gnd cell_6t
Xbit_r157_c21 bl[21] br[21] wl[157] vdd gnd cell_6t
Xbit_r158_c21 bl[21] br[21] wl[158] vdd gnd cell_6t
Xbit_r159_c21 bl[21] br[21] wl[159] vdd gnd cell_6t
Xbit_r160_c21 bl[21] br[21] wl[160] vdd gnd cell_6t
Xbit_r161_c21 bl[21] br[21] wl[161] vdd gnd cell_6t
Xbit_r162_c21 bl[21] br[21] wl[162] vdd gnd cell_6t
Xbit_r163_c21 bl[21] br[21] wl[163] vdd gnd cell_6t
Xbit_r164_c21 bl[21] br[21] wl[164] vdd gnd cell_6t
Xbit_r165_c21 bl[21] br[21] wl[165] vdd gnd cell_6t
Xbit_r166_c21 bl[21] br[21] wl[166] vdd gnd cell_6t
Xbit_r167_c21 bl[21] br[21] wl[167] vdd gnd cell_6t
Xbit_r168_c21 bl[21] br[21] wl[168] vdd gnd cell_6t
Xbit_r169_c21 bl[21] br[21] wl[169] vdd gnd cell_6t
Xbit_r170_c21 bl[21] br[21] wl[170] vdd gnd cell_6t
Xbit_r171_c21 bl[21] br[21] wl[171] vdd gnd cell_6t
Xbit_r172_c21 bl[21] br[21] wl[172] vdd gnd cell_6t
Xbit_r173_c21 bl[21] br[21] wl[173] vdd gnd cell_6t
Xbit_r174_c21 bl[21] br[21] wl[174] vdd gnd cell_6t
Xbit_r175_c21 bl[21] br[21] wl[175] vdd gnd cell_6t
Xbit_r176_c21 bl[21] br[21] wl[176] vdd gnd cell_6t
Xbit_r177_c21 bl[21] br[21] wl[177] vdd gnd cell_6t
Xbit_r178_c21 bl[21] br[21] wl[178] vdd gnd cell_6t
Xbit_r179_c21 bl[21] br[21] wl[179] vdd gnd cell_6t
Xbit_r180_c21 bl[21] br[21] wl[180] vdd gnd cell_6t
Xbit_r181_c21 bl[21] br[21] wl[181] vdd gnd cell_6t
Xbit_r182_c21 bl[21] br[21] wl[182] vdd gnd cell_6t
Xbit_r183_c21 bl[21] br[21] wl[183] vdd gnd cell_6t
Xbit_r184_c21 bl[21] br[21] wl[184] vdd gnd cell_6t
Xbit_r185_c21 bl[21] br[21] wl[185] vdd gnd cell_6t
Xbit_r186_c21 bl[21] br[21] wl[186] vdd gnd cell_6t
Xbit_r187_c21 bl[21] br[21] wl[187] vdd gnd cell_6t
Xbit_r188_c21 bl[21] br[21] wl[188] vdd gnd cell_6t
Xbit_r189_c21 bl[21] br[21] wl[189] vdd gnd cell_6t
Xbit_r190_c21 bl[21] br[21] wl[190] vdd gnd cell_6t
Xbit_r191_c21 bl[21] br[21] wl[191] vdd gnd cell_6t
Xbit_r192_c21 bl[21] br[21] wl[192] vdd gnd cell_6t
Xbit_r193_c21 bl[21] br[21] wl[193] vdd gnd cell_6t
Xbit_r194_c21 bl[21] br[21] wl[194] vdd gnd cell_6t
Xbit_r195_c21 bl[21] br[21] wl[195] vdd gnd cell_6t
Xbit_r196_c21 bl[21] br[21] wl[196] vdd gnd cell_6t
Xbit_r197_c21 bl[21] br[21] wl[197] vdd gnd cell_6t
Xbit_r198_c21 bl[21] br[21] wl[198] vdd gnd cell_6t
Xbit_r199_c21 bl[21] br[21] wl[199] vdd gnd cell_6t
Xbit_r200_c21 bl[21] br[21] wl[200] vdd gnd cell_6t
Xbit_r201_c21 bl[21] br[21] wl[201] vdd gnd cell_6t
Xbit_r202_c21 bl[21] br[21] wl[202] vdd gnd cell_6t
Xbit_r203_c21 bl[21] br[21] wl[203] vdd gnd cell_6t
Xbit_r204_c21 bl[21] br[21] wl[204] vdd gnd cell_6t
Xbit_r205_c21 bl[21] br[21] wl[205] vdd gnd cell_6t
Xbit_r206_c21 bl[21] br[21] wl[206] vdd gnd cell_6t
Xbit_r207_c21 bl[21] br[21] wl[207] vdd gnd cell_6t
Xbit_r208_c21 bl[21] br[21] wl[208] vdd gnd cell_6t
Xbit_r209_c21 bl[21] br[21] wl[209] vdd gnd cell_6t
Xbit_r210_c21 bl[21] br[21] wl[210] vdd gnd cell_6t
Xbit_r211_c21 bl[21] br[21] wl[211] vdd gnd cell_6t
Xbit_r212_c21 bl[21] br[21] wl[212] vdd gnd cell_6t
Xbit_r213_c21 bl[21] br[21] wl[213] vdd gnd cell_6t
Xbit_r214_c21 bl[21] br[21] wl[214] vdd gnd cell_6t
Xbit_r215_c21 bl[21] br[21] wl[215] vdd gnd cell_6t
Xbit_r216_c21 bl[21] br[21] wl[216] vdd gnd cell_6t
Xbit_r217_c21 bl[21] br[21] wl[217] vdd gnd cell_6t
Xbit_r218_c21 bl[21] br[21] wl[218] vdd gnd cell_6t
Xbit_r219_c21 bl[21] br[21] wl[219] vdd gnd cell_6t
Xbit_r220_c21 bl[21] br[21] wl[220] vdd gnd cell_6t
Xbit_r221_c21 bl[21] br[21] wl[221] vdd gnd cell_6t
Xbit_r222_c21 bl[21] br[21] wl[222] vdd gnd cell_6t
Xbit_r223_c21 bl[21] br[21] wl[223] vdd gnd cell_6t
Xbit_r224_c21 bl[21] br[21] wl[224] vdd gnd cell_6t
Xbit_r225_c21 bl[21] br[21] wl[225] vdd gnd cell_6t
Xbit_r226_c21 bl[21] br[21] wl[226] vdd gnd cell_6t
Xbit_r227_c21 bl[21] br[21] wl[227] vdd gnd cell_6t
Xbit_r228_c21 bl[21] br[21] wl[228] vdd gnd cell_6t
Xbit_r229_c21 bl[21] br[21] wl[229] vdd gnd cell_6t
Xbit_r230_c21 bl[21] br[21] wl[230] vdd gnd cell_6t
Xbit_r231_c21 bl[21] br[21] wl[231] vdd gnd cell_6t
Xbit_r232_c21 bl[21] br[21] wl[232] vdd gnd cell_6t
Xbit_r233_c21 bl[21] br[21] wl[233] vdd gnd cell_6t
Xbit_r234_c21 bl[21] br[21] wl[234] vdd gnd cell_6t
Xbit_r235_c21 bl[21] br[21] wl[235] vdd gnd cell_6t
Xbit_r236_c21 bl[21] br[21] wl[236] vdd gnd cell_6t
Xbit_r237_c21 bl[21] br[21] wl[237] vdd gnd cell_6t
Xbit_r238_c21 bl[21] br[21] wl[238] vdd gnd cell_6t
Xbit_r239_c21 bl[21] br[21] wl[239] vdd gnd cell_6t
Xbit_r240_c21 bl[21] br[21] wl[240] vdd gnd cell_6t
Xbit_r241_c21 bl[21] br[21] wl[241] vdd gnd cell_6t
Xbit_r242_c21 bl[21] br[21] wl[242] vdd gnd cell_6t
Xbit_r243_c21 bl[21] br[21] wl[243] vdd gnd cell_6t
Xbit_r244_c21 bl[21] br[21] wl[244] vdd gnd cell_6t
Xbit_r245_c21 bl[21] br[21] wl[245] vdd gnd cell_6t
Xbit_r246_c21 bl[21] br[21] wl[246] vdd gnd cell_6t
Xbit_r247_c21 bl[21] br[21] wl[247] vdd gnd cell_6t
Xbit_r248_c21 bl[21] br[21] wl[248] vdd gnd cell_6t
Xbit_r249_c21 bl[21] br[21] wl[249] vdd gnd cell_6t
Xbit_r250_c21 bl[21] br[21] wl[250] vdd gnd cell_6t
Xbit_r251_c21 bl[21] br[21] wl[251] vdd gnd cell_6t
Xbit_r252_c21 bl[21] br[21] wl[252] vdd gnd cell_6t
Xbit_r253_c21 bl[21] br[21] wl[253] vdd gnd cell_6t
Xbit_r254_c21 bl[21] br[21] wl[254] vdd gnd cell_6t
Xbit_r255_c21 bl[21] br[21] wl[255] vdd gnd cell_6t
Xbit_r0_c22 bl[22] br[22] wl[0] vdd gnd cell_6t
Xbit_r1_c22 bl[22] br[22] wl[1] vdd gnd cell_6t
Xbit_r2_c22 bl[22] br[22] wl[2] vdd gnd cell_6t
Xbit_r3_c22 bl[22] br[22] wl[3] vdd gnd cell_6t
Xbit_r4_c22 bl[22] br[22] wl[4] vdd gnd cell_6t
Xbit_r5_c22 bl[22] br[22] wl[5] vdd gnd cell_6t
Xbit_r6_c22 bl[22] br[22] wl[6] vdd gnd cell_6t
Xbit_r7_c22 bl[22] br[22] wl[7] vdd gnd cell_6t
Xbit_r8_c22 bl[22] br[22] wl[8] vdd gnd cell_6t
Xbit_r9_c22 bl[22] br[22] wl[9] vdd gnd cell_6t
Xbit_r10_c22 bl[22] br[22] wl[10] vdd gnd cell_6t
Xbit_r11_c22 bl[22] br[22] wl[11] vdd gnd cell_6t
Xbit_r12_c22 bl[22] br[22] wl[12] vdd gnd cell_6t
Xbit_r13_c22 bl[22] br[22] wl[13] vdd gnd cell_6t
Xbit_r14_c22 bl[22] br[22] wl[14] vdd gnd cell_6t
Xbit_r15_c22 bl[22] br[22] wl[15] vdd gnd cell_6t
Xbit_r16_c22 bl[22] br[22] wl[16] vdd gnd cell_6t
Xbit_r17_c22 bl[22] br[22] wl[17] vdd gnd cell_6t
Xbit_r18_c22 bl[22] br[22] wl[18] vdd gnd cell_6t
Xbit_r19_c22 bl[22] br[22] wl[19] vdd gnd cell_6t
Xbit_r20_c22 bl[22] br[22] wl[20] vdd gnd cell_6t
Xbit_r21_c22 bl[22] br[22] wl[21] vdd gnd cell_6t
Xbit_r22_c22 bl[22] br[22] wl[22] vdd gnd cell_6t
Xbit_r23_c22 bl[22] br[22] wl[23] vdd gnd cell_6t
Xbit_r24_c22 bl[22] br[22] wl[24] vdd gnd cell_6t
Xbit_r25_c22 bl[22] br[22] wl[25] vdd gnd cell_6t
Xbit_r26_c22 bl[22] br[22] wl[26] vdd gnd cell_6t
Xbit_r27_c22 bl[22] br[22] wl[27] vdd gnd cell_6t
Xbit_r28_c22 bl[22] br[22] wl[28] vdd gnd cell_6t
Xbit_r29_c22 bl[22] br[22] wl[29] vdd gnd cell_6t
Xbit_r30_c22 bl[22] br[22] wl[30] vdd gnd cell_6t
Xbit_r31_c22 bl[22] br[22] wl[31] vdd gnd cell_6t
Xbit_r32_c22 bl[22] br[22] wl[32] vdd gnd cell_6t
Xbit_r33_c22 bl[22] br[22] wl[33] vdd gnd cell_6t
Xbit_r34_c22 bl[22] br[22] wl[34] vdd gnd cell_6t
Xbit_r35_c22 bl[22] br[22] wl[35] vdd gnd cell_6t
Xbit_r36_c22 bl[22] br[22] wl[36] vdd gnd cell_6t
Xbit_r37_c22 bl[22] br[22] wl[37] vdd gnd cell_6t
Xbit_r38_c22 bl[22] br[22] wl[38] vdd gnd cell_6t
Xbit_r39_c22 bl[22] br[22] wl[39] vdd gnd cell_6t
Xbit_r40_c22 bl[22] br[22] wl[40] vdd gnd cell_6t
Xbit_r41_c22 bl[22] br[22] wl[41] vdd gnd cell_6t
Xbit_r42_c22 bl[22] br[22] wl[42] vdd gnd cell_6t
Xbit_r43_c22 bl[22] br[22] wl[43] vdd gnd cell_6t
Xbit_r44_c22 bl[22] br[22] wl[44] vdd gnd cell_6t
Xbit_r45_c22 bl[22] br[22] wl[45] vdd gnd cell_6t
Xbit_r46_c22 bl[22] br[22] wl[46] vdd gnd cell_6t
Xbit_r47_c22 bl[22] br[22] wl[47] vdd gnd cell_6t
Xbit_r48_c22 bl[22] br[22] wl[48] vdd gnd cell_6t
Xbit_r49_c22 bl[22] br[22] wl[49] vdd gnd cell_6t
Xbit_r50_c22 bl[22] br[22] wl[50] vdd gnd cell_6t
Xbit_r51_c22 bl[22] br[22] wl[51] vdd gnd cell_6t
Xbit_r52_c22 bl[22] br[22] wl[52] vdd gnd cell_6t
Xbit_r53_c22 bl[22] br[22] wl[53] vdd gnd cell_6t
Xbit_r54_c22 bl[22] br[22] wl[54] vdd gnd cell_6t
Xbit_r55_c22 bl[22] br[22] wl[55] vdd gnd cell_6t
Xbit_r56_c22 bl[22] br[22] wl[56] vdd gnd cell_6t
Xbit_r57_c22 bl[22] br[22] wl[57] vdd gnd cell_6t
Xbit_r58_c22 bl[22] br[22] wl[58] vdd gnd cell_6t
Xbit_r59_c22 bl[22] br[22] wl[59] vdd gnd cell_6t
Xbit_r60_c22 bl[22] br[22] wl[60] vdd gnd cell_6t
Xbit_r61_c22 bl[22] br[22] wl[61] vdd gnd cell_6t
Xbit_r62_c22 bl[22] br[22] wl[62] vdd gnd cell_6t
Xbit_r63_c22 bl[22] br[22] wl[63] vdd gnd cell_6t
Xbit_r64_c22 bl[22] br[22] wl[64] vdd gnd cell_6t
Xbit_r65_c22 bl[22] br[22] wl[65] vdd gnd cell_6t
Xbit_r66_c22 bl[22] br[22] wl[66] vdd gnd cell_6t
Xbit_r67_c22 bl[22] br[22] wl[67] vdd gnd cell_6t
Xbit_r68_c22 bl[22] br[22] wl[68] vdd gnd cell_6t
Xbit_r69_c22 bl[22] br[22] wl[69] vdd gnd cell_6t
Xbit_r70_c22 bl[22] br[22] wl[70] vdd gnd cell_6t
Xbit_r71_c22 bl[22] br[22] wl[71] vdd gnd cell_6t
Xbit_r72_c22 bl[22] br[22] wl[72] vdd gnd cell_6t
Xbit_r73_c22 bl[22] br[22] wl[73] vdd gnd cell_6t
Xbit_r74_c22 bl[22] br[22] wl[74] vdd gnd cell_6t
Xbit_r75_c22 bl[22] br[22] wl[75] vdd gnd cell_6t
Xbit_r76_c22 bl[22] br[22] wl[76] vdd gnd cell_6t
Xbit_r77_c22 bl[22] br[22] wl[77] vdd gnd cell_6t
Xbit_r78_c22 bl[22] br[22] wl[78] vdd gnd cell_6t
Xbit_r79_c22 bl[22] br[22] wl[79] vdd gnd cell_6t
Xbit_r80_c22 bl[22] br[22] wl[80] vdd gnd cell_6t
Xbit_r81_c22 bl[22] br[22] wl[81] vdd gnd cell_6t
Xbit_r82_c22 bl[22] br[22] wl[82] vdd gnd cell_6t
Xbit_r83_c22 bl[22] br[22] wl[83] vdd gnd cell_6t
Xbit_r84_c22 bl[22] br[22] wl[84] vdd gnd cell_6t
Xbit_r85_c22 bl[22] br[22] wl[85] vdd gnd cell_6t
Xbit_r86_c22 bl[22] br[22] wl[86] vdd gnd cell_6t
Xbit_r87_c22 bl[22] br[22] wl[87] vdd gnd cell_6t
Xbit_r88_c22 bl[22] br[22] wl[88] vdd gnd cell_6t
Xbit_r89_c22 bl[22] br[22] wl[89] vdd gnd cell_6t
Xbit_r90_c22 bl[22] br[22] wl[90] vdd gnd cell_6t
Xbit_r91_c22 bl[22] br[22] wl[91] vdd gnd cell_6t
Xbit_r92_c22 bl[22] br[22] wl[92] vdd gnd cell_6t
Xbit_r93_c22 bl[22] br[22] wl[93] vdd gnd cell_6t
Xbit_r94_c22 bl[22] br[22] wl[94] vdd gnd cell_6t
Xbit_r95_c22 bl[22] br[22] wl[95] vdd gnd cell_6t
Xbit_r96_c22 bl[22] br[22] wl[96] vdd gnd cell_6t
Xbit_r97_c22 bl[22] br[22] wl[97] vdd gnd cell_6t
Xbit_r98_c22 bl[22] br[22] wl[98] vdd gnd cell_6t
Xbit_r99_c22 bl[22] br[22] wl[99] vdd gnd cell_6t
Xbit_r100_c22 bl[22] br[22] wl[100] vdd gnd cell_6t
Xbit_r101_c22 bl[22] br[22] wl[101] vdd gnd cell_6t
Xbit_r102_c22 bl[22] br[22] wl[102] vdd gnd cell_6t
Xbit_r103_c22 bl[22] br[22] wl[103] vdd gnd cell_6t
Xbit_r104_c22 bl[22] br[22] wl[104] vdd gnd cell_6t
Xbit_r105_c22 bl[22] br[22] wl[105] vdd gnd cell_6t
Xbit_r106_c22 bl[22] br[22] wl[106] vdd gnd cell_6t
Xbit_r107_c22 bl[22] br[22] wl[107] vdd gnd cell_6t
Xbit_r108_c22 bl[22] br[22] wl[108] vdd gnd cell_6t
Xbit_r109_c22 bl[22] br[22] wl[109] vdd gnd cell_6t
Xbit_r110_c22 bl[22] br[22] wl[110] vdd gnd cell_6t
Xbit_r111_c22 bl[22] br[22] wl[111] vdd gnd cell_6t
Xbit_r112_c22 bl[22] br[22] wl[112] vdd gnd cell_6t
Xbit_r113_c22 bl[22] br[22] wl[113] vdd gnd cell_6t
Xbit_r114_c22 bl[22] br[22] wl[114] vdd gnd cell_6t
Xbit_r115_c22 bl[22] br[22] wl[115] vdd gnd cell_6t
Xbit_r116_c22 bl[22] br[22] wl[116] vdd gnd cell_6t
Xbit_r117_c22 bl[22] br[22] wl[117] vdd gnd cell_6t
Xbit_r118_c22 bl[22] br[22] wl[118] vdd gnd cell_6t
Xbit_r119_c22 bl[22] br[22] wl[119] vdd gnd cell_6t
Xbit_r120_c22 bl[22] br[22] wl[120] vdd gnd cell_6t
Xbit_r121_c22 bl[22] br[22] wl[121] vdd gnd cell_6t
Xbit_r122_c22 bl[22] br[22] wl[122] vdd gnd cell_6t
Xbit_r123_c22 bl[22] br[22] wl[123] vdd gnd cell_6t
Xbit_r124_c22 bl[22] br[22] wl[124] vdd gnd cell_6t
Xbit_r125_c22 bl[22] br[22] wl[125] vdd gnd cell_6t
Xbit_r126_c22 bl[22] br[22] wl[126] vdd gnd cell_6t
Xbit_r127_c22 bl[22] br[22] wl[127] vdd gnd cell_6t
Xbit_r128_c22 bl[22] br[22] wl[128] vdd gnd cell_6t
Xbit_r129_c22 bl[22] br[22] wl[129] vdd gnd cell_6t
Xbit_r130_c22 bl[22] br[22] wl[130] vdd gnd cell_6t
Xbit_r131_c22 bl[22] br[22] wl[131] vdd gnd cell_6t
Xbit_r132_c22 bl[22] br[22] wl[132] vdd gnd cell_6t
Xbit_r133_c22 bl[22] br[22] wl[133] vdd gnd cell_6t
Xbit_r134_c22 bl[22] br[22] wl[134] vdd gnd cell_6t
Xbit_r135_c22 bl[22] br[22] wl[135] vdd gnd cell_6t
Xbit_r136_c22 bl[22] br[22] wl[136] vdd gnd cell_6t
Xbit_r137_c22 bl[22] br[22] wl[137] vdd gnd cell_6t
Xbit_r138_c22 bl[22] br[22] wl[138] vdd gnd cell_6t
Xbit_r139_c22 bl[22] br[22] wl[139] vdd gnd cell_6t
Xbit_r140_c22 bl[22] br[22] wl[140] vdd gnd cell_6t
Xbit_r141_c22 bl[22] br[22] wl[141] vdd gnd cell_6t
Xbit_r142_c22 bl[22] br[22] wl[142] vdd gnd cell_6t
Xbit_r143_c22 bl[22] br[22] wl[143] vdd gnd cell_6t
Xbit_r144_c22 bl[22] br[22] wl[144] vdd gnd cell_6t
Xbit_r145_c22 bl[22] br[22] wl[145] vdd gnd cell_6t
Xbit_r146_c22 bl[22] br[22] wl[146] vdd gnd cell_6t
Xbit_r147_c22 bl[22] br[22] wl[147] vdd gnd cell_6t
Xbit_r148_c22 bl[22] br[22] wl[148] vdd gnd cell_6t
Xbit_r149_c22 bl[22] br[22] wl[149] vdd gnd cell_6t
Xbit_r150_c22 bl[22] br[22] wl[150] vdd gnd cell_6t
Xbit_r151_c22 bl[22] br[22] wl[151] vdd gnd cell_6t
Xbit_r152_c22 bl[22] br[22] wl[152] vdd gnd cell_6t
Xbit_r153_c22 bl[22] br[22] wl[153] vdd gnd cell_6t
Xbit_r154_c22 bl[22] br[22] wl[154] vdd gnd cell_6t
Xbit_r155_c22 bl[22] br[22] wl[155] vdd gnd cell_6t
Xbit_r156_c22 bl[22] br[22] wl[156] vdd gnd cell_6t
Xbit_r157_c22 bl[22] br[22] wl[157] vdd gnd cell_6t
Xbit_r158_c22 bl[22] br[22] wl[158] vdd gnd cell_6t
Xbit_r159_c22 bl[22] br[22] wl[159] vdd gnd cell_6t
Xbit_r160_c22 bl[22] br[22] wl[160] vdd gnd cell_6t
Xbit_r161_c22 bl[22] br[22] wl[161] vdd gnd cell_6t
Xbit_r162_c22 bl[22] br[22] wl[162] vdd gnd cell_6t
Xbit_r163_c22 bl[22] br[22] wl[163] vdd gnd cell_6t
Xbit_r164_c22 bl[22] br[22] wl[164] vdd gnd cell_6t
Xbit_r165_c22 bl[22] br[22] wl[165] vdd gnd cell_6t
Xbit_r166_c22 bl[22] br[22] wl[166] vdd gnd cell_6t
Xbit_r167_c22 bl[22] br[22] wl[167] vdd gnd cell_6t
Xbit_r168_c22 bl[22] br[22] wl[168] vdd gnd cell_6t
Xbit_r169_c22 bl[22] br[22] wl[169] vdd gnd cell_6t
Xbit_r170_c22 bl[22] br[22] wl[170] vdd gnd cell_6t
Xbit_r171_c22 bl[22] br[22] wl[171] vdd gnd cell_6t
Xbit_r172_c22 bl[22] br[22] wl[172] vdd gnd cell_6t
Xbit_r173_c22 bl[22] br[22] wl[173] vdd gnd cell_6t
Xbit_r174_c22 bl[22] br[22] wl[174] vdd gnd cell_6t
Xbit_r175_c22 bl[22] br[22] wl[175] vdd gnd cell_6t
Xbit_r176_c22 bl[22] br[22] wl[176] vdd gnd cell_6t
Xbit_r177_c22 bl[22] br[22] wl[177] vdd gnd cell_6t
Xbit_r178_c22 bl[22] br[22] wl[178] vdd gnd cell_6t
Xbit_r179_c22 bl[22] br[22] wl[179] vdd gnd cell_6t
Xbit_r180_c22 bl[22] br[22] wl[180] vdd gnd cell_6t
Xbit_r181_c22 bl[22] br[22] wl[181] vdd gnd cell_6t
Xbit_r182_c22 bl[22] br[22] wl[182] vdd gnd cell_6t
Xbit_r183_c22 bl[22] br[22] wl[183] vdd gnd cell_6t
Xbit_r184_c22 bl[22] br[22] wl[184] vdd gnd cell_6t
Xbit_r185_c22 bl[22] br[22] wl[185] vdd gnd cell_6t
Xbit_r186_c22 bl[22] br[22] wl[186] vdd gnd cell_6t
Xbit_r187_c22 bl[22] br[22] wl[187] vdd gnd cell_6t
Xbit_r188_c22 bl[22] br[22] wl[188] vdd gnd cell_6t
Xbit_r189_c22 bl[22] br[22] wl[189] vdd gnd cell_6t
Xbit_r190_c22 bl[22] br[22] wl[190] vdd gnd cell_6t
Xbit_r191_c22 bl[22] br[22] wl[191] vdd gnd cell_6t
Xbit_r192_c22 bl[22] br[22] wl[192] vdd gnd cell_6t
Xbit_r193_c22 bl[22] br[22] wl[193] vdd gnd cell_6t
Xbit_r194_c22 bl[22] br[22] wl[194] vdd gnd cell_6t
Xbit_r195_c22 bl[22] br[22] wl[195] vdd gnd cell_6t
Xbit_r196_c22 bl[22] br[22] wl[196] vdd gnd cell_6t
Xbit_r197_c22 bl[22] br[22] wl[197] vdd gnd cell_6t
Xbit_r198_c22 bl[22] br[22] wl[198] vdd gnd cell_6t
Xbit_r199_c22 bl[22] br[22] wl[199] vdd gnd cell_6t
Xbit_r200_c22 bl[22] br[22] wl[200] vdd gnd cell_6t
Xbit_r201_c22 bl[22] br[22] wl[201] vdd gnd cell_6t
Xbit_r202_c22 bl[22] br[22] wl[202] vdd gnd cell_6t
Xbit_r203_c22 bl[22] br[22] wl[203] vdd gnd cell_6t
Xbit_r204_c22 bl[22] br[22] wl[204] vdd gnd cell_6t
Xbit_r205_c22 bl[22] br[22] wl[205] vdd gnd cell_6t
Xbit_r206_c22 bl[22] br[22] wl[206] vdd gnd cell_6t
Xbit_r207_c22 bl[22] br[22] wl[207] vdd gnd cell_6t
Xbit_r208_c22 bl[22] br[22] wl[208] vdd gnd cell_6t
Xbit_r209_c22 bl[22] br[22] wl[209] vdd gnd cell_6t
Xbit_r210_c22 bl[22] br[22] wl[210] vdd gnd cell_6t
Xbit_r211_c22 bl[22] br[22] wl[211] vdd gnd cell_6t
Xbit_r212_c22 bl[22] br[22] wl[212] vdd gnd cell_6t
Xbit_r213_c22 bl[22] br[22] wl[213] vdd gnd cell_6t
Xbit_r214_c22 bl[22] br[22] wl[214] vdd gnd cell_6t
Xbit_r215_c22 bl[22] br[22] wl[215] vdd gnd cell_6t
Xbit_r216_c22 bl[22] br[22] wl[216] vdd gnd cell_6t
Xbit_r217_c22 bl[22] br[22] wl[217] vdd gnd cell_6t
Xbit_r218_c22 bl[22] br[22] wl[218] vdd gnd cell_6t
Xbit_r219_c22 bl[22] br[22] wl[219] vdd gnd cell_6t
Xbit_r220_c22 bl[22] br[22] wl[220] vdd gnd cell_6t
Xbit_r221_c22 bl[22] br[22] wl[221] vdd gnd cell_6t
Xbit_r222_c22 bl[22] br[22] wl[222] vdd gnd cell_6t
Xbit_r223_c22 bl[22] br[22] wl[223] vdd gnd cell_6t
Xbit_r224_c22 bl[22] br[22] wl[224] vdd gnd cell_6t
Xbit_r225_c22 bl[22] br[22] wl[225] vdd gnd cell_6t
Xbit_r226_c22 bl[22] br[22] wl[226] vdd gnd cell_6t
Xbit_r227_c22 bl[22] br[22] wl[227] vdd gnd cell_6t
Xbit_r228_c22 bl[22] br[22] wl[228] vdd gnd cell_6t
Xbit_r229_c22 bl[22] br[22] wl[229] vdd gnd cell_6t
Xbit_r230_c22 bl[22] br[22] wl[230] vdd gnd cell_6t
Xbit_r231_c22 bl[22] br[22] wl[231] vdd gnd cell_6t
Xbit_r232_c22 bl[22] br[22] wl[232] vdd gnd cell_6t
Xbit_r233_c22 bl[22] br[22] wl[233] vdd gnd cell_6t
Xbit_r234_c22 bl[22] br[22] wl[234] vdd gnd cell_6t
Xbit_r235_c22 bl[22] br[22] wl[235] vdd gnd cell_6t
Xbit_r236_c22 bl[22] br[22] wl[236] vdd gnd cell_6t
Xbit_r237_c22 bl[22] br[22] wl[237] vdd gnd cell_6t
Xbit_r238_c22 bl[22] br[22] wl[238] vdd gnd cell_6t
Xbit_r239_c22 bl[22] br[22] wl[239] vdd gnd cell_6t
Xbit_r240_c22 bl[22] br[22] wl[240] vdd gnd cell_6t
Xbit_r241_c22 bl[22] br[22] wl[241] vdd gnd cell_6t
Xbit_r242_c22 bl[22] br[22] wl[242] vdd gnd cell_6t
Xbit_r243_c22 bl[22] br[22] wl[243] vdd gnd cell_6t
Xbit_r244_c22 bl[22] br[22] wl[244] vdd gnd cell_6t
Xbit_r245_c22 bl[22] br[22] wl[245] vdd gnd cell_6t
Xbit_r246_c22 bl[22] br[22] wl[246] vdd gnd cell_6t
Xbit_r247_c22 bl[22] br[22] wl[247] vdd gnd cell_6t
Xbit_r248_c22 bl[22] br[22] wl[248] vdd gnd cell_6t
Xbit_r249_c22 bl[22] br[22] wl[249] vdd gnd cell_6t
Xbit_r250_c22 bl[22] br[22] wl[250] vdd gnd cell_6t
Xbit_r251_c22 bl[22] br[22] wl[251] vdd gnd cell_6t
Xbit_r252_c22 bl[22] br[22] wl[252] vdd gnd cell_6t
Xbit_r253_c22 bl[22] br[22] wl[253] vdd gnd cell_6t
Xbit_r254_c22 bl[22] br[22] wl[254] vdd gnd cell_6t
Xbit_r255_c22 bl[22] br[22] wl[255] vdd gnd cell_6t
Xbit_r0_c23 bl[23] br[23] wl[0] vdd gnd cell_6t
Xbit_r1_c23 bl[23] br[23] wl[1] vdd gnd cell_6t
Xbit_r2_c23 bl[23] br[23] wl[2] vdd gnd cell_6t
Xbit_r3_c23 bl[23] br[23] wl[3] vdd gnd cell_6t
Xbit_r4_c23 bl[23] br[23] wl[4] vdd gnd cell_6t
Xbit_r5_c23 bl[23] br[23] wl[5] vdd gnd cell_6t
Xbit_r6_c23 bl[23] br[23] wl[6] vdd gnd cell_6t
Xbit_r7_c23 bl[23] br[23] wl[7] vdd gnd cell_6t
Xbit_r8_c23 bl[23] br[23] wl[8] vdd gnd cell_6t
Xbit_r9_c23 bl[23] br[23] wl[9] vdd gnd cell_6t
Xbit_r10_c23 bl[23] br[23] wl[10] vdd gnd cell_6t
Xbit_r11_c23 bl[23] br[23] wl[11] vdd gnd cell_6t
Xbit_r12_c23 bl[23] br[23] wl[12] vdd gnd cell_6t
Xbit_r13_c23 bl[23] br[23] wl[13] vdd gnd cell_6t
Xbit_r14_c23 bl[23] br[23] wl[14] vdd gnd cell_6t
Xbit_r15_c23 bl[23] br[23] wl[15] vdd gnd cell_6t
Xbit_r16_c23 bl[23] br[23] wl[16] vdd gnd cell_6t
Xbit_r17_c23 bl[23] br[23] wl[17] vdd gnd cell_6t
Xbit_r18_c23 bl[23] br[23] wl[18] vdd gnd cell_6t
Xbit_r19_c23 bl[23] br[23] wl[19] vdd gnd cell_6t
Xbit_r20_c23 bl[23] br[23] wl[20] vdd gnd cell_6t
Xbit_r21_c23 bl[23] br[23] wl[21] vdd gnd cell_6t
Xbit_r22_c23 bl[23] br[23] wl[22] vdd gnd cell_6t
Xbit_r23_c23 bl[23] br[23] wl[23] vdd gnd cell_6t
Xbit_r24_c23 bl[23] br[23] wl[24] vdd gnd cell_6t
Xbit_r25_c23 bl[23] br[23] wl[25] vdd gnd cell_6t
Xbit_r26_c23 bl[23] br[23] wl[26] vdd gnd cell_6t
Xbit_r27_c23 bl[23] br[23] wl[27] vdd gnd cell_6t
Xbit_r28_c23 bl[23] br[23] wl[28] vdd gnd cell_6t
Xbit_r29_c23 bl[23] br[23] wl[29] vdd gnd cell_6t
Xbit_r30_c23 bl[23] br[23] wl[30] vdd gnd cell_6t
Xbit_r31_c23 bl[23] br[23] wl[31] vdd gnd cell_6t
Xbit_r32_c23 bl[23] br[23] wl[32] vdd gnd cell_6t
Xbit_r33_c23 bl[23] br[23] wl[33] vdd gnd cell_6t
Xbit_r34_c23 bl[23] br[23] wl[34] vdd gnd cell_6t
Xbit_r35_c23 bl[23] br[23] wl[35] vdd gnd cell_6t
Xbit_r36_c23 bl[23] br[23] wl[36] vdd gnd cell_6t
Xbit_r37_c23 bl[23] br[23] wl[37] vdd gnd cell_6t
Xbit_r38_c23 bl[23] br[23] wl[38] vdd gnd cell_6t
Xbit_r39_c23 bl[23] br[23] wl[39] vdd gnd cell_6t
Xbit_r40_c23 bl[23] br[23] wl[40] vdd gnd cell_6t
Xbit_r41_c23 bl[23] br[23] wl[41] vdd gnd cell_6t
Xbit_r42_c23 bl[23] br[23] wl[42] vdd gnd cell_6t
Xbit_r43_c23 bl[23] br[23] wl[43] vdd gnd cell_6t
Xbit_r44_c23 bl[23] br[23] wl[44] vdd gnd cell_6t
Xbit_r45_c23 bl[23] br[23] wl[45] vdd gnd cell_6t
Xbit_r46_c23 bl[23] br[23] wl[46] vdd gnd cell_6t
Xbit_r47_c23 bl[23] br[23] wl[47] vdd gnd cell_6t
Xbit_r48_c23 bl[23] br[23] wl[48] vdd gnd cell_6t
Xbit_r49_c23 bl[23] br[23] wl[49] vdd gnd cell_6t
Xbit_r50_c23 bl[23] br[23] wl[50] vdd gnd cell_6t
Xbit_r51_c23 bl[23] br[23] wl[51] vdd gnd cell_6t
Xbit_r52_c23 bl[23] br[23] wl[52] vdd gnd cell_6t
Xbit_r53_c23 bl[23] br[23] wl[53] vdd gnd cell_6t
Xbit_r54_c23 bl[23] br[23] wl[54] vdd gnd cell_6t
Xbit_r55_c23 bl[23] br[23] wl[55] vdd gnd cell_6t
Xbit_r56_c23 bl[23] br[23] wl[56] vdd gnd cell_6t
Xbit_r57_c23 bl[23] br[23] wl[57] vdd gnd cell_6t
Xbit_r58_c23 bl[23] br[23] wl[58] vdd gnd cell_6t
Xbit_r59_c23 bl[23] br[23] wl[59] vdd gnd cell_6t
Xbit_r60_c23 bl[23] br[23] wl[60] vdd gnd cell_6t
Xbit_r61_c23 bl[23] br[23] wl[61] vdd gnd cell_6t
Xbit_r62_c23 bl[23] br[23] wl[62] vdd gnd cell_6t
Xbit_r63_c23 bl[23] br[23] wl[63] vdd gnd cell_6t
Xbit_r64_c23 bl[23] br[23] wl[64] vdd gnd cell_6t
Xbit_r65_c23 bl[23] br[23] wl[65] vdd gnd cell_6t
Xbit_r66_c23 bl[23] br[23] wl[66] vdd gnd cell_6t
Xbit_r67_c23 bl[23] br[23] wl[67] vdd gnd cell_6t
Xbit_r68_c23 bl[23] br[23] wl[68] vdd gnd cell_6t
Xbit_r69_c23 bl[23] br[23] wl[69] vdd gnd cell_6t
Xbit_r70_c23 bl[23] br[23] wl[70] vdd gnd cell_6t
Xbit_r71_c23 bl[23] br[23] wl[71] vdd gnd cell_6t
Xbit_r72_c23 bl[23] br[23] wl[72] vdd gnd cell_6t
Xbit_r73_c23 bl[23] br[23] wl[73] vdd gnd cell_6t
Xbit_r74_c23 bl[23] br[23] wl[74] vdd gnd cell_6t
Xbit_r75_c23 bl[23] br[23] wl[75] vdd gnd cell_6t
Xbit_r76_c23 bl[23] br[23] wl[76] vdd gnd cell_6t
Xbit_r77_c23 bl[23] br[23] wl[77] vdd gnd cell_6t
Xbit_r78_c23 bl[23] br[23] wl[78] vdd gnd cell_6t
Xbit_r79_c23 bl[23] br[23] wl[79] vdd gnd cell_6t
Xbit_r80_c23 bl[23] br[23] wl[80] vdd gnd cell_6t
Xbit_r81_c23 bl[23] br[23] wl[81] vdd gnd cell_6t
Xbit_r82_c23 bl[23] br[23] wl[82] vdd gnd cell_6t
Xbit_r83_c23 bl[23] br[23] wl[83] vdd gnd cell_6t
Xbit_r84_c23 bl[23] br[23] wl[84] vdd gnd cell_6t
Xbit_r85_c23 bl[23] br[23] wl[85] vdd gnd cell_6t
Xbit_r86_c23 bl[23] br[23] wl[86] vdd gnd cell_6t
Xbit_r87_c23 bl[23] br[23] wl[87] vdd gnd cell_6t
Xbit_r88_c23 bl[23] br[23] wl[88] vdd gnd cell_6t
Xbit_r89_c23 bl[23] br[23] wl[89] vdd gnd cell_6t
Xbit_r90_c23 bl[23] br[23] wl[90] vdd gnd cell_6t
Xbit_r91_c23 bl[23] br[23] wl[91] vdd gnd cell_6t
Xbit_r92_c23 bl[23] br[23] wl[92] vdd gnd cell_6t
Xbit_r93_c23 bl[23] br[23] wl[93] vdd gnd cell_6t
Xbit_r94_c23 bl[23] br[23] wl[94] vdd gnd cell_6t
Xbit_r95_c23 bl[23] br[23] wl[95] vdd gnd cell_6t
Xbit_r96_c23 bl[23] br[23] wl[96] vdd gnd cell_6t
Xbit_r97_c23 bl[23] br[23] wl[97] vdd gnd cell_6t
Xbit_r98_c23 bl[23] br[23] wl[98] vdd gnd cell_6t
Xbit_r99_c23 bl[23] br[23] wl[99] vdd gnd cell_6t
Xbit_r100_c23 bl[23] br[23] wl[100] vdd gnd cell_6t
Xbit_r101_c23 bl[23] br[23] wl[101] vdd gnd cell_6t
Xbit_r102_c23 bl[23] br[23] wl[102] vdd gnd cell_6t
Xbit_r103_c23 bl[23] br[23] wl[103] vdd gnd cell_6t
Xbit_r104_c23 bl[23] br[23] wl[104] vdd gnd cell_6t
Xbit_r105_c23 bl[23] br[23] wl[105] vdd gnd cell_6t
Xbit_r106_c23 bl[23] br[23] wl[106] vdd gnd cell_6t
Xbit_r107_c23 bl[23] br[23] wl[107] vdd gnd cell_6t
Xbit_r108_c23 bl[23] br[23] wl[108] vdd gnd cell_6t
Xbit_r109_c23 bl[23] br[23] wl[109] vdd gnd cell_6t
Xbit_r110_c23 bl[23] br[23] wl[110] vdd gnd cell_6t
Xbit_r111_c23 bl[23] br[23] wl[111] vdd gnd cell_6t
Xbit_r112_c23 bl[23] br[23] wl[112] vdd gnd cell_6t
Xbit_r113_c23 bl[23] br[23] wl[113] vdd gnd cell_6t
Xbit_r114_c23 bl[23] br[23] wl[114] vdd gnd cell_6t
Xbit_r115_c23 bl[23] br[23] wl[115] vdd gnd cell_6t
Xbit_r116_c23 bl[23] br[23] wl[116] vdd gnd cell_6t
Xbit_r117_c23 bl[23] br[23] wl[117] vdd gnd cell_6t
Xbit_r118_c23 bl[23] br[23] wl[118] vdd gnd cell_6t
Xbit_r119_c23 bl[23] br[23] wl[119] vdd gnd cell_6t
Xbit_r120_c23 bl[23] br[23] wl[120] vdd gnd cell_6t
Xbit_r121_c23 bl[23] br[23] wl[121] vdd gnd cell_6t
Xbit_r122_c23 bl[23] br[23] wl[122] vdd gnd cell_6t
Xbit_r123_c23 bl[23] br[23] wl[123] vdd gnd cell_6t
Xbit_r124_c23 bl[23] br[23] wl[124] vdd gnd cell_6t
Xbit_r125_c23 bl[23] br[23] wl[125] vdd gnd cell_6t
Xbit_r126_c23 bl[23] br[23] wl[126] vdd gnd cell_6t
Xbit_r127_c23 bl[23] br[23] wl[127] vdd gnd cell_6t
Xbit_r128_c23 bl[23] br[23] wl[128] vdd gnd cell_6t
Xbit_r129_c23 bl[23] br[23] wl[129] vdd gnd cell_6t
Xbit_r130_c23 bl[23] br[23] wl[130] vdd gnd cell_6t
Xbit_r131_c23 bl[23] br[23] wl[131] vdd gnd cell_6t
Xbit_r132_c23 bl[23] br[23] wl[132] vdd gnd cell_6t
Xbit_r133_c23 bl[23] br[23] wl[133] vdd gnd cell_6t
Xbit_r134_c23 bl[23] br[23] wl[134] vdd gnd cell_6t
Xbit_r135_c23 bl[23] br[23] wl[135] vdd gnd cell_6t
Xbit_r136_c23 bl[23] br[23] wl[136] vdd gnd cell_6t
Xbit_r137_c23 bl[23] br[23] wl[137] vdd gnd cell_6t
Xbit_r138_c23 bl[23] br[23] wl[138] vdd gnd cell_6t
Xbit_r139_c23 bl[23] br[23] wl[139] vdd gnd cell_6t
Xbit_r140_c23 bl[23] br[23] wl[140] vdd gnd cell_6t
Xbit_r141_c23 bl[23] br[23] wl[141] vdd gnd cell_6t
Xbit_r142_c23 bl[23] br[23] wl[142] vdd gnd cell_6t
Xbit_r143_c23 bl[23] br[23] wl[143] vdd gnd cell_6t
Xbit_r144_c23 bl[23] br[23] wl[144] vdd gnd cell_6t
Xbit_r145_c23 bl[23] br[23] wl[145] vdd gnd cell_6t
Xbit_r146_c23 bl[23] br[23] wl[146] vdd gnd cell_6t
Xbit_r147_c23 bl[23] br[23] wl[147] vdd gnd cell_6t
Xbit_r148_c23 bl[23] br[23] wl[148] vdd gnd cell_6t
Xbit_r149_c23 bl[23] br[23] wl[149] vdd gnd cell_6t
Xbit_r150_c23 bl[23] br[23] wl[150] vdd gnd cell_6t
Xbit_r151_c23 bl[23] br[23] wl[151] vdd gnd cell_6t
Xbit_r152_c23 bl[23] br[23] wl[152] vdd gnd cell_6t
Xbit_r153_c23 bl[23] br[23] wl[153] vdd gnd cell_6t
Xbit_r154_c23 bl[23] br[23] wl[154] vdd gnd cell_6t
Xbit_r155_c23 bl[23] br[23] wl[155] vdd gnd cell_6t
Xbit_r156_c23 bl[23] br[23] wl[156] vdd gnd cell_6t
Xbit_r157_c23 bl[23] br[23] wl[157] vdd gnd cell_6t
Xbit_r158_c23 bl[23] br[23] wl[158] vdd gnd cell_6t
Xbit_r159_c23 bl[23] br[23] wl[159] vdd gnd cell_6t
Xbit_r160_c23 bl[23] br[23] wl[160] vdd gnd cell_6t
Xbit_r161_c23 bl[23] br[23] wl[161] vdd gnd cell_6t
Xbit_r162_c23 bl[23] br[23] wl[162] vdd gnd cell_6t
Xbit_r163_c23 bl[23] br[23] wl[163] vdd gnd cell_6t
Xbit_r164_c23 bl[23] br[23] wl[164] vdd gnd cell_6t
Xbit_r165_c23 bl[23] br[23] wl[165] vdd gnd cell_6t
Xbit_r166_c23 bl[23] br[23] wl[166] vdd gnd cell_6t
Xbit_r167_c23 bl[23] br[23] wl[167] vdd gnd cell_6t
Xbit_r168_c23 bl[23] br[23] wl[168] vdd gnd cell_6t
Xbit_r169_c23 bl[23] br[23] wl[169] vdd gnd cell_6t
Xbit_r170_c23 bl[23] br[23] wl[170] vdd gnd cell_6t
Xbit_r171_c23 bl[23] br[23] wl[171] vdd gnd cell_6t
Xbit_r172_c23 bl[23] br[23] wl[172] vdd gnd cell_6t
Xbit_r173_c23 bl[23] br[23] wl[173] vdd gnd cell_6t
Xbit_r174_c23 bl[23] br[23] wl[174] vdd gnd cell_6t
Xbit_r175_c23 bl[23] br[23] wl[175] vdd gnd cell_6t
Xbit_r176_c23 bl[23] br[23] wl[176] vdd gnd cell_6t
Xbit_r177_c23 bl[23] br[23] wl[177] vdd gnd cell_6t
Xbit_r178_c23 bl[23] br[23] wl[178] vdd gnd cell_6t
Xbit_r179_c23 bl[23] br[23] wl[179] vdd gnd cell_6t
Xbit_r180_c23 bl[23] br[23] wl[180] vdd gnd cell_6t
Xbit_r181_c23 bl[23] br[23] wl[181] vdd gnd cell_6t
Xbit_r182_c23 bl[23] br[23] wl[182] vdd gnd cell_6t
Xbit_r183_c23 bl[23] br[23] wl[183] vdd gnd cell_6t
Xbit_r184_c23 bl[23] br[23] wl[184] vdd gnd cell_6t
Xbit_r185_c23 bl[23] br[23] wl[185] vdd gnd cell_6t
Xbit_r186_c23 bl[23] br[23] wl[186] vdd gnd cell_6t
Xbit_r187_c23 bl[23] br[23] wl[187] vdd gnd cell_6t
Xbit_r188_c23 bl[23] br[23] wl[188] vdd gnd cell_6t
Xbit_r189_c23 bl[23] br[23] wl[189] vdd gnd cell_6t
Xbit_r190_c23 bl[23] br[23] wl[190] vdd gnd cell_6t
Xbit_r191_c23 bl[23] br[23] wl[191] vdd gnd cell_6t
Xbit_r192_c23 bl[23] br[23] wl[192] vdd gnd cell_6t
Xbit_r193_c23 bl[23] br[23] wl[193] vdd gnd cell_6t
Xbit_r194_c23 bl[23] br[23] wl[194] vdd gnd cell_6t
Xbit_r195_c23 bl[23] br[23] wl[195] vdd gnd cell_6t
Xbit_r196_c23 bl[23] br[23] wl[196] vdd gnd cell_6t
Xbit_r197_c23 bl[23] br[23] wl[197] vdd gnd cell_6t
Xbit_r198_c23 bl[23] br[23] wl[198] vdd gnd cell_6t
Xbit_r199_c23 bl[23] br[23] wl[199] vdd gnd cell_6t
Xbit_r200_c23 bl[23] br[23] wl[200] vdd gnd cell_6t
Xbit_r201_c23 bl[23] br[23] wl[201] vdd gnd cell_6t
Xbit_r202_c23 bl[23] br[23] wl[202] vdd gnd cell_6t
Xbit_r203_c23 bl[23] br[23] wl[203] vdd gnd cell_6t
Xbit_r204_c23 bl[23] br[23] wl[204] vdd gnd cell_6t
Xbit_r205_c23 bl[23] br[23] wl[205] vdd gnd cell_6t
Xbit_r206_c23 bl[23] br[23] wl[206] vdd gnd cell_6t
Xbit_r207_c23 bl[23] br[23] wl[207] vdd gnd cell_6t
Xbit_r208_c23 bl[23] br[23] wl[208] vdd gnd cell_6t
Xbit_r209_c23 bl[23] br[23] wl[209] vdd gnd cell_6t
Xbit_r210_c23 bl[23] br[23] wl[210] vdd gnd cell_6t
Xbit_r211_c23 bl[23] br[23] wl[211] vdd gnd cell_6t
Xbit_r212_c23 bl[23] br[23] wl[212] vdd gnd cell_6t
Xbit_r213_c23 bl[23] br[23] wl[213] vdd gnd cell_6t
Xbit_r214_c23 bl[23] br[23] wl[214] vdd gnd cell_6t
Xbit_r215_c23 bl[23] br[23] wl[215] vdd gnd cell_6t
Xbit_r216_c23 bl[23] br[23] wl[216] vdd gnd cell_6t
Xbit_r217_c23 bl[23] br[23] wl[217] vdd gnd cell_6t
Xbit_r218_c23 bl[23] br[23] wl[218] vdd gnd cell_6t
Xbit_r219_c23 bl[23] br[23] wl[219] vdd gnd cell_6t
Xbit_r220_c23 bl[23] br[23] wl[220] vdd gnd cell_6t
Xbit_r221_c23 bl[23] br[23] wl[221] vdd gnd cell_6t
Xbit_r222_c23 bl[23] br[23] wl[222] vdd gnd cell_6t
Xbit_r223_c23 bl[23] br[23] wl[223] vdd gnd cell_6t
Xbit_r224_c23 bl[23] br[23] wl[224] vdd gnd cell_6t
Xbit_r225_c23 bl[23] br[23] wl[225] vdd gnd cell_6t
Xbit_r226_c23 bl[23] br[23] wl[226] vdd gnd cell_6t
Xbit_r227_c23 bl[23] br[23] wl[227] vdd gnd cell_6t
Xbit_r228_c23 bl[23] br[23] wl[228] vdd gnd cell_6t
Xbit_r229_c23 bl[23] br[23] wl[229] vdd gnd cell_6t
Xbit_r230_c23 bl[23] br[23] wl[230] vdd gnd cell_6t
Xbit_r231_c23 bl[23] br[23] wl[231] vdd gnd cell_6t
Xbit_r232_c23 bl[23] br[23] wl[232] vdd gnd cell_6t
Xbit_r233_c23 bl[23] br[23] wl[233] vdd gnd cell_6t
Xbit_r234_c23 bl[23] br[23] wl[234] vdd gnd cell_6t
Xbit_r235_c23 bl[23] br[23] wl[235] vdd gnd cell_6t
Xbit_r236_c23 bl[23] br[23] wl[236] vdd gnd cell_6t
Xbit_r237_c23 bl[23] br[23] wl[237] vdd gnd cell_6t
Xbit_r238_c23 bl[23] br[23] wl[238] vdd gnd cell_6t
Xbit_r239_c23 bl[23] br[23] wl[239] vdd gnd cell_6t
Xbit_r240_c23 bl[23] br[23] wl[240] vdd gnd cell_6t
Xbit_r241_c23 bl[23] br[23] wl[241] vdd gnd cell_6t
Xbit_r242_c23 bl[23] br[23] wl[242] vdd gnd cell_6t
Xbit_r243_c23 bl[23] br[23] wl[243] vdd gnd cell_6t
Xbit_r244_c23 bl[23] br[23] wl[244] vdd gnd cell_6t
Xbit_r245_c23 bl[23] br[23] wl[245] vdd gnd cell_6t
Xbit_r246_c23 bl[23] br[23] wl[246] vdd gnd cell_6t
Xbit_r247_c23 bl[23] br[23] wl[247] vdd gnd cell_6t
Xbit_r248_c23 bl[23] br[23] wl[248] vdd gnd cell_6t
Xbit_r249_c23 bl[23] br[23] wl[249] vdd gnd cell_6t
Xbit_r250_c23 bl[23] br[23] wl[250] vdd gnd cell_6t
Xbit_r251_c23 bl[23] br[23] wl[251] vdd gnd cell_6t
Xbit_r252_c23 bl[23] br[23] wl[252] vdd gnd cell_6t
Xbit_r253_c23 bl[23] br[23] wl[253] vdd gnd cell_6t
Xbit_r254_c23 bl[23] br[23] wl[254] vdd gnd cell_6t
Xbit_r255_c23 bl[23] br[23] wl[255] vdd gnd cell_6t
Xbit_r0_c24 bl[24] br[24] wl[0] vdd gnd cell_6t
Xbit_r1_c24 bl[24] br[24] wl[1] vdd gnd cell_6t
Xbit_r2_c24 bl[24] br[24] wl[2] vdd gnd cell_6t
Xbit_r3_c24 bl[24] br[24] wl[3] vdd gnd cell_6t
Xbit_r4_c24 bl[24] br[24] wl[4] vdd gnd cell_6t
Xbit_r5_c24 bl[24] br[24] wl[5] vdd gnd cell_6t
Xbit_r6_c24 bl[24] br[24] wl[6] vdd gnd cell_6t
Xbit_r7_c24 bl[24] br[24] wl[7] vdd gnd cell_6t
Xbit_r8_c24 bl[24] br[24] wl[8] vdd gnd cell_6t
Xbit_r9_c24 bl[24] br[24] wl[9] vdd gnd cell_6t
Xbit_r10_c24 bl[24] br[24] wl[10] vdd gnd cell_6t
Xbit_r11_c24 bl[24] br[24] wl[11] vdd gnd cell_6t
Xbit_r12_c24 bl[24] br[24] wl[12] vdd gnd cell_6t
Xbit_r13_c24 bl[24] br[24] wl[13] vdd gnd cell_6t
Xbit_r14_c24 bl[24] br[24] wl[14] vdd gnd cell_6t
Xbit_r15_c24 bl[24] br[24] wl[15] vdd gnd cell_6t
Xbit_r16_c24 bl[24] br[24] wl[16] vdd gnd cell_6t
Xbit_r17_c24 bl[24] br[24] wl[17] vdd gnd cell_6t
Xbit_r18_c24 bl[24] br[24] wl[18] vdd gnd cell_6t
Xbit_r19_c24 bl[24] br[24] wl[19] vdd gnd cell_6t
Xbit_r20_c24 bl[24] br[24] wl[20] vdd gnd cell_6t
Xbit_r21_c24 bl[24] br[24] wl[21] vdd gnd cell_6t
Xbit_r22_c24 bl[24] br[24] wl[22] vdd gnd cell_6t
Xbit_r23_c24 bl[24] br[24] wl[23] vdd gnd cell_6t
Xbit_r24_c24 bl[24] br[24] wl[24] vdd gnd cell_6t
Xbit_r25_c24 bl[24] br[24] wl[25] vdd gnd cell_6t
Xbit_r26_c24 bl[24] br[24] wl[26] vdd gnd cell_6t
Xbit_r27_c24 bl[24] br[24] wl[27] vdd gnd cell_6t
Xbit_r28_c24 bl[24] br[24] wl[28] vdd gnd cell_6t
Xbit_r29_c24 bl[24] br[24] wl[29] vdd gnd cell_6t
Xbit_r30_c24 bl[24] br[24] wl[30] vdd gnd cell_6t
Xbit_r31_c24 bl[24] br[24] wl[31] vdd gnd cell_6t
Xbit_r32_c24 bl[24] br[24] wl[32] vdd gnd cell_6t
Xbit_r33_c24 bl[24] br[24] wl[33] vdd gnd cell_6t
Xbit_r34_c24 bl[24] br[24] wl[34] vdd gnd cell_6t
Xbit_r35_c24 bl[24] br[24] wl[35] vdd gnd cell_6t
Xbit_r36_c24 bl[24] br[24] wl[36] vdd gnd cell_6t
Xbit_r37_c24 bl[24] br[24] wl[37] vdd gnd cell_6t
Xbit_r38_c24 bl[24] br[24] wl[38] vdd gnd cell_6t
Xbit_r39_c24 bl[24] br[24] wl[39] vdd gnd cell_6t
Xbit_r40_c24 bl[24] br[24] wl[40] vdd gnd cell_6t
Xbit_r41_c24 bl[24] br[24] wl[41] vdd gnd cell_6t
Xbit_r42_c24 bl[24] br[24] wl[42] vdd gnd cell_6t
Xbit_r43_c24 bl[24] br[24] wl[43] vdd gnd cell_6t
Xbit_r44_c24 bl[24] br[24] wl[44] vdd gnd cell_6t
Xbit_r45_c24 bl[24] br[24] wl[45] vdd gnd cell_6t
Xbit_r46_c24 bl[24] br[24] wl[46] vdd gnd cell_6t
Xbit_r47_c24 bl[24] br[24] wl[47] vdd gnd cell_6t
Xbit_r48_c24 bl[24] br[24] wl[48] vdd gnd cell_6t
Xbit_r49_c24 bl[24] br[24] wl[49] vdd gnd cell_6t
Xbit_r50_c24 bl[24] br[24] wl[50] vdd gnd cell_6t
Xbit_r51_c24 bl[24] br[24] wl[51] vdd gnd cell_6t
Xbit_r52_c24 bl[24] br[24] wl[52] vdd gnd cell_6t
Xbit_r53_c24 bl[24] br[24] wl[53] vdd gnd cell_6t
Xbit_r54_c24 bl[24] br[24] wl[54] vdd gnd cell_6t
Xbit_r55_c24 bl[24] br[24] wl[55] vdd gnd cell_6t
Xbit_r56_c24 bl[24] br[24] wl[56] vdd gnd cell_6t
Xbit_r57_c24 bl[24] br[24] wl[57] vdd gnd cell_6t
Xbit_r58_c24 bl[24] br[24] wl[58] vdd gnd cell_6t
Xbit_r59_c24 bl[24] br[24] wl[59] vdd gnd cell_6t
Xbit_r60_c24 bl[24] br[24] wl[60] vdd gnd cell_6t
Xbit_r61_c24 bl[24] br[24] wl[61] vdd gnd cell_6t
Xbit_r62_c24 bl[24] br[24] wl[62] vdd gnd cell_6t
Xbit_r63_c24 bl[24] br[24] wl[63] vdd gnd cell_6t
Xbit_r64_c24 bl[24] br[24] wl[64] vdd gnd cell_6t
Xbit_r65_c24 bl[24] br[24] wl[65] vdd gnd cell_6t
Xbit_r66_c24 bl[24] br[24] wl[66] vdd gnd cell_6t
Xbit_r67_c24 bl[24] br[24] wl[67] vdd gnd cell_6t
Xbit_r68_c24 bl[24] br[24] wl[68] vdd gnd cell_6t
Xbit_r69_c24 bl[24] br[24] wl[69] vdd gnd cell_6t
Xbit_r70_c24 bl[24] br[24] wl[70] vdd gnd cell_6t
Xbit_r71_c24 bl[24] br[24] wl[71] vdd gnd cell_6t
Xbit_r72_c24 bl[24] br[24] wl[72] vdd gnd cell_6t
Xbit_r73_c24 bl[24] br[24] wl[73] vdd gnd cell_6t
Xbit_r74_c24 bl[24] br[24] wl[74] vdd gnd cell_6t
Xbit_r75_c24 bl[24] br[24] wl[75] vdd gnd cell_6t
Xbit_r76_c24 bl[24] br[24] wl[76] vdd gnd cell_6t
Xbit_r77_c24 bl[24] br[24] wl[77] vdd gnd cell_6t
Xbit_r78_c24 bl[24] br[24] wl[78] vdd gnd cell_6t
Xbit_r79_c24 bl[24] br[24] wl[79] vdd gnd cell_6t
Xbit_r80_c24 bl[24] br[24] wl[80] vdd gnd cell_6t
Xbit_r81_c24 bl[24] br[24] wl[81] vdd gnd cell_6t
Xbit_r82_c24 bl[24] br[24] wl[82] vdd gnd cell_6t
Xbit_r83_c24 bl[24] br[24] wl[83] vdd gnd cell_6t
Xbit_r84_c24 bl[24] br[24] wl[84] vdd gnd cell_6t
Xbit_r85_c24 bl[24] br[24] wl[85] vdd gnd cell_6t
Xbit_r86_c24 bl[24] br[24] wl[86] vdd gnd cell_6t
Xbit_r87_c24 bl[24] br[24] wl[87] vdd gnd cell_6t
Xbit_r88_c24 bl[24] br[24] wl[88] vdd gnd cell_6t
Xbit_r89_c24 bl[24] br[24] wl[89] vdd gnd cell_6t
Xbit_r90_c24 bl[24] br[24] wl[90] vdd gnd cell_6t
Xbit_r91_c24 bl[24] br[24] wl[91] vdd gnd cell_6t
Xbit_r92_c24 bl[24] br[24] wl[92] vdd gnd cell_6t
Xbit_r93_c24 bl[24] br[24] wl[93] vdd gnd cell_6t
Xbit_r94_c24 bl[24] br[24] wl[94] vdd gnd cell_6t
Xbit_r95_c24 bl[24] br[24] wl[95] vdd gnd cell_6t
Xbit_r96_c24 bl[24] br[24] wl[96] vdd gnd cell_6t
Xbit_r97_c24 bl[24] br[24] wl[97] vdd gnd cell_6t
Xbit_r98_c24 bl[24] br[24] wl[98] vdd gnd cell_6t
Xbit_r99_c24 bl[24] br[24] wl[99] vdd gnd cell_6t
Xbit_r100_c24 bl[24] br[24] wl[100] vdd gnd cell_6t
Xbit_r101_c24 bl[24] br[24] wl[101] vdd gnd cell_6t
Xbit_r102_c24 bl[24] br[24] wl[102] vdd gnd cell_6t
Xbit_r103_c24 bl[24] br[24] wl[103] vdd gnd cell_6t
Xbit_r104_c24 bl[24] br[24] wl[104] vdd gnd cell_6t
Xbit_r105_c24 bl[24] br[24] wl[105] vdd gnd cell_6t
Xbit_r106_c24 bl[24] br[24] wl[106] vdd gnd cell_6t
Xbit_r107_c24 bl[24] br[24] wl[107] vdd gnd cell_6t
Xbit_r108_c24 bl[24] br[24] wl[108] vdd gnd cell_6t
Xbit_r109_c24 bl[24] br[24] wl[109] vdd gnd cell_6t
Xbit_r110_c24 bl[24] br[24] wl[110] vdd gnd cell_6t
Xbit_r111_c24 bl[24] br[24] wl[111] vdd gnd cell_6t
Xbit_r112_c24 bl[24] br[24] wl[112] vdd gnd cell_6t
Xbit_r113_c24 bl[24] br[24] wl[113] vdd gnd cell_6t
Xbit_r114_c24 bl[24] br[24] wl[114] vdd gnd cell_6t
Xbit_r115_c24 bl[24] br[24] wl[115] vdd gnd cell_6t
Xbit_r116_c24 bl[24] br[24] wl[116] vdd gnd cell_6t
Xbit_r117_c24 bl[24] br[24] wl[117] vdd gnd cell_6t
Xbit_r118_c24 bl[24] br[24] wl[118] vdd gnd cell_6t
Xbit_r119_c24 bl[24] br[24] wl[119] vdd gnd cell_6t
Xbit_r120_c24 bl[24] br[24] wl[120] vdd gnd cell_6t
Xbit_r121_c24 bl[24] br[24] wl[121] vdd gnd cell_6t
Xbit_r122_c24 bl[24] br[24] wl[122] vdd gnd cell_6t
Xbit_r123_c24 bl[24] br[24] wl[123] vdd gnd cell_6t
Xbit_r124_c24 bl[24] br[24] wl[124] vdd gnd cell_6t
Xbit_r125_c24 bl[24] br[24] wl[125] vdd gnd cell_6t
Xbit_r126_c24 bl[24] br[24] wl[126] vdd gnd cell_6t
Xbit_r127_c24 bl[24] br[24] wl[127] vdd gnd cell_6t
Xbit_r128_c24 bl[24] br[24] wl[128] vdd gnd cell_6t
Xbit_r129_c24 bl[24] br[24] wl[129] vdd gnd cell_6t
Xbit_r130_c24 bl[24] br[24] wl[130] vdd gnd cell_6t
Xbit_r131_c24 bl[24] br[24] wl[131] vdd gnd cell_6t
Xbit_r132_c24 bl[24] br[24] wl[132] vdd gnd cell_6t
Xbit_r133_c24 bl[24] br[24] wl[133] vdd gnd cell_6t
Xbit_r134_c24 bl[24] br[24] wl[134] vdd gnd cell_6t
Xbit_r135_c24 bl[24] br[24] wl[135] vdd gnd cell_6t
Xbit_r136_c24 bl[24] br[24] wl[136] vdd gnd cell_6t
Xbit_r137_c24 bl[24] br[24] wl[137] vdd gnd cell_6t
Xbit_r138_c24 bl[24] br[24] wl[138] vdd gnd cell_6t
Xbit_r139_c24 bl[24] br[24] wl[139] vdd gnd cell_6t
Xbit_r140_c24 bl[24] br[24] wl[140] vdd gnd cell_6t
Xbit_r141_c24 bl[24] br[24] wl[141] vdd gnd cell_6t
Xbit_r142_c24 bl[24] br[24] wl[142] vdd gnd cell_6t
Xbit_r143_c24 bl[24] br[24] wl[143] vdd gnd cell_6t
Xbit_r144_c24 bl[24] br[24] wl[144] vdd gnd cell_6t
Xbit_r145_c24 bl[24] br[24] wl[145] vdd gnd cell_6t
Xbit_r146_c24 bl[24] br[24] wl[146] vdd gnd cell_6t
Xbit_r147_c24 bl[24] br[24] wl[147] vdd gnd cell_6t
Xbit_r148_c24 bl[24] br[24] wl[148] vdd gnd cell_6t
Xbit_r149_c24 bl[24] br[24] wl[149] vdd gnd cell_6t
Xbit_r150_c24 bl[24] br[24] wl[150] vdd gnd cell_6t
Xbit_r151_c24 bl[24] br[24] wl[151] vdd gnd cell_6t
Xbit_r152_c24 bl[24] br[24] wl[152] vdd gnd cell_6t
Xbit_r153_c24 bl[24] br[24] wl[153] vdd gnd cell_6t
Xbit_r154_c24 bl[24] br[24] wl[154] vdd gnd cell_6t
Xbit_r155_c24 bl[24] br[24] wl[155] vdd gnd cell_6t
Xbit_r156_c24 bl[24] br[24] wl[156] vdd gnd cell_6t
Xbit_r157_c24 bl[24] br[24] wl[157] vdd gnd cell_6t
Xbit_r158_c24 bl[24] br[24] wl[158] vdd gnd cell_6t
Xbit_r159_c24 bl[24] br[24] wl[159] vdd gnd cell_6t
Xbit_r160_c24 bl[24] br[24] wl[160] vdd gnd cell_6t
Xbit_r161_c24 bl[24] br[24] wl[161] vdd gnd cell_6t
Xbit_r162_c24 bl[24] br[24] wl[162] vdd gnd cell_6t
Xbit_r163_c24 bl[24] br[24] wl[163] vdd gnd cell_6t
Xbit_r164_c24 bl[24] br[24] wl[164] vdd gnd cell_6t
Xbit_r165_c24 bl[24] br[24] wl[165] vdd gnd cell_6t
Xbit_r166_c24 bl[24] br[24] wl[166] vdd gnd cell_6t
Xbit_r167_c24 bl[24] br[24] wl[167] vdd gnd cell_6t
Xbit_r168_c24 bl[24] br[24] wl[168] vdd gnd cell_6t
Xbit_r169_c24 bl[24] br[24] wl[169] vdd gnd cell_6t
Xbit_r170_c24 bl[24] br[24] wl[170] vdd gnd cell_6t
Xbit_r171_c24 bl[24] br[24] wl[171] vdd gnd cell_6t
Xbit_r172_c24 bl[24] br[24] wl[172] vdd gnd cell_6t
Xbit_r173_c24 bl[24] br[24] wl[173] vdd gnd cell_6t
Xbit_r174_c24 bl[24] br[24] wl[174] vdd gnd cell_6t
Xbit_r175_c24 bl[24] br[24] wl[175] vdd gnd cell_6t
Xbit_r176_c24 bl[24] br[24] wl[176] vdd gnd cell_6t
Xbit_r177_c24 bl[24] br[24] wl[177] vdd gnd cell_6t
Xbit_r178_c24 bl[24] br[24] wl[178] vdd gnd cell_6t
Xbit_r179_c24 bl[24] br[24] wl[179] vdd gnd cell_6t
Xbit_r180_c24 bl[24] br[24] wl[180] vdd gnd cell_6t
Xbit_r181_c24 bl[24] br[24] wl[181] vdd gnd cell_6t
Xbit_r182_c24 bl[24] br[24] wl[182] vdd gnd cell_6t
Xbit_r183_c24 bl[24] br[24] wl[183] vdd gnd cell_6t
Xbit_r184_c24 bl[24] br[24] wl[184] vdd gnd cell_6t
Xbit_r185_c24 bl[24] br[24] wl[185] vdd gnd cell_6t
Xbit_r186_c24 bl[24] br[24] wl[186] vdd gnd cell_6t
Xbit_r187_c24 bl[24] br[24] wl[187] vdd gnd cell_6t
Xbit_r188_c24 bl[24] br[24] wl[188] vdd gnd cell_6t
Xbit_r189_c24 bl[24] br[24] wl[189] vdd gnd cell_6t
Xbit_r190_c24 bl[24] br[24] wl[190] vdd gnd cell_6t
Xbit_r191_c24 bl[24] br[24] wl[191] vdd gnd cell_6t
Xbit_r192_c24 bl[24] br[24] wl[192] vdd gnd cell_6t
Xbit_r193_c24 bl[24] br[24] wl[193] vdd gnd cell_6t
Xbit_r194_c24 bl[24] br[24] wl[194] vdd gnd cell_6t
Xbit_r195_c24 bl[24] br[24] wl[195] vdd gnd cell_6t
Xbit_r196_c24 bl[24] br[24] wl[196] vdd gnd cell_6t
Xbit_r197_c24 bl[24] br[24] wl[197] vdd gnd cell_6t
Xbit_r198_c24 bl[24] br[24] wl[198] vdd gnd cell_6t
Xbit_r199_c24 bl[24] br[24] wl[199] vdd gnd cell_6t
Xbit_r200_c24 bl[24] br[24] wl[200] vdd gnd cell_6t
Xbit_r201_c24 bl[24] br[24] wl[201] vdd gnd cell_6t
Xbit_r202_c24 bl[24] br[24] wl[202] vdd gnd cell_6t
Xbit_r203_c24 bl[24] br[24] wl[203] vdd gnd cell_6t
Xbit_r204_c24 bl[24] br[24] wl[204] vdd gnd cell_6t
Xbit_r205_c24 bl[24] br[24] wl[205] vdd gnd cell_6t
Xbit_r206_c24 bl[24] br[24] wl[206] vdd gnd cell_6t
Xbit_r207_c24 bl[24] br[24] wl[207] vdd gnd cell_6t
Xbit_r208_c24 bl[24] br[24] wl[208] vdd gnd cell_6t
Xbit_r209_c24 bl[24] br[24] wl[209] vdd gnd cell_6t
Xbit_r210_c24 bl[24] br[24] wl[210] vdd gnd cell_6t
Xbit_r211_c24 bl[24] br[24] wl[211] vdd gnd cell_6t
Xbit_r212_c24 bl[24] br[24] wl[212] vdd gnd cell_6t
Xbit_r213_c24 bl[24] br[24] wl[213] vdd gnd cell_6t
Xbit_r214_c24 bl[24] br[24] wl[214] vdd gnd cell_6t
Xbit_r215_c24 bl[24] br[24] wl[215] vdd gnd cell_6t
Xbit_r216_c24 bl[24] br[24] wl[216] vdd gnd cell_6t
Xbit_r217_c24 bl[24] br[24] wl[217] vdd gnd cell_6t
Xbit_r218_c24 bl[24] br[24] wl[218] vdd gnd cell_6t
Xbit_r219_c24 bl[24] br[24] wl[219] vdd gnd cell_6t
Xbit_r220_c24 bl[24] br[24] wl[220] vdd gnd cell_6t
Xbit_r221_c24 bl[24] br[24] wl[221] vdd gnd cell_6t
Xbit_r222_c24 bl[24] br[24] wl[222] vdd gnd cell_6t
Xbit_r223_c24 bl[24] br[24] wl[223] vdd gnd cell_6t
Xbit_r224_c24 bl[24] br[24] wl[224] vdd gnd cell_6t
Xbit_r225_c24 bl[24] br[24] wl[225] vdd gnd cell_6t
Xbit_r226_c24 bl[24] br[24] wl[226] vdd gnd cell_6t
Xbit_r227_c24 bl[24] br[24] wl[227] vdd gnd cell_6t
Xbit_r228_c24 bl[24] br[24] wl[228] vdd gnd cell_6t
Xbit_r229_c24 bl[24] br[24] wl[229] vdd gnd cell_6t
Xbit_r230_c24 bl[24] br[24] wl[230] vdd gnd cell_6t
Xbit_r231_c24 bl[24] br[24] wl[231] vdd gnd cell_6t
Xbit_r232_c24 bl[24] br[24] wl[232] vdd gnd cell_6t
Xbit_r233_c24 bl[24] br[24] wl[233] vdd gnd cell_6t
Xbit_r234_c24 bl[24] br[24] wl[234] vdd gnd cell_6t
Xbit_r235_c24 bl[24] br[24] wl[235] vdd gnd cell_6t
Xbit_r236_c24 bl[24] br[24] wl[236] vdd gnd cell_6t
Xbit_r237_c24 bl[24] br[24] wl[237] vdd gnd cell_6t
Xbit_r238_c24 bl[24] br[24] wl[238] vdd gnd cell_6t
Xbit_r239_c24 bl[24] br[24] wl[239] vdd gnd cell_6t
Xbit_r240_c24 bl[24] br[24] wl[240] vdd gnd cell_6t
Xbit_r241_c24 bl[24] br[24] wl[241] vdd gnd cell_6t
Xbit_r242_c24 bl[24] br[24] wl[242] vdd gnd cell_6t
Xbit_r243_c24 bl[24] br[24] wl[243] vdd gnd cell_6t
Xbit_r244_c24 bl[24] br[24] wl[244] vdd gnd cell_6t
Xbit_r245_c24 bl[24] br[24] wl[245] vdd gnd cell_6t
Xbit_r246_c24 bl[24] br[24] wl[246] vdd gnd cell_6t
Xbit_r247_c24 bl[24] br[24] wl[247] vdd gnd cell_6t
Xbit_r248_c24 bl[24] br[24] wl[248] vdd gnd cell_6t
Xbit_r249_c24 bl[24] br[24] wl[249] vdd gnd cell_6t
Xbit_r250_c24 bl[24] br[24] wl[250] vdd gnd cell_6t
Xbit_r251_c24 bl[24] br[24] wl[251] vdd gnd cell_6t
Xbit_r252_c24 bl[24] br[24] wl[252] vdd gnd cell_6t
Xbit_r253_c24 bl[24] br[24] wl[253] vdd gnd cell_6t
Xbit_r254_c24 bl[24] br[24] wl[254] vdd gnd cell_6t
Xbit_r255_c24 bl[24] br[24] wl[255] vdd gnd cell_6t
Xbit_r0_c25 bl[25] br[25] wl[0] vdd gnd cell_6t
Xbit_r1_c25 bl[25] br[25] wl[1] vdd gnd cell_6t
Xbit_r2_c25 bl[25] br[25] wl[2] vdd gnd cell_6t
Xbit_r3_c25 bl[25] br[25] wl[3] vdd gnd cell_6t
Xbit_r4_c25 bl[25] br[25] wl[4] vdd gnd cell_6t
Xbit_r5_c25 bl[25] br[25] wl[5] vdd gnd cell_6t
Xbit_r6_c25 bl[25] br[25] wl[6] vdd gnd cell_6t
Xbit_r7_c25 bl[25] br[25] wl[7] vdd gnd cell_6t
Xbit_r8_c25 bl[25] br[25] wl[8] vdd gnd cell_6t
Xbit_r9_c25 bl[25] br[25] wl[9] vdd gnd cell_6t
Xbit_r10_c25 bl[25] br[25] wl[10] vdd gnd cell_6t
Xbit_r11_c25 bl[25] br[25] wl[11] vdd gnd cell_6t
Xbit_r12_c25 bl[25] br[25] wl[12] vdd gnd cell_6t
Xbit_r13_c25 bl[25] br[25] wl[13] vdd gnd cell_6t
Xbit_r14_c25 bl[25] br[25] wl[14] vdd gnd cell_6t
Xbit_r15_c25 bl[25] br[25] wl[15] vdd gnd cell_6t
Xbit_r16_c25 bl[25] br[25] wl[16] vdd gnd cell_6t
Xbit_r17_c25 bl[25] br[25] wl[17] vdd gnd cell_6t
Xbit_r18_c25 bl[25] br[25] wl[18] vdd gnd cell_6t
Xbit_r19_c25 bl[25] br[25] wl[19] vdd gnd cell_6t
Xbit_r20_c25 bl[25] br[25] wl[20] vdd gnd cell_6t
Xbit_r21_c25 bl[25] br[25] wl[21] vdd gnd cell_6t
Xbit_r22_c25 bl[25] br[25] wl[22] vdd gnd cell_6t
Xbit_r23_c25 bl[25] br[25] wl[23] vdd gnd cell_6t
Xbit_r24_c25 bl[25] br[25] wl[24] vdd gnd cell_6t
Xbit_r25_c25 bl[25] br[25] wl[25] vdd gnd cell_6t
Xbit_r26_c25 bl[25] br[25] wl[26] vdd gnd cell_6t
Xbit_r27_c25 bl[25] br[25] wl[27] vdd gnd cell_6t
Xbit_r28_c25 bl[25] br[25] wl[28] vdd gnd cell_6t
Xbit_r29_c25 bl[25] br[25] wl[29] vdd gnd cell_6t
Xbit_r30_c25 bl[25] br[25] wl[30] vdd gnd cell_6t
Xbit_r31_c25 bl[25] br[25] wl[31] vdd gnd cell_6t
Xbit_r32_c25 bl[25] br[25] wl[32] vdd gnd cell_6t
Xbit_r33_c25 bl[25] br[25] wl[33] vdd gnd cell_6t
Xbit_r34_c25 bl[25] br[25] wl[34] vdd gnd cell_6t
Xbit_r35_c25 bl[25] br[25] wl[35] vdd gnd cell_6t
Xbit_r36_c25 bl[25] br[25] wl[36] vdd gnd cell_6t
Xbit_r37_c25 bl[25] br[25] wl[37] vdd gnd cell_6t
Xbit_r38_c25 bl[25] br[25] wl[38] vdd gnd cell_6t
Xbit_r39_c25 bl[25] br[25] wl[39] vdd gnd cell_6t
Xbit_r40_c25 bl[25] br[25] wl[40] vdd gnd cell_6t
Xbit_r41_c25 bl[25] br[25] wl[41] vdd gnd cell_6t
Xbit_r42_c25 bl[25] br[25] wl[42] vdd gnd cell_6t
Xbit_r43_c25 bl[25] br[25] wl[43] vdd gnd cell_6t
Xbit_r44_c25 bl[25] br[25] wl[44] vdd gnd cell_6t
Xbit_r45_c25 bl[25] br[25] wl[45] vdd gnd cell_6t
Xbit_r46_c25 bl[25] br[25] wl[46] vdd gnd cell_6t
Xbit_r47_c25 bl[25] br[25] wl[47] vdd gnd cell_6t
Xbit_r48_c25 bl[25] br[25] wl[48] vdd gnd cell_6t
Xbit_r49_c25 bl[25] br[25] wl[49] vdd gnd cell_6t
Xbit_r50_c25 bl[25] br[25] wl[50] vdd gnd cell_6t
Xbit_r51_c25 bl[25] br[25] wl[51] vdd gnd cell_6t
Xbit_r52_c25 bl[25] br[25] wl[52] vdd gnd cell_6t
Xbit_r53_c25 bl[25] br[25] wl[53] vdd gnd cell_6t
Xbit_r54_c25 bl[25] br[25] wl[54] vdd gnd cell_6t
Xbit_r55_c25 bl[25] br[25] wl[55] vdd gnd cell_6t
Xbit_r56_c25 bl[25] br[25] wl[56] vdd gnd cell_6t
Xbit_r57_c25 bl[25] br[25] wl[57] vdd gnd cell_6t
Xbit_r58_c25 bl[25] br[25] wl[58] vdd gnd cell_6t
Xbit_r59_c25 bl[25] br[25] wl[59] vdd gnd cell_6t
Xbit_r60_c25 bl[25] br[25] wl[60] vdd gnd cell_6t
Xbit_r61_c25 bl[25] br[25] wl[61] vdd gnd cell_6t
Xbit_r62_c25 bl[25] br[25] wl[62] vdd gnd cell_6t
Xbit_r63_c25 bl[25] br[25] wl[63] vdd gnd cell_6t
Xbit_r64_c25 bl[25] br[25] wl[64] vdd gnd cell_6t
Xbit_r65_c25 bl[25] br[25] wl[65] vdd gnd cell_6t
Xbit_r66_c25 bl[25] br[25] wl[66] vdd gnd cell_6t
Xbit_r67_c25 bl[25] br[25] wl[67] vdd gnd cell_6t
Xbit_r68_c25 bl[25] br[25] wl[68] vdd gnd cell_6t
Xbit_r69_c25 bl[25] br[25] wl[69] vdd gnd cell_6t
Xbit_r70_c25 bl[25] br[25] wl[70] vdd gnd cell_6t
Xbit_r71_c25 bl[25] br[25] wl[71] vdd gnd cell_6t
Xbit_r72_c25 bl[25] br[25] wl[72] vdd gnd cell_6t
Xbit_r73_c25 bl[25] br[25] wl[73] vdd gnd cell_6t
Xbit_r74_c25 bl[25] br[25] wl[74] vdd gnd cell_6t
Xbit_r75_c25 bl[25] br[25] wl[75] vdd gnd cell_6t
Xbit_r76_c25 bl[25] br[25] wl[76] vdd gnd cell_6t
Xbit_r77_c25 bl[25] br[25] wl[77] vdd gnd cell_6t
Xbit_r78_c25 bl[25] br[25] wl[78] vdd gnd cell_6t
Xbit_r79_c25 bl[25] br[25] wl[79] vdd gnd cell_6t
Xbit_r80_c25 bl[25] br[25] wl[80] vdd gnd cell_6t
Xbit_r81_c25 bl[25] br[25] wl[81] vdd gnd cell_6t
Xbit_r82_c25 bl[25] br[25] wl[82] vdd gnd cell_6t
Xbit_r83_c25 bl[25] br[25] wl[83] vdd gnd cell_6t
Xbit_r84_c25 bl[25] br[25] wl[84] vdd gnd cell_6t
Xbit_r85_c25 bl[25] br[25] wl[85] vdd gnd cell_6t
Xbit_r86_c25 bl[25] br[25] wl[86] vdd gnd cell_6t
Xbit_r87_c25 bl[25] br[25] wl[87] vdd gnd cell_6t
Xbit_r88_c25 bl[25] br[25] wl[88] vdd gnd cell_6t
Xbit_r89_c25 bl[25] br[25] wl[89] vdd gnd cell_6t
Xbit_r90_c25 bl[25] br[25] wl[90] vdd gnd cell_6t
Xbit_r91_c25 bl[25] br[25] wl[91] vdd gnd cell_6t
Xbit_r92_c25 bl[25] br[25] wl[92] vdd gnd cell_6t
Xbit_r93_c25 bl[25] br[25] wl[93] vdd gnd cell_6t
Xbit_r94_c25 bl[25] br[25] wl[94] vdd gnd cell_6t
Xbit_r95_c25 bl[25] br[25] wl[95] vdd gnd cell_6t
Xbit_r96_c25 bl[25] br[25] wl[96] vdd gnd cell_6t
Xbit_r97_c25 bl[25] br[25] wl[97] vdd gnd cell_6t
Xbit_r98_c25 bl[25] br[25] wl[98] vdd gnd cell_6t
Xbit_r99_c25 bl[25] br[25] wl[99] vdd gnd cell_6t
Xbit_r100_c25 bl[25] br[25] wl[100] vdd gnd cell_6t
Xbit_r101_c25 bl[25] br[25] wl[101] vdd gnd cell_6t
Xbit_r102_c25 bl[25] br[25] wl[102] vdd gnd cell_6t
Xbit_r103_c25 bl[25] br[25] wl[103] vdd gnd cell_6t
Xbit_r104_c25 bl[25] br[25] wl[104] vdd gnd cell_6t
Xbit_r105_c25 bl[25] br[25] wl[105] vdd gnd cell_6t
Xbit_r106_c25 bl[25] br[25] wl[106] vdd gnd cell_6t
Xbit_r107_c25 bl[25] br[25] wl[107] vdd gnd cell_6t
Xbit_r108_c25 bl[25] br[25] wl[108] vdd gnd cell_6t
Xbit_r109_c25 bl[25] br[25] wl[109] vdd gnd cell_6t
Xbit_r110_c25 bl[25] br[25] wl[110] vdd gnd cell_6t
Xbit_r111_c25 bl[25] br[25] wl[111] vdd gnd cell_6t
Xbit_r112_c25 bl[25] br[25] wl[112] vdd gnd cell_6t
Xbit_r113_c25 bl[25] br[25] wl[113] vdd gnd cell_6t
Xbit_r114_c25 bl[25] br[25] wl[114] vdd gnd cell_6t
Xbit_r115_c25 bl[25] br[25] wl[115] vdd gnd cell_6t
Xbit_r116_c25 bl[25] br[25] wl[116] vdd gnd cell_6t
Xbit_r117_c25 bl[25] br[25] wl[117] vdd gnd cell_6t
Xbit_r118_c25 bl[25] br[25] wl[118] vdd gnd cell_6t
Xbit_r119_c25 bl[25] br[25] wl[119] vdd gnd cell_6t
Xbit_r120_c25 bl[25] br[25] wl[120] vdd gnd cell_6t
Xbit_r121_c25 bl[25] br[25] wl[121] vdd gnd cell_6t
Xbit_r122_c25 bl[25] br[25] wl[122] vdd gnd cell_6t
Xbit_r123_c25 bl[25] br[25] wl[123] vdd gnd cell_6t
Xbit_r124_c25 bl[25] br[25] wl[124] vdd gnd cell_6t
Xbit_r125_c25 bl[25] br[25] wl[125] vdd gnd cell_6t
Xbit_r126_c25 bl[25] br[25] wl[126] vdd gnd cell_6t
Xbit_r127_c25 bl[25] br[25] wl[127] vdd gnd cell_6t
Xbit_r128_c25 bl[25] br[25] wl[128] vdd gnd cell_6t
Xbit_r129_c25 bl[25] br[25] wl[129] vdd gnd cell_6t
Xbit_r130_c25 bl[25] br[25] wl[130] vdd gnd cell_6t
Xbit_r131_c25 bl[25] br[25] wl[131] vdd gnd cell_6t
Xbit_r132_c25 bl[25] br[25] wl[132] vdd gnd cell_6t
Xbit_r133_c25 bl[25] br[25] wl[133] vdd gnd cell_6t
Xbit_r134_c25 bl[25] br[25] wl[134] vdd gnd cell_6t
Xbit_r135_c25 bl[25] br[25] wl[135] vdd gnd cell_6t
Xbit_r136_c25 bl[25] br[25] wl[136] vdd gnd cell_6t
Xbit_r137_c25 bl[25] br[25] wl[137] vdd gnd cell_6t
Xbit_r138_c25 bl[25] br[25] wl[138] vdd gnd cell_6t
Xbit_r139_c25 bl[25] br[25] wl[139] vdd gnd cell_6t
Xbit_r140_c25 bl[25] br[25] wl[140] vdd gnd cell_6t
Xbit_r141_c25 bl[25] br[25] wl[141] vdd gnd cell_6t
Xbit_r142_c25 bl[25] br[25] wl[142] vdd gnd cell_6t
Xbit_r143_c25 bl[25] br[25] wl[143] vdd gnd cell_6t
Xbit_r144_c25 bl[25] br[25] wl[144] vdd gnd cell_6t
Xbit_r145_c25 bl[25] br[25] wl[145] vdd gnd cell_6t
Xbit_r146_c25 bl[25] br[25] wl[146] vdd gnd cell_6t
Xbit_r147_c25 bl[25] br[25] wl[147] vdd gnd cell_6t
Xbit_r148_c25 bl[25] br[25] wl[148] vdd gnd cell_6t
Xbit_r149_c25 bl[25] br[25] wl[149] vdd gnd cell_6t
Xbit_r150_c25 bl[25] br[25] wl[150] vdd gnd cell_6t
Xbit_r151_c25 bl[25] br[25] wl[151] vdd gnd cell_6t
Xbit_r152_c25 bl[25] br[25] wl[152] vdd gnd cell_6t
Xbit_r153_c25 bl[25] br[25] wl[153] vdd gnd cell_6t
Xbit_r154_c25 bl[25] br[25] wl[154] vdd gnd cell_6t
Xbit_r155_c25 bl[25] br[25] wl[155] vdd gnd cell_6t
Xbit_r156_c25 bl[25] br[25] wl[156] vdd gnd cell_6t
Xbit_r157_c25 bl[25] br[25] wl[157] vdd gnd cell_6t
Xbit_r158_c25 bl[25] br[25] wl[158] vdd gnd cell_6t
Xbit_r159_c25 bl[25] br[25] wl[159] vdd gnd cell_6t
Xbit_r160_c25 bl[25] br[25] wl[160] vdd gnd cell_6t
Xbit_r161_c25 bl[25] br[25] wl[161] vdd gnd cell_6t
Xbit_r162_c25 bl[25] br[25] wl[162] vdd gnd cell_6t
Xbit_r163_c25 bl[25] br[25] wl[163] vdd gnd cell_6t
Xbit_r164_c25 bl[25] br[25] wl[164] vdd gnd cell_6t
Xbit_r165_c25 bl[25] br[25] wl[165] vdd gnd cell_6t
Xbit_r166_c25 bl[25] br[25] wl[166] vdd gnd cell_6t
Xbit_r167_c25 bl[25] br[25] wl[167] vdd gnd cell_6t
Xbit_r168_c25 bl[25] br[25] wl[168] vdd gnd cell_6t
Xbit_r169_c25 bl[25] br[25] wl[169] vdd gnd cell_6t
Xbit_r170_c25 bl[25] br[25] wl[170] vdd gnd cell_6t
Xbit_r171_c25 bl[25] br[25] wl[171] vdd gnd cell_6t
Xbit_r172_c25 bl[25] br[25] wl[172] vdd gnd cell_6t
Xbit_r173_c25 bl[25] br[25] wl[173] vdd gnd cell_6t
Xbit_r174_c25 bl[25] br[25] wl[174] vdd gnd cell_6t
Xbit_r175_c25 bl[25] br[25] wl[175] vdd gnd cell_6t
Xbit_r176_c25 bl[25] br[25] wl[176] vdd gnd cell_6t
Xbit_r177_c25 bl[25] br[25] wl[177] vdd gnd cell_6t
Xbit_r178_c25 bl[25] br[25] wl[178] vdd gnd cell_6t
Xbit_r179_c25 bl[25] br[25] wl[179] vdd gnd cell_6t
Xbit_r180_c25 bl[25] br[25] wl[180] vdd gnd cell_6t
Xbit_r181_c25 bl[25] br[25] wl[181] vdd gnd cell_6t
Xbit_r182_c25 bl[25] br[25] wl[182] vdd gnd cell_6t
Xbit_r183_c25 bl[25] br[25] wl[183] vdd gnd cell_6t
Xbit_r184_c25 bl[25] br[25] wl[184] vdd gnd cell_6t
Xbit_r185_c25 bl[25] br[25] wl[185] vdd gnd cell_6t
Xbit_r186_c25 bl[25] br[25] wl[186] vdd gnd cell_6t
Xbit_r187_c25 bl[25] br[25] wl[187] vdd gnd cell_6t
Xbit_r188_c25 bl[25] br[25] wl[188] vdd gnd cell_6t
Xbit_r189_c25 bl[25] br[25] wl[189] vdd gnd cell_6t
Xbit_r190_c25 bl[25] br[25] wl[190] vdd gnd cell_6t
Xbit_r191_c25 bl[25] br[25] wl[191] vdd gnd cell_6t
Xbit_r192_c25 bl[25] br[25] wl[192] vdd gnd cell_6t
Xbit_r193_c25 bl[25] br[25] wl[193] vdd gnd cell_6t
Xbit_r194_c25 bl[25] br[25] wl[194] vdd gnd cell_6t
Xbit_r195_c25 bl[25] br[25] wl[195] vdd gnd cell_6t
Xbit_r196_c25 bl[25] br[25] wl[196] vdd gnd cell_6t
Xbit_r197_c25 bl[25] br[25] wl[197] vdd gnd cell_6t
Xbit_r198_c25 bl[25] br[25] wl[198] vdd gnd cell_6t
Xbit_r199_c25 bl[25] br[25] wl[199] vdd gnd cell_6t
Xbit_r200_c25 bl[25] br[25] wl[200] vdd gnd cell_6t
Xbit_r201_c25 bl[25] br[25] wl[201] vdd gnd cell_6t
Xbit_r202_c25 bl[25] br[25] wl[202] vdd gnd cell_6t
Xbit_r203_c25 bl[25] br[25] wl[203] vdd gnd cell_6t
Xbit_r204_c25 bl[25] br[25] wl[204] vdd gnd cell_6t
Xbit_r205_c25 bl[25] br[25] wl[205] vdd gnd cell_6t
Xbit_r206_c25 bl[25] br[25] wl[206] vdd gnd cell_6t
Xbit_r207_c25 bl[25] br[25] wl[207] vdd gnd cell_6t
Xbit_r208_c25 bl[25] br[25] wl[208] vdd gnd cell_6t
Xbit_r209_c25 bl[25] br[25] wl[209] vdd gnd cell_6t
Xbit_r210_c25 bl[25] br[25] wl[210] vdd gnd cell_6t
Xbit_r211_c25 bl[25] br[25] wl[211] vdd gnd cell_6t
Xbit_r212_c25 bl[25] br[25] wl[212] vdd gnd cell_6t
Xbit_r213_c25 bl[25] br[25] wl[213] vdd gnd cell_6t
Xbit_r214_c25 bl[25] br[25] wl[214] vdd gnd cell_6t
Xbit_r215_c25 bl[25] br[25] wl[215] vdd gnd cell_6t
Xbit_r216_c25 bl[25] br[25] wl[216] vdd gnd cell_6t
Xbit_r217_c25 bl[25] br[25] wl[217] vdd gnd cell_6t
Xbit_r218_c25 bl[25] br[25] wl[218] vdd gnd cell_6t
Xbit_r219_c25 bl[25] br[25] wl[219] vdd gnd cell_6t
Xbit_r220_c25 bl[25] br[25] wl[220] vdd gnd cell_6t
Xbit_r221_c25 bl[25] br[25] wl[221] vdd gnd cell_6t
Xbit_r222_c25 bl[25] br[25] wl[222] vdd gnd cell_6t
Xbit_r223_c25 bl[25] br[25] wl[223] vdd gnd cell_6t
Xbit_r224_c25 bl[25] br[25] wl[224] vdd gnd cell_6t
Xbit_r225_c25 bl[25] br[25] wl[225] vdd gnd cell_6t
Xbit_r226_c25 bl[25] br[25] wl[226] vdd gnd cell_6t
Xbit_r227_c25 bl[25] br[25] wl[227] vdd gnd cell_6t
Xbit_r228_c25 bl[25] br[25] wl[228] vdd gnd cell_6t
Xbit_r229_c25 bl[25] br[25] wl[229] vdd gnd cell_6t
Xbit_r230_c25 bl[25] br[25] wl[230] vdd gnd cell_6t
Xbit_r231_c25 bl[25] br[25] wl[231] vdd gnd cell_6t
Xbit_r232_c25 bl[25] br[25] wl[232] vdd gnd cell_6t
Xbit_r233_c25 bl[25] br[25] wl[233] vdd gnd cell_6t
Xbit_r234_c25 bl[25] br[25] wl[234] vdd gnd cell_6t
Xbit_r235_c25 bl[25] br[25] wl[235] vdd gnd cell_6t
Xbit_r236_c25 bl[25] br[25] wl[236] vdd gnd cell_6t
Xbit_r237_c25 bl[25] br[25] wl[237] vdd gnd cell_6t
Xbit_r238_c25 bl[25] br[25] wl[238] vdd gnd cell_6t
Xbit_r239_c25 bl[25] br[25] wl[239] vdd gnd cell_6t
Xbit_r240_c25 bl[25] br[25] wl[240] vdd gnd cell_6t
Xbit_r241_c25 bl[25] br[25] wl[241] vdd gnd cell_6t
Xbit_r242_c25 bl[25] br[25] wl[242] vdd gnd cell_6t
Xbit_r243_c25 bl[25] br[25] wl[243] vdd gnd cell_6t
Xbit_r244_c25 bl[25] br[25] wl[244] vdd gnd cell_6t
Xbit_r245_c25 bl[25] br[25] wl[245] vdd gnd cell_6t
Xbit_r246_c25 bl[25] br[25] wl[246] vdd gnd cell_6t
Xbit_r247_c25 bl[25] br[25] wl[247] vdd gnd cell_6t
Xbit_r248_c25 bl[25] br[25] wl[248] vdd gnd cell_6t
Xbit_r249_c25 bl[25] br[25] wl[249] vdd gnd cell_6t
Xbit_r250_c25 bl[25] br[25] wl[250] vdd gnd cell_6t
Xbit_r251_c25 bl[25] br[25] wl[251] vdd gnd cell_6t
Xbit_r252_c25 bl[25] br[25] wl[252] vdd gnd cell_6t
Xbit_r253_c25 bl[25] br[25] wl[253] vdd gnd cell_6t
Xbit_r254_c25 bl[25] br[25] wl[254] vdd gnd cell_6t
Xbit_r255_c25 bl[25] br[25] wl[255] vdd gnd cell_6t
Xbit_r0_c26 bl[26] br[26] wl[0] vdd gnd cell_6t
Xbit_r1_c26 bl[26] br[26] wl[1] vdd gnd cell_6t
Xbit_r2_c26 bl[26] br[26] wl[2] vdd gnd cell_6t
Xbit_r3_c26 bl[26] br[26] wl[3] vdd gnd cell_6t
Xbit_r4_c26 bl[26] br[26] wl[4] vdd gnd cell_6t
Xbit_r5_c26 bl[26] br[26] wl[5] vdd gnd cell_6t
Xbit_r6_c26 bl[26] br[26] wl[6] vdd gnd cell_6t
Xbit_r7_c26 bl[26] br[26] wl[7] vdd gnd cell_6t
Xbit_r8_c26 bl[26] br[26] wl[8] vdd gnd cell_6t
Xbit_r9_c26 bl[26] br[26] wl[9] vdd gnd cell_6t
Xbit_r10_c26 bl[26] br[26] wl[10] vdd gnd cell_6t
Xbit_r11_c26 bl[26] br[26] wl[11] vdd gnd cell_6t
Xbit_r12_c26 bl[26] br[26] wl[12] vdd gnd cell_6t
Xbit_r13_c26 bl[26] br[26] wl[13] vdd gnd cell_6t
Xbit_r14_c26 bl[26] br[26] wl[14] vdd gnd cell_6t
Xbit_r15_c26 bl[26] br[26] wl[15] vdd gnd cell_6t
Xbit_r16_c26 bl[26] br[26] wl[16] vdd gnd cell_6t
Xbit_r17_c26 bl[26] br[26] wl[17] vdd gnd cell_6t
Xbit_r18_c26 bl[26] br[26] wl[18] vdd gnd cell_6t
Xbit_r19_c26 bl[26] br[26] wl[19] vdd gnd cell_6t
Xbit_r20_c26 bl[26] br[26] wl[20] vdd gnd cell_6t
Xbit_r21_c26 bl[26] br[26] wl[21] vdd gnd cell_6t
Xbit_r22_c26 bl[26] br[26] wl[22] vdd gnd cell_6t
Xbit_r23_c26 bl[26] br[26] wl[23] vdd gnd cell_6t
Xbit_r24_c26 bl[26] br[26] wl[24] vdd gnd cell_6t
Xbit_r25_c26 bl[26] br[26] wl[25] vdd gnd cell_6t
Xbit_r26_c26 bl[26] br[26] wl[26] vdd gnd cell_6t
Xbit_r27_c26 bl[26] br[26] wl[27] vdd gnd cell_6t
Xbit_r28_c26 bl[26] br[26] wl[28] vdd gnd cell_6t
Xbit_r29_c26 bl[26] br[26] wl[29] vdd gnd cell_6t
Xbit_r30_c26 bl[26] br[26] wl[30] vdd gnd cell_6t
Xbit_r31_c26 bl[26] br[26] wl[31] vdd gnd cell_6t
Xbit_r32_c26 bl[26] br[26] wl[32] vdd gnd cell_6t
Xbit_r33_c26 bl[26] br[26] wl[33] vdd gnd cell_6t
Xbit_r34_c26 bl[26] br[26] wl[34] vdd gnd cell_6t
Xbit_r35_c26 bl[26] br[26] wl[35] vdd gnd cell_6t
Xbit_r36_c26 bl[26] br[26] wl[36] vdd gnd cell_6t
Xbit_r37_c26 bl[26] br[26] wl[37] vdd gnd cell_6t
Xbit_r38_c26 bl[26] br[26] wl[38] vdd gnd cell_6t
Xbit_r39_c26 bl[26] br[26] wl[39] vdd gnd cell_6t
Xbit_r40_c26 bl[26] br[26] wl[40] vdd gnd cell_6t
Xbit_r41_c26 bl[26] br[26] wl[41] vdd gnd cell_6t
Xbit_r42_c26 bl[26] br[26] wl[42] vdd gnd cell_6t
Xbit_r43_c26 bl[26] br[26] wl[43] vdd gnd cell_6t
Xbit_r44_c26 bl[26] br[26] wl[44] vdd gnd cell_6t
Xbit_r45_c26 bl[26] br[26] wl[45] vdd gnd cell_6t
Xbit_r46_c26 bl[26] br[26] wl[46] vdd gnd cell_6t
Xbit_r47_c26 bl[26] br[26] wl[47] vdd gnd cell_6t
Xbit_r48_c26 bl[26] br[26] wl[48] vdd gnd cell_6t
Xbit_r49_c26 bl[26] br[26] wl[49] vdd gnd cell_6t
Xbit_r50_c26 bl[26] br[26] wl[50] vdd gnd cell_6t
Xbit_r51_c26 bl[26] br[26] wl[51] vdd gnd cell_6t
Xbit_r52_c26 bl[26] br[26] wl[52] vdd gnd cell_6t
Xbit_r53_c26 bl[26] br[26] wl[53] vdd gnd cell_6t
Xbit_r54_c26 bl[26] br[26] wl[54] vdd gnd cell_6t
Xbit_r55_c26 bl[26] br[26] wl[55] vdd gnd cell_6t
Xbit_r56_c26 bl[26] br[26] wl[56] vdd gnd cell_6t
Xbit_r57_c26 bl[26] br[26] wl[57] vdd gnd cell_6t
Xbit_r58_c26 bl[26] br[26] wl[58] vdd gnd cell_6t
Xbit_r59_c26 bl[26] br[26] wl[59] vdd gnd cell_6t
Xbit_r60_c26 bl[26] br[26] wl[60] vdd gnd cell_6t
Xbit_r61_c26 bl[26] br[26] wl[61] vdd gnd cell_6t
Xbit_r62_c26 bl[26] br[26] wl[62] vdd gnd cell_6t
Xbit_r63_c26 bl[26] br[26] wl[63] vdd gnd cell_6t
Xbit_r64_c26 bl[26] br[26] wl[64] vdd gnd cell_6t
Xbit_r65_c26 bl[26] br[26] wl[65] vdd gnd cell_6t
Xbit_r66_c26 bl[26] br[26] wl[66] vdd gnd cell_6t
Xbit_r67_c26 bl[26] br[26] wl[67] vdd gnd cell_6t
Xbit_r68_c26 bl[26] br[26] wl[68] vdd gnd cell_6t
Xbit_r69_c26 bl[26] br[26] wl[69] vdd gnd cell_6t
Xbit_r70_c26 bl[26] br[26] wl[70] vdd gnd cell_6t
Xbit_r71_c26 bl[26] br[26] wl[71] vdd gnd cell_6t
Xbit_r72_c26 bl[26] br[26] wl[72] vdd gnd cell_6t
Xbit_r73_c26 bl[26] br[26] wl[73] vdd gnd cell_6t
Xbit_r74_c26 bl[26] br[26] wl[74] vdd gnd cell_6t
Xbit_r75_c26 bl[26] br[26] wl[75] vdd gnd cell_6t
Xbit_r76_c26 bl[26] br[26] wl[76] vdd gnd cell_6t
Xbit_r77_c26 bl[26] br[26] wl[77] vdd gnd cell_6t
Xbit_r78_c26 bl[26] br[26] wl[78] vdd gnd cell_6t
Xbit_r79_c26 bl[26] br[26] wl[79] vdd gnd cell_6t
Xbit_r80_c26 bl[26] br[26] wl[80] vdd gnd cell_6t
Xbit_r81_c26 bl[26] br[26] wl[81] vdd gnd cell_6t
Xbit_r82_c26 bl[26] br[26] wl[82] vdd gnd cell_6t
Xbit_r83_c26 bl[26] br[26] wl[83] vdd gnd cell_6t
Xbit_r84_c26 bl[26] br[26] wl[84] vdd gnd cell_6t
Xbit_r85_c26 bl[26] br[26] wl[85] vdd gnd cell_6t
Xbit_r86_c26 bl[26] br[26] wl[86] vdd gnd cell_6t
Xbit_r87_c26 bl[26] br[26] wl[87] vdd gnd cell_6t
Xbit_r88_c26 bl[26] br[26] wl[88] vdd gnd cell_6t
Xbit_r89_c26 bl[26] br[26] wl[89] vdd gnd cell_6t
Xbit_r90_c26 bl[26] br[26] wl[90] vdd gnd cell_6t
Xbit_r91_c26 bl[26] br[26] wl[91] vdd gnd cell_6t
Xbit_r92_c26 bl[26] br[26] wl[92] vdd gnd cell_6t
Xbit_r93_c26 bl[26] br[26] wl[93] vdd gnd cell_6t
Xbit_r94_c26 bl[26] br[26] wl[94] vdd gnd cell_6t
Xbit_r95_c26 bl[26] br[26] wl[95] vdd gnd cell_6t
Xbit_r96_c26 bl[26] br[26] wl[96] vdd gnd cell_6t
Xbit_r97_c26 bl[26] br[26] wl[97] vdd gnd cell_6t
Xbit_r98_c26 bl[26] br[26] wl[98] vdd gnd cell_6t
Xbit_r99_c26 bl[26] br[26] wl[99] vdd gnd cell_6t
Xbit_r100_c26 bl[26] br[26] wl[100] vdd gnd cell_6t
Xbit_r101_c26 bl[26] br[26] wl[101] vdd gnd cell_6t
Xbit_r102_c26 bl[26] br[26] wl[102] vdd gnd cell_6t
Xbit_r103_c26 bl[26] br[26] wl[103] vdd gnd cell_6t
Xbit_r104_c26 bl[26] br[26] wl[104] vdd gnd cell_6t
Xbit_r105_c26 bl[26] br[26] wl[105] vdd gnd cell_6t
Xbit_r106_c26 bl[26] br[26] wl[106] vdd gnd cell_6t
Xbit_r107_c26 bl[26] br[26] wl[107] vdd gnd cell_6t
Xbit_r108_c26 bl[26] br[26] wl[108] vdd gnd cell_6t
Xbit_r109_c26 bl[26] br[26] wl[109] vdd gnd cell_6t
Xbit_r110_c26 bl[26] br[26] wl[110] vdd gnd cell_6t
Xbit_r111_c26 bl[26] br[26] wl[111] vdd gnd cell_6t
Xbit_r112_c26 bl[26] br[26] wl[112] vdd gnd cell_6t
Xbit_r113_c26 bl[26] br[26] wl[113] vdd gnd cell_6t
Xbit_r114_c26 bl[26] br[26] wl[114] vdd gnd cell_6t
Xbit_r115_c26 bl[26] br[26] wl[115] vdd gnd cell_6t
Xbit_r116_c26 bl[26] br[26] wl[116] vdd gnd cell_6t
Xbit_r117_c26 bl[26] br[26] wl[117] vdd gnd cell_6t
Xbit_r118_c26 bl[26] br[26] wl[118] vdd gnd cell_6t
Xbit_r119_c26 bl[26] br[26] wl[119] vdd gnd cell_6t
Xbit_r120_c26 bl[26] br[26] wl[120] vdd gnd cell_6t
Xbit_r121_c26 bl[26] br[26] wl[121] vdd gnd cell_6t
Xbit_r122_c26 bl[26] br[26] wl[122] vdd gnd cell_6t
Xbit_r123_c26 bl[26] br[26] wl[123] vdd gnd cell_6t
Xbit_r124_c26 bl[26] br[26] wl[124] vdd gnd cell_6t
Xbit_r125_c26 bl[26] br[26] wl[125] vdd gnd cell_6t
Xbit_r126_c26 bl[26] br[26] wl[126] vdd gnd cell_6t
Xbit_r127_c26 bl[26] br[26] wl[127] vdd gnd cell_6t
Xbit_r128_c26 bl[26] br[26] wl[128] vdd gnd cell_6t
Xbit_r129_c26 bl[26] br[26] wl[129] vdd gnd cell_6t
Xbit_r130_c26 bl[26] br[26] wl[130] vdd gnd cell_6t
Xbit_r131_c26 bl[26] br[26] wl[131] vdd gnd cell_6t
Xbit_r132_c26 bl[26] br[26] wl[132] vdd gnd cell_6t
Xbit_r133_c26 bl[26] br[26] wl[133] vdd gnd cell_6t
Xbit_r134_c26 bl[26] br[26] wl[134] vdd gnd cell_6t
Xbit_r135_c26 bl[26] br[26] wl[135] vdd gnd cell_6t
Xbit_r136_c26 bl[26] br[26] wl[136] vdd gnd cell_6t
Xbit_r137_c26 bl[26] br[26] wl[137] vdd gnd cell_6t
Xbit_r138_c26 bl[26] br[26] wl[138] vdd gnd cell_6t
Xbit_r139_c26 bl[26] br[26] wl[139] vdd gnd cell_6t
Xbit_r140_c26 bl[26] br[26] wl[140] vdd gnd cell_6t
Xbit_r141_c26 bl[26] br[26] wl[141] vdd gnd cell_6t
Xbit_r142_c26 bl[26] br[26] wl[142] vdd gnd cell_6t
Xbit_r143_c26 bl[26] br[26] wl[143] vdd gnd cell_6t
Xbit_r144_c26 bl[26] br[26] wl[144] vdd gnd cell_6t
Xbit_r145_c26 bl[26] br[26] wl[145] vdd gnd cell_6t
Xbit_r146_c26 bl[26] br[26] wl[146] vdd gnd cell_6t
Xbit_r147_c26 bl[26] br[26] wl[147] vdd gnd cell_6t
Xbit_r148_c26 bl[26] br[26] wl[148] vdd gnd cell_6t
Xbit_r149_c26 bl[26] br[26] wl[149] vdd gnd cell_6t
Xbit_r150_c26 bl[26] br[26] wl[150] vdd gnd cell_6t
Xbit_r151_c26 bl[26] br[26] wl[151] vdd gnd cell_6t
Xbit_r152_c26 bl[26] br[26] wl[152] vdd gnd cell_6t
Xbit_r153_c26 bl[26] br[26] wl[153] vdd gnd cell_6t
Xbit_r154_c26 bl[26] br[26] wl[154] vdd gnd cell_6t
Xbit_r155_c26 bl[26] br[26] wl[155] vdd gnd cell_6t
Xbit_r156_c26 bl[26] br[26] wl[156] vdd gnd cell_6t
Xbit_r157_c26 bl[26] br[26] wl[157] vdd gnd cell_6t
Xbit_r158_c26 bl[26] br[26] wl[158] vdd gnd cell_6t
Xbit_r159_c26 bl[26] br[26] wl[159] vdd gnd cell_6t
Xbit_r160_c26 bl[26] br[26] wl[160] vdd gnd cell_6t
Xbit_r161_c26 bl[26] br[26] wl[161] vdd gnd cell_6t
Xbit_r162_c26 bl[26] br[26] wl[162] vdd gnd cell_6t
Xbit_r163_c26 bl[26] br[26] wl[163] vdd gnd cell_6t
Xbit_r164_c26 bl[26] br[26] wl[164] vdd gnd cell_6t
Xbit_r165_c26 bl[26] br[26] wl[165] vdd gnd cell_6t
Xbit_r166_c26 bl[26] br[26] wl[166] vdd gnd cell_6t
Xbit_r167_c26 bl[26] br[26] wl[167] vdd gnd cell_6t
Xbit_r168_c26 bl[26] br[26] wl[168] vdd gnd cell_6t
Xbit_r169_c26 bl[26] br[26] wl[169] vdd gnd cell_6t
Xbit_r170_c26 bl[26] br[26] wl[170] vdd gnd cell_6t
Xbit_r171_c26 bl[26] br[26] wl[171] vdd gnd cell_6t
Xbit_r172_c26 bl[26] br[26] wl[172] vdd gnd cell_6t
Xbit_r173_c26 bl[26] br[26] wl[173] vdd gnd cell_6t
Xbit_r174_c26 bl[26] br[26] wl[174] vdd gnd cell_6t
Xbit_r175_c26 bl[26] br[26] wl[175] vdd gnd cell_6t
Xbit_r176_c26 bl[26] br[26] wl[176] vdd gnd cell_6t
Xbit_r177_c26 bl[26] br[26] wl[177] vdd gnd cell_6t
Xbit_r178_c26 bl[26] br[26] wl[178] vdd gnd cell_6t
Xbit_r179_c26 bl[26] br[26] wl[179] vdd gnd cell_6t
Xbit_r180_c26 bl[26] br[26] wl[180] vdd gnd cell_6t
Xbit_r181_c26 bl[26] br[26] wl[181] vdd gnd cell_6t
Xbit_r182_c26 bl[26] br[26] wl[182] vdd gnd cell_6t
Xbit_r183_c26 bl[26] br[26] wl[183] vdd gnd cell_6t
Xbit_r184_c26 bl[26] br[26] wl[184] vdd gnd cell_6t
Xbit_r185_c26 bl[26] br[26] wl[185] vdd gnd cell_6t
Xbit_r186_c26 bl[26] br[26] wl[186] vdd gnd cell_6t
Xbit_r187_c26 bl[26] br[26] wl[187] vdd gnd cell_6t
Xbit_r188_c26 bl[26] br[26] wl[188] vdd gnd cell_6t
Xbit_r189_c26 bl[26] br[26] wl[189] vdd gnd cell_6t
Xbit_r190_c26 bl[26] br[26] wl[190] vdd gnd cell_6t
Xbit_r191_c26 bl[26] br[26] wl[191] vdd gnd cell_6t
Xbit_r192_c26 bl[26] br[26] wl[192] vdd gnd cell_6t
Xbit_r193_c26 bl[26] br[26] wl[193] vdd gnd cell_6t
Xbit_r194_c26 bl[26] br[26] wl[194] vdd gnd cell_6t
Xbit_r195_c26 bl[26] br[26] wl[195] vdd gnd cell_6t
Xbit_r196_c26 bl[26] br[26] wl[196] vdd gnd cell_6t
Xbit_r197_c26 bl[26] br[26] wl[197] vdd gnd cell_6t
Xbit_r198_c26 bl[26] br[26] wl[198] vdd gnd cell_6t
Xbit_r199_c26 bl[26] br[26] wl[199] vdd gnd cell_6t
Xbit_r200_c26 bl[26] br[26] wl[200] vdd gnd cell_6t
Xbit_r201_c26 bl[26] br[26] wl[201] vdd gnd cell_6t
Xbit_r202_c26 bl[26] br[26] wl[202] vdd gnd cell_6t
Xbit_r203_c26 bl[26] br[26] wl[203] vdd gnd cell_6t
Xbit_r204_c26 bl[26] br[26] wl[204] vdd gnd cell_6t
Xbit_r205_c26 bl[26] br[26] wl[205] vdd gnd cell_6t
Xbit_r206_c26 bl[26] br[26] wl[206] vdd gnd cell_6t
Xbit_r207_c26 bl[26] br[26] wl[207] vdd gnd cell_6t
Xbit_r208_c26 bl[26] br[26] wl[208] vdd gnd cell_6t
Xbit_r209_c26 bl[26] br[26] wl[209] vdd gnd cell_6t
Xbit_r210_c26 bl[26] br[26] wl[210] vdd gnd cell_6t
Xbit_r211_c26 bl[26] br[26] wl[211] vdd gnd cell_6t
Xbit_r212_c26 bl[26] br[26] wl[212] vdd gnd cell_6t
Xbit_r213_c26 bl[26] br[26] wl[213] vdd gnd cell_6t
Xbit_r214_c26 bl[26] br[26] wl[214] vdd gnd cell_6t
Xbit_r215_c26 bl[26] br[26] wl[215] vdd gnd cell_6t
Xbit_r216_c26 bl[26] br[26] wl[216] vdd gnd cell_6t
Xbit_r217_c26 bl[26] br[26] wl[217] vdd gnd cell_6t
Xbit_r218_c26 bl[26] br[26] wl[218] vdd gnd cell_6t
Xbit_r219_c26 bl[26] br[26] wl[219] vdd gnd cell_6t
Xbit_r220_c26 bl[26] br[26] wl[220] vdd gnd cell_6t
Xbit_r221_c26 bl[26] br[26] wl[221] vdd gnd cell_6t
Xbit_r222_c26 bl[26] br[26] wl[222] vdd gnd cell_6t
Xbit_r223_c26 bl[26] br[26] wl[223] vdd gnd cell_6t
Xbit_r224_c26 bl[26] br[26] wl[224] vdd gnd cell_6t
Xbit_r225_c26 bl[26] br[26] wl[225] vdd gnd cell_6t
Xbit_r226_c26 bl[26] br[26] wl[226] vdd gnd cell_6t
Xbit_r227_c26 bl[26] br[26] wl[227] vdd gnd cell_6t
Xbit_r228_c26 bl[26] br[26] wl[228] vdd gnd cell_6t
Xbit_r229_c26 bl[26] br[26] wl[229] vdd gnd cell_6t
Xbit_r230_c26 bl[26] br[26] wl[230] vdd gnd cell_6t
Xbit_r231_c26 bl[26] br[26] wl[231] vdd gnd cell_6t
Xbit_r232_c26 bl[26] br[26] wl[232] vdd gnd cell_6t
Xbit_r233_c26 bl[26] br[26] wl[233] vdd gnd cell_6t
Xbit_r234_c26 bl[26] br[26] wl[234] vdd gnd cell_6t
Xbit_r235_c26 bl[26] br[26] wl[235] vdd gnd cell_6t
Xbit_r236_c26 bl[26] br[26] wl[236] vdd gnd cell_6t
Xbit_r237_c26 bl[26] br[26] wl[237] vdd gnd cell_6t
Xbit_r238_c26 bl[26] br[26] wl[238] vdd gnd cell_6t
Xbit_r239_c26 bl[26] br[26] wl[239] vdd gnd cell_6t
Xbit_r240_c26 bl[26] br[26] wl[240] vdd gnd cell_6t
Xbit_r241_c26 bl[26] br[26] wl[241] vdd gnd cell_6t
Xbit_r242_c26 bl[26] br[26] wl[242] vdd gnd cell_6t
Xbit_r243_c26 bl[26] br[26] wl[243] vdd gnd cell_6t
Xbit_r244_c26 bl[26] br[26] wl[244] vdd gnd cell_6t
Xbit_r245_c26 bl[26] br[26] wl[245] vdd gnd cell_6t
Xbit_r246_c26 bl[26] br[26] wl[246] vdd gnd cell_6t
Xbit_r247_c26 bl[26] br[26] wl[247] vdd gnd cell_6t
Xbit_r248_c26 bl[26] br[26] wl[248] vdd gnd cell_6t
Xbit_r249_c26 bl[26] br[26] wl[249] vdd gnd cell_6t
Xbit_r250_c26 bl[26] br[26] wl[250] vdd gnd cell_6t
Xbit_r251_c26 bl[26] br[26] wl[251] vdd gnd cell_6t
Xbit_r252_c26 bl[26] br[26] wl[252] vdd gnd cell_6t
Xbit_r253_c26 bl[26] br[26] wl[253] vdd gnd cell_6t
Xbit_r254_c26 bl[26] br[26] wl[254] vdd gnd cell_6t
Xbit_r255_c26 bl[26] br[26] wl[255] vdd gnd cell_6t
Xbit_r0_c27 bl[27] br[27] wl[0] vdd gnd cell_6t
Xbit_r1_c27 bl[27] br[27] wl[1] vdd gnd cell_6t
Xbit_r2_c27 bl[27] br[27] wl[2] vdd gnd cell_6t
Xbit_r3_c27 bl[27] br[27] wl[3] vdd gnd cell_6t
Xbit_r4_c27 bl[27] br[27] wl[4] vdd gnd cell_6t
Xbit_r5_c27 bl[27] br[27] wl[5] vdd gnd cell_6t
Xbit_r6_c27 bl[27] br[27] wl[6] vdd gnd cell_6t
Xbit_r7_c27 bl[27] br[27] wl[7] vdd gnd cell_6t
Xbit_r8_c27 bl[27] br[27] wl[8] vdd gnd cell_6t
Xbit_r9_c27 bl[27] br[27] wl[9] vdd gnd cell_6t
Xbit_r10_c27 bl[27] br[27] wl[10] vdd gnd cell_6t
Xbit_r11_c27 bl[27] br[27] wl[11] vdd gnd cell_6t
Xbit_r12_c27 bl[27] br[27] wl[12] vdd gnd cell_6t
Xbit_r13_c27 bl[27] br[27] wl[13] vdd gnd cell_6t
Xbit_r14_c27 bl[27] br[27] wl[14] vdd gnd cell_6t
Xbit_r15_c27 bl[27] br[27] wl[15] vdd gnd cell_6t
Xbit_r16_c27 bl[27] br[27] wl[16] vdd gnd cell_6t
Xbit_r17_c27 bl[27] br[27] wl[17] vdd gnd cell_6t
Xbit_r18_c27 bl[27] br[27] wl[18] vdd gnd cell_6t
Xbit_r19_c27 bl[27] br[27] wl[19] vdd gnd cell_6t
Xbit_r20_c27 bl[27] br[27] wl[20] vdd gnd cell_6t
Xbit_r21_c27 bl[27] br[27] wl[21] vdd gnd cell_6t
Xbit_r22_c27 bl[27] br[27] wl[22] vdd gnd cell_6t
Xbit_r23_c27 bl[27] br[27] wl[23] vdd gnd cell_6t
Xbit_r24_c27 bl[27] br[27] wl[24] vdd gnd cell_6t
Xbit_r25_c27 bl[27] br[27] wl[25] vdd gnd cell_6t
Xbit_r26_c27 bl[27] br[27] wl[26] vdd gnd cell_6t
Xbit_r27_c27 bl[27] br[27] wl[27] vdd gnd cell_6t
Xbit_r28_c27 bl[27] br[27] wl[28] vdd gnd cell_6t
Xbit_r29_c27 bl[27] br[27] wl[29] vdd gnd cell_6t
Xbit_r30_c27 bl[27] br[27] wl[30] vdd gnd cell_6t
Xbit_r31_c27 bl[27] br[27] wl[31] vdd gnd cell_6t
Xbit_r32_c27 bl[27] br[27] wl[32] vdd gnd cell_6t
Xbit_r33_c27 bl[27] br[27] wl[33] vdd gnd cell_6t
Xbit_r34_c27 bl[27] br[27] wl[34] vdd gnd cell_6t
Xbit_r35_c27 bl[27] br[27] wl[35] vdd gnd cell_6t
Xbit_r36_c27 bl[27] br[27] wl[36] vdd gnd cell_6t
Xbit_r37_c27 bl[27] br[27] wl[37] vdd gnd cell_6t
Xbit_r38_c27 bl[27] br[27] wl[38] vdd gnd cell_6t
Xbit_r39_c27 bl[27] br[27] wl[39] vdd gnd cell_6t
Xbit_r40_c27 bl[27] br[27] wl[40] vdd gnd cell_6t
Xbit_r41_c27 bl[27] br[27] wl[41] vdd gnd cell_6t
Xbit_r42_c27 bl[27] br[27] wl[42] vdd gnd cell_6t
Xbit_r43_c27 bl[27] br[27] wl[43] vdd gnd cell_6t
Xbit_r44_c27 bl[27] br[27] wl[44] vdd gnd cell_6t
Xbit_r45_c27 bl[27] br[27] wl[45] vdd gnd cell_6t
Xbit_r46_c27 bl[27] br[27] wl[46] vdd gnd cell_6t
Xbit_r47_c27 bl[27] br[27] wl[47] vdd gnd cell_6t
Xbit_r48_c27 bl[27] br[27] wl[48] vdd gnd cell_6t
Xbit_r49_c27 bl[27] br[27] wl[49] vdd gnd cell_6t
Xbit_r50_c27 bl[27] br[27] wl[50] vdd gnd cell_6t
Xbit_r51_c27 bl[27] br[27] wl[51] vdd gnd cell_6t
Xbit_r52_c27 bl[27] br[27] wl[52] vdd gnd cell_6t
Xbit_r53_c27 bl[27] br[27] wl[53] vdd gnd cell_6t
Xbit_r54_c27 bl[27] br[27] wl[54] vdd gnd cell_6t
Xbit_r55_c27 bl[27] br[27] wl[55] vdd gnd cell_6t
Xbit_r56_c27 bl[27] br[27] wl[56] vdd gnd cell_6t
Xbit_r57_c27 bl[27] br[27] wl[57] vdd gnd cell_6t
Xbit_r58_c27 bl[27] br[27] wl[58] vdd gnd cell_6t
Xbit_r59_c27 bl[27] br[27] wl[59] vdd gnd cell_6t
Xbit_r60_c27 bl[27] br[27] wl[60] vdd gnd cell_6t
Xbit_r61_c27 bl[27] br[27] wl[61] vdd gnd cell_6t
Xbit_r62_c27 bl[27] br[27] wl[62] vdd gnd cell_6t
Xbit_r63_c27 bl[27] br[27] wl[63] vdd gnd cell_6t
Xbit_r64_c27 bl[27] br[27] wl[64] vdd gnd cell_6t
Xbit_r65_c27 bl[27] br[27] wl[65] vdd gnd cell_6t
Xbit_r66_c27 bl[27] br[27] wl[66] vdd gnd cell_6t
Xbit_r67_c27 bl[27] br[27] wl[67] vdd gnd cell_6t
Xbit_r68_c27 bl[27] br[27] wl[68] vdd gnd cell_6t
Xbit_r69_c27 bl[27] br[27] wl[69] vdd gnd cell_6t
Xbit_r70_c27 bl[27] br[27] wl[70] vdd gnd cell_6t
Xbit_r71_c27 bl[27] br[27] wl[71] vdd gnd cell_6t
Xbit_r72_c27 bl[27] br[27] wl[72] vdd gnd cell_6t
Xbit_r73_c27 bl[27] br[27] wl[73] vdd gnd cell_6t
Xbit_r74_c27 bl[27] br[27] wl[74] vdd gnd cell_6t
Xbit_r75_c27 bl[27] br[27] wl[75] vdd gnd cell_6t
Xbit_r76_c27 bl[27] br[27] wl[76] vdd gnd cell_6t
Xbit_r77_c27 bl[27] br[27] wl[77] vdd gnd cell_6t
Xbit_r78_c27 bl[27] br[27] wl[78] vdd gnd cell_6t
Xbit_r79_c27 bl[27] br[27] wl[79] vdd gnd cell_6t
Xbit_r80_c27 bl[27] br[27] wl[80] vdd gnd cell_6t
Xbit_r81_c27 bl[27] br[27] wl[81] vdd gnd cell_6t
Xbit_r82_c27 bl[27] br[27] wl[82] vdd gnd cell_6t
Xbit_r83_c27 bl[27] br[27] wl[83] vdd gnd cell_6t
Xbit_r84_c27 bl[27] br[27] wl[84] vdd gnd cell_6t
Xbit_r85_c27 bl[27] br[27] wl[85] vdd gnd cell_6t
Xbit_r86_c27 bl[27] br[27] wl[86] vdd gnd cell_6t
Xbit_r87_c27 bl[27] br[27] wl[87] vdd gnd cell_6t
Xbit_r88_c27 bl[27] br[27] wl[88] vdd gnd cell_6t
Xbit_r89_c27 bl[27] br[27] wl[89] vdd gnd cell_6t
Xbit_r90_c27 bl[27] br[27] wl[90] vdd gnd cell_6t
Xbit_r91_c27 bl[27] br[27] wl[91] vdd gnd cell_6t
Xbit_r92_c27 bl[27] br[27] wl[92] vdd gnd cell_6t
Xbit_r93_c27 bl[27] br[27] wl[93] vdd gnd cell_6t
Xbit_r94_c27 bl[27] br[27] wl[94] vdd gnd cell_6t
Xbit_r95_c27 bl[27] br[27] wl[95] vdd gnd cell_6t
Xbit_r96_c27 bl[27] br[27] wl[96] vdd gnd cell_6t
Xbit_r97_c27 bl[27] br[27] wl[97] vdd gnd cell_6t
Xbit_r98_c27 bl[27] br[27] wl[98] vdd gnd cell_6t
Xbit_r99_c27 bl[27] br[27] wl[99] vdd gnd cell_6t
Xbit_r100_c27 bl[27] br[27] wl[100] vdd gnd cell_6t
Xbit_r101_c27 bl[27] br[27] wl[101] vdd gnd cell_6t
Xbit_r102_c27 bl[27] br[27] wl[102] vdd gnd cell_6t
Xbit_r103_c27 bl[27] br[27] wl[103] vdd gnd cell_6t
Xbit_r104_c27 bl[27] br[27] wl[104] vdd gnd cell_6t
Xbit_r105_c27 bl[27] br[27] wl[105] vdd gnd cell_6t
Xbit_r106_c27 bl[27] br[27] wl[106] vdd gnd cell_6t
Xbit_r107_c27 bl[27] br[27] wl[107] vdd gnd cell_6t
Xbit_r108_c27 bl[27] br[27] wl[108] vdd gnd cell_6t
Xbit_r109_c27 bl[27] br[27] wl[109] vdd gnd cell_6t
Xbit_r110_c27 bl[27] br[27] wl[110] vdd gnd cell_6t
Xbit_r111_c27 bl[27] br[27] wl[111] vdd gnd cell_6t
Xbit_r112_c27 bl[27] br[27] wl[112] vdd gnd cell_6t
Xbit_r113_c27 bl[27] br[27] wl[113] vdd gnd cell_6t
Xbit_r114_c27 bl[27] br[27] wl[114] vdd gnd cell_6t
Xbit_r115_c27 bl[27] br[27] wl[115] vdd gnd cell_6t
Xbit_r116_c27 bl[27] br[27] wl[116] vdd gnd cell_6t
Xbit_r117_c27 bl[27] br[27] wl[117] vdd gnd cell_6t
Xbit_r118_c27 bl[27] br[27] wl[118] vdd gnd cell_6t
Xbit_r119_c27 bl[27] br[27] wl[119] vdd gnd cell_6t
Xbit_r120_c27 bl[27] br[27] wl[120] vdd gnd cell_6t
Xbit_r121_c27 bl[27] br[27] wl[121] vdd gnd cell_6t
Xbit_r122_c27 bl[27] br[27] wl[122] vdd gnd cell_6t
Xbit_r123_c27 bl[27] br[27] wl[123] vdd gnd cell_6t
Xbit_r124_c27 bl[27] br[27] wl[124] vdd gnd cell_6t
Xbit_r125_c27 bl[27] br[27] wl[125] vdd gnd cell_6t
Xbit_r126_c27 bl[27] br[27] wl[126] vdd gnd cell_6t
Xbit_r127_c27 bl[27] br[27] wl[127] vdd gnd cell_6t
Xbit_r128_c27 bl[27] br[27] wl[128] vdd gnd cell_6t
Xbit_r129_c27 bl[27] br[27] wl[129] vdd gnd cell_6t
Xbit_r130_c27 bl[27] br[27] wl[130] vdd gnd cell_6t
Xbit_r131_c27 bl[27] br[27] wl[131] vdd gnd cell_6t
Xbit_r132_c27 bl[27] br[27] wl[132] vdd gnd cell_6t
Xbit_r133_c27 bl[27] br[27] wl[133] vdd gnd cell_6t
Xbit_r134_c27 bl[27] br[27] wl[134] vdd gnd cell_6t
Xbit_r135_c27 bl[27] br[27] wl[135] vdd gnd cell_6t
Xbit_r136_c27 bl[27] br[27] wl[136] vdd gnd cell_6t
Xbit_r137_c27 bl[27] br[27] wl[137] vdd gnd cell_6t
Xbit_r138_c27 bl[27] br[27] wl[138] vdd gnd cell_6t
Xbit_r139_c27 bl[27] br[27] wl[139] vdd gnd cell_6t
Xbit_r140_c27 bl[27] br[27] wl[140] vdd gnd cell_6t
Xbit_r141_c27 bl[27] br[27] wl[141] vdd gnd cell_6t
Xbit_r142_c27 bl[27] br[27] wl[142] vdd gnd cell_6t
Xbit_r143_c27 bl[27] br[27] wl[143] vdd gnd cell_6t
Xbit_r144_c27 bl[27] br[27] wl[144] vdd gnd cell_6t
Xbit_r145_c27 bl[27] br[27] wl[145] vdd gnd cell_6t
Xbit_r146_c27 bl[27] br[27] wl[146] vdd gnd cell_6t
Xbit_r147_c27 bl[27] br[27] wl[147] vdd gnd cell_6t
Xbit_r148_c27 bl[27] br[27] wl[148] vdd gnd cell_6t
Xbit_r149_c27 bl[27] br[27] wl[149] vdd gnd cell_6t
Xbit_r150_c27 bl[27] br[27] wl[150] vdd gnd cell_6t
Xbit_r151_c27 bl[27] br[27] wl[151] vdd gnd cell_6t
Xbit_r152_c27 bl[27] br[27] wl[152] vdd gnd cell_6t
Xbit_r153_c27 bl[27] br[27] wl[153] vdd gnd cell_6t
Xbit_r154_c27 bl[27] br[27] wl[154] vdd gnd cell_6t
Xbit_r155_c27 bl[27] br[27] wl[155] vdd gnd cell_6t
Xbit_r156_c27 bl[27] br[27] wl[156] vdd gnd cell_6t
Xbit_r157_c27 bl[27] br[27] wl[157] vdd gnd cell_6t
Xbit_r158_c27 bl[27] br[27] wl[158] vdd gnd cell_6t
Xbit_r159_c27 bl[27] br[27] wl[159] vdd gnd cell_6t
Xbit_r160_c27 bl[27] br[27] wl[160] vdd gnd cell_6t
Xbit_r161_c27 bl[27] br[27] wl[161] vdd gnd cell_6t
Xbit_r162_c27 bl[27] br[27] wl[162] vdd gnd cell_6t
Xbit_r163_c27 bl[27] br[27] wl[163] vdd gnd cell_6t
Xbit_r164_c27 bl[27] br[27] wl[164] vdd gnd cell_6t
Xbit_r165_c27 bl[27] br[27] wl[165] vdd gnd cell_6t
Xbit_r166_c27 bl[27] br[27] wl[166] vdd gnd cell_6t
Xbit_r167_c27 bl[27] br[27] wl[167] vdd gnd cell_6t
Xbit_r168_c27 bl[27] br[27] wl[168] vdd gnd cell_6t
Xbit_r169_c27 bl[27] br[27] wl[169] vdd gnd cell_6t
Xbit_r170_c27 bl[27] br[27] wl[170] vdd gnd cell_6t
Xbit_r171_c27 bl[27] br[27] wl[171] vdd gnd cell_6t
Xbit_r172_c27 bl[27] br[27] wl[172] vdd gnd cell_6t
Xbit_r173_c27 bl[27] br[27] wl[173] vdd gnd cell_6t
Xbit_r174_c27 bl[27] br[27] wl[174] vdd gnd cell_6t
Xbit_r175_c27 bl[27] br[27] wl[175] vdd gnd cell_6t
Xbit_r176_c27 bl[27] br[27] wl[176] vdd gnd cell_6t
Xbit_r177_c27 bl[27] br[27] wl[177] vdd gnd cell_6t
Xbit_r178_c27 bl[27] br[27] wl[178] vdd gnd cell_6t
Xbit_r179_c27 bl[27] br[27] wl[179] vdd gnd cell_6t
Xbit_r180_c27 bl[27] br[27] wl[180] vdd gnd cell_6t
Xbit_r181_c27 bl[27] br[27] wl[181] vdd gnd cell_6t
Xbit_r182_c27 bl[27] br[27] wl[182] vdd gnd cell_6t
Xbit_r183_c27 bl[27] br[27] wl[183] vdd gnd cell_6t
Xbit_r184_c27 bl[27] br[27] wl[184] vdd gnd cell_6t
Xbit_r185_c27 bl[27] br[27] wl[185] vdd gnd cell_6t
Xbit_r186_c27 bl[27] br[27] wl[186] vdd gnd cell_6t
Xbit_r187_c27 bl[27] br[27] wl[187] vdd gnd cell_6t
Xbit_r188_c27 bl[27] br[27] wl[188] vdd gnd cell_6t
Xbit_r189_c27 bl[27] br[27] wl[189] vdd gnd cell_6t
Xbit_r190_c27 bl[27] br[27] wl[190] vdd gnd cell_6t
Xbit_r191_c27 bl[27] br[27] wl[191] vdd gnd cell_6t
Xbit_r192_c27 bl[27] br[27] wl[192] vdd gnd cell_6t
Xbit_r193_c27 bl[27] br[27] wl[193] vdd gnd cell_6t
Xbit_r194_c27 bl[27] br[27] wl[194] vdd gnd cell_6t
Xbit_r195_c27 bl[27] br[27] wl[195] vdd gnd cell_6t
Xbit_r196_c27 bl[27] br[27] wl[196] vdd gnd cell_6t
Xbit_r197_c27 bl[27] br[27] wl[197] vdd gnd cell_6t
Xbit_r198_c27 bl[27] br[27] wl[198] vdd gnd cell_6t
Xbit_r199_c27 bl[27] br[27] wl[199] vdd gnd cell_6t
Xbit_r200_c27 bl[27] br[27] wl[200] vdd gnd cell_6t
Xbit_r201_c27 bl[27] br[27] wl[201] vdd gnd cell_6t
Xbit_r202_c27 bl[27] br[27] wl[202] vdd gnd cell_6t
Xbit_r203_c27 bl[27] br[27] wl[203] vdd gnd cell_6t
Xbit_r204_c27 bl[27] br[27] wl[204] vdd gnd cell_6t
Xbit_r205_c27 bl[27] br[27] wl[205] vdd gnd cell_6t
Xbit_r206_c27 bl[27] br[27] wl[206] vdd gnd cell_6t
Xbit_r207_c27 bl[27] br[27] wl[207] vdd gnd cell_6t
Xbit_r208_c27 bl[27] br[27] wl[208] vdd gnd cell_6t
Xbit_r209_c27 bl[27] br[27] wl[209] vdd gnd cell_6t
Xbit_r210_c27 bl[27] br[27] wl[210] vdd gnd cell_6t
Xbit_r211_c27 bl[27] br[27] wl[211] vdd gnd cell_6t
Xbit_r212_c27 bl[27] br[27] wl[212] vdd gnd cell_6t
Xbit_r213_c27 bl[27] br[27] wl[213] vdd gnd cell_6t
Xbit_r214_c27 bl[27] br[27] wl[214] vdd gnd cell_6t
Xbit_r215_c27 bl[27] br[27] wl[215] vdd gnd cell_6t
Xbit_r216_c27 bl[27] br[27] wl[216] vdd gnd cell_6t
Xbit_r217_c27 bl[27] br[27] wl[217] vdd gnd cell_6t
Xbit_r218_c27 bl[27] br[27] wl[218] vdd gnd cell_6t
Xbit_r219_c27 bl[27] br[27] wl[219] vdd gnd cell_6t
Xbit_r220_c27 bl[27] br[27] wl[220] vdd gnd cell_6t
Xbit_r221_c27 bl[27] br[27] wl[221] vdd gnd cell_6t
Xbit_r222_c27 bl[27] br[27] wl[222] vdd gnd cell_6t
Xbit_r223_c27 bl[27] br[27] wl[223] vdd gnd cell_6t
Xbit_r224_c27 bl[27] br[27] wl[224] vdd gnd cell_6t
Xbit_r225_c27 bl[27] br[27] wl[225] vdd gnd cell_6t
Xbit_r226_c27 bl[27] br[27] wl[226] vdd gnd cell_6t
Xbit_r227_c27 bl[27] br[27] wl[227] vdd gnd cell_6t
Xbit_r228_c27 bl[27] br[27] wl[228] vdd gnd cell_6t
Xbit_r229_c27 bl[27] br[27] wl[229] vdd gnd cell_6t
Xbit_r230_c27 bl[27] br[27] wl[230] vdd gnd cell_6t
Xbit_r231_c27 bl[27] br[27] wl[231] vdd gnd cell_6t
Xbit_r232_c27 bl[27] br[27] wl[232] vdd gnd cell_6t
Xbit_r233_c27 bl[27] br[27] wl[233] vdd gnd cell_6t
Xbit_r234_c27 bl[27] br[27] wl[234] vdd gnd cell_6t
Xbit_r235_c27 bl[27] br[27] wl[235] vdd gnd cell_6t
Xbit_r236_c27 bl[27] br[27] wl[236] vdd gnd cell_6t
Xbit_r237_c27 bl[27] br[27] wl[237] vdd gnd cell_6t
Xbit_r238_c27 bl[27] br[27] wl[238] vdd gnd cell_6t
Xbit_r239_c27 bl[27] br[27] wl[239] vdd gnd cell_6t
Xbit_r240_c27 bl[27] br[27] wl[240] vdd gnd cell_6t
Xbit_r241_c27 bl[27] br[27] wl[241] vdd gnd cell_6t
Xbit_r242_c27 bl[27] br[27] wl[242] vdd gnd cell_6t
Xbit_r243_c27 bl[27] br[27] wl[243] vdd gnd cell_6t
Xbit_r244_c27 bl[27] br[27] wl[244] vdd gnd cell_6t
Xbit_r245_c27 bl[27] br[27] wl[245] vdd gnd cell_6t
Xbit_r246_c27 bl[27] br[27] wl[246] vdd gnd cell_6t
Xbit_r247_c27 bl[27] br[27] wl[247] vdd gnd cell_6t
Xbit_r248_c27 bl[27] br[27] wl[248] vdd gnd cell_6t
Xbit_r249_c27 bl[27] br[27] wl[249] vdd gnd cell_6t
Xbit_r250_c27 bl[27] br[27] wl[250] vdd gnd cell_6t
Xbit_r251_c27 bl[27] br[27] wl[251] vdd gnd cell_6t
Xbit_r252_c27 bl[27] br[27] wl[252] vdd gnd cell_6t
Xbit_r253_c27 bl[27] br[27] wl[253] vdd gnd cell_6t
Xbit_r254_c27 bl[27] br[27] wl[254] vdd gnd cell_6t
Xbit_r255_c27 bl[27] br[27] wl[255] vdd gnd cell_6t
Xbit_r0_c28 bl[28] br[28] wl[0] vdd gnd cell_6t
Xbit_r1_c28 bl[28] br[28] wl[1] vdd gnd cell_6t
Xbit_r2_c28 bl[28] br[28] wl[2] vdd gnd cell_6t
Xbit_r3_c28 bl[28] br[28] wl[3] vdd gnd cell_6t
Xbit_r4_c28 bl[28] br[28] wl[4] vdd gnd cell_6t
Xbit_r5_c28 bl[28] br[28] wl[5] vdd gnd cell_6t
Xbit_r6_c28 bl[28] br[28] wl[6] vdd gnd cell_6t
Xbit_r7_c28 bl[28] br[28] wl[7] vdd gnd cell_6t
Xbit_r8_c28 bl[28] br[28] wl[8] vdd gnd cell_6t
Xbit_r9_c28 bl[28] br[28] wl[9] vdd gnd cell_6t
Xbit_r10_c28 bl[28] br[28] wl[10] vdd gnd cell_6t
Xbit_r11_c28 bl[28] br[28] wl[11] vdd gnd cell_6t
Xbit_r12_c28 bl[28] br[28] wl[12] vdd gnd cell_6t
Xbit_r13_c28 bl[28] br[28] wl[13] vdd gnd cell_6t
Xbit_r14_c28 bl[28] br[28] wl[14] vdd gnd cell_6t
Xbit_r15_c28 bl[28] br[28] wl[15] vdd gnd cell_6t
Xbit_r16_c28 bl[28] br[28] wl[16] vdd gnd cell_6t
Xbit_r17_c28 bl[28] br[28] wl[17] vdd gnd cell_6t
Xbit_r18_c28 bl[28] br[28] wl[18] vdd gnd cell_6t
Xbit_r19_c28 bl[28] br[28] wl[19] vdd gnd cell_6t
Xbit_r20_c28 bl[28] br[28] wl[20] vdd gnd cell_6t
Xbit_r21_c28 bl[28] br[28] wl[21] vdd gnd cell_6t
Xbit_r22_c28 bl[28] br[28] wl[22] vdd gnd cell_6t
Xbit_r23_c28 bl[28] br[28] wl[23] vdd gnd cell_6t
Xbit_r24_c28 bl[28] br[28] wl[24] vdd gnd cell_6t
Xbit_r25_c28 bl[28] br[28] wl[25] vdd gnd cell_6t
Xbit_r26_c28 bl[28] br[28] wl[26] vdd gnd cell_6t
Xbit_r27_c28 bl[28] br[28] wl[27] vdd gnd cell_6t
Xbit_r28_c28 bl[28] br[28] wl[28] vdd gnd cell_6t
Xbit_r29_c28 bl[28] br[28] wl[29] vdd gnd cell_6t
Xbit_r30_c28 bl[28] br[28] wl[30] vdd gnd cell_6t
Xbit_r31_c28 bl[28] br[28] wl[31] vdd gnd cell_6t
Xbit_r32_c28 bl[28] br[28] wl[32] vdd gnd cell_6t
Xbit_r33_c28 bl[28] br[28] wl[33] vdd gnd cell_6t
Xbit_r34_c28 bl[28] br[28] wl[34] vdd gnd cell_6t
Xbit_r35_c28 bl[28] br[28] wl[35] vdd gnd cell_6t
Xbit_r36_c28 bl[28] br[28] wl[36] vdd gnd cell_6t
Xbit_r37_c28 bl[28] br[28] wl[37] vdd gnd cell_6t
Xbit_r38_c28 bl[28] br[28] wl[38] vdd gnd cell_6t
Xbit_r39_c28 bl[28] br[28] wl[39] vdd gnd cell_6t
Xbit_r40_c28 bl[28] br[28] wl[40] vdd gnd cell_6t
Xbit_r41_c28 bl[28] br[28] wl[41] vdd gnd cell_6t
Xbit_r42_c28 bl[28] br[28] wl[42] vdd gnd cell_6t
Xbit_r43_c28 bl[28] br[28] wl[43] vdd gnd cell_6t
Xbit_r44_c28 bl[28] br[28] wl[44] vdd gnd cell_6t
Xbit_r45_c28 bl[28] br[28] wl[45] vdd gnd cell_6t
Xbit_r46_c28 bl[28] br[28] wl[46] vdd gnd cell_6t
Xbit_r47_c28 bl[28] br[28] wl[47] vdd gnd cell_6t
Xbit_r48_c28 bl[28] br[28] wl[48] vdd gnd cell_6t
Xbit_r49_c28 bl[28] br[28] wl[49] vdd gnd cell_6t
Xbit_r50_c28 bl[28] br[28] wl[50] vdd gnd cell_6t
Xbit_r51_c28 bl[28] br[28] wl[51] vdd gnd cell_6t
Xbit_r52_c28 bl[28] br[28] wl[52] vdd gnd cell_6t
Xbit_r53_c28 bl[28] br[28] wl[53] vdd gnd cell_6t
Xbit_r54_c28 bl[28] br[28] wl[54] vdd gnd cell_6t
Xbit_r55_c28 bl[28] br[28] wl[55] vdd gnd cell_6t
Xbit_r56_c28 bl[28] br[28] wl[56] vdd gnd cell_6t
Xbit_r57_c28 bl[28] br[28] wl[57] vdd gnd cell_6t
Xbit_r58_c28 bl[28] br[28] wl[58] vdd gnd cell_6t
Xbit_r59_c28 bl[28] br[28] wl[59] vdd gnd cell_6t
Xbit_r60_c28 bl[28] br[28] wl[60] vdd gnd cell_6t
Xbit_r61_c28 bl[28] br[28] wl[61] vdd gnd cell_6t
Xbit_r62_c28 bl[28] br[28] wl[62] vdd gnd cell_6t
Xbit_r63_c28 bl[28] br[28] wl[63] vdd gnd cell_6t
Xbit_r64_c28 bl[28] br[28] wl[64] vdd gnd cell_6t
Xbit_r65_c28 bl[28] br[28] wl[65] vdd gnd cell_6t
Xbit_r66_c28 bl[28] br[28] wl[66] vdd gnd cell_6t
Xbit_r67_c28 bl[28] br[28] wl[67] vdd gnd cell_6t
Xbit_r68_c28 bl[28] br[28] wl[68] vdd gnd cell_6t
Xbit_r69_c28 bl[28] br[28] wl[69] vdd gnd cell_6t
Xbit_r70_c28 bl[28] br[28] wl[70] vdd gnd cell_6t
Xbit_r71_c28 bl[28] br[28] wl[71] vdd gnd cell_6t
Xbit_r72_c28 bl[28] br[28] wl[72] vdd gnd cell_6t
Xbit_r73_c28 bl[28] br[28] wl[73] vdd gnd cell_6t
Xbit_r74_c28 bl[28] br[28] wl[74] vdd gnd cell_6t
Xbit_r75_c28 bl[28] br[28] wl[75] vdd gnd cell_6t
Xbit_r76_c28 bl[28] br[28] wl[76] vdd gnd cell_6t
Xbit_r77_c28 bl[28] br[28] wl[77] vdd gnd cell_6t
Xbit_r78_c28 bl[28] br[28] wl[78] vdd gnd cell_6t
Xbit_r79_c28 bl[28] br[28] wl[79] vdd gnd cell_6t
Xbit_r80_c28 bl[28] br[28] wl[80] vdd gnd cell_6t
Xbit_r81_c28 bl[28] br[28] wl[81] vdd gnd cell_6t
Xbit_r82_c28 bl[28] br[28] wl[82] vdd gnd cell_6t
Xbit_r83_c28 bl[28] br[28] wl[83] vdd gnd cell_6t
Xbit_r84_c28 bl[28] br[28] wl[84] vdd gnd cell_6t
Xbit_r85_c28 bl[28] br[28] wl[85] vdd gnd cell_6t
Xbit_r86_c28 bl[28] br[28] wl[86] vdd gnd cell_6t
Xbit_r87_c28 bl[28] br[28] wl[87] vdd gnd cell_6t
Xbit_r88_c28 bl[28] br[28] wl[88] vdd gnd cell_6t
Xbit_r89_c28 bl[28] br[28] wl[89] vdd gnd cell_6t
Xbit_r90_c28 bl[28] br[28] wl[90] vdd gnd cell_6t
Xbit_r91_c28 bl[28] br[28] wl[91] vdd gnd cell_6t
Xbit_r92_c28 bl[28] br[28] wl[92] vdd gnd cell_6t
Xbit_r93_c28 bl[28] br[28] wl[93] vdd gnd cell_6t
Xbit_r94_c28 bl[28] br[28] wl[94] vdd gnd cell_6t
Xbit_r95_c28 bl[28] br[28] wl[95] vdd gnd cell_6t
Xbit_r96_c28 bl[28] br[28] wl[96] vdd gnd cell_6t
Xbit_r97_c28 bl[28] br[28] wl[97] vdd gnd cell_6t
Xbit_r98_c28 bl[28] br[28] wl[98] vdd gnd cell_6t
Xbit_r99_c28 bl[28] br[28] wl[99] vdd gnd cell_6t
Xbit_r100_c28 bl[28] br[28] wl[100] vdd gnd cell_6t
Xbit_r101_c28 bl[28] br[28] wl[101] vdd gnd cell_6t
Xbit_r102_c28 bl[28] br[28] wl[102] vdd gnd cell_6t
Xbit_r103_c28 bl[28] br[28] wl[103] vdd gnd cell_6t
Xbit_r104_c28 bl[28] br[28] wl[104] vdd gnd cell_6t
Xbit_r105_c28 bl[28] br[28] wl[105] vdd gnd cell_6t
Xbit_r106_c28 bl[28] br[28] wl[106] vdd gnd cell_6t
Xbit_r107_c28 bl[28] br[28] wl[107] vdd gnd cell_6t
Xbit_r108_c28 bl[28] br[28] wl[108] vdd gnd cell_6t
Xbit_r109_c28 bl[28] br[28] wl[109] vdd gnd cell_6t
Xbit_r110_c28 bl[28] br[28] wl[110] vdd gnd cell_6t
Xbit_r111_c28 bl[28] br[28] wl[111] vdd gnd cell_6t
Xbit_r112_c28 bl[28] br[28] wl[112] vdd gnd cell_6t
Xbit_r113_c28 bl[28] br[28] wl[113] vdd gnd cell_6t
Xbit_r114_c28 bl[28] br[28] wl[114] vdd gnd cell_6t
Xbit_r115_c28 bl[28] br[28] wl[115] vdd gnd cell_6t
Xbit_r116_c28 bl[28] br[28] wl[116] vdd gnd cell_6t
Xbit_r117_c28 bl[28] br[28] wl[117] vdd gnd cell_6t
Xbit_r118_c28 bl[28] br[28] wl[118] vdd gnd cell_6t
Xbit_r119_c28 bl[28] br[28] wl[119] vdd gnd cell_6t
Xbit_r120_c28 bl[28] br[28] wl[120] vdd gnd cell_6t
Xbit_r121_c28 bl[28] br[28] wl[121] vdd gnd cell_6t
Xbit_r122_c28 bl[28] br[28] wl[122] vdd gnd cell_6t
Xbit_r123_c28 bl[28] br[28] wl[123] vdd gnd cell_6t
Xbit_r124_c28 bl[28] br[28] wl[124] vdd gnd cell_6t
Xbit_r125_c28 bl[28] br[28] wl[125] vdd gnd cell_6t
Xbit_r126_c28 bl[28] br[28] wl[126] vdd gnd cell_6t
Xbit_r127_c28 bl[28] br[28] wl[127] vdd gnd cell_6t
Xbit_r128_c28 bl[28] br[28] wl[128] vdd gnd cell_6t
Xbit_r129_c28 bl[28] br[28] wl[129] vdd gnd cell_6t
Xbit_r130_c28 bl[28] br[28] wl[130] vdd gnd cell_6t
Xbit_r131_c28 bl[28] br[28] wl[131] vdd gnd cell_6t
Xbit_r132_c28 bl[28] br[28] wl[132] vdd gnd cell_6t
Xbit_r133_c28 bl[28] br[28] wl[133] vdd gnd cell_6t
Xbit_r134_c28 bl[28] br[28] wl[134] vdd gnd cell_6t
Xbit_r135_c28 bl[28] br[28] wl[135] vdd gnd cell_6t
Xbit_r136_c28 bl[28] br[28] wl[136] vdd gnd cell_6t
Xbit_r137_c28 bl[28] br[28] wl[137] vdd gnd cell_6t
Xbit_r138_c28 bl[28] br[28] wl[138] vdd gnd cell_6t
Xbit_r139_c28 bl[28] br[28] wl[139] vdd gnd cell_6t
Xbit_r140_c28 bl[28] br[28] wl[140] vdd gnd cell_6t
Xbit_r141_c28 bl[28] br[28] wl[141] vdd gnd cell_6t
Xbit_r142_c28 bl[28] br[28] wl[142] vdd gnd cell_6t
Xbit_r143_c28 bl[28] br[28] wl[143] vdd gnd cell_6t
Xbit_r144_c28 bl[28] br[28] wl[144] vdd gnd cell_6t
Xbit_r145_c28 bl[28] br[28] wl[145] vdd gnd cell_6t
Xbit_r146_c28 bl[28] br[28] wl[146] vdd gnd cell_6t
Xbit_r147_c28 bl[28] br[28] wl[147] vdd gnd cell_6t
Xbit_r148_c28 bl[28] br[28] wl[148] vdd gnd cell_6t
Xbit_r149_c28 bl[28] br[28] wl[149] vdd gnd cell_6t
Xbit_r150_c28 bl[28] br[28] wl[150] vdd gnd cell_6t
Xbit_r151_c28 bl[28] br[28] wl[151] vdd gnd cell_6t
Xbit_r152_c28 bl[28] br[28] wl[152] vdd gnd cell_6t
Xbit_r153_c28 bl[28] br[28] wl[153] vdd gnd cell_6t
Xbit_r154_c28 bl[28] br[28] wl[154] vdd gnd cell_6t
Xbit_r155_c28 bl[28] br[28] wl[155] vdd gnd cell_6t
Xbit_r156_c28 bl[28] br[28] wl[156] vdd gnd cell_6t
Xbit_r157_c28 bl[28] br[28] wl[157] vdd gnd cell_6t
Xbit_r158_c28 bl[28] br[28] wl[158] vdd gnd cell_6t
Xbit_r159_c28 bl[28] br[28] wl[159] vdd gnd cell_6t
Xbit_r160_c28 bl[28] br[28] wl[160] vdd gnd cell_6t
Xbit_r161_c28 bl[28] br[28] wl[161] vdd gnd cell_6t
Xbit_r162_c28 bl[28] br[28] wl[162] vdd gnd cell_6t
Xbit_r163_c28 bl[28] br[28] wl[163] vdd gnd cell_6t
Xbit_r164_c28 bl[28] br[28] wl[164] vdd gnd cell_6t
Xbit_r165_c28 bl[28] br[28] wl[165] vdd gnd cell_6t
Xbit_r166_c28 bl[28] br[28] wl[166] vdd gnd cell_6t
Xbit_r167_c28 bl[28] br[28] wl[167] vdd gnd cell_6t
Xbit_r168_c28 bl[28] br[28] wl[168] vdd gnd cell_6t
Xbit_r169_c28 bl[28] br[28] wl[169] vdd gnd cell_6t
Xbit_r170_c28 bl[28] br[28] wl[170] vdd gnd cell_6t
Xbit_r171_c28 bl[28] br[28] wl[171] vdd gnd cell_6t
Xbit_r172_c28 bl[28] br[28] wl[172] vdd gnd cell_6t
Xbit_r173_c28 bl[28] br[28] wl[173] vdd gnd cell_6t
Xbit_r174_c28 bl[28] br[28] wl[174] vdd gnd cell_6t
Xbit_r175_c28 bl[28] br[28] wl[175] vdd gnd cell_6t
Xbit_r176_c28 bl[28] br[28] wl[176] vdd gnd cell_6t
Xbit_r177_c28 bl[28] br[28] wl[177] vdd gnd cell_6t
Xbit_r178_c28 bl[28] br[28] wl[178] vdd gnd cell_6t
Xbit_r179_c28 bl[28] br[28] wl[179] vdd gnd cell_6t
Xbit_r180_c28 bl[28] br[28] wl[180] vdd gnd cell_6t
Xbit_r181_c28 bl[28] br[28] wl[181] vdd gnd cell_6t
Xbit_r182_c28 bl[28] br[28] wl[182] vdd gnd cell_6t
Xbit_r183_c28 bl[28] br[28] wl[183] vdd gnd cell_6t
Xbit_r184_c28 bl[28] br[28] wl[184] vdd gnd cell_6t
Xbit_r185_c28 bl[28] br[28] wl[185] vdd gnd cell_6t
Xbit_r186_c28 bl[28] br[28] wl[186] vdd gnd cell_6t
Xbit_r187_c28 bl[28] br[28] wl[187] vdd gnd cell_6t
Xbit_r188_c28 bl[28] br[28] wl[188] vdd gnd cell_6t
Xbit_r189_c28 bl[28] br[28] wl[189] vdd gnd cell_6t
Xbit_r190_c28 bl[28] br[28] wl[190] vdd gnd cell_6t
Xbit_r191_c28 bl[28] br[28] wl[191] vdd gnd cell_6t
Xbit_r192_c28 bl[28] br[28] wl[192] vdd gnd cell_6t
Xbit_r193_c28 bl[28] br[28] wl[193] vdd gnd cell_6t
Xbit_r194_c28 bl[28] br[28] wl[194] vdd gnd cell_6t
Xbit_r195_c28 bl[28] br[28] wl[195] vdd gnd cell_6t
Xbit_r196_c28 bl[28] br[28] wl[196] vdd gnd cell_6t
Xbit_r197_c28 bl[28] br[28] wl[197] vdd gnd cell_6t
Xbit_r198_c28 bl[28] br[28] wl[198] vdd gnd cell_6t
Xbit_r199_c28 bl[28] br[28] wl[199] vdd gnd cell_6t
Xbit_r200_c28 bl[28] br[28] wl[200] vdd gnd cell_6t
Xbit_r201_c28 bl[28] br[28] wl[201] vdd gnd cell_6t
Xbit_r202_c28 bl[28] br[28] wl[202] vdd gnd cell_6t
Xbit_r203_c28 bl[28] br[28] wl[203] vdd gnd cell_6t
Xbit_r204_c28 bl[28] br[28] wl[204] vdd gnd cell_6t
Xbit_r205_c28 bl[28] br[28] wl[205] vdd gnd cell_6t
Xbit_r206_c28 bl[28] br[28] wl[206] vdd gnd cell_6t
Xbit_r207_c28 bl[28] br[28] wl[207] vdd gnd cell_6t
Xbit_r208_c28 bl[28] br[28] wl[208] vdd gnd cell_6t
Xbit_r209_c28 bl[28] br[28] wl[209] vdd gnd cell_6t
Xbit_r210_c28 bl[28] br[28] wl[210] vdd gnd cell_6t
Xbit_r211_c28 bl[28] br[28] wl[211] vdd gnd cell_6t
Xbit_r212_c28 bl[28] br[28] wl[212] vdd gnd cell_6t
Xbit_r213_c28 bl[28] br[28] wl[213] vdd gnd cell_6t
Xbit_r214_c28 bl[28] br[28] wl[214] vdd gnd cell_6t
Xbit_r215_c28 bl[28] br[28] wl[215] vdd gnd cell_6t
Xbit_r216_c28 bl[28] br[28] wl[216] vdd gnd cell_6t
Xbit_r217_c28 bl[28] br[28] wl[217] vdd gnd cell_6t
Xbit_r218_c28 bl[28] br[28] wl[218] vdd gnd cell_6t
Xbit_r219_c28 bl[28] br[28] wl[219] vdd gnd cell_6t
Xbit_r220_c28 bl[28] br[28] wl[220] vdd gnd cell_6t
Xbit_r221_c28 bl[28] br[28] wl[221] vdd gnd cell_6t
Xbit_r222_c28 bl[28] br[28] wl[222] vdd gnd cell_6t
Xbit_r223_c28 bl[28] br[28] wl[223] vdd gnd cell_6t
Xbit_r224_c28 bl[28] br[28] wl[224] vdd gnd cell_6t
Xbit_r225_c28 bl[28] br[28] wl[225] vdd gnd cell_6t
Xbit_r226_c28 bl[28] br[28] wl[226] vdd gnd cell_6t
Xbit_r227_c28 bl[28] br[28] wl[227] vdd gnd cell_6t
Xbit_r228_c28 bl[28] br[28] wl[228] vdd gnd cell_6t
Xbit_r229_c28 bl[28] br[28] wl[229] vdd gnd cell_6t
Xbit_r230_c28 bl[28] br[28] wl[230] vdd gnd cell_6t
Xbit_r231_c28 bl[28] br[28] wl[231] vdd gnd cell_6t
Xbit_r232_c28 bl[28] br[28] wl[232] vdd gnd cell_6t
Xbit_r233_c28 bl[28] br[28] wl[233] vdd gnd cell_6t
Xbit_r234_c28 bl[28] br[28] wl[234] vdd gnd cell_6t
Xbit_r235_c28 bl[28] br[28] wl[235] vdd gnd cell_6t
Xbit_r236_c28 bl[28] br[28] wl[236] vdd gnd cell_6t
Xbit_r237_c28 bl[28] br[28] wl[237] vdd gnd cell_6t
Xbit_r238_c28 bl[28] br[28] wl[238] vdd gnd cell_6t
Xbit_r239_c28 bl[28] br[28] wl[239] vdd gnd cell_6t
Xbit_r240_c28 bl[28] br[28] wl[240] vdd gnd cell_6t
Xbit_r241_c28 bl[28] br[28] wl[241] vdd gnd cell_6t
Xbit_r242_c28 bl[28] br[28] wl[242] vdd gnd cell_6t
Xbit_r243_c28 bl[28] br[28] wl[243] vdd gnd cell_6t
Xbit_r244_c28 bl[28] br[28] wl[244] vdd gnd cell_6t
Xbit_r245_c28 bl[28] br[28] wl[245] vdd gnd cell_6t
Xbit_r246_c28 bl[28] br[28] wl[246] vdd gnd cell_6t
Xbit_r247_c28 bl[28] br[28] wl[247] vdd gnd cell_6t
Xbit_r248_c28 bl[28] br[28] wl[248] vdd gnd cell_6t
Xbit_r249_c28 bl[28] br[28] wl[249] vdd gnd cell_6t
Xbit_r250_c28 bl[28] br[28] wl[250] vdd gnd cell_6t
Xbit_r251_c28 bl[28] br[28] wl[251] vdd gnd cell_6t
Xbit_r252_c28 bl[28] br[28] wl[252] vdd gnd cell_6t
Xbit_r253_c28 bl[28] br[28] wl[253] vdd gnd cell_6t
Xbit_r254_c28 bl[28] br[28] wl[254] vdd gnd cell_6t
Xbit_r255_c28 bl[28] br[28] wl[255] vdd gnd cell_6t
Xbit_r0_c29 bl[29] br[29] wl[0] vdd gnd cell_6t
Xbit_r1_c29 bl[29] br[29] wl[1] vdd gnd cell_6t
Xbit_r2_c29 bl[29] br[29] wl[2] vdd gnd cell_6t
Xbit_r3_c29 bl[29] br[29] wl[3] vdd gnd cell_6t
Xbit_r4_c29 bl[29] br[29] wl[4] vdd gnd cell_6t
Xbit_r5_c29 bl[29] br[29] wl[5] vdd gnd cell_6t
Xbit_r6_c29 bl[29] br[29] wl[6] vdd gnd cell_6t
Xbit_r7_c29 bl[29] br[29] wl[7] vdd gnd cell_6t
Xbit_r8_c29 bl[29] br[29] wl[8] vdd gnd cell_6t
Xbit_r9_c29 bl[29] br[29] wl[9] vdd gnd cell_6t
Xbit_r10_c29 bl[29] br[29] wl[10] vdd gnd cell_6t
Xbit_r11_c29 bl[29] br[29] wl[11] vdd gnd cell_6t
Xbit_r12_c29 bl[29] br[29] wl[12] vdd gnd cell_6t
Xbit_r13_c29 bl[29] br[29] wl[13] vdd gnd cell_6t
Xbit_r14_c29 bl[29] br[29] wl[14] vdd gnd cell_6t
Xbit_r15_c29 bl[29] br[29] wl[15] vdd gnd cell_6t
Xbit_r16_c29 bl[29] br[29] wl[16] vdd gnd cell_6t
Xbit_r17_c29 bl[29] br[29] wl[17] vdd gnd cell_6t
Xbit_r18_c29 bl[29] br[29] wl[18] vdd gnd cell_6t
Xbit_r19_c29 bl[29] br[29] wl[19] vdd gnd cell_6t
Xbit_r20_c29 bl[29] br[29] wl[20] vdd gnd cell_6t
Xbit_r21_c29 bl[29] br[29] wl[21] vdd gnd cell_6t
Xbit_r22_c29 bl[29] br[29] wl[22] vdd gnd cell_6t
Xbit_r23_c29 bl[29] br[29] wl[23] vdd gnd cell_6t
Xbit_r24_c29 bl[29] br[29] wl[24] vdd gnd cell_6t
Xbit_r25_c29 bl[29] br[29] wl[25] vdd gnd cell_6t
Xbit_r26_c29 bl[29] br[29] wl[26] vdd gnd cell_6t
Xbit_r27_c29 bl[29] br[29] wl[27] vdd gnd cell_6t
Xbit_r28_c29 bl[29] br[29] wl[28] vdd gnd cell_6t
Xbit_r29_c29 bl[29] br[29] wl[29] vdd gnd cell_6t
Xbit_r30_c29 bl[29] br[29] wl[30] vdd gnd cell_6t
Xbit_r31_c29 bl[29] br[29] wl[31] vdd gnd cell_6t
Xbit_r32_c29 bl[29] br[29] wl[32] vdd gnd cell_6t
Xbit_r33_c29 bl[29] br[29] wl[33] vdd gnd cell_6t
Xbit_r34_c29 bl[29] br[29] wl[34] vdd gnd cell_6t
Xbit_r35_c29 bl[29] br[29] wl[35] vdd gnd cell_6t
Xbit_r36_c29 bl[29] br[29] wl[36] vdd gnd cell_6t
Xbit_r37_c29 bl[29] br[29] wl[37] vdd gnd cell_6t
Xbit_r38_c29 bl[29] br[29] wl[38] vdd gnd cell_6t
Xbit_r39_c29 bl[29] br[29] wl[39] vdd gnd cell_6t
Xbit_r40_c29 bl[29] br[29] wl[40] vdd gnd cell_6t
Xbit_r41_c29 bl[29] br[29] wl[41] vdd gnd cell_6t
Xbit_r42_c29 bl[29] br[29] wl[42] vdd gnd cell_6t
Xbit_r43_c29 bl[29] br[29] wl[43] vdd gnd cell_6t
Xbit_r44_c29 bl[29] br[29] wl[44] vdd gnd cell_6t
Xbit_r45_c29 bl[29] br[29] wl[45] vdd gnd cell_6t
Xbit_r46_c29 bl[29] br[29] wl[46] vdd gnd cell_6t
Xbit_r47_c29 bl[29] br[29] wl[47] vdd gnd cell_6t
Xbit_r48_c29 bl[29] br[29] wl[48] vdd gnd cell_6t
Xbit_r49_c29 bl[29] br[29] wl[49] vdd gnd cell_6t
Xbit_r50_c29 bl[29] br[29] wl[50] vdd gnd cell_6t
Xbit_r51_c29 bl[29] br[29] wl[51] vdd gnd cell_6t
Xbit_r52_c29 bl[29] br[29] wl[52] vdd gnd cell_6t
Xbit_r53_c29 bl[29] br[29] wl[53] vdd gnd cell_6t
Xbit_r54_c29 bl[29] br[29] wl[54] vdd gnd cell_6t
Xbit_r55_c29 bl[29] br[29] wl[55] vdd gnd cell_6t
Xbit_r56_c29 bl[29] br[29] wl[56] vdd gnd cell_6t
Xbit_r57_c29 bl[29] br[29] wl[57] vdd gnd cell_6t
Xbit_r58_c29 bl[29] br[29] wl[58] vdd gnd cell_6t
Xbit_r59_c29 bl[29] br[29] wl[59] vdd gnd cell_6t
Xbit_r60_c29 bl[29] br[29] wl[60] vdd gnd cell_6t
Xbit_r61_c29 bl[29] br[29] wl[61] vdd gnd cell_6t
Xbit_r62_c29 bl[29] br[29] wl[62] vdd gnd cell_6t
Xbit_r63_c29 bl[29] br[29] wl[63] vdd gnd cell_6t
Xbit_r64_c29 bl[29] br[29] wl[64] vdd gnd cell_6t
Xbit_r65_c29 bl[29] br[29] wl[65] vdd gnd cell_6t
Xbit_r66_c29 bl[29] br[29] wl[66] vdd gnd cell_6t
Xbit_r67_c29 bl[29] br[29] wl[67] vdd gnd cell_6t
Xbit_r68_c29 bl[29] br[29] wl[68] vdd gnd cell_6t
Xbit_r69_c29 bl[29] br[29] wl[69] vdd gnd cell_6t
Xbit_r70_c29 bl[29] br[29] wl[70] vdd gnd cell_6t
Xbit_r71_c29 bl[29] br[29] wl[71] vdd gnd cell_6t
Xbit_r72_c29 bl[29] br[29] wl[72] vdd gnd cell_6t
Xbit_r73_c29 bl[29] br[29] wl[73] vdd gnd cell_6t
Xbit_r74_c29 bl[29] br[29] wl[74] vdd gnd cell_6t
Xbit_r75_c29 bl[29] br[29] wl[75] vdd gnd cell_6t
Xbit_r76_c29 bl[29] br[29] wl[76] vdd gnd cell_6t
Xbit_r77_c29 bl[29] br[29] wl[77] vdd gnd cell_6t
Xbit_r78_c29 bl[29] br[29] wl[78] vdd gnd cell_6t
Xbit_r79_c29 bl[29] br[29] wl[79] vdd gnd cell_6t
Xbit_r80_c29 bl[29] br[29] wl[80] vdd gnd cell_6t
Xbit_r81_c29 bl[29] br[29] wl[81] vdd gnd cell_6t
Xbit_r82_c29 bl[29] br[29] wl[82] vdd gnd cell_6t
Xbit_r83_c29 bl[29] br[29] wl[83] vdd gnd cell_6t
Xbit_r84_c29 bl[29] br[29] wl[84] vdd gnd cell_6t
Xbit_r85_c29 bl[29] br[29] wl[85] vdd gnd cell_6t
Xbit_r86_c29 bl[29] br[29] wl[86] vdd gnd cell_6t
Xbit_r87_c29 bl[29] br[29] wl[87] vdd gnd cell_6t
Xbit_r88_c29 bl[29] br[29] wl[88] vdd gnd cell_6t
Xbit_r89_c29 bl[29] br[29] wl[89] vdd gnd cell_6t
Xbit_r90_c29 bl[29] br[29] wl[90] vdd gnd cell_6t
Xbit_r91_c29 bl[29] br[29] wl[91] vdd gnd cell_6t
Xbit_r92_c29 bl[29] br[29] wl[92] vdd gnd cell_6t
Xbit_r93_c29 bl[29] br[29] wl[93] vdd gnd cell_6t
Xbit_r94_c29 bl[29] br[29] wl[94] vdd gnd cell_6t
Xbit_r95_c29 bl[29] br[29] wl[95] vdd gnd cell_6t
Xbit_r96_c29 bl[29] br[29] wl[96] vdd gnd cell_6t
Xbit_r97_c29 bl[29] br[29] wl[97] vdd gnd cell_6t
Xbit_r98_c29 bl[29] br[29] wl[98] vdd gnd cell_6t
Xbit_r99_c29 bl[29] br[29] wl[99] vdd gnd cell_6t
Xbit_r100_c29 bl[29] br[29] wl[100] vdd gnd cell_6t
Xbit_r101_c29 bl[29] br[29] wl[101] vdd gnd cell_6t
Xbit_r102_c29 bl[29] br[29] wl[102] vdd gnd cell_6t
Xbit_r103_c29 bl[29] br[29] wl[103] vdd gnd cell_6t
Xbit_r104_c29 bl[29] br[29] wl[104] vdd gnd cell_6t
Xbit_r105_c29 bl[29] br[29] wl[105] vdd gnd cell_6t
Xbit_r106_c29 bl[29] br[29] wl[106] vdd gnd cell_6t
Xbit_r107_c29 bl[29] br[29] wl[107] vdd gnd cell_6t
Xbit_r108_c29 bl[29] br[29] wl[108] vdd gnd cell_6t
Xbit_r109_c29 bl[29] br[29] wl[109] vdd gnd cell_6t
Xbit_r110_c29 bl[29] br[29] wl[110] vdd gnd cell_6t
Xbit_r111_c29 bl[29] br[29] wl[111] vdd gnd cell_6t
Xbit_r112_c29 bl[29] br[29] wl[112] vdd gnd cell_6t
Xbit_r113_c29 bl[29] br[29] wl[113] vdd gnd cell_6t
Xbit_r114_c29 bl[29] br[29] wl[114] vdd gnd cell_6t
Xbit_r115_c29 bl[29] br[29] wl[115] vdd gnd cell_6t
Xbit_r116_c29 bl[29] br[29] wl[116] vdd gnd cell_6t
Xbit_r117_c29 bl[29] br[29] wl[117] vdd gnd cell_6t
Xbit_r118_c29 bl[29] br[29] wl[118] vdd gnd cell_6t
Xbit_r119_c29 bl[29] br[29] wl[119] vdd gnd cell_6t
Xbit_r120_c29 bl[29] br[29] wl[120] vdd gnd cell_6t
Xbit_r121_c29 bl[29] br[29] wl[121] vdd gnd cell_6t
Xbit_r122_c29 bl[29] br[29] wl[122] vdd gnd cell_6t
Xbit_r123_c29 bl[29] br[29] wl[123] vdd gnd cell_6t
Xbit_r124_c29 bl[29] br[29] wl[124] vdd gnd cell_6t
Xbit_r125_c29 bl[29] br[29] wl[125] vdd gnd cell_6t
Xbit_r126_c29 bl[29] br[29] wl[126] vdd gnd cell_6t
Xbit_r127_c29 bl[29] br[29] wl[127] vdd gnd cell_6t
Xbit_r128_c29 bl[29] br[29] wl[128] vdd gnd cell_6t
Xbit_r129_c29 bl[29] br[29] wl[129] vdd gnd cell_6t
Xbit_r130_c29 bl[29] br[29] wl[130] vdd gnd cell_6t
Xbit_r131_c29 bl[29] br[29] wl[131] vdd gnd cell_6t
Xbit_r132_c29 bl[29] br[29] wl[132] vdd gnd cell_6t
Xbit_r133_c29 bl[29] br[29] wl[133] vdd gnd cell_6t
Xbit_r134_c29 bl[29] br[29] wl[134] vdd gnd cell_6t
Xbit_r135_c29 bl[29] br[29] wl[135] vdd gnd cell_6t
Xbit_r136_c29 bl[29] br[29] wl[136] vdd gnd cell_6t
Xbit_r137_c29 bl[29] br[29] wl[137] vdd gnd cell_6t
Xbit_r138_c29 bl[29] br[29] wl[138] vdd gnd cell_6t
Xbit_r139_c29 bl[29] br[29] wl[139] vdd gnd cell_6t
Xbit_r140_c29 bl[29] br[29] wl[140] vdd gnd cell_6t
Xbit_r141_c29 bl[29] br[29] wl[141] vdd gnd cell_6t
Xbit_r142_c29 bl[29] br[29] wl[142] vdd gnd cell_6t
Xbit_r143_c29 bl[29] br[29] wl[143] vdd gnd cell_6t
Xbit_r144_c29 bl[29] br[29] wl[144] vdd gnd cell_6t
Xbit_r145_c29 bl[29] br[29] wl[145] vdd gnd cell_6t
Xbit_r146_c29 bl[29] br[29] wl[146] vdd gnd cell_6t
Xbit_r147_c29 bl[29] br[29] wl[147] vdd gnd cell_6t
Xbit_r148_c29 bl[29] br[29] wl[148] vdd gnd cell_6t
Xbit_r149_c29 bl[29] br[29] wl[149] vdd gnd cell_6t
Xbit_r150_c29 bl[29] br[29] wl[150] vdd gnd cell_6t
Xbit_r151_c29 bl[29] br[29] wl[151] vdd gnd cell_6t
Xbit_r152_c29 bl[29] br[29] wl[152] vdd gnd cell_6t
Xbit_r153_c29 bl[29] br[29] wl[153] vdd gnd cell_6t
Xbit_r154_c29 bl[29] br[29] wl[154] vdd gnd cell_6t
Xbit_r155_c29 bl[29] br[29] wl[155] vdd gnd cell_6t
Xbit_r156_c29 bl[29] br[29] wl[156] vdd gnd cell_6t
Xbit_r157_c29 bl[29] br[29] wl[157] vdd gnd cell_6t
Xbit_r158_c29 bl[29] br[29] wl[158] vdd gnd cell_6t
Xbit_r159_c29 bl[29] br[29] wl[159] vdd gnd cell_6t
Xbit_r160_c29 bl[29] br[29] wl[160] vdd gnd cell_6t
Xbit_r161_c29 bl[29] br[29] wl[161] vdd gnd cell_6t
Xbit_r162_c29 bl[29] br[29] wl[162] vdd gnd cell_6t
Xbit_r163_c29 bl[29] br[29] wl[163] vdd gnd cell_6t
Xbit_r164_c29 bl[29] br[29] wl[164] vdd gnd cell_6t
Xbit_r165_c29 bl[29] br[29] wl[165] vdd gnd cell_6t
Xbit_r166_c29 bl[29] br[29] wl[166] vdd gnd cell_6t
Xbit_r167_c29 bl[29] br[29] wl[167] vdd gnd cell_6t
Xbit_r168_c29 bl[29] br[29] wl[168] vdd gnd cell_6t
Xbit_r169_c29 bl[29] br[29] wl[169] vdd gnd cell_6t
Xbit_r170_c29 bl[29] br[29] wl[170] vdd gnd cell_6t
Xbit_r171_c29 bl[29] br[29] wl[171] vdd gnd cell_6t
Xbit_r172_c29 bl[29] br[29] wl[172] vdd gnd cell_6t
Xbit_r173_c29 bl[29] br[29] wl[173] vdd gnd cell_6t
Xbit_r174_c29 bl[29] br[29] wl[174] vdd gnd cell_6t
Xbit_r175_c29 bl[29] br[29] wl[175] vdd gnd cell_6t
Xbit_r176_c29 bl[29] br[29] wl[176] vdd gnd cell_6t
Xbit_r177_c29 bl[29] br[29] wl[177] vdd gnd cell_6t
Xbit_r178_c29 bl[29] br[29] wl[178] vdd gnd cell_6t
Xbit_r179_c29 bl[29] br[29] wl[179] vdd gnd cell_6t
Xbit_r180_c29 bl[29] br[29] wl[180] vdd gnd cell_6t
Xbit_r181_c29 bl[29] br[29] wl[181] vdd gnd cell_6t
Xbit_r182_c29 bl[29] br[29] wl[182] vdd gnd cell_6t
Xbit_r183_c29 bl[29] br[29] wl[183] vdd gnd cell_6t
Xbit_r184_c29 bl[29] br[29] wl[184] vdd gnd cell_6t
Xbit_r185_c29 bl[29] br[29] wl[185] vdd gnd cell_6t
Xbit_r186_c29 bl[29] br[29] wl[186] vdd gnd cell_6t
Xbit_r187_c29 bl[29] br[29] wl[187] vdd gnd cell_6t
Xbit_r188_c29 bl[29] br[29] wl[188] vdd gnd cell_6t
Xbit_r189_c29 bl[29] br[29] wl[189] vdd gnd cell_6t
Xbit_r190_c29 bl[29] br[29] wl[190] vdd gnd cell_6t
Xbit_r191_c29 bl[29] br[29] wl[191] vdd gnd cell_6t
Xbit_r192_c29 bl[29] br[29] wl[192] vdd gnd cell_6t
Xbit_r193_c29 bl[29] br[29] wl[193] vdd gnd cell_6t
Xbit_r194_c29 bl[29] br[29] wl[194] vdd gnd cell_6t
Xbit_r195_c29 bl[29] br[29] wl[195] vdd gnd cell_6t
Xbit_r196_c29 bl[29] br[29] wl[196] vdd gnd cell_6t
Xbit_r197_c29 bl[29] br[29] wl[197] vdd gnd cell_6t
Xbit_r198_c29 bl[29] br[29] wl[198] vdd gnd cell_6t
Xbit_r199_c29 bl[29] br[29] wl[199] vdd gnd cell_6t
Xbit_r200_c29 bl[29] br[29] wl[200] vdd gnd cell_6t
Xbit_r201_c29 bl[29] br[29] wl[201] vdd gnd cell_6t
Xbit_r202_c29 bl[29] br[29] wl[202] vdd gnd cell_6t
Xbit_r203_c29 bl[29] br[29] wl[203] vdd gnd cell_6t
Xbit_r204_c29 bl[29] br[29] wl[204] vdd gnd cell_6t
Xbit_r205_c29 bl[29] br[29] wl[205] vdd gnd cell_6t
Xbit_r206_c29 bl[29] br[29] wl[206] vdd gnd cell_6t
Xbit_r207_c29 bl[29] br[29] wl[207] vdd gnd cell_6t
Xbit_r208_c29 bl[29] br[29] wl[208] vdd gnd cell_6t
Xbit_r209_c29 bl[29] br[29] wl[209] vdd gnd cell_6t
Xbit_r210_c29 bl[29] br[29] wl[210] vdd gnd cell_6t
Xbit_r211_c29 bl[29] br[29] wl[211] vdd gnd cell_6t
Xbit_r212_c29 bl[29] br[29] wl[212] vdd gnd cell_6t
Xbit_r213_c29 bl[29] br[29] wl[213] vdd gnd cell_6t
Xbit_r214_c29 bl[29] br[29] wl[214] vdd gnd cell_6t
Xbit_r215_c29 bl[29] br[29] wl[215] vdd gnd cell_6t
Xbit_r216_c29 bl[29] br[29] wl[216] vdd gnd cell_6t
Xbit_r217_c29 bl[29] br[29] wl[217] vdd gnd cell_6t
Xbit_r218_c29 bl[29] br[29] wl[218] vdd gnd cell_6t
Xbit_r219_c29 bl[29] br[29] wl[219] vdd gnd cell_6t
Xbit_r220_c29 bl[29] br[29] wl[220] vdd gnd cell_6t
Xbit_r221_c29 bl[29] br[29] wl[221] vdd gnd cell_6t
Xbit_r222_c29 bl[29] br[29] wl[222] vdd gnd cell_6t
Xbit_r223_c29 bl[29] br[29] wl[223] vdd gnd cell_6t
Xbit_r224_c29 bl[29] br[29] wl[224] vdd gnd cell_6t
Xbit_r225_c29 bl[29] br[29] wl[225] vdd gnd cell_6t
Xbit_r226_c29 bl[29] br[29] wl[226] vdd gnd cell_6t
Xbit_r227_c29 bl[29] br[29] wl[227] vdd gnd cell_6t
Xbit_r228_c29 bl[29] br[29] wl[228] vdd gnd cell_6t
Xbit_r229_c29 bl[29] br[29] wl[229] vdd gnd cell_6t
Xbit_r230_c29 bl[29] br[29] wl[230] vdd gnd cell_6t
Xbit_r231_c29 bl[29] br[29] wl[231] vdd gnd cell_6t
Xbit_r232_c29 bl[29] br[29] wl[232] vdd gnd cell_6t
Xbit_r233_c29 bl[29] br[29] wl[233] vdd gnd cell_6t
Xbit_r234_c29 bl[29] br[29] wl[234] vdd gnd cell_6t
Xbit_r235_c29 bl[29] br[29] wl[235] vdd gnd cell_6t
Xbit_r236_c29 bl[29] br[29] wl[236] vdd gnd cell_6t
Xbit_r237_c29 bl[29] br[29] wl[237] vdd gnd cell_6t
Xbit_r238_c29 bl[29] br[29] wl[238] vdd gnd cell_6t
Xbit_r239_c29 bl[29] br[29] wl[239] vdd gnd cell_6t
Xbit_r240_c29 bl[29] br[29] wl[240] vdd gnd cell_6t
Xbit_r241_c29 bl[29] br[29] wl[241] vdd gnd cell_6t
Xbit_r242_c29 bl[29] br[29] wl[242] vdd gnd cell_6t
Xbit_r243_c29 bl[29] br[29] wl[243] vdd gnd cell_6t
Xbit_r244_c29 bl[29] br[29] wl[244] vdd gnd cell_6t
Xbit_r245_c29 bl[29] br[29] wl[245] vdd gnd cell_6t
Xbit_r246_c29 bl[29] br[29] wl[246] vdd gnd cell_6t
Xbit_r247_c29 bl[29] br[29] wl[247] vdd gnd cell_6t
Xbit_r248_c29 bl[29] br[29] wl[248] vdd gnd cell_6t
Xbit_r249_c29 bl[29] br[29] wl[249] vdd gnd cell_6t
Xbit_r250_c29 bl[29] br[29] wl[250] vdd gnd cell_6t
Xbit_r251_c29 bl[29] br[29] wl[251] vdd gnd cell_6t
Xbit_r252_c29 bl[29] br[29] wl[252] vdd gnd cell_6t
Xbit_r253_c29 bl[29] br[29] wl[253] vdd gnd cell_6t
Xbit_r254_c29 bl[29] br[29] wl[254] vdd gnd cell_6t
Xbit_r255_c29 bl[29] br[29] wl[255] vdd gnd cell_6t
Xbit_r0_c30 bl[30] br[30] wl[0] vdd gnd cell_6t
Xbit_r1_c30 bl[30] br[30] wl[1] vdd gnd cell_6t
Xbit_r2_c30 bl[30] br[30] wl[2] vdd gnd cell_6t
Xbit_r3_c30 bl[30] br[30] wl[3] vdd gnd cell_6t
Xbit_r4_c30 bl[30] br[30] wl[4] vdd gnd cell_6t
Xbit_r5_c30 bl[30] br[30] wl[5] vdd gnd cell_6t
Xbit_r6_c30 bl[30] br[30] wl[6] vdd gnd cell_6t
Xbit_r7_c30 bl[30] br[30] wl[7] vdd gnd cell_6t
Xbit_r8_c30 bl[30] br[30] wl[8] vdd gnd cell_6t
Xbit_r9_c30 bl[30] br[30] wl[9] vdd gnd cell_6t
Xbit_r10_c30 bl[30] br[30] wl[10] vdd gnd cell_6t
Xbit_r11_c30 bl[30] br[30] wl[11] vdd gnd cell_6t
Xbit_r12_c30 bl[30] br[30] wl[12] vdd gnd cell_6t
Xbit_r13_c30 bl[30] br[30] wl[13] vdd gnd cell_6t
Xbit_r14_c30 bl[30] br[30] wl[14] vdd gnd cell_6t
Xbit_r15_c30 bl[30] br[30] wl[15] vdd gnd cell_6t
Xbit_r16_c30 bl[30] br[30] wl[16] vdd gnd cell_6t
Xbit_r17_c30 bl[30] br[30] wl[17] vdd gnd cell_6t
Xbit_r18_c30 bl[30] br[30] wl[18] vdd gnd cell_6t
Xbit_r19_c30 bl[30] br[30] wl[19] vdd gnd cell_6t
Xbit_r20_c30 bl[30] br[30] wl[20] vdd gnd cell_6t
Xbit_r21_c30 bl[30] br[30] wl[21] vdd gnd cell_6t
Xbit_r22_c30 bl[30] br[30] wl[22] vdd gnd cell_6t
Xbit_r23_c30 bl[30] br[30] wl[23] vdd gnd cell_6t
Xbit_r24_c30 bl[30] br[30] wl[24] vdd gnd cell_6t
Xbit_r25_c30 bl[30] br[30] wl[25] vdd gnd cell_6t
Xbit_r26_c30 bl[30] br[30] wl[26] vdd gnd cell_6t
Xbit_r27_c30 bl[30] br[30] wl[27] vdd gnd cell_6t
Xbit_r28_c30 bl[30] br[30] wl[28] vdd gnd cell_6t
Xbit_r29_c30 bl[30] br[30] wl[29] vdd gnd cell_6t
Xbit_r30_c30 bl[30] br[30] wl[30] vdd gnd cell_6t
Xbit_r31_c30 bl[30] br[30] wl[31] vdd gnd cell_6t
Xbit_r32_c30 bl[30] br[30] wl[32] vdd gnd cell_6t
Xbit_r33_c30 bl[30] br[30] wl[33] vdd gnd cell_6t
Xbit_r34_c30 bl[30] br[30] wl[34] vdd gnd cell_6t
Xbit_r35_c30 bl[30] br[30] wl[35] vdd gnd cell_6t
Xbit_r36_c30 bl[30] br[30] wl[36] vdd gnd cell_6t
Xbit_r37_c30 bl[30] br[30] wl[37] vdd gnd cell_6t
Xbit_r38_c30 bl[30] br[30] wl[38] vdd gnd cell_6t
Xbit_r39_c30 bl[30] br[30] wl[39] vdd gnd cell_6t
Xbit_r40_c30 bl[30] br[30] wl[40] vdd gnd cell_6t
Xbit_r41_c30 bl[30] br[30] wl[41] vdd gnd cell_6t
Xbit_r42_c30 bl[30] br[30] wl[42] vdd gnd cell_6t
Xbit_r43_c30 bl[30] br[30] wl[43] vdd gnd cell_6t
Xbit_r44_c30 bl[30] br[30] wl[44] vdd gnd cell_6t
Xbit_r45_c30 bl[30] br[30] wl[45] vdd gnd cell_6t
Xbit_r46_c30 bl[30] br[30] wl[46] vdd gnd cell_6t
Xbit_r47_c30 bl[30] br[30] wl[47] vdd gnd cell_6t
Xbit_r48_c30 bl[30] br[30] wl[48] vdd gnd cell_6t
Xbit_r49_c30 bl[30] br[30] wl[49] vdd gnd cell_6t
Xbit_r50_c30 bl[30] br[30] wl[50] vdd gnd cell_6t
Xbit_r51_c30 bl[30] br[30] wl[51] vdd gnd cell_6t
Xbit_r52_c30 bl[30] br[30] wl[52] vdd gnd cell_6t
Xbit_r53_c30 bl[30] br[30] wl[53] vdd gnd cell_6t
Xbit_r54_c30 bl[30] br[30] wl[54] vdd gnd cell_6t
Xbit_r55_c30 bl[30] br[30] wl[55] vdd gnd cell_6t
Xbit_r56_c30 bl[30] br[30] wl[56] vdd gnd cell_6t
Xbit_r57_c30 bl[30] br[30] wl[57] vdd gnd cell_6t
Xbit_r58_c30 bl[30] br[30] wl[58] vdd gnd cell_6t
Xbit_r59_c30 bl[30] br[30] wl[59] vdd gnd cell_6t
Xbit_r60_c30 bl[30] br[30] wl[60] vdd gnd cell_6t
Xbit_r61_c30 bl[30] br[30] wl[61] vdd gnd cell_6t
Xbit_r62_c30 bl[30] br[30] wl[62] vdd gnd cell_6t
Xbit_r63_c30 bl[30] br[30] wl[63] vdd gnd cell_6t
Xbit_r64_c30 bl[30] br[30] wl[64] vdd gnd cell_6t
Xbit_r65_c30 bl[30] br[30] wl[65] vdd gnd cell_6t
Xbit_r66_c30 bl[30] br[30] wl[66] vdd gnd cell_6t
Xbit_r67_c30 bl[30] br[30] wl[67] vdd gnd cell_6t
Xbit_r68_c30 bl[30] br[30] wl[68] vdd gnd cell_6t
Xbit_r69_c30 bl[30] br[30] wl[69] vdd gnd cell_6t
Xbit_r70_c30 bl[30] br[30] wl[70] vdd gnd cell_6t
Xbit_r71_c30 bl[30] br[30] wl[71] vdd gnd cell_6t
Xbit_r72_c30 bl[30] br[30] wl[72] vdd gnd cell_6t
Xbit_r73_c30 bl[30] br[30] wl[73] vdd gnd cell_6t
Xbit_r74_c30 bl[30] br[30] wl[74] vdd gnd cell_6t
Xbit_r75_c30 bl[30] br[30] wl[75] vdd gnd cell_6t
Xbit_r76_c30 bl[30] br[30] wl[76] vdd gnd cell_6t
Xbit_r77_c30 bl[30] br[30] wl[77] vdd gnd cell_6t
Xbit_r78_c30 bl[30] br[30] wl[78] vdd gnd cell_6t
Xbit_r79_c30 bl[30] br[30] wl[79] vdd gnd cell_6t
Xbit_r80_c30 bl[30] br[30] wl[80] vdd gnd cell_6t
Xbit_r81_c30 bl[30] br[30] wl[81] vdd gnd cell_6t
Xbit_r82_c30 bl[30] br[30] wl[82] vdd gnd cell_6t
Xbit_r83_c30 bl[30] br[30] wl[83] vdd gnd cell_6t
Xbit_r84_c30 bl[30] br[30] wl[84] vdd gnd cell_6t
Xbit_r85_c30 bl[30] br[30] wl[85] vdd gnd cell_6t
Xbit_r86_c30 bl[30] br[30] wl[86] vdd gnd cell_6t
Xbit_r87_c30 bl[30] br[30] wl[87] vdd gnd cell_6t
Xbit_r88_c30 bl[30] br[30] wl[88] vdd gnd cell_6t
Xbit_r89_c30 bl[30] br[30] wl[89] vdd gnd cell_6t
Xbit_r90_c30 bl[30] br[30] wl[90] vdd gnd cell_6t
Xbit_r91_c30 bl[30] br[30] wl[91] vdd gnd cell_6t
Xbit_r92_c30 bl[30] br[30] wl[92] vdd gnd cell_6t
Xbit_r93_c30 bl[30] br[30] wl[93] vdd gnd cell_6t
Xbit_r94_c30 bl[30] br[30] wl[94] vdd gnd cell_6t
Xbit_r95_c30 bl[30] br[30] wl[95] vdd gnd cell_6t
Xbit_r96_c30 bl[30] br[30] wl[96] vdd gnd cell_6t
Xbit_r97_c30 bl[30] br[30] wl[97] vdd gnd cell_6t
Xbit_r98_c30 bl[30] br[30] wl[98] vdd gnd cell_6t
Xbit_r99_c30 bl[30] br[30] wl[99] vdd gnd cell_6t
Xbit_r100_c30 bl[30] br[30] wl[100] vdd gnd cell_6t
Xbit_r101_c30 bl[30] br[30] wl[101] vdd gnd cell_6t
Xbit_r102_c30 bl[30] br[30] wl[102] vdd gnd cell_6t
Xbit_r103_c30 bl[30] br[30] wl[103] vdd gnd cell_6t
Xbit_r104_c30 bl[30] br[30] wl[104] vdd gnd cell_6t
Xbit_r105_c30 bl[30] br[30] wl[105] vdd gnd cell_6t
Xbit_r106_c30 bl[30] br[30] wl[106] vdd gnd cell_6t
Xbit_r107_c30 bl[30] br[30] wl[107] vdd gnd cell_6t
Xbit_r108_c30 bl[30] br[30] wl[108] vdd gnd cell_6t
Xbit_r109_c30 bl[30] br[30] wl[109] vdd gnd cell_6t
Xbit_r110_c30 bl[30] br[30] wl[110] vdd gnd cell_6t
Xbit_r111_c30 bl[30] br[30] wl[111] vdd gnd cell_6t
Xbit_r112_c30 bl[30] br[30] wl[112] vdd gnd cell_6t
Xbit_r113_c30 bl[30] br[30] wl[113] vdd gnd cell_6t
Xbit_r114_c30 bl[30] br[30] wl[114] vdd gnd cell_6t
Xbit_r115_c30 bl[30] br[30] wl[115] vdd gnd cell_6t
Xbit_r116_c30 bl[30] br[30] wl[116] vdd gnd cell_6t
Xbit_r117_c30 bl[30] br[30] wl[117] vdd gnd cell_6t
Xbit_r118_c30 bl[30] br[30] wl[118] vdd gnd cell_6t
Xbit_r119_c30 bl[30] br[30] wl[119] vdd gnd cell_6t
Xbit_r120_c30 bl[30] br[30] wl[120] vdd gnd cell_6t
Xbit_r121_c30 bl[30] br[30] wl[121] vdd gnd cell_6t
Xbit_r122_c30 bl[30] br[30] wl[122] vdd gnd cell_6t
Xbit_r123_c30 bl[30] br[30] wl[123] vdd gnd cell_6t
Xbit_r124_c30 bl[30] br[30] wl[124] vdd gnd cell_6t
Xbit_r125_c30 bl[30] br[30] wl[125] vdd gnd cell_6t
Xbit_r126_c30 bl[30] br[30] wl[126] vdd gnd cell_6t
Xbit_r127_c30 bl[30] br[30] wl[127] vdd gnd cell_6t
Xbit_r128_c30 bl[30] br[30] wl[128] vdd gnd cell_6t
Xbit_r129_c30 bl[30] br[30] wl[129] vdd gnd cell_6t
Xbit_r130_c30 bl[30] br[30] wl[130] vdd gnd cell_6t
Xbit_r131_c30 bl[30] br[30] wl[131] vdd gnd cell_6t
Xbit_r132_c30 bl[30] br[30] wl[132] vdd gnd cell_6t
Xbit_r133_c30 bl[30] br[30] wl[133] vdd gnd cell_6t
Xbit_r134_c30 bl[30] br[30] wl[134] vdd gnd cell_6t
Xbit_r135_c30 bl[30] br[30] wl[135] vdd gnd cell_6t
Xbit_r136_c30 bl[30] br[30] wl[136] vdd gnd cell_6t
Xbit_r137_c30 bl[30] br[30] wl[137] vdd gnd cell_6t
Xbit_r138_c30 bl[30] br[30] wl[138] vdd gnd cell_6t
Xbit_r139_c30 bl[30] br[30] wl[139] vdd gnd cell_6t
Xbit_r140_c30 bl[30] br[30] wl[140] vdd gnd cell_6t
Xbit_r141_c30 bl[30] br[30] wl[141] vdd gnd cell_6t
Xbit_r142_c30 bl[30] br[30] wl[142] vdd gnd cell_6t
Xbit_r143_c30 bl[30] br[30] wl[143] vdd gnd cell_6t
Xbit_r144_c30 bl[30] br[30] wl[144] vdd gnd cell_6t
Xbit_r145_c30 bl[30] br[30] wl[145] vdd gnd cell_6t
Xbit_r146_c30 bl[30] br[30] wl[146] vdd gnd cell_6t
Xbit_r147_c30 bl[30] br[30] wl[147] vdd gnd cell_6t
Xbit_r148_c30 bl[30] br[30] wl[148] vdd gnd cell_6t
Xbit_r149_c30 bl[30] br[30] wl[149] vdd gnd cell_6t
Xbit_r150_c30 bl[30] br[30] wl[150] vdd gnd cell_6t
Xbit_r151_c30 bl[30] br[30] wl[151] vdd gnd cell_6t
Xbit_r152_c30 bl[30] br[30] wl[152] vdd gnd cell_6t
Xbit_r153_c30 bl[30] br[30] wl[153] vdd gnd cell_6t
Xbit_r154_c30 bl[30] br[30] wl[154] vdd gnd cell_6t
Xbit_r155_c30 bl[30] br[30] wl[155] vdd gnd cell_6t
Xbit_r156_c30 bl[30] br[30] wl[156] vdd gnd cell_6t
Xbit_r157_c30 bl[30] br[30] wl[157] vdd gnd cell_6t
Xbit_r158_c30 bl[30] br[30] wl[158] vdd gnd cell_6t
Xbit_r159_c30 bl[30] br[30] wl[159] vdd gnd cell_6t
Xbit_r160_c30 bl[30] br[30] wl[160] vdd gnd cell_6t
Xbit_r161_c30 bl[30] br[30] wl[161] vdd gnd cell_6t
Xbit_r162_c30 bl[30] br[30] wl[162] vdd gnd cell_6t
Xbit_r163_c30 bl[30] br[30] wl[163] vdd gnd cell_6t
Xbit_r164_c30 bl[30] br[30] wl[164] vdd gnd cell_6t
Xbit_r165_c30 bl[30] br[30] wl[165] vdd gnd cell_6t
Xbit_r166_c30 bl[30] br[30] wl[166] vdd gnd cell_6t
Xbit_r167_c30 bl[30] br[30] wl[167] vdd gnd cell_6t
Xbit_r168_c30 bl[30] br[30] wl[168] vdd gnd cell_6t
Xbit_r169_c30 bl[30] br[30] wl[169] vdd gnd cell_6t
Xbit_r170_c30 bl[30] br[30] wl[170] vdd gnd cell_6t
Xbit_r171_c30 bl[30] br[30] wl[171] vdd gnd cell_6t
Xbit_r172_c30 bl[30] br[30] wl[172] vdd gnd cell_6t
Xbit_r173_c30 bl[30] br[30] wl[173] vdd gnd cell_6t
Xbit_r174_c30 bl[30] br[30] wl[174] vdd gnd cell_6t
Xbit_r175_c30 bl[30] br[30] wl[175] vdd gnd cell_6t
Xbit_r176_c30 bl[30] br[30] wl[176] vdd gnd cell_6t
Xbit_r177_c30 bl[30] br[30] wl[177] vdd gnd cell_6t
Xbit_r178_c30 bl[30] br[30] wl[178] vdd gnd cell_6t
Xbit_r179_c30 bl[30] br[30] wl[179] vdd gnd cell_6t
Xbit_r180_c30 bl[30] br[30] wl[180] vdd gnd cell_6t
Xbit_r181_c30 bl[30] br[30] wl[181] vdd gnd cell_6t
Xbit_r182_c30 bl[30] br[30] wl[182] vdd gnd cell_6t
Xbit_r183_c30 bl[30] br[30] wl[183] vdd gnd cell_6t
Xbit_r184_c30 bl[30] br[30] wl[184] vdd gnd cell_6t
Xbit_r185_c30 bl[30] br[30] wl[185] vdd gnd cell_6t
Xbit_r186_c30 bl[30] br[30] wl[186] vdd gnd cell_6t
Xbit_r187_c30 bl[30] br[30] wl[187] vdd gnd cell_6t
Xbit_r188_c30 bl[30] br[30] wl[188] vdd gnd cell_6t
Xbit_r189_c30 bl[30] br[30] wl[189] vdd gnd cell_6t
Xbit_r190_c30 bl[30] br[30] wl[190] vdd gnd cell_6t
Xbit_r191_c30 bl[30] br[30] wl[191] vdd gnd cell_6t
Xbit_r192_c30 bl[30] br[30] wl[192] vdd gnd cell_6t
Xbit_r193_c30 bl[30] br[30] wl[193] vdd gnd cell_6t
Xbit_r194_c30 bl[30] br[30] wl[194] vdd gnd cell_6t
Xbit_r195_c30 bl[30] br[30] wl[195] vdd gnd cell_6t
Xbit_r196_c30 bl[30] br[30] wl[196] vdd gnd cell_6t
Xbit_r197_c30 bl[30] br[30] wl[197] vdd gnd cell_6t
Xbit_r198_c30 bl[30] br[30] wl[198] vdd gnd cell_6t
Xbit_r199_c30 bl[30] br[30] wl[199] vdd gnd cell_6t
Xbit_r200_c30 bl[30] br[30] wl[200] vdd gnd cell_6t
Xbit_r201_c30 bl[30] br[30] wl[201] vdd gnd cell_6t
Xbit_r202_c30 bl[30] br[30] wl[202] vdd gnd cell_6t
Xbit_r203_c30 bl[30] br[30] wl[203] vdd gnd cell_6t
Xbit_r204_c30 bl[30] br[30] wl[204] vdd gnd cell_6t
Xbit_r205_c30 bl[30] br[30] wl[205] vdd gnd cell_6t
Xbit_r206_c30 bl[30] br[30] wl[206] vdd gnd cell_6t
Xbit_r207_c30 bl[30] br[30] wl[207] vdd gnd cell_6t
Xbit_r208_c30 bl[30] br[30] wl[208] vdd gnd cell_6t
Xbit_r209_c30 bl[30] br[30] wl[209] vdd gnd cell_6t
Xbit_r210_c30 bl[30] br[30] wl[210] vdd gnd cell_6t
Xbit_r211_c30 bl[30] br[30] wl[211] vdd gnd cell_6t
Xbit_r212_c30 bl[30] br[30] wl[212] vdd gnd cell_6t
Xbit_r213_c30 bl[30] br[30] wl[213] vdd gnd cell_6t
Xbit_r214_c30 bl[30] br[30] wl[214] vdd gnd cell_6t
Xbit_r215_c30 bl[30] br[30] wl[215] vdd gnd cell_6t
Xbit_r216_c30 bl[30] br[30] wl[216] vdd gnd cell_6t
Xbit_r217_c30 bl[30] br[30] wl[217] vdd gnd cell_6t
Xbit_r218_c30 bl[30] br[30] wl[218] vdd gnd cell_6t
Xbit_r219_c30 bl[30] br[30] wl[219] vdd gnd cell_6t
Xbit_r220_c30 bl[30] br[30] wl[220] vdd gnd cell_6t
Xbit_r221_c30 bl[30] br[30] wl[221] vdd gnd cell_6t
Xbit_r222_c30 bl[30] br[30] wl[222] vdd gnd cell_6t
Xbit_r223_c30 bl[30] br[30] wl[223] vdd gnd cell_6t
Xbit_r224_c30 bl[30] br[30] wl[224] vdd gnd cell_6t
Xbit_r225_c30 bl[30] br[30] wl[225] vdd gnd cell_6t
Xbit_r226_c30 bl[30] br[30] wl[226] vdd gnd cell_6t
Xbit_r227_c30 bl[30] br[30] wl[227] vdd gnd cell_6t
Xbit_r228_c30 bl[30] br[30] wl[228] vdd gnd cell_6t
Xbit_r229_c30 bl[30] br[30] wl[229] vdd gnd cell_6t
Xbit_r230_c30 bl[30] br[30] wl[230] vdd gnd cell_6t
Xbit_r231_c30 bl[30] br[30] wl[231] vdd gnd cell_6t
Xbit_r232_c30 bl[30] br[30] wl[232] vdd gnd cell_6t
Xbit_r233_c30 bl[30] br[30] wl[233] vdd gnd cell_6t
Xbit_r234_c30 bl[30] br[30] wl[234] vdd gnd cell_6t
Xbit_r235_c30 bl[30] br[30] wl[235] vdd gnd cell_6t
Xbit_r236_c30 bl[30] br[30] wl[236] vdd gnd cell_6t
Xbit_r237_c30 bl[30] br[30] wl[237] vdd gnd cell_6t
Xbit_r238_c30 bl[30] br[30] wl[238] vdd gnd cell_6t
Xbit_r239_c30 bl[30] br[30] wl[239] vdd gnd cell_6t
Xbit_r240_c30 bl[30] br[30] wl[240] vdd gnd cell_6t
Xbit_r241_c30 bl[30] br[30] wl[241] vdd gnd cell_6t
Xbit_r242_c30 bl[30] br[30] wl[242] vdd gnd cell_6t
Xbit_r243_c30 bl[30] br[30] wl[243] vdd gnd cell_6t
Xbit_r244_c30 bl[30] br[30] wl[244] vdd gnd cell_6t
Xbit_r245_c30 bl[30] br[30] wl[245] vdd gnd cell_6t
Xbit_r246_c30 bl[30] br[30] wl[246] vdd gnd cell_6t
Xbit_r247_c30 bl[30] br[30] wl[247] vdd gnd cell_6t
Xbit_r248_c30 bl[30] br[30] wl[248] vdd gnd cell_6t
Xbit_r249_c30 bl[30] br[30] wl[249] vdd gnd cell_6t
Xbit_r250_c30 bl[30] br[30] wl[250] vdd gnd cell_6t
Xbit_r251_c30 bl[30] br[30] wl[251] vdd gnd cell_6t
Xbit_r252_c30 bl[30] br[30] wl[252] vdd gnd cell_6t
Xbit_r253_c30 bl[30] br[30] wl[253] vdd gnd cell_6t
Xbit_r254_c30 bl[30] br[30] wl[254] vdd gnd cell_6t
Xbit_r255_c30 bl[30] br[30] wl[255] vdd gnd cell_6t
Xbit_r0_c31 bl[31] br[31] wl[0] vdd gnd cell_6t
Xbit_r1_c31 bl[31] br[31] wl[1] vdd gnd cell_6t
Xbit_r2_c31 bl[31] br[31] wl[2] vdd gnd cell_6t
Xbit_r3_c31 bl[31] br[31] wl[3] vdd gnd cell_6t
Xbit_r4_c31 bl[31] br[31] wl[4] vdd gnd cell_6t
Xbit_r5_c31 bl[31] br[31] wl[5] vdd gnd cell_6t
Xbit_r6_c31 bl[31] br[31] wl[6] vdd gnd cell_6t
Xbit_r7_c31 bl[31] br[31] wl[7] vdd gnd cell_6t
Xbit_r8_c31 bl[31] br[31] wl[8] vdd gnd cell_6t
Xbit_r9_c31 bl[31] br[31] wl[9] vdd gnd cell_6t
Xbit_r10_c31 bl[31] br[31] wl[10] vdd gnd cell_6t
Xbit_r11_c31 bl[31] br[31] wl[11] vdd gnd cell_6t
Xbit_r12_c31 bl[31] br[31] wl[12] vdd gnd cell_6t
Xbit_r13_c31 bl[31] br[31] wl[13] vdd gnd cell_6t
Xbit_r14_c31 bl[31] br[31] wl[14] vdd gnd cell_6t
Xbit_r15_c31 bl[31] br[31] wl[15] vdd gnd cell_6t
Xbit_r16_c31 bl[31] br[31] wl[16] vdd gnd cell_6t
Xbit_r17_c31 bl[31] br[31] wl[17] vdd gnd cell_6t
Xbit_r18_c31 bl[31] br[31] wl[18] vdd gnd cell_6t
Xbit_r19_c31 bl[31] br[31] wl[19] vdd gnd cell_6t
Xbit_r20_c31 bl[31] br[31] wl[20] vdd gnd cell_6t
Xbit_r21_c31 bl[31] br[31] wl[21] vdd gnd cell_6t
Xbit_r22_c31 bl[31] br[31] wl[22] vdd gnd cell_6t
Xbit_r23_c31 bl[31] br[31] wl[23] vdd gnd cell_6t
Xbit_r24_c31 bl[31] br[31] wl[24] vdd gnd cell_6t
Xbit_r25_c31 bl[31] br[31] wl[25] vdd gnd cell_6t
Xbit_r26_c31 bl[31] br[31] wl[26] vdd gnd cell_6t
Xbit_r27_c31 bl[31] br[31] wl[27] vdd gnd cell_6t
Xbit_r28_c31 bl[31] br[31] wl[28] vdd gnd cell_6t
Xbit_r29_c31 bl[31] br[31] wl[29] vdd gnd cell_6t
Xbit_r30_c31 bl[31] br[31] wl[30] vdd gnd cell_6t
Xbit_r31_c31 bl[31] br[31] wl[31] vdd gnd cell_6t
Xbit_r32_c31 bl[31] br[31] wl[32] vdd gnd cell_6t
Xbit_r33_c31 bl[31] br[31] wl[33] vdd gnd cell_6t
Xbit_r34_c31 bl[31] br[31] wl[34] vdd gnd cell_6t
Xbit_r35_c31 bl[31] br[31] wl[35] vdd gnd cell_6t
Xbit_r36_c31 bl[31] br[31] wl[36] vdd gnd cell_6t
Xbit_r37_c31 bl[31] br[31] wl[37] vdd gnd cell_6t
Xbit_r38_c31 bl[31] br[31] wl[38] vdd gnd cell_6t
Xbit_r39_c31 bl[31] br[31] wl[39] vdd gnd cell_6t
Xbit_r40_c31 bl[31] br[31] wl[40] vdd gnd cell_6t
Xbit_r41_c31 bl[31] br[31] wl[41] vdd gnd cell_6t
Xbit_r42_c31 bl[31] br[31] wl[42] vdd gnd cell_6t
Xbit_r43_c31 bl[31] br[31] wl[43] vdd gnd cell_6t
Xbit_r44_c31 bl[31] br[31] wl[44] vdd gnd cell_6t
Xbit_r45_c31 bl[31] br[31] wl[45] vdd gnd cell_6t
Xbit_r46_c31 bl[31] br[31] wl[46] vdd gnd cell_6t
Xbit_r47_c31 bl[31] br[31] wl[47] vdd gnd cell_6t
Xbit_r48_c31 bl[31] br[31] wl[48] vdd gnd cell_6t
Xbit_r49_c31 bl[31] br[31] wl[49] vdd gnd cell_6t
Xbit_r50_c31 bl[31] br[31] wl[50] vdd gnd cell_6t
Xbit_r51_c31 bl[31] br[31] wl[51] vdd gnd cell_6t
Xbit_r52_c31 bl[31] br[31] wl[52] vdd gnd cell_6t
Xbit_r53_c31 bl[31] br[31] wl[53] vdd gnd cell_6t
Xbit_r54_c31 bl[31] br[31] wl[54] vdd gnd cell_6t
Xbit_r55_c31 bl[31] br[31] wl[55] vdd gnd cell_6t
Xbit_r56_c31 bl[31] br[31] wl[56] vdd gnd cell_6t
Xbit_r57_c31 bl[31] br[31] wl[57] vdd gnd cell_6t
Xbit_r58_c31 bl[31] br[31] wl[58] vdd gnd cell_6t
Xbit_r59_c31 bl[31] br[31] wl[59] vdd gnd cell_6t
Xbit_r60_c31 bl[31] br[31] wl[60] vdd gnd cell_6t
Xbit_r61_c31 bl[31] br[31] wl[61] vdd gnd cell_6t
Xbit_r62_c31 bl[31] br[31] wl[62] vdd gnd cell_6t
Xbit_r63_c31 bl[31] br[31] wl[63] vdd gnd cell_6t
Xbit_r64_c31 bl[31] br[31] wl[64] vdd gnd cell_6t
Xbit_r65_c31 bl[31] br[31] wl[65] vdd gnd cell_6t
Xbit_r66_c31 bl[31] br[31] wl[66] vdd gnd cell_6t
Xbit_r67_c31 bl[31] br[31] wl[67] vdd gnd cell_6t
Xbit_r68_c31 bl[31] br[31] wl[68] vdd gnd cell_6t
Xbit_r69_c31 bl[31] br[31] wl[69] vdd gnd cell_6t
Xbit_r70_c31 bl[31] br[31] wl[70] vdd gnd cell_6t
Xbit_r71_c31 bl[31] br[31] wl[71] vdd gnd cell_6t
Xbit_r72_c31 bl[31] br[31] wl[72] vdd gnd cell_6t
Xbit_r73_c31 bl[31] br[31] wl[73] vdd gnd cell_6t
Xbit_r74_c31 bl[31] br[31] wl[74] vdd gnd cell_6t
Xbit_r75_c31 bl[31] br[31] wl[75] vdd gnd cell_6t
Xbit_r76_c31 bl[31] br[31] wl[76] vdd gnd cell_6t
Xbit_r77_c31 bl[31] br[31] wl[77] vdd gnd cell_6t
Xbit_r78_c31 bl[31] br[31] wl[78] vdd gnd cell_6t
Xbit_r79_c31 bl[31] br[31] wl[79] vdd gnd cell_6t
Xbit_r80_c31 bl[31] br[31] wl[80] vdd gnd cell_6t
Xbit_r81_c31 bl[31] br[31] wl[81] vdd gnd cell_6t
Xbit_r82_c31 bl[31] br[31] wl[82] vdd gnd cell_6t
Xbit_r83_c31 bl[31] br[31] wl[83] vdd gnd cell_6t
Xbit_r84_c31 bl[31] br[31] wl[84] vdd gnd cell_6t
Xbit_r85_c31 bl[31] br[31] wl[85] vdd gnd cell_6t
Xbit_r86_c31 bl[31] br[31] wl[86] vdd gnd cell_6t
Xbit_r87_c31 bl[31] br[31] wl[87] vdd gnd cell_6t
Xbit_r88_c31 bl[31] br[31] wl[88] vdd gnd cell_6t
Xbit_r89_c31 bl[31] br[31] wl[89] vdd gnd cell_6t
Xbit_r90_c31 bl[31] br[31] wl[90] vdd gnd cell_6t
Xbit_r91_c31 bl[31] br[31] wl[91] vdd gnd cell_6t
Xbit_r92_c31 bl[31] br[31] wl[92] vdd gnd cell_6t
Xbit_r93_c31 bl[31] br[31] wl[93] vdd gnd cell_6t
Xbit_r94_c31 bl[31] br[31] wl[94] vdd gnd cell_6t
Xbit_r95_c31 bl[31] br[31] wl[95] vdd gnd cell_6t
Xbit_r96_c31 bl[31] br[31] wl[96] vdd gnd cell_6t
Xbit_r97_c31 bl[31] br[31] wl[97] vdd gnd cell_6t
Xbit_r98_c31 bl[31] br[31] wl[98] vdd gnd cell_6t
Xbit_r99_c31 bl[31] br[31] wl[99] vdd gnd cell_6t
Xbit_r100_c31 bl[31] br[31] wl[100] vdd gnd cell_6t
Xbit_r101_c31 bl[31] br[31] wl[101] vdd gnd cell_6t
Xbit_r102_c31 bl[31] br[31] wl[102] vdd gnd cell_6t
Xbit_r103_c31 bl[31] br[31] wl[103] vdd gnd cell_6t
Xbit_r104_c31 bl[31] br[31] wl[104] vdd gnd cell_6t
Xbit_r105_c31 bl[31] br[31] wl[105] vdd gnd cell_6t
Xbit_r106_c31 bl[31] br[31] wl[106] vdd gnd cell_6t
Xbit_r107_c31 bl[31] br[31] wl[107] vdd gnd cell_6t
Xbit_r108_c31 bl[31] br[31] wl[108] vdd gnd cell_6t
Xbit_r109_c31 bl[31] br[31] wl[109] vdd gnd cell_6t
Xbit_r110_c31 bl[31] br[31] wl[110] vdd gnd cell_6t
Xbit_r111_c31 bl[31] br[31] wl[111] vdd gnd cell_6t
Xbit_r112_c31 bl[31] br[31] wl[112] vdd gnd cell_6t
Xbit_r113_c31 bl[31] br[31] wl[113] vdd gnd cell_6t
Xbit_r114_c31 bl[31] br[31] wl[114] vdd gnd cell_6t
Xbit_r115_c31 bl[31] br[31] wl[115] vdd gnd cell_6t
Xbit_r116_c31 bl[31] br[31] wl[116] vdd gnd cell_6t
Xbit_r117_c31 bl[31] br[31] wl[117] vdd gnd cell_6t
Xbit_r118_c31 bl[31] br[31] wl[118] vdd gnd cell_6t
Xbit_r119_c31 bl[31] br[31] wl[119] vdd gnd cell_6t
Xbit_r120_c31 bl[31] br[31] wl[120] vdd gnd cell_6t
Xbit_r121_c31 bl[31] br[31] wl[121] vdd gnd cell_6t
Xbit_r122_c31 bl[31] br[31] wl[122] vdd gnd cell_6t
Xbit_r123_c31 bl[31] br[31] wl[123] vdd gnd cell_6t
Xbit_r124_c31 bl[31] br[31] wl[124] vdd gnd cell_6t
Xbit_r125_c31 bl[31] br[31] wl[125] vdd gnd cell_6t
Xbit_r126_c31 bl[31] br[31] wl[126] vdd gnd cell_6t
Xbit_r127_c31 bl[31] br[31] wl[127] vdd gnd cell_6t
Xbit_r128_c31 bl[31] br[31] wl[128] vdd gnd cell_6t
Xbit_r129_c31 bl[31] br[31] wl[129] vdd gnd cell_6t
Xbit_r130_c31 bl[31] br[31] wl[130] vdd gnd cell_6t
Xbit_r131_c31 bl[31] br[31] wl[131] vdd gnd cell_6t
Xbit_r132_c31 bl[31] br[31] wl[132] vdd gnd cell_6t
Xbit_r133_c31 bl[31] br[31] wl[133] vdd gnd cell_6t
Xbit_r134_c31 bl[31] br[31] wl[134] vdd gnd cell_6t
Xbit_r135_c31 bl[31] br[31] wl[135] vdd gnd cell_6t
Xbit_r136_c31 bl[31] br[31] wl[136] vdd gnd cell_6t
Xbit_r137_c31 bl[31] br[31] wl[137] vdd gnd cell_6t
Xbit_r138_c31 bl[31] br[31] wl[138] vdd gnd cell_6t
Xbit_r139_c31 bl[31] br[31] wl[139] vdd gnd cell_6t
Xbit_r140_c31 bl[31] br[31] wl[140] vdd gnd cell_6t
Xbit_r141_c31 bl[31] br[31] wl[141] vdd gnd cell_6t
Xbit_r142_c31 bl[31] br[31] wl[142] vdd gnd cell_6t
Xbit_r143_c31 bl[31] br[31] wl[143] vdd gnd cell_6t
Xbit_r144_c31 bl[31] br[31] wl[144] vdd gnd cell_6t
Xbit_r145_c31 bl[31] br[31] wl[145] vdd gnd cell_6t
Xbit_r146_c31 bl[31] br[31] wl[146] vdd gnd cell_6t
Xbit_r147_c31 bl[31] br[31] wl[147] vdd gnd cell_6t
Xbit_r148_c31 bl[31] br[31] wl[148] vdd gnd cell_6t
Xbit_r149_c31 bl[31] br[31] wl[149] vdd gnd cell_6t
Xbit_r150_c31 bl[31] br[31] wl[150] vdd gnd cell_6t
Xbit_r151_c31 bl[31] br[31] wl[151] vdd gnd cell_6t
Xbit_r152_c31 bl[31] br[31] wl[152] vdd gnd cell_6t
Xbit_r153_c31 bl[31] br[31] wl[153] vdd gnd cell_6t
Xbit_r154_c31 bl[31] br[31] wl[154] vdd gnd cell_6t
Xbit_r155_c31 bl[31] br[31] wl[155] vdd gnd cell_6t
Xbit_r156_c31 bl[31] br[31] wl[156] vdd gnd cell_6t
Xbit_r157_c31 bl[31] br[31] wl[157] vdd gnd cell_6t
Xbit_r158_c31 bl[31] br[31] wl[158] vdd gnd cell_6t
Xbit_r159_c31 bl[31] br[31] wl[159] vdd gnd cell_6t
Xbit_r160_c31 bl[31] br[31] wl[160] vdd gnd cell_6t
Xbit_r161_c31 bl[31] br[31] wl[161] vdd gnd cell_6t
Xbit_r162_c31 bl[31] br[31] wl[162] vdd gnd cell_6t
Xbit_r163_c31 bl[31] br[31] wl[163] vdd gnd cell_6t
Xbit_r164_c31 bl[31] br[31] wl[164] vdd gnd cell_6t
Xbit_r165_c31 bl[31] br[31] wl[165] vdd gnd cell_6t
Xbit_r166_c31 bl[31] br[31] wl[166] vdd gnd cell_6t
Xbit_r167_c31 bl[31] br[31] wl[167] vdd gnd cell_6t
Xbit_r168_c31 bl[31] br[31] wl[168] vdd gnd cell_6t
Xbit_r169_c31 bl[31] br[31] wl[169] vdd gnd cell_6t
Xbit_r170_c31 bl[31] br[31] wl[170] vdd gnd cell_6t
Xbit_r171_c31 bl[31] br[31] wl[171] vdd gnd cell_6t
Xbit_r172_c31 bl[31] br[31] wl[172] vdd gnd cell_6t
Xbit_r173_c31 bl[31] br[31] wl[173] vdd gnd cell_6t
Xbit_r174_c31 bl[31] br[31] wl[174] vdd gnd cell_6t
Xbit_r175_c31 bl[31] br[31] wl[175] vdd gnd cell_6t
Xbit_r176_c31 bl[31] br[31] wl[176] vdd gnd cell_6t
Xbit_r177_c31 bl[31] br[31] wl[177] vdd gnd cell_6t
Xbit_r178_c31 bl[31] br[31] wl[178] vdd gnd cell_6t
Xbit_r179_c31 bl[31] br[31] wl[179] vdd gnd cell_6t
Xbit_r180_c31 bl[31] br[31] wl[180] vdd gnd cell_6t
Xbit_r181_c31 bl[31] br[31] wl[181] vdd gnd cell_6t
Xbit_r182_c31 bl[31] br[31] wl[182] vdd gnd cell_6t
Xbit_r183_c31 bl[31] br[31] wl[183] vdd gnd cell_6t
Xbit_r184_c31 bl[31] br[31] wl[184] vdd gnd cell_6t
Xbit_r185_c31 bl[31] br[31] wl[185] vdd gnd cell_6t
Xbit_r186_c31 bl[31] br[31] wl[186] vdd gnd cell_6t
Xbit_r187_c31 bl[31] br[31] wl[187] vdd gnd cell_6t
Xbit_r188_c31 bl[31] br[31] wl[188] vdd gnd cell_6t
Xbit_r189_c31 bl[31] br[31] wl[189] vdd gnd cell_6t
Xbit_r190_c31 bl[31] br[31] wl[190] vdd gnd cell_6t
Xbit_r191_c31 bl[31] br[31] wl[191] vdd gnd cell_6t
Xbit_r192_c31 bl[31] br[31] wl[192] vdd gnd cell_6t
Xbit_r193_c31 bl[31] br[31] wl[193] vdd gnd cell_6t
Xbit_r194_c31 bl[31] br[31] wl[194] vdd gnd cell_6t
Xbit_r195_c31 bl[31] br[31] wl[195] vdd gnd cell_6t
Xbit_r196_c31 bl[31] br[31] wl[196] vdd gnd cell_6t
Xbit_r197_c31 bl[31] br[31] wl[197] vdd gnd cell_6t
Xbit_r198_c31 bl[31] br[31] wl[198] vdd gnd cell_6t
Xbit_r199_c31 bl[31] br[31] wl[199] vdd gnd cell_6t
Xbit_r200_c31 bl[31] br[31] wl[200] vdd gnd cell_6t
Xbit_r201_c31 bl[31] br[31] wl[201] vdd gnd cell_6t
Xbit_r202_c31 bl[31] br[31] wl[202] vdd gnd cell_6t
Xbit_r203_c31 bl[31] br[31] wl[203] vdd gnd cell_6t
Xbit_r204_c31 bl[31] br[31] wl[204] vdd gnd cell_6t
Xbit_r205_c31 bl[31] br[31] wl[205] vdd gnd cell_6t
Xbit_r206_c31 bl[31] br[31] wl[206] vdd gnd cell_6t
Xbit_r207_c31 bl[31] br[31] wl[207] vdd gnd cell_6t
Xbit_r208_c31 bl[31] br[31] wl[208] vdd gnd cell_6t
Xbit_r209_c31 bl[31] br[31] wl[209] vdd gnd cell_6t
Xbit_r210_c31 bl[31] br[31] wl[210] vdd gnd cell_6t
Xbit_r211_c31 bl[31] br[31] wl[211] vdd gnd cell_6t
Xbit_r212_c31 bl[31] br[31] wl[212] vdd gnd cell_6t
Xbit_r213_c31 bl[31] br[31] wl[213] vdd gnd cell_6t
Xbit_r214_c31 bl[31] br[31] wl[214] vdd gnd cell_6t
Xbit_r215_c31 bl[31] br[31] wl[215] vdd gnd cell_6t
Xbit_r216_c31 bl[31] br[31] wl[216] vdd gnd cell_6t
Xbit_r217_c31 bl[31] br[31] wl[217] vdd gnd cell_6t
Xbit_r218_c31 bl[31] br[31] wl[218] vdd gnd cell_6t
Xbit_r219_c31 bl[31] br[31] wl[219] vdd gnd cell_6t
Xbit_r220_c31 bl[31] br[31] wl[220] vdd gnd cell_6t
Xbit_r221_c31 bl[31] br[31] wl[221] vdd gnd cell_6t
Xbit_r222_c31 bl[31] br[31] wl[222] vdd gnd cell_6t
Xbit_r223_c31 bl[31] br[31] wl[223] vdd gnd cell_6t
Xbit_r224_c31 bl[31] br[31] wl[224] vdd gnd cell_6t
Xbit_r225_c31 bl[31] br[31] wl[225] vdd gnd cell_6t
Xbit_r226_c31 bl[31] br[31] wl[226] vdd gnd cell_6t
Xbit_r227_c31 bl[31] br[31] wl[227] vdd gnd cell_6t
Xbit_r228_c31 bl[31] br[31] wl[228] vdd gnd cell_6t
Xbit_r229_c31 bl[31] br[31] wl[229] vdd gnd cell_6t
Xbit_r230_c31 bl[31] br[31] wl[230] vdd gnd cell_6t
Xbit_r231_c31 bl[31] br[31] wl[231] vdd gnd cell_6t
Xbit_r232_c31 bl[31] br[31] wl[232] vdd gnd cell_6t
Xbit_r233_c31 bl[31] br[31] wl[233] vdd gnd cell_6t
Xbit_r234_c31 bl[31] br[31] wl[234] vdd gnd cell_6t
Xbit_r235_c31 bl[31] br[31] wl[235] vdd gnd cell_6t
Xbit_r236_c31 bl[31] br[31] wl[236] vdd gnd cell_6t
Xbit_r237_c31 bl[31] br[31] wl[237] vdd gnd cell_6t
Xbit_r238_c31 bl[31] br[31] wl[238] vdd gnd cell_6t
Xbit_r239_c31 bl[31] br[31] wl[239] vdd gnd cell_6t
Xbit_r240_c31 bl[31] br[31] wl[240] vdd gnd cell_6t
Xbit_r241_c31 bl[31] br[31] wl[241] vdd gnd cell_6t
Xbit_r242_c31 bl[31] br[31] wl[242] vdd gnd cell_6t
Xbit_r243_c31 bl[31] br[31] wl[243] vdd gnd cell_6t
Xbit_r244_c31 bl[31] br[31] wl[244] vdd gnd cell_6t
Xbit_r245_c31 bl[31] br[31] wl[245] vdd gnd cell_6t
Xbit_r246_c31 bl[31] br[31] wl[246] vdd gnd cell_6t
Xbit_r247_c31 bl[31] br[31] wl[247] vdd gnd cell_6t
Xbit_r248_c31 bl[31] br[31] wl[248] vdd gnd cell_6t
Xbit_r249_c31 bl[31] br[31] wl[249] vdd gnd cell_6t
Xbit_r250_c31 bl[31] br[31] wl[250] vdd gnd cell_6t
Xbit_r251_c31 bl[31] br[31] wl[251] vdd gnd cell_6t
Xbit_r252_c31 bl[31] br[31] wl[252] vdd gnd cell_6t
Xbit_r253_c31 bl[31] br[31] wl[253] vdd gnd cell_6t
Xbit_r254_c31 bl[31] br[31] wl[254] vdd gnd cell_6t
Xbit_r255_c31 bl[31] br[31] wl[255] vdd gnd cell_6t
Xbit_r0_c32 bl[32] br[32] wl[0] vdd gnd cell_6t
Xbit_r1_c32 bl[32] br[32] wl[1] vdd gnd cell_6t
Xbit_r2_c32 bl[32] br[32] wl[2] vdd gnd cell_6t
Xbit_r3_c32 bl[32] br[32] wl[3] vdd gnd cell_6t
Xbit_r4_c32 bl[32] br[32] wl[4] vdd gnd cell_6t
Xbit_r5_c32 bl[32] br[32] wl[5] vdd gnd cell_6t
Xbit_r6_c32 bl[32] br[32] wl[6] vdd gnd cell_6t
Xbit_r7_c32 bl[32] br[32] wl[7] vdd gnd cell_6t
Xbit_r8_c32 bl[32] br[32] wl[8] vdd gnd cell_6t
Xbit_r9_c32 bl[32] br[32] wl[9] vdd gnd cell_6t
Xbit_r10_c32 bl[32] br[32] wl[10] vdd gnd cell_6t
Xbit_r11_c32 bl[32] br[32] wl[11] vdd gnd cell_6t
Xbit_r12_c32 bl[32] br[32] wl[12] vdd gnd cell_6t
Xbit_r13_c32 bl[32] br[32] wl[13] vdd gnd cell_6t
Xbit_r14_c32 bl[32] br[32] wl[14] vdd gnd cell_6t
Xbit_r15_c32 bl[32] br[32] wl[15] vdd gnd cell_6t
Xbit_r16_c32 bl[32] br[32] wl[16] vdd gnd cell_6t
Xbit_r17_c32 bl[32] br[32] wl[17] vdd gnd cell_6t
Xbit_r18_c32 bl[32] br[32] wl[18] vdd gnd cell_6t
Xbit_r19_c32 bl[32] br[32] wl[19] vdd gnd cell_6t
Xbit_r20_c32 bl[32] br[32] wl[20] vdd gnd cell_6t
Xbit_r21_c32 bl[32] br[32] wl[21] vdd gnd cell_6t
Xbit_r22_c32 bl[32] br[32] wl[22] vdd gnd cell_6t
Xbit_r23_c32 bl[32] br[32] wl[23] vdd gnd cell_6t
Xbit_r24_c32 bl[32] br[32] wl[24] vdd gnd cell_6t
Xbit_r25_c32 bl[32] br[32] wl[25] vdd gnd cell_6t
Xbit_r26_c32 bl[32] br[32] wl[26] vdd gnd cell_6t
Xbit_r27_c32 bl[32] br[32] wl[27] vdd gnd cell_6t
Xbit_r28_c32 bl[32] br[32] wl[28] vdd gnd cell_6t
Xbit_r29_c32 bl[32] br[32] wl[29] vdd gnd cell_6t
Xbit_r30_c32 bl[32] br[32] wl[30] vdd gnd cell_6t
Xbit_r31_c32 bl[32] br[32] wl[31] vdd gnd cell_6t
Xbit_r32_c32 bl[32] br[32] wl[32] vdd gnd cell_6t
Xbit_r33_c32 bl[32] br[32] wl[33] vdd gnd cell_6t
Xbit_r34_c32 bl[32] br[32] wl[34] vdd gnd cell_6t
Xbit_r35_c32 bl[32] br[32] wl[35] vdd gnd cell_6t
Xbit_r36_c32 bl[32] br[32] wl[36] vdd gnd cell_6t
Xbit_r37_c32 bl[32] br[32] wl[37] vdd gnd cell_6t
Xbit_r38_c32 bl[32] br[32] wl[38] vdd gnd cell_6t
Xbit_r39_c32 bl[32] br[32] wl[39] vdd gnd cell_6t
Xbit_r40_c32 bl[32] br[32] wl[40] vdd gnd cell_6t
Xbit_r41_c32 bl[32] br[32] wl[41] vdd gnd cell_6t
Xbit_r42_c32 bl[32] br[32] wl[42] vdd gnd cell_6t
Xbit_r43_c32 bl[32] br[32] wl[43] vdd gnd cell_6t
Xbit_r44_c32 bl[32] br[32] wl[44] vdd gnd cell_6t
Xbit_r45_c32 bl[32] br[32] wl[45] vdd gnd cell_6t
Xbit_r46_c32 bl[32] br[32] wl[46] vdd gnd cell_6t
Xbit_r47_c32 bl[32] br[32] wl[47] vdd gnd cell_6t
Xbit_r48_c32 bl[32] br[32] wl[48] vdd gnd cell_6t
Xbit_r49_c32 bl[32] br[32] wl[49] vdd gnd cell_6t
Xbit_r50_c32 bl[32] br[32] wl[50] vdd gnd cell_6t
Xbit_r51_c32 bl[32] br[32] wl[51] vdd gnd cell_6t
Xbit_r52_c32 bl[32] br[32] wl[52] vdd gnd cell_6t
Xbit_r53_c32 bl[32] br[32] wl[53] vdd gnd cell_6t
Xbit_r54_c32 bl[32] br[32] wl[54] vdd gnd cell_6t
Xbit_r55_c32 bl[32] br[32] wl[55] vdd gnd cell_6t
Xbit_r56_c32 bl[32] br[32] wl[56] vdd gnd cell_6t
Xbit_r57_c32 bl[32] br[32] wl[57] vdd gnd cell_6t
Xbit_r58_c32 bl[32] br[32] wl[58] vdd gnd cell_6t
Xbit_r59_c32 bl[32] br[32] wl[59] vdd gnd cell_6t
Xbit_r60_c32 bl[32] br[32] wl[60] vdd gnd cell_6t
Xbit_r61_c32 bl[32] br[32] wl[61] vdd gnd cell_6t
Xbit_r62_c32 bl[32] br[32] wl[62] vdd gnd cell_6t
Xbit_r63_c32 bl[32] br[32] wl[63] vdd gnd cell_6t
Xbit_r64_c32 bl[32] br[32] wl[64] vdd gnd cell_6t
Xbit_r65_c32 bl[32] br[32] wl[65] vdd gnd cell_6t
Xbit_r66_c32 bl[32] br[32] wl[66] vdd gnd cell_6t
Xbit_r67_c32 bl[32] br[32] wl[67] vdd gnd cell_6t
Xbit_r68_c32 bl[32] br[32] wl[68] vdd gnd cell_6t
Xbit_r69_c32 bl[32] br[32] wl[69] vdd gnd cell_6t
Xbit_r70_c32 bl[32] br[32] wl[70] vdd gnd cell_6t
Xbit_r71_c32 bl[32] br[32] wl[71] vdd gnd cell_6t
Xbit_r72_c32 bl[32] br[32] wl[72] vdd gnd cell_6t
Xbit_r73_c32 bl[32] br[32] wl[73] vdd gnd cell_6t
Xbit_r74_c32 bl[32] br[32] wl[74] vdd gnd cell_6t
Xbit_r75_c32 bl[32] br[32] wl[75] vdd gnd cell_6t
Xbit_r76_c32 bl[32] br[32] wl[76] vdd gnd cell_6t
Xbit_r77_c32 bl[32] br[32] wl[77] vdd gnd cell_6t
Xbit_r78_c32 bl[32] br[32] wl[78] vdd gnd cell_6t
Xbit_r79_c32 bl[32] br[32] wl[79] vdd gnd cell_6t
Xbit_r80_c32 bl[32] br[32] wl[80] vdd gnd cell_6t
Xbit_r81_c32 bl[32] br[32] wl[81] vdd gnd cell_6t
Xbit_r82_c32 bl[32] br[32] wl[82] vdd gnd cell_6t
Xbit_r83_c32 bl[32] br[32] wl[83] vdd gnd cell_6t
Xbit_r84_c32 bl[32] br[32] wl[84] vdd gnd cell_6t
Xbit_r85_c32 bl[32] br[32] wl[85] vdd gnd cell_6t
Xbit_r86_c32 bl[32] br[32] wl[86] vdd gnd cell_6t
Xbit_r87_c32 bl[32] br[32] wl[87] vdd gnd cell_6t
Xbit_r88_c32 bl[32] br[32] wl[88] vdd gnd cell_6t
Xbit_r89_c32 bl[32] br[32] wl[89] vdd gnd cell_6t
Xbit_r90_c32 bl[32] br[32] wl[90] vdd gnd cell_6t
Xbit_r91_c32 bl[32] br[32] wl[91] vdd gnd cell_6t
Xbit_r92_c32 bl[32] br[32] wl[92] vdd gnd cell_6t
Xbit_r93_c32 bl[32] br[32] wl[93] vdd gnd cell_6t
Xbit_r94_c32 bl[32] br[32] wl[94] vdd gnd cell_6t
Xbit_r95_c32 bl[32] br[32] wl[95] vdd gnd cell_6t
Xbit_r96_c32 bl[32] br[32] wl[96] vdd gnd cell_6t
Xbit_r97_c32 bl[32] br[32] wl[97] vdd gnd cell_6t
Xbit_r98_c32 bl[32] br[32] wl[98] vdd gnd cell_6t
Xbit_r99_c32 bl[32] br[32] wl[99] vdd gnd cell_6t
Xbit_r100_c32 bl[32] br[32] wl[100] vdd gnd cell_6t
Xbit_r101_c32 bl[32] br[32] wl[101] vdd gnd cell_6t
Xbit_r102_c32 bl[32] br[32] wl[102] vdd gnd cell_6t
Xbit_r103_c32 bl[32] br[32] wl[103] vdd gnd cell_6t
Xbit_r104_c32 bl[32] br[32] wl[104] vdd gnd cell_6t
Xbit_r105_c32 bl[32] br[32] wl[105] vdd gnd cell_6t
Xbit_r106_c32 bl[32] br[32] wl[106] vdd gnd cell_6t
Xbit_r107_c32 bl[32] br[32] wl[107] vdd gnd cell_6t
Xbit_r108_c32 bl[32] br[32] wl[108] vdd gnd cell_6t
Xbit_r109_c32 bl[32] br[32] wl[109] vdd gnd cell_6t
Xbit_r110_c32 bl[32] br[32] wl[110] vdd gnd cell_6t
Xbit_r111_c32 bl[32] br[32] wl[111] vdd gnd cell_6t
Xbit_r112_c32 bl[32] br[32] wl[112] vdd gnd cell_6t
Xbit_r113_c32 bl[32] br[32] wl[113] vdd gnd cell_6t
Xbit_r114_c32 bl[32] br[32] wl[114] vdd gnd cell_6t
Xbit_r115_c32 bl[32] br[32] wl[115] vdd gnd cell_6t
Xbit_r116_c32 bl[32] br[32] wl[116] vdd gnd cell_6t
Xbit_r117_c32 bl[32] br[32] wl[117] vdd gnd cell_6t
Xbit_r118_c32 bl[32] br[32] wl[118] vdd gnd cell_6t
Xbit_r119_c32 bl[32] br[32] wl[119] vdd gnd cell_6t
Xbit_r120_c32 bl[32] br[32] wl[120] vdd gnd cell_6t
Xbit_r121_c32 bl[32] br[32] wl[121] vdd gnd cell_6t
Xbit_r122_c32 bl[32] br[32] wl[122] vdd gnd cell_6t
Xbit_r123_c32 bl[32] br[32] wl[123] vdd gnd cell_6t
Xbit_r124_c32 bl[32] br[32] wl[124] vdd gnd cell_6t
Xbit_r125_c32 bl[32] br[32] wl[125] vdd gnd cell_6t
Xbit_r126_c32 bl[32] br[32] wl[126] vdd gnd cell_6t
Xbit_r127_c32 bl[32] br[32] wl[127] vdd gnd cell_6t
Xbit_r128_c32 bl[32] br[32] wl[128] vdd gnd cell_6t
Xbit_r129_c32 bl[32] br[32] wl[129] vdd gnd cell_6t
Xbit_r130_c32 bl[32] br[32] wl[130] vdd gnd cell_6t
Xbit_r131_c32 bl[32] br[32] wl[131] vdd gnd cell_6t
Xbit_r132_c32 bl[32] br[32] wl[132] vdd gnd cell_6t
Xbit_r133_c32 bl[32] br[32] wl[133] vdd gnd cell_6t
Xbit_r134_c32 bl[32] br[32] wl[134] vdd gnd cell_6t
Xbit_r135_c32 bl[32] br[32] wl[135] vdd gnd cell_6t
Xbit_r136_c32 bl[32] br[32] wl[136] vdd gnd cell_6t
Xbit_r137_c32 bl[32] br[32] wl[137] vdd gnd cell_6t
Xbit_r138_c32 bl[32] br[32] wl[138] vdd gnd cell_6t
Xbit_r139_c32 bl[32] br[32] wl[139] vdd gnd cell_6t
Xbit_r140_c32 bl[32] br[32] wl[140] vdd gnd cell_6t
Xbit_r141_c32 bl[32] br[32] wl[141] vdd gnd cell_6t
Xbit_r142_c32 bl[32] br[32] wl[142] vdd gnd cell_6t
Xbit_r143_c32 bl[32] br[32] wl[143] vdd gnd cell_6t
Xbit_r144_c32 bl[32] br[32] wl[144] vdd gnd cell_6t
Xbit_r145_c32 bl[32] br[32] wl[145] vdd gnd cell_6t
Xbit_r146_c32 bl[32] br[32] wl[146] vdd gnd cell_6t
Xbit_r147_c32 bl[32] br[32] wl[147] vdd gnd cell_6t
Xbit_r148_c32 bl[32] br[32] wl[148] vdd gnd cell_6t
Xbit_r149_c32 bl[32] br[32] wl[149] vdd gnd cell_6t
Xbit_r150_c32 bl[32] br[32] wl[150] vdd gnd cell_6t
Xbit_r151_c32 bl[32] br[32] wl[151] vdd gnd cell_6t
Xbit_r152_c32 bl[32] br[32] wl[152] vdd gnd cell_6t
Xbit_r153_c32 bl[32] br[32] wl[153] vdd gnd cell_6t
Xbit_r154_c32 bl[32] br[32] wl[154] vdd gnd cell_6t
Xbit_r155_c32 bl[32] br[32] wl[155] vdd gnd cell_6t
Xbit_r156_c32 bl[32] br[32] wl[156] vdd gnd cell_6t
Xbit_r157_c32 bl[32] br[32] wl[157] vdd gnd cell_6t
Xbit_r158_c32 bl[32] br[32] wl[158] vdd gnd cell_6t
Xbit_r159_c32 bl[32] br[32] wl[159] vdd gnd cell_6t
Xbit_r160_c32 bl[32] br[32] wl[160] vdd gnd cell_6t
Xbit_r161_c32 bl[32] br[32] wl[161] vdd gnd cell_6t
Xbit_r162_c32 bl[32] br[32] wl[162] vdd gnd cell_6t
Xbit_r163_c32 bl[32] br[32] wl[163] vdd gnd cell_6t
Xbit_r164_c32 bl[32] br[32] wl[164] vdd gnd cell_6t
Xbit_r165_c32 bl[32] br[32] wl[165] vdd gnd cell_6t
Xbit_r166_c32 bl[32] br[32] wl[166] vdd gnd cell_6t
Xbit_r167_c32 bl[32] br[32] wl[167] vdd gnd cell_6t
Xbit_r168_c32 bl[32] br[32] wl[168] vdd gnd cell_6t
Xbit_r169_c32 bl[32] br[32] wl[169] vdd gnd cell_6t
Xbit_r170_c32 bl[32] br[32] wl[170] vdd gnd cell_6t
Xbit_r171_c32 bl[32] br[32] wl[171] vdd gnd cell_6t
Xbit_r172_c32 bl[32] br[32] wl[172] vdd gnd cell_6t
Xbit_r173_c32 bl[32] br[32] wl[173] vdd gnd cell_6t
Xbit_r174_c32 bl[32] br[32] wl[174] vdd gnd cell_6t
Xbit_r175_c32 bl[32] br[32] wl[175] vdd gnd cell_6t
Xbit_r176_c32 bl[32] br[32] wl[176] vdd gnd cell_6t
Xbit_r177_c32 bl[32] br[32] wl[177] vdd gnd cell_6t
Xbit_r178_c32 bl[32] br[32] wl[178] vdd gnd cell_6t
Xbit_r179_c32 bl[32] br[32] wl[179] vdd gnd cell_6t
Xbit_r180_c32 bl[32] br[32] wl[180] vdd gnd cell_6t
Xbit_r181_c32 bl[32] br[32] wl[181] vdd gnd cell_6t
Xbit_r182_c32 bl[32] br[32] wl[182] vdd gnd cell_6t
Xbit_r183_c32 bl[32] br[32] wl[183] vdd gnd cell_6t
Xbit_r184_c32 bl[32] br[32] wl[184] vdd gnd cell_6t
Xbit_r185_c32 bl[32] br[32] wl[185] vdd gnd cell_6t
Xbit_r186_c32 bl[32] br[32] wl[186] vdd gnd cell_6t
Xbit_r187_c32 bl[32] br[32] wl[187] vdd gnd cell_6t
Xbit_r188_c32 bl[32] br[32] wl[188] vdd gnd cell_6t
Xbit_r189_c32 bl[32] br[32] wl[189] vdd gnd cell_6t
Xbit_r190_c32 bl[32] br[32] wl[190] vdd gnd cell_6t
Xbit_r191_c32 bl[32] br[32] wl[191] vdd gnd cell_6t
Xbit_r192_c32 bl[32] br[32] wl[192] vdd gnd cell_6t
Xbit_r193_c32 bl[32] br[32] wl[193] vdd gnd cell_6t
Xbit_r194_c32 bl[32] br[32] wl[194] vdd gnd cell_6t
Xbit_r195_c32 bl[32] br[32] wl[195] vdd gnd cell_6t
Xbit_r196_c32 bl[32] br[32] wl[196] vdd gnd cell_6t
Xbit_r197_c32 bl[32] br[32] wl[197] vdd gnd cell_6t
Xbit_r198_c32 bl[32] br[32] wl[198] vdd gnd cell_6t
Xbit_r199_c32 bl[32] br[32] wl[199] vdd gnd cell_6t
Xbit_r200_c32 bl[32] br[32] wl[200] vdd gnd cell_6t
Xbit_r201_c32 bl[32] br[32] wl[201] vdd gnd cell_6t
Xbit_r202_c32 bl[32] br[32] wl[202] vdd gnd cell_6t
Xbit_r203_c32 bl[32] br[32] wl[203] vdd gnd cell_6t
Xbit_r204_c32 bl[32] br[32] wl[204] vdd gnd cell_6t
Xbit_r205_c32 bl[32] br[32] wl[205] vdd gnd cell_6t
Xbit_r206_c32 bl[32] br[32] wl[206] vdd gnd cell_6t
Xbit_r207_c32 bl[32] br[32] wl[207] vdd gnd cell_6t
Xbit_r208_c32 bl[32] br[32] wl[208] vdd gnd cell_6t
Xbit_r209_c32 bl[32] br[32] wl[209] vdd gnd cell_6t
Xbit_r210_c32 bl[32] br[32] wl[210] vdd gnd cell_6t
Xbit_r211_c32 bl[32] br[32] wl[211] vdd gnd cell_6t
Xbit_r212_c32 bl[32] br[32] wl[212] vdd gnd cell_6t
Xbit_r213_c32 bl[32] br[32] wl[213] vdd gnd cell_6t
Xbit_r214_c32 bl[32] br[32] wl[214] vdd gnd cell_6t
Xbit_r215_c32 bl[32] br[32] wl[215] vdd gnd cell_6t
Xbit_r216_c32 bl[32] br[32] wl[216] vdd gnd cell_6t
Xbit_r217_c32 bl[32] br[32] wl[217] vdd gnd cell_6t
Xbit_r218_c32 bl[32] br[32] wl[218] vdd gnd cell_6t
Xbit_r219_c32 bl[32] br[32] wl[219] vdd gnd cell_6t
Xbit_r220_c32 bl[32] br[32] wl[220] vdd gnd cell_6t
Xbit_r221_c32 bl[32] br[32] wl[221] vdd gnd cell_6t
Xbit_r222_c32 bl[32] br[32] wl[222] vdd gnd cell_6t
Xbit_r223_c32 bl[32] br[32] wl[223] vdd gnd cell_6t
Xbit_r224_c32 bl[32] br[32] wl[224] vdd gnd cell_6t
Xbit_r225_c32 bl[32] br[32] wl[225] vdd gnd cell_6t
Xbit_r226_c32 bl[32] br[32] wl[226] vdd gnd cell_6t
Xbit_r227_c32 bl[32] br[32] wl[227] vdd gnd cell_6t
Xbit_r228_c32 bl[32] br[32] wl[228] vdd gnd cell_6t
Xbit_r229_c32 bl[32] br[32] wl[229] vdd gnd cell_6t
Xbit_r230_c32 bl[32] br[32] wl[230] vdd gnd cell_6t
Xbit_r231_c32 bl[32] br[32] wl[231] vdd gnd cell_6t
Xbit_r232_c32 bl[32] br[32] wl[232] vdd gnd cell_6t
Xbit_r233_c32 bl[32] br[32] wl[233] vdd gnd cell_6t
Xbit_r234_c32 bl[32] br[32] wl[234] vdd gnd cell_6t
Xbit_r235_c32 bl[32] br[32] wl[235] vdd gnd cell_6t
Xbit_r236_c32 bl[32] br[32] wl[236] vdd gnd cell_6t
Xbit_r237_c32 bl[32] br[32] wl[237] vdd gnd cell_6t
Xbit_r238_c32 bl[32] br[32] wl[238] vdd gnd cell_6t
Xbit_r239_c32 bl[32] br[32] wl[239] vdd gnd cell_6t
Xbit_r240_c32 bl[32] br[32] wl[240] vdd gnd cell_6t
Xbit_r241_c32 bl[32] br[32] wl[241] vdd gnd cell_6t
Xbit_r242_c32 bl[32] br[32] wl[242] vdd gnd cell_6t
Xbit_r243_c32 bl[32] br[32] wl[243] vdd gnd cell_6t
Xbit_r244_c32 bl[32] br[32] wl[244] vdd gnd cell_6t
Xbit_r245_c32 bl[32] br[32] wl[245] vdd gnd cell_6t
Xbit_r246_c32 bl[32] br[32] wl[246] vdd gnd cell_6t
Xbit_r247_c32 bl[32] br[32] wl[247] vdd gnd cell_6t
Xbit_r248_c32 bl[32] br[32] wl[248] vdd gnd cell_6t
Xbit_r249_c32 bl[32] br[32] wl[249] vdd gnd cell_6t
Xbit_r250_c32 bl[32] br[32] wl[250] vdd gnd cell_6t
Xbit_r251_c32 bl[32] br[32] wl[251] vdd gnd cell_6t
Xbit_r252_c32 bl[32] br[32] wl[252] vdd gnd cell_6t
Xbit_r253_c32 bl[32] br[32] wl[253] vdd gnd cell_6t
Xbit_r254_c32 bl[32] br[32] wl[254] vdd gnd cell_6t
Xbit_r255_c32 bl[32] br[32] wl[255] vdd gnd cell_6t
Xbit_r0_c33 bl[33] br[33] wl[0] vdd gnd cell_6t
Xbit_r1_c33 bl[33] br[33] wl[1] vdd gnd cell_6t
Xbit_r2_c33 bl[33] br[33] wl[2] vdd gnd cell_6t
Xbit_r3_c33 bl[33] br[33] wl[3] vdd gnd cell_6t
Xbit_r4_c33 bl[33] br[33] wl[4] vdd gnd cell_6t
Xbit_r5_c33 bl[33] br[33] wl[5] vdd gnd cell_6t
Xbit_r6_c33 bl[33] br[33] wl[6] vdd gnd cell_6t
Xbit_r7_c33 bl[33] br[33] wl[7] vdd gnd cell_6t
Xbit_r8_c33 bl[33] br[33] wl[8] vdd gnd cell_6t
Xbit_r9_c33 bl[33] br[33] wl[9] vdd gnd cell_6t
Xbit_r10_c33 bl[33] br[33] wl[10] vdd gnd cell_6t
Xbit_r11_c33 bl[33] br[33] wl[11] vdd gnd cell_6t
Xbit_r12_c33 bl[33] br[33] wl[12] vdd gnd cell_6t
Xbit_r13_c33 bl[33] br[33] wl[13] vdd gnd cell_6t
Xbit_r14_c33 bl[33] br[33] wl[14] vdd gnd cell_6t
Xbit_r15_c33 bl[33] br[33] wl[15] vdd gnd cell_6t
Xbit_r16_c33 bl[33] br[33] wl[16] vdd gnd cell_6t
Xbit_r17_c33 bl[33] br[33] wl[17] vdd gnd cell_6t
Xbit_r18_c33 bl[33] br[33] wl[18] vdd gnd cell_6t
Xbit_r19_c33 bl[33] br[33] wl[19] vdd gnd cell_6t
Xbit_r20_c33 bl[33] br[33] wl[20] vdd gnd cell_6t
Xbit_r21_c33 bl[33] br[33] wl[21] vdd gnd cell_6t
Xbit_r22_c33 bl[33] br[33] wl[22] vdd gnd cell_6t
Xbit_r23_c33 bl[33] br[33] wl[23] vdd gnd cell_6t
Xbit_r24_c33 bl[33] br[33] wl[24] vdd gnd cell_6t
Xbit_r25_c33 bl[33] br[33] wl[25] vdd gnd cell_6t
Xbit_r26_c33 bl[33] br[33] wl[26] vdd gnd cell_6t
Xbit_r27_c33 bl[33] br[33] wl[27] vdd gnd cell_6t
Xbit_r28_c33 bl[33] br[33] wl[28] vdd gnd cell_6t
Xbit_r29_c33 bl[33] br[33] wl[29] vdd gnd cell_6t
Xbit_r30_c33 bl[33] br[33] wl[30] vdd gnd cell_6t
Xbit_r31_c33 bl[33] br[33] wl[31] vdd gnd cell_6t
Xbit_r32_c33 bl[33] br[33] wl[32] vdd gnd cell_6t
Xbit_r33_c33 bl[33] br[33] wl[33] vdd gnd cell_6t
Xbit_r34_c33 bl[33] br[33] wl[34] vdd gnd cell_6t
Xbit_r35_c33 bl[33] br[33] wl[35] vdd gnd cell_6t
Xbit_r36_c33 bl[33] br[33] wl[36] vdd gnd cell_6t
Xbit_r37_c33 bl[33] br[33] wl[37] vdd gnd cell_6t
Xbit_r38_c33 bl[33] br[33] wl[38] vdd gnd cell_6t
Xbit_r39_c33 bl[33] br[33] wl[39] vdd gnd cell_6t
Xbit_r40_c33 bl[33] br[33] wl[40] vdd gnd cell_6t
Xbit_r41_c33 bl[33] br[33] wl[41] vdd gnd cell_6t
Xbit_r42_c33 bl[33] br[33] wl[42] vdd gnd cell_6t
Xbit_r43_c33 bl[33] br[33] wl[43] vdd gnd cell_6t
Xbit_r44_c33 bl[33] br[33] wl[44] vdd gnd cell_6t
Xbit_r45_c33 bl[33] br[33] wl[45] vdd gnd cell_6t
Xbit_r46_c33 bl[33] br[33] wl[46] vdd gnd cell_6t
Xbit_r47_c33 bl[33] br[33] wl[47] vdd gnd cell_6t
Xbit_r48_c33 bl[33] br[33] wl[48] vdd gnd cell_6t
Xbit_r49_c33 bl[33] br[33] wl[49] vdd gnd cell_6t
Xbit_r50_c33 bl[33] br[33] wl[50] vdd gnd cell_6t
Xbit_r51_c33 bl[33] br[33] wl[51] vdd gnd cell_6t
Xbit_r52_c33 bl[33] br[33] wl[52] vdd gnd cell_6t
Xbit_r53_c33 bl[33] br[33] wl[53] vdd gnd cell_6t
Xbit_r54_c33 bl[33] br[33] wl[54] vdd gnd cell_6t
Xbit_r55_c33 bl[33] br[33] wl[55] vdd gnd cell_6t
Xbit_r56_c33 bl[33] br[33] wl[56] vdd gnd cell_6t
Xbit_r57_c33 bl[33] br[33] wl[57] vdd gnd cell_6t
Xbit_r58_c33 bl[33] br[33] wl[58] vdd gnd cell_6t
Xbit_r59_c33 bl[33] br[33] wl[59] vdd gnd cell_6t
Xbit_r60_c33 bl[33] br[33] wl[60] vdd gnd cell_6t
Xbit_r61_c33 bl[33] br[33] wl[61] vdd gnd cell_6t
Xbit_r62_c33 bl[33] br[33] wl[62] vdd gnd cell_6t
Xbit_r63_c33 bl[33] br[33] wl[63] vdd gnd cell_6t
Xbit_r64_c33 bl[33] br[33] wl[64] vdd gnd cell_6t
Xbit_r65_c33 bl[33] br[33] wl[65] vdd gnd cell_6t
Xbit_r66_c33 bl[33] br[33] wl[66] vdd gnd cell_6t
Xbit_r67_c33 bl[33] br[33] wl[67] vdd gnd cell_6t
Xbit_r68_c33 bl[33] br[33] wl[68] vdd gnd cell_6t
Xbit_r69_c33 bl[33] br[33] wl[69] vdd gnd cell_6t
Xbit_r70_c33 bl[33] br[33] wl[70] vdd gnd cell_6t
Xbit_r71_c33 bl[33] br[33] wl[71] vdd gnd cell_6t
Xbit_r72_c33 bl[33] br[33] wl[72] vdd gnd cell_6t
Xbit_r73_c33 bl[33] br[33] wl[73] vdd gnd cell_6t
Xbit_r74_c33 bl[33] br[33] wl[74] vdd gnd cell_6t
Xbit_r75_c33 bl[33] br[33] wl[75] vdd gnd cell_6t
Xbit_r76_c33 bl[33] br[33] wl[76] vdd gnd cell_6t
Xbit_r77_c33 bl[33] br[33] wl[77] vdd gnd cell_6t
Xbit_r78_c33 bl[33] br[33] wl[78] vdd gnd cell_6t
Xbit_r79_c33 bl[33] br[33] wl[79] vdd gnd cell_6t
Xbit_r80_c33 bl[33] br[33] wl[80] vdd gnd cell_6t
Xbit_r81_c33 bl[33] br[33] wl[81] vdd gnd cell_6t
Xbit_r82_c33 bl[33] br[33] wl[82] vdd gnd cell_6t
Xbit_r83_c33 bl[33] br[33] wl[83] vdd gnd cell_6t
Xbit_r84_c33 bl[33] br[33] wl[84] vdd gnd cell_6t
Xbit_r85_c33 bl[33] br[33] wl[85] vdd gnd cell_6t
Xbit_r86_c33 bl[33] br[33] wl[86] vdd gnd cell_6t
Xbit_r87_c33 bl[33] br[33] wl[87] vdd gnd cell_6t
Xbit_r88_c33 bl[33] br[33] wl[88] vdd gnd cell_6t
Xbit_r89_c33 bl[33] br[33] wl[89] vdd gnd cell_6t
Xbit_r90_c33 bl[33] br[33] wl[90] vdd gnd cell_6t
Xbit_r91_c33 bl[33] br[33] wl[91] vdd gnd cell_6t
Xbit_r92_c33 bl[33] br[33] wl[92] vdd gnd cell_6t
Xbit_r93_c33 bl[33] br[33] wl[93] vdd gnd cell_6t
Xbit_r94_c33 bl[33] br[33] wl[94] vdd gnd cell_6t
Xbit_r95_c33 bl[33] br[33] wl[95] vdd gnd cell_6t
Xbit_r96_c33 bl[33] br[33] wl[96] vdd gnd cell_6t
Xbit_r97_c33 bl[33] br[33] wl[97] vdd gnd cell_6t
Xbit_r98_c33 bl[33] br[33] wl[98] vdd gnd cell_6t
Xbit_r99_c33 bl[33] br[33] wl[99] vdd gnd cell_6t
Xbit_r100_c33 bl[33] br[33] wl[100] vdd gnd cell_6t
Xbit_r101_c33 bl[33] br[33] wl[101] vdd gnd cell_6t
Xbit_r102_c33 bl[33] br[33] wl[102] vdd gnd cell_6t
Xbit_r103_c33 bl[33] br[33] wl[103] vdd gnd cell_6t
Xbit_r104_c33 bl[33] br[33] wl[104] vdd gnd cell_6t
Xbit_r105_c33 bl[33] br[33] wl[105] vdd gnd cell_6t
Xbit_r106_c33 bl[33] br[33] wl[106] vdd gnd cell_6t
Xbit_r107_c33 bl[33] br[33] wl[107] vdd gnd cell_6t
Xbit_r108_c33 bl[33] br[33] wl[108] vdd gnd cell_6t
Xbit_r109_c33 bl[33] br[33] wl[109] vdd gnd cell_6t
Xbit_r110_c33 bl[33] br[33] wl[110] vdd gnd cell_6t
Xbit_r111_c33 bl[33] br[33] wl[111] vdd gnd cell_6t
Xbit_r112_c33 bl[33] br[33] wl[112] vdd gnd cell_6t
Xbit_r113_c33 bl[33] br[33] wl[113] vdd gnd cell_6t
Xbit_r114_c33 bl[33] br[33] wl[114] vdd gnd cell_6t
Xbit_r115_c33 bl[33] br[33] wl[115] vdd gnd cell_6t
Xbit_r116_c33 bl[33] br[33] wl[116] vdd gnd cell_6t
Xbit_r117_c33 bl[33] br[33] wl[117] vdd gnd cell_6t
Xbit_r118_c33 bl[33] br[33] wl[118] vdd gnd cell_6t
Xbit_r119_c33 bl[33] br[33] wl[119] vdd gnd cell_6t
Xbit_r120_c33 bl[33] br[33] wl[120] vdd gnd cell_6t
Xbit_r121_c33 bl[33] br[33] wl[121] vdd gnd cell_6t
Xbit_r122_c33 bl[33] br[33] wl[122] vdd gnd cell_6t
Xbit_r123_c33 bl[33] br[33] wl[123] vdd gnd cell_6t
Xbit_r124_c33 bl[33] br[33] wl[124] vdd gnd cell_6t
Xbit_r125_c33 bl[33] br[33] wl[125] vdd gnd cell_6t
Xbit_r126_c33 bl[33] br[33] wl[126] vdd gnd cell_6t
Xbit_r127_c33 bl[33] br[33] wl[127] vdd gnd cell_6t
Xbit_r128_c33 bl[33] br[33] wl[128] vdd gnd cell_6t
Xbit_r129_c33 bl[33] br[33] wl[129] vdd gnd cell_6t
Xbit_r130_c33 bl[33] br[33] wl[130] vdd gnd cell_6t
Xbit_r131_c33 bl[33] br[33] wl[131] vdd gnd cell_6t
Xbit_r132_c33 bl[33] br[33] wl[132] vdd gnd cell_6t
Xbit_r133_c33 bl[33] br[33] wl[133] vdd gnd cell_6t
Xbit_r134_c33 bl[33] br[33] wl[134] vdd gnd cell_6t
Xbit_r135_c33 bl[33] br[33] wl[135] vdd gnd cell_6t
Xbit_r136_c33 bl[33] br[33] wl[136] vdd gnd cell_6t
Xbit_r137_c33 bl[33] br[33] wl[137] vdd gnd cell_6t
Xbit_r138_c33 bl[33] br[33] wl[138] vdd gnd cell_6t
Xbit_r139_c33 bl[33] br[33] wl[139] vdd gnd cell_6t
Xbit_r140_c33 bl[33] br[33] wl[140] vdd gnd cell_6t
Xbit_r141_c33 bl[33] br[33] wl[141] vdd gnd cell_6t
Xbit_r142_c33 bl[33] br[33] wl[142] vdd gnd cell_6t
Xbit_r143_c33 bl[33] br[33] wl[143] vdd gnd cell_6t
Xbit_r144_c33 bl[33] br[33] wl[144] vdd gnd cell_6t
Xbit_r145_c33 bl[33] br[33] wl[145] vdd gnd cell_6t
Xbit_r146_c33 bl[33] br[33] wl[146] vdd gnd cell_6t
Xbit_r147_c33 bl[33] br[33] wl[147] vdd gnd cell_6t
Xbit_r148_c33 bl[33] br[33] wl[148] vdd gnd cell_6t
Xbit_r149_c33 bl[33] br[33] wl[149] vdd gnd cell_6t
Xbit_r150_c33 bl[33] br[33] wl[150] vdd gnd cell_6t
Xbit_r151_c33 bl[33] br[33] wl[151] vdd gnd cell_6t
Xbit_r152_c33 bl[33] br[33] wl[152] vdd gnd cell_6t
Xbit_r153_c33 bl[33] br[33] wl[153] vdd gnd cell_6t
Xbit_r154_c33 bl[33] br[33] wl[154] vdd gnd cell_6t
Xbit_r155_c33 bl[33] br[33] wl[155] vdd gnd cell_6t
Xbit_r156_c33 bl[33] br[33] wl[156] vdd gnd cell_6t
Xbit_r157_c33 bl[33] br[33] wl[157] vdd gnd cell_6t
Xbit_r158_c33 bl[33] br[33] wl[158] vdd gnd cell_6t
Xbit_r159_c33 bl[33] br[33] wl[159] vdd gnd cell_6t
Xbit_r160_c33 bl[33] br[33] wl[160] vdd gnd cell_6t
Xbit_r161_c33 bl[33] br[33] wl[161] vdd gnd cell_6t
Xbit_r162_c33 bl[33] br[33] wl[162] vdd gnd cell_6t
Xbit_r163_c33 bl[33] br[33] wl[163] vdd gnd cell_6t
Xbit_r164_c33 bl[33] br[33] wl[164] vdd gnd cell_6t
Xbit_r165_c33 bl[33] br[33] wl[165] vdd gnd cell_6t
Xbit_r166_c33 bl[33] br[33] wl[166] vdd gnd cell_6t
Xbit_r167_c33 bl[33] br[33] wl[167] vdd gnd cell_6t
Xbit_r168_c33 bl[33] br[33] wl[168] vdd gnd cell_6t
Xbit_r169_c33 bl[33] br[33] wl[169] vdd gnd cell_6t
Xbit_r170_c33 bl[33] br[33] wl[170] vdd gnd cell_6t
Xbit_r171_c33 bl[33] br[33] wl[171] vdd gnd cell_6t
Xbit_r172_c33 bl[33] br[33] wl[172] vdd gnd cell_6t
Xbit_r173_c33 bl[33] br[33] wl[173] vdd gnd cell_6t
Xbit_r174_c33 bl[33] br[33] wl[174] vdd gnd cell_6t
Xbit_r175_c33 bl[33] br[33] wl[175] vdd gnd cell_6t
Xbit_r176_c33 bl[33] br[33] wl[176] vdd gnd cell_6t
Xbit_r177_c33 bl[33] br[33] wl[177] vdd gnd cell_6t
Xbit_r178_c33 bl[33] br[33] wl[178] vdd gnd cell_6t
Xbit_r179_c33 bl[33] br[33] wl[179] vdd gnd cell_6t
Xbit_r180_c33 bl[33] br[33] wl[180] vdd gnd cell_6t
Xbit_r181_c33 bl[33] br[33] wl[181] vdd gnd cell_6t
Xbit_r182_c33 bl[33] br[33] wl[182] vdd gnd cell_6t
Xbit_r183_c33 bl[33] br[33] wl[183] vdd gnd cell_6t
Xbit_r184_c33 bl[33] br[33] wl[184] vdd gnd cell_6t
Xbit_r185_c33 bl[33] br[33] wl[185] vdd gnd cell_6t
Xbit_r186_c33 bl[33] br[33] wl[186] vdd gnd cell_6t
Xbit_r187_c33 bl[33] br[33] wl[187] vdd gnd cell_6t
Xbit_r188_c33 bl[33] br[33] wl[188] vdd gnd cell_6t
Xbit_r189_c33 bl[33] br[33] wl[189] vdd gnd cell_6t
Xbit_r190_c33 bl[33] br[33] wl[190] vdd gnd cell_6t
Xbit_r191_c33 bl[33] br[33] wl[191] vdd gnd cell_6t
Xbit_r192_c33 bl[33] br[33] wl[192] vdd gnd cell_6t
Xbit_r193_c33 bl[33] br[33] wl[193] vdd gnd cell_6t
Xbit_r194_c33 bl[33] br[33] wl[194] vdd gnd cell_6t
Xbit_r195_c33 bl[33] br[33] wl[195] vdd gnd cell_6t
Xbit_r196_c33 bl[33] br[33] wl[196] vdd gnd cell_6t
Xbit_r197_c33 bl[33] br[33] wl[197] vdd gnd cell_6t
Xbit_r198_c33 bl[33] br[33] wl[198] vdd gnd cell_6t
Xbit_r199_c33 bl[33] br[33] wl[199] vdd gnd cell_6t
Xbit_r200_c33 bl[33] br[33] wl[200] vdd gnd cell_6t
Xbit_r201_c33 bl[33] br[33] wl[201] vdd gnd cell_6t
Xbit_r202_c33 bl[33] br[33] wl[202] vdd gnd cell_6t
Xbit_r203_c33 bl[33] br[33] wl[203] vdd gnd cell_6t
Xbit_r204_c33 bl[33] br[33] wl[204] vdd gnd cell_6t
Xbit_r205_c33 bl[33] br[33] wl[205] vdd gnd cell_6t
Xbit_r206_c33 bl[33] br[33] wl[206] vdd gnd cell_6t
Xbit_r207_c33 bl[33] br[33] wl[207] vdd gnd cell_6t
Xbit_r208_c33 bl[33] br[33] wl[208] vdd gnd cell_6t
Xbit_r209_c33 bl[33] br[33] wl[209] vdd gnd cell_6t
Xbit_r210_c33 bl[33] br[33] wl[210] vdd gnd cell_6t
Xbit_r211_c33 bl[33] br[33] wl[211] vdd gnd cell_6t
Xbit_r212_c33 bl[33] br[33] wl[212] vdd gnd cell_6t
Xbit_r213_c33 bl[33] br[33] wl[213] vdd gnd cell_6t
Xbit_r214_c33 bl[33] br[33] wl[214] vdd gnd cell_6t
Xbit_r215_c33 bl[33] br[33] wl[215] vdd gnd cell_6t
Xbit_r216_c33 bl[33] br[33] wl[216] vdd gnd cell_6t
Xbit_r217_c33 bl[33] br[33] wl[217] vdd gnd cell_6t
Xbit_r218_c33 bl[33] br[33] wl[218] vdd gnd cell_6t
Xbit_r219_c33 bl[33] br[33] wl[219] vdd gnd cell_6t
Xbit_r220_c33 bl[33] br[33] wl[220] vdd gnd cell_6t
Xbit_r221_c33 bl[33] br[33] wl[221] vdd gnd cell_6t
Xbit_r222_c33 bl[33] br[33] wl[222] vdd gnd cell_6t
Xbit_r223_c33 bl[33] br[33] wl[223] vdd gnd cell_6t
Xbit_r224_c33 bl[33] br[33] wl[224] vdd gnd cell_6t
Xbit_r225_c33 bl[33] br[33] wl[225] vdd gnd cell_6t
Xbit_r226_c33 bl[33] br[33] wl[226] vdd gnd cell_6t
Xbit_r227_c33 bl[33] br[33] wl[227] vdd gnd cell_6t
Xbit_r228_c33 bl[33] br[33] wl[228] vdd gnd cell_6t
Xbit_r229_c33 bl[33] br[33] wl[229] vdd gnd cell_6t
Xbit_r230_c33 bl[33] br[33] wl[230] vdd gnd cell_6t
Xbit_r231_c33 bl[33] br[33] wl[231] vdd gnd cell_6t
Xbit_r232_c33 bl[33] br[33] wl[232] vdd gnd cell_6t
Xbit_r233_c33 bl[33] br[33] wl[233] vdd gnd cell_6t
Xbit_r234_c33 bl[33] br[33] wl[234] vdd gnd cell_6t
Xbit_r235_c33 bl[33] br[33] wl[235] vdd gnd cell_6t
Xbit_r236_c33 bl[33] br[33] wl[236] vdd gnd cell_6t
Xbit_r237_c33 bl[33] br[33] wl[237] vdd gnd cell_6t
Xbit_r238_c33 bl[33] br[33] wl[238] vdd gnd cell_6t
Xbit_r239_c33 bl[33] br[33] wl[239] vdd gnd cell_6t
Xbit_r240_c33 bl[33] br[33] wl[240] vdd gnd cell_6t
Xbit_r241_c33 bl[33] br[33] wl[241] vdd gnd cell_6t
Xbit_r242_c33 bl[33] br[33] wl[242] vdd gnd cell_6t
Xbit_r243_c33 bl[33] br[33] wl[243] vdd gnd cell_6t
Xbit_r244_c33 bl[33] br[33] wl[244] vdd gnd cell_6t
Xbit_r245_c33 bl[33] br[33] wl[245] vdd gnd cell_6t
Xbit_r246_c33 bl[33] br[33] wl[246] vdd gnd cell_6t
Xbit_r247_c33 bl[33] br[33] wl[247] vdd gnd cell_6t
Xbit_r248_c33 bl[33] br[33] wl[248] vdd gnd cell_6t
Xbit_r249_c33 bl[33] br[33] wl[249] vdd gnd cell_6t
Xbit_r250_c33 bl[33] br[33] wl[250] vdd gnd cell_6t
Xbit_r251_c33 bl[33] br[33] wl[251] vdd gnd cell_6t
Xbit_r252_c33 bl[33] br[33] wl[252] vdd gnd cell_6t
Xbit_r253_c33 bl[33] br[33] wl[253] vdd gnd cell_6t
Xbit_r254_c33 bl[33] br[33] wl[254] vdd gnd cell_6t
Xbit_r255_c33 bl[33] br[33] wl[255] vdd gnd cell_6t
Xbit_r0_c34 bl[34] br[34] wl[0] vdd gnd cell_6t
Xbit_r1_c34 bl[34] br[34] wl[1] vdd gnd cell_6t
Xbit_r2_c34 bl[34] br[34] wl[2] vdd gnd cell_6t
Xbit_r3_c34 bl[34] br[34] wl[3] vdd gnd cell_6t
Xbit_r4_c34 bl[34] br[34] wl[4] vdd gnd cell_6t
Xbit_r5_c34 bl[34] br[34] wl[5] vdd gnd cell_6t
Xbit_r6_c34 bl[34] br[34] wl[6] vdd gnd cell_6t
Xbit_r7_c34 bl[34] br[34] wl[7] vdd gnd cell_6t
Xbit_r8_c34 bl[34] br[34] wl[8] vdd gnd cell_6t
Xbit_r9_c34 bl[34] br[34] wl[9] vdd gnd cell_6t
Xbit_r10_c34 bl[34] br[34] wl[10] vdd gnd cell_6t
Xbit_r11_c34 bl[34] br[34] wl[11] vdd gnd cell_6t
Xbit_r12_c34 bl[34] br[34] wl[12] vdd gnd cell_6t
Xbit_r13_c34 bl[34] br[34] wl[13] vdd gnd cell_6t
Xbit_r14_c34 bl[34] br[34] wl[14] vdd gnd cell_6t
Xbit_r15_c34 bl[34] br[34] wl[15] vdd gnd cell_6t
Xbit_r16_c34 bl[34] br[34] wl[16] vdd gnd cell_6t
Xbit_r17_c34 bl[34] br[34] wl[17] vdd gnd cell_6t
Xbit_r18_c34 bl[34] br[34] wl[18] vdd gnd cell_6t
Xbit_r19_c34 bl[34] br[34] wl[19] vdd gnd cell_6t
Xbit_r20_c34 bl[34] br[34] wl[20] vdd gnd cell_6t
Xbit_r21_c34 bl[34] br[34] wl[21] vdd gnd cell_6t
Xbit_r22_c34 bl[34] br[34] wl[22] vdd gnd cell_6t
Xbit_r23_c34 bl[34] br[34] wl[23] vdd gnd cell_6t
Xbit_r24_c34 bl[34] br[34] wl[24] vdd gnd cell_6t
Xbit_r25_c34 bl[34] br[34] wl[25] vdd gnd cell_6t
Xbit_r26_c34 bl[34] br[34] wl[26] vdd gnd cell_6t
Xbit_r27_c34 bl[34] br[34] wl[27] vdd gnd cell_6t
Xbit_r28_c34 bl[34] br[34] wl[28] vdd gnd cell_6t
Xbit_r29_c34 bl[34] br[34] wl[29] vdd gnd cell_6t
Xbit_r30_c34 bl[34] br[34] wl[30] vdd gnd cell_6t
Xbit_r31_c34 bl[34] br[34] wl[31] vdd gnd cell_6t
Xbit_r32_c34 bl[34] br[34] wl[32] vdd gnd cell_6t
Xbit_r33_c34 bl[34] br[34] wl[33] vdd gnd cell_6t
Xbit_r34_c34 bl[34] br[34] wl[34] vdd gnd cell_6t
Xbit_r35_c34 bl[34] br[34] wl[35] vdd gnd cell_6t
Xbit_r36_c34 bl[34] br[34] wl[36] vdd gnd cell_6t
Xbit_r37_c34 bl[34] br[34] wl[37] vdd gnd cell_6t
Xbit_r38_c34 bl[34] br[34] wl[38] vdd gnd cell_6t
Xbit_r39_c34 bl[34] br[34] wl[39] vdd gnd cell_6t
Xbit_r40_c34 bl[34] br[34] wl[40] vdd gnd cell_6t
Xbit_r41_c34 bl[34] br[34] wl[41] vdd gnd cell_6t
Xbit_r42_c34 bl[34] br[34] wl[42] vdd gnd cell_6t
Xbit_r43_c34 bl[34] br[34] wl[43] vdd gnd cell_6t
Xbit_r44_c34 bl[34] br[34] wl[44] vdd gnd cell_6t
Xbit_r45_c34 bl[34] br[34] wl[45] vdd gnd cell_6t
Xbit_r46_c34 bl[34] br[34] wl[46] vdd gnd cell_6t
Xbit_r47_c34 bl[34] br[34] wl[47] vdd gnd cell_6t
Xbit_r48_c34 bl[34] br[34] wl[48] vdd gnd cell_6t
Xbit_r49_c34 bl[34] br[34] wl[49] vdd gnd cell_6t
Xbit_r50_c34 bl[34] br[34] wl[50] vdd gnd cell_6t
Xbit_r51_c34 bl[34] br[34] wl[51] vdd gnd cell_6t
Xbit_r52_c34 bl[34] br[34] wl[52] vdd gnd cell_6t
Xbit_r53_c34 bl[34] br[34] wl[53] vdd gnd cell_6t
Xbit_r54_c34 bl[34] br[34] wl[54] vdd gnd cell_6t
Xbit_r55_c34 bl[34] br[34] wl[55] vdd gnd cell_6t
Xbit_r56_c34 bl[34] br[34] wl[56] vdd gnd cell_6t
Xbit_r57_c34 bl[34] br[34] wl[57] vdd gnd cell_6t
Xbit_r58_c34 bl[34] br[34] wl[58] vdd gnd cell_6t
Xbit_r59_c34 bl[34] br[34] wl[59] vdd gnd cell_6t
Xbit_r60_c34 bl[34] br[34] wl[60] vdd gnd cell_6t
Xbit_r61_c34 bl[34] br[34] wl[61] vdd gnd cell_6t
Xbit_r62_c34 bl[34] br[34] wl[62] vdd gnd cell_6t
Xbit_r63_c34 bl[34] br[34] wl[63] vdd gnd cell_6t
Xbit_r64_c34 bl[34] br[34] wl[64] vdd gnd cell_6t
Xbit_r65_c34 bl[34] br[34] wl[65] vdd gnd cell_6t
Xbit_r66_c34 bl[34] br[34] wl[66] vdd gnd cell_6t
Xbit_r67_c34 bl[34] br[34] wl[67] vdd gnd cell_6t
Xbit_r68_c34 bl[34] br[34] wl[68] vdd gnd cell_6t
Xbit_r69_c34 bl[34] br[34] wl[69] vdd gnd cell_6t
Xbit_r70_c34 bl[34] br[34] wl[70] vdd gnd cell_6t
Xbit_r71_c34 bl[34] br[34] wl[71] vdd gnd cell_6t
Xbit_r72_c34 bl[34] br[34] wl[72] vdd gnd cell_6t
Xbit_r73_c34 bl[34] br[34] wl[73] vdd gnd cell_6t
Xbit_r74_c34 bl[34] br[34] wl[74] vdd gnd cell_6t
Xbit_r75_c34 bl[34] br[34] wl[75] vdd gnd cell_6t
Xbit_r76_c34 bl[34] br[34] wl[76] vdd gnd cell_6t
Xbit_r77_c34 bl[34] br[34] wl[77] vdd gnd cell_6t
Xbit_r78_c34 bl[34] br[34] wl[78] vdd gnd cell_6t
Xbit_r79_c34 bl[34] br[34] wl[79] vdd gnd cell_6t
Xbit_r80_c34 bl[34] br[34] wl[80] vdd gnd cell_6t
Xbit_r81_c34 bl[34] br[34] wl[81] vdd gnd cell_6t
Xbit_r82_c34 bl[34] br[34] wl[82] vdd gnd cell_6t
Xbit_r83_c34 bl[34] br[34] wl[83] vdd gnd cell_6t
Xbit_r84_c34 bl[34] br[34] wl[84] vdd gnd cell_6t
Xbit_r85_c34 bl[34] br[34] wl[85] vdd gnd cell_6t
Xbit_r86_c34 bl[34] br[34] wl[86] vdd gnd cell_6t
Xbit_r87_c34 bl[34] br[34] wl[87] vdd gnd cell_6t
Xbit_r88_c34 bl[34] br[34] wl[88] vdd gnd cell_6t
Xbit_r89_c34 bl[34] br[34] wl[89] vdd gnd cell_6t
Xbit_r90_c34 bl[34] br[34] wl[90] vdd gnd cell_6t
Xbit_r91_c34 bl[34] br[34] wl[91] vdd gnd cell_6t
Xbit_r92_c34 bl[34] br[34] wl[92] vdd gnd cell_6t
Xbit_r93_c34 bl[34] br[34] wl[93] vdd gnd cell_6t
Xbit_r94_c34 bl[34] br[34] wl[94] vdd gnd cell_6t
Xbit_r95_c34 bl[34] br[34] wl[95] vdd gnd cell_6t
Xbit_r96_c34 bl[34] br[34] wl[96] vdd gnd cell_6t
Xbit_r97_c34 bl[34] br[34] wl[97] vdd gnd cell_6t
Xbit_r98_c34 bl[34] br[34] wl[98] vdd gnd cell_6t
Xbit_r99_c34 bl[34] br[34] wl[99] vdd gnd cell_6t
Xbit_r100_c34 bl[34] br[34] wl[100] vdd gnd cell_6t
Xbit_r101_c34 bl[34] br[34] wl[101] vdd gnd cell_6t
Xbit_r102_c34 bl[34] br[34] wl[102] vdd gnd cell_6t
Xbit_r103_c34 bl[34] br[34] wl[103] vdd gnd cell_6t
Xbit_r104_c34 bl[34] br[34] wl[104] vdd gnd cell_6t
Xbit_r105_c34 bl[34] br[34] wl[105] vdd gnd cell_6t
Xbit_r106_c34 bl[34] br[34] wl[106] vdd gnd cell_6t
Xbit_r107_c34 bl[34] br[34] wl[107] vdd gnd cell_6t
Xbit_r108_c34 bl[34] br[34] wl[108] vdd gnd cell_6t
Xbit_r109_c34 bl[34] br[34] wl[109] vdd gnd cell_6t
Xbit_r110_c34 bl[34] br[34] wl[110] vdd gnd cell_6t
Xbit_r111_c34 bl[34] br[34] wl[111] vdd gnd cell_6t
Xbit_r112_c34 bl[34] br[34] wl[112] vdd gnd cell_6t
Xbit_r113_c34 bl[34] br[34] wl[113] vdd gnd cell_6t
Xbit_r114_c34 bl[34] br[34] wl[114] vdd gnd cell_6t
Xbit_r115_c34 bl[34] br[34] wl[115] vdd gnd cell_6t
Xbit_r116_c34 bl[34] br[34] wl[116] vdd gnd cell_6t
Xbit_r117_c34 bl[34] br[34] wl[117] vdd gnd cell_6t
Xbit_r118_c34 bl[34] br[34] wl[118] vdd gnd cell_6t
Xbit_r119_c34 bl[34] br[34] wl[119] vdd gnd cell_6t
Xbit_r120_c34 bl[34] br[34] wl[120] vdd gnd cell_6t
Xbit_r121_c34 bl[34] br[34] wl[121] vdd gnd cell_6t
Xbit_r122_c34 bl[34] br[34] wl[122] vdd gnd cell_6t
Xbit_r123_c34 bl[34] br[34] wl[123] vdd gnd cell_6t
Xbit_r124_c34 bl[34] br[34] wl[124] vdd gnd cell_6t
Xbit_r125_c34 bl[34] br[34] wl[125] vdd gnd cell_6t
Xbit_r126_c34 bl[34] br[34] wl[126] vdd gnd cell_6t
Xbit_r127_c34 bl[34] br[34] wl[127] vdd gnd cell_6t
Xbit_r128_c34 bl[34] br[34] wl[128] vdd gnd cell_6t
Xbit_r129_c34 bl[34] br[34] wl[129] vdd gnd cell_6t
Xbit_r130_c34 bl[34] br[34] wl[130] vdd gnd cell_6t
Xbit_r131_c34 bl[34] br[34] wl[131] vdd gnd cell_6t
Xbit_r132_c34 bl[34] br[34] wl[132] vdd gnd cell_6t
Xbit_r133_c34 bl[34] br[34] wl[133] vdd gnd cell_6t
Xbit_r134_c34 bl[34] br[34] wl[134] vdd gnd cell_6t
Xbit_r135_c34 bl[34] br[34] wl[135] vdd gnd cell_6t
Xbit_r136_c34 bl[34] br[34] wl[136] vdd gnd cell_6t
Xbit_r137_c34 bl[34] br[34] wl[137] vdd gnd cell_6t
Xbit_r138_c34 bl[34] br[34] wl[138] vdd gnd cell_6t
Xbit_r139_c34 bl[34] br[34] wl[139] vdd gnd cell_6t
Xbit_r140_c34 bl[34] br[34] wl[140] vdd gnd cell_6t
Xbit_r141_c34 bl[34] br[34] wl[141] vdd gnd cell_6t
Xbit_r142_c34 bl[34] br[34] wl[142] vdd gnd cell_6t
Xbit_r143_c34 bl[34] br[34] wl[143] vdd gnd cell_6t
Xbit_r144_c34 bl[34] br[34] wl[144] vdd gnd cell_6t
Xbit_r145_c34 bl[34] br[34] wl[145] vdd gnd cell_6t
Xbit_r146_c34 bl[34] br[34] wl[146] vdd gnd cell_6t
Xbit_r147_c34 bl[34] br[34] wl[147] vdd gnd cell_6t
Xbit_r148_c34 bl[34] br[34] wl[148] vdd gnd cell_6t
Xbit_r149_c34 bl[34] br[34] wl[149] vdd gnd cell_6t
Xbit_r150_c34 bl[34] br[34] wl[150] vdd gnd cell_6t
Xbit_r151_c34 bl[34] br[34] wl[151] vdd gnd cell_6t
Xbit_r152_c34 bl[34] br[34] wl[152] vdd gnd cell_6t
Xbit_r153_c34 bl[34] br[34] wl[153] vdd gnd cell_6t
Xbit_r154_c34 bl[34] br[34] wl[154] vdd gnd cell_6t
Xbit_r155_c34 bl[34] br[34] wl[155] vdd gnd cell_6t
Xbit_r156_c34 bl[34] br[34] wl[156] vdd gnd cell_6t
Xbit_r157_c34 bl[34] br[34] wl[157] vdd gnd cell_6t
Xbit_r158_c34 bl[34] br[34] wl[158] vdd gnd cell_6t
Xbit_r159_c34 bl[34] br[34] wl[159] vdd gnd cell_6t
Xbit_r160_c34 bl[34] br[34] wl[160] vdd gnd cell_6t
Xbit_r161_c34 bl[34] br[34] wl[161] vdd gnd cell_6t
Xbit_r162_c34 bl[34] br[34] wl[162] vdd gnd cell_6t
Xbit_r163_c34 bl[34] br[34] wl[163] vdd gnd cell_6t
Xbit_r164_c34 bl[34] br[34] wl[164] vdd gnd cell_6t
Xbit_r165_c34 bl[34] br[34] wl[165] vdd gnd cell_6t
Xbit_r166_c34 bl[34] br[34] wl[166] vdd gnd cell_6t
Xbit_r167_c34 bl[34] br[34] wl[167] vdd gnd cell_6t
Xbit_r168_c34 bl[34] br[34] wl[168] vdd gnd cell_6t
Xbit_r169_c34 bl[34] br[34] wl[169] vdd gnd cell_6t
Xbit_r170_c34 bl[34] br[34] wl[170] vdd gnd cell_6t
Xbit_r171_c34 bl[34] br[34] wl[171] vdd gnd cell_6t
Xbit_r172_c34 bl[34] br[34] wl[172] vdd gnd cell_6t
Xbit_r173_c34 bl[34] br[34] wl[173] vdd gnd cell_6t
Xbit_r174_c34 bl[34] br[34] wl[174] vdd gnd cell_6t
Xbit_r175_c34 bl[34] br[34] wl[175] vdd gnd cell_6t
Xbit_r176_c34 bl[34] br[34] wl[176] vdd gnd cell_6t
Xbit_r177_c34 bl[34] br[34] wl[177] vdd gnd cell_6t
Xbit_r178_c34 bl[34] br[34] wl[178] vdd gnd cell_6t
Xbit_r179_c34 bl[34] br[34] wl[179] vdd gnd cell_6t
Xbit_r180_c34 bl[34] br[34] wl[180] vdd gnd cell_6t
Xbit_r181_c34 bl[34] br[34] wl[181] vdd gnd cell_6t
Xbit_r182_c34 bl[34] br[34] wl[182] vdd gnd cell_6t
Xbit_r183_c34 bl[34] br[34] wl[183] vdd gnd cell_6t
Xbit_r184_c34 bl[34] br[34] wl[184] vdd gnd cell_6t
Xbit_r185_c34 bl[34] br[34] wl[185] vdd gnd cell_6t
Xbit_r186_c34 bl[34] br[34] wl[186] vdd gnd cell_6t
Xbit_r187_c34 bl[34] br[34] wl[187] vdd gnd cell_6t
Xbit_r188_c34 bl[34] br[34] wl[188] vdd gnd cell_6t
Xbit_r189_c34 bl[34] br[34] wl[189] vdd gnd cell_6t
Xbit_r190_c34 bl[34] br[34] wl[190] vdd gnd cell_6t
Xbit_r191_c34 bl[34] br[34] wl[191] vdd gnd cell_6t
Xbit_r192_c34 bl[34] br[34] wl[192] vdd gnd cell_6t
Xbit_r193_c34 bl[34] br[34] wl[193] vdd gnd cell_6t
Xbit_r194_c34 bl[34] br[34] wl[194] vdd gnd cell_6t
Xbit_r195_c34 bl[34] br[34] wl[195] vdd gnd cell_6t
Xbit_r196_c34 bl[34] br[34] wl[196] vdd gnd cell_6t
Xbit_r197_c34 bl[34] br[34] wl[197] vdd gnd cell_6t
Xbit_r198_c34 bl[34] br[34] wl[198] vdd gnd cell_6t
Xbit_r199_c34 bl[34] br[34] wl[199] vdd gnd cell_6t
Xbit_r200_c34 bl[34] br[34] wl[200] vdd gnd cell_6t
Xbit_r201_c34 bl[34] br[34] wl[201] vdd gnd cell_6t
Xbit_r202_c34 bl[34] br[34] wl[202] vdd gnd cell_6t
Xbit_r203_c34 bl[34] br[34] wl[203] vdd gnd cell_6t
Xbit_r204_c34 bl[34] br[34] wl[204] vdd gnd cell_6t
Xbit_r205_c34 bl[34] br[34] wl[205] vdd gnd cell_6t
Xbit_r206_c34 bl[34] br[34] wl[206] vdd gnd cell_6t
Xbit_r207_c34 bl[34] br[34] wl[207] vdd gnd cell_6t
Xbit_r208_c34 bl[34] br[34] wl[208] vdd gnd cell_6t
Xbit_r209_c34 bl[34] br[34] wl[209] vdd gnd cell_6t
Xbit_r210_c34 bl[34] br[34] wl[210] vdd gnd cell_6t
Xbit_r211_c34 bl[34] br[34] wl[211] vdd gnd cell_6t
Xbit_r212_c34 bl[34] br[34] wl[212] vdd gnd cell_6t
Xbit_r213_c34 bl[34] br[34] wl[213] vdd gnd cell_6t
Xbit_r214_c34 bl[34] br[34] wl[214] vdd gnd cell_6t
Xbit_r215_c34 bl[34] br[34] wl[215] vdd gnd cell_6t
Xbit_r216_c34 bl[34] br[34] wl[216] vdd gnd cell_6t
Xbit_r217_c34 bl[34] br[34] wl[217] vdd gnd cell_6t
Xbit_r218_c34 bl[34] br[34] wl[218] vdd gnd cell_6t
Xbit_r219_c34 bl[34] br[34] wl[219] vdd gnd cell_6t
Xbit_r220_c34 bl[34] br[34] wl[220] vdd gnd cell_6t
Xbit_r221_c34 bl[34] br[34] wl[221] vdd gnd cell_6t
Xbit_r222_c34 bl[34] br[34] wl[222] vdd gnd cell_6t
Xbit_r223_c34 bl[34] br[34] wl[223] vdd gnd cell_6t
Xbit_r224_c34 bl[34] br[34] wl[224] vdd gnd cell_6t
Xbit_r225_c34 bl[34] br[34] wl[225] vdd gnd cell_6t
Xbit_r226_c34 bl[34] br[34] wl[226] vdd gnd cell_6t
Xbit_r227_c34 bl[34] br[34] wl[227] vdd gnd cell_6t
Xbit_r228_c34 bl[34] br[34] wl[228] vdd gnd cell_6t
Xbit_r229_c34 bl[34] br[34] wl[229] vdd gnd cell_6t
Xbit_r230_c34 bl[34] br[34] wl[230] vdd gnd cell_6t
Xbit_r231_c34 bl[34] br[34] wl[231] vdd gnd cell_6t
Xbit_r232_c34 bl[34] br[34] wl[232] vdd gnd cell_6t
Xbit_r233_c34 bl[34] br[34] wl[233] vdd gnd cell_6t
Xbit_r234_c34 bl[34] br[34] wl[234] vdd gnd cell_6t
Xbit_r235_c34 bl[34] br[34] wl[235] vdd gnd cell_6t
Xbit_r236_c34 bl[34] br[34] wl[236] vdd gnd cell_6t
Xbit_r237_c34 bl[34] br[34] wl[237] vdd gnd cell_6t
Xbit_r238_c34 bl[34] br[34] wl[238] vdd gnd cell_6t
Xbit_r239_c34 bl[34] br[34] wl[239] vdd gnd cell_6t
Xbit_r240_c34 bl[34] br[34] wl[240] vdd gnd cell_6t
Xbit_r241_c34 bl[34] br[34] wl[241] vdd gnd cell_6t
Xbit_r242_c34 bl[34] br[34] wl[242] vdd gnd cell_6t
Xbit_r243_c34 bl[34] br[34] wl[243] vdd gnd cell_6t
Xbit_r244_c34 bl[34] br[34] wl[244] vdd gnd cell_6t
Xbit_r245_c34 bl[34] br[34] wl[245] vdd gnd cell_6t
Xbit_r246_c34 bl[34] br[34] wl[246] vdd gnd cell_6t
Xbit_r247_c34 bl[34] br[34] wl[247] vdd gnd cell_6t
Xbit_r248_c34 bl[34] br[34] wl[248] vdd gnd cell_6t
Xbit_r249_c34 bl[34] br[34] wl[249] vdd gnd cell_6t
Xbit_r250_c34 bl[34] br[34] wl[250] vdd gnd cell_6t
Xbit_r251_c34 bl[34] br[34] wl[251] vdd gnd cell_6t
Xbit_r252_c34 bl[34] br[34] wl[252] vdd gnd cell_6t
Xbit_r253_c34 bl[34] br[34] wl[253] vdd gnd cell_6t
Xbit_r254_c34 bl[34] br[34] wl[254] vdd gnd cell_6t
Xbit_r255_c34 bl[34] br[34] wl[255] vdd gnd cell_6t
Xbit_r0_c35 bl[35] br[35] wl[0] vdd gnd cell_6t
Xbit_r1_c35 bl[35] br[35] wl[1] vdd gnd cell_6t
Xbit_r2_c35 bl[35] br[35] wl[2] vdd gnd cell_6t
Xbit_r3_c35 bl[35] br[35] wl[3] vdd gnd cell_6t
Xbit_r4_c35 bl[35] br[35] wl[4] vdd gnd cell_6t
Xbit_r5_c35 bl[35] br[35] wl[5] vdd gnd cell_6t
Xbit_r6_c35 bl[35] br[35] wl[6] vdd gnd cell_6t
Xbit_r7_c35 bl[35] br[35] wl[7] vdd gnd cell_6t
Xbit_r8_c35 bl[35] br[35] wl[8] vdd gnd cell_6t
Xbit_r9_c35 bl[35] br[35] wl[9] vdd gnd cell_6t
Xbit_r10_c35 bl[35] br[35] wl[10] vdd gnd cell_6t
Xbit_r11_c35 bl[35] br[35] wl[11] vdd gnd cell_6t
Xbit_r12_c35 bl[35] br[35] wl[12] vdd gnd cell_6t
Xbit_r13_c35 bl[35] br[35] wl[13] vdd gnd cell_6t
Xbit_r14_c35 bl[35] br[35] wl[14] vdd gnd cell_6t
Xbit_r15_c35 bl[35] br[35] wl[15] vdd gnd cell_6t
Xbit_r16_c35 bl[35] br[35] wl[16] vdd gnd cell_6t
Xbit_r17_c35 bl[35] br[35] wl[17] vdd gnd cell_6t
Xbit_r18_c35 bl[35] br[35] wl[18] vdd gnd cell_6t
Xbit_r19_c35 bl[35] br[35] wl[19] vdd gnd cell_6t
Xbit_r20_c35 bl[35] br[35] wl[20] vdd gnd cell_6t
Xbit_r21_c35 bl[35] br[35] wl[21] vdd gnd cell_6t
Xbit_r22_c35 bl[35] br[35] wl[22] vdd gnd cell_6t
Xbit_r23_c35 bl[35] br[35] wl[23] vdd gnd cell_6t
Xbit_r24_c35 bl[35] br[35] wl[24] vdd gnd cell_6t
Xbit_r25_c35 bl[35] br[35] wl[25] vdd gnd cell_6t
Xbit_r26_c35 bl[35] br[35] wl[26] vdd gnd cell_6t
Xbit_r27_c35 bl[35] br[35] wl[27] vdd gnd cell_6t
Xbit_r28_c35 bl[35] br[35] wl[28] vdd gnd cell_6t
Xbit_r29_c35 bl[35] br[35] wl[29] vdd gnd cell_6t
Xbit_r30_c35 bl[35] br[35] wl[30] vdd gnd cell_6t
Xbit_r31_c35 bl[35] br[35] wl[31] vdd gnd cell_6t
Xbit_r32_c35 bl[35] br[35] wl[32] vdd gnd cell_6t
Xbit_r33_c35 bl[35] br[35] wl[33] vdd gnd cell_6t
Xbit_r34_c35 bl[35] br[35] wl[34] vdd gnd cell_6t
Xbit_r35_c35 bl[35] br[35] wl[35] vdd gnd cell_6t
Xbit_r36_c35 bl[35] br[35] wl[36] vdd gnd cell_6t
Xbit_r37_c35 bl[35] br[35] wl[37] vdd gnd cell_6t
Xbit_r38_c35 bl[35] br[35] wl[38] vdd gnd cell_6t
Xbit_r39_c35 bl[35] br[35] wl[39] vdd gnd cell_6t
Xbit_r40_c35 bl[35] br[35] wl[40] vdd gnd cell_6t
Xbit_r41_c35 bl[35] br[35] wl[41] vdd gnd cell_6t
Xbit_r42_c35 bl[35] br[35] wl[42] vdd gnd cell_6t
Xbit_r43_c35 bl[35] br[35] wl[43] vdd gnd cell_6t
Xbit_r44_c35 bl[35] br[35] wl[44] vdd gnd cell_6t
Xbit_r45_c35 bl[35] br[35] wl[45] vdd gnd cell_6t
Xbit_r46_c35 bl[35] br[35] wl[46] vdd gnd cell_6t
Xbit_r47_c35 bl[35] br[35] wl[47] vdd gnd cell_6t
Xbit_r48_c35 bl[35] br[35] wl[48] vdd gnd cell_6t
Xbit_r49_c35 bl[35] br[35] wl[49] vdd gnd cell_6t
Xbit_r50_c35 bl[35] br[35] wl[50] vdd gnd cell_6t
Xbit_r51_c35 bl[35] br[35] wl[51] vdd gnd cell_6t
Xbit_r52_c35 bl[35] br[35] wl[52] vdd gnd cell_6t
Xbit_r53_c35 bl[35] br[35] wl[53] vdd gnd cell_6t
Xbit_r54_c35 bl[35] br[35] wl[54] vdd gnd cell_6t
Xbit_r55_c35 bl[35] br[35] wl[55] vdd gnd cell_6t
Xbit_r56_c35 bl[35] br[35] wl[56] vdd gnd cell_6t
Xbit_r57_c35 bl[35] br[35] wl[57] vdd gnd cell_6t
Xbit_r58_c35 bl[35] br[35] wl[58] vdd gnd cell_6t
Xbit_r59_c35 bl[35] br[35] wl[59] vdd gnd cell_6t
Xbit_r60_c35 bl[35] br[35] wl[60] vdd gnd cell_6t
Xbit_r61_c35 bl[35] br[35] wl[61] vdd gnd cell_6t
Xbit_r62_c35 bl[35] br[35] wl[62] vdd gnd cell_6t
Xbit_r63_c35 bl[35] br[35] wl[63] vdd gnd cell_6t
Xbit_r64_c35 bl[35] br[35] wl[64] vdd gnd cell_6t
Xbit_r65_c35 bl[35] br[35] wl[65] vdd gnd cell_6t
Xbit_r66_c35 bl[35] br[35] wl[66] vdd gnd cell_6t
Xbit_r67_c35 bl[35] br[35] wl[67] vdd gnd cell_6t
Xbit_r68_c35 bl[35] br[35] wl[68] vdd gnd cell_6t
Xbit_r69_c35 bl[35] br[35] wl[69] vdd gnd cell_6t
Xbit_r70_c35 bl[35] br[35] wl[70] vdd gnd cell_6t
Xbit_r71_c35 bl[35] br[35] wl[71] vdd gnd cell_6t
Xbit_r72_c35 bl[35] br[35] wl[72] vdd gnd cell_6t
Xbit_r73_c35 bl[35] br[35] wl[73] vdd gnd cell_6t
Xbit_r74_c35 bl[35] br[35] wl[74] vdd gnd cell_6t
Xbit_r75_c35 bl[35] br[35] wl[75] vdd gnd cell_6t
Xbit_r76_c35 bl[35] br[35] wl[76] vdd gnd cell_6t
Xbit_r77_c35 bl[35] br[35] wl[77] vdd gnd cell_6t
Xbit_r78_c35 bl[35] br[35] wl[78] vdd gnd cell_6t
Xbit_r79_c35 bl[35] br[35] wl[79] vdd gnd cell_6t
Xbit_r80_c35 bl[35] br[35] wl[80] vdd gnd cell_6t
Xbit_r81_c35 bl[35] br[35] wl[81] vdd gnd cell_6t
Xbit_r82_c35 bl[35] br[35] wl[82] vdd gnd cell_6t
Xbit_r83_c35 bl[35] br[35] wl[83] vdd gnd cell_6t
Xbit_r84_c35 bl[35] br[35] wl[84] vdd gnd cell_6t
Xbit_r85_c35 bl[35] br[35] wl[85] vdd gnd cell_6t
Xbit_r86_c35 bl[35] br[35] wl[86] vdd gnd cell_6t
Xbit_r87_c35 bl[35] br[35] wl[87] vdd gnd cell_6t
Xbit_r88_c35 bl[35] br[35] wl[88] vdd gnd cell_6t
Xbit_r89_c35 bl[35] br[35] wl[89] vdd gnd cell_6t
Xbit_r90_c35 bl[35] br[35] wl[90] vdd gnd cell_6t
Xbit_r91_c35 bl[35] br[35] wl[91] vdd gnd cell_6t
Xbit_r92_c35 bl[35] br[35] wl[92] vdd gnd cell_6t
Xbit_r93_c35 bl[35] br[35] wl[93] vdd gnd cell_6t
Xbit_r94_c35 bl[35] br[35] wl[94] vdd gnd cell_6t
Xbit_r95_c35 bl[35] br[35] wl[95] vdd gnd cell_6t
Xbit_r96_c35 bl[35] br[35] wl[96] vdd gnd cell_6t
Xbit_r97_c35 bl[35] br[35] wl[97] vdd gnd cell_6t
Xbit_r98_c35 bl[35] br[35] wl[98] vdd gnd cell_6t
Xbit_r99_c35 bl[35] br[35] wl[99] vdd gnd cell_6t
Xbit_r100_c35 bl[35] br[35] wl[100] vdd gnd cell_6t
Xbit_r101_c35 bl[35] br[35] wl[101] vdd gnd cell_6t
Xbit_r102_c35 bl[35] br[35] wl[102] vdd gnd cell_6t
Xbit_r103_c35 bl[35] br[35] wl[103] vdd gnd cell_6t
Xbit_r104_c35 bl[35] br[35] wl[104] vdd gnd cell_6t
Xbit_r105_c35 bl[35] br[35] wl[105] vdd gnd cell_6t
Xbit_r106_c35 bl[35] br[35] wl[106] vdd gnd cell_6t
Xbit_r107_c35 bl[35] br[35] wl[107] vdd gnd cell_6t
Xbit_r108_c35 bl[35] br[35] wl[108] vdd gnd cell_6t
Xbit_r109_c35 bl[35] br[35] wl[109] vdd gnd cell_6t
Xbit_r110_c35 bl[35] br[35] wl[110] vdd gnd cell_6t
Xbit_r111_c35 bl[35] br[35] wl[111] vdd gnd cell_6t
Xbit_r112_c35 bl[35] br[35] wl[112] vdd gnd cell_6t
Xbit_r113_c35 bl[35] br[35] wl[113] vdd gnd cell_6t
Xbit_r114_c35 bl[35] br[35] wl[114] vdd gnd cell_6t
Xbit_r115_c35 bl[35] br[35] wl[115] vdd gnd cell_6t
Xbit_r116_c35 bl[35] br[35] wl[116] vdd gnd cell_6t
Xbit_r117_c35 bl[35] br[35] wl[117] vdd gnd cell_6t
Xbit_r118_c35 bl[35] br[35] wl[118] vdd gnd cell_6t
Xbit_r119_c35 bl[35] br[35] wl[119] vdd gnd cell_6t
Xbit_r120_c35 bl[35] br[35] wl[120] vdd gnd cell_6t
Xbit_r121_c35 bl[35] br[35] wl[121] vdd gnd cell_6t
Xbit_r122_c35 bl[35] br[35] wl[122] vdd gnd cell_6t
Xbit_r123_c35 bl[35] br[35] wl[123] vdd gnd cell_6t
Xbit_r124_c35 bl[35] br[35] wl[124] vdd gnd cell_6t
Xbit_r125_c35 bl[35] br[35] wl[125] vdd gnd cell_6t
Xbit_r126_c35 bl[35] br[35] wl[126] vdd gnd cell_6t
Xbit_r127_c35 bl[35] br[35] wl[127] vdd gnd cell_6t
Xbit_r128_c35 bl[35] br[35] wl[128] vdd gnd cell_6t
Xbit_r129_c35 bl[35] br[35] wl[129] vdd gnd cell_6t
Xbit_r130_c35 bl[35] br[35] wl[130] vdd gnd cell_6t
Xbit_r131_c35 bl[35] br[35] wl[131] vdd gnd cell_6t
Xbit_r132_c35 bl[35] br[35] wl[132] vdd gnd cell_6t
Xbit_r133_c35 bl[35] br[35] wl[133] vdd gnd cell_6t
Xbit_r134_c35 bl[35] br[35] wl[134] vdd gnd cell_6t
Xbit_r135_c35 bl[35] br[35] wl[135] vdd gnd cell_6t
Xbit_r136_c35 bl[35] br[35] wl[136] vdd gnd cell_6t
Xbit_r137_c35 bl[35] br[35] wl[137] vdd gnd cell_6t
Xbit_r138_c35 bl[35] br[35] wl[138] vdd gnd cell_6t
Xbit_r139_c35 bl[35] br[35] wl[139] vdd gnd cell_6t
Xbit_r140_c35 bl[35] br[35] wl[140] vdd gnd cell_6t
Xbit_r141_c35 bl[35] br[35] wl[141] vdd gnd cell_6t
Xbit_r142_c35 bl[35] br[35] wl[142] vdd gnd cell_6t
Xbit_r143_c35 bl[35] br[35] wl[143] vdd gnd cell_6t
Xbit_r144_c35 bl[35] br[35] wl[144] vdd gnd cell_6t
Xbit_r145_c35 bl[35] br[35] wl[145] vdd gnd cell_6t
Xbit_r146_c35 bl[35] br[35] wl[146] vdd gnd cell_6t
Xbit_r147_c35 bl[35] br[35] wl[147] vdd gnd cell_6t
Xbit_r148_c35 bl[35] br[35] wl[148] vdd gnd cell_6t
Xbit_r149_c35 bl[35] br[35] wl[149] vdd gnd cell_6t
Xbit_r150_c35 bl[35] br[35] wl[150] vdd gnd cell_6t
Xbit_r151_c35 bl[35] br[35] wl[151] vdd gnd cell_6t
Xbit_r152_c35 bl[35] br[35] wl[152] vdd gnd cell_6t
Xbit_r153_c35 bl[35] br[35] wl[153] vdd gnd cell_6t
Xbit_r154_c35 bl[35] br[35] wl[154] vdd gnd cell_6t
Xbit_r155_c35 bl[35] br[35] wl[155] vdd gnd cell_6t
Xbit_r156_c35 bl[35] br[35] wl[156] vdd gnd cell_6t
Xbit_r157_c35 bl[35] br[35] wl[157] vdd gnd cell_6t
Xbit_r158_c35 bl[35] br[35] wl[158] vdd gnd cell_6t
Xbit_r159_c35 bl[35] br[35] wl[159] vdd gnd cell_6t
Xbit_r160_c35 bl[35] br[35] wl[160] vdd gnd cell_6t
Xbit_r161_c35 bl[35] br[35] wl[161] vdd gnd cell_6t
Xbit_r162_c35 bl[35] br[35] wl[162] vdd gnd cell_6t
Xbit_r163_c35 bl[35] br[35] wl[163] vdd gnd cell_6t
Xbit_r164_c35 bl[35] br[35] wl[164] vdd gnd cell_6t
Xbit_r165_c35 bl[35] br[35] wl[165] vdd gnd cell_6t
Xbit_r166_c35 bl[35] br[35] wl[166] vdd gnd cell_6t
Xbit_r167_c35 bl[35] br[35] wl[167] vdd gnd cell_6t
Xbit_r168_c35 bl[35] br[35] wl[168] vdd gnd cell_6t
Xbit_r169_c35 bl[35] br[35] wl[169] vdd gnd cell_6t
Xbit_r170_c35 bl[35] br[35] wl[170] vdd gnd cell_6t
Xbit_r171_c35 bl[35] br[35] wl[171] vdd gnd cell_6t
Xbit_r172_c35 bl[35] br[35] wl[172] vdd gnd cell_6t
Xbit_r173_c35 bl[35] br[35] wl[173] vdd gnd cell_6t
Xbit_r174_c35 bl[35] br[35] wl[174] vdd gnd cell_6t
Xbit_r175_c35 bl[35] br[35] wl[175] vdd gnd cell_6t
Xbit_r176_c35 bl[35] br[35] wl[176] vdd gnd cell_6t
Xbit_r177_c35 bl[35] br[35] wl[177] vdd gnd cell_6t
Xbit_r178_c35 bl[35] br[35] wl[178] vdd gnd cell_6t
Xbit_r179_c35 bl[35] br[35] wl[179] vdd gnd cell_6t
Xbit_r180_c35 bl[35] br[35] wl[180] vdd gnd cell_6t
Xbit_r181_c35 bl[35] br[35] wl[181] vdd gnd cell_6t
Xbit_r182_c35 bl[35] br[35] wl[182] vdd gnd cell_6t
Xbit_r183_c35 bl[35] br[35] wl[183] vdd gnd cell_6t
Xbit_r184_c35 bl[35] br[35] wl[184] vdd gnd cell_6t
Xbit_r185_c35 bl[35] br[35] wl[185] vdd gnd cell_6t
Xbit_r186_c35 bl[35] br[35] wl[186] vdd gnd cell_6t
Xbit_r187_c35 bl[35] br[35] wl[187] vdd gnd cell_6t
Xbit_r188_c35 bl[35] br[35] wl[188] vdd gnd cell_6t
Xbit_r189_c35 bl[35] br[35] wl[189] vdd gnd cell_6t
Xbit_r190_c35 bl[35] br[35] wl[190] vdd gnd cell_6t
Xbit_r191_c35 bl[35] br[35] wl[191] vdd gnd cell_6t
Xbit_r192_c35 bl[35] br[35] wl[192] vdd gnd cell_6t
Xbit_r193_c35 bl[35] br[35] wl[193] vdd gnd cell_6t
Xbit_r194_c35 bl[35] br[35] wl[194] vdd gnd cell_6t
Xbit_r195_c35 bl[35] br[35] wl[195] vdd gnd cell_6t
Xbit_r196_c35 bl[35] br[35] wl[196] vdd gnd cell_6t
Xbit_r197_c35 bl[35] br[35] wl[197] vdd gnd cell_6t
Xbit_r198_c35 bl[35] br[35] wl[198] vdd gnd cell_6t
Xbit_r199_c35 bl[35] br[35] wl[199] vdd gnd cell_6t
Xbit_r200_c35 bl[35] br[35] wl[200] vdd gnd cell_6t
Xbit_r201_c35 bl[35] br[35] wl[201] vdd gnd cell_6t
Xbit_r202_c35 bl[35] br[35] wl[202] vdd gnd cell_6t
Xbit_r203_c35 bl[35] br[35] wl[203] vdd gnd cell_6t
Xbit_r204_c35 bl[35] br[35] wl[204] vdd gnd cell_6t
Xbit_r205_c35 bl[35] br[35] wl[205] vdd gnd cell_6t
Xbit_r206_c35 bl[35] br[35] wl[206] vdd gnd cell_6t
Xbit_r207_c35 bl[35] br[35] wl[207] vdd gnd cell_6t
Xbit_r208_c35 bl[35] br[35] wl[208] vdd gnd cell_6t
Xbit_r209_c35 bl[35] br[35] wl[209] vdd gnd cell_6t
Xbit_r210_c35 bl[35] br[35] wl[210] vdd gnd cell_6t
Xbit_r211_c35 bl[35] br[35] wl[211] vdd gnd cell_6t
Xbit_r212_c35 bl[35] br[35] wl[212] vdd gnd cell_6t
Xbit_r213_c35 bl[35] br[35] wl[213] vdd gnd cell_6t
Xbit_r214_c35 bl[35] br[35] wl[214] vdd gnd cell_6t
Xbit_r215_c35 bl[35] br[35] wl[215] vdd gnd cell_6t
Xbit_r216_c35 bl[35] br[35] wl[216] vdd gnd cell_6t
Xbit_r217_c35 bl[35] br[35] wl[217] vdd gnd cell_6t
Xbit_r218_c35 bl[35] br[35] wl[218] vdd gnd cell_6t
Xbit_r219_c35 bl[35] br[35] wl[219] vdd gnd cell_6t
Xbit_r220_c35 bl[35] br[35] wl[220] vdd gnd cell_6t
Xbit_r221_c35 bl[35] br[35] wl[221] vdd gnd cell_6t
Xbit_r222_c35 bl[35] br[35] wl[222] vdd gnd cell_6t
Xbit_r223_c35 bl[35] br[35] wl[223] vdd gnd cell_6t
Xbit_r224_c35 bl[35] br[35] wl[224] vdd gnd cell_6t
Xbit_r225_c35 bl[35] br[35] wl[225] vdd gnd cell_6t
Xbit_r226_c35 bl[35] br[35] wl[226] vdd gnd cell_6t
Xbit_r227_c35 bl[35] br[35] wl[227] vdd gnd cell_6t
Xbit_r228_c35 bl[35] br[35] wl[228] vdd gnd cell_6t
Xbit_r229_c35 bl[35] br[35] wl[229] vdd gnd cell_6t
Xbit_r230_c35 bl[35] br[35] wl[230] vdd gnd cell_6t
Xbit_r231_c35 bl[35] br[35] wl[231] vdd gnd cell_6t
Xbit_r232_c35 bl[35] br[35] wl[232] vdd gnd cell_6t
Xbit_r233_c35 bl[35] br[35] wl[233] vdd gnd cell_6t
Xbit_r234_c35 bl[35] br[35] wl[234] vdd gnd cell_6t
Xbit_r235_c35 bl[35] br[35] wl[235] vdd gnd cell_6t
Xbit_r236_c35 bl[35] br[35] wl[236] vdd gnd cell_6t
Xbit_r237_c35 bl[35] br[35] wl[237] vdd gnd cell_6t
Xbit_r238_c35 bl[35] br[35] wl[238] vdd gnd cell_6t
Xbit_r239_c35 bl[35] br[35] wl[239] vdd gnd cell_6t
Xbit_r240_c35 bl[35] br[35] wl[240] vdd gnd cell_6t
Xbit_r241_c35 bl[35] br[35] wl[241] vdd gnd cell_6t
Xbit_r242_c35 bl[35] br[35] wl[242] vdd gnd cell_6t
Xbit_r243_c35 bl[35] br[35] wl[243] vdd gnd cell_6t
Xbit_r244_c35 bl[35] br[35] wl[244] vdd gnd cell_6t
Xbit_r245_c35 bl[35] br[35] wl[245] vdd gnd cell_6t
Xbit_r246_c35 bl[35] br[35] wl[246] vdd gnd cell_6t
Xbit_r247_c35 bl[35] br[35] wl[247] vdd gnd cell_6t
Xbit_r248_c35 bl[35] br[35] wl[248] vdd gnd cell_6t
Xbit_r249_c35 bl[35] br[35] wl[249] vdd gnd cell_6t
Xbit_r250_c35 bl[35] br[35] wl[250] vdd gnd cell_6t
Xbit_r251_c35 bl[35] br[35] wl[251] vdd gnd cell_6t
Xbit_r252_c35 bl[35] br[35] wl[252] vdd gnd cell_6t
Xbit_r253_c35 bl[35] br[35] wl[253] vdd gnd cell_6t
Xbit_r254_c35 bl[35] br[35] wl[254] vdd gnd cell_6t
Xbit_r255_c35 bl[35] br[35] wl[255] vdd gnd cell_6t
Xbit_r0_c36 bl[36] br[36] wl[0] vdd gnd cell_6t
Xbit_r1_c36 bl[36] br[36] wl[1] vdd gnd cell_6t
Xbit_r2_c36 bl[36] br[36] wl[2] vdd gnd cell_6t
Xbit_r3_c36 bl[36] br[36] wl[3] vdd gnd cell_6t
Xbit_r4_c36 bl[36] br[36] wl[4] vdd gnd cell_6t
Xbit_r5_c36 bl[36] br[36] wl[5] vdd gnd cell_6t
Xbit_r6_c36 bl[36] br[36] wl[6] vdd gnd cell_6t
Xbit_r7_c36 bl[36] br[36] wl[7] vdd gnd cell_6t
Xbit_r8_c36 bl[36] br[36] wl[8] vdd gnd cell_6t
Xbit_r9_c36 bl[36] br[36] wl[9] vdd gnd cell_6t
Xbit_r10_c36 bl[36] br[36] wl[10] vdd gnd cell_6t
Xbit_r11_c36 bl[36] br[36] wl[11] vdd gnd cell_6t
Xbit_r12_c36 bl[36] br[36] wl[12] vdd gnd cell_6t
Xbit_r13_c36 bl[36] br[36] wl[13] vdd gnd cell_6t
Xbit_r14_c36 bl[36] br[36] wl[14] vdd gnd cell_6t
Xbit_r15_c36 bl[36] br[36] wl[15] vdd gnd cell_6t
Xbit_r16_c36 bl[36] br[36] wl[16] vdd gnd cell_6t
Xbit_r17_c36 bl[36] br[36] wl[17] vdd gnd cell_6t
Xbit_r18_c36 bl[36] br[36] wl[18] vdd gnd cell_6t
Xbit_r19_c36 bl[36] br[36] wl[19] vdd gnd cell_6t
Xbit_r20_c36 bl[36] br[36] wl[20] vdd gnd cell_6t
Xbit_r21_c36 bl[36] br[36] wl[21] vdd gnd cell_6t
Xbit_r22_c36 bl[36] br[36] wl[22] vdd gnd cell_6t
Xbit_r23_c36 bl[36] br[36] wl[23] vdd gnd cell_6t
Xbit_r24_c36 bl[36] br[36] wl[24] vdd gnd cell_6t
Xbit_r25_c36 bl[36] br[36] wl[25] vdd gnd cell_6t
Xbit_r26_c36 bl[36] br[36] wl[26] vdd gnd cell_6t
Xbit_r27_c36 bl[36] br[36] wl[27] vdd gnd cell_6t
Xbit_r28_c36 bl[36] br[36] wl[28] vdd gnd cell_6t
Xbit_r29_c36 bl[36] br[36] wl[29] vdd gnd cell_6t
Xbit_r30_c36 bl[36] br[36] wl[30] vdd gnd cell_6t
Xbit_r31_c36 bl[36] br[36] wl[31] vdd gnd cell_6t
Xbit_r32_c36 bl[36] br[36] wl[32] vdd gnd cell_6t
Xbit_r33_c36 bl[36] br[36] wl[33] vdd gnd cell_6t
Xbit_r34_c36 bl[36] br[36] wl[34] vdd gnd cell_6t
Xbit_r35_c36 bl[36] br[36] wl[35] vdd gnd cell_6t
Xbit_r36_c36 bl[36] br[36] wl[36] vdd gnd cell_6t
Xbit_r37_c36 bl[36] br[36] wl[37] vdd gnd cell_6t
Xbit_r38_c36 bl[36] br[36] wl[38] vdd gnd cell_6t
Xbit_r39_c36 bl[36] br[36] wl[39] vdd gnd cell_6t
Xbit_r40_c36 bl[36] br[36] wl[40] vdd gnd cell_6t
Xbit_r41_c36 bl[36] br[36] wl[41] vdd gnd cell_6t
Xbit_r42_c36 bl[36] br[36] wl[42] vdd gnd cell_6t
Xbit_r43_c36 bl[36] br[36] wl[43] vdd gnd cell_6t
Xbit_r44_c36 bl[36] br[36] wl[44] vdd gnd cell_6t
Xbit_r45_c36 bl[36] br[36] wl[45] vdd gnd cell_6t
Xbit_r46_c36 bl[36] br[36] wl[46] vdd gnd cell_6t
Xbit_r47_c36 bl[36] br[36] wl[47] vdd gnd cell_6t
Xbit_r48_c36 bl[36] br[36] wl[48] vdd gnd cell_6t
Xbit_r49_c36 bl[36] br[36] wl[49] vdd gnd cell_6t
Xbit_r50_c36 bl[36] br[36] wl[50] vdd gnd cell_6t
Xbit_r51_c36 bl[36] br[36] wl[51] vdd gnd cell_6t
Xbit_r52_c36 bl[36] br[36] wl[52] vdd gnd cell_6t
Xbit_r53_c36 bl[36] br[36] wl[53] vdd gnd cell_6t
Xbit_r54_c36 bl[36] br[36] wl[54] vdd gnd cell_6t
Xbit_r55_c36 bl[36] br[36] wl[55] vdd gnd cell_6t
Xbit_r56_c36 bl[36] br[36] wl[56] vdd gnd cell_6t
Xbit_r57_c36 bl[36] br[36] wl[57] vdd gnd cell_6t
Xbit_r58_c36 bl[36] br[36] wl[58] vdd gnd cell_6t
Xbit_r59_c36 bl[36] br[36] wl[59] vdd gnd cell_6t
Xbit_r60_c36 bl[36] br[36] wl[60] vdd gnd cell_6t
Xbit_r61_c36 bl[36] br[36] wl[61] vdd gnd cell_6t
Xbit_r62_c36 bl[36] br[36] wl[62] vdd gnd cell_6t
Xbit_r63_c36 bl[36] br[36] wl[63] vdd gnd cell_6t
Xbit_r64_c36 bl[36] br[36] wl[64] vdd gnd cell_6t
Xbit_r65_c36 bl[36] br[36] wl[65] vdd gnd cell_6t
Xbit_r66_c36 bl[36] br[36] wl[66] vdd gnd cell_6t
Xbit_r67_c36 bl[36] br[36] wl[67] vdd gnd cell_6t
Xbit_r68_c36 bl[36] br[36] wl[68] vdd gnd cell_6t
Xbit_r69_c36 bl[36] br[36] wl[69] vdd gnd cell_6t
Xbit_r70_c36 bl[36] br[36] wl[70] vdd gnd cell_6t
Xbit_r71_c36 bl[36] br[36] wl[71] vdd gnd cell_6t
Xbit_r72_c36 bl[36] br[36] wl[72] vdd gnd cell_6t
Xbit_r73_c36 bl[36] br[36] wl[73] vdd gnd cell_6t
Xbit_r74_c36 bl[36] br[36] wl[74] vdd gnd cell_6t
Xbit_r75_c36 bl[36] br[36] wl[75] vdd gnd cell_6t
Xbit_r76_c36 bl[36] br[36] wl[76] vdd gnd cell_6t
Xbit_r77_c36 bl[36] br[36] wl[77] vdd gnd cell_6t
Xbit_r78_c36 bl[36] br[36] wl[78] vdd gnd cell_6t
Xbit_r79_c36 bl[36] br[36] wl[79] vdd gnd cell_6t
Xbit_r80_c36 bl[36] br[36] wl[80] vdd gnd cell_6t
Xbit_r81_c36 bl[36] br[36] wl[81] vdd gnd cell_6t
Xbit_r82_c36 bl[36] br[36] wl[82] vdd gnd cell_6t
Xbit_r83_c36 bl[36] br[36] wl[83] vdd gnd cell_6t
Xbit_r84_c36 bl[36] br[36] wl[84] vdd gnd cell_6t
Xbit_r85_c36 bl[36] br[36] wl[85] vdd gnd cell_6t
Xbit_r86_c36 bl[36] br[36] wl[86] vdd gnd cell_6t
Xbit_r87_c36 bl[36] br[36] wl[87] vdd gnd cell_6t
Xbit_r88_c36 bl[36] br[36] wl[88] vdd gnd cell_6t
Xbit_r89_c36 bl[36] br[36] wl[89] vdd gnd cell_6t
Xbit_r90_c36 bl[36] br[36] wl[90] vdd gnd cell_6t
Xbit_r91_c36 bl[36] br[36] wl[91] vdd gnd cell_6t
Xbit_r92_c36 bl[36] br[36] wl[92] vdd gnd cell_6t
Xbit_r93_c36 bl[36] br[36] wl[93] vdd gnd cell_6t
Xbit_r94_c36 bl[36] br[36] wl[94] vdd gnd cell_6t
Xbit_r95_c36 bl[36] br[36] wl[95] vdd gnd cell_6t
Xbit_r96_c36 bl[36] br[36] wl[96] vdd gnd cell_6t
Xbit_r97_c36 bl[36] br[36] wl[97] vdd gnd cell_6t
Xbit_r98_c36 bl[36] br[36] wl[98] vdd gnd cell_6t
Xbit_r99_c36 bl[36] br[36] wl[99] vdd gnd cell_6t
Xbit_r100_c36 bl[36] br[36] wl[100] vdd gnd cell_6t
Xbit_r101_c36 bl[36] br[36] wl[101] vdd gnd cell_6t
Xbit_r102_c36 bl[36] br[36] wl[102] vdd gnd cell_6t
Xbit_r103_c36 bl[36] br[36] wl[103] vdd gnd cell_6t
Xbit_r104_c36 bl[36] br[36] wl[104] vdd gnd cell_6t
Xbit_r105_c36 bl[36] br[36] wl[105] vdd gnd cell_6t
Xbit_r106_c36 bl[36] br[36] wl[106] vdd gnd cell_6t
Xbit_r107_c36 bl[36] br[36] wl[107] vdd gnd cell_6t
Xbit_r108_c36 bl[36] br[36] wl[108] vdd gnd cell_6t
Xbit_r109_c36 bl[36] br[36] wl[109] vdd gnd cell_6t
Xbit_r110_c36 bl[36] br[36] wl[110] vdd gnd cell_6t
Xbit_r111_c36 bl[36] br[36] wl[111] vdd gnd cell_6t
Xbit_r112_c36 bl[36] br[36] wl[112] vdd gnd cell_6t
Xbit_r113_c36 bl[36] br[36] wl[113] vdd gnd cell_6t
Xbit_r114_c36 bl[36] br[36] wl[114] vdd gnd cell_6t
Xbit_r115_c36 bl[36] br[36] wl[115] vdd gnd cell_6t
Xbit_r116_c36 bl[36] br[36] wl[116] vdd gnd cell_6t
Xbit_r117_c36 bl[36] br[36] wl[117] vdd gnd cell_6t
Xbit_r118_c36 bl[36] br[36] wl[118] vdd gnd cell_6t
Xbit_r119_c36 bl[36] br[36] wl[119] vdd gnd cell_6t
Xbit_r120_c36 bl[36] br[36] wl[120] vdd gnd cell_6t
Xbit_r121_c36 bl[36] br[36] wl[121] vdd gnd cell_6t
Xbit_r122_c36 bl[36] br[36] wl[122] vdd gnd cell_6t
Xbit_r123_c36 bl[36] br[36] wl[123] vdd gnd cell_6t
Xbit_r124_c36 bl[36] br[36] wl[124] vdd gnd cell_6t
Xbit_r125_c36 bl[36] br[36] wl[125] vdd gnd cell_6t
Xbit_r126_c36 bl[36] br[36] wl[126] vdd gnd cell_6t
Xbit_r127_c36 bl[36] br[36] wl[127] vdd gnd cell_6t
Xbit_r128_c36 bl[36] br[36] wl[128] vdd gnd cell_6t
Xbit_r129_c36 bl[36] br[36] wl[129] vdd gnd cell_6t
Xbit_r130_c36 bl[36] br[36] wl[130] vdd gnd cell_6t
Xbit_r131_c36 bl[36] br[36] wl[131] vdd gnd cell_6t
Xbit_r132_c36 bl[36] br[36] wl[132] vdd gnd cell_6t
Xbit_r133_c36 bl[36] br[36] wl[133] vdd gnd cell_6t
Xbit_r134_c36 bl[36] br[36] wl[134] vdd gnd cell_6t
Xbit_r135_c36 bl[36] br[36] wl[135] vdd gnd cell_6t
Xbit_r136_c36 bl[36] br[36] wl[136] vdd gnd cell_6t
Xbit_r137_c36 bl[36] br[36] wl[137] vdd gnd cell_6t
Xbit_r138_c36 bl[36] br[36] wl[138] vdd gnd cell_6t
Xbit_r139_c36 bl[36] br[36] wl[139] vdd gnd cell_6t
Xbit_r140_c36 bl[36] br[36] wl[140] vdd gnd cell_6t
Xbit_r141_c36 bl[36] br[36] wl[141] vdd gnd cell_6t
Xbit_r142_c36 bl[36] br[36] wl[142] vdd gnd cell_6t
Xbit_r143_c36 bl[36] br[36] wl[143] vdd gnd cell_6t
Xbit_r144_c36 bl[36] br[36] wl[144] vdd gnd cell_6t
Xbit_r145_c36 bl[36] br[36] wl[145] vdd gnd cell_6t
Xbit_r146_c36 bl[36] br[36] wl[146] vdd gnd cell_6t
Xbit_r147_c36 bl[36] br[36] wl[147] vdd gnd cell_6t
Xbit_r148_c36 bl[36] br[36] wl[148] vdd gnd cell_6t
Xbit_r149_c36 bl[36] br[36] wl[149] vdd gnd cell_6t
Xbit_r150_c36 bl[36] br[36] wl[150] vdd gnd cell_6t
Xbit_r151_c36 bl[36] br[36] wl[151] vdd gnd cell_6t
Xbit_r152_c36 bl[36] br[36] wl[152] vdd gnd cell_6t
Xbit_r153_c36 bl[36] br[36] wl[153] vdd gnd cell_6t
Xbit_r154_c36 bl[36] br[36] wl[154] vdd gnd cell_6t
Xbit_r155_c36 bl[36] br[36] wl[155] vdd gnd cell_6t
Xbit_r156_c36 bl[36] br[36] wl[156] vdd gnd cell_6t
Xbit_r157_c36 bl[36] br[36] wl[157] vdd gnd cell_6t
Xbit_r158_c36 bl[36] br[36] wl[158] vdd gnd cell_6t
Xbit_r159_c36 bl[36] br[36] wl[159] vdd gnd cell_6t
Xbit_r160_c36 bl[36] br[36] wl[160] vdd gnd cell_6t
Xbit_r161_c36 bl[36] br[36] wl[161] vdd gnd cell_6t
Xbit_r162_c36 bl[36] br[36] wl[162] vdd gnd cell_6t
Xbit_r163_c36 bl[36] br[36] wl[163] vdd gnd cell_6t
Xbit_r164_c36 bl[36] br[36] wl[164] vdd gnd cell_6t
Xbit_r165_c36 bl[36] br[36] wl[165] vdd gnd cell_6t
Xbit_r166_c36 bl[36] br[36] wl[166] vdd gnd cell_6t
Xbit_r167_c36 bl[36] br[36] wl[167] vdd gnd cell_6t
Xbit_r168_c36 bl[36] br[36] wl[168] vdd gnd cell_6t
Xbit_r169_c36 bl[36] br[36] wl[169] vdd gnd cell_6t
Xbit_r170_c36 bl[36] br[36] wl[170] vdd gnd cell_6t
Xbit_r171_c36 bl[36] br[36] wl[171] vdd gnd cell_6t
Xbit_r172_c36 bl[36] br[36] wl[172] vdd gnd cell_6t
Xbit_r173_c36 bl[36] br[36] wl[173] vdd gnd cell_6t
Xbit_r174_c36 bl[36] br[36] wl[174] vdd gnd cell_6t
Xbit_r175_c36 bl[36] br[36] wl[175] vdd gnd cell_6t
Xbit_r176_c36 bl[36] br[36] wl[176] vdd gnd cell_6t
Xbit_r177_c36 bl[36] br[36] wl[177] vdd gnd cell_6t
Xbit_r178_c36 bl[36] br[36] wl[178] vdd gnd cell_6t
Xbit_r179_c36 bl[36] br[36] wl[179] vdd gnd cell_6t
Xbit_r180_c36 bl[36] br[36] wl[180] vdd gnd cell_6t
Xbit_r181_c36 bl[36] br[36] wl[181] vdd gnd cell_6t
Xbit_r182_c36 bl[36] br[36] wl[182] vdd gnd cell_6t
Xbit_r183_c36 bl[36] br[36] wl[183] vdd gnd cell_6t
Xbit_r184_c36 bl[36] br[36] wl[184] vdd gnd cell_6t
Xbit_r185_c36 bl[36] br[36] wl[185] vdd gnd cell_6t
Xbit_r186_c36 bl[36] br[36] wl[186] vdd gnd cell_6t
Xbit_r187_c36 bl[36] br[36] wl[187] vdd gnd cell_6t
Xbit_r188_c36 bl[36] br[36] wl[188] vdd gnd cell_6t
Xbit_r189_c36 bl[36] br[36] wl[189] vdd gnd cell_6t
Xbit_r190_c36 bl[36] br[36] wl[190] vdd gnd cell_6t
Xbit_r191_c36 bl[36] br[36] wl[191] vdd gnd cell_6t
Xbit_r192_c36 bl[36] br[36] wl[192] vdd gnd cell_6t
Xbit_r193_c36 bl[36] br[36] wl[193] vdd gnd cell_6t
Xbit_r194_c36 bl[36] br[36] wl[194] vdd gnd cell_6t
Xbit_r195_c36 bl[36] br[36] wl[195] vdd gnd cell_6t
Xbit_r196_c36 bl[36] br[36] wl[196] vdd gnd cell_6t
Xbit_r197_c36 bl[36] br[36] wl[197] vdd gnd cell_6t
Xbit_r198_c36 bl[36] br[36] wl[198] vdd gnd cell_6t
Xbit_r199_c36 bl[36] br[36] wl[199] vdd gnd cell_6t
Xbit_r200_c36 bl[36] br[36] wl[200] vdd gnd cell_6t
Xbit_r201_c36 bl[36] br[36] wl[201] vdd gnd cell_6t
Xbit_r202_c36 bl[36] br[36] wl[202] vdd gnd cell_6t
Xbit_r203_c36 bl[36] br[36] wl[203] vdd gnd cell_6t
Xbit_r204_c36 bl[36] br[36] wl[204] vdd gnd cell_6t
Xbit_r205_c36 bl[36] br[36] wl[205] vdd gnd cell_6t
Xbit_r206_c36 bl[36] br[36] wl[206] vdd gnd cell_6t
Xbit_r207_c36 bl[36] br[36] wl[207] vdd gnd cell_6t
Xbit_r208_c36 bl[36] br[36] wl[208] vdd gnd cell_6t
Xbit_r209_c36 bl[36] br[36] wl[209] vdd gnd cell_6t
Xbit_r210_c36 bl[36] br[36] wl[210] vdd gnd cell_6t
Xbit_r211_c36 bl[36] br[36] wl[211] vdd gnd cell_6t
Xbit_r212_c36 bl[36] br[36] wl[212] vdd gnd cell_6t
Xbit_r213_c36 bl[36] br[36] wl[213] vdd gnd cell_6t
Xbit_r214_c36 bl[36] br[36] wl[214] vdd gnd cell_6t
Xbit_r215_c36 bl[36] br[36] wl[215] vdd gnd cell_6t
Xbit_r216_c36 bl[36] br[36] wl[216] vdd gnd cell_6t
Xbit_r217_c36 bl[36] br[36] wl[217] vdd gnd cell_6t
Xbit_r218_c36 bl[36] br[36] wl[218] vdd gnd cell_6t
Xbit_r219_c36 bl[36] br[36] wl[219] vdd gnd cell_6t
Xbit_r220_c36 bl[36] br[36] wl[220] vdd gnd cell_6t
Xbit_r221_c36 bl[36] br[36] wl[221] vdd gnd cell_6t
Xbit_r222_c36 bl[36] br[36] wl[222] vdd gnd cell_6t
Xbit_r223_c36 bl[36] br[36] wl[223] vdd gnd cell_6t
Xbit_r224_c36 bl[36] br[36] wl[224] vdd gnd cell_6t
Xbit_r225_c36 bl[36] br[36] wl[225] vdd gnd cell_6t
Xbit_r226_c36 bl[36] br[36] wl[226] vdd gnd cell_6t
Xbit_r227_c36 bl[36] br[36] wl[227] vdd gnd cell_6t
Xbit_r228_c36 bl[36] br[36] wl[228] vdd gnd cell_6t
Xbit_r229_c36 bl[36] br[36] wl[229] vdd gnd cell_6t
Xbit_r230_c36 bl[36] br[36] wl[230] vdd gnd cell_6t
Xbit_r231_c36 bl[36] br[36] wl[231] vdd gnd cell_6t
Xbit_r232_c36 bl[36] br[36] wl[232] vdd gnd cell_6t
Xbit_r233_c36 bl[36] br[36] wl[233] vdd gnd cell_6t
Xbit_r234_c36 bl[36] br[36] wl[234] vdd gnd cell_6t
Xbit_r235_c36 bl[36] br[36] wl[235] vdd gnd cell_6t
Xbit_r236_c36 bl[36] br[36] wl[236] vdd gnd cell_6t
Xbit_r237_c36 bl[36] br[36] wl[237] vdd gnd cell_6t
Xbit_r238_c36 bl[36] br[36] wl[238] vdd gnd cell_6t
Xbit_r239_c36 bl[36] br[36] wl[239] vdd gnd cell_6t
Xbit_r240_c36 bl[36] br[36] wl[240] vdd gnd cell_6t
Xbit_r241_c36 bl[36] br[36] wl[241] vdd gnd cell_6t
Xbit_r242_c36 bl[36] br[36] wl[242] vdd gnd cell_6t
Xbit_r243_c36 bl[36] br[36] wl[243] vdd gnd cell_6t
Xbit_r244_c36 bl[36] br[36] wl[244] vdd gnd cell_6t
Xbit_r245_c36 bl[36] br[36] wl[245] vdd gnd cell_6t
Xbit_r246_c36 bl[36] br[36] wl[246] vdd gnd cell_6t
Xbit_r247_c36 bl[36] br[36] wl[247] vdd gnd cell_6t
Xbit_r248_c36 bl[36] br[36] wl[248] vdd gnd cell_6t
Xbit_r249_c36 bl[36] br[36] wl[249] vdd gnd cell_6t
Xbit_r250_c36 bl[36] br[36] wl[250] vdd gnd cell_6t
Xbit_r251_c36 bl[36] br[36] wl[251] vdd gnd cell_6t
Xbit_r252_c36 bl[36] br[36] wl[252] vdd gnd cell_6t
Xbit_r253_c36 bl[36] br[36] wl[253] vdd gnd cell_6t
Xbit_r254_c36 bl[36] br[36] wl[254] vdd gnd cell_6t
Xbit_r255_c36 bl[36] br[36] wl[255] vdd gnd cell_6t
Xbit_r0_c37 bl[37] br[37] wl[0] vdd gnd cell_6t
Xbit_r1_c37 bl[37] br[37] wl[1] vdd gnd cell_6t
Xbit_r2_c37 bl[37] br[37] wl[2] vdd gnd cell_6t
Xbit_r3_c37 bl[37] br[37] wl[3] vdd gnd cell_6t
Xbit_r4_c37 bl[37] br[37] wl[4] vdd gnd cell_6t
Xbit_r5_c37 bl[37] br[37] wl[5] vdd gnd cell_6t
Xbit_r6_c37 bl[37] br[37] wl[6] vdd gnd cell_6t
Xbit_r7_c37 bl[37] br[37] wl[7] vdd gnd cell_6t
Xbit_r8_c37 bl[37] br[37] wl[8] vdd gnd cell_6t
Xbit_r9_c37 bl[37] br[37] wl[9] vdd gnd cell_6t
Xbit_r10_c37 bl[37] br[37] wl[10] vdd gnd cell_6t
Xbit_r11_c37 bl[37] br[37] wl[11] vdd gnd cell_6t
Xbit_r12_c37 bl[37] br[37] wl[12] vdd gnd cell_6t
Xbit_r13_c37 bl[37] br[37] wl[13] vdd gnd cell_6t
Xbit_r14_c37 bl[37] br[37] wl[14] vdd gnd cell_6t
Xbit_r15_c37 bl[37] br[37] wl[15] vdd gnd cell_6t
Xbit_r16_c37 bl[37] br[37] wl[16] vdd gnd cell_6t
Xbit_r17_c37 bl[37] br[37] wl[17] vdd gnd cell_6t
Xbit_r18_c37 bl[37] br[37] wl[18] vdd gnd cell_6t
Xbit_r19_c37 bl[37] br[37] wl[19] vdd gnd cell_6t
Xbit_r20_c37 bl[37] br[37] wl[20] vdd gnd cell_6t
Xbit_r21_c37 bl[37] br[37] wl[21] vdd gnd cell_6t
Xbit_r22_c37 bl[37] br[37] wl[22] vdd gnd cell_6t
Xbit_r23_c37 bl[37] br[37] wl[23] vdd gnd cell_6t
Xbit_r24_c37 bl[37] br[37] wl[24] vdd gnd cell_6t
Xbit_r25_c37 bl[37] br[37] wl[25] vdd gnd cell_6t
Xbit_r26_c37 bl[37] br[37] wl[26] vdd gnd cell_6t
Xbit_r27_c37 bl[37] br[37] wl[27] vdd gnd cell_6t
Xbit_r28_c37 bl[37] br[37] wl[28] vdd gnd cell_6t
Xbit_r29_c37 bl[37] br[37] wl[29] vdd gnd cell_6t
Xbit_r30_c37 bl[37] br[37] wl[30] vdd gnd cell_6t
Xbit_r31_c37 bl[37] br[37] wl[31] vdd gnd cell_6t
Xbit_r32_c37 bl[37] br[37] wl[32] vdd gnd cell_6t
Xbit_r33_c37 bl[37] br[37] wl[33] vdd gnd cell_6t
Xbit_r34_c37 bl[37] br[37] wl[34] vdd gnd cell_6t
Xbit_r35_c37 bl[37] br[37] wl[35] vdd gnd cell_6t
Xbit_r36_c37 bl[37] br[37] wl[36] vdd gnd cell_6t
Xbit_r37_c37 bl[37] br[37] wl[37] vdd gnd cell_6t
Xbit_r38_c37 bl[37] br[37] wl[38] vdd gnd cell_6t
Xbit_r39_c37 bl[37] br[37] wl[39] vdd gnd cell_6t
Xbit_r40_c37 bl[37] br[37] wl[40] vdd gnd cell_6t
Xbit_r41_c37 bl[37] br[37] wl[41] vdd gnd cell_6t
Xbit_r42_c37 bl[37] br[37] wl[42] vdd gnd cell_6t
Xbit_r43_c37 bl[37] br[37] wl[43] vdd gnd cell_6t
Xbit_r44_c37 bl[37] br[37] wl[44] vdd gnd cell_6t
Xbit_r45_c37 bl[37] br[37] wl[45] vdd gnd cell_6t
Xbit_r46_c37 bl[37] br[37] wl[46] vdd gnd cell_6t
Xbit_r47_c37 bl[37] br[37] wl[47] vdd gnd cell_6t
Xbit_r48_c37 bl[37] br[37] wl[48] vdd gnd cell_6t
Xbit_r49_c37 bl[37] br[37] wl[49] vdd gnd cell_6t
Xbit_r50_c37 bl[37] br[37] wl[50] vdd gnd cell_6t
Xbit_r51_c37 bl[37] br[37] wl[51] vdd gnd cell_6t
Xbit_r52_c37 bl[37] br[37] wl[52] vdd gnd cell_6t
Xbit_r53_c37 bl[37] br[37] wl[53] vdd gnd cell_6t
Xbit_r54_c37 bl[37] br[37] wl[54] vdd gnd cell_6t
Xbit_r55_c37 bl[37] br[37] wl[55] vdd gnd cell_6t
Xbit_r56_c37 bl[37] br[37] wl[56] vdd gnd cell_6t
Xbit_r57_c37 bl[37] br[37] wl[57] vdd gnd cell_6t
Xbit_r58_c37 bl[37] br[37] wl[58] vdd gnd cell_6t
Xbit_r59_c37 bl[37] br[37] wl[59] vdd gnd cell_6t
Xbit_r60_c37 bl[37] br[37] wl[60] vdd gnd cell_6t
Xbit_r61_c37 bl[37] br[37] wl[61] vdd gnd cell_6t
Xbit_r62_c37 bl[37] br[37] wl[62] vdd gnd cell_6t
Xbit_r63_c37 bl[37] br[37] wl[63] vdd gnd cell_6t
Xbit_r64_c37 bl[37] br[37] wl[64] vdd gnd cell_6t
Xbit_r65_c37 bl[37] br[37] wl[65] vdd gnd cell_6t
Xbit_r66_c37 bl[37] br[37] wl[66] vdd gnd cell_6t
Xbit_r67_c37 bl[37] br[37] wl[67] vdd gnd cell_6t
Xbit_r68_c37 bl[37] br[37] wl[68] vdd gnd cell_6t
Xbit_r69_c37 bl[37] br[37] wl[69] vdd gnd cell_6t
Xbit_r70_c37 bl[37] br[37] wl[70] vdd gnd cell_6t
Xbit_r71_c37 bl[37] br[37] wl[71] vdd gnd cell_6t
Xbit_r72_c37 bl[37] br[37] wl[72] vdd gnd cell_6t
Xbit_r73_c37 bl[37] br[37] wl[73] vdd gnd cell_6t
Xbit_r74_c37 bl[37] br[37] wl[74] vdd gnd cell_6t
Xbit_r75_c37 bl[37] br[37] wl[75] vdd gnd cell_6t
Xbit_r76_c37 bl[37] br[37] wl[76] vdd gnd cell_6t
Xbit_r77_c37 bl[37] br[37] wl[77] vdd gnd cell_6t
Xbit_r78_c37 bl[37] br[37] wl[78] vdd gnd cell_6t
Xbit_r79_c37 bl[37] br[37] wl[79] vdd gnd cell_6t
Xbit_r80_c37 bl[37] br[37] wl[80] vdd gnd cell_6t
Xbit_r81_c37 bl[37] br[37] wl[81] vdd gnd cell_6t
Xbit_r82_c37 bl[37] br[37] wl[82] vdd gnd cell_6t
Xbit_r83_c37 bl[37] br[37] wl[83] vdd gnd cell_6t
Xbit_r84_c37 bl[37] br[37] wl[84] vdd gnd cell_6t
Xbit_r85_c37 bl[37] br[37] wl[85] vdd gnd cell_6t
Xbit_r86_c37 bl[37] br[37] wl[86] vdd gnd cell_6t
Xbit_r87_c37 bl[37] br[37] wl[87] vdd gnd cell_6t
Xbit_r88_c37 bl[37] br[37] wl[88] vdd gnd cell_6t
Xbit_r89_c37 bl[37] br[37] wl[89] vdd gnd cell_6t
Xbit_r90_c37 bl[37] br[37] wl[90] vdd gnd cell_6t
Xbit_r91_c37 bl[37] br[37] wl[91] vdd gnd cell_6t
Xbit_r92_c37 bl[37] br[37] wl[92] vdd gnd cell_6t
Xbit_r93_c37 bl[37] br[37] wl[93] vdd gnd cell_6t
Xbit_r94_c37 bl[37] br[37] wl[94] vdd gnd cell_6t
Xbit_r95_c37 bl[37] br[37] wl[95] vdd gnd cell_6t
Xbit_r96_c37 bl[37] br[37] wl[96] vdd gnd cell_6t
Xbit_r97_c37 bl[37] br[37] wl[97] vdd gnd cell_6t
Xbit_r98_c37 bl[37] br[37] wl[98] vdd gnd cell_6t
Xbit_r99_c37 bl[37] br[37] wl[99] vdd gnd cell_6t
Xbit_r100_c37 bl[37] br[37] wl[100] vdd gnd cell_6t
Xbit_r101_c37 bl[37] br[37] wl[101] vdd gnd cell_6t
Xbit_r102_c37 bl[37] br[37] wl[102] vdd gnd cell_6t
Xbit_r103_c37 bl[37] br[37] wl[103] vdd gnd cell_6t
Xbit_r104_c37 bl[37] br[37] wl[104] vdd gnd cell_6t
Xbit_r105_c37 bl[37] br[37] wl[105] vdd gnd cell_6t
Xbit_r106_c37 bl[37] br[37] wl[106] vdd gnd cell_6t
Xbit_r107_c37 bl[37] br[37] wl[107] vdd gnd cell_6t
Xbit_r108_c37 bl[37] br[37] wl[108] vdd gnd cell_6t
Xbit_r109_c37 bl[37] br[37] wl[109] vdd gnd cell_6t
Xbit_r110_c37 bl[37] br[37] wl[110] vdd gnd cell_6t
Xbit_r111_c37 bl[37] br[37] wl[111] vdd gnd cell_6t
Xbit_r112_c37 bl[37] br[37] wl[112] vdd gnd cell_6t
Xbit_r113_c37 bl[37] br[37] wl[113] vdd gnd cell_6t
Xbit_r114_c37 bl[37] br[37] wl[114] vdd gnd cell_6t
Xbit_r115_c37 bl[37] br[37] wl[115] vdd gnd cell_6t
Xbit_r116_c37 bl[37] br[37] wl[116] vdd gnd cell_6t
Xbit_r117_c37 bl[37] br[37] wl[117] vdd gnd cell_6t
Xbit_r118_c37 bl[37] br[37] wl[118] vdd gnd cell_6t
Xbit_r119_c37 bl[37] br[37] wl[119] vdd gnd cell_6t
Xbit_r120_c37 bl[37] br[37] wl[120] vdd gnd cell_6t
Xbit_r121_c37 bl[37] br[37] wl[121] vdd gnd cell_6t
Xbit_r122_c37 bl[37] br[37] wl[122] vdd gnd cell_6t
Xbit_r123_c37 bl[37] br[37] wl[123] vdd gnd cell_6t
Xbit_r124_c37 bl[37] br[37] wl[124] vdd gnd cell_6t
Xbit_r125_c37 bl[37] br[37] wl[125] vdd gnd cell_6t
Xbit_r126_c37 bl[37] br[37] wl[126] vdd gnd cell_6t
Xbit_r127_c37 bl[37] br[37] wl[127] vdd gnd cell_6t
Xbit_r128_c37 bl[37] br[37] wl[128] vdd gnd cell_6t
Xbit_r129_c37 bl[37] br[37] wl[129] vdd gnd cell_6t
Xbit_r130_c37 bl[37] br[37] wl[130] vdd gnd cell_6t
Xbit_r131_c37 bl[37] br[37] wl[131] vdd gnd cell_6t
Xbit_r132_c37 bl[37] br[37] wl[132] vdd gnd cell_6t
Xbit_r133_c37 bl[37] br[37] wl[133] vdd gnd cell_6t
Xbit_r134_c37 bl[37] br[37] wl[134] vdd gnd cell_6t
Xbit_r135_c37 bl[37] br[37] wl[135] vdd gnd cell_6t
Xbit_r136_c37 bl[37] br[37] wl[136] vdd gnd cell_6t
Xbit_r137_c37 bl[37] br[37] wl[137] vdd gnd cell_6t
Xbit_r138_c37 bl[37] br[37] wl[138] vdd gnd cell_6t
Xbit_r139_c37 bl[37] br[37] wl[139] vdd gnd cell_6t
Xbit_r140_c37 bl[37] br[37] wl[140] vdd gnd cell_6t
Xbit_r141_c37 bl[37] br[37] wl[141] vdd gnd cell_6t
Xbit_r142_c37 bl[37] br[37] wl[142] vdd gnd cell_6t
Xbit_r143_c37 bl[37] br[37] wl[143] vdd gnd cell_6t
Xbit_r144_c37 bl[37] br[37] wl[144] vdd gnd cell_6t
Xbit_r145_c37 bl[37] br[37] wl[145] vdd gnd cell_6t
Xbit_r146_c37 bl[37] br[37] wl[146] vdd gnd cell_6t
Xbit_r147_c37 bl[37] br[37] wl[147] vdd gnd cell_6t
Xbit_r148_c37 bl[37] br[37] wl[148] vdd gnd cell_6t
Xbit_r149_c37 bl[37] br[37] wl[149] vdd gnd cell_6t
Xbit_r150_c37 bl[37] br[37] wl[150] vdd gnd cell_6t
Xbit_r151_c37 bl[37] br[37] wl[151] vdd gnd cell_6t
Xbit_r152_c37 bl[37] br[37] wl[152] vdd gnd cell_6t
Xbit_r153_c37 bl[37] br[37] wl[153] vdd gnd cell_6t
Xbit_r154_c37 bl[37] br[37] wl[154] vdd gnd cell_6t
Xbit_r155_c37 bl[37] br[37] wl[155] vdd gnd cell_6t
Xbit_r156_c37 bl[37] br[37] wl[156] vdd gnd cell_6t
Xbit_r157_c37 bl[37] br[37] wl[157] vdd gnd cell_6t
Xbit_r158_c37 bl[37] br[37] wl[158] vdd gnd cell_6t
Xbit_r159_c37 bl[37] br[37] wl[159] vdd gnd cell_6t
Xbit_r160_c37 bl[37] br[37] wl[160] vdd gnd cell_6t
Xbit_r161_c37 bl[37] br[37] wl[161] vdd gnd cell_6t
Xbit_r162_c37 bl[37] br[37] wl[162] vdd gnd cell_6t
Xbit_r163_c37 bl[37] br[37] wl[163] vdd gnd cell_6t
Xbit_r164_c37 bl[37] br[37] wl[164] vdd gnd cell_6t
Xbit_r165_c37 bl[37] br[37] wl[165] vdd gnd cell_6t
Xbit_r166_c37 bl[37] br[37] wl[166] vdd gnd cell_6t
Xbit_r167_c37 bl[37] br[37] wl[167] vdd gnd cell_6t
Xbit_r168_c37 bl[37] br[37] wl[168] vdd gnd cell_6t
Xbit_r169_c37 bl[37] br[37] wl[169] vdd gnd cell_6t
Xbit_r170_c37 bl[37] br[37] wl[170] vdd gnd cell_6t
Xbit_r171_c37 bl[37] br[37] wl[171] vdd gnd cell_6t
Xbit_r172_c37 bl[37] br[37] wl[172] vdd gnd cell_6t
Xbit_r173_c37 bl[37] br[37] wl[173] vdd gnd cell_6t
Xbit_r174_c37 bl[37] br[37] wl[174] vdd gnd cell_6t
Xbit_r175_c37 bl[37] br[37] wl[175] vdd gnd cell_6t
Xbit_r176_c37 bl[37] br[37] wl[176] vdd gnd cell_6t
Xbit_r177_c37 bl[37] br[37] wl[177] vdd gnd cell_6t
Xbit_r178_c37 bl[37] br[37] wl[178] vdd gnd cell_6t
Xbit_r179_c37 bl[37] br[37] wl[179] vdd gnd cell_6t
Xbit_r180_c37 bl[37] br[37] wl[180] vdd gnd cell_6t
Xbit_r181_c37 bl[37] br[37] wl[181] vdd gnd cell_6t
Xbit_r182_c37 bl[37] br[37] wl[182] vdd gnd cell_6t
Xbit_r183_c37 bl[37] br[37] wl[183] vdd gnd cell_6t
Xbit_r184_c37 bl[37] br[37] wl[184] vdd gnd cell_6t
Xbit_r185_c37 bl[37] br[37] wl[185] vdd gnd cell_6t
Xbit_r186_c37 bl[37] br[37] wl[186] vdd gnd cell_6t
Xbit_r187_c37 bl[37] br[37] wl[187] vdd gnd cell_6t
Xbit_r188_c37 bl[37] br[37] wl[188] vdd gnd cell_6t
Xbit_r189_c37 bl[37] br[37] wl[189] vdd gnd cell_6t
Xbit_r190_c37 bl[37] br[37] wl[190] vdd gnd cell_6t
Xbit_r191_c37 bl[37] br[37] wl[191] vdd gnd cell_6t
Xbit_r192_c37 bl[37] br[37] wl[192] vdd gnd cell_6t
Xbit_r193_c37 bl[37] br[37] wl[193] vdd gnd cell_6t
Xbit_r194_c37 bl[37] br[37] wl[194] vdd gnd cell_6t
Xbit_r195_c37 bl[37] br[37] wl[195] vdd gnd cell_6t
Xbit_r196_c37 bl[37] br[37] wl[196] vdd gnd cell_6t
Xbit_r197_c37 bl[37] br[37] wl[197] vdd gnd cell_6t
Xbit_r198_c37 bl[37] br[37] wl[198] vdd gnd cell_6t
Xbit_r199_c37 bl[37] br[37] wl[199] vdd gnd cell_6t
Xbit_r200_c37 bl[37] br[37] wl[200] vdd gnd cell_6t
Xbit_r201_c37 bl[37] br[37] wl[201] vdd gnd cell_6t
Xbit_r202_c37 bl[37] br[37] wl[202] vdd gnd cell_6t
Xbit_r203_c37 bl[37] br[37] wl[203] vdd gnd cell_6t
Xbit_r204_c37 bl[37] br[37] wl[204] vdd gnd cell_6t
Xbit_r205_c37 bl[37] br[37] wl[205] vdd gnd cell_6t
Xbit_r206_c37 bl[37] br[37] wl[206] vdd gnd cell_6t
Xbit_r207_c37 bl[37] br[37] wl[207] vdd gnd cell_6t
Xbit_r208_c37 bl[37] br[37] wl[208] vdd gnd cell_6t
Xbit_r209_c37 bl[37] br[37] wl[209] vdd gnd cell_6t
Xbit_r210_c37 bl[37] br[37] wl[210] vdd gnd cell_6t
Xbit_r211_c37 bl[37] br[37] wl[211] vdd gnd cell_6t
Xbit_r212_c37 bl[37] br[37] wl[212] vdd gnd cell_6t
Xbit_r213_c37 bl[37] br[37] wl[213] vdd gnd cell_6t
Xbit_r214_c37 bl[37] br[37] wl[214] vdd gnd cell_6t
Xbit_r215_c37 bl[37] br[37] wl[215] vdd gnd cell_6t
Xbit_r216_c37 bl[37] br[37] wl[216] vdd gnd cell_6t
Xbit_r217_c37 bl[37] br[37] wl[217] vdd gnd cell_6t
Xbit_r218_c37 bl[37] br[37] wl[218] vdd gnd cell_6t
Xbit_r219_c37 bl[37] br[37] wl[219] vdd gnd cell_6t
Xbit_r220_c37 bl[37] br[37] wl[220] vdd gnd cell_6t
Xbit_r221_c37 bl[37] br[37] wl[221] vdd gnd cell_6t
Xbit_r222_c37 bl[37] br[37] wl[222] vdd gnd cell_6t
Xbit_r223_c37 bl[37] br[37] wl[223] vdd gnd cell_6t
Xbit_r224_c37 bl[37] br[37] wl[224] vdd gnd cell_6t
Xbit_r225_c37 bl[37] br[37] wl[225] vdd gnd cell_6t
Xbit_r226_c37 bl[37] br[37] wl[226] vdd gnd cell_6t
Xbit_r227_c37 bl[37] br[37] wl[227] vdd gnd cell_6t
Xbit_r228_c37 bl[37] br[37] wl[228] vdd gnd cell_6t
Xbit_r229_c37 bl[37] br[37] wl[229] vdd gnd cell_6t
Xbit_r230_c37 bl[37] br[37] wl[230] vdd gnd cell_6t
Xbit_r231_c37 bl[37] br[37] wl[231] vdd gnd cell_6t
Xbit_r232_c37 bl[37] br[37] wl[232] vdd gnd cell_6t
Xbit_r233_c37 bl[37] br[37] wl[233] vdd gnd cell_6t
Xbit_r234_c37 bl[37] br[37] wl[234] vdd gnd cell_6t
Xbit_r235_c37 bl[37] br[37] wl[235] vdd gnd cell_6t
Xbit_r236_c37 bl[37] br[37] wl[236] vdd gnd cell_6t
Xbit_r237_c37 bl[37] br[37] wl[237] vdd gnd cell_6t
Xbit_r238_c37 bl[37] br[37] wl[238] vdd gnd cell_6t
Xbit_r239_c37 bl[37] br[37] wl[239] vdd gnd cell_6t
Xbit_r240_c37 bl[37] br[37] wl[240] vdd gnd cell_6t
Xbit_r241_c37 bl[37] br[37] wl[241] vdd gnd cell_6t
Xbit_r242_c37 bl[37] br[37] wl[242] vdd gnd cell_6t
Xbit_r243_c37 bl[37] br[37] wl[243] vdd gnd cell_6t
Xbit_r244_c37 bl[37] br[37] wl[244] vdd gnd cell_6t
Xbit_r245_c37 bl[37] br[37] wl[245] vdd gnd cell_6t
Xbit_r246_c37 bl[37] br[37] wl[246] vdd gnd cell_6t
Xbit_r247_c37 bl[37] br[37] wl[247] vdd gnd cell_6t
Xbit_r248_c37 bl[37] br[37] wl[248] vdd gnd cell_6t
Xbit_r249_c37 bl[37] br[37] wl[249] vdd gnd cell_6t
Xbit_r250_c37 bl[37] br[37] wl[250] vdd gnd cell_6t
Xbit_r251_c37 bl[37] br[37] wl[251] vdd gnd cell_6t
Xbit_r252_c37 bl[37] br[37] wl[252] vdd gnd cell_6t
Xbit_r253_c37 bl[37] br[37] wl[253] vdd gnd cell_6t
Xbit_r254_c37 bl[37] br[37] wl[254] vdd gnd cell_6t
Xbit_r255_c37 bl[37] br[37] wl[255] vdd gnd cell_6t
Xbit_r0_c38 bl[38] br[38] wl[0] vdd gnd cell_6t
Xbit_r1_c38 bl[38] br[38] wl[1] vdd gnd cell_6t
Xbit_r2_c38 bl[38] br[38] wl[2] vdd gnd cell_6t
Xbit_r3_c38 bl[38] br[38] wl[3] vdd gnd cell_6t
Xbit_r4_c38 bl[38] br[38] wl[4] vdd gnd cell_6t
Xbit_r5_c38 bl[38] br[38] wl[5] vdd gnd cell_6t
Xbit_r6_c38 bl[38] br[38] wl[6] vdd gnd cell_6t
Xbit_r7_c38 bl[38] br[38] wl[7] vdd gnd cell_6t
Xbit_r8_c38 bl[38] br[38] wl[8] vdd gnd cell_6t
Xbit_r9_c38 bl[38] br[38] wl[9] vdd gnd cell_6t
Xbit_r10_c38 bl[38] br[38] wl[10] vdd gnd cell_6t
Xbit_r11_c38 bl[38] br[38] wl[11] vdd gnd cell_6t
Xbit_r12_c38 bl[38] br[38] wl[12] vdd gnd cell_6t
Xbit_r13_c38 bl[38] br[38] wl[13] vdd gnd cell_6t
Xbit_r14_c38 bl[38] br[38] wl[14] vdd gnd cell_6t
Xbit_r15_c38 bl[38] br[38] wl[15] vdd gnd cell_6t
Xbit_r16_c38 bl[38] br[38] wl[16] vdd gnd cell_6t
Xbit_r17_c38 bl[38] br[38] wl[17] vdd gnd cell_6t
Xbit_r18_c38 bl[38] br[38] wl[18] vdd gnd cell_6t
Xbit_r19_c38 bl[38] br[38] wl[19] vdd gnd cell_6t
Xbit_r20_c38 bl[38] br[38] wl[20] vdd gnd cell_6t
Xbit_r21_c38 bl[38] br[38] wl[21] vdd gnd cell_6t
Xbit_r22_c38 bl[38] br[38] wl[22] vdd gnd cell_6t
Xbit_r23_c38 bl[38] br[38] wl[23] vdd gnd cell_6t
Xbit_r24_c38 bl[38] br[38] wl[24] vdd gnd cell_6t
Xbit_r25_c38 bl[38] br[38] wl[25] vdd gnd cell_6t
Xbit_r26_c38 bl[38] br[38] wl[26] vdd gnd cell_6t
Xbit_r27_c38 bl[38] br[38] wl[27] vdd gnd cell_6t
Xbit_r28_c38 bl[38] br[38] wl[28] vdd gnd cell_6t
Xbit_r29_c38 bl[38] br[38] wl[29] vdd gnd cell_6t
Xbit_r30_c38 bl[38] br[38] wl[30] vdd gnd cell_6t
Xbit_r31_c38 bl[38] br[38] wl[31] vdd gnd cell_6t
Xbit_r32_c38 bl[38] br[38] wl[32] vdd gnd cell_6t
Xbit_r33_c38 bl[38] br[38] wl[33] vdd gnd cell_6t
Xbit_r34_c38 bl[38] br[38] wl[34] vdd gnd cell_6t
Xbit_r35_c38 bl[38] br[38] wl[35] vdd gnd cell_6t
Xbit_r36_c38 bl[38] br[38] wl[36] vdd gnd cell_6t
Xbit_r37_c38 bl[38] br[38] wl[37] vdd gnd cell_6t
Xbit_r38_c38 bl[38] br[38] wl[38] vdd gnd cell_6t
Xbit_r39_c38 bl[38] br[38] wl[39] vdd gnd cell_6t
Xbit_r40_c38 bl[38] br[38] wl[40] vdd gnd cell_6t
Xbit_r41_c38 bl[38] br[38] wl[41] vdd gnd cell_6t
Xbit_r42_c38 bl[38] br[38] wl[42] vdd gnd cell_6t
Xbit_r43_c38 bl[38] br[38] wl[43] vdd gnd cell_6t
Xbit_r44_c38 bl[38] br[38] wl[44] vdd gnd cell_6t
Xbit_r45_c38 bl[38] br[38] wl[45] vdd gnd cell_6t
Xbit_r46_c38 bl[38] br[38] wl[46] vdd gnd cell_6t
Xbit_r47_c38 bl[38] br[38] wl[47] vdd gnd cell_6t
Xbit_r48_c38 bl[38] br[38] wl[48] vdd gnd cell_6t
Xbit_r49_c38 bl[38] br[38] wl[49] vdd gnd cell_6t
Xbit_r50_c38 bl[38] br[38] wl[50] vdd gnd cell_6t
Xbit_r51_c38 bl[38] br[38] wl[51] vdd gnd cell_6t
Xbit_r52_c38 bl[38] br[38] wl[52] vdd gnd cell_6t
Xbit_r53_c38 bl[38] br[38] wl[53] vdd gnd cell_6t
Xbit_r54_c38 bl[38] br[38] wl[54] vdd gnd cell_6t
Xbit_r55_c38 bl[38] br[38] wl[55] vdd gnd cell_6t
Xbit_r56_c38 bl[38] br[38] wl[56] vdd gnd cell_6t
Xbit_r57_c38 bl[38] br[38] wl[57] vdd gnd cell_6t
Xbit_r58_c38 bl[38] br[38] wl[58] vdd gnd cell_6t
Xbit_r59_c38 bl[38] br[38] wl[59] vdd gnd cell_6t
Xbit_r60_c38 bl[38] br[38] wl[60] vdd gnd cell_6t
Xbit_r61_c38 bl[38] br[38] wl[61] vdd gnd cell_6t
Xbit_r62_c38 bl[38] br[38] wl[62] vdd gnd cell_6t
Xbit_r63_c38 bl[38] br[38] wl[63] vdd gnd cell_6t
Xbit_r64_c38 bl[38] br[38] wl[64] vdd gnd cell_6t
Xbit_r65_c38 bl[38] br[38] wl[65] vdd gnd cell_6t
Xbit_r66_c38 bl[38] br[38] wl[66] vdd gnd cell_6t
Xbit_r67_c38 bl[38] br[38] wl[67] vdd gnd cell_6t
Xbit_r68_c38 bl[38] br[38] wl[68] vdd gnd cell_6t
Xbit_r69_c38 bl[38] br[38] wl[69] vdd gnd cell_6t
Xbit_r70_c38 bl[38] br[38] wl[70] vdd gnd cell_6t
Xbit_r71_c38 bl[38] br[38] wl[71] vdd gnd cell_6t
Xbit_r72_c38 bl[38] br[38] wl[72] vdd gnd cell_6t
Xbit_r73_c38 bl[38] br[38] wl[73] vdd gnd cell_6t
Xbit_r74_c38 bl[38] br[38] wl[74] vdd gnd cell_6t
Xbit_r75_c38 bl[38] br[38] wl[75] vdd gnd cell_6t
Xbit_r76_c38 bl[38] br[38] wl[76] vdd gnd cell_6t
Xbit_r77_c38 bl[38] br[38] wl[77] vdd gnd cell_6t
Xbit_r78_c38 bl[38] br[38] wl[78] vdd gnd cell_6t
Xbit_r79_c38 bl[38] br[38] wl[79] vdd gnd cell_6t
Xbit_r80_c38 bl[38] br[38] wl[80] vdd gnd cell_6t
Xbit_r81_c38 bl[38] br[38] wl[81] vdd gnd cell_6t
Xbit_r82_c38 bl[38] br[38] wl[82] vdd gnd cell_6t
Xbit_r83_c38 bl[38] br[38] wl[83] vdd gnd cell_6t
Xbit_r84_c38 bl[38] br[38] wl[84] vdd gnd cell_6t
Xbit_r85_c38 bl[38] br[38] wl[85] vdd gnd cell_6t
Xbit_r86_c38 bl[38] br[38] wl[86] vdd gnd cell_6t
Xbit_r87_c38 bl[38] br[38] wl[87] vdd gnd cell_6t
Xbit_r88_c38 bl[38] br[38] wl[88] vdd gnd cell_6t
Xbit_r89_c38 bl[38] br[38] wl[89] vdd gnd cell_6t
Xbit_r90_c38 bl[38] br[38] wl[90] vdd gnd cell_6t
Xbit_r91_c38 bl[38] br[38] wl[91] vdd gnd cell_6t
Xbit_r92_c38 bl[38] br[38] wl[92] vdd gnd cell_6t
Xbit_r93_c38 bl[38] br[38] wl[93] vdd gnd cell_6t
Xbit_r94_c38 bl[38] br[38] wl[94] vdd gnd cell_6t
Xbit_r95_c38 bl[38] br[38] wl[95] vdd gnd cell_6t
Xbit_r96_c38 bl[38] br[38] wl[96] vdd gnd cell_6t
Xbit_r97_c38 bl[38] br[38] wl[97] vdd gnd cell_6t
Xbit_r98_c38 bl[38] br[38] wl[98] vdd gnd cell_6t
Xbit_r99_c38 bl[38] br[38] wl[99] vdd gnd cell_6t
Xbit_r100_c38 bl[38] br[38] wl[100] vdd gnd cell_6t
Xbit_r101_c38 bl[38] br[38] wl[101] vdd gnd cell_6t
Xbit_r102_c38 bl[38] br[38] wl[102] vdd gnd cell_6t
Xbit_r103_c38 bl[38] br[38] wl[103] vdd gnd cell_6t
Xbit_r104_c38 bl[38] br[38] wl[104] vdd gnd cell_6t
Xbit_r105_c38 bl[38] br[38] wl[105] vdd gnd cell_6t
Xbit_r106_c38 bl[38] br[38] wl[106] vdd gnd cell_6t
Xbit_r107_c38 bl[38] br[38] wl[107] vdd gnd cell_6t
Xbit_r108_c38 bl[38] br[38] wl[108] vdd gnd cell_6t
Xbit_r109_c38 bl[38] br[38] wl[109] vdd gnd cell_6t
Xbit_r110_c38 bl[38] br[38] wl[110] vdd gnd cell_6t
Xbit_r111_c38 bl[38] br[38] wl[111] vdd gnd cell_6t
Xbit_r112_c38 bl[38] br[38] wl[112] vdd gnd cell_6t
Xbit_r113_c38 bl[38] br[38] wl[113] vdd gnd cell_6t
Xbit_r114_c38 bl[38] br[38] wl[114] vdd gnd cell_6t
Xbit_r115_c38 bl[38] br[38] wl[115] vdd gnd cell_6t
Xbit_r116_c38 bl[38] br[38] wl[116] vdd gnd cell_6t
Xbit_r117_c38 bl[38] br[38] wl[117] vdd gnd cell_6t
Xbit_r118_c38 bl[38] br[38] wl[118] vdd gnd cell_6t
Xbit_r119_c38 bl[38] br[38] wl[119] vdd gnd cell_6t
Xbit_r120_c38 bl[38] br[38] wl[120] vdd gnd cell_6t
Xbit_r121_c38 bl[38] br[38] wl[121] vdd gnd cell_6t
Xbit_r122_c38 bl[38] br[38] wl[122] vdd gnd cell_6t
Xbit_r123_c38 bl[38] br[38] wl[123] vdd gnd cell_6t
Xbit_r124_c38 bl[38] br[38] wl[124] vdd gnd cell_6t
Xbit_r125_c38 bl[38] br[38] wl[125] vdd gnd cell_6t
Xbit_r126_c38 bl[38] br[38] wl[126] vdd gnd cell_6t
Xbit_r127_c38 bl[38] br[38] wl[127] vdd gnd cell_6t
Xbit_r128_c38 bl[38] br[38] wl[128] vdd gnd cell_6t
Xbit_r129_c38 bl[38] br[38] wl[129] vdd gnd cell_6t
Xbit_r130_c38 bl[38] br[38] wl[130] vdd gnd cell_6t
Xbit_r131_c38 bl[38] br[38] wl[131] vdd gnd cell_6t
Xbit_r132_c38 bl[38] br[38] wl[132] vdd gnd cell_6t
Xbit_r133_c38 bl[38] br[38] wl[133] vdd gnd cell_6t
Xbit_r134_c38 bl[38] br[38] wl[134] vdd gnd cell_6t
Xbit_r135_c38 bl[38] br[38] wl[135] vdd gnd cell_6t
Xbit_r136_c38 bl[38] br[38] wl[136] vdd gnd cell_6t
Xbit_r137_c38 bl[38] br[38] wl[137] vdd gnd cell_6t
Xbit_r138_c38 bl[38] br[38] wl[138] vdd gnd cell_6t
Xbit_r139_c38 bl[38] br[38] wl[139] vdd gnd cell_6t
Xbit_r140_c38 bl[38] br[38] wl[140] vdd gnd cell_6t
Xbit_r141_c38 bl[38] br[38] wl[141] vdd gnd cell_6t
Xbit_r142_c38 bl[38] br[38] wl[142] vdd gnd cell_6t
Xbit_r143_c38 bl[38] br[38] wl[143] vdd gnd cell_6t
Xbit_r144_c38 bl[38] br[38] wl[144] vdd gnd cell_6t
Xbit_r145_c38 bl[38] br[38] wl[145] vdd gnd cell_6t
Xbit_r146_c38 bl[38] br[38] wl[146] vdd gnd cell_6t
Xbit_r147_c38 bl[38] br[38] wl[147] vdd gnd cell_6t
Xbit_r148_c38 bl[38] br[38] wl[148] vdd gnd cell_6t
Xbit_r149_c38 bl[38] br[38] wl[149] vdd gnd cell_6t
Xbit_r150_c38 bl[38] br[38] wl[150] vdd gnd cell_6t
Xbit_r151_c38 bl[38] br[38] wl[151] vdd gnd cell_6t
Xbit_r152_c38 bl[38] br[38] wl[152] vdd gnd cell_6t
Xbit_r153_c38 bl[38] br[38] wl[153] vdd gnd cell_6t
Xbit_r154_c38 bl[38] br[38] wl[154] vdd gnd cell_6t
Xbit_r155_c38 bl[38] br[38] wl[155] vdd gnd cell_6t
Xbit_r156_c38 bl[38] br[38] wl[156] vdd gnd cell_6t
Xbit_r157_c38 bl[38] br[38] wl[157] vdd gnd cell_6t
Xbit_r158_c38 bl[38] br[38] wl[158] vdd gnd cell_6t
Xbit_r159_c38 bl[38] br[38] wl[159] vdd gnd cell_6t
Xbit_r160_c38 bl[38] br[38] wl[160] vdd gnd cell_6t
Xbit_r161_c38 bl[38] br[38] wl[161] vdd gnd cell_6t
Xbit_r162_c38 bl[38] br[38] wl[162] vdd gnd cell_6t
Xbit_r163_c38 bl[38] br[38] wl[163] vdd gnd cell_6t
Xbit_r164_c38 bl[38] br[38] wl[164] vdd gnd cell_6t
Xbit_r165_c38 bl[38] br[38] wl[165] vdd gnd cell_6t
Xbit_r166_c38 bl[38] br[38] wl[166] vdd gnd cell_6t
Xbit_r167_c38 bl[38] br[38] wl[167] vdd gnd cell_6t
Xbit_r168_c38 bl[38] br[38] wl[168] vdd gnd cell_6t
Xbit_r169_c38 bl[38] br[38] wl[169] vdd gnd cell_6t
Xbit_r170_c38 bl[38] br[38] wl[170] vdd gnd cell_6t
Xbit_r171_c38 bl[38] br[38] wl[171] vdd gnd cell_6t
Xbit_r172_c38 bl[38] br[38] wl[172] vdd gnd cell_6t
Xbit_r173_c38 bl[38] br[38] wl[173] vdd gnd cell_6t
Xbit_r174_c38 bl[38] br[38] wl[174] vdd gnd cell_6t
Xbit_r175_c38 bl[38] br[38] wl[175] vdd gnd cell_6t
Xbit_r176_c38 bl[38] br[38] wl[176] vdd gnd cell_6t
Xbit_r177_c38 bl[38] br[38] wl[177] vdd gnd cell_6t
Xbit_r178_c38 bl[38] br[38] wl[178] vdd gnd cell_6t
Xbit_r179_c38 bl[38] br[38] wl[179] vdd gnd cell_6t
Xbit_r180_c38 bl[38] br[38] wl[180] vdd gnd cell_6t
Xbit_r181_c38 bl[38] br[38] wl[181] vdd gnd cell_6t
Xbit_r182_c38 bl[38] br[38] wl[182] vdd gnd cell_6t
Xbit_r183_c38 bl[38] br[38] wl[183] vdd gnd cell_6t
Xbit_r184_c38 bl[38] br[38] wl[184] vdd gnd cell_6t
Xbit_r185_c38 bl[38] br[38] wl[185] vdd gnd cell_6t
Xbit_r186_c38 bl[38] br[38] wl[186] vdd gnd cell_6t
Xbit_r187_c38 bl[38] br[38] wl[187] vdd gnd cell_6t
Xbit_r188_c38 bl[38] br[38] wl[188] vdd gnd cell_6t
Xbit_r189_c38 bl[38] br[38] wl[189] vdd gnd cell_6t
Xbit_r190_c38 bl[38] br[38] wl[190] vdd gnd cell_6t
Xbit_r191_c38 bl[38] br[38] wl[191] vdd gnd cell_6t
Xbit_r192_c38 bl[38] br[38] wl[192] vdd gnd cell_6t
Xbit_r193_c38 bl[38] br[38] wl[193] vdd gnd cell_6t
Xbit_r194_c38 bl[38] br[38] wl[194] vdd gnd cell_6t
Xbit_r195_c38 bl[38] br[38] wl[195] vdd gnd cell_6t
Xbit_r196_c38 bl[38] br[38] wl[196] vdd gnd cell_6t
Xbit_r197_c38 bl[38] br[38] wl[197] vdd gnd cell_6t
Xbit_r198_c38 bl[38] br[38] wl[198] vdd gnd cell_6t
Xbit_r199_c38 bl[38] br[38] wl[199] vdd gnd cell_6t
Xbit_r200_c38 bl[38] br[38] wl[200] vdd gnd cell_6t
Xbit_r201_c38 bl[38] br[38] wl[201] vdd gnd cell_6t
Xbit_r202_c38 bl[38] br[38] wl[202] vdd gnd cell_6t
Xbit_r203_c38 bl[38] br[38] wl[203] vdd gnd cell_6t
Xbit_r204_c38 bl[38] br[38] wl[204] vdd gnd cell_6t
Xbit_r205_c38 bl[38] br[38] wl[205] vdd gnd cell_6t
Xbit_r206_c38 bl[38] br[38] wl[206] vdd gnd cell_6t
Xbit_r207_c38 bl[38] br[38] wl[207] vdd gnd cell_6t
Xbit_r208_c38 bl[38] br[38] wl[208] vdd gnd cell_6t
Xbit_r209_c38 bl[38] br[38] wl[209] vdd gnd cell_6t
Xbit_r210_c38 bl[38] br[38] wl[210] vdd gnd cell_6t
Xbit_r211_c38 bl[38] br[38] wl[211] vdd gnd cell_6t
Xbit_r212_c38 bl[38] br[38] wl[212] vdd gnd cell_6t
Xbit_r213_c38 bl[38] br[38] wl[213] vdd gnd cell_6t
Xbit_r214_c38 bl[38] br[38] wl[214] vdd gnd cell_6t
Xbit_r215_c38 bl[38] br[38] wl[215] vdd gnd cell_6t
Xbit_r216_c38 bl[38] br[38] wl[216] vdd gnd cell_6t
Xbit_r217_c38 bl[38] br[38] wl[217] vdd gnd cell_6t
Xbit_r218_c38 bl[38] br[38] wl[218] vdd gnd cell_6t
Xbit_r219_c38 bl[38] br[38] wl[219] vdd gnd cell_6t
Xbit_r220_c38 bl[38] br[38] wl[220] vdd gnd cell_6t
Xbit_r221_c38 bl[38] br[38] wl[221] vdd gnd cell_6t
Xbit_r222_c38 bl[38] br[38] wl[222] vdd gnd cell_6t
Xbit_r223_c38 bl[38] br[38] wl[223] vdd gnd cell_6t
Xbit_r224_c38 bl[38] br[38] wl[224] vdd gnd cell_6t
Xbit_r225_c38 bl[38] br[38] wl[225] vdd gnd cell_6t
Xbit_r226_c38 bl[38] br[38] wl[226] vdd gnd cell_6t
Xbit_r227_c38 bl[38] br[38] wl[227] vdd gnd cell_6t
Xbit_r228_c38 bl[38] br[38] wl[228] vdd gnd cell_6t
Xbit_r229_c38 bl[38] br[38] wl[229] vdd gnd cell_6t
Xbit_r230_c38 bl[38] br[38] wl[230] vdd gnd cell_6t
Xbit_r231_c38 bl[38] br[38] wl[231] vdd gnd cell_6t
Xbit_r232_c38 bl[38] br[38] wl[232] vdd gnd cell_6t
Xbit_r233_c38 bl[38] br[38] wl[233] vdd gnd cell_6t
Xbit_r234_c38 bl[38] br[38] wl[234] vdd gnd cell_6t
Xbit_r235_c38 bl[38] br[38] wl[235] vdd gnd cell_6t
Xbit_r236_c38 bl[38] br[38] wl[236] vdd gnd cell_6t
Xbit_r237_c38 bl[38] br[38] wl[237] vdd gnd cell_6t
Xbit_r238_c38 bl[38] br[38] wl[238] vdd gnd cell_6t
Xbit_r239_c38 bl[38] br[38] wl[239] vdd gnd cell_6t
Xbit_r240_c38 bl[38] br[38] wl[240] vdd gnd cell_6t
Xbit_r241_c38 bl[38] br[38] wl[241] vdd gnd cell_6t
Xbit_r242_c38 bl[38] br[38] wl[242] vdd gnd cell_6t
Xbit_r243_c38 bl[38] br[38] wl[243] vdd gnd cell_6t
Xbit_r244_c38 bl[38] br[38] wl[244] vdd gnd cell_6t
Xbit_r245_c38 bl[38] br[38] wl[245] vdd gnd cell_6t
Xbit_r246_c38 bl[38] br[38] wl[246] vdd gnd cell_6t
Xbit_r247_c38 bl[38] br[38] wl[247] vdd gnd cell_6t
Xbit_r248_c38 bl[38] br[38] wl[248] vdd gnd cell_6t
Xbit_r249_c38 bl[38] br[38] wl[249] vdd gnd cell_6t
Xbit_r250_c38 bl[38] br[38] wl[250] vdd gnd cell_6t
Xbit_r251_c38 bl[38] br[38] wl[251] vdd gnd cell_6t
Xbit_r252_c38 bl[38] br[38] wl[252] vdd gnd cell_6t
Xbit_r253_c38 bl[38] br[38] wl[253] vdd gnd cell_6t
Xbit_r254_c38 bl[38] br[38] wl[254] vdd gnd cell_6t
Xbit_r255_c38 bl[38] br[38] wl[255] vdd gnd cell_6t
Xbit_r0_c39 bl[39] br[39] wl[0] vdd gnd cell_6t
Xbit_r1_c39 bl[39] br[39] wl[1] vdd gnd cell_6t
Xbit_r2_c39 bl[39] br[39] wl[2] vdd gnd cell_6t
Xbit_r3_c39 bl[39] br[39] wl[3] vdd gnd cell_6t
Xbit_r4_c39 bl[39] br[39] wl[4] vdd gnd cell_6t
Xbit_r5_c39 bl[39] br[39] wl[5] vdd gnd cell_6t
Xbit_r6_c39 bl[39] br[39] wl[6] vdd gnd cell_6t
Xbit_r7_c39 bl[39] br[39] wl[7] vdd gnd cell_6t
Xbit_r8_c39 bl[39] br[39] wl[8] vdd gnd cell_6t
Xbit_r9_c39 bl[39] br[39] wl[9] vdd gnd cell_6t
Xbit_r10_c39 bl[39] br[39] wl[10] vdd gnd cell_6t
Xbit_r11_c39 bl[39] br[39] wl[11] vdd gnd cell_6t
Xbit_r12_c39 bl[39] br[39] wl[12] vdd gnd cell_6t
Xbit_r13_c39 bl[39] br[39] wl[13] vdd gnd cell_6t
Xbit_r14_c39 bl[39] br[39] wl[14] vdd gnd cell_6t
Xbit_r15_c39 bl[39] br[39] wl[15] vdd gnd cell_6t
Xbit_r16_c39 bl[39] br[39] wl[16] vdd gnd cell_6t
Xbit_r17_c39 bl[39] br[39] wl[17] vdd gnd cell_6t
Xbit_r18_c39 bl[39] br[39] wl[18] vdd gnd cell_6t
Xbit_r19_c39 bl[39] br[39] wl[19] vdd gnd cell_6t
Xbit_r20_c39 bl[39] br[39] wl[20] vdd gnd cell_6t
Xbit_r21_c39 bl[39] br[39] wl[21] vdd gnd cell_6t
Xbit_r22_c39 bl[39] br[39] wl[22] vdd gnd cell_6t
Xbit_r23_c39 bl[39] br[39] wl[23] vdd gnd cell_6t
Xbit_r24_c39 bl[39] br[39] wl[24] vdd gnd cell_6t
Xbit_r25_c39 bl[39] br[39] wl[25] vdd gnd cell_6t
Xbit_r26_c39 bl[39] br[39] wl[26] vdd gnd cell_6t
Xbit_r27_c39 bl[39] br[39] wl[27] vdd gnd cell_6t
Xbit_r28_c39 bl[39] br[39] wl[28] vdd gnd cell_6t
Xbit_r29_c39 bl[39] br[39] wl[29] vdd gnd cell_6t
Xbit_r30_c39 bl[39] br[39] wl[30] vdd gnd cell_6t
Xbit_r31_c39 bl[39] br[39] wl[31] vdd gnd cell_6t
Xbit_r32_c39 bl[39] br[39] wl[32] vdd gnd cell_6t
Xbit_r33_c39 bl[39] br[39] wl[33] vdd gnd cell_6t
Xbit_r34_c39 bl[39] br[39] wl[34] vdd gnd cell_6t
Xbit_r35_c39 bl[39] br[39] wl[35] vdd gnd cell_6t
Xbit_r36_c39 bl[39] br[39] wl[36] vdd gnd cell_6t
Xbit_r37_c39 bl[39] br[39] wl[37] vdd gnd cell_6t
Xbit_r38_c39 bl[39] br[39] wl[38] vdd gnd cell_6t
Xbit_r39_c39 bl[39] br[39] wl[39] vdd gnd cell_6t
Xbit_r40_c39 bl[39] br[39] wl[40] vdd gnd cell_6t
Xbit_r41_c39 bl[39] br[39] wl[41] vdd gnd cell_6t
Xbit_r42_c39 bl[39] br[39] wl[42] vdd gnd cell_6t
Xbit_r43_c39 bl[39] br[39] wl[43] vdd gnd cell_6t
Xbit_r44_c39 bl[39] br[39] wl[44] vdd gnd cell_6t
Xbit_r45_c39 bl[39] br[39] wl[45] vdd gnd cell_6t
Xbit_r46_c39 bl[39] br[39] wl[46] vdd gnd cell_6t
Xbit_r47_c39 bl[39] br[39] wl[47] vdd gnd cell_6t
Xbit_r48_c39 bl[39] br[39] wl[48] vdd gnd cell_6t
Xbit_r49_c39 bl[39] br[39] wl[49] vdd gnd cell_6t
Xbit_r50_c39 bl[39] br[39] wl[50] vdd gnd cell_6t
Xbit_r51_c39 bl[39] br[39] wl[51] vdd gnd cell_6t
Xbit_r52_c39 bl[39] br[39] wl[52] vdd gnd cell_6t
Xbit_r53_c39 bl[39] br[39] wl[53] vdd gnd cell_6t
Xbit_r54_c39 bl[39] br[39] wl[54] vdd gnd cell_6t
Xbit_r55_c39 bl[39] br[39] wl[55] vdd gnd cell_6t
Xbit_r56_c39 bl[39] br[39] wl[56] vdd gnd cell_6t
Xbit_r57_c39 bl[39] br[39] wl[57] vdd gnd cell_6t
Xbit_r58_c39 bl[39] br[39] wl[58] vdd gnd cell_6t
Xbit_r59_c39 bl[39] br[39] wl[59] vdd gnd cell_6t
Xbit_r60_c39 bl[39] br[39] wl[60] vdd gnd cell_6t
Xbit_r61_c39 bl[39] br[39] wl[61] vdd gnd cell_6t
Xbit_r62_c39 bl[39] br[39] wl[62] vdd gnd cell_6t
Xbit_r63_c39 bl[39] br[39] wl[63] vdd gnd cell_6t
Xbit_r64_c39 bl[39] br[39] wl[64] vdd gnd cell_6t
Xbit_r65_c39 bl[39] br[39] wl[65] vdd gnd cell_6t
Xbit_r66_c39 bl[39] br[39] wl[66] vdd gnd cell_6t
Xbit_r67_c39 bl[39] br[39] wl[67] vdd gnd cell_6t
Xbit_r68_c39 bl[39] br[39] wl[68] vdd gnd cell_6t
Xbit_r69_c39 bl[39] br[39] wl[69] vdd gnd cell_6t
Xbit_r70_c39 bl[39] br[39] wl[70] vdd gnd cell_6t
Xbit_r71_c39 bl[39] br[39] wl[71] vdd gnd cell_6t
Xbit_r72_c39 bl[39] br[39] wl[72] vdd gnd cell_6t
Xbit_r73_c39 bl[39] br[39] wl[73] vdd gnd cell_6t
Xbit_r74_c39 bl[39] br[39] wl[74] vdd gnd cell_6t
Xbit_r75_c39 bl[39] br[39] wl[75] vdd gnd cell_6t
Xbit_r76_c39 bl[39] br[39] wl[76] vdd gnd cell_6t
Xbit_r77_c39 bl[39] br[39] wl[77] vdd gnd cell_6t
Xbit_r78_c39 bl[39] br[39] wl[78] vdd gnd cell_6t
Xbit_r79_c39 bl[39] br[39] wl[79] vdd gnd cell_6t
Xbit_r80_c39 bl[39] br[39] wl[80] vdd gnd cell_6t
Xbit_r81_c39 bl[39] br[39] wl[81] vdd gnd cell_6t
Xbit_r82_c39 bl[39] br[39] wl[82] vdd gnd cell_6t
Xbit_r83_c39 bl[39] br[39] wl[83] vdd gnd cell_6t
Xbit_r84_c39 bl[39] br[39] wl[84] vdd gnd cell_6t
Xbit_r85_c39 bl[39] br[39] wl[85] vdd gnd cell_6t
Xbit_r86_c39 bl[39] br[39] wl[86] vdd gnd cell_6t
Xbit_r87_c39 bl[39] br[39] wl[87] vdd gnd cell_6t
Xbit_r88_c39 bl[39] br[39] wl[88] vdd gnd cell_6t
Xbit_r89_c39 bl[39] br[39] wl[89] vdd gnd cell_6t
Xbit_r90_c39 bl[39] br[39] wl[90] vdd gnd cell_6t
Xbit_r91_c39 bl[39] br[39] wl[91] vdd gnd cell_6t
Xbit_r92_c39 bl[39] br[39] wl[92] vdd gnd cell_6t
Xbit_r93_c39 bl[39] br[39] wl[93] vdd gnd cell_6t
Xbit_r94_c39 bl[39] br[39] wl[94] vdd gnd cell_6t
Xbit_r95_c39 bl[39] br[39] wl[95] vdd gnd cell_6t
Xbit_r96_c39 bl[39] br[39] wl[96] vdd gnd cell_6t
Xbit_r97_c39 bl[39] br[39] wl[97] vdd gnd cell_6t
Xbit_r98_c39 bl[39] br[39] wl[98] vdd gnd cell_6t
Xbit_r99_c39 bl[39] br[39] wl[99] vdd gnd cell_6t
Xbit_r100_c39 bl[39] br[39] wl[100] vdd gnd cell_6t
Xbit_r101_c39 bl[39] br[39] wl[101] vdd gnd cell_6t
Xbit_r102_c39 bl[39] br[39] wl[102] vdd gnd cell_6t
Xbit_r103_c39 bl[39] br[39] wl[103] vdd gnd cell_6t
Xbit_r104_c39 bl[39] br[39] wl[104] vdd gnd cell_6t
Xbit_r105_c39 bl[39] br[39] wl[105] vdd gnd cell_6t
Xbit_r106_c39 bl[39] br[39] wl[106] vdd gnd cell_6t
Xbit_r107_c39 bl[39] br[39] wl[107] vdd gnd cell_6t
Xbit_r108_c39 bl[39] br[39] wl[108] vdd gnd cell_6t
Xbit_r109_c39 bl[39] br[39] wl[109] vdd gnd cell_6t
Xbit_r110_c39 bl[39] br[39] wl[110] vdd gnd cell_6t
Xbit_r111_c39 bl[39] br[39] wl[111] vdd gnd cell_6t
Xbit_r112_c39 bl[39] br[39] wl[112] vdd gnd cell_6t
Xbit_r113_c39 bl[39] br[39] wl[113] vdd gnd cell_6t
Xbit_r114_c39 bl[39] br[39] wl[114] vdd gnd cell_6t
Xbit_r115_c39 bl[39] br[39] wl[115] vdd gnd cell_6t
Xbit_r116_c39 bl[39] br[39] wl[116] vdd gnd cell_6t
Xbit_r117_c39 bl[39] br[39] wl[117] vdd gnd cell_6t
Xbit_r118_c39 bl[39] br[39] wl[118] vdd gnd cell_6t
Xbit_r119_c39 bl[39] br[39] wl[119] vdd gnd cell_6t
Xbit_r120_c39 bl[39] br[39] wl[120] vdd gnd cell_6t
Xbit_r121_c39 bl[39] br[39] wl[121] vdd gnd cell_6t
Xbit_r122_c39 bl[39] br[39] wl[122] vdd gnd cell_6t
Xbit_r123_c39 bl[39] br[39] wl[123] vdd gnd cell_6t
Xbit_r124_c39 bl[39] br[39] wl[124] vdd gnd cell_6t
Xbit_r125_c39 bl[39] br[39] wl[125] vdd gnd cell_6t
Xbit_r126_c39 bl[39] br[39] wl[126] vdd gnd cell_6t
Xbit_r127_c39 bl[39] br[39] wl[127] vdd gnd cell_6t
Xbit_r128_c39 bl[39] br[39] wl[128] vdd gnd cell_6t
Xbit_r129_c39 bl[39] br[39] wl[129] vdd gnd cell_6t
Xbit_r130_c39 bl[39] br[39] wl[130] vdd gnd cell_6t
Xbit_r131_c39 bl[39] br[39] wl[131] vdd gnd cell_6t
Xbit_r132_c39 bl[39] br[39] wl[132] vdd gnd cell_6t
Xbit_r133_c39 bl[39] br[39] wl[133] vdd gnd cell_6t
Xbit_r134_c39 bl[39] br[39] wl[134] vdd gnd cell_6t
Xbit_r135_c39 bl[39] br[39] wl[135] vdd gnd cell_6t
Xbit_r136_c39 bl[39] br[39] wl[136] vdd gnd cell_6t
Xbit_r137_c39 bl[39] br[39] wl[137] vdd gnd cell_6t
Xbit_r138_c39 bl[39] br[39] wl[138] vdd gnd cell_6t
Xbit_r139_c39 bl[39] br[39] wl[139] vdd gnd cell_6t
Xbit_r140_c39 bl[39] br[39] wl[140] vdd gnd cell_6t
Xbit_r141_c39 bl[39] br[39] wl[141] vdd gnd cell_6t
Xbit_r142_c39 bl[39] br[39] wl[142] vdd gnd cell_6t
Xbit_r143_c39 bl[39] br[39] wl[143] vdd gnd cell_6t
Xbit_r144_c39 bl[39] br[39] wl[144] vdd gnd cell_6t
Xbit_r145_c39 bl[39] br[39] wl[145] vdd gnd cell_6t
Xbit_r146_c39 bl[39] br[39] wl[146] vdd gnd cell_6t
Xbit_r147_c39 bl[39] br[39] wl[147] vdd gnd cell_6t
Xbit_r148_c39 bl[39] br[39] wl[148] vdd gnd cell_6t
Xbit_r149_c39 bl[39] br[39] wl[149] vdd gnd cell_6t
Xbit_r150_c39 bl[39] br[39] wl[150] vdd gnd cell_6t
Xbit_r151_c39 bl[39] br[39] wl[151] vdd gnd cell_6t
Xbit_r152_c39 bl[39] br[39] wl[152] vdd gnd cell_6t
Xbit_r153_c39 bl[39] br[39] wl[153] vdd gnd cell_6t
Xbit_r154_c39 bl[39] br[39] wl[154] vdd gnd cell_6t
Xbit_r155_c39 bl[39] br[39] wl[155] vdd gnd cell_6t
Xbit_r156_c39 bl[39] br[39] wl[156] vdd gnd cell_6t
Xbit_r157_c39 bl[39] br[39] wl[157] vdd gnd cell_6t
Xbit_r158_c39 bl[39] br[39] wl[158] vdd gnd cell_6t
Xbit_r159_c39 bl[39] br[39] wl[159] vdd gnd cell_6t
Xbit_r160_c39 bl[39] br[39] wl[160] vdd gnd cell_6t
Xbit_r161_c39 bl[39] br[39] wl[161] vdd gnd cell_6t
Xbit_r162_c39 bl[39] br[39] wl[162] vdd gnd cell_6t
Xbit_r163_c39 bl[39] br[39] wl[163] vdd gnd cell_6t
Xbit_r164_c39 bl[39] br[39] wl[164] vdd gnd cell_6t
Xbit_r165_c39 bl[39] br[39] wl[165] vdd gnd cell_6t
Xbit_r166_c39 bl[39] br[39] wl[166] vdd gnd cell_6t
Xbit_r167_c39 bl[39] br[39] wl[167] vdd gnd cell_6t
Xbit_r168_c39 bl[39] br[39] wl[168] vdd gnd cell_6t
Xbit_r169_c39 bl[39] br[39] wl[169] vdd gnd cell_6t
Xbit_r170_c39 bl[39] br[39] wl[170] vdd gnd cell_6t
Xbit_r171_c39 bl[39] br[39] wl[171] vdd gnd cell_6t
Xbit_r172_c39 bl[39] br[39] wl[172] vdd gnd cell_6t
Xbit_r173_c39 bl[39] br[39] wl[173] vdd gnd cell_6t
Xbit_r174_c39 bl[39] br[39] wl[174] vdd gnd cell_6t
Xbit_r175_c39 bl[39] br[39] wl[175] vdd gnd cell_6t
Xbit_r176_c39 bl[39] br[39] wl[176] vdd gnd cell_6t
Xbit_r177_c39 bl[39] br[39] wl[177] vdd gnd cell_6t
Xbit_r178_c39 bl[39] br[39] wl[178] vdd gnd cell_6t
Xbit_r179_c39 bl[39] br[39] wl[179] vdd gnd cell_6t
Xbit_r180_c39 bl[39] br[39] wl[180] vdd gnd cell_6t
Xbit_r181_c39 bl[39] br[39] wl[181] vdd gnd cell_6t
Xbit_r182_c39 bl[39] br[39] wl[182] vdd gnd cell_6t
Xbit_r183_c39 bl[39] br[39] wl[183] vdd gnd cell_6t
Xbit_r184_c39 bl[39] br[39] wl[184] vdd gnd cell_6t
Xbit_r185_c39 bl[39] br[39] wl[185] vdd gnd cell_6t
Xbit_r186_c39 bl[39] br[39] wl[186] vdd gnd cell_6t
Xbit_r187_c39 bl[39] br[39] wl[187] vdd gnd cell_6t
Xbit_r188_c39 bl[39] br[39] wl[188] vdd gnd cell_6t
Xbit_r189_c39 bl[39] br[39] wl[189] vdd gnd cell_6t
Xbit_r190_c39 bl[39] br[39] wl[190] vdd gnd cell_6t
Xbit_r191_c39 bl[39] br[39] wl[191] vdd gnd cell_6t
Xbit_r192_c39 bl[39] br[39] wl[192] vdd gnd cell_6t
Xbit_r193_c39 bl[39] br[39] wl[193] vdd gnd cell_6t
Xbit_r194_c39 bl[39] br[39] wl[194] vdd gnd cell_6t
Xbit_r195_c39 bl[39] br[39] wl[195] vdd gnd cell_6t
Xbit_r196_c39 bl[39] br[39] wl[196] vdd gnd cell_6t
Xbit_r197_c39 bl[39] br[39] wl[197] vdd gnd cell_6t
Xbit_r198_c39 bl[39] br[39] wl[198] vdd gnd cell_6t
Xbit_r199_c39 bl[39] br[39] wl[199] vdd gnd cell_6t
Xbit_r200_c39 bl[39] br[39] wl[200] vdd gnd cell_6t
Xbit_r201_c39 bl[39] br[39] wl[201] vdd gnd cell_6t
Xbit_r202_c39 bl[39] br[39] wl[202] vdd gnd cell_6t
Xbit_r203_c39 bl[39] br[39] wl[203] vdd gnd cell_6t
Xbit_r204_c39 bl[39] br[39] wl[204] vdd gnd cell_6t
Xbit_r205_c39 bl[39] br[39] wl[205] vdd gnd cell_6t
Xbit_r206_c39 bl[39] br[39] wl[206] vdd gnd cell_6t
Xbit_r207_c39 bl[39] br[39] wl[207] vdd gnd cell_6t
Xbit_r208_c39 bl[39] br[39] wl[208] vdd gnd cell_6t
Xbit_r209_c39 bl[39] br[39] wl[209] vdd gnd cell_6t
Xbit_r210_c39 bl[39] br[39] wl[210] vdd gnd cell_6t
Xbit_r211_c39 bl[39] br[39] wl[211] vdd gnd cell_6t
Xbit_r212_c39 bl[39] br[39] wl[212] vdd gnd cell_6t
Xbit_r213_c39 bl[39] br[39] wl[213] vdd gnd cell_6t
Xbit_r214_c39 bl[39] br[39] wl[214] vdd gnd cell_6t
Xbit_r215_c39 bl[39] br[39] wl[215] vdd gnd cell_6t
Xbit_r216_c39 bl[39] br[39] wl[216] vdd gnd cell_6t
Xbit_r217_c39 bl[39] br[39] wl[217] vdd gnd cell_6t
Xbit_r218_c39 bl[39] br[39] wl[218] vdd gnd cell_6t
Xbit_r219_c39 bl[39] br[39] wl[219] vdd gnd cell_6t
Xbit_r220_c39 bl[39] br[39] wl[220] vdd gnd cell_6t
Xbit_r221_c39 bl[39] br[39] wl[221] vdd gnd cell_6t
Xbit_r222_c39 bl[39] br[39] wl[222] vdd gnd cell_6t
Xbit_r223_c39 bl[39] br[39] wl[223] vdd gnd cell_6t
Xbit_r224_c39 bl[39] br[39] wl[224] vdd gnd cell_6t
Xbit_r225_c39 bl[39] br[39] wl[225] vdd gnd cell_6t
Xbit_r226_c39 bl[39] br[39] wl[226] vdd gnd cell_6t
Xbit_r227_c39 bl[39] br[39] wl[227] vdd gnd cell_6t
Xbit_r228_c39 bl[39] br[39] wl[228] vdd gnd cell_6t
Xbit_r229_c39 bl[39] br[39] wl[229] vdd gnd cell_6t
Xbit_r230_c39 bl[39] br[39] wl[230] vdd gnd cell_6t
Xbit_r231_c39 bl[39] br[39] wl[231] vdd gnd cell_6t
Xbit_r232_c39 bl[39] br[39] wl[232] vdd gnd cell_6t
Xbit_r233_c39 bl[39] br[39] wl[233] vdd gnd cell_6t
Xbit_r234_c39 bl[39] br[39] wl[234] vdd gnd cell_6t
Xbit_r235_c39 bl[39] br[39] wl[235] vdd gnd cell_6t
Xbit_r236_c39 bl[39] br[39] wl[236] vdd gnd cell_6t
Xbit_r237_c39 bl[39] br[39] wl[237] vdd gnd cell_6t
Xbit_r238_c39 bl[39] br[39] wl[238] vdd gnd cell_6t
Xbit_r239_c39 bl[39] br[39] wl[239] vdd gnd cell_6t
Xbit_r240_c39 bl[39] br[39] wl[240] vdd gnd cell_6t
Xbit_r241_c39 bl[39] br[39] wl[241] vdd gnd cell_6t
Xbit_r242_c39 bl[39] br[39] wl[242] vdd gnd cell_6t
Xbit_r243_c39 bl[39] br[39] wl[243] vdd gnd cell_6t
Xbit_r244_c39 bl[39] br[39] wl[244] vdd gnd cell_6t
Xbit_r245_c39 bl[39] br[39] wl[245] vdd gnd cell_6t
Xbit_r246_c39 bl[39] br[39] wl[246] vdd gnd cell_6t
Xbit_r247_c39 bl[39] br[39] wl[247] vdd gnd cell_6t
Xbit_r248_c39 bl[39] br[39] wl[248] vdd gnd cell_6t
Xbit_r249_c39 bl[39] br[39] wl[249] vdd gnd cell_6t
Xbit_r250_c39 bl[39] br[39] wl[250] vdd gnd cell_6t
Xbit_r251_c39 bl[39] br[39] wl[251] vdd gnd cell_6t
Xbit_r252_c39 bl[39] br[39] wl[252] vdd gnd cell_6t
Xbit_r253_c39 bl[39] br[39] wl[253] vdd gnd cell_6t
Xbit_r254_c39 bl[39] br[39] wl[254] vdd gnd cell_6t
Xbit_r255_c39 bl[39] br[39] wl[255] vdd gnd cell_6t
Xbit_r0_c40 bl[40] br[40] wl[0] vdd gnd cell_6t
Xbit_r1_c40 bl[40] br[40] wl[1] vdd gnd cell_6t
Xbit_r2_c40 bl[40] br[40] wl[2] vdd gnd cell_6t
Xbit_r3_c40 bl[40] br[40] wl[3] vdd gnd cell_6t
Xbit_r4_c40 bl[40] br[40] wl[4] vdd gnd cell_6t
Xbit_r5_c40 bl[40] br[40] wl[5] vdd gnd cell_6t
Xbit_r6_c40 bl[40] br[40] wl[6] vdd gnd cell_6t
Xbit_r7_c40 bl[40] br[40] wl[7] vdd gnd cell_6t
Xbit_r8_c40 bl[40] br[40] wl[8] vdd gnd cell_6t
Xbit_r9_c40 bl[40] br[40] wl[9] vdd gnd cell_6t
Xbit_r10_c40 bl[40] br[40] wl[10] vdd gnd cell_6t
Xbit_r11_c40 bl[40] br[40] wl[11] vdd gnd cell_6t
Xbit_r12_c40 bl[40] br[40] wl[12] vdd gnd cell_6t
Xbit_r13_c40 bl[40] br[40] wl[13] vdd gnd cell_6t
Xbit_r14_c40 bl[40] br[40] wl[14] vdd gnd cell_6t
Xbit_r15_c40 bl[40] br[40] wl[15] vdd gnd cell_6t
Xbit_r16_c40 bl[40] br[40] wl[16] vdd gnd cell_6t
Xbit_r17_c40 bl[40] br[40] wl[17] vdd gnd cell_6t
Xbit_r18_c40 bl[40] br[40] wl[18] vdd gnd cell_6t
Xbit_r19_c40 bl[40] br[40] wl[19] vdd gnd cell_6t
Xbit_r20_c40 bl[40] br[40] wl[20] vdd gnd cell_6t
Xbit_r21_c40 bl[40] br[40] wl[21] vdd gnd cell_6t
Xbit_r22_c40 bl[40] br[40] wl[22] vdd gnd cell_6t
Xbit_r23_c40 bl[40] br[40] wl[23] vdd gnd cell_6t
Xbit_r24_c40 bl[40] br[40] wl[24] vdd gnd cell_6t
Xbit_r25_c40 bl[40] br[40] wl[25] vdd gnd cell_6t
Xbit_r26_c40 bl[40] br[40] wl[26] vdd gnd cell_6t
Xbit_r27_c40 bl[40] br[40] wl[27] vdd gnd cell_6t
Xbit_r28_c40 bl[40] br[40] wl[28] vdd gnd cell_6t
Xbit_r29_c40 bl[40] br[40] wl[29] vdd gnd cell_6t
Xbit_r30_c40 bl[40] br[40] wl[30] vdd gnd cell_6t
Xbit_r31_c40 bl[40] br[40] wl[31] vdd gnd cell_6t
Xbit_r32_c40 bl[40] br[40] wl[32] vdd gnd cell_6t
Xbit_r33_c40 bl[40] br[40] wl[33] vdd gnd cell_6t
Xbit_r34_c40 bl[40] br[40] wl[34] vdd gnd cell_6t
Xbit_r35_c40 bl[40] br[40] wl[35] vdd gnd cell_6t
Xbit_r36_c40 bl[40] br[40] wl[36] vdd gnd cell_6t
Xbit_r37_c40 bl[40] br[40] wl[37] vdd gnd cell_6t
Xbit_r38_c40 bl[40] br[40] wl[38] vdd gnd cell_6t
Xbit_r39_c40 bl[40] br[40] wl[39] vdd gnd cell_6t
Xbit_r40_c40 bl[40] br[40] wl[40] vdd gnd cell_6t
Xbit_r41_c40 bl[40] br[40] wl[41] vdd gnd cell_6t
Xbit_r42_c40 bl[40] br[40] wl[42] vdd gnd cell_6t
Xbit_r43_c40 bl[40] br[40] wl[43] vdd gnd cell_6t
Xbit_r44_c40 bl[40] br[40] wl[44] vdd gnd cell_6t
Xbit_r45_c40 bl[40] br[40] wl[45] vdd gnd cell_6t
Xbit_r46_c40 bl[40] br[40] wl[46] vdd gnd cell_6t
Xbit_r47_c40 bl[40] br[40] wl[47] vdd gnd cell_6t
Xbit_r48_c40 bl[40] br[40] wl[48] vdd gnd cell_6t
Xbit_r49_c40 bl[40] br[40] wl[49] vdd gnd cell_6t
Xbit_r50_c40 bl[40] br[40] wl[50] vdd gnd cell_6t
Xbit_r51_c40 bl[40] br[40] wl[51] vdd gnd cell_6t
Xbit_r52_c40 bl[40] br[40] wl[52] vdd gnd cell_6t
Xbit_r53_c40 bl[40] br[40] wl[53] vdd gnd cell_6t
Xbit_r54_c40 bl[40] br[40] wl[54] vdd gnd cell_6t
Xbit_r55_c40 bl[40] br[40] wl[55] vdd gnd cell_6t
Xbit_r56_c40 bl[40] br[40] wl[56] vdd gnd cell_6t
Xbit_r57_c40 bl[40] br[40] wl[57] vdd gnd cell_6t
Xbit_r58_c40 bl[40] br[40] wl[58] vdd gnd cell_6t
Xbit_r59_c40 bl[40] br[40] wl[59] vdd gnd cell_6t
Xbit_r60_c40 bl[40] br[40] wl[60] vdd gnd cell_6t
Xbit_r61_c40 bl[40] br[40] wl[61] vdd gnd cell_6t
Xbit_r62_c40 bl[40] br[40] wl[62] vdd gnd cell_6t
Xbit_r63_c40 bl[40] br[40] wl[63] vdd gnd cell_6t
Xbit_r64_c40 bl[40] br[40] wl[64] vdd gnd cell_6t
Xbit_r65_c40 bl[40] br[40] wl[65] vdd gnd cell_6t
Xbit_r66_c40 bl[40] br[40] wl[66] vdd gnd cell_6t
Xbit_r67_c40 bl[40] br[40] wl[67] vdd gnd cell_6t
Xbit_r68_c40 bl[40] br[40] wl[68] vdd gnd cell_6t
Xbit_r69_c40 bl[40] br[40] wl[69] vdd gnd cell_6t
Xbit_r70_c40 bl[40] br[40] wl[70] vdd gnd cell_6t
Xbit_r71_c40 bl[40] br[40] wl[71] vdd gnd cell_6t
Xbit_r72_c40 bl[40] br[40] wl[72] vdd gnd cell_6t
Xbit_r73_c40 bl[40] br[40] wl[73] vdd gnd cell_6t
Xbit_r74_c40 bl[40] br[40] wl[74] vdd gnd cell_6t
Xbit_r75_c40 bl[40] br[40] wl[75] vdd gnd cell_6t
Xbit_r76_c40 bl[40] br[40] wl[76] vdd gnd cell_6t
Xbit_r77_c40 bl[40] br[40] wl[77] vdd gnd cell_6t
Xbit_r78_c40 bl[40] br[40] wl[78] vdd gnd cell_6t
Xbit_r79_c40 bl[40] br[40] wl[79] vdd gnd cell_6t
Xbit_r80_c40 bl[40] br[40] wl[80] vdd gnd cell_6t
Xbit_r81_c40 bl[40] br[40] wl[81] vdd gnd cell_6t
Xbit_r82_c40 bl[40] br[40] wl[82] vdd gnd cell_6t
Xbit_r83_c40 bl[40] br[40] wl[83] vdd gnd cell_6t
Xbit_r84_c40 bl[40] br[40] wl[84] vdd gnd cell_6t
Xbit_r85_c40 bl[40] br[40] wl[85] vdd gnd cell_6t
Xbit_r86_c40 bl[40] br[40] wl[86] vdd gnd cell_6t
Xbit_r87_c40 bl[40] br[40] wl[87] vdd gnd cell_6t
Xbit_r88_c40 bl[40] br[40] wl[88] vdd gnd cell_6t
Xbit_r89_c40 bl[40] br[40] wl[89] vdd gnd cell_6t
Xbit_r90_c40 bl[40] br[40] wl[90] vdd gnd cell_6t
Xbit_r91_c40 bl[40] br[40] wl[91] vdd gnd cell_6t
Xbit_r92_c40 bl[40] br[40] wl[92] vdd gnd cell_6t
Xbit_r93_c40 bl[40] br[40] wl[93] vdd gnd cell_6t
Xbit_r94_c40 bl[40] br[40] wl[94] vdd gnd cell_6t
Xbit_r95_c40 bl[40] br[40] wl[95] vdd gnd cell_6t
Xbit_r96_c40 bl[40] br[40] wl[96] vdd gnd cell_6t
Xbit_r97_c40 bl[40] br[40] wl[97] vdd gnd cell_6t
Xbit_r98_c40 bl[40] br[40] wl[98] vdd gnd cell_6t
Xbit_r99_c40 bl[40] br[40] wl[99] vdd gnd cell_6t
Xbit_r100_c40 bl[40] br[40] wl[100] vdd gnd cell_6t
Xbit_r101_c40 bl[40] br[40] wl[101] vdd gnd cell_6t
Xbit_r102_c40 bl[40] br[40] wl[102] vdd gnd cell_6t
Xbit_r103_c40 bl[40] br[40] wl[103] vdd gnd cell_6t
Xbit_r104_c40 bl[40] br[40] wl[104] vdd gnd cell_6t
Xbit_r105_c40 bl[40] br[40] wl[105] vdd gnd cell_6t
Xbit_r106_c40 bl[40] br[40] wl[106] vdd gnd cell_6t
Xbit_r107_c40 bl[40] br[40] wl[107] vdd gnd cell_6t
Xbit_r108_c40 bl[40] br[40] wl[108] vdd gnd cell_6t
Xbit_r109_c40 bl[40] br[40] wl[109] vdd gnd cell_6t
Xbit_r110_c40 bl[40] br[40] wl[110] vdd gnd cell_6t
Xbit_r111_c40 bl[40] br[40] wl[111] vdd gnd cell_6t
Xbit_r112_c40 bl[40] br[40] wl[112] vdd gnd cell_6t
Xbit_r113_c40 bl[40] br[40] wl[113] vdd gnd cell_6t
Xbit_r114_c40 bl[40] br[40] wl[114] vdd gnd cell_6t
Xbit_r115_c40 bl[40] br[40] wl[115] vdd gnd cell_6t
Xbit_r116_c40 bl[40] br[40] wl[116] vdd gnd cell_6t
Xbit_r117_c40 bl[40] br[40] wl[117] vdd gnd cell_6t
Xbit_r118_c40 bl[40] br[40] wl[118] vdd gnd cell_6t
Xbit_r119_c40 bl[40] br[40] wl[119] vdd gnd cell_6t
Xbit_r120_c40 bl[40] br[40] wl[120] vdd gnd cell_6t
Xbit_r121_c40 bl[40] br[40] wl[121] vdd gnd cell_6t
Xbit_r122_c40 bl[40] br[40] wl[122] vdd gnd cell_6t
Xbit_r123_c40 bl[40] br[40] wl[123] vdd gnd cell_6t
Xbit_r124_c40 bl[40] br[40] wl[124] vdd gnd cell_6t
Xbit_r125_c40 bl[40] br[40] wl[125] vdd gnd cell_6t
Xbit_r126_c40 bl[40] br[40] wl[126] vdd gnd cell_6t
Xbit_r127_c40 bl[40] br[40] wl[127] vdd gnd cell_6t
Xbit_r128_c40 bl[40] br[40] wl[128] vdd gnd cell_6t
Xbit_r129_c40 bl[40] br[40] wl[129] vdd gnd cell_6t
Xbit_r130_c40 bl[40] br[40] wl[130] vdd gnd cell_6t
Xbit_r131_c40 bl[40] br[40] wl[131] vdd gnd cell_6t
Xbit_r132_c40 bl[40] br[40] wl[132] vdd gnd cell_6t
Xbit_r133_c40 bl[40] br[40] wl[133] vdd gnd cell_6t
Xbit_r134_c40 bl[40] br[40] wl[134] vdd gnd cell_6t
Xbit_r135_c40 bl[40] br[40] wl[135] vdd gnd cell_6t
Xbit_r136_c40 bl[40] br[40] wl[136] vdd gnd cell_6t
Xbit_r137_c40 bl[40] br[40] wl[137] vdd gnd cell_6t
Xbit_r138_c40 bl[40] br[40] wl[138] vdd gnd cell_6t
Xbit_r139_c40 bl[40] br[40] wl[139] vdd gnd cell_6t
Xbit_r140_c40 bl[40] br[40] wl[140] vdd gnd cell_6t
Xbit_r141_c40 bl[40] br[40] wl[141] vdd gnd cell_6t
Xbit_r142_c40 bl[40] br[40] wl[142] vdd gnd cell_6t
Xbit_r143_c40 bl[40] br[40] wl[143] vdd gnd cell_6t
Xbit_r144_c40 bl[40] br[40] wl[144] vdd gnd cell_6t
Xbit_r145_c40 bl[40] br[40] wl[145] vdd gnd cell_6t
Xbit_r146_c40 bl[40] br[40] wl[146] vdd gnd cell_6t
Xbit_r147_c40 bl[40] br[40] wl[147] vdd gnd cell_6t
Xbit_r148_c40 bl[40] br[40] wl[148] vdd gnd cell_6t
Xbit_r149_c40 bl[40] br[40] wl[149] vdd gnd cell_6t
Xbit_r150_c40 bl[40] br[40] wl[150] vdd gnd cell_6t
Xbit_r151_c40 bl[40] br[40] wl[151] vdd gnd cell_6t
Xbit_r152_c40 bl[40] br[40] wl[152] vdd gnd cell_6t
Xbit_r153_c40 bl[40] br[40] wl[153] vdd gnd cell_6t
Xbit_r154_c40 bl[40] br[40] wl[154] vdd gnd cell_6t
Xbit_r155_c40 bl[40] br[40] wl[155] vdd gnd cell_6t
Xbit_r156_c40 bl[40] br[40] wl[156] vdd gnd cell_6t
Xbit_r157_c40 bl[40] br[40] wl[157] vdd gnd cell_6t
Xbit_r158_c40 bl[40] br[40] wl[158] vdd gnd cell_6t
Xbit_r159_c40 bl[40] br[40] wl[159] vdd gnd cell_6t
Xbit_r160_c40 bl[40] br[40] wl[160] vdd gnd cell_6t
Xbit_r161_c40 bl[40] br[40] wl[161] vdd gnd cell_6t
Xbit_r162_c40 bl[40] br[40] wl[162] vdd gnd cell_6t
Xbit_r163_c40 bl[40] br[40] wl[163] vdd gnd cell_6t
Xbit_r164_c40 bl[40] br[40] wl[164] vdd gnd cell_6t
Xbit_r165_c40 bl[40] br[40] wl[165] vdd gnd cell_6t
Xbit_r166_c40 bl[40] br[40] wl[166] vdd gnd cell_6t
Xbit_r167_c40 bl[40] br[40] wl[167] vdd gnd cell_6t
Xbit_r168_c40 bl[40] br[40] wl[168] vdd gnd cell_6t
Xbit_r169_c40 bl[40] br[40] wl[169] vdd gnd cell_6t
Xbit_r170_c40 bl[40] br[40] wl[170] vdd gnd cell_6t
Xbit_r171_c40 bl[40] br[40] wl[171] vdd gnd cell_6t
Xbit_r172_c40 bl[40] br[40] wl[172] vdd gnd cell_6t
Xbit_r173_c40 bl[40] br[40] wl[173] vdd gnd cell_6t
Xbit_r174_c40 bl[40] br[40] wl[174] vdd gnd cell_6t
Xbit_r175_c40 bl[40] br[40] wl[175] vdd gnd cell_6t
Xbit_r176_c40 bl[40] br[40] wl[176] vdd gnd cell_6t
Xbit_r177_c40 bl[40] br[40] wl[177] vdd gnd cell_6t
Xbit_r178_c40 bl[40] br[40] wl[178] vdd gnd cell_6t
Xbit_r179_c40 bl[40] br[40] wl[179] vdd gnd cell_6t
Xbit_r180_c40 bl[40] br[40] wl[180] vdd gnd cell_6t
Xbit_r181_c40 bl[40] br[40] wl[181] vdd gnd cell_6t
Xbit_r182_c40 bl[40] br[40] wl[182] vdd gnd cell_6t
Xbit_r183_c40 bl[40] br[40] wl[183] vdd gnd cell_6t
Xbit_r184_c40 bl[40] br[40] wl[184] vdd gnd cell_6t
Xbit_r185_c40 bl[40] br[40] wl[185] vdd gnd cell_6t
Xbit_r186_c40 bl[40] br[40] wl[186] vdd gnd cell_6t
Xbit_r187_c40 bl[40] br[40] wl[187] vdd gnd cell_6t
Xbit_r188_c40 bl[40] br[40] wl[188] vdd gnd cell_6t
Xbit_r189_c40 bl[40] br[40] wl[189] vdd gnd cell_6t
Xbit_r190_c40 bl[40] br[40] wl[190] vdd gnd cell_6t
Xbit_r191_c40 bl[40] br[40] wl[191] vdd gnd cell_6t
Xbit_r192_c40 bl[40] br[40] wl[192] vdd gnd cell_6t
Xbit_r193_c40 bl[40] br[40] wl[193] vdd gnd cell_6t
Xbit_r194_c40 bl[40] br[40] wl[194] vdd gnd cell_6t
Xbit_r195_c40 bl[40] br[40] wl[195] vdd gnd cell_6t
Xbit_r196_c40 bl[40] br[40] wl[196] vdd gnd cell_6t
Xbit_r197_c40 bl[40] br[40] wl[197] vdd gnd cell_6t
Xbit_r198_c40 bl[40] br[40] wl[198] vdd gnd cell_6t
Xbit_r199_c40 bl[40] br[40] wl[199] vdd gnd cell_6t
Xbit_r200_c40 bl[40] br[40] wl[200] vdd gnd cell_6t
Xbit_r201_c40 bl[40] br[40] wl[201] vdd gnd cell_6t
Xbit_r202_c40 bl[40] br[40] wl[202] vdd gnd cell_6t
Xbit_r203_c40 bl[40] br[40] wl[203] vdd gnd cell_6t
Xbit_r204_c40 bl[40] br[40] wl[204] vdd gnd cell_6t
Xbit_r205_c40 bl[40] br[40] wl[205] vdd gnd cell_6t
Xbit_r206_c40 bl[40] br[40] wl[206] vdd gnd cell_6t
Xbit_r207_c40 bl[40] br[40] wl[207] vdd gnd cell_6t
Xbit_r208_c40 bl[40] br[40] wl[208] vdd gnd cell_6t
Xbit_r209_c40 bl[40] br[40] wl[209] vdd gnd cell_6t
Xbit_r210_c40 bl[40] br[40] wl[210] vdd gnd cell_6t
Xbit_r211_c40 bl[40] br[40] wl[211] vdd gnd cell_6t
Xbit_r212_c40 bl[40] br[40] wl[212] vdd gnd cell_6t
Xbit_r213_c40 bl[40] br[40] wl[213] vdd gnd cell_6t
Xbit_r214_c40 bl[40] br[40] wl[214] vdd gnd cell_6t
Xbit_r215_c40 bl[40] br[40] wl[215] vdd gnd cell_6t
Xbit_r216_c40 bl[40] br[40] wl[216] vdd gnd cell_6t
Xbit_r217_c40 bl[40] br[40] wl[217] vdd gnd cell_6t
Xbit_r218_c40 bl[40] br[40] wl[218] vdd gnd cell_6t
Xbit_r219_c40 bl[40] br[40] wl[219] vdd gnd cell_6t
Xbit_r220_c40 bl[40] br[40] wl[220] vdd gnd cell_6t
Xbit_r221_c40 bl[40] br[40] wl[221] vdd gnd cell_6t
Xbit_r222_c40 bl[40] br[40] wl[222] vdd gnd cell_6t
Xbit_r223_c40 bl[40] br[40] wl[223] vdd gnd cell_6t
Xbit_r224_c40 bl[40] br[40] wl[224] vdd gnd cell_6t
Xbit_r225_c40 bl[40] br[40] wl[225] vdd gnd cell_6t
Xbit_r226_c40 bl[40] br[40] wl[226] vdd gnd cell_6t
Xbit_r227_c40 bl[40] br[40] wl[227] vdd gnd cell_6t
Xbit_r228_c40 bl[40] br[40] wl[228] vdd gnd cell_6t
Xbit_r229_c40 bl[40] br[40] wl[229] vdd gnd cell_6t
Xbit_r230_c40 bl[40] br[40] wl[230] vdd gnd cell_6t
Xbit_r231_c40 bl[40] br[40] wl[231] vdd gnd cell_6t
Xbit_r232_c40 bl[40] br[40] wl[232] vdd gnd cell_6t
Xbit_r233_c40 bl[40] br[40] wl[233] vdd gnd cell_6t
Xbit_r234_c40 bl[40] br[40] wl[234] vdd gnd cell_6t
Xbit_r235_c40 bl[40] br[40] wl[235] vdd gnd cell_6t
Xbit_r236_c40 bl[40] br[40] wl[236] vdd gnd cell_6t
Xbit_r237_c40 bl[40] br[40] wl[237] vdd gnd cell_6t
Xbit_r238_c40 bl[40] br[40] wl[238] vdd gnd cell_6t
Xbit_r239_c40 bl[40] br[40] wl[239] vdd gnd cell_6t
Xbit_r240_c40 bl[40] br[40] wl[240] vdd gnd cell_6t
Xbit_r241_c40 bl[40] br[40] wl[241] vdd gnd cell_6t
Xbit_r242_c40 bl[40] br[40] wl[242] vdd gnd cell_6t
Xbit_r243_c40 bl[40] br[40] wl[243] vdd gnd cell_6t
Xbit_r244_c40 bl[40] br[40] wl[244] vdd gnd cell_6t
Xbit_r245_c40 bl[40] br[40] wl[245] vdd gnd cell_6t
Xbit_r246_c40 bl[40] br[40] wl[246] vdd gnd cell_6t
Xbit_r247_c40 bl[40] br[40] wl[247] vdd gnd cell_6t
Xbit_r248_c40 bl[40] br[40] wl[248] vdd gnd cell_6t
Xbit_r249_c40 bl[40] br[40] wl[249] vdd gnd cell_6t
Xbit_r250_c40 bl[40] br[40] wl[250] vdd gnd cell_6t
Xbit_r251_c40 bl[40] br[40] wl[251] vdd gnd cell_6t
Xbit_r252_c40 bl[40] br[40] wl[252] vdd gnd cell_6t
Xbit_r253_c40 bl[40] br[40] wl[253] vdd gnd cell_6t
Xbit_r254_c40 bl[40] br[40] wl[254] vdd gnd cell_6t
Xbit_r255_c40 bl[40] br[40] wl[255] vdd gnd cell_6t
Xbit_r0_c41 bl[41] br[41] wl[0] vdd gnd cell_6t
Xbit_r1_c41 bl[41] br[41] wl[1] vdd gnd cell_6t
Xbit_r2_c41 bl[41] br[41] wl[2] vdd gnd cell_6t
Xbit_r3_c41 bl[41] br[41] wl[3] vdd gnd cell_6t
Xbit_r4_c41 bl[41] br[41] wl[4] vdd gnd cell_6t
Xbit_r5_c41 bl[41] br[41] wl[5] vdd gnd cell_6t
Xbit_r6_c41 bl[41] br[41] wl[6] vdd gnd cell_6t
Xbit_r7_c41 bl[41] br[41] wl[7] vdd gnd cell_6t
Xbit_r8_c41 bl[41] br[41] wl[8] vdd gnd cell_6t
Xbit_r9_c41 bl[41] br[41] wl[9] vdd gnd cell_6t
Xbit_r10_c41 bl[41] br[41] wl[10] vdd gnd cell_6t
Xbit_r11_c41 bl[41] br[41] wl[11] vdd gnd cell_6t
Xbit_r12_c41 bl[41] br[41] wl[12] vdd gnd cell_6t
Xbit_r13_c41 bl[41] br[41] wl[13] vdd gnd cell_6t
Xbit_r14_c41 bl[41] br[41] wl[14] vdd gnd cell_6t
Xbit_r15_c41 bl[41] br[41] wl[15] vdd gnd cell_6t
Xbit_r16_c41 bl[41] br[41] wl[16] vdd gnd cell_6t
Xbit_r17_c41 bl[41] br[41] wl[17] vdd gnd cell_6t
Xbit_r18_c41 bl[41] br[41] wl[18] vdd gnd cell_6t
Xbit_r19_c41 bl[41] br[41] wl[19] vdd gnd cell_6t
Xbit_r20_c41 bl[41] br[41] wl[20] vdd gnd cell_6t
Xbit_r21_c41 bl[41] br[41] wl[21] vdd gnd cell_6t
Xbit_r22_c41 bl[41] br[41] wl[22] vdd gnd cell_6t
Xbit_r23_c41 bl[41] br[41] wl[23] vdd gnd cell_6t
Xbit_r24_c41 bl[41] br[41] wl[24] vdd gnd cell_6t
Xbit_r25_c41 bl[41] br[41] wl[25] vdd gnd cell_6t
Xbit_r26_c41 bl[41] br[41] wl[26] vdd gnd cell_6t
Xbit_r27_c41 bl[41] br[41] wl[27] vdd gnd cell_6t
Xbit_r28_c41 bl[41] br[41] wl[28] vdd gnd cell_6t
Xbit_r29_c41 bl[41] br[41] wl[29] vdd gnd cell_6t
Xbit_r30_c41 bl[41] br[41] wl[30] vdd gnd cell_6t
Xbit_r31_c41 bl[41] br[41] wl[31] vdd gnd cell_6t
Xbit_r32_c41 bl[41] br[41] wl[32] vdd gnd cell_6t
Xbit_r33_c41 bl[41] br[41] wl[33] vdd gnd cell_6t
Xbit_r34_c41 bl[41] br[41] wl[34] vdd gnd cell_6t
Xbit_r35_c41 bl[41] br[41] wl[35] vdd gnd cell_6t
Xbit_r36_c41 bl[41] br[41] wl[36] vdd gnd cell_6t
Xbit_r37_c41 bl[41] br[41] wl[37] vdd gnd cell_6t
Xbit_r38_c41 bl[41] br[41] wl[38] vdd gnd cell_6t
Xbit_r39_c41 bl[41] br[41] wl[39] vdd gnd cell_6t
Xbit_r40_c41 bl[41] br[41] wl[40] vdd gnd cell_6t
Xbit_r41_c41 bl[41] br[41] wl[41] vdd gnd cell_6t
Xbit_r42_c41 bl[41] br[41] wl[42] vdd gnd cell_6t
Xbit_r43_c41 bl[41] br[41] wl[43] vdd gnd cell_6t
Xbit_r44_c41 bl[41] br[41] wl[44] vdd gnd cell_6t
Xbit_r45_c41 bl[41] br[41] wl[45] vdd gnd cell_6t
Xbit_r46_c41 bl[41] br[41] wl[46] vdd gnd cell_6t
Xbit_r47_c41 bl[41] br[41] wl[47] vdd gnd cell_6t
Xbit_r48_c41 bl[41] br[41] wl[48] vdd gnd cell_6t
Xbit_r49_c41 bl[41] br[41] wl[49] vdd gnd cell_6t
Xbit_r50_c41 bl[41] br[41] wl[50] vdd gnd cell_6t
Xbit_r51_c41 bl[41] br[41] wl[51] vdd gnd cell_6t
Xbit_r52_c41 bl[41] br[41] wl[52] vdd gnd cell_6t
Xbit_r53_c41 bl[41] br[41] wl[53] vdd gnd cell_6t
Xbit_r54_c41 bl[41] br[41] wl[54] vdd gnd cell_6t
Xbit_r55_c41 bl[41] br[41] wl[55] vdd gnd cell_6t
Xbit_r56_c41 bl[41] br[41] wl[56] vdd gnd cell_6t
Xbit_r57_c41 bl[41] br[41] wl[57] vdd gnd cell_6t
Xbit_r58_c41 bl[41] br[41] wl[58] vdd gnd cell_6t
Xbit_r59_c41 bl[41] br[41] wl[59] vdd gnd cell_6t
Xbit_r60_c41 bl[41] br[41] wl[60] vdd gnd cell_6t
Xbit_r61_c41 bl[41] br[41] wl[61] vdd gnd cell_6t
Xbit_r62_c41 bl[41] br[41] wl[62] vdd gnd cell_6t
Xbit_r63_c41 bl[41] br[41] wl[63] vdd gnd cell_6t
Xbit_r64_c41 bl[41] br[41] wl[64] vdd gnd cell_6t
Xbit_r65_c41 bl[41] br[41] wl[65] vdd gnd cell_6t
Xbit_r66_c41 bl[41] br[41] wl[66] vdd gnd cell_6t
Xbit_r67_c41 bl[41] br[41] wl[67] vdd gnd cell_6t
Xbit_r68_c41 bl[41] br[41] wl[68] vdd gnd cell_6t
Xbit_r69_c41 bl[41] br[41] wl[69] vdd gnd cell_6t
Xbit_r70_c41 bl[41] br[41] wl[70] vdd gnd cell_6t
Xbit_r71_c41 bl[41] br[41] wl[71] vdd gnd cell_6t
Xbit_r72_c41 bl[41] br[41] wl[72] vdd gnd cell_6t
Xbit_r73_c41 bl[41] br[41] wl[73] vdd gnd cell_6t
Xbit_r74_c41 bl[41] br[41] wl[74] vdd gnd cell_6t
Xbit_r75_c41 bl[41] br[41] wl[75] vdd gnd cell_6t
Xbit_r76_c41 bl[41] br[41] wl[76] vdd gnd cell_6t
Xbit_r77_c41 bl[41] br[41] wl[77] vdd gnd cell_6t
Xbit_r78_c41 bl[41] br[41] wl[78] vdd gnd cell_6t
Xbit_r79_c41 bl[41] br[41] wl[79] vdd gnd cell_6t
Xbit_r80_c41 bl[41] br[41] wl[80] vdd gnd cell_6t
Xbit_r81_c41 bl[41] br[41] wl[81] vdd gnd cell_6t
Xbit_r82_c41 bl[41] br[41] wl[82] vdd gnd cell_6t
Xbit_r83_c41 bl[41] br[41] wl[83] vdd gnd cell_6t
Xbit_r84_c41 bl[41] br[41] wl[84] vdd gnd cell_6t
Xbit_r85_c41 bl[41] br[41] wl[85] vdd gnd cell_6t
Xbit_r86_c41 bl[41] br[41] wl[86] vdd gnd cell_6t
Xbit_r87_c41 bl[41] br[41] wl[87] vdd gnd cell_6t
Xbit_r88_c41 bl[41] br[41] wl[88] vdd gnd cell_6t
Xbit_r89_c41 bl[41] br[41] wl[89] vdd gnd cell_6t
Xbit_r90_c41 bl[41] br[41] wl[90] vdd gnd cell_6t
Xbit_r91_c41 bl[41] br[41] wl[91] vdd gnd cell_6t
Xbit_r92_c41 bl[41] br[41] wl[92] vdd gnd cell_6t
Xbit_r93_c41 bl[41] br[41] wl[93] vdd gnd cell_6t
Xbit_r94_c41 bl[41] br[41] wl[94] vdd gnd cell_6t
Xbit_r95_c41 bl[41] br[41] wl[95] vdd gnd cell_6t
Xbit_r96_c41 bl[41] br[41] wl[96] vdd gnd cell_6t
Xbit_r97_c41 bl[41] br[41] wl[97] vdd gnd cell_6t
Xbit_r98_c41 bl[41] br[41] wl[98] vdd gnd cell_6t
Xbit_r99_c41 bl[41] br[41] wl[99] vdd gnd cell_6t
Xbit_r100_c41 bl[41] br[41] wl[100] vdd gnd cell_6t
Xbit_r101_c41 bl[41] br[41] wl[101] vdd gnd cell_6t
Xbit_r102_c41 bl[41] br[41] wl[102] vdd gnd cell_6t
Xbit_r103_c41 bl[41] br[41] wl[103] vdd gnd cell_6t
Xbit_r104_c41 bl[41] br[41] wl[104] vdd gnd cell_6t
Xbit_r105_c41 bl[41] br[41] wl[105] vdd gnd cell_6t
Xbit_r106_c41 bl[41] br[41] wl[106] vdd gnd cell_6t
Xbit_r107_c41 bl[41] br[41] wl[107] vdd gnd cell_6t
Xbit_r108_c41 bl[41] br[41] wl[108] vdd gnd cell_6t
Xbit_r109_c41 bl[41] br[41] wl[109] vdd gnd cell_6t
Xbit_r110_c41 bl[41] br[41] wl[110] vdd gnd cell_6t
Xbit_r111_c41 bl[41] br[41] wl[111] vdd gnd cell_6t
Xbit_r112_c41 bl[41] br[41] wl[112] vdd gnd cell_6t
Xbit_r113_c41 bl[41] br[41] wl[113] vdd gnd cell_6t
Xbit_r114_c41 bl[41] br[41] wl[114] vdd gnd cell_6t
Xbit_r115_c41 bl[41] br[41] wl[115] vdd gnd cell_6t
Xbit_r116_c41 bl[41] br[41] wl[116] vdd gnd cell_6t
Xbit_r117_c41 bl[41] br[41] wl[117] vdd gnd cell_6t
Xbit_r118_c41 bl[41] br[41] wl[118] vdd gnd cell_6t
Xbit_r119_c41 bl[41] br[41] wl[119] vdd gnd cell_6t
Xbit_r120_c41 bl[41] br[41] wl[120] vdd gnd cell_6t
Xbit_r121_c41 bl[41] br[41] wl[121] vdd gnd cell_6t
Xbit_r122_c41 bl[41] br[41] wl[122] vdd gnd cell_6t
Xbit_r123_c41 bl[41] br[41] wl[123] vdd gnd cell_6t
Xbit_r124_c41 bl[41] br[41] wl[124] vdd gnd cell_6t
Xbit_r125_c41 bl[41] br[41] wl[125] vdd gnd cell_6t
Xbit_r126_c41 bl[41] br[41] wl[126] vdd gnd cell_6t
Xbit_r127_c41 bl[41] br[41] wl[127] vdd gnd cell_6t
Xbit_r128_c41 bl[41] br[41] wl[128] vdd gnd cell_6t
Xbit_r129_c41 bl[41] br[41] wl[129] vdd gnd cell_6t
Xbit_r130_c41 bl[41] br[41] wl[130] vdd gnd cell_6t
Xbit_r131_c41 bl[41] br[41] wl[131] vdd gnd cell_6t
Xbit_r132_c41 bl[41] br[41] wl[132] vdd gnd cell_6t
Xbit_r133_c41 bl[41] br[41] wl[133] vdd gnd cell_6t
Xbit_r134_c41 bl[41] br[41] wl[134] vdd gnd cell_6t
Xbit_r135_c41 bl[41] br[41] wl[135] vdd gnd cell_6t
Xbit_r136_c41 bl[41] br[41] wl[136] vdd gnd cell_6t
Xbit_r137_c41 bl[41] br[41] wl[137] vdd gnd cell_6t
Xbit_r138_c41 bl[41] br[41] wl[138] vdd gnd cell_6t
Xbit_r139_c41 bl[41] br[41] wl[139] vdd gnd cell_6t
Xbit_r140_c41 bl[41] br[41] wl[140] vdd gnd cell_6t
Xbit_r141_c41 bl[41] br[41] wl[141] vdd gnd cell_6t
Xbit_r142_c41 bl[41] br[41] wl[142] vdd gnd cell_6t
Xbit_r143_c41 bl[41] br[41] wl[143] vdd gnd cell_6t
Xbit_r144_c41 bl[41] br[41] wl[144] vdd gnd cell_6t
Xbit_r145_c41 bl[41] br[41] wl[145] vdd gnd cell_6t
Xbit_r146_c41 bl[41] br[41] wl[146] vdd gnd cell_6t
Xbit_r147_c41 bl[41] br[41] wl[147] vdd gnd cell_6t
Xbit_r148_c41 bl[41] br[41] wl[148] vdd gnd cell_6t
Xbit_r149_c41 bl[41] br[41] wl[149] vdd gnd cell_6t
Xbit_r150_c41 bl[41] br[41] wl[150] vdd gnd cell_6t
Xbit_r151_c41 bl[41] br[41] wl[151] vdd gnd cell_6t
Xbit_r152_c41 bl[41] br[41] wl[152] vdd gnd cell_6t
Xbit_r153_c41 bl[41] br[41] wl[153] vdd gnd cell_6t
Xbit_r154_c41 bl[41] br[41] wl[154] vdd gnd cell_6t
Xbit_r155_c41 bl[41] br[41] wl[155] vdd gnd cell_6t
Xbit_r156_c41 bl[41] br[41] wl[156] vdd gnd cell_6t
Xbit_r157_c41 bl[41] br[41] wl[157] vdd gnd cell_6t
Xbit_r158_c41 bl[41] br[41] wl[158] vdd gnd cell_6t
Xbit_r159_c41 bl[41] br[41] wl[159] vdd gnd cell_6t
Xbit_r160_c41 bl[41] br[41] wl[160] vdd gnd cell_6t
Xbit_r161_c41 bl[41] br[41] wl[161] vdd gnd cell_6t
Xbit_r162_c41 bl[41] br[41] wl[162] vdd gnd cell_6t
Xbit_r163_c41 bl[41] br[41] wl[163] vdd gnd cell_6t
Xbit_r164_c41 bl[41] br[41] wl[164] vdd gnd cell_6t
Xbit_r165_c41 bl[41] br[41] wl[165] vdd gnd cell_6t
Xbit_r166_c41 bl[41] br[41] wl[166] vdd gnd cell_6t
Xbit_r167_c41 bl[41] br[41] wl[167] vdd gnd cell_6t
Xbit_r168_c41 bl[41] br[41] wl[168] vdd gnd cell_6t
Xbit_r169_c41 bl[41] br[41] wl[169] vdd gnd cell_6t
Xbit_r170_c41 bl[41] br[41] wl[170] vdd gnd cell_6t
Xbit_r171_c41 bl[41] br[41] wl[171] vdd gnd cell_6t
Xbit_r172_c41 bl[41] br[41] wl[172] vdd gnd cell_6t
Xbit_r173_c41 bl[41] br[41] wl[173] vdd gnd cell_6t
Xbit_r174_c41 bl[41] br[41] wl[174] vdd gnd cell_6t
Xbit_r175_c41 bl[41] br[41] wl[175] vdd gnd cell_6t
Xbit_r176_c41 bl[41] br[41] wl[176] vdd gnd cell_6t
Xbit_r177_c41 bl[41] br[41] wl[177] vdd gnd cell_6t
Xbit_r178_c41 bl[41] br[41] wl[178] vdd gnd cell_6t
Xbit_r179_c41 bl[41] br[41] wl[179] vdd gnd cell_6t
Xbit_r180_c41 bl[41] br[41] wl[180] vdd gnd cell_6t
Xbit_r181_c41 bl[41] br[41] wl[181] vdd gnd cell_6t
Xbit_r182_c41 bl[41] br[41] wl[182] vdd gnd cell_6t
Xbit_r183_c41 bl[41] br[41] wl[183] vdd gnd cell_6t
Xbit_r184_c41 bl[41] br[41] wl[184] vdd gnd cell_6t
Xbit_r185_c41 bl[41] br[41] wl[185] vdd gnd cell_6t
Xbit_r186_c41 bl[41] br[41] wl[186] vdd gnd cell_6t
Xbit_r187_c41 bl[41] br[41] wl[187] vdd gnd cell_6t
Xbit_r188_c41 bl[41] br[41] wl[188] vdd gnd cell_6t
Xbit_r189_c41 bl[41] br[41] wl[189] vdd gnd cell_6t
Xbit_r190_c41 bl[41] br[41] wl[190] vdd gnd cell_6t
Xbit_r191_c41 bl[41] br[41] wl[191] vdd gnd cell_6t
Xbit_r192_c41 bl[41] br[41] wl[192] vdd gnd cell_6t
Xbit_r193_c41 bl[41] br[41] wl[193] vdd gnd cell_6t
Xbit_r194_c41 bl[41] br[41] wl[194] vdd gnd cell_6t
Xbit_r195_c41 bl[41] br[41] wl[195] vdd gnd cell_6t
Xbit_r196_c41 bl[41] br[41] wl[196] vdd gnd cell_6t
Xbit_r197_c41 bl[41] br[41] wl[197] vdd gnd cell_6t
Xbit_r198_c41 bl[41] br[41] wl[198] vdd gnd cell_6t
Xbit_r199_c41 bl[41] br[41] wl[199] vdd gnd cell_6t
Xbit_r200_c41 bl[41] br[41] wl[200] vdd gnd cell_6t
Xbit_r201_c41 bl[41] br[41] wl[201] vdd gnd cell_6t
Xbit_r202_c41 bl[41] br[41] wl[202] vdd gnd cell_6t
Xbit_r203_c41 bl[41] br[41] wl[203] vdd gnd cell_6t
Xbit_r204_c41 bl[41] br[41] wl[204] vdd gnd cell_6t
Xbit_r205_c41 bl[41] br[41] wl[205] vdd gnd cell_6t
Xbit_r206_c41 bl[41] br[41] wl[206] vdd gnd cell_6t
Xbit_r207_c41 bl[41] br[41] wl[207] vdd gnd cell_6t
Xbit_r208_c41 bl[41] br[41] wl[208] vdd gnd cell_6t
Xbit_r209_c41 bl[41] br[41] wl[209] vdd gnd cell_6t
Xbit_r210_c41 bl[41] br[41] wl[210] vdd gnd cell_6t
Xbit_r211_c41 bl[41] br[41] wl[211] vdd gnd cell_6t
Xbit_r212_c41 bl[41] br[41] wl[212] vdd gnd cell_6t
Xbit_r213_c41 bl[41] br[41] wl[213] vdd gnd cell_6t
Xbit_r214_c41 bl[41] br[41] wl[214] vdd gnd cell_6t
Xbit_r215_c41 bl[41] br[41] wl[215] vdd gnd cell_6t
Xbit_r216_c41 bl[41] br[41] wl[216] vdd gnd cell_6t
Xbit_r217_c41 bl[41] br[41] wl[217] vdd gnd cell_6t
Xbit_r218_c41 bl[41] br[41] wl[218] vdd gnd cell_6t
Xbit_r219_c41 bl[41] br[41] wl[219] vdd gnd cell_6t
Xbit_r220_c41 bl[41] br[41] wl[220] vdd gnd cell_6t
Xbit_r221_c41 bl[41] br[41] wl[221] vdd gnd cell_6t
Xbit_r222_c41 bl[41] br[41] wl[222] vdd gnd cell_6t
Xbit_r223_c41 bl[41] br[41] wl[223] vdd gnd cell_6t
Xbit_r224_c41 bl[41] br[41] wl[224] vdd gnd cell_6t
Xbit_r225_c41 bl[41] br[41] wl[225] vdd gnd cell_6t
Xbit_r226_c41 bl[41] br[41] wl[226] vdd gnd cell_6t
Xbit_r227_c41 bl[41] br[41] wl[227] vdd gnd cell_6t
Xbit_r228_c41 bl[41] br[41] wl[228] vdd gnd cell_6t
Xbit_r229_c41 bl[41] br[41] wl[229] vdd gnd cell_6t
Xbit_r230_c41 bl[41] br[41] wl[230] vdd gnd cell_6t
Xbit_r231_c41 bl[41] br[41] wl[231] vdd gnd cell_6t
Xbit_r232_c41 bl[41] br[41] wl[232] vdd gnd cell_6t
Xbit_r233_c41 bl[41] br[41] wl[233] vdd gnd cell_6t
Xbit_r234_c41 bl[41] br[41] wl[234] vdd gnd cell_6t
Xbit_r235_c41 bl[41] br[41] wl[235] vdd gnd cell_6t
Xbit_r236_c41 bl[41] br[41] wl[236] vdd gnd cell_6t
Xbit_r237_c41 bl[41] br[41] wl[237] vdd gnd cell_6t
Xbit_r238_c41 bl[41] br[41] wl[238] vdd gnd cell_6t
Xbit_r239_c41 bl[41] br[41] wl[239] vdd gnd cell_6t
Xbit_r240_c41 bl[41] br[41] wl[240] vdd gnd cell_6t
Xbit_r241_c41 bl[41] br[41] wl[241] vdd gnd cell_6t
Xbit_r242_c41 bl[41] br[41] wl[242] vdd gnd cell_6t
Xbit_r243_c41 bl[41] br[41] wl[243] vdd gnd cell_6t
Xbit_r244_c41 bl[41] br[41] wl[244] vdd gnd cell_6t
Xbit_r245_c41 bl[41] br[41] wl[245] vdd gnd cell_6t
Xbit_r246_c41 bl[41] br[41] wl[246] vdd gnd cell_6t
Xbit_r247_c41 bl[41] br[41] wl[247] vdd gnd cell_6t
Xbit_r248_c41 bl[41] br[41] wl[248] vdd gnd cell_6t
Xbit_r249_c41 bl[41] br[41] wl[249] vdd gnd cell_6t
Xbit_r250_c41 bl[41] br[41] wl[250] vdd gnd cell_6t
Xbit_r251_c41 bl[41] br[41] wl[251] vdd gnd cell_6t
Xbit_r252_c41 bl[41] br[41] wl[252] vdd gnd cell_6t
Xbit_r253_c41 bl[41] br[41] wl[253] vdd gnd cell_6t
Xbit_r254_c41 bl[41] br[41] wl[254] vdd gnd cell_6t
Xbit_r255_c41 bl[41] br[41] wl[255] vdd gnd cell_6t
Xbit_r0_c42 bl[42] br[42] wl[0] vdd gnd cell_6t
Xbit_r1_c42 bl[42] br[42] wl[1] vdd gnd cell_6t
Xbit_r2_c42 bl[42] br[42] wl[2] vdd gnd cell_6t
Xbit_r3_c42 bl[42] br[42] wl[3] vdd gnd cell_6t
Xbit_r4_c42 bl[42] br[42] wl[4] vdd gnd cell_6t
Xbit_r5_c42 bl[42] br[42] wl[5] vdd gnd cell_6t
Xbit_r6_c42 bl[42] br[42] wl[6] vdd gnd cell_6t
Xbit_r7_c42 bl[42] br[42] wl[7] vdd gnd cell_6t
Xbit_r8_c42 bl[42] br[42] wl[8] vdd gnd cell_6t
Xbit_r9_c42 bl[42] br[42] wl[9] vdd gnd cell_6t
Xbit_r10_c42 bl[42] br[42] wl[10] vdd gnd cell_6t
Xbit_r11_c42 bl[42] br[42] wl[11] vdd gnd cell_6t
Xbit_r12_c42 bl[42] br[42] wl[12] vdd gnd cell_6t
Xbit_r13_c42 bl[42] br[42] wl[13] vdd gnd cell_6t
Xbit_r14_c42 bl[42] br[42] wl[14] vdd gnd cell_6t
Xbit_r15_c42 bl[42] br[42] wl[15] vdd gnd cell_6t
Xbit_r16_c42 bl[42] br[42] wl[16] vdd gnd cell_6t
Xbit_r17_c42 bl[42] br[42] wl[17] vdd gnd cell_6t
Xbit_r18_c42 bl[42] br[42] wl[18] vdd gnd cell_6t
Xbit_r19_c42 bl[42] br[42] wl[19] vdd gnd cell_6t
Xbit_r20_c42 bl[42] br[42] wl[20] vdd gnd cell_6t
Xbit_r21_c42 bl[42] br[42] wl[21] vdd gnd cell_6t
Xbit_r22_c42 bl[42] br[42] wl[22] vdd gnd cell_6t
Xbit_r23_c42 bl[42] br[42] wl[23] vdd gnd cell_6t
Xbit_r24_c42 bl[42] br[42] wl[24] vdd gnd cell_6t
Xbit_r25_c42 bl[42] br[42] wl[25] vdd gnd cell_6t
Xbit_r26_c42 bl[42] br[42] wl[26] vdd gnd cell_6t
Xbit_r27_c42 bl[42] br[42] wl[27] vdd gnd cell_6t
Xbit_r28_c42 bl[42] br[42] wl[28] vdd gnd cell_6t
Xbit_r29_c42 bl[42] br[42] wl[29] vdd gnd cell_6t
Xbit_r30_c42 bl[42] br[42] wl[30] vdd gnd cell_6t
Xbit_r31_c42 bl[42] br[42] wl[31] vdd gnd cell_6t
Xbit_r32_c42 bl[42] br[42] wl[32] vdd gnd cell_6t
Xbit_r33_c42 bl[42] br[42] wl[33] vdd gnd cell_6t
Xbit_r34_c42 bl[42] br[42] wl[34] vdd gnd cell_6t
Xbit_r35_c42 bl[42] br[42] wl[35] vdd gnd cell_6t
Xbit_r36_c42 bl[42] br[42] wl[36] vdd gnd cell_6t
Xbit_r37_c42 bl[42] br[42] wl[37] vdd gnd cell_6t
Xbit_r38_c42 bl[42] br[42] wl[38] vdd gnd cell_6t
Xbit_r39_c42 bl[42] br[42] wl[39] vdd gnd cell_6t
Xbit_r40_c42 bl[42] br[42] wl[40] vdd gnd cell_6t
Xbit_r41_c42 bl[42] br[42] wl[41] vdd gnd cell_6t
Xbit_r42_c42 bl[42] br[42] wl[42] vdd gnd cell_6t
Xbit_r43_c42 bl[42] br[42] wl[43] vdd gnd cell_6t
Xbit_r44_c42 bl[42] br[42] wl[44] vdd gnd cell_6t
Xbit_r45_c42 bl[42] br[42] wl[45] vdd gnd cell_6t
Xbit_r46_c42 bl[42] br[42] wl[46] vdd gnd cell_6t
Xbit_r47_c42 bl[42] br[42] wl[47] vdd gnd cell_6t
Xbit_r48_c42 bl[42] br[42] wl[48] vdd gnd cell_6t
Xbit_r49_c42 bl[42] br[42] wl[49] vdd gnd cell_6t
Xbit_r50_c42 bl[42] br[42] wl[50] vdd gnd cell_6t
Xbit_r51_c42 bl[42] br[42] wl[51] vdd gnd cell_6t
Xbit_r52_c42 bl[42] br[42] wl[52] vdd gnd cell_6t
Xbit_r53_c42 bl[42] br[42] wl[53] vdd gnd cell_6t
Xbit_r54_c42 bl[42] br[42] wl[54] vdd gnd cell_6t
Xbit_r55_c42 bl[42] br[42] wl[55] vdd gnd cell_6t
Xbit_r56_c42 bl[42] br[42] wl[56] vdd gnd cell_6t
Xbit_r57_c42 bl[42] br[42] wl[57] vdd gnd cell_6t
Xbit_r58_c42 bl[42] br[42] wl[58] vdd gnd cell_6t
Xbit_r59_c42 bl[42] br[42] wl[59] vdd gnd cell_6t
Xbit_r60_c42 bl[42] br[42] wl[60] vdd gnd cell_6t
Xbit_r61_c42 bl[42] br[42] wl[61] vdd gnd cell_6t
Xbit_r62_c42 bl[42] br[42] wl[62] vdd gnd cell_6t
Xbit_r63_c42 bl[42] br[42] wl[63] vdd gnd cell_6t
Xbit_r64_c42 bl[42] br[42] wl[64] vdd gnd cell_6t
Xbit_r65_c42 bl[42] br[42] wl[65] vdd gnd cell_6t
Xbit_r66_c42 bl[42] br[42] wl[66] vdd gnd cell_6t
Xbit_r67_c42 bl[42] br[42] wl[67] vdd gnd cell_6t
Xbit_r68_c42 bl[42] br[42] wl[68] vdd gnd cell_6t
Xbit_r69_c42 bl[42] br[42] wl[69] vdd gnd cell_6t
Xbit_r70_c42 bl[42] br[42] wl[70] vdd gnd cell_6t
Xbit_r71_c42 bl[42] br[42] wl[71] vdd gnd cell_6t
Xbit_r72_c42 bl[42] br[42] wl[72] vdd gnd cell_6t
Xbit_r73_c42 bl[42] br[42] wl[73] vdd gnd cell_6t
Xbit_r74_c42 bl[42] br[42] wl[74] vdd gnd cell_6t
Xbit_r75_c42 bl[42] br[42] wl[75] vdd gnd cell_6t
Xbit_r76_c42 bl[42] br[42] wl[76] vdd gnd cell_6t
Xbit_r77_c42 bl[42] br[42] wl[77] vdd gnd cell_6t
Xbit_r78_c42 bl[42] br[42] wl[78] vdd gnd cell_6t
Xbit_r79_c42 bl[42] br[42] wl[79] vdd gnd cell_6t
Xbit_r80_c42 bl[42] br[42] wl[80] vdd gnd cell_6t
Xbit_r81_c42 bl[42] br[42] wl[81] vdd gnd cell_6t
Xbit_r82_c42 bl[42] br[42] wl[82] vdd gnd cell_6t
Xbit_r83_c42 bl[42] br[42] wl[83] vdd gnd cell_6t
Xbit_r84_c42 bl[42] br[42] wl[84] vdd gnd cell_6t
Xbit_r85_c42 bl[42] br[42] wl[85] vdd gnd cell_6t
Xbit_r86_c42 bl[42] br[42] wl[86] vdd gnd cell_6t
Xbit_r87_c42 bl[42] br[42] wl[87] vdd gnd cell_6t
Xbit_r88_c42 bl[42] br[42] wl[88] vdd gnd cell_6t
Xbit_r89_c42 bl[42] br[42] wl[89] vdd gnd cell_6t
Xbit_r90_c42 bl[42] br[42] wl[90] vdd gnd cell_6t
Xbit_r91_c42 bl[42] br[42] wl[91] vdd gnd cell_6t
Xbit_r92_c42 bl[42] br[42] wl[92] vdd gnd cell_6t
Xbit_r93_c42 bl[42] br[42] wl[93] vdd gnd cell_6t
Xbit_r94_c42 bl[42] br[42] wl[94] vdd gnd cell_6t
Xbit_r95_c42 bl[42] br[42] wl[95] vdd gnd cell_6t
Xbit_r96_c42 bl[42] br[42] wl[96] vdd gnd cell_6t
Xbit_r97_c42 bl[42] br[42] wl[97] vdd gnd cell_6t
Xbit_r98_c42 bl[42] br[42] wl[98] vdd gnd cell_6t
Xbit_r99_c42 bl[42] br[42] wl[99] vdd gnd cell_6t
Xbit_r100_c42 bl[42] br[42] wl[100] vdd gnd cell_6t
Xbit_r101_c42 bl[42] br[42] wl[101] vdd gnd cell_6t
Xbit_r102_c42 bl[42] br[42] wl[102] vdd gnd cell_6t
Xbit_r103_c42 bl[42] br[42] wl[103] vdd gnd cell_6t
Xbit_r104_c42 bl[42] br[42] wl[104] vdd gnd cell_6t
Xbit_r105_c42 bl[42] br[42] wl[105] vdd gnd cell_6t
Xbit_r106_c42 bl[42] br[42] wl[106] vdd gnd cell_6t
Xbit_r107_c42 bl[42] br[42] wl[107] vdd gnd cell_6t
Xbit_r108_c42 bl[42] br[42] wl[108] vdd gnd cell_6t
Xbit_r109_c42 bl[42] br[42] wl[109] vdd gnd cell_6t
Xbit_r110_c42 bl[42] br[42] wl[110] vdd gnd cell_6t
Xbit_r111_c42 bl[42] br[42] wl[111] vdd gnd cell_6t
Xbit_r112_c42 bl[42] br[42] wl[112] vdd gnd cell_6t
Xbit_r113_c42 bl[42] br[42] wl[113] vdd gnd cell_6t
Xbit_r114_c42 bl[42] br[42] wl[114] vdd gnd cell_6t
Xbit_r115_c42 bl[42] br[42] wl[115] vdd gnd cell_6t
Xbit_r116_c42 bl[42] br[42] wl[116] vdd gnd cell_6t
Xbit_r117_c42 bl[42] br[42] wl[117] vdd gnd cell_6t
Xbit_r118_c42 bl[42] br[42] wl[118] vdd gnd cell_6t
Xbit_r119_c42 bl[42] br[42] wl[119] vdd gnd cell_6t
Xbit_r120_c42 bl[42] br[42] wl[120] vdd gnd cell_6t
Xbit_r121_c42 bl[42] br[42] wl[121] vdd gnd cell_6t
Xbit_r122_c42 bl[42] br[42] wl[122] vdd gnd cell_6t
Xbit_r123_c42 bl[42] br[42] wl[123] vdd gnd cell_6t
Xbit_r124_c42 bl[42] br[42] wl[124] vdd gnd cell_6t
Xbit_r125_c42 bl[42] br[42] wl[125] vdd gnd cell_6t
Xbit_r126_c42 bl[42] br[42] wl[126] vdd gnd cell_6t
Xbit_r127_c42 bl[42] br[42] wl[127] vdd gnd cell_6t
Xbit_r128_c42 bl[42] br[42] wl[128] vdd gnd cell_6t
Xbit_r129_c42 bl[42] br[42] wl[129] vdd gnd cell_6t
Xbit_r130_c42 bl[42] br[42] wl[130] vdd gnd cell_6t
Xbit_r131_c42 bl[42] br[42] wl[131] vdd gnd cell_6t
Xbit_r132_c42 bl[42] br[42] wl[132] vdd gnd cell_6t
Xbit_r133_c42 bl[42] br[42] wl[133] vdd gnd cell_6t
Xbit_r134_c42 bl[42] br[42] wl[134] vdd gnd cell_6t
Xbit_r135_c42 bl[42] br[42] wl[135] vdd gnd cell_6t
Xbit_r136_c42 bl[42] br[42] wl[136] vdd gnd cell_6t
Xbit_r137_c42 bl[42] br[42] wl[137] vdd gnd cell_6t
Xbit_r138_c42 bl[42] br[42] wl[138] vdd gnd cell_6t
Xbit_r139_c42 bl[42] br[42] wl[139] vdd gnd cell_6t
Xbit_r140_c42 bl[42] br[42] wl[140] vdd gnd cell_6t
Xbit_r141_c42 bl[42] br[42] wl[141] vdd gnd cell_6t
Xbit_r142_c42 bl[42] br[42] wl[142] vdd gnd cell_6t
Xbit_r143_c42 bl[42] br[42] wl[143] vdd gnd cell_6t
Xbit_r144_c42 bl[42] br[42] wl[144] vdd gnd cell_6t
Xbit_r145_c42 bl[42] br[42] wl[145] vdd gnd cell_6t
Xbit_r146_c42 bl[42] br[42] wl[146] vdd gnd cell_6t
Xbit_r147_c42 bl[42] br[42] wl[147] vdd gnd cell_6t
Xbit_r148_c42 bl[42] br[42] wl[148] vdd gnd cell_6t
Xbit_r149_c42 bl[42] br[42] wl[149] vdd gnd cell_6t
Xbit_r150_c42 bl[42] br[42] wl[150] vdd gnd cell_6t
Xbit_r151_c42 bl[42] br[42] wl[151] vdd gnd cell_6t
Xbit_r152_c42 bl[42] br[42] wl[152] vdd gnd cell_6t
Xbit_r153_c42 bl[42] br[42] wl[153] vdd gnd cell_6t
Xbit_r154_c42 bl[42] br[42] wl[154] vdd gnd cell_6t
Xbit_r155_c42 bl[42] br[42] wl[155] vdd gnd cell_6t
Xbit_r156_c42 bl[42] br[42] wl[156] vdd gnd cell_6t
Xbit_r157_c42 bl[42] br[42] wl[157] vdd gnd cell_6t
Xbit_r158_c42 bl[42] br[42] wl[158] vdd gnd cell_6t
Xbit_r159_c42 bl[42] br[42] wl[159] vdd gnd cell_6t
Xbit_r160_c42 bl[42] br[42] wl[160] vdd gnd cell_6t
Xbit_r161_c42 bl[42] br[42] wl[161] vdd gnd cell_6t
Xbit_r162_c42 bl[42] br[42] wl[162] vdd gnd cell_6t
Xbit_r163_c42 bl[42] br[42] wl[163] vdd gnd cell_6t
Xbit_r164_c42 bl[42] br[42] wl[164] vdd gnd cell_6t
Xbit_r165_c42 bl[42] br[42] wl[165] vdd gnd cell_6t
Xbit_r166_c42 bl[42] br[42] wl[166] vdd gnd cell_6t
Xbit_r167_c42 bl[42] br[42] wl[167] vdd gnd cell_6t
Xbit_r168_c42 bl[42] br[42] wl[168] vdd gnd cell_6t
Xbit_r169_c42 bl[42] br[42] wl[169] vdd gnd cell_6t
Xbit_r170_c42 bl[42] br[42] wl[170] vdd gnd cell_6t
Xbit_r171_c42 bl[42] br[42] wl[171] vdd gnd cell_6t
Xbit_r172_c42 bl[42] br[42] wl[172] vdd gnd cell_6t
Xbit_r173_c42 bl[42] br[42] wl[173] vdd gnd cell_6t
Xbit_r174_c42 bl[42] br[42] wl[174] vdd gnd cell_6t
Xbit_r175_c42 bl[42] br[42] wl[175] vdd gnd cell_6t
Xbit_r176_c42 bl[42] br[42] wl[176] vdd gnd cell_6t
Xbit_r177_c42 bl[42] br[42] wl[177] vdd gnd cell_6t
Xbit_r178_c42 bl[42] br[42] wl[178] vdd gnd cell_6t
Xbit_r179_c42 bl[42] br[42] wl[179] vdd gnd cell_6t
Xbit_r180_c42 bl[42] br[42] wl[180] vdd gnd cell_6t
Xbit_r181_c42 bl[42] br[42] wl[181] vdd gnd cell_6t
Xbit_r182_c42 bl[42] br[42] wl[182] vdd gnd cell_6t
Xbit_r183_c42 bl[42] br[42] wl[183] vdd gnd cell_6t
Xbit_r184_c42 bl[42] br[42] wl[184] vdd gnd cell_6t
Xbit_r185_c42 bl[42] br[42] wl[185] vdd gnd cell_6t
Xbit_r186_c42 bl[42] br[42] wl[186] vdd gnd cell_6t
Xbit_r187_c42 bl[42] br[42] wl[187] vdd gnd cell_6t
Xbit_r188_c42 bl[42] br[42] wl[188] vdd gnd cell_6t
Xbit_r189_c42 bl[42] br[42] wl[189] vdd gnd cell_6t
Xbit_r190_c42 bl[42] br[42] wl[190] vdd gnd cell_6t
Xbit_r191_c42 bl[42] br[42] wl[191] vdd gnd cell_6t
Xbit_r192_c42 bl[42] br[42] wl[192] vdd gnd cell_6t
Xbit_r193_c42 bl[42] br[42] wl[193] vdd gnd cell_6t
Xbit_r194_c42 bl[42] br[42] wl[194] vdd gnd cell_6t
Xbit_r195_c42 bl[42] br[42] wl[195] vdd gnd cell_6t
Xbit_r196_c42 bl[42] br[42] wl[196] vdd gnd cell_6t
Xbit_r197_c42 bl[42] br[42] wl[197] vdd gnd cell_6t
Xbit_r198_c42 bl[42] br[42] wl[198] vdd gnd cell_6t
Xbit_r199_c42 bl[42] br[42] wl[199] vdd gnd cell_6t
Xbit_r200_c42 bl[42] br[42] wl[200] vdd gnd cell_6t
Xbit_r201_c42 bl[42] br[42] wl[201] vdd gnd cell_6t
Xbit_r202_c42 bl[42] br[42] wl[202] vdd gnd cell_6t
Xbit_r203_c42 bl[42] br[42] wl[203] vdd gnd cell_6t
Xbit_r204_c42 bl[42] br[42] wl[204] vdd gnd cell_6t
Xbit_r205_c42 bl[42] br[42] wl[205] vdd gnd cell_6t
Xbit_r206_c42 bl[42] br[42] wl[206] vdd gnd cell_6t
Xbit_r207_c42 bl[42] br[42] wl[207] vdd gnd cell_6t
Xbit_r208_c42 bl[42] br[42] wl[208] vdd gnd cell_6t
Xbit_r209_c42 bl[42] br[42] wl[209] vdd gnd cell_6t
Xbit_r210_c42 bl[42] br[42] wl[210] vdd gnd cell_6t
Xbit_r211_c42 bl[42] br[42] wl[211] vdd gnd cell_6t
Xbit_r212_c42 bl[42] br[42] wl[212] vdd gnd cell_6t
Xbit_r213_c42 bl[42] br[42] wl[213] vdd gnd cell_6t
Xbit_r214_c42 bl[42] br[42] wl[214] vdd gnd cell_6t
Xbit_r215_c42 bl[42] br[42] wl[215] vdd gnd cell_6t
Xbit_r216_c42 bl[42] br[42] wl[216] vdd gnd cell_6t
Xbit_r217_c42 bl[42] br[42] wl[217] vdd gnd cell_6t
Xbit_r218_c42 bl[42] br[42] wl[218] vdd gnd cell_6t
Xbit_r219_c42 bl[42] br[42] wl[219] vdd gnd cell_6t
Xbit_r220_c42 bl[42] br[42] wl[220] vdd gnd cell_6t
Xbit_r221_c42 bl[42] br[42] wl[221] vdd gnd cell_6t
Xbit_r222_c42 bl[42] br[42] wl[222] vdd gnd cell_6t
Xbit_r223_c42 bl[42] br[42] wl[223] vdd gnd cell_6t
Xbit_r224_c42 bl[42] br[42] wl[224] vdd gnd cell_6t
Xbit_r225_c42 bl[42] br[42] wl[225] vdd gnd cell_6t
Xbit_r226_c42 bl[42] br[42] wl[226] vdd gnd cell_6t
Xbit_r227_c42 bl[42] br[42] wl[227] vdd gnd cell_6t
Xbit_r228_c42 bl[42] br[42] wl[228] vdd gnd cell_6t
Xbit_r229_c42 bl[42] br[42] wl[229] vdd gnd cell_6t
Xbit_r230_c42 bl[42] br[42] wl[230] vdd gnd cell_6t
Xbit_r231_c42 bl[42] br[42] wl[231] vdd gnd cell_6t
Xbit_r232_c42 bl[42] br[42] wl[232] vdd gnd cell_6t
Xbit_r233_c42 bl[42] br[42] wl[233] vdd gnd cell_6t
Xbit_r234_c42 bl[42] br[42] wl[234] vdd gnd cell_6t
Xbit_r235_c42 bl[42] br[42] wl[235] vdd gnd cell_6t
Xbit_r236_c42 bl[42] br[42] wl[236] vdd gnd cell_6t
Xbit_r237_c42 bl[42] br[42] wl[237] vdd gnd cell_6t
Xbit_r238_c42 bl[42] br[42] wl[238] vdd gnd cell_6t
Xbit_r239_c42 bl[42] br[42] wl[239] vdd gnd cell_6t
Xbit_r240_c42 bl[42] br[42] wl[240] vdd gnd cell_6t
Xbit_r241_c42 bl[42] br[42] wl[241] vdd gnd cell_6t
Xbit_r242_c42 bl[42] br[42] wl[242] vdd gnd cell_6t
Xbit_r243_c42 bl[42] br[42] wl[243] vdd gnd cell_6t
Xbit_r244_c42 bl[42] br[42] wl[244] vdd gnd cell_6t
Xbit_r245_c42 bl[42] br[42] wl[245] vdd gnd cell_6t
Xbit_r246_c42 bl[42] br[42] wl[246] vdd gnd cell_6t
Xbit_r247_c42 bl[42] br[42] wl[247] vdd gnd cell_6t
Xbit_r248_c42 bl[42] br[42] wl[248] vdd gnd cell_6t
Xbit_r249_c42 bl[42] br[42] wl[249] vdd gnd cell_6t
Xbit_r250_c42 bl[42] br[42] wl[250] vdd gnd cell_6t
Xbit_r251_c42 bl[42] br[42] wl[251] vdd gnd cell_6t
Xbit_r252_c42 bl[42] br[42] wl[252] vdd gnd cell_6t
Xbit_r253_c42 bl[42] br[42] wl[253] vdd gnd cell_6t
Xbit_r254_c42 bl[42] br[42] wl[254] vdd gnd cell_6t
Xbit_r255_c42 bl[42] br[42] wl[255] vdd gnd cell_6t
Xbit_r0_c43 bl[43] br[43] wl[0] vdd gnd cell_6t
Xbit_r1_c43 bl[43] br[43] wl[1] vdd gnd cell_6t
Xbit_r2_c43 bl[43] br[43] wl[2] vdd gnd cell_6t
Xbit_r3_c43 bl[43] br[43] wl[3] vdd gnd cell_6t
Xbit_r4_c43 bl[43] br[43] wl[4] vdd gnd cell_6t
Xbit_r5_c43 bl[43] br[43] wl[5] vdd gnd cell_6t
Xbit_r6_c43 bl[43] br[43] wl[6] vdd gnd cell_6t
Xbit_r7_c43 bl[43] br[43] wl[7] vdd gnd cell_6t
Xbit_r8_c43 bl[43] br[43] wl[8] vdd gnd cell_6t
Xbit_r9_c43 bl[43] br[43] wl[9] vdd gnd cell_6t
Xbit_r10_c43 bl[43] br[43] wl[10] vdd gnd cell_6t
Xbit_r11_c43 bl[43] br[43] wl[11] vdd gnd cell_6t
Xbit_r12_c43 bl[43] br[43] wl[12] vdd gnd cell_6t
Xbit_r13_c43 bl[43] br[43] wl[13] vdd gnd cell_6t
Xbit_r14_c43 bl[43] br[43] wl[14] vdd gnd cell_6t
Xbit_r15_c43 bl[43] br[43] wl[15] vdd gnd cell_6t
Xbit_r16_c43 bl[43] br[43] wl[16] vdd gnd cell_6t
Xbit_r17_c43 bl[43] br[43] wl[17] vdd gnd cell_6t
Xbit_r18_c43 bl[43] br[43] wl[18] vdd gnd cell_6t
Xbit_r19_c43 bl[43] br[43] wl[19] vdd gnd cell_6t
Xbit_r20_c43 bl[43] br[43] wl[20] vdd gnd cell_6t
Xbit_r21_c43 bl[43] br[43] wl[21] vdd gnd cell_6t
Xbit_r22_c43 bl[43] br[43] wl[22] vdd gnd cell_6t
Xbit_r23_c43 bl[43] br[43] wl[23] vdd gnd cell_6t
Xbit_r24_c43 bl[43] br[43] wl[24] vdd gnd cell_6t
Xbit_r25_c43 bl[43] br[43] wl[25] vdd gnd cell_6t
Xbit_r26_c43 bl[43] br[43] wl[26] vdd gnd cell_6t
Xbit_r27_c43 bl[43] br[43] wl[27] vdd gnd cell_6t
Xbit_r28_c43 bl[43] br[43] wl[28] vdd gnd cell_6t
Xbit_r29_c43 bl[43] br[43] wl[29] vdd gnd cell_6t
Xbit_r30_c43 bl[43] br[43] wl[30] vdd gnd cell_6t
Xbit_r31_c43 bl[43] br[43] wl[31] vdd gnd cell_6t
Xbit_r32_c43 bl[43] br[43] wl[32] vdd gnd cell_6t
Xbit_r33_c43 bl[43] br[43] wl[33] vdd gnd cell_6t
Xbit_r34_c43 bl[43] br[43] wl[34] vdd gnd cell_6t
Xbit_r35_c43 bl[43] br[43] wl[35] vdd gnd cell_6t
Xbit_r36_c43 bl[43] br[43] wl[36] vdd gnd cell_6t
Xbit_r37_c43 bl[43] br[43] wl[37] vdd gnd cell_6t
Xbit_r38_c43 bl[43] br[43] wl[38] vdd gnd cell_6t
Xbit_r39_c43 bl[43] br[43] wl[39] vdd gnd cell_6t
Xbit_r40_c43 bl[43] br[43] wl[40] vdd gnd cell_6t
Xbit_r41_c43 bl[43] br[43] wl[41] vdd gnd cell_6t
Xbit_r42_c43 bl[43] br[43] wl[42] vdd gnd cell_6t
Xbit_r43_c43 bl[43] br[43] wl[43] vdd gnd cell_6t
Xbit_r44_c43 bl[43] br[43] wl[44] vdd gnd cell_6t
Xbit_r45_c43 bl[43] br[43] wl[45] vdd gnd cell_6t
Xbit_r46_c43 bl[43] br[43] wl[46] vdd gnd cell_6t
Xbit_r47_c43 bl[43] br[43] wl[47] vdd gnd cell_6t
Xbit_r48_c43 bl[43] br[43] wl[48] vdd gnd cell_6t
Xbit_r49_c43 bl[43] br[43] wl[49] vdd gnd cell_6t
Xbit_r50_c43 bl[43] br[43] wl[50] vdd gnd cell_6t
Xbit_r51_c43 bl[43] br[43] wl[51] vdd gnd cell_6t
Xbit_r52_c43 bl[43] br[43] wl[52] vdd gnd cell_6t
Xbit_r53_c43 bl[43] br[43] wl[53] vdd gnd cell_6t
Xbit_r54_c43 bl[43] br[43] wl[54] vdd gnd cell_6t
Xbit_r55_c43 bl[43] br[43] wl[55] vdd gnd cell_6t
Xbit_r56_c43 bl[43] br[43] wl[56] vdd gnd cell_6t
Xbit_r57_c43 bl[43] br[43] wl[57] vdd gnd cell_6t
Xbit_r58_c43 bl[43] br[43] wl[58] vdd gnd cell_6t
Xbit_r59_c43 bl[43] br[43] wl[59] vdd gnd cell_6t
Xbit_r60_c43 bl[43] br[43] wl[60] vdd gnd cell_6t
Xbit_r61_c43 bl[43] br[43] wl[61] vdd gnd cell_6t
Xbit_r62_c43 bl[43] br[43] wl[62] vdd gnd cell_6t
Xbit_r63_c43 bl[43] br[43] wl[63] vdd gnd cell_6t
Xbit_r64_c43 bl[43] br[43] wl[64] vdd gnd cell_6t
Xbit_r65_c43 bl[43] br[43] wl[65] vdd gnd cell_6t
Xbit_r66_c43 bl[43] br[43] wl[66] vdd gnd cell_6t
Xbit_r67_c43 bl[43] br[43] wl[67] vdd gnd cell_6t
Xbit_r68_c43 bl[43] br[43] wl[68] vdd gnd cell_6t
Xbit_r69_c43 bl[43] br[43] wl[69] vdd gnd cell_6t
Xbit_r70_c43 bl[43] br[43] wl[70] vdd gnd cell_6t
Xbit_r71_c43 bl[43] br[43] wl[71] vdd gnd cell_6t
Xbit_r72_c43 bl[43] br[43] wl[72] vdd gnd cell_6t
Xbit_r73_c43 bl[43] br[43] wl[73] vdd gnd cell_6t
Xbit_r74_c43 bl[43] br[43] wl[74] vdd gnd cell_6t
Xbit_r75_c43 bl[43] br[43] wl[75] vdd gnd cell_6t
Xbit_r76_c43 bl[43] br[43] wl[76] vdd gnd cell_6t
Xbit_r77_c43 bl[43] br[43] wl[77] vdd gnd cell_6t
Xbit_r78_c43 bl[43] br[43] wl[78] vdd gnd cell_6t
Xbit_r79_c43 bl[43] br[43] wl[79] vdd gnd cell_6t
Xbit_r80_c43 bl[43] br[43] wl[80] vdd gnd cell_6t
Xbit_r81_c43 bl[43] br[43] wl[81] vdd gnd cell_6t
Xbit_r82_c43 bl[43] br[43] wl[82] vdd gnd cell_6t
Xbit_r83_c43 bl[43] br[43] wl[83] vdd gnd cell_6t
Xbit_r84_c43 bl[43] br[43] wl[84] vdd gnd cell_6t
Xbit_r85_c43 bl[43] br[43] wl[85] vdd gnd cell_6t
Xbit_r86_c43 bl[43] br[43] wl[86] vdd gnd cell_6t
Xbit_r87_c43 bl[43] br[43] wl[87] vdd gnd cell_6t
Xbit_r88_c43 bl[43] br[43] wl[88] vdd gnd cell_6t
Xbit_r89_c43 bl[43] br[43] wl[89] vdd gnd cell_6t
Xbit_r90_c43 bl[43] br[43] wl[90] vdd gnd cell_6t
Xbit_r91_c43 bl[43] br[43] wl[91] vdd gnd cell_6t
Xbit_r92_c43 bl[43] br[43] wl[92] vdd gnd cell_6t
Xbit_r93_c43 bl[43] br[43] wl[93] vdd gnd cell_6t
Xbit_r94_c43 bl[43] br[43] wl[94] vdd gnd cell_6t
Xbit_r95_c43 bl[43] br[43] wl[95] vdd gnd cell_6t
Xbit_r96_c43 bl[43] br[43] wl[96] vdd gnd cell_6t
Xbit_r97_c43 bl[43] br[43] wl[97] vdd gnd cell_6t
Xbit_r98_c43 bl[43] br[43] wl[98] vdd gnd cell_6t
Xbit_r99_c43 bl[43] br[43] wl[99] vdd gnd cell_6t
Xbit_r100_c43 bl[43] br[43] wl[100] vdd gnd cell_6t
Xbit_r101_c43 bl[43] br[43] wl[101] vdd gnd cell_6t
Xbit_r102_c43 bl[43] br[43] wl[102] vdd gnd cell_6t
Xbit_r103_c43 bl[43] br[43] wl[103] vdd gnd cell_6t
Xbit_r104_c43 bl[43] br[43] wl[104] vdd gnd cell_6t
Xbit_r105_c43 bl[43] br[43] wl[105] vdd gnd cell_6t
Xbit_r106_c43 bl[43] br[43] wl[106] vdd gnd cell_6t
Xbit_r107_c43 bl[43] br[43] wl[107] vdd gnd cell_6t
Xbit_r108_c43 bl[43] br[43] wl[108] vdd gnd cell_6t
Xbit_r109_c43 bl[43] br[43] wl[109] vdd gnd cell_6t
Xbit_r110_c43 bl[43] br[43] wl[110] vdd gnd cell_6t
Xbit_r111_c43 bl[43] br[43] wl[111] vdd gnd cell_6t
Xbit_r112_c43 bl[43] br[43] wl[112] vdd gnd cell_6t
Xbit_r113_c43 bl[43] br[43] wl[113] vdd gnd cell_6t
Xbit_r114_c43 bl[43] br[43] wl[114] vdd gnd cell_6t
Xbit_r115_c43 bl[43] br[43] wl[115] vdd gnd cell_6t
Xbit_r116_c43 bl[43] br[43] wl[116] vdd gnd cell_6t
Xbit_r117_c43 bl[43] br[43] wl[117] vdd gnd cell_6t
Xbit_r118_c43 bl[43] br[43] wl[118] vdd gnd cell_6t
Xbit_r119_c43 bl[43] br[43] wl[119] vdd gnd cell_6t
Xbit_r120_c43 bl[43] br[43] wl[120] vdd gnd cell_6t
Xbit_r121_c43 bl[43] br[43] wl[121] vdd gnd cell_6t
Xbit_r122_c43 bl[43] br[43] wl[122] vdd gnd cell_6t
Xbit_r123_c43 bl[43] br[43] wl[123] vdd gnd cell_6t
Xbit_r124_c43 bl[43] br[43] wl[124] vdd gnd cell_6t
Xbit_r125_c43 bl[43] br[43] wl[125] vdd gnd cell_6t
Xbit_r126_c43 bl[43] br[43] wl[126] vdd gnd cell_6t
Xbit_r127_c43 bl[43] br[43] wl[127] vdd gnd cell_6t
Xbit_r128_c43 bl[43] br[43] wl[128] vdd gnd cell_6t
Xbit_r129_c43 bl[43] br[43] wl[129] vdd gnd cell_6t
Xbit_r130_c43 bl[43] br[43] wl[130] vdd gnd cell_6t
Xbit_r131_c43 bl[43] br[43] wl[131] vdd gnd cell_6t
Xbit_r132_c43 bl[43] br[43] wl[132] vdd gnd cell_6t
Xbit_r133_c43 bl[43] br[43] wl[133] vdd gnd cell_6t
Xbit_r134_c43 bl[43] br[43] wl[134] vdd gnd cell_6t
Xbit_r135_c43 bl[43] br[43] wl[135] vdd gnd cell_6t
Xbit_r136_c43 bl[43] br[43] wl[136] vdd gnd cell_6t
Xbit_r137_c43 bl[43] br[43] wl[137] vdd gnd cell_6t
Xbit_r138_c43 bl[43] br[43] wl[138] vdd gnd cell_6t
Xbit_r139_c43 bl[43] br[43] wl[139] vdd gnd cell_6t
Xbit_r140_c43 bl[43] br[43] wl[140] vdd gnd cell_6t
Xbit_r141_c43 bl[43] br[43] wl[141] vdd gnd cell_6t
Xbit_r142_c43 bl[43] br[43] wl[142] vdd gnd cell_6t
Xbit_r143_c43 bl[43] br[43] wl[143] vdd gnd cell_6t
Xbit_r144_c43 bl[43] br[43] wl[144] vdd gnd cell_6t
Xbit_r145_c43 bl[43] br[43] wl[145] vdd gnd cell_6t
Xbit_r146_c43 bl[43] br[43] wl[146] vdd gnd cell_6t
Xbit_r147_c43 bl[43] br[43] wl[147] vdd gnd cell_6t
Xbit_r148_c43 bl[43] br[43] wl[148] vdd gnd cell_6t
Xbit_r149_c43 bl[43] br[43] wl[149] vdd gnd cell_6t
Xbit_r150_c43 bl[43] br[43] wl[150] vdd gnd cell_6t
Xbit_r151_c43 bl[43] br[43] wl[151] vdd gnd cell_6t
Xbit_r152_c43 bl[43] br[43] wl[152] vdd gnd cell_6t
Xbit_r153_c43 bl[43] br[43] wl[153] vdd gnd cell_6t
Xbit_r154_c43 bl[43] br[43] wl[154] vdd gnd cell_6t
Xbit_r155_c43 bl[43] br[43] wl[155] vdd gnd cell_6t
Xbit_r156_c43 bl[43] br[43] wl[156] vdd gnd cell_6t
Xbit_r157_c43 bl[43] br[43] wl[157] vdd gnd cell_6t
Xbit_r158_c43 bl[43] br[43] wl[158] vdd gnd cell_6t
Xbit_r159_c43 bl[43] br[43] wl[159] vdd gnd cell_6t
Xbit_r160_c43 bl[43] br[43] wl[160] vdd gnd cell_6t
Xbit_r161_c43 bl[43] br[43] wl[161] vdd gnd cell_6t
Xbit_r162_c43 bl[43] br[43] wl[162] vdd gnd cell_6t
Xbit_r163_c43 bl[43] br[43] wl[163] vdd gnd cell_6t
Xbit_r164_c43 bl[43] br[43] wl[164] vdd gnd cell_6t
Xbit_r165_c43 bl[43] br[43] wl[165] vdd gnd cell_6t
Xbit_r166_c43 bl[43] br[43] wl[166] vdd gnd cell_6t
Xbit_r167_c43 bl[43] br[43] wl[167] vdd gnd cell_6t
Xbit_r168_c43 bl[43] br[43] wl[168] vdd gnd cell_6t
Xbit_r169_c43 bl[43] br[43] wl[169] vdd gnd cell_6t
Xbit_r170_c43 bl[43] br[43] wl[170] vdd gnd cell_6t
Xbit_r171_c43 bl[43] br[43] wl[171] vdd gnd cell_6t
Xbit_r172_c43 bl[43] br[43] wl[172] vdd gnd cell_6t
Xbit_r173_c43 bl[43] br[43] wl[173] vdd gnd cell_6t
Xbit_r174_c43 bl[43] br[43] wl[174] vdd gnd cell_6t
Xbit_r175_c43 bl[43] br[43] wl[175] vdd gnd cell_6t
Xbit_r176_c43 bl[43] br[43] wl[176] vdd gnd cell_6t
Xbit_r177_c43 bl[43] br[43] wl[177] vdd gnd cell_6t
Xbit_r178_c43 bl[43] br[43] wl[178] vdd gnd cell_6t
Xbit_r179_c43 bl[43] br[43] wl[179] vdd gnd cell_6t
Xbit_r180_c43 bl[43] br[43] wl[180] vdd gnd cell_6t
Xbit_r181_c43 bl[43] br[43] wl[181] vdd gnd cell_6t
Xbit_r182_c43 bl[43] br[43] wl[182] vdd gnd cell_6t
Xbit_r183_c43 bl[43] br[43] wl[183] vdd gnd cell_6t
Xbit_r184_c43 bl[43] br[43] wl[184] vdd gnd cell_6t
Xbit_r185_c43 bl[43] br[43] wl[185] vdd gnd cell_6t
Xbit_r186_c43 bl[43] br[43] wl[186] vdd gnd cell_6t
Xbit_r187_c43 bl[43] br[43] wl[187] vdd gnd cell_6t
Xbit_r188_c43 bl[43] br[43] wl[188] vdd gnd cell_6t
Xbit_r189_c43 bl[43] br[43] wl[189] vdd gnd cell_6t
Xbit_r190_c43 bl[43] br[43] wl[190] vdd gnd cell_6t
Xbit_r191_c43 bl[43] br[43] wl[191] vdd gnd cell_6t
Xbit_r192_c43 bl[43] br[43] wl[192] vdd gnd cell_6t
Xbit_r193_c43 bl[43] br[43] wl[193] vdd gnd cell_6t
Xbit_r194_c43 bl[43] br[43] wl[194] vdd gnd cell_6t
Xbit_r195_c43 bl[43] br[43] wl[195] vdd gnd cell_6t
Xbit_r196_c43 bl[43] br[43] wl[196] vdd gnd cell_6t
Xbit_r197_c43 bl[43] br[43] wl[197] vdd gnd cell_6t
Xbit_r198_c43 bl[43] br[43] wl[198] vdd gnd cell_6t
Xbit_r199_c43 bl[43] br[43] wl[199] vdd gnd cell_6t
Xbit_r200_c43 bl[43] br[43] wl[200] vdd gnd cell_6t
Xbit_r201_c43 bl[43] br[43] wl[201] vdd gnd cell_6t
Xbit_r202_c43 bl[43] br[43] wl[202] vdd gnd cell_6t
Xbit_r203_c43 bl[43] br[43] wl[203] vdd gnd cell_6t
Xbit_r204_c43 bl[43] br[43] wl[204] vdd gnd cell_6t
Xbit_r205_c43 bl[43] br[43] wl[205] vdd gnd cell_6t
Xbit_r206_c43 bl[43] br[43] wl[206] vdd gnd cell_6t
Xbit_r207_c43 bl[43] br[43] wl[207] vdd gnd cell_6t
Xbit_r208_c43 bl[43] br[43] wl[208] vdd gnd cell_6t
Xbit_r209_c43 bl[43] br[43] wl[209] vdd gnd cell_6t
Xbit_r210_c43 bl[43] br[43] wl[210] vdd gnd cell_6t
Xbit_r211_c43 bl[43] br[43] wl[211] vdd gnd cell_6t
Xbit_r212_c43 bl[43] br[43] wl[212] vdd gnd cell_6t
Xbit_r213_c43 bl[43] br[43] wl[213] vdd gnd cell_6t
Xbit_r214_c43 bl[43] br[43] wl[214] vdd gnd cell_6t
Xbit_r215_c43 bl[43] br[43] wl[215] vdd gnd cell_6t
Xbit_r216_c43 bl[43] br[43] wl[216] vdd gnd cell_6t
Xbit_r217_c43 bl[43] br[43] wl[217] vdd gnd cell_6t
Xbit_r218_c43 bl[43] br[43] wl[218] vdd gnd cell_6t
Xbit_r219_c43 bl[43] br[43] wl[219] vdd gnd cell_6t
Xbit_r220_c43 bl[43] br[43] wl[220] vdd gnd cell_6t
Xbit_r221_c43 bl[43] br[43] wl[221] vdd gnd cell_6t
Xbit_r222_c43 bl[43] br[43] wl[222] vdd gnd cell_6t
Xbit_r223_c43 bl[43] br[43] wl[223] vdd gnd cell_6t
Xbit_r224_c43 bl[43] br[43] wl[224] vdd gnd cell_6t
Xbit_r225_c43 bl[43] br[43] wl[225] vdd gnd cell_6t
Xbit_r226_c43 bl[43] br[43] wl[226] vdd gnd cell_6t
Xbit_r227_c43 bl[43] br[43] wl[227] vdd gnd cell_6t
Xbit_r228_c43 bl[43] br[43] wl[228] vdd gnd cell_6t
Xbit_r229_c43 bl[43] br[43] wl[229] vdd gnd cell_6t
Xbit_r230_c43 bl[43] br[43] wl[230] vdd gnd cell_6t
Xbit_r231_c43 bl[43] br[43] wl[231] vdd gnd cell_6t
Xbit_r232_c43 bl[43] br[43] wl[232] vdd gnd cell_6t
Xbit_r233_c43 bl[43] br[43] wl[233] vdd gnd cell_6t
Xbit_r234_c43 bl[43] br[43] wl[234] vdd gnd cell_6t
Xbit_r235_c43 bl[43] br[43] wl[235] vdd gnd cell_6t
Xbit_r236_c43 bl[43] br[43] wl[236] vdd gnd cell_6t
Xbit_r237_c43 bl[43] br[43] wl[237] vdd gnd cell_6t
Xbit_r238_c43 bl[43] br[43] wl[238] vdd gnd cell_6t
Xbit_r239_c43 bl[43] br[43] wl[239] vdd gnd cell_6t
Xbit_r240_c43 bl[43] br[43] wl[240] vdd gnd cell_6t
Xbit_r241_c43 bl[43] br[43] wl[241] vdd gnd cell_6t
Xbit_r242_c43 bl[43] br[43] wl[242] vdd gnd cell_6t
Xbit_r243_c43 bl[43] br[43] wl[243] vdd gnd cell_6t
Xbit_r244_c43 bl[43] br[43] wl[244] vdd gnd cell_6t
Xbit_r245_c43 bl[43] br[43] wl[245] vdd gnd cell_6t
Xbit_r246_c43 bl[43] br[43] wl[246] vdd gnd cell_6t
Xbit_r247_c43 bl[43] br[43] wl[247] vdd gnd cell_6t
Xbit_r248_c43 bl[43] br[43] wl[248] vdd gnd cell_6t
Xbit_r249_c43 bl[43] br[43] wl[249] vdd gnd cell_6t
Xbit_r250_c43 bl[43] br[43] wl[250] vdd gnd cell_6t
Xbit_r251_c43 bl[43] br[43] wl[251] vdd gnd cell_6t
Xbit_r252_c43 bl[43] br[43] wl[252] vdd gnd cell_6t
Xbit_r253_c43 bl[43] br[43] wl[253] vdd gnd cell_6t
Xbit_r254_c43 bl[43] br[43] wl[254] vdd gnd cell_6t
Xbit_r255_c43 bl[43] br[43] wl[255] vdd gnd cell_6t
Xbit_r0_c44 bl[44] br[44] wl[0] vdd gnd cell_6t
Xbit_r1_c44 bl[44] br[44] wl[1] vdd gnd cell_6t
Xbit_r2_c44 bl[44] br[44] wl[2] vdd gnd cell_6t
Xbit_r3_c44 bl[44] br[44] wl[3] vdd gnd cell_6t
Xbit_r4_c44 bl[44] br[44] wl[4] vdd gnd cell_6t
Xbit_r5_c44 bl[44] br[44] wl[5] vdd gnd cell_6t
Xbit_r6_c44 bl[44] br[44] wl[6] vdd gnd cell_6t
Xbit_r7_c44 bl[44] br[44] wl[7] vdd gnd cell_6t
Xbit_r8_c44 bl[44] br[44] wl[8] vdd gnd cell_6t
Xbit_r9_c44 bl[44] br[44] wl[9] vdd gnd cell_6t
Xbit_r10_c44 bl[44] br[44] wl[10] vdd gnd cell_6t
Xbit_r11_c44 bl[44] br[44] wl[11] vdd gnd cell_6t
Xbit_r12_c44 bl[44] br[44] wl[12] vdd gnd cell_6t
Xbit_r13_c44 bl[44] br[44] wl[13] vdd gnd cell_6t
Xbit_r14_c44 bl[44] br[44] wl[14] vdd gnd cell_6t
Xbit_r15_c44 bl[44] br[44] wl[15] vdd gnd cell_6t
Xbit_r16_c44 bl[44] br[44] wl[16] vdd gnd cell_6t
Xbit_r17_c44 bl[44] br[44] wl[17] vdd gnd cell_6t
Xbit_r18_c44 bl[44] br[44] wl[18] vdd gnd cell_6t
Xbit_r19_c44 bl[44] br[44] wl[19] vdd gnd cell_6t
Xbit_r20_c44 bl[44] br[44] wl[20] vdd gnd cell_6t
Xbit_r21_c44 bl[44] br[44] wl[21] vdd gnd cell_6t
Xbit_r22_c44 bl[44] br[44] wl[22] vdd gnd cell_6t
Xbit_r23_c44 bl[44] br[44] wl[23] vdd gnd cell_6t
Xbit_r24_c44 bl[44] br[44] wl[24] vdd gnd cell_6t
Xbit_r25_c44 bl[44] br[44] wl[25] vdd gnd cell_6t
Xbit_r26_c44 bl[44] br[44] wl[26] vdd gnd cell_6t
Xbit_r27_c44 bl[44] br[44] wl[27] vdd gnd cell_6t
Xbit_r28_c44 bl[44] br[44] wl[28] vdd gnd cell_6t
Xbit_r29_c44 bl[44] br[44] wl[29] vdd gnd cell_6t
Xbit_r30_c44 bl[44] br[44] wl[30] vdd gnd cell_6t
Xbit_r31_c44 bl[44] br[44] wl[31] vdd gnd cell_6t
Xbit_r32_c44 bl[44] br[44] wl[32] vdd gnd cell_6t
Xbit_r33_c44 bl[44] br[44] wl[33] vdd gnd cell_6t
Xbit_r34_c44 bl[44] br[44] wl[34] vdd gnd cell_6t
Xbit_r35_c44 bl[44] br[44] wl[35] vdd gnd cell_6t
Xbit_r36_c44 bl[44] br[44] wl[36] vdd gnd cell_6t
Xbit_r37_c44 bl[44] br[44] wl[37] vdd gnd cell_6t
Xbit_r38_c44 bl[44] br[44] wl[38] vdd gnd cell_6t
Xbit_r39_c44 bl[44] br[44] wl[39] vdd gnd cell_6t
Xbit_r40_c44 bl[44] br[44] wl[40] vdd gnd cell_6t
Xbit_r41_c44 bl[44] br[44] wl[41] vdd gnd cell_6t
Xbit_r42_c44 bl[44] br[44] wl[42] vdd gnd cell_6t
Xbit_r43_c44 bl[44] br[44] wl[43] vdd gnd cell_6t
Xbit_r44_c44 bl[44] br[44] wl[44] vdd gnd cell_6t
Xbit_r45_c44 bl[44] br[44] wl[45] vdd gnd cell_6t
Xbit_r46_c44 bl[44] br[44] wl[46] vdd gnd cell_6t
Xbit_r47_c44 bl[44] br[44] wl[47] vdd gnd cell_6t
Xbit_r48_c44 bl[44] br[44] wl[48] vdd gnd cell_6t
Xbit_r49_c44 bl[44] br[44] wl[49] vdd gnd cell_6t
Xbit_r50_c44 bl[44] br[44] wl[50] vdd gnd cell_6t
Xbit_r51_c44 bl[44] br[44] wl[51] vdd gnd cell_6t
Xbit_r52_c44 bl[44] br[44] wl[52] vdd gnd cell_6t
Xbit_r53_c44 bl[44] br[44] wl[53] vdd gnd cell_6t
Xbit_r54_c44 bl[44] br[44] wl[54] vdd gnd cell_6t
Xbit_r55_c44 bl[44] br[44] wl[55] vdd gnd cell_6t
Xbit_r56_c44 bl[44] br[44] wl[56] vdd gnd cell_6t
Xbit_r57_c44 bl[44] br[44] wl[57] vdd gnd cell_6t
Xbit_r58_c44 bl[44] br[44] wl[58] vdd gnd cell_6t
Xbit_r59_c44 bl[44] br[44] wl[59] vdd gnd cell_6t
Xbit_r60_c44 bl[44] br[44] wl[60] vdd gnd cell_6t
Xbit_r61_c44 bl[44] br[44] wl[61] vdd gnd cell_6t
Xbit_r62_c44 bl[44] br[44] wl[62] vdd gnd cell_6t
Xbit_r63_c44 bl[44] br[44] wl[63] vdd gnd cell_6t
Xbit_r64_c44 bl[44] br[44] wl[64] vdd gnd cell_6t
Xbit_r65_c44 bl[44] br[44] wl[65] vdd gnd cell_6t
Xbit_r66_c44 bl[44] br[44] wl[66] vdd gnd cell_6t
Xbit_r67_c44 bl[44] br[44] wl[67] vdd gnd cell_6t
Xbit_r68_c44 bl[44] br[44] wl[68] vdd gnd cell_6t
Xbit_r69_c44 bl[44] br[44] wl[69] vdd gnd cell_6t
Xbit_r70_c44 bl[44] br[44] wl[70] vdd gnd cell_6t
Xbit_r71_c44 bl[44] br[44] wl[71] vdd gnd cell_6t
Xbit_r72_c44 bl[44] br[44] wl[72] vdd gnd cell_6t
Xbit_r73_c44 bl[44] br[44] wl[73] vdd gnd cell_6t
Xbit_r74_c44 bl[44] br[44] wl[74] vdd gnd cell_6t
Xbit_r75_c44 bl[44] br[44] wl[75] vdd gnd cell_6t
Xbit_r76_c44 bl[44] br[44] wl[76] vdd gnd cell_6t
Xbit_r77_c44 bl[44] br[44] wl[77] vdd gnd cell_6t
Xbit_r78_c44 bl[44] br[44] wl[78] vdd gnd cell_6t
Xbit_r79_c44 bl[44] br[44] wl[79] vdd gnd cell_6t
Xbit_r80_c44 bl[44] br[44] wl[80] vdd gnd cell_6t
Xbit_r81_c44 bl[44] br[44] wl[81] vdd gnd cell_6t
Xbit_r82_c44 bl[44] br[44] wl[82] vdd gnd cell_6t
Xbit_r83_c44 bl[44] br[44] wl[83] vdd gnd cell_6t
Xbit_r84_c44 bl[44] br[44] wl[84] vdd gnd cell_6t
Xbit_r85_c44 bl[44] br[44] wl[85] vdd gnd cell_6t
Xbit_r86_c44 bl[44] br[44] wl[86] vdd gnd cell_6t
Xbit_r87_c44 bl[44] br[44] wl[87] vdd gnd cell_6t
Xbit_r88_c44 bl[44] br[44] wl[88] vdd gnd cell_6t
Xbit_r89_c44 bl[44] br[44] wl[89] vdd gnd cell_6t
Xbit_r90_c44 bl[44] br[44] wl[90] vdd gnd cell_6t
Xbit_r91_c44 bl[44] br[44] wl[91] vdd gnd cell_6t
Xbit_r92_c44 bl[44] br[44] wl[92] vdd gnd cell_6t
Xbit_r93_c44 bl[44] br[44] wl[93] vdd gnd cell_6t
Xbit_r94_c44 bl[44] br[44] wl[94] vdd gnd cell_6t
Xbit_r95_c44 bl[44] br[44] wl[95] vdd gnd cell_6t
Xbit_r96_c44 bl[44] br[44] wl[96] vdd gnd cell_6t
Xbit_r97_c44 bl[44] br[44] wl[97] vdd gnd cell_6t
Xbit_r98_c44 bl[44] br[44] wl[98] vdd gnd cell_6t
Xbit_r99_c44 bl[44] br[44] wl[99] vdd gnd cell_6t
Xbit_r100_c44 bl[44] br[44] wl[100] vdd gnd cell_6t
Xbit_r101_c44 bl[44] br[44] wl[101] vdd gnd cell_6t
Xbit_r102_c44 bl[44] br[44] wl[102] vdd gnd cell_6t
Xbit_r103_c44 bl[44] br[44] wl[103] vdd gnd cell_6t
Xbit_r104_c44 bl[44] br[44] wl[104] vdd gnd cell_6t
Xbit_r105_c44 bl[44] br[44] wl[105] vdd gnd cell_6t
Xbit_r106_c44 bl[44] br[44] wl[106] vdd gnd cell_6t
Xbit_r107_c44 bl[44] br[44] wl[107] vdd gnd cell_6t
Xbit_r108_c44 bl[44] br[44] wl[108] vdd gnd cell_6t
Xbit_r109_c44 bl[44] br[44] wl[109] vdd gnd cell_6t
Xbit_r110_c44 bl[44] br[44] wl[110] vdd gnd cell_6t
Xbit_r111_c44 bl[44] br[44] wl[111] vdd gnd cell_6t
Xbit_r112_c44 bl[44] br[44] wl[112] vdd gnd cell_6t
Xbit_r113_c44 bl[44] br[44] wl[113] vdd gnd cell_6t
Xbit_r114_c44 bl[44] br[44] wl[114] vdd gnd cell_6t
Xbit_r115_c44 bl[44] br[44] wl[115] vdd gnd cell_6t
Xbit_r116_c44 bl[44] br[44] wl[116] vdd gnd cell_6t
Xbit_r117_c44 bl[44] br[44] wl[117] vdd gnd cell_6t
Xbit_r118_c44 bl[44] br[44] wl[118] vdd gnd cell_6t
Xbit_r119_c44 bl[44] br[44] wl[119] vdd gnd cell_6t
Xbit_r120_c44 bl[44] br[44] wl[120] vdd gnd cell_6t
Xbit_r121_c44 bl[44] br[44] wl[121] vdd gnd cell_6t
Xbit_r122_c44 bl[44] br[44] wl[122] vdd gnd cell_6t
Xbit_r123_c44 bl[44] br[44] wl[123] vdd gnd cell_6t
Xbit_r124_c44 bl[44] br[44] wl[124] vdd gnd cell_6t
Xbit_r125_c44 bl[44] br[44] wl[125] vdd gnd cell_6t
Xbit_r126_c44 bl[44] br[44] wl[126] vdd gnd cell_6t
Xbit_r127_c44 bl[44] br[44] wl[127] vdd gnd cell_6t
Xbit_r128_c44 bl[44] br[44] wl[128] vdd gnd cell_6t
Xbit_r129_c44 bl[44] br[44] wl[129] vdd gnd cell_6t
Xbit_r130_c44 bl[44] br[44] wl[130] vdd gnd cell_6t
Xbit_r131_c44 bl[44] br[44] wl[131] vdd gnd cell_6t
Xbit_r132_c44 bl[44] br[44] wl[132] vdd gnd cell_6t
Xbit_r133_c44 bl[44] br[44] wl[133] vdd gnd cell_6t
Xbit_r134_c44 bl[44] br[44] wl[134] vdd gnd cell_6t
Xbit_r135_c44 bl[44] br[44] wl[135] vdd gnd cell_6t
Xbit_r136_c44 bl[44] br[44] wl[136] vdd gnd cell_6t
Xbit_r137_c44 bl[44] br[44] wl[137] vdd gnd cell_6t
Xbit_r138_c44 bl[44] br[44] wl[138] vdd gnd cell_6t
Xbit_r139_c44 bl[44] br[44] wl[139] vdd gnd cell_6t
Xbit_r140_c44 bl[44] br[44] wl[140] vdd gnd cell_6t
Xbit_r141_c44 bl[44] br[44] wl[141] vdd gnd cell_6t
Xbit_r142_c44 bl[44] br[44] wl[142] vdd gnd cell_6t
Xbit_r143_c44 bl[44] br[44] wl[143] vdd gnd cell_6t
Xbit_r144_c44 bl[44] br[44] wl[144] vdd gnd cell_6t
Xbit_r145_c44 bl[44] br[44] wl[145] vdd gnd cell_6t
Xbit_r146_c44 bl[44] br[44] wl[146] vdd gnd cell_6t
Xbit_r147_c44 bl[44] br[44] wl[147] vdd gnd cell_6t
Xbit_r148_c44 bl[44] br[44] wl[148] vdd gnd cell_6t
Xbit_r149_c44 bl[44] br[44] wl[149] vdd gnd cell_6t
Xbit_r150_c44 bl[44] br[44] wl[150] vdd gnd cell_6t
Xbit_r151_c44 bl[44] br[44] wl[151] vdd gnd cell_6t
Xbit_r152_c44 bl[44] br[44] wl[152] vdd gnd cell_6t
Xbit_r153_c44 bl[44] br[44] wl[153] vdd gnd cell_6t
Xbit_r154_c44 bl[44] br[44] wl[154] vdd gnd cell_6t
Xbit_r155_c44 bl[44] br[44] wl[155] vdd gnd cell_6t
Xbit_r156_c44 bl[44] br[44] wl[156] vdd gnd cell_6t
Xbit_r157_c44 bl[44] br[44] wl[157] vdd gnd cell_6t
Xbit_r158_c44 bl[44] br[44] wl[158] vdd gnd cell_6t
Xbit_r159_c44 bl[44] br[44] wl[159] vdd gnd cell_6t
Xbit_r160_c44 bl[44] br[44] wl[160] vdd gnd cell_6t
Xbit_r161_c44 bl[44] br[44] wl[161] vdd gnd cell_6t
Xbit_r162_c44 bl[44] br[44] wl[162] vdd gnd cell_6t
Xbit_r163_c44 bl[44] br[44] wl[163] vdd gnd cell_6t
Xbit_r164_c44 bl[44] br[44] wl[164] vdd gnd cell_6t
Xbit_r165_c44 bl[44] br[44] wl[165] vdd gnd cell_6t
Xbit_r166_c44 bl[44] br[44] wl[166] vdd gnd cell_6t
Xbit_r167_c44 bl[44] br[44] wl[167] vdd gnd cell_6t
Xbit_r168_c44 bl[44] br[44] wl[168] vdd gnd cell_6t
Xbit_r169_c44 bl[44] br[44] wl[169] vdd gnd cell_6t
Xbit_r170_c44 bl[44] br[44] wl[170] vdd gnd cell_6t
Xbit_r171_c44 bl[44] br[44] wl[171] vdd gnd cell_6t
Xbit_r172_c44 bl[44] br[44] wl[172] vdd gnd cell_6t
Xbit_r173_c44 bl[44] br[44] wl[173] vdd gnd cell_6t
Xbit_r174_c44 bl[44] br[44] wl[174] vdd gnd cell_6t
Xbit_r175_c44 bl[44] br[44] wl[175] vdd gnd cell_6t
Xbit_r176_c44 bl[44] br[44] wl[176] vdd gnd cell_6t
Xbit_r177_c44 bl[44] br[44] wl[177] vdd gnd cell_6t
Xbit_r178_c44 bl[44] br[44] wl[178] vdd gnd cell_6t
Xbit_r179_c44 bl[44] br[44] wl[179] vdd gnd cell_6t
Xbit_r180_c44 bl[44] br[44] wl[180] vdd gnd cell_6t
Xbit_r181_c44 bl[44] br[44] wl[181] vdd gnd cell_6t
Xbit_r182_c44 bl[44] br[44] wl[182] vdd gnd cell_6t
Xbit_r183_c44 bl[44] br[44] wl[183] vdd gnd cell_6t
Xbit_r184_c44 bl[44] br[44] wl[184] vdd gnd cell_6t
Xbit_r185_c44 bl[44] br[44] wl[185] vdd gnd cell_6t
Xbit_r186_c44 bl[44] br[44] wl[186] vdd gnd cell_6t
Xbit_r187_c44 bl[44] br[44] wl[187] vdd gnd cell_6t
Xbit_r188_c44 bl[44] br[44] wl[188] vdd gnd cell_6t
Xbit_r189_c44 bl[44] br[44] wl[189] vdd gnd cell_6t
Xbit_r190_c44 bl[44] br[44] wl[190] vdd gnd cell_6t
Xbit_r191_c44 bl[44] br[44] wl[191] vdd gnd cell_6t
Xbit_r192_c44 bl[44] br[44] wl[192] vdd gnd cell_6t
Xbit_r193_c44 bl[44] br[44] wl[193] vdd gnd cell_6t
Xbit_r194_c44 bl[44] br[44] wl[194] vdd gnd cell_6t
Xbit_r195_c44 bl[44] br[44] wl[195] vdd gnd cell_6t
Xbit_r196_c44 bl[44] br[44] wl[196] vdd gnd cell_6t
Xbit_r197_c44 bl[44] br[44] wl[197] vdd gnd cell_6t
Xbit_r198_c44 bl[44] br[44] wl[198] vdd gnd cell_6t
Xbit_r199_c44 bl[44] br[44] wl[199] vdd gnd cell_6t
Xbit_r200_c44 bl[44] br[44] wl[200] vdd gnd cell_6t
Xbit_r201_c44 bl[44] br[44] wl[201] vdd gnd cell_6t
Xbit_r202_c44 bl[44] br[44] wl[202] vdd gnd cell_6t
Xbit_r203_c44 bl[44] br[44] wl[203] vdd gnd cell_6t
Xbit_r204_c44 bl[44] br[44] wl[204] vdd gnd cell_6t
Xbit_r205_c44 bl[44] br[44] wl[205] vdd gnd cell_6t
Xbit_r206_c44 bl[44] br[44] wl[206] vdd gnd cell_6t
Xbit_r207_c44 bl[44] br[44] wl[207] vdd gnd cell_6t
Xbit_r208_c44 bl[44] br[44] wl[208] vdd gnd cell_6t
Xbit_r209_c44 bl[44] br[44] wl[209] vdd gnd cell_6t
Xbit_r210_c44 bl[44] br[44] wl[210] vdd gnd cell_6t
Xbit_r211_c44 bl[44] br[44] wl[211] vdd gnd cell_6t
Xbit_r212_c44 bl[44] br[44] wl[212] vdd gnd cell_6t
Xbit_r213_c44 bl[44] br[44] wl[213] vdd gnd cell_6t
Xbit_r214_c44 bl[44] br[44] wl[214] vdd gnd cell_6t
Xbit_r215_c44 bl[44] br[44] wl[215] vdd gnd cell_6t
Xbit_r216_c44 bl[44] br[44] wl[216] vdd gnd cell_6t
Xbit_r217_c44 bl[44] br[44] wl[217] vdd gnd cell_6t
Xbit_r218_c44 bl[44] br[44] wl[218] vdd gnd cell_6t
Xbit_r219_c44 bl[44] br[44] wl[219] vdd gnd cell_6t
Xbit_r220_c44 bl[44] br[44] wl[220] vdd gnd cell_6t
Xbit_r221_c44 bl[44] br[44] wl[221] vdd gnd cell_6t
Xbit_r222_c44 bl[44] br[44] wl[222] vdd gnd cell_6t
Xbit_r223_c44 bl[44] br[44] wl[223] vdd gnd cell_6t
Xbit_r224_c44 bl[44] br[44] wl[224] vdd gnd cell_6t
Xbit_r225_c44 bl[44] br[44] wl[225] vdd gnd cell_6t
Xbit_r226_c44 bl[44] br[44] wl[226] vdd gnd cell_6t
Xbit_r227_c44 bl[44] br[44] wl[227] vdd gnd cell_6t
Xbit_r228_c44 bl[44] br[44] wl[228] vdd gnd cell_6t
Xbit_r229_c44 bl[44] br[44] wl[229] vdd gnd cell_6t
Xbit_r230_c44 bl[44] br[44] wl[230] vdd gnd cell_6t
Xbit_r231_c44 bl[44] br[44] wl[231] vdd gnd cell_6t
Xbit_r232_c44 bl[44] br[44] wl[232] vdd gnd cell_6t
Xbit_r233_c44 bl[44] br[44] wl[233] vdd gnd cell_6t
Xbit_r234_c44 bl[44] br[44] wl[234] vdd gnd cell_6t
Xbit_r235_c44 bl[44] br[44] wl[235] vdd gnd cell_6t
Xbit_r236_c44 bl[44] br[44] wl[236] vdd gnd cell_6t
Xbit_r237_c44 bl[44] br[44] wl[237] vdd gnd cell_6t
Xbit_r238_c44 bl[44] br[44] wl[238] vdd gnd cell_6t
Xbit_r239_c44 bl[44] br[44] wl[239] vdd gnd cell_6t
Xbit_r240_c44 bl[44] br[44] wl[240] vdd gnd cell_6t
Xbit_r241_c44 bl[44] br[44] wl[241] vdd gnd cell_6t
Xbit_r242_c44 bl[44] br[44] wl[242] vdd gnd cell_6t
Xbit_r243_c44 bl[44] br[44] wl[243] vdd gnd cell_6t
Xbit_r244_c44 bl[44] br[44] wl[244] vdd gnd cell_6t
Xbit_r245_c44 bl[44] br[44] wl[245] vdd gnd cell_6t
Xbit_r246_c44 bl[44] br[44] wl[246] vdd gnd cell_6t
Xbit_r247_c44 bl[44] br[44] wl[247] vdd gnd cell_6t
Xbit_r248_c44 bl[44] br[44] wl[248] vdd gnd cell_6t
Xbit_r249_c44 bl[44] br[44] wl[249] vdd gnd cell_6t
Xbit_r250_c44 bl[44] br[44] wl[250] vdd gnd cell_6t
Xbit_r251_c44 bl[44] br[44] wl[251] vdd gnd cell_6t
Xbit_r252_c44 bl[44] br[44] wl[252] vdd gnd cell_6t
Xbit_r253_c44 bl[44] br[44] wl[253] vdd gnd cell_6t
Xbit_r254_c44 bl[44] br[44] wl[254] vdd gnd cell_6t
Xbit_r255_c44 bl[44] br[44] wl[255] vdd gnd cell_6t
Xbit_r0_c45 bl[45] br[45] wl[0] vdd gnd cell_6t
Xbit_r1_c45 bl[45] br[45] wl[1] vdd gnd cell_6t
Xbit_r2_c45 bl[45] br[45] wl[2] vdd gnd cell_6t
Xbit_r3_c45 bl[45] br[45] wl[3] vdd gnd cell_6t
Xbit_r4_c45 bl[45] br[45] wl[4] vdd gnd cell_6t
Xbit_r5_c45 bl[45] br[45] wl[5] vdd gnd cell_6t
Xbit_r6_c45 bl[45] br[45] wl[6] vdd gnd cell_6t
Xbit_r7_c45 bl[45] br[45] wl[7] vdd gnd cell_6t
Xbit_r8_c45 bl[45] br[45] wl[8] vdd gnd cell_6t
Xbit_r9_c45 bl[45] br[45] wl[9] vdd gnd cell_6t
Xbit_r10_c45 bl[45] br[45] wl[10] vdd gnd cell_6t
Xbit_r11_c45 bl[45] br[45] wl[11] vdd gnd cell_6t
Xbit_r12_c45 bl[45] br[45] wl[12] vdd gnd cell_6t
Xbit_r13_c45 bl[45] br[45] wl[13] vdd gnd cell_6t
Xbit_r14_c45 bl[45] br[45] wl[14] vdd gnd cell_6t
Xbit_r15_c45 bl[45] br[45] wl[15] vdd gnd cell_6t
Xbit_r16_c45 bl[45] br[45] wl[16] vdd gnd cell_6t
Xbit_r17_c45 bl[45] br[45] wl[17] vdd gnd cell_6t
Xbit_r18_c45 bl[45] br[45] wl[18] vdd gnd cell_6t
Xbit_r19_c45 bl[45] br[45] wl[19] vdd gnd cell_6t
Xbit_r20_c45 bl[45] br[45] wl[20] vdd gnd cell_6t
Xbit_r21_c45 bl[45] br[45] wl[21] vdd gnd cell_6t
Xbit_r22_c45 bl[45] br[45] wl[22] vdd gnd cell_6t
Xbit_r23_c45 bl[45] br[45] wl[23] vdd gnd cell_6t
Xbit_r24_c45 bl[45] br[45] wl[24] vdd gnd cell_6t
Xbit_r25_c45 bl[45] br[45] wl[25] vdd gnd cell_6t
Xbit_r26_c45 bl[45] br[45] wl[26] vdd gnd cell_6t
Xbit_r27_c45 bl[45] br[45] wl[27] vdd gnd cell_6t
Xbit_r28_c45 bl[45] br[45] wl[28] vdd gnd cell_6t
Xbit_r29_c45 bl[45] br[45] wl[29] vdd gnd cell_6t
Xbit_r30_c45 bl[45] br[45] wl[30] vdd gnd cell_6t
Xbit_r31_c45 bl[45] br[45] wl[31] vdd gnd cell_6t
Xbit_r32_c45 bl[45] br[45] wl[32] vdd gnd cell_6t
Xbit_r33_c45 bl[45] br[45] wl[33] vdd gnd cell_6t
Xbit_r34_c45 bl[45] br[45] wl[34] vdd gnd cell_6t
Xbit_r35_c45 bl[45] br[45] wl[35] vdd gnd cell_6t
Xbit_r36_c45 bl[45] br[45] wl[36] vdd gnd cell_6t
Xbit_r37_c45 bl[45] br[45] wl[37] vdd gnd cell_6t
Xbit_r38_c45 bl[45] br[45] wl[38] vdd gnd cell_6t
Xbit_r39_c45 bl[45] br[45] wl[39] vdd gnd cell_6t
Xbit_r40_c45 bl[45] br[45] wl[40] vdd gnd cell_6t
Xbit_r41_c45 bl[45] br[45] wl[41] vdd gnd cell_6t
Xbit_r42_c45 bl[45] br[45] wl[42] vdd gnd cell_6t
Xbit_r43_c45 bl[45] br[45] wl[43] vdd gnd cell_6t
Xbit_r44_c45 bl[45] br[45] wl[44] vdd gnd cell_6t
Xbit_r45_c45 bl[45] br[45] wl[45] vdd gnd cell_6t
Xbit_r46_c45 bl[45] br[45] wl[46] vdd gnd cell_6t
Xbit_r47_c45 bl[45] br[45] wl[47] vdd gnd cell_6t
Xbit_r48_c45 bl[45] br[45] wl[48] vdd gnd cell_6t
Xbit_r49_c45 bl[45] br[45] wl[49] vdd gnd cell_6t
Xbit_r50_c45 bl[45] br[45] wl[50] vdd gnd cell_6t
Xbit_r51_c45 bl[45] br[45] wl[51] vdd gnd cell_6t
Xbit_r52_c45 bl[45] br[45] wl[52] vdd gnd cell_6t
Xbit_r53_c45 bl[45] br[45] wl[53] vdd gnd cell_6t
Xbit_r54_c45 bl[45] br[45] wl[54] vdd gnd cell_6t
Xbit_r55_c45 bl[45] br[45] wl[55] vdd gnd cell_6t
Xbit_r56_c45 bl[45] br[45] wl[56] vdd gnd cell_6t
Xbit_r57_c45 bl[45] br[45] wl[57] vdd gnd cell_6t
Xbit_r58_c45 bl[45] br[45] wl[58] vdd gnd cell_6t
Xbit_r59_c45 bl[45] br[45] wl[59] vdd gnd cell_6t
Xbit_r60_c45 bl[45] br[45] wl[60] vdd gnd cell_6t
Xbit_r61_c45 bl[45] br[45] wl[61] vdd gnd cell_6t
Xbit_r62_c45 bl[45] br[45] wl[62] vdd gnd cell_6t
Xbit_r63_c45 bl[45] br[45] wl[63] vdd gnd cell_6t
Xbit_r64_c45 bl[45] br[45] wl[64] vdd gnd cell_6t
Xbit_r65_c45 bl[45] br[45] wl[65] vdd gnd cell_6t
Xbit_r66_c45 bl[45] br[45] wl[66] vdd gnd cell_6t
Xbit_r67_c45 bl[45] br[45] wl[67] vdd gnd cell_6t
Xbit_r68_c45 bl[45] br[45] wl[68] vdd gnd cell_6t
Xbit_r69_c45 bl[45] br[45] wl[69] vdd gnd cell_6t
Xbit_r70_c45 bl[45] br[45] wl[70] vdd gnd cell_6t
Xbit_r71_c45 bl[45] br[45] wl[71] vdd gnd cell_6t
Xbit_r72_c45 bl[45] br[45] wl[72] vdd gnd cell_6t
Xbit_r73_c45 bl[45] br[45] wl[73] vdd gnd cell_6t
Xbit_r74_c45 bl[45] br[45] wl[74] vdd gnd cell_6t
Xbit_r75_c45 bl[45] br[45] wl[75] vdd gnd cell_6t
Xbit_r76_c45 bl[45] br[45] wl[76] vdd gnd cell_6t
Xbit_r77_c45 bl[45] br[45] wl[77] vdd gnd cell_6t
Xbit_r78_c45 bl[45] br[45] wl[78] vdd gnd cell_6t
Xbit_r79_c45 bl[45] br[45] wl[79] vdd gnd cell_6t
Xbit_r80_c45 bl[45] br[45] wl[80] vdd gnd cell_6t
Xbit_r81_c45 bl[45] br[45] wl[81] vdd gnd cell_6t
Xbit_r82_c45 bl[45] br[45] wl[82] vdd gnd cell_6t
Xbit_r83_c45 bl[45] br[45] wl[83] vdd gnd cell_6t
Xbit_r84_c45 bl[45] br[45] wl[84] vdd gnd cell_6t
Xbit_r85_c45 bl[45] br[45] wl[85] vdd gnd cell_6t
Xbit_r86_c45 bl[45] br[45] wl[86] vdd gnd cell_6t
Xbit_r87_c45 bl[45] br[45] wl[87] vdd gnd cell_6t
Xbit_r88_c45 bl[45] br[45] wl[88] vdd gnd cell_6t
Xbit_r89_c45 bl[45] br[45] wl[89] vdd gnd cell_6t
Xbit_r90_c45 bl[45] br[45] wl[90] vdd gnd cell_6t
Xbit_r91_c45 bl[45] br[45] wl[91] vdd gnd cell_6t
Xbit_r92_c45 bl[45] br[45] wl[92] vdd gnd cell_6t
Xbit_r93_c45 bl[45] br[45] wl[93] vdd gnd cell_6t
Xbit_r94_c45 bl[45] br[45] wl[94] vdd gnd cell_6t
Xbit_r95_c45 bl[45] br[45] wl[95] vdd gnd cell_6t
Xbit_r96_c45 bl[45] br[45] wl[96] vdd gnd cell_6t
Xbit_r97_c45 bl[45] br[45] wl[97] vdd gnd cell_6t
Xbit_r98_c45 bl[45] br[45] wl[98] vdd gnd cell_6t
Xbit_r99_c45 bl[45] br[45] wl[99] vdd gnd cell_6t
Xbit_r100_c45 bl[45] br[45] wl[100] vdd gnd cell_6t
Xbit_r101_c45 bl[45] br[45] wl[101] vdd gnd cell_6t
Xbit_r102_c45 bl[45] br[45] wl[102] vdd gnd cell_6t
Xbit_r103_c45 bl[45] br[45] wl[103] vdd gnd cell_6t
Xbit_r104_c45 bl[45] br[45] wl[104] vdd gnd cell_6t
Xbit_r105_c45 bl[45] br[45] wl[105] vdd gnd cell_6t
Xbit_r106_c45 bl[45] br[45] wl[106] vdd gnd cell_6t
Xbit_r107_c45 bl[45] br[45] wl[107] vdd gnd cell_6t
Xbit_r108_c45 bl[45] br[45] wl[108] vdd gnd cell_6t
Xbit_r109_c45 bl[45] br[45] wl[109] vdd gnd cell_6t
Xbit_r110_c45 bl[45] br[45] wl[110] vdd gnd cell_6t
Xbit_r111_c45 bl[45] br[45] wl[111] vdd gnd cell_6t
Xbit_r112_c45 bl[45] br[45] wl[112] vdd gnd cell_6t
Xbit_r113_c45 bl[45] br[45] wl[113] vdd gnd cell_6t
Xbit_r114_c45 bl[45] br[45] wl[114] vdd gnd cell_6t
Xbit_r115_c45 bl[45] br[45] wl[115] vdd gnd cell_6t
Xbit_r116_c45 bl[45] br[45] wl[116] vdd gnd cell_6t
Xbit_r117_c45 bl[45] br[45] wl[117] vdd gnd cell_6t
Xbit_r118_c45 bl[45] br[45] wl[118] vdd gnd cell_6t
Xbit_r119_c45 bl[45] br[45] wl[119] vdd gnd cell_6t
Xbit_r120_c45 bl[45] br[45] wl[120] vdd gnd cell_6t
Xbit_r121_c45 bl[45] br[45] wl[121] vdd gnd cell_6t
Xbit_r122_c45 bl[45] br[45] wl[122] vdd gnd cell_6t
Xbit_r123_c45 bl[45] br[45] wl[123] vdd gnd cell_6t
Xbit_r124_c45 bl[45] br[45] wl[124] vdd gnd cell_6t
Xbit_r125_c45 bl[45] br[45] wl[125] vdd gnd cell_6t
Xbit_r126_c45 bl[45] br[45] wl[126] vdd gnd cell_6t
Xbit_r127_c45 bl[45] br[45] wl[127] vdd gnd cell_6t
Xbit_r128_c45 bl[45] br[45] wl[128] vdd gnd cell_6t
Xbit_r129_c45 bl[45] br[45] wl[129] vdd gnd cell_6t
Xbit_r130_c45 bl[45] br[45] wl[130] vdd gnd cell_6t
Xbit_r131_c45 bl[45] br[45] wl[131] vdd gnd cell_6t
Xbit_r132_c45 bl[45] br[45] wl[132] vdd gnd cell_6t
Xbit_r133_c45 bl[45] br[45] wl[133] vdd gnd cell_6t
Xbit_r134_c45 bl[45] br[45] wl[134] vdd gnd cell_6t
Xbit_r135_c45 bl[45] br[45] wl[135] vdd gnd cell_6t
Xbit_r136_c45 bl[45] br[45] wl[136] vdd gnd cell_6t
Xbit_r137_c45 bl[45] br[45] wl[137] vdd gnd cell_6t
Xbit_r138_c45 bl[45] br[45] wl[138] vdd gnd cell_6t
Xbit_r139_c45 bl[45] br[45] wl[139] vdd gnd cell_6t
Xbit_r140_c45 bl[45] br[45] wl[140] vdd gnd cell_6t
Xbit_r141_c45 bl[45] br[45] wl[141] vdd gnd cell_6t
Xbit_r142_c45 bl[45] br[45] wl[142] vdd gnd cell_6t
Xbit_r143_c45 bl[45] br[45] wl[143] vdd gnd cell_6t
Xbit_r144_c45 bl[45] br[45] wl[144] vdd gnd cell_6t
Xbit_r145_c45 bl[45] br[45] wl[145] vdd gnd cell_6t
Xbit_r146_c45 bl[45] br[45] wl[146] vdd gnd cell_6t
Xbit_r147_c45 bl[45] br[45] wl[147] vdd gnd cell_6t
Xbit_r148_c45 bl[45] br[45] wl[148] vdd gnd cell_6t
Xbit_r149_c45 bl[45] br[45] wl[149] vdd gnd cell_6t
Xbit_r150_c45 bl[45] br[45] wl[150] vdd gnd cell_6t
Xbit_r151_c45 bl[45] br[45] wl[151] vdd gnd cell_6t
Xbit_r152_c45 bl[45] br[45] wl[152] vdd gnd cell_6t
Xbit_r153_c45 bl[45] br[45] wl[153] vdd gnd cell_6t
Xbit_r154_c45 bl[45] br[45] wl[154] vdd gnd cell_6t
Xbit_r155_c45 bl[45] br[45] wl[155] vdd gnd cell_6t
Xbit_r156_c45 bl[45] br[45] wl[156] vdd gnd cell_6t
Xbit_r157_c45 bl[45] br[45] wl[157] vdd gnd cell_6t
Xbit_r158_c45 bl[45] br[45] wl[158] vdd gnd cell_6t
Xbit_r159_c45 bl[45] br[45] wl[159] vdd gnd cell_6t
Xbit_r160_c45 bl[45] br[45] wl[160] vdd gnd cell_6t
Xbit_r161_c45 bl[45] br[45] wl[161] vdd gnd cell_6t
Xbit_r162_c45 bl[45] br[45] wl[162] vdd gnd cell_6t
Xbit_r163_c45 bl[45] br[45] wl[163] vdd gnd cell_6t
Xbit_r164_c45 bl[45] br[45] wl[164] vdd gnd cell_6t
Xbit_r165_c45 bl[45] br[45] wl[165] vdd gnd cell_6t
Xbit_r166_c45 bl[45] br[45] wl[166] vdd gnd cell_6t
Xbit_r167_c45 bl[45] br[45] wl[167] vdd gnd cell_6t
Xbit_r168_c45 bl[45] br[45] wl[168] vdd gnd cell_6t
Xbit_r169_c45 bl[45] br[45] wl[169] vdd gnd cell_6t
Xbit_r170_c45 bl[45] br[45] wl[170] vdd gnd cell_6t
Xbit_r171_c45 bl[45] br[45] wl[171] vdd gnd cell_6t
Xbit_r172_c45 bl[45] br[45] wl[172] vdd gnd cell_6t
Xbit_r173_c45 bl[45] br[45] wl[173] vdd gnd cell_6t
Xbit_r174_c45 bl[45] br[45] wl[174] vdd gnd cell_6t
Xbit_r175_c45 bl[45] br[45] wl[175] vdd gnd cell_6t
Xbit_r176_c45 bl[45] br[45] wl[176] vdd gnd cell_6t
Xbit_r177_c45 bl[45] br[45] wl[177] vdd gnd cell_6t
Xbit_r178_c45 bl[45] br[45] wl[178] vdd gnd cell_6t
Xbit_r179_c45 bl[45] br[45] wl[179] vdd gnd cell_6t
Xbit_r180_c45 bl[45] br[45] wl[180] vdd gnd cell_6t
Xbit_r181_c45 bl[45] br[45] wl[181] vdd gnd cell_6t
Xbit_r182_c45 bl[45] br[45] wl[182] vdd gnd cell_6t
Xbit_r183_c45 bl[45] br[45] wl[183] vdd gnd cell_6t
Xbit_r184_c45 bl[45] br[45] wl[184] vdd gnd cell_6t
Xbit_r185_c45 bl[45] br[45] wl[185] vdd gnd cell_6t
Xbit_r186_c45 bl[45] br[45] wl[186] vdd gnd cell_6t
Xbit_r187_c45 bl[45] br[45] wl[187] vdd gnd cell_6t
Xbit_r188_c45 bl[45] br[45] wl[188] vdd gnd cell_6t
Xbit_r189_c45 bl[45] br[45] wl[189] vdd gnd cell_6t
Xbit_r190_c45 bl[45] br[45] wl[190] vdd gnd cell_6t
Xbit_r191_c45 bl[45] br[45] wl[191] vdd gnd cell_6t
Xbit_r192_c45 bl[45] br[45] wl[192] vdd gnd cell_6t
Xbit_r193_c45 bl[45] br[45] wl[193] vdd gnd cell_6t
Xbit_r194_c45 bl[45] br[45] wl[194] vdd gnd cell_6t
Xbit_r195_c45 bl[45] br[45] wl[195] vdd gnd cell_6t
Xbit_r196_c45 bl[45] br[45] wl[196] vdd gnd cell_6t
Xbit_r197_c45 bl[45] br[45] wl[197] vdd gnd cell_6t
Xbit_r198_c45 bl[45] br[45] wl[198] vdd gnd cell_6t
Xbit_r199_c45 bl[45] br[45] wl[199] vdd gnd cell_6t
Xbit_r200_c45 bl[45] br[45] wl[200] vdd gnd cell_6t
Xbit_r201_c45 bl[45] br[45] wl[201] vdd gnd cell_6t
Xbit_r202_c45 bl[45] br[45] wl[202] vdd gnd cell_6t
Xbit_r203_c45 bl[45] br[45] wl[203] vdd gnd cell_6t
Xbit_r204_c45 bl[45] br[45] wl[204] vdd gnd cell_6t
Xbit_r205_c45 bl[45] br[45] wl[205] vdd gnd cell_6t
Xbit_r206_c45 bl[45] br[45] wl[206] vdd gnd cell_6t
Xbit_r207_c45 bl[45] br[45] wl[207] vdd gnd cell_6t
Xbit_r208_c45 bl[45] br[45] wl[208] vdd gnd cell_6t
Xbit_r209_c45 bl[45] br[45] wl[209] vdd gnd cell_6t
Xbit_r210_c45 bl[45] br[45] wl[210] vdd gnd cell_6t
Xbit_r211_c45 bl[45] br[45] wl[211] vdd gnd cell_6t
Xbit_r212_c45 bl[45] br[45] wl[212] vdd gnd cell_6t
Xbit_r213_c45 bl[45] br[45] wl[213] vdd gnd cell_6t
Xbit_r214_c45 bl[45] br[45] wl[214] vdd gnd cell_6t
Xbit_r215_c45 bl[45] br[45] wl[215] vdd gnd cell_6t
Xbit_r216_c45 bl[45] br[45] wl[216] vdd gnd cell_6t
Xbit_r217_c45 bl[45] br[45] wl[217] vdd gnd cell_6t
Xbit_r218_c45 bl[45] br[45] wl[218] vdd gnd cell_6t
Xbit_r219_c45 bl[45] br[45] wl[219] vdd gnd cell_6t
Xbit_r220_c45 bl[45] br[45] wl[220] vdd gnd cell_6t
Xbit_r221_c45 bl[45] br[45] wl[221] vdd gnd cell_6t
Xbit_r222_c45 bl[45] br[45] wl[222] vdd gnd cell_6t
Xbit_r223_c45 bl[45] br[45] wl[223] vdd gnd cell_6t
Xbit_r224_c45 bl[45] br[45] wl[224] vdd gnd cell_6t
Xbit_r225_c45 bl[45] br[45] wl[225] vdd gnd cell_6t
Xbit_r226_c45 bl[45] br[45] wl[226] vdd gnd cell_6t
Xbit_r227_c45 bl[45] br[45] wl[227] vdd gnd cell_6t
Xbit_r228_c45 bl[45] br[45] wl[228] vdd gnd cell_6t
Xbit_r229_c45 bl[45] br[45] wl[229] vdd gnd cell_6t
Xbit_r230_c45 bl[45] br[45] wl[230] vdd gnd cell_6t
Xbit_r231_c45 bl[45] br[45] wl[231] vdd gnd cell_6t
Xbit_r232_c45 bl[45] br[45] wl[232] vdd gnd cell_6t
Xbit_r233_c45 bl[45] br[45] wl[233] vdd gnd cell_6t
Xbit_r234_c45 bl[45] br[45] wl[234] vdd gnd cell_6t
Xbit_r235_c45 bl[45] br[45] wl[235] vdd gnd cell_6t
Xbit_r236_c45 bl[45] br[45] wl[236] vdd gnd cell_6t
Xbit_r237_c45 bl[45] br[45] wl[237] vdd gnd cell_6t
Xbit_r238_c45 bl[45] br[45] wl[238] vdd gnd cell_6t
Xbit_r239_c45 bl[45] br[45] wl[239] vdd gnd cell_6t
Xbit_r240_c45 bl[45] br[45] wl[240] vdd gnd cell_6t
Xbit_r241_c45 bl[45] br[45] wl[241] vdd gnd cell_6t
Xbit_r242_c45 bl[45] br[45] wl[242] vdd gnd cell_6t
Xbit_r243_c45 bl[45] br[45] wl[243] vdd gnd cell_6t
Xbit_r244_c45 bl[45] br[45] wl[244] vdd gnd cell_6t
Xbit_r245_c45 bl[45] br[45] wl[245] vdd gnd cell_6t
Xbit_r246_c45 bl[45] br[45] wl[246] vdd gnd cell_6t
Xbit_r247_c45 bl[45] br[45] wl[247] vdd gnd cell_6t
Xbit_r248_c45 bl[45] br[45] wl[248] vdd gnd cell_6t
Xbit_r249_c45 bl[45] br[45] wl[249] vdd gnd cell_6t
Xbit_r250_c45 bl[45] br[45] wl[250] vdd gnd cell_6t
Xbit_r251_c45 bl[45] br[45] wl[251] vdd gnd cell_6t
Xbit_r252_c45 bl[45] br[45] wl[252] vdd gnd cell_6t
Xbit_r253_c45 bl[45] br[45] wl[253] vdd gnd cell_6t
Xbit_r254_c45 bl[45] br[45] wl[254] vdd gnd cell_6t
Xbit_r255_c45 bl[45] br[45] wl[255] vdd gnd cell_6t
Xbit_r0_c46 bl[46] br[46] wl[0] vdd gnd cell_6t
Xbit_r1_c46 bl[46] br[46] wl[1] vdd gnd cell_6t
Xbit_r2_c46 bl[46] br[46] wl[2] vdd gnd cell_6t
Xbit_r3_c46 bl[46] br[46] wl[3] vdd gnd cell_6t
Xbit_r4_c46 bl[46] br[46] wl[4] vdd gnd cell_6t
Xbit_r5_c46 bl[46] br[46] wl[5] vdd gnd cell_6t
Xbit_r6_c46 bl[46] br[46] wl[6] vdd gnd cell_6t
Xbit_r7_c46 bl[46] br[46] wl[7] vdd gnd cell_6t
Xbit_r8_c46 bl[46] br[46] wl[8] vdd gnd cell_6t
Xbit_r9_c46 bl[46] br[46] wl[9] vdd gnd cell_6t
Xbit_r10_c46 bl[46] br[46] wl[10] vdd gnd cell_6t
Xbit_r11_c46 bl[46] br[46] wl[11] vdd gnd cell_6t
Xbit_r12_c46 bl[46] br[46] wl[12] vdd gnd cell_6t
Xbit_r13_c46 bl[46] br[46] wl[13] vdd gnd cell_6t
Xbit_r14_c46 bl[46] br[46] wl[14] vdd gnd cell_6t
Xbit_r15_c46 bl[46] br[46] wl[15] vdd gnd cell_6t
Xbit_r16_c46 bl[46] br[46] wl[16] vdd gnd cell_6t
Xbit_r17_c46 bl[46] br[46] wl[17] vdd gnd cell_6t
Xbit_r18_c46 bl[46] br[46] wl[18] vdd gnd cell_6t
Xbit_r19_c46 bl[46] br[46] wl[19] vdd gnd cell_6t
Xbit_r20_c46 bl[46] br[46] wl[20] vdd gnd cell_6t
Xbit_r21_c46 bl[46] br[46] wl[21] vdd gnd cell_6t
Xbit_r22_c46 bl[46] br[46] wl[22] vdd gnd cell_6t
Xbit_r23_c46 bl[46] br[46] wl[23] vdd gnd cell_6t
Xbit_r24_c46 bl[46] br[46] wl[24] vdd gnd cell_6t
Xbit_r25_c46 bl[46] br[46] wl[25] vdd gnd cell_6t
Xbit_r26_c46 bl[46] br[46] wl[26] vdd gnd cell_6t
Xbit_r27_c46 bl[46] br[46] wl[27] vdd gnd cell_6t
Xbit_r28_c46 bl[46] br[46] wl[28] vdd gnd cell_6t
Xbit_r29_c46 bl[46] br[46] wl[29] vdd gnd cell_6t
Xbit_r30_c46 bl[46] br[46] wl[30] vdd gnd cell_6t
Xbit_r31_c46 bl[46] br[46] wl[31] vdd gnd cell_6t
Xbit_r32_c46 bl[46] br[46] wl[32] vdd gnd cell_6t
Xbit_r33_c46 bl[46] br[46] wl[33] vdd gnd cell_6t
Xbit_r34_c46 bl[46] br[46] wl[34] vdd gnd cell_6t
Xbit_r35_c46 bl[46] br[46] wl[35] vdd gnd cell_6t
Xbit_r36_c46 bl[46] br[46] wl[36] vdd gnd cell_6t
Xbit_r37_c46 bl[46] br[46] wl[37] vdd gnd cell_6t
Xbit_r38_c46 bl[46] br[46] wl[38] vdd gnd cell_6t
Xbit_r39_c46 bl[46] br[46] wl[39] vdd gnd cell_6t
Xbit_r40_c46 bl[46] br[46] wl[40] vdd gnd cell_6t
Xbit_r41_c46 bl[46] br[46] wl[41] vdd gnd cell_6t
Xbit_r42_c46 bl[46] br[46] wl[42] vdd gnd cell_6t
Xbit_r43_c46 bl[46] br[46] wl[43] vdd gnd cell_6t
Xbit_r44_c46 bl[46] br[46] wl[44] vdd gnd cell_6t
Xbit_r45_c46 bl[46] br[46] wl[45] vdd gnd cell_6t
Xbit_r46_c46 bl[46] br[46] wl[46] vdd gnd cell_6t
Xbit_r47_c46 bl[46] br[46] wl[47] vdd gnd cell_6t
Xbit_r48_c46 bl[46] br[46] wl[48] vdd gnd cell_6t
Xbit_r49_c46 bl[46] br[46] wl[49] vdd gnd cell_6t
Xbit_r50_c46 bl[46] br[46] wl[50] vdd gnd cell_6t
Xbit_r51_c46 bl[46] br[46] wl[51] vdd gnd cell_6t
Xbit_r52_c46 bl[46] br[46] wl[52] vdd gnd cell_6t
Xbit_r53_c46 bl[46] br[46] wl[53] vdd gnd cell_6t
Xbit_r54_c46 bl[46] br[46] wl[54] vdd gnd cell_6t
Xbit_r55_c46 bl[46] br[46] wl[55] vdd gnd cell_6t
Xbit_r56_c46 bl[46] br[46] wl[56] vdd gnd cell_6t
Xbit_r57_c46 bl[46] br[46] wl[57] vdd gnd cell_6t
Xbit_r58_c46 bl[46] br[46] wl[58] vdd gnd cell_6t
Xbit_r59_c46 bl[46] br[46] wl[59] vdd gnd cell_6t
Xbit_r60_c46 bl[46] br[46] wl[60] vdd gnd cell_6t
Xbit_r61_c46 bl[46] br[46] wl[61] vdd gnd cell_6t
Xbit_r62_c46 bl[46] br[46] wl[62] vdd gnd cell_6t
Xbit_r63_c46 bl[46] br[46] wl[63] vdd gnd cell_6t
Xbit_r64_c46 bl[46] br[46] wl[64] vdd gnd cell_6t
Xbit_r65_c46 bl[46] br[46] wl[65] vdd gnd cell_6t
Xbit_r66_c46 bl[46] br[46] wl[66] vdd gnd cell_6t
Xbit_r67_c46 bl[46] br[46] wl[67] vdd gnd cell_6t
Xbit_r68_c46 bl[46] br[46] wl[68] vdd gnd cell_6t
Xbit_r69_c46 bl[46] br[46] wl[69] vdd gnd cell_6t
Xbit_r70_c46 bl[46] br[46] wl[70] vdd gnd cell_6t
Xbit_r71_c46 bl[46] br[46] wl[71] vdd gnd cell_6t
Xbit_r72_c46 bl[46] br[46] wl[72] vdd gnd cell_6t
Xbit_r73_c46 bl[46] br[46] wl[73] vdd gnd cell_6t
Xbit_r74_c46 bl[46] br[46] wl[74] vdd gnd cell_6t
Xbit_r75_c46 bl[46] br[46] wl[75] vdd gnd cell_6t
Xbit_r76_c46 bl[46] br[46] wl[76] vdd gnd cell_6t
Xbit_r77_c46 bl[46] br[46] wl[77] vdd gnd cell_6t
Xbit_r78_c46 bl[46] br[46] wl[78] vdd gnd cell_6t
Xbit_r79_c46 bl[46] br[46] wl[79] vdd gnd cell_6t
Xbit_r80_c46 bl[46] br[46] wl[80] vdd gnd cell_6t
Xbit_r81_c46 bl[46] br[46] wl[81] vdd gnd cell_6t
Xbit_r82_c46 bl[46] br[46] wl[82] vdd gnd cell_6t
Xbit_r83_c46 bl[46] br[46] wl[83] vdd gnd cell_6t
Xbit_r84_c46 bl[46] br[46] wl[84] vdd gnd cell_6t
Xbit_r85_c46 bl[46] br[46] wl[85] vdd gnd cell_6t
Xbit_r86_c46 bl[46] br[46] wl[86] vdd gnd cell_6t
Xbit_r87_c46 bl[46] br[46] wl[87] vdd gnd cell_6t
Xbit_r88_c46 bl[46] br[46] wl[88] vdd gnd cell_6t
Xbit_r89_c46 bl[46] br[46] wl[89] vdd gnd cell_6t
Xbit_r90_c46 bl[46] br[46] wl[90] vdd gnd cell_6t
Xbit_r91_c46 bl[46] br[46] wl[91] vdd gnd cell_6t
Xbit_r92_c46 bl[46] br[46] wl[92] vdd gnd cell_6t
Xbit_r93_c46 bl[46] br[46] wl[93] vdd gnd cell_6t
Xbit_r94_c46 bl[46] br[46] wl[94] vdd gnd cell_6t
Xbit_r95_c46 bl[46] br[46] wl[95] vdd gnd cell_6t
Xbit_r96_c46 bl[46] br[46] wl[96] vdd gnd cell_6t
Xbit_r97_c46 bl[46] br[46] wl[97] vdd gnd cell_6t
Xbit_r98_c46 bl[46] br[46] wl[98] vdd gnd cell_6t
Xbit_r99_c46 bl[46] br[46] wl[99] vdd gnd cell_6t
Xbit_r100_c46 bl[46] br[46] wl[100] vdd gnd cell_6t
Xbit_r101_c46 bl[46] br[46] wl[101] vdd gnd cell_6t
Xbit_r102_c46 bl[46] br[46] wl[102] vdd gnd cell_6t
Xbit_r103_c46 bl[46] br[46] wl[103] vdd gnd cell_6t
Xbit_r104_c46 bl[46] br[46] wl[104] vdd gnd cell_6t
Xbit_r105_c46 bl[46] br[46] wl[105] vdd gnd cell_6t
Xbit_r106_c46 bl[46] br[46] wl[106] vdd gnd cell_6t
Xbit_r107_c46 bl[46] br[46] wl[107] vdd gnd cell_6t
Xbit_r108_c46 bl[46] br[46] wl[108] vdd gnd cell_6t
Xbit_r109_c46 bl[46] br[46] wl[109] vdd gnd cell_6t
Xbit_r110_c46 bl[46] br[46] wl[110] vdd gnd cell_6t
Xbit_r111_c46 bl[46] br[46] wl[111] vdd gnd cell_6t
Xbit_r112_c46 bl[46] br[46] wl[112] vdd gnd cell_6t
Xbit_r113_c46 bl[46] br[46] wl[113] vdd gnd cell_6t
Xbit_r114_c46 bl[46] br[46] wl[114] vdd gnd cell_6t
Xbit_r115_c46 bl[46] br[46] wl[115] vdd gnd cell_6t
Xbit_r116_c46 bl[46] br[46] wl[116] vdd gnd cell_6t
Xbit_r117_c46 bl[46] br[46] wl[117] vdd gnd cell_6t
Xbit_r118_c46 bl[46] br[46] wl[118] vdd gnd cell_6t
Xbit_r119_c46 bl[46] br[46] wl[119] vdd gnd cell_6t
Xbit_r120_c46 bl[46] br[46] wl[120] vdd gnd cell_6t
Xbit_r121_c46 bl[46] br[46] wl[121] vdd gnd cell_6t
Xbit_r122_c46 bl[46] br[46] wl[122] vdd gnd cell_6t
Xbit_r123_c46 bl[46] br[46] wl[123] vdd gnd cell_6t
Xbit_r124_c46 bl[46] br[46] wl[124] vdd gnd cell_6t
Xbit_r125_c46 bl[46] br[46] wl[125] vdd gnd cell_6t
Xbit_r126_c46 bl[46] br[46] wl[126] vdd gnd cell_6t
Xbit_r127_c46 bl[46] br[46] wl[127] vdd gnd cell_6t
Xbit_r128_c46 bl[46] br[46] wl[128] vdd gnd cell_6t
Xbit_r129_c46 bl[46] br[46] wl[129] vdd gnd cell_6t
Xbit_r130_c46 bl[46] br[46] wl[130] vdd gnd cell_6t
Xbit_r131_c46 bl[46] br[46] wl[131] vdd gnd cell_6t
Xbit_r132_c46 bl[46] br[46] wl[132] vdd gnd cell_6t
Xbit_r133_c46 bl[46] br[46] wl[133] vdd gnd cell_6t
Xbit_r134_c46 bl[46] br[46] wl[134] vdd gnd cell_6t
Xbit_r135_c46 bl[46] br[46] wl[135] vdd gnd cell_6t
Xbit_r136_c46 bl[46] br[46] wl[136] vdd gnd cell_6t
Xbit_r137_c46 bl[46] br[46] wl[137] vdd gnd cell_6t
Xbit_r138_c46 bl[46] br[46] wl[138] vdd gnd cell_6t
Xbit_r139_c46 bl[46] br[46] wl[139] vdd gnd cell_6t
Xbit_r140_c46 bl[46] br[46] wl[140] vdd gnd cell_6t
Xbit_r141_c46 bl[46] br[46] wl[141] vdd gnd cell_6t
Xbit_r142_c46 bl[46] br[46] wl[142] vdd gnd cell_6t
Xbit_r143_c46 bl[46] br[46] wl[143] vdd gnd cell_6t
Xbit_r144_c46 bl[46] br[46] wl[144] vdd gnd cell_6t
Xbit_r145_c46 bl[46] br[46] wl[145] vdd gnd cell_6t
Xbit_r146_c46 bl[46] br[46] wl[146] vdd gnd cell_6t
Xbit_r147_c46 bl[46] br[46] wl[147] vdd gnd cell_6t
Xbit_r148_c46 bl[46] br[46] wl[148] vdd gnd cell_6t
Xbit_r149_c46 bl[46] br[46] wl[149] vdd gnd cell_6t
Xbit_r150_c46 bl[46] br[46] wl[150] vdd gnd cell_6t
Xbit_r151_c46 bl[46] br[46] wl[151] vdd gnd cell_6t
Xbit_r152_c46 bl[46] br[46] wl[152] vdd gnd cell_6t
Xbit_r153_c46 bl[46] br[46] wl[153] vdd gnd cell_6t
Xbit_r154_c46 bl[46] br[46] wl[154] vdd gnd cell_6t
Xbit_r155_c46 bl[46] br[46] wl[155] vdd gnd cell_6t
Xbit_r156_c46 bl[46] br[46] wl[156] vdd gnd cell_6t
Xbit_r157_c46 bl[46] br[46] wl[157] vdd gnd cell_6t
Xbit_r158_c46 bl[46] br[46] wl[158] vdd gnd cell_6t
Xbit_r159_c46 bl[46] br[46] wl[159] vdd gnd cell_6t
Xbit_r160_c46 bl[46] br[46] wl[160] vdd gnd cell_6t
Xbit_r161_c46 bl[46] br[46] wl[161] vdd gnd cell_6t
Xbit_r162_c46 bl[46] br[46] wl[162] vdd gnd cell_6t
Xbit_r163_c46 bl[46] br[46] wl[163] vdd gnd cell_6t
Xbit_r164_c46 bl[46] br[46] wl[164] vdd gnd cell_6t
Xbit_r165_c46 bl[46] br[46] wl[165] vdd gnd cell_6t
Xbit_r166_c46 bl[46] br[46] wl[166] vdd gnd cell_6t
Xbit_r167_c46 bl[46] br[46] wl[167] vdd gnd cell_6t
Xbit_r168_c46 bl[46] br[46] wl[168] vdd gnd cell_6t
Xbit_r169_c46 bl[46] br[46] wl[169] vdd gnd cell_6t
Xbit_r170_c46 bl[46] br[46] wl[170] vdd gnd cell_6t
Xbit_r171_c46 bl[46] br[46] wl[171] vdd gnd cell_6t
Xbit_r172_c46 bl[46] br[46] wl[172] vdd gnd cell_6t
Xbit_r173_c46 bl[46] br[46] wl[173] vdd gnd cell_6t
Xbit_r174_c46 bl[46] br[46] wl[174] vdd gnd cell_6t
Xbit_r175_c46 bl[46] br[46] wl[175] vdd gnd cell_6t
Xbit_r176_c46 bl[46] br[46] wl[176] vdd gnd cell_6t
Xbit_r177_c46 bl[46] br[46] wl[177] vdd gnd cell_6t
Xbit_r178_c46 bl[46] br[46] wl[178] vdd gnd cell_6t
Xbit_r179_c46 bl[46] br[46] wl[179] vdd gnd cell_6t
Xbit_r180_c46 bl[46] br[46] wl[180] vdd gnd cell_6t
Xbit_r181_c46 bl[46] br[46] wl[181] vdd gnd cell_6t
Xbit_r182_c46 bl[46] br[46] wl[182] vdd gnd cell_6t
Xbit_r183_c46 bl[46] br[46] wl[183] vdd gnd cell_6t
Xbit_r184_c46 bl[46] br[46] wl[184] vdd gnd cell_6t
Xbit_r185_c46 bl[46] br[46] wl[185] vdd gnd cell_6t
Xbit_r186_c46 bl[46] br[46] wl[186] vdd gnd cell_6t
Xbit_r187_c46 bl[46] br[46] wl[187] vdd gnd cell_6t
Xbit_r188_c46 bl[46] br[46] wl[188] vdd gnd cell_6t
Xbit_r189_c46 bl[46] br[46] wl[189] vdd gnd cell_6t
Xbit_r190_c46 bl[46] br[46] wl[190] vdd gnd cell_6t
Xbit_r191_c46 bl[46] br[46] wl[191] vdd gnd cell_6t
Xbit_r192_c46 bl[46] br[46] wl[192] vdd gnd cell_6t
Xbit_r193_c46 bl[46] br[46] wl[193] vdd gnd cell_6t
Xbit_r194_c46 bl[46] br[46] wl[194] vdd gnd cell_6t
Xbit_r195_c46 bl[46] br[46] wl[195] vdd gnd cell_6t
Xbit_r196_c46 bl[46] br[46] wl[196] vdd gnd cell_6t
Xbit_r197_c46 bl[46] br[46] wl[197] vdd gnd cell_6t
Xbit_r198_c46 bl[46] br[46] wl[198] vdd gnd cell_6t
Xbit_r199_c46 bl[46] br[46] wl[199] vdd gnd cell_6t
Xbit_r200_c46 bl[46] br[46] wl[200] vdd gnd cell_6t
Xbit_r201_c46 bl[46] br[46] wl[201] vdd gnd cell_6t
Xbit_r202_c46 bl[46] br[46] wl[202] vdd gnd cell_6t
Xbit_r203_c46 bl[46] br[46] wl[203] vdd gnd cell_6t
Xbit_r204_c46 bl[46] br[46] wl[204] vdd gnd cell_6t
Xbit_r205_c46 bl[46] br[46] wl[205] vdd gnd cell_6t
Xbit_r206_c46 bl[46] br[46] wl[206] vdd gnd cell_6t
Xbit_r207_c46 bl[46] br[46] wl[207] vdd gnd cell_6t
Xbit_r208_c46 bl[46] br[46] wl[208] vdd gnd cell_6t
Xbit_r209_c46 bl[46] br[46] wl[209] vdd gnd cell_6t
Xbit_r210_c46 bl[46] br[46] wl[210] vdd gnd cell_6t
Xbit_r211_c46 bl[46] br[46] wl[211] vdd gnd cell_6t
Xbit_r212_c46 bl[46] br[46] wl[212] vdd gnd cell_6t
Xbit_r213_c46 bl[46] br[46] wl[213] vdd gnd cell_6t
Xbit_r214_c46 bl[46] br[46] wl[214] vdd gnd cell_6t
Xbit_r215_c46 bl[46] br[46] wl[215] vdd gnd cell_6t
Xbit_r216_c46 bl[46] br[46] wl[216] vdd gnd cell_6t
Xbit_r217_c46 bl[46] br[46] wl[217] vdd gnd cell_6t
Xbit_r218_c46 bl[46] br[46] wl[218] vdd gnd cell_6t
Xbit_r219_c46 bl[46] br[46] wl[219] vdd gnd cell_6t
Xbit_r220_c46 bl[46] br[46] wl[220] vdd gnd cell_6t
Xbit_r221_c46 bl[46] br[46] wl[221] vdd gnd cell_6t
Xbit_r222_c46 bl[46] br[46] wl[222] vdd gnd cell_6t
Xbit_r223_c46 bl[46] br[46] wl[223] vdd gnd cell_6t
Xbit_r224_c46 bl[46] br[46] wl[224] vdd gnd cell_6t
Xbit_r225_c46 bl[46] br[46] wl[225] vdd gnd cell_6t
Xbit_r226_c46 bl[46] br[46] wl[226] vdd gnd cell_6t
Xbit_r227_c46 bl[46] br[46] wl[227] vdd gnd cell_6t
Xbit_r228_c46 bl[46] br[46] wl[228] vdd gnd cell_6t
Xbit_r229_c46 bl[46] br[46] wl[229] vdd gnd cell_6t
Xbit_r230_c46 bl[46] br[46] wl[230] vdd gnd cell_6t
Xbit_r231_c46 bl[46] br[46] wl[231] vdd gnd cell_6t
Xbit_r232_c46 bl[46] br[46] wl[232] vdd gnd cell_6t
Xbit_r233_c46 bl[46] br[46] wl[233] vdd gnd cell_6t
Xbit_r234_c46 bl[46] br[46] wl[234] vdd gnd cell_6t
Xbit_r235_c46 bl[46] br[46] wl[235] vdd gnd cell_6t
Xbit_r236_c46 bl[46] br[46] wl[236] vdd gnd cell_6t
Xbit_r237_c46 bl[46] br[46] wl[237] vdd gnd cell_6t
Xbit_r238_c46 bl[46] br[46] wl[238] vdd gnd cell_6t
Xbit_r239_c46 bl[46] br[46] wl[239] vdd gnd cell_6t
Xbit_r240_c46 bl[46] br[46] wl[240] vdd gnd cell_6t
Xbit_r241_c46 bl[46] br[46] wl[241] vdd gnd cell_6t
Xbit_r242_c46 bl[46] br[46] wl[242] vdd gnd cell_6t
Xbit_r243_c46 bl[46] br[46] wl[243] vdd gnd cell_6t
Xbit_r244_c46 bl[46] br[46] wl[244] vdd gnd cell_6t
Xbit_r245_c46 bl[46] br[46] wl[245] vdd gnd cell_6t
Xbit_r246_c46 bl[46] br[46] wl[246] vdd gnd cell_6t
Xbit_r247_c46 bl[46] br[46] wl[247] vdd gnd cell_6t
Xbit_r248_c46 bl[46] br[46] wl[248] vdd gnd cell_6t
Xbit_r249_c46 bl[46] br[46] wl[249] vdd gnd cell_6t
Xbit_r250_c46 bl[46] br[46] wl[250] vdd gnd cell_6t
Xbit_r251_c46 bl[46] br[46] wl[251] vdd gnd cell_6t
Xbit_r252_c46 bl[46] br[46] wl[252] vdd gnd cell_6t
Xbit_r253_c46 bl[46] br[46] wl[253] vdd gnd cell_6t
Xbit_r254_c46 bl[46] br[46] wl[254] vdd gnd cell_6t
Xbit_r255_c46 bl[46] br[46] wl[255] vdd gnd cell_6t
Xbit_r0_c47 bl[47] br[47] wl[0] vdd gnd cell_6t
Xbit_r1_c47 bl[47] br[47] wl[1] vdd gnd cell_6t
Xbit_r2_c47 bl[47] br[47] wl[2] vdd gnd cell_6t
Xbit_r3_c47 bl[47] br[47] wl[3] vdd gnd cell_6t
Xbit_r4_c47 bl[47] br[47] wl[4] vdd gnd cell_6t
Xbit_r5_c47 bl[47] br[47] wl[5] vdd gnd cell_6t
Xbit_r6_c47 bl[47] br[47] wl[6] vdd gnd cell_6t
Xbit_r7_c47 bl[47] br[47] wl[7] vdd gnd cell_6t
Xbit_r8_c47 bl[47] br[47] wl[8] vdd gnd cell_6t
Xbit_r9_c47 bl[47] br[47] wl[9] vdd gnd cell_6t
Xbit_r10_c47 bl[47] br[47] wl[10] vdd gnd cell_6t
Xbit_r11_c47 bl[47] br[47] wl[11] vdd gnd cell_6t
Xbit_r12_c47 bl[47] br[47] wl[12] vdd gnd cell_6t
Xbit_r13_c47 bl[47] br[47] wl[13] vdd gnd cell_6t
Xbit_r14_c47 bl[47] br[47] wl[14] vdd gnd cell_6t
Xbit_r15_c47 bl[47] br[47] wl[15] vdd gnd cell_6t
Xbit_r16_c47 bl[47] br[47] wl[16] vdd gnd cell_6t
Xbit_r17_c47 bl[47] br[47] wl[17] vdd gnd cell_6t
Xbit_r18_c47 bl[47] br[47] wl[18] vdd gnd cell_6t
Xbit_r19_c47 bl[47] br[47] wl[19] vdd gnd cell_6t
Xbit_r20_c47 bl[47] br[47] wl[20] vdd gnd cell_6t
Xbit_r21_c47 bl[47] br[47] wl[21] vdd gnd cell_6t
Xbit_r22_c47 bl[47] br[47] wl[22] vdd gnd cell_6t
Xbit_r23_c47 bl[47] br[47] wl[23] vdd gnd cell_6t
Xbit_r24_c47 bl[47] br[47] wl[24] vdd gnd cell_6t
Xbit_r25_c47 bl[47] br[47] wl[25] vdd gnd cell_6t
Xbit_r26_c47 bl[47] br[47] wl[26] vdd gnd cell_6t
Xbit_r27_c47 bl[47] br[47] wl[27] vdd gnd cell_6t
Xbit_r28_c47 bl[47] br[47] wl[28] vdd gnd cell_6t
Xbit_r29_c47 bl[47] br[47] wl[29] vdd gnd cell_6t
Xbit_r30_c47 bl[47] br[47] wl[30] vdd gnd cell_6t
Xbit_r31_c47 bl[47] br[47] wl[31] vdd gnd cell_6t
Xbit_r32_c47 bl[47] br[47] wl[32] vdd gnd cell_6t
Xbit_r33_c47 bl[47] br[47] wl[33] vdd gnd cell_6t
Xbit_r34_c47 bl[47] br[47] wl[34] vdd gnd cell_6t
Xbit_r35_c47 bl[47] br[47] wl[35] vdd gnd cell_6t
Xbit_r36_c47 bl[47] br[47] wl[36] vdd gnd cell_6t
Xbit_r37_c47 bl[47] br[47] wl[37] vdd gnd cell_6t
Xbit_r38_c47 bl[47] br[47] wl[38] vdd gnd cell_6t
Xbit_r39_c47 bl[47] br[47] wl[39] vdd gnd cell_6t
Xbit_r40_c47 bl[47] br[47] wl[40] vdd gnd cell_6t
Xbit_r41_c47 bl[47] br[47] wl[41] vdd gnd cell_6t
Xbit_r42_c47 bl[47] br[47] wl[42] vdd gnd cell_6t
Xbit_r43_c47 bl[47] br[47] wl[43] vdd gnd cell_6t
Xbit_r44_c47 bl[47] br[47] wl[44] vdd gnd cell_6t
Xbit_r45_c47 bl[47] br[47] wl[45] vdd gnd cell_6t
Xbit_r46_c47 bl[47] br[47] wl[46] vdd gnd cell_6t
Xbit_r47_c47 bl[47] br[47] wl[47] vdd gnd cell_6t
Xbit_r48_c47 bl[47] br[47] wl[48] vdd gnd cell_6t
Xbit_r49_c47 bl[47] br[47] wl[49] vdd gnd cell_6t
Xbit_r50_c47 bl[47] br[47] wl[50] vdd gnd cell_6t
Xbit_r51_c47 bl[47] br[47] wl[51] vdd gnd cell_6t
Xbit_r52_c47 bl[47] br[47] wl[52] vdd gnd cell_6t
Xbit_r53_c47 bl[47] br[47] wl[53] vdd gnd cell_6t
Xbit_r54_c47 bl[47] br[47] wl[54] vdd gnd cell_6t
Xbit_r55_c47 bl[47] br[47] wl[55] vdd gnd cell_6t
Xbit_r56_c47 bl[47] br[47] wl[56] vdd gnd cell_6t
Xbit_r57_c47 bl[47] br[47] wl[57] vdd gnd cell_6t
Xbit_r58_c47 bl[47] br[47] wl[58] vdd gnd cell_6t
Xbit_r59_c47 bl[47] br[47] wl[59] vdd gnd cell_6t
Xbit_r60_c47 bl[47] br[47] wl[60] vdd gnd cell_6t
Xbit_r61_c47 bl[47] br[47] wl[61] vdd gnd cell_6t
Xbit_r62_c47 bl[47] br[47] wl[62] vdd gnd cell_6t
Xbit_r63_c47 bl[47] br[47] wl[63] vdd gnd cell_6t
Xbit_r64_c47 bl[47] br[47] wl[64] vdd gnd cell_6t
Xbit_r65_c47 bl[47] br[47] wl[65] vdd gnd cell_6t
Xbit_r66_c47 bl[47] br[47] wl[66] vdd gnd cell_6t
Xbit_r67_c47 bl[47] br[47] wl[67] vdd gnd cell_6t
Xbit_r68_c47 bl[47] br[47] wl[68] vdd gnd cell_6t
Xbit_r69_c47 bl[47] br[47] wl[69] vdd gnd cell_6t
Xbit_r70_c47 bl[47] br[47] wl[70] vdd gnd cell_6t
Xbit_r71_c47 bl[47] br[47] wl[71] vdd gnd cell_6t
Xbit_r72_c47 bl[47] br[47] wl[72] vdd gnd cell_6t
Xbit_r73_c47 bl[47] br[47] wl[73] vdd gnd cell_6t
Xbit_r74_c47 bl[47] br[47] wl[74] vdd gnd cell_6t
Xbit_r75_c47 bl[47] br[47] wl[75] vdd gnd cell_6t
Xbit_r76_c47 bl[47] br[47] wl[76] vdd gnd cell_6t
Xbit_r77_c47 bl[47] br[47] wl[77] vdd gnd cell_6t
Xbit_r78_c47 bl[47] br[47] wl[78] vdd gnd cell_6t
Xbit_r79_c47 bl[47] br[47] wl[79] vdd gnd cell_6t
Xbit_r80_c47 bl[47] br[47] wl[80] vdd gnd cell_6t
Xbit_r81_c47 bl[47] br[47] wl[81] vdd gnd cell_6t
Xbit_r82_c47 bl[47] br[47] wl[82] vdd gnd cell_6t
Xbit_r83_c47 bl[47] br[47] wl[83] vdd gnd cell_6t
Xbit_r84_c47 bl[47] br[47] wl[84] vdd gnd cell_6t
Xbit_r85_c47 bl[47] br[47] wl[85] vdd gnd cell_6t
Xbit_r86_c47 bl[47] br[47] wl[86] vdd gnd cell_6t
Xbit_r87_c47 bl[47] br[47] wl[87] vdd gnd cell_6t
Xbit_r88_c47 bl[47] br[47] wl[88] vdd gnd cell_6t
Xbit_r89_c47 bl[47] br[47] wl[89] vdd gnd cell_6t
Xbit_r90_c47 bl[47] br[47] wl[90] vdd gnd cell_6t
Xbit_r91_c47 bl[47] br[47] wl[91] vdd gnd cell_6t
Xbit_r92_c47 bl[47] br[47] wl[92] vdd gnd cell_6t
Xbit_r93_c47 bl[47] br[47] wl[93] vdd gnd cell_6t
Xbit_r94_c47 bl[47] br[47] wl[94] vdd gnd cell_6t
Xbit_r95_c47 bl[47] br[47] wl[95] vdd gnd cell_6t
Xbit_r96_c47 bl[47] br[47] wl[96] vdd gnd cell_6t
Xbit_r97_c47 bl[47] br[47] wl[97] vdd gnd cell_6t
Xbit_r98_c47 bl[47] br[47] wl[98] vdd gnd cell_6t
Xbit_r99_c47 bl[47] br[47] wl[99] vdd gnd cell_6t
Xbit_r100_c47 bl[47] br[47] wl[100] vdd gnd cell_6t
Xbit_r101_c47 bl[47] br[47] wl[101] vdd gnd cell_6t
Xbit_r102_c47 bl[47] br[47] wl[102] vdd gnd cell_6t
Xbit_r103_c47 bl[47] br[47] wl[103] vdd gnd cell_6t
Xbit_r104_c47 bl[47] br[47] wl[104] vdd gnd cell_6t
Xbit_r105_c47 bl[47] br[47] wl[105] vdd gnd cell_6t
Xbit_r106_c47 bl[47] br[47] wl[106] vdd gnd cell_6t
Xbit_r107_c47 bl[47] br[47] wl[107] vdd gnd cell_6t
Xbit_r108_c47 bl[47] br[47] wl[108] vdd gnd cell_6t
Xbit_r109_c47 bl[47] br[47] wl[109] vdd gnd cell_6t
Xbit_r110_c47 bl[47] br[47] wl[110] vdd gnd cell_6t
Xbit_r111_c47 bl[47] br[47] wl[111] vdd gnd cell_6t
Xbit_r112_c47 bl[47] br[47] wl[112] vdd gnd cell_6t
Xbit_r113_c47 bl[47] br[47] wl[113] vdd gnd cell_6t
Xbit_r114_c47 bl[47] br[47] wl[114] vdd gnd cell_6t
Xbit_r115_c47 bl[47] br[47] wl[115] vdd gnd cell_6t
Xbit_r116_c47 bl[47] br[47] wl[116] vdd gnd cell_6t
Xbit_r117_c47 bl[47] br[47] wl[117] vdd gnd cell_6t
Xbit_r118_c47 bl[47] br[47] wl[118] vdd gnd cell_6t
Xbit_r119_c47 bl[47] br[47] wl[119] vdd gnd cell_6t
Xbit_r120_c47 bl[47] br[47] wl[120] vdd gnd cell_6t
Xbit_r121_c47 bl[47] br[47] wl[121] vdd gnd cell_6t
Xbit_r122_c47 bl[47] br[47] wl[122] vdd gnd cell_6t
Xbit_r123_c47 bl[47] br[47] wl[123] vdd gnd cell_6t
Xbit_r124_c47 bl[47] br[47] wl[124] vdd gnd cell_6t
Xbit_r125_c47 bl[47] br[47] wl[125] vdd gnd cell_6t
Xbit_r126_c47 bl[47] br[47] wl[126] vdd gnd cell_6t
Xbit_r127_c47 bl[47] br[47] wl[127] vdd gnd cell_6t
Xbit_r128_c47 bl[47] br[47] wl[128] vdd gnd cell_6t
Xbit_r129_c47 bl[47] br[47] wl[129] vdd gnd cell_6t
Xbit_r130_c47 bl[47] br[47] wl[130] vdd gnd cell_6t
Xbit_r131_c47 bl[47] br[47] wl[131] vdd gnd cell_6t
Xbit_r132_c47 bl[47] br[47] wl[132] vdd gnd cell_6t
Xbit_r133_c47 bl[47] br[47] wl[133] vdd gnd cell_6t
Xbit_r134_c47 bl[47] br[47] wl[134] vdd gnd cell_6t
Xbit_r135_c47 bl[47] br[47] wl[135] vdd gnd cell_6t
Xbit_r136_c47 bl[47] br[47] wl[136] vdd gnd cell_6t
Xbit_r137_c47 bl[47] br[47] wl[137] vdd gnd cell_6t
Xbit_r138_c47 bl[47] br[47] wl[138] vdd gnd cell_6t
Xbit_r139_c47 bl[47] br[47] wl[139] vdd gnd cell_6t
Xbit_r140_c47 bl[47] br[47] wl[140] vdd gnd cell_6t
Xbit_r141_c47 bl[47] br[47] wl[141] vdd gnd cell_6t
Xbit_r142_c47 bl[47] br[47] wl[142] vdd gnd cell_6t
Xbit_r143_c47 bl[47] br[47] wl[143] vdd gnd cell_6t
Xbit_r144_c47 bl[47] br[47] wl[144] vdd gnd cell_6t
Xbit_r145_c47 bl[47] br[47] wl[145] vdd gnd cell_6t
Xbit_r146_c47 bl[47] br[47] wl[146] vdd gnd cell_6t
Xbit_r147_c47 bl[47] br[47] wl[147] vdd gnd cell_6t
Xbit_r148_c47 bl[47] br[47] wl[148] vdd gnd cell_6t
Xbit_r149_c47 bl[47] br[47] wl[149] vdd gnd cell_6t
Xbit_r150_c47 bl[47] br[47] wl[150] vdd gnd cell_6t
Xbit_r151_c47 bl[47] br[47] wl[151] vdd gnd cell_6t
Xbit_r152_c47 bl[47] br[47] wl[152] vdd gnd cell_6t
Xbit_r153_c47 bl[47] br[47] wl[153] vdd gnd cell_6t
Xbit_r154_c47 bl[47] br[47] wl[154] vdd gnd cell_6t
Xbit_r155_c47 bl[47] br[47] wl[155] vdd gnd cell_6t
Xbit_r156_c47 bl[47] br[47] wl[156] vdd gnd cell_6t
Xbit_r157_c47 bl[47] br[47] wl[157] vdd gnd cell_6t
Xbit_r158_c47 bl[47] br[47] wl[158] vdd gnd cell_6t
Xbit_r159_c47 bl[47] br[47] wl[159] vdd gnd cell_6t
Xbit_r160_c47 bl[47] br[47] wl[160] vdd gnd cell_6t
Xbit_r161_c47 bl[47] br[47] wl[161] vdd gnd cell_6t
Xbit_r162_c47 bl[47] br[47] wl[162] vdd gnd cell_6t
Xbit_r163_c47 bl[47] br[47] wl[163] vdd gnd cell_6t
Xbit_r164_c47 bl[47] br[47] wl[164] vdd gnd cell_6t
Xbit_r165_c47 bl[47] br[47] wl[165] vdd gnd cell_6t
Xbit_r166_c47 bl[47] br[47] wl[166] vdd gnd cell_6t
Xbit_r167_c47 bl[47] br[47] wl[167] vdd gnd cell_6t
Xbit_r168_c47 bl[47] br[47] wl[168] vdd gnd cell_6t
Xbit_r169_c47 bl[47] br[47] wl[169] vdd gnd cell_6t
Xbit_r170_c47 bl[47] br[47] wl[170] vdd gnd cell_6t
Xbit_r171_c47 bl[47] br[47] wl[171] vdd gnd cell_6t
Xbit_r172_c47 bl[47] br[47] wl[172] vdd gnd cell_6t
Xbit_r173_c47 bl[47] br[47] wl[173] vdd gnd cell_6t
Xbit_r174_c47 bl[47] br[47] wl[174] vdd gnd cell_6t
Xbit_r175_c47 bl[47] br[47] wl[175] vdd gnd cell_6t
Xbit_r176_c47 bl[47] br[47] wl[176] vdd gnd cell_6t
Xbit_r177_c47 bl[47] br[47] wl[177] vdd gnd cell_6t
Xbit_r178_c47 bl[47] br[47] wl[178] vdd gnd cell_6t
Xbit_r179_c47 bl[47] br[47] wl[179] vdd gnd cell_6t
Xbit_r180_c47 bl[47] br[47] wl[180] vdd gnd cell_6t
Xbit_r181_c47 bl[47] br[47] wl[181] vdd gnd cell_6t
Xbit_r182_c47 bl[47] br[47] wl[182] vdd gnd cell_6t
Xbit_r183_c47 bl[47] br[47] wl[183] vdd gnd cell_6t
Xbit_r184_c47 bl[47] br[47] wl[184] vdd gnd cell_6t
Xbit_r185_c47 bl[47] br[47] wl[185] vdd gnd cell_6t
Xbit_r186_c47 bl[47] br[47] wl[186] vdd gnd cell_6t
Xbit_r187_c47 bl[47] br[47] wl[187] vdd gnd cell_6t
Xbit_r188_c47 bl[47] br[47] wl[188] vdd gnd cell_6t
Xbit_r189_c47 bl[47] br[47] wl[189] vdd gnd cell_6t
Xbit_r190_c47 bl[47] br[47] wl[190] vdd gnd cell_6t
Xbit_r191_c47 bl[47] br[47] wl[191] vdd gnd cell_6t
Xbit_r192_c47 bl[47] br[47] wl[192] vdd gnd cell_6t
Xbit_r193_c47 bl[47] br[47] wl[193] vdd gnd cell_6t
Xbit_r194_c47 bl[47] br[47] wl[194] vdd gnd cell_6t
Xbit_r195_c47 bl[47] br[47] wl[195] vdd gnd cell_6t
Xbit_r196_c47 bl[47] br[47] wl[196] vdd gnd cell_6t
Xbit_r197_c47 bl[47] br[47] wl[197] vdd gnd cell_6t
Xbit_r198_c47 bl[47] br[47] wl[198] vdd gnd cell_6t
Xbit_r199_c47 bl[47] br[47] wl[199] vdd gnd cell_6t
Xbit_r200_c47 bl[47] br[47] wl[200] vdd gnd cell_6t
Xbit_r201_c47 bl[47] br[47] wl[201] vdd gnd cell_6t
Xbit_r202_c47 bl[47] br[47] wl[202] vdd gnd cell_6t
Xbit_r203_c47 bl[47] br[47] wl[203] vdd gnd cell_6t
Xbit_r204_c47 bl[47] br[47] wl[204] vdd gnd cell_6t
Xbit_r205_c47 bl[47] br[47] wl[205] vdd gnd cell_6t
Xbit_r206_c47 bl[47] br[47] wl[206] vdd gnd cell_6t
Xbit_r207_c47 bl[47] br[47] wl[207] vdd gnd cell_6t
Xbit_r208_c47 bl[47] br[47] wl[208] vdd gnd cell_6t
Xbit_r209_c47 bl[47] br[47] wl[209] vdd gnd cell_6t
Xbit_r210_c47 bl[47] br[47] wl[210] vdd gnd cell_6t
Xbit_r211_c47 bl[47] br[47] wl[211] vdd gnd cell_6t
Xbit_r212_c47 bl[47] br[47] wl[212] vdd gnd cell_6t
Xbit_r213_c47 bl[47] br[47] wl[213] vdd gnd cell_6t
Xbit_r214_c47 bl[47] br[47] wl[214] vdd gnd cell_6t
Xbit_r215_c47 bl[47] br[47] wl[215] vdd gnd cell_6t
Xbit_r216_c47 bl[47] br[47] wl[216] vdd gnd cell_6t
Xbit_r217_c47 bl[47] br[47] wl[217] vdd gnd cell_6t
Xbit_r218_c47 bl[47] br[47] wl[218] vdd gnd cell_6t
Xbit_r219_c47 bl[47] br[47] wl[219] vdd gnd cell_6t
Xbit_r220_c47 bl[47] br[47] wl[220] vdd gnd cell_6t
Xbit_r221_c47 bl[47] br[47] wl[221] vdd gnd cell_6t
Xbit_r222_c47 bl[47] br[47] wl[222] vdd gnd cell_6t
Xbit_r223_c47 bl[47] br[47] wl[223] vdd gnd cell_6t
Xbit_r224_c47 bl[47] br[47] wl[224] vdd gnd cell_6t
Xbit_r225_c47 bl[47] br[47] wl[225] vdd gnd cell_6t
Xbit_r226_c47 bl[47] br[47] wl[226] vdd gnd cell_6t
Xbit_r227_c47 bl[47] br[47] wl[227] vdd gnd cell_6t
Xbit_r228_c47 bl[47] br[47] wl[228] vdd gnd cell_6t
Xbit_r229_c47 bl[47] br[47] wl[229] vdd gnd cell_6t
Xbit_r230_c47 bl[47] br[47] wl[230] vdd gnd cell_6t
Xbit_r231_c47 bl[47] br[47] wl[231] vdd gnd cell_6t
Xbit_r232_c47 bl[47] br[47] wl[232] vdd gnd cell_6t
Xbit_r233_c47 bl[47] br[47] wl[233] vdd gnd cell_6t
Xbit_r234_c47 bl[47] br[47] wl[234] vdd gnd cell_6t
Xbit_r235_c47 bl[47] br[47] wl[235] vdd gnd cell_6t
Xbit_r236_c47 bl[47] br[47] wl[236] vdd gnd cell_6t
Xbit_r237_c47 bl[47] br[47] wl[237] vdd gnd cell_6t
Xbit_r238_c47 bl[47] br[47] wl[238] vdd gnd cell_6t
Xbit_r239_c47 bl[47] br[47] wl[239] vdd gnd cell_6t
Xbit_r240_c47 bl[47] br[47] wl[240] vdd gnd cell_6t
Xbit_r241_c47 bl[47] br[47] wl[241] vdd gnd cell_6t
Xbit_r242_c47 bl[47] br[47] wl[242] vdd gnd cell_6t
Xbit_r243_c47 bl[47] br[47] wl[243] vdd gnd cell_6t
Xbit_r244_c47 bl[47] br[47] wl[244] vdd gnd cell_6t
Xbit_r245_c47 bl[47] br[47] wl[245] vdd gnd cell_6t
Xbit_r246_c47 bl[47] br[47] wl[246] vdd gnd cell_6t
Xbit_r247_c47 bl[47] br[47] wl[247] vdd gnd cell_6t
Xbit_r248_c47 bl[47] br[47] wl[248] vdd gnd cell_6t
Xbit_r249_c47 bl[47] br[47] wl[249] vdd gnd cell_6t
Xbit_r250_c47 bl[47] br[47] wl[250] vdd gnd cell_6t
Xbit_r251_c47 bl[47] br[47] wl[251] vdd gnd cell_6t
Xbit_r252_c47 bl[47] br[47] wl[252] vdd gnd cell_6t
Xbit_r253_c47 bl[47] br[47] wl[253] vdd gnd cell_6t
Xbit_r254_c47 bl[47] br[47] wl[254] vdd gnd cell_6t
Xbit_r255_c47 bl[47] br[47] wl[255] vdd gnd cell_6t
Xbit_r0_c48 bl[48] br[48] wl[0] vdd gnd cell_6t
Xbit_r1_c48 bl[48] br[48] wl[1] vdd gnd cell_6t
Xbit_r2_c48 bl[48] br[48] wl[2] vdd gnd cell_6t
Xbit_r3_c48 bl[48] br[48] wl[3] vdd gnd cell_6t
Xbit_r4_c48 bl[48] br[48] wl[4] vdd gnd cell_6t
Xbit_r5_c48 bl[48] br[48] wl[5] vdd gnd cell_6t
Xbit_r6_c48 bl[48] br[48] wl[6] vdd gnd cell_6t
Xbit_r7_c48 bl[48] br[48] wl[7] vdd gnd cell_6t
Xbit_r8_c48 bl[48] br[48] wl[8] vdd gnd cell_6t
Xbit_r9_c48 bl[48] br[48] wl[9] vdd gnd cell_6t
Xbit_r10_c48 bl[48] br[48] wl[10] vdd gnd cell_6t
Xbit_r11_c48 bl[48] br[48] wl[11] vdd gnd cell_6t
Xbit_r12_c48 bl[48] br[48] wl[12] vdd gnd cell_6t
Xbit_r13_c48 bl[48] br[48] wl[13] vdd gnd cell_6t
Xbit_r14_c48 bl[48] br[48] wl[14] vdd gnd cell_6t
Xbit_r15_c48 bl[48] br[48] wl[15] vdd gnd cell_6t
Xbit_r16_c48 bl[48] br[48] wl[16] vdd gnd cell_6t
Xbit_r17_c48 bl[48] br[48] wl[17] vdd gnd cell_6t
Xbit_r18_c48 bl[48] br[48] wl[18] vdd gnd cell_6t
Xbit_r19_c48 bl[48] br[48] wl[19] vdd gnd cell_6t
Xbit_r20_c48 bl[48] br[48] wl[20] vdd gnd cell_6t
Xbit_r21_c48 bl[48] br[48] wl[21] vdd gnd cell_6t
Xbit_r22_c48 bl[48] br[48] wl[22] vdd gnd cell_6t
Xbit_r23_c48 bl[48] br[48] wl[23] vdd gnd cell_6t
Xbit_r24_c48 bl[48] br[48] wl[24] vdd gnd cell_6t
Xbit_r25_c48 bl[48] br[48] wl[25] vdd gnd cell_6t
Xbit_r26_c48 bl[48] br[48] wl[26] vdd gnd cell_6t
Xbit_r27_c48 bl[48] br[48] wl[27] vdd gnd cell_6t
Xbit_r28_c48 bl[48] br[48] wl[28] vdd gnd cell_6t
Xbit_r29_c48 bl[48] br[48] wl[29] vdd gnd cell_6t
Xbit_r30_c48 bl[48] br[48] wl[30] vdd gnd cell_6t
Xbit_r31_c48 bl[48] br[48] wl[31] vdd gnd cell_6t
Xbit_r32_c48 bl[48] br[48] wl[32] vdd gnd cell_6t
Xbit_r33_c48 bl[48] br[48] wl[33] vdd gnd cell_6t
Xbit_r34_c48 bl[48] br[48] wl[34] vdd gnd cell_6t
Xbit_r35_c48 bl[48] br[48] wl[35] vdd gnd cell_6t
Xbit_r36_c48 bl[48] br[48] wl[36] vdd gnd cell_6t
Xbit_r37_c48 bl[48] br[48] wl[37] vdd gnd cell_6t
Xbit_r38_c48 bl[48] br[48] wl[38] vdd gnd cell_6t
Xbit_r39_c48 bl[48] br[48] wl[39] vdd gnd cell_6t
Xbit_r40_c48 bl[48] br[48] wl[40] vdd gnd cell_6t
Xbit_r41_c48 bl[48] br[48] wl[41] vdd gnd cell_6t
Xbit_r42_c48 bl[48] br[48] wl[42] vdd gnd cell_6t
Xbit_r43_c48 bl[48] br[48] wl[43] vdd gnd cell_6t
Xbit_r44_c48 bl[48] br[48] wl[44] vdd gnd cell_6t
Xbit_r45_c48 bl[48] br[48] wl[45] vdd gnd cell_6t
Xbit_r46_c48 bl[48] br[48] wl[46] vdd gnd cell_6t
Xbit_r47_c48 bl[48] br[48] wl[47] vdd gnd cell_6t
Xbit_r48_c48 bl[48] br[48] wl[48] vdd gnd cell_6t
Xbit_r49_c48 bl[48] br[48] wl[49] vdd gnd cell_6t
Xbit_r50_c48 bl[48] br[48] wl[50] vdd gnd cell_6t
Xbit_r51_c48 bl[48] br[48] wl[51] vdd gnd cell_6t
Xbit_r52_c48 bl[48] br[48] wl[52] vdd gnd cell_6t
Xbit_r53_c48 bl[48] br[48] wl[53] vdd gnd cell_6t
Xbit_r54_c48 bl[48] br[48] wl[54] vdd gnd cell_6t
Xbit_r55_c48 bl[48] br[48] wl[55] vdd gnd cell_6t
Xbit_r56_c48 bl[48] br[48] wl[56] vdd gnd cell_6t
Xbit_r57_c48 bl[48] br[48] wl[57] vdd gnd cell_6t
Xbit_r58_c48 bl[48] br[48] wl[58] vdd gnd cell_6t
Xbit_r59_c48 bl[48] br[48] wl[59] vdd gnd cell_6t
Xbit_r60_c48 bl[48] br[48] wl[60] vdd gnd cell_6t
Xbit_r61_c48 bl[48] br[48] wl[61] vdd gnd cell_6t
Xbit_r62_c48 bl[48] br[48] wl[62] vdd gnd cell_6t
Xbit_r63_c48 bl[48] br[48] wl[63] vdd gnd cell_6t
Xbit_r64_c48 bl[48] br[48] wl[64] vdd gnd cell_6t
Xbit_r65_c48 bl[48] br[48] wl[65] vdd gnd cell_6t
Xbit_r66_c48 bl[48] br[48] wl[66] vdd gnd cell_6t
Xbit_r67_c48 bl[48] br[48] wl[67] vdd gnd cell_6t
Xbit_r68_c48 bl[48] br[48] wl[68] vdd gnd cell_6t
Xbit_r69_c48 bl[48] br[48] wl[69] vdd gnd cell_6t
Xbit_r70_c48 bl[48] br[48] wl[70] vdd gnd cell_6t
Xbit_r71_c48 bl[48] br[48] wl[71] vdd gnd cell_6t
Xbit_r72_c48 bl[48] br[48] wl[72] vdd gnd cell_6t
Xbit_r73_c48 bl[48] br[48] wl[73] vdd gnd cell_6t
Xbit_r74_c48 bl[48] br[48] wl[74] vdd gnd cell_6t
Xbit_r75_c48 bl[48] br[48] wl[75] vdd gnd cell_6t
Xbit_r76_c48 bl[48] br[48] wl[76] vdd gnd cell_6t
Xbit_r77_c48 bl[48] br[48] wl[77] vdd gnd cell_6t
Xbit_r78_c48 bl[48] br[48] wl[78] vdd gnd cell_6t
Xbit_r79_c48 bl[48] br[48] wl[79] vdd gnd cell_6t
Xbit_r80_c48 bl[48] br[48] wl[80] vdd gnd cell_6t
Xbit_r81_c48 bl[48] br[48] wl[81] vdd gnd cell_6t
Xbit_r82_c48 bl[48] br[48] wl[82] vdd gnd cell_6t
Xbit_r83_c48 bl[48] br[48] wl[83] vdd gnd cell_6t
Xbit_r84_c48 bl[48] br[48] wl[84] vdd gnd cell_6t
Xbit_r85_c48 bl[48] br[48] wl[85] vdd gnd cell_6t
Xbit_r86_c48 bl[48] br[48] wl[86] vdd gnd cell_6t
Xbit_r87_c48 bl[48] br[48] wl[87] vdd gnd cell_6t
Xbit_r88_c48 bl[48] br[48] wl[88] vdd gnd cell_6t
Xbit_r89_c48 bl[48] br[48] wl[89] vdd gnd cell_6t
Xbit_r90_c48 bl[48] br[48] wl[90] vdd gnd cell_6t
Xbit_r91_c48 bl[48] br[48] wl[91] vdd gnd cell_6t
Xbit_r92_c48 bl[48] br[48] wl[92] vdd gnd cell_6t
Xbit_r93_c48 bl[48] br[48] wl[93] vdd gnd cell_6t
Xbit_r94_c48 bl[48] br[48] wl[94] vdd gnd cell_6t
Xbit_r95_c48 bl[48] br[48] wl[95] vdd gnd cell_6t
Xbit_r96_c48 bl[48] br[48] wl[96] vdd gnd cell_6t
Xbit_r97_c48 bl[48] br[48] wl[97] vdd gnd cell_6t
Xbit_r98_c48 bl[48] br[48] wl[98] vdd gnd cell_6t
Xbit_r99_c48 bl[48] br[48] wl[99] vdd gnd cell_6t
Xbit_r100_c48 bl[48] br[48] wl[100] vdd gnd cell_6t
Xbit_r101_c48 bl[48] br[48] wl[101] vdd gnd cell_6t
Xbit_r102_c48 bl[48] br[48] wl[102] vdd gnd cell_6t
Xbit_r103_c48 bl[48] br[48] wl[103] vdd gnd cell_6t
Xbit_r104_c48 bl[48] br[48] wl[104] vdd gnd cell_6t
Xbit_r105_c48 bl[48] br[48] wl[105] vdd gnd cell_6t
Xbit_r106_c48 bl[48] br[48] wl[106] vdd gnd cell_6t
Xbit_r107_c48 bl[48] br[48] wl[107] vdd gnd cell_6t
Xbit_r108_c48 bl[48] br[48] wl[108] vdd gnd cell_6t
Xbit_r109_c48 bl[48] br[48] wl[109] vdd gnd cell_6t
Xbit_r110_c48 bl[48] br[48] wl[110] vdd gnd cell_6t
Xbit_r111_c48 bl[48] br[48] wl[111] vdd gnd cell_6t
Xbit_r112_c48 bl[48] br[48] wl[112] vdd gnd cell_6t
Xbit_r113_c48 bl[48] br[48] wl[113] vdd gnd cell_6t
Xbit_r114_c48 bl[48] br[48] wl[114] vdd gnd cell_6t
Xbit_r115_c48 bl[48] br[48] wl[115] vdd gnd cell_6t
Xbit_r116_c48 bl[48] br[48] wl[116] vdd gnd cell_6t
Xbit_r117_c48 bl[48] br[48] wl[117] vdd gnd cell_6t
Xbit_r118_c48 bl[48] br[48] wl[118] vdd gnd cell_6t
Xbit_r119_c48 bl[48] br[48] wl[119] vdd gnd cell_6t
Xbit_r120_c48 bl[48] br[48] wl[120] vdd gnd cell_6t
Xbit_r121_c48 bl[48] br[48] wl[121] vdd gnd cell_6t
Xbit_r122_c48 bl[48] br[48] wl[122] vdd gnd cell_6t
Xbit_r123_c48 bl[48] br[48] wl[123] vdd gnd cell_6t
Xbit_r124_c48 bl[48] br[48] wl[124] vdd gnd cell_6t
Xbit_r125_c48 bl[48] br[48] wl[125] vdd gnd cell_6t
Xbit_r126_c48 bl[48] br[48] wl[126] vdd gnd cell_6t
Xbit_r127_c48 bl[48] br[48] wl[127] vdd gnd cell_6t
Xbit_r128_c48 bl[48] br[48] wl[128] vdd gnd cell_6t
Xbit_r129_c48 bl[48] br[48] wl[129] vdd gnd cell_6t
Xbit_r130_c48 bl[48] br[48] wl[130] vdd gnd cell_6t
Xbit_r131_c48 bl[48] br[48] wl[131] vdd gnd cell_6t
Xbit_r132_c48 bl[48] br[48] wl[132] vdd gnd cell_6t
Xbit_r133_c48 bl[48] br[48] wl[133] vdd gnd cell_6t
Xbit_r134_c48 bl[48] br[48] wl[134] vdd gnd cell_6t
Xbit_r135_c48 bl[48] br[48] wl[135] vdd gnd cell_6t
Xbit_r136_c48 bl[48] br[48] wl[136] vdd gnd cell_6t
Xbit_r137_c48 bl[48] br[48] wl[137] vdd gnd cell_6t
Xbit_r138_c48 bl[48] br[48] wl[138] vdd gnd cell_6t
Xbit_r139_c48 bl[48] br[48] wl[139] vdd gnd cell_6t
Xbit_r140_c48 bl[48] br[48] wl[140] vdd gnd cell_6t
Xbit_r141_c48 bl[48] br[48] wl[141] vdd gnd cell_6t
Xbit_r142_c48 bl[48] br[48] wl[142] vdd gnd cell_6t
Xbit_r143_c48 bl[48] br[48] wl[143] vdd gnd cell_6t
Xbit_r144_c48 bl[48] br[48] wl[144] vdd gnd cell_6t
Xbit_r145_c48 bl[48] br[48] wl[145] vdd gnd cell_6t
Xbit_r146_c48 bl[48] br[48] wl[146] vdd gnd cell_6t
Xbit_r147_c48 bl[48] br[48] wl[147] vdd gnd cell_6t
Xbit_r148_c48 bl[48] br[48] wl[148] vdd gnd cell_6t
Xbit_r149_c48 bl[48] br[48] wl[149] vdd gnd cell_6t
Xbit_r150_c48 bl[48] br[48] wl[150] vdd gnd cell_6t
Xbit_r151_c48 bl[48] br[48] wl[151] vdd gnd cell_6t
Xbit_r152_c48 bl[48] br[48] wl[152] vdd gnd cell_6t
Xbit_r153_c48 bl[48] br[48] wl[153] vdd gnd cell_6t
Xbit_r154_c48 bl[48] br[48] wl[154] vdd gnd cell_6t
Xbit_r155_c48 bl[48] br[48] wl[155] vdd gnd cell_6t
Xbit_r156_c48 bl[48] br[48] wl[156] vdd gnd cell_6t
Xbit_r157_c48 bl[48] br[48] wl[157] vdd gnd cell_6t
Xbit_r158_c48 bl[48] br[48] wl[158] vdd gnd cell_6t
Xbit_r159_c48 bl[48] br[48] wl[159] vdd gnd cell_6t
Xbit_r160_c48 bl[48] br[48] wl[160] vdd gnd cell_6t
Xbit_r161_c48 bl[48] br[48] wl[161] vdd gnd cell_6t
Xbit_r162_c48 bl[48] br[48] wl[162] vdd gnd cell_6t
Xbit_r163_c48 bl[48] br[48] wl[163] vdd gnd cell_6t
Xbit_r164_c48 bl[48] br[48] wl[164] vdd gnd cell_6t
Xbit_r165_c48 bl[48] br[48] wl[165] vdd gnd cell_6t
Xbit_r166_c48 bl[48] br[48] wl[166] vdd gnd cell_6t
Xbit_r167_c48 bl[48] br[48] wl[167] vdd gnd cell_6t
Xbit_r168_c48 bl[48] br[48] wl[168] vdd gnd cell_6t
Xbit_r169_c48 bl[48] br[48] wl[169] vdd gnd cell_6t
Xbit_r170_c48 bl[48] br[48] wl[170] vdd gnd cell_6t
Xbit_r171_c48 bl[48] br[48] wl[171] vdd gnd cell_6t
Xbit_r172_c48 bl[48] br[48] wl[172] vdd gnd cell_6t
Xbit_r173_c48 bl[48] br[48] wl[173] vdd gnd cell_6t
Xbit_r174_c48 bl[48] br[48] wl[174] vdd gnd cell_6t
Xbit_r175_c48 bl[48] br[48] wl[175] vdd gnd cell_6t
Xbit_r176_c48 bl[48] br[48] wl[176] vdd gnd cell_6t
Xbit_r177_c48 bl[48] br[48] wl[177] vdd gnd cell_6t
Xbit_r178_c48 bl[48] br[48] wl[178] vdd gnd cell_6t
Xbit_r179_c48 bl[48] br[48] wl[179] vdd gnd cell_6t
Xbit_r180_c48 bl[48] br[48] wl[180] vdd gnd cell_6t
Xbit_r181_c48 bl[48] br[48] wl[181] vdd gnd cell_6t
Xbit_r182_c48 bl[48] br[48] wl[182] vdd gnd cell_6t
Xbit_r183_c48 bl[48] br[48] wl[183] vdd gnd cell_6t
Xbit_r184_c48 bl[48] br[48] wl[184] vdd gnd cell_6t
Xbit_r185_c48 bl[48] br[48] wl[185] vdd gnd cell_6t
Xbit_r186_c48 bl[48] br[48] wl[186] vdd gnd cell_6t
Xbit_r187_c48 bl[48] br[48] wl[187] vdd gnd cell_6t
Xbit_r188_c48 bl[48] br[48] wl[188] vdd gnd cell_6t
Xbit_r189_c48 bl[48] br[48] wl[189] vdd gnd cell_6t
Xbit_r190_c48 bl[48] br[48] wl[190] vdd gnd cell_6t
Xbit_r191_c48 bl[48] br[48] wl[191] vdd gnd cell_6t
Xbit_r192_c48 bl[48] br[48] wl[192] vdd gnd cell_6t
Xbit_r193_c48 bl[48] br[48] wl[193] vdd gnd cell_6t
Xbit_r194_c48 bl[48] br[48] wl[194] vdd gnd cell_6t
Xbit_r195_c48 bl[48] br[48] wl[195] vdd gnd cell_6t
Xbit_r196_c48 bl[48] br[48] wl[196] vdd gnd cell_6t
Xbit_r197_c48 bl[48] br[48] wl[197] vdd gnd cell_6t
Xbit_r198_c48 bl[48] br[48] wl[198] vdd gnd cell_6t
Xbit_r199_c48 bl[48] br[48] wl[199] vdd gnd cell_6t
Xbit_r200_c48 bl[48] br[48] wl[200] vdd gnd cell_6t
Xbit_r201_c48 bl[48] br[48] wl[201] vdd gnd cell_6t
Xbit_r202_c48 bl[48] br[48] wl[202] vdd gnd cell_6t
Xbit_r203_c48 bl[48] br[48] wl[203] vdd gnd cell_6t
Xbit_r204_c48 bl[48] br[48] wl[204] vdd gnd cell_6t
Xbit_r205_c48 bl[48] br[48] wl[205] vdd gnd cell_6t
Xbit_r206_c48 bl[48] br[48] wl[206] vdd gnd cell_6t
Xbit_r207_c48 bl[48] br[48] wl[207] vdd gnd cell_6t
Xbit_r208_c48 bl[48] br[48] wl[208] vdd gnd cell_6t
Xbit_r209_c48 bl[48] br[48] wl[209] vdd gnd cell_6t
Xbit_r210_c48 bl[48] br[48] wl[210] vdd gnd cell_6t
Xbit_r211_c48 bl[48] br[48] wl[211] vdd gnd cell_6t
Xbit_r212_c48 bl[48] br[48] wl[212] vdd gnd cell_6t
Xbit_r213_c48 bl[48] br[48] wl[213] vdd gnd cell_6t
Xbit_r214_c48 bl[48] br[48] wl[214] vdd gnd cell_6t
Xbit_r215_c48 bl[48] br[48] wl[215] vdd gnd cell_6t
Xbit_r216_c48 bl[48] br[48] wl[216] vdd gnd cell_6t
Xbit_r217_c48 bl[48] br[48] wl[217] vdd gnd cell_6t
Xbit_r218_c48 bl[48] br[48] wl[218] vdd gnd cell_6t
Xbit_r219_c48 bl[48] br[48] wl[219] vdd gnd cell_6t
Xbit_r220_c48 bl[48] br[48] wl[220] vdd gnd cell_6t
Xbit_r221_c48 bl[48] br[48] wl[221] vdd gnd cell_6t
Xbit_r222_c48 bl[48] br[48] wl[222] vdd gnd cell_6t
Xbit_r223_c48 bl[48] br[48] wl[223] vdd gnd cell_6t
Xbit_r224_c48 bl[48] br[48] wl[224] vdd gnd cell_6t
Xbit_r225_c48 bl[48] br[48] wl[225] vdd gnd cell_6t
Xbit_r226_c48 bl[48] br[48] wl[226] vdd gnd cell_6t
Xbit_r227_c48 bl[48] br[48] wl[227] vdd gnd cell_6t
Xbit_r228_c48 bl[48] br[48] wl[228] vdd gnd cell_6t
Xbit_r229_c48 bl[48] br[48] wl[229] vdd gnd cell_6t
Xbit_r230_c48 bl[48] br[48] wl[230] vdd gnd cell_6t
Xbit_r231_c48 bl[48] br[48] wl[231] vdd gnd cell_6t
Xbit_r232_c48 bl[48] br[48] wl[232] vdd gnd cell_6t
Xbit_r233_c48 bl[48] br[48] wl[233] vdd gnd cell_6t
Xbit_r234_c48 bl[48] br[48] wl[234] vdd gnd cell_6t
Xbit_r235_c48 bl[48] br[48] wl[235] vdd gnd cell_6t
Xbit_r236_c48 bl[48] br[48] wl[236] vdd gnd cell_6t
Xbit_r237_c48 bl[48] br[48] wl[237] vdd gnd cell_6t
Xbit_r238_c48 bl[48] br[48] wl[238] vdd gnd cell_6t
Xbit_r239_c48 bl[48] br[48] wl[239] vdd gnd cell_6t
Xbit_r240_c48 bl[48] br[48] wl[240] vdd gnd cell_6t
Xbit_r241_c48 bl[48] br[48] wl[241] vdd gnd cell_6t
Xbit_r242_c48 bl[48] br[48] wl[242] vdd gnd cell_6t
Xbit_r243_c48 bl[48] br[48] wl[243] vdd gnd cell_6t
Xbit_r244_c48 bl[48] br[48] wl[244] vdd gnd cell_6t
Xbit_r245_c48 bl[48] br[48] wl[245] vdd gnd cell_6t
Xbit_r246_c48 bl[48] br[48] wl[246] vdd gnd cell_6t
Xbit_r247_c48 bl[48] br[48] wl[247] vdd gnd cell_6t
Xbit_r248_c48 bl[48] br[48] wl[248] vdd gnd cell_6t
Xbit_r249_c48 bl[48] br[48] wl[249] vdd gnd cell_6t
Xbit_r250_c48 bl[48] br[48] wl[250] vdd gnd cell_6t
Xbit_r251_c48 bl[48] br[48] wl[251] vdd gnd cell_6t
Xbit_r252_c48 bl[48] br[48] wl[252] vdd gnd cell_6t
Xbit_r253_c48 bl[48] br[48] wl[253] vdd gnd cell_6t
Xbit_r254_c48 bl[48] br[48] wl[254] vdd gnd cell_6t
Xbit_r255_c48 bl[48] br[48] wl[255] vdd gnd cell_6t
Xbit_r0_c49 bl[49] br[49] wl[0] vdd gnd cell_6t
Xbit_r1_c49 bl[49] br[49] wl[1] vdd gnd cell_6t
Xbit_r2_c49 bl[49] br[49] wl[2] vdd gnd cell_6t
Xbit_r3_c49 bl[49] br[49] wl[3] vdd gnd cell_6t
Xbit_r4_c49 bl[49] br[49] wl[4] vdd gnd cell_6t
Xbit_r5_c49 bl[49] br[49] wl[5] vdd gnd cell_6t
Xbit_r6_c49 bl[49] br[49] wl[6] vdd gnd cell_6t
Xbit_r7_c49 bl[49] br[49] wl[7] vdd gnd cell_6t
Xbit_r8_c49 bl[49] br[49] wl[8] vdd gnd cell_6t
Xbit_r9_c49 bl[49] br[49] wl[9] vdd gnd cell_6t
Xbit_r10_c49 bl[49] br[49] wl[10] vdd gnd cell_6t
Xbit_r11_c49 bl[49] br[49] wl[11] vdd gnd cell_6t
Xbit_r12_c49 bl[49] br[49] wl[12] vdd gnd cell_6t
Xbit_r13_c49 bl[49] br[49] wl[13] vdd gnd cell_6t
Xbit_r14_c49 bl[49] br[49] wl[14] vdd gnd cell_6t
Xbit_r15_c49 bl[49] br[49] wl[15] vdd gnd cell_6t
Xbit_r16_c49 bl[49] br[49] wl[16] vdd gnd cell_6t
Xbit_r17_c49 bl[49] br[49] wl[17] vdd gnd cell_6t
Xbit_r18_c49 bl[49] br[49] wl[18] vdd gnd cell_6t
Xbit_r19_c49 bl[49] br[49] wl[19] vdd gnd cell_6t
Xbit_r20_c49 bl[49] br[49] wl[20] vdd gnd cell_6t
Xbit_r21_c49 bl[49] br[49] wl[21] vdd gnd cell_6t
Xbit_r22_c49 bl[49] br[49] wl[22] vdd gnd cell_6t
Xbit_r23_c49 bl[49] br[49] wl[23] vdd gnd cell_6t
Xbit_r24_c49 bl[49] br[49] wl[24] vdd gnd cell_6t
Xbit_r25_c49 bl[49] br[49] wl[25] vdd gnd cell_6t
Xbit_r26_c49 bl[49] br[49] wl[26] vdd gnd cell_6t
Xbit_r27_c49 bl[49] br[49] wl[27] vdd gnd cell_6t
Xbit_r28_c49 bl[49] br[49] wl[28] vdd gnd cell_6t
Xbit_r29_c49 bl[49] br[49] wl[29] vdd gnd cell_6t
Xbit_r30_c49 bl[49] br[49] wl[30] vdd gnd cell_6t
Xbit_r31_c49 bl[49] br[49] wl[31] vdd gnd cell_6t
Xbit_r32_c49 bl[49] br[49] wl[32] vdd gnd cell_6t
Xbit_r33_c49 bl[49] br[49] wl[33] vdd gnd cell_6t
Xbit_r34_c49 bl[49] br[49] wl[34] vdd gnd cell_6t
Xbit_r35_c49 bl[49] br[49] wl[35] vdd gnd cell_6t
Xbit_r36_c49 bl[49] br[49] wl[36] vdd gnd cell_6t
Xbit_r37_c49 bl[49] br[49] wl[37] vdd gnd cell_6t
Xbit_r38_c49 bl[49] br[49] wl[38] vdd gnd cell_6t
Xbit_r39_c49 bl[49] br[49] wl[39] vdd gnd cell_6t
Xbit_r40_c49 bl[49] br[49] wl[40] vdd gnd cell_6t
Xbit_r41_c49 bl[49] br[49] wl[41] vdd gnd cell_6t
Xbit_r42_c49 bl[49] br[49] wl[42] vdd gnd cell_6t
Xbit_r43_c49 bl[49] br[49] wl[43] vdd gnd cell_6t
Xbit_r44_c49 bl[49] br[49] wl[44] vdd gnd cell_6t
Xbit_r45_c49 bl[49] br[49] wl[45] vdd gnd cell_6t
Xbit_r46_c49 bl[49] br[49] wl[46] vdd gnd cell_6t
Xbit_r47_c49 bl[49] br[49] wl[47] vdd gnd cell_6t
Xbit_r48_c49 bl[49] br[49] wl[48] vdd gnd cell_6t
Xbit_r49_c49 bl[49] br[49] wl[49] vdd gnd cell_6t
Xbit_r50_c49 bl[49] br[49] wl[50] vdd gnd cell_6t
Xbit_r51_c49 bl[49] br[49] wl[51] vdd gnd cell_6t
Xbit_r52_c49 bl[49] br[49] wl[52] vdd gnd cell_6t
Xbit_r53_c49 bl[49] br[49] wl[53] vdd gnd cell_6t
Xbit_r54_c49 bl[49] br[49] wl[54] vdd gnd cell_6t
Xbit_r55_c49 bl[49] br[49] wl[55] vdd gnd cell_6t
Xbit_r56_c49 bl[49] br[49] wl[56] vdd gnd cell_6t
Xbit_r57_c49 bl[49] br[49] wl[57] vdd gnd cell_6t
Xbit_r58_c49 bl[49] br[49] wl[58] vdd gnd cell_6t
Xbit_r59_c49 bl[49] br[49] wl[59] vdd gnd cell_6t
Xbit_r60_c49 bl[49] br[49] wl[60] vdd gnd cell_6t
Xbit_r61_c49 bl[49] br[49] wl[61] vdd gnd cell_6t
Xbit_r62_c49 bl[49] br[49] wl[62] vdd gnd cell_6t
Xbit_r63_c49 bl[49] br[49] wl[63] vdd gnd cell_6t
Xbit_r64_c49 bl[49] br[49] wl[64] vdd gnd cell_6t
Xbit_r65_c49 bl[49] br[49] wl[65] vdd gnd cell_6t
Xbit_r66_c49 bl[49] br[49] wl[66] vdd gnd cell_6t
Xbit_r67_c49 bl[49] br[49] wl[67] vdd gnd cell_6t
Xbit_r68_c49 bl[49] br[49] wl[68] vdd gnd cell_6t
Xbit_r69_c49 bl[49] br[49] wl[69] vdd gnd cell_6t
Xbit_r70_c49 bl[49] br[49] wl[70] vdd gnd cell_6t
Xbit_r71_c49 bl[49] br[49] wl[71] vdd gnd cell_6t
Xbit_r72_c49 bl[49] br[49] wl[72] vdd gnd cell_6t
Xbit_r73_c49 bl[49] br[49] wl[73] vdd gnd cell_6t
Xbit_r74_c49 bl[49] br[49] wl[74] vdd gnd cell_6t
Xbit_r75_c49 bl[49] br[49] wl[75] vdd gnd cell_6t
Xbit_r76_c49 bl[49] br[49] wl[76] vdd gnd cell_6t
Xbit_r77_c49 bl[49] br[49] wl[77] vdd gnd cell_6t
Xbit_r78_c49 bl[49] br[49] wl[78] vdd gnd cell_6t
Xbit_r79_c49 bl[49] br[49] wl[79] vdd gnd cell_6t
Xbit_r80_c49 bl[49] br[49] wl[80] vdd gnd cell_6t
Xbit_r81_c49 bl[49] br[49] wl[81] vdd gnd cell_6t
Xbit_r82_c49 bl[49] br[49] wl[82] vdd gnd cell_6t
Xbit_r83_c49 bl[49] br[49] wl[83] vdd gnd cell_6t
Xbit_r84_c49 bl[49] br[49] wl[84] vdd gnd cell_6t
Xbit_r85_c49 bl[49] br[49] wl[85] vdd gnd cell_6t
Xbit_r86_c49 bl[49] br[49] wl[86] vdd gnd cell_6t
Xbit_r87_c49 bl[49] br[49] wl[87] vdd gnd cell_6t
Xbit_r88_c49 bl[49] br[49] wl[88] vdd gnd cell_6t
Xbit_r89_c49 bl[49] br[49] wl[89] vdd gnd cell_6t
Xbit_r90_c49 bl[49] br[49] wl[90] vdd gnd cell_6t
Xbit_r91_c49 bl[49] br[49] wl[91] vdd gnd cell_6t
Xbit_r92_c49 bl[49] br[49] wl[92] vdd gnd cell_6t
Xbit_r93_c49 bl[49] br[49] wl[93] vdd gnd cell_6t
Xbit_r94_c49 bl[49] br[49] wl[94] vdd gnd cell_6t
Xbit_r95_c49 bl[49] br[49] wl[95] vdd gnd cell_6t
Xbit_r96_c49 bl[49] br[49] wl[96] vdd gnd cell_6t
Xbit_r97_c49 bl[49] br[49] wl[97] vdd gnd cell_6t
Xbit_r98_c49 bl[49] br[49] wl[98] vdd gnd cell_6t
Xbit_r99_c49 bl[49] br[49] wl[99] vdd gnd cell_6t
Xbit_r100_c49 bl[49] br[49] wl[100] vdd gnd cell_6t
Xbit_r101_c49 bl[49] br[49] wl[101] vdd gnd cell_6t
Xbit_r102_c49 bl[49] br[49] wl[102] vdd gnd cell_6t
Xbit_r103_c49 bl[49] br[49] wl[103] vdd gnd cell_6t
Xbit_r104_c49 bl[49] br[49] wl[104] vdd gnd cell_6t
Xbit_r105_c49 bl[49] br[49] wl[105] vdd gnd cell_6t
Xbit_r106_c49 bl[49] br[49] wl[106] vdd gnd cell_6t
Xbit_r107_c49 bl[49] br[49] wl[107] vdd gnd cell_6t
Xbit_r108_c49 bl[49] br[49] wl[108] vdd gnd cell_6t
Xbit_r109_c49 bl[49] br[49] wl[109] vdd gnd cell_6t
Xbit_r110_c49 bl[49] br[49] wl[110] vdd gnd cell_6t
Xbit_r111_c49 bl[49] br[49] wl[111] vdd gnd cell_6t
Xbit_r112_c49 bl[49] br[49] wl[112] vdd gnd cell_6t
Xbit_r113_c49 bl[49] br[49] wl[113] vdd gnd cell_6t
Xbit_r114_c49 bl[49] br[49] wl[114] vdd gnd cell_6t
Xbit_r115_c49 bl[49] br[49] wl[115] vdd gnd cell_6t
Xbit_r116_c49 bl[49] br[49] wl[116] vdd gnd cell_6t
Xbit_r117_c49 bl[49] br[49] wl[117] vdd gnd cell_6t
Xbit_r118_c49 bl[49] br[49] wl[118] vdd gnd cell_6t
Xbit_r119_c49 bl[49] br[49] wl[119] vdd gnd cell_6t
Xbit_r120_c49 bl[49] br[49] wl[120] vdd gnd cell_6t
Xbit_r121_c49 bl[49] br[49] wl[121] vdd gnd cell_6t
Xbit_r122_c49 bl[49] br[49] wl[122] vdd gnd cell_6t
Xbit_r123_c49 bl[49] br[49] wl[123] vdd gnd cell_6t
Xbit_r124_c49 bl[49] br[49] wl[124] vdd gnd cell_6t
Xbit_r125_c49 bl[49] br[49] wl[125] vdd gnd cell_6t
Xbit_r126_c49 bl[49] br[49] wl[126] vdd gnd cell_6t
Xbit_r127_c49 bl[49] br[49] wl[127] vdd gnd cell_6t
Xbit_r128_c49 bl[49] br[49] wl[128] vdd gnd cell_6t
Xbit_r129_c49 bl[49] br[49] wl[129] vdd gnd cell_6t
Xbit_r130_c49 bl[49] br[49] wl[130] vdd gnd cell_6t
Xbit_r131_c49 bl[49] br[49] wl[131] vdd gnd cell_6t
Xbit_r132_c49 bl[49] br[49] wl[132] vdd gnd cell_6t
Xbit_r133_c49 bl[49] br[49] wl[133] vdd gnd cell_6t
Xbit_r134_c49 bl[49] br[49] wl[134] vdd gnd cell_6t
Xbit_r135_c49 bl[49] br[49] wl[135] vdd gnd cell_6t
Xbit_r136_c49 bl[49] br[49] wl[136] vdd gnd cell_6t
Xbit_r137_c49 bl[49] br[49] wl[137] vdd gnd cell_6t
Xbit_r138_c49 bl[49] br[49] wl[138] vdd gnd cell_6t
Xbit_r139_c49 bl[49] br[49] wl[139] vdd gnd cell_6t
Xbit_r140_c49 bl[49] br[49] wl[140] vdd gnd cell_6t
Xbit_r141_c49 bl[49] br[49] wl[141] vdd gnd cell_6t
Xbit_r142_c49 bl[49] br[49] wl[142] vdd gnd cell_6t
Xbit_r143_c49 bl[49] br[49] wl[143] vdd gnd cell_6t
Xbit_r144_c49 bl[49] br[49] wl[144] vdd gnd cell_6t
Xbit_r145_c49 bl[49] br[49] wl[145] vdd gnd cell_6t
Xbit_r146_c49 bl[49] br[49] wl[146] vdd gnd cell_6t
Xbit_r147_c49 bl[49] br[49] wl[147] vdd gnd cell_6t
Xbit_r148_c49 bl[49] br[49] wl[148] vdd gnd cell_6t
Xbit_r149_c49 bl[49] br[49] wl[149] vdd gnd cell_6t
Xbit_r150_c49 bl[49] br[49] wl[150] vdd gnd cell_6t
Xbit_r151_c49 bl[49] br[49] wl[151] vdd gnd cell_6t
Xbit_r152_c49 bl[49] br[49] wl[152] vdd gnd cell_6t
Xbit_r153_c49 bl[49] br[49] wl[153] vdd gnd cell_6t
Xbit_r154_c49 bl[49] br[49] wl[154] vdd gnd cell_6t
Xbit_r155_c49 bl[49] br[49] wl[155] vdd gnd cell_6t
Xbit_r156_c49 bl[49] br[49] wl[156] vdd gnd cell_6t
Xbit_r157_c49 bl[49] br[49] wl[157] vdd gnd cell_6t
Xbit_r158_c49 bl[49] br[49] wl[158] vdd gnd cell_6t
Xbit_r159_c49 bl[49] br[49] wl[159] vdd gnd cell_6t
Xbit_r160_c49 bl[49] br[49] wl[160] vdd gnd cell_6t
Xbit_r161_c49 bl[49] br[49] wl[161] vdd gnd cell_6t
Xbit_r162_c49 bl[49] br[49] wl[162] vdd gnd cell_6t
Xbit_r163_c49 bl[49] br[49] wl[163] vdd gnd cell_6t
Xbit_r164_c49 bl[49] br[49] wl[164] vdd gnd cell_6t
Xbit_r165_c49 bl[49] br[49] wl[165] vdd gnd cell_6t
Xbit_r166_c49 bl[49] br[49] wl[166] vdd gnd cell_6t
Xbit_r167_c49 bl[49] br[49] wl[167] vdd gnd cell_6t
Xbit_r168_c49 bl[49] br[49] wl[168] vdd gnd cell_6t
Xbit_r169_c49 bl[49] br[49] wl[169] vdd gnd cell_6t
Xbit_r170_c49 bl[49] br[49] wl[170] vdd gnd cell_6t
Xbit_r171_c49 bl[49] br[49] wl[171] vdd gnd cell_6t
Xbit_r172_c49 bl[49] br[49] wl[172] vdd gnd cell_6t
Xbit_r173_c49 bl[49] br[49] wl[173] vdd gnd cell_6t
Xbit_r174_c49 bl[49] br[49] wl[174] vdd gnd cell_6t
Xbit_r175_c49 bl[49] br[49] wl[175] vdd gnd cell_6t
Xbit_r176_c49 bl[49] br[49] wl[176] vdd gnd cell_6t
Xbit_r177_c49 bl[49] br[49] wl[177] vdd gnd cell_6t
Xbit_r178_c49 bl[49] br[49] wl[178] vdd gnd cell_6t
Xbit_r179_c49 bl[49] br[49] wl[179] vdd gnd cell_6t
Xbit_r180_c49 bl[49] br[49] wl[180] vdd gnd cell_6t
Xbit_r181_c49 bl[49] br[49] wl[181] vdd gnd cell_6t
Xbit_r182_c49 bl[49] br[49] wl[182] vdd gnd cell_6t
Xbit_r183_c49 bl[49] br[49] wl[183] vdd gnd cell_6t
Xbit_r184_c49 bl[49] br[49] wl[184] vdd gnd cell_6t
Xbit_r185_c49 bl[49] br[49] wl[185] vdd gnd cell_6t
Xbit_r186_c49 bl[49] br[49] wl[186] vdd gnd cell_6t
Xbit_r187_c49 bl[49] br[49] wl[187] vdd gnd cell_6t
Xbit_r188_c49 bl[49] br[49] wl[188] vdd gnd cell_6t
Xbit_r189_c49 bl[49] br[49] wl[189] vdd gnd cell_6t
Xbit_r190_c49 bl[49] br[49] wl[190] vdd gnd cell_6t
Xbit_r191_c49 bl[49] br[49] wl[191] vdd gnd cell_6t
Xbit_r192_c49 bl[49] br[49] wl[192] vdd gnd cell_6t
Xbit_r193_c49 bl[49] br[49] wl[193] vdd gnd cell_6t
Xbit_r194_c49 bl[49] br[49] wl[194] vdd gnd cell_6t
Xbit_r195_c49 bl[49] br[49] wl[195] vdd gnd cell_6t
Xbit_r196_c49 bl[49] br[49] wl[196] vdd gnd cell_6t
Xbit_r197_c49 bl[49] br[49] wl[197] vdd gnd cell_6t
Xbit_r198_c49 bl[49] br[49] wl[198] vdd gnd cell_6t
Xbit_r199_c49 bl[49] br[49] wl[199] vdd gnd cell_6t
Xbit_r200_c49 bl[49] br[49] wl[200] vdd gnd cell_6t
Xbit_r201_c49 bl[49] br[49] wl[201] vdd gnd cell_6t
Xbit_r202_c49 bl[49] br[49] wl[202] vdd gnd cell_6t
Xbit_r203_c49 bl[49] br[49] wl[203] vdd gnd cell_6t
Xbit_r204_c49 bl[49] br[49] wl[204] vdd gnd cell_6t
Xbit_r205_c49 bl[49] br[49] wl[205] vdd gnd cell_6t
Xbit_r206_c49 bl[49] br[49] wl[206] vdd gnd cell_6t
Xbit_r207_c49 bl[49] br[49] wl[207] vdd gnd cell_6t
Xbit_r208_c49 bl[49] br[49] wl[208] vdd gnd cell_6t
Xbit_r209_c49 bl[49] br[49] wl[209] vdd gnd cell_6t
Xbit_r210_c49 bl[49] br[49] wl[210] vdd gnd cell_6t
Xbit_r211_c49 bl[49] br[49] wl[211] vdd gnd cell_6t
Xbit_r212_c49 bl[49] br[49] wl[212] vdd gnd cell_6t
Xbit_r213_c49 bl[49] br[49] wl[213] vdd gnd cell_6t
Xbit_r214_c49 bl[49] br[49] wl[214] vdd gnd cell_6t
Xbit_r215_c49 bl[49] br[49] wl[215] vdd gnd cell_6t
Xbit_r216_c49 bl[49] br[49] wl[216] vdd gnd cell_6t
Xbit_r217_c49 bl[49] br[49] wl[217] vdd gnd cell_6t
Xbit_r218_c49 bl[49] br[49] wl[218] vdd gnd cell_6t
Xbit_r219_c49 bl[49] br[49] wl[219] vdd gnd cell_6t
Xbit_r220_c49 bl[49] br[49] wl[220] vdd gnd cell_6t
Xbit_r221_c49 bl[49] br[49] wl[221] vdd gnd cell_6t
Xbit_r222_c49 bl[49] br[49] wl[222] vdd gnd cell_6t
Xbit_r223_c49 bl[49] br[49] wl[223] vdd gnd cell_6t
Xbit_r224_c49 bl[49] br[49] wl[224] vdd gnd cell_6t
Xbit_r225_c49 bl[49] br[49] wl[225] vdd gnd cell_6t
Xbit_r226_c49 bl[49] br[49] wl[226] vdd gnd cell_6t
Xbit_r227_c49 bl[49] br[49] wl[227] vdd gnd cell_6t
Xbit_r228_c49 bl[49] br[49] wl[228] vdd gnd cell_6t
Xbit_r229_c49 bl[49] br[49] wl[229] vdd gnd cell_6t
Xbit_r230_c49 bl[49] br[49] wl[230] vdd gnd cell_6t
Xbit_r231_c49 bl[49] br[49] wl[231] vdd gnd cell_6t
Xbit_r232_c49 bl[49] br[49] wl[232] vdd gnd cell_6t
Xbit_r233_c49 bl[49] br[49] wl[233] vdd gnd cell_6t
Xbit_r234_c49 bl[49] br[49] wl[234] vdd gnd cell_6t
Xbit_r235_c49 bl[49] br[49] wl[235] vdd gnd cell_6t
Xbit_r236_c49 bl[49] br[49] wl[236] vdd gnd cell_6t
Xbit_r237_c49 bl[49] br[49] wl[237] vdd gnd cell_6t
Xbit_r238_c49 bl[49] br[49] wl[238] vdd gnd cell_6t
Xbit_r239_c49 bl[49] br[49] wl[239] vdd gnd cell_6t
Xbit_r240_c49 bl[49] br[49] wl[240] vdd gnd cell_6t
Xbit_r241_c49 bl[49] br[49] wl[241] vdd gnd cell_6t
Xbit_r242_c49 bl[49] br[49] wl[242] vdd gnd cell_6t
Xbit_r243_c49 bl[49] br[49] wl[243] vdd gnd cell_6t
Xbit_r244_c49 bl[49] br[49] wl[244] vdd gnd cell_6t
Xbit_r245_c49 bl[49] br[49] wl[245] vdd gnd cell_6t
Xbit_r246_c49 bl[49] br[49] wl[246] vdd gnd cell_6t
Xbit_r247_c49 bl[49] br[49] wl[247] vdd gnd cell_6t
Xbit_r248_c49 bl[49] br[49] wl[248] vdd gnd cell_6t
Xbit_r249_c49 bl[49] br[49] wl[249] vdd gnd cell_6t
Xbit_r250_c49 bl[49] br[49] wl[250] vdd gnd cell_6t
Xbit_r251_c49 bl[49] br[49] wl[251] vdd gnd cell_6t
Xbit_r252_c49 bl[49] br[49] wl[252] vdd gnd cell_6t
Xbit_r253_c49 bl[49] br[49] wl[253] vdd gnd cell_6t
Xbit_r254_c49 bl[49] br[49] wl[254] vdd gnd cell_6t
Xbit_r255_c49 bl[49] br[49] wl[255] vdd gnd cell_6t
Xbit_r0_c50 bl[50] br[50] wl[0] vdd gnd cell_6t
Xbit_r1_c50 bl[50] br[50] wl[1] vdd gnd cell_6t
Xbit_r2_c50 bl[50] br[50] wl[2] vdd gnd cell_6t
Xbit_r3_c50 bl[50] br[50] wl[3] vdd gnd cell_6t
Xbit_r4_c50 bl[50] br[50] wl[4] vdd gnd cell_6t
Xbit_r5_c50 bl[50] br[50] wl[5] vdd gnd cell_6t
Xbit_r6_c50 bl[50] br[50] wl[6] vdd gnd cell_6t
Xbit_r7_c50 bl[50] br[50] wl[7] vdd gnd cell_6t
Xbit_r8_c50 bl[50] br[50] wl[8] vdd gnd cell_6t
Xbit_r9_c50 bl[50] br[50] wl[9] vdd gnd cell_6t
Xbit_r10_c50 bl[50] br[50] wl[10] vdd gnd cell_6t
Xbit_r11_c50 bl[50] br[50] wl[11] vdd gnd cell_6t
Xbit_r12_c50 bl[50] br[50] wl[12] vdd gnd cell_6t
Xbit_r13_c50 bl[50] br[50] wl[13] vdd gnd cell_6t
Xbit_r14_c50 bl[50] br[50] wl[14] vdd gnd cell_6t
Xbit_r15_c50 bl[50] br[50] wl[15] vdd gnd cell_6t
Xbit_r16_c50 bl[50] br[50] wl[16] vdd gnd cell_6t
Xbit_r17_c50 bl[50] br[50] wl[17] vdd gnd cell_6t
Xbit_r18_c50 bl[50] br[50] wl[18] vdd gnd cell_6t
Xbit_r19_c50 bl[50] br[50] wl[19] vdd gnd cell_6t
Xbit_r20_c50 bl[50] br[50] wl[20] vdd gnd cell_6t
Xbit_r21_c50 bl[50] br[50] wl[21] vdd gnd cell_6t
Xbit_r22_c50 bl[50] br[50] wl[22] vdd gnd cell_6t
Xbit_r23_c50 bl[50] br[50] wl[23] vdd gnd cell_6t
Xbit_r24_c50 bl[50] br[50] wl[24] vdd gnd cell_6t
Xbit_r25_c50 bl[50] br[50] wl[25] vdd gnd cell_6t
Xbit_r26_c50 bl[50] br[50] wl[26] vdd gnd cell_6t
Xbit_r27_c50 bl[50] br[50] wl[27] vdd gnd cell_6t
Xbit_r28_c50 bl[50] br[50] wl[28] vdd gnd cell_6t
Xbit_r29_c50 bl[50] br[50] wl[29] vdd gnd cell_6t
Xbit_r30_c50 bl[50] br[50] wl[30] vdd gnd cell_6t
Xbit_r31_c50 bl[50] br[50] wl[31] vdd gnd cell_6t
Xbit_r32_c50 bl[50] br[50] wl[32] vdd gnd cell_6t
Xbit_r33_c50 bl[50] br[50] wl[33] vdd gnd cell_6t
Xbit_r34_c50 bl[50] br[50] wl[34] vdd gnd cell_6t
Xbit_r35_c50 bl[50] br[50] wl[35] vdd gnd cell_6t
Xbit_r36_c50 bl[50] br[50] wl[36] vdd gnd cell_6t
Xbit_r37_c50 bl[50] br[50] wl[37] vdd gnd cell_6t
Xbit_r38_c50 bl[50] br[50] wl[38] vdd gnd cell_6t
Xbit_r39_c50 bl[50] br[50] wl[39] vdd gnd cell_6t
Xbit_r40_c50 bl[50] br[50] wl[40] vdd gnd cell_6t
Xbit_r41_c50 bl[50] br[50] wl[41] vdd gnd cell_6t
Xbit_r42_c50 bl[50] br[50] wl[42] vdd gnd cell_6t
Xbit_r43_c50 bl[50] br[50] wl[43] vdd gnd cell_6t
Xbit_r44_c50 bl[50] br[50] wl[44] vdd gnd cell_6t
Xbit_r45_c50 bl[50] br[50] wl[45] vdd gnd cell_6t
Xbit_r46_c50 bl[50] br[50] wl[46] vdd gnd cell_6t
Xbit_r47_c50 bl[50] br[50] wl[47] vdd gnd cell_6t
Xbit_r48_c50 bl[50] br[50] wl[48] vdd gnd cell_6t
Xbit_r49_c50 bl[50] br[50] wl[49] vdd gnd cell_6t
Xbit_r50_c50 bl[50] br[50] wl[50] vdd gnd cell_6t
Xbit_r51_c50 bl[50] br[50] wl[51] vdd gnd cell_6t
Xbit_r52_c50 bl[50] br[50] wl[52] vdd gnd cell_6t
Xbit_r53_c50 bl[50] br[50] wl[53] vdd gnd cell_6t
Xbit_r54_c50 bl[50] br[50] wl[54] vdd gnd cell_6t
Xbit_r55_c50 bl[50] br[50] wl[55] vdd gnd cell_6t
Xbit_r56_c50 bl[50] br[50] wl[56] vdd gnd cell_6t
Xbit_r57_c50 bl[50] br[50] wl[57] vdd gnd cell_6t
Xbit_r58_c50 bl[50] br[50] wl[58] vdd gnd cell_6t
Xbit_r59_c50 bl[50] br[50] wl[59] vdd gnd cell_6t
Xbit_r60_c50 bl[50] br[50] wl[60] vdd gnd cell_6t
Xbit_r61_c50 bl[50] br[50] wl[61] vdd gnd cell_6t
Xbit_r62_c50 bl[50] br[50] wl[62] vdd gnd cell_6t
Xbit_r63_c50 bl[50] br[50] wl[63] vdd gnd cell_6t
Xbit_r64_c50 bl[50] br[50] wl[64] vdd gnd cell_6t
Xbit_r65_c50 bl[50] br[50] wl[65] vdd gnd cell_6t
Xbit_r66_c50 bl[50] br[50] wl[66] vdd gnd cell_6t
Xbit_r67_c50 bl[50] br[50] wl[67] vdd gnd cell_6t
Xbit_r68_c50 bl[50] br[50] wl[68] vdd gnd cell_6t
Xbit_r69_c50 bl[50] br[50] wl[69] vdd gnd cell_6t
Xbit_r70_c50 bl[50] br[50] wl[70] vdd gnd cell_6t
Xbit_r71_c50 bl[50] br[50] wl[71] vdd gnd cell_6t
Xbit_r72_c50 bl[50] br[50] wl[72] vdd gnd cell_6t
Xbit_r73_c50 bl[50] br[50] wl[73] vdd gnd cell_6t
Xbit_r74_c50 bl[50] br[50] wl[74] vdd gnd cell_6t
Xbit_r75_c50 bl[50] br[50] wl[75] vdd gnd cell_6t
Xbit_r76_c50 bl[50] br[50] wl[76] vdd gnd cell_6t
Xbit_r77_c50 bl[50] br[50] wl[77] vdd gnd cell_6t
Xbit_r78_c50 bl[50] br[50] wl[78] vdd gnd cell_6t
Xbit_r79_c50 bl[50] br[50] wl[79] vdd gnd cell_6t
Xbit_r80_c50 bl[50] br[50] wl[80] vdd gnd cell_6t
Xbit_r81_c50 bl[50] br[50] wl[81] vdd gnd cell_6t
Xbit_r82_c50 bl[50] br[50] wl[82] vdd gnd cell_6t
Xbit_r83_c50 bl[50] br[50] wl[83] vdd gnd cell_6t
Xbit_r84_c50 bl[50] br[50] wl[84] vdd gnd cell_6t
Xbit_r85_c50 bl[50] br[50] wl[85] vdd gnd cell_6t
Xbit_r86_c50 bl[50] br[50] wl[86] vdd gnd cell_6t
Xbit_r87_c50 bl[50] br[50] wl[87] vdd gnd cell_6t
Xbit_r88_c50 bl[50] br[50] wl[88] vdd gnd cell_6t
Xbit_r89_c50 bl[50] br[50] wl[89] vdd gnd cell_6t
Xbit_r90_c50 bl[50] br[50] wl[90] vdd gnd cell_6t
Xbit_r91_c50 bl[50] br[50] wl[91] vdd gnd cell_6t
Xbit_r92_c50 bl[50] br[50] wl[92] vdd gnd cell_6t
Xbit_r93_c50 bl[50] br[50] wl[93] vdd gnd cell_6t
Xbit_r94_c50 bl[50] br[50] wl[94] vdd gnd cell_6t
Xbit_r95_c50 bl[50] br[50] wl[95] vdd gnd cell_6t
Xbit_r96_c50 bl[50] br[50] wl[96] vdd gnd cell_6t
Xbit_r97_c50 bl[50] br[50] wl[97] vdd gnd cell_6t
Xbit_r98_c50 bl[50] br[50] wl[98] vdd gnd cell_6t
Xbit_r99_c50 bl[50] br[50] wl[99] vdd gnd cell_6t
Xbit_r100_c50 bl[50] br[50] wl[100] vdd gnd cell_6t
Xbit_r101_c50 bl[50] br[50] wl[101] vdd gnd cell_6t
Xbit_r102_c50 bl[50] br[50] wl[102] vdd gnd cell_6t
Xbit_r103_c50 bl[50] br[50] wl[103] vdd gnd cell_6t
Xbit_r104_c50 bl[50] br[50] wl[104] vdd gnd cell_6t
Xbit_r105_c50 bl[50] br[50] wl[105] vdd gnd cell_6t
Xbit_r106_c50 bl[50] br[50] wl[106] vdd gnd cell_6t
Xbit_r107_c50 bl[50] br[50] wl[107] vdd gnd cell_6t
Xbit_r108_c50 bl[50] br[50] wl[108] vdd gnd cell_6t
Xbit_r109_c50 bl[50] br[50] wl[109] vdd gnd cell_6t
Xbit_r110_c50 bl[50] br[50] wl[110] vdd gnd cell_6t
Xbit_r111_c50 bl[50] br[50] wl[111] vdd gnd cell_6t
Xbit_r112_c50 bl[50] br[50] wl[112] vdd gnd cell_6t
Xbit_r113_c50 bl[50] br[50] wl[113] vdd gnd cell_6t
Xbit_r114_c50 bl[50] br[50] wl[114] vdd gnd cell_6t
Xbit_r115_c50 bl[50] br[50] wl[115] vdd gnd cell_6t
Xbit_r116_c50 bl[50] br[50] wl[116] vdd gnd cell_6t
Xbit_r117_c50 bl[50] br[50] wl[117] vdd gnd cell_6t
Xbit_r118_c50 bl[50] br[50] wl[118] vdd gnd cell_6t
Xbit_r119_c50 bl[50] br[50] wl[119] vdd gnd cell_6t
Xbit_r120_c50 bl[50] br[50] wl[120] vdd gnd cell_6t
Xbit_r121_c50 bl[50] br[50] wl[121] vdd gnd cell_6t
Xbit_r122_c50 bl[50] br[50] wl[122] vdd gnd cell_6t
Xbit_r123_c50 bl[50] br[50] wl[123] vdd gnd cell_6t
Xbit_r124_c50 bl[50] br[50] wl[124] vdd gnd cell_6t
Xbit_r125_c50 bl[50] br[50] wl[125] vdd gnd cell_6t
Xbit_r126_c50 bl[50] br[50] wl[126] vdd gnd cell_6t
Xbit_r127_c50 bl[50] br[50] wl[127] vdd gnd cell_6t
Xbit_r128_c50 bl[50] br[50] wl[128] vdd gnd cell_6t
Xbit_r129_c50 bl[50] br[50] wl[129] vdd gnd cell_6t
Xbit_r130_c50 bl[50] br[50] wl[130] vdd gnd cell_6t
Xbit_r131_c50 bl[50] br[50] wl[131] vdd gnd cell_6t
Xbit_r132_c50 bl[50] br[50] wl[132] vdd gnd cell_6t
Xbit_r133_c50 bl[50] br[50] wl[133] vdd gnd cell_6t
Xbit_r134_c50 bl[50] br[50] wl[134] vdd gnd cell_6t
Xbit_r135_c50 bl[50] br[50] wl[135] vdd gnd cell_6t
Xbit_r136_c50 bl[50] br[50] wl[136] vdd gnd cell_6t
Xbit_r137_c50 bl[50] br[50] wl[137] vdd gnd cell_6t
Xbit_r138_c50 bl[50] br[50] wl[138] vdd gnd cell_6t
Xbit_r139_c50 bl[50] br[50] wl[139] vdd gnd cell_6t
Xbit_r140_c50 bl[50] br[50] wl[140] vdd gnd cell_6t
Xbit_r141_c50 bl[50] br[50] wl[141] vdd gnd cell_6t
Xbit_r142_c50 bl[50] br[50] wl[142] vdd gnd cell_6t
Xbit_r143_c50 bl[50] br[50] wl[143] vdd gnd cell_6t
Xbit_r144_c50 bl[50] br[50] wl[144] vdd gnd cell_6t
Xbit_r145_c50 bl[50] br[50] wl[145] vdd gnd cell_6t
Xbit_r146_c50 bl[50] br[50] wl[146] vdd gnd cell_6t
Xbit_r147_c50 bl[50] br[50] wl[147] vdd gnd cell_6t
Xbit_r148_c50 bl[50] br[50] wl[148] vdd gnd cell_6t
Xbit_r149_c50 bl[50] br[50] wl[149] vdd gnd cell_6t
Xbit_r150_c50 bl[50] br[50] wl[150] vdd gnd cell_6t
Xbit_r151_c50 bl[50] br[50] wl[151] vdd gnd cell_6t
Xbit_r152_c50 bl[50] br[50] wl[152] vdd gnd cell_6t
Xbit_r153_c50 bl[50] br[50] wl[153] vdd gnd cell_6t
Xbit_r154_c50 bl[50] br[50] wl[154] vdd gnd cell_6t
Xbit_r155_c50 bl[50] br[50] wl[155] vdd gnd cell_6t
Xbit_r156_c50 bl[50] br[50] wl[156] vdd gnd cell_6t
Xbit_r157_c50 bl[50] br[50] wl[157] vdd gnd cell_6t
Xbit_r158_c50 bl[50] br[50] wl[158] vdd gnd cell_6t
Xbit_r159_c50 bl[50] br[50] wl[159] vdd gnd cell_6t
Xbit_r160_c50 bl[50] br[50] wl[160] vdd gnd cell_6t
Xbit_r161_c50 bl[50] br[50] wl[161] vdd gnd cell_6t
Xbit_r162_c50 bl[50] br[50] wl[162] vdd gnd cell_6t
Xbit_r163_c50 bl[50] br[50] wl[163] vdd gnd cell_6t
Xbit_r164_c50 bl[50] br[50] wl[164] vdd gnd cell_6t
Xbit_r165_c50 bl[50] br[50] wl[165] vdd gnd cell_6t
Xbit_r166_c50 bl[50] br[50] wl[166] vdd gnd cell_6t
Xbit_r167_c50 bl[50] br[50] wl[167] vdd gnd cell_6t
Xbit_r168_c50 bl[50] br[50] wl[168] vdd gnd cell_6t
Xbit_r169_c50 bl[50] br[50] wl[169] vdd gnd cell_6t
Xbit_r170_c50 bl[50] br[50] wl[170] vdd gnd cell_6t
Xbit_r171_c50 bl[50] br[50] wl[171] vdd gnd cell_6t
Xbit_r172_c50 bl[50] br[50] wl[172] vdd gnd cell_6t
Xbit_r173_c50 bl[50] br[50] wl[173] vdd gnd cell_6t
Xbit_r174_c50 bl[50] br[50] wl[174] vdd gnd cell_6t
Xbit_r175_c50 bl[50] br[50] wl[175] vdd gnd cell_6t
Xbit_r176_c50 bl[50] br[50] wl[176] vdd gnd cell_6t
Xbit_r177_c50 bl[50] br[50] wl[177] vdd gnd cell_6t
Xbit_r178_c50 bl[50] br[50] wl[178] vdd gnd cell_6t
Xbit_r179_c50 bl[50] br[50] wl[179] vdd gnd cell_6t
Xbit_r180_c50 bl[50] br[50] wl[180] vdd gnd cell_6t
Xbit_r181_c50 bl[50] br[50] wl[181] vdd gnd cell_6t
Xbit_r182_c50 bl[50] br[50] wl[182] vdd gnd cell_6t
Xbit_r183_c50 bl[50] br[50] wl[183] vdd gnd cell_6t
Xbit_r184_c50 bl[50] br[50] wl[184] vdd gnd cell_6t
Xbit_r185_c50 bl[50] br[50] wl[185] vdd gnd cell_6t
Xbit_r186_c50 bl[50] br[50] wl[186] vdd gnd cell_6t
Xbit_r187_c50 bl[50] br[50] wl[187] vdd gnd cell_6t
Xbit_r188_c50 bl[50] br[50] wl[188] vdd gnd cell_6t
Xbit_r189_c50 bl[50] br[50] wl[189] vdd gnd cell_6t
Xbit_r190_c50 bl[50] br[50] wl[190] vdd gnd cell_6t
Xbit_r191_c50 bl[50] br[50] wl[191] vdd gnd cell_6t
Xbit_r192_c50 bl[50] br[50] wl[192] vdd gnd cell_6t
Xbit_r193_c50 bl[50] br[50] wl[193] vdd gnd cell_6t
Xbit_r194_c50 bl[50] br[50] wl[194] vdd gnd cell_6t
Xbit_r195_c50 bl[50] br[50] wl[195] vdd gnd cell_6t
Xbit_r196_c50 bl[50] br[50] wl[196] vdd gnd cell_6t
Xbit_r197_c50 bl[50] br[50] wl[197] vdd gnd cell_6t
Xbit_r198_c50 bl[50] br[50] wl[198] vdd gnd cell_6t
Xbit_r199_c50 bl[50] br[50] wl[199] vdd gnd cell_6t
Xbit_r200_c50 bl[50] br[50] wl[200] vdd gnd cell_6t
Xbit_r201_c50 bl[50] br[50] wl[201] vdd gnd cell_6t
Xbit_r202_c50 bl[50] br[50] wl[202] vdd gnd cell_6t
Xbit_r203_c50 bl[50] br[50] wl[203] vdd gnd cell_6t
Xbit_r204_c50 bl[50] br[50] wl[204] vdd gnd cell_6t
Xbit_r205_c50 bl[50] br[50] wl[205] vdd gnd cell_6t
Xbit_r206_c50 bl[50] br[50] wl[206] vdd gnd cell_6t
Xbit_r207_c50 bl[50] br[50] wl[207] vdd gnd cell_6t
Xbit_r208_c50 bl[50] br[50] wl[208] vdd gnd cell_6t
Xbit_r209_c50 bl[50] br[50] wl[209] vdd gnd cell_6t
Xbit_r210_c50 bl[50] br[50] wl[210] vdd gnd cell_6t
Xbit_r211_c50 bl[50] br[50] wl[211] vdd gnd cell_6t
Xbit_r212_c50 bl[50] br[50] wl[212] vdd gnd cell_6t
Xbit_r213_c50 bl[50] br[50] wl[213] vdd gnd cell_6t
Xbit_r214_c50 bl[50] br[50] wl[214] vdd gnd cell_6t
Xbit_r215_c50 bl[50] br[50] wl[215] vdd gnd cell_6t
Xbit_r216_c50 bl[50] br[50] wl[216] vdd gnd cell_6t
Xbit_r217_c50 bl[50] br[50] wl[217] vdd gnd cell_6t
Xbit_r218_c50 bl[50] br[50] wl[218] vdd gnd cell_6t
Xbit_r219_c50 bl[50] br[50] wl[219] vdd gnd cell_6t
Xbit_r220_c50 bl[50] br[50] wl[220] vdd gnd cell_6t
Xbit_r221_c50 bl[50] br[50] wl[221] vdd gnd cell_6t
Xbit_r222_c50 bl[50] br[50] wl[222] vdd gnd cell_6t
Xbit_r223_c50 bl[50] br[50] wl[223] vdd gnd cell_6t
Xbit_r224_c50 bl[50] br[50] wl[224] vdd gnd cell_6t
Xbit_r225_c50 bl[50] br[50] wl[225] vdd gnd cell_6t
Xbit_r226_c50 bl[50] br[50] wl[226] vdd gnd cell_6t
Xbit_r227_c50 bl[50] br[50] wl[227] vdd gnd cell_6t
Xbit_r228_c50 bl[50] br[50] wl[228] vdd gnd cell_6t
Xbit_r229_c50 bl[50] br[50] wl[229] vdd gnd cell_6t
Xbit_r230_c50 bl[50] br[50] wl[230] vdd gnd cell_6t
Xbit_r231_c50 bl[50] br[50] wl[231] vdd gnd cell_6t
Xbit_r232_c50 bl[50] br[50] wl[232] vdd gnd cell_6t
Xbit_r233_c50 bl[50] br[50] wl[233] vdd gnd cell_6t
Xbit_r234_c50 bl[50] br[50] wl[234] vdd gnd cell_6t
Xbit_r235_c50 bl[50] br[50] wl[235] vdd gnd cell_6t
Xbit_r236_c50 bl[50] br[50] wl[236] vdd gnd cell_6t
Xbit_r237_c50 bl[50] br[50] wl[237] vdd gnd cell_6t
Xbit_r238_c50 bl[50] br[50] wl[238] vdd gnd cell_6t
Xbit_r239_c50 bl[50] br[50] wl[239] vdd gnd cell_6t
Xbit_r240_c50 bl[50] br[50] wl[240] vdd gnd cell_6t
Xbit_r241_c50 bl[50] br[50] wl[241] vdd gnd cell_6t
Xbit_r242_c50 bl[50] br[50] wl[242] vdd gnd cell_6t
Xbit_r243_c50 bl[50] br[50] wl[243] vdd gnd cell_6t
Xbit_r244_c50 bl[50] br[50] wl[244] vdd gnd cell_6t
Xbit_r245_c50 bl[50] br[50] wl[245] vdd gnd cell_6t
Xbit_r246_c50 bl[50] br[50] wl[246] vdd gnd cell_6t
Xbit_r247_c50 bl[50] br[50] wl[247] vdd gnd cell_6t
Xbit_r248_c50 bl[50] br[50] wl[248] vdd gnd cell_6t
Xbit_r249_c50 bl[50] br[50] wl[249] vdd gnd cell_6t
Xbit_r250_c50 bl[50] br[50] wl[250] vdd gnd cell_6t
Xbit_r251_c50 bl[50] br[50] wl[251] vdd gnd cell_6t
Xbit_r252_c50 bl[50] br[50] wl[252] vdd gnd cell_6t
Xbit_r253_c50 bl[50] br[50] wl[253] vdd gnd cell_6t
Xbit_r254_c50 bl[50] br[50] wl[254] vdd gnd cell_6t
Xbit_r255_c50 bl[50] br[50] wl[255] vdd gnd cell_6t
Xbit_r0_c51 bl[51] br[51] wl[0] vdd gnd cell_6t
Xbit_r1_c51 bl[51] br[51] wl[1] vdd gnd cell_6t
Xbit_r2_c51 bl[51] br[51] wl[2] vdd gnd cell_6t
Xbit_r3_c51 bl[51] br[51] wl[3] vdd gnd cell_6t
Xbit_r4_c51 bl[51] br[51] wl[4] vdd gnd cell_6t
Xbit_r5_c51 bl[51] br[51] wl[5] vdd gnd cell_6t
Xbit_r6_c51 bl[51] br[51] wl[6] vdd gnd cell_6t
Xbit_r7_c51 bl[51] br[51] wl[7] vdd gnd cell_6t
Xbit_r8_c51 bl[51] br[51] wl[8] vdd gnd cell_6t
Xbit_r9_c51 bl[51] br[51] wl[9] vdd gnd cell_6t
Xbit_r10_c51 bl[51] br[51] wl[10] vdd gnd cell_6t
Xbit_r11_c51 bl[51] br[51] wl[11] vdd gnd cell_6t
Xbit_r12_c51 bl[51] br[51] wl[12] vdd gnd cell_6t
Xbit_r13_c51 bl[51] br[51] wl[13] vdd gnd cell_6t
Xbit_r14_c51 bl[51] br[51] wl[14] vdd gnd cell_6t
Xbit_r15_c51 bl[51] br[51] wl[15] vdd gnd cell_6t
Xbit_r16_c51 bl[51] br[51] wl[16] vdd gnd cell_6t
Xbit_r17_c51 bl[51] br[51] wl[17] vdd gnd cell_6t
Xbit_r18_c51 bl[51] br[51] wl[18] vdd gnd cell_6t
Xbit_r19_c51 bl[51] br[51] wl[19] vdd gnd cell_6t
Xbit_r20_c51 bl[51] br[51] wl[20] vdd gnd cell_6t
Xbit_r21_c51 bl[51] br[51] wl[21] vdd gnd cell_6t
Xbit_r22_c51 bl[51] br[51] wl[22] vdd gnd cell_6t
Xbit_r23_c51 bl[51] br[51] wl[23] vdd gnd cell_6t
Xbit_r24_c51 bl[51] br[51] wl[24] vdd gnd cell_6t
Xbit_r25_c51 bl[51] br[51] wl[25] vdd gnd cell_6t
Xbit_r26_c51 bl[51] br[51] wl[26] vdd gnd cell_6t
Xbit_r27_c51 bl[51] br[51] wl[27] vdd gnd cell_6t
Xbit_r28_c51 bl[51] br[51] wl[28] vdd gnd cell_6t
Xbit_r29_c51 bl[51] br[51] wl[29] vdd gnd cell_6t
Xbit_r30_c51 bl[51] br[51] wl[30] vdd gnd cell_6t
Xbit_r31_c51 bl[51] br[51] wl[31] vdd gnd cell_6t
Xbit_r32_c51 bl[51] br[51] wl[32] vdd gnd cell_6t
Xbit_r33_c51 bl[51] br[51] wl[33] vdd gnd cell_6t
Xbit_r34_c51 bl[51] br[51] wl[34] vdd gnd cell_6t
Xbit_r35_c51 bl[51] br[51] wl[35] vdd gnd cell_6t
Xbit_r36_c51 bl[51] br[51] wl[36] vdd gnd cell_6t
Xbit_r37_c51 bl[51] br[51] wl[37] vdd gnd cell_6t
Xbit_r38_c51 bl[51] br[51] wl[38] vdd gnd cell_6t
Xbit_r39_c51 bl[51] br[51] wl[39] vdd gnd cell_6t
Xbit_r40_c51 bl[51] br[51] wl[40] vdd gnd cell_6t
Xbit_r41_c51 bl[51] br[51] wl[41] vdd gnd cell_6t
Xbit_r42_c51 bl[51] br[51] wl[42] vdd gnd cell_6t
Xbit_r43_c51 bl[51] br[51] wl[43] vdd gnd cell_6t
Xbit_r44_c51 bl[51] br[51] wl[44] vdd gnd cell_6t
Xbit_r45_c51 bl[51] br[51] wl[45] vdd gnd cell_6t
Xbit_r46_c51 bl[51] br[51] wl[46] vdd gnd cell_6t
Xbit_r47_c51 bl[51] br[51] wl[47] vdd gnd cell_6t
Xbit_r48_c51 bl[51] br[51] wl[48] vdd gnd cell_6t
Xbit_r49_c51 bl[51] br[51] wl[49] vdd gnd cell_6t
Xbit_r50_c51 bl[51] br[51] wl[50] vdd gnd cell_6t
Xbit_r51_c51 bl[51] br[51] wl[51] vdd gnd cell_6t
Xbit_r52_c51 bl[51] br[51] wl[52] vdd gnd cell_6t
Xbit_r53_c51 bl[51] br[51] wl[53] vdd gnd cell_6t
Xbit_r54_c51 bl[51] br[51] wl[54] vdd gnd cell_6t
Xbit_r55_c51 bl[51] br[51] wl[55] vdd gnd cell_6t
Xbit_r56_c51 bl[51] br[51] wl[56] vdd gnd cell_6t
Xbit_r57_c51 bl[51] br[51] wl[57] vdd gnd cell_6t
Xbit_r58_c51 bl[51] br[51] wl[58] vdd gnd cell_6t
Xbit_r59_c51 bl[51] br[51] wl[59] vdd gnd cell_6t
Xbit_r60_c51 bl[51] br[51] wl[60] vdd gnd cell_6t
Xbit_r61_c51 bl[51] br[51] wl[61] vdd gnd cell_6t
Xbit_r62_c51 bl[51] br[51] wl[62] vdd gnd cell_6t
Xbit_r63_c51 bl[51] br[51] wl[63] vdd gnd cell_6t
Xbit_r64_c51 bl[51] br[51] wl[64] vdd gnd cell_6t
Xbit_r65_c51 bl[51] br[51] wl[65] vdd gnd cell_6t
Xbit_r66_c51 bl[51] br[51] wl[66] vdd gnd cell_6t
Xbit_r67_c51 bl[51] br[51] wl[67] vdd gnd cell_6t
Xbit_r68_c51 bl[51] br[51] wl[68] vdd gnd cell_6t
Xbit_r69_c51 bl[51] br[51] wl[69] vdd gnd cell_6t
Xbit_r70_c51 bl[51] br[51] wl[70] vdd gnd cell_6t
Xbit_r71_c51 bl[51] br[51] wl[71] vdd gnd cell_6t
Xbit_r72_c51 bl[51] br[51] wl[72] vdd gnd cell_6t
Xbit_r73_c51 bl[51] br[51] wl[73] vdd gnd cell_6t
Xbit_r74_c51 bl[51] br[51] wl[74] vdd gnd cell_6t
Xbit_r75_c51 bl[51] br[51] wl[75] vdd gnd cell_6t
Xbit_r76_c51 bl[51] br[51] wl[76] vdd gnd cell_6t
Xbit_r77_c51 bl[51] br[51] wl[77] vdd gnd cell_6t
Xbit_r78_c51 bl[51] br[51] wl[78] vdd gnd cell_6t
Xbit_r79_c51 bl[51] br[51] wl[79] vdd gnd cell_6t
Xbit_r80_c51 bl[51] br[51] wl[80] vdd gnd cell_6t
Xbit_r81_c51 bl[51] br[51] wl[81] vdd gnd cell_6t
Xbit_r82_c51 bl[51] br[51] wl[82] vdd gnd cell_6t
Xbit_r83_c51 bl[51] br[51] wl[83] vdd gnd cell_6t
Xbit_r84_c51 bl[51] br[51] wl[84] vdd gnd cell_6t
Xbit_r85_c51 bl[51] br[51] wl[85] vdd gnd cell_6t
Xbit_r86_c51 bl[51] br[51] wl[86] vdd gnd cell_6t
Xbit_r87_c51 bl[51] br[51] wl[87] vdd gnd cell_6t
Xbit_r88_c51 bl[51] br[51] wl[88] vdd gnd cell_6t
Xbit_r89_c51 bl[51] br[51] wl[89] vdd gnd cell_6t
Xbit_r90_c51 bl[51] br[51] wl[90] vdd gnd cell_6t
Xbit_r91_c51 bl[51] br[51] wl[91] vdd gnd cell_6t
Xbit_r92_c51 bl[51] br[51] wl[92] vdd gnd cell_6t
Xbit_r93_c51 bl[51] br[51] wl[93] vdd gnd cell_6t
Xbit_r94_c51 bl[51] br[51] wl[94] vdd gnd cell_6t
Xbit_r95_c51 bl[51] br[51] wl[95] vdd gnd cell_6t
Xbit_r96_c51 bl[51] br[51] wl[96] vdd gnd cell_6t
Xbit_r97_c51 bl[51] br[51] wl[97] vdd gnd cell_6t
Xbit_r98_c51 bl[51] br[51] wl[98] vdd gnd cell_6t
Xbit_r99_c51 bl[51] br[51] wl[99] vdd gnd cell_6t
Xbit_r100_c51 bl[51] br[51] wl[100] vdd gnd cell_6t
Xbit_r101_c51 bl[51] br[51] wl[101] vdd gnd cell_6t
Xbit_r102_c51 bl[51] br[51] wl[102] vdd gnd cell_6t
Xbit_r103_c51 bl[51] br[51] wl[103] vdd gnd cell_6t
Xbit_r104_c51 bl[51] br[51] wl[104] vdd gnd cell_6t
Xbit_r105_c51 bl[51] br[51] wl[105] vdd gnd cell_6t
Xbit_r106_c51 bl[51] br[51] wl[106] vdd gnd cell_6t
Xbit_r107_c51 bl[51] br[51] wl[107] vdd gnd cell_6t
Xbit_r108_c51 bl[51] br[51] wl[108] vdd gnd cell_6t
Xbit_r109_c51 bl[51] br[51] wl[109] vdd gnd cell_6t
Xbit_r110_c51 bl[51] br[51] wl[110] vdd gnd cell_6t
Xbit_r111_c51 bl[51] br[51] wl[111] vdd gnd cell_6t
Xbit_r112_c51 bl[51] br[51] wl[112] vdd gnd cell_6t
Xbit_r113_c51 bl[51] br[51] wl[113] vdd gnd cell_6t
Xbit_r114_c51 bl[51] br[51] wl[114] vdd gnd cell_6t
Xbit_r115_c51 bl[51] br[51] wl[115] vdd gnd cell_6t
Xbit_r116_c51 bl[51] br[51] wl[116] vdd gnd cell_6t
Xbit_r117_c51 bl[51] br[51] wl[117] vdd gnd cell_6t
Xbit_r118_c51 bl[51] br[51] wl[118] vdd gnd cell_6t
Xbit_r119_c51 bl[51] br[51] wl[119] vdd gnd cell_6t
Xbit_r120_c51 bl[51] br[51] wl[120] vdd gnd cell_6t
Xbit_r121_c51 bl[51] br[51] wl[121] vdd gnd cell_6t
Xbit_r122_c51 bl[51] br[51] wl[122] vdd gnd cell_6t
Xbit_r123_c51 bl[51] br[51] wl[123] vdd gnd cell_6t
Xbit_r124_c51 bl[51] br[51] wl[124] vdd gnd cell_6t
Xbit_r125_c51 bl[51] br[51] wl[125] vdd gnd cell_6t
Xbit_r126_c51 bl[51] br[51] wl[126] vdd gnd cell_6t
Xbit_r127_c51 bl[51] br[51] wl[127] vdd gnd cell_6t
Xbit_r128_c51 bl[51] br[51] wl[128] vdd gnd cell_6t
Xbit_r129_c51 bl[51] br[51] wl[129] vdd gnd cell_6t
Xbit_r130_c51 bl[51] br[51] wl[130] vdd gnd cell_6t
Xbit_r131_c51 bl[51] br[51] wl[131] vdd gnd cell_6t
Xbit_r132_c51 bl[51] br[51] wl[132] vdd gnd cell_6t
Xbit_r133_c51 bl[51] br[51] wl[133] vdd gnd cell_6t
Xbit_r134_c51 bl[51] br[51] wl[134] vdd gnd cell_6t
Xbit_r135_c51 bl[51] br[51] wl[135] vdd gnd cell_6t
Xbit_r136_c51 bl[51] br[51] wl[136] vdd gnd cell_6t
Xbit_r137_c51 bl[51] br[51] wl[137] vdd gnd cell_6t
Xbit_r138_c51 bl[51] br[51] wl[138] vdd gnd cell_6t
Xbit_r139_c51 bl[51] br[51] wl[139] vdd gnd cell_6t
Xbit_r140_c51 bl[51] br[51] wl[140] vdd gnd cell_6t
Xbit_r141_c51 bl[51] br[51] wl[141] vdd gnd cell_6t
Xbit_r142_c51 bl[51] br[51] wl[142] vdd gnd cell_6t
Xbit_r143_c51 bl[51] br[51] wl[143] vdd gnd cell_6t
Xbit_r144_c51 bl[51] br[51] wl[144] vdd gnd cell_6t
Xbit_r145_c51 bl[51] br[51] wl[145] vdd gnd cell_6t
Xbit_r146_c51 bl[51] br[51] wl[146] vdd gnd cell_6t
Xbit_r147_c51 bl[51] br[51] wl[147] vdd gnd cell_6t
Xbit_r148_c51 bl[51] br[51] wl[148] vdd gnd cell_6t
Xbit_r149_c51 bl[51] br[51] wl[149] vdd gnd cell_6t
Xbit_r150_c51 bl[51] br[51] wl[150] vdd gnd cell_6t
Xbit_r151_c51 bl[51] br[51] wl[151] vdd gnd cell_6t
Xbit_r152_c51 bl[51] br[51] wl[152] vdd gnd cell_6t
Xbit_r153_c51 bl[51] br[51] wl[153] vdd gnd cell_6t
Xbit_r154_c51 bl[51] br[51] wl[154] vdd gnd cell_6t
Xbit_r155_c51 bl[51] br[51] wl[155] vdd gnd cell_6t
Xbit_r156_c51 bl[51] br[51] wl[156] vdd gnd cell_6t
Xbit_r157_c51 bl[51] br[51] wl[157] vdd gnd cell_6t
Xbit_r158_c51 bl[51] br[51] wl[158] vdd gnd cell_6t
Xbit_r159_c51 bl[51] br[51] wl[159] vdd gnd cell_6t
Xbit_r160_c51 bl[51] br[51] wl[160] vdd gnd cell_6t
Xbit_r161_c51 bl[51] br[51] wl[161] vdd gnd cell_6t
Xbit_r162_c51 bl[51] br[51] wl[162] vdd gnd cell_6t
Xbit_r163_c51 bl[51] br[51] wl[163] vdd gnd cell_6t
Xbit_r164_c51 bl[51] br[51] wl[164] vdd gnd cell_6t
Xbit_r165_c51 bl[51] br[51] wl[165] vdd gnd cell_6t
Xbit_r166_c51 bl[51] br[51] wl[166] vdd gnd cell_6t
Xbit_r167_c51 bl[51] br[51] wl[167] vdd gnd cell_6t
Xbit_r168_c51 bl[51] br[51] wl[168] vdd gnd cell_6t
Xbit_r169_c51 bl[51] br[51] wl[169] vdd gnd cell_6t
Xbit_r170_c51 bl[51] br[51] wl[170] vdd gnd cell_6t
Xbit_r171_c51 bl[51] br[51] wl[171] vdd gnd cell_6t
Xbit_r172_c51 bl[51] br[51] wl[172] vdd gnd cell_6t
Xbit_r173_c51 bl[51] br[51] wl[173] vdd gnd cell_6t
Xbit_r174_c51 bl[51] br[51] wl[174] vdd gnd cell_6t
Xbit_r175_c51 bl[51] br[51] wl[175] vdd gnd cell_6t
Xbit_r176_c51 bl[51] br[51] wl[176] vdd gnd cell_6t
Xbit_r177_c51 bl[51] br[51] wl[177] vdd gnd cell_6t
Xbit_r178_c51 bl[51] br[51] wl[178] vdd gnd cell_6t
Xbit_r179_c51 bl[51] br[51] wl[179] vdd gnd cell_6t
Xbit_r180_c51 bl[51] br[51] wl[180] vdd gnd cell_6t
Xbit_r181_c51 bl[51] br[51] wl[181] vdd gnd cell_6t
Xbit_r182_c51 bl[51] br[51] wl[182] vdd gnd cell_6t
Xbit_r183_c51 bl[51] br[51] wl[183] vdd gnd cell_6t
Xbit_r184_c51 bl[51] br[51] wl[184] vdd gnd cell_6t
Xbit_r185_c51 bl[51] br[51] wl[185] vdd gnd cell_6t
Xbit_r186_c51 bl[51] br[51] wl[186] vdd gnd cell_6t
Xbit_r187_c51 bl[51] br[51] wl[187] vdd gnd cell_6t
Xbit_r188_c51 bl[51] br[51] wl[188] vdd gnd cell_6t
Xbit_r189_c51 bl[51] br[51] wl[189] vdd gnd cell_6t
Xbit_r190_c51 bl[51] br[51] wl[190] vdd gnd cell_6t
Xbit_r191_c51 bl[51] br[51] wl[191] vdd gnd cell_6t
Xbit_r192_c51 bl[51] br[51] wl[192] vdd gnd cell_6t
Xbit_r193_c51 bl[51] br[51] wl[193] vdd gnd cell_6t
Xbit_r194_c51 bl[51] br[51] wl[194] vdd gnd cell_6t
Xbit_r195_c51 bl[51] br[51] wl[195] vdd gnd cell_6t
Xbit_r196_c51 bl[51] br[51] wl[196] vdd gnd cell_6t
Xbit_r197_c51 bl[51] br[51] wl[197] vdd gnd cell_6t
Xbit_r198_c51 bl[51] br[51] wl[198] vdd gnd cell_6t
Xbit_r199_c51 bl[51] br[51] wl[199] vdd gnd cell_6t
Xbit_r200_c51 bl[51] br[51] wl[200] vdd gnd cell_6t
Xbit_r201_c51 bl[51] br[51] wl[201] vdd gnd cell_6t
Xbit_r202_c51 bl[51] br[51] wl[202] vdd gnd cell_6t
Xbit_r203_c51 bl[51] br[51] wl[203] vdd gnd cell_6t
Xbit_r204_c51 bl[51] br[51] wl[204] vdd gnd cell_6t
Xbit_r205_c51 bl[51] br[51] wl[205] vdd gnd cell_6t
Xbit_r206_c51 bl[51] br[51] wl[206] vdd gnd cell_6t
Xbit_r207_c51 bl[51] br[51] wl[207] vdd gnd cell_6t
Xbit_r208_c51 bl[51] br[51] wl[208] vdd gnd cell_6t
Xbit_r209_c51 bl[51] br[51] wl[209] vdd gnd cell_6t
Xbit_r210_c51 bl[51] br[51] wl[210] vdd gnd cell_6t
Xbit_r211_c51 bl[51] br[51] wl[211] vdd gnd cell_6t
Xbit_r212_c51 bl[51] br[51] wl[212] vdd gnd cell_6t
Xbit_r213_c51 bl[51] br[51] wl[213] vdd gnd cell_6t
Xbit_r214_c51 bl[51] br[51] wl[214] vdd gnd cell_6t
Xbit_r215_c51 bl[51] br[51] wl[215] vdd gnd cell_6t
Xbit_r216_c51 bl[51] br[51] wl[216] vdd gnd cell_6t
Xbit_r217_c51 bl[51] br[51] wl[217] vdd gnd cell_6t
Xbit_r218_c51 bl[51] br[51] wl[218] vdd gnd cell_6t
Xbit_r219_c51 bl[51] br[51] wl[219] vdd gnd cell_6t
Xbit_r220_c51 bl[51] br[51] wl[220] vdd gnd cell_6t
Xbit_r221_c51 bl[51] br[51] wl[221] vdd gnd cell_6t
Xbit_r222_c51 bl[51] br[51] wl[222] vdd gnd cell_6t
Xbit_r223_c51 bl[51] br[51] wl[223] vdd gnd cell_6t
Xbit_r224_c51 bl[51] br[51] wl[224] vdd gnd cell_6t
Xbit_r225_c51 bl[51] br[51] wl[225] vdd gnd cell_6t
Xbit_r226_c51 bl[51] br[51] wl[226] vdd gnd cell_6t
Xbit_r227_c51 bl[51] br[51] wl[227] vdd gnd cell_6t
Xbit_r228_c51 bl[51] br[51] wl[228] vdd gnd cell_6t
Xbit_r229_c51 bl[51] br[51] wl[229] vdd gnd cell_6t
Xbit_r230_c51 bl[51] br[51] wl[230] vdd gnd cell_6t
Xbit_r231_c51 bl[51] br[51] wl[231] vdd gnd cell_6t
Xbit_r232_c51 bl[51] br[51] wl[232] vdd gnd cell_6t
Xbit_r233_c51 bl[51] br[51] wl[233] vdd gnd cell_6t
Xbit_r234_c51 bl[51] br[51] wl[234] vdd gnd cell_6t
Xbit_r235_c51 bl[51] br[51] wl[235] vdd gnd cell_6t
Xbit_r236_c51 bl[51] br[51] wl[236] vdd gnd cell_6t
Xbit_r237_c51 bl[51] br[51] wl[237] vdd gnd cell_6t
Xbit_r238_c51 bl[51] br[51] wl[238] vdd gnd cell_6t
Xbit_r239_c51 bl[51] br[51] wl[239] vdd gnd cell_6t
Xbit_r240_c51 bl[51] br[51] wl[240] vdd gnd cell_6t
Xbit_r241_c51 bl[51] br[51] wl[241] vdd gnd cell_6t
Xbit_r242_c51 bl[51] br[51] wl[242] vdd gnd cell_6t
Xbit_r243_c51 bl[51] br[51] wl[243] vdd gnd cell_6t
Xbit_r244_c51 bl[51] br[51] wl[244] vdd gnd cell_6t
Xbit_r245_c51 bl[51] br[51] wl[245] vdd gnd cell_6t
Xbit_r246_c51 bl[51] br[51] wl[246] vdd gnd cell_6t
Xbit_r247_c51 bl[51] br[51] wl[247] vdd gnd cell_6t
Xbit_r248_c51 bl[51] br[51] wl[248] vdd gnd cell_6t
Xbit_r249_c51 bl[51] br[51] wl[249] vdd gnd cell_6t
Xbit_r250_c51 bl[51] br[51] wl[250] vdd gnd cell_6t
Xbit_r251_c51 bl[51] br[51] wl[251] vdd gnd cell_6t
Xbit_r252_c51 bl[51] br[51] wl[252] vdd gnd cell_6t
Xbit_r253_c51 bl[51] br[51] wl[253] vdd gnd cell_6t
Xbit_r254_c51 bl[51] br[51] wl[254] vdd gnd cell_6t
Xbit_r255_c51 bl[51] br[51] wl[255] vdd gnd cell_6t
Xbit_r0_c52 bl[52] br[52] wl[0] vdd gnd cell_6t
Xbit_r1_c52 bl[52] br[52] wl[1] vdd gnd cell_6t
Xbit_r2_c52 bl[52] br[52] wl[2] vdd gnd cell_6t
Xbit_r3_c52 bl[52] br[52] wl[3] vdd gnd cell_6t
Xbit_r4_c52 bl[52] br[52] wl[4] vdd gnd cell_6t
Xbit_r5_c52 bl[52] br[52] wl[5] vdd gnd cell_6t
Xbit_r6_c52 bl[52] br[52] wl[6] vdd gnd cell_6t
Xbit_r7_c52 bl[52] br[52] wl[7] vdd gnd cell_6t
Xbit_r8_c52 bl[52] br[52] wl[8] vdd gnd cell_6t
Xbit_r9_c52 bl[52] br[52] wl[9] vdd gnd cell_6t
Xbit_r10_c52 bl[52] br[52] wl[10] vdd gnd cell_6t
Xbit_r11_c52 bl[52] br[52] wl[11] vdd gnd cell_6t
Xbit_r12_c52 bl[52] br[52] wl[12] vdd gnd cell_6t
Xbit_r13_c52 bl[52] br[52] wl[13] vdd gnd cell_6t
Xbit_r14_c52 bl[52] br[52] wl[14] vdd gnd cell_6t
Xbit_r15_c52 bl[52] br[52] wl[15] vdd gnd cell_6t
Xbit_r16_c52 bl[52] br[52] wl[16] vdd gnd cell_6t
Xbit_r17_c52 bl[52] br[52] wl[17] vdd gnd cell_6t
Xbit_r18_c52 bl[52] br[52] wl[18] vdd gnd cell_6t
Xbit_r19_c52 bl[52] br[52] wl[19] vdd gnd cell_6t
Xbit_r20_c52 bl[52] br[52] wl[20] vdd gnd cell_6t
Xbit_r21_c52 bl[52] br[52] wl[21] vdd gnd cell_6t
Xbit_r22_c52 bl[52] br[52] wl[22] vdd gnd cell_6t
Xbit_r23_c52 bl[52] br[52] wl[23] vdd gnd cell_6t
Xbit_r24_c52 bl[52] br[52] wl[24] vdd gnd cell_6t
Xbit_r25_c52 bl[52] br[52] wl[25] vdd gnd cell_6t
Xbit_r26_c52 bl[52] br[52] wl[26] vdd gnd cell_6t
Xbit_r27_c52 bl[52] br[52] wl[27] vdd gnd cell_6t
Xbit_r28_c52 bl[52] br[52] wl[28] vdd gnd cell_6t
Xbit_r29_c52 bl[52] br[52] wl[29] vdd gnd cell_6t
Xbit_r30_c52 bl[52] br[52] wl[30] vdd gnd cell_6t
Xbit_r31_c52 bl[52] br[52] wl[31] vdd gnd cell_6t
Xbit_r32_c52 bl[52] br[52] wl[32] vdd gnd cell_6t
Xbit_r33_c52 bl[52] br[52] wl[33] vdd gnd cell_6t
Xbit_r34_c52 bl[52] br[52] wl[34] vdd gnd cell_6t
Xbit_r35_c52 bl[52] br[52] wl[35] vdd gnd cell_6t
Xbit_r36_c52 bl[52] br[52] wl[36] vdd gnd cell_6t
Xbit_r37_c52 bl[52] br[52] wl[37] vdd gnd cell_6t
Xbit_r38_c52 bl[52] br[52] wl[38] vdd gnd cell_6t
Xbit_r39_c52 bl[52] br[52] wl[39] vdd gnd cell_6t
Xbit_r40_c52 bl[52] br[52] wl[40] vdd gnd cell_6t
Xbit_r41_c52 bl[52] br[52] wl[41] vdd gnd cell_6t
Xbit_r42_c52 bl[52] br[52] wl[42] vdd gnd cell_6t
Xbit_r43_c52 bl[52] br[52] wl[43] vdd gnd cell_6t
Xbit_r44_c52 bl[52] br[52] wl[44] vdd gnd cell_6t
Xbit_r45_c52 bl[52] br[52] wl[45] vdd gnd cell_6t
Xbit_r46_c52 bl[52] br[52] wl[46] vdd gnd cell_6t
Xbit_r47_c52 bl[52] br[52] wl[47] vdd gnd cell_6t
Xbit_r48_c52 bl[52] br[52] wl[48] vdd gnd cell_6t
Xbit_r49_c52 bl[52] br[52] wl[49] vdd gnd cell_6t
Xbit_r50_c52 bl[52] br[52] wl[50] vdd gnd cell_6t
Xbit_r51_c52 bl[52] br[52] wl[51] vdd gnd cell_6t
Xbit_r52_c52 bl[52] br[52] wl[52] vdd gnd cell_6t
Xbit_r53_c52 bl[52] br[52] wl[53] vdd gnd cell_6t
Xbit_r54_c52 bl[52] br[52] wl[54] vdd gnd cell_6t
Xbit_r55_c52 bl[52] br[52] wl[55] vdd gnd cell_6t
Xbit_r56_c52 bl[52] br[52] wl[56] vdd gnd cell_6t
Xbit_r57_c52 bl[52] br[52] wl[57] vdd gnd cell_6t
Xbit_r58_c52 bl[52] br[52] wl[58] vdd gnd cell_6t
Xbit_r59_c52 bl[52] br[52] wl[59] vdd gnd cell_6t
Xbit_r60_c52 bl[52] br[52] wl[60] vdd gnd cell_6t
Xbit_r61_c52 bl[52] br[52] wl[61] vdd gnd cell_6t
Xbit_r62_c52 bl[52] br[52] wl[62] vdd gnd cell_6t
Xbit_r63_c52 bl[52] br[52] wl[63] vdd gnd cell_6t
Xbit_r64_c52 bl[52] br[52] wl[64] vdd gnd cell_6t
Xbit_r65_c52 bl[52] br[52] wl[65] vdd gnd cell_6t
Xbit_r66_c52 bl[52] br[52] wl[66] vdd gnd cell_6t
Xbit_r67_c52 bl[52] br[52] wl[67] vdd gnd cell_6t
Xbit_r68_c52 bl[52] br[52] wl[68] vdd gnd cell_6t
Xbit_r69_c52 bl[52] br[52] wl[69] vdd gnd cell_6t
Xbit_r70_c52 bl[52] br[52] wl[70] vdd gnd cell_6t
Xbit_r71_c52 bl[52] br[52] wl[71] vdd gnd cell_6t
Xbit_r72_c52 bl[52] br[52] wl[72] vdd gnd cell_6t
Xbit_r73_c52 bl[52] br[52] wl[73] vdd gnd cell_6t
Xbit_r74_c52 bl[52] br[52] wl[74] vdd gnd cell_6t
Xbit_r75_c52 bl[52] br[52] wl[75] vdd gnd cell_6t
Xbit_r76_c52 bl[52] br[52] wl[76] vdd gnd cell_6t
Xbit_r77_c52 bl[52] br[52] wl[77] vdd gnd cell_6t
Xbit_r78_c52 bl[52] br[52] wl[78] vdd gnd cell_6t
Xbit_r79_c52 bl[52] br[52] wl[79] vdd gnd cell_6t
Xbit_r80_c52 bl[52] br[52] wl[80] vdd gnd cell_6t
Xbit_r81_c52 bl[52] br[52] wl[81] vdd gnd cell_6t
Xbit_r82_c52 bl[52] br[52] wl[82] vdd gnd cell_6t
Xbit_r83_c52 bl[52] br[52] wl[83] vdd gnd cell_6t
Xbit_r84_c52 bl[52] br[52] wl[84] vdd gnd cell_6t
Xbit_r85_c52 bl[52] br[52] wl[85] vdd gnd cell_6t
Xbit_r86_c52 bl[52] br[52] wl[86] vdd gnd cell_6t
Xbit_r87_c52 bl[52] br[52] wl[87] vdd gnd cell_6t
Xbit_r88_c52 bl[52] br[52] wl[88] vdd gnd cell_6t
Xbit_r89_c52 bl[52] br[52] wl[89] vdd gnd cell_6t
Xbit_r90_c52 bl[52] br[52] wl[90] vdd gnd cell_6t
Xbit_r91_c52 bl[52] br[52] wl[91] vdd gnd cell_6t
Xbit_r92_c52 bl[52] br[52] wl[92] vdd gnd cell_6t
Xbit_r93_c52 bl[52] br[52] wl[93] vdd gnd cell_6t
Xbit_r94_c52 bl[52] br[52] wl[94] vdd gnd cell_6t
Xbit_r95_c52 bl[52] br[52] wl[95] vdd gnd cell_6t
Xbit_r96_c52 bl[52] br[52] wl[96] vdd gnd cell_6t
Xbit_r97_c52 bl[52] br[52] wl[97] vdd gnd cell_6t
Xbit_r98_c52 bl[52] br[52] wl[98] vdd gnd cell_6t
Xbit_r99_c52 bl[52] br[52] wl[99] vdd gnd cell_6t
Xbit_r100_c52 bl[52] br[52] wl[100] vdd gnd cell_6t
Xbit_r101_c52 bl[52] br[52] wl[101] vdd gnd cell_6t
Xbit_r102_c52 bl[52] br[52] wl[102] vdd gnd cell_6t
Xbit_r103_c52 bl[52] br[52] wl[103] vdd gnd cell_6t
Xbit_r104_c52 bl[52] br[52] wl[104] vdd gnd cell_6t
Xbit_r105_c52 bl[52] br[52] wl[105] vdd gnd cell_6t
Xbit_r106_c52 bl[52] br[52] wl[106] vdd gnd cell_6t
Xbit_r107_c52 bl[52] br[52] wl[107] vdd gnd cell_6t
Xbit_r108_c52 bl[52] br[52] wl[108] vdd gnd cell_6t
Xbit_r109_c52 bl[52] br[52] wl[109] vdd gnd cell_6t
Xbit_r110_c52 bl[52] br[52] wl[110] vdd gnd cell_6t
Xbit_r111_c52 bl[52] br[52] wl[111] vdd gnd cell_6t
Xbit_r112_c52 bl[52] br[52] wl[112] vdd gnd cell_6t
Xbit_r113_c52 bl[52] br[52] wl[113] vdd gnd cell_6t
Xbit_r114_c52 bl[52] br[52] wl[114] vdd gnd cell_6t
Xbit_r115_c52 bl[52] br[52] wl[115] vdd gnd cell_6t
Xbit_r116_c52 bl[52] br[52] wl[116] vdd gnd cell_6t
Xbit_r117_c52 bl[52] br[52] wl[117] vdd gnd cell_6t
Xbit_r118_c52 bl[52] br[52] wl[118] vdd gnd cell_6t
Xbit_r119_c52 bl[52] br[52] wl[119] vdd gnd cell_6t
Xbit_r120_c52 bl[52] br[52] wl[120] vdd gnd cell_6t
Xbit_r121_c52 bl[52] br[52] wl[121] vdd gnd cell_6t
Xbit_r122_c52 bl[52] br[52] wl[122] vdd gnd cell_6t
Xbit_r123_c52 bl[52] br[52] wl[123] vdd gnd cell_6t
Xbit_r124_c52 bl[52] br[52] wl[124] vdd gnd cell_6t
Xbit_r125_c52 bl[52] br[52] wl[125] vdd gnd cell_6t
Xbit_r126_c52 bl[52] br[52] wl[126] vdd gnd cell_6t
Xbit_r127_c52 bl[52] br[52] wl[127] vdd gnd cell_6t
Xbit_r128_c52 bl[52] br[52] wl[128] vdd gnd cell_6t
Xbit_r129_c52 bl[52] br[52] wl[129] vdd gnd cell_6t
Xbit_r130_c52 bl[52] br[52] wl[130] vdd gnd cell_6t
Xbit_r131_c52 bl[52] br[52] wl[131] vdd gnd cell_6t
Xbit_r132_c52 bl[52] br[52] wl[132] vdd gnd cell_6t
Xbit_r133_c52 bl[52] br[52] wl[133] vdd gnd cell_6t
Xbit_r134_c52 bl[52] br[52] wl[134] vdd gnd cell_6t
Xbit_r135_c52 bl[52] br[52] wl[135] vdd gnd cell_6t
Xbit_r136_c52 bl[52] br[52] wl[136] vdd gnd cell_6t
Xbit_r137_c52 bl[52] br[52] wl[137] vdd gnd cell_6t
Xbit_r138_c52 bl[52] br[52] wl[138] vdd gnd cell_6t
Xbit_r139_c52 bl[52] br[52] wl[139] vdd gnd cell_6t
Xbit_r140_c52 bl[52] br[52] wl[140] vdd gnd cell_6t
Xbit_r141_c52 bl[52] br[52] wl[141] vdd gnd cell_6t
Xbit_r142_c52 bl[52] br[52] wl[142] vdd gnd cell_6t
Xbit_r143_c52 bl[52] br[52] wl[143] vdd gnd cell_6t
Xbit_r144_c52 bl[52] br[52] wl[144] vdd gnd cell_6t
Xbit_r145_c52 bl[52] br[52] wl[145] vdd gnd cell_6t
Xbit_r146_c52 bl[52] br[52] wl[146] vdd gnd cell_6t
Xbit_r147_c52 bl[52] br[52] wl[147] vdd gnd cell_6t
Xbit_r148_c52 bl[52] br[52] wl[148] vdd gnd cell_6t
Xbit_r149_c52 bl[52] br[52] wl[149] vdd gnd cell_6t
Xbit_r150_c52 bl[52] br[52] wl[150] vdd gnd cell_6t
Xbit_r151_c52 bl[52] br[52] wl[151] vdd gnd cell_6t
Xbit_r152_c52 bl[52] br[52] wl[152] vdd gnd cell_6t
Xbit_r153_c52 bl[52] br[52] wl[153] vdd gnd cell_6t
Xbit_r154_c52 bl[52] br[52] wl[154] vdd gnd cell_6t
Xbit_r155_c52 bl[52] br[52] wl[155] vdd gnd cell_6t
Xbit_r156_c52 bl[52] br[52] wl[156] vdd gnd cell_6t
Xbit_r157_c52 bl[52] br[52] wl[157] vdd gnd cell_6t
Xbit_r158_c52 bl[52] br[52] wl[158] vdd gnd cell_6t
Xbit_r159_c52 bl[52] br[52] wl[159] vdd gnd cell_6t
Xbit_r160_c52 bl[52] br[52] wl[160] vdd gnd cell_6t
Xbit_r161_c52 bl[52] br[52] wl[161] vdd gnd cell_6t
Xbit_r162_c52 bl[52] br[52] wl[162] vdd gnd cell_6t
Xbit_r163_c52 bl[52] br[52] wl[163] vdd gnd cell_6t
Xbit_r164_c52 bl[52] br[52] wl[164] vdd gnd cell_6t
Xbit_r165_c52 bl[52] br[52] wl[165] vdd gnd cell_6t
Xbit_r166_c52 bl[52] br[52] wl[166] vdd gnd cell_6t
Xbit_r167_c52 bl[52] br[52] wl[167] vdd gnd cell_6t
Xbit_r168_c52 bl[52] br[52] wl[168] vdd gnd cell_6t
Xbit_r169_c52 bl[52] br[52] wl[169] vdd gnd cell_6t
Xbit_r170_c52 bl[52] br[52] wl[170] vdd gnd cell_6t
Xbit_r171_c52 bl[52] br[52] wl[171] vdd gnd cell_6t
Xbit_r172_c52 bl[52] br[52] wl[172] vdd gnd cell_6t
Xbit_r173_c52 bl[52] br[52] wl[173] vdd gnd cell_6t
Xbit_r174_c52 bl[52] br[52] wl[174] vdd gnd cell_6t
Xbit_r175_c52 bl[52] br[52] wl[175] vdd gnd cell_6t
Xbit_r176_c52 bl[52] br[52] wl[176] vdd gnd cell_6t
Xbit_r177_c52 bl[52] br[52] wl[177] vdd gnd cell_6t
Xbit_r178_c52 bl[52] br[52] wl[178] vdd gnd cell_6t
Xbit_r179_c52 bl[52] br[52] wl[179] vdd gnd cell_6t
Xbit_r180_c52 bl[52] br[52] wl[180] vdd gnd cell_6t
Xbit_r181_c52 bl[52] br[52] wl[181] vdd gnd cell_6t
Xbit_r182_c52 bl[52] br[52] wl[182] vdd gnd cell_6t
Xbit_r183_c52 bl[52] br[52] wl[183] vdd gnd cell_6t
Xbit_r184_c52 bl[52] br[52] wl[184] vdd gnd cell_6t
Xbit_r185_c52 bl[52] br[52] wl[185] vdd gnd cell_6t
Xbit_r186_c52 bl[52] br[52] wl[186] vdd gnd cell_6t
Xbit_r187_c52 bl[52] br[52] wl[187] vdd gnd cell_6t
Xbit_r188_c52 bl[52] br[52] wl[188] vdd gnd cell_6t
Xbit_r189_c52 bl[52] br[52] wl[189] vdd gnd cell_6t
Xbit_r190_c52 bl[52] br[52] wl[190] vdd gnd cell_6t
Xbit_r191_c52 bl[52] br[52] wl[191] vdd gnd cell_6t
Xbit_r192_c52 bl[52] br[52] wl[192] vdd gnd cell_6t
Xbit_r193_c52 bl[52] br[52] wl[193] vdd gnd cell_6t
Xbit_r194_c52 bl[52] br[52] wl[194] vdd gnd cell_6t
Xbit_r195_c52 bl[52] br[52] wl[195] vdd gnd cell_6t
Xbit_r196_c52 bl[52] br[52] wl[196] vdd gnd cell_6t
Xbit_r197_c52 bl[52] br[52] wl[197] vdd gnd cell_6t
Xbit_r198_c52 bl[52] br[52] wl[198] vdd gnd cell_6t
Xbit_r199_c52 bl[52] br[52] wl[199] vdd gnd cell_6t
Xbit_r200_c52 bl[52] br[52] wl[200] vdd gnd cell_6t
Xbit_r201_c52 bl[52] br[52] wl[201] vdd gnd cell_6t
Xbit_r202_c52 bl[52] br[52] wl[202] vdd gnd cell_6t
Xbit_r203_c52 bl[52] br[52] wl[203] vdd gnd cell_6t
Xbit_r204_c52 bl[52] br[52] wl[204] vdd gnd cell_6t
Xbit_r205_c52 bl[52] br[52] wl[205] vdd gnd cell_6t
Xbit_r206_c52 bl[52] br[52] wl[206] vdd gnd cell_6t
Xbit_r207_c52 bl[52] br[52] wl[207] vdd gnd cell_6t
Xbit_r208_c52 bl[52] br[52] wl[208] vdd gnd cell_6t
Xbit_r209_c52 bl[52] br[52] wl[209] vdd gnd cell_6t
Xbit_r210_c52 bl[52] br[52] wl[210] vdd gnd cell_6t
Xbit_r211_c52 bl[52] br[52] wl[211] vdd gnd cell_6t
Xbit_r212_c52 bl[52] br[52] wl[212] vdd gnd cell_6t
Xbit_r213_c52 bl[52] br[52] wl[213] vdd gnd cell_6t
Xbit_r214_c52 bl[52] br[52] wl[214] vdd gnd cell_6t
Xbit_r215_c52 bl[52] br[52] wl[215] vdd gnd cell_6t
Xbit_r216_c52 bl[52] br[52] wl[216] vdd gnd cell_6t
Xbit_r217_c52 bl[52] br[52] wl[217] vdd gnd cell_6t
Xbit_r218_c52 bl[52] br[52] wl[218] vdd gnd cell_6t
Xbit_r219_c52 bl[52] br[52] wl[219] vdd gnd cell_6t
Xbit_r220_c52 bl[52] br[52] wl[220] vdd gnd cell_6t
Xbit_r221_c52 bl[52] br[52] wl[221] vdd gnd cell_6t
Xbit_r222_c52 bl[52] br[52] wl[222] vdd gnd cell_6t
Xbit_r223_c52 bl[52] br[52] wl[223] vdd gnd cell_6t
Xbit_r224_c52 bl[52] br[52] wl[224] vdd gnd cell_6t
Xbit_r225_c52 bl[52] br[52] wl[225] vdd gnd cell_6t
Xbit_r226_c52 bl[52] br[52] wl[226] vdd gnd cell_6t
Xbit_r227_c52 bl[52] br[52] wl[227] vdd gnd cell_6t
Xbit_r228_c52 bl[52] br[52] wl[228] vdd gnd cell_6t
Xbit_r229_c52 bl[52] br[52] wl[229] vdd gnd cell_6t
Xbit_r230_c52 bl[52] br[52] wl[230] vdd gnd cell_6t
Xbit_r231_c52 bl[52] br[52] wl[231] vdd gnd cell_6t
Xbit_r232_c52 bl[52] br[52] wl[232] vdd gnd cell_6t
Xbit_r233_c52 bl[52] br[52] wl[233] vdd gnd cell_6t
Xbit_r234_c52 bl[52] br[52] wl[234] vdd gnd cell_6t
Xbit_r235_c52 bl[52] br[52] wl[235] vdd gnd cell_6t
Xbit_r236_c52 bl[52] br[52] wl[236] vdd gnd cell_6t
Xbit_r237_c52 bl[52] br[52] wl[237] vdd gnd cell_6t
Xbit_r238_c52 bl[52] br[52] wl[238] vdd gnd cell_6t
Xbit_r239_c52 bl[52] br[52] wl[239] vdd gnd cell_6t
Xbit_r240_c52 bl[52] br[52] wl[240] vdd gnd cell_6t
Xbit_r241_c52 bl[52] br[52] wl[241] vdd gnd cell_6t
Xbit_r242_c52 bl[52] br[52] wl[242] vdd gnd cell_6t
Xbit_r243_c52 bl[52] br[52] wl[243] vdd gnd cell_6t
Xbit_r244_c52 bl[52] br[52] wl[244] vdd gnd cell_6t
Xbit_r245_c52 bl[52] br[52] wl[245] vdd gnd cell_6t
Xbit_r246_c52 bl[52] br[52] wl[246] vdd gnd cell_6t
Xbit_r247_c52 bl[52] br[52] wl[247] vdd gnd cell_6t
Xbit_r248_c52 bl[52] br[52] wl[248] vdd gnd cell_6t
Xbit_r249_c52 bl[52] br[52] wl[249] vdd gnd cell_6t
Xbit_r250_c52 bl[52] br[52] wl[250] vdd gnd cell_6t
Xbit_r251_c52 bl[52] br[52] wl[251] vdd gnd cell_6t
Xbit_r252_c52 bl[52] br[52] wl[252] vdd gnd cell_6t
Xbit_r253_c52 bl[52] br[52] wl[253] vdd gnd cell_6t
Xbit_r254_c52 bl[52] br[52] wl[254] vdd gnd cell_6t
Xbit_r255_c52 bl[52] br[52] wl[255] vdd gnd cell_6t
Xbit_r0_c53 bl[53] br[53] wl[0] vdd gnd cell_6t
Xbit_r1_c53 bl[53] br[53] wl[1] vdd gnd cell_6t
Xbit_r2_c53 bl[53] br[53] wl[2] vdd gnd cell_6t
Xbit_r3_c53 bl[53] br[53] wl[3] vdd gnd cell_6t
Xbit_r4_c53 bl[53] br[53] wl[4] vdd gnd cell_6t
Xbit_r5_c53 bl[53] br[53] wl[5] vdd gnd cell_6t
Xbit_r6_c53 bl[53] br[53] wl[6] vdd gnd cell_6t
Xbit_r7_c53 bl[53] br[53] wl[7] vdd gnd cell_6t
Xbit_r8_c53 bl[53] br[53] wl[8] vdd gnd cell_6t
Xbit_r9_c53 bl[53] br[53] wl[9] vdd gnd cell_6t
Xbit_r10_c53 bl[53] br[53] wl[10] vdd gnd cell_6t
Xbit_r11_c53 bl[53] br[53] wl[11] vdd gnd cell_6t
Xbit_r12_c53 bl[53] br[53] wl[12] vdd gnd cell_6t
Xbit_r13_c53 bl[53] br[53] wl[13] vdd gnd cell_6t
Xbit_r14_c53 bl[53] br[53] wl[14] vdd gnd cell_6t
Xbit_r15_c53 bl[53] br[53] wl[15] vdd gnd cell_6t
Xbit_r16_c53 bl[53] br[53] wl[16] vdd gnd cell_6t
Xbit_r17_c53 bl[53] br[53] wl[17] vdd gnd cell_6t
Xbit_r18_c53 bl[53] br[53] wl[18] vdd gnd cell_6t
Xbit_r19_c53 bl[53] br[53] wl[19] vdd gnd cell_6t
Xbit_r20_c53 bl[53] br[53] wl[20] vdd gnd cell_6t
Xbit_r21_c53 bl[53] br[53] wl[21] vdd gnd cell_6t
Xbit_r22_c53 bl[53] br[53] wl[22] vdd gnd cell_6t
Xbit_r23_c53 bl[53] br[53] wl[23] vdd gnd cell_6t
Xbit_r24_c53 bl[53] br[53] wl[24] vdd gnd cell_6t
Xbit_r25_c53 bl[53] br[53] wl[25] vdd gnd cell_6t
Xbit_r26_c53 bl[53] br[53] wl[26] vdd gnd cell_6t
Xbit_r27_c53 bl[53] br[53] wl[27] vdd gnd cell_6t
Xbit_r28_c53 bl[53] br[53] wl[28] vdd gnd cell_6t
Xbit_r29_c53 bl[53] br[53] wl[29] vdd gnd cell_6t
Xbit_r30_c53 bl[53] br[53] wl[30] vdd gnd cell_6t
Xbit_r31_c53 bl[53] br[53] wl[31] vdd gnd cell_6t
Xbit_r32_c53 bl[53] br[53] wl[32] vdd gnd cell_6t
Xbit_r33_c53 bl[53] br[53] wl[33] vdd gnd cell_6t
Xbit_r34_c53 bl[53] br[53] wl[34] vdd gnd cell_6t
Xbit_r35_c53 bl[53] br[53] wl[35] vdd gnd cell_6t
Xbit_r36_c53 bl[53] br[53] wl[36] vdd gnd cell_6t
Xbit_r37_c53 bl[53] br[53] wl[37] vdd gnd cell_6t
Xbit_r38_c53 bl[53] br[53] wl[38] vdd gnd cell_6t
Xbit_r39_c53 bl[53] br[53] wl[39] vdd gnd cell_6t
Xbit_r40_c53 bl[53] br[53] wl[40] vdd gnd cell_6t
Xbit_r41_c53 bl[53] br[53] wl[41] vdd gnd cell_6t
Xbit_r42_c53 bl[53] br[53] wl[42] vdd gnd cell_6t
Xbit_r43_c53 bl[53] br[53] wl[43] vdd gnd cell_6t
Xbit_r44_c53 bl[53] br[53] wl[44] vdd gnd cell_6t
Xbit_r45_c53 bl[53] br[53] wl[45] vdd gnd cell_6t
Xbit_r46_c53 bl[53] br[53] wl[46] vdd gnd cell_6t
Xbit_r47_c53 bl[53] br[53] wl[47] vdd gnd cell_6t
Xbit_r48_c53 bl[53] br[53] wl[48] vdd gnd cell_6t
Xbit_r49_c53 bl[53] br[53] wl[49] vdd gnd cell_6t
Xbit_r50_c53 bl[53] br[53] wl[50] vdd gnd cell_6t
Xbit_r51_c53 bl[53] br[53] wl[51] vdd gnd cell_6t
Xbit_r52_c53 bl[53] br[53] wl[52] vdd gnd cell_6t
Xbit_r53_c53 bl[53] br[53] wl[53] vdd gnd cell_6t
Xbit_r54_c53 bl[53] br[53] wl[54] vdd gnd cell_6t
Xbit_r55_c53 bl[53] br[53] wl[55] vdd gnd cell_6t
Xbit_r56_c53 bl[53] br[53] wl[56] vdd gnd cell_6t
Xbit_r57_c53 bl[53] br[53] wl[57] vdd gnd cell_6t
Xbit_r58_c53 bl[53] br[53] wl[58] vdd gnd cell_6t
Xbit_r59_c53 bl[53] br[53] wl[59] vdd gnd cell_6t
Xbit_r60_c53 bl[53] br[53] wl[60] vdd gnd cell_6t
Xbit_r61_c53 bl[53] br[53] wl[61] vdd gnd cell_6t
Xbit_r62_c53 bl[53] br[53] wl[62] vdd gnd cell_6t
Xbit_r63_c53 bl[53] br[53] wl[63] vdd gnd cell_6t
Xbit_r64_c53 bl[53] br[53] wl[64] vdd gnd cell_6t
Xbit_r65_c53 bl[53] br[53] wl[65] vdd gnd cell_6t
Xbit_r66_c53 bl[53] br[53] wl[66] vdd gnd cell_6t
Xbit_r67_c53 bl[53] br[53] wl[67] vdd gnd cell_6t
Xbit_r68_c53 bl[53] br[53] wl[68] vdd gnd cell_6t
Xbit_r69_c53 bl[53] br[53] wl[69] vdd gnd cell_6t
Xbit_r70_c53 bl[53] br[53] wl[70] vdd gnd cell_6t
Xbit_r71_c53 bl[53] br[53] wl[71] vdd gnd cell_6t
Xbit_r72_c53 bl[53] br[53] wl[72] vdd gnd cell_6t
Xbit_r73_c53 bl[53] br[53] wl[73] vdd gnd cell_6t
Xbit_r74_c53 bl[53] br[53] wl[74] vdd gnd cell_6t
Xbit_r75_c53 bl[53] br[53] wl[75] vdd gnd cell_6t
Xbit_r76_c53 bl[53] br[53] wl[76] vdd gnd cell_6t
Xbit_r77_c53 bl[53] br[53] wl[77] vdd gnd cell_6t
Xbit_r78_c53 bl[53] br[53] wl[78] vdd gnd cell_6t
Xbit_r79_c53 bl[53] br[53] wl[79] vdd gnd cell_6t
Xbit_r80_c53 bl[53] br[53] wl[80] vdd gnd cell_6t
Xbit_r81_c53 bl[53] br[53] wl[81] vdd gnd cell_6t
Xbit_r82_c53 bl[53] br[53] wl[82] vdd gnd cell_6t
Xbit_r83_c53 bl[53] br[53] wl[83] vdd gnd cell_6t
Xbit_r84_c53 bl[53] br[53] wl[84] vdd gnd cell_6t
Xbit_r85_c53 bl[53] br[53] wl[85] vdd gnd cell_6t
Xbit_r86_c53 bl[53] br[53] wl[86] vdd gnd cell_6t
Xbit_r87_c53 bl[53] br[53] wl[87] vdd gnd cell_6t
Xbit_r88_c53 bl[53] br[53] wl[88] vdd gnd cell_6t
Xbit_r89_c53 bl[53] br[53] wl[89] vdd gnd cell_6t
Xbit_r90_c53 bl[53] br[53] wl[90] vdd gnd cell_6t
Xbit_r91_c53 bl[53] br[53] wl[91] vdd gnd cell_6t
Xbit_r92_c53 bl[53] br[53] wl[92] vdd gnd cell_6t
Xbit_r93_c53 bl[53] br[53] wl[93] vdd gnd cell_6t
Xbit_r94_c53 bl[53] br[53] wl[94] vdd gnd cell_6t
Xbit_r95_c53 bl[53] br[53] wl[95] vdd gnd cell_6t
Xbit_r96_c53 bl[53] br[53] wl[96] vdd gnd cell_6t
Xbit_r97_c53 bl[53] br[53] wl[97] vdd gnd cell_6t
Xbit_r98_c53 bl[53] br[53] wl[98] vdd gnd cell_6t
Xbit_r99_c53 bl[53] br[53] wl[99] vdd gnd cell_6t
Xbit_r100_c53 bl[53] br[53] wl[100] vdd gnd cell_6t
Xbit_r101_c53 bl[53] br[53] wl[101] vdd gnd cell_6t
Xbit_r102_c53 bl[53] br[53] wl[102] vdd gnd cell_6t
Xbit_r103_c53 bl[53] br[53] wl[103] vdd gnd cell_6t
Xbit_r104_c53 bl[53] br[53] wl[104] vdd gnd cell_6t
Xbit_r105_c53 bl[53] br[53] wl[105] vdd gnd cell_6t
Xbit_r106_c53 bl[53] br[53] wl[106] vdd gnd cell_6t
Xbit_r107_c53 bl[53] br[53] wl[107] vdd gnd cell_6t
Xbit_r108_c53 bl[53] br[53] wl[108] vdd gnd cell_6t
Xbit_r109_c53 bl[53] br[53] wl[109] vdd gnd cell_6t
Xbit_r110_c53 bl[53] br[53] wl[110] vdd gnd cell_6t
Xbit_r111_c53 bl[53] br[53] wl[111] vdd gnd cell_6t
Xbit_r112_c53 bl[53] br[53] wl[112] vdd gnd cell_6t
Xbit_r113_c53 bl[53] br[53] wl[113] vdd gnd cell_6t
Xbit_r114_c53 bl[53] br[53] wl[114] vdd gnd cell_6t
Xbit_r115_c53 bl[53] br[53] wl[115] vdd gnd cell_6t
Xbit_r116_c53 bl[53] br[53] wl[116] vdd gnd cell_6t
Xbit_r117_c53 bl[53] br[53] wl[117] vdd gnd cell_6t
Xbit_r118_c53 bl[53] br[53] wl[118] vdd gnd cell_6t
Xbit_r119_c53 bl[53] br[53] wl[119] vdd gnd cell_6t
Xbit_r120_c53 bl[53] br[53] wl[120] vdd gnd cell_6t
Xbit_r121_c53 bl[53] br[53] wl[121] vdd gnd cell_6t
Xbit_r122_c53 bl[53] br[53] wl[122] vdd gnd cell_6t
Xbit_r123_c53 bl[53] br[53] wl[123] vdd gnd cell_6t
Xbit_r124_c53 bl[53] br[53] wl[124] vdd gnd cell_6t
Xbit_r125_c53 bl[53] br[53] wl[125] vdd gnd cell_6t
Xbit_r126_c53 bl[53] br[53] wl[126] vdd gnd cell_6t
Xbit_r127_c53 bl[53] br[53] wl[127] vdd gnd cell_6t
Xbit_r128_c53 bl[53] br[53] wl[128] vdd gnd cell_6t
Xbit_r129_c53 bl[53] br[53] wl[129] vdd gnd cell_6t
Xbit_r130_c53 bl[53] br[53] wl[130] vdd gnd cell_6t
Xbit_r131_c53 bl[53] br[53] wl[131] vdd gnd cell_6t
Xbit_r132_c53 bl[53] br[53] wl[132] vdd gnd cell_6t
Xbit_r133_c53 bl[53] br[53] wl[133] vdd gnd cell_6t
Xbit_r134_c53 bl[53] br[53] wl[134] vdd gnd cell_6t
Xbit_r135_c53 bl[53] br[53] wl[135] vdd gnd cell_6t
Xbit_r136_c53 bl[53] br[53] wl[136] vdd gnd cell_6t
Xbit_r137_c53 bl[53] br[53] wl[137] vdd gnd cell_6t
Xbit_r138_c53 bl[53] br[53] wl[138] vdd gnd cell_6t
Xbit_r139_c53 bl[53] br[53] wl[139] vdd gnd cell_6t
Xbit_r140_c53 bl[53] br[53] wl[140] vdd gnd cell_6t
Xbit_r141_c53 bl[53] br[53] wl[141] vdd gnd cell_6t
Xbit_r142_c53 bl[53] br[53] wl[142] vdd gnd cell_6t
Xbit_r143_c53 bl[53] br[53] wl[143] vdd gnd cell_6t
Xbit_r144_c53 bl[53] br[53] wl[144] vdd gnd cell_6t
Xbit_r145_c53 bl[53] br[53] wl[145] vdd gnd cell_6t
Xbit_r146_c53 bl[53] br[53] wl[146] vdd gnd cell_6t
Xbit_r147_c53 bl[53] br[53] wl[147] vdd gnd cell_6t
Xbit_r148_c53 bl[53] br[53] wl[148] vdd gnd cell_6t
Xbit_r149_c53 bl[53] br[53] wl[149] vdd gnd cell_6t
Xbit_r150_c53 bl[53] br[53] wl[150] vdd gnd cell_6t
Xbit_r151_c53 bl[53] br[53] wl[151] vdd gnd cell_6t
Xbit_r152_c53 bl[53] br[53] wl[152] vdd gnd cell_6t
Xbit_r153_c53 bl[53] br[53] wl[153] vdd gnd cell_6t
Xbit_r154_c53 bl[53] br[53] wl[154] vdd gnd cell_6t
Xbit_r155_c53 bl[53] br[53] wl[155] vdd gnd cell_6t
Xbit_r156_c53 bl[53] br[53] wl[156] vdd gnd cell_6t
Xbit_r157_c53 bl[53] br[53] wl[157] vdd gnd cell_6t
Xbit_r158_c53 bl[53] br[53] wl[158] vdd gnd cell_6t
Xbit_r159_c53 bl[53] br[53] wl[159] vdd gnd cell_6t
Xbit_r160_c53 bl[53] br[53] wl[160] vdd gnd cell_6t
Xbit_r161_c53 bl[53] br[53] wl[161] vdd gnd cell_6t
Xbit_r162_c53 bl[53] br[53] wl[162] vdd gnd cell_6t
Xbit_r163_c53 bl[53] br[53] wl[163] vdd gnd cell_6t
Xbit_r164_c53 bl[53] br[53] wl[164] vdd gnd cell_6t
Xbit_r165_c53 bl[53] br[53] wl[165] vdd gnd cell_6t
Xbit_r166_c53 bl[53] br[53] wl[166] vdd gnd cell_6t
Xbit_r167_c53 bl[53] br[53] wl[167] vdd gnd cell_6t
Xbit_r168_c53 bl[53] br[53] wl[168] vdd gnd cell_6t
Xbit_r169_c53 bl[53] br[53] wl[169] vdd gnd cell_6t
Xbit_r170_c53 bl[53] br[53] wl[170] vdd gnd cell_6t
Xbit_r171_c53 bl[53] br[53] wl[171] vdd gnd cell_6t
Xbit_r172_c53 bl[53] br[53] wl[172] vdd gnd cell_6t
Xbit_r173_c53 bl[53] br[53] wl[173] vdd gnd cell_6t
Xbit_r174_c53 bl[53] br[53] wl[174] vdd gnd cell_6t
Xbit_r175_c53 bl[53] br[53] wl[175] vdd gnd cell_6t
Xbit_r176_c53 bl[53] br[53] wl[176] vdd gnd cell_6t
Xbit_r177_c53 bl[53] br[53] wl[177] vdd gnd cell_6t
Xbit_r178_c53 bl[53] br[53] wl[178] vdd gnd cell_6t
Xbit_r179_c53 bl[53] br[53] wl[179] vdd gnd cell_6t
Xbit_r180_c53 bl[53] br[53] wl[180] vdd gnd cell_6t
Xbit_r181_c53 bl[53] br[53] wl[181] vdd gnd cell_6t
Xbit_r182_c53 bl[53] br[53] wl[182] vdd gnd cell_6t
Xbit_r183_c53 bl[53] br[53] wl[183] vdd gnd cell_6t
Xbit_r184_c53 bl[53] br[53] wl[184] vdd gnd cell_6t
Xbit_r185_c53 bl[53] br[53] wl[185] vdd gnd cell_6t
Xbit_r186_c53 bl[53] br[53] wl[186] vdd gnd cell_6t
Xbit_r187_c53 bl[53] br[53] wl[187] vdd gnd cell_6t
Xbit_r188_c53 bl[53] br[53] wl[188] vdd gnd cell_6t
Xbit_r189_c53 bl[53] br[53] wl[189] vdd gnd cell_6t
Xbit_r190_c53 bl[53] br[53] wl[190] vdd gnd cell_6t
Xbit_r191_c53 bl[53] br[53] wl[191] vdd gnd cell_6t
Xbit_r192_c53 bl[53] br[53] wl[192] vdd gnd cell_6t
Xbit_r193_c53 bl[53] br[53] wl[193] vdd gnd cell_6t
Xbit_r194_c53 bl[53] br[53] wl[194] vdd gnd cell_6t
Xbit_r195_c53 bl[53] br[53] wl[195] vdd gnd cell_6t
Xbit_r196_c53 bl[53] br[53] wl[196] vdd gnd cell_6t
Xbit_r197_c53 bl[53] br[53] wl[197] vdd gnd cell_6t
Xbit_r198_c53 bl[53] br[53] wl[198] vdd gnd cell_6t
Xbit_r199_c53 bl[53] br[53] wl[199] vdd gnd cell_6t
Xbit_r200_c53 bl[53] br[53] wl[200] vdd gnd cell_6t
Xbit_r201_c53 bl[53] br[53] wl[201] vdd gnd cell_6t
Xbit_r202_c53 bl[53] br[53] wl[202] vdd gnd cell_6t
Xbit_r203_c53 bl[53] br[53] wl[203] vdd gnd cell_6t
Xbit_r204_c53 bl[53] br[53] wl[204] vdd gnd cell_6t
Xbit_r205_c53 bl[53] br[53] wl[205] vdd gnd cell_6t
Xbit_r206_c53 bl[53] br[53] wl[206] vdd gnd cell_6t
Xbit_r207_c53 bl[53] br[53] wl[207] vdd gnd cell_6t
Xbit_r208_c53 bl[53] br[53] wl[208] vdd gnd cell_6t
Xbit_r209_c53 bl[53] br[53] wl[209] vdd gnd cell_6t
Xbit_r210_c53 bl[53] br[53] wl[210] vdd gnd cell_6t
Xbit_r211_c53 bl[53] br[53] wl[211] vdd gnd cell_6t
Xbit_r212_c53 bl[53] br[53] wl[212] vdd gnd cell_6t
Xbit_r213_c53 bl[53] br[53] wl[213] vdd gnd cell_6t
Xbit_r214_c53 bl[53] br[53] wl[214] vdd gnd cell_6t
Xbit_r215_c53 bl[53] br[53] wl[215] vdd gnd cell_6t
Xbit_r216_c53 bl[53] br[53] wl[216] vdd gnd cell_6t
Xbit_r217_c53 bl[53] br[53] wl[217] vdd gnd cell_6t
Xbit_r218_c53 bl[53] br[53] wl[218] vdd gnd cell_6t
Xbit_r219_c53 bl[53] br[53] wl[219] vdd gnd cell_6t
Xbit_r220_c53 bl[53] br[53] wl[220] vdd gnd cell_6t
Xbit_r221_c53 bl[53] br[53] wl[221] vdd gnd cell_6t
Xbit_r222_c53 bl[53] br[53] wl[222] vdd gnd cell_6t
Xbit_r223_c53 bl[53] br[53] wl[223] vdd gnd cell_6t
Xbit_r224_c53 bl[53] br[53] wl[224] vdd gnd cell_6t
Xbit_r225_c53 bl[53] br[53] wl[225] vdd gnd cell_6t
Xbit_r226_c53 bl[53] br[53] wl[226] vdd gnd cell_6t
Xbit_r227_c53 bl[53] br[53] wl[227] vdd gnd cell_6t
Xbit_r228_c53 bl[53] br[53] wl[228] vdd gnd cell_6t
Xbit_r229_c53 bl[53] br[53] wl[229] vdd gnd cell_6t
Xbit_r230_c53 bl[53] br[53] wl[230] vdd gnd cell_6t
Xbit_r231_c53 bl[53] br[53] wl[231] vdd gnd cell_6t
Xbit_r232_c53 bl[53] br[53] wl[232] vdd gnd cell_6t
Xbit_r233_c53 bl[53] br[53] wl[233] vdd gnd cell_6t
Xbit_r234_c53 bl[53] br[53] wl[234] vdd gnd cell_6t
Xbit_r235_c53 bl[53] br[53] wl[235] vdd gnd cell_6t
Xbit_r236_c53 bl[53] br[53] wl[236] vdd gnd cell_6t
Xbit_r237_c53 bl[53] br[53] wl[237] vdd gnd cell_6t
Xbit_r238_c53 bl[53] br[53] wl[238] vdd gnd cell_6t
Xbit_r239_c53 bl[53] br[53] wl[239] vdd gnd cell_6t
Xbit_r240_c53 bl[53] br[53] wl[240] vdd gnd cell_6t
Xbit_r241_c53 bl[53] br[53] wl[241] vdd gnd cell_6t
Xbit_r242_c53 bl[53] br[53] wl[242] vdd gnd cell_6t
Xbit_r243_c53 bl[53] br[53] wl[243] vdd gnd cell_6t
Xbit_r244_c53 bl[53] br[53] wl[244] vdd gnd cell_6t
Xbit_r245_c53 bl[53] br[53] wl[245] vdd gnd cell_6t
Xbit_r246_c53 bl[53] br[53] wl[246] vdd gnd cell_6t
Xbit_r247_c53 bl[53] br[53] wl[247] vdd gnd cell_6t
Xbit_r248_c53 bl[53] br[53] wl[248] vdd gnd cell_6t
Xbit_r249_c53 bl[53] br[53] wl[249] vdd gnd cell_6t
Xbit_r250_c53 bl[53] br[53] wl[250] vdd gnd cell_6t
Xbit_r251_c53 bl[53] br[53] wl[251] vdd gnd cell_6t
Xbit_r252_c53 bl[53] br[53] wl[252] vdd gnd cell_6t
Xbit_r253_c53 bl[53] br[53] wl[253] vdd gnd cell_6t
Xbit_r254_c53 bl[53] br[53] wl[254] vdd gnd cell_6t
Xbit_r255_c53 bl[53] br[53] wl[255] vdd gnd cell_6t
Xbit_r0_c54 bl[54] br[54] wl[0] vdd gnd cell_6t
Xbit_r1_c54 bl[54] br[54] wl[1] vdd gnd cell_6t
Xbit_r2_c54 bl[54] br[54] wl[2] vdd gnd cell_6t
Xbit_r3_c54 bl[54] br[54] wl[3] vdd gnd cell_6t
Xbit_r4_c54 bl[54] br[54] wl[4] vdd gnd cell_6t
Xbit_r5_c54 bl[54] br[54] wl[5] vdd gnd cell_6t
Xbit_r6_c54 bl[54] br[54] wl[6] vdd gnd cell_6t
Xbit_r7_c54 bl[54] br[54] wl[7] vdd gnd cell_6t
Xbit_r8_c54 bl[54] br[54] wl[8] vdd gnd cell_6t
Xbit_r9_c54 bl[54] br[54] wl[9] vdd gnd cell_6t
Xbit_r10_c54 bl[54] br[54] wl[10] vdd gnd cell_6t
Xbit_r11_c54 bl[54] br[54] wl[11] vdd gnd cell_6t
Xbit_r12_c54 bl[54] br[54] wl[12] vdd gnd cell_6t
Xbit_r13_c54 bl[54] br[54] wl[13] vdd gnd cell_6t
Xbit_r14_c54 bl[54] br[54] wl[14] vdd gnd cell_6t
Xbit_r15_c54 bl[54] br[54] wl[15] vdd gnd cell_6t
Xbit_r16_c54 bl[54] br[54] wl[16] vdd gnd cell_6t
Xbit_r17_c54 bl[54] br[54] wl[17] vdd gnd cell_6t
Xbit_r18_c54 bl[54] br[54] wl[18] vdd gnd cell_6t
Xbit_r19_c54 bl[54] br[54] wl[19] vdd gnd cell_6t
Xbit_r20_c54 bl[54] br[54] wl[20] vdd gnd cell_6t
Xbit_r21_c54 bl[54] br[54] wl[21] vdd gnd cell_6t
Xbit_r22_c54 bl[54] br[54] wl[22] vdd gnd cell_6t
Xbit_r23_c54 bl[54] br[54] wl[23] vdd gnd cell_6t
Xbit_r24_c54 bl[54] br[54] wl[24] vdd gnd cell_6t
Xbit_r25_c54 bl[54] br[54] wl[25] vdd gnd cell_6t
Xbit_r26_c54 bl[54] br[54] wl[26] vdd gnd cell_6t
Xbit_r27_c54 bl[54] br[54] wl[27] vdd gnd cell_6t
Xbit_r28_c54 bl[54] br[54] wl[28] vdd gnd cell_6t
Xbit_r29_c54 bl[54] br[54] wl[29] vdd gnd cell_6t
Xbit_r30_c54 bl[54] br[54] wl[30] vdd gnd cell_6t
Xbit_r31_c54 bl[54] br[54] wl[31] vdd gnd cell_6t
Xbit_r32_c54 bl[54] br[54] wl[32] vdd gnd cell_6t
Xbit_r33_c54 bl[54] br[54] wl[33] vdd gnd cell_6t
Xbit_r34_c54 bl[54] br[54] wl[34] vdd gnd cell_6t
Xbit_r35_c54 bl[54] br[54] wl[35] vdd gnd cell_6t
Xbit_r36_c54 bl[54] br[54] wl[36] vdd gnd cell_6t
Xbit_r37_c54 bl[54] br[54] wl[37] vdd gnd cell_6t
Xbit_r38_c54 bl[54] br[54] wl[38] vdd gnd cell_6t
Xbit_r39_c54 bl[54] br[54] wl[39] vdd gnd cell_6t
Xbit_r40_c54 bl[54] br[54] wl[40] vdd gnd cell_6t
Xbit_r41_c54 bl[54] br[54] wl[41] vdd gnd cell_6t
Xbit_r42_c54 bl[54] br[54] wl[42] vdd gnd cell_6t
Xbit_r43_c54 bl[54] br[54] wl[43] vdd gnd cell_6t
Xbit_r44_c54 bl[54] br[54] wl[44] vdd gnd cell_6t
Xbit_r45_c54 bl[54] br[54] wl[45] vdd gnd cell_6t
Xbit_r46_c54 bl[54] br[54] wl[46] vdd gnd cell_6t
Xbit_r47_c54 bl[54] br[54] wl[47] vdd gnd cell_6t
Xbit_r48_c54 bl[54] br[54] wl[48] vdd gnd cell_6t
Xbit_r49_c54 bl[54] br[54] wl[49] vdd gnd cell_6t
Xbit_r50_c54 bl[54] br[54] wl[50] vdd gnd cell_6t
Xbit_r51_c54 bl[54] br[54] wl[51] vdd gnd cell_6t
Xbit_r52_c54 bl[54] br[54] wl[52] vdd gnd cell_6t
Xbit_r53_c54 bl[54] br[54] wl[53] vdd gnd cell_6t
Xbit_r54_c54 bl[54] br[54] wl[54] vdd gnd cell_6t
Xbit_r55_c54 bl[54] br[54] wl[55] vdd gnd cell_6t
Xbit_r56_c54 bl[54] br[54] wl[56] vdd gnd cell_6t
Xbit_r57_c54 bl[54] br[54] wl[57] vdd gnd cell_6t
Xbit_r58_c54 bl[54] br[54] wl[58] vdd gnd cell_6t
Xbit_r59_c54 bl[54] br[54] wl[59] vdd gnd cell_6t
Xbit_r60_c54 bl[54] br[54] wl[60] vdd gnd cell_6t
Xbit_r61_c54 bl[54] br[54] wl[61] vdd gnd cell_6t
Xbit_r62_c54 bl[54] br[54] wl[62] vdd gnd cell_6t
Xbit_r63_c54 bl[54] br[54] wl[63] vdd gnd cell_6t
Xbit_r64_c54 bl[54] br[54] wl[64] vdd gnd cell_6t
Xbit_r65_c54 bl[54] br[54] wl[65] vdd gnd cell_6t
Xbit_r66_c54 bl[54] br[54] wl[66] vdd gnd cell_6t
Xbit_r67_c54 bl[54] br[54] wl[67] vdd gnd cell_6t
Xbit_r68_c54 bl[54] br[54] wl[68] vdd gnd cell_6t
Xbit_r69_c54 bl[54] br[54] wl[69] vdd gnd cell_6t
Xbit_r70_c54 bl[54] br[54] wl[70] vdd gnd cell_6t
Xbit_r71_c54 bl[54] br[54] wl[71] vdd gnd cell_6t
Xbit_r72_c54 bl[54] br[54] wl[72] vdd gnd cell_6t
Xbit_r73_c54 bl[54] br[54] wl[73] vdd gnd cell_6t
Xbit_r74_c54 bl[54] br[54] wl[74] vdd gnd cell_6t
Xbit_r75_c54 bl[54] br[54] wl[75] vdd gnd cell_6t
Xbit_r76_c54 bl[54] br[54] wl[76] vdd gnd cell_6t
Xbit_r77_c54 bl[54] br[54] wl[77] vdd gnd cell_6t
Xbit_r78_c54 bl[54] br[54] wl[78] vdd gnd cell_6t
Xbit_r79_c54 bl[54] br[54] wl[79] vdd gnd cell_6t
Xbit_r80_c54 bl[54] br[54] wl[80] vdd gnd cell_6t
Xbit_r81_c54 bl[54] br[54] wl[81] vdd gnd cell_6t
Xbit_r82_c54 bl[54] br[54] wl[82] vdd gnd cell_6t
Xbit_r83_c54 bl[54] br[54] wl[83] vdd gnd cell_6t
Xbit_r84_c54 bl[54] br[54] wl[84] vdd gnd cell_6t
Xbit_r85_c54 bl[54] br[54] wl[85] vdd gnd cell_6t
Xbit_r86_c54 bl[54] br[54] wl[86] vdd gnd cell_6t
Xbit_r87_c54 bl[54] br[54] wl[87] vdd gnd cell_6t
Xbit_r88_c54 bl[54] br[54] wl[88] vdd gnd cell_6t
Xbit_r89_c54 bl[54] br[54] wl[89] vdd gnd cell_6t
Xbit_r90_c54 bl[54] br[54] wl[90] vdd gnd cell_6t
Xbit_r91_c54 bl[54] br[54] wl[91] vdd gnd cell_6t
Xbit_r92_c54 bl[54] br[54] wl[92] vdd gnd cell_6t
Xbit_r93_c54 bl[54] br[54] wl[93] vdd gnd cell_6t
Xbit_r94_c54 bl[54] br[54] wl[94] vdd gnd cell_6t
Xbit_r95_c54 bl[54] br[54] wl[95] vdd gnd cell_6t
Xbit_r96_c54 bl[54] br[54] wl[96] vdd gnd cell_6t
Xbit_r97_c54 bl[54] br[54] wl[97] vdd gnd cell_6t
Xbit_r98_c54 bl[54] br[54] wl[98] vdd gnd cell_6t
Xbit_r99_c54 bl[54] br[54] wl[99] vdd gnd cell_6t
Xbit_r100_c54 bl[54] br[54] wl[100] vdd gnd cell_6t
Xbit_r101_c54 bl[54] br[54] wl[101] vdd gnd cell_6t
Xbit_r102_c54 bl[54] br[54] wl[102] vdd gnd cell_6t
Xbit_r103_c54 bl[54] br[54] wl[103] vdd gnd cell_6t
Xbit_r104_c54 bl[54] br[54] wl[104] vdd gnd cell_6t
Xbit_r105_c54 bl[54] br[54] wl[105] vdd gnd cell_6t
Xbit_r106_c54 bl[54] br[54] wl[106] vdd gnd cell_6t
Xbit_r107_c54 bl[54] br[54] wl[107] vdd gnd cell_6t
Xbit_r108_c54 bl[54] br[54] wl[108] vdd gnd cell_6t
Xbit_r109_c54 bl[54] br[54] wl[109] vdd gnd cell_6t
Xbit_r110_c54 bl[54] br[54] wl[110] vdd gnd cell_6t
Xbit_r111_c54 bl[54] br[54] wl[111] vdd gnd cell_6t
Xbit_r112_c54 bl[54] br[54] wl[112] vdd gnd cell_6t
Xbit_r113_c54 bl[54] br[54] wl[113] vdd gnd cell_6t
Xbit_r114_c54 bl[54] br[54] wl[114] vdd gnd cell_6t
Xbit_r115_c54 bl[54] br[54] wl[115] vdd gnd cell_6t
Xbit_r116_c54 bl[54] br[54] wl[116] vdd gnd cell_6t
Xbit_r117_c54 bl[54] br[54] wl[117] vdd gnd cell_6t
Xbit_r118_c54 bl[54] br[54] wl[118] vdd gnd cell_6t
Xbit_r119_c54 bl[54] br[54] wl[119] vdd gnd cell_6t
Xbit_r120_c54 bl[54] br[54] wl[120] vdd gnd cell_6t
Xbit_r121_c54 bl[54] br[54] wl[121] vdd gnd cell_6t
Xbit_r122_c54 bl[54] br[54] wl[122] vdd gnd cell_6t
Xbit_r123_c54 bl[54] br[54] wl[123] vdd gnd cell_6t
Xbit_r124_c54 bl[54] br[54] wl[124] vdd gnd cell_6t
Xbit_r125_c54 bl[54] br[54] wl[125] vdd gnd cell_6t
Xbit_r126_c54 bl[54] br[54] wl[126] vdd gnd cell_6t
Xbit_r127_c54 bl[54] br[54] wl[127] vdd gnd cell_6t
Xbit_r128_c54 bl[54] br[54] wl[128] vdd gnd cell_6t
Xbit_r129_c54 bl[54] br[54] wl[129] vdd gnd cell_6t
Xbit_r130_c54 bl[54] br[54] wl[130] vdd gnd cell_6t
Xbit_r131_c54 bl[54] br[54] wl[131] vdd gnd cell_6t
Xbit_r132_c54 bl[54] br[54] wl[132] vdd gnd cell_6t
Xbit_r133_c54 bl[54] br[54] wl[133] vdd gnd cell_6t
Xbit_r134_c54 bl[54] br[54] wl[134] vdd gnd cell_6t
Xbit_r135_c54 bl[54] br[54] wl[135] vdd gnd cell_6t
Xbit_r136_c54 bl[54] br[54] wl[136] vdd gnd cell_6t
Xbit_r137_c54 bl[54] br[54] wl[137] vdd gnd cell_6t
Xbit_r138_c54 bl[54] br[54] wl[138] vdd gnd cell_6t
Xbit_r139_c54 bl[54] br[54] wl[139] vdd gnd cell_6t
Xbit_r140_c54 bl[54] br[54] wl[140] vdd gnd cell_6t
Xbit_r141_c54 bl[54] br[54] wl[141] vdd gnd cell_6t
Xbit_r142_c54 bl[54] br[54] wl[142] vdd gnd cell_6t
Xbit_r143_c54 bl[54] br[54] wl[143] vdd gnd cell_6t
Xbit_r144_c54 bl[54] br[54] wl[144] vdd gnd cell_6t
Xbit_r145_c54 bl[54] br[54] wl[145] vdd gnd cell_6t
Xbit_r146_c54 bl[54] br[54] wl[146] vdd gnd cell_6t
Xbit_r147_c54 bl[54] br[54] wl[147] vdd gnd cell_6t
Xbit_r148_c54 bl[54] br[54] wl[148] vdd gnd cell_6t
Xbit_r149_c54 bl[54] br[54] wl[149] vdd gnd cell_6t
Xbit_r150_c54 bl[54] br[54] wl[150] vdd gnd cell_6t
Xbit_r151_c54 bl[54] br[54] wl[151] vdd gnd cell_6t
Xbit_r152_c54 bl[54] br[54] wl[152] vdd gnd cell_6t
Xbit_r153_c54 bl[54] br[54] wl[153] vdd gnd cell_6t
Xbit_r154_c54 bl[54] br[54] wl[154] vdd gnd cell_6t
Xbit_r155_c54 bl[54] br[54] wl[155] vdd gnd cell_6t
Xbit_r156_c54 bl[54] br[54] wl[156] vdd gnd cell_6t
Xbit_r157_c54 bl[54] br[54] wl[157] vdd gnd cell_6t
Xbit_r158_c54 bl[54] br[54] wl[158] vdd gnd cell_6t
Xbit_r159_c54 bl[54] br[54] wl[159] vdd gnd cell_6t
Xbit_r160_c54 bl[54] br[54] wl[160] vdd gnd cell_6t
Xbit_r161_c54 bl[54] br[54] wl[161] vdd gnd cell_6t
Xbit_r162_c54 bl[54] br[54] wl[162] vdd gnd cell_6t
Xbit_r163_c54 bl[54] br[54] wl[163] vdd gnd cell_6t
Xbit_r164_c54 bl[54] br[54] wl[164] vdd gnd cell_6t
Xbit_r165_c54 bl[54] br[54] wl[165] vdd gnd cell_6t
Xbit_r166_c54 bl[54] br[54] wl[166] vdd gnd cell_6t
Xbit_r167_c54 bl[54] br[54] wl[167] vdd gnd cell_6t
Xbit_r168_c54 bl[54] br[54] wl[168] vdd gnd cell_6t
Xbit_r169_c54 bl[54] br[54] wl[169] vdd gnd cell_6t
Xbit_r170_c54 bl[54] br[54] wl[170] vdd gnd cell_6t
Xbit_r171_c54 bl[54] br[54] wl[171] vdd gnd cell_6t
Xbit_r172_c54 bl[54] br[54] wl[172] vdd gnd cell_6t
Xbit_r173_c54 bl[54] br[54] wl[173] vdd gnd cell_6t
Xbit_r174_c54 bl[54] br[54] wl[174] vdd gnd cell_6t
Xbit_r175_c54 bl[54] br[54] wl[175] vdd gnd cell_6t
Xbit_r176_c54 bl[54] br[54] wl[176] vdd gnd cell_6t
Xbit_r177_c54 bl[54] br[54] wl[177] vdd gnd cell_6t
Xbit_r178_c54 bl[54] br[54] wl[178] vdd gnd cell_6t
Xbit_r179_c54 bl[54] br[54] wl[179] vdd gnd cell_6t
Xbit_r180_c54 bl[54] br[54] wl[180] vdd gnd cell_6t
Xbit_r181_c54 bl[54] br[54] wl[181] vdd gnd cell_6t
Xbit_r182_c54 bl[54] br[54] wl[182] vdd gnd cell_6t
Xbit_r183_c54 bl[54] br[54] wl[183] vdd gnd cell_6t
Xbit_r184_c54 bl[54] br[54] wl[184] vdd gnd cell_6t
Xbit_r185_c54 bl[54] br[54] wl[185] vdd gnd cell_6t
Xbit_r186_c54 bl[54] br[54] wl[186] vdd gnd cell_6t
Xbit_r187_c54 bl[54] br[54] wl[187] vdd gnd cell_6t
Xbit_r188_c54 bl[54] br[54] wl[188] vdd gnd cell_6t
Xbit_r189_c54 bl[54] br[54] wl[189] vdd gnd cell_6t
Xbit_r190_c54 bl[54] br[54] wl[190] vdd gnd cell_6t
Xbit_r191_c54 bl[54] br[54] wl[191] vdd gnd cell_6t
Xbit_r192_c54 bl[54] br[54] wl[192] vdd gnd cell_6t
Xbit_r193_c54 bl[54] br[54] wl[193] vdd gnd cell_6t
Xbit_r194_c54 bl[54] br[54] wl[194] vdd gnd cell_6t
Xbit_r195_c54 bl[54] br[54] wl[195] vdd gnd cell_6t
Xbit_r196_c54 bl[54] br[54] wl[196] vdd gnd cell_6t
Xbit_r197_c54 bl[54] br[54] wl[197] vdd gnd cell_6t
Xbit_r198_c54 bl[54] br[54] wl[198] vdd gnd cell_6t
Xbit_r199_c54 bl[54] br[54] wl[199] vdd gnd cell_6t
Xbit_r200_c54 bl[54] br[54] wl[200] vdd gnd cell_6t
Xbit_r201_c54 bl[54] br[54] wl[201] vdd gnd cell_6t
Xbit_r202_c54 bl[54] br[54] wl[202] vdd gnd cell_6t
Xbit_r203_c54 bl[54] br[54] wl[203] vdd gnd cell_6t
Xbit_r204_c54 bl[54] br[54] wl[204] vdd gnd cell_6t
Xbit_r205_c54 bl[54] br[54] wl[205] vdd gnd cell_6t
Xbit_r206_c54 bl[54] br[54] wl[206] vdd gnd cell_6t
Xbit_r207_c54 bl[54] br[54] wl[207] vdd gnd cell_6t
Xbit_r208_c54 bl[54] br[54] wl[208] vdd gnd cell_6t
Xbit_r209_c54 bl[54] br[54] wl[209] vdd gnd cell_6t
Xbit_r210_c54 bl[54] br[54] wl[210] vdd gnd cell_6t
Xbit_r211_c54 bl[54] br[54] wl[211] vdd gnd cell_6t
Xbit_r212_c54 bl[54] br[54] wl[212] vdd gnd cell_6t
Xbit_r213_c54 bl[54] br[54] wl[213] vdd gnd cell_6t
Xbit_r214_c54 bl[54] br[54] wl[214] vdd gnd cell_6t
Xbit_r215_c54 bl[54] br[54] wl[215] vdd gnd cell_6t
Xbit_r216_c54 bl[54] br[54] wl[216] vdd gnd cell_6t
Xbit_r217_c54 bl[54] br[54] wl[217] vdd gnd cell_6t
Xbit_r218_c54 bl[54] br[54] wl[218] vdd gnd cell_6t
Xbit_r219_c54 bl[54] br[54] wl[219] vdd gnd cell_6t
Xbit_r220_c54 bl[54] br[54] wl[220] vdd gnd cell_6t
Xbit_r221_c54 bl[54] br[54] wl[221] vdd gnd cell_6t
Xbit_r222_c54 bl[54] br[54] wl[222] vdd gnd cell_6t
Xbit_r223_c54 bl[54] br[54] wl[223] vdd gnd cell_6t
Xbit_r224_c54 bl[54] br[54] wl[224] vdd gnd cell_6t
Xbit_r225_c54 bl[54] br[54] wl[225] vdd gnd cell_6t
Xbit_r226_c54 bl[54] br[54] wl[226] vdd gnd cell_6t
Xbit_r227_c54 bl[54] br[54] wl[227] vdd gnd cell_6t
Xbit_r228_c54 bl[54] br[54] wl[228] vdd gnd cell_6t
Xbit_r229_c54 bl[54] br[54] wl[229] vdd gnd cell_6t
Xbit_r230_c54 bl[54] br[54] wl[230] vdd gnd cell_6t
Xbit_r231_c54 bl[54] br[54] wl[231] vdd gnd cell_6t
Xbit_r232_c54 bl[54] br[54] wl[232] vdd gnd cell_6t
Xbit_r233_c54 bl[54] br[54] wl[233] vdd gnd cell_6t
Xbit_r234_c54 bl[54] br[54] wl[234] vdd gnd cell_6t
Xbit_r235_c54 bl[54] br[54] wl[235] vdd gnd cell_6t
Xbit_r236_c54 bl[54] br[54] wl[236] vdd gnd cell_6t
Xbit_r237_c54 bl[54] br[54] wl[237] vdd gnd cell_6t
Xbit_r238_c54 bl[54] br[54] wl[238] vdd gnd cell_6t
Xbit_r239_c54 bl[54] br[54] wl[239] vdd gnd cell_6t
Xbit_r240_c54 bl[54] br[54] wl[240] vdd gnd cell_6t
Xbit_r241_c54 bl[54] br[54] wl[241] vdd gnd cell_6t
Xbit_r242_c54 bl[54] br[54] wl[242] vdd gnd cell_6t
Xbit_r243_c54 bl[54] br[54] wl[243] vdd gnd cell_6t
Xbit_r244_c54 bl[54] br[54] wl[244] vdd gnd cell_6t
Xbit_r245_c54 bl[54] br[54] wl[245] vdd gnd cell_6t
Xbit_r246_c54 bl[54] br[54] wl[246] vdd gnd cell_6t
Xbit_r247_c54 bl[54] br[54] wl[247] vdd gnd cell_6t
Xbit_r248_c54 bl[54] br[54] wl[248] vdd gnd cell_6t
Xbit_r249_c54 bl[54] br[54] wl[249] vdd gnd cell_6t
Xbit_r250_c54 bl[54] br[54] wl[250] vdd gnd cell_6t
Xbit_r251_c54 bl[54] br[54] wl[251] vdd gnd cell_6t
Xbit_r252_c54 bl[54] br[54] wl[252] vdd gnd cell_6t
Xbit_r253_c54 bl[54] br[54] wl[253] vdd gnd cell_6t
Xbit_r254_c54 bl[54] br[54] wl[254] vdd gnd cell_6t
Xbit_r255_c54 bl[54] br[54] wl[255] vdd gnd cell_6t
Xbit_r0_c55 bl[55] br[55] wl[0] vdd gnd cell_6t
Xbit_r1_c55 bl[55] br[55] wl[1] vdd gnd cell_6t
Xbit_r2_c55 bl[55] br[55] wl[2] vdd gnd cell_6t
Xbit_r3_c55 bl[55] br[55] wl[3] vdd gnd cell_6t
Xbit_r4_c55 bl[55] br[55] wl[4] vdd gnd cell_6t
Xbit_r5_c55 bl[55] br[55] wl[5] vdd gnd cell_6t
Xbit_r6_c55 bl[55] br[55] wl[6] vdd gnd cell_6t
Xbit_r7_c55 bl[55] br[55] wl[7] vdd gnd cell_6t
Xbit_r8_c55 bl[55] br[55] wl[8] vdd gnd cell_6t
Xbit_r9_c55 bl[55] br[55] wl[9] vdd gnd cell_6t
Xbit_r10_c55 bl[55] br[55] wl[10] vdd gnd cell_6t
Xbit_r11_c55 bl[55] br[55] wl[11] vdd gnd cell_6t
Xbit_r12_c55 bl[55] br[55] wl[12] vdd gnd cell_6t
Xbit_r13_c55 bl[55] br[55] wl[13] vdd gnd cell_6t
Xbit_r14_c55 bl[55] br[55] wl[14] vdd gnd cell_6t
Xbit_r15_c55 bl[55] br[55] wl[15] vdd gnd cell_6t
Xbit_r16_c55 bl[55] br[55] wl[16] vdd gnd cell_6t
Xbit_r17_c55 bl[55] br[55] wl[17] vdd gnd cell_6t
Xbit_r18_c55 bl[55] br[55] wl[18] vdd gnd cell_6t
Xbit_r19_c55 bl[55] br[55] wl[19] vdd gnd cell_6t
Xbit_r20_c55 bl[55] br[55] wl[20] vdd gnd cell_6t
Xbit_r21_c55 bl[55] br[55] wl[21] vdd gnd cell_6t
Xbit_r22_c55 bl[55] br[55] wl[22] vdd gnd cell_6t
Xbit_r23_c55 bl[55] br[55] wl[23] vdd gnd cell_6t
Xbit_r24_c55 bl[55] br[55] wl[24] vdd gnd cell_6t
Xbit_r25_c55 bl[55] br[55] wl[25] vdd gnd cell_6t
Xbit_r26_c55 bl[55] br[55] wl[26] vdd gnd cell_6t
Xbit_r27_c55 bl[55] br[55] wl[27] vdd gnd cell_6t
Xbit_r28_c55 bl[55] br[55] wl[28] vdd gnd cell_6t
Xbit_r29_c55 bl[55] br[55] wl[29] vdd gnd cell_6t
Xbit_r30_c55 bl[55] br[55] wl[30] vdd gnd cell_6t
Xbit_r31_c55 bl[55] br[55] wl[31] vdd gnd cell_6t
Xbit_r32_c55 bl[55] br[55] wl[32] vdd gnd cell_6t
Xbit_r33_c55 bl[55] br[55] wl[33] vdd gnd cell_6t
Xbit_r34_c55 bl[55] br[55] wl[34] vdd gnd cell_6t
Xbit_r35_c55 bl[55] br[55] wl[35] vdd gnd cell_6t
Xbit_r36_c55 bl[55] br[55] wl[36] vdd gnd cell_6t
Xbit_r37_c55 bl[55] br[55] wl[37] vdd gnd cell_6t
Xbit_r38_c55 bl[55] br[55] wl[38] vdd gnd cell_6t
Xbit_r39_c55 bl[55] br[55] wl[39] vdd gnd cell_6t
Xbit_r40_c55 bl[55] br[55] wl[40] vdd gnd cell_6t
Xbit_r41_c55 bl[55] br[55] wl[41] vdd gnd cell_6t
Xbit_r42_c55 bl[55] br[55] wl[42] vdd gnd cell_6t
Xbit_r43_c55 bl[55] br[55] wl[43] vdd gnd cell_6t
Xbit_r44_c55 bl[55] br[55] wl[44] vdd gnd cell_6t
Xbit_r45_c55 bl[55] br[55] wl[45] vdd gnd cell_6t
Xbit_r46_c55 bl[55] br[55] wl[46] vdd gnd cell_6t
Xbit_r47_c55 bl[55] br[55] wl[47] vdd gnd cell_6t
Xbit_r48_c55 bl[55] br[55] wl[48] vdd gnd cell_6t
Xbit_r49_c55 bl[55] br[55] wl[49] vdd gnd cell_6t
Xbit_r50_c55 bl[55] br[55] wl[50] vdd gnd cell_6t
Xbit_r51_c55 bl[55] br[55] wl[51] vdd gnd cell_6t
Xbit_r52_c55 bl[55] br[55] wl[52] vdd gnd cell_6t
Xbit_r53_c55 bl[55] br[55] wl[53] vdd gnd cell_6t
Xbit_r54_c55 bl[55] br[55] wl[54] vdd gnd cell_6t
Xbit_r55_c55 bl[55] br[55] wl[55] vdd gnd cell_6t
Xbit_r56_c55 bl[55] br[55] wl[56] vdd gnd cell_6t
Xbit_r57_c55 bl[55] br[55] wl[57] vdd gnd cell_6t
Xbit_r58_c55 bl[55] br[55] wl[58] vdd gnd cell_6t
Xbit_r59_c55 bl[55] br[55] wl[59] vdd gnd cell_6t
Xbit_r60_c55 bl[55] br[55] wl[60] vdd gnd cell_6t
Xbit_r61_c55 bl[55] br[55] wl[61] vdd gnd cell_6t
Xbit_r62_c55 bl[55] br[55] wl[62] vdd gnd cell_6t
Xbit_r63_c55 bl[55] br[55] wl[63] vdd gnd cell_6t
Xbit_r64_c55 bl[55] br[55] wl[64] vdd gnd cell_6t
Xbit_r65_c55 bl[55] br[55] wl[65] vdd gnd cell_6t
Xbit_r66_c55 bl[55] br[55] wl[66] vdd gnd cell_6t
Xbit_r67_c55 bl[55] br[55] wl[67] vdd gnd cell_6t
Xbit_r68_c55 bl[55] br[55] wl[68] vdd gnd cell_6t
Xbit_r69_c55 bl[55] br[55] wl[69] vdd gnd cell_6t
Xbit_r70_c55 bl[55] br[55] wl[70] vdd gnd cell_6t
Xbit_r71_c55 bl[55] br[55] wl[71] vdd gnd cell_6t
Xbit_r72_c55 bl[55] br[55] wl[72] vdd gnd cell_6t
Xbit_r73_c55 bl[55] br[55] wl[73] vdd gnd cell_6t
Xbit_r74_c55 bl[55] br[55] wl[74] vdd gnd cell_6t
Xbit_r75_c55 bl[55] br[55] wl[75] vdd gnd cell_6t
Xbit_r76_c55 bl[55] br[55] wl[76] vdd gnd cell_6t
Xbit_r77_c55 bl[55] br[55] wl[77] vdd gnd cell_6t
Xbit_r78_c55 bl[55] br[55] wl[78] vdd gnd cell_6t
Xbit_r79_c55 bl[55] br[55] wl[79] vdd gnd cell_6t
Xbit_r80_c55 bl[55] br[55] wl[80] vdd gnd cell_6t
Xbit_r81_c55 bl[55] br[55] wl[81] vdd gnd cell_6t
Xbit_r82_c55 bl[55] br[55] wl[82] vdd gnd cell_6t
Xbit_r83_c55 bl[55] br[55] wl[83] vdd gnd cell_6t
Xbit_r84_c55 bl[55] br[55] wl[84] vdd gnd cell_6t
Xbit_r85_c55 bl[55] br[55] wl[85] vdd gnd cell_6t
Xbit_r86_c55 bl[55] br[55] wl[86] vdd gnd cell_6t
Xbit_r87_c55 bl[55] br[55] wl[87] vdd gnd cell_6t
Xbit_r88_c55 bl[55] br[55] wl[88] vdd gnd cell_6t
Xbit_r89_c55 bl[55] br[55] wl[89] vdd gnd cell_6t
Xbit_r90_c55 bl[55] br[55] wl[90] vdd gnd cell_6t
Xbit_r91_c55 bl[55] br[55] wl[91] vdd gnd cell_6t
Xbit_r92_c55 bl[55] br[55] wl[92] vdd gnd cell_6t
Xbit_r93_c55 bl[55] br[55] wl[93] vdd gnd cell_6t
Xbit_r94_c55 bl[55] br[55] wl[94] vdd gnd cell_6t
Xbit_r95_c55 bl[55] br[55] wl[95] vdd gnd cell_6t
Xbit_r96_c55 bl[55] br[55] wl[96] vdd gnd cell_6t
Xbit_r97_c55 bl[55] br[55] wl[97] vdd gnd cell_6t
Xbit_r98_c55 bl[55] br[55] wl[98] vdd gnd cell_6t
Xbit_r99_c55 bl[55] br[55] wl[99] vdd gnd cell_6t
Xbit_r100_c55 bl[55] br[55] wl[100] vdd gnd cell_6t
Xbit_r101_c55 bl[55] br[55] wl[101] vdd gnd cell_6t
Xbit_r102_c55 bl[55] br[55] wl[102] vdd gnd cell_6t
Xbit_r103_c55 bl[55] br[55] wl[103] vdd gnd cell_6t
Xbit_r104_c55 bl[55] br[55] wl[104] vdd gnd cell_6t
Xbit_r105_c55 bl[55] br[55] wl[105] vdd gnd cell_6t
Xbit_r106_c55 bl[55] br[55] wl[106] vdd gnd cell_6t
Xbit_r107_c55 bl[55] br[55] wl[107] vdd gnd cell_6t
Xbit_r108_c55 bl[55] br[55] wl[108] vdd gnd cell_6t
Xbit_r109_c55 bl[55] br[55] wl[109] vdd gnd cell_6t
Xbit_r110_c55 bl[55] br[55] wl[110] vdd gnd cell_6t
Xbit_r111_c55 bl[55] br[55] wl[111] vdd gnd cell_6t
Xbit_r112_c55 bl[55] br[55] wl[112] vdd gnd cell_6t
Xbit_r113_c55 bl[55] br[55] wl[113] vdd gnd cell_6t
Xbit_r114_c55 bl[55] br[55] wl[114] vdd gnd cell_6t
Xbit_r115_c55 bl[55] br[55] wl[115] vdd gnd cell_6t
Xbit_r116_c55 bl[55] br[55] wl[116] vdd gnd cell_6t
Xbit_r117_c55 bl[55] br[55] wl[117] vdd gnd cell_6t
Xbit_r118_c55 bl[55] br[55] wl[118] vdd gnd cell_6t
Xbit_r119_c55 bl[55] br[55] wl[119] vdd gnd cell_6t
Xbit_r120_c55 bl[55] br[55] wl[120] vdd gnd cell_6t
Xbit_r121_c55 bl[55] br[55] wl[121] vdd gnd cell_6t
Xbit_r122_c55 bl[55] br[55] wl[122] vdd gnd cell_6t
Xbit_r123_c55 bl[55] br[55] wl[123] vdd gnd cell_6t
Xbit_r124_c55 bl[55] br[55] wl[124] vdd gnd cell_6t
Xbit_r125_c55 bl[55] br[55] wl[125] vdd gnd cell_6t
Xbit_r126_c55 bl[55] br[55] wl[126] vdd gnd cell_6t
Xbit_r127_c55 bl[55] br[55] wl[127] vdd gnd cell_6t
Xbit_r128_c55 bl[55] br[55] wl[128] vdd gnd cell_6t
Xbit_r129_c55 bl[55] br[55] wl[129] vdd gnd cell_6t
Xbit_r130_c55 bl[55] br[55] wl[130] vdd gnd cell_6t
Xbit_r131_c55 bl[55] br[55] wl[131] vdd gnd cell_6t
Xbit_r132_c55 bl[55] br[55] wl[132] vdd gnd cell_6t
Xbit_r133_c55 bl[55] br[55] wl[133] vdd gnd cell_6t
Xbit_r134_c55 bl[55] br[55] wl[134] vdd gnd cell_6t
Xbit_r135_c55 bl[55] br[55] wl[135] vdd gnd cell_6t
Xbit_r136_c55 bl[55] br[55] wl[136] vdd gnd cell_6t
Xbit_r137_c55 bl[55] br[55] wl[137] vdd gnd cell_6t
Xbit_r138_c55 bl[55] br[55] wl[138] vdd gnd cell_6t
Xbit_r139_c55 bl[55] br[55] wl[139] vdd gnd cell_6t
Xbit_r140_c55 bl[55] br[55] wl[140] vdd gnd cell_6t
Xbit_r141_c55 bl[55] br[55] wl[141] vdd gnd cell_6t
Xbit_r142_c55 bl[55] br[55] wl[142] vdd gnd cell_6t
Xbit_r143_c55 bl[55] br[55] wl[143] vdd gnd cell_6t
Xbit_r144_c55 bl[55] br[55] wl[144] vdd gnd cell_6t
Xbit_r145_c55 bl[55] br[55] wl[145] vdd gnd cell_6t
Xbit_r146_c55 bl[55] br[55] wl[146] vdd gnd cell_6t
Xbit_r147_c55 bl[55] br[55] wl[147] vdd gnd cell_6t
Xbit_r148_c55 bl[55] br[55] wl[148] vdd gnd cell_6t
Xbit_r149_c55 bl[55] br[55] wl[149] vdd gnd cell_6t
Xbit_r150_c55 bl[55] br[55] wl[150] vdd gnd cell_6t
Xbit_r151_c55 bl[55] br[55] wl[151] vdd gnd cell_6t
Xbit_r152_c55 bl[55] br[55] wl[152] vdd gnd cell_6t
Xbit_r153_c55 bl[55] br[55] wl[153] vdd gnd cell_6t
Xbit_r154_c55 bl[55] br[55] wl[154] vdd gnd cell_6t
Xbit_r155_c55 bl[55] br[55] wl[155] vdd gnd cell_6t
Xbit_r156_c55 bl[55] br[55] wl[156] vdd gnd cell_6t
Xbit_r157_c55 bl[55] br[55] wl[157] vdd gnd cell_6t
Xbit_r158_c55 bl[55] br[55] wl[158] vdd gnd cell_6t
Xbit_r159_c55 bl[55] br[55] wl[159] vdd gnd cell_6t
Xbit_r160_c55 bl[55] br[55] wl[160] vdd gnd cell_6t
Xbit_r161_c55 bl[55] br[55] wl[161] vdd gnd cell_6t
Xbit_r162_c55 bl[55] br[55] wl[162] vdd gnd cell_6t
Xbit_r163_c55 bl[55] br[55] wl[163] vdd gnd cell_6t
Xbit_r164_c55 bl[55] br[55] wl[164] vdd gnd cell_6t
Xbit_r165_c55 bl[55] br[55] wl[165] vdd gnd cell_6t
Xbit_r166_c55 bl[55] br[55] wl[166] vdd gnd cell_6t
Xbit_r167_c55 bl[55] br[55] wl[167] vdd gnd cell_6t
Xbit_r168_c55 bl[55] br[55] wl[168] vdd gnd cell_6t
Xbit_r169_c55 bl[55] br[55] wl[169] vdd gnd cell_6t
Xbit_r170_c55 bl[55] br[55] wl[170] vdd gnd cell_6t
Xbit_r171_c55 bl[55] br[55] wl[171] vdd gnd cell_6t
Xbit_r172_c55 bl[55] br[55] wl[172] vdd gnd cell_6t
Xbit_r173_c55 bl[55] br[55] wl[173] vdd gnd cell_6t
Xbit_r174_c55 bl[55] br[55] wl[174] vdd gnd cell_6t
Xbit_r175_c55 bl[55] br[55] wl[175] vdd gnd cell_6t
Xbit_r176_c55 bl[55] br[55] wl[176] vdd gnd cell_6t
Xbit_r177_c55 bl[55] br[55] wl[177] vdd gnd cell_6t
Xbit_r178_c55 bl[55] br[55] wl[178] vdd gnd cell_6t
Xbit_r179_c55 bl[55] br[55] wl[179] vdd gnd cell_6t
Xbit_r180_c55 bl[55] br[55] wl[180] vdd gnd cell_6t
Xbit_r181_c55 bl[55] br[55] wl[181] vdd gnd cell_6t
Xbit_r182_c55 bl[55] br[55] wl[182] vdd gnd cell_6t
Xbit_r183_c55 bl[55] br[55] wl[183] vdd gnd cell_6t
Xbit_r184_c55 bl[55] br[55] wl[184] vdd gnd cell_6t
Xbit_r185_c55 bl[55] br[55] wl[185] vdd gnd cell_6t
Xbit_r186_c55 bl[55] br[55] wl[186] vdd gnd cell_6t
Xbit_r187_c55 bl[55] br[55] wl[187] vdd gnd cell_6t
Xbit_r188_c55 bl[55] br[55] wl[188] vdd gnd cell_6t
Xbit_r189_c55 bl[55] br[55] wl[189] vdd gnd cell_6t
Xbit_r190_c55 bl[55] br[55] wl[190] vdd gnd cell_6t
Xbit_r191_c55 bl[55] br[55] wl[191] vdd gnd cell_6t
Xbit_r192_c55 bl[55] br[55] wl[192] vdd gnd cell_6t
Xbit_r193_c55 bl[55] br[55] wl[193] vdd gnd cell_6t
Xbit_r194_c55 bl[55] br[55] wl[194] vdd gnd cell_6t
Xbit_r195_c55 bl[55] br[55] wl[195] vdd gnd cell_6t
Xbit_r196_c55 bl[55] br[55] wl[196] vdd gnd cell_6t
Xbit_r197_c55 bl[55] br[55] wl[197] vdd gnd cell_6t
Xbit_r198_c55 bl[55] br[55] wl[198] vdd gnd cell_6t
Xbit_r199_c55 bl[55] br[55] wl[199] vdd gnd cell_6t
Xbit_r200_c55 bl[55] br[55] wl[200] vdd gnd cell_6t
Xbit_r201_c55 bl[55] br[55] wl[201] vdd gnd cell_6t
Xbit_r202_c55 bl[55] br[55] wl[202] vdd gnd cell_6t
Xbit_r203_c55 bl[55] br[55] wl[203] vdd gnd cell_6t
Xbit_r204_c55 bl[55] br[55] wl[204] vdd gnd cell_6t
Xbit_r205_c55 bl[55] br[55] wl[205] vdd gnd cell_6t
Xbit_r206_c55 bl[55] br[55] wl[206] vdd gnd cell_6t
Xbit_r207_c55 bl[55] br[55] wl[207] vdd gnd cell_6t
Xbit_r208_c55 bl[55] br[55] wl[208] vdd gnd cell_6t
Xbit_r209_c55 bl[55] br[55] wl[209] vdd gnd cell_6t
Xbit_r210_c55 bl[55] br[55] wl[210] vdd gnd cell_6t
Xbit_r211_c55 bl[55] br[55] wl[211] vdd gnd cell_6t
Xbit_r212_c55 bl[55] br[55] wl[212] vdd gnd cell_6t
Xbit_r213_c55 bl[55] br[55] wl[213] vdd gnd cell_6t
Xbit_r214_c55 bl[55] br[55] wl[214] vdd gnd cell_6t
Xbit_r215_c55 bl[55] br[55] wl[215] vdd gnd cell_6t
Xbit_r216_c55 bl[55] br[55] wl[216] vdd gnd cell_6t
Xbit_r217_c55 bl[55] br[55] wl[217] vdd gnd cell_6t
Xbit_r218_c55 bl[55] br[55] wl[218] vdd gnd cell_6t
Xbit_r219_c55 bl[55] br[55] wl[219] vdd gnd cell_6t
Xbit_r220_c55 bl[55] br[55] wl[220] vdd gnd cell_6t
Xbit_r221_c55 bl[55] br[55] wl[221] vdd gnd cell_6t
Xbit_r222_c55 bl[55] br[55] wl[222] vdd gnd cell_6t
Xbit_r223_c55 bl[55] br[55] wl[223] vdd gnd cell_6t
Xbit_r224_c55 bl[55] br[55] wl[224] vdd gnd cell_6t
Xbit_r225_c55 bl[55] br[55] wl[225] vdd gnd cell_6t
Xbit_r226_c55 bl[55] br[55] wl[226] vdd gnd cell_6t
Xbit_r227_c55 bl[55] br[55] wl[227] vdd gnd cell_6t
Xbit_r228_c55 bl[55] br[55] wl[228] vdd gnd cell_6t
Xbit_r229_c55 bl[55] br[55] wl[229] vdd gnd cell_6t
Xbit_r230_c55 bl[55] br[55] wl[230] vdd gnd cell_6t
Xbit_r231_c55 bl[55] br[55] wl[231] vdd gnd cell_6t
Xbit_r232_c55 bl[55] br[55] wl[232] vdd gnd cell_6t
Xbit_r233_c55 bl[55] br[55] wl[233] vdd gnd cell_6t
Xbit_r234_c55 bl[55] br[55] wl[234] vdd gnd cell_6t
Xbit_r235_c55 bl[55] br[55] wl[235] vdd gnd cell_6t
Xbit_r236_c55 bl[55] br[55] wl[236] vdd gnd cell_6t
Xbit_r237_c55 bl[55] br[55] wl[237] vdd gnd cell_6t
Xbit_r238_c55 bl[55] br[55] wl[238] vdd gnd cell_6t
Xbit_r239_c55 bl[55] br[55] wl[239] vdd gnd cell_6t
Xbit_r240_c55 bl[55] br[55] wl[240] vdd gnd cell_6t
Xbit_r241_c55 bl[55] br[55] wl[241] vdd gnd cell_6t
Xbit_r242_c55 bl[55] br[55] wl[242] vdd gnd cell_6t
Xbit_r243_c55 bl[55] br[55] wl[243] vdd gnd cell_6t
Xbit_r244_c55 bl[55] br[55] wl[244] vdd gnd cell_6t
Xbit_r245_c55 bl[55] br[55] wl[245] vdd gnd cell_6t
Xbit_r246_c55 bl[55] br[55] wl[246] vdd gnd cell_6t
Xbit_r247_c55 bl[55] br[55] wl[247] vdd gnd cell_6t
Xbit_r248_c55 bl[55] br[55] wl[248] vdd gnd cell_6t
Xbit_r249_c55 bl[55] br[55] wl[249] vdd gnd cell_6t
Xbit_r250_c55 bl[55] br[55] wl[250] vdd gnd cell_6t
Xbit_r251_c55 bl[55] br[55] wl[251] vdd gnd cell_6t
Xbit_r252_c55 bl[55] br[55] wl[252] vdd gnd cell_6t
Xbit_r253_c55 bl[55] br[55] wl[253] vdd gnd cell_6t
Xbit_r254_c55 bl[55] br[55] wl[254] vdd gnd cell_6t
Xbit_r255_c55 bl[55] br[55] wl[255] vdd gnd cell_6t
Xbit_r0_c56 bl[56] br[56] wl[0] vdd gnd cell_6t
Xbit_r1_c56 bl[56] br[56] wl[1] vdd gnd cell_6t
Xbit_r2_c56 bl[56] br[56] wl[2] vdd gnd cell_6t
Xbit_r3_c56 bl[56] br[56] wl[3] vdd gnd cell_6t
Xbit_r4_c56 bl[56] br[56] wl[4] vdd gnd cell_6t
Xbit_r5_c56 bl[56] br[56] wl[5] vdd gnd cell_6t
Xbit_r6_c56 bl[56] br[56] wl[6] vdd gnd cell_6t
Xbit_r7_c56 bl[56] br[56] wl[7] vdd gnd cell_6t
Xbit_r8_c56 bl[56] br[56] wl[8] vdd gnd cell_6t
Xbit_r9_c56 bl[56] br[56] wl[9] vdd gnd cell_6t
Xbit_r10_c56 bl[56] br[56] wl[10] vdd gnd cell_6t
Xbit_r11_c56 bl[56] br[56] wl[11] vdd gnd cell_6t
Xbit_r12_c56 bl[56] br[56] wl[12] vdd gnd cell_6t
Xbit_r13_c56 bl[56] br[56] wl[13] vdd gnd cell_6t
Xbit_r14_c56 bl[56] br[56] wl[14] vdd gnd cell_6t
Xbit_r15_c56 bl[56] br[56] wl[15] vdd gnd cell_6t
Xbit_r16_c56 bl[56] br[56] wl[16] vdd gnd cell_6t
Xbit_r17_c56 bl[56] br[56] wl[17] vdd gnd cell_6t
Xbit_r18_c56 bl[56] br[56] wl[18] vdd gnd cell_6t
Xbit_r19_c56 bl[56] br[56] wl[19] vdd gnd cell_6t
Xbit_r20_c56 bl[56] br[56] wl[20] vdd gnd cell_6t
Xbit_r21_c56 bl[56] br[56] wl[21] vdd gnd cell_6t
Xbit_r22_c56 bl[56] br[56] wl[22] vdd gnd cell_6t
Xbit_r23_c56 bl[56] br[56] wl[23] vdd gnd cell_6t
Xbit_r24_c56 bl[56] br[56] wl[24] vdd gnd cell_6t
Xbit_r25_c56 bl[56] br[56] wl[25] vdd gnd cell_6t
Xbit_r26_c56 bl[56] br[56] wl[26] vdd gnd cell_6t
Xbit_r27_c56 bl[56] br[56] wl[27] vdd gnd cell_6t
Xbit_r28_c56 bl[56] br[56] wl[28] vdd gnd cell_6t
Xbit_r29_c56 bl[56] br[56] wl[29] vdd gnd cell_6t
Xbit_r30_c56 bl[56] br[56] wl[30] vdd gnd cell_6t
Xbit_r31_c56 bl[56] br[56] wl[31] vdd gnd cell_6t
Xbit_r32_c56 bl[56] br[56] wl[32] vdd gnd cell_6t
Xbit_r33_c56 bl[56] br[56] wl[33] vdd gnd cell_6t
Xbit_r34_c56 bl[56] br[56] wl[34] vdd gnd cell_6t
Xbit_r35_c56 bl[56] br[56] wl[35] vdd gnd cell_6t
Xbit_r36_c56 bl[56] br[56] wl[36] vdd gnd cell_6t
Xbit_r37_c56 bl[56] br[56] wl[37] vdd gnd cell_6t
Xbit_r38_c56 bl[56] br[56] wl[38] vdd gnd cell_6t
Xbit_r39_c56 bl[56] br[56] wl[39] vdd gnd cell_6t
Xbit_r40_c56 bl[56] br[56] wl[40] vdd gnd cell_6t
Xbit_r41_c56 bl[56] br[56] wl[41] vdd gnd cell_6t
Xbit_r42_c56 bl[56] br[56] wl[42] vdd gnd cell_6t
Xbit_r43_c56 bl[56] br[56] wl[43] vdd gnd cell_6t
Xbit_r44_c56 bl[56] br[56] wl[44] vdd gnd cell_6t
Xbit_r45_c56 bl[56] br[56] wl[45] vdd gnd cell_6t
Xbit_r46_c56 bl[56] br[56] wl[46] vdd gnd cell_6t
Xbit_r47_c56 bl[56] br[56] wl[47] vdd gnd cell_6t
Xbit_r48_c56 bl[56] br[56] wl[48] vdd gnd cell_6t
Xbit_r49_c56 bl[56] br[56] wl[49] vdd gnd cell_6t
Xbit_r50_c56 bl[56] br[56] wl[50] vdd gnd cell_6t
Xbit_r51_c56 bl[56] br[56] wl[51] vdd gnd cell_6t
Xbit_r52_c56 bl[56] br[56] wl[52] vdd gnd cell_6t
Xbit_r53_c56 bl[56] br[56] wl[53] vdd gnd cell_6t
Xbit_r54_c56 bl[56] br[56] wl[54] vdd gnd cell_6t
Xbit_r55_c56 bl[56] br[56] wl[55] vdd gnd cell_6t
Xbit_r56_c56 bl[56] br[56] wl[56] vdd gnd cell_6t
Xbit_r57_c56 bl[56] br[56] wl[57] vdd gnd cell_6t
Xbit_r58_c56 bl[56] br[56] wl[58] vdd gnd cell_6t
Xbit_r59_c56 bl[56] br[56] wl[59] vdd gnd cell_6t
Xbit_r60_c56 bl[56] br[56] wl[60] vdd gnd cell_6t
Xbit_r61_c56 bl[56] br[56] wl[61] vdd gnd cell_6t
Xbit_r62_c56 bl[56] br[56] wl[62] vdd gnd cell_6t
Xbit_r63_c56 bl[56] br[56] wl[63] vdd gnd cell_6t
Xbit_r64_c56 bl[56] br[56] wl[64] vdd gnd cell_6t
Xbit_r65_c56 bl[56] br[56] wl[65] vdd gnd cell_6t
Xbit_r66_c56 bl[56] br[56] wl[66] vdd gnd cell_6t
Xbit_r67_c56 bl[56] br[56] wl[67] vdd gnd cell_6t
Xbit_r68_c56 bl[56] br[56] wl[68] vdd gnd cell_6t
Xbit_r69_c56 bl[56] br[56] wl[69] vdd gnd cell_6t
Xbit_r70_c56 bl[56] br[56] wl[70] vdd gnd cell_6t
Xbit_r71_c56 bl[56] br[56] wl[71] vdd gnd cell_6t
Xbit_r72_c56 bl[56] br[56] wl[72] vdd gnd cell_6t
Xbit_r73_c56 bl[56] br[56] wl[73] vdd gnd cell_6t
Xbit_r74_c56 bl[56] br[56] wl[74] vdd gnd cell_6t
Xbit_r75_c56 bl[56] br[56] wl[75] vdd gnd cell_6t
Xbit_r76_c56 bl[56] br[56] wl[76] vdd gnd cell_6t
Xbit_r77_c56 bl[56] br[56] wl[77] vdd gnd cell_6t
Xbit_r78_c56 bl[56] br[56] wl[78] vdd gnd cell_6t
Xbit_r79_c56 bl[56] br[56] wl[79] vdd gnd cell_6t
Xbit_r80_c56 bl[56] br[56] wl[80] vdd gnd cell_6t
Xbit_r81_c56 bl[56] br[56] wl[81] vdd gnd cell_6t
Xbit_r82_c56 bl[56] br[56] wl[82] vdd gnd cell_6t
Xbit_r83_c56 bl[56] br[56] wl[83] vdd gnd cell_6t
Xbit_r84_c56 bl[56] br[56] wl[84] vdd gnd cell_6t
Xbit_r85_c56 bl[56] br[56] wl[85] vdd gnd cell_6t
Xbit_r86_c56 bl[56] br[56] wl[86] vdd gnd cell_6t
Xbit_r87_c56 bl[56] br[56] wl[87] vdd gnd cell_6t
Xbit_r88_c56 bl[56] br[56] wl[88] vdd gnd cell_6t
Xbit_r89_c56 bl[56] br[56] wl[89] vdd gnd cell_6t
Xbit_r90_c56 bl[56] br[56] wl[90] vdd gnd cell_6t
Xbit_r91_c56 bl[56] br[56] wl[91] vdd gnd cell_6t
Xbit_r92_c56 bl[56] br[56] wl[92] vdd gnd cell_6t
Xbit_r93_c56 bl[56] br[56] wl[93] vdd gnd cell_6t
Xbit_r94_c56 bl[56] br[56] wl[94] vdd gnd cell_6t
Xbit_r95_c56 bl[56] br[56] wl[95] vdd gnd cell_6t
Xbit_r96_c56 bl[56] br[56] wl[96] vdd gnd cell_6t
Xbit_r97_c56 bl[56] br[56] wl[97] vdd gnd cell_6t
Xbit_r98_c56 bl[56] br[56] wl[98] vdd gnd cell_6t
Xbit_r99_c56 bl[56] br[56] wl[99] vdd gnd cell_6t
Xbit_r100_c56 bl[56] br[56] wl[100] vdd gnd cell_6t
Xbit_r101_c56 bl[56] br[56] wl[101] vdd gnd cell_6t
Xbit_r102_c56 bl[56] br[56] wl[102] vdd gnd cell_6t
Xbit_r103_c56 bl[56] br[56] wl[103] vdd gnd cell_6t
Xbit_r104_c56 bl[56] br[56] wl[104] vdd gnd cell_6t
Xbit_r105_c56 bl[56] br[56] wl[105] vdd gnd cell_6t
Xbit_r106_c56 bl[56] br[56] wl[106] vdd gnd cell_6t
Xbit_r107_c56 bl[56] br[56] wl[107] vdd gnd cell_6t
Xbit_r108_c56 bl[56] br[56] wl[108] vdd gnd cell_6t
Xbit_r109_c56 bl[56] br[56] wl[109] vdd gnd cell_6t
Xbit_r110_c56 bl[56] br[56] wl[110] vdd gnd cell_6t
Xbit_r111_c56 bl[56] br[56] wl[111] vdd gnd cell_6t
Xbit_r112_c56 bl[56] br[56] wl[112] vdd gnd cell_6t
Xbit_r113_c56 bl[56] br[56] wl[113] vdd gnd cell_6t
Xbit_r114_c56 bl[56] br[56] wl[114] vdd gnd cell_6t
Xbit_r115_c56 bl[56] br[56] wl[115] vdd gnd cell_6t
Xbit_r116_c56 bl[56] br[56] wl[116] vdd gnd cell_6t
Xbit_r117_c56 bl[56] br[56] wl[117] vdd gnd cell_6t
Xbit_r118_c56 bl[56] br[56] wl[118] vdd gnd cell_6t
Xbit_r119_c56 bl[56] br[56] wl[119] vdd gnd cell_6t
Xbit_r120_c56 bl[56] br[56] wl[120] vdd gnd cell_6t
Xbit_r121_c56 bl[56] br[56] wl[121] vdd gnd cell_6t
Xbit_r122_c56 bl[56] br[56] wl[122] vdd gnd cell_6t
Xbit_r123_c56 bl[56] br[56] wl[123] vdd gnd cell_6t
Xbit_r124_c56 bl[56] br[56] wl[124] vdd gnd cell_6t
Xbit_r125_c56 bl[56] br[56] wl[125] vdd gnd cell_6t
Xbit_r126_c56 bl[56] br[56] wl[126] vdd gnd cell_6t
Xbit_r127_c56 bl[56] br[56] wl[127] vdd gnd cell_6t
Xbit_r128_c56 bl[56] br[56] wl[128] vdd gnd cell_6t
Xbit_r129_c56 bl[56] br[56] wl[129] vdd gnd cell_6t
Xbit_r130_c56 bl[56] br[56] wl[130] vdd gnd cell_6t
Xbit_r131_c56 bl[56] br[56] wl[131] vdd gnd cell_6t
Xbit_r132_c56 bl[56] br[56] wl[132] vdd gnd cell_6t
Xbit_r133_c56 bl[56] br[56] wl[133] vdd gnd cell_6t
Xbit_r134_c56 bl[56] br[56] wl[134] vdd gnd cell_6t
Xbit_r135_c56 bl[56] br[56] wl[135] vdd gnd cell_6t
Xbit_r136_c56 bl[56] br[56] wl[136] vdd gnd cell_6t
Xbit_r137_c56 bl[56] br[56] wl[137] vdd gnd cell_6t
Xbit_r138_c56 bl[56] br[56] wl[138] vdd gnd cell_6t
Xbit_r139_c56 bl[56] br[56] wl[139] vdd gnd cell_6t
Xbit_r140_c56 bl[56] br[56] wl[140] vdd gnd cell_6t
Xbit_r141_c56 bl[56] br[56] wl[141] vdd gnd cell_6t
Xbit_r142_c56 bl[56] br[56] wl[142] vdd gnd cell_6t
Xbit_r143_c56 bl[56] br[56] wl[143] vdd gnd cell_6t
Xbit_r144_c56 bl[56] br[56] wl[144] vdd gnd cell_6t
Xbit_r145_c56 bl[56] br[56] wl[145] vdd gnd cell_6t
Xbit_r146_c56 bl[56] br[56] wl[146] vdd gnd cell_6t
Xbit_r147_c56 bl[56] br[56] wl[147] vdd gnd cell_6t
Xbit_r148_c56 bl[56] br[56] wl[148] vdd gnd cell_6t
Xbit_r149_c56 bl[56] br[56] wl[149] vdd gnd cell_6t
Xbit_r150_c56 bl[56] br[56] wl[150] vdd gnd cell_6t
Xbit_r151_c56 bl[56] br[56] wl[151] vdd gnd cell_6t
Xbit_r152_c56 bl[56] br[56] wl[152] vdd gnd cell_6t
Xbit_r153_c56 bl[56] br[56] wl[153] vdd gnd cell_6t
Xbit_r154_c56 bl[56] br[56] wl[154] vdd gnd cell_6t
Xbit_r155_c56 bl[56] br[56] wl[155] vdd gnd cell_6t
Xbit_r156_c56 bl[56] br[56] wl[156] vdd gnd cell_6t
Xbit_r157_c56 bl[56] br[56] wl[157] vdd gnd cell_6t
Xbit_r158_c56 bl[56] br[56] wl[158] vdd gnd cell_6t
Xbit_r159_c56 bl[56] br[56] wl[159] vdd gnd cell_6t
Xbit_r160_c56 bl[56] br[56] wl[160] vdd gnd cell_6t
Xbit_r161_c56 bl[56] br[56] wl[161] vdd gnd cell_6t
Xbit_r162_c56 bl[56] br[56] wl[162] vdd gnd cell_6t
Xbit_r163_c56 bl[56] br[56] wl[163] vdd gnd cell_6t
Xbit_r164_c56 bl[56] br[56] wl[164] vdd gnd cell_6t
Xbit_r165_c56 bl[56] br[56] wl[165] vdd gnd cell_6t
Xbit_r166_c56 bl[56] br[56] wl[166] vdd gnd cell_6t
Xbit_r167_c56 bl[56] br[56] wl[167] vdd gnd cell_6t
Xbit_r168_c56 bl[56] br[56] wl[168] vdd gnd cell_6t
Xbit_r169_c56 bl[56] br[56] wl[169] vdd gnd cell_6t
Xbit_r170_c56 bl[56] br[56] wl[170] vdd gnd cell_6t
Xbit_r171_c56 bl[56] br[56] wl[171] vdd gnd cell_6t
Xbit_r172_c56 bl[56] br[56] wl[172] vdd gnd cell_6t
Xbit_r173_c56 bl[56] br[56] wl[173] vdd gnd cell_6t
Xbit_r174_c56 bl[56] br[56] wl[174] vdd gnd cell_6t
Xbit_r175_c56 bl[56] br[56] wl[175] vdd gnd cell_6t
Xbit_r176_c56 bl[56] br[56] wl[176] vdd gnd cell_6t
Xbit_r177_c56 bl[56] br[56] wl[177] vdd gnd cell_6t
Xbit_r178_c56 bl[56] br[56] wl[178] vdd gnd cell_6t
Xbit_r179_c56 bl[56] br[56] wl[179] vdd gnd cell_6t
Xbit_r180_c56 bl[56] br[56] wl[180] vdd gnd cell_6t
Xbit_r181_c56 bl[56] br[56] wl[181] vdd gnd cell_6t
Xbit_r182_c56 bl[56] br[56] wl[182] vdd gnd cell_6t
Xbit_r183_c56 bl[56] br[56] wl[183] vdd gnd cell_6t
Xbit_r184_c56 bl[56] br[56] wl[184] vdd gnd cell_6t
Xbit_r185_c56 bl[56] br[56] wl[185] vdd gnd cell_6t
Xbit_r186_c56 bl[56] br[56] wl[186] vdd gnd cell_6t
Xbit_r187_c56 bl[56] br[56] wl[187] vdd gnd cell_6t
Xbit_r188_c56 bl[56] br[56] wl[188] vdd gnd cell_6t
Xbit_r189_c56 bl[56] br[56] wl[189] vdd gnd cell_6t
Xbit_r190_c56 bl[56] br[56] wl[190] vdd gnd cell_6t
Xbit_r191_c56 bl[56] br[56] wl[191] vdd gnd cell_6t
Xbit_r192_c56 bl[56] br[56] wl[192] vdd gnd cell_6t
Xbit_r193_c56 bl[56] br[56] wl[193] vdd gnd cell_6t
Xbit_r194_c56 bl[56] br[56] wl[194] vdd gnd cell_6t
Xbit_r195_c56 bl[56] br[56] wl[195] vdd gnd cell_6t
Xbit_r196_c56 bl[56] br[56] wl[196] vdd gnd cell_6t
Xbit_r197_c56 bl[56] br[56] wl[197] vdd gnd cell_6t
Xbit_r198_c56 bl[56] br[56] wl[198] vdd gnd cell_6t
Xbit_r199_c56 bl[56] br[56] wl[199] vdd gnd cell_6t
Xbit_r200_c56 bl[56] br[56] wl[200] vdd gnd cell_6t
Xbit_r201_c56 bl[56] br[56] wl[201] vdd gnd cell_6t
Xbit_r202_c56 bl[56] br[56] wl[202] vdd gnd cell_6t
Xbit_r203_c56 bl[56] br[56] wl[203] vdd gnd cell_6t
Xbit_r204_c56 bl[56] br[56] wl[204] vdd gnd cell_6t
Xbit_r205_c56 bl[56] br[56] wl[205] vdd gnd cell_6t
Xbit_r206_c56 bl[56] br[56] wl[206] vdd gnd cell_6t
Xbit_r207_c56 bl[56] br[56] wl[207] vdd gnd cell_6t
Xbit_r208_c56 bl[56] br[56] wl[208] vdd gnd cell_6t
Xbit_r209_c56 bl[56] br[56] wl[209] vdd gnd cell_6t
Xbit_r210_c56 bl[56] br[56] wl[210] vdd gnd cell_6t
Xbit_r211_c56 bl[56] br[56] wl[211] vdd gnd cell_6t
Xbit_r212_c56 bl[56] br[56] wl[212] vdd gnd cell_6t
Xbit_r213_c56 bl[56] br[56] wl[213] vdd gnd cell_6t
Xbit_r214_c56 bl[56] br[56] wl[214] vdd gnd cell_6t
Xbit_r215_c56 bl[56] br[56] wl[215] vdd gnd cell_6t
Xbit_r216_c56 bl[56] br[56] wl[216] vdd gnd cell_6t
Xbit_r217_c56 bl[56] br[56] wl[217] vdd gnd cell_6t
Xbit_r218_c56 bl[56] br[56] wl[218] vdd gnd cell_6t
Xbit_r219_c56 bl[56] br[56] wl[219] vdd gnd cell_6t
Xbit_r220_c56 bl[56] br[56] wl[220] vdd gnd cell_6t
Xbit_r221_c56 bl[56] br[56] wl[221] vdd gnd cell_6t
Xbit_r222_c56 bl[56] br[56] wl[222] vdd gnd cell_6t
Xbit_r223_c56 bl[56] br[56] wl[223] vdd gnd cell_6t
Xbit_r224_c56 bl[56] br[56] wl[224] vdd gnd cell_6t
Xbit_r225_c56 bl[56] br[56] wl[225] vdd gnd cell_6t
Xbit_r226_c56 bl[56] br[56] wl[226] vdd gnd cell_6t
Xbit_r227_c56 bl[56] br[56] wl[227] vdd gnd cell_6t
Xbit_r228_c56 bl[56] br[56] wl[228] vdd gnd cell_6t
Xbit_r229_c56 bl[56] br[56] wl[229] vdd gnd cell_6t
Xbit_r230_c56 bl[56] br[56] wl[230] vdd gnd cell_6t
Xbit_r231_c56 bl[56] br[56] wl[231] vdd gnd cell_6t
Xbit_r232_c56 bl[56] br[56] wl[232] vdd gnd cell_6t
Xbit_r233_c56 bl[56] br[56] wl[233] vdd gnd cell_6t
Xbit_r234_c56 bl[56] br[56] wl[234] vdd gnd cell_6t
Xbit_r235_c56 bl[56] br[56] wl[235] vdd gnd cell_6t
Xbit_r236_c56 bl[56] br[56] wl[236] vdd gnd cell_6t
Xbit_r237_c56 bl[56] br[56] wl[237] vdd gnd cell_6t
Xbit_r238_c56 bl[56] br[56] wl[238] vdd gnd cell_6t
Xbit_r239_c56 bl[56] br[56] wl[239] vdd gnd cell_6t
Xbit_r240_c56 bl[56] br[56] wl[240] vdd gnd cell_6t
Xbit_r241_c56 bl[56] br[56] wl[241] vdd gnd cell_6t
Xbit_r242_c56 bl[56] br[56] wl[242] vdd gnd cell_6t
Xbit_r243_c56 bl[56] br[56] wl[243] vdd gnd cell_6t
Xbit_r244_c56 bl[56] br[56] wl[244] vdd gnd cell_6t
Xbit_r245_c56 bl[56] br[56] wl[245] vdd gnd cell_6t
Xbit_r246_c56 bl[56] br[56] wl[246] vdd gnd cell_6t
Xbit_r247_c56 bl[56] br[56] wl[247] vdd gnd cell_6t
Xbit_r248_c56 bl[56] br[56] wl[248] vdd gnd cell_6t
Xbit_r249_c56 bl[56] br[56] wl[249] vdd gnd cell_6t
Xbit_r250_c56 bl[56] br[56] wl[250] vdd gnd cell_6t
Xbit_r251_c56 bl[56] br[56] wl[251] vdd gnd cell_6t
Xbit_r252_c56 bl[56] br[56] wl[252] vdd gnd cell_6t
Xbit_r253_c56 bl[56] br[56] wl[253] vdd gnd cell_6t
Xbit_r254_c56 bl[56] br[56] wl[254] vdd gnd cell_6t
Xbit_r255_c56 bl[56] br[56] wl[255] vdd gnd cell_6t
Xbit_r0_c57 bl[57] br[57] wl[0] vdd gnd cell_6t
Xbit_r1_c57 bl[57] br[57] wl[1] vdd gnd cell_6t
Xbit_r2_c57 bl[57] br[57] wl[2] vdd gnd cell_6t
Xbit_r3_c57 bl[57] br[57] wl[3] vdd gnd cell_6t
Xbit_r4_c57 bl[57] br[57] wl[4] vdd gnd cell_6t
Xbit_r5_c57 bl[57] br[57] wl[5] vdd gnd cell_6t
Xbit_r6_c57 bl[57] br[57] wl[6] vdd gnd cell_6t
Xbit_r7_c57 bl[57] br[57] wl[7] vdd gnd cell_6t
Xbit_r8_c57 bl[57] br[57] wl[8] vdd gnd cell_6t
Xbit_r9_c57 bl[57] br[57] wl[9] vdd gnd cell_6t
Xbit_r10_c57 bl[57] br[57] wl[10] vdd gnd cell_6t
Xbit_r11_c57 bl[57] br[57] wl[11] vdd gnd cell_6t
Xbit_r12_c57 bl[57] br[57] wl[12] vdd gnd cell_6t
Xbit_r13_c57 bl[57] br[57] wl[13] vdd gnd cell_6t
Xbit_r14_c57 bl[57] br[57] wl[14] vdd gnd cell_6t
Xbit_r15_c57 bl[57] br[57] wl[15] vdd gnd cell_6t
Xbit_r16_c57 bl[57] br[57] wl[16] vdd gnd cell_6t
Xbit_r17_c57 bl[57] br[57] wl[17] vdd gnd cell_6t
Xbit_r18_c57 bl[57] br[57] wl[18] vdd gnd cell_6t
Xbit_r19_c57 bl[57] br[57] wl[19] vdd gnd cell_6t
Xbit_r20_c57 bl[57] br[57] wl[20] vdd gnd cell_6t
Xbit_r21_c57 bl[57] br[57] wl[21] vdd gnd cell_6t
Xbit_r22_c57 bl[57] br[57] wl[22] vdd gnd cell_6t
Xbit_r23_c57 bl[57] br[57] wl[23] vdd gnd cell_6t
Xbit_r24_c57 bl[57] br[57] wl[24] vdd gnd cell_6t
Xbit_r25_c57 bl[57] br[57] wl[25] vdd gnd cell_6t
Xbit_r26_c57 bl[57] br[57] wl[26] vdd gnd cell_6t
Xbit_r27_c57 bl[57] br[57] wl[27] vdd gnd cell_6t
Xbit_r28_c57 bl[57] br[57] wl[28] vdd gnd cell_6t
Xbit_r29_c57 bl[57] br[57] wl[29] vdd gnd cell_6t
Xbit_r30_c57 bl[57] br[57] wl[30] vdd gnd cell_6t
Xbit_r31_c57 bl[57] br[57] wl[31] vdd gnd cell_6t
Xbit_r32_c57 bl[57] br[57] wl[32] vdd gnd cell_6t
Xbit_r33_c57 bl[57] br[57] wl[33] vdd gnd cell_6t
Xbit_r34_c57 bl[57] br[57] wl[34] vdd gnd cell_6t
Xbit_r35_c57 bl[57] br[57] wl[35] vdd gnd cell_6t
Xbit_r36_c57 bl[57] br[57] wl[36] vdd gnd cell_6t
Xbit_r37_c57 bl[57] br[57] wl[37] vdd gnd cell_6t
Xbit_r38_c57 bl[57] br[57] wl[38] vdd gnd cell_6t
Xbit_r39_c57 bl[57] br[57] wl[39] vdd gnd cell_6t
Xbit_r40_c57 bl[57] br[57] wl[40] vdd gnd cell_6t
Xbit_r41_c57 bl[57] br[57] wl[41] vdd gnd cell_6t
Xbit_r42_c57 bl[57] br[57] wl[42] vdd gnd cell_6t
Xbit_r43_c57 bl[57] br[57] wl[43] vdd gnd cell_6t
Xbit_r44_c57 bl[57] br[57] wl[44] vdd gnd cell_6t
Xbit_r45_c57 bl[57] br[57] wl[45] vdd gnd cell_6t
Xbit_r46_c57 bl[57] br[57] wl[46] vdd gnd cell_6t
Xbit_r47_c57 bl[57] br[57] wl[47] vdd gnd cell_6t
Xbit_r48_c57 bl[57] br[57] wl[48] vdd gnd cell_6t
Xbit_r49_c57 bl[57] br[57] wl[49] vdd gnd cell_6t
Xbit_r50_c57 bl[57] br[57] wl[50] vdd gnd cell_6t
Xbit_r51_c57 bl[57] br[57] wl[51] vdd gnd cell_6t
Xbit_r52_c57 bl[57] br[57] wl[52] vdd gnd cell_6t
Xbit_r53_c57 bl[57] br[57] wl[53] vdd gnd cell_6t
Xbit_r54_c57 bl[57] br[57] wl[54] vdd gnd cell_6t
Xbit_r55_c57 bl[57] br[57] wl[55] vdd gnd cell_6t
Xbit_r56_c57 bl[57] br[57] wl[56] vdd gnd cell_6t
Xbit_r57_c57 bl[57] br[57] wl[57] vdd gnd cell_6t
Xbit_r58_c57 bl[57] br[57] wl[58] vdd gnd cell_6t
Xbit_r59_c57 bl[57] br[57] wl[59] vdd gnd cell_6t
Xbit_r60_c57 bl[57] br[57] wl[60] vdd gnd cell_6t
Xbit_r61_c57 bl[57] br[57] wl[61] vdd gnd cell_6t
Xbit_r62_c57 bl[57] br[57] wl[62] vdd gnd cell_6t
Xbit_r63_c57 bl[57] br[57] wl[63] vdd gnd cell_6t
Xbit_r64_c57 bl[57] br[57] wl[64] vdd gnd cell_6t
Xbit_r65_c57 bl[57] br[57] wl[65] vdd gnd cell_6t
Xbit_r66_c57 bl[57] br[57] wl[66] vdd gnd cell_6t
Xbit_r67_c57 bl[57] br[57] wl[67] vdd gnd cell_6t
Xbit_r68_c57 bl[57] br[57] wl[68] vdd gnd cell_6t
Xbit_r69_c57 bl[57] br[57] wl[69] vdd gnd cell_6t
Xbit_r70_c57 bl[57] br[57] wl[70] vdd gnd cell_6t
Xbit_r71_c57 bl[57] br[57] wl[71] vdd gnd cell_6t
Xbit_r72_c57 bl[57] br[57] wl[72] vdd gnd cell_6t
Xbit_r73_c57 bl[57] br[57] wl[73] vdd gnd cell_6t
Xbit_r74_c57 bl[57] br[57] wl[74] vdd gnd cell_6t
Xbit_r75_c57 bl[57] br[57] wl[75] vdd gnd cell_6t
Xbit_r76_c57 bl[57] br[57] wl[76] vdd gnd cell_6t
Xbit_r77_c57 bl[57] br[57] wl[77] vdd gnd cell_6t
Xbit_r78_c57 bl[57] br[57] wl[78] vdd gnd cell_6t
Xbit_r79_c57 bl[57] br[57] wl[79] vdd gnd cell_6t
Xbit_r80_c57 bl[57] br[57] wl[80] vdd gnd cell_6t
Xbit_r81_c57 bl[57] br[57] wl[81] vdd gnd cell_6t
Xbit_r82_c57 bl[57] br[57] wl[82] vdd gnd cell_6t
Xbit_r83_c57 bl[57] br[57] wl[83] vdd gnd cell_6t
Xbit_r84_c57 bl[57] br[57] wl[84] vdd gnd cell_6t
Xbit_r85_c57 bl[57] br[57] wl[85] vdd gnd cell_6t
Xbit_r86_c57 bl[57] br[57] wl[86] vdd gnd cell_6t
Xbit_r87_c57 bl[57] br[57] wl[87] vdd gnd cell_6t
Xbit_r88_c57 bl[57] br[57] wl[88] vdd gnd cell_6t
Xbit_r89_c57 bl[57] br[57] wl[89] vdd gnd cell_6t
Xbit_r90_c57 bl[57] br[57] wl[90] vdd gnd cell_6t
Xbit_r91_c57 bl[57] br[57] wl[91] vdd gnd cell_6t
Xbit_r92_c57 bl[57] br[57] wl[92] vdd gnd cell_6t
Xbit_r93_c57 bl[57] br[57] wl[93] vdd gnd cell_6t
Xbit_r94_c57 bl[57] br[57] wl[94] vdd gnd cell_6t
Xbit_r95_c57 bl[57] br[57] wl[95] vdd gnd cell_6t
Xbit_r96_c57 bl[57] br[57] wl[96] vdd gnd cell_6t
Xbit_r97_c57 bl[57] br[57] wl[97] vdd gnd cell_6t
Xbit_r98_c57 bl[57] br[57] wl[98] vdd gnd cell_6t
Xbit_r99_c57 bl[57] br[57] wl[99] vdd gnd cell_6t
Xbit_r100_c57 bl[57] br[57] wl[100] vdd gnd cell_6t
Xbit_r101_c57 bl[57] br[57] wl[101] vdd gnd cell_6t
Xbit_r102_c57 bl[57] br[57] wl[102] vdd gnd cell_6t
Xbit_r103_c57 bl[57] br[57] wl[103] vdd gnd cell_6t
Xbit_r104_c57 bl[57] br[57] wl[104] vdd gnd cell_6t
Xbit_r105_c57 bl[57] br[57] wl[105] vdd gnd cell_6t
Xbit_r106_c57 bl[57] br[57] wl[106] vdd gnd cell_6t
Xbit_r107_c57 bl[57] br[57] wl[107] vdd gnd cell_6t
Xbit_r108_c57 bl[57] br[57] wl[108] vdd gnd cell_6t
Xbit_r109_c57 bl[57] br[57] wl[109] vdd gnd cell_6t
Xbit_r110_c57 bl[57] br[57] wl[110] vdd gnd cell_6t
Xbit_r111_c57 bl[57] br[57] wl[111] vdd gnd cell_6t
Xbit_r112_c57 bl[57] br[57] wl[112] vdd gnd cell_6t
Xbit_r113_c57 bl[57] br[57] wl[113] vdd gnd cell_6t
Xbit_r114_c57 bl[57] br[57] wl[114] vdd gnd cell_6t
Xbit_r115_c57 bl[57] br[57] wl[115] vdd gnd cell_6t
Xbit_r116_c57 bl[57] br[57] wl[116] vdd gnd cell_6t
Xbit_r117_c57 bl[57] br[57] wl[117] vdd gnd cell_6t
Xbit_r118_c57 bl[57] br[57] wl[118] vdd gnd cell_6t
Xbit_r119_c57 bl[57] br[57] wl[119] vdd gnd cell_6t
Xbit_r120_c57 bl[57] br[57] wl[120] vdd gnd cell_6t
Xbit_r121_c57 bl[57] br[57] wl[121] vdd gnd cell_6t
Xbit_r122_c57 bl[57] br[57] wl[122] vdd gnd cell_6t
Xbit_r123_c57 bl[57] br[57] wl[123] vdd gnd cell_6t
Xbit_r124_c57 bl[57] br[57] wl[124] vdd gnd cell_6t
Xbit_r125_c57 bl[57] br[57] wl[125] vdd gnd cell_6t
Xbit_r126_c57 bl[57] br[57] wl[126] vdd gnd cell_6t
Xbit_r127_c57 bl[57] br[57] wl[127] vdd gnd cell_6t
Xbit_r128_c57 bl[57] br[57] wl[128] vdd gnd cell_6t
Xbit_r129_c57 bl[57] br[57] wl[129] vdd gnd cell_6t
Xbit_r130_c57 bl[57] br[57] wl[130] vdd gnd cell_6t
Xbit_r131_c57 bl[57] br[57] wl[131] vdd gnd cell_6t
Xbit_r132_c57 bl[57] br[57] wl[132] vdd gnd cell_6t
Xbit_r133_c57 bl[57] br[57] wl[133] vdd gnd cell_6t
Xbit_r134_c57 bl[57] br[57] wl[134] vdd gnd cell_6t
Xbit_r135_c57 bl[57] br[57] wl[135] vdd gnd cell_6t
Xbit_r136_c57 bl[57] br[57] wl[136] vdd gnd cell_6t
Xbit_r137_c57 bl[57] br[57] wl[137] vdd gnd cell_6t
Xbit_r138_c57 bl[57] br[57] wl[138] vdd gnd cell_6t
Xbit_r139_c57 bl[57] br[57] wl[139] vdd gnd cell_6t
Xbit_r140_c57 bl[57] br[57] wl[140] vdd gnd cell_6t
Xbit_r141_c57 bl[57] br[57] wl[141] vdd gnd cell_6t
Xbit_r142_c57 bl[57] br[57] wl[142] vdd gnd cell_6t
Xbit_r143_c57 bl[57] br[57] wl[143] vdd gnd cell_6t
Xbit_r144_c57 bl[57] br[57] wl[144] vdd gnd cell_6t
Xbit_r145_c57 bl[57] br[57] wl[145] vdd gnd cell_6t
Xbit_r146_c57 bl[57] br[57] wl[146] vdd gnd cell_6t
Xbit_r147_c57 bl[57] br[57] wl[147] vdd gnd cell_6t
Xbit_r148_c57 bl[57] br[57] wl[148] vdd gnd cell_6t
Xbit_r149_c57 bl[57] br[57] wl[149] vdd gnd cell_6t
Xbit_r150_c57 bl[57] br[57] wl[150] vdd gnd cell_6t
Xbit_r151_c57 bl[57] br[57] wl[151] vdd gnd cell_6t
Xbit_r152_c57 bl[57] br[57] wl[152] vdd gnd cell_6t
Xbit_r153_c57 bl[57] br[57] wl[153] vdd gnd cell_6t
Xbit_r154_c57 bl[57] br[57] wl[154] vdd gnd cell_6t
Xbit_r155_c57 bl[57] br[57] wl[155] vdd gnd cell_6t
Xbit_r156_c57 bl[57] br[57] wl[156] vdd gnd cell_6t
Xbit_r157_c57 bl[57] br[57] wl[157] vdd gnd cell_6t
Xbit_r158_c57 bl[57] br[57] wl[158] vdd gnd cell_6t
Xbit_r159_c57 bl[57] br[57] wl[159] vdd gnd cell_6t
Xbit_r160_c57 bl[57] br[57] wl[160] vdd gnd cell_6t
Xbit_r161_c57 bl[57] br[57] wl[161] vdd gnd cell_6t
Xbit_r162_c57 bl[57] br[57] wl[162] vdd gnd cell_6t
Xbit_r163_c57 bl[57] br[57] wl[163] vdd gnd cell_6t
Xbit_r164_c57 bl[57] br[57] wl[164] vdd gnd cell_6t
Xbit_r165_c57 bl[57] br[57] wl[165] vdd gnd cell_6t
Xbit_r166_c57 bl[57] br[57] wl[166] vdd gnd cell_6t
Xbit_r167_c57 bl[57] br[57] wl[167] vdd gnd cell_6t
Xbit_r168_c57 bl[57] br[57] wl[168] vdd gnd cell_6t
Xbit_r169_c57 bl[57] br[57] wl[169] vdd gnd cell_6t
Xbit_r170_c57 bl[57] br[57] wl[170] vdd gnd cell_6t
Xbit_r171_c57 bl[57] br[57] wl[171] vdd gnd cell_6t
Xbit_r172_c57 bl[57] br[57] wl[172] vdd gnd cell_6t
Xbit_r173_c57 bl[57] br[57] wl[173] vdd gnd cell_6t
Xbit_r174_c57 bl[57] br[57] wl[174] vdd gnd cell_6t
Xbit_r175_c57 bl[57] br[57] wl[175] vdd gnd cell_6t
Xbit_r176_c57 bl[57] br[57] wl[176] vdd gnd cell_6t
Xbit_r177_c57 bl[57] br[57] wl[177] vdd gnd cell_6t
Xbit_r178_c57 bl[57] br[57] wl[178] vdd gnd cell_6t
Xbit_r179_c57 bl[57] br[57] wl[179] vdd gnd cell_6t
Xbit_r180_c57 bl[57] br[57] wl[180] vdd gnd cell_6t
Xbit_r181_c57 bl[57] br[57] wl[181] vdd gnd cell_6t
Xbit_r182_c57 bl[57] br[57] wl[182] vdd gnd cell_6t
Xbit_r183_c57 bl[57] br[57] wl[183] vdd gnd cell_6t
Xbit_r184_c57 bl[57] br[57] wl[184] vdd gnd cell_6t
Xbit_r185_c57 bl[57] br[57] wl[185] vdd gnd cell_6t
Xbit_r186_c57 bl[57] br[57] wl[186] vdd gnd cell_6t
Xbit_r187_c57 bl[57] br[57] wl[187] vdd gnd cell_6t
Xbit_r188_c57 bl[57] br[57] wl[188] vdd gnd cell_6t
Xbit_r189_c57 bl[57] br[57] wl[189] vdd gnd cell_6t
Xbit_r190_c57 bl[57] br[57] wl[190] vdd gnd cell_6t
Xbit_r191_c57 bl[57] br[57] wl[191] vdd gnd cell_6t
Xbit_r192_c57 bl[57] br[57] wl[192] vdd gnd cell_6t
Xbit_r193_c57 bl[57] br[57] wl[193] vdd gnd cell_6t
Xbit_r194_c57 bl[57] br[57] wl[194] vdd gnd cell_6t
Xbit_r195_c57 bl[57] br[57] wl[195] vdd gnd cell_6t
Xbit_r196_c57 bl[57] br[57] wl[196] vdd gnd cell_6t
Xbit_r197_c57 bl[57] br[57] wl[197] vdd gnd cell_6t
Xbit_r198_c57 bl[57] br[57] wl[198] vdd gnd cell_6t
Xbit_r199_c57 bl[57] br[57] wl[199] vdd gnd cell_6t
Xbit_r200_c57 bl[57] br[57] wl[200] vdd gnd cell_6t
Xbit_r201_c57 bl[57] br[57] wl[201] vdd gnd cell_6t
Xbit_r202_c57 bl[57] br[57] wl[202] vdd gnd cell_6t
Xbit_r203_c57 bl[57] br[57] wl[203] vdd gnd cell_6t
Xbit_r204_c57 bl[57] br[57] wl[204] vdd gnd cell_6t
Xbit_r205_c57 bl[57] br[57] wl[205] vdd gnd cell_6t
Xbit_r206_c57 bl[57] br[57] wl[206] vdd gnd cell_6t
Xbit_r207_c57 bl[57] br[57] wl[207] vdd gnd cell_6t
Xbit_r208_c57 bl[57] br[57] wl[208] vdd gnd cell_6t
Xbit_r209_c57 bl[57] br[57] wl[209] vdd gnd cell_6t
Xbit_r210_c57 bl[57] br[57] wl[210] vdd gnd cell_6t
Xbit_r211_c57 bl[57] br[57] wl[211] vdd gnd cell_6t
Xbit_r212_c57 bl[57] br[57] wl[212] vdd gnd cell_6t
Xbit_r213_c57 bl[57] br[57] wl[213] vdd gnd cell_6t
Xbit_r214_c57 bl[57] br[57] wl[214] vdd gnd cell_6t
Xbit_r215_c57 bl[57] br[57] wl[215] vdd gnd cell_6t
Xbit_r216_c57 bl[57] br[57] wl[216] vdd gnd cell_6t
Xbit_r217_c57 bl[57] br[57] wl[217] vdd gnd cell_6t
Xbit_r218_c57 bl[57] br[57] wl[218] vdd gnd cell_6t
Xbit_r219_c57 bl[57] br[57] wl[219] vdd gnd cell_6t
Xbit_r220_c57 bl[57] br[57] wl[220] vdd gnd cell_6t
Xbit_r221_c57 bl[57] br[57] wl[221] vdd gnd cell_6t
Xbit_r222_c57 bl[57] br[57] wl[222] vdd gnd cell_6t
Xbit_r223_c57 bl[57] br[57] wl[223] vdd gnd cell_6t
Xbit_r224_c57 bl[57] br[57] wl[224] vdd gnd cell_6t
Xbit_r225_c57 bl[57] br[57] wl[225] vdd gnd cell_6t
Xbit_r226_c57 bl[57] br[57] wl[226] vdd gnd cell_6t
Xbit_r227_c57 bl[57] br[57] wl[227] vdd gnd cell_6t
Xbit_r228_c57 bl[57] br[57] wl[228] vdd gnd cell_6t
Xbit_r229_c57 bl[57] br[57] wl[229] vdd gnd cell_6t
Xbit_r230_c57 bl[57] br[57] wl[230] vdd gnd cell_6t
Xbit_r231_c57 bl[57] br[57] wl[231] vdd gnd cell_6t
Xbit_r232_c57 bl[57] br[57] wl[232] vdd gnd cell_6t
Xbit_r233_c57 bl[57] br[57] wl[233] vdd gnd cell_6t
Xbit_r234_c57 bl[57] br[57] wl[234] vdd gnd cell_6t
Xbit_r235_c57 bl[57] br[57] wl[235] vdd gnd cell_6t
Xbit_r236_c57 bl[57] br[57] wl[236] vdd gnd cell_6t
Xbit_r237_c57 bl[57] br[57] wl[237] vdd gnd cell_6t
Xbit_r238_c57 bl[57] br[57] wl[238] vdd gnd cell_6t
Xbit_r239_c57 bl[57] br[57] wl[239] vdd gnd cell_6t
Xbit_r240_c57 bl[57] br[57] wl[240] vdd gnd cell_6t
Xbit_r241_c57 bl[57] br[57] wl[241] vdd gnd cell_6t
Xbit_r242_c57 bl[57] br[57] wl[242] vdd gnd cell_6t
Xbit_r243_c57 bl[57] br[57] wl[243] vdd gnd cell_6t
Xbit_r244_c57 bl[57] br[57] wl[244] vdd gnd cell_6t
Xbit_r245_c57 bl[57] br[57] wl[245] vdd gnd cell_6t
Xbit_r246_c57 bl[57] br[57] wl[246] vdd gnd cell_6t
Xbit_r247_c57 bl[57] br[57] wl[247] vdd gnd cell_6t
Xbit_r248_c57 bl[57] br[57] wl[248] vdd gnd cell_6t
Xbit_r249_c57 bl[57] br[57] wl[249] vdd gnd cell_6t
Xbit_r250_c57 bl[57] br[57] wl[250] vdd gnd cell_6t
Xbit_r251_c57 bl[57] br[57] wl[251] vdd gnd cell_6t
Xbit_r252_c57 bl[57] br[57] wl[252] vdd gnd cell_6t
Xbit_r253_c57 bl[57] br[57] wl[253] vdd gnd cell_6t
Xbit_r254_c57 bl[57] br[57] wl[254] vdd gnd cell_6t
Xbit_r255_c57 bl[57] br[57] wl[255] vdd gnd cell_6t
Xbit_r0_c58 bl[58] br[58] wl[0] vdd gnd cell_6t
Xbit_r1_c58 bl[58] br[58] wl[1] vdd gnd cell_6t
Xbit_r2_c58 bl[58] br[58] wl[2] vdd gnd cell_6t
Xbit_r3_c58 bl[58] br[58] wl[3] vdd gnd cell_6t
Xbit_r4_c58 bl[58] br[58] wl[4] vdd gnd cell_6t
Xbit_r5_c58 bl[58] br[58] wl[5] vdd gnd cell_6t
Xbit_r6_c58 bl[58] br[58] wl[6] vdd gnd cell_6t
Xbit_r7_c58 bl[58] br[58] wl[7] vdd gnd cell_6t
Xbit_r8_c58 bl[58] br[58] wl[8] vdd gnd cell_6t
Xbit_r9_c58 bl[58] br[58] wl[9] vdd gnd cell_6t
Xbit_r10_c58 bl[58] br[58] wl[10] vdd gnd cell_6t
Xbit_r11_c58 bl[58] br[58] wl[11] vdd gnd cell_6t
Xbit_r12_c58 bl[58] br[58] wl[12] vdd gnd cell_6t
Xbit_r13_c58 bl[58] br[58] wl[13] vdd gnd cell_6t
Xbit_r14_c58 bl[58] br[58] wl[14] vdd gnd cell_6t
Xbit_r15_c58 bl[58] br[58] wl[15] vdd gnd cell_6t
Xbit_r16_c58 bl[58] br[58] wl[16] vdd gnd cell_6t
Xbit_r17_c58 bl[58] br[58] wl[17] vdd gnd cell_6t
Xbit_r18_c58 bl[58] br[58] wl[18] vdd gnd cell_6t
Xbit_r19_c58 bl[58] br[58] wl[19] vdd gnd cell_6t
Xbit_r20_c58 bl[58] br[58] wl[20] vdd gnd cell_6t
Xbit_r21_c58 bl[58] br[58] wl[21] vdd gnd cell_6t
Xbit_r22_c58 bl[58] br[58] wl[22] vdd gnd cell_6t
Xbit_r23_c58 bl[58] br[58] wl[23] vdd gnd cell_6t
Xbit_r24_c58 bl[58] br[58] wl[24] vdd gnd cell_6t
Xbit_r25_c58 bl[58] br[58] wl[25] vdd gnd cell_6t
Xbit_r26_c58 bl[58] br[58] wl[26] vdd gnd cell_6t
Xbit_r27_c58 bl[58] br[58] wl[27] vdd gnd cell_6t
Xbit_r28_c58 bl[58] br[58] wl[28] vdd gnd cell_6t
Xbit_r29_c58 bl[58] br[58] wl[29] vdd gnd cell_6t
Xbit_r30_c58 bl[58] br[58] wl[30] vdd gnd cell_6t
Xbit_r31_c58 bl[58] br[58] wl[31] vdd gnd cell_6t
Xbit_r32_c58 bl[58] br[58] wl[32] vdd gnd cell_6t
Xbit_r33_c58 bl[58] br[58] wl[33] vdd gnd cell_6t
Xbit_r34_c58 bl[58] br[58] wl[34] vdd gnd cell_6t
Xbit_r35_c58 bl[58] br[58] wl[35] vdd gnd cell_6t
Xbit_r36_c58 bl[58] br[58] wl[36] vdd gnd cell_6t
Xbit_r37_c58 bl[58] br[58] wl[37] vdd gnd cell_6t
Xbit_r38_c58 bl[58] br[58] wl[38] vdd gnd cell_6t
Xbit_r39_c58 bl[58] br[58] wl[39] vdd gnd cell_6t
Xbit_r40_c58 bl[58] br[58] wl[40] vdd gnd cell_6t
Xbit_r41_c58 bl[58] br[58] wl[41] vdd gnd cell_6t
Xbit_r42_c58 bl[58] br[58] wl[42] vdd gnd cell_6t
Xbit_r43_c58 bl[58] br[58] wl[43] vdd gnd cell_6t
Xbit_r44_c58 bl[58] br[58] wl[44] vdd gnd cell_6t
Xbit_r45_c58 bl[58] br[58] wl[45] vdd gnd cell_6t
Xbit_r46_c58 bl[58] br[58] wl[46] vdd gnd cell_6t
Xbit_r47_c58 bl[58] br[58] wl[47] vdd gnd cell_6t
Xbit_r48_c58 bl[58] br[58] wl[48] vdd gnd cell_6t
Xbit_r49_c58 bl[58] br[58] wl[49] vdd gnd cell_6t
Xbit_r50_c58 bl[58] br[58] wl[50] vdd gnd cell_6t
Xbit_r51_c58 bl[58] br[58] wl[51] vdd gnd cell_6t
Xbit_r52_c58 bl[58] br[58] wl[52] vdd gnd cell_6t
Xbit_r53_c58 bl[58] br[58] wl[53] vdd gnd cell_6t
Xbit_r54_c58 bl[58] br[58] wl[54] vdd gnd cell_6t
Xbit_r55_c58 bl[58] br[58] wl[55] vdd gnd cell_6t
Xbit_r56_c58 bl[58] br[58] wl[56] vdd gnd cell_6t
Xbit_r57_c58 bl[58] br[58] wl[57] vdd gnd cell_6t
Xbit_r58_c58 bl[58] br[58] wl[58] vdd gnd cell_6t
Xbit_r59_c58 bl[58] br[58] wl[59] vdd gnd cell_6t
Xbit_r60_c58 bl[58] br[58] wl[60] vdd gnd cell_6t
Xbit_r61_c58 bl[58] br[58] wl[61] vdd gnd cell_6t
Xbit_r62_c58 bl[58] br[58] wl[62] vdd gnd cell_6t
Xbit_r63_c58 bl[58] br[58] wl[63] vdd gnd cell_6t
Xbit_r64_c58 bl[58] br[58] wl[64] vdd gnd cell_6t
Xbit_r65_c58 bl[58] br[58] wl[65] vdd gnd cell_6t
Xbit_r66_c58 bl[58] br[58] wl[66] vdd gnd cell_6t
Xbit_r67_c58 bl[58] br[58] wl[67] vdd gnd cell_6t
Xbit_r68_c58 bl[58] br[58] wl[68] vdd gnd cell_6t
Xbit_r69_c58 bl[58] br[58] wl[69] vdd gnd cell_6t
Xbit_r70_c58 bl[58] br[58] wl[70] vdd gnd cell_6t
Xbit_r71_c58 bl[58] br[58] wl[71] vdd gnd cell_6t
Xbit_r72_c58 bl[58] br[58] wl[72] vdd gnd cell_6t
Xbit_r73_c58 bl[58] br[58] wl[73] vdd gnd cell_6t
Xbit_r74_c58 bl[58] br[58] wl[74] vdd gnd cell_6t
Xbit_r75_c58 bl[58] br[58] wl[75] vdd gnd cell_6t
Xbit_r76_c58 bl[58] br[58] wl[76] vdd gnd cell_6t
Xbit_r77_c58 bl[58] br[58] wl[77] vdd gnd cell_6t
Xbit_r78_c58 bl[58] br[58] wl[78] vdd gnd cell_6t
Xbit_r79_c58 bl[58] br[58] wl[79] vdd gnd cell_6t
Xbit_r80_c58 bl[58] br[58] wl[80] vdd gnd cell_6t
Xbit_r81_c58 bl[58] br[58] wl[81] vdd gnd cell_6t
Xbit_r82_c58 bl[58] br[58] wl[82] vdd gnd cell_6t
Xbit_r83_c58 bl[58] br[58] wl[83] vdd gnd cell_6t
Xbit_r84_c58 bl[58] br[58] wl[84] vdd gnd cell_6t
Xbit_r85_c58 bl[58] br[58] wl[85] vdd gnd cell_6t
Xbit_r86_c58 bl[58] br[58] wl[86] vdd gnd cell_6t
Xbit_r87_c58 bl[58] br[58] wl[87] vdd gnd cell_6t
Xbit_r88_c58 bl[58] br[58] wl[88] vdd gnd cell_6t
Xbit_r89_c58 bl[58] br[58] wl[89] vdd gnd cell_6t
Xbit_r90_c58 bl[58] br[58] wl[90] vdd gnd cell_6t
Xbit_r91_c58 bl[58] br[58] wl[91] vdd gnd cell_6t
Xbit_r92_c58 bl[58] br[58] wl[92] vdd gnd cell_6t
Xbit_r93_c58 bl[58] br[58] wl[93] vdd gnd cell_6t
Xbit_r94_c58 bl[58] br[58] wl[94] vdd gnd cell_6t
Xbit_r95_c58 bl[58] br[58] wl[95] vdd gnd cell_6t
Xbit_r96_c58 bl[58] br[58] wl[96] vdd gnd cell_6t
Xbit_r97_c58 bl[58] br[58] wl[97] vdd gnd cell_6t
Xbit_r98_c58 bl[58] br[58] wl[98] vdd gnd cell_6t
Xbit_r99_c58 bl[58] br[58] wl[99] vdd gnd cell_6t
Xbit_r100_c58 bl[58] br[58] wl[100] vdd gnd cell_6t
Xbit_r101_c58 bl[58] br[58] wl[101] vdd gnd cell_6t
Xbit_r102_c58 bl[58] br[58] wl[102] vdd gnd cell_6t
Xbit_r103_c58 bl[58] br[58] wl[103] vdd gnd cell_6t
Xbit_r104_c58 bl[58] br[58] wl[104] vdd gnd cell_6t
Xbit_r105_c58 bl[58] br[58] wl[105] vdd gnd cell_6t
Xbit_r106_c58 bl[58] br[58] wl[106] vdd gnd cell_6t
Xbit_r107_c58 bl[58] br[58] wl[107] vdd gnd cell_6t
Xbit_r108_c58 bl[58] br[58] wl[108] vdd gnd cell_6t
Xbit_r109_c58 bl[58] br[58] wl[109] vdd gnd cell_6t
Xbit_r110_c58 bl[58] br[58] wl[110] vdd gnd cell_6t
Xbit_r111_c58 bl[58] br[58] wl[111] vdd gnd cell_6t
Xbit_r112_c58 bl[58] br[58] wl[112] vdd gnd cell_6t
Xbit_r113_c58 bl[58] br[58] wl[113] vdd gnd cell_6t
Xbit_r114_c58 bl[58] br[58] wl[114] vdd gnd cell_6t
Xbit_r115_c58 bl[58] br[58] wl[115] vdd gnd cell_6t
Xbit_r116_c58 bl[58] br[58] wl[116] vdd gnd cell_6t
Xbit_r117_c58 bl[58] br[58] wl[117] vdd gnd cell_6t
Xbit_r118_c58 bl[58] br[58] wl[118] vdd gnd cell_6t
Xbit_r119_c58 bl[58] br[58] wl[119] vdd gnd cell_6t
Xbit_r120_c58 bl[58] br[58] wl[120] vdd gnd cell_6t
Xbit_r121_c58 bl[58] br[58] wl[121] vdd gnd cell_6t
Xbit_r122_c58 bl[58] br[58] wl[122] vdd gnd cell_6t
Xbit_r123_c58 bl[58] br[58] wl[123] vdd gnd cell_6t
Xbit_r124_c58 bl[58] br[58] wl[124] vdd gnd cell_6t
Xbit_r125_c58 bl[58] br[58] wl[125] vdd gnd cell_6t
Xbit_r126_c58 bl[58] br[58] wl[126] vdd gnd cell_6t
Xbit_r127_c58 bl[58] br[58] wl[127] vdd gnd cell_6t
Xbit_r128_c58 bl[58] br[58] wl[128] vdd gnd cell_6t
Xbit_r129_c58 bl[58] br[58] wl[129] vdd gnd cell_6t
Xbit_r130_c58 bl[58] br[58] wl[130] vdd gnd cell_6t
Xbit_r131_c58 bl[58] br[58] wl[131] vdd gnd cell_6t
Xbit_r132_c58 bl[58] br[58] wl[132] vdd gnd cell_6t
Xbit_r133_c58 bl[58] br[58] wl[133] vdd gnd cell_6t
Xbit_r134_c58 bl[58] br[58] wl[134] vdd gnd cell_6t
Xbit_r135_c58 bl[58] br[58] wl[135] vdd gnd cell_6t
Xbit_r136_c58 bl[58] br[58] wl[136] vdd gnd cell_6t
Xbit_r137_c58 bl[58] br[58] wl[137] vdd gnd cell_6t
Xbit_r138_c58 bl[58] br[58] wl[138] vdd gnd cell_6t
Xbit_r139_c58 bl[58] br[58] wl[139] vdd gnd cell_6t
Xbit_r140_c58 bl[58] br[58] wl[140] vdd gnd cell_6t
Xbit_r141_c58 bl[58] br[58] wl[141] vdd gnd cell_6t
Xbit_r142_c58 bl[58] br[58] wl[142] vdd gnd cell_6t
Xbit_r143_c58 bl[58] br[58] wl[143] vdd gnd cell_6t
Xbit_r144_c58 bl[58] br[58] wl[144] vdd gnd cell_6t
Xbit_r145_c58 bl[58] br[58] wl[145] vdd gnd cell_6t
Xbit_r146_c58 bl[58] br[58] wl[146] vdd gnd cell_6t
Xbit_r147_c58 bl[58] br[58] wl[147] vdd gnd cell_6t
Xbit_r148_c58 bl[58] br[58] wl[148] vdd gnd cell_6t
Xbit_r149_c58 bl[58] br[58] wl[149] vdd gnd cell_6t
Xbit_r150_c58 bl[58] br[58] wl[150] vdd gnd cell_6t
Xbit_r151_c58 bl[58] br[58] wl[151] vdd gnd cell_6t
Xbit_r152_c58 bl[58] br[58] wl[152] vdd gnd cell_6t
Xbit_r153_c58 bl[58] br[58] wl[153] vdd gnd cell_6t
Xbit_r154_c58 bl[58] br[58] wl[154] vdd gnd cell_6t
Xbit_r155_c58 bl[58] br[58] wl[155] vdd gnd cell_6t
Xbit_r156_c58 bl[58] br[58] wl[156] vdd gnd cell_6t
Xbit_r157_c58 bl[58] br[58] wl[157] vdd gnd cell_6t
Xbit_r158_c58 bl[58] br[58] wl[158] vdd gnd cell_6t
Xbit_r159_c58 bl[58] br[58] wl[159] vdd gnd cell_6t
Xbit_r160_c58 bl[58] br[58] wl[160] vdd gnd cell_6t
Xbit_r161_c58 bl[58] br[58] wl[161] vdd gnd cell_6t
Xbit_r162_c58 bl[58] br[58] wl[162] vdd gnd cell_6t
Xbit_r163_c58 bl[58] br[58] wl[163] vdd gnd cell_6t
Xbit_r164_c58 bl[58] br[58] wl[164] vdd gnd cell_6t
Xbit_r165_c58 bl[58] br[58] wl[165] vdd gnd cell_6t
Xbit_r166_c58 bl[58] br[58] wl[166] vdd gnd cell_6t
Xbit_r167_c58 bl[58] br[58] wl[167] vdd gnd cell_6t
Xbit_r168_c58 bl[58] br[58] wl[168] vdd gnd cell_6t
Xbit_r169_c58 bl[58] br[58] wl[169] vdd gnd cell_6t
Xbit_r170_c58 bl[58] br[58] wl[170] vdd gnd cell_6t
Xbit_r171_c58 bl[58] br[58] wl[171] vdd gnd cell_6t
Xbit_r172_c58 bl[58] br[58] wl[172] vdd gnd cell_6t
Xbit_r173_c58 bl[58] br[58] wl[173] vdd gnd cell_6t
Xbit_r174_c58 bl[58] br[58] wl[174] vdd gnd cell_6t
Xbit_r175_c58 bl[58] br[58] wl[175] vdd gnd cell_6t
Xbit_r176_c58 bl[58] br[58] wl[176] vdd gnd cell_6t
Xbit_r177_c58 bl[58] br[58] wl[177] vdd gnd cell_6t
Xbit_r178_c58 bl[58] br[58] wl[178] vdd gnd cell_6t
Xbit_r179_c58 bl[58] br[58] wl[179] vdd gnd cell_6t
Xbit_r180_c58 bl[58] br[58] wl[180] vdd gnd cell_6t
Xbit_r181_c58 bl[58] br[58] wl[181] vdd gnd cell_6t
Xbit_r182_c58 bl[58] br[58] wl[182] vdd gnd cell_6t
Xbit_r183_c58 bl[58] br[58] wl[183] vdd gnd cell_6t
Xbit_r184_c58 bl[58] br[58] wl[184] vdd gnd cell_6t
Xbit_r185_c58 bl[58] br[58] wl[185] vdd gnd cell_6t
Xbit_r186_c58 bl[58] br[58] wl[186] vdd gnd cell_6t
Xbit_r187_c58 bl[58] br[58] wl[187] vdd gnd cell_6t
Xbit_r188_c58 bl[58] br[58] wl[188] vdd gnd cell_6t
Xbit_r189_c58 bl[58] br[58] wl[189] vdd gnd cell_6t
Xbit_r190_c58 bl[58] br[58] wl[190] vdd gnd cell_6t
Xbit_r191_c58 bl[58] br[58] wl[191] vdd gnd cell_6t
Xbit_r192_c58 bl[58] br[58] wl[192] vdd gnd cell_6t
Xbit_r193_c58 bl[58] br[58] wl[193] vdd gnd cell_6t
Xbit_r194_c58 bl[58] br[58] wl[194] vdd gnd cell_6t
Xbit_r195_c58 bl[58] br[58] wl[195] vdd gnd cell_6t
Xbit_r196_c58 bl[58] br[58] wl[196] vdd gnd cell_6t
Xbit_r197_c58 bl[58] br[58] wl[197] vdd gnd cell_6t
Xbit_r198_c58 bl[58] br[58] wl[198] vdd gnd cell_6t
Xbit_r199_c58 bl[58] br[58] wl[199] vdd gnd cell_6t
Xbit_r200_c58 bl[58] br[58] wl[200] vdd gnd cell_6t
Xbit_r201_c58 bl[58] br[58] wl[201] vdd gnd cell_6t
Xbit_r202_c58 bl[58] br[58] wl[202] vdd gnd cell_6t
Xbit_r203_c58 bl[58] br[58] wl[203] vdd gnd cell_6t
Xbit_r204_c58 bl[58] br[58] wl[204] vdd gnd cell_6t
Xbit_r205_c58 bl[58] br[58] wl[205] vdd gnd cell_6t
Xbit_r206_c58 bl[58] br[58] wl[206] vdd gnd cell_6t
Xbit_r207_c58 bl[58] br[58] wl[207] vdd gnd cell_6t
Xbit_r208_c58 bl[58] br[58] wl[208] vdd gnd cell_6t
Xbit_r209_c58 bl[58] br[58] wl[209] vdd gnd cell_6t
Xbit_r210_c58 bl[58] br[58] wl[210] vdd gnd cell_6t
Xbit_r211_c58 bl[58] br[58] wl[211] vdd gnd cell_6t
Xbit_r212_c58 bl[58] br[58] wl[212] vdd gnd cell_6t
Xbit_r213_c58 bl[58] br[58] wl[213] vdd gnd cell_6t
Xbit_r214_c58 bl[58] br[58] wl[214] vdd gnd cell_6t
Xbit_r215_c58 bl[58] br[58] wl[215] vdd gnd cell_6t
Xbit_r216_c58 bl[58] br[58] wl[216] vdd gnd cell_6t
Xbit_r217_c58 bl[58] br[58] wl[217] vdd gnd cell_6t
Xbit_r218_c58 bl[58] br[58] wl[218] vdd gnd cell_6t
Xbit_r219_c58 bl[58] br[58] wl[219] vdd gnd cell_6t
Xbit_r220_c58 bl[58] br[58] wl[220] vdd gnd cell_6t
Xbit_r221_c58 bl[58] br[58] wl[221] vdd gnd cell_6t
Xbit_r222_c58 bl[58] br[58] wl[222] vdd gnd cell_6t
Xbit_r223_c58 bl[58] br[58] wl[223] vdd gnd cell_6t
Xbit_r224_c58 bl[58] br[58] wl[224] vdd gnd cell_6t
Xbit_r225_c58 bl[58] br[58] wl[225] vdd gnd cell_6t
Xbit_r226_c58 bl[58] br[58] wl[226] vdd gnd cell_6t
Xbit_r227_c58 bl[58] br[58] wl[227] vdd gnd cell_6t
Xbit_r228_c58 bl[58] br[58] wl[228] vdd gnd cell_6t
Xbit_r229_c58 bl[58] br[58] wl[229] vdd gnd cell_6t
Xbit_r230_c58 bl[58] br[58] wl[230] vdd gnd cell_6t
Xbit_r231_c58 bl[58] br[58] wl[231] vdd gnd cell_6t
Xbit_r232_c58 bl[58] br[58] wl[232] vdd gnd cell_6t
Xbit_r233_c58 bl[58] br[58] wl[233] vdd gnd cell_6t
Xbit_r234_c58 bl[58] br[58] wl[234] vdd gnd cell_6t
Xbit_r235_c58 bl[58] br[58] wl[235] vdd gnd cell_6t
Xbit_r236_c58 bl[58] br[58] wl[236] vdd gnd cell_6t
Xbit_r237_c58 bl[58] br[58] wl[237] vdd gnd cell_6t
Xbit_r238_c58 bl[58] br[58] wl[238] vdd gnd cell_6t
Xbit_r239_c58 bl[58] br[58] wl[239] vdd gnd cell_6t
Xbit_r240_c58 bl[58] br[58] wl[240] vdd gnd cell_6t
Xbit_r241_c58 bl[58] br[58] wl[241] vdd gnd cell_6t
Xbit_r242_c58 bl[58] br[58] wl[242] vdd gnd cell_6t
Xbit_r243_c58 bl[58] br[58] wl[243] vdd gnd cell_6t
Xbit_r244_c58 bl[58] br[58] wl[244] vdd gnd cell_6t
Xbit_r245_c58 bl[58] br[58] wl[245] vdd gnd cell_6t
Xbit_r246_c58 bl[58] br[58] wl[246] vdd gnd cell_6t
Xbit_r247_c58 bl[58] br[58] wl[247] vdd gnd cell_6t
Xbit_r248_c58 bl[58] br[58] wl[248] vdd gnd cell_6t
Xbit_r249_c58 bl[58] br[58] wl[249] vdd gnd cell_6t
Xbit_r250_c58 bl[58] br[58] wl[250] vdd gnd cell_6t
Xbit_r251_c58 bl[58] br[58] wl[251] vdd gnd cell_6t
Xbit_r252_c58 bl[58] br[58] wl[252] vdd gnd cell_6t
Xbit_r253_c58 bl[58] br[58] wl[253] vdd gnd cell_6t
Xbit_r254_c58 bl[58] br[58] wl[254] vdd gnd cell_6t
Xbit_r255_c58 bl[58] br[58] wl[255] vdd gnd cell_6t
Xbit_r0_c59 bl[59] br[59] wl[0] vdd gnd cell_6t
Xbit_r1_c59 bl[59] br[59] wl[1] vdd gnd cell_6t
Xbit_r2_c59 bl[59] br[59] wl[2] vdd gnd cell_6t
Xbit_r3_c59 bl[59] br[59] wl[3] vdd gnd cell_6t
Xbit_r4_c59 bl[59] br[59] wl[4] vdd gnd cell_6t
Xbit_r5_c59 bl[59] br[59] wl[5] vdd gnd cell_6t
Xbit_r6_c59 bl[59] br[59] wl[6] vdd gnd cell_6t
Xbit_r7_c59 bl[59] br[59] wl[7] vdd gnd cell_6t
Xbit_r8_c59 bl[59] br[59] wl[8] vdd gnd cell_6t
Xbit_r9_c59 bl[59] br[59] wl[9] vdd gnd cell_6t
Xbit_r10_c59 bl[59] br[59] wl[10] vdd gnd cell_6t
Xbit_r11_c59 bl[59] br[59] wl[11] vdd gnd cell_6t
Xbit_r12_c59 bl[59] br[59] wl[12] vdd gnd cell_6t
Xbit_r13_c59 bl[59] br[59] wl[13] vdd gnd cell_6t
Xbit_r14_c59 bl[59] br[59] wl[14] vdd gnd cell_6t
Xbit_r15_c59 bl[59] br[59] wl[15] vdd gnd cell_6t
Xbit_r16_c59 bl[59] br[59] wl[16] vdd gnd cell_6t
Xbit_r17_c59 bl[59] br[59] wl[17] vdd gnd cell_6t
Xbit_r18_c59 bl[59] br[59] wl[18] vdd gnd cell_6t
Xbit_r19_c59 bl[59] br[59] wl[19] vdd gnd cell_6t
Xbit_r20_c59 bl[59] br[59] wl[20] vdd gnd cell_6t
Xbit_r21_c59 bl[59] br[59] wl[21] vdd gnd cell_6t
Xbit_r22_c59 bl[59] br[59] wl[22] vdd gnd cell_6t
Xbit_r23_c59 bl[59] br[59] wl[23] vdd gnd cell_6t
Xbit_r24_c59 bl[59] br[59] wl[24] vdd gnd cell_6t
Xbit_r25_c59 bl[59] br[59] wl[25] vdd gnd cell_6t
Xbit_r26_c59 bl[59] br[59] wl[26] vdd gnd cell_6t
Xbit_r27_c59 bl[59] br[59] wl[27] vdd gnd cell_6t
Xbit_r28_c59 bl[59] br[59] wl[28] vdd gnd cell_6t
Xbit_r29_c59 bl[59] br[59] wl[29] vdd gnd cell_6t
Xbit_r30_c59 bl[59] br[59] wl[30] vdd gnd cell_6t
Xbit_r31_c59 bl[59] br[59] wl[31] vdd gnd cell_6t
Xbit_r32_c59 bl[59] br[59] wl[32] vdd gnd cell_6t
Xbit_r33_c59 bl[59] br[59] wl[33] vdd gnd cell_6t
Xbit_r34_c59 bl[59] br[59] wl[34] vdd gnd cell_6t
Xbit_r35_c59 bl[59] br[59] wl[35] vdd gnd cell_6t
Xbit_r36_c59 bl[59] br[59] wl[36] vdd gnd cell_6t
Xbit_r37_c59 bl[59] br[59] wl[37] vdd gnd cell_6t
Xbit_r38_c59 bl[59] br[59] wl[38] vdd gnd cell_6t
Xbit_r39_c59 bl[59] br[59] wl[39] vdd gnd cell_6t
Xbit_r40_c59 bl[59] br[59] wl[40] vdd gnd cell_6t
Xbit_r41_c59 bl[59] br[59] wl[41] vdd gnd cell_6t
Xbit_r42_c59 bl[59] br[59] wl[42] vdd gnd cell_6t
Xbit_r43_c59 bl[59] br[59] wl[43] vdd gnd cell_6t
Xbit_r44_c59 bl[59] br[59] wl[44] vdd gnd cell_6t
Xbit_r45_c59 bl[59] br[59] wl[45] vdd gnd cell_6t
Xbit_r46_c59 bl[59] br[59] wl[46] vdd gnd cell_6t
Xbit_r47_c59 bl[59] br[59] wl[47] vdd gnd cell_6t
Xbit_r48_c59 bl[59] br[59] wl[48] vdd gnd cell_6t
Xbit_r49_c59 bl[59] br[59] wl[49] vdd gnd cell_6t
Xbit_r50_c59 bl[59] br[59] wl[50] vdd gnd cell_6t
Xbit_r51_c59 bl[59] br[59] wl[51] vdd gnd cell_6t
Xbit_r52_c59 bl[59] br[59] wl[52] vdd gnd cell_6t
Xbit_r53_c59 bl[59] br[59] wl[53] vdd gnd cell_6t
Xbit_r54_c59 bl[59] br[59] wl[54] vdd gnd cell_6t
Xbit_r55_c59 bl[59] br[59] wl[55] vdd gnd cell_6t
Xbit_r56_c59 bl[59] br[59] wl[56] vdd gnd cell_6t
Xbit_r57_c59 bl[59] br[59] wl[57] vdd gnd cell_6t
Xbit_r58_c59 bl[59] br[59] wl[58] vdd gnd cell_6t
Xbit_r59_c59 bl[59] br[59] wl[59] vdd gnd cell_6t
Xbit_r60_c59 bl[59] br[59] wl[60] vdd gnd cell_6t
Xbit_r61_c59 bl[59] br[59] wl[61] vdd gnd cell_6t
Xbit_r62_c59 bl[59] br[59] wl[62] vdd gnd cell_6t
Xbit_r63_c59 bl[59] br[59] wl[63] vdd gnd cell_6t
Xbit_r64_c59 bl[59] br[59] wl[64] vdd gnd cell_6t
Xbit_r65_c59 bl[59] br[59] wl[65] vdd gnd cell_6t
Xbit_r66_c59 bl[59] br[59] wl[66] vdd gnd cell_6t
Xbit_r67_c59 bl[59] br[59] wl[67] vdd gnd cell_6t
Xbit_r68_c59 bl[59] br[59] wl[68] vdd gnd cell_6t
Xbit_r69_c59 bl[59] br[59] wl[69] vdd gnd cell_6t
Xbit_r70_c59 bl[59] br[59] wl[70] vdd gnd cell_6t
Xbit_r71_c59 bl[59] br[59] wl[71] vdd gnd cell_6t
Xbit_r72_c59 bl[59] br[59] wl[72] vdd gnd cell_6t
Xbit_r73_c59 bl[59] br[59] wl[73] vdd gnd cell_6t
Xbit_r74_c59 bl[59] br[59] wl[74] vdd gnd cell_6t
Xbit_r75_c59 bl[59] br[59] wl[75] vdd gnd cell_6t
Xbit_r76_c59 bl[59] br[59] wl[76] vdd gnd cell_6t
Xbit_r77_c59 bl[59] br[59] wl[77] vdd gnd cell_6t
Xbit_r78_c59 bl[59] br[59] wl[78] vdd gnd cell_6t
Xbit_r79_c59 bl[59] br[59] wl[79] vdd gnd cell_6t
Xbit_r80_c59 bl[59] br[59] wl[80] vdd gnd cell_6t
Xbit_r81_c59 bl[59] br[59] wl[81] vdd gnd cell_6t
Xbit_r82_c59 bl[59] br[59] wl[82] vdd gnd cell_6t
Xbit_r83_c59 bl[59] br[59] wl[83] vdd gnd cell_6t
Xbit_r84_c59 bl[59] br[59] wl[84] vdd gnd cell_6t
Xbit_r85_c59 bl[59] br[59] wl[85] vdd gnd cell_6t
Xbit_r86_c59 bl[59] br[59] wl[86] vdd gnd cell_6t
Xbit_r87_c59 bl[59] br[59] wl[87] vdd gnd cell_6t
Xbit_r88_c59 bl[59] br[59] wl[88] vdd gnd cell_6t
Xbit_r89_c59 bl[59] br[59] wl[89] vdd gnd cell_6t
Xbit_r90_c59 bl[59] br[59] wl[90] vdd gnd cell_6t
Xbit_r91_c59 bl[59] br[59] wl[91] vdd gnd cell_6t
Xbit_r92_c59 bl[59] br[59] wl[92] vdd gnd cell_6t
Xbit_r93_c59 bl[59] br[59] wl[93] vdd gnd cell_6t
Xbit_r94_c59 bl[59] br[59] wl[94] vdd gnd cell_6t
Xbit_r95_c59 bl[59] br[59] wl[95] vdd gnd cell_6t
Xbit_r96_c59 bl[59] br[59] wl[96] vdd gnd cell_6t
Xbit_r97_c59 bl[59] br[59] wl[97] vdd gnd cell_6t
Xbit_r98_c59 bl[59] br[59] wl[98] vdd gnd cell_6t
Xbit_r99_c59 bl[59] br[59] wl[99] vdd gnd cell_6t
Xbit_r100_c59 bl[59] br[59] wl[100] vdd gnd cell_6t
Xbit_r101_c59 bl[59] br[59] wl[101] vdd gnd cell_6t
Xbit_r102_c59 bl[59] br[59] wl[102] vdd gnd cell_6t
Xbit_r103_c59 bl[59] br[59] wl[103] vdd gnd cell_6t
Xbit_r104_c59 bl[59] br[59] wl[104] vdd gnd cell_6t
Xbit_r105_c59 bl[59] br[59] wl[105] vdd gnd cell_6t
Xbit_r106_c59 bl[59] br[59] wl[106] vdd gnd cell_6t
Xbit_r107_c59 bl[59] br[59] wl[107] vdd gnd cell_6t
Xbit_r108_c59 bl[59] br[59] wl[108] vdd gnd cell_6t
Xbit_r109_c59 bl[59] br[59] wl[109] vdd gnd cell_6t
Xbit_r110_c59 bl[59] br[59] wl[110] vdd gnd cell_6t
Xbit_r111_c59 bl[59] br[59] wl[111] vdd gnd cell_6t
Xbit_r112_c59 bl[59] br[59] wl[112] vdd gnd cell_6t
Xbit_r113_c59 bl[59] br[59] wl[113] vdd gnd cell_6t
Xbit_r114_c59 bl[59] br[59] wl[114] vdd gnd cell_6t
Xbit_r115_c59 bl[59] br[59] wl[115] vdd gnd cell_6t
Xbit_r116_c59 bl[59] br[59] wl[116] vdd gnd cell_6t
Xbit_r117_c59 bl[59] br[59] wl[117] vdd gnd cell_6t
Xbit_r118_c59 bl[59] br[59] wl[118] vdd gnd cell_6t
Xbit_r119_c59 bl[59] br[59] wl[119] vdd gnd cell_6t
Xbit_r120_c59 bl[59] br[59] wl[120] vdd gnd cell_6t
Xbit_r121_c59 bl[59] br[59] wl[121] vdd gnd cell_6t
Xbit_r122_c59 bl[59] br[59] wl[122] vdd gnd cell_6t
Xbit_r123_c59 bl[59] br[59] wl[123] vdd gnd cell_6t
Xbit_r124_c59 bl[59] br[59] wl[124] vdd gnd cell_6t
Xbit_r125_c59 bl[59] br[59] wl[125] vdd gnd cell_6t
Xbit_r126_c59 bl[59] br[59] wl[126] vdd gnd cell_6t
Xbit_r127_c59 bl[59] br[59] wl[127] vdd gnd cell_6t
Xbit_r128_c59 bl[59] br[59] wl[128] vdd gnd cell_6t
Xbit_r129_c59 bl[59] br[59] wl[129] vdd gnd cell_6t
Xbit_r130_c59 bl[59] br[59] wl[130] vdd gnd cell_6t
Xbit_r131_c59 bl[59] br[59] wl[131] vdd gnd cell_6t
Xbit_r132_c59 bl[59] br[59] wl[132] vdd gnd cell_6t
Xbit_r133_c59 bl[59] br[59] wl[133] vdd gnd cell_6t
Xbit_r134_c59 bl[59] br[59] wl[134] vdd gnd cell_6t
Xbit_r135_c59 bl[59] br[59] wl[135] vdd gnd cell_6t
Xbit_r136_c59 bl[59] br[59] wl[136] vdd gnd cell_6t
Xbit_r137_c59 bl[59] br[59] wl[137] vdd gnd cell_6t
Xbit_r138_c59 bl[59] br[59] wl[138] vdd gnd cell_6t
Xbit_r139_c59 bl[59] br[59] wl[139] vdd gnd cell_6t
Xbit_r140_c59 bl[59] br[59] wl[140] vdd gnd cell_6t
Xbit_r141_c59 bl[59] br[59] wl[141] vdd gnd cell_6t
Xbit_r142_c59 bl[59] br[59] wl[142] vdd gnd cell_6t
Xbit_r143_c59 bl[59] br[59] wl[143] vdd gnd cell_6t
Xbit_r144_c59 bl[59] br[59] wl[144] vdd gnd cell_6t
Xbit_r145_c59 bl[59] br[59] wl[145] vdd gnd cell_6t
Xbit_r146_c59 bl[59] br[59] wl[146] vdd gnd cell_6t
Xbit_r147_c59 bl[59] br[59] wl[147] vdd gnd cell_6t
Xbit_r148_c59 bl[59] br[59] wl[148] vdd gnd cell_6t
Xbit_r149_c59 bl[59] br[59] wl[149] vdd gnd cell_6t
Xbit_r150_c59 bl[59] br[59] wl[150] vdd gnd cell_6t
Xbit_r151_c59 bl[59] br[59] wl[151] vdd gnd cell_6t
Xbit_r152_c59 bl[59] br[59] wl[152] vdd gnd cell_6t
Xbit_r153_c59 bl[59] br[59] wl[153] vdd gnd cell_6t
Xbit_r154_c59 bl[59] br[59] wl[154] vdd gnd cell_6t
Xbit_r155_c59 bl[59] br[59] wl[155] vdd gnd cell_6t
Xbit_r156_c59 bl[59] br[59] wl[156] vdd gnd cell_6t
Xbit_r157_c59 bl[59] br[59] wl[157] vdd gnd cell_6t
Xbit_r158_c59 bl[59] br[59] wl[158] vdd gnd cell_6t
Xbit_r159_c59 bl[59] br[59] wl[159] vdd gnd cell_6t
Xbit_r160_c59 bl[59] br[59] wl[160] vdd gnd cell_6t
Xbit_r161_c59 bl[59] br[59] wl[161] vdd gnd cell_6t
Xbit_r162_c59 bl[59] br[59] wl[162] vdd gnd cell_6t
Xbit_r163_c59 bl[59] br[59] wl[163] vdd gnd cell_6t
Xbit_r164_c59 bl[59] br[59] wl[164] vdd gnd cell_6t
Xbit_r165_c59 bl[59] br[59] wl[165] vdd gnd cell_6t
Xbit_r166_c59 bl[59] br[59] wl[166] vdd gnd cell_6t
Xbit_r167_c59 bl[59] br[59] wl[167] vdd gnd cell_6t
Xbit_r168_c59 bl[59] br[59] wl[168] vdd gnd cell_6t
Xbit_r169_c59 bl[59] br[59] wl[169] vdd gnd cell_6t
Xbit_r170_c59 bl[59] br[59] wl[170] vdd gnd cell_6t
Xbit_r171_c59 bl[59] br[59] wl[171] vdd gnd cell_6t
Xbit_r172_c59 bl[59] br[59] wl[172] vdd gnd cell_6t
Xbit_r173_c59 bl[59] br[59] wl[173] vdd gnd cell_6t
Xbit_r174_c59 bl[59] br[59] wl[174] vdd gnd cell_6t
Xbit_r175_c59 bl[59] br[59] wl[175] vdd gnd cell_6t
Xbit_r176_c59 bl[59] br[59] wl[176] vdd gnd cell_6t
Xbit_r177_c59 bl[59] br[59] wl[177] vdd gnd cell_6t
Xbit_r178_c59 bl[59] br[59] wl[178] vdd gnd cell_6t
Xbit_r179_c59 bl[59] br[59] wl[179] vdd gnd cell_6t
Xbit_r180_c59 bl[59] br[59] wl[180] vdd gnd cell_6t
Xbit_r181_c59 bl[59] br[59] wl[181] vdd gnd cell_6t
Xbit_r182_c59 bl[59] br[59] wl[182] vdd gnd cell_6t
Xbit_r183_c59 bl[59] br[59] wl[183] vdd gnd cell_6t
Xbit_r184_c59 bl[59] br[59] wl[184] vdd gnd cell_6t
Xbit_r185_c59 bl[59] br[59] wl[185] vdd gnd cell_6t
Xbit_r186_c59 bl[59] br[59] wl[186] vdd gnd cell_6t
Xbit_r187_c59 bl[59] br[59] wl[187] vdd gnd cell_6t
Xbit_r188_c59 bl[59] br[59] wl[188] vdd gnd cell_6t
Xbit_r189_c59 bl[59] br[59] wl[189] vdd gnd cell_6t
Xbit_r190_c59 bl[59] br[59] wl[190] vdd gnd cell_6t
Xbit_r191_c59 bl[59] br[59] wl[191] vdd gnd cell_6t
Xbit_r192_c59 bl[59] br[59] wl[192] vdd gnd cell_6t
Xbit_r193_c59 bl[59] br[59] wl[193] vdd gnd cell_6t
Xbit_r194_c59 bl[59] br[59] wl[194] vdd gnd cell_6t
Xbit_r195_c59 bl[59] br[59] wl[195] vdd gnd cell_6t
Xbit_r196_c59 bl[59] br[59] wl[196] vdd gnd cell_6t
Xbit_r197_c59 bl[59] br[59] wl[197] vdd gnd cell_6t
Xbit_r198_c59 bl[59] br[59] wl[198] vdd gnd cell_6t
Xbit_r199_c59 bl[59] br[59] wl[199] vdd gnd cell_6t
Xbit_r200_c59 bl[59] br[59] wl[200] vdd gnd cell_6t
Xbit_r201_c59 bl[59] br[59] wl[201] vdd gnd cell_6t
Xbit_r202_c59 bl[59] br[59] wl[202] vdd gnd cell_6t
Xbit_r203_c59 bl[59] br[59] wl[203] vdd gnd cell_6t
Xbit_r204_c59 bl[59] br[59] wl[204] vdd gnd cell_6t
Xbit_r205_c59 bl[59] br[59] wl[205] vdd gnd cell_6t
Xbit_r206_c59 bl[59] br[59] wl[206] vdd gnd cell_6t
Xbit_r207_c59 bl[59] br[59] wl[207] vdd gnd cell_6t
Xbit_r208_c59 bl[59] br[59] wl[208] vdd gnd cell_6t
Xbit_r209_c59 bl[59] br[59] wl[209] vdd gnd cell_6t
Xbit_r210_c59 bl[59] br[59] wl[210] vdd gnd cell_6t
Xbit_r211_c59 bl[59] br[59] wl[211] vdd gnd cell_6t
Xbit_r212_c59 bl[59] br[59] wl[212] vdd gnd cell_6t
Xbit_r213_c59 bl[59] br[59] wl[213] vdd gnd cell_6t
Xbit_r214_c59 bl[59] br[59] wl[214] vdd gnd cell_6t
Xbit_r215_c59 bl[59] br[59] wl[215] vdd gnd cell_6t
Xbit_r216_c59 bl[59] br[59] wl[216] vdd gnd cell_6t
Xbit_r217_c59 bl[59] br[59] wl[217] vdd gnd cell_6t
Xbit_r218_c59 bl[59] br[59] wl[218] vdd gnd cell_6t
Xbit_r219_c59 bl[59] br[59] wl[219] vdd gnd cell_6t
Xbit_r220_c59 bl[59] br[59] wl[220] vdd gnd cell_6t
Xbit_r221_c59 bl[59] br[59] wl[221] vdd gnd cell_6t
Xbit_r222_c59 bl[59] br[59] wl[222] vdd gnd cell_6t
Xbit_r223_c59 bl[59] br[59] wl[223] vdd gnd cell_6t
Xbit_r224_c59 bl[59] br[59] wl[224] vdd gnd cell_6t
Xbit_r225_c59 bl[59] br[59] wl[225] vdd gnd cell_6t
Xbit_r226_c59 bl[59] br[59] wl[226] vdd gnd cell_6t
Xbit_r227_c59 bl[59] br[59] wl[227] vdd gnd cell_6t
Xbit_r228_c59 bl[59] br[59] wl[228] vdd gnd cell_6t
Xbit_r229_c59 bl[59] br[59] wl[229] vdd gnd cell_6t
Xbit_r230_c59 bl[59] br[59] wl[230] vdd gnd cell_6t
Xbit_r231_c59 bl[59] br[59] wl[231] vdd gnd cell_6t
Xbit_r232_c59 bl[59] br[59] wl[232] vdd gnd cell_6t
Xbit_r233_c59 bl[59] br[59] wl[233] vdd gnd cell_6t
Xbit_r234_c59 bl[59] br[59] wl[234] vdd gnd cell_6t
Xbit_r235_c59 bl[59] br[59] wl[235] vdd gnd cell_6t
Xbit_r236_c59 bl[59] br[59] wl[236] vdd gnd cell_6t
Xbit_r237_c59 bl[59] br[59] wl[237] vdd gnd cell_6t
Xbit_r238_c59 bl[59] br[59] wl[238] vdd gnd cell_6t
Xbit_r239_c59 bl[59] br[59] wl[239] vdd gnd cell_6t
Xbit_r240_c59 bl[59] br[59] wl[240] vdd gnd cell_6t
Xbit_r241_c59 bl[59] br[59] wl[241] vdd gnd cell_6t
Xbit_r242_c59 bl[59] br[59] wl[242] vdd gnd cell_6t
Xbit_r243_c59 bl[59] br[59] wl[243] vdd gnd cell_6t
Xbit_r244_c59 bl[59] br[59] wl[244] vdd gnd cell_6t
Xbit_r245_c59 bl[59] br[59] wl[245] vdd gnd cell_6t
Xbit_r246_c59 bl[59] br[59] wl[246] vdd gnd cell_6t
Xbit_r247_c59 bl[59] br[59] wl[247] vdd gnd cell_6t
Xbit_r248_c59 bl[59] br[59] wl[248] vdd gnd cell_6t
Xbit_r249_c59 bl[59] br[59] wl[249] vdd gnd cell_6t
Xbit_r250_c59 bl[59] br[59] wl[250] vdd gnd cell_6t
Xbit_r251_c59 bl[59] br[59] wl[251] vdd gnd cell_6t
Xbit_r252_c59 bl[59] br[59] wl[252] vdd gnd cell_6t
Xbit_r253_c59 bl[59] br[59] wl[253] vdd gnd cell_6t
Xbit_r254_c59 bl[59] br[59] wl[254] vdd gnd cell_6t
Xbit_r255_c59 bl[59] br[59] wl[255] vdd gnd cell_6t
Xbit_r0_c60 bl[60] br[60] wl[0] vdd gnd cell_6t
Xbit_r1_c60 bl[60] br[60] wl[1] vdd gnd cell_6t
Xbit_r2_c60 bl[60] br[60] wl[2] vdd gnd cell_6t
Xbit_r3_c60 bl[60] br[60] wl[3] vdd gnd cell_6t
Xbit_r4_c60 bl[60] br[60] wl[4] vdd gnd cell_6t
Xbit_r5_c60 bl[60] br[60] wl[5] vdd gnd cell_6t
Xbit_r6_c60 bl[60] br[60] wl[6] vdd gnd cell_6t
Xbit_r7_c60 bl[60] br[60] wl[7] vdd gnd cell_6t
Xbit_r8_c60 bl[60] br[60] wl[8] vdd gnd cell_6t
Xbit_r9_c60 bl[60] br[60] wl[9] vdd gnd cell_6t
Xbit_r10_c60 bl[60] br[60] wl[10] vdd gnd cell_6t
Xbit_r11_c60 bl[60] br[60] wl[11] vdd gnd cell_6t
Xbit_r12_c60 bl[60] br[60] wl[12] vdd gnd cell_6t
Xbit_r13_c60 bl[60] br[60] wl[13] vdd gnd cell_6t
Xbit_r14_c60 bl[60] br[60] wl[14] vdd gnd cell_6t
Xbit_r15_c60 bl[60] br[60] wl[15] vdd gnd cell_6t
Xbit_r16_c60 bl[60] br[60] wl[16] vdd gnd cell_6t
Xbit_r17_c60 bl[60] br[60] wl[17] vdd gnd cell_6t
Xbit_r18_c60 bl[60] br[60] wl[18] vdd gnd cell_6t
Xbit_r19_c60 bl[60] br[60] wl[19] vdd gnd cell_6t
Xbit_r20_c60 bl[60] br[60] wl[20] vdd gnd cell_6t
Xbit_r21_c60 bl[60] br[60] wl[21] vdd gnd cell_6t
Xbit_r22_c60 bl[60] br[60] wl[22] vdd gnd cell_6t
Xbit_r23_c60 bl[60] br[60] wl[23] vdd gnd cell_6t
Xbit_r24_c60 bl[60] br[60] wl[24] vdd gnd cell_6t
Xbit_r25_c60 bl[60] br[60] wl[25] vdd gnd cell_6t
Xbit_r26_c60 bl[60] br[60] wl[26] vdd gnd cell_6t
Xbit_r27_c60 bl[60] br[60] wl[27] vdd gnd cell_6t
Xbit_r28_c60 bl[60] br[60] wl[28] vdd gnd cell_6t
Xbit_r29_c60 bl[60] br[60] wl[29] vdd gnd cell_6t
Xbit_r30_c60 bl[60] br[60] wl[30] vdd gnd cell_6t
Xbit_r31_c60 bl[60] br[60] wl[31] vdd gnd cell_6t
Xbit_r32_c60 bl[60] br[60] wl[32] vdd gnd cell_6t
Xbit_r33_c60 bl[60] br[60] wl[33] vdd gnd cell_6t
Xbit_r34_c60 bl[60] br[60] wl[34] vdd gnd cell_6t
Xbit_r35_c60 bl[60] br[60] wl[35] vdd gnd cell_6t
Xbit_r36_c60 bl[60] br[60] wl[36] vdd gnd cell_6t
Xbit_r37_c60 bl[60] br[60] wl[37] vdd gnd cell_6t
Xbit_r38_c60 bl[60] br[60] wl[38] vdd gnd cell_6t
Xbit_r39_c60 bl[60] br[60] wl[39] vdd gnd cell_6t
Xbit_r40_c60 bl[60] br[60] wl[40] vdd gnd cell_6t
Xbit_r41_c60 bl[60] br[60] wl[41] vdd gnd cell_6t
Xbit_r42_c60 bl[60] br[60] wl[42] vdd gnd cell_6t
Xbit_r43_c60 bl[60] br[60] wl[43] vdd gnd cell_6t
Xbit_r44_c60 bl[60] br[60] wl[44] vdd gnd cell_6t
Xbit_r45_c60 bl[60] br[60] wl[45] vdd gnd cell_6t
Xbit_r46_c60 bl[60] br[60] wl[46] vdd gnd cell_6t
Xbit_r47_c60 bl[60] br[60] wl[47] vdd gnd cell_6t
Xbit_r48_c60 bl[60] br[60] wl[48] vdd gnd cell_6t
Xbit_r49_c60 bl[60] br[60] wl[49] vdd gnd cell_6t
Xbit_r50_c60 bl[60] br[60] wl[50] vdd gnd cell_6t
Xbit_r51_c60 bl[60] br[60] wl[51] vdd gnd cell_6t
Xbit_r52_c60 bl[60] br[60] wl[52] vdd gnd cell_6t
Xbit_r53_c60 bl[60] br[60] wl[53] vdd gnd cell_6t
Xbit_r54_c60 bl[60] br[60] wl[54] vdd gnd cell_6t
Xbit_r55_c60 bl[60] br[60] wl[55] vdd gnd cell_6t
Xbit_r56_c60 bl[60] br[60] wl[56] vdd gnd cell_6t
Xbit_r57_c60 bl[60] br[60] wl[57] vdd gnd cell_6t
Xbit_r58_c60 bl[60] br[60] wl[58] vdd gnd cell_6t
Xbit_r59_c60 bl[60] br[60] wl[59] vdd gnd cell_6t
Xbit_r60_c60 bl[60] br[60] wl[60] vdd gnd cell_6t
Xbit_r61_c60 bl[60] br[60] wl[61] vdd gnd cell_6t
Xbit_r62_c60 bl[60] br[60] wl[62] vdd gnd cell_6t
Xbit_r63_c60 bl[60] br[60] wl[63] vdd gnd cell_6t
Xbit_r64_c60 bl[60] br[60] wl[64] vdd gnd cell_6t
Xbit_r65_c60 bl[60] br[60] wl[65] vdd gnd cell_6t
Xbit_r66_c60 bl[60] br[60] wl[66] vdd gnd cell_6t
Xbit_r67_c60 bl[60] br[60] wl[67] vdd gnd cell_6t
Xbit_r68_c60 bl[60] br[60] wl[68] vdd gnd cell_6t
Xbit_r69_c60 bl[60] br[60] wl[69] vdd gnd cell_6t
Xbit_r70_c60 bl[60] br[60] wl[70] vdd gnd cell_6t
Xbit_r71_c60 bl[60] br[60] wl[71] vdd gnd cell_6t
Xbit_r72_c60 bl[60] br[60] wl[72] vdd gnd cell_6t
Xbit_r73_c60 bl[60] br[60] wl[73] vdd gnd cell_6t
Xbit_r74_c60 bl[60] br[60] wl[74] vdd gnd cell_6t
Xbit_r75_c60 bl[60] br[60] wl[75] vdd gnd cell_6t
Xbit_r76_c60 bl[60] br[60] wl[76] vdd gnd cell_6t
Xbit_r77_c60 bl[60] br[60] wl[77] vdd gnd cell_6t
Xbit_r78_c60 bl[60] br[60] wl[78] vdd gnd cell_6t
Xbit_r79_c60 bl[60] br[60] wl[79] vdd gnd cell_6t
Xbit_r80_c60 bl[60] br[60] wl[80] vdd gnd cell_6t
Xbit_r81_c60 bl[60] br[60] wl[81] vdd gnd cell_6t
Xbit_r82_c60 bl[60] br[60] wl[82] vdd gnd cell_6t
Xbit_r83_c60 bl[60] br[60] wl[83] vdd gnd cell_6t
Xbit_r84_c60 bl[60] br[60] wl[84] vdd gnd cell_6t
Xbit_r85_c60 bl[60] br[60] wl[85] vdd gnd cell_6t
Xbit_r86_c60 bl[60] br[60] wl[86] vdd gnd cell_6t
Xbit_r87_c60 bl[60] br[60] wl[87] vdd gnd cell_6t
Xbit_r88_c60 bl[60] br[60] wl[88] vdd gnd cell_6t
Xbit_r89_c60 bl[60] br[60] wl[89] vdd gnd cell_6t
Xbit_r90_c60 bl[60] br[60] wl[90] vdd gnd cell_6t
Xbit_r91_c60 bl[60] br[60] wl[91] vdd gnd cell_6t
Xbit_r92_c60 bl[60] br[60] wl[92] vdd gnd cell_6t
Xbit_r93_c60 bl[60] br[60] wl[93] vdd gnd cell_6t
Xbit_r94_c60 bl[60] br[60] wl[94] vdd gnd cell_6t
Xbit_r95_c60 bl[60] br[60] wl[95] vdd gnd cell_6t
Xbit_r96_c60 bl[60] br[60] wl[96] vdd gnd cell_6t
Xbit_r97_c60 bl[60] br[60] wl[97] vdd gnd cell_6t
Xbit_r98_c60 bl[60] br[60] wl[98] vdd gnd cell_6t
Xbit_r99_c60 bl[60] br[60] wl[99] vdd gnd cell_6t
Xbit_r100_c60 bl[60] br[60] wl[100] vdd gnd cell_6t
Xbit_r101_c60 bl[60] br[60] wl[101] vdd gnd cell_6t
Xbit_r102_c60 bl[60] br[60] wl[102] vdd gnd cell_6t
Xbit_r103_c60 bl[60] br[60] wl[103] vdd gnd cell_6t
Xbit_r104_c60 bl[60] br[60] wl[104] vdd gnd cell_6t
Xbit_r105_c60 bl[60] br[60] wl[105] vdd gnd cell_6t
Xbit_r106_c60 bl[60] br[60] wl[106] vdd gnd cell_6t
Xbit_r107_c60 bl[60] br[60] wl[107] vdd gnd cell_6t
Xbit_r108_c60 bl[60] br[60] wl[108] vdd gnd cell_6t
Xbit_r109_c60 bl[60] br[60] wl[109] vdd gnd cell_6t
Xbit_r110_c60 bl[60] br[60] wl[110] vdd gnd cell_6t
Xbit_r111_c60 bl[60] br[60] wl[111] vdd gnd cell_6t
Xbit_r112_c60 bl[60] br[60] wl[112] vdd gnd cell_6t
Xbit_r113_c60 bl[60] br[60] wl[113] vdd gnd cell_6t
Xbit_r114_c60 bl[60] br[60] wl[114] vdd gnd cell_6t
Xbit_r115_c60 bl[60] br[60] wl[115] vdd gnd cell_6t
Xbit_r116_c60 bl[60] br[60] wl[116] vdd gnd cell_6t
Xbit_r117_c60 bl[60] br[60] wl[117] vdd gnd cell_6t
Xbit_r118_c60 bl[60] br[60] wl[118] vdd gnd cell_6t
Xbit_r119_c60 bl[60] br[60] wl[119] vdd gnd cell_6t
Xbit_r120_c60 bl[60] br[60] wl[120] vdd gnd cell_6t
Xbit_r121_c60 bl[60] br[60] wl[121] vdd gnd cell_6t
Xbit_r122_c60 bl[60] br[60] wl[122] vdd gnd cell_6t
Xbit_r123_c60 bl[60] br[60] wl[123] vdd gnd cell_6t
Xbit_r124_c60 bl[60] br[60] wl[124] vdd gnd cell_6t
Xbit_r125_c60 bl[60] br[60] wl[125] vdd gnd cell_6t
Xbit_r126_c60 bl[60] br[60] wl[126] vdd gnd cell_6t
Xbit_r127_c60 bl[60] br[60] wl[127] vdd gnd cell_6t
Xbit_r128_c60 bl[60] br[60] wl[128] vdd gnd cell_6t
Xbit_r129_c60 bl[60] br[60] wl[129] vdd gnd cell_6t
Xbit_r130_c60 bl[60] br[60] wl[130] vdd gnd cell_6t
Xbit_r131_c60 bl[60] br[60] wl[131] vdd gnd cell_6t
Xbit_r132_c60 bl[60] br[60] wl[132] vdd gnd cell_6t
Xbit_r133_c60 bl[60] br[60] wl[133] vdd gnd cell_6t
Xbit_r134_c60 bl[60] br[60] wl[134] vdd gnd cell_6t
Xbit_r135_c60 bl[60] br[60] wl[135] vdd gnd cell_6t
Xbit_r136_c60 bl[60] br[60] wl[136] vdd gnd cell_6t
Xbit_r137_c60 bl[60] br[60] wl[137] vdd gnd cell_6t
Xbit_r138_c60 bl[60] br[60] wl[138] vdd gnd cell_6t
Xbit_r139_c60 bl[60] br[60] wl[139] vdd gnd cell_6t
Xbit_r140_c60 bl[60] br[60] wl[140] vdd gnd cell_6t
Xbit_r141_c60 bl[60] br[60] wl[141] vdd gnd cell_6t
Xbit_r142_c60 bl[60] br[60] wl[142] vdd gnd cell_6t
Xbit_r143_c60 bl[60] br[60] wl[143] vdd gnd cell_6t
Xbit_r144_c60 bl[60] br[60] wl[144] vdd gnd cell_6t
Xbit_r145_c60 bl[60] br[60] wl[145] vdd gnd cell_6t
Xbit_r146_c60 bl[60] br[60] wl[146] vdd gnd cell_6t
Xbit_r147_c60 bl[60] br[60] wl[147] vdd gnd cell_6t
Xbit_r148_c60 bl[60] br[60] wl[148] vdd gnd cell_6t
Xbit_r149_c60 bl[60] br[60] wl[149] vdd gnd cell_6t
Xbit_r150_c60 bl[60] br[60] wl[150] vdd gnd cell_6t
Xbit_r151_c60 bl[60] br[60] wl[151] vdd gnd cell_6t
Xbit_r152_c60 bl[60] br[60] wl[152] vdd gnd cell_6t
Xbit_r153_c60 bl[60] br[60] wl[153] vdd gnd cell_6t
Xbit_r154_c60 bl[60] br[60] wl[154] vdd gnd cell_6t
Xbit_r155_c60 bl[60] br[60] wl[155] vdd gnd cell_6t
Xbit_r156_c60 bl[60] br[60] wl[156] vdd gnd cell_6t
Xbit_r157_c60 bl[60] br[60] wl[157] vdd gnd cell_6t
Xbit_r158_c60 bl[60] br[60] wl[158] vdd gnd cell_6t
Xbit_r159_c60 bl[60] br[60] wl[159] vdd gnd cell_6t
Xbit_r160_c60 bl[60] br[60] wl[160] vdd gnd cell_6t
Xbit_r161_c60 bl[60] br[60] wl[161] vdd gnd cell_6t
Xbit_r162_c60 bl[60] br[60] wl[162] vdd gnd cell_6t
Xbit_r163_c60 bl[60] br[60] wl[163] vdd gnd cell_6t
Xbit_r164_c60 bl[60] br[60] wl[164] vdd gnd cell_6t
Xbit_r165_c60 bl[60] br[60] wl[165] vdd gnd cell_6t
Xbit_r166_c60 bl[60] br[60] wl[166] vdd gnd cell_6t
Xbit_r167_c60 bl[60] br[60] wl[167] vdd gnd cell_6t
Xbit_r168_c60 bl[60] br[60] wl[168] vdd gnd cell_6t
Xbit_r169_c60 bl[60] br[60] wl[169] vdd gnd cell_6t
Xbit_r170_c60 bl[60] br[60] wl[170] vdd gnd cell_6t
Xbit_r171_c60 bl[60] br[60] wl[171] vdd gnd cell_6t
Xbit_r172_c60 bl[60] br[60] wl[172] vdd gnd cell_6t
Xbit_r173_c60 bl[60] br[60] wl[173] vdd gnd cell_6t
Xbit_r174_c60 bl[60] br[60] wl[174] vdd gnd cell_6t
Xbit_r175_c60 bl[60] br[60] wl[175] vdd gnd cell_6t
Xbit_r176_c60 bl[60] br[60] wl[176] vdd gnd cell_6t
Xbit_r177_c60 bl[60] br[60] wl[177] vdd gnd cell_6t
Xbit_r178_c60 bl[60] br[60] wl[178] vdd gnd cell_6t
Xbit_r179_c60 bl[60] br[60] wl[179] vdd gnd cell_6t
Xbit_r180_c60 bl[60] br[60] wl[180] vdd gnd cell_6t
Xbit_r181_c60 bl[60] br[60] wl[181] vdd gnd cell_6t
Xbit_r182_c60 bl[60] br[60] wl[182] vdd gnd cell_6t
Xbit_r183_c60 bl[60] br[60] wl[183] vdd gnd cell_6t
Xbit_r184_c60 bl[60] br[60] wl[184] vdd gnd cell_6t
Xbit_r185_c60 bl[60] br[60] wl[185] vdd gnd cell_6t
Xbit_r186_c60 bl[60] br[60] wl[186] vdd gnd cell_6t
Xbit_r187_c60 bl[60] br[60] wl[187] vdd gnd cell_6t
Xbit_r188_c60 bl[60] br[60] wl[188] vdd gnd cell_6t
Xbit_r189_c60 bl[60] br[60] wl[189] vdd gnd cell_6t
Xbit_r190_c60 bl[60] br[60] wl[190] vdd gnd cell_6t
Xbit_r191_c60 bl[60] br[60] wl[191] vdd gnd cell_6t
Xbit_r192_c60 bl[60] br[60] wl[192] vdd gnd cell_6t
Xbit_r193_c60 bl[60] br[60] wl[193] vdd gnd cell_6t
Xbit_r194_c60 bl[60] br[60] wl[194] vdd gnd cell_6t
Xbit_r195_c60 bl[60] br[60] wl[195] vdd gnd cell_6t
Xbit_r196_c60 bl[60] br[60] wl[196] vdd gnd cell_6t
Xbit_r197_c60 bl[60] br[60] wl[197] vdd gnd cell_6t
Xbit_r198_c60 bl[60] br[60] wl[198] vdd gnd cell_6t
Xbit_r199_c60 bl[60] br[60] wl[199] vdd gnd cell_6t
Xbit_r200_c60 bl[60] br[60] wl[200] vdd gnd cell_6t
Xbit_r201_c60 bl[60] br[60] wl[201] vdd gnd cell_6t
Xbit_r202_c60 bl[60] br[60] wl[202] vdd gnd cell_6t
Xbit_r203_c60 bl[60] br[60] wl[203] vdd gnd cell_6t
Xbit_r204_c60 bl[60] br[60] wl[204] vdd gnd cell_6t
Xbit_r205_c60 bl[60] br[60] wl[205] vdd gnd cell_6t
Xbit_r206_c60 bl[60] br[60] wl[206] vdd gnd cell_6t
Xbit_r207_c60 bl[60] br[60] wl[207] vdd gnd cell_6t
Xbit_r208_c60 bl[60] br[60] wl[208] vdd gnd cell_6t
Xbit_r209_c60 bl[60] br[60] wl[209] vdd gnd cell_6t
Xbit_r210_c60 bl[60] br[60] wl[210] vdd gnd cell_6t
Xbit_r211_c60 bl[60] br[60] wl[211] vdd gnd cell_6t
Xbit_r212_c60 bl[60] br[60] wl[212] vdd gnd cell_6t
Xbit_r213_c60 bl[60] br[60] wl[213] vdd gnd cell_6t
Xbit_r214_c60 bl[60] br[60] wl[214] vdd gnd cell_6t
Xbit_r215_c60 bl[60] br[60] wl[215] vdd gnd cell_6t
Xbit_r216_c60 bl[60] br[60] wl[216] vdd gnd cell_6t
Xbit_r217_c60 bl[60] br[60] wl[217] vdd gnd cell_6t
Xbit_r218_c60 bl[60] br[60] wl[218] vdd gnd cell_6t
Xbit_r219_c60 bl[60] br[60] wl[219] vdd gnd cell_6t
Xbit_r220_c60 bl[60] br[60] wl[220] vdd gnd cell_6t
Xbit_r221_c60 bl[60] br[60] wl[221] vdd gnd cell_6t
Xbit_r222_c60 bl[60] br[60] wl[222] vdd gnd cell_6t
Xbit_r223_c60 bl[60] br[60] wl[223] vdd gnd cell_6t
Xbit_r224_c60 bl[60] br[60] wl[224] vdd gnd cell_6t
Xbit_r225_c60 bl[60] br[60] wl[225] vdd gnd cell_6t
Xbit_r226_c60 bl[60] br[60] wl[226] vdd gnd cell_6t
Xbit_r227_c60 bl[60] br[60] wl[227] vdd gnd cell_6t
Xbit_r228_c60 bl[60] br[60] wl[228] vdd gnd cell_6t
Xbit_r229_c60 bl[60] br[60] wl[229] vdd gnd cell_6t
Xbit_r230_c60 bl[60] br[60] wl[230] vdd gnd cell_6t
Xbit_r231_c60 bl[60] br[60] wl[231] vdd gnd cell_6t
Xbit_r232_c60 bl[60] br[60] wl[232] vdd gnd cell_6t
Xbit_r233_c60 bl[60] br[60] wl[233] vdd gnd cell_6t
Xbit_r234_c60 bl[60] br[60] wl[234] vdd gnd cell_6t
Xbit_r235_c60 bl[60] br[60] wl[235] vdd gnd cell_6t
Xbit_r236_c60 bl[60] br[60] wl[236] vdd gnd cell_6t
Xbit_r237_c60 bl[60] br[60] wl[237] vdd gnd cell_6t
Xbit_r238_c60 bl[60] br[60] wl[238] vdd gnd cell_6t
Xbit_r239_c60 bl[60] br[60] wl[239] vdd gnd cell_6t
Xbit_r240_c60 bl[60] br[60] wl[240] vdd gnd cell_6t
Xbit_r241_c60 bl[60] br[60] wl[241] vdd gnd cell_6t
Xbit_r242_c60 bl[60] br[60] wl[242] vdd gnd cell_6t
Xbit_r243_c60 bl[60] br[60] wl[243] vdd gnd cell_6t
Xbit_r244_c60 bl[60] br[60] wl[244] vdd gnd cell_6t
Xbit_r245_c60 bl[60] br[60] wl[245] vdd gnd cell_6t
Xbit_r246_c60 bl[60] br[60] wl[246] vdd gnd cell_6t
Xbit_r247_c60 bl[60] br[60] wl[247] vdd gnd cell_6t
Xbit_r248_c60 bl[60] br[60] wl[248] vdd gnd cell_6t
Xbit_r249_c60 bl[60] br[60] wl[249] vdd gnd cell_6t
Xbit_r250_c60 bl[60] br[60] wl[250] vdd gnd cell_6t
Xbit_r251_c60 bl[60] br[60] wl[251] vdd gnd cell_6t
Xbit_r252_c60 bl[60] br[60] wl[252] vdd gnd cell_6t
Xbit_r253_c60 bl[60] br[60] wl[253] vdd gnd cell_6t
Xbit_r254_c60 bl[60] br[60] wl[254] vdd gnd cell_6t
Xbit_r255_c60 bl[60] br[60] wl[255] vdd gnd cell_6t
Xbit_r0_c61 bl[61] br[61] wl[0] vdd gnd cell_6t
Xbit_r1_c61 bl[61] br[61] wl[1] vdd gnd cell_6t
Xbit_r2_c61 bl[61] br[61] wl[2] vdd gnd cell_6t
Xbit_r3_c61 bl[61] br[61] wl[3] vdd gnd cell_6t
Xbit_r4_c61 bl[61] br[61] wl[4] vdd gnd cell_6t
Xbit_r5_c61 bl[61] br[61] wl[5] vdd gnd cell_6t
Xbit_r6_c61 bl[61] br[61] wl[6] vdd gnd cell_6t
Xbit_r7_c61 bl[61] br[61] wl[7] vdd gnd cell_6t
Xbit_r8_c61 bl[61] br[61] wl[8] vdd gnd cell_6t
Xbit_r9_c61 bl[61] br[61] wl[9] vdd gnd cell_6t
Xbit_r10_c61 bl[61] br[61] wl[10] vdd gnd cell_6t
Xbit_r11_c61 bl[61] br[61] wl[11] vdd gnd cell_6t
Xbit_r12_c61 bl[61] br[61] wl[12] vdd gnd cell_6t
Xbit_r13_c61 bl[61] br[61] wl[13] vdd gnd cell_6t
Xbit_r14_c61 bl[61] br[61] wl[14] vdd gnd cell_6t
Xbit_r15_c61 bl[61] br[61] wl[15] vdd gnd cell_6t
Xbit_r16_c61 bl[61] br[61] wl[16] vdd gnd cell_6t
Xbit_r17_c61 bl[61] br[61] wl[17] vdd gnd cell_6t
Xbit_r18_c61 bl[61] br[61] wl[18] vdd gnd cell_6t
Xbit_r19_c61 bl[61] br[61] wl[19] vdd gnd cell_6t
Xbit_r20_c61 bl[61] br[61] wl[20] vdd gnd cell_6t
Xbit_r21_c61 bl[61] br[61] wl[21] vdd gnd cell_6t
Xbit_r22_c61 bl[61] br[61] wl[22] vdd gnd cell_6t
Xbit_r23_c61 bl[61] br[61] wl[23] vdd gnd cell_6t
Xbit_r24_c61 bl[61] br[61] wl[24] vdd gnd cell_6t
Xbit_r25_c61 bl[61] br[61] wl[25] vdd gnd cell_6t
Xbit_r26_c61 bl[61] br[61] wl[26] vdd gnd cell_6t
Xbit_r27_c61 bl[61] br[61] wl[27] vdd gnd cell_6t
Xbit_r28_c61 bl[61] br[61] wl[28] vdd gnd cell_6t
Xbit_r29_c61 bl[61] br[61] wl[29] vdd gnd cell_6t
Xbit_r30_c61 bl[61] br[61] wl[30] vdd gnd cell_6t
Xbit_r31_c61 bl[61] br[61] wl[31] vdd gnd cell_6t
Xbit_r32_c61 bl[61] br[61] wl[32] vdd gnd cell_6t
Xbit_r33_c61 bl[61] br[61] wl[33] vdd gnd cell_6t
Xbit_r34_c61 bl[61] br[61] wl[34] vdd gnd cell_6t
Xbit_r35_c61 bl[61] br[61] wl[35] vdd gnd cell_6t
Xbit_r36_c61 bl[61] br[61] wl[36] vdd gnd cell_6t
Xbit_r37_c61 bl[61] br[61] wl[37] vdd gnd cell_6t
Xbit_r38_c61 bl[61] br[61] wl[38] vdd gnd cell_6t
Xbit_r39_c61 bl[61] br[61] wl[39] vdd gnd cell_6t
Xbit_r40_c61 bl[61] br[61] wl[40] vdd gnd cell_6t
Xbit_r41_c61 bl[61] br[61] wl[41] vdd gnd cell_6t
Xbit_r42_c61 bl[61] br[61] wl[42] vdd gnd cell_6t
Xbit_r43_c61 bl[61] br[61] wl[43] vdd gnd cell_6t
Xbit_r44_c61 bl[61] br[61] wl[44] vdd gnd cell_6t
Xbit_r45_c61 bl[61] br[61] wl[45] vdd gnd cell_6t
Xbit_r46_c61 bl[61] br[61] wl[46] vdd gnd cell_6t
Xbit_r47_c61 bl[61] br[61] wl[47] vdd gnd cell_6t
Xbit_r48_c61 bl[61] br[61] wl[48] vdd gnd cell_6t
Xbit_r49_c61 bl[61] br[61] wl[49] vdd gnd cell_6t
Xbit_r50_c61 bl[61] br[61] wl[50] vdd gnd cell_6t
Xbit_r51_c61 bl[61] br[61] wl[51] vdd gnd cell_6t
Xbit_r52_c61 bl[61] br[61] wl[52] vdd gnd cell_6t
Xbit_r53_c61 bl[61] br[61] wl[53] vdd gnd cell_6t
Xbit_r54_c61 bl[61] br[61] wl[54] vdd gnd cell_6t
Xbit_r55_c61 bl[61] br[61] wl[55] vdd gnd cell_6t
Xbit_r56_c61 bl[61] br[61] wl[56] vdd gnd cell_6t
Xbit_r57_c61 bl[61] br[61] wl[57] vdd gnd cell_6t
Xbit_r58_c61 bl[61] br[61] wl[58] vdd gnd cell_6t
Xbit_r59_c61 bl[61] br[61] wl[59] vdd gnd cell_6t
Xbit_r60_c61 bl[61] br[61] wl[60] vdd gnd cell_6t
Xbit_r61_c61 bl[61] br[61] wl[61] vdd gnd cell_6t
Xbit_r62_c61 bl[61] br[61] wl[62] vdd gnd cell_6t
Xbit_r63_c61 bl[61] br[61] wl[63] vdd gnd cell_6t
Xbit_r64_c61 bl[61] br[61] wl[64] vdd gnd cell_6t
Xbit_r65_c61 bl[61] br[61] wl[65] vdd gnd cell_6t
Xbit_r66_c61 bl[61] br[61] wl[66] vdd gnd cell_6t
Xbit_r67_c61 bl[61] br[61] wl[67] vdd gnd cell_6t
Xbit_r68_c61 bl[61] br[61] wl[68] vdd gnd cell_6t
Xbit_r69_c61 bl[61] br[61] wl[69] vdd gnd cell_6t
Xbit_r70_c61 bl[61] br[61] wl[70] vdd gnd cell_6t
Xbit_r71_c61 bl[61] br[61] wl[71] vdd gnd cell_6t
Xbit_r72_c61 bl[61] br[61] wl[72] vdd gnd cell_6t
Xbit_r73_c61 bl[61] br[61] wl[73] vdd gnd cell_6t
Xbit_r74_c61 bl[61] br[61] wl[74] vdd gnd cell_6t
Xbit_r75_c61 bl[61] br[61] wl[75] vdd gnd cell_6t
Xbit_r76_c61 bl[61] br[61] wl[76] vdd gnd cell_6t
Xbit_r77_c61 bl[61] br[61] wl[77] vdd gnd cell_6t
Xbit_r78_c61 bl[61] br[61] wl[78] vdd gnd cell_6t
Xbit_r79_c61 bl[61] br[61] wl[79] vdd gnd cell_6t
Xbit_r80_c61 bl[61] br[61] wl[80] vdd gnd cell_6t
Xbit_r81_c61 bl[61] br[61] wl[81] vdd gnd cell_6t
Xbit_r82_c61 bl[61] br[61] wl[82] vdd gnd cell_6t
Xbit_r83_c61 bl[61] br[61] wl[83] vdd gnd cell_6t
Xbit_r84_c61 bl[61] br[61] wl[84] vdd gnd cell_6t
Xbit_r85_c61 bl[61] br[61] wl[85] vdd gnd cell_6t
Xbit_r86_c61 bl[61] br[61] wl[86] vdd gnd cell_6t
Xbit_r87_c61 bl[61] br[61] wl[87] vdd gnd cell_6t
Xbit_r88_c61 bl[61] br[61] wl[88] vdd gnd cell_6t
Xbit_r89_c61 bl[61] br[61] wl[89] vdd gnd cell_6t
Xbit_r90_c61 bl[61] br[61] wl[90] vdd gnd cell_6t
Xbit_r91_c61 bl[61] br[61] wl[91] vdd gnd cell_6t
Xbit_r92_c61 bl[61] br[61] wl[92] vdd gnd cell_6t
Xbit_r93_c61 bl[61] br[61] wl[93] vdd gnd cell_6t
Xbit_r94_c61 bl[61] br[61] wl[94] vdd gnd cell_6t
Xbit_r95_c61 bl[61] br[61] wl[95] vdd gnd cell_6t
Xbit_r96_c61 bl[61] br[61] wl[96] vdd gnd cell_6t
Xbit_r97_c61 bl[61] br[61] wl[97] vdd gnd cell_6t
Xbit_r98_c61 bl[61] br[61] wl[98] vdd gnd cell_6t
Xbit_r99_c61 bl[61] br[61] wl[99] vdd gnd cell_6t
Xbit_r100_c61 bl[61] br[61] wl[100] vdd gnd cell_6t
Xbit_r101_c61 bl[61] br[61] wl[101] vdd gnd cell_6t
Xbit_r102_c61 bl[61] br[61] wl[102] vdd gnd cell_6t
Xbit_r103_c61 bl[61] br[61] wl[103] vdd gnd cell_6t
Xbit_r104_c61 bl[61] br[61] wl[104] vdd gnd cell_6t
Xbit_r105_c61 bl[61] br[61] wl[105] vdd gnd cell_6t
Xbit_r106_c61 bl[61] br[61] wl[106] vdd gnd cell_6t
Xbit_r107_c61 bl[61] br[61] wl[107] vdd gnd cell_6t
Xbit_r108_c61 bl[61] br[61] wl[108] vdd gnd cell_6t
Xbit_r109_c61 bl[61] br[61] wl[109] vdd gnd cell_6t
Xbit_r110_c61 bl[61] br[61] wl[110] vdd gnd cell_6t
Xbit_r111_c61 bl[61] br[61] wl[111] vdd gnd cell_6t
Xbit_r112_c61 bl[61] br[61] wl[112] vdd gnd cell_6t
Xbit_r113_c61 bl[61] br[61] wl[113] vdd gnd cell_6t
Xbit_r114_c61 bl[61] br[61] wl[114] vdd gnd cell_6t
Xbit_r115_c61 bl[61] br[61] wl[115] vdd gnd cell_6t
Xbit_r116_c61 bl[61] br[61] wl[116] vdd gnd cell_6t
Xbit_r117_c61 bl[61] br[61] wl[117] vdd gnd cell_6t
Xbit_r118_c61 bl[61] br[61] wl[118] vdd gnd cell_6t
Xbit_r119_c61 bl[61] br[61] wl[119] vdd gnd cell_6t
Xbit_r120_c61 bl[61] br[61] wl[120] vdd gnd cell_6t
Xbit_r121_c61 bl[61] br[61] wl[121] vdd gnd cell_6t
Xbit_r122_c61 bl[61] br[61] wl[122] vdd gnd cell_6t
Xbit_r123_c61 bl[61] br[61] wl[123] vdd gnd cell_6t
Xbit_r124_c61 bl[61] br[61] wl[124] vdd gnd cell_6t
Xbit_r125_c61 bl[61] br[61] wl[125] vdd gnd cell_6t
Xbit_r126_c61 bl[61] br[61] wl[126] vdd gnd cell_6t
Xbit_r127_c61 bl[61] br[61] wl[127] vdd gnd cell_6t
Xbit_r128_c61 bl[61] br[61] wl[128] vdd gnd cell_6t
Xbit_r129_c61 bl[61] br[61] wl[129] vdd gnd cell_6t
Xbit_r130_c61 bl[61] br[61] wl[130] vdd gnd cell_6t
Xbit_r131_c61 bl[61] br[61] wl[131] vdd gnd cell_6t
Xbit_r132_c61 bl[61] br[61] wl[132] vdd gnd cell_6t
Xbit_r133_c61 bl[61] br[61] wl[133] vdd gnd cell_6t
Xbit_r134_c61 bl[61] br[61] wl[134] vdd gnd cell_6t
Xbit_r135_c61 bl[61] br[61] wl[135] vdd gnd cell_6t
Xbit_r136_c61 bl[61] br[61] wl[136] vdd gnd cell_6t
Xbit_r137_c61 bl[61] br[61] wl[137] vdd gnd cell_6t
Xbit_r138_c61 bl[61] br[61] wl[138] vdd gnd cell_6t
Xbit_r139_c61 bl[61] br[61] wl[139] vdd gnd cell_6t
Xbit_r140_c61 bl[61] br[61] wl[140] vdd gnd cell_6t
Xbit_r141_c61 bl[61] br[61] wl[141] vdd gnd cell_6t
Xbit_r142_c61 bl[61] br[61] wl[142] vdd gnd cell_6t
Xbit_r143_c61 bl[61] br[61] wl[143] vdd gnd cell_6t
Xbit_r144_c61 bl[61] br[61] wl[144] vdd gnd cell_6t
Xbit_r145_c61 bl[61] br[61] wl[145] vdd gnd cell_6t
Xbit_r146_c61 bl[61] br[61] wl[146] vdd gnd cell_6t
Xbit_r147_c61 bl[61] br[61] wl[147] vdd gnd cell_6t
Xbit_r148_c61 bl[61] br[61] wl[148] vdd gnd cell_6t
Xbit_r149_c61 bl[61] br[61] wl[149] vdd gnd cell_6t
Xbit_r150_c61 bl[61] br[61] wl[150] vdd gnd cell_6t
Xbit_r151_c61 bl[61] br[61] wl[151] vdd gnd cell_6t
Xbit_r152_c61 bl[61] br[61] wl[152] vdd gnd cell_6t
Xbit_r153_c61 bl[61] br[61] wl[153] vdd gnd cell_6t
Xbit_r154_c61 bl[61] br[61] wl[154] vdd gnd cell_6t
Xbit_r155_c61 bl[61] br[61] wl[155] vdd gnd cell_6t
Xbit_r156_c61 bl[61] br[61] wl[156] vdd gnd cell_6t
Xbit_r157_c61 bl[61] br[61] wl[157] vdd gnd cell_6t
Xbit_r158_c61 bl[61] br[61] wl[158] vdd gnd cell_6t
Xbit_r159_c61 bl[61] br[61] wl[159] vdd gnd cell_6t
Xbit_r160_c61 bl[61] br[61] wl[160] vdd gnd cell_6t
Xbit_r161_c61 bl[61] br[61] wl[161] vdd gnd cell_6t
Xbit_r162_c61 bl[61] br[61] wl[162] vdd gnd cell_6t
Xbit_r163_c61 bl[61] br[61] wl[163] vdd gnd cell_6t
Xbit_r164_c61 bl[61] br[61] wl[164] vdd gnd cell_6t
Xbit_r165_c61 bl[61] br[61] wl[165] vdd gnd cell_6t
Xbit_r166_c61 bl[61] br[61] wl[166] vdd gnd cell_6t
Xbit_r167_c61 bl[61] br[61] wl[167] vdd gnd cell_6t
Xbit_r168_c61 bl[61] br[61] wl[168] vdd gnd cell_6t
Xbit_r169_c61 bl[61] br[61] wl[169] vdd gnd cell_6t
Xbit_r170_c61 bl[61] br[61] wl[170] vdd gnd cell_6t
Xbit_r171_c61 bl[61] br[61] wl[171] vdd gnd cell_6t
Xbit_r172_c61 bl[61] br[61] wl[172] vdd gnd cell_6t
Xbit_r173_c61 bl[61] br[61] wl[173] vdd gnd cell_6t
Xbit_r174_c61 bl[61] br[61] wl[174] vdd gnd cell_6t
Xbit_r175_c61 bl[61] br[61] wl[175] vdd gnd cell_6t
Xbit_r176_c61 bl[61] br[61] wl[176] vdd gnd cell_6t
Xbit_r177_c61 bl[61] br[61] wl[177] vdd gnd cell_6t
Xbit_r178_c61 bl[61] br[61] wl[178] vdd gnd cell_6t
Xbit_r179_c61 bl[61] br[61] wl[179] vdd gnd cell_6t
Xbit_r180_c61 bl[61] br[61] wl[180] vdd gnd cell_6t
Xbit_r181_c61 bl[61] br[61] wl[181] vdd gnd cell_6t
Xbit_r182_c61 bl[61] br[61] wl[182] vdd gnd cell_6t
Xbit_r183_c61 bl[61] br[61] wl[183] vdd gnd cell_6t
Xbit_r184_c61 bl[61] br[61] wl[184] vdd gnd cell_6t
Xbit_r185_c61 bl[61] br[61] wl[185] vdd gnd cell_6t
Xbit_r186_c61 bl[61] br[61] wl[186] vdd gnd cell_6t
Xbit_r187_c61 bl[61] br[61] wl[187] vdd gnd cell_6t
Xbit_r188_c61 bl[61] br[61] wl[188] vdd gnd cell_6t
Xbit_r189_c61 bl[61] br[61] wl[189] vdd gnd cell_6t
Xbit_r190_c61 bl[61] br[61] wl[190] vdd gnd cell_6t
Xbit_r191_c61 bl[61] br[61] wl[191] vdd gnd cell_6t
Xbit_r192_c61 bl[61] br[61] wl[192] vdd gnd cell_6t
Xbit_r193_c61 bl[61] br[61] wl[193] vdd gnd cell_6t
Xbit_r194_c61 bl[61] br[61] wl[194] vdd gnd cell_6t
Xbit_r195_c61 bl[61] br[61] wl[195] vdd gnd cell_6t
Xbit_r196_c61 bl[61] br[61] wl[196] vdd gnd cell_6t
Xbit_r197_c61 bl[61] br[61] wl[197] vdd gnd cell_6t
Xbit_r198_c61 bl[61] br[61] wl[198] vdd gnd cell_6t
Xbit_r199_c61 bl[61] br[61] wl[199] vdd gnd cell_6t
Xbit_r200_c61 bl[61] br[61] wl[200] vdd gnd cell_6t
Xbit_r201_c61 bl[61] br[61] wl[201] vdd gnd cell_6t
Xbit_r202_c61 bl[61] br[61] wl[202] vdd gnd cell_6t
Xbit_r203_c61 bl[61] br[61] wl[203] vdd gnd cell_6t
Xbit_r204_c61 bl[61] br[61] wl[204] vdd gnd cell_6t
Xbit_r205_c61 bl[61] br[61] wl[205] vdd gnd cell_6t
Xbit_r206_c61 bl[61] br[61] wl[206] vdd gnd cell_6t
Xbit_r207_c61 bl[61] br[61] wl[207] vdd gnd cell_6t
Xbit_r208_c61 bl[61] br[61] wl[208] vdd gnd cell_6t
Xbit_r209_c61 bl[61] br[61] wl[209] vdd gnd cell_6t
Xbit_r210_c61 bl[61] br[61] wl[210] vdd gnd cell_6t
Xbit_r211_c61 bl[61] br[61] wl[211] vdd gnd cell_6t
Xbit_r212_c61 bl[61] br[61] wl[212] vdd gnd cell_6t
Xbit_r213_c61 bl[61] br[61] wl[213] vdd gnd cell_6t
Xbit_r214_c61 bl[61] br[61] wl[214] vdd gnd cell_6t
Xbit_r215_c61 bl[61] br[61] wl[215] vdd gnd cell_6t
Xbit_r216_c61 bl[61] br[61] wl[216] vdd gnd cell_6t
Xbit_r217_c61 bl[61] br[61] wl[217] vdd gnd cell_6t
Xbit_r218_c61 bl[61] br[61] wl[218] vdd gnd cell_6t
Xbit_r219_c61 bl[61] br[61] wl[219] vdd gnd cell_6t
Xbit_r220_c61 bl[61] br[61] wl[220] vdd gnd cell_6t
Xbit_r221_c61 bl[61] br[61] wl[221] vdd gnd cell_6t
Xbit_r222_c61 bl[61] br[61] wl[222] vdd gnd cell_6t
Xbit_r223_c61 bl[61] br[61] wl[223] vdd gnd cell_6t
Xbit_r224_c61 bl[61] br[61] wl[224] vdd gnd cell_6t
Xbit_r225_c61 bl[61] br[61] wl[225] vdd gnd cell_6t
Xbit_r226_c61 bl[61] br[61] wl[226] vdd gnd cell_6t
Xbit_r227_c61 bl[61] br[61] wl[227] vdd gnd cell_6t
Xbit_r228_c61 bl[61] br[61] wl[228] vdd gnd cell_6t
Xbit_r229_c61 bl[61] br[61] wl[229] vdd gnd cell_6t
Xbit_r230_c61 bl[61] br[61] wl[230] vdd gnd cell_6t
Xbit_r231_c61 bl[61] br[61] wl[231] vdd gnd cell_6t
Xbit_r232_c61 bl[61] br[61] wl[232] vdd gnd cell_6t
Xbit_r233_c61 bl[61] br[61] wl[233] vdd gnd cell_6t
Xbit_r234_c61 bl[61] br[61] wl[234] vdd gnd cell_6t
Xbit_r235_c61 bl[61] br[61] wl[235] vdd gnd cell_6t
Xbit_r236_c61 bl[61] br[61] wl[236] vdd gnd cell_6t
Xbit_r237_c61 bl[61] br[61] wl[237] vdd gnd cell_6t
Xbit_r238_c61 bl[61] br[61] wl[238] vdd gnd cell_6t
Xbit_r239_c61 bl[61] br[61] wl[239] vdd gnd cell_6t
Xbit_r240_c61 bl[61] br[61] wl[240] vdd gnd cell_6t
Xbit_r241_c61 bl[61] br[61] wl[241] vdd gnd cell_6t
Xbit_r242_c61 bl[61] br[61] wl[242] vdd gnd cell_6t
Xbit_r243_c61 bl[61] br[61] wl[243] vdd gnd cell_6t
Xbit_r244_c61 bl[61] br[61] wl[244] vdd gnd cell_6t
Xbit_r245_c61 bl[61] br[61] wl[245] vdd gnd cell_6t
Xbit_r246_c61 bl[61] br[61] wl[246] vdd gnd cell_6t
Xbit_r247_c61 bl[61] br[61] wl[247] vdd gnd cell_6t
Xbit_r248_c61 bl[61] br[61] wl[248] vdd gnd cell_6t
Xbit_r249_c61 bl[61] br[61] wl[249] vdd gnd cell_6t
Xbit_r250_c61 bl[61] br[61] wl[250] vdd gnd cell_6t
Xbit_r251_c61 bl[61] br[61] wl[251] vdd gnd cell_6t
Xbit_r252_c61 bl[61] br[61] wl[252] vdd gnd cell_6t
Xbit_r253_c61 bl[61] br[61] wl[253] vdd gnd cell_6t
Xbit_r254_c61 bl[61] br[61] wl[254] vdd gnd cell_6t
Xbit_r255_c61 bl[61] br[61] wl[255] vdd gnd cell_6t
Xbit_r0_c62 bl[62] br[62] wl[0] vdd gnd cell_6t
Xbit_r1_c62 bl[62] br[62] wl[1] vdd gnd cell_6t
Xbit_r2_c62 bl[62] br[62] wl[2] vdd gnd cell_6t
Xbit_r3_c62 bl[62] br[62] wl[3] vdd gnd cell_6t
Xbit_r4_c62 bl[62] br[62] wl[4] vdd gnd cell_6t
Xbit_r5_c62 bl[62] br[62] wl[5] vdd gnd cell_6t
Xbit_r6_c62 bl[62] br[62] wl[6] vdd gnd cell_6t
Xbit_r7_c62 bl[62] br[62] wl[7] vdd gnd cell_6t
Xbit_r8_c62 bl[62] br[62] wl[8] vdd gnd cell_6t
Xbit_r9_c62 bl[62] br[62] wl[9] vdd gnd cell_6t
Xbit_r10_c62 bl[62] br[62] wl[10] vdd gnd cell_6t
Xbit_r11_c62 bl[62] br[62] wl[11] vdd gnd cell_6t
Xbit_r12_c62 bl[62] br[62] wl[12] vdd gnd cell_6t
Xbit_r13_c62 bl[62] br[62] wl[13] vdd gnd cell_6t
Xbit_r14_c62 bl[62] br[62] wl[14] vdd gnd cell_6t
Xbit_r15_c62 bl[62] br[62] wl[15] vdd gnd cell_6t
Xbit_r16_c62 bl[62] br[62] wl[16] vdd gnd cell_6t
Xbit_r17_c62 bl[62] br[62] wl[17] vdd gnd cell_6t
Xbit_r18_c62 bl[62] br[62] wl[18] vdd gnd cell_6t
Xbit_r19_c62 bl[62] br[62] wl[19] vdd gnd cell_6t
Xbit_r20_c62 bl[62] br[62] wl[20] vdd gnd cell_6t
Xbit_r21_c62 bl[62] br[62] wl[21] vdd gnd cell_6t
Xbit_r22_c62 bl[62] br[62] wl[22] vdd gnd cell_6t
Xbit_r23_c62 bl[62] br[62] wl[23] vdd gnd cell_6t
Xbit_r24_c62 bl[62] br[62] wl[24] vdd gnd cell_6t
Xbit_r25_c62 bl[62] br[62] wl[25] vdd gnd cell_6t
Xbit_r26_c62 bl[62] br[62] wl[26] vdd gnd cell_6t
Xbit_r27_c62 bl[62] br[62] wl[27] vdd gnd cell_6t
Xbit_r28_c62 bl[62] br[62] wl[28] vdd gnd cell_6t
Xbit_r29_c62 bl[62] br[62] wl[29] vdd gnd cell_6t
Xbit_r30_c62 bl[62] br[62] wl[30] vdd gnd cell_6t
Xbit_r31_c62 bl[62] br[62] wl[31] vdd gnd cell_6t
Xbit_r32_c62 bl[62] br[62] wl[32] vdd gnd cell_6t
Xbit_r33_c62 bl[62] br[62] wl[33] vdd gnd cell_6t
Xbit_r34_c62 bl[62] br[62] wl[34] vdd gnd cell_6t
Xbit_r35_c62 bl[62] br[62] wl[35] vdd gnd cell_6t
Xbit_r36_c62 bl[62] br[62] wl[36] vdd gnd cell_6t
Xbit_r37_c62 bl[62] br[62] wl[37] vdd gnd cell_6t
Xbit_r38_c62 bl[62] br[62] wl[38] vdd gnd cell_6t
Xbit_r39_c62 bl[62] br[62] wl[39] vdd gnd cell_6t
Xbit_r40_c62 bl[62] br[62] wl[40] vdd gnd cell_6t
Xbit_r41_c62 bl[62] br[62] wl[41] vdd gnd cell_6t
Xbit_r42_c62 bl[62] br[62] wl[42] vdd gnd cell_6t
Xbit_r43_c62 bl[62] br[62] wl[43] vdd gnd cell_6t
Xbit_r44_c62 bl[62] br[62] wl[44] vdd gnd cell_6t
Xbit_r45_c62 bl[62] br[62] wl[45] vdd gnd cell_6t
Xbit_r46_c62 bl[62] br[62] wl[46] vdd gnd cell_6t
Xbit_r47_c62 bl[62] br[62] wl[47] vdd gnd cell_6t
Xbit_r48_c62 bl[62] br[62] wl[48] vdd gnd cell_6t
Xbit_r49_c62 bl[62] br[62] wl[49] vdd gnd cell_6t
Xbit_r50_c62 bl[62] br[62] wl[50] vdd gnd cell_6t
Xbit_r51_c62 bl[62] br[62] wl[51] vdd gnd cell_6t
Xbit_r52_c62 bl[62] br[62] wl[52] vdd gnd cell_6t
Xbit_r53_c62 bl[62] br[62] wl[53] vdd gnd cell_6t
Xbit_r54_c62 bl[62] br[62] wl[54] vdd gnd cell_6t
Xbit_r55_c62 bl[62] br[62] wl[55] vdd gnd cell_6t
Xbit_r56_c62 bl[62] br[62] wl[56] vdd gnd cell_6t
Xbit_r57_c62 bl[62] br[62] wl[57] vdd gnd cell_6t
Xbit_r58_c62 bl[62] br[62] wl[58] vdd gnd cell_6t
Xbit_r59_c62 bl[62] br[62] wl[59] vdd gnd cell_6t
Xbit_r60_c62 bl[62] br[62] wl[60] vdd gnd cell_6t
Xbit_r61_c62 bl[62] br[62] wl[61] vdd gnd cell_6t
Xbit_r62_c62 bl[62] br[62] wl[62] vdd gnd cell_6t
Xbit_r63_c62 bl[62] br[62] wl[63] vdd gnd cell_6t
Xbit_r64_c62 bl[62] br[62] wl[64] vdd gnd cell_6t
Xbit_r65_c62 bl[62] br[62] wl[65] vdd gnd cell_6t
Xbit_r66_c62 bl[62] br[62] wl[66] vdd gnd cell_6t
Xbit_r67_c62 bl[62] br[62] wl[67] vdd gnd cell_6t
Xbit_r68_c62 bl[62] br[62] wl[68] vdd gnd cell_6t
Xbit_r69_c62 bl[62] br[62] wl[69] vdd gnd cell_6t
Xbit_r70_c62 bl[62] br[62] wl[70] vdd gnd cell_6t
Xbit_r71_c62 bl[62] br[62] wl[71] vdd gnd cell_6t
Xbit_r72_c62 bl[62] br[62] wl[72] vdd gnd cell_6t
Xbit_r73_c62 bl[62] br[62] wl[73] vdd gnd cell_6t
Xbit_r74_c62 bl[62] br[62] wl[74] vdd gnd cell_6t
Xbit_r75_c62 bl[62] br[62] wl[75] vdd gnd cell_6t
Xbit_r76_c62 bl[62] br[62] wl[76] vdd gnd cell_6t
Xbit_r77_c62 bl[62] br[62] wl[77] vdd gnd cell_6t
Xbit_r78_c62 bl[62] br[62] wl[78] vdd gnd cell_6t
Xbit_r79_c62 bl[62] br[62] wl[79] vdd gnd cell_6t
Xbit_r80_c62 bl[62] br[62] wl[80] vdd gnd cell_6t
Xbit_r81_c62 bl[62] br[62] wl[81] vdd gnd cell_6t
Xbit_r82_c62 bl[62] br[62] wl[82] vdd gnd cell_6t
Xbit_r83_c62 bl[62] br[62] wl[83] vdd gnd cell_6t
Xbit_r84_c62 bl[62] br[62] wl[84] vdd gnd cell_6t
Xbit_r85_c62 bl[62] br[62] wl[85] vdd gnd cell_6t
Xbit_r86_c62 bl[62] br[62] wl[86] vdd gnd cell_6t
Xbit_r87_c62 bl[62] br[62] wl[87] vdd gnd cell_6t
Xbit_r88_c62 bl[62] br[62] wl[88] vdd gnd cell_6t
Xbit_r89_c62 bl[62] br[62] wl[89] vdd gnd cell_6t
Xbit_r90_c62 bl[62] br[62] wl[90] vdd gnd cell_6t
Xbit_r91_c62 bl[62] br[62] wl[91] vdd gnd cell_6t
Xbit_r92_c62 bl[62] br[62] wl[92] vdd gnd cell_6t
Xbit_r93_c62 bl[62] br[62] wl[93] vdd gnd cell_6t
Xbit_r94_c62 bl[62] br[62] wl[94] vdd gnd cell_6t
Xbit_r95_c62 bl[62] br[62] wl[95] vdd gnd cell_6t
Xbit_r96_c62 bl[62] br[62] wl[96] vdd gnd cell_6t
Xbit_r97_c62 bl[62] br[62] wl[97] vdd gnd cell_6t
Xbit_r98_c62 bl[62] br[62] wl[98] vdd gnd cell_6t
Xbit_r99_c62 bl[62] br[62] wl[99] vdd gnd cell_6t
Xbit_r100_c62 bl[62] br[62] wl[100] vdd gnd cell_6t
Xbit_r101_c62 bl[62] br[62] wl[101] vdd gnd cell_6t
Xbit_r102_c62 bl[62] br[62] wl[102] vdd gnd cell_6t
Xbit_r103_c62 bl[62] br[62] wl[103] vdd gnd cell_6t
Xbit_r104_c62 bl[62] br[62] wl[104] vdd gnd cell_6t
Xbit_r105_c62 bl[62] br[62] wl[105] vdd gnd cell_6t
Xbit_r106_c62 bl[62] br[62] wl[106] vdd gnd cell_6t
Xbit_r107_c62 bl[62] br[62] wl[107] vdd gnd cell_6t
Xbit_r108_c62 bl[62] br[62] wl[108] vdd gnd cell_6t
Xbit_r109_c62 bl[62] br[62] wl[109] vdd gnd cell_6t
Xbit_r110_c62 bl[62] br[62] wl[110] vdd gnd cell_6t
Xbit_r111_c62 bl[62] br[62] wl[111] vdd gnd cell_6t
Xbit_r112_c62 bl[62] br[62] wl[112] vdd gnd cell_6t
Xbit_r113_c62 bl[62] br[62] wl[113] vdd gnd cell_6t
Xbit_r114_c62 bl[62] br[62] wl[114] vdd gnd cell_6t
Xbit_r115_c62 bl[62] br[62] wl[115] vdd gnd cell_6t
Xbit_r116_c62 bl[62] br[62] wl[116] vdd gnd cell_6t
Xbit_r117_c62 bl[62] br[62] wl[117] vdd gnd cell_6t
Xbit_r118_c62 bl[62] br[62] wl[118] vdd gnd cell_6t
Xbit_r119_c62 bl[62] br[62] wl[119] vdd gnd cell_6t
Xbit_r120_c62 bl[62] br[62] wl[120] vdd gnd cell_6t
Xbit_r121_c62 bl[62] br[62] wl[121] vdd gnd cell_6t
Xbit_r122_c62 bl[62] br[62] wl[122] vdd gnd cell_6t
Xbit_r123_c62 bl[62] br[62] wl[123] vdd gnd cell_6t
Xbit_r124_c62 bl[62] br[62] wl[124] vdd gnd cell_6t
Xbit_r125_c62 bl[62] br[62] wl[125] vdd gnd cell_6t
Xbit_r126_c62 bl[62] br[62] wl[126] vdd gnd cell_6t
Xbit_r127_c62 bl[62] br[62] wl[127] vdd gnd cell_6t
Xbit_r128_c62 bl[62] br[62] wl[128] vdd gnd cell_6t
Xbit_r129_c62 bl[62] br[62] wl[129] vdd gnd cell_6t
Xbit_r130_c62 bl[62] br[62] wl[130] vdd gnd cell_6t
Xbit_r131_c62 bl[62] br[62] wl[131] vdd gnd cell_6t
Xbit_r132_c62 bl[62] br[62] wl[132] vdd gnd cell_6t
Xbit_r133_c62 bl[62] br[62] wl[133] vdd gnd cell_6t
Xbit_r134_c62 bl[62] br[62] wl[134] vdd gnd cell_6t
Xbit_r135_c62 bl[62] br[62] wl[135] vdd gnd cell_6t
Xbit_r136_c62 bl[62] br[62] wl[136] vdd gnd cell_6t
Xbit_r137_c62 bl[62] br[62] wl[137] vdd gnd cell_6t
Xbit_r138_c62 bl[62] br[62] wl[138] vdd gnd cell_6t
Xbit_r139_c62 bl[62] br[62] wl[139] vdd gnd cell_6t
Xbit_r140_c62 bl[62] br[62] wl[140] vdd gnd cell_6t
Xbit_r141_c62 bl[62] br[62] wl[141] vdd gnd cell_6t
Xbit_r142_c62 bl[62] br[62] wl[142] vdd gnd cell_6t
Xbit_r143_c62 bl[62] br[62] wl[143] vdd gnd cell_6t
Xbit_r144_c62 bl[62] br[62] wl[144] vdd gnd cell_6t
Xbit_r145_c62 bl[62] br[62] wl[145] vdd gnd cell_6t
Xbit_r146_c62 bl[62] br[62] wl[146] vdd gnd cell_6t
Xbit_r147_c62 bl[62] br[62] wl[147] vdd gnd cell_6t
Xbit_r148_c62 bl[62] br[62] wl[148] vdd gnd cell_6t
Xbit_r149_c62 bl[62] br[62] wl[149] vdd gnd cell_6t
Xbit_r150_c62 bl[62] br[62] wl[150] vdd gnd cell_6t
Xbit_r151_c62 bl[62] br[62] wl[151] vdd gnd cell_6t
Xbit_r152_c62 bl[62] br[62] wl[152] vdd gnd cell_6t
Xbit_r153_c62 bl[62] br[62] wl[153] vdd gnd cell_6t
Xbit_r154_c62 bl[62] br[62] wl[154] vdd gnd cell_6t
Xbit_r155_c62 bl[62] br[62] wl[155] vdd gnd cell_6t
Xbit_r156_c62 bl[62] br[62] wl[156] vdd gnd cell_6t
Xbit_r157_c62 bl[62] br[62] wl[157] vdd gnd cell_6t
Xbit_r158_c62 bl[62] br[62] wl[158] vdd gnd cell_6t
Xbit_r159_c62 bl[62] br[62] wl[159] vdd gnd cell_6t
Xbit_r160_c62 bl[62] br[62] wl[160] vdd gnd cell_6t
Xbit_r161_c62 bl[62] br[62] wl[161] vdd gnd cell_6t
Xbit_r162_c62 bl[62] br[62] wl[162] vdd gnd cell_6t
Xbit_r163_c62 bl[62] br[62] wl[163] vdd gnd cell_6t
Xbit_r164_c62 bl[62] br[62] wl[164] vdd gnd cell_6t
Xbit_r165_c62 bl[62] br[62] wl[165] vdd gnd cell_6t
Xbit_r166_c62 bl[62] br[62] wl[166] vdd gnd cell_6t
Xbit_r167_c62 bl[62] br[62] wl[167] vdd gnd cell_6t
Xbit_r168_c62 bl[62] br[62] wl[168] vdd gnd cell_6t
Xbit_r169_c62 bl[62] br[62] wl[169] vdd gnd cell_6t
Xbit_r170_c62 bl[62] br[62] wl[170] vdd gnd cell_6t
Xbit_r171_c62 bl[62] br[62] wl[171] vdd gnd cell_6t
Xbit_r172_c62 bl[62] br[62] wl[172] vdd gnd cell_6t
Xbit_r173_c62 bl[62] br[62] wl[173] vdd gnd cell_6t
Xbit_r174_c62 bl[62] br[62] wl[174] vdd gnd cell_6t
Xbit_r175_c62 bl[62] br[62] wl[175] vdd gnd cell_6t
Xbit_r176_c62 bl[62] br[62] wl[176] vdd gnd cell_6t
Xbit_r177_c62 bl[62] br[62] wl[177] vdd gnd cell_6t
Xbit_r178_c62 bl[62] br[62] wl[178] vdd gnd cell_6t
Xbit_r179_c62 bl[62] br[62] wl[179] vdd gnd cell_6t
Xbit_r180_c62 bl[62] br[62] wl[180] vdd gnd cell_6t
Xbit_r181_c62 bl[62] br[62] wl[181] vdd gnd cell_6t
Xbit_r182_c62 bl[62] br[62] wl[182] vdd gnd cell_6t
Xbit_r183_c62 bl[62] br[62] wl[183] vdd gnd cell_6t
Xbit_r184_c62 bl[62] br[62] wl[184] vdd gnd cell_6t
Xbit_r185_c62 bl[62] br[62] wl[185] vdd gnd cell_6t
Xbit_r186_c62 bl[62] br[62] wl[186] vdd gnd cell_6t
Xbit_r187_c62 bl[62] br[62] wl[187] vdd gnd cell_6t
Xbit_r188_c62 bl[62] br[62] wl[188] vdd gnd cell_6t
Xbit_r189_c62 bl[62] br[62] wl[189] vdd gnd cell_6t
Xbit_r190_c62 bl[62] br[62] wl[190] vdd gnd cell_6t
Xbit_r191_c62 bl[62] br[62] wl[191] vdd gnd cell_6t
Xbit_r192_c62 bl[62] br[62] wl[192] vdd gnd cell_6t
Xbit_r193_c62 bl[62] br[62] wl[193] vdd gnd cell_6t
Xbit_r194_c62 bl[62] br[62] wl[194] vdd gnd cell_6t
Xbit_r195_c62 bl[62] br[62] wl[195] vdd gnd cell_6t
Xbit_r196_c62 bl[62] br[62] wl[196] vdd gnd cell_6t
Xbit_r197_c62 bl[62] br[62] wl[197] vdd gnd cell_6t
Xbit_r198_c62 bl[62] br[62] wl[198] vdd gnd cell_6t
Xbit_r199_c62 bl[62] br[62] wl[199] vdd gnd cell_6t
Xbit_r200_c62 bl[62] br[62] wl[200] vdd gnd cell_6t
Xbit_r201_c62 bl[62] br[62] wl[201] vdd gnd cell_6t
Xbit_r202_c62 bl[62] br[62] wl[202] vdd gnd cell_6t
Xbit_r203_c62 bl[62] br[62] wl[203] vdd gnd cell_6t
Xbit_r204_c62 bl[62] br[62] wl[204] vdd gnd cell_6t
Xbit_r205_c62 bl[62] br[62] wl[205] vdd gnd cell_6t
Xbit_r206_c62 bl[62] br[62] wl[206] vdd gnd cell_6t
Xbit_r207_c62 bl[62] br[62] wl[207] vdd gnd cell_6t
Xbit_r208_c62 bl[62] br[62] wl[208] vdd gnd cell_6t
Xbit_r209_c62 bl[62] br[62] wl[209] vdd gnd cell_6t
Xbit_r210_c62 bl[62] br[62] wl[210] vdd gnd cell_6t
Xbit_r211_c62 bl[62] br[62] wl[211] vdd gnd cell_6t
Xbit_r212_c62 bl[62] br[62] wl[212] vdd gnd cell_6t
Xbit_r213_c62 bl[62] br[62] wl[213] vdd gnd cell_6t
Xbit_r214_c62 bl[62] br[62] wl[214] vdd gnd cell_6t
Xbit_r215_c62 bl[62] br[62] wl[215] vdd gnd cell_6t
Xbit_r216_c62 bl[62] br[62] wl[216] vdd gnd cell_6t
Xbit_r217_c62 bl[62] br[62] wl[217] vdd gnd cell_6t
Xbit_r218_c62 bl[62] br[62] wl[218] vdd gnd cell_6t
Xbit_r219_c62 bl[62] br[62] wl[219] vdd gnd cell_6t
Xbit_r220_c62 bl[62] br[62] wl[220] vdd gnd cell_6t
Xbit_r221_c62 bl[62] br[62] wl[221] vdd gnd cell_6t
Xbit_r222_c62 bl[62] br[62] wl[222] vdd gnd cell_6t
Xbit_r223_c62 bl[62] br[62] wl[223] vdd gnd cell_6t
Xbit_r224_c62 bl[62] br[62] wl[224] vdd gnd cell_6t
Xbit_r225_c62 bl[62] br[62] wl[225] vdd gnd cell_6t
Xbit_r226_c62 bl[62] br[62] wl[226] vdd gnd cell_6t
Xbit_r227_c62 bl[62] br[62] wl[227] vdd gnd cell_6t
Xbit_r228_c62 bl[62] br[62] wl[228] vdd gnd cell_6t
Xbit_r229_c62 bl[62] br[62] wl[229] vdd gnd cell_6t
Xbit_r230_c62 bl[62] br[62] wl[230] vdd gnd cell_6t
Xbit_r231_c62 bl[62] br[62] wl[231] vdd gnd cell_6t
Xbit_r232_c62 bl[62] br[62] wl[232] vdd gnd cell_6t
Xbit_r233_c62 bl[62] br[62] wl[233] vdd gnd cell_6t
Xbit_r234_c62 bl[62] br[62] wl[234] vdd gnd cell_6t
Xbit_r235_c62 bl[62] br[62] wl[235] vdd gnd cell_6t
Xbit_r236_c62 bl[62] br[62] wl[236] vdd gnd cell_6t
Xbit_r237_c62 bl[62] br[62] wl[237] vdd gnd cell_6t
Xbit_r238_c62 bl[62] br[62] wl[238] vdd gnd cell_6t
Xbit_r239_c62 bl[62] br[62] wl[239] vdd gnd cell_6t
Xbit_r240_c62 bl[62] br[62] wl[240] vdd gnd cell_6t
Xbit_r241_c62 bl[62] br[62] wl[241] vdd gnd cell_6t
Xbit_r242_c62 bl[62] br[62] wl[242] vdd gnd cell_6t
Xbit_r243_c62 bl[62] br[62] wl[243] vdd gnd cell_6t
Xbit_r244_c62 bl[62] br[62] wl[244] vdd gnd cell_6t
Xbit_r245_c62 bl[62] br[62] wl[245] vdd gnd cell_6t
Xbit_r246_c62 bl[62] br[62] wl[246] vdd gnd cell_6t
Xbit_r247_c62 bl[62] br[62] wl[247] vdd gnd cell_6t
Xbit_r248_c62 bl[62] br[62] wl[248] vdd gnd cell_6t
Xbit_r249_c62 bl[62] br[62] wl[249] vdd gnd cell_6t
Xbit_r250_c62 bl[62] br[62] wl[250] vdd gnd cell_6t
Xbit_r251_c62 bl[62] br[62] wl[251] vdd gnd cell_6t
Xbit_r252_c62 bl[62] br[62] wl[252] vdd gnd cell_6t
Xbit_r253_c62 bl[62] br[62] wl[253] vdd gnd cell_6t
Xbit_r254_c62 bl[62] br[62] wl[254] vdd gnd cell_6t
Xbit_r255_c62 bl[62] br[62] wl[255] vdd gnd cell_6t
Xbit_r0_c63 bl[63] br[63] wl[0] vdd gnd cell_6t
Xbit_r1_c63 bl[63] br[63] wl[1] vdd gnd cell_6t
Xbit_r2_c63 bl[63] br[63] wl[2] vdd gnd cell_6t
Xbit_r3_c63 bl[63] br[63] wl[3] vdd gnd cell_6t
Xbit_r4_c63 bl[63] br[63] wl[4] vdd gnd cell_6t
Xbit_r5_c63 bl[63] br[63] wl[5] vdd gnd cell_6t
Xbit_r6_c63 bl[63] br[63] wl[6] vdd gnd cell_6t
Xbit_r7_c63 bl[63] br[63] wl[7] vdd gnd cell_6t
Xbit_r8_c63 bl[63] br[63] wl[8] vdd gnd cell_6t
Xbit_r9_c63 bl[63] br[63] wl[9] vdd gnd cell_6t
Xbit_r10_c63 bl[63] br[63] wl[10] vdd gnd cell_6t
Xbit_r11_c63 bl[63] br[63] wl[11] vdd gnd cell_6t
Xbit_r12_c63 bl[63] br[63] wl[12] vdd gnd cell_6t
Xbit_r13_c63 bl[63] br[63] wl[13] vdd gnd cell_6t
Xbit_r14_c63 bl[63] br[63] wl[14] vdd gnd cell_6t
Xbit_r15_c63 bl[63] br[63] wl[15] vdd gnd cell_6t
Xbit_r16_c63 bl[63] br[63] wl[16] vdd gnd cell_6t
Xbit_r17_c63 bl[63] br[63] wl[17] vdd gnd cell_6t
Xbit_r18_c63 bl[63] br[63] wl[18] vdd gnd cell_6t
Xbit_r19_c63 bl[63] br[63] wl[19] vdd gnd cell_6t
Xbit_r20_c63 bl[63] br[63] wl[20] vdd gnd cell_6t
Xbit_r21_c63 bl[63] br[63] wl[21] vdd gnd cell_6t
Xbit_r22_c63 bl[63] br[63] wl[22] vdd gnd cell_6t
Xbit_r23_c63 bl[63] br[63] wl[23] vdd gnd cell_6t
Xbit_r24_c63 bl[63] br[63] wl[24] vdd gnd cell_6t
Xbit_r25_c63 bl[63] br[63] wl[25] vdd gnd cell_6t
Xbit_r26_c63 bl[63] br[63] wl[26] vdd gnd cell_6t
Xbit_r27_c63 bl[63] br[63] wl[27] vdd gnd cell_6t
Xbit_r28_c63 bl[63] br[63] wl[28] vdd gnd cell_6t
Xbit_r29_c63 bl[63] br[63] wl[29] vdd gnd cell_6t
Xbit_r30_c63 bl[63] br[63] wl[30] vdd gnd cell_6t
Xbit_r31_c63 bl[63] br[63] wl[31] vdd gnd cell_6t
Xbit_r32_c63 bl[63] br[63] wl[32] vdd gnd cell_6t
Xbit_r33_c63 bl[63] br[63] wl[33] vdd gnd cell_6t
Xbit_r34_c63 bl[63] br[63] wl[34] vdd gnd cell_6t
Xbit_r35_c63 bl[63] br[63] wl[35] vdd gnd cell_6t
Xbit_r36_c63 bl[63] br[63] wl[36] vdd gnd cell_6t
Xbit_r37_c63 bl[63] br[63] wl[37] vdd gnd cell_6t
Xbit_r38_c63 bl[63] br[63] wl[38] vdd gnd cell_6t
Xbit_r39_c63 bl[63] br[63] wl[39] vdd gnd cell_6t
Xbit_r40_c63 bl[63] br[63] wl[40] vdd gnd cell_6t
Xbit_r41_c63 bl[63] br[63] wl[41] vdd gnd cell_6t
Xbit_r42_c63 bl[63] br[63] wl[42] vdd gnd cell_6t
Xbit_r43_c63 bl[63] br[63] wl[43] vdd gnd cell_6t
Xbit_r44_c63 bl[63] br[63] wl[44] vdd gnd cell_6t
Xbit_r45_c63 bl[63] br[63] wl[45] vdd gnd cell_6t
Xbit_r46_c63 bl[63] br[63] wl[46] vdd gnd cell_6t
Xbit_r47_c63 bl[63] br[63] wl[47] vdd gnd cell_6t
Xbit_r48_c63 bl[63] br[63] wl[48] vdd gnd cell_6t
Xbit_r49_c63 bl[63] br[63] wl[49] vdd gnd cell_6t
Xbit_r50_c63 bl[63] br[63] wl[50] vdd gnd cell_6t
Xbit_r51_c63 bl[63] br[63] wl[51] vdd gnd cell_6t
Xbit_r52_c63 bl[63] br[63] wl[52] vdd gnd cell_6t
Xbit_r53_c63 bl[63] br[63] wl[53] vdd gnd cell_6t
Xbit_r54_c63 bl[63] br[63] wl[54] vdd gnd cell_6t
Xbit_r55_c63 bl[63] br[63] wl[55] vdd gnd cell_6t
Xbit_r56_c63 bl[63] br[63] wl[56] vdd gnd cell_6t
Xbit_r57_c63 bl[63] br[63] wl[57] vdd gnd cell_6t
Xbit_r58_c63 bl[63] br[63] wl[58] vdd gnd cell_6t
Xbit_r59_c63 bl[63] br[63] wl[59] vdd gnd cell_6t
Xbit_r60_c63 bl[63] br[63] wl[60] vdd gnd cell_6t
Xbit_r61_c63 bl[63] br[63] wl[61] vdd gnd cell_6t
Xbit_r62_c63 bl[63] br[63] wl[62] vdd gnd cell_6t
Xbit_r63_c63 bl[63] br[63] wl[63] vdd gnd cell_6t
Xbit_r64_c63 bl[63] br[63] wl[64] vdd gnd cell_6t
Xbit_r65_c63 bl[63] br[63] wl[65] vdd gnd cell_6t
Xbit_r66_c63 bl[63] br[63] wl[66] vdd gnd cell_6t
Xbit_r67_c63 bl[63] br[63] wl[67] vdd gnd cell_6t
Xbit_r68_c63 bl[63] br[63] wl[68] vdd gnd cell_6t
Xbit_r69_c63 bl[63] br[63] wl[69] vdd gnd cell_6t
Xbit_r70_c63 bl[63] br[63] wl[70] vdd gnd cell_6t
Xbit_r71_c63 bl[63] br[63] wl[71] vdd gnd cell_6t
Xbit_r72_c63 bl[63] br[63] wl[72] vdd gnd cell_6t
Xbit_r73_c63 bl[63] br[63] wl[73] vdd gnd cell_6t
Xbit_r74_c63 bl[63] br[63] wl[74] vdd gnd cell_6t
Xbit_r75_c63 bl[63] br[63] wl[75] vdd gnd cell_6t
Xbit_r76_c63 bl[63] br[63] wl[76] vdd gnd cell_6t
Xbit_r77_c63 bl[63] br[63] wl[77] vdd gnd cell_6t
Xbit_r78_c63 bl[63] br[63] wl[78] vdd gnd cell_6t
Xbit_r79_c63 bl[63] br[63] wl[79] vdd gnd cell_6t
Xbit_r80_c63 bl[63] br[63] wl[80] vdd gnd cell_6t
Xbit_r81_c63 bl[63] br[63] wl[81] vdd gnd cell_6t
Xbit_r82_c63 bl[63] br[63] wl[82] vdd gnd cell_6t
Xbit_r83_c63 bl[63] br[63] wl[83] vdd gnd cell_6t
Xbit_r84_c63 bl[63] br[63] wl[84] vdd gnd cell_6t
Xbit_r85_c63 bl[63] br[63] wl[85] vdd gnd cell_6t
Xbit_r86_c63 bl[63] br[63] wl[86] vdd gnd cell_6t
Xbit_r87_c63 bl[63] br[63] wl[87] vdd gnd cell_6t
Xbit_r88_c63 bl[63] br[63] wl[88] vdd gnd cell_6t
Xbit_r89_c63 bl[63] br[63] wl[89] vdd gnd cell_6t
Xbit_r90_c63 bl[63] br[63] wl[90] vdd gnd cell_6t
Xbit_r91_c63 bl[63] br[63] wl[91] vdd gnd cell_6t
Xbit_r92_c63 bl[63] br[63] wl[92] vdd gnd cell_6t
Xbit_r93_c63 bl[63] br[63] wl[93] vdd gnd cell_6t
Xbit_r94_c63 bl[63] br[63] wl[94] vdd gnd cell_6t
Xbit_r95_c63 bl[63] br[63] wl[95] vdd gnd cell_6t
Xbit_r96_c63 bl[63] br[63] wl[96] vdd gnd cell_6t
Xbit_r97_c63 bl[63] br[63] wl[97] vdd gnd cell_6t
Xbit_r98_c63 bl[63] br[63] wl[98] vdd gnd cell_6t
Xbit_r99_c63 bl[63] br[63] wl[99] vdd gnd cell_6t
Xbit_r100_c63 bl[63] br[63] wl[100] vdd gnd cell_6t
Xbit_r101_c63 bl[63] br[63] wl[101] vdd gnd cell_6t
Xbit_r102_c63 bl[63] br[63] wl[102] vdd gnd cell_6t
Xbit_r103_c63 bl[63] br[63] wl[103] vdd gnd cell_6t
Xbit_r104_c63 bl[63] br[63] wl[104] vdd gnd cell_6t
Xbit_r105_c63 bl[63] br[63] wl[105] vdd gnd cell_6t
Xbit_r106_c63 bl[63] br[63] wl[106] vdd gnd cell_6t
Xbit_r107_c63 bl[63] br[63] wl[107] vdd gnd cell_6t
Xbit_r108_c63 bl[63] br[63] wl[108] vdd gnd cell_6t
Xbit_r109_c63 bl[63] br[63] wl[109] vdd gnd cell_6t
Xbit_r110_c63 bl[63] br[63] wl[110] vdd gnd cell_6t
Xbit_r111_c63 bl[63] br[63] wl[111] vdd gnd cell_6t
Xbit_r112_c63 bl[63] br[63] wl[112] vdd gnd cell_6t
Xbit_r113_c63 bl[63] br[63] wl[113] vdd gnd cell_6t
Xbit_r114_c63 bl[63] br[63] wl[114] vdd gnd cell_6t
Xbit_r115_c63 bl[63] br[63] wl[115] vdd gnd cell_6t
Xbit_r116_c63 bl[63] br[63] wl[116] vdd gnd cell_6t
Xbit_r117_c63 bl[63] br[63] wl[117] vdd gnd cell_6t
Xbit_r118_c63 bl[63] br[63] wl[118] vdd gnd cell_6t
Xbit_r119_c63 bl[63] br[63] wl[119] vdd gnd cell_6t
Xbit_r120_c63 bl[63] br[63] wl[120] vdd gnd cell_6t
Xbit_r121_c63 bl[63] br[63] wl[121] vdd gnd cell_6t
Xbit_r122_c63 bl[63] br[63] wl[122] vdd gnd cell_6t
Xbit_r123_c63 bl[63] br[63] wl[123] vdd gnd cell_6t
Xbit_r124_c63 bl[63] br[63] wl[124] vdd gnd cell_6t
Xbit_r125_c63 bl[63] br[63] wl[125] vdd gnd cell_6t
Xbit_r126_c63 bl[63] br[63] wl[126] vdd gnd cell_6t
Xbit_r127_c63 bl[63] br[63] wl[127] vdd gnd cell_6t
Xbit_r128_c63 bl[63] br[63] wl[128] vdd gnd cell_6t
Xbit_r129_c63 bl[63] br[63] wl[129] vdd gnd cell_6t
Xbit_r130_c63 bl[63] br[63] wl[130] vdd gnd cell_6t
Xbit_r131_c63 bl[63] br[63] wl[131] vdd gnd cell_6t
Xbit_r132_c63 bl[63] br[63] wl[132] vdd gnd cell_6t
Xbit_r133_c63 bl[63] br[63] wl[133] vdd gnd cell_6t
Xbit_r134_c63 bl[63] br[63] wl[134] vdd gnd cell_6t
Xbit_r135_c63 bl[63] br[63] wl[135] vdd gnd cell_6t
Xbit_r136_c63 bl[63] br[63] wl[136] vdd gnd cell_6t
Xbit_r137_c63 bl[63] br[63] wl[137] vdd gnd cell_6t
Xbit_r138_c63 bl[63] br[63] wl[138] vdd gnd cell_6t
Xbit_r139_c63 bl[63] br[63] wl[139] vdd gnd cell_6t
Xbit_r140_c63 bl[63] br[63] wl[140] vdd gnd cell_6t
Xbit_r141_c63 bl[63] br[63] wl[141] vdd gnd cell_6t
Xbit_r142_c63 bl[63] br[63] wl[142] vdd gnd cell_6t
Xbit_r143_c63 bl[63] br[63] wl[143] vdd gnd cell_6t
Xbit_r144_c63 bl[63] br[63] wl[144] vdd gnd cell_6t
Xbit_r145_c63 bl[63] br[63] wl[145] vdd gnd cell_6t
Xbit_r146_c63 bl[63] br[63] wl[146] vdd gnd cell_6t
Xbit_r147_c63 bl[63] br[63] wl[147] vdd gnd cell_6t
Xbit_r148_c63 bl[63] br[63] wl[148] vdd gnd cell_6t
Xbit_r149_c63 bl[63] br[63] wl[149] vdd gnd cell_6t
Xbit_r150_c63 bl[63] br[63] wl[150] vdd gnd cell_6t
Xbit_r151_c63 bl[63] br[63] wl[151] vdd gnd cell_6t
Xbit_r152_c63 bl[63] br[63] wl[152] vdd gnd cell_6t
Xbit_r153_c63 bl[63] br[63] wl[153] vdd gnd cell_6t
Xbit_r154_c63 bl[63] br[63] wl[154] vdd gnd cell_6t
Xbit_r155_c63 bl[63] br[63] wl[155] vdd gnd cell_6t
Xbit_r156_c63 bl[63] br[63] wl[156] vdd gnd cell_6t
Xbit_r157_c63 bl[63] br[63] wl[157] vdd gnd cell_6t
Xbit_r158_c63 bl[63] br[63] wl[158] vdd gnd cell_6t
Xbit_r159_c63 bl[63] br[63] wl[159] vdd gnd cell_6t
Xbit_r160_c63 bl[63] br[63] wl[160] vdd gnd cell_6t
Xbit_r161_c63 bl[63] br[63] wl[161] vdd gnd cell_6t
Xbit_r162_c63 bl[63] br[63] wl[162] vdd gnd cell_6t
Xbit_r163_c63 bl[63] br[63] wl[163] vdd gnd cell_6t
Xbit_r164_c63 bl[63] br[63] wl[164] vdd gnd cell_6t
Xbit_r165_c63 bl[63] br[63] wl[165] vdd gnd cell_6t
Xbit_r166_c63 bl[63] br[63] wl[166] vdd gnd cell_6t
Xbit_r167_c63 bl[63] br[63] wl[167] vdd gnd cell_6t
Xbit_r168_c63 bl[63] br[63] wl[168] vdd gnd cell_6t
Xbit_r169_c63 bl[63] br[63] wl[169] vdd gnd cell_6t
Xbit_r170_c63 bl[63] br[63] wl[170] vdd gnd cell_6t
Xbit_r171_c63 bl[63] br[63] wl[171] vdd gnd cell_6t
Xbit_r172_c63 bl[63] br[63] wl[172] vdd gnd cell_6t
Xbit_r173_c63 bl[63] br[63] wl[173] vdd gnd cell_6t
Xbit_r174_c63 bl[63] br[63] wl[174] vdd gnd cell_6t
Xbit_r175_c63 bl[63] br[63] wl[175] vdd gnd cell_6t
Xbit_r176_c63 bl[63] br[63] wl[176] vdd gnd cell_6t
Xbit_r177_c63 bl[63] br[63] wl[177] vdd gnd cell_6t
Xbit_r178_c63 bl[63] br[63] wl[178] vdd gnd cell_6t
Xbit_r179_c63 bl[63] br[63] wl[179] vdd gnd cell_6t
Xbit_r180_c63 bl[63] br[63] wl[180] vdd gnd cell_6t
Xbit_r181_c63 bl[63] br[63] wl[181] vdd gnd cell_6t
Xbit_r182_c63 bl[63] br[63] wl[182] vdd gnd cell_6t
Xbit_r183_c63 bl[63] br[63] wl[183] vdd gnd cell_6t
Xbit_r184_c63 bl[63] br[63] wl[184] vdd gnd cell_6t
Xbit_r185_c63 bl[63] br[63] wl[185] vdd gnd cell_6t
Xbit_r186_c63 bl[63] br[63] wl[186] vdd gnd cell_6t
Xbit_r187_c63 bl[63] br[63] wl[187] vdd gnd cell_6t
Xbit_r188_c63 bl[63] br[63] wl[188] vdd gnd cell_6t
Xbit_r189_c63 bl[63] br[63] wl[189] vdd gnd cell_6t
Xbit_r190_c63 bl[63] br[63] wl[190] vdd gnd cell_6t
Xbit_r191_c63 bl[63] br[63] wl[191] vdd gnd cell_6t
Xbit_r192_c63 bl[63] br[63] wl[192] vdd gnd cell_6t
Xbit_r193_c63 bl[63] br[63] wl[193] vdd gnd cell_6t
Xbit_r194_c63 bl[63] br[63] wl[194] vdd gnd cell_6t
Xbit_r195_c63 bl[63] br[63] wl[195] vdd gnd cell_6t
Xbit_r196_c63 bl[63] br[63] wl[196] vdd gnd cell_6t
Xbit_r197_c63 bl[63] br[63] wl[197] vdd gnd cell_6t
Xbit_r198_c63 bl[63] br[63] wl[198] vdd gnd cell_6t
Xbit_r199_c63 bl[63] br[63] wl[199] vdd gnd cell_6t
Xbit_r200_c63 bl[63] br[63] wl[200] vdd gnd cell_6t
Xbit_r201_c63 bl[63] br[63] wl[201] vdd gnd cell_6t
Xbit_r202_c63 bl[63] br[63] wl[202] vdd gnd cell_6t
Xbit_r203_c63 bl[63] br[63] wl[203] vdd gnd cell_6t
Xbit_r204_c63 bl[63] br[63] wl[204] vdd gnd cell_6t
Xbit_r205_c63 bl[63] br[63] wl[205] vdd gnd cell_6t
Xbit_r206_c63 bl[63] br[63] wl[206] vdd gnd cell_6t
Xbit_r207_c63 bl[63] br[63] wl[207] vdd gnd cell_6t
Xbit_r208_c63 bl[63] br[63] wl[208] vdd gnd cell_6t
Xbit_r209_c63 bl[63] br[63] wl[209] vdd gnd cell_6t
Xbit_r210_c63 bl[63] br[63] wl[210] vdd gnd cell_6t
Xbit_r211_c63 bl[63] br[63] wl[211] vdd gnd cell_6t
Xbit_r212_c63 bl[63] br[63] wl[212] vdd gnd cell_6t
Xbit_r213_c63 bl[63] br[63] wl[213] vdd gnd cell_6t
Xbit_r214_c63 bl[63] br[63] wl[214] vdd gnd cell_6t
Xbit_r215_c63 bl[63] br[63] wl[215] vdd gnd cell_6t
Xbit_r216_c63 bl[63] br[63] wl[216] vdd gnd cell_6t
Xbit_r217_c63 bl[63] br[63] wl[217] vdd gnd cell_6t
Xbit_r218_c63 bl[63] br[63] wl[218] vdd gnd cell_6t
Xbit_r219_c63 bl[63] br[63] wl[219] vdd gnd cell_6t
Xbit_r220_c63 bl[63] br[63] wl[220] vdd gnd cell_6t
Xbit_r221_c63 bl[63] br[63] wl[221] vdd gnd cell_6t
Xbit_r222_c63 bl[63] br[63] wl[222] vdd gnd cell_6t
Xbit_r223_c63 bl[63] br[63] wl[223] vdd gnd cell_6t
Xbit_r224_c63 bl[63] br[63] wl[224] vdd gnd cell_6t
Xbit_r225_c63 bl[63] br[63] wl[225] vdd gnd cell_6t
Xbit_r226_c63 bl[63] br[63] wl[226] vdd gnd cell_6t
Xbit_r227_c63 bl[63] br[63] wl[227] vdd gnd cell_6t
Xbit_r228_c63 bl[63] br[63] wl[228] vdd gnd cell_6t
Xbit_r229_c63 bl[63] br[63] wl[229] vdd gnd cell_6t
Xbit_r230_c63 bl[63] br[63] wl[230] vdd gnd cell_6t
Xbit_r231_c63 bl[63] br[63] wl[231] vdd gnd cell_6t
Xbit_r232_c63 bl[63] br[63] wl[232] vdd gnd cell_6t
Xbit_r233_c63 bl[63] br[63] wl[233] vdd gnd cell_6t
Xbit_r234_c63 bl[63] br[63] wl[234] vdd gnd cell_6t
Xbit_r235_c63 bl[63] br[63] wl[235] vdd gnd cell_6t
Xbit_r236_c63 bl[63] br[63] wl[236] vdd gnd cell_6t
Xbit_r237_c63 bl[63] br[63] wl[237] vdd gnd cell_6t
Xbit_r238_c63 bl[63] br[63] wl[238] vdd gnd cell_6t
Xbit_r239_c63 bl[63] br[63] wl[239] vdd gnd cell_6t
Xbit_r240_c63 bl[63] br[63] wl[240] vdd gnd cell_6t
Xbit_r241_c63 bl[63] br[63] wl[241] vdd gnd cell_6t
Xbit_r242_c63 bl[63] br[63] wl[242] vdd gnd cell_6t
Xbit_r243_c63 bl[63] br[63] wl[243] vdd gnd cell_6t
Xbit_r244_c63 bl[63] br[63] wl[244] vdd gnd cell_6t
Xbit_r245_c63 bl[63] br[63] wl[245] vdd gnd cell_6t
Xbit_r246_c63 bl[63] br[63] wl[246] vdd gnd cell_6t
Xbit_r247_c63 bl[63] br[63] wl[247] vdd gnd cell_6t
Xbit_r248_c63 bl[63] br[63] wl[248] vdd gnd cell_6t
Xbit_r249_c63 bl[63] br[63] wl[249] vdd gnd cell_6t
Xbit_r250_c63 bl[63] br[63] wl[250] vdd gnd cell_6t
Xbit_r251_c63 bl[63] br[63] wl[251] vdd gnd cell_6t
Xbit_r252_c63 bl[63] br[63] wl[252] vdd gnd cell_6t
Xbit_r253_c63 bl[63] br[63] wl[253] vdd gnd cell_6t
Xbit_r254_c63 bl[63] br[63] wl[254] vdd gnd cell_6t
Xbit_r255_c63 bl[63] br[63] wl[255] vdd gnd cell_6t
Xbit_r0_c64 bl[64] br[64] wl[0] vdd gnd cell_6t
Xbit_r1_c64 bl[64] br[64] wl[1] vdd gnd cell_6t
Xbit_r2_c64 bl[64] br[64] wl[2] vdd gnd cell_6t
Xbit_r3_c64 bl[64] br[64] wl[3] vdd gnd cell_6t
Xbit_r4_c64 bl[64] br[64] wl[4] vdd gnd cell_6t
Xbit_r5_c64 bl[64] br[64] wl[5] vdd gnd cell_6t
Xbit_r6_c64 bl[64] br[64] wl[6] vdd gnd cell_6t
Xbit_r7_c64 bl[64] br[64] wl[7] vdd gnd cell_6t
Xbit_r8_c64 bl[64] br[64] wl[8] vdd gnd cell_6t
Xbit_r9_c64 bl[64] br[64] wl[9] vdd gnd cell_6t
Xbit_r10_c64 bl[64] br[64] wl[10] vdd gnd cell_6t
Xbit_r11_c64 bl[64] br[64] wl[11] vdd gnd cell_6t
Xbit_r12_c64 bl[64] br[64] wl[12] vdd gnd cell_6t
Xbit_r13_c64 bl[64] br[64] wl[13] vdd gnd cell_6t
Xbit_r14_c64 bl[64] br[64] wl[14] vdd gnd cell_6t
Xbit_r15_c64 bl[64] br[64] wl[15] vdd gnd cell_6t
Xbit_r16_c64 bl[64] br[64] wl[16] vdd gnd cell_6t
Xbit_r17_c64 bl[64] br[64] wl[17] vdd gnd cell_6t
Xbit_r18_c64 bl[64] br[64] wl[18] vdd gnd cell_6t
Xbit_r19_c64 bl[64] br[64] wl[19] vdd gnd cell_6t
Xbit_r20_c64 bl[64] br[64] wl[20] vdd gnd cell_6t
Xbit_r21_c64 bl[64] br[64] wl[21] vdd gnd cell_6t
Xbit_r22_c64 bl[64] br[64] wl[22] vdd gnd cell_6t
Xbit_r23_c64 bl[64] br[64] wl[23] vdd gnd cell_6t
Xbit_r24_c64 bl[64] br[64] wl[24] vdd gnd cell_6t
Xbit_r25_c64 bl[64] br[64] wl[25] vdd gnd cell_6t
Xbit_r26_c64 bl[64] br[64] wl[26] vdd gnd cell_6t
Xbit_r27_c64 bl[64] br[64] wl[27] vdd gnd cell_6t
Xbit_r28_c64 bl[64] br[64] wl[28] vdd gnd cell_6t
Xbit_r29_c64 bl[64] br[64] wl[29] vdd gnd cell_6t
Xbit_r30_c64 bl[64] br[64] wl[30] vdd gnd cell_6t
Xbit_r31_c64 bl[64] br[64] wl[31] vdd gnd cell_6t
Xbit_r32_c64 bl[64] br[64] wl[32] vdd gnd cell_6t
Xbit_r33_c64 bl[64] br[64] wl[33] vdd gnd cell_6t
Xbit_r34_c64 bl[64] br[64] wl[34] vdd gnd cell_6t
Xbit_r35_c64 bl[64] br[64] wl[35] vdd gnd cell_6t
Xbit_r36_c64 bl[64] br[64] wl[36] vdd gnd cell_6t
Xbit_r37_c64 bl[64] br[64] wl[37] vdd gnd cell_6t
Xbit_r38_c64 bl[64] br[64] wl[38] vdd gnd cell_6t
Xbit_r39_c64 bl[64] br[64] wl[39] vdd gnd cell_6t
Xbit_r40_c64 bl[64] br[64] wl[40] vdd gnd cell_6t
Xbit_r41_c64 bl[64] br[64] wl[41] vdd gnd cell_6t
Xbit_r42_c64 bl[64] br[64] wl[42] vdd gnd cell_6t
Xbit_r43_c64 bl[64] br[64] wl[43] vdd gnd cell_6t
Xbit_r44_c64 bl[64] br[64] wl[44] vdd gnd cell_6t
Xbit_r45_c64 bl[64] br[64] wl[45] vdd gnd cell_6t
Xbit_r46_c64 bl[64] br[64] wl[46] vdd gnd cell_6t
Xbit_r47_c64 bl[64] br[64] wl[47] vdd gnd cell_6t
Xbit_r48_c64 bl[64] br[64] wl[48] vdd gnd cell_6t
Xbit_r49_c64 bl[64] br[64] wl[49] vdd gnd cell_6t
Xbit_r50_c64 bl[64] br[64] wl[50] vdd gnd cell_6t
Xbit_r51_c64 bl[64] br[64] wl[51] vdd gnd cell_6t
Xbit_r52_c64 bl[64] br[64] wl[52] vdd gnd cell_6t
Xbit_r53_c64 bl[64] br[64] wl[53] vdd gnd cell_6t
Xbit_r54_c64 bl[64] br[64] wl[54] vdd gnd cell_6t
Xbit_r55_c64 bl[64] br[64] wl[55] vdd gnd cell_6t
Xbit_r56_c64 bl[64] br[64] wl[56] vdd gnd cell_6t
Xbit_r57_c64 bl[64] br[64] wl[57] vdd gnd cell_6t
Xbit_r58_c64 bl[64] br[64] wl[58] vdd gnd cell_6t
Xbit_r59_c64 bl[64] br[64] wl[59] vdd gnd cell_6t
Xbit_r60_c64 bl[64] br[64] wl[60] vdd gnd cell_6t
Xbit_r61_c64 bl[64] br[64] wl[61] vdd gnd cell_6t
Xbit_r62_c64 bl[64] br[64] wl[62] vdd gnd cell_6t
Xbit_r63_c64 bl[64] br[64] wl[63] vdd gnd cell_6t
Xbit_r64_c64 bl[64] br[64] wl[64] vdd gnd cell_6t
Xbit_r65_c64 bl[64] br[64] wl[65] vdd gnd cell_6t
Xbit_r66_c64 bl[64] br[64] wl[66] vdd gnd cell_6t
Xbit_r67_c64 bl[64] br[64] wl[67] vdd gnd cell_6t
Xbit_r68_c64 bl[64] br[64] wl[68] vdd gnd cell_6t
Xbit_r69_c64 bl[64] br[64] wl[69] vdd gnd cell_6t
Xbit_r70_c64 bl[64] br[64] wl[70] vdd gnd cell_6t
Xbit_r71_c64 bl[64] br[64] wl[71] vdd gnd cell_6t
Xbit_r72_c64 bl[64] br[64] wl[72] vdd gnd cell_6t
Xbit_r73_c64 bl[64] br[64] wl[73] vdd gnd cell_6t
Xbit_r74_c64 bl[64] br[64] wl[74] vdd gnd cell_6t
Xbit_r75_c64 bl[64] br[64] wl[75] vdd gnd cell_6t
Xbit_r76_c64 bl[64] br[64] wl[76] vdd gnd cell_6t
Xbit_r77_c64 bl[64] br[64] wl[77] vdd gnd cell_6t
Xbit_r78_c64 bl[64] br[64] wl[78] vdd gnd cell_6t
Xbit_r79_c64 bl[64] br[64] wl[79] vdd gnd cell_6t
Xbit_r80_c64 bl[64] br[64] wl[80] vdd gnd cell_6t
Xbit_r81_c64 bl[64] br[64] wl[81] vdd gnd cell_6t
Xbit_r82_c64 bl[64] br[64] wl[82] vdd gnd cell_6t
Xbit_r83_c64 bl[64] br[64] wl[83] vdd gnd cell_6t
Xbit_r84_c64 bl[64] br[64] wl[84] vdd gnd cell_6t
Xbit_r85_c64 bl[64] br[64] wl[85] vdd gnd cell_6t
Xbit_r86_c64 bl[64] br[64] wl[86] vdd gnd cell_6t
Xbit_r87_c64 bl[64] br[64] wl[87] vdd gnd cell_6t
Xbit_r88_c64 bl[64] br[64] wl[88] vdd gnd cell_6t
Xbit_r89_c64 bl[64] br[64] wl[89] vdd gnd cell_6t
Xbit_r90_c64 bl[64] br[64] wl[90] vdd gnd cell_6t
Xbit_r91_c64 bl[64] br[64] wl[91] vdd gnd cell_6t
Xbit_r92_c64 bl[64] br[64] wl[92] vdd gnd cell_6t
Xbit_r93_c64 bl[64] br[64] wl[93] vdd gnd cell_6t
Xbit_r94_c64 bl[64] br[64] wl[94] vdd gnd cell_6t
Xbit_r95_c64 bl[64] br[64] wl[95] vdd gnd cell_6t
Xbit_r96_c64 bl[64] br[64] wl[96] vdd gnd cell_6t
Xbit_r97_c64 bl[64] br[64] wl[97] vdd gnd cell_6t
Xbit_r98_c64 bl[64] br[64] wl[98] vdd gnd cell_6t
Xbit_r99_c64 bl[64] br[64] wl[99] vdd gnd cell_6t
Xbit_r100_c64 bl[64] br[64] wl[100] vdd gnd cell_6t
Xbit_r101_c64 bl[64] br[64] wl[101] vdd gnd cell_6t
Xbit_r102_c64 bl[64] br[64] wl[102] vdd gnd cell_6t
Xbit_r103_c64 bl[64] br[64] wl[103] vdd gnd cell_6t
Xbit_r104_c64 bl[64] br[64] wl[104] vdd gnd cell_6t
Xbit_r105_c64 bl[64] br[64] wl[105] vdd gnd cell_6t
Xbit_r106_c64 bl[64] br[64] wl[106] vdd gnd cell_6t
Xbit_r107_c64 bl[64] br[64] wl[107] vdd gnd cell_6t
Xbit_r108_c64 bl[64] br[64] wl[108] vdd gnd cell_6t
Xbit_r109_c64 bl[64] br[64] wl[109] vdd gnd cell_6t
Xbit_r110_c64 bl[64] br[64] wl[110] vdd gnd cell_6t
Xbit_r111_c64 bl[64] br[64] wl[111] vdd gnd cell_6t
Xbit_r112_c64 bl[64] br[64] wl[112] vdd gnd cell_6t
Xbit_r113_c64 bl[64] br[64] wl[113] vdd gnd cell_6t
Xbit_r114_c64 bl[64] br[64] wl[114] vdd gnd cell_6t
Xbit_r115_c64 bl[64] br[64] wl[115] vdd gnd cell_6t
Xbit_r116_c64 bl[64] br[64] wl[116] vdd gnd cell_6t
Xbit_r117_c64 bl[64] br[64] wl[117] vdd gnd cell_6t
Xbit_r118_c64 bl[64] br[64] wl[118] vdd gnd cell_6t
Xbit_r119_c64 bl[64] br[64] wl[119] vdd gnd cell_6t
Xbit_r120_c64 bl[64] br[64] wl[120] vdd gnd cell_6t
Xbit_r121_c64 bl[64] br[64] wl[121] vdd gnd cell_6t
Xbit_r122_c64 bl[64] br[64] wl[122] vdd gnd cell_6t
Xbit_r123_c64 bl[64] br[64] wl[123] vdd gnd cell_6t
Xbit_r124_c64 bl[64] br[64] wl[124] vdd gnd cell_6t
Xbit_r125_c64 bl[64] br[64] wl[125] vdd gnd cell_6t
Xbit_r126_c64 bl[64] br[64] wl[126] vdd gnd cell_6t
Xbit_r127_c64 bl[64] br[64] wl[127] vdd gnd cell_6t
Xbit_r128_c64 bl[64] br[64] wl[128] vdd gnd cell_6t
Xbit_r129_c64 bl[64] br[64] wl[129] vdd gnd cell_6t
Xbit_r130_c64 bl[64] br[64] wl[130] vdd gnd cell_6t
Xbit_r131_c64 bl[64] br[64] wl[131] vdd gnd cell_6t
Xbit_r132_c64 bl[64] br[64] wl[132] vdd gnd cell_6t
Xbit_r133_c64 bl[64] br[64] wl[133] vdd gnd cell_6t
Xbit_r134_c64 bl[64] br[64] wl[134] vdd gnd cell_6t
Xbit_r135_c64 bl[64] br[64] wl[135] vdd gnd cell_6t
Xbit_r136_c64 bl[64] br[64] wl[136] vdd gnd cell_6t
Xbit_r137_c64 bl[64] br[64] wl[137] vdd gnd cell_6t
Xbit_r138_c64 bl[64] br[64] wl[138] vdd gnd cell_6t
Xbit_r139_c64 bl[64] br[64] wl[139] vdd gnd cell_6t
Xbit_r140_c64 bl[64] br[64] wl[140] vdd gnd cell_6t
Xbit_r141_c64 bl[64] br[64] wl[141] vdd gnd cell_6t
Xbit_r142_c64 bl[64] br[64] wl[142] vdd gnd cell_6t
Xbit_r143_c64 bl[64] br[64] wl[143] vdd gnd cell_6t
Xbit_r144_c64 bl[64] br[64] wl[144] vdd gnd cell_6t
Xbit_r145_c64 bl[64] br[64] wl[145] vdd gnd cell_6t
Xbit_r146_c64 bl[64] br[64] wl[146] vdd gnd cell_6t
Xbit_r147_c64 bl[64] br[64] wl[147] vdd gnd cell_6t
Xbit_r148_c64 bl[64] br[64] wl[148] vdd gnd cell_6t
Xbit_r149_c64 bl[64] br[64] wl[149] vdd gnd cell_6t
Xbit_r150_c64 bl[64] br[64] wl[150] vdd gnd cell_6t
Xbit_r151_c64 bl[64] br[64] wl[151] vdd gnd cell_6t
Xbit_r152_c64 bl[64] br[64] wl[152] vdd gnd cell_6t
Xbit_r153_c64 bl[64] br[64] wl[153] vdd gnd cell_6t
Xbit_r154_c64 bl[64] br[64] wl[154] vdd gnd cell_6t
Xbit_r155_c64 bl[64] br[64] wl[155] vdd gnd cell_6t
Xbit_r156_c64 bl[64] br[64] wl[156] vdd gnd cell_6t
Xbit_r157_c64 bl[64] br[64] wl[157] vdd gnd cell_6t
Xbit_r158_c64 bl[64] br[64] wl[158] vdd gnd cell_6t
Xbit_r159_c64 bl[64] br[64] wl[159] vdd gnd cell_6t
Xbit_r160_c64 bl[64] br[64] wl[160] vdd gnd cell_6t
Xbit_r161_c64 bl[64] br[64] wl[161] vdd gnd cell_6t
Xbit_r162_c64 bl[64] br[64] wl[162] vdd gnd cell_6t
Xbit_r163_c64 bl[64] br[64] wl[163] vdd gnd cell_6t
Xbit_r164_c64 bl[64] br[64] wl[164] vdd gnd cell_6t
Xbit_r165_c64 bl[64] br[64] wl[165] vdd gnd cell_6t
Xbit_r166_c64 bl[64] br[64] wl[166] vdd gnd cell_6t
Xbit_r167_c64 bl[64] br[64] wl[167] vdd gnd cell_6t
Xbit_r168_c64 bl[64] br[64] wl[168] vdd gnd cell_6t
Xbit_r169_c64 bl[64] br[64] wl[169] vdd gnd cell_6t
Xbit_r170_c64 bl[64] br[64] wl[170] vdd gnd cell_6t
Xbit_r171_c64 bl[64] br[64] wl[171] vdd gnd cell_6t
Xbit_r172_c64 bl[64] br[64] wl[172] vdd gnd cell_6t
Xbit_r173_c64 bl[64] br[64] wl[173] vdd gnd cell_6t
Xbit_r174_c64 bl[64] br[64] wl[174] vdd gnd cell_6t
Xbit_r175_c64 bl[64] br[64] wl[175] vdd gnd cell_6t
Xbit_r176_c64 bl[64] br[64] wl[176] vdd gnd cell_6t
Xbit_r177_c64 bl[64] br[64] wl[177] vdd gnd cell_6t
Xbit_r178_c64 bl[64] br[64] wl[178] vdd gnd cell_6t
Xbit_r179_c64 bl[64] br[64] wl[179] vdd gnd cell_6t
Xbit_r180_c64 bl[64] br[64] wl[180] vdd gnd cell_6t
Xbit_r181_c64 bl[64] br[64] wl[181] vdd gnd cell_6t
Xbit_r182_c64 bl[64] br[64] wl[182] vdd gnd cell_6t
Xbit_r183_c64 bl[64] br[64] wl[183] vdd gnd cell_6t
Xbit_r184_c64 bl[64] br[64] wl[184] vdd gnd cell_6t
Xbit_r185_c64 bl[64] br[64] wl[185] vdd gnd cell_6t
Xbit_r186_c64 bl[64] br[64] wl[186] vdd gnd cell_6t
Xbit_r187_c64 bl[64] br[64] wl[187] vdd gnd cell_6t
Xbit_r188_c64 bl[64] br[64] wl[188] vdd gnd cell_6t
Xbit_r189_c64 bl[64] br[64] wl[189] vdd gnd cell_6t
Xbit_r190_c64 bl[64] br[64] wl[190] vdd gnd cell_6t
Xbit_r191_c64 bl[64] br[64] wl[191] vdd gnd cell_6t
Xbit_r192_c64 bl[64] br[64] wl[192] vdd gnd cell_6t
Xbit_r193_c64 bl[64] br[64] wl[193] vdd gnd cell_6t
Xbit_r194_c64 bl[64] br[64] wl[194] vdd gnd cell_6t
Xbit_r195_c64 bl[64] br[64] wl[195] vdd gnd cell_6t
Xbit_r196_c64 bl[64] br[64] wl[196] vdd gnd cell_6t
Xbit_r197_c64 bl[64] br[64] wl[197] vdd gnd cell_6t
Xbit_r198_c64 bl[64] br[64] wl[198] vdd gnd cell_6t
Xbit_r199_c64 bl[64] br[64] wl[199] vdd gnd cell_6t
Xbit_r200_c64 bl[64] br[64] wl[200] vdd gnd cell_6t
Xbit_r201_c64 bl[64] br[64] wl[201] vdd gnd cell_6t
Xbit_r202_c64 bl[64] br[64] wl[202] vdd gnd cell_6t
Xbit_r203_c64 bl[64] br[64] wl[203] vdd gnd cell_6t
Xbit_r204_c64 bl[64] br[64] wl[204] vdd gnd cell_6t
Xbit_r205_c64 bl[64] br[64] wl[205] vdd gnd cell_6t
Xbit_r206_c64 bl[64] br[64] wl[206] vdd gnd cell_6t
Xbit_r207_c64 bl[64] br[64] wl[207] vdd gnd cell_6t
Xbit_r208_c64 bl[64] br[64] wl[208] vdd gnd cell_6t
Xbit_r209_c64 bl[64] br[64] wl[209] vdd gnd cell_6t
Xbit_r210_c64 bl[64] br[64] wl[210] vdd gnd cell_6t
Xbit_r211_c64 bl[64] br[64] wl[211] vdd gnd cell_6t
Xbit_r212_c64 bl[64] br[64] wl[212] vdd gnd cell_6t
Xbit_r213_c64 bl[64] br[64] wl[213] vdd gnd cell_6t
Xbit_r214_c64 bl[64] br[64] wl[214] vdd gnd cell_6t
Xbit_r215_c64 bl[64] br[64] wl[215] vdd gnd cell_6t
Xbit_r216_c64 bl[64] br[64] wl[216] vdd gnd cell_6t
Xbit_r217_c64 bl[64] br[64] wl[217] vdd gnd cell_6t
Xbit_r218_c64 bl[64] br[64] wl[218] vdd gnd cell_6t
Xbit_r219_c64 bl[64] br[64] wl[219] vdd gnd cell_6t
Xbit_r220_c64 bl[64] br[64] wl[220] vdd gnd cell_6t
Xbit_r221_c64 bl[64] br[64] wl[221] vdd gnd cell_6t
Xbit_r222_c64 bl[64] br[64] wl[222] vdd gnd cell_6t
Xbit_r223_c64 bl[64] br[64] wl[223] vdd gnd cell_6t
Xbit_r224_c64 bl[64] br[64] wl[224] vdd gnd cell_6t
Xbit_r225_c64 bl[64] br[64] wl[225] vdd gnd cell_6t
Xbit_r226_c64 bl[64] br[64] wl[226] vdd gnd cell_6t
Xbit_r227_c64 bl[64] br[64] wl[227] vdd gnd cell_6t
Xbit_r228_c64 bl[64] br[64] wl[228] vdd gnd cell_6t
Xbit_r229_c64 bl[64] br[64] wl[229] vdd gnd cell_6t
Xbit_r230_c64 bl[64] br[64] wl[230] vdd gnd cell_6t
Xbit_r231_c64 bl[64] br[64] wl[231] vdd gnd cell_6t
Xbit_r232_c64 bl[64] br[64] wl[232] vdd gnd cell_6t
Xbit_r233_c64 bl[64] br[64] wl[233] vdd gnd cell_6t
Xbit_r234_c64 bl[64] br[64] wl[234] vdd gnd cell_6t
Xbit_r235_c64 bl[64] br[64] wl[235] vdd gnd cell_6t
Xbit_r236_c64 bl[64] br[64] wl[236] vdd gnd cell_6t
Xbit_r237_c64 bl[64] br[64] wl[237] vdd gnd cell_6t
Xbit_r238_c64 bl[64] br[64] wl[238] vdd gnd cell_6t
Xbit_r239_c64 bl[64] br[64] wl[239] vdd gnd cell_6t
Xbit_r240_c64 bl[64] br[64] wl[240] vdd gnd cell_6t
Xbit_r241_c64 bl[64] br[64] wl[241] vdd gnd cell_6t
Xbit_r242_c64 bl[64] br[64] wl[242] vdd gnd cell_6t
Xbit_r243_c64 bl[64] br[64] wl[243] vdd gnd cell_6t
Xbit_r244_c64 bl[64] br[64] wl[244] vdd gnd cell_6t
Xbit_r245_c64 bl[64] br[64] wl[245] vdd gnd cell_6t
Xbit_r246_c64 bl[64] br[64] wl[246] vdd gnd cell_6t
Xbit_r247_c64 bl[64] br[64] wl[247] vdd gnd cell_6t
Xbit_r248_c64 bl[64] br[64] wl[248] vdd gnd cell_6t
Xbit_r249_c64 bl[64] br[64] wl[249] vdd gnd cell_6t
Xbit_r250_c64 bl[64] br[64] wl[250] vdd gnd cell_6t
Xbit_r251_c64 bl[64] br[64] wl[251] vdd gnd cell_6t
Xbit_r252_c64 bl[64] br[64] wl[252] vdd gnd cell_6t
Xbit_r253_c64 bl[64] br[64] wl[253] vdd gnd cell_6t
Xbit_r254_c64 bl[64] br[64] wl[254] vdd gnd cell_6t
Xbit_r255_c64 bl[64] br[64] wl[255] vdd gnd cell_6t
Xbit_r0_c65 bl[65] br[65] wl[0] vdd gnd cell_6t
Xbit_r1_c65 bl[65] br[65] wl[1] vdd gnd cell_6t
Xbit_r2_c65 bl[65] br[65] wl[2] vdd gnd cell_6t
Xbit_r3_c65 bl[65] br[65] wl[3] vdd gnd cell_6t
Xbit_r4_c65 bl[65] br[65] wl[4] vdd gnd cell_6t
Xbit_r5_c65 bl[65] br[65] wl[5] vdd gnd cell_6t
Xbit_r6_c65 bl[65] br[65] wl[6] vdd gnd cell_6t
Xbit_r7_c65 bl[65] br[65] wl[7] vdd gnd cell_6t
Xbit_r8_c65 bl[65] br[65] wl[8] vdd gnd cell_6t
Xbit_r9_c65 bl[65] br[65] wl[9] vdd gnd cell_6t
Xbit_r10_c65 bl[65] br[65] wl[10] vdd gnd cell_6t
Xbit_r11_c65 bl[65] br[65] wl[11] vdd gnd cell_6t
Xbit_r12_c65 bl[65] br[65] wl[12] vdd gnd cell_6t
Xbit_r13_c65 bl[65] br[65] wl[13] vdd gnd cell_6t
Xbit_r14_c65 bl[65] br[65] wl[14] vdd gnd cell_6t
Xbit_r15_c65 bl[65] br[65] wl[15] vdd gnd cell_6t
Xbit_r16_c65 bl[65] br[65] wl[16] vdd gnd cell_6t
Xbit_r17_c65 bl[65] br[65] wl[17] vdd gnd cell_6t
Xbit_r18_c65 bl[65] br[65] wl[18] vdd gnd cell_6t
Xbit_r19_c65 bl[65] br[65] wl[19] vdd gnd cell_6t
Xbit_r20_c65 bl[65] br[65] wl[20] vdd gnd cell_6t
Xbit_r21_c65 bl[65] br[65] wl[21] vdd gnd cell_6t
Xbit_r22_c65 bl[65] br[65] wl[22] vdd gnd cell_6t
Xbit_r23_c65 bl[65] br[65] wl[23] vdd gnd cell_6t
Xbit_r24_c65 bl[65] br[65] wl[24] vdd gnd cell_6t
Xbit_r25_c65 bl[65] br[65] wl[25] vdd gnd cell_6t
Xbit_r26_c65 bl[65] br[65] wl[26] vdd gnd cell_6t
Xbit_r27_c65 bl[65] br[65] wl[27] vdd gnd cell_6t
Xbit_r28_c65 bl[65] br[65] wl[28] vdd gnd cell_6t
Xbit_r29_c65 bl[65] br[65] wl[29] vdd gnd cell_6t
Xbit_r30_c65 bl[65] br[65] wl[30] vdd gnd cell_6t
Xbit_r31_c65 bl[65] br[65] wl[31] vdd gnd cell_6t
Xbit_r32_c65 bl[65] br[65] wl[32] vdd gnd cell_6t
Xbit_r33_c65 bl[65] br[65] wl[33] vdd gnd cell_6t
Xbit_r34_c65 bl[65] br[65] wl[34] vdd gnd cell_6t
Xbit_r35_c65 bl[65] br[65] wl[35] vdd gnd cell_6t
Xbit_r36_c65 bl[65] br[65] wl[36] vdd gnd cell_6t
Xbit_r37_c65 bl[65] br[65] wl[37] vdd gnd cell_6t
Xbit_r38_c65 bl[65] br[65] wl[38] vdd gnd cell_6t
Xbit_r39_c65 bl[65] br[65] wl[39] vdd gnd cell_6t
Xbit_r40_c65 bl[65] br[65] wl[40] vdd gnd cell_6t
Xbit_r41_c65 bl[65] br[65] wl[41] vdd gnd cell_6t
Xbit_r42_c65 bl[65] br[65] wl[42] vdd gnd cell_6t
Xbit_r43_c65 bl[65] br[65] wl[43] vdd gnd cell_6t
Xbit_r44_c65 bl[65] br[65] wl[44] vdd gnd cell_6t
Xbit_r45_c65 bl[65] br[65] wl[45] vdd gnd cell_6t
Xbit_r46_c65 bl[65] br[65] wl[46] vdd gnd cell_6t
Xbit_r47_c65 bl[65] br[65] wl[47] vdd gnd cell_6t
Xbit_r48_c65 bl[65] br[65] wl[48] vdd gnd cell_6t
Xbit_r49_c65 bl[65] br[65] wl[49] vdd gnd cell_6t
Xbit_r50_c65 bl[65] br[65] wl[50] vdd gnd cell_6t
Xbit_r51_c65 bl[65] br[65] wl[51] vdd gnd cell_6t
Xbit_r52_c65 bl[65] br[65] wl[52] vdd gnd cell_6t
Xbit_r53_c65 bl[65] br[65] wl[53] vdd gnd cell_6t
Xbit_r54_c65 bl[65] br[65] wl[54] vdd gnd cell_6t
Xbit_r55_c65 bl[65] br[65] wl[55] vdd gnd cell_6t
Xbit_r56_c65 bl[65] br[65] wl[56] vdd gnd cell_6t
Xbit_r57_c65 bl[65] br[65] wl[57] vdd gnd cell_6t
Xbit_r58_c65 bl[65] br[65] wl[58] vdd gnd cell_6t
Xbit_r59_c65 bl[65] br[65] wl[59] vdd gnd cell_6t
Xbit_r60_c65 bl[65] br[65] wl[60] vdd gnd cell_6t
Xbit_r61_c65 bl[65] br[65] wl[61] vdd gnd cell_6t
Xbit_r62_c65 bl[65] br[65] wl[62] vdd gnd cell_6t
Xbit_r63_c65 bl[65] br[65] wl[63] vdd gnd cell_6t
Xbit_r64_c65 bl[65] br[65] wl[64] vdd gnd cell_6t
Xbit_r65_c65 bl[65] br[65] wl[65] vdd gnd cell_6t
Xbit_r66_c65 bl[65] br[65] wl[66] vdd gnd cell_6t
Xbit_r67_c65 bl[65] br[65] wl[67] vdd gnd cell_6t
Xbit_r68_c65 bl[65] br[65] wl[68] vdd gnd cell_6t
Xbit_r69_c65 bl[65] br[65] wl[69] vdd gnd cell_6t
Xbit_r70_c65 bl[65] br[65] wl[70] vdd gnd cell_6t
Xbit_r71_c65 bl[65] br[65] wl[71] vdd gnd cell_6t
Xbit_r72_c65 bl[65] br[65] wl[72] vdd gnd cell_6t
Xbit_r73_c65 bl[65] br[65] wl[73] vdd gnd cell_6t
Xbit_r74_c65 bl[65] br[65] wl[74] vdd gnd cell_6t
Xbit_r75_c65 bl[65] br[65] wl[75] vdd gnd cell_6t
Xbit_r76_c65 bl[65] br[65] wl[76] vdd gnd cell_6t
Xbit_r77_c65 bl[65] br[65] wl[77] vdd gnd cell_6t
Xbit_r78_c65 bl[65] br[65] wl[78] vdd gnd cell_6t
Xbit_r79_c65 bl[65] br[65] wl[79] vdd gnd cell_6t
Xbit_r80_c65 bl[65] br[65] wl[80] vdd gnd cell_6t
Xbit_r81_c65 bl[65] br[65] wl[81] vdd gnd cell_6t
Xbit_r82_c65 bl[65] br[65] wl[82] vdd gnd cell_6t
Xbit_r83_c65 bl[65] br[65] wl[83] vdd gnd cell_6t
Xbit_r84_c65 bl[65] br[65] wl[84] vdd gnd cell_6t
Xbit_r85_c65 bl[65] br[65] wl[85] vdd gnd cell_6t
Xbit_r86_c65 bl[65] br[65] wl[86] vdd gnd cell_6t
Xbit_r87_c65 bl[65] br[65] wl[87] vdd gnd cell_6t
Xbit_r88_c65 bl[65] br[65] wl[88] vdd gnd cell_6t
Xbit_r89_c65 bl[65] br[65] wl[89] vdd gnd cell_6t
Xbit_r90_c65 bl[65] br[65] wl[90] vdd gnd cell_6t
Xbit_r91_c65 bl[65] br[65] wl[91] vdd gnd cell_6t
Xbit_r92_c65 bl[65] br[65] wl[92] vdd gnd cell_6t
Xbit_r93_c65 bl[65] br[65] wl[93] vdd gnd cell_6t
Xbit_r94_c65 bl[65] br[65] wl[94] vdd gnd cell_6t
Xbit_r95_c65 bl[65] br[65] wl[95] vdd gnd cell_6t
Xbit_r96_c65 bl[65] br[65] wl[96] vdd gnd cell_6t
Xbit_r97_c65 bl[65] br[65] wl[97] vdd gnd cell_6t
Xbit_r98_c65 bl[65] br[65] wl[98] vdd gnd cell_6t
Xbit_r99_c65 bl[65] br[65] wl[99] vdd gnd cell_6t
Xbit_r100_c65 bl[65] br[65] wl[100] vdd gnd cell_6t
Xbit_r101_c65 bl[65] br[65] wl[101] vdd gnd cell_6t
Xbit_r102_c65 bl[65] br[65] wl[102] vdd gnd cell_6t
Xbit_r103_c65 bl[65] br[65] wl[103] vdd gnd cell_6t
Xbit_r104_c65 bl[65] br[65] wl[104] vdd gnd cell_6t
Xbit_r105_c65 bl[65] br[65] wl[105] vdd gnd cell_6t
Xbit_r106_c65 bl[65] br[65] wl[106] vdd gnd cell_6t
Xbit_r107_c65 bl[65] br[65] wl[107] vdd gnd cell_6t
Xbit_r108_c65 bl[65] br[65] wl[108] vdd gnd cell_6t
Xbit_r109_c65 bl[65] br[65] wl[109] vdd gnd cell_6t
Xbit_r110_c65 bl[65] br[65] wl[110] vdd gnd cell_6t
Xbit_r111_c65 bl[65] br[65] wl[111] vdd gnd cell_6t
Xbit_r112_c65 bl[65] br[65] wl[112] vdd gnd cell_6t
Xbit_r113_c65 bl[65] br[65] wl[113] vdd gnd cell_6t
Xbit_r114_c65 bl[65] br[65] wl[114] vdd gnd cell_6t
Xbit_r115_c65 bl[65] br[65] wl[115] vdd gnd cell_6t
Xbit_r116_c65 bl[65] br[65] wl[116] vdd gnd cell_6t
Xbit_r117_c65 bl[65] br[65] wl[117] vdd gnd cell_6t
Xbit_r118_c65 bl[65] br[65] wl[118] vdd gnd cell_6t
Xbit_r119_c65 bl[65] br[65] wl[119] vdd gnd cell_6t
Xbit_r120_c65 bl[65] br[65] wl[120] vdd gnd cell_6t
Xbit_r121_c65 bl[65] br[65] wl[121] vdd gnd cell_6t
Xbit_r122_c65 bl[65] br[65] wl[122] vdd gnd cell_6t
Xbit_r123_c65 bl[65] br[65] wl[123] vdd gnd cell_6t
Xbit_r124_c65 bl[65] br[65] wl[124] vdd gnd cell_6t
Xbit_r125_c65 bl[65] br[65] wl[125] vdd gnd cell_6t
Xbit_r126_c65 bl[65] br[65] wl[126] vdd gnd cell_6t
Xbit_r127_c65 bl[65] br[65] wl[127] vdd gnd cell_6t
Xbit_r128_c65 bl[65] br[65] wl[128] vdd gnd cell_6t
Xbit_r129_c65 bl[65] br[65] wl[129] vdd gnd cell_6t
Xbit_r130_c65 bl[65] br[65] wl[130] vdd gnd cell_6t
Xbit_r131_c65 bl[65] br[65] wl[131] vdd gnd cell_6t
Xbit_r132_c65 bl[65] br[65] wl[132] vdd gnd cell_6t
Xbit_r133_c65 bl[65] br[65] wl[133] vdd gnd cell_6t
Xbit_r134_c65 bl[65] br[65] wl[134] vdd gnd cell_6t
Xbit_r135_c65 bl[65] br[65] wl[135] vdd gnd cell_6t
Xbit_r136_c65 bl[65] br[65] wl[136] vdd gnd cell_6t
Xbit_r137_c65 bl[65] br[65] wl[137] vdd gnd cell_6t
Xbit_r138_c65 bl[65] br[65] wl[138] vdd gnd cell_6t
Xbit_r139_c65 bl[65] br[65] wl[139] vdd gnd cell_6t
Xbit_r140_c65 bl[65] br[65] wl[140] vdd gnd cell_6t
Xbit_r141_c65 bl[65] br[65] wl[141] vdd gnd cell_6t
Xbit_r142_c65 bl[65] br[65] wl[142] vdd gnd cell_6t
Xbit_r143_c65 bl[65] br[65] wl[143] vdd gnd cell_6t
Xbit_r144_c65 bl[65] br[65] wl[144] vdd gnd cell_6t
Xbit_r145_c65 bl[65] br[65] wl[145] vdd gnd cell_6t
Xbit_r146_c65 bl[65] br[65] wl[146] vdd gnd cell_6t
Xbit_r147_c65 bl[65] br[65] wl[147] vdd gnd cell_6t
Xbit_r148_c65 bl[65] br[65] wl[148] vdd gnd cell_6t
Xbit_r149_c65 bl[65] br[65] wl[149] vdd gnd cell_6t
Xbit_r150_c65 bl[65] br[65] wl[150] vdd gnd cell_6t
Xbit_r151_c65 bl[65] br[65] wl[151] vdd gnd cell_6t
Xbit_r152_c65 bl[65] br[65] wl[152] vdd gnd cell_6t
Xbit_r153_c65 bl[65] br[65] wl[153] vdd gnd cell_6t
Xbit_r154_c65 bl[65] br[65] wl[154] vdd gnd cell_6t
Xbit_r155_c65 bl[65] br[65] wl[155] vdd gnd cell_6t
Xbit_r156_c65 bl[65] br[65] wl[156] vdd gnd cell_6t
Xbit_r157_c65 bl[65] br[65] wl[157] vdd gnd cell_6t
Xbit_r158_c65 bl[65] br[65] wl[158] vdd gnd cell_6t
Xbit_r159_c65 bl[65] br[65] wl[159] vdd gnd cell_6t
Xbit_r160_c65 bl[65] br[65] wl[160] vdd gnd cell_6t
Xbit_r161_c65 bl[65] br[65] wl[161] vdd gnd cell_6t
Xbit_r162_c65 bl[65] br[65] wl[162] vdd gnd cell_6t
Xbit_r163_c65 bl[65] br[65] wl[163] vdd gnd cell_6t
Xbit_r164_c65 bl[65] br[65] wl[164] vdd gnd cell_6t
Xbit_r165_c65 bl[65] br[65] wl[165] vdd gnd cell_6t
Xbit_r166_c65 bl[65] br[65] wl[166] vdd gnd cell_6t
Xbit_r167_c65 bl[65] br[65] wl[167] vdd gnd cell_6t
Xbit_r168_c65 bl[65] br[65] wl[168] vdd gnd cell_6t
Xbit_r169_c65 bl[65] br[65] wl[169] vdd gnd cell_6t
Xbit_r170_c65 bl[65] br[65] wl[170] vdd gnd cell_6t
Xbit_r171_c65 bl[65] br[65] wl[171] vdd gnd cell_6t
Xbit_r172_c65 bl[65] br[65] wl[172] vdd gnd cell_6t
Xbit_r173_c65 bl[65] br[65] wl[173] vdd gnd cell_6t
Xbit_r174_c65 bl[65] br[65] wl[174] vdd gnd cell_6t
Xbit_r175_c65 bl[65] br[65] wl[175] vdd gnd cell_6t
Xbit_r176_c65 bl[65] br[65] wl[176] vdd gnd cell_6t
Xbit_r177_c65 bl[65] br[65] wl[177] vdd gnd cell_6t
Xbit_r178_c65 bl[65] br[65] wl[178] vdd gnd cell_6t
Xbit_r179_c65 bl[65] br[65] wl[179] vdd gnd cell_6t
Xbit_r180_c65 bl[65] br[65] wl[180] vdd gnd cell_6t
Xbit_r181_c65 bl[65] br[65] wl[181] vdd gnd cell_6t
Xbit_r182_c65 bl[65] br[65] wl[182] vdd gnd cell_6t
Xbit_r183_c65 bl[65] br[65] wl[183] vdd gnd cell_6t
Xbit_r184_c65 bl[65] br[65] wl[184] vdd gnd cell_6t
Xbit_r185_c65 bl[65] br[65] wl[185] vdd gnd cell_6t
Xbit_r186_c65 bl[65] br[65] wl[186] vdd gnd cell_6t
Xbit_r187_c65 bl[65] br[65] wl[187] vdd gnd cell_6t
Xbit_r188_c65 bl[65] br[65] wl[188] vdd gnd cell_6t
Xbit_r189_c65 bl[65] br[65] wl[189] vdd gnd cell_6t
Xbit_r190_c65 bl[65] br[65] wl[190] vdd gnd cell_6t
Xbit_r191_c65 bl[65] br[65] wl[191] vdd gnd cell_6t
Xbit_r192_c65 bl[65] br[65] wl[192] vdd gnd cell_6t
Xbit_r193_c65 bl[65] br[65] wl[193] vdd gnd cell_6t
Xbit_r194_c65 bl[65] br[65] wl[194] vdd gnd cell_6t
Xbit_r195_c65 bl[65] br[65] wl[195] vdd gnd cell_6t
Xbit_r196_c65 bl[65] br[65] wl[196] vdd gnd cell_6t
Xbit_r197_c65 bl[65] br[65] wl[197] vdd gnd cell_6t
Xbit_r198_c65 bl[65] br[65] wl[198] vdd gnd cell_6t
Xbit_r199_c65 bl[65] br[65] wl[199] vdd gnd cell_6t
Xbit_r200_c65 bl[65] br[65] wl[200] vdd gnd cell_6t
Xbit_r201_c65 bl[65] br[65] wl[201] vdd gnd cell_6t
Xbit_r202_c65 bl[65] br[65] wl[202] vdd gnd cell_6t
Xbit_r203_c65 bl[65] br[65] wl[203] vdd gnd cell_6t
Xbit_r204_c65 bl[65] br[65] wl[204] vdd gnd cell_6t
Xbit_r205_c65 bl[65] br[65] wl[205] vdd gnd cell_6t
Xbit_r206_c65 bl[65] br[65] wl[206] vdd gnd cell_6t
Xbit_r207_c65 bl[65] br[65] wl[207] vdd gnd cell_6t
Xbit_r208_c65 bl[65] br[65] wl[208] vdd gnd cell_6t
Xbit_r209_c65 bl[65] br[65] wl[209] vdd gnd cell_6t
Xbit_r210_c65 bl[65] br[65] wl[210] vdd gnd cell_6t
Xbit_r211_c65 bl[65] br[65] wl[211] vdd gnd cell_6t
Xbit_r212_c65 bl[65] br[65] wl[212] vdd gnd cell_6t
Xbit_r213_c65 bl[65] br[65] wl[213] vdd gnd cell_6t
Xbit_r214_c65 bl[65] br[65] wl[214] vdd gnd cell_6t
Xbit_r215_c65 bl[65] br[65] wl[215] vdd gnd cell_6t
Xbit_r216_c65 bl[65] br[65] wl[216] vdd gnd cell_6t
Xbit_r217_c65 bl[65] br[65] wl[217] vdd gnd cell_6t
Xbit_r218_c65 bl[65] br[65] wl[218] vdd gnd cell_6t
Xbit_r219_c65 bl[65] br[65] wl[219] vdd gnd cell_6t
Xbit_r220_c65 bl[65] br[65] wl[220] vdd gnd cell_6t
Xbit_r221_c65 bl[65] br[65] wl[221] vdd gnd cell_6t
Xbit_r222_c65 bl[65] br[65] wl[222] vdd gnd cell_6t
Xbit_r223_c65 bl[65] br[65] wl[223] vdd gnd cell_6t
Xbit_r224_c65 bl[65] br[65] wl[224] vdd gnd cell_6t
Xbit_r225_c65 bl[65] br[65] wl[225] vdd gnd cell_6t
Xbit_r226_c65 bl[65] br[65] wl[226] vdd gnd cell_6t
Xbit_r227_c65 bl[65] br[65] wl[227] vdd gnd cell_6t
Xbit_r228_c65 bl[65] br[65] wl[228] vdd gnd cell_6t
Xbit_r229_c65 bl[65] br[65] wl[229] vdd gnd cell_6t
Xbit_r230_c65 bl[65] br[65] wl[230] vdd gnd cell_6t
Xbit_r231_c65 bl[65] br[65] wl[231] vdd gnd cell_6t
Xbit_r232_c65 bl[65] br[65] wl[232] vdd gnd cell_6t
Xbit_r233_c65 bl[65] br[65] wl[233] vdd gnd cell_6t
Xbit_r234_c65 bl[65] br[65] wl[234] vdd gnd cell_6t
Xbit_r235_c65 bl[65] br[65] wl[235] vdd gnd cell_6t
Xbit_r236_c65 bl[65] br[65] wl[236] vdd gnd cell_6t
Xbit_r237_c65 bl[65] br[65] wl[237] vdd gnd cell_6t
Xbit_r238_c65 bl[65] br[65] wl[238] vdd gnd cell_6t
Xbit_r239_c65 bl[65] br[65] wl[239] vdd gnd cell_6t
Xbit_r240_c65 bl[65] br[65] wl[240] vdd gnd cell_6t
Xbit_r241_c65 bl[65] br[65] wl[241] vdd gnd cell_6t
Xbit_r242_c65 bl[65] br[65] wl[242] vdd gnd cell_6t
Xbit_r243_c65 bl[65] br[65] wl[243] vdd gnd cell_6t
Xbit_r244_c65 bl[65] br[65] wl[244] vdd gnd cell_6t
Xbit_r245_c65 bl[65] br[65] wl[245] vdd gnd cell_6t
Xbit_r246_c65 bl[65] br[65] wl[246] vdd gnd cell_6t
Xbit_r247_c65 bl[65] br[65] wl[247] vdd gnd cell_6t
Xbit_r248_c65 bl[65] br[65] wl[248] vdd gnd cell_6t
Xbit_r249_c65 bl[65] br[65] wl[249] vdd gnd cell_6t
Xbit_r250_c65 bl[65] br[65] wl[250] vdd gnd cell_6t
Xbit_r251_c65 bl[65] br[65] wl[251] vdd gnd cell_6t
Xbit_r252_c65 bl[65] br[65] wl[252] vdd gnd cell_6t
Xbit_r253_c65 bl[65] br[65] wl[253] vdd gnd cell_6t
Xbit_r254_c65 bl[65] br[65] wl[254] vdd gnd cell_6t
Xbit_r255_c65 bl[65] br[65] wl[255] vdd gnd cell_6t
Xbit_r0_c66 bl[66] br[66] wl[0] vdd gnd cell_6t
Xbit_r1_c66 bl[66] br[66] wl[1] vdd gnd cell_6t
Xbit_r2_c66 bl[66] br[66] wl[2] vdd gnd cell_6t
Xbit_r3_c66 bl[66] br[66] wl[3] vdd gnd cell_6t
Xbit_r4_c66 bl[66] br[66] wl[4] vdd gnd cell_6t
Xbit_r5_c66 bl[66] br[66] wl[5] vdd gnd cell_6t
Xbit_r6_c66 bl[66] br[66] wl[6] vdd gnd cell_6t
Xbit_r7_c66 bl[66] br[66] wl[7] vdd gnd cell_6t
Xbit_r8_c66 bl[66] br[66] wl[8] vdd gnd cell_6t
Xbit_r9_c66 bl[66] br[66] wl[9] vdd gnd cell_6t
Xbit_r10_c66 bl[66] br[66] wl[10] vdd gnd cell_6t
Xbit_r11_c66 bl[66] br[66] wl[11] vdd gnd cell_6t
Xbit_r12_c66 bl[66] br[66] wl[12] vdd gnd cell_6t
Xbit_r13_c66 bl[66] br[66] wl[13] vdd gnd cell_6t
Xbit_r14_c66 bl[66] br[66] wl[14] vdd gnd cell_6t
Xbit_r15_c66 bl[66] br[66] wl[15] vdd gnd cell_6t
Xbit_r16_c66 bl[66] br[66] wl[16] vdd gnd cell_6t
Xbit_r17_c66 bl[66] br[66] wl[17] vdd gnd cell_6t
Xbit_r18_c66 bl[66] br[66] wl[18] vdd gnd cell_6t
Xbit_r19_c66 bl[66] br[66] wl[19] vdd gnd cell_6t
Xbit_r20_c66 bl[66] br[66] wl[20] vdd gnd cell_6t
Xbit_r21_c66 bl[66] br[66] wl[21] vdd gnd cell_6t
Xbit_r22_c66 bl[66] br[66] wl[22] vdd gnd cell_6t
Xbit_r23_c66 bl[66] br[66] wl[23] vdd gnd cell_6t
Xbit_r24_c66 bl[66] br[66] wl[24] vdd gnd cell_6t
Xbit_r25_c66 bl[66] br[66] wl[25] vdd gnd cell_6t
Xbit_r26_c66 bl[66] br[66] wl[26] vdd gnd cell_6t
Xbit_r27_c66 bl[66] br[66] wl[27] vdd gnd cell_6t
Xbit_r28_c66 bl[66] br[66] wl[28] vdd gnd cell_6t
Xbit_r29_c66 bl[66] br[66] wl[29] vdd gnd cell_6t
Xbit_r30_c66 bl[66] br[66] wl[30] vdd gnd cell_6t
Xbit_r31_c66 bl[66] br[66] wl[31] vdd gnd cell_6t
Xbit_r32_c66 bl[66] br[66] wl[32] vdd gnd cell_6t
Xbit_r33_c66 bl[66] br[66] wl[33] vdd gnd cell_6t
Xbit_r34_c66 bl[66] br[66] wl[34] vdd gnd cell_6t
Xbit_r35_c66 bl[66] br[66] wl[35] vdd gnd cell_6t
Xbit_r36_c66 bl[66] br[66] wl[36] vdd gnd cell_6t
Xbit_r37_c66 bl[66] br[66] wl[37] vdd gnd cell_6t
Xbit_r38_c66 bl[66] br[66] wl[38] vdd gnd cell_6t
Xbit_r39_c66 bl[66] br[66] wl[39] vdd gnd cell_6t
Xbit_r40_c66 bl[66] br[66] wl[40] vdd gnd cell_6t
Xbit_r41_c66 bl[66] br[66] wl[41] vdd gnd cell_6t
Xbit_r42_c66 bl[66] br[66] wl[42] vdd gnd cell_6t
Xbit_r43_c66 bl[66] br[66] wl[43] vdd gnd cell_6t
Xbit_r44_c66 bl[66] br[66] wl[44] vdd gnd cell_6t
Xbit_r45_c66 bl[66] br[66] wl[45] vdd gnd cell_6t
Xbit_r46_c66 bl[66] br[66] wl[46] vdd gnd cell_6t
Xbit_r47_c66 bl[66] br[66] wl[47] vdd gnd cell_6t
Xbit_r48_c66 bl[66] br[66] wl[48] vdd gnd cell_6t
Xbit_r49_c66 bl[66] br[66] wl[49] vdd gnd cell_6t
Xbit_r50_c66 bl[66] br[66] wl[50] vdd gnd cell_6t
Xbit_r51_c66 bl[66] br[66] wl[51] vdd gnd cell_6t
Xbit_r52_c66 bl[66] br[66] wl[52] vdd gnd cell_6t
Xbit_r53_c66 bl[66] br[66] wl[53] vdd gnd cell_6t
Xbit_r54_c66 bl[66] br[66] wl[54] vdd gnd cell_6t
Xbit_r55_c66 bl[66] br[66] wl[55] vdd gnd cell_6t
Xbit_r56_c66 bl[66] br[66] wl[56] vdd gnd cell_6t
Xbit_r57_c66 bl[66] br[66] wl[57] vdd gnd cell_6t
Xbit_r58_c66 bl[66] br[66] wl[58] vdd gnd cell_6t
Xbit_r59_c66 bl[66] br[66] wl[59] vdd gnd cell_6t
Xbit_r60_c66 bl[66] br[66] wl[60] vdd gnd cell_6t
Xbit_r61_c66 bl[66] br[66] wl[61] vdd gnd cell_6t
Xbit_r62_c66 bl[66] br[66] wl[62] vdd gnd cell_6t
Xbit_r63_c66 bl[66] br[66] wl[63] vdd gnd cell_6t
Xbit_r64_c66 bl[66] br[66] wl[64] vdd gnd cell_6t
Xbit_r65_c66 bl[66] br[66] wl[65] vdd gnd cell_6t
Xbit_r66_c66 bl[66] br[66] wl[66] vdd gnd cell_6t
Xbit_r67_c66 bl[66] br[66] wl[67] vdd gnd cell_6t
Xbit_r68_c66 bl[66] br[66] wl[68] vdd gnd cell_6t
Xbit_r69_c66 bl[66] br[66] wl[69] vdd gnd cell_6t
Xbit_r70_c66 bl[66] br[66] wl[70] vdd gnd cell_6t
Xbit_r71_c66 bl[66] br[66] wl[71] vdd gnd cell_6t
Xbit_r72_c66 bl[66] br[66] wl[72] vdd gnd cell_6t
Xbit_r73_c66 bl[66] br[66] wl[73] vdd gnd cell_6t
Xbit_r74_c66 bl[66] br[66] wl[74] vdd gnd cell_6t
Xbit_r75_c66 bl[66] br[66] wl[75] vdd gnd cell_6t
Xbit_r76_c66 bl[66] br[66] wl[76] vdd gnd cell_6t
Xbit_r77_c66 bl[66] br[66] wl[77] vdd gnd cell_6t
Xbit_r78_c66 bl[66] br[66] wl[78] vdd gnd cell_6t
Xbit_r79_c66 bl[66] br[66] wl[79] vdd gnd cell_6t
Xbit_r80_c66 bl[66] br[66] wl[80] vdd gnd cell_6t
Xbit_r81_c66 bl[66] br[66] wl[81] vdd gnd cell_6t
Xbit_r82_c66 bl[66] br[66] wl[82] vdd gnd cell_6t
Xbit_r83_c66 bl[66] br[66] wl[83] vdd gnd cell_6t
Xbit_r84_c66 bl[66] br[66] wl[84] vdd gnd cell_6t
Xbit_r85_c66 bl[66] br[66] wl[85] vdd gnd cell_6t
Xbit_r86_c66 bl[66] br[66] wl[86] vdd gnd cell_6t
Xbit_r87_c66 bl[66] br[66] wl[87] vdd gnd cell_6t
Xbit_r88_c66 bl[66] br[66] wl[88] vdd gnd cell_6t
Xbit_r89_c66 bl[66] br[66] wl[89] vdd gnd cell_6t
Xbit_r90_c66 bl[66] br[66] wl[90] vdd gnd cell_6t
Xbit_r91_c66 bl[66] br[66] wl[91] vdd gnd cell_6t
Xbit_r92_c66 bl[66] br[66] wl[92] vdd gnd cell_6t
Xbit_r93_c66 bl[66] br[66] wl[93] vdd gnd cell_6t
Xbit_r94_c66 bl[66] br[66] wl[94] vdd gnd cell_6t
Xbit_r95_c66 bl[66] br[66] wl[95] vdd gnd cell_6t
Xbit_r96_c66 bl[66] br[66] wl[96] vdd gnd cell_6t
Xbit_r97_c66 bl[66] br[66] wl[97] vdd gnd cell_6t
Xbit_r98_c66 bl[66] br[66] wl[98] vdd gnd cell_6t
Xbit_r99_c66 bl[66] br[66] wl[99] vdd gnd cell_6t
Xbit_r100_c66 bl[66] br[66] wl[100] vdd gnd cell_6t
Xbit_r101_c66 bl[66] br[66] wl[101] vdd gnd cell_6t
Xbit_r102_c66 bl[66] br[66] wl[102] vdd gnd cell_6t
Xbit_r103_c66 bl[66] br[66] wl[103] vdd gnd cell_6t
Xbit_r104_c66 bl[66] br[66] wl[104] vdd gnd cell_6t
Xbit_r105_c66 bl[66] br[66] wl[105] vdd gnd cell_6t
Xbit_r106_c66 bl[66] br[66] wl[106] vdd gnd cell_6t
Xbit_r107_c66 bl[66] br[66] wl[107] vdd gnd cell_6t
Xbit_r108_c66 bl[66] br[66] wl[108] vdd gnd cell_6t
Xbit_r109_c66 bl[66] br[66] wl[109] vdd gnd cell_6t
Xbit_r110_c66 bl[66] br[66] wl[110] vdd gnd cell_6t
Xbit_r111_c66 bl[66] br[66] wl[111] vdd gnd cell_6t
Xbit_r112_c66 bl[66] br[66] wl[112] vdd gnd cell_6t
Xbit_r113_c66 bl[66] br[66] wl[113] vdd gnd cell_6t
Xbit_r114_c66 bl[66] br[66] wl[114] vdd gnd cell_6t
Xbit_r115_c66 bl[66] br[66] wl[115] vdd gnd cell_6t
Xbit_r116_c66 bl[66] br[66] wl[116] vdd gnd cell_6t
Xbit_r117_c66 bl[66] br[66] wl[117] vdd gnd cell_6t
Xbit_r118_c66 bl[66] br[66] wl[118] vdd gnd cell_6t
Xbit_r119_c66 bl[66] br[66] wl[119] vdd gnd cell_6t
Xbit_r120_c66 bl[66] br[66] wl[120] vdd gnd cell_6t
Xbit_r121_c66 bl[66] br[66] wl[121] vdd gnd cell_6t
Xbit_r122_c66 bl[66] br[66] wl[122] vdd gnd cell_6t
Xbit_r123_c66 bl[66] br[66] wl[123] vdd gnd cell_6t
Xbit_r124_c66 bl[66] br[66] wl[124] vdd gnd cell_6t
Xbit_r125_c66 bl[66] br[66] wl[125] vdd gnd cell_6t
Xbit_r126_c66 bl[66] br[66] wl[126] vdd gnd cell_6t
Xbit_r127_c66 bl[66] br[66] wl[127] vdd gnd cell_6t
Xbit_r128_c66 bl[66] br[66] wl[128] vdd gnd cell_6t
Xbit_r129_c66 bl[66] br[66] wl[129] vdd gnd cell_6t
Xbit_r130_c66 bl[66] br[66] wl[130] vdd gnd cell_6t
Xbit_r131_c66 bl[66] br[66] wl[131] vdd gnd cell_6t
Xbit_r132_c66 bl[66] br[66] wl[132] vdd gnd cell_6t
Xbit_r133_c66 bl[66] br[66] wl[133] vdd gnd cell_6t
Xbit_r134_c66 bl[66] br[66] wl[134] vdd gnd cell_6t
Xbit_r135_c66 bl[66] br[66] wl[135] vdd gnd cell_6t
Xbit_r136_c66 bl[66] br[66] wl[136] vdd gnd cell_6t
Xbit_r137_c66 bl[66] br[66] wl[137] vdd gnd cell_6t
Xbit_r138_c66 bl[66] br[66] wl[138] vdd gnd cell_6t
Xbit_r139_c66 bl[66] br[66] wl[139] vdd gnd cell_6t
Xbit_r140_c66 bl[66] br[66] wl[140] vdd gnd cell_6t
Xbit_r141_c66 bl[66] br[66] wl[141] vdd gnd cell_6t
Xbit_r142_c66 bl[66] br[66] wl[142] vdd gnd cell_6t
Xbit_r143_c66 bl[66] br[66] wl[143] vdd gnd cell_6t
Xbit_r144_c66 bl[66] br[66] wl[144] vdd gnd cell_6t
Xbit_r145_c66 bl[66] br[66] wl[145] vdd gnd cell_6t
Xbit_r146_c66 bl[66] br[66] wl[146] vdd gnd cell_6t
Xbit_r147_c66 bl[66] br[66] wl[147] vdd gnd cell_6t
Xbit_r148_c66 bl[66] br[66] wl[148] vdd gnd cell_6t
Xbit_r149_c66 bl[66] br[66] wl[149] vdd gnd cell_6t
Xbit_r150_c66 bl[66] br[66] wl[150] vdd gnd cell_6t
Xbit_r151_c66 bl[66] br[66] wl[151] vdd gnd cell_6t
Xbit_r152_c66 bl[66] br[66] wl[152] vdd gnd cell_6t
Xbit_r153_c66 bl[66] br[66] wl[153] vdd gnd cell_6t
Xbit_r154_c66 bl[66] br[66] wl[154] vdd gnd cell_6t
Xbit_r155_c66 bl[66] br[66] wl[155] vdd gnd cell_6t
Xbit_r156_c66 bl[66] br[66] wl[156] vdd gnd cell_6t
Xbit_r157_c66 bl[66] br[66] wl[157] vdd gnd cell_6t
Xbit_r158_c66 bl[66] br[66] wl[158] vdd gnd cell_6t
Xbit_r159_c66 bl[66] br[66] wl[159] vdd gnd cell_6t
Xbit_r160_c66 bl[66] br[66] wl[160] vdd gnd cell_6t
Xbit_r161_c66 bl[66] br[66] wl[161] vdd gnd cell_6t
Xbit_r162_c66 bl[66] br[66] wl[162] vdd gnd cell_6t
Xbit_r163_c66 bl[66] br[66] wl[163] vdd gnd cell_6t
Xbit_r164_c66 bl[66] br[66] wl[164] vdd gnd cell_6t
Xbit_r165_c66 bl[66] br[66] wl[165] vdd gnd cell_6t
Xbit_r166_c66 bl[66] br[66] wl[166] vdd gnd cell_6t
Xbit_r167_c66 bl[66] br[66] wl[167] vdd gnd cell_6t
Xbit_r168_c66 bl[66] br[66] wl[168] vdd gnd cell_6t
Xbit_r169_c66 bl[66] br[66] wl[169] vdd gnd cell_6t
Xbit_r170_c66 bl[66] br[66] wl[170] vdd gnd cell_6t
Xbit_r171_c66 bl[66] br[66] wl[171] vdd gnd cell_6t
Xbit_r172_c66 bl[66] br[66] wl[172] vdd gnd cell_6t
Xbit_r173_c66 bl[66] br[66] wl[173] vdd gnd cell_6t
Xbit_r174_c66 bl[66] br[66] wl[174] vdd gnd cell_6t
Xbit_r175_c66 bl[66] br[66] wl[175] vdd gnd cell_6t
Xbit_r176_c66 bl[66] br[66] wl[176] vdd gnd cell_6t
Xbit_r177_c66 bl[66] br[66] wl[177] vdd gnd cell_6t
Xbit_r178_c66 bl[66] br[66] wl[178] vdd gnd cell_6t
Xbit_r179_c66 bl[66] br[66] wl[179] vdd gnd cell_6t
Xbit_r180_c66 bl[66] br[66] wl[180] vdd gnd cell_6t
Xbit_r181_c66 bl[66] br[66] wl[181] vdd gnd cell_6t
Xbit_r182_c66 bl[66] br[66] wl[182] vdd gnd cell_6t
Xbit_r183_c66 bl[66] br[66] wl[183] vdd gnd cell_6t
Xbit_r184_c66 bl[66] br[66] wl[184] vdd gnd cell_6t
Xbit_r185_c66 bl[66] br[66] wl[185] vdd gnd cell_6t
Xbit_r186_c66 bl[66] br[66] wl[186] vdd gnd cell_6t
Xbit_r187_c66 bl[66] br[66] wl[187] vdd gnd cell_6t
Xbit_r188_c66 bl[66] br[66] wl[188] vdd gnd cell_6t
Xbit_r189_c66 bl[66] br[66] wl[189] vdd gnd cell_6t
Xbit_r190_c66 bl[66] br[66] wl[190] vdd gnd cell_6t
Xbit_r191_c66 bl[66] br[66] wl[191] vdd gnd cell_6t
Xbit_r192_c66 bl[66] br[66] wl[192] vdd gnd cell_6t
Xbit_r193_c66 bl[66] br[66] wl[193] vdd gnd cell_6t
Xbit_r194_c66 bl[66] br[66] wl[194] vdd gnd cell_6t
Xbit_r195_c66 bl[66] br[66] wl[195] vdd gnd cell_6t
Xbit_r196_c66 bl[66] br[66] wl[196] vdd gnd cell_6t
Xbit_r197_c66 bl[66] br[66] wl[197] vdd gnd cell_6t
Xbit_r198_c66 bl[66] br[66] wl[198] vdd gnd cell_6t
Xbit_r199_c66 bl[66] br[66] wl[199] vdd gnd cell_6t
Xbit_r200_c66 bl[66] br[66] wl[200] vdd gnd cell_6t
Xbit_r201_c66 bl[66] br[66] wl[201] vdd gnd cell_6t
Xbit_r202_c66 bl[66] br[66] wl[202] vdd gnd cell_6t
Xbit_r203_c66 bl[66] br[66] wl[203] vdd gnd cell_6t
Xbit_r204_c66 bl[66] br[66] wl[204] vdd gnd cell_6t
Xbit_r205_c66 bl[66] br[66] wl[205] vdd gnd cell_6t
Xbit_r206_c66 bl[66] br[66] wl[206] vdd gnd cell_6t
Xbit_r207_c66 bl[66] br[66] wl[207] vdd gnd cell_6t
Xbit_r208_c66 bl[66] br[66] wl[208] vdd gnd cell_6t
Xbit_r209_c66 bl[66] br[66] wl[209] vdd gnd cell_6t
Xbit_r210_c66 bl[66] br[66] wl[210] vdd gnd cell_6t
Xbit_r211_c66 bl[66] br[66] wl[211] vdd gnd cell_6t
Xbit_r212_c66 bl[66] br[66] wl[212] vdd gnd cell_6t
Xbit_r213_c66 bl[66] br[66] wl[213] vdd gnd cell_6t
Xbit_r214_c66 bl[66] br[66] wl[214] vdd gnd cell_6t
Xbit_r215_c66 bl[66] br[66] wl[215] vdd gnd cell_6t
Xbit_r216_c66 bl[66] br[66] wl[216] vdd gnd cell_6t
Xbit_r217_c66 bl[66] br[66] wl[217] vdd gnd cell_6t
Xbit_r218_c66 bl[66] br[66] wl[218] vdd gnd cell_6t
Xbit_r219_c66 bl[66] br[66] wl[219] vdd gnd cell_6t
Xbit_r220_c66 bl[66] br[66] wl[220] vdd gnd cell_6t
Xbit_r221_c66 bl[66] br[66] wl[221] vdd gnd cell_6t
Xbit_r222_c66 bl[66] br[66] wl[222] vdd gnd cell_6t
Xbit_r223_c66 bl[66] br[66] wl[223] vdd gnd cell_6t
Xbit_r224_c66 bl[66] br[66] wl[224] vdd gnd cell_6t
Xbit_r225_c66 bl[66] br[66] wl[225] vdd gnd cell_6t
Xbit_r226_c66 bl[66] br[66] wl[226] vdd gnd cell_6t
Xbit_r227_c66 bl[66] br[66] wl[227] vdd gnd cell_6t
Xbit_r228_c66 bl[66] br[66] wl[228] vdd gnd cell_6t
Xbit_r229_c66 bl[66] br[66] wl[229] vdd gnd cell_6t
Xbit_r230_c66 bl[66] br[66] wl[230] vdd gnd cell_6t
Xbit_r231_c66 bl[66] br[66] wl[231] vdd gnd cell_6t
Xbit_r232_c66 bl[66] br[66] wl[232] vdd gnd cell_6t
Xbit_r233_c66 bl[66] br[66] wl[233] vdd gnd cell_6t
Xbit_r234_c66 bl[66] br[66] wl[234] vdd gnd cell_6t
Xbit_r235_c66 bl[66] br[66] wl[235] vdd gnd cell_6t
Xbit_r236_c66 bl[66] br[66] wl[236] vdd gnd cell_6t
Xbit_r237_c66 bl[66] br[66] wl[237] vdd gnd cell_6t
Xbit_r238_c66 bl[66] br[66] wl[238] vdd gnd cell_6t
Xbit_r239_c66 bl[66] br[66] wl[239] vdd gnd cell_6t
Xbit_r240_c66 bl[66] br[66] wl[240] vdd gnd cell_6t
Xbit_r241_c66 bl[66] br[66] wl[241] vdd gnd cell_6t
Xbit_r242_c66 bl[66] br[66] wl[242] vdd gnd cell_6t
Xbit_r243_c66 bl[66] br[66] wl[243] vdd gnd cell_6t
Xbit_r244_c66 bl[66] br[66] wl[244] vdd gnd cell_6t
Xbit_r245_c66 bl[66] br[66] wl[245] vdd gnd cell_6t
Xbit_r246_c66 bl[66] br[66] wl[246] vdd gnd cell_6t
Xbit_r247_c66 bl[66] br[66] wl[247] vdd gnd cell_6t
Xbit_r248_c66 bl[66] br[66] wl[248] vdd gnd cell_6t
Xbit_r249_c66 bl[66] br[66] wl[249] vdd gnd cell_6t
Xbit_r250_c66 bl[66] br[66] wl[250] vdd gnd cell_6t
Xbit_r251_c66 bl[66] br[66] wl[251] vdd gnd cell_6t
Xbit_r252_c66 bl[66] br[66] wl[252] vdd gnd cell_6t
Xbit_r253_c66 bl[66] br[66] wl[253] vdd gnd cell_6t
Xbit_r254_c66 bl[66] br[66] wl[254] vdd gnd cell_6t
Xbit_r255_c66 bl[66] br[66] wl[255] vdd gnd cell_6t
Xbit_r0_c67 bl[67] br[67] wl[0] vdd gnd cell_6t
Xbit_r1_c67 bl[67] br[67] wl[1] vdd gnd cell_6t
Xbit_r2_c67 bl[67] br[67] wl[2] vdd gnd cell_6t
Xbit_r3_c67 bl[67] br[67] wl[3] vdd gnd cell_6t
Xbit_r4_c67 bl[67] br[67] wl[4] vdd gnd cell_6t
Xbit_r5_c67 bl[67] br[67] wl[5] vdd gnd cell_6t
Xbit_r6_c67 bl[67] br[67] wl[6] vdd gnd cell_6t
Xbit_r7_c67 bl[67] br[67] wl[7] vdd gnd cell_6t
Xbit_r8_c67 bl[67] br[67] wl[8] vdd gnd cell_6t
Xbit_r9_c67 bl[67] br[67] wl[9] vdd gnd cell_6t
Xbit_r10_c67 bl[67] br[67] wl[10] vdd gnd cell_6t
Xbit_r11_c67 bl[67] br[67] wl[11] vdd gnd cell_6t
Xbit_r12_c67 bl[67] br[67] wl[12] vdd gnd cell_6t
Xbit_r13_c67 bl[67] br[67] wl[13] vdd gnd cell_6t
Xbit_r14_c67 bl[67] br[67] wl[14] vdd gnd cell_6t
Xbit_r15_c67 bl[67] br[67] wl[15] vdd gnd cell_6t
Xbit_r16_c67 bl[67] br[67] wl[16] vdd gnd cell_6t
Xbit_r17_c67 bl[67] br[67] wl[17] vdd gnd cell_6t
Xbit_r18_c67 bl[67] br[67] wl[18] vdd gnd cell_6t
Xbit_r19_c67 bl[67] br[67] wl[19] vdd gnd cell_6t
Xbit_r20_c67 bl[67] br[67] wl[20] vdd gnd cell_6t
Xbit_r21_c67 bl[67] br[67] wl[21] vdd gnd cell_6t
Xbit_r22_c67 bl[67] br[67] wl[22] vdd gnd cell_6t
Xbit_r23_c67 bl[67] br[67] wl[23] vdd gnd cell_6t
Xbit_r24_c67 bl[67] br[67] wl[24] vdd gnd cell_6t
Xbit_r25_c67 bl[67] br[67] wl[25] vdd gnd cell_6t
Xbit_r26_c67 bl[67] br[67] wl[26] vdd gnd cell_6t
Xbit_r27_c67 bl[67] br[67] wl[27] vdd gnd cell_6t
Xbit_r28_c67 bl[67] br[67] wl[28] vdd gnd cell_6t
Xbit_r29_c67 bl[67] br[67] wl[29] vdd gnd cell_6t
Xbit_r30_c67 bl[67] br[67] wl[30] vdd gnd cell_6t
Xbit_r31_c67 bl[67] br[67] wl[31] vdd gnd cell_6t
Xbit_r32_c67 bl[67] br[67] wl[32] vdd gnd cell_6t
Xbit_r33_c67 bl[67] br[67] wl[33] vdd gnd cell_6t
Xbit_r34_c67 bl[67] br[67] wl[34] vdd gnd cell_6t
Xbit_r35_c67 bl[67] br[67] wl[35] vdd gnd cell_6t
Xbit_r36_c67 bl[67] br[67] wl[36] vdd gnd cell_6t
Xbit_r37_c67 bl[67] br[67] wl[37] vdd gnd cell_6t
Xbit_r38_c67 bl[67] br[67] wl[38] vdd gnd cell_6t
Xbit_r39_c67 bl[67] br[67] wl[39] vdd gnd cell_6t
Xbit_r40_c67 bl[67] br[67] wl[40] vdd gnd cell_6t
Xbit_r41_c67 bl[67] br[67] wl[41] vdd gnd cell_6t
Xbit_r42_c67 bl[67] br[67] wl[42] vdd gnd cell_6t
Xbit_r43_c67 bl[67] br[67] wl[43] vdd gnd cell_6t
Xbit_r44_c67 bl[67] br[67] wl[44] vdd gnd cell_6t
Xbit_r45_c67 bl[67] br[67] wl[45] vdd gnd cell_6t
Xbit_r46_c67 bl[67] br[67] wl[46] vdd gnd cell_6t
Xbit_r47_c67 bl[67] br[67] wl[47] vdd gnd cell_6t
Xbit_r48_c67 bl[67] br[67] wl[48] vdd gnd cell_6t
Xbit_r49_c67 bl[67] br[67] wl[49] vdd gnd cell_6t
Xbit_r50_c67 bl[67] br[67] wl[50] vdd gnd cell_6t
Xbit_r51_c67 bl[67] br[67] wl[51] vdd gnd cell_6t
Xbit_r52_c67 bl[67] br[67] wl[52] vdd gnd cell_6t
Xbit_r53_c67 bl[67] br[67] wl[53] vdd gnd cell_6t
Xbit_r54_c67 bl[67] br[67] wl[54] vdd gnd cell_6t
Xbit_r55_c67 bl[67] br[67] wl[55] vdd gnd cell_6t
Xbit_r56_c67 bl[67] br[67] wl[56] vdd gnd cell_6t
Xbit_r57_c67 bl[67] br[67] wl[57] vdd gnd cell_6t
Xbit_r58_c67 bl[67] br[67] wl[58] vdd gnd cell_6t
Xbit_r59_c67 bl[67] br[67] wl[59] vdd gnd cell_6t
Xbit_r60_c67 bl[67] br[67] wl[60] vdd gnd cell_6t
Xbit_r61_c67 bl[67] br[67] wl[61] vdd gnd cell_6t
Xbit_r62_c67 bl[67] br[67] wl[62] vdd gnd cell_6t
Xbit_r63_c67 bl[67] br[67] wl[63] vdd gnd cell_6t
Xbit_r64_c67 bl[67] br[67] wl[64] vdd gnd cell_6t
Xbit_r65_c67 bl[67] br[67] wl[65] vdd gnd cell_6t
Xbit_r66_c67 bl[67] br[67] wl[66] vdd gnd cell_6t
Xbit_r67_c67 bl[67] br[67] wl[67] vdd gnd cell_6t
Xbit_r68_c67 bl[67] br[67] wl[68] vdd gnd cell_6t
Xbit_r69_c67 bl[67] br[67] wl[69] vdd gnd cell_6t
Xbit_r70_c67 bl[67] br[67] wl[70] vdd gnd cell_6t
Xbit_r71_c67 bl[67] br[67] wl[71] vdd gnd cell_6t
Xbit_r72_c67 bl[67] br[67] wl[72] vdd gnd cell_6t
Xbit_r73_c67 bl[67] br[67] wl[73] vdd gnd cell_6t
Xbit_r74_c67 bl[67] br[67] wl[74] vdd gnd cell_6t
Xbit_r75_c67 bl[67] br[67] wl[75] vdd gnd cell_6t
Xbit_r76_c67 bl[67] br[67] wl[76] vdd gnd cell_6t
Xbit_r77_c67 bl[67] br[67] wl[77] vdd gnd cell_6t
Xbit_r78_c67 bl[67] br[67] wl[78] vdd gnd cell_6t
Xbit_r79_c67 bl[67] br[67] wl[79] vdd gnd cell_6t
Xbit_r80_c67 bl[67] br[67] wl[80] vdd gnd cell_6t
Xbit_r81_c67 bl[67] br[67] wl[81] vdd gnd cell_6t
Xbit_r82_c67 bl[67] br[67] wl[82] vdd gnd cell_6t
Xbit_r83_c67 bl[67] br[67] wl[83] vdd gnd cell_6t
Xbit_r84_c67 bl[67] br[67] wl[84] vdd gnd cell_6t
Xbit_r85_c67 bl[67] br[67] wl[85] vdd gnd cell_6t
Xbit_r86_c67 bl[67] br[67] wl[86] vdd gnd cell_6t
Xbit_r87_c67 bl[67] br[67] wl[87] vdd gnd cell_6t
Xbit_r88_c67 bl[67] br[67] wl[88] vdd gnd cell_6t
Xbit_r89_c67 bl[67] br[67] wl[89] vdd gnd cell_6t
Xbit_r90_c67 bl[67] br[67] wl[90] vdd gnd cell_6t
Xbit_r91_c67 bl[67] br[67] wl[91] vdd gnd cell_6t
Xbit_r92_c67 bl[67] br[67] wl[92] vdd gnd cell_6t
Xbit_r93_c67 bl[67] br[67] wl[93] vdd gnd cell_6t
Xbit_r94_c67 bl[67] br[67] wl[94] vdd gnd cell_6t
Xbit_r95_c67 bl[67] br[67] wl[95] vdd gnd cell_6t
Xbit_r96_c67 bl[67] br[67] wl[96] vdd gnd cell_6t
Xbit_r97_c67 bl[67] br[67] wl[97] vdd gnd cell_6t
Xbit_r98_c67 bl[67] br[67] wl[98] vdd gnd cell_6t
Xbit_r99_c67 bl[67] br[67] wl[99] vdd gnd cell_6t
Xbit_r100_c67 bl[67] br[67] wl[100] vdd gnd cell_6t
Xbit_r101_c67 bl[67] br[67] wl[101] vdd gnd cell_6t
Xbit_r102_c67 bl[67] br[67] wl[102] vdd gnd cell_6t
Xbit_r103_c67 bl[67] br[67] wl[103] vdd gnd cell_6t
Xbit_r104_c67 bl[67] br[67] wl[104] vdd gnd cell_6t
Xbit_r105_c67 bl[67] br[67] wl[105] vdd gnd cell_6t
Xbit_r106_c67 bl[67] br[67] wl[106] vdd gnd cell_6t
Xbit_r107_c67 bl[67] br[67] wl[107] vdd gnd cell_6t
Xbit_r108_c67 bl[67] br[67] wl[108] vdd gnd cell_6t
Xbit_r109_c67 bl[67] br[67] wl[109] vdd gnd cell_6t
Xbit_r110_c67 bl[67] br[67] wl[110] vdd gnd cell_6t
Xbit_r111_c67 bl[67] br[67] wl[111] vdd gnd cell_6t
Xbit_r112_c67 bl[67] br[67] wl[112] vdd gnd cell_6t
Xbit_r113_c67 bl[67] br[67] wl[113] vdd gnd cell_6t
Xbit_r114_c67 bl[67] br[67] wl[114] vdd gnd cell_6t
Xbit_r115_c67 bl[67] br[67] wl[115] vdd gnd cell_6t
Xbit_r116_c67 bl[67] br[67] wl[116] vdd gnd cell_6t
Xbit_r117_c67 bl[67] br[67] wl[117] vdd gnd cell_6t
Xbit_r118_c67 bl[67] br[67] wl[118] vdd gnd cell_6t
Xbit_r119_c67 bl[67] br[67] wl[119] vdd gnd cell_6t
Xbit_r120_c67 bl[67] br[67] wl[120] vdd gnd cell_6t
Xbit_r121_c67 bl[67] br[67] wl[121] vdd gnd cell_6t
Xbit_r122_c67 bl[67] br[67] wl[122] vdd gnd cell_6t
Xbit_r123_c67 bl[67] br[67] wl[123] vdd gnd cell_6t
Xbit_r124_c67 bl[67] br[67] wl[124] vdd gnd cell_6t
Xbit_r125_c67 bl[67] br[67] wl[125] vdd gnd cell_6t
Xbit_r126_c67 bl[67] br[67] wl[126] vdd gnd cell_6t
Xbit_r127_c67 bl[67] br[67] wl[127] vdd gnd cell_6t
Xbit_r128_c67 bl[67] br[67] wl[128] vdd gnd cell_6t
Xbit_r129_c67 bl[67] br[67] wl[129] vdd gnd cell_6t
Xbit_r130_c67 bl[67] br[67] wl[130] vdd gnd cell_6t
Xbit_r131_c67 bl[67] br[67] wl[131] vdd gnd cell_6t
Xbit_r132_c67 bl[67] br[67] wl[132] vdd gnd cell_6t
Xbit_r133_c67 bl[67] br[67] wl[133] vdd gnd cell_6t
Xbit_r134_c67 bl[67] br[67] wl[134] vdd gnd cell_6t
Xbit_r135_c67 bl[67] br[67] wl[135] vdd gnd cell_6t
Xbit_r136_c67 bl[67] br[67] wl[136] vdd gnd cell_6t
Xbit_r137_c67 bl[67] br[67] wl[137] vdd gnd cell_6t
Xbit_r138_c67 bl[67] br[67] wl[138] vdd gnd cell_6t
Xbit_r139_c67 bl[67] br[67] wl[139] vdd gnd cell_6t
Xbit_r140_c67 bl[67] br[67] wl[140] vdd gnd cell_6t
Xbit_r141_c67 bl[67] br[67] wl[141] vdd gnd cell_6t
Xbit_r142_c67 bl[67] br[67] wl[142] vdd gnd cell_6t
Xbit_r143_c67 bl[67] br[67] wl[143] vdd gnd cell_6t
Xbit_r144_c67 bl[67] br[67] wl[144] vdd gnd cell_6t
Xbit_r145_c67 bl[67] br[67] wl[145] vdd gnd cell_6t
Xbit_r146_c67 bl[67] br[67] wl[146] vdd gnd cell_6t
Xbit_r147_c67 bl[67] br[67] wl[147] vdd gnd cell_6t
Xbit_r148_c67 bl[67] br[67] wl[148] vdd gnd cell_6t
Xbit_r149_c67 bl[67] br[67] wl[149] vdd gnd cell_6t
Xbit_r150_c67 bl[67] br[67] wl[150] vdd gnd cell_6t
Xbit_r151_c67 bl[67] br[67] wl[151] vdd gnd cell_6t
Xbit_r152_c67 bl[67] br[67] wl[152] vdd gnd cell_6t
Xbit_r153_c67 bl[67] br[67] wl[153] vdd gnd cell_6t
Xbit_r154_c67 bl[67] br[67] wl[154] vdd gnd cell_6t
Xbit_r155_c67 bl[67] br[67] wl[155] vdd gnd cell_6t
Xbit_r156_c67 bl[67] br[67] wl[156] vdd gnd cell_6t
Xbit_r157_c67 bl[67] br[67] wl[157] vdd gnd cell_6t
Xbit_r158_c67 bl[67] br[67] wl[158] vdd gnd cell_6t
Xbit_r159_c67 bl[67] br[67] wl[159] vdd gnd cell_6t
Xbit_r160_c67 bl[67] br[67] wl[160] vdd gnd cell_6t
Xbit_r161_c67 bl[67] br[67] wl[161] vdd gnd cell_6t
Xbit_r162_c67 bl[67] br[67] wl[162] vdd gnd cell_6t
Xbit_r163_c67 bl[67] br[67] wl[163] vdd gnd cell_6t
Xbit_r164_c67 bl[67] br[67] wl[164] vdd gnd cell_6t
Xbit_r165_c67 bl[67] br[67] wl[165] vdd gnd cell_6t
Xbit_r166_c67 bl[67] br[67] wl[166] vdd gnd cell_6t
Xbit_r167_c67 bl[67] br[67] wl[167] vdd gnd cell_6t
Xbit_r168_c67 bl[67] br[67] wl[168] vdd gnd cell_6t
Xbit_r169_c67 bl[67] br[67] wl[169] vdd gnd cell_6t
Xbit_r170_c67 bl[67] br[67] wl[170] vdd gnd cell_6t
Xbit_r171_c67 bl[67] br[67] wl[171] vdd gnd cell_6t
Xbit_r172_c67 bl[67] br[67] wl[172] vdd gnd cell_6t
Xbit_r173_c67 bl[67] br[67] wl[173] vdd gnd cell_6t
Xbit_r174_c67 bl[67] br[67] wl[174] vdd gnd cell_6t
Xbit_r175_c67 bl[67] br[67] wl[175] vdd gnd cell_6t
Xbit_r176_c67 bl[67] br[67] wl[176] vdd gnd cell_6t
Xbit_r177_c67 bl[67] br[67] wl[177] vdd gnd cell_6t
Xbit_r178_c67 bl[67] br[67] wl[178] vdd gnd cell_6t
Xbit_r179_c67 bl[67] br[67] wl[179] vdd gnd cell_6t
Xbit_r180_c67 bl[67] br[67] wl[180] vdd gnd cell_6t
Xbit_r181_c67 bl[67] br[67] wl[181] vdd gnd cell_6t
Xbit_r182_c67 bl[67] br[67] wl[182] vdd gnd cell_6t
Xbit_r183_c67 bl[67] br[67] wl[183] vdd gnd cell_6t
Xbit_r184_c67 bl[67] br[67] wl[184] vdd gnd cell_6t
Xbit_r185_c67 bl[67] br[67] wl[185] vdd gnd cell_6t
Xbit_r186_c67 bl[67] br[67] wl[186] vdd gnd cell_6t
Xbit_r187_c67 bl[67] br[67] wl[187] vdd gnd cell_6t
Xbit_r188_c67 bl[67] br[67] wl[188] vdd gnd cell_6t
Xbit_r189_c67 bl[67] br[67] wl[189] vdd gnd cell_6t
Xbit_r190_c67 bl[67] br[67] wl[190] vdd gnd cell_6t
Xbit_r191_c67 bl[67] br[67] wl[191] vdd gnd cell_6t
Xbit_r192_c67 bl[67] br[67] wl[192] vdd gnd cell_6t
Xbit_r193_c67 bl[67] br[67] wl[193] vdd gnd cell_6t
Xbit_r194_c67 bl[67] br[67] wl[194] vdd gnd cell_6t
Xbit_r195_c67 bl[67] br[67] wl[195] vdd gnd cell_6t
Xbit_r196_c67 bl[67] br[67] wl[196] vdd gnd cell_6t
Xbit_r197_c67 bl[67] br[67] wl[197] vdd gnd cell_6t
Xbit_r198_c67 bl[67] br[67] wl[198] vdd gnd cell_6t
Xbit_r199_c67 bl[67] br[67] wl[199] vdd gnd cell_6t
Xbit_r200_c67 bl[67] br[67] wl[200] vdd gnd cell_6t
Xbit_r201_c67 bl[67] br[67] wl[201] vdd gnd cell_6t
Xbit_r202_c67 bl[67] br[67] wl[202] vdd gnd cell_6t
Xbit_r203_c67 bl[67] br[67] wl[203] vdd gnd cell_6t
Xbit_r204_c67 bl[67] br[67] wl[204] vdd gnd cell_6t
Xbit_r205_c67 bl[67] br[67] wl[205] vdd gnd cell_6t
Xbit_r206_c67 bl[67] br[67] wl[206] vdd gnd cell_6t
Xbit_r207_c67 bl[67] br[67] wl[207] vdd gnd cell_6t
Xbit_r208_c67 bl[67] br[67] wl[208] vdd gnd cell_6t
Xbit_r209_c67 bl[67] br[67] wl[209] vdd gnd cell_6t
Xbit_r210_c67 bl[67] br[67] wl[210] vdd gnd cell_6t
Xbit_r211_c67 bl[67] br[67] wl[211] vdd gnd cell_6t
Xbit_r212_c67 bl[67] br[67] wl[212] vdd gnd cell_6t
Xbit_r213_c67 bl[67] br[67] wl[213] vdd gnd cell_6t
Xbit_r214_c67 bl[67] br[67] wl[214] vdd gnd cell_6t
Xbit_r215_c67 bl[67] br[67] wl[215] vdd gnd cell_6t
Xbit_r216_c67 bl[67] br[67] wl[216] vdd gnd cell_6t
Xbit_r217_c67 bl[67] br[67] wl[217] vdd gnd cell_6t
Xbit_r218_c67 bl[67] br[67] wl[218] vdd gnd cell_6t
Xbit_r219_c67 bl[67] br[67] wl[219] vdd gnd cell_6t
Xbit_r220_c67 bl[67] br[67] wl[220] vdd gnd cell_6t
Xbit_r221_c67 bl[67] br[67] wl[221] vdd gnd cell_6t
Xbit_r222_c67 bl[67] br[67] wl[222] vdd gnd cell_6t
Xbit_r223_c67 bl[67] br[67] wl[223] vdd gnd cell_6t
Xbit_r224_c67 bl[67] br[67] wl[224] vdd gnd cell_6t
Xbit_r225_c67 bl[67] br[67] wl[225] vdd gnd cell_6t
Xbit_r226_c67 bl[67] br[67] wl[226] vdd gnd cell_6t
Xbit_r227_c67 bl[67] br[67] wl[227] vdd gnd cell_6t
Xbit_r228_c67 bl[67] br[67] wl[228] vdd gnd cell_6t
Xbit_r229_c67 bl[67] br[67] wl[229] vdd gnd cell_6t
Xbit_r230_c67 bl[67] br[67] wl[230] vdd gnd cell_6t
Xbit_r231_c67 bl[67] br[67] wl[231] vdd gnd cell_6t
Xbit_r232_c67 bl[67] br[67] wl[232] vdd gnd cell_6t
Xbit_r233_c67 bl[67] br[67] wl[233] vdd gnd cell_6t
Xbit_r234_c67 bl[67] br[67] wl[234] vdd gnd cell_6t
Xbit_r235_c67 bl[67] br[67] wl[235] vdd gnd cell_6t
Xbit_r236_c67 bl[67] br[67] wl[236] vdd gnd cell_6t
Xbit_r237_c67 bl[67] br[67] wl[237] vdd gnd cell_6t
Xbit_r238_c67 bl[67] br[67] wl[238] vdd gnd cell_6t
Xbit_r239_c67 bl[67] br[67] wl[239] vdd gnd cell_6t
Xbit_r240_c67 bl[67] br[67] wl[240] vdd gnd cell_6t
Xbit_r241_c67 bl[67] br[67] wl[241] vdd gnd cell_6t
Xbit_r242_c67 bl[67] br[67] wl[242] vdd gnd cell_6t
Xbit_r243_c67 bl[67] br[67] wl[243] vdd gnd cell_6t
Xbit_r244_c67 bl[67] br[67] wl[244] vdd gnd cell_6t
Xbit_r245_c67 bl[67] br[67] wl[245] vdd gnd cell_6t
Xbit_r246_c67 bl[67] br[67] wl[246] vdd gnd cell_6t
Xbit_r247_c67 bl[67] br[67] wl[247] vdd gnd cell_6t
Xbit_r248_c67 bl[67] br[67] wl[248] vdd gnd cell_6t
Xbit_r249_c67 bl[67] br[67] wl[249] vdd gnd cell_6t
Xbit_r250_c67 bl[67] br[67] wl[250] vdd gnd cell_6t
Xbit_r251_c67 bl[67] br[67] wl[251] vdd gnd cell_6t
Xbit_r252_c67 bl[67] br[67] wl[252] vdd gnd cell_6t
Xbit_r253_c67 bl[67] br[67] wl[253] vdd gnd cell_6t
Xbit_r254_c67 bl[67] br[67] wl[254] vdd gnd cell_6t
Xbit_r255_c67 bl[67] br[67] wl[255] vdd gnd cell_6t
Xbit_r0_c68 bl[68] br[68] wl[0] vdd gnd cell_6t
Xbit_r1_c68 bl[68] br[68] wl[1] vdd gnd cell_6t
Xbit_r2_c68 bl[68] br[68] wl[2] vdd gnd cell_6t
Xbit_r3_c68 bl[68] br[68] wl[3] vdd gnd cell_6t
Xbit_r4_c68 bl[68] br[68] wl[4] vdd gnd cell_6t
Xbit_r5_c68 bl[68] br[68] wl[5] vdd gnd cell_6t
Xbit_r6_c68 bl[68] br[68] wl[6] vdd gnd cell_6t
Xbit_r7_c68 bl[68] br[68] wl[7] vdd gnd cell_6t
Xbit_r8_c68 bl[68] br[68] wl[8] vdd gnd cell_6t
Xbit_r9_c68 bl[68] br[68] wl[9] vdd gnd cell_6t
Xbit_r10_c68 bl[68] br[68] wl[10] vdd gnd cell_6t
Xbit_r11_c68 bl[68] br[68] wl[11] vdd gnd cell_6t
Xbit_r12_c68 bl[68] br[68] wl[12] vdd gnd cell_6t
Xbit_r13_c68 bl[68] br[68] wl[13] vdd gnd cell_6t
Xbit_r14_c68 bl[68] br[68] wl[14] vdd gnd cell_6t
Xbit_r15_c68 bl[68] br[68] wl[15] vdd gnd cell_6t
Xbit_r16_c68 bl[68] br[68] wl[16] vdd gnd cell_6t
Xbit_r17_c68 bl[68] br[68] wl[17] vdd gnd cell_6t
Xbit_r18_c68 bl[68] br[68] wl[18] vdd gnd cell_6t
Xbit_r19_c68 bl[68] br[68] wl[19] vdd gnd cell_6t
Xbit_r20_c68 bl[68] br[68] wl[20] vdd gnd cell_6t
Xbit_r21_c68 bl[68] br[68] wl[21] vdd gnd cell_6t
Xbit_r22_c68 bl[68] br[68] wl[22] vdd gnd cell_6t
Xbit_r23_c68 bl[68] br[68] wl[23] vdd gnd cell_6t
Xbit_r24_c68 bl[68] br[68] wl[24] vdd gnd cell_6t
Xbit_r25_c68 bl[68] br[68] wl[25] vdd gnd cell_6t
Xbit_r26_c68 bl[68] br[68] wl[26] vdd gnd cell_6t
Xbit_r27_c68 bl[68] br[68] wl[27] vdd gnd cell_6t
Xbit_r28_c68 bl[68] br[68] wl[28] vdd gnd cell_6t
Xbit_r29_c68 bl[68] br[68] wl[29] vdd gnd cell_6t
Xbit_r30_c68 bl[68] br[68] wl[30] vdd gnd cell_6t
Xbit_r31_c68 bl[68] br[68] wl[31] vdd gnd cell_6t
Xbit_r32_c68 bl[68] br[68] wl[32] vdd gnd cell_6t
Xbit_r33_c68 bl[68] br[68] wl[33] vdd gnd cell_6t
Xbit_r34_c68 bl[68] br[68] wl[34] vdd gnd cell_6t
Xbit_r35_c68 bl[68] br[68] wl[35] vdd gnd cell_6t
Xbit_r36_c68 bl[68] br[68] wl[36] vdd gnd cell_6t
Xbit_r37_c68 bl[68] br[68] wl[37] vdd gnd cell_6t
Xbit_r38_c68 bl[68] br[68] wl[38] vdd gnd cell_6t
Xbit_r39_c68 bl[68] br[68] wl[39] vdd gnd cell_6t
Xbit_r40_c68 bl[68] br[68] wl[40] vdd gnd cell_6t
Xbit_r41_c68 bl[68] br[68] wl[41] vdd gnd cell_6t
Xbit_r42_c68 bl[68] br[68] wl[42] vdd gnd cell_6t
Xbit_r43_c68 bl[68] br[68] wl[43] vdd gnd cell_6t
Xbit_r44_c68 bl[68] br[68] wl[44] vdd gnd cell_6t
Xbit_r45_c68 bl[68] br[68] wl[45] vdd gnd cell_6t
Xbit_r46_c68 bl[68] br[68] wl[46] vdd gnd cell_6t
Xbit_r47_c68 bl[68] br[68] wl[47] vdd gnd cell_6t
Xbit_r48_c68 bl[68] br[68] wl[48] vdd gnd cell_6t
Xbit_r49_c68 bl[68] br[68] wl[49] vdd gnd cell_6t
Xbit_r50_c68 bl[68] br[68] wl[50] vdd gnd cell_6t
Xbit_r51_c68 bl[68] br[68] wl[51] vdd gnd cell_6t
Xbit_r52_c68 bl[68] br[68] wl[52] vdd gnd cell_6t
Xbit_r53_c68 bl[68] br[68] wl[53] vdd gnd cell_6t
Xbit_r54_c68 bl[68] br[68] wl[54] vdd gnd cell_6t
Xbit_r55_c68 bl[68] br[68] wl[55] vdd gnd cell_6t
Xbit_r56_c68 bl[68] br[68] wl[56] vdd gnd cell_6t
Xbit_r57_c68 bl[68] br[68] wl[57] vdd gnd cell_6t
Xbit_r58_c68 bl[68] br[68] wl[58] vdd gnd cell_6t
Xbit_r59_c68 bl[68] br[68] wl[59] vdd gnd cell_6t
Xbit_r60_c68 bl[68] br[68] wl[60] vdd gnd cell_6t
Xbit_r61_c68 bl[68] br[68] wl[61] vdd gnd cell_6t
Xbit_r62_c68 bl[68] br[68] wl[62] vdd gnd cell_6t
Xbit_r63_c68 bl[68] br[68] wl[63] vdd gnd cell_6t
Xbit_r64_c68 bl[68] br[68] wl[64] vdd gnd cell_6t
Xbit_r65_c68 bl[68] br[68] wl[65] vdd gnd cell_6t
Xbit_r66_c68 bl[68] br[68] wl[66] vdd gnd cell_6t
Xbit_r67_c68 bl[68] br[68] wl[67] vdd gnd cell_6t
Xbit_r68_c68 bl[68] br[68] wl[68] vdd gnd cell_6t
Xbit_r69_c68 bl[68] br[68] wl[69] vdd gnd cell_6t
Xbit_r70_c68 bl[68] br[68] wl[70] vdd gnd cell_6t
Xbit_r71_c68 bl[68] br[68] wl[71] vdd gnd cell_6t
Xbit_r72_c68 bl[68] br[68] wl[72] vdd gnd cell_6t
Xbit_r73_c68 bl[68] br[68] wl[73] vdd gnd cell_6t
Xbit_r74_c68 bl[68] br[68] wl[74] vdd gnd cell_6t
Xbit_r75_c68 bl[68] br[68] wl[75] vdd gnd cell_6t
Xbit_r76_c68 bl[68] br[68] wl[76] vdd gnd cell_6t
Xbit_r77_c68 bl[68] br[68] wl[77] vdd gnd cell_6t
Xbit_r78_c68 bl[68] br[68] wl[78] vdd gnd cell_6t
Xbit_r79_c68 bl[68] br[68] wl[79] vdd gnd cell_6t
Xbit_r80_c68 bl[68] br[68] wl[80] vdd gnd cell_6t
Xbit_r81_c68 bl[68] br[68] wl[81] vdd gnd cell_6t
Xbit_r82_c68 bl[68] br[68] wl[82] vdd gnd cell_6t
Xbit_r83_c68 bl[68] br[68] wl[83] vdd gnd cell_6t
Xbit_r84_c68 bl[68] br[68] wl[84] vdd gnd cell_6t
Xbit_r85_c68 bl[68] br[68] wl[85] vdd gnd cell_6t
Xbit_r86_c68 bl[68] br[68] wl[86] vdd gnd cell_6t
Xbit_r87_c68 bl[68] br[68] wl[87] vdd gnd cell_6t
Xbit_r88_c68 bl[68] br[68] wl[88] vdd gnd cell_6t
Xbit_r89_c68 bl[68] br[68] wl[89] vdd gnd cell_6t
Xbit_r90_c68 bl[68] br[68] wl[90] vdd gnd cell_6t
Xbit_r91_c68 bl[68] br[68] wl[91] vdd gnd cell_6t
Xbit_r92_c68 bl[68] br[68] wl[92] vdd gnd cell_6t
Xbit_r93_c68 bl[68] br[68] wl[93] vdd gnd cell_6t
Xbit_r94_c68 bl[68] br[68] wl[94] vdd gnd cell_6t
Xbit_r95_c68 bl[68] br[68] wl[95] vdd gnd cell_6t
Xbit_r96_c68 bl[68] br[68] wl[96] vdd gnd cell_6t
Xbit_r97_c68 bl[68] br[68] wl[97] vdd gnd cell_6t
Xbit_r98_c68 bl[68] br[68] wl[98] vdd gnd cell_6t
Xbit_r99_c68 bl[68] br[68] wl[99] vdd gnd cell_6t
Xbit_r100_c68 bl[68] br[68] wl[100] vdd gnd cell_6t
Xbit_r101_c68 bl[68] br[68] wl[101] vdd gnd cell_6t
Xbit_r102_c68 bl[68] br[68] wl[102] vdd gnd cell_6t
Xbit_r103_c68 bl[68] br[68] wl[103] vdd gnd cell_6t
Xbit_r104_c68 bl[68] br[68] wl[104] vdd gnd cell_6t
Xbit_r105_c68 bl[68] br[68] wl[105] vdd gnd cell_6t
Xbit_r106_c68 bl[68] br[68] wl[106] vdd gnd cell_6t
Xbit_r107_c68 bl[68] br[68] wl[107] vdd gnd cell_6t
Xbit_r108_c68 bl[68] br[68] wl[108] vdd gnd cell_6t
Xbit_r109_c68 bl[68] br[68] wl[109] vdd gnd cell_6t
Xbit_r110_c68 bl[68] br[68] wl[110] vdd gnd cell_6t
Xbit_r111_c68 bl[68] br[68] wl[111] vdd gnd cell_6t
Xbit_r112_c68 bl[68] br[68] wl[112] vdd gnd cell_6t
Xbit_r113_c68 bl[68] br[68] wl[113] vdd gnd cell_6t
Xbit_r114_c68 bl[68] br[68] wl[114] vdd gnd cell_6t
Xbit_r115_c68 bl[68] br[68] wl[115] vdd gnd cell_6t
Xbit_r116_c68 bl[68] br[68] wl[116] vdd gnd cell_6t
Xbit_r117_c68 bl[68] br[68] wl[117] vdd gnd cell_6t
Xbit_r118_c68 bl[68] br[68] wl[118] vdd gnd cell_6t
Xbit_r119_c68 bl[68] br[68] wl[119] vdd gnd cell_6t
Xbit_r120_c68 bl[68] br[68] wl[120] vdd gnd cell_6t
Xbit_r121_c68 bl[68] br[68] wl[121] vdd gnd cell_6t
Xbit_r122_c68 bl[68] br[68] wl[122] vdd gnd cell_6t
Xbit_r123_c68 bl[68] br[68] wl[123] vdd gnd cell_6t
Xbit_r124_c68 bl[68] br[68] wl[124] vdd gnd cell_6t
Xbit_r125_c68 bl[68] br[68] wl[125] vdd gnd cell_6t
Xbit_r126_c68 bl[68] br[68] wl[126] vdd gnd cell_6t
Xbit_r127_c68 bl[68] br[68] wl[127] vdd gnd cell_6t
Xbit_r128_c68 bl[68] br[68] wl[128] vdd gnd cell_6t
Xbit_r129_c68 bl[68] br[68] wl[129] vdd gnd cell_6t
Xbit_r130_c68 bl[68] br[68] wl[130] vdd gnd cell_6t
Xbit_r131_c68 bl[68] br[68] wl[131] vdd gnd cell_6t
Xbit_r132_c68 bl[68] br[68] wl[132] vdd gnd cell_6t
Xbit_r133_c68 bl[68] br[68] wl[133] vdd gnd cell_6t
Xbit_r134_c68 bl[68] br[68] wl[134] vdd gnd cell_6t
Xbit_r135_c68 bl[68] br[68] wl[135] vdd gnd cell_6t
Xbit_r136_c68 bl[68] br[68] wl[136] vdd gnd cell_6t
Xbit_r137_c68 bl[68] br[68] wl[137] vdd gnd cell_6t
Xbit_r138_c68 bl[68] br[68] wl[138] vdd gnd cell_6t
Xbit_r139_c68 bl[68] br[68] wl[139] vdd gnd cell_6t
Xbit_r140_c68 bl[68] br[68] wl[140] vdd gnd cell_6t
Xbit_r141_c68 bl[68] br[68] wl[141] vdd gnd cell_6t
Xbit_r142_c68 bl[68] br[68] wl[142] vdd gnd cell_6t
Xbit_r143_c68 bl[68] br[68] wl[143] vdd gnd cell_6t
Xbit_r144_c68 bl[68] br[68] wl[144] vdd gnd cell_6t
Xbit_r145_c68 bl[68] br[68] wl[145] vdd gnd cell_6t
Xbit_r146_c68 bl[68] br[68] wl[146] vdd gnd cell_6t
Xbit_r147_c68 bl[68] br[68] wl[147] vdd gnd cell_6t
Xbit_r148_c68 bl[68] br[68] wl[148] vdd gnd cell_6t
Xbit_r149_c68 bl[68] br[68] wl[149] vdd gnd cell_6t
Xbit_r150_c68 bl[68] br[68] wl[150] vdd gnd cell_6t
Xbit_r151_c68 bl[68] br[68] wl[151] vdd gnd cell_6t
Xbit_r152_c68 bl[68] br[68] wl[152] vdd gnd cell_6t
Xbit_r153_c68 bl[68] br[68] wl[153] vdd gnd cell_6t
Xbit_r154_c68 bl[68] br[68] wl[154] vdd gnd cell_6t
Xbit_r155_c68 bl[68] br[68] wl[155] vdd gnd cell_6t
Xbit_r156_c68 bl[68] br[68] wl[156] vdd gnd cell_6t
Xbit_r157_c68 bl[68] br[68] wl[157] vdd gnd cell_6t
Xbit_r158_c68 bl[68] br[68] wl[158] vdd gnd cell_6t
Xbit_r159_c68 bl[68] br[68] wl[159] vdd gnd cell_6t
Xbit_r160_c68 bl[68] br[68] wl[160] vdd gnd cell_6t
Xbit_r161_c68 bl[68] br[68] wl[161] vdd gnd cell_6t
Xbit_r162_c68 bl[68] br[68] wl[162] vdd gnd cell_6t
Xbit_r163_c68 bl[68] br[68] wl[163] vdd gnd cell_6t
Xbit_r164_c68 bl[68] br[68] wl[164] vdd gnd cell_6t
Xbit_r165_c68 bl[68] br[68] wl[165] vdd gnd cell_6t
Xbit_r166_c68 bl[68] br[68] wl[166] vdd gnd cell_6t
Xbit_r167_c68 bl[68] br[68] wl[167] vdd gnd cell_6t
Xbit_r168_c68 bl[68] br[68] wl[168] vdd gnd cell_6t
Xbit_r169_c68 bl[68] br[68] wl[169] vdd gnd cell_6t
Xbit_r170_c68 bl[68] br[68] wl[170] vdd gnd cell_6t
Xbit_r171_c68 bl[68] br[68] wl[171] vdd gnd cell_6t
Xbit_r172_c68 bl[68] br[68] wl[172] vdd gnd cell_6t
Xbit_r173_c68 bl[68] br[68] wl[173] vdd gnd cell_6t
Xbit_r174_c68 bl[68] br[68] wl[174] vdd gnd cell_6t
Xbit_r175_c68 bl[68] br[68] wl[175] vdd gnd cell_6t
Xbit_r176_c68 bl[68] br[68] wl[176] vdd gnd cell_6t
Xbit_r177_c68 bl[68] br[68] wl[177] vdd gnd cell_6t
Xbit_r178_c68 bl[68] br[68] wl[178] vdd gnd cell_6t
Xbit_r179_c68 bl[68] br[68] wl[179] vdd gnd cell_6t
Xbit_r180_c68 bl[68] br[68] wl[180] vdd gnd cell_6t
Xbit_r181_c68 bl[68] br[68] wl[181] vdd gnd cell_6t
Xbit_r182_c68 bl[68] br[68] wl[182] vdd gnd cell_6t
Xbit_r183_c68 bl[68] br[68] wl[183] vdd gnd cell_6t
Xbit_r184_c68 bl[68] br[68] wl[184] vdd gnd cell_6t
Xbit_r185_c68 bl[68] br[68] wl[185] vdd gnd cell_6t
Xbit_r186_c68 bl[68] br[68] wl[186] vdd gnd cell_6t
Xbit_r187_c68 bl[68] br[68] wl[187] vdd gnd cell_6t
Xbit_r188_c68 bl[68] br[68] wl[188] vdd gnd cell_6t
Xbit_r189_c68 bl[68] br[68] wl[189] vdd gnd cell_6t
Xbit_r190_c68 bl[68] br[68] wl[190] vdd gnd cell_6t
Xbit_r191_c68 bl[68] br[68] wl[191] vdd gnd cell_6t
Xbit_r192_c68 bl[68] br[68] wl[192] vdd gnd cell_6t
Xbit_r193_c68 bl[68] br[68] wl[193] vdd gnd cell_6t
Xbit_r194_c68 bl[68] br[68] wl[194] vdd gnd cell_6t
Xbit_r195_c68 bl[68] br[68] wl[195] vdd gnd cell_6t
Xbit_r196_c68 bl[68] br[68] wl[196] vdd gnd cell_6t
Xbit_r197_c68 bl[68] br[68] wl[197] vdd gnd cell_6t
Xbit_r198_c68 bl[68] br[68] wl[198] vdd gnd cell_6t
Xbit_r199_c68 bl[68] br[68] wl[199] vdd gnd cell_6t
Xbit_r200_c68 bl[68] br[68] wl[200] vdd gnd cell_6t
Xbit_r201_c68 bl[68] br[68] wl[201] vdd gnd cell_6t
Xbit_r202_c68 bl[68] br[68] wl[202] vdd gnd cell_6t
Xbit_r203_c68 bl[68] br[68] wl[203] vdd gnd cell_6t
Xbit_r204_c68 bl[68] br[68] wl[204] vdd gnd cell_6t
Xbit_r205_c68 bl[68] br[68] wl[205] vdd gnd cell_6t
Xbit_r206_c68 bl[68] br[68] wl[206] vdd gnd cell_6t
Xbit_r207_c68 bl[68] br[68] wl[207] vdd gnd cell_6t
Xbit_r208_c68 bl[68] br[68] wl[208] vdd gnd cell_6t
Xbit_r209_c68 bl[68] br[68] wl[209] vdd gnd cell_6t
Xbit_r210_c68 bl[68] br[68] wl[210] vdd gnd cell_6t
Xbit_r211_c68 bl[68] br[68] wl[211] vdd gnd cell_6t
Xbit_r212_c68 bl[68] br[68] wl[212] vdd gnd cell_6t
Xbit_r213_c68 bl[68] br[68] wl[213] vdd gnd cell_6t
Xbit_r214_c68 bl[68] br[68] wl[214] vdd gnd cell_6t
Xbit_r215_c68 bl[68] br[68] wl[215] vdd gnd cell_6t
Xbit_r216_c68 bl[68] br[68] wl[216] vdd gnd cell_6t
Xbit_r217_c68 bl[68] br[68] wl[217] vdd gnd cell_6t
Xbit_r218_c68 bl[68] br[68] wl[218] vdd gnd cell_6t
Xbit_r219_c68 bl[68] br[68] wl[219] vdd gnd cell_6t
Xbit_r220_c68 bl[68] br[68] wl[220] vdd gnd cell_6t
Xbit_r221_c68 bl[68] br[68] wl[221] vdd gnd cell_6t
Xbit_r222_c68 bl[68] br[68] wl[222] vdd gnd cell_6t
Xbit_r223_c68 bl[68] br[68] wl[223] vdd gnd cell_6t
Xbit_r224_c68 bl[68] br[68] wl[224] vdd gnd cell_6t
Xbit_r225_c68 bl[68] br[68] wl[225] vdd gnd cell_6t
Xbit_r226_c68 bl[68] br[68] wl[226] vdd gnd cell_6t
Xbit_r227_c68 bl[68] br[68] wl[227] vdd gnd cell_6t
Xbit_r228_c68 bl[68] br[68] wl[228] vdd gnd cell_6t
Xbit_r229_c68 bl[68] br[68] wl[229] vdd gnd cell_6t
Xbit_r230_c68 bl[68] br[68] wl[230] vdd gnd cell_6t
Xbit_r231_c68 bl[68] br[68] wl[231] vdd gnd cell_6t
Xbit_r232_c68 bl[68] br[68] wl[232] vdd gnd cell_6t
Xbit_r233_c68 bl[68] br[68] wl[233] vdd gnd cell_6t
Xbit_r234_c68 bl[68] br[68] wl[234] vdd gnd cell_6t
Xbit_r235_c68 bl[68] br[68] wl[235] vdd gnd cell_6t
Xbit_r236_c68 bl[68] br[68] wl[236] vdd gnd cell_6t
Xbit_r237_c68 bl[68] br[68] wl[237] vdd gnd cell_6t
Xbit_r238_c68 bl[68] br[68] wl[238] vdd gnd cell_6t
Xbit_r239_c68 bl[68] br[68] wl[239] vdd gnd cell_6t
Xbit_r240_c68 bl[68] br[68] wl[240] vdd gnd cell_6t
Xbit_r241_c68 bl[68] br[68] wl[241] vdd gnd cell_6t
Xbit_r242_c68 bl[68] br[68] wl[242] vdd gnd cell_6t
Xbit_r243_c68 bl[68] br[68] wl[243] vdd gnd cell_6t
Xbit_r244_c68 bl[68] br[68] wl[244] vdd gnd cell_6t
Xbit_r245_c68 bl[68] br[68] wl[245] vdd gnd cell_6t
Xbit_r246_c68 bl[68] br[68] wl[246] vdd gnd cell_6t
Xbit_r247_c68 bl[68] br[68] wl[247] vdd gnd cell_6t
Xbit_r248_c68 bl[68] br[68] wl[248] vdd gnd cell_6t
Xbit_r249_c68 bl[68] br[68] wl[249] vdd gnd cell_6t
Xbit_r250_c68 bl[68] br[68] wl[250] vdd gnd cell_6t
Xbit_r251_c68 bl[68] br[68] wl[251] vdd gnd cell_6t
Xbit_r252_c68 bl[68] br[68] wl[252] vdd gnd cell_6t
Xbit_r253_c68 bl[68] br[68] wl[253] vdd gnd cell_6t
Xbit_r254_c68 bl[68] br[68] wl[254] vdd gnd cell_6t
Xbit_r255_c68 bl[68] br[68] wl[255] vdd gnd cell_6t
Xbit_r0_c69 bl[69] br[69] wl[0] vdd gnd cell_6t
Xbit_r1_c69 bl[69] br[69] wl[1] vdd gnd cell_6t
Xbit_r2_c69 bl[69] br[69] wl[2] vdd gnd cell_6t
Xbit_r3_c69 bl[69] br[69] wl[3] vdd gnd cell_6t
Xbit_r4_c69 bl[69] br[69] wl[4] vdd gnd cell_6t
Xbit_r5_c69 bl[69] br[69] wl[5] vdd gnd cell_6t
Xbit_r6_c69 bl[69] br[69] wl[6] vdd gnd cell_6t
Xbit_r7_c69 bl[69] br[69] wl[7] vdd gnd cell_6t
Xbit_r8_c69 bl[69] br[69] wl[8] vdd gnd cell_6t
Xbit_r9_c69 bl[69] br[69] wl[9] vdd gnd cell_6t
Xbit_r10_c69 bl[69] br[69] wl[10] vdd gnd cell_6t
Xbit_r11_c69 bl[69] br[69] wl[11] vdd gnd cell_6t
Xbit_r12_c69 bl[69] br[69] wl[12] vdd gnd cell_6t
Xbit_r13_c69 bl[69] br[69] wl[13] vdd gnd cell_6t
Xbit_r14_c69 bl[69] br[69] wl[14] vdd gnd cell_6t
Xbit_r15_c69 bl[69] br[69] wl[15] vdd gnd cell_6t
Xbit_r16_c69 bl[69] br[69] wl[16] vdd gnd cell_6t
Xbit_r17_c69 bl[69] br[69] wl[17] vdd gnd cell_6t
Xbit_r18_c69 bl[69] br[69] wl[18] vdd gnd cell_6t
Xbit_r19_c69 bl[69] br[69] wl[19] vdd gnd cell_6t
Xbit_r20_c69 bl[69] br[69] wl[20] vdd gnd cell_6t
Xbit_r21_c69 bl[69] br[69] wl[21] vdd gnd cell_6t
Xbit_r22_c69 bl[69] br[69] wl[22] vdd gnd cell_6t
Xbit_r23_c69 bl[69] br[69] wl[23] vdd gnd cell_6t
Xbit_r24_c69 bl[69] br[69] wl[24] vdd gnd cell_6t
Xbit_r25_c69 bl[69] br[69] wl[25] vdd gnd cell_6t
Xbit_r26_c69 bl[69] br[69] wl[26] vdd gnd cell_6t
Xbit_r27_c69 bl[69] br[69] wl[27] vdd gnd cell_6t
Xbit_r28_c69 bl[69] br[69] wl[28] vdd gnd cell_6t
Xbit_r29_c69 bl[69] br[69] wl[29] vdd gnd cell_6t
Xbit_r30_c69 bl[69] br[69] wl[30] vdd gnd cell_6t
Xbit_r31_c69 bl[69] br[69] wl[31] vdd gnd cell_6t
Xbit_r32_c69 bl[69] br[69] wl[32] vdd gnd cell_6t
Xbit_r33_c69 bl[69] br[69] wl[33] vdd gnd cell_6t
Xbit_r34_c69 bl[69] br[69] wl[34] vdd gnd cell_6t
Xbit_r35_c69 bl[69] br[69] wl[35] vdd gnd cell_6t
Xbit_r36_c69 bl[69] br[69] wl[36] vdd gnd cell_6t
Xbit_r37_c69 bl[69] br[69] wl[37] vdd gnd cell_6t
Xbit_r38_c69 bl[69] br[69] wl[38] vdd gnd cell_6t
Xbit_r39_c69 bl[69] br[69] wl[39] vdd gnd cell_6t
Xbit_r40_c69 bl[69] br[69] wl[40] vdd gnd cell_6t
Xbit_r41_c69 bl[69] br[69] wl[41] vdd gnd cell_6t
Xbit_r42_c69 bl[69] br[69] wl[42] vdd gnd cell_6t
Xbit_r43_c69 bl[69] br[69] wl[43] vdd gnd cell_6t
Xbit_r44_c69 bl[69] br[69] wl[44] vdd gnd cell_6t
Xbit_r45_c69 bl[69] br[69] wl[45] vdd gnd cell_6t
Xbit_r46_c69 bl[69] br[69] wl[46] vdd gnd cell_6t
Xbit_r47_c69 bl[69] br[69] wl[47] vdd gnd cell_6t
Xbit_r48_c69 bl[69] br[69] wl[48] vdd gnd cell_6t
Xbit_r49_c69 bl[69] br[69] wl[49] vdd gnd cell_6t
Xbit_r50_c69 bl[69] br[69] wl[50] vdd gnd cell_6t
Xbit_r51_c69 bl[69] br[69] wl[51] vdd gnd cell_6t
Xbit_r52_c69 bl[69] br[69] wl[52] vdd gnd cell_6t
Xbit_r53_c69 bl[69] br[69] wl[53] vdd gnd cell_6t
Xbit_r54_c69 bl[69] br[69] wl[54] vdd gnd cell_6t
Xbit_r55_c69 bl[69] br[69] wl[55] vdd gnd cell_6t
Xbit_r56_c69 bl[69] br[69] wl[56] vdd gnd cell_6t
Xbit_r57_c69 bl[69] br[69] wl[57] vdd gnd cell_6t
Xbit_r58_c69 bl[69] br[69] wl[58] vdd gnd cell_6t
Xbit_r59_c69 bl[69] br[69] wl[59] vdd gnd cell_6t
Xbit_r60_c69 bl[69] br[69] wl[60] vdd gnd cell_6t
Xbit_r61_c69 bl[69] br[69] wl[61] vdd gnd cell_6t
Xbit_r62_c69 bl[69] br[69] wl[62] vdd gnd cell_6t
Xbit_r63_c69 bl[69] br[69] wl[63] vdd gnd cell_6t
Xbit_r64_c69 bl[69] br[69] wl[64] vdd gnd cell_6t
Xbit_r65_c69 bl[69] br[69] wl[65] vdd gnd cell_6t
Xbit_r66_c69 bl[69] br[69] wl[66] vdd gnd cell_6t
Xbit_r67_c69 bl[69] br[69] wl[67] vdd gnd cell_6t
Xbit_r68_c69 bl[69] br[69] wl[68] vdd gnd cell_6t
Xbit_r69_c69 bl[69] br[69] wl[69] vdd gnd cell_6t
Xbit_r70_c69 bl[69] br[69] wl[70] vdd gnd cell_6t
Xbit_r71_c69 bl[69] br[69] wl[71] vdd gnd cell_6t
Xbit_r72_c69 bl[69] br[69] wl[72] vdd gnd cell_6t
Xbit_r73_c69 bl[69] br[69] wl[73] vdd gnd cell_6t
Xbit_r74_c69 bl[69] br[69] wl[74] vdd gnd cell_6t
Xbit_r75_c69 bl[69] br[69] wl[75] vdd gnd cell_6t
Xbit_r76_c69 bl[69] br[69] wl[76] vdd gnd cell_6t
Xbit_r77_c69 bl[69] br[69] wl[77] vdd gnd cell_6t
Xbit_r78_c69 bl[69] br[69] wl[78] vdd gnd cell_6t
Xbit_r79_c69 bl[69] br[69] wl[79] vdd gnd cell_6t
Xbit_r80_c69 bl[69] br[69] wl[80] vdd gnd cell_6t
Xbit_r81_c69 bl[69] br[69] wl[81] vdd gnd cell_6t
Xbit_r82_c69 bl[69] br[69] wl[82] vdd gnd cell_6t
Xbit_r83_c69 bl[69] br[69] wl[83] vdd gnd cell_6t
Xbit_r84_c69 bl[69] br[69] wl[84] vdd gnd cell_6t
Xbit_r85_c69 bl[69] br[69] wl[85] vdd gnd cell_6t
Xbit_r86_c69 bl[69] br[69] wl[86] vdd gnd cell_6t
Xbit_r87_c69 bl[69] br[69] wl[87] vdd gnd cell_6t
Xbit_r88_c69 bl[69] br[69] wl[88] vdd gnd cell_6t
Xbit_r89_c69 bl[69] br[69] wl[89] vdd gnd cell_6t
Xbit_r90_c69 bl[69] br[69] wl[90] vdd gnd cell_6t
Xbit_r91_c69 bl[69] br[69] wl[91] vdd gnd cell_6t
Xbit_r92_c69 bl[69] br[69] wl[92] vdd gnd cell_6t
Xbit_r93_c69 bl[69] br[69] wl[93] vdd gnd cell_6t
Xbit_r94_c69 bl[69] br[69] wl[94] vdd gnd cell_6t
Xbit_r95_c69 bl[69] br[69] wl[95] vdd gnd cell_6t
Xbit_r96_c69 bl[69] br[69] wl[96] vdd gnd cell_6t
Xbit_r97_c69 bl[69] br[69] wl[97] vdd gnd cell_6t
Xbit_r98_c69 bl[69] br[69] wl[98] vdd gnd cell_6t
Xbit_r99_c69 bl[69] br[69] wl[99] vdd gnd cell_6t
Xbit_r100_c69 bl[69] br[69] wl[100] vdd gnd cell_6t
Xbit_r101_c69 bl[69] br[69] wl[101] vdd gnd cell_6t
Xbit_r102_c69 bl[69] br[69] wl[102] vdd gnd cell_6t
Xbit_r103_c69 bl[69] br[69] wl[103] vdd gnd cell_6t
Xbit_r104_c69 bl[69] br[69] wl[104] vdd gnd cell_6t
Xbit_r105_c69 bl[69] br[69] wl[105] vdd gnd cell_6t
Xbit_r106_c69 bl[69] br[69] wl[106] vdd gnd cell_6t
Xbit_r107_c69 bl[69] br[69] wl[107] vdd gnd cell_6t
Xbit_r108_c69 bl[69] br[69] wl[108] vdd gnd cell_6t
Xbit_r109_c69 bl[69] br[69] wl[109] vdd gnd cell_6t
Xbit_r110_c69 bl[69] br[69] wl[110] vdd gnd cell_6t
Xbit_r111_c69 bl[69] br[69] wl[111] vdd gnd cell_6t
Xbit_r112_c69 bl[69] br[69] wl[112] vdd gnd cell_6t
Xbit_r113_c69 bl[69] br[69] wl[113] vdd gnd cell_6t
Xbit_r114_c69 bl[69] br[69] wl[114] vdd gnd cell_6t
Xbit_r115_c69 bl[69] br[69] wl[115] vdd gnd cell_6t
Xbit_r116_c69 bl[69] br[69] wl[116] vdd gnd cell_6t
Xbit_r117_c69 bl[69] br[69] wl[117] vdd gnd cell_6t
Xbit_r118_c69 bl[69] br[69] wl[118] vdd gnd cell_6t
Xbit_r119_c69 bl[69] br[69] wl[119] vdd gnd cell_6t
Xbit_r120_c69 bl[69] br[69] wl[120] vdd gnd cell_6t
Xbit_r121_c69 bl[69] br[69] wl[121] vdd gnd cell_6t
Xbit_r122_c69 bl[69] br[69] wl[122] vdd gnd cell_6t
Xbit_r123_c69 bl[69] br[69] wl[123] vdd gnd cell_6t
Xbit_r124_c69 bl[69] br[69] wl[124] vdd gnd cell_6t
Xbit_r125_c69 bl[69] br[69] wl[125] vdd gnd cell_6t
Xbit_r126_c69 bl[69] br[69] wl[126] vdd gnd cell_6t
Xbit_r127_c69 bl[69] br[69] wl[127] vdd gnd cell_6t
Xbit_r128_c69 bl[69] br[69] wl[128] vdd gnd cell_6t
Xbit_r129_c69 bl[69] br[69] wl[129] vdd gnd cell_6t
Xbit_r130_c69 bl[69] br[69] wl[130] vdd gnd cell_6t
Xbit_r131_c69 bl[69] br[69] wl[131] vdd gnd cell_6t
Xbit_r132_c69 bl[69] br[69] wl[132] vdd gnd cell_6t
Xbit_r133_c69 bl[69] br[69] wl[133] vdd gnd cell_6t
Xbit_r134_c69 bl[69] br[69] wl[134] vdd gnd cell_6t
Xbit_r135_c69 bl[69] br[69] wl[135] vdd gnd cell_6t
Xbit_r136_c69 bl[69] br[69] wl[136] vdd gnd cell_6t
Xbit_r137_c69 bl[69] br[69] wl[137] vdd gnd cell_6t
Xbit_r138_c69 bl[69] br[69] wl[138] vdd gnd cell_6t
Xbit_r139_c69 bl[69] br[69] wl[139] vdd gnd cell_6t
Xbit_r140_c69 bl[69] br[69] wl[140] vdd gnd cell_6t
Xbit_r141_c69 bl[69] br[69] wl[141] vdd gnd cell_6t
Xbit_r142_c69 bl[69] br[69] wl[142] vdd gnd cell_6t
Xbit_r143_c69 bl[69] br[69] wl[143] vdd gnd cell_6t
Xbit_r144_c69 bl[69] br[69] wl[144] vdd gnd cell_6t
Xbit_r145_c69 bl[69] br[69] wl[145] vdd gnd cell_6t
Xbit_r146_c69 bl[69] br[69] wl[146] vdd gnd cell_6t
Xbit_r147_c69 bl[69] br[69] wl[147] vdd gnd cell_6t
Xbit_r148_c69 bl[69] br[69] wl[148] vdd gnd cell_6t
Xbit_r149_c69 bl[69] br[69] wl[149] vdd gnd cell_6t
Xbit_r150_c69 bl[69] br[69] wl[150] vdd gnd cell_6t
Xbit_r151_c69 bl[69] br[69] wl[151] vdd gnd cell_6t
Xbit_r152_c69 bl[69] br[69] wl[152] vdd gnd cell_6t
Xbit_r153_c69 bl[69] br[69] wl[153] vdd gnd cell_6t
Xbit_r154_c69 bl[69] br[69] wl[154] vdd gnd cell_6t
Xbit_r155_c69 bl[69] br[69] wl[155] vdd gnd cell_6t
Xbit_r156_c69 bl[69] br[69] wl[156] vdd gnd cell_6t
Xbit_r157_c69 bl[69] br[69] wl[157] vdd gnd cell_6t
Xbit_r158_c69 bl[69] br[69] wl[158] vdd gnd cell_6t
Xbit_r159_c69 bl[69] br[69] wl[159] vdd gnd cell_6t
Xbit_r160_c69 bl[69] br[69] wl[160] vdd gnd cell_6t
Xbit_r161_c69 bl[69] br[69] wl[161] vdd gnd cell_6t
Xbit_r162_c69 bl[69] br[69] wl[162] vdd gnd cell_6t
Xbit_r163_c69 bl[69] br[69] wl[163] vdd gnd cell_6t
Xbit_r164_c69 bl[69] br[69] wl[164] vdd gnd cell_6t
Xbit_r165_c69 bl[69] br[69] wl[165] vdd gnd cell_6t
Xbit_r166_c69 bl[69] br[69] wl[166] vdd gnd cell_6t
Xbit_r167_c69 bl[69] br[69] wl[167] vdd gnd cell_6t
Xbit_r168_c69 bl[69] br[69] wl[168] vdd gnd cell_6t
Xbit_r169_c69 bl[69] br[69] wl[169] vdd gnd cell_6t
Xbit_r170_c69 bl[69] br[69] wl[170] vdd gnd cell_6t
Xbit_r171_c69 bl[69] br[69] wl[171] vdd gnd cell_6t
Xbit_r172_c69 bl[69] br[69] wl[172] vdd gnd cell_6t
Xbit_r173_c69 bl[69] br[69] wl[173] vdd gnd cell_6t
Xbit_r174_c69 bl[69] br[69] wl[174] vdd gnd cell_6t
Xbit_r175_c69 bl[69] br[69] wl[175] vdd gnd cell_6t
Xbit_r176_c69 bl[69] br[69] wl[176] vdd gnd cell_6t
Xbit_r177_c69 bl[69] br[69] wl[177] vdd gnd cell_6t
Xbit_r178_c69 bl[69] br[69] wl[178] vdd gnd cell_6t
Xbit_r179_c69 bl[69] br[69] wl[179] vdd gnd cell_6t
Xbit_r180_c69 bl[69] br[69] wl[180] vdd gnd cell_6t
Xbit_r181_c69 bl[69] br[69] wl[181] vdd gnd cell_6t
Xbit_r182_c69 bl[69] br[69] wl[182] vdd gnd cell_6t
Xbit_r183_c69 bl[69] br[69] wl[183] vdd gnd cell_6t
Xbit_r184_c69 bl[69] br[69] wl[184] vdd gnd cell_6t
Xbit_r185_c69 bl[69] br[69] wl[185] vdd gnd cell_6t
Xbit_r186_c69 bl[69] br[69] wl[186] vdd gnd cell_6t
Xbit_r187_c69 bl[69] br[69] wl[187] vdd gnd cell_6t
Xbit_r188_c69 bl[69] br[69] wl[188] vdd gnd cell_6t
Xbit_r189_c69 bl[69] br[69] wl[189] vdd gnd cell_6t
Xbit_r190_c69 bl[69] br[69] wl[190] vdd gnd cell_6t
Xbit_r191_c69 bl[69] br[69] wl[191] vdd gnd cell_6t
Xbit_r192_c69 bl[69] br[69] wl[192] vdd gnd cell_6t
Xbit_r193_c69 bl[69] br[69] wl[193] vdd gnd cell_6t
Xbit_r194_c69 bl[69] br[69] wl[194] vdd gnd cell_6t
Xbit_r195_c69 bl[69] br[69] wl[195] vdd gnd cell_6t
Xbit_r196_c69 bl[69] br[69] wl[196] vdd gnd cell_6t
Xbit_r197_c69 bl[69] br[69] wl[197] vdd gnd cell_6t
Xbit_r198_c69 bl[69] br[69] wl[198] vdd gnd cell_6t
Xbit_r199_c69 bl[69] br[69] wl[199] vdd gnd cell_6t
Xbit_r200_c69 bl[69] br[69] wl[200] vdd gnd cell_6t
Xbit_r201_c69 bl[69] br[69] wl[201] vdd gnd cell_6t
Xbit_r202_c69 bl[69] br[69] wl[202] vdd gnd cell_6t
Xbit_r203_c69 bl[69] br[69] wl[203] vdd gnd cell_6t
Xbit_r204_c69 bl[69] br[69] wl[204] vdd gnd cell_6t
Xbit_r205_c69 bl[69] br[69] wl[205] vdd gnd cell_6t
Xbit_r206_c69 bl[69] br[69] wl[206] vdd gnd cell_6t
Xbit_r207_c69 bl[69] br[69] wl[207] vdd gnd cell_6t
Xbit_r208_c69 bl[69] br[69] wl[208] vdd gnd cell_6t
Xbit_r209_c69 bl[69] br[69] wl[209] vdd gnd cell_6t
Xbit_r210_c69 bl[69] br[69] wl[210] vdd gnd cell_6t
Xbit_r211_c69 bl[69] br[69] wl[211] vdd gnd cell_6t
Xbit_r212_c69 bl[69] br[69] wl[212] vdd gnd cell_6t
Xbit_r213_c69 bl[69] br[69] wl[213] vdd gnd cell_6t
Xbit_r214_c69 bl[69] br[69] wl[214] vdd gnd cell_6t
Xbit_r215_c69 bl[69] br[69] wl[215] vdd gnd cell_6t
Xbit_r216_c69 bl[69] br[69] wl[216] vdd gnd cell_6t
Xbit_r217_c69 bl[69] br[69] wl[217] vdd gnd cell_6t
Xbit_r218_c69 bl[69] br[69] wl[218] vdd gnd cell_6t
Xbit_r219_c69 bl[69] br[69] wl[219] vdd gnd cell_6t
Xbit_r220_c69 bl[69] br[69] wl[220] vdd gnd cell_6t
Xbit_r221_c69 bl[69] br[69] wl[221] vdd gnd cell_6t
Xbit_r222_c69 bl[69] br[69] wl[222] vdd gnd cell_6t
Xbit_r223_c69 bl[69] br[69] wl[223] vdd gnd cell_6t
Xbit_r224_c69 bl[69] br[69] wl[224] vdd gnd cell_6t
Xbit_r225_c69 bl[69] br[69] wl[225] vdd gnd cell_6t
Xbit_r226_c69 bl[69] br[69] wl[226] vdd gnd cell_6t
Xbit_r227_c69 bl[69] br[69] wl[227] vdd gnd cell_6t
Xbit_r228_c69 bl[69] br[69] wl[228] vdd gnd cell_6t
Xbit_r229_c69 bl[69] br[69] wl[229] vdd gnd cell_6t
Xbit_r230_c69 bl[69] br[69] wl[230] vdd gnd cell_6t
Xbit_r231_c69 bl[69] br[69] wl[231] vdd gnd cell_6t
Xbit_r232_c69 bl[69] br[69] wl[232] vdd gnd cell_6t
Xbit_r233_c69 bl[69] br[69] wl[233] vdd gnd cell_6t
Xbit_r234_c69 bl[69] br[69] wl[234] vdd gnd cell_6t
Xbit_r235_c69 bl[69] br[69] wl[235] vdd gnd cell_6t
Xbit_r236_c69 bl[69] br[69] wl[236] vdd gnd cell_6t
Xbit_r237_c69 bl[69] br[69] wl[237] vdd gnd cell_6t
Xbit_r238_c69 bl[69] br[69] wl[238] vdd gnd cell_6t
Xbit_r239_c69 bl[69] br[69] wl[239] vdd gnd cell_6t
Xbit_r240_c69 bl[69] br[69] wl[240] vdd gnd cell_6t
Xbit_r241_c69 bl[69] br[69] wl[241] vdd gnd cell_6t
Xbit_r242_c69 bl[69] br[69] wl[242] vdd gnd cell_6t
Xbit_r243_c69 bl[69] br[69] wl[243] vdd gnd cell_6t
Xbit_r244_c69 bl[69] br[69] wl[244] vdd gnd cell_6t
Xbit_r245_c69 bl[69] br[69] wl[245] vdd gnd cell_6t
Xbit_r246_c69 bl[69] br[69] wl[246] vdd gnd cell_6t
Xbit_r247_c69 bl[69] br[69] wl[247] vdd gnd cell_6t
Xbit_r248_c69 bl[69] br[69] wl[248] vdd gnd cell_6t
Xbit_r249_c69 bl[69] br[69] wl[249] vdd gnd cell_6t
Xbit_r250_c69 bl[69] br[69] wl[250] vdd gnd cell_6t
Xbit_r251_c69 bl[69] br[69] wl[251] vdd gnd cell_6t
Xbit_r252_c69 bl[69] br[69] wl[252] vdd gnd cell_6t
Xbit_r253_c69 bl[69] br[69] wl[253] vdd gnd cell_6t
Xbit_r254_c69 bl[69] br[69] wl[254] vdd gnd cell_6t
Xbit_r255_c69 bl[69] br[69] wl[255] vdd gnd cell_6t
Xbit_r0_c70 bl[70] br[70] wl[0] vdd gnd cell_6t
Xbit_r1_c70 bl[70] br[70] wl[1] vdd gnd cell_6t
Xbit_r2_c70 bl[70] br[70] wl[2] vdd gnd cell_6t
Xbit_r3_c70 bl[70] br[70] wl[3] vdd gnd cell_6t
Xbit_r4_c70 bl[70] br[70] wl[4] vdd gnd cell_6t
Xbit_r5_c70 bl[70] br[70] wl[5] vdd gnd cell_6t
Xbit_r6_c70 bl[70] br[70] wl[6] vdd gnd cell_6t
Xbit_r7_c70 bl[70] br[70] wl[7] vdd gnd cell_6t
Xbit_r8_c70 bl[70] br[70] wl[8] vdd gnd cell_6t
Xbit_r9_c70 bl[70] br[70] wl[9] vdd gnd cell_6t
Xbit_r10_c70 bl[70] br[70] wl[10] vdd gnd cell_6t
Xbit_r11_c70 bl[70] br[70] wl[11] vdd gnd cell_6t
Xbit_r12_c70 bl[70] br[70] wl[12] vdd gnd cell_6t
Xbit_r13_c70 bl[70] br[70] wl[13] vdd gnd cell_6t
Xbit_r14_c70 bl[70] br[70] wl[14] vdd gnd cell_6t
Xbit_r15_c70 bl[70] br[70] wl[15] vdd gnd cell_6t
Xbit_r16_c70 bl[70] br[70] wl[16] vdd gnd cell_6t
Xbit_r17_c70 bl[70] br[70] wl[17] vdd gnd cell_6t
Xbit_r18_c70 bl[70] br[70] wl[18] vdd gnd cell_6t
Xbit_r19_c70 bl[70] br[70] wl[19] vdd gnd cell_6t
Xbit_r20_c70 bl[70] br[70] wl[20] vdd gnd cell_6t
Xbit_r21_c70 bl[70] br[70] wl[21] vdd gnd cell_6t
Xbit_r22_c70 bl[70] br[70] wl[22] vdd gnd cell_6t
Xbit_r23_c70 bl[70] br[70] wl[23] vdd gnd cell_6t
Xbit_r24_c70 bl[70] br[70] wl[24] vdd gnd cell_6t
Xbit_r25_c70 bl[70] br[70] wl[25] vdd gnd cell_6t
Xbit_r26_c70 bl[70] br[70] wl[26] vdd gnd cell_6t
Xbit_r27_c70 bl[70] br[70] wl[27] vdd gnd cell_6t
Xbit_r28_c70 bl[70] br[70] wl[28] vdd gnd cell_6t
Xbit_r29_c70 bl[70] br[70] wl[29] vdd gnd cell_6t
Xbit_r30_c70 bl[70] br[70] wl[30] vdd gnd cell_6t
Xbit_r31_c70 bl[70] br[70] wl[31] vdd gnd cell_6t
Xbit_r32_c70 bl[70] br[70] wl[32] vdd gnd cell_6t
Xbit_r33_c70 bl[70] br[70] wl[33] vdd gnd cell_6t
Xbit_r34_c70 bl[70] br[70] wl[34] vdd gnd cell_6t
Xbit_r35_c70 bl[70] br[70] wl[35] vdd gnd cell_6t
Xbit_r36_c70 bl[70] br[70] wl[36] vdd gnd cell_6t
Xbit_r37_c70 bl[70] br[70] wl[37] vdd gnd cell_6t
Xbit_r38_c70 bl[70] br[70] wl[38] vdd gnd cell_6t
Xbit_r39_c70 bl[70] br[70] wl[39] vdd gnd cell_6t
Xbit_r40_c70 bl[70] br[70] wl[40] vdd gnd cell_6t
Xbit_r41_c70 bl[70] br[70] wl[41] vdd gnd cell_6t
Xbit_r42_c70 bl[70] br[70] wl[42] vdd gnd cell_6t
Xbit_r43_c70 bl[70] br[70] wl[43] vdd gnd cell_6t
Xbit_r44_c70 bl[70] br[70] wl[44] vdd gnd cell_6t
Xbit_r45_c70 bl[70] br[70] wl[45] vdd gnd cell_6t
Xbit_r46_c70 bl[70] br[70] wl[46] vdd gnd cell_6t
Xbit_r47_c70 bl[70] br[70] wl[47] vdd gnd cell_6t
Xbit_r48_c70 bl[70] br[70] wl[48] vdd gnd cell_6t
Xbit_r49_c70 bl[70] br[70] wl[49] vdd gnd cell_6t
Xbit_r50_c70 bl[70] br[70] wl[50] vdd gnd cell_6t
Xbit_r51_c70 bl[70] br[70] wl[51] vdd gnd cell_6t
Xbit_r52_c70 bl[70] br[70] wl[52] vdd gnd cell_6t
Xbit_r53_c70 bl[70] br[70] wl[53] vdd gnd cell_6t
Xbit_r54_c70 bl[70] br[70] wl[54] vdd gnd cell_6t
Xbit_r55_c70 bl[70] br[70] wl[55] vdd gnd cell_6t
Xbit_r56_c70 bl[70] br[70] wl[56] vdd gnd cell_6t
Xbit_r57_c70 bl[70] br[70] wl[57] vdd gnd cell_6t
Xbit_r58_c70 bl[70] br[70] wl[58] vdd gnd cell_6t
Xbit_r59_c70 bl[70] br[70] wl[59] vdd gnd cell_6t
Xbit_r60_c70 bl[70] br[70] wl[60] vdd gnd cell_6t
Xbit_r61_c70 bl[70] br[70] wl[61] vdd gnd cell_6t
Xbit_r62_c70 bl[70] br[70] wl[62] vdd gnd cell_6t
Xbit_r63_c70 bl[70] br[70] wl[63] vdd gnd cell_6t
Xbit_r64_c70 bl[70] br[70] wl[64] vdd gnd cell_6t
Xbit_r65_c70 bl[70] br[70] wl[65] vdd gnd cell_6t
Xbit_r66_c70 bl[70] br[70] wl[66] vdd gnd cell_6t
Xbit_r67_c70 bl[70] br[70] wl[67] vdd gnd cell_6t
Xbit_r68_c70 bl[70] br[70] wl[68] vdd gnd cell_6t
Xbit_r69_c70 bl[70] br[70] wl[69] vdd gnd cell_6t
Xbit_r70_c70 bl[70] br[70] wl[70] vdd gnd cell_6t
Xbit_r71_c70 bl[70] br[70] wl[71] vdd gnd cell_6t
Xbit_r72_c70 bl[70] br[70] wl[72] vdd gnd cell_6t
Xbit_r73_c70 bl[70] br[70] wl[73] vdd gnd cell_6t
Xbit_r74_c70 bl[70] br[70] wl[74] vdd gnd cell_6t
Xbit_r75_c70 bl[70] br[70] wl[75] vdd gnd cell_6t
Xbit_r76_c70 bl[70] br[70] wl[76] vdd gnd cell_6t
Xbit_r77_c70 bl[70] br[70] wl[77] vdd gnd cell_6t
Xbit_r78_c70 bl[70] br[70] wl[78] vdd gnd cell_6t
Xbit_r79_c70 bl[70] br[70] wl[79] vdd gnd cell_6t
Xbit_r80_c70 bl[70] br[70] wl[80] vdd gnd cell_6t
Xbit_r81_c70 bl[70] br[70] wl[81] vdd gnd cell_6t
Xbit_r82_c70 bl[70] br[70] wl[82] vdd gnd cell_6t
Xbit_r83_c70 bl[70] br[70] wl[83] vdd gnd cell_6t
Xbit_r84_c70 bl[70] br[70] wl[84] vdd gnd cell_6t
Xbit_r85_c70 bl[70] br[70] wl[85] vdd gnd cell_6t
Xbit_r86_c70 bl[70] br[70] wl[86] vdd gnd cell_6t
Xbit_r87_c70 bl[70] br[70] wl[87] vdd gnd cell_6t
Xbit_r88_c70 bl[70] br[70] wl[88] vdd gnd cell_6t
Xbit_r89_c70 bl[70] br[70] wl[89] vdd gnd cell_6t
Xbit_r90_c70 bl[70] br[70] wl[90] vdd gnd cell_6t
Xbit_r91_c70 bl[70] br[70] wl[91] vdd gnd cell_6t
Xbit_r92_c70 bl[70] br[70] wl[92] vdd gnd cell_6t
Xbit_r93_c70 bl[70] br[70] wl[93] vdd gnd cell_6t
Xbit_r94_c70 bl[70] br[70] wl[94] vdd gnd cell_6t
Xbit_r95_c70 bl[70] br[70] wl[95] vdd gnd cell_6t
Xbit_r96_c70 bl[70] br[70] wl[96] vdd gnd cell_6t
Xbit_r97_c70 bl[70] br[70] wl[97] vdd gnd cell_6t
Xbit_r98_c70 bl[70] br[70] wl[98] vdd gnd cell_6t
Xbit_r99_c70 bl[70] br[70] wl[99] vdd gnd cell_6t
Xbit_r100_c70 bl[70] br[70] wl[100] vdd gnd cell_6t
Xbit_r101_c70 bl[70] br[70] wl[101] vdd gnd cell_6t
Xbit_r102_c70 bl[70] br[70] wl[102] vdd gnd cell_6t
Xbit_r103_c70 bl[70] br[70] wl[103] vdd gnd cell_6t
Xbit_r104_c70 bl[70] br[70] wl[104] vdd gnd cell_6t
Xbit_r105_c70 bl[70] br[70] wl[105] vdd gnd cell_6t
Xbit_r106_c70 bl[70] br[70] wl[106] vdd gnd cell_6t
Xbit_r107_c70 bl[70] br[70] wl[107] vdd gnd cell_6t
Xbit_r108_c70 bl[70] br[70] wl[108] vdd gnd cell_6t
Xbit_r109_c70 bl[70] br[70] wl[109] vdd gnd cell_6t
Xbit_r110_c70 bl[70] br[70] wl[110] vdd gnd cell_6t
Xbit_r111_c70 bl[70] br[70] wl[111] vdd gnd cell_6t
Xbit_r112_c70 bl[70] br[70] wl[112] vdd gnd cell_6t
Xbit_r113_c70 bl[70] br[70] wl[113] vdd gnd cell_6t
Xbit_r114_c70 bl[70] br[70] wl[114] vdd gnd cell_6t
Xbit_r115_c70 bl[70] br[70] wl[115] vdd gnd cell_6t
Xbit_r116_c70 bl[70] br[70] wl[116] vdd gnd cell_6t
Xbit_r117_c70 bl[70] br[70] wl[117] vdd gnd cell_6t
Xbit_r118_c70 bl[70] br[70] wl[118] vdd gnd cell_6t
Xbit_r119_c70 bl[70] br[70] wl[119] vdd gnd cell_6t
Xbit_r120_c70 bl[70] br[70] wl[120] vdd gnd cell_6t
Xbit_r121_c70 bl[70] br[70] wl[121] vdd gnd cell_6t
Xbit_r122_c70 bl[70] br[70] wl[122] vdd gnd cell_6t
Xbit_r123_c70 bl[70] br[70] wl[123] vdd gnd cell_6t
Xbit_r124_c70 bl[70] br[70] wl[124] vdd gnd cell_6t
Xbit_r125_c70 bl[70] br[70] wl[125] vdd gnd cell_6t
Xbit_r126_c70 bl[70] br[70] wl[126] vdd gnd cell_6t
Xbit_r127_c70 bl[70] br[70] wl[127] vdd gnd cell_6t
Xbit_r128_c70 bl[70] br[70] wl[128] vdd gnd cell_6t
Xbit_r129_c70 bl[70] br[70] wl[129] vdd gnd cell_6t
Xbit_r130_c70 bl[70] br[70] wl[130] vdd gnd cell_6t
Xbit_r131_c70 bl[70] br[70] wl[131] vdd gnd cell_6t
Xbit_r132_c70 bl[70] br[70] wl[132] vdd gnd cell_6t
Xbit_r133_c70 bl[70] br[70] wl[133] vdd gnd cell_6t
Xbit_r134_c70 bl[70] br[70] wl[134] vdd gnd cell_6t
Xbit_r135_c70 bl[70] br[70] wl[135] vdd gnd cell_6t
Xbit_r136_c70 bl[70] br[70] wl[136] vdd gnd cell_6t
Xbit_r137_c70 bl[70] br[70] wl[137] vdd gnd cell_6t
Xbit_r138_c70 bl[70] br[70] wl[138] vdd gnd cell_6t
Xbit_r139_c70 bl[70] br[70] wl[139] vdd gnd cell_6t
Xbit_r140_c70 bl[70] br[70] wl[140] vdd gnd cell_6t
Xbit_r141_c70 bl[70] br[70] wl[141] vdd gnd cell_6t
Xbit_r142_c70 bl[70] br[70] wl[142] vdd gnd cell_6t
Xbit_r143_c70 bl[70] br[70] wl[143] vdd gnd cell_6t
Xbit_r144_c70 bl[70] br[70] wl[144] vdd gnd cell_6t
Xbit_r145_c70 bl[70] br[70] wl[145] vdd gnd cell_6t
Xbit_r146_c70 bl[70] br[70] wl[146] vdd gnd cell_6t
Xbit_r147_c70 bl[70] br[70] wl[147] vdd gnd cell_6t
Xbit_r148_c70 bl[70] br[70] wl[148] vdd gnd cell_6t
Xbit_r149_c70 bl[70] br[70] wl[149] vdd gnd cell_6t
Xbit_r150_c70 bl[70] br[70] wl[150] vdd gnd cell_6t
Xbit_r151_c70 bl[70] br[70] wl[151] vdd gnd cell_6t
Xbit_r152_c70 bl[70] br[70] wl[152] vdd gnd cell_6t
Xbit_r153_c70 bl[70] br[70] wl[153] vdd gnd cell_6t
Xbit_r154_c70 bl[70] br[70] wl[154] vdd gnd cell_6t
Xbit_r155_c70 bl[70] br[70] wl[155] vdd gnd cell_6t
Xbit_r156_c70 bl[70] br[70] wl[156] vdd gnd cell_6t
Xbit_r157_c70 bl[70] br[70] wl[157] vdd gnd cell_6t
Xbit_r158_c70 bl[70] br[70] wl[158] vdd gnd cell_6t
Xbit_r159_c70 bl[70] br[70] wl[159] vdd gnd cell_6t
Xbit_r160_c70 bl[70] br[70] wl[160] vdd gnd cell_6t
Xbit_r161_c70 bl[70] br[70] wl[161] vdd gnd cell_6t
Xbit_r162_c70 bl[70] br[70] wl[162] vdd gnd cell_6t
Xbit_r163_c70 bl[70] br[70] wl[163] vdd gnd cell_6t
Xbit_r164_c70 bl[70] br[70] wl[164] vdd gnd cell_6t
Xbit_r165_c70 bl[70] br[70] wl[165] vdd gnd cell_6t
Xbit_r166_c70 bl[70] br[70] wl[166] vdd gnd cell_6t
Xbit_r167_c70 bl[70] br[70] wl[167] vdd gnd cell_6t
Xbit_r168_c70 bl[70] br[70] wl[168] vdd gnd cell_6t
Xbit_r169_c70 bl[70] br[70] wl[169] vdd gnd cell_6t
Xbit_r170_c70 bl[70] br[70] wl[170] vdd gnd cell_6t
Xbit_r171_c70 bl[70] br[70] wl[171] vdd gnd cell_6t
Xbit_r172_c70 bl[70] br[70] wl[172] vdd gnd cell_6t
Xbit_r173_c70 bl[70] br[70] wl[173] vdd gnd cell_6t
Xbit_r174_c70 bl[70] br[70] wl[174] vdd gnd cell_6t
Xbit_r175_c70 bl[70] br[70] wl[175] vdd gnd cell_6t
Xbit_r176_c70 bl[70] br[70] wl[176] vdd gnd cell_6t
Xbit_r177_c70 bl[70] br[70] wl[177] vdd gnd cell_6t
Xbit_r178_c70 bl[70] br[70] wl[178] vdd gnd cell_6t
Xbit_r179_c70 bl[70] br[70] wl[179] vdd gnd cell_6t
Xbit_r180_c70 bl[70] br[70] wl[180] vdd gnd cell_6t
Xbit_r181_c70 bl[70] br[70] wl[181] vdd gnd cell_6t
Xbit_r182_c70 bl[70] br[70] wl[182] vdd gnd cell_6t
Xbit_r183_c70 bl[70] br[70] wl[183] vdd gnd cell_6t
Xbit_r184_c70 bl[70] br[70] wl[184] vdd gnd cell_6t
Xbit_r185_c70 bl[70] br[70] wl[185] vdd gnd cell_6t
Xbit_r186_c70 bl[70] br[70] wl[186] vdd gnd cell_6t
Xbit_r187_c70 bl[70] br[70] wl[187] vdd gnd cell_6t
Xbit_r188_c70 bl[70] br[70] wl[188] vdd gnd cell_6t
Xbit_r189_c70 bl[70] br[70] wl[189] vdd gnd cell_6t
Xbit_r190_c70 bl[70] br[70] wl[190] vdd gnd cell_6t
Xbit_r191_c70 bl[70] br[70] wl[191] vdd gnd cell_6t
Xbit_r192_c70 bl[70] br[70] wl[192] vdd gnd cell_6t
Xbit_r193_c70 bl[70] br[70] wl[193] vdd gnd cell_6t
Xbit_r194_c70 bl[70] br[70] wl[194] vdd gnd cell_6t
Xbit_r195_c70 bl[70] br[70] wl[195] vdd gnd cell_6t
Xbit_r196_c70 bl[70] br[70] wl[196] vdd gnd cell_6t
Xbit_r197_c70 bl[70] br[70] wl[197] vdd gnd cell_6t
Xbit_r198_c70 bl[70] br[70] wl[198] vdd gnd cell_6t
Xbit_r199_c70 bl[70] br[70] wl[199] vdd gnd cell_6t
Xbit_r200_c70 bl[70] br[70] wl[200] vdd gnd cell_6t
Xbit_r201_c70 bl[70] br[70] wl[201] vdd gnd cell_6t
Xbit_r202_c70 bl[70] br[70] wl[202] vdd gnd cell_6t
Xbit_r203_c70 bl[70] br[70] wl[203] vdd gnd cell_6t
Xbit_r204_c70 bl[70] br[70] wl[204] vdd gnd cell_6t
Xbit_r205_c70 bl[70] br[70] wl[205] vdd gnd cell_6t
Xbit_r206_c70 bl[70] br[70] wl[206] vdd gnd cell_6t
Xbit_r207_c70 bl[70] br[70] wl[207] vdd gnd cell_6t
Xbit_r208_c70 bl[70] br[70] wl[208] vdd gnd cell_6t
Xbit_r209_c70 bl[70] br[70] wl[209] vdd gnd cell_6t
Xbit_r210_c70 bl[70] br[70] wl[210] vdd gnd cell_6t
Xbit_r211_c70 bl[70] br[70] wl[211] vdd gnd cell_6t
Xbit_r212_c70 bl[70] br[70] wl[212] vdd gnd cell_6t
Xbit_r213_c70 bl[70] br[70] wl[213] vdd gnd cell_6t
Xbit_r214_c70 bl[70] br[70] wl[214] vdd gnd cell_6t
Xbit_r215_c70 bl[70] br[70] wl[215] vdd gnd cell_6t
Xbit_r216_c70 bl[70] br[70] wl[216] vdd gnd cell_6t
Xbit_r217_c70 bl[70] br[70] wl[217] vdd gnd cell_6t
Xbit_r218_c70 bl[70] br[70] wl[218] vdd gnd cell_6t
Xbit_r219_c70 bl[70] br[70] wl[219] vdd gnd cell_6t
Xbit_r220_c70 bl[70] br[70] wl[220] vdd gnd cell_6t
Xbit_r221_c70 bl[70] br[70] wl[221] vdd gnd cell_6t
Xbit_r222_c70 bl[70] br[70] wl[222] vdd gnd cell_6t
Xbit_r223_c70 bl[70] br[70] wl[223] vdd gnd cell_6t
Xbit_r224_c70 bl[70] br[70] wl[224] vdd gnd cell_6t
Xbit_r225_c70 bl[70] br[70] wl[225] vdd gnd cell_6t
Xbit_r226_c70 bl[70] br[70] wl[226] vdd gnd cell_6t
Xbit_r227_c70 bl[70] br[70] wl[227] vdd gnd cell_6t
Xbit_r228_c70 bl[70] br[70] wl[228] vdd gnd cell_6t
Xbit_r229_c70 bl[70] br[70] wl[229] vdd gnd cell_6t
Xbit_r230_c70 bl[70] br[70] wl[230] vdd gnd cell_6t
Xbit_r231_c70 bl[70] br[70] wl[231] vdd gnd cell_6t
Xbit_r232_c70 bl[70] br[70] wl[232] vdd gnd cell_6t
Xbit_r233_c70 bl[70] br[70] wl[233] vdd gnd cell_6t
Xbit_r234_c70 bl[70] br[70] wl[234] vdd gnd cell_6t
Xbit_r235_c70 bl[70] br[70] wl[235] vdd gnd cell_6t
Xbit_r236_c70 bl[70] br[70] wl[236] vdd gnd cell_6t
Xbit_r237_c70 bl[70] br[70] wl[237] vdd gnd cell_6t
Xbit_r238_c70 bl[70] br[70] wl[238] vdd gnd cell_6t
Xbit_r239_c70 bl[70] br[70] wl[239] vdd gnd cell_6t
Xbit_r240_c70 bl[70] br[70] wl[240] vdd gnd cell_6t
Xbit_r241_c70 bl[70] br[70] wl[241] vdd gnd cell_6t
Xbit_r242_c70 bl[70] br[70] wl[242] vdd gnd cell_6t
Xbit_r243_c70 bl[70] br[70] wl[243] vdd gnd cell_6t
Xbit_r244_c70 bl[70] br[70] wl[244] vdd gnd cell_6t
Xbit_r245_c70 bl[70] br[70] wl[245] vdd gnd cell_6t
Xbit_r246_c70 bl[70] br[70] wl[246] vdd gnd cell_6t
Xbit_r247_c70 bl[70] br[70] wl[247] vdd gnd cell_6t
Xbit_r248_c70 bl[70] br[70] wl[248] vdd gnd cell_6t
Xbit_r249_c70 bl[70] br[70] wl[249] vdd gnd cell_6t
Xbit_r250_c70 bl[70] br[70] wl[250] vdd gnd cell_6t
Xbit_r251_c70 bl[70] br[70] wl[251] vdd gnd cell_6t
Xbit_r252_c70 bl[70] br[70] wl[252] vdd gnd cell_6t
Xbit_r253_c70 bl[70] br[70] wl[253] vdd gnd cell_6t
Xbit_r254_c70 bl[70] br[70] wl[254] vdd gnd cell_6t
Xbit_r255_c70 bl[70] br[70] wl[255] vdd gnd cell_6t
Xbit_r0_c71 bl[71] br[71] wl[0] vdd gnd cell_6t
Xbit_r1_c71 bl[71] br[71] wl[1] vdd gnd cell_6t
Xbit_r2_c71 bl[71] br[71] wl[2] vdd gnd cell_6t
Xbit_r3_c71 bl[71] br[71] wl[3] vdd gnd cell_6t
Xbit_r4_c71 bl[71] br[71] wl[4] vdd gnd cell_6t
Xbit_r5_c71 bl[71] br[71] wl[5] vdd gnd cell_6t
Xbit_r6_c71 bl[71] br[71] wl[6] vdd gnd cell_6t
Xbit_r7_c71 bl[71] br[71] wl[7] vdd gnd cell_6t
Xbit_r8_c71 bl[71] br[71] wl[8] vdd gnd cell_6t
Xbit_r9_c71 bl[71] br[71] wl[9] vdd gnd cell_6t
Xbit_r10_c71 bl[71] br[71] wl[10] vdd gnd cell_6t
Xbit_r11_c71 bl[71] br[71] wl[11] vdd gnd cell_6t
Xbit_r12_c71 bl[71] br[71] wl[12] vdd gnd cell_6t
Xbit_r13_c71 bl[71] br[71] wl[13] vdd gnd cell_6t
Xbit_r14_c71 bl[71] br[71] wl[14] vdd gnd cell_6t
Xbit_r15_c71 bl[71] br[71] wl[15] vdd gnd cell_6t
Xbit_r16_c71 bl[71] br[71] wl[16] vdd gnd cell_6t
Xbit_r17_c71 bl[71] br[71] wl[17] vdd gnd cell_6t
Xbit_r18_c71 bl[71] br[71] wl[18] vdd gnd cell_6t
Xbit_r19_c71 bl[71] br[71] wl[19] vdd gnd cell_6t
Xbit_r20_c71 bl[71] br[71] wl[20] vdd gnd cell_6t
Xbit_r21_c71 bl[71] br[71] wl[21] vdd gnd cell_6t
Xbit_r22_c71 bl[71] br[71] wl[22] vdd gnd cell_6t
Xbit_r23_c71 bl[71] br[71] wl[23] vdd gnd cell_6t
Xbit_r24_c71 bl[71] br[71] wl[24] vdd gnd cell_6t
Xbit_r25_c71 bl[71] br[71] wl[25] vdd gnd cell_6t
Xbit_r26_c71 bl[71] br[71] wl[26] vdd gnd cell_6t
Xbit_r27_c71 bl[71] br[71] wl[27] vdd gnd cell_6t
Xbit_r28_c71 bl[71] br[71] wl[28] vdd gnd cell_6t
Xbit_r29_c71 bl[71] br[71] wl[29] vdd gnd cell_6t
Xbit_r30_c71 bl[71] br[71] wl[30] vdd gnd cell_6t
Xbit_r31_c71 bl[71] br[71] wl[31] vdd gnd cell_6t
Xbit_r32_c71 bl[71] br[71] wl[32] vdd gnd cell_6t
Xbit_r33_c71 bl[71] br[71] wl[33] vdd gnd cell_6t
Xbit_r34_c71 bl[71] br[71] wl[34] vdd gnd cell_6t
Xbit_r35_c71 bl[71] br[71] wl[35] vdd gnd cell_6t
Xbit_r36_c71 bl[71] br[71] wl[36] vdd gnd cell_6t
Xbit_r37_c71 bl[71] br[71] wl[37] vdd gnd cell_6t
Xbit_r38_c71 bl[71] br[71] wl[38] vdd gnd cell_6t
Xbit_r39_c71 bl[71] br[71] wl[39] vdd gnd cell_6t
Xbit_r40_c71 bl[71] br[71] wl[40] vdd gnd cell_6t
Xbit_r41_c71 bl[71] br[71] wl[41] vdd gnd cell_6t
Xbit_r42_c71 bl[71] br[71] wl[42] vdd gnd cell_6t
Xbit_r43_c71 bl[71] br[71] wl[43] vdd gnd cell_6t
Xbit_r44_c71 bl[71] br[71] wl[44] vdd gnd cell_6t
Xbit_r45_c71 bl[71] br[71] wl[45] vdd gnd cell_6t
Xbit_r46_c71 bl[71] br[71] wl[46] vdd gnd cell_6t
Xbit_r47_c71 bl[71] br[71] wl[47] vdd gnd cell_6t
Xbit_r48_c71 bl[71] br[71] wl[48] vdd gnd cell_6t
Xbit_r49_c71 bl[71] br[71] wl[49] vdd gnd cell_6t
Xbit_r50_c71 bl[71] br[71] wl[50] vdd gnd cell_6t
Xbit_r51_c71 bl[71] br[71] wl[51] vdd gnd cell_6t
Xbit_r52_c71 bl[71] br[71] wl[52] vdd gnd cell_6t
Xbit_r53_c71 bl[71] br[71] wl[53] vdd gnd cell_6t
Xbit_r54_c71 bl[71] br[71] wl[54] vdd gnd cell_6t
Xbit_r55_c71 bl[71] br[71] wl[55] vdd gnd cell_6t
Xbit_r56_c71 bl[71] br[71] wl[56] vdd gnd cell_6t
Xbit_r57_c71 bl[71] br[71] wl[57] vdd gnd cell_6t
Xbit_r58_c71 bl[71] br[71] wl[58] vdd gnd cell_6t
Xbit_r59_c71 bl[71] br[71] wl[59] vdd gnd cell_6t
Xbit_r60_c71 bl[71] br[71] wl[60] vdd gnd cell_6t
Xbit_r61_c71 bl[71] br[71] wl[61] vdd gnd cell_6t
Xbit_r62_c71 bl[71] br[71] wl[62] vdd gnd cell_6t
Xbit_r63_c71 bl[71] br[71] wl[63] vdd gnd cell_6t
Xbit_r64_c71 bl[71] br[71] wl[64] vdd gnd cell_6t
Xbit_r65_c71 bl[71] br[71] wl[65] vdd gnd cell_6t
Xbit_r66_c71 bl[71] br[71] wl[66] vdd gnd cell_6t
Xbit_r67_c71 bl[71] br[71] wl[67] vdd gnd cell_6t
Xbit_r68_c71 bl[71] br[71] wl[68] vdd gnd cell_6t
Xbit_r69_c71 bl[71] br[71] wl[69] vdd gnd cell_6t
Xbit_r70_c71 bl[71] br[71] wl[70] vdd gnd cell_6t
Xbit_r71_c71 bl[71] br[71] wl[71] vdd gnd cell_6t
Xbit_r72_c71 bl[71] br[71] wl[72] vdd gnd cell_6t
Xbit_r73_c71 bl[71] br[71] wl[73] vdd gnd cell_6t
Xbit_r74_c71 bl[71] br[71] wl[74] vdd gnd cell_6t
Xbit_r75_c71 bl[71] br[71] wl[75] vdd gnd cell_6t
Xbit_r76_c71 bl[71] br[71] wl[76] vdd gnd cell_6t
Xbit_r77_c71 bl[71] br[71] wl[77] vdd gnd cell_6t
Xbit_r78_c71 bl[71] br[71] wl[78] vdd gnd cell_6t
Xbit_r79_c71 bl[71] br[71] wl[79] vdd gnd cell_6t
Xbit_r80_c71 bl[71] br[71] wl[80] vdd gnd cell_6t
Xbit_r81_c71 bl[71] br[71] wl[81] vdd gnd cell_6t
Xbit_r82_c71 bl[71] br[71] wl[82] vdd gnd cell_6t
Xbit_r83_c71 bl[71] br[71] wl[83] vdd gnd cell_6t
Xbit_r84_c71 bl[71] br[71] wl[84] vdd gnd cell_6t
Xbit_r85_c71 bl[71] br[71] wl[85] vdd gnd cell_6t
Xbit_r86_c71 bl[71] br[71] wl[86] vdd gnd cell_6t
Xbit_r87_c71 bl[71] br[71] wl[87] vdd gnd cell_6t
Xbit_r88_c71 bl[71] br[71] wl[88] vdd gnd cell_6t
Xbit_r89_c71 bl[71] br[71] wl[89] vdd gnd cell_6t
Xbit_r90_c71 bl[71] br[71] wl[90] vdd gnd cell_6t
Xbit_r91_c71 bl[71] br[71] wl[91] vdd gnd cell_6t
Xbit_r92_c71 bl[71] br[71] wl[92] vdd gnd cell_6t
Xbit_r93_c71 bl[71] br[71] wl[93] vdd gnd cell_6t
Xbit_r94_c71 bl[71] br[71] wl[94] vdd gnd cell_6t
Xbit_r95_c71 bl[71] br[71] wl[95] vdd gnd cell_6t
Xbit_r96_c71 bl[71] br[71] wl[96] vdd gnd cell_6t
Xbit_r97_c71 bl[71] br[71] wl[97] vdd gnd cell_6t
Xbit_r98_c71 bl[71] br[71] wl[98] vdd gnd cell_6t
Xbit_r99_c71 bl[71] br[71] wl[99] vdd gnd cell_6t
Xbit_r100_c71 bl[71] br[71] wl[100] vdd gnd cell_6t
Xbit_r101_c71 bl[71] br[71] wl[101] vdd gnd cell_6t
Xbit_r102_c71 bl[71] br[71] wl[102] vdd gnd cell_6t
Xbit_r103_c71 bl[71] br[71] wl[103] vdd gnd cell_6t
Xbit_r104_c71 bl[71] br[71] wl[104] vdd gnd cell_6t
Xbit_r105_c71 bl[71] br[71] wl[105] vdd gnd cell_6t
Xbit_r106_c71 bl[71] br[71] wl[106] vdd gnd cell_6t
Xbit_r107_c71 bl[71] br[71] wl[107] vdd gnd cell_6t
Xbit_r108_c71 bl[71] br[71] wl[108] vdd gnd cell_6t
Xbit_r109_c71 bl[71] br[71] wl[109] vdd gnd cell_6t
Xbit_r110_c71 bl[71] br[71] wl[110] vdd gnd cell_6t
Xbit_r111_c71 bl[71] br[71] wl[111] vdd gnd cell_6t
Xbit_r112_c71 bl[71] br[71] wl[112] vdd gnd cell_6t
Xbit_r113_c71 bl[71] br[71] wl[113] vdd gnd cell_6t
Xbit_r114_c71 bl[71] br[71] wl[114] vdd gnd cell_6t
Xbit_r115_c71 bl[71] br[71] wl[115] vdd gnd cell_6t
Xbit_r116_c71 bl[71] br[71] wl[116] vdd gnd cell_6t
Xbit_r117_c71 bl[71] br[71] wl[117] vdd gnd cell_6t
Xbit_r118_c71 bl[71] br[71] wl[118] vdd gnd cell_6t
Xbit_r119_c71 bl[71] br[71] wl[119] vdd gnd cell_6t
Xbit_r120_c71 bl[71] br[71] wl[120] vdd gnd cell_6t
Xbit_r121_c71 bl[71] br[71] wl[121] vdd gnd cell_6t
Xbit_r122_c71 bl[71] br[71] wl[122] vdd gnd cell_6t
Xbit_r123_c71 bl[71] br[71] wl[123] vdd gnd cell_6t
Xbit_r124_c71 bl[71] br[71] wl[124] vdd gnd cell_6t
Xbit_r125_c71 bl[71] br[71] wl[125] vdd gnd cell_6t
Xbit_r126_c71 bl[71] br[71] wl[126] vdd gnd cell_6t
Xbit_r127_c71 bl[71] br[71] wl[127] vdd gnd cell_6t
Xbit_r128_c71 bl[71] br[71] wl[128] vdd gnd cell_6t
Xbit_r129_c71 bl[71] br[71] wl[129] vdd gnd cell_6t
Xbit_r130_c71 bl[71] br[71] wl[130] vdd gnd cell_6t
Xbit_r131_c71 bl[71] br[71] wl[131] vdd gnd cell_6t
Xbit_r132_c71 bl[71] br[71] wl[132] vdd gnd cell_6t
Xbit_r133_c71 bl[71] br[71] wl[133] vdd gnd cell_6t
Xbit_r134_c71 bl[71] br[71] wl[134] vdd gnd cell_6t
Xbit_r135_c71 bl[71] br[71] wl[135] vdd gnd cell_6t
Xbit_r136_c71 bl[71] br[71] wl[136] vdd gnd cell_6t
Xbit_r137_c71 bl[71] br[71] wl[137] vdd gnd cell_6t
Xbit_r138_c71 bl[71] br[71] wl[138] vdd gnd cell_6t
Xbit_r139_c71 bl[71] br[71] wl[139] vdd gnd cell_6t
Xbit_r140_c71 bl[71] br[71] wl[140] vdd gnd cell_6t
Xbit_r141_c71 bl[71] br[71] wl[141] vdd gnd cell_6t
Xbit_r142_c71 bl[71] br[71] wl[142] vdd gnd cell_6t
Xbit_r143_c71 bl[71] br[71] wl[143] vdd gnd cell_6t
Xbit_r144_c71 bl[71] br[71] wl[144] vdd gnd cell_6t
Xbit_r145_c71 bl[71] br[71] wl[145] vdd gnd cell_6t
Xbit_r146_c71 bl[71] br[71] wl[146] vdd gnd cell_6t
Xbit_r147_c71 bl[71] br[71] wl[147] vdd gnd cell_6t
Xbit_r148_c71 bl[71] br[71] wl[148] vdd gnd cell_6t
Xbit_r149_c71 bl[71] br[71] wl[149] vdd gnd cell_6t
Xbit_r150_c71 bl[71] br[71] wl[150] vdd gnd cell_6t
Xbit_r151_c71 bl[71] br[71] wl[151] vdd gnd cell_6t
Xbit_r152_c71 bl[71] br[71] wl[152] vdd gnd cell_6t
Xbit_r153_c71 bl[71] br[71] wl[153] vdd gnd cell_6t
Xbit_r154_c71 bl[71] br[71] wl[154] vdd gnd cell_6t
Xbit_r155_c71 bl[71] br[71] wl[155] vdd gnd cell_6t
Xbit_r156_c71 bl[71] br[71] wl[156] vdd gnd cell_6t
Xbit_r157_c71 bl[71] br[71] wl[157] vdd gnd cell_6t
Xbit_r158_c71 bl[71] br[71] wl[158] vdd gnd cell_6t
Xbit_r159_c71 bl[71] br[71] wl[159] vdd gnd cell_6t
Xbit_r160_c71 bl[71] br[71] wl[160] vdd gnd cell_6t
Xbit_r161_c71 bl[71] br[71] wl[161] vdd gnd cell_6t
Xbit_r162_c71 bl[71] br[71] wl[162] vdd gnd cell_6t
Xbit_r163_c71 bl[71] br[71] wl[163] vdd gnd cell_6t
Xbit_r164_c71 bl[71] br[71] wl[164] vdd gnd cell_6t
Xbit_r165_c71 bl[71] br[71] wl[165] vdd gnd cell_6t
Xbit_r166_c71 bl[71] br[71] wl[166] vdd gnd cell_6t
Xbit_r167_c71 bl[71] br[71] wl[167] vdd gnd cell_6t
Xbit_r168_c71 bl[71] br[71] wl[168] vdd gnd cell_6t
Xbit_r169_c71 bl[71] br[71] wl[169] vdd gnd cell_6t
Xbit_r170_c71 bl[71] br[71] wl[170] vdd gnd cell_6t
Xbit_r171_c71 bl[71] br[71] wl[171] vdd gnd cell_6t
Xbit_r172_c71 bl[71] br[71] wl[172] vdd gnd cell_6t
Xbit_r173_c71 bl[71] br[71] wl[173] vdd gnd cell_6t
Xbit_r174_c71 bl[71] br[71] wl[174] vdd gnd cell_6t
Xbit_r175_c71 bl[71] br[71] wl[175] vdd gnd cell_6t
Xbit_r176_c71 bl[71] br[71] wl[176] vdd gnd cell_6t
Xbit_r177_c71 bl[71] br[71] wl[177] vdd gnd cell_6t
Xbit_r178_c71 bl[71] br[71] wl[178] vdd gnd cell_6t
Xbit_r179_c71 bl[71] br[71] wl[179] vdd gnd cell_6t
Xbit_r180_c71 bl[71] br[71] wl[180] vdd gnd cell_6t
Xbit_r181_c71 bl[71] br[71] wl[181] vdd gnd cell_6t
Xbit_r182_c71 bl[71] br[71] wl[182] vdd gnd cell_6t
Xbit_r183_c71 bl[71] br[71] wl[183] vdd gnd cell_6t
Xbit_r184_c71 bl[71] br[71] wl[184] vdd gnd cell_6t
Xbit_r185_c71 bl[71] br[71] wl[185] vdd gnd cell_6t
Xbit_r186_c71 bl[71] br[71] wl[186] vdd gnd cell_6t
Xbit_r187_c71 bl[71] br[71] wl[187] vdd gnd cell_6t
Xbit_r188_c71 bl[71] br[71] wl[188] vdd gnd cell_6t
Xbit_r189_c71 bl[71] br[71] wl[189] vdd gnd cell_6t
Xbit_r190_c71 bl[71] br[71] wl[190] vdd gnd cell_6t
Xbit_r191_c71 bl[71] br[71] wl[191] vdd gnd cell_6t
Xbit_r192_c71 bl[71] br[71] wl[192] vdd gnd cell_6t
Xbit_r193_c71 bl[71] br[71] wl[193] vdd gnd cell_6t
Xbit_r194_c71 bl[71] br[71] wl[194] vdd gnd cell_6t
Xbit_r195_c71 bl[71] br[71] wl[195] vdd gnd cell_6t
Xbit_r196_c71 bl[71] br[71] wl[196] vdd gnd cell_6t
Xbit_r197_c71 bl[71] br[71] wl[197] vdd gnd cell_6t
Xbit_r198_c71 bl[71] br[71] wl[198] vdd gnd cell_6t
Xbit_r199_c71 bl[71] br[71] wl[199] vdd gnd cell_6t
Xbit_r200_c71 bl[71] br[71] wl[200] vdd gnd cell_6t
Xbit_r201_c71 bl[71] br[71] wl[201] vdd gnd cell_6t
Xbit_r202_c71 bl[71] br[71] wl[202] vdd gnd cell_6t
Xbit_r203_c71 bl[71] br[71] wl[203] vdd gnd cell_6t
Xbit_r204_c71 bl[71] br[71] wl[204] vdd gnd cell_6t
Xbit_r205_c71 bl[71] br[71] wl[205] vdd gnd cell_6t
Xbit_r206_c71 bl[71] br[71] wl[206] vdd gnd cell_6t
Xbit_r207_c71 bl[71] br[71] wl[207] vdd gnd cell_6t
Xbit_r208_c71 bl[71] br[71] wl[208] vdd gnd cell_6t
Xbit_r209_c71 bl[71] br[71] wl[209] vdd gnd cell_6t
Xbit_r210_c71 bl[71] br[71] wl[210] vdd gnd cell_6t
Xbit_r211_c71 bl[71] br[71] wl[211] vdd gnd cell_6t
Xbit_r212_c71 bl[71] br[71] wl[212] vdd gnd cell_6t
Xbit_r213_c71 bl[71] br[71] wl[213] vdd gnd cell_6t
Xbit_r214_c71 bl[71] br[71] wl[214] vdd gnd cell_6t
Xbit_r215_c71 bl[71] br[71] wl[215] vdd gnd cell_6t
Xbit_r216_c71 bl[71] br[71] wl[216] vdd gnd cell_6t
Xbit_r217_c71 bl[71] br[71] wl[217] vdd gnd cell_6t
Xbit_r218_c71 bl[71] br[71] wl[218] vdd gnd cell_6t
Xbit_r219_c71 bl[71] br[71] wl[219] vdd gnd cell_6t
Xbit_r220_c71 bl[71] br[71] wl[220] vdd gnd cell_6t
Xbit_r221_c71 bl[71] br[71] wl[221] vdd gnd cell_6t
Xbit_r222_c71 bl[71] br[71] wl[222] vdd gnd cell_6t
Xbit_r223_c71 bl[71] br[71] wl[223] vdd gnd cell_6t
Xbit_r224_c71 bl[71] br[71] wl[224] vdd gnd cell_6t
Xbit_r225_c71 bl[71] br[71] wl[225] vdd gnd cell_6t
Xbit_r226_c71 bl[71] br[71] wl[226] vdd gnd cell_6t
Xbit_r227_c71 bl[71] br[71] wl[227] vdd gnd cell_6t
Xbit_r228_c71 bl[71] br[71] wl[228] vdd gnd cell_6t
Xbit_r229_c71 bl[71] br[71] wl[229] vdd gnd cell_6t
Xbit_r230_c71 bl[71] br[71] wl[230] vdd gnd cell_6t
Xbit_r231_c71 bl[71] br[71] wl[231] vdd gnd cell_6t
Xbit_r232_c71 bl[71] br[71] wl[232] vdd gnd cell_6t
Xbit_r233_c71 bl[71] br[71] wl[233] vdd gnd cell_6t
Xbit_r234_c71 bl[71] br[71] wl[234] vdd gnd cell_6t
Xbit_r235_c71 bl[71] br[71] wl[235] vdd gnd cell_6t
Xbit_r236_c71 bl[71] br[71] wl[236] vdd gnd cell_6t
Xbit_r237_c71 bl[71] br[71] wl[237] vdd gnd cell_6t
Xbit_r238_c71 bl[71] br[71] wl[238] vdd gnd cell_6t
Xbit_r239_c71 bl[71] br[71] wl[239] vdd gnd cell_6t
Xbit_r240_c71 bl[71] br[71] wl[240] vdd gnd cell_6t
Xbit_r241_c71 bl[71] br[71] wl[241] vdd gnd cell_6t
Xbit_r242_c71 bl[71] br[71] wl[242] vdd gnd cell_6t
Xbit_r243_c71 bl[71] br[71] wl[243] vdd gnd cell_6t
Xbit_r244_c71 bl[71] br[71] wl[244] vdd gnd cell_6t
Xbit_r245_c71 bl[71] br[71] wl[245] vdd gnd cell_6t
Xbit_r246_c71 bl[71] br[71] wl[246] vdd gnd cell_6t
Xbit_r247_c71 bl[71] br[71] wl[247] vdd gnd cell_6t
Xbit_r248_c71 bl[71] br[71] wl[248] vdd gnd cell_6t
Xbit_r249_c71 bl[71] br[71] wl[249] vdd gnd cell_6t
Xbit_r250_c71 bl[71] br[71] wl[250] vdd gnd cell_6t
Xbit_r251_c71 bl[71] br[71] wl[251] vdd gnd cell_6t
Xbit_r252_c71 bl[71] br[71] wl[252] vdd gnd cell_6t
Xbit_r253_c71 bl[71] br[71] wl[253] vdd gnd cell_6t
Xbit_r254_c71 bl[71] br[71] wl[254] vdd gnd cell_6t
Xbit_r255_c71 bl[71] br[71] wl[255] vdd gnd cell_6t
Xbit_r0_c72 bl[72] br[72] wl[0] vdd gnd cell_6t
Xbit_r1_c72 bl[72] br[72] wl[1] vdd gnd cell_6t
Xbit_r2_c72 bl[72] br[72] wl[2] vdd gnd cell_6t
Xbit_r3_c72 bl[72] br[72] wl[3] vdd gnd cell_6t
Xbit_r4_c72 bl[72] br[72] wl[4] vdd gnd cell_6t
Xbit_r5_c72 bl[72] br[72] wl[5] vdd gnd cell_6t
Xbit_r6_c72 bl[72] br[72] wl[6] vdd gnd cell_6t
Xbit_r7_c72 bl[72] br[72] wl[7] vdd gnd cell_6t
Xbit_r8_c72 bl[72] br[72] wl[8] vdd gnd cell_6t
Xbit_r9_c72 bl[72] br[72] wl[9] vdd gnd cell_6t
Xbit_r10_c72 bl[72] br[72] wl[10] vdd gnd cell_6t
Xbit_r11_c72 bl[72] br[72] wl[11] vdd gnd cell_6t
Xbit_r12_c72 bl[72] br[72] wl[12] vdd gnd cell_6t
Xbit_r13_c72 bl[72] br[72] wl[13] vdd gnd cell_6t
Xbit_r14_c72 bl[72] br[72] wl[14] vdd gnd cell_6t
Xbit_r15_c72 bl[72] br[72] wl[15] vdd gnd cell_6t
Xbit_r16_c72 bl[72] br[72] wl[16] vdd gnd cell_6t
Xbit_r17_c72 bl[72] br[72] wl[17] vdd gnd cell_6t
Xbit_r18_c72 bl[72] br[72] wl[18] vdd gnd cell_6t
Xbit_r19_c72 bl[72] br[72] wl[19] vdd gnd cell_6t
Xbit_r20_c72 bl[72] br[72] wl[20] vdd gnd cell_6t
Xbit_r21_c72 bl[72] br[72] wl[21] vdd gnd cell_6t
Xbit_r22_c72 bl[72] br[72] wl[22] vdd gnd cell_6t
Xbit_r23_c72 bl[72] br[72] wl[23] vdd gnd cell_6t
Xbit_r24_c72 bl[72] br[72] wl[24] vdd gnd cell_6t
Xbit_r25_c72 bl[72] br[72] wl[25] vdd gnd cell_6t
Xbit_r26_c72 bl[72] br[72] wl[26] vdd gnd cell_6t
Xbit_r27_c72 bl[72] br[72] wl[27] vdd gnd cell_6t
Xbit_r28_c72 bl[72] br[72] wl[28] vdd gnd cell_6t
Xbit_r29_c72 bl[72] br[72] wl[29] vdd gnd cell_6t
Xbit_r30_c72 bl[72] br[72] wl[30] vdd gnd cell_6t
Xbit_r31_c72 bl[72] br[72] wl[31] vdd gnd cell_6t
Xbit_r32_c72 bl[72] br[72] wl[32] vdd gnd cell_6t
Xbit_r33_c72 bl[72] br[72] wl[33] vdd gnd cell_6t
Xbit_r34_c72 bl[72] br[72] wl[34] vdd gnd cell_6t
Xbit_r35_c72 bl[72] br[72] wl[35] vdd gnd cell_6t
Xbit_r36_c72 bl[72] br[72] wl[36] vdd gnd cell_6t
Xbit_r37_c72 bl[72] br[72] wl[37] vdd gnd cell_6t
Xbit_r38_c72 bl[72] br[72] wl[38] vdd gnd cell_6t
Xbit_r39_c72 bl[72] br[72] wl[39] vdd gnd cell_6t
Xbit_r40_c72 bl[72] br[72] wl[40] vdd gnd cell_6t
Xbit_r41_c72 bl[72] br[72] wl[41] vdd gnd cell_6t
Xbit_r42_c72 bl[72] br[72] wl[42] vdd gnd cell_6t
Xbit_r43_c72 bl[72] br[72] wl[43] vdd gnd cell_6t
Xbit_r44_c72 bl[72] br[72] wl[44] vdd gnd cell_6t
Xbit_r45_c72 bl[72] br[72] wl[45] vdd gnd cell_6t
Xbit_r46_c72 bl[72] br[72] wl[46] vdd gnd cell_6t
Xbit_r47_c72 bl[72] br[72] wl[47] vdd gnd cell_6t
Xbit_r48_c72 bl[72] br[72] wl[48] vdd gnd cell_6t
Xbit_r49_c72 bl[72] br[72] wl[49] vdd gnd cell_6t
Xbit_r50_c72 bl[72] br[72] wl[50] vdd gnd cell_6t
Xbit_r51_c72 bl[72] br[72] wl[51] vdd gnd cell_6t
Xbit_r52_c72 bl[72] br[72] wl[52] vdd gnd cell_6t
Xbit_r53_c72 bl[72] br[72] wl[53] vdd gnd cell_6t
Xbit_r54_c72 bl[72] br[72] wl[54] vdd gnd cell_6t
Xbit_r55_c72 bl[72] br[72] wl[55] vdd gnd cell_6t
Xbit_r56_c72 bl[72] br[72] wl[56] vdd gnd cell_6t
Xbit_r57_c72 bl[72] br[72] wl[57] vdd gnd cell_6t
Xbit_r58_c72 bl[72] br[72] wl[58] vdd gnd cell_6t
Xbit_r59_c72 bl[72] br[72] wl[59] vdd gnd cell_6t
Xbit_r60_c72 bl[72] br[72] wl[60] vdd gnd cell_6t
Xbit_r61_c72 bl[72] br[72] wl[61] vdd gnd cell_6t
Xbit_r62_c72 bl[72] br[72] wl[62] vdd gnd cell_6t
Xbit_r63_c72 bl[72] br[72] wl[63] vdd gnd cell_6t
Xbit_r64_c72 bl[72] br[72] wl[64] vdd gnd cell_6t
Xbit_r65_c72 bl[72] br[72] wl[65] vdd gnd cell_6t
Xbit_r66_c72 bl[72] br[72] wl[66] vdd gnd cell_6t
Xbit_r67_c72 bl[72] br[72] wl[67] vdd gnd cell_6t
Xbit_r68_c72 bl[72] br[72] wl[68] vdd gnd cell_6t
Xbit_r69_c72 bl[72] br[72] wl[69] vdd gnd cell_6t
Xbit_r70_c72 bl[72] br[72] wl[70] vdd gnd cell_6t
Xbit_r71_c72 bl[72] br[72] wl[71] vdd gnd cell_6t
Xbit_r72_c72 bl[72] br[72] wl[72] vdd gnd cell_6t
Xbit_r73_c72 bl[72] br[72] wl[73] vdd gnd cell_6t
Xbit_r74_c72 bl[72] br[72] wl[74] vdd gnd cell_6t
Xbit_r75_c72 bl[72] br[72] wl[75] vdd gnd cell_6t
Xbit_r76_c72 bl[72] br[72] wl[76] vdd gnd cell_6t
Xbit_r77_c72 bl[72] br[72] wl[77] vdd gnd cell_6t
Xbit_r78_c72 bl[72] br[72] wl[78] vdd gnd cell_6t
Xbit_r79_c72 bl[72] br[72] wl[79] vdd gnd cell_6t
Xbit_r80_c72 bl[72] br[72] wl[80] vdd gnd cell_6t
Xbit_r81_c72 bl[72] br[72] wl[81] vdd gnd cell_6t
Xbit_r82_c72 bl[72] br[72] wl[82] vdd gnd cell_6t
Xbit_r83_c72 bl[72] br[72] wl[83] vdd gnd cell_6t
Xbit_r84_c72 bl[72] br[72] wl[84] vdd gnd cell_6t
Xbit_r85_c72 bl[72] br[72] wl[85] vdd gnd cell_6t
Xbit_r86_c72 bl[72] br[72] wl[86] vdd gnd cell_6t
Xbit_r87_c72 bl[72] br[72] wl[87] vdd gnd cell_6t
Xbit_r88_c72 bl[72] br[72] wl[88] vdd gnd cell_6t
Xbit_r89_c72 bl[72] br[72] wl[89] vdd gnd cell_6t
Xbit_r90_c72 bl[72] br[72] wl[90] vdd gnd cell_6t
Xbit_r91_c72 bl[72] br[72] wl[91] vdd gnd cell_6t
Xbit_r92_c72 bl[72] br[72] wl[92] vdd gnd cell_6t
Xbit_r93_c72 bl[72] br[72] wl[93] vdd gnd cell_6t
Xbit_r94_c72 bl[72] br[72] wl[94] vdd gnd cell_6t
Xbit_r95_c72 bl[72] br[72] wl[95] vdd gnd cell_6t
Xbit_r96_c72 bl[72] br[72] wl[96] vdd gnd cell_6t
Xbit_r97_c72 bl[72] br[72] wl[97] vdd gnd cell_6t
Xbit_r98_c72 bl[72] br[72] wl[98] vdd gnd cell_6t
Xbit_r99_c72 bl[72] br[72] wl[99] vdd gnd cell_6t
Xbit_r100_c72 bl[72] br[72] wl[100] vdd gnd cell_6t
Xbit_r101_c72 bl[72] br[72] wl[101] vdd gnd cell_6t
Xbit_r102_c72 bl[72] br[72] wl[102] vdd gnd cell_6t
Xbit_r103_c72 bl[72] br[72] wl[103] vdd gnd cell_6t
Xbit_r104_c72 bl[72] br[72] wl[104] vdd gnd cell_6t
Xbit_r105_c72 bl[72] br[72] wl[105] vdd gnd cell_6t
Xbit_r106_c72 bl[72] br[72] wl[106] vdd gnd cell_6t
Xbit_r107_c72 bl[72] br[72] wl[107] vdd gnd cell_6t
Xbit_r108_c72 bl[72] br[72] wl[108] vdd gnd cell_6t
Xbit_r109_c72 bl[72] br[72] wl[109] vdd gnd cell_6t
Xbit_r110_c72 bl[72] br[72] wl[110] vdd gnd cell_6t
Xbit_r111_c72 bl[72] br[72] wl[111] vdd gnd cell_6t
Xbit_r112_c72 bl[72] br[72] wl[112] vdd gnd cell_6t
Xbit_r113_c72 bl[72] br[72] wl[113] vdd gnd cell_6t
Xbit_r114_c72 bl[72] br[72] wl[114] vdd gnd cell_6t
Xbit_r115_c72 bl[72] br[72] wl[115] vdd gnd cell_6t
Xbit_r116_c72 bl[72] br[72] wl[116] vdd gnd cell_6t
Xbit_r117_c72 bl[72] br[72] wl[117] vdd gnd cell_6t
Xbit_r118_c72 bl[72] br[72] wl[118] vdd gnd cell_6t
Xbit_r119_c72 bl[72] br[72] wl[119] vdd gnd cell_6t
Xbit_r120_c72 bl[72] br[72] wl[120] vdd gnd cell_6t
Xbit_r121_c72 bl[72] br[72] wl[121] vdd gnd cell_6t
Xbit_r122_c72 bl[72] br[72] wl[122] vdd gnd cell_6t
Xbit_r123_c72 bl[72] br[72] wl[123] vdd gnd cell_6t
Xbit_r124_c72 bl[72] br[72] wl[124] vdd gnd cell_6t
Xbit_r125_c72 bl[72] br[72] wl[125] vdd gnd cell_6t
Xbit_r126_c72 bl[72] br[72] wl[126] vdd gnd cell_6t
Xbit_r127_c72 bl[72] br[72] wl[127] vdd gnd cell_6t
Xbit_r128_c72 bl[72] br[72] wl[128] vdd gnd cell_6t
Xbit_r129_c72 bl[72] br[72] wl[129] vdd gnd cell_6t
Xbit_r130_c72 bl[72] br[72] wl[130] vdd gnd cell_6t
Xbit_r131_c72 bl[72] br[72] wl[131] vdd gnd cell_6t
Xbit_r132_c72 bl[72] br[72] wl[132] vdd gnd cell_6t
Xbit_r133_c72 bl[72] br[72] wl[133] vdd gnd cell_6t
Xbit_r134_c72 bl[72] br[72] wl[134] vdd gnd cell_6t
Xbit_r135_c72 bl[72] br[72] wl[135] vdd gnd cell_6t
Xbit_r136_c72 bl[72] br[72] wl[136] vdd gnd cell_6t
Xbit_r137_c72 bl[72] br[72] wl[137] vdd gnd cell_6t
Xbit_r138_c72 bl[72] br[72] wl[138] vdd gnd cell_6t
Xbit_r139_c72 bl[72] br[72] wl[139] vdd gnd cell_6t
Xbit_r140_c72 bl[72] br[72] wl[140] vdd gnd cell_6t
Xbit_r141_c72 bl[72] br[72] wl[141] vdd gnd cell_6t
Xbit_r142_c72 bl[72] br[72] wl[142] vdd gnd cell_6t
Xbit_r143_c72 bl[72] br[72] wl[143] vdd gnd cell_6t
Xbit_r144_c72 bl[72] br[72] wl[144] vdd gnd cell_6t
Xbit_r145_c72 bl[72] br[72] wl[145] vdd gnd cell_6t
Xbit_r146_c72 bl[72] br[72] wl[146] vdd gnd cell_6t
Xbit_r147_c72 bl[72] br[72] wl[147] vdd gnd cell_6t
Xbit_r148_c72 bl[72] br[72] wl[148] vdd gnd cell_6t
Xbit_r149_c72 bl[72] br[72] wl[149] vdd gnd cell_6t
Xbit_r150_c72 bl[72] br[72] wl[150] vdd gnd cell_6t
Xbit_r151_c72 bl[72] br[72] wl[151] vdd gnd cell_6t
Xbit_r152_c72 bl[72] br[72] wl[152] vdd gnd cell_6t
Xbit_r153_c72 bl[72] br[72] wl[153] vdd gnd cell_6t
Xbit_r154_c72 bl[72] br[72] wl[154] vdd gnd cell_6t
Xbit_r155_c72 bl[72] br[72] wl[155] vdd gnd cell_6t
Xbit_r156_c72 bl[72] br[72] wl[156] vdd gnd cell_6t
Xbit_r157_c72 bl[72] br[72] wl[157] vdd gnd cell_6t
Xbit_r158_c72 bl[72] br[72] wl[158] vdd gnd cell_6t
Xbit_r159_c72 bl[72] br[72] wl[159] vdd gnd cell_6t
Xbit_r160_c72 bl[72] br[72] wl[160] vdd gnd cell_6t
Xbit_r161_c72 bl[72] br[72] wl[161] vdd gnd cell_6t
Xbit_r162_c72 bl[72] br[72] wl[162] vdd gnd cell_6t
Xbit_r163_c72 bl[72] br[72] wl[163] vdd gnd cell_6t
Xbit_r164_c72 bl[72] br[72] wl[164] vdd gnd cell_6t
Xbit_r165_c72 bl[72] br[72] wl[165] vdd gnd cell_6t
Xbit_r166_c72 bl[72] br[72] wl[166] vdd gnd cell_6t
Xbit_r167_c72 bl[72] br[72] wl[167] vdd gnd cell_6t
Xbit_r168_c72 bl[72] br[72] wl[168] vdd gnd cell_6t
Xbit_r169_c72 bl[72] br[72] wl[169] vdd gnd cell_6t
Xbit_r170_c72 bl[72] br[72] wl[170] vdd gnd cell_6t
Xbit_r171_c72 bl[72] br[72] wl[171] vdd gnd cell_6t
Xbit_r172_c72 bl[72] br[72] wl[172] vdd gnd cell_6t
Xbit_r173_c72 bl[72] br[72] wl[173] vdd gnd cell_6t
Xbit_r174_c72 bl[72] br[72] wl[174] vdd gnd cell_6t
Xbit_r175_c72 bl[72] br[72] wl[175] vdd gnd cell_6t
Xbit_r176_c72 bl[72] br[72] wl[176] vdd gnd cell_6t
Xbit_r177_c72 bl[72] br[72] wl[177] vdd gnd cell_6t
Xbit_r178_c72 bl[72] br[72] wl[178] vdd gnd cell_6t
Xbit_r179_c72 bl[72] br[72] wl[179] vdd gnd cell_6t
Xbit_r180_c72 bl[72] br[72] wl[180] vdd gnd cell_6t
Xbit_r181_c72 bl[72] br[72] wl[181] vdd gnd cell_6t
Xbit_r182_c72 bl[72] br[72] wl[182] vdd gnd cell_6t
Xbit_r183_c72 bl[72] br[72] wl[183] vdd gnd cell_6t
Xbit_r184_c72 bl[72] br[72] wl[184] vdd gnd cell_6t
Xbit_r185_c72 bl[72] br[72] wl[185] vdd gnd cell_6t
Xbit_r186_c72 bl[72] br[72] wl[186] vdd gnd cell_6t
Xbit_r187_c72 bl[72] br[72] wl[187] vdd gnd cell_6t
Xbit_r188_c72 bl[72] br[72] wl[188] vdd gnd cell_6t
Xbit_r189_c72 bl[72] br[72] wl[189] vdd gnd cell_6t
Xbit_r190_c72 bl[72] br[72] wl[190] vdd gnd cell_6t
Xbit_r191_c72 bl[72] br[72] wl[191] vdd gnd cell_6t
Xbit_r192_c72 bl[72] br[72] wl[192] vdd gnd cell_6t
Xbit_r193_c72 bl[72] br[72] wl[193] vdd gnd cell_6t
Xbit_r194_c72 bl[72] br[72] wl[194] vdd gnd cell_6t
Xbit_r195_c72 bl[72] br[72] wl[195] vdd gnd cell_6t
Xbit_r196_c72 bl[72] br[72] wl[196] vdd gnd cell_6t
Xbit_r197_c72 bl[72] br[72] wl[197] vdd gnd cell_6t
Xbit_r198_c72 bl[72] br[72] wl[198] vdd gnd cell_6t
Xbit_r199_c72 bl[72] br[72] wl[199] vdd gnd cell_6t
Xbit_r200_c72 bl[72] br[72] wl[200] vdd gnd cell_6t
Xbit_r201_c72 bl[72] br[72] wl[201] vdd gnd cell_6t
Xbit_r202_c72 bl[72] br[72] wl[202] vdd gnd cell_6t
Xbit_r203_c72 bl[72] br[72] wl[203] vdd gnd cell_6t
Xbit_r204_c72 bl[72] br[72] wl[204] vdd gnd cell_6t
Xbit_r205_c72 bl[72] br[72] wl[205] vdd gnd cell_6t
Xbit_r206_c72 bl[72] br[72] wl[206] vdd gnd cell_6t
Xbit_r207_c72 bl[72] br[72] wl[207] vdd gnd cell_6t
Xbit_r208_c72 bl[72] br[72] wl[208] vdd gnd cell_6t
Xbit_r209_c72 bl[72] br[72] wl[209] vdd gnd cell_6t
Xbit_r210_c72 bl[72] br[72] wl[210] vdd gnd cell_6t
Xbit_r211_c72 bl[72] br[72] wl[211] vdd gnd cell_6t
Xbit_r212_c72 bl[72] br[72] wl[212] vdd gnd cell_6t
Xbit_r213_c72 bl[72] br[72] wl[213] vdd gnd cell_6t
Xbit_r214_c72 bl[72] br[72] wl[214] vdd gnd cell_6t
Xbit_r215_c72 bl[72] br[72] wl[215] vdd gnd cell_6t
Xbit_r216_c72 bl[72] br[72] wl[216] vdd gnd cell_6t
Xbit_r217_c72 bl[72] br[72] wl[217] vdd gnd cell_6t
Xbit_r218_c72 bl[72] br[72] wl[218] vdd gnd cell_6t
Xbit_r219_c72 bl[72] br[72] wl[219] vdd gnd cell_6t
Xbit_r220_c72 bl[72] br[72] wl[220] vdd gnd cell_6t
Xbit_r221_c72 bl[72] br[72] wl[221] vdd gnd cell_6t
Xbit_r222_c72 bl[72] br[72] wl[222] vdd gnd cell_6t
Xbit_r223_c72 bl[72] br[72] wl[223] vdd gnd cell_6t
Xbit_r224_c72 bl[72] br[72] wl[224] vdd gnd cell_6t
Xbit_r225_c72 bl[72] br[72] wl[225] vdd gnd cell_6t
Xbit_r226_c72 bl[72] br[72] wl[226] vdd gnd cell_6t
Xbit_r227_c72 bl[72] br[72] wl[227] vdd gnd cell_6t
Xbit_r228_c72 bl[72] br[72] wl[228] vdd gnd cell_6t
Xbit_r229_c72 bl[72] br[72] wl[229] vdd gnd cell_6t
Xbit_r230_c72 bl[72] br[72] wl[230] vdd gnd cell_6t
Xbit_r231_c72 bl[72] br[72] wl[231] vdd gnd cell_6t
Xbit_r232_c72 bl[72] br[72] wl[232] vdd gnd cell_6t
Xbit_r233_c72 bl[72] br[72] wl[233] vdd gnd cell_6t
Xbit_r234_c72 bl[72] br[72] wl[234] vdd gnd cell_6t
Xbit_r235_c72 bl[72] br[72] wl[235] vdd gnd cell_6t
Xbit_r236_c72 bl[72] br[72] wl[236] vdd gnd cell_6t
Xbit_r237_c72 bl[72] br[72] wl[237] vdd gnd cell_6t
Xbit_r238_c72 bl[72] br[72] wl[238] vdd gnd cell_6t
Xbit_r239_c72 bl[72] br[72] wl[239] vdd gnd cell_6t
Xbit_r240_c72 bl[72] br[72] wl[240] vdd gnd cell_6t
Xbit_r241_c72 bl[72] br[72] wl[241] vdd gnd cell_6t
Xbit_r242_c72 bl[72] br[72] wl[242] vdd gnd cell_6t
Xbit_r243_c72 bl[72] br[72] wl[243] vdd gnd cell_6t
Xbit_r244_c72 bl[72] br[72] wl[244] vdd gnd cell_6t
Xbit_r245_c72 bl[72] br[72] wl[245] vdd gnd cell_6t
Xbit_r246_c72 bl[72] br[72] wl[246] vdd gnd cell_6t
Xbit_r247_c72 bl[72] br[72] wl[247] vdd gnd cell_6t
Xbit_r248_c72 bl[72] br[72] wl[248] vdd gnd cell_6t
Xbit_r249_c72 bl[72] br[72] wl[249] vdd gnd cell_6t
Xbit_r250_c72 bl[72] br[72] wl[250] vdd gnd cell_6t
Xbit_r251_c72 bl[72] br[72] wl[251] vdd gnd cell_6t
Xbit_r252_c72 bl[72] br[72] wl[252] vdd gnd cell_6t
Xbit_r253_c72 bl[72] br[72] wl[253] vdd gnd cell_6t
Xbit_r254_c72 bl[72] br[72] wl[254] vdd gnd cell_6t
Xbit_r255_c72 bl[72] br[72] wl[255] vdd gnd cell_6t
Xbit_r0_c73 bl[73] br[73] wl[0] vdd gnd cell_6t
Xbit_r1_c73 bl[73] br[73] wl[1] vdd gnd cell_6t
Xbit_r2_c73 bl[73] br[73] wl[2] vdd gnd cell_6t
Xbit_r3_c73 bl[73] br[73] wl[3] vdd gnd cell_6t
Xbit_r4_c73 bl[73] br[73] wl[4] vdd gnd cell_6t
Xbit_r5_c73 bl[73] br[73] wl[5] vdd gnd cell_6t
Xbit_r6_c73 bl[73] br[73] wl[6] vdd gnd cell_6t
Xbit_r7_c73 bl[73] br[73] wl[7] vdd gnd cell_6t
Xbit_r8_c73 bl[73] br[73] wl[8] vdd gnd cell_6t
Xbit_r9_c73 bl[73] br[73] wl[9] vdd gnd cell_6t
Xbit_r10_c73 bl[73] br[73] wl[10] vdd gnd cell_6t
Xbit_r11_c73 bl[73] br[73] wl[11] vdd gnd cell_6t
Xbit_r12_c73 bl[73] br[73] wl[12] vdd gnd cell_6t
Xbit_r13_c73 bl[73] br[73] wl[13] vdd gnd cell_6t
Xbit_r14_c73 bl[73] br[73] wl[14] vdd gnd cell_6t
Xbit_r15_c73 bl[73] br[73] wl[15] vdd gnd cell_6t
Xbit_r16_c73 bl[73] br[73] wl[16] vdd gnd cell_6t
Xbit_r17_c73 bl[73] br[73] wl[17] vdd gnd cell_6t
Xbit_r18_c73 bl[73] br[73] wl[18] vdd gnd cell_6t
Xbit_r19_c73 bl[73] br[73] wl[19] vdd gnd cell_6t
Xbit_r20_c73 bl[73] br[73] wl[20] vdd gnd cell_6t
Xbit_r21_c73 bl[73] br[73] wl[21] vdd gnd cell_6t
Xbit_r22_c73 bl[73] br[73] wl[22] vdd gnd cell_6t
Xbit_r23_c73 bl[73] br[73] wl[23] vdd gnd cell_6t
Xbit_r24_c73 bl[73] br[73] wl[24] vdd gnd cell_6t
Xbit_r25_c73 bl[73] br[73] wl[25] vdd gnd cell_6t
Xbit_r26_c73 bl[73] br[73] wl[26] vdd gnd cell_6t
Xbit_r27_c73 bl[73] br[73] wl[27] vdd gnd cell_6t
Xbit_r28_c73 bl[73] br[73] wl[28] vdd gnd cell_6t
Xbit_r29_c73 bl[73] br[73] wl[29] vdd gnd cell_6t
Xbit_r30_c73 bl[73] br[73] wl[30] vdd gnd cell_6t
Xbit_r31_c73 bl[73] br[73] wl[31] vdd gnd cell_6t
Xbit_r32_c73 bl[73] br[73] wl[32] vdd gnd cell_6t
Xbit_r33_c73 bl[73] br[73] wl[33] vdd gnd cell_6t
Xbit_r34_c73 bl[73] br[73] wl[34] vdd gnd cell_6t
Xbit_r35_c73 bl[73] br[73] wl[35] vdd gnd cell_6t
Xbit_r36_c73 bl[73] br[73] wl[36] vdd gnd cell_6t
Xbit_r37_c73 bl[73] br[73] wl[37] vdd gnd cell_6t
Xbit_r38_c73 bl[73] br[73] wl[38] vdd gnd cell_6t
Xbit_r39_c73 bl[73] br[73] wl[39] vdd gnd cell_6t
Xbit_r40_c73 bl[73] br[73] wl[40] vdd gnd cell_6t
Xbit_r41_c73 bl[73] br[73] wl[41] vdd gnd cell_6t
Xbit_r42_c73 bl[73] br[73] wl[42] vdd gnd cell_6t
Xbit_r43_c73 bl[73] br[73] wl[43] vdd gnd cell_6t
Xbit_r44_c73 bl[73] br[73] wl[44] vdd gnd cell_6t
Xbit_r45_c73 bl[73] br[73] wl[45] vdd gnd cell_6t
Xbit_r46_c73 bl[73] br[73] wl[46] vdd gnd cell_6t
Xbit_r47_c73 bl[73] br[73] wl[47] vdd gnd cell_6t
Xbit_r48_c73 bl[73] br[73] wl[48] vdd gnd cell_6t
Xbit_r49_c73 bl[73] br[73] wl[49] vdd gnd cell_6t
Xbit_r50_c73 bl[73] br[73] wl[50] vdd gnd cell_6t
Xbit_r51_c73 bl[73] br[73] wl[51] vdd gnd cell_6t
Xbit_r52_c73 bl[73] br[73] wl[52] vdd gnd cell_6t
Xbit_r53_c73 bl[73] br[73] wl[53] vdd gnd cell_6t
Xbit_r54_c73 bl[73] br[73] wl[54] vdd gnd cell_6t
Xbit_r55_c73 bl[73] br[73] wl[55] vdd gnd cell_6t
Xbit_r56_c73 bl[73] br[73] wl[56] vdd gnd cell_6t
Xbit_r57_c73 bl[73] br[73] wl[57] vdd gnd cell_6t
Xbit_r58_c73 bl[73] br[73] wl[58] vdd gnd cell_6t
Xbit_r59_c73 bl[73] br[73] wl[59] vdd gnd cell_6t
Xbit_r60_c73 bl[73] br[73] wl[60] vdd gnd cell_6t
Xbit_r61_c73 bl[73] br[73] wl[61] vdd gnd cell_6t
Xbit_r62_c73 bl[73] br[73] wl[62] vdd gnd cell_6t
Xbit_r63_c73 bl[73] br[73] wl[63] vdd gnd cell_6t
Xbit_r64_c73 bl[73] br[73] wl[64] vdd gnd cell_6t
Xbit_r65_c73 bl[73] br[73] wl[65] vdd gnd cell_6t
Xbit_r66_c73 bl[73] br[73] wl[66] vdd gnd cell_6t
Xbit_r67_c73 bl[73] br[73] wl[67] vdd gnd cell_6t
Xbit_r68_c73 bl[73] br[73] wl[68] vdd gnd cell_6t
Xbit_r69_c73 bl[73] br[73] wl[69] vdd gnd cell_6t
Xbit_r70_c73 bl[73] br[73] wl[70] vdd gnd cell_6t
Xbit_r71_c73 bl[73] br[73] wl[71] vdd gnd cell_6t
Xbit_r72_c73 bl[73] br[73] wl[72] vdd gnd cell_6t
Xbit_r73_c73 bl[73] br[73] wl[73] vdd gnd cell_6t
Xbit_r74_c73 bl[73] br[73] wl[74] vdd gnd cell_6t
Xbit_r75_c73 bl[73] br[73] wl[75] vdd gnd cell_6t
Xbit_r76_c73 bl[73] br[73] wl[76] vdd gnd cell_6t
Xbit_r77_c73 bl[73] br[73] wl[77] vdd gnd cell_6t
Xbit_r78_c73 bl[73] br[73] wl[78] vdd gnd cell_6t
Xbit_r79_c73 bl[73] br[73] wl[79] vdd gnd cell_6t
Xbit_r80_c73 bl[73] br[73] wl[80] vdd gnd cell_6t
Xbit_r81_c73 bl[73] br[73] wl[81] vdd gnd cell_6t
Xbit_r82_c73 bl[73] br[73] wl[82] vdd gnd cell_6t
Xbit_r83_c73 bl[73] br[73] wl[83] vdd gnd cell_6t
Xbit_r84_c73 bl[73] br[73] wl[84] vdd gnd cell_6t
Xbit_r85_c73 bl[73] br[73] wl[85] vdd gnd cell_6t
Xbit_r86_c73 bl[73] br[73] wl[86] vdd gnd cell_6t
Xbit_r87_c73 bl[73] br[73] wl[87] vdd gnd cell_6t
Xbit_r88_c73 bl[73] br[73] wl[88] vdd gnd cell_6t
Xbit_r89_c73 bl[73] br[73] wl[89] vdd gnd cell_6t
Xbit_r90_c73 bl[73] br[73] wl[90] vdd gnd cell_6t
Xbit_r91_c73 bl[73] br[73] wl[91] vdd gnd cell_6t
Xbit_r92_c73 bl[73] br[73] wl[92] vdd gnd cell_6t
Xbit_r93_c73 bl[73] br[73] wl[93] vdd gnd cell_6t
Xbit_r94_c73 bl[73] br[73] wl[94] vdd gnd cell_6t
Xbit_r95_c73 bl[73] br[73] wl[95] vdd gnd cell_6t
Xbit_r96_c73 bl[73] br[73] wl[96] vdd gnd cell_6t
Xbit_r97_c73 bl[73] br[73] wl[97] vdd gnd cell_6t
Xbit_r98_c73 bl[73] br[73] wl[98] vdd gnd cell_6t
Xbit_r99_c73 bl[73] br[73] wl[99] vdd gnd cell_6t
Xbit_r100_c73 bl[73] br[73] wl[100] vdd gnd cell_6t
Xbit_r101_c73 bl[73] br[73] wl[101] vdd gnd cell_6t
Xbit_r102_c73 bl[73] br[73] wl[102] vdd gnd cell_6t
Xbit_r103_c73 bl[73] br[73] wl[103] vdd gnd cell_6t
Xbit_r104_c73 bl[73] br[73] wl[104] vdd gnd cell_6t
Xbit_r105_c73 bl[73] br[73] wl[105] vdd gnd cell_6t
Xbit_r106_c73 bl[73] br[73] wl[106] vdd gnd cell_6t
Xbit_r107_c73 bl[73] br[73] wl[107] vdd gnd cell_6t
Xbit_r108_c73 bl[73] br[73] wl[108] vdd gnd cell_6t
Xbit_r109_c73 bl[73] br[73] wl[109] vdd gnd cell_6t
Xbit_r110_c73 bl[73] br[73] wl[110] vdd gnd cell_6t
Xbit_r111_c73 bl[73] br[73] wl[111] vdd gnd cell_6t
Xbit_r112_c73 bl[73] br[73] wl[112] vdd gnd cell_6t
Xbit_r113_c73 bl[73] br[73] wl[113] vdd gnd cell_6t
Xbit_r114_c73 bl[73] br[73] wl[114] vdd gnd cell_6t
Xbit_r115_c73 bl[73] br[73] wl[115] vdd gnd cell_6t
Xbit_r116_c73 bl[73] br[73] wl[116] vdd gnd cell_6t
Xbit_r117_c73 bl[73] br[73] wl[117] vdd gnd cell_6t
Xbit_r118_c73 bl[73] br[73] wl[118] vdd gnd cell_6t
Xbit_r119_c73 bl[73] br[73] wl[119] vdd gnd cell_6t
Xbit_r120_c73 bl[73] br[73] wl[120] vdd gnd cell_6t
Xbit_r121_c73 bl[73] br[73] wl[121] vdd gnd cell_6t
Xbit_r122_c73 bl[73] br[73] wl[122] vdd gnd cell_6t
Xbit_r123_c73 bl[73] br[73] wl[123] vdd gnd cell_6t
Xbit_r124_c73 bl[73] br[73] wl[124] vdd gnd cell_6t
Xbit_r125_c73 bl[73] br[73] wl[125] vdd gnd cell_6t
Xbit_r126_c73 bl[73] br[73] wl[126] vdd gnd cell_6t
Xbit_r127_c73 bl[73] br[73] wl[127] vdd gnd cell_6t
Xbit_r128_c73 bl[73] br[73] wl[128] vdd gnd cell_6t
Xbit_r129_c73 bl[73] br[73] wl[129] vdd gnd cell_6t
Xbit_r130_c73 bl[73] br[73] wl[130] vdd gnd cell_6t
Xbit_r131_c73 bl[73] br[73] wl[131] vdd gnd cell_6t
Xbit_r132_c73 bl[73] br[73] wl[132] vdd gnd cell_6t
Xbit_r133_c73 bl[73] br[73] wl[133] vdd gnd cell_6t
Xbit_r134_c73 bl[73] br[73] wl[134] vdd gnd cell_6t
Xbit_r135_c73 bl[73] br[73] wl[135] vdd gnd cell_6t
Xbit_r136_c73 bl[73] br[73] wl[136] vdd gnd cell_6t
Xbit_r137_c73 bl[73] br[73] wl[137] vdd gnd cell_6t
Xbit_r138_c73 bl[73] br[73] wl[138] vdd gnd cell_6t
Xbit_r139_c73 bl[73] br[73] wl[139] vdd gnd cell_6t
Xbit_r140_c73 bl[73] br[73] wl[140] vdd gnd cell_6t
Xbit_r141_c73 bl[73] br[73] wl[141] vdd gnd cell_6t
Xbit_r142_c73 bl[73] br[73] wl[142] vdd gnd cell_6t
Xbit_r143_c73 bl[73] br[73] wl[143] vdd gnd cell_6t
Xbit_r144_c73 bl[73] br[73] wl[144] vdd gnd cell_6t
Xbit_r145_c73 bl[73] br[73] wl[145] vdd gnd cell_6t
Xbit_r146_c73 bl[73] br[73] wl[146] vdd gnd cell_6t
Xbit_r147_c73 bl[73] br[73] wl[147] vdd gnd cell_6t
Xbit_r148_c73 bl[73] br[73] wl[148] vdd gnd cell_6t
Xbit_r149_c73 bl[73] br[73] wl[149] vdd gnd cell_6t
Xbit_r150_c73 bl[73] br[73] wl[150] vdd gnd cell_6t
Xbit_r151_c73 bl[73] br[73] wl[151] vdd gnd cell_6t
Xbit_r152_c73 bl[73] br[73] wl[152] vdd gnd cell_6t
Xbit_r153_c73 bl[73] br[73] wl[153] vdd gnd cell_6t
Xbit_r154_c73 bl[73] br[73] wl[154] vdd gnd cell_6t
Xbit_r155_c73 bl[73] br[73] wl[155] vdd gnd cell_6t
Xbit_r156_c73 bl[73] br[73] wl[156] vdd gnd cell_6t
Xbit_r157_c73 bl[73] br[73] wl[157] vdd gnd cell_6t
Xbit_r158_c73 bl[73] br[73] wl[158] vdd gnd cell_6t
Xbit_r159_c73 bl[73] br[73] wl[159] vdd gnd cell_6t
Xbit_r160_c73 bl[73] br[73] wl[160] vdd gnd cell_6t
Xbit_r161_c73 bl[73] br[73] wl[161] vdd gnd cell_6t
Xbit_r162_c73 bl[73] br[73] wl[162] vdd gnd cell_6t
Xbit_r163_c73 bl[73] br[73] wl[163] vdd gnd cell_6t
Xbit_r164_c73 bl[73] br[73] wl[164] vdd gnd cell_6t
Xbit_r165_c73 bl[73] br[73] wl[165] vdd gnd cell_6t
Xbit_r166_c73 bl[73] br[73] wl[166] vdd gnd cell_6t
Xbit_r167_c73 bl[73] br[73] wl[167] vdd gnd cell_6t
Xbit_r168_c73 bl[73] br[73] wl[168] vdd gnd cell_6t
Xbit_r169_c73 bl[73] br[73] wl[169] vdd gnd cell_6t
Xbit_r170_c73 bl[73] br[73] wl[170] vdd gnd cell_6t
Xbit_r171_c73 bl[73] br[73] wl[171] vdd gnd cell_6t
Xbit_r172_c73 bl[73] br[73] wl[172] vdd gnd cell_6t
Xbit_r173_c73 bl[73] br[73] wl[173] vdd gnd cell_6t
Xbit_r174_c73 bl[73] br[73] wl[174] vdd gnd cell_6t
Xbit_r175_c73 bl[73] br[73] wl[175] vdd gnd cell_6t
Xbit_r176_c73 bl[73] br[73] wl[176] vdd gnd cell_6t
Xbit_r177_c73 bl[73] br[73] wl[177] vdd gnd cell_6t
Xbit_r178_c73 bl[73] br[73] wl[178] vdd gnd cell_6t
Xbit_r179_c73 bl[73] br[73] wl[179] vdd gnd cell_6t
Xbit_r180_c73 bl[73] br[73] wl[180] vdd gnd cell_6t
Xbit_r181_c73 bl[73] br[73] wl[181] vdd gnd cell_6t
Xbit_r182_c73 bl[73] br[73] wl[182] vdd gnd cell_6t
Xbit_r183_c73 bl[73] br[73] wl[183] vdd gnd cell_6t
Xbit_r184_c73 bl[73] br[73] wl[184] vdd gnd cell_6t
Xbit_r185_c73 bl[73] br[73] wl[185] vdd gnd cell_6t
Xbit_r186_c73 bl[73] br[73] wl[186] vdd gnd cell_6t
Xbit_r187_c73 bl[73] br[73] wl[187] vdd gnd cell_6t
Xbit_r188_c73 bl[73] br[73] wl[188] vdd gnd cell_6t
Xbit_r189_c73 bl[73] br[73] wl[189] vdd gnd cell_6t
Xbit_r190_c73 bl[73] br[73] wl[190] vdd gnd cell_6t
Xbit_r191_c73 bl[73] br[73] wl[191] vdd gnd cell_6t
Xbit_r192_c73 bl[73] br[73] wl[192] vdd gnd cell_6t
Xbit_r193_c73 bl[73] br[73] wl[193] vdd gnd cell_6t
Xbit_r194_c73 bl[73] br[73] wl[194] vdd gnd cell_6t
Xbit_r195_c73 bl[73] br[73] wl[195] vdd gnd cell_6t
Xbit_r196_c73 bl[73] br[73] wl[196] vdd gnd cell_6t
Xbit_r197_c73 bl[73] br[73] wl[197] vdd gnd cell_6t
Xbit_r198_c73 bl[73] br[73] wl[198] vdd gnd cell_6t
Xbit_r199_c73 bl[73] br[73] wl[199] vdd gnd cell_6t
Xbit_r200_c73 bl[73] br[73] wl[200] vdd gnd cell_6t
Xbit_r201_c73 bl[73] br[73] wl[201] vdd gnd cell_6t
Xbit_r202_c73 bl[73] br[73] wl[202] vdd gnd cell_6t
Xbit_r203_c73 bl[73] br[73] wl[203] vdd gnd cell_6t
Xbit_r204_c73 bl[73] br[73] wl[204] vdd gnd cell_6t
Xbit_r205_c73 bl[73] br[73] wl[205] vdd gnd cell_6t
Xbit_r206_c73 bl[73] br[73] wl[206] vdd gnd cell_6t
Xbit_r207_c73 bl[73] br[73] wl[207] vdd gnd cell_6t
Xbit_r208_c73 bl[73] br[73] wl[208] vdd gnd cell_6t
Xbit_r209_c73 bl[73] br[73] wl[209] vdd gnd cell_6t
Xbit_r210_c73 bl[73] br[73] wl[210] vdd gnd cell_6t
Xbit_r211_c73 bl[73] br[73] wl[211] vdd gnd cell_6t
Xbit_r212_c73 bl[73] br[73] wl[212] vdd gnd cell_6t
Xbit_r213_c73 bl[73] br[73] wl[213] vdd gnd cell_6t
Xbit_r214_c73 bl[73] br[73] wl[214] vdd gnd cell_6t
Xbit_r215_c73 bl[73] br[73] wl[215] vdd gnd cell_6t
Xbit_r216_c73 bl[73] br[73] wl[216] vdd gnd cell_6t
Xbit_r217_c73 bl[73] br[73] wl[217] vdd gnd cell_6t
Xbit_r218_c73 bl[73] br[73] wl[218] vdd gnd cell_6t
Xbit_r219_c73 bl[73] br[73] wl[219] vdd gnd cell_6t
Xbit_r220_c73 bl[73] br[73] wl[220] vdd gnd cell_6t
Xbit_r221_c73 bl[73] br[73] wl[221] vdd gnd cell_6t
Xbit_r222_c73 bl[73] br[73] wl[222] vdd gnd cell_6t
Xbit_r223_c73 bl[73] br[73] wl[223] vdd gnd cell_6t
Xbit_r224_c73 bl[73] br[73] wl[224] vdd gnd cell_6t
Xbit_r225_c73 bl[73] br[73] wl[225] vdd gnd cell_6t
Xbit_r226_c73 bl[73] br[73] wl[226] vdd gnd cell_6t
Xbit_r227_c73 bl[73] br[73] wl[227] vdd gnd cell_6t
Xbit_r228_c73 bl[73] br[73] wl[228] vdd gnd cell_6t
Xbit_r229_c73 bl[73] br[73] wl[229] vdd gnd cell_6t
Xbit_r230_c73 bl[73] br[73] wl[230] vdd gnd cell_6t
Xbit_r231_c73 bl[73] br[73] wl[231] vdd gnd cell_6t
Xbit_r232_c73 bl[73] br[73] wl[232] vdd gnd cell_6t
Xbit_r233_c73 bl[73] br[73] wl[233] vdd gnd cell_6t
Xbit_r234_c73 bl[73] br[73] wl[234] vdd gnd cell_6t
Xbit_r235_c73 bl[73] br[73] wl[235] vdd gnd cell_6t
Xbit_r236_c73 bl[73] br[73] wl[236] vdd gnd cell_6t
Xbit_r237_c73 bl[73] br[73] wl[237] vdd gnd cell_6t
Xbit_r238_c73 bl[73] br[73] wl[238] vdd gnd cell_6t
Xbit_r239_c73 bl[73] br[73] wl[239] vdd gnd cell_6t
Xbit_r240_c73 bl[73] br[73] wl[240] vdd gnd cell_6t
Xbit_r241_c73 bl[73] br[73] wl[241] vdd gnd cell_6t
Xbit_r242_c73 bl[73] br[73] wl[242] vdd gnd cell_6t
Xbit_r243_c73 bl[73] br[73] wl[243] vdd gnd cell_6t
Xbit_r244_c73 bl[73] br[73] wl[244] vdd gnd cell_6t
Xbit_r245_c73 bl[73] br[73] wl[245] vdd gnd cell_6t
Xbit_r246_c73 bl[73] br[73] wl[246] vdd gnd cell_6t
Xbit_r247_c73 bl[73] br[73] wl[247] vdd gnd cell_6t
Xbit_r248_c73 bl[73] br[73] wl[248] vdd gnd cell_6t
Xbit_r249_c73 bl[73] br[73] wl[249] vdd gnd cell_6t
Xbit_r250_c73 bl[73] br[73] wl[250] vdd gnd cell_6t
Xbit_r251_c73 bl[73] br[73] wl[251] vdd gnd cell_6t
Xbit_r252_c73 bl[73] br[73] wl[252] vdd gnd cell_6t
Xbit_r253_c73 bl[73] br[73] wl[253] vdd gnd cell_6t
Xbit_r254_c73 bl[73] br[73] wl[254] vdd gnd cell_6t
Xbit_r255_c73 bl[73] br[73] wl[255] vdd gnd cell_6t
Xbit_r0_c74 bl[74] br[74] wl[0] vdd gnd cell_6t
Xbit_r1_c74 bl[74] br[74] wl[1] vdd gnd cell_6t
Xbit_r2_c74 bl[74] br[74] wl[2] vdd gnd cell_6t
Xbit_r3_c74 bl[74] br[74] wl[3] vdd gnd cell_6t
Xbit_r4_c74 bl[74] br[74] wl[4] vdd gnd cell_6t
Xbit_r5_c74 bl[74] br[74] wl[5] vdd gnd cell_6t
Xbit_r6_c74 bl[74] br[74] wl[6] vdd gnd cell_6t
Xbit_r7_c74 bl[74] br[74] wl[7] vdd gnd cell_6t
Xbit_r8_c74 bl[74] br[74] wl[8] vdd gnd cell_6t
Xbit_r9_c74 bl[74] br[74] wl[9] vdd gnd cell_6t
Xbit_r10_c74 bl[74] br[74] wl[10] vdd gnd cell_6t
Xbit_r11_c74 bl[74] br[74] wl[11] vdd gnd cell_6t
Xbit_r12_c74 bl[74] br[74] wl[12] vdd gnd cell_6t
Xbit_r13_c74 bl[74] br[74] wl[13] vdd gnd cell_6t
Xbit_r14_c74 bl[74] br[74] wl[14] vdd gnd cell_6t
Xbit_r15_c74 bl[74] br[74] wl[15] vdd gnd cell_6t
Xbit_r16_c74 bl[74] br[74] wl[16] vdd gnd cell_6t
Xbit_r17_c74 bl[74] br[74] wl[17] vdd gnd cell_6t
Xbit_r18_c74 bl[74] br[74] wl[18] vdd gnd cell_6t
Xbit_r19_c74 bl[74] br[74] wl[19] vdd gnd cell_6t
Xbit_r20_c74 bl[74] br[74] wl[20] vdd gnd cell_6t
Xbit_r21_c74 bl[74] br[74] wl[21] vdd gnd cell_6t
Xbit_r22_c74 bl[74] br[74] wl[22] vdd gnd cell_6t
Xbit_r23_c74 bl[74] br[74] wl[23] vdd gnd cell_6t
Xbit_r24_c74 bl[74] br[74] wl[24] vdd gnd cell_6t
Xbit_r25_c74 bl[74] br[74] wl[25] vdd gnd cell_6t
Xbit_r26_c74 bl[74] br[74] wl[26] vdd gnd cell_6t
Xbit_r27_c74 bl[74] br[74] wl[27] vdd gnd cell_6t
Xbit_r28_c74 bl[74] br[74] wl[28] vdd gnd cell_6t
Xbit_r29_c74 bl[74] br[74] wl[29] vdd gnd cell_6t
Xbit_r30_c74 bl[74] br[74] wl[30] vdd gnd cell_6t
Xbit_r31_c74 bl[74] br[74] wl[31] vdd gnd cell_6t
Xbit_r32_c74 bl[74] br[74] wl[32] vdd gnd cell_6t
Xbit_r33_c74 bl[74] br[74] wl[33] vdd gnd cell_6t
Xbit_r34_c74 bl[74] br[74] wl[34] vdd gnd cell_6t
Xbit_r35_c74 bl[74] br[74] wl[35] vdd gnd cell_6t
Xbit_r36_c74 bl[74] br[74] wl[36] vdd gnd cell_6t
Xbit_r37_c74 bl[74] br[74] wl[37] vdd gnd cell_6t
Xbit_r38_c74 bl[74] br[74] wl[38] vdd gnd cell_6t
Xbit_r39_c74 bl[74] br[74] wl[39] vdd gnd cell_6t
Xbit_r40_c74 bl[74] br[74] wl[40] vdd gnd cell_6t
Xbit_r41_c74 bl[74] br[74] wl[41] vdd gnd cell_6t
Xbit_r42_c74 bl[74] br[74] wl[42] vdd gnd cell_6t
Xbit_r43_c74 bl[74] br[74] wl[43] vdd gnd cell_6t
Xbit_r44_c74 bl[74] br[74] wl[44] vdd gnd cell_6t
Xbit_r45_c74 bl[74] br[74] wl[45] vdd gnd cell_6t
Xbit_r46_c74 bl[74] br[74] wl[46] vdd gnd cell_6t
Xbit_r47_c74 bl[74] br[74] wl[47] vdd gnd cell_6t
Xbit_r48_c74 bl[74] br[74] wl[48] vdd gnd cell_6t
Xbit_r49_c74 bl[74] br[74] wl[49] vdd gnd cell_6t
Xbit_r50_c74 bl[74] br[74] wl[50] vdd gnd cell_6t
Xbit_r51_c74 bl[74] br[74] wl[51] vdd gnd cell_6t
Xbit_r52_c74 bl[74] br[74] wl[52] vdd gnd cell_6t
Xbit_r53_c74 bl[74] br[74] wl[53] vdd gnd cell_6t
Xbit_r54_c74 bl[74] br[74] wl[54] vdd gnd cell_6t
Xbit_r55_c74 bl[74] br[74] wl[55] vdd gnd cell_6t
Xbit_r56_c74 bl[74] br[74] wl[56] vdd gnd cell_6t
Xbit_r57_c74 bl[74] br[74] wl[57] vdd gnd cell_6t
Xbit_r58_c74 bl[74] br[74] wl[58] vdd gnd cell_6t
Xbit_r59_c74 bl[74] br[74] wl[59] vdd gnd cell_6t
Xbit_r60_c74 bl[74] br[74] wl[60] vdd gnd cell_6t
Xbit_r61_c74 bl[74] br[74] wl[61] vdd gnd cell_6t
Xbit_r62_c74 bl[74] br[74] wl[62] vdd gnd cell_6t
Xbit_r63_c74 bl[74] br[74] wl[63] vdd gnd cell_6t
Xbit_r64_c74 bl[74] br[74] wl[64] vdd gnd cell_6t
Xbit_r65_c74 bl[74] br[74] wl[65] vdd gnd cell_6t
Xbit_r66_c74 bl[74] br[74] wl[66] vdd gnd cell_6t
Xbit_r67_c74 bl[74] br[74] wl[67] vdd gnd cell_6t
Xbit_r68_c74 bl[74] br[74] wl[68] vdd gnd cell_6t
Xbit_r69_c74 bl[74] br[74] wl[69] vdd gnd cell_6t
Xbit_r70_c74 bl[74] br[74] wl[70] vdd gnd cell_6t
Xbit_r71_c74 bl[74] br[74] wl[71] vdd gnd cell_6t
Xbit_r72_c74 bl[74] br[74] wl[72] vdd gnd cell_6t
Xbit_r73_c74 bl[74] br[74] wl[73] vdd gnd cell_6t
Xbit_r74_c74 bl[74] br[74] wl[74] vdd gnd cell_6t
Xbit_r75_c74 bl[74] br[74] wl[75] vdd gnd cell_6t
Xbit_r76_c74 bl[74] br[74] wl[76] vdd gnd cell_6t
Xbit_r77_c74 bl[74] br[74] wl[77] vdd gnd cell_6t
Xbit_r78_c74 bl[74] br[74] wl[78] vdd gnd cell_6t
Xbit_r79_c74 bl[74] br[74] wl[79] vdd gnd cell_6t
Xbit_r80_c74 bl[74] br[74] wl[80] vdd gnd cell_6t
Xbit_r81_c74 bl[74] br[74] wl[81] vdd gnd cell_6t
Xbit_r82_c74 bl[74] br[74] wl[82] vdd gnd cell_6t
Xbit_r83_c74 bl[74] br[74] wl[83] vdd gnd cell_6t
Xbit_r84_c74 bl[74] br[74] wl[84] vdd gnd cell_6t
Xbit_r85_c74 bl[74] br[74] wl[85] vdd gnd cell_6t
Xbit_r86_c74 bl[74] br[74] wl[86] vdd gnd cell_6t
Xbit_r87_c74 bl[74] br[74] wl[87] vdd gnd cell_6t
Xbit_r88_c74 bl[74] br[74] wl[88] vdd gnd cell_6t
Xbit_r89_c74 bl[74] br[74] wl[89] vdd gnd cell_6t
Xbit_r90_c74 bl[74] br[74] wl[90] vdd gnd cell_6t
Xbit_r91_c74 bl[74] br[74] wl[91] vdd gnd cell_6t
Xbit_r92_c74 bl[74] br[74] wl[92] vdd gnd cell_6t
Xbit_r93_c74 bl[74] br[74] wl[93] vdd gnd cell_6t
Xbit_r94_c74 bl[74] br[74] wl[94] vdd gnd cell_6t
Xbit_r95_c74 bl[74] br[74] wl[95] vdd gnd cell_6t
Xbit_r96_c74 bl[74] br[74] wl[96] vdd gnd cell_6t
Xbit_r97_c74 bl[74] br[74] wl[97] vdd gnd cell_6t
Xbit_r98_c74 bl[74] br[74] wl[98] vdd gnd cell_6t
Xbit_r99_c74 bl[74] br[74] wl[99] vdd gnd cell_6t
Xbit_r100_c74 bl[74] br[74] wl[100] vdd gnd cell_6t
Xbit_r101_c74 bl[74] br[74] wl[101] vdd gnd cell_6t
Xbit_r102_c74 bl[74] br[74] wl[102] vdd gnd cell_6t
Xbit_r103_c74 bl[74] br[74] wl[103] vdd gnd cell_6t
Xbit_r104_c74 bl[74] br[74] wl[104] vdd gnd cell_6t
Xbit_r105_c74 bl[74] br[74] wl[105] vdd gnd cell_6t
Xbit_r106_c74 bl[74] br[74] wl[106] vdd gnd cell_6t
Xbit_r107_c74 bl[74] br[74] wl[107] vdd gnd cell_6t
Xbit_r108_c74 bl[74] br[74] wl[108] vdd gnd cell_6t
Xbit_r109_c74 bl[74] br[74] wl[109] vdd gnd cell_6t
Xbit_r110_c74 bl[74] br[74] wl[110] vdd gnd cell_6t
Xbit_r111_c74 bl[74] br[74] wl[111] vdd gnd cell_6t
Xbit_r112_c74 bl[74] br[74] wl[112] vdd gnd cell_6t
Xbit_r113_c74 bl[74] br[74] wl[113] vdd gnd cell_6t
Xbit_r114_c74 bl[74] br[74] wl[114] vdd gnd cell_6t
Xbit_r115_c74 bl[74] br[74] wl[115] vdd gnd cell_6t
Xbit_r116_c74 bl[74] br[74] wl[116] vdd gnd cell_6t
Xbit_r117_c74 bl[74] br[74] wl[117] vdd gnd cell_6t
Xbit_r118_c74 bl[74] br[74] wl[118] vdd gnd cell_6t
Xbit_r119_c74 bl[74] br[74] wl[119] vdd gnd cell_6t
Xbit_r120_c74 bl[74] br[74] wl[120] vdd gnd cell_6t
Xbit_r121_c74 bl[74] br[74] wl[121] vdd gnd cell_6t
Xbit_r122_c74 bl[74] br[74] wl[122] vdd gnd cell_6t
Xbit_r123_c74 bl[74] br[74] wl[123] vdd gnd cell_6t
Xbit_r124_c74 bl[74] br[74] wl[124] vdd gnd cell_6t
Xbit_r125_c74 bl[74] br[74] wl[125] vdd gnd cell_6t
Xbit_r126_c74 bl[74] br[74] wl[126] vdd gnd cell_6t
Xbit_r127_c74 bl[74] br[74] wl[127] vdd gnd cell_6t
Xbit_r128_c74 bl[74] br[74] wl[128] vdd gnd cell_6t
Xbit_r129_c74 bl[74] br[74] wl[129] vdd gnd cell_6t
Xbit_r130_c74 bl[74] br[74] wl[130] vdd gnd cell_6t
Xbit_r131_c74 bl[74] br[74] wl[131] vdd gnd cell_6t
Xbit_r132_c74 bl[74] br[74] wl[132] vdd gnd cell_6t
Xbit_r133_c74 bl[74] br[74] wl[133] vdd gnd cell_6t
Xbit_r134_c74 bl[74] br[74] wl[134] vdd gnd cell_6t
Xbit_r135_c74 bl[74] br[74] wl[135] vdd gnd cell_6t
Xbit_r136_c74 bl[74] br[74] wl[136] vdd gnd cell_6t
Xbit_r137_c74 bl[74] br[74] wl[137] vdd gnd cell_6t
Xbit_r138_c74 bl[74] br[74] wl[138] vdd gnd cell_6t
Xbit_r139_c74 bl[74] br[74] wl[139] vdd gnd cell_6t
Xbit_r140_c74 bl[74] br[74] wl[140] vdd gnd cell_6t
Xbit_r141_c74 bl[74] br[74] wl[141] vdd gnd cell_6t
Xbit_r142_c74 bl[74] br[74] wl[142] vdd gnd cell_6t
Xbit_r143_c74 bl[74] br[74] wl[143] vdd gnd cell_6t
Xbit_r144_c74 bl[74] br[74] wl[144] vdd gnd cell_6t
Xbit_r145_c74 bl[74] br[74] wl[145] vdd gnd cell_6t
Xbit_r146_c74 bl[74] br[74] wl[146] vdd gnd cell_6t
Xbit_r147_c74 bl[74] br[74] wl[147] vdd gnd cell_6t
Xbit_r148_c74 bl[74] br[74] wl[148] vdd gnd cell_6t
Xbit_r149_c74 bl[74] br[74] wl[149] vdd gnd cell_6t
Xbit_r150_c74 bl[74] br[74] wl[150] vdd gnd cell_6t
Xbit_r151_c74 bl[74] br[74] wl[151] vdd gnd cell_6t
Xbit_r152_c74 bl[74] br[74] wl[152] vdd gnd cell_6t
Xbit_r153_c74 bl[74] br[74] wl[153] vdd gnd cell_6t
Xbit_r154_c74 bl[74] br[74] wl[154] vdd gnd cell_6t
Xbit_r155_c74 bl[74] br[74] wl[155] vdd gnd cell_6t
Xbit_r156_c74 bl[74] br[74] wl[156] vdd gnd cell_6t
Xbit_r157_c74 bl[74] br[74] wl[157] vdd gnd cell_6t
Xbit_r158_c74 bl[74] br[74] wl[158] vdd gnd cell_6t
Xbit_r159_c74 bl[74] br[74] wl[159] vdd gnd cell_6t
Xbit_r160_c74 bl[74] br[74] wl[160] vdd gnd cell_6t
Xbit_r161_c74 bl[74] br[74] wl[161] vdd gnd cell_6t
Xbit_r162_c74 bl[74] br[74] wl[162] vdd gnd cell_6t
Xbit_r163_c74 bl[74] br[74] wl[163] vdd gnd cell_6t
Xbit_r164_c74 bl[74] br[74] wl[164] vdd gnd cell_6t
Xbit_r165_c74 bl[74] br[74] wl[165] vdd gnd cell_6t
Xbit_r166_c74 bl[74] br[74] wl[166] vdd gnd cell_6t
Xbit_r167_c74 bl[74] br[74] wl[167] vdd gnd cell_6t
Xbit_r168_c74 bl[74] br[74] wl[168] vdd gnd cell_6t
Xbit_r169_c74 bl[74] br[74] wl[169] vdd gnd cell_6t
Xbit_r170_c74 bl[74] br[74] wl[170] vdd gnd cell_6t
Xbit_r171_c74 bl[74] br[74] wl[171] vdd gnd cell_6t
Xbit_r172_c74 bl[74] br[74] wl[172] vdd gnd cell_6t
Xbit_r173_c74 bl[74] br[74] wl[173] vdd gnd cell_6t
Xbit_r174_c74 bl[74] br[74] wl[174] vdd gnd cell_6t
Xbit_r175_c74 bl[74] br[74] wl[175] vdd gnd cell_6t
Xbit_r176_c74 bl[74] br[74] wl[176] vdd gnd cell_6t
Xbit_r177_c74 bl[74] br[74] wl[177] vdd gnd cell_6t
Xbit_r178_c74 bl[74] br[74] wl[178] vdd gnd cell_6t
Xbit_r179_c74 bl[74] br[74] wl[179] vdd gnd cell_6t
Xbit_r180_c74 bl[74] br[74] wl[180] vdd gnd cell_6t
Xbit_r181_c74 bl[74] br[74] wl[181] vdd gnd cell_6t
Xbit_r182_c74 bl[74] br[74] wl[182] vdd gnd cell_6t
Xbit_r183_c74 bl[74] br[74] wl[183] vdd gnd cell_6t
Xbit_r184_c74 bl[74] br[74] wl[184] vdd gnd cell_6t
Xbit_r185_c74 bl[74] br[74] wl[185] vdd gnd cell_6t
Xbit_r186_c74 bl[74] br[74] wl[186] vdd gnd cell_6t
Xbit_r187_c74 bl[74] br[74] wl[187] vdd gnd cell_6t
Xbit_r188_c74 bl[74] br[74] wl[188] vdd gnd cell_6t
Xbit_r189_c74 bl[74] br[74] wl[189] vdd gnd cell_6t
Xbit_r190_c74 bl[74] br[74] wl[190] vdd gnd cell_6t
Xbit_r191_c74 bl[74] br[74] wl[191] vdd gnd cell_6t
Xbit_r192_c74 bl[74] br[74] wl[192] vdd gnd cell_6t
Xbit_r193_c74 bl[74] br[74] wl[193] vdd gnd cell_6t
Xbit_r194_c74 bl[74] br[74] wl[194] vdd gnd cell_6t
Xbit_r195_c74 bl[74] br[74] wl[195] vdd gnd cell_6t
Xbit_r196_c74 bl[74] br[74] wl[196] vdd gnd cell_6t
Xbit_r197_c74 bl[74] br[74] wl[197] vdd gnd cell_6t
Xbit_r198_c74 bl[74] br[74] wl[198] vdd gnd cell_6t
Xbit_r199_c74 bl[74] br[74] wl[199] vdd gnd cell_6t
Xbit_r200_c74 bl[74] br[74] wl[200] vdd gnd cell_6t
Xbit_r201_c74 bl[74] br[74] wl[201] vdd gnd cell_6t
Xbit_r202_c74 bl[74] br[74] wl[202] vdd gnd cell_6t
Xbit_r203_c74 bl[74] br[74] wl[203] vdd gnd cell_6t
Xbit_r204_c74 bl[74] br[74] wl[204] vdd gnd cell_6t
Xbit_r205_c74 bl[74] br[74] wl[205] vdd gnd cell_6t
Xbit_r206_c74 bl[74] br[74] wl[206] vdd gnd cell_6t
Xbit_r207_c74 bl[74] br[74] wl[207] vdd gnd cell_6t
Xbit_r208_c74 bl[74] br[74] wl[208] vdd gnd cell_6t
Xbit_r209_c74 bl[74] br[74] wl[209] vdd gnd cell_6t
Xbit_r210_c74 bl[74] br[74] wl[210] vdd gnd cell_6t
Xbit_r211_c74 bl[74] br[74] wl[211] vdd gnd cell_6t
Xbit_r212_c74 bl[74] br[74] wl[212] vdd gnd cell_6t
Xbit_r213_c74 bl[74] br[74] wl[213] vdd gnd cell_6t
Xbit_r214_c74 bl[74] br[74] wl[214] vdd gnd cell_6t
Xbit_r215_c74 bl[74] br[74] wl[215] vdd gnd cell_6t
Xbit_r216_c74 bl[74] br[74] wl[216] vdd gnd cell_6t
Xbit_r217_c74 bl[74] br[74] wl[217] vdd gnd cell_6t
Xbit_r218_c74 bl[74] br[74] wl[218] vdd gnd cell_6t
Xbit_r219_c74 bl[74] br[74] wl[219] vdd gnd cell_6t
Xbit_r220_c74 bl[74] br[74] wl[220] vdd gnd cell_6t
Xbit_r221_c74 bl[74] br[74] wl[221] vdd gnd cell_6t
Xbit_r222_c74 bl[74] br[74] wl[222] vdd gnd cell_6t
Xbit_r223_c74 bl[74] br[74] wl[223] vdd gnd cell_6t
Xbit_r224_c74 bl[74] br[74] wl[224] vdd gnd cell_6t
Xbit_r225_c74 bl[74] br[74] wl[225] vdd gnd cell_6t
Xbit_r226_c74 bl[74] br[74] wl[226] vdd gnd cell_6t
Xbit_r227_c74 bl[74] br[74] wl[227] vdd gnd cell_6t
Xbit_r228_c74 bl[74] br[74] wl[228] vdd gnd cell_6t
Xbit_r229_c74 bl[74] br[74] wl[229] vdd gnd cell_6t
Xbit_r230_c74 bl[74] br[74] wl[230] vdd gnd cell_6t
Xbit_r231_c74 bl[74] br[74] wl[231] vdd gnd cell_6t
Xbit_r232_c74 bl[74] br[74] wl[232] vdd gnd cell_6t
Xbit_r233_c74 bl[74] br[74] wl[233] vdd gnd cell_6t
Xbit_r234_c74 bl[74] br[74] wl[234] vdd gnd cell_6t
Xbit_r235_c74 bl[74] br[74] wl[235] vdd gnd cell_6t
Xbit_r236_c74 bl[74] br[74] wl[236] vdd gnd cell_6t
Xbit_r237_c74 bl[74] br[74] wl[237] vdd gnd cell_6t
Xbit_r238_c74 bl[74] br[74] wl[238] vdd gnd cell_6t
Xbit_r239_c74 bl[74] br[74] wl[239] vdd gnd cell_6t
Xbit_r240_c74 bl[74] br[74] wl[240] vdd gnd cell_6t
Xbit_r241_c74 bl[74] br[74] wl[241] vdd gnd cell_6t
Xbit_r242_c74 bl[74] br[74] wl[242] vdd gnd cell_6t
Xbit_r243_c74 bl[74] br[74] wl[243] vdd gnd cell_6t
Xbit_r244_c74 bl[74] br[74] wl[244] vdd gnd cell_6t
Xbit_r245_c74 bl[74] br[74] wl[245] vdd gnd cell_6t
Xbit_r246_c74 bl[74] br[74] wl[246] vdd gnd cell_6t
Xbit_r247_c74 bl[74] br[74] wl[247] vdd gnd cell_6t
Xbit_r248_c74 bl[74] br[74] wl[248] vdd gnd cell_6t
Xbit_r249_c74 bl[74] br[74] wl[249] vdd gnd cell_6t
Xbit_r250_c74 bl[74] br[74] wl[250] vdd gnd cell_6t
Xbit_r251_c74 bl[74] br[74] wl[251] vdd gnd cell_6t
Xbit_r252_c74 bl[74] br[74] wl[252] vdd gnd cell_6t
Xbit_r253_c74 bl[74] br[74] wl[253] vdd gnd cell_6t
Xbit_r254_c74 bl[74] br[74] wl[254] vdd gnd cell_6t
Xbit_r255_c74 bl[74] br[74] wl[255] vdd gnd cell_6t
Xbit_r0_c75 bl[75] br[75] wl[0] vdd gnd cell_6t
Xbit_r1_c75 bl[75] br[75] wl[1] vdd gnd cell_6t
Xbit_r2_c75 bl[75] br[75] wl[2] vdd gnd cell_6t
Xbit_r3_c75 bl[75] br[75] wl[3] vdd gnd cell_6t
Xbit_r4_c75 bl[75] br[75] wl[4] vdd gnd cell_6t
Xbit_r5_c75 bl[75] br[75] wl[5] vdd gnd cell_6t
Xbit_r6_c75 bl[75] br[75] wl[6] vdd gnd cell_6t
Xbit_r7_c75 bl[75] br[75] wl[7] vdd gnd cell_6t
Xbit_r8_c75 bl[75] br[75] wl[8] vdd gnd cell_6t
Xbit_r9_c75 bl[75] br[75] wl[9] vdd gnd cell_6t
Xbit_r10_c75 bl[75] br[75] wl[10] vdd gnd cell_6t
Xbit_r11_c75 bl[75] br[75] wl[11] vdd gnd cell_6t
Xbit_r12_c75 bl[75] br[75] wl[12] vdd gnd cell_6t
Xbit_r13_c75 bl[75] br[75] wl[13] vdd gnd cell_6t
Xbit_r14_c75 bl[75] br[75] wl[14] vdd gnd cell_6t
Xbit_r15_c75 bl[75] br[75] wl[15] vdd gnd cell_6t
Xbit_r16_c75 bl[75] br[75] wl[16] vdd gnd cell_6t
Xbit_r17_c75 bl[75] br[75] wl[17] vdd gnd cell_6t
Xbit_r18_c75 bl[75] br[75] wl[18] vdd gnd cell_6t
Xbit_r19_c75 bl[75] br[75] wl[19] vdd gnd cell_6t
Xbit_r20_c75 bl[75] br[75] wl[20] vdd gnd cell_6t
Xbit_r21_c75 bl[75] br[75] wl[21] vdd gnd cell_6t
Xbit_r22_c75 bl[75] br[75] wl[22] vdd gnd cell_6t
Xbit_r23_c75 bl[75] br[75] wl[23] vdd gnd cell_6t
Xbit_r24_c75 bl[75] br[75] wl[24] vdd gnd cell_6t
Xbit_r25_c75 bl[75] br[75] wl[25] vdd gnd cell_6t
Xbit_r26_c75 bl[75] br[75] wl[26] vdd gnd cell_6t
Xbit_r27_c75 bl[75] br[75] wl[27] vdd gnd cell_6t
Xbit_r28_c75 bl[75] br[75] wl[28] vdd gnd cell_6t
Xbit_r29_c75 bl[75] br[75] wl[29] vdd gnd cell_6t
Xbit_r30_c75 bl[75] br[75] wl[30] vdd gnd cell_6t
Xbit_r31_c75 bl[75] br[75] wl[31] vdd gnd cell_6t
Xbit_r32_c75 bl[75] br[75] wl[32] vdd gnd cell_6t
Xbit_r33_c75 bl[75] br[75] wl[33] vdd gnd cell_6t
Xbit_r34_c75 bl[75] br[75] wl[34] vdd gnd cell_6t
Xbit_r35_c75 bl[75] br[75] wl[35] vdd gnd cell_6t
Xbit_r36_c75 bl[75] br[75] wl[36] vdd gnd cell_6t
Xbit_r37_c75 bl[75] br[75] wl[37] vdd gnd cell_6t
Xbit_r38_c75 bl[75] br[75] wl[38] vdd gnd cell_6t
Xbit_r39_c75 bl[75] br[75] wl[39] vdd gnd cell_6t
Xbit_r40_c75 bl[75] br[75] wl[40] vdd gnd cell_6t
Xbit_r41_c75 bl[75] br[75] wl[41] vdd gnd cell_6t
Xbit_r42_c75 bl[75] br[75] wl[42] vdd gnd cell_6t
Xbit_r43_c75 bl[75] br[75] wl[43] vdd gnd cell_6t
Xbit_r44_c75 bl[75] br[75] wl[44] vdd gnd cell_6t
Xbit_r45_c75 bl[75] br[75] wl[45] vdd gnd cell_6t
Xbit_r46_c75 bl[75] br[75] wl[46] vdd gnd cell_6t
Xbit_r47_c75 bl[75] br[75] wl[47] vdd gnd cell_6t
Xbit_r48_c75 bl[75] br[75] wl[48] vdd gnd cell_6t
Xbit_r49_c75 bl[75] br[75] wl[49] vdd gnd cell_6t
Xbit_r50_c75 bl[75] br[75] wl[50] vdd gnd cell_6t
Xbit_r51_c75 bl[75] br[75] wl[51] vdd gnd cell_6t
Xbit_r52_c75 bl[75] br[75] wl[52] vdd gnd cell_6t
Xbit_r53_c75 bl[75] br[75] wl[53] vdd gnd cell_6t
Xbit_r54_c75 bl[75] br[75] wl[54] vdd gnd cell_6t
Xbit_r55_c75 bl[75] br[75] wl[55] vdd gnd cell_6t
Xbit_r56_c75 bl[75] br[75] wl[56] vdd gnd cell_6t
Xbit_r57_c75 bl[75] br[75] wl[57] vdd gnd cell_6t
Xbit_r58_c75 bl[75] br[75] wl[58] vdd gnd cell_6t
Xbit_r59_c75 bl[75] br[75] wl[59] vdd gnd cell_6t
Xbit_r60_c75 bl[75] br[75] wl[60] vdd gnd cell_6t
Xbit_r61_c75 bl[75] br[75] wl[61] vdd gnd cell_6t
Xbit_r62_c75 bl[75] br[75] wl[62] vdd gnd cell_6t
Xbit_r63_c75 bl[75] br[75] wl[63] vdd gnd cell_6t
Xbit_r64_c75 bl[75] br[75] wl[64] vdd gnd cell_6t
Xbit_r65_c75 bl[75] br[75] wl[65] vdd gnd cell_6t
Xbit_r66_c75 bl[75] br[75] wl[66] vdd gnd cell_6t
Xbit_r67_c75 bl[75] br[75] wl[67] vdd gnd cell_6t
Xbit_r68_c75 bl[75] br[75] wl[68] vdd gnd cell_6t
Xbit_r69_c75 bl[75] br[75] wl[69] vdd gnd cell_6t
Xbit_r70_c75 bl[75] br[75] wl[70] vdd gnd cell_6t
Xbit_r71_c75 bl[75] br[75] wl[71] vdd gnd cell_6t
Xbit_r72_c75 bl[75] br[75] wl[72] vdd gnd cell_6t
Xbit_r73_c75 bl[75] br[75] wl[73] vdd gnd cell_6t
Xbit_r74_c75 bl[75] br[75] wl[74] vdd gnd cell_6t
Xbit_r75_c75 bl[75] br[75] wl[75] vdd gnd cell_6t
Xbit_r76_c75 bl[75] br[75] wl[76] vdd gnd cell_6t
Xbit_r77_c75 bl[75] br[75] wl[77] vdd gnd cell_6t
Xbit_r78_c75 bl[75] br[75] wl[78] vdd gnd cell_6t
Xbit_r79_c75 bl[75] br[75] wl[79] vdd gnd cell_6t
Xbit_r80_c75 bl[75] br[75] wl[80] vdd gnd cell_6t
Xbit_r81_c75 bl[75] br[75] wl[81] vdd gnd cell_6t
Xbit_r82_c75 bl[75] br[75] wl[82] vdd gnd cell_6t
Xbit_r83_c75 bl[75] br[75] wl[83] vdd gnd cell_6t
Xbit_r84_c75 bl[75] br[75] wl[84] vdd gnd cell_6t
Xbit_r85_c75 bl[75] br[75] wl[85] vdd gnd cell_6t
Xbit_r86_c75 bl[75] br[75] wl[86] vdd gnd cell_6t
Xbit_r87_c75 bl[75] br[75] wl[87] vdd gnd cell_6t
Xbit_r88_c75 bl[75] br[75] wl[88] vdd gnd cell_6t
Xbit_r89_c75 bl[75] br[75] wl[89] vdd gnd cell_6t
Xbit_r90_c75 bl[75] br[75] wl[90] vdd gnd cell_6t
Xbit_r91_c75 bl[75] br[75] wl[91] vdd gnd cell_6t
Xbit_r92_c75 bl[75] br[75] wl[92] vdd gnd cell_6t
Xbit_r93_c75 bl[75] br[75] wl[93] vdd gnd cell_6t
Xbit_r94_c75 bl[75] br[75] wl[94] vdd gnd cell_6t
Xbit_r95_c75 bl[75] br[75] wl[95] vdd gnd cell_6t
Xbit_r96_c75 bl[75] br[75] wl[96] vdd gnd cell_6t
Xbit_r97_c75 bl[75] br[75] wl[97] vdd gnd cell_6t
Xbit_r98_c75 bl[75] br[75] wl[98] vdd gnd cell_6t
Xbit_r99_c75 bl[75] br[75] wl[99] vdd gnd cell_6t
Xbit_r100_c75 bl[75] br[75] wl[100] vdd gnd cell_6t
Xbit_r101_c75 bl[75] br[75] wl[101] vdd gnd cell_6t
Xbit_r102_c75 bl[75] br[75] wl[102] vdd gnd cell_6t
Xbit_r103_c75 bl[75] br[75] wl[103] vdd gnd cell_6t
Xbit_r104_c75 bl[75] br[75] wl[104] vdd gnd cell_6t
Xbit_r105_c75 bl[75] br[75] wl[105] vdd gnd cell_6t
Xbit_r106_c75 bl[75] br[75] wl[106] vdd gnd cell_6t
Xbit_r107_c75 bl[75] br[75] wl[107] vdd gnd cell_6t
Xbit_r108_c75 bl[75] br[75] wl[108] vdd gnd cell_6t
Xbit_r109_c75 bl[75] br[75] wl[109] vdd gnd cell_6t
Xbit_r110_c75 bl[75] br[75] wl[110] vdd gnd cell_6t
Xbit_r111_c75 bl[75] br[75] wl[111] vdd gnd cell_6t
Xbit_r112_c75 bl[75] br[75] wl[112] vdd gnd cell_6t
Xbit_r113_c75 bl[75] br[75] wl[113] vdd gnd cell_6t
Xbit_r114_c75 bl[75] br[75] wl[114] vdd gnd cell_6t
Xbit_r115_c75 bl[75] br[75] wl[115] vdd gnd cell_6t
Xbit_r116_c75 bl[75] br[75] wl[116] vdd gnd cell_6t
Xbit_r117_c75 bl[75] br[75] wl[117] vdd gnd cell_6t
Xbit_r118_c75 bl[75] br[75] wl[118] vdd gnd cell_6t
Xbit_r119_c75 bl[75] br[75] wl[119] vdd gnd cell_6t
Xbit_r120_c75 bl[75] br[75] wl[120] vdd gnd cell_6t
Xbit_r121_c75 bl[75] br[75] wl[121] vdd gnd cell_6t
Xbit_r122_c75 bl[75] br[75] wl[122] vdd gnd cell_6t
Xbit_r123_c75 bl[75] br[75] wl[123] vdd gnd cell_6t
Xbit_r124_c75 bl[75] br[75] wl[124] vdd gnd cell_6t
Xbit_r125_c75 bl[75] br[75] wl[125] vdd gnd cell_6t
Xbit_r126_c75 bl[75] br[75] wl[126] vdd gnd cell_6t
Xbit_r127_c75 bl[75] br[75] wl[127] vdd gnd cell_6t
Xbit_r128_c75 bl[75] br[75] wl[128] vdd gnd cell_6t
Xbit_r129_c75 bl[75] br[75] wl[129] vdd gnd cell_6t
Xbit_r130_c75 bl[75] br[75] wl[130] vdd gnd cell_6t
Xbit_r131_c75 bl[75] br[75] wl[131] vdd gnd cell_6t
Xbit_r132_c75 bl[75] br[75] wl[132] vdd gnd cell_6t
Xbit_r133_c75 bl[75] br[75] wl[133] vdd gnd cell_6t
Xbit_r134_c75 bl[75] br[75] wl[134] vdd gnd cell_6t
Xbit_r135_c75 bl[75] br[75] wl[135] vdd gnd cell_6t
Xbit_r136_c75 bl[75] br[75] wl[136] vdd gnd cell_6t
Xbit_r137_c75 bl[75] br[75] wl[137] vdd gnd cell_6t
Xbit_r138_c75 bl[75] br[75] wl[138] vdd gnd cell_6t
Xbit_r139_c75 bl[75] br[75] wl[139] vdd gnd cell_6t
Xbit_r140_c75 bl[75] br[75] wl[140] vdd gnd cell_6t
Xbit_r141_c75 bl[75] br[75] wl[141] vdd gnd cell_6t
Xbit_r142_c75 bl[75] br[75] wl[142] vdd gnd cell_6t
Xbit_r143_c75 bl[75] br[75] wl[143] vdd gnd cell_6t
Xbit_r144_c75 bl[75] br[75] wl[144] vdd gnd cell_6t
Xbit_r145_c75 bl[75] br[75] wl[145] vdd gnd cell_6t
Xbit_r146_c75 bl[75] br[75] wl[146] vdd gnd cell_6t
Xbit_r147_c75 bl[75] br[75] wl[147] vdd gnd cell_6t
Xbit_r148_c75 bl[75] br[75] wl[148] vdd gnd cell_6t
Xbit_r149_c75 bl[75] br[75] wl[149] vdd gnd cell_6t
Xbit_r150_c75 bl[75] br[75] wl[150] vdd gnd cell_6t
Xbit_r151_c75 bl[75] br[75] wl[151] vdd gnd cell_6t
Xbit_r152_c75 bl[75] br[75] wl[152] vdd gnd cell_6t
Xbit_r153_c75 bl[75] br[75] wl[153] vdd gnd cell_6t
Xbit_r154_c75 bl[75] br[75] wl[154] vdd gnd cell_6t
Xbit_r155_c75 bl[75] br[75] wl[155] vdd gnd cell_6t
Xbit_r156_c75 bl[75] br[75] wl[156] vdd gnd cell_6t
Xbit_r157_c75 bl[75] br[75] wl[157] vdd gnd cell_6t
Xbit_r158_c75 bl[75] br[75] wl[158] vdd gnd cell_6t
Xbit_r159_c75 bl[75] br[75] wl[159] vdd gnd cell_6t
Xbit_r160_c75 bl[75] br[75] wl[160] vdd gnd cell_6t
Xbit_r161_c75 bl[75] br[75] wl[161] vdd gnd cell_6t
Xbit_r162_c75 bl[75] br[75] wl[162] vdd gnd cell_6t
Xbit_r163_c75 bl[75] br[75] wl[163] vdd gnd cell_6t
Xbit_r164_c75 bl[75] br[75] wl[164] vdd gnd cell_6t
Xbit_r165_c75 bl[75] br[75] wl[165] vdd gnd cell_6t
Xbit_r166_c75 bl[75] br[75] wl[166] vdd gnd cell_6t
Xbit_r167_c75 bl[75] br[75] wl[167] vdd gnd cell_6t
Xbit_r168_c75 bl[75] br[75] wl[168] vdd gnd cell_6t
Xbit_r169_c75 bl[75] br[75] wl[169] vdd gnd cell_6t
Xbit_r170_c75 bl[75] br[75] wl[170] vdd gnd cell_6t
Xbit_r171_c75 bl[75] br[75] wl[171] vdd gnd cell_6t
Xbit_r172_c75 bl[75] br[75] wl[172] vdd gnd cell_6t
Xbit_r173_c75 bl[75] br[75] wl[173] vdd gnd cell_6t
Xbit_r174_c75 bl[75] br[75] wl[174] vdd gnd cell_6t
Xbit_r175_c75 bl[75] br[75] wl[175] vdd gnd cell_6t
Xbit_r176_c75 bl[75] br[75] wl[176] vdd gnd cell_6t
Xbit_r177_c75 bl[75] br[75] wl[177] vdd gnd cell_6t
Xbit_r178_c75 bl[75] br[75] wl[178] vdd gnd cell_6t
Xbit_r179_c75 bl[75] br[75] wl[179] vdd gnd cell_6t
Xbit_r180_c75 bl[75] br[75] wl[180] vdd gnd cell_6t
Xbit_r181_c75 bl[75] br[75] wl[181] vdd gnd cell_6t
Xbit_r182_c75 bl[75] br[75] wl[182] vdd gnd cell_6t
Xbit_r183_c75 bl[75] br[75] wl[183] vdd gnd cell_6t
Xbit_r184_c75 bl[75] br[75] wl[184] vdd gnd cell_6t
Xbit_r185_c75 bl[75] br[75] wl[185] vdd gnd cell_6t
Xbit_r186_c75 bl[75] br[75] wl[186] vdd gnd cell_6t
Xbit_r187_c75 bl[75] br[75] wl[187] vdd gnd cell_6t
Xbit_r188_c75 bl[75] br[75] wl[188] vdd gnd cell_6t
Xbit_r189_c75 bl[75] br[75] wl[189] vdd gnd cell_6t
Xbit_r190_c75 bl[75] br[75] wl[190] vdd gnd cell_6t
Xbit_r191_c75 bl[75] br[75] wl[191] vdd gnd cell_6t
Xbit_r192_c75 bl[75] br[75] wl[192] vdd gnd cell_6t
Xbit_r193_c75 bl[75] br[75] wl[193] vdd gnd cell_6t
Xbit_r194_c75 bl[75] br[75] wl[194] vdd gnd cell_6t
Xbit_r195_c75 bl[75] br[75] wl[195] vdd gnd cell_6t
Xbit_r196_c75 bl[75] br[75] wl[196] vdd gnd cell_6t
Xbit_r197_c75 bl[75] br[75] wl[197] vdd gnd cell_6t
Xbit_r198_c75 bl[75] br[75] wl[198] vdd gnd cell_6t
Xbit_r199_c75 bl[75] br[75] wl[199] vdd gnd cell_6t
Xbit_r200_c75 bl[75] br[75] wl[200] vdd gnd cell_6t
Xbit_r201_c75 bl[75] br[75] wl[201] vdd gnd cell_6t
Xbit_r202_c75 bl[75] br[75] wl[202] vdd gnd cell_6t
Xbit_r203_c75 bl[75] br[75] wl[203] vdd gnd cell_6t
Xbit_r204_c75 bl[75] br[75] wl[204] vdd gnd cell_6t
Xbit_r205_c75 bl[75] br[75] wl[205] vdd gnd cell_6t
Xbit_r206_c75 bl[75] br[75] wl[206] vdd gnd cell_6t
Xbit_r207_c75 bl[75] br[75] wl[207] vdd gnd cell_6t
Xbit_r208_c75 bl[75] br[75] wl[208] vdd gnd cell_6t
Xbit_r209_c75 bl[75] br[75] wl[209] vdd gnd cell_6t
Xbit_r210_c75 bl[75] br[75] wl[210] vdd gnd cell_6t
Xbit_r211_c75 bl[75] br[75] wl[211] vdd gnd cell_6t
Xbit_r212_c75 bl[75] br[75] wl[212] vdd gnd cell_6t
Xbit_r213_c75 bl[75] br[75] wl[213] vdd gnd cell_6t
Xbit_r214_c75 bl[75] br[75] wl[214] vdd gnd cell_6t
Xbit_r215_c75 bl[75] br[75] wl[215] vdd gnd cell_6t
Xbit_r216_c75 bl[75] br[75] wl[216] vdd gnd cell_6t
Xbit_r217_c75 bl[75] br[75] wl[217] vdd gnd cell_6t
Xbit_r218_c75 bl[75] br[75] wl[218] vdd gnd cell_6t
Xbit_r219_c75 bl[75] br[75] wl[219] vdd gnd cell_6t
Xbit_r220_c75 bl[75] br[75] wl[220] vdd gnd cell_6t
Xbit_r221_c75 bl[75] br[75] wl[221] vdd gnd cell_6t
Xbit_r222_c75 bl[75] br[75] wl[222] vdd gnd cell_6t
Xbit_r223_c75 bl[75] br[75] wl[223] vdd gnd cell_6t
Xbit_r224_c75 bl[75] br[75] wl[224] vdd gnd cell_6t
Xbit_r225_c75 bl[75] br[75] wl[225] vdd gnd cell_6t
Xbit_r226_c75 bl[75] br[75] wl[226] vdd gnd cell_6t
Xbit_r227_c75 bl[75] br[75] wl[227] vdd gnd cell_6t
Xbit_r228_c75 bl[75] br[75] wl[228] vdd gnd cell_6t
Xbit_r229_c75 bl[75] br[75] wl[229] vdd gnd cell_6t
Xbit_r230_c75 bl[75] br[75] wl[230] vdd gnd cell_6t
Xbit_r231_c75 bl[75] br[75] wl[231] vdd gnd cell_6t
Xbit_r232_c75 bl[75] br[75] wl[232] vdd gnd cell_6t
Xbit_r233_c75 bl[75] br[75] wl[233] vdd gnd cell_6t
Xbit_r234_c75 bl[75] br[75] wl[234] vdd gnd cell_6t
Xbit_r235_c75 bl[75] br[75] wl[235] vdd gnd cell_6t
Xbit_r236_c75 bl[75] br[75] wl[236] vdd gnd cell_6t
Xbit_r237_c75 bl[75] br[75] wl[237] vdd gnd cell_6t
Xbit_r238_c75 bl[75] br[75] wl[238] vdd gnd cell_6t
Xbit_r239_c75 bl[75] br[75] wl[239] vdd gnd cell_6t
Xbit_r240_c75 bl[75] br[75] wl[240] vdd gnd cell_6t
Xbit_r241_c75 bl[75] br[75] wl[241] vdd gnd cell_6t
Xbit_r242_c75 bl[75] br[75] wl[242] vdd gnd cell_6t
Xbit_r243_c75 bl[75] br[75] wl[243] vdd gnd cell_6t
Xbit_r244_c75 bl[75] br[75] wl[244] vdd gnd cell_6t
Xbit_r245_c75 bl[75] br[75] wl[245] vdd gnd cell_6t
Xbit_r246_c75 bl[75] br[75] wl[246] vdd gnd cell_6t
Xbit_r247_c75 bl[75] br[75] wl[247] vdd gnd cell_6t
Xbit_r248_c75 bl[75] br[75] wl[248] vdd gnd cell_6t
Xbit_r249_c75 bl[75] br[75] wl[249] vdd gnd cell_6t
Xbit_r250_c75 bl[75] br[75] wl[250] vdd gnd cell_6t
Xbit_r251_c75 bl[75] br[75] wl[251] vdd gnd cell_6t
Xbit_r252_c75 bl[75] br[75] wl[252] vdd gnd cell_6t
Xbit_r253_c75 bl[75] br[75] wl[253] vdd gnd cell_6t
Xbit_r254_c75 bl[75] br[75] wl[254] vdd gnd cell_6t
Xbit_r255_c75 bl[75] br[75] wl[255] vdd gnd cell_6t
Xbit_r0_c76 bl[76] br[76] wl[0] vdd gnd cell_6t
Xbit_r1_c76 bl[76] br[76] wl[1] vdd gnd cell_6t
Xbit_r2_c76 bl[76] br[76] wl[2] vdd gnd cell_6t
Xbit_r3_c76 bl[76] br[76] wl[3] vdd gnd cell_6t
Xbit_r4_c76 bl[76] br[76] wl[4] vdd gnd cell_6t
Xbit_r5_c76 bl[76] br[76] wl[5] vdd gnd cell_6t
Xbit_r6_c76 bl[76] br[76] wl[6] vdd gnd cell_6t
Xbit_r7_c76 bl[76] br[76] wl[7] vdd gnd cell_6t
Xbit_r8_c76 bl[76] br[76] wl[8] vdd gnd cell_6t
Xbit_r9_c76 bl[76] br[76] wl[9] vdd gnd cell_6t
Xbit_r10_c76 bl[76] br[76] wl[10] vdd gnd cell_6t
Xbit_r11_c76 bl[76] br[76] wl[11] vdd gnd cell_6t
Xbit_r12_c76 bl[76] br[76] wl[12] vdd gnd cell_6t
Xbit_r13_c76 bl[76] br[76] wl[13] vdd gnd cell_6t
Xbit_r14_c76 bl[76] br[76] wl[14] vdd gnd cell_6t
Xbit_r15_c76 bl[76] br[76] wl[15] vdd gnd cell_6t
Xbit_r16_c76 bl[76] br[76] wl[16] vdd gnd cell_6t
Xbit_r17_c76 bl[76] br[76] wl[17] vdd gnd cell_6t
Xbit_r18_c76 bl[76] br[76] wl[18] vdd gnd cell_6t
Xbit_r19_c76 bl[76] br[76] wl[19] vdd gnd cell_6t
Xbit_r20_c76 bl[76] br[76] wl[20] vdd gnd cell_6t
Xbit_r21_c76 bl[76] br[76] wl[21] vdd gnd cell_6t
Xbit_r22_c76 bl[76] br[76] wl[22] vdd gnd cell_6t
Xbit_r23_c76 bl[76] br[76] wl[23] vdd gnd cell_6t
Xbit_r24_c76 bl[76] br[76] wl[24] vdd gnd cell_6t
Xbit_r25_c76 bl[76] br[76] wl[25] vdd gnd cell_6t
Xbit_r26_c76 bl[76] br[76] wl[26] vdd gnd cell_6t
Xbit_r27_c76 bl[76] br[76] wl[27] vdd gnd cell_6t
Xbit_r28_c76 bl[76] br[76] wl[28] vdd gnd cell_6t
Xbit_r29_c76 bl[76] br[76] wl[29] vdd gnd cell_6t
Xbit_r30_c76 bl[76] br[76] wl[30] vdd gnd cell_6t
Xbit_r31_c76 bl[76] br[76] wl[31] vdd gnd cell_6t
Xbit_r32_c76 bl[76] br[76] wl[32] vdd gnd cell_6t
Xbit_r33_c76 bl[76] br[76] wl[33] vdd gnd cell_6t
Xbit_r34_c76 bl[76] br[76] wl[34] vdd gnd cell_6t
Xbit_r35_c76 bl[76] br[76] wl[35] vdd gnd cell_6t
Xbit_r36_c76 bl[76] br[76] wl[36] vdd gnd cell_6t
Xbit_r37_c76 bl[76] br[76] wl[37] vdd gnd cell_6t
Xbit_r38_c76 bl[76] br[76] wl[38] vdd gnd cell_6t
Xbit_r39_c76 bl[76] br[76] wl[39] vdd gnd cell_6t
Xbit_r40_c76 bl[76] br[76] wl[40] vdd gnd cell_6t
Xbit_r41_c76 bl[76] br[76] wl[41] vdd gnd cell_6t
Xbit_r42_c76 bl[76] br[76] wl[42] vdd gnd cell_6t
Xbit_r43_c76 bl[76] br[76] wl[43] vdd gnd cell_6t
Xbit_r44_c76 bl[76] br[76] wl[44] vdd gnd cell_6t
Xbit_r45_c76 bl[76] br[76] wl[45] vdd gnd cell_6t
Xbit_r46_c76 bl[76] br[76] wl[46] vdd gnd cell_6t
Xbit_r47_c76 bl[76] br[76] wl[47] vdd gnd cell_6t
Xbit_r48_c76 bl[76] br[76] wl[48] vdd gnd cell_6t
Xbit_r49_c76 bl[76] br[76] wl[49] vdd gnd cell_6t
Xbit_r50_c76 bl[76] br[76] wl[50] vdd gnd cell_6t
Xbit_r51_c76 bl[76] br[76] wl[51] vdd gnd cell_6t
Xbit_r52_c76 bl[76] br[76] wl[52] vdd gnd cell_6t
Xbit_r53_c76 bl[76] br[76] wl[53] vdd gnd cell_6t
Xbit_r54_c76 bl[76] br[76] wl[54] vdd gnd cell_6t
Xbit_r55_c76 bl[76] br[76] wl[55] vdd gnd cell_6t
Xbit_r56_c76 bl[76] br[76] wl[56] vdd gnd cell_6t
Xbit_r57_c76 bl[76] br[76] wl[57] vdd gnd cell_6t
Xbit_r58_c76 bl[76] br[76] wl[58] vdd gnd cell_6t
Xbit_r59_c76 bl[76] br[76] wl[59] vdd gnd cell_6t
Xbit_r60_c76 bl[76] br[76] wl[60] vdd gnd cell_6t
Xbit_r61_c76 bl[76] br[76] wl[61] vdd gnd cell_6t
Xbit_r62_c76 bl[76] br[76] wl[62] vdd gnd cell_6t
Xbit_r63_c76 bl[76] br[76] wl[63] vdd gnd cell_6t
Xbit_r64_c76 bl[76] br[76] wl[64] vdd gnd cell_6t
Xbit_r65_c76 bl[76] br[76] wl[65] vdd gnd cell_6t
Xbit_r66_c76 bl[76] br[76] wl[66] vdd gnd cell_6t
Xbit_r67_c76 bl[76] br[76] wl[67] vdd gnd cell_6t
Xbit_r68_c76 bl[76] br[76] wl[68] vdd gnd cell_6t
Xbit_r69_c76 bl[76] br[76] wl[69] vdd gnd cell_6t
Xbit_r70_c76 bl[76] br[76] wl[70] vdd gnd cell_6t
Xbit_r71_c76 bl[76] br[76] wl[71] vdd gnd cell_6t
Xbit_r72_c76 bl[76] br[76] wl[72] vdd gnd cell_6t
Xbit_r73_c76 bl[76] br[76] wl[73] vdd gnd cell_6t
Xbit_r74_c76 bl[76] br[76] wl[74] vdd gnd cell_6t
Xbit_r75_c76 bl[76] br[76] wl[75] vdd gnd cell_6t
Xbit_r76_c76 bl[76] br[76] wl[76] vdd gnd cell_6t
Xbit_r77_c76 bl[76] br[76] wl[77] vdd gnd cell_6t
Xbit_r78_c76 bl[76] br[76] wl[78] vdd gnd cell_6t
Xbit_r79_c76 bl[76] br[76] wl[79] vdd gnd cell_6t
Xbit_r80_c76 bl[76] br[76] wl[80] vdd gnd cell_6t
Xbit_r81_c76 bl[76] br[76] wl[81] vdd gnd cell_6t
Xbit_r82_c76 bl[76] br[76] wl[82] vdd gnd cell_6t
Xbit_r83_c76 bl[76] br[76] wl[83] vdd gnd cell_6t
Xbit_r84_c76 bl[76] br[76] wl[84] vdd gnd cell_6t
Xbit_r85_c76 bl[76] br[76] wl[85] vdd gnd cell_6t
Xbit_r86_c76 bl[76] br[76] wl[86] vdd gnd cell_6t
Xbit_r87_c76 bl[76] br[76] wl[87] vdd gnd cell_6t
Xbit_r88_c76 bl[76] br[76] wl[88] vdd gnd cell_6t
Xbit_r89_c76 bl[76] br[76] wl[89] vdd gnd cell_6t
Xbit_r90_c76 bl[76] br[76] wl[90] vdd gnd cell_6t
Xbit_r91_c76 bl[76] br[76] wl[91] vdd gnd cell_6t
Xbit_r92_c76 bl[76] br[76] wl[92] vdd gnd cell_6t
Xbit_r93_c76 bl[76] br[76] wl[93] vdd gnd cell_6t
Xbit_r94_c76 bl[76] br[76] wl[94] vdd gnd cell_6t
Xbit_r95_c76 bl[76] br[76] wl[95] vdd gnd cell_6t
Xbit_r96_c76 bl[76] br[76] wl[96] vdd gnd cell_6t
Xbit_r97_c76 bl[76] br[76] wl[97] vdd gnd cell_6t
Xbit_r98_c76 bl[76] br[76] wl[98] vdd gnd cell_6t
Xbit_r99_c76 bl[76] br[76] wl[99] vdd gnd cell_6t
Xbit_r100_c76 bl[76] br[76] wl[100] vdd gnd cell_6t
Xbit_r101_c76 bl[76] br[76] wl[101] vdd gnd cell_6t
Xbit_r102_c76 bl[76] br[76] wl[102] vdd gnd cell_6t
Xbit_r103_c76 bl[76] br[76] wl[103] vdd gnd cell_6t
Xbit_r104_c76 bl[76] br[76] wl[104] vdd gnd cell_6t
Xbit_r105_c76 bl[76] br[76] wl[105] vdd gnd cell_6t
Xbit_r106_c76 bl[76] br[76] wl[106] vdd gnd cell_6t
Xbit_r107_c76 bl[76] br[76] wl[107] vdd gnd cell_6t
Xbit_r108_c76 bl[76] br[76] wl[108] vdd gnd cell_6t
Xbit_r109_c76 bl[76] br[76] wl[109] vdd gnd cell_6t
Xbit_r110_c76 bl[76] br[76] wl[110] vdd gnd cell_6t
Xbit_r111_c76 bl[76] br[76] wl[111] vdd gnd cell_6t
Xbit_r112_c76 bl[76] br[76] wl[112] vdd gnd cell_6t
Xbit_r113_c76 bl[76] br[76] wl[113] vdd gnd cell_6t
Xbit_r114_c76 bl[76] br[76] wl[114] vdd gnd cell_6t
Xbit_r115_c76 bl[76] br[76] wl[115] vdd gnd cell_6t
Xbit_r116_c76 bl[76] br[76] wl[116] vdd gnd cell_6t
Xbit_r117_c76 bl[76] br[76] wl[117] vdd gnd cell_6t
Xbit_r118_c76 bl[76] br[76] wl[118] vdd gnd cell_6t
Xbit_r119_c76 bl[76] br[76] wl[119] vdd gnd cell_6t
Xbit_r120_c76 bl[76] br[76] wl[120] vdd gnd cell_6t
Xbit_r121_c76 bl[76] br[76] wl[121] vdd gnd cell_6t
Xbit_r122_c76 bl[76] br[76] wl[122] vdd gnd cell_6t
Xbit_r123_c76 bl[76] br[76] wl[123] vdd gnd cell_6t
Xbit_r124_c76 bl[76] br[76] wl[124] vdd gnd cell_6t
Xbit_r125_c76 bl[76] br[76] wl[125] vdd gnd cell_6t
Xbit_r126_c76 bl[76] br[76] wl[126] vdd gnd cell_6t
Xbit_r127_c76 bl[76] br[76] wl[127] vdd gnd cell_6t
Xbit_r128_c76 bl[76] br[76] wl[128] vdd gnd cell_6t
Xbit_r129_c76 bl[76] br[76] wl[129] vdd gnd cell_6t
Xbit_r130_c76 bl[76] br[76] wl[130] vdd gnd cell_6t
Xbit_r131_c76 bl[76] br[76] wl[131] vdd gnd cell_6t
Xbit_r132_c76 bl[76] br[76] wl[132] vdd gnd cell_6t
Xbit_r133_c76 bl[76] br[76] wl[133] vdd gnd cell_6t
Xbit_r134_c76 bl[76] br[76] wl[134] vdd gnd cell_6t
Xbit_r135_c76 bl[76] br[76] wl[135] vdd gnd cell_6t
Xbit_r136_c76 bl[76] br[76] wl[136] vdd gnd cell_6t
Xbit_r137_c76 bl[76] br[76] wl[137] vdd gnd cell_6t
Xbit_r138_c76 bl[76] br[76] wl[138] vdd gnd cell_6t
Xbit_r139_c76 bl[76] br[76] wl[139] vdd gnd cell_6t
Xbit_r140_c76 bl[76] br[76] wl[140] vdd gnd cell_6t
Xbit_r141_c76 bl[76] br[76] wl[141] vdd gnd cell_6t
Xbit_r142_c76 bl[76] br[76] wl[142] vdd gnd cell_6t
Xbit_r143_c76 bl[76] br[76] wl[143] vdd gnd cell_6t
Xbit_r144_c76 bl[76] br[76] wl[144] vdd gnd cell_6t
Xbit_r145_c76 bl[76] br[76] wl[145] vdd gnd cell_6t
Xbit_r146_c76 bl[76] br[76] wl[146] vdd gnd cell_6t
Xbit_r147_c76 bl[76] br[76] wl[147] vdd gnd cell_6t
Xbit_r148_c76 bl[76] br[76] wl[148] vdd gnd cell_6t
Xbit_r149_c76 bl[76] br[76] wl[149] vdd gnd cell_6t
Xbit_r150_c76 bl[76] br[76] wl[150] vdd gnd cell_6t
Xbit_r151_c76 bl[76] br[76] wl[151] vdd gnd cell_6t
Xbit_r152_c76 bl[76] br[76] wl[152] vdd gnd cell_6t
Xbit_r153_c76 bl[76] br[76] wl[153] vdd gnd cell_6t
Xbit_r154_c76 bl[76] br[76] wl[154] vdd gnd cell_6t
Xbit_r155_c76 bl[76] br[76] wl[155] vdd gnd cell_6t
Xbit_r156_c76 bl[76] br[76] wl[156] vdd gnd cell_6t
Xbit_r157_c76 bl[76] br[76] wl[157] vdd gnd cell_6t
Xbit_r158_c76 bl[76] br[76] wl[158] vdd gnd cell_6t
Xbit_r159_c76 bl[76] br[76] wl[159] vdd gnd cell_6t
Xbit_r160_c76 bl[76] br[76] wl[160] vdd gnd cell_6t
Xbit_r161_c76 bl[76] br[76] wl[161] vdd gnd cell_6t
Xbit_r162_c76 bl[76] br[76] wl[162] vdd gnd cell_6t
Xbit_r163_c76 bl[76] br[76] wl[163] vdd gnd cell_6t
Xbit_r164_c76 bl[76] br[76] wl[164] vdd gnd cell_6t
Xbit_r165_c76 bl[76] br[76] wl[165] vdd gnd cell_6t
Xbit_r166_c76 bl[76] br[76] wl[166] vdd gnd cell_6t
Xbit_r167_c76 bl[76] br[76] wl[167] vdd gnd cell_6t
Xbit_r168_c76 bl[76] br[76] wl[168] vdd gnd cell_6t
Xbit_r169_c76 bl[76] br[76] wl[169] vdd gnd cell_6t
Xbit_r170_c76 bl[76] br[76] wl[170] vdd gnd cell_6t
Xbit_r171_c76 bl[76] br[76] wl[171] vdd gnd cell_6t
Xbit_r172_c76 bl[76] br[76] wl[172] vdd gnd cell_6t
Xbit_r173_c76 bl[76] br[76] wl[173] vdd gnd cell_6t
Xbit_r174_c76 bl[76] br[76] wl[174] vdd gnd cell_6t
Xbit_r175_c76 bl[76] br[76] wl[175] vdd gnd cell_6t
Xbit_r176_c76 bl[76] br[76] wl[176] vdd gnd cell_6t
Xbit_r177_c76 bl[76] br[76] wl[177] vdd gnd cell_6t
Xbit_r178_c76 bl[76] br[76] wl[178] vdd gnd cell_6t
Xbit_r179_c76 bl[76] br[76] wl[179] vdd gnd cell_6t
Xbit_r180_c76 bl[76] br[76] wl[180] vdd gnd cell_6t
Xbit_r181_c76 bl[76] br[76] wl[181] vdd gnd cell_6t
Xbit_r182_c76 bl[76] br[76] wl[182] vdd gnd cell_6t
Xbit_r183_c76 bl[76] br[76] wl[183] vdd gnd cell_6t
Xbit_r184_c76 bl[76] br[76] wl[184] vdd gnd cell_6t
Xbit_r185_c76 bl[76] br[76] wl[185] vdd gnd cell_6t
Xbit_r186_c76 bl[76] br[76] wl[186] vdd gnd cell_6t
Xbit_r187_c76 bl[76] br[76] wl[187] vdd gnd cell_6t
Xbit_r188_c76 bl[76] br[76] wl[188] vdd gnd cell_6t
Xbit_r189_c76 bl[76] br[76] wl[189] vdd gnd cell_6t
Xbit_r190_c76 bl[76] br[76] wl[190] vdd gnd cell_6t
Xbit_r191_c76 bl[76] br[76] wl[191] vdd gnd cell_6t
Xbit_r192_c76 bl[76] br[76] wl[192] vdd gnd cell_6t
Xbit_r193_c76 bl[76] br[76] wl[193] vdd gnd cell_6t
Xbit_r194_c76 bl[76] br[76] wl[194] vdd gnd cell_6t
Xbit_r195_c76 bl[76] br[76] wl[195] vdd gnd cell_6t
Xbit_r196_c76 bl[76] br[76] wl[196] vdd gnd cell_6t
Xbit_r197_c76 bl[76] br[76] wl[197] vdd gnd cell_6t
Xbit_r198_c76 bl[76] br[76] wl[198] vdd gnd cell_6t
Xbit_r199_c76 bl[76] br[76] wl[199] vdd gnd cell_6t
Xbit_r200_c76 bl[76] br[76] wl[200] vdd gnd cell_6t
Xbit_r201_c76 bl[76] br[76] wl[201] vdd gnd cell_6t
Xbit_r202_c76 bl[76] br[76] wl[202] vdd gnd cell_6t
Xbit_r203_c76 bl[76] br[76] wl[203] vdd gnd cell_6t
Xbit_r204_c76 bl[76] br[76] wl[204] vdd gnd cell_6t
Xbit_r205_c76 bl[76] br[76] wl[205] vdd gnd cell_6t
Xbit_r206_c76 bl[76] br[76] wl[206] vdd gnd cell_6t
Xbit_r207_c76 bl[76] br[76] wl[207] vdd gnd cell_6t
Xbit_r208_c76 bl[76] br[76] wl[208] vdd gnd cell_6t
Xbit_r209_c76 bl[76] br[76] wl[209] vdd gnd cell_6t
Xbit_r210_c76 bl[76] br[76] wl[210] vdd gnd cell_6t
Xbit_r211_c76 bl[76] br[76] wl[211] vdd gnd cell_6t
Xbit_r212_c76 bl[76] br[76] wl[212] vdd gnd cell_6t
Xbit_r213_c76 bl[76] br[76] wl[213] vdd gnd cell_6t
Xbit_r214_c76 bl[76] br[76] wl[214] vdd gnd cell_6t
Xbit_r215_c76 bl[76] br[76] wl[215] vdd gnd cell_6t
Xbit_r216_c76 bl[76] br[76] wl[216] vdd gnd cell_6t
Xbit_r217_c76 bl[76] br[76] wl[217] vdd gnd cell_6t
Xbit_r218_c76 bl[76] br[76] wl[218] vdd gnd cell_6t
Xbit_r219_c76 bl[76] br[76] wl[219] vdd gnd cell_6t
Xbit_r220_c76 bl[76] br[76] wl[220] vdd gnd cell_6t
Xbit_r221_c76 bl[76] br[76] wl[221] vdd gnd cell_6t
Xbit_r222_c76 bl[76] br[76] wl[222] vdd gnd cell_6t
Xbit_r223_c76 bl[76] br[76] wl[223] vdd gnd cell_6t
Xbit_r224_c76 bl[76] br[76] wl[224] vdd gnd cell_6t
Xbit_r225_c76 bl[76] br[76] wl[225] vdd gnd cell_6t
Xbit_r226_c76 bl[76] br[76] wl[226] vdd gnd cell_6t
Xbit_r227_c76 bl[76] br[76] wl[227] vdd gnd cell_6t
Xbit_r228_c76 bl[76] br[76] wl[228] vdd gnd cell_6t
Xbit_r229_c76 bl[76] br[76] wl[229] vdd gnd cell_6t
Xbit_r230_c76 bl[76] br[76] wl[230] vdd gnd cell_6t
Xbit_r231_c76 bl[76] br[76] wl[231] vdd gnd cell_6t
Xbit_r232_c76 bl[76] br[76] wl[232] vdd gnd cell_6t
Xbit_r233_c76 bl[76] br[76] wl[233] vdd gnd cell_6t
Xbit_r234_c76 bl[76] br[76] wl[234] vdd gnd cell_6t
Xbit_r235_c76 bl[76] br[76] wl[235] vdd gnd cell_6t
Xbit_r236_c76 bl[76] br[76] wl[236] vdd gnd cell_6t
Xbit_r237_c76 bl[76] br[76] wl[237] vdd gnd cell_6t
Xbit_r238_c76 bl[76] br[76] wl[238] vdd gnd cell_6t
Xbit_r239_c76 bl[76] br[76] wl[239] vdd gnd cell_6t
Xbit_r240_c76 bl[76] br[76] wl[240] vdd gnd cell_6t
Xbit_r241_c76 bl[76] br[76] wl[241] vdd gnd cell_6t
Xbit_r242_c76 bl[76] br[76] wl[242] vdd gnd cell_6t
Xbit_r243_c76 bl[76] br[76] wl[243] vdd gnd cell_6t
Xbit_r244_c76 bl[76] br[76] wl[244] vdd gnd cell_6t
Xbit_r245_c76 bl[76] br[76] wl[245] vdd gnd cell_6t
Xbit_r246_c76 bl[76] br[76] wl[246] vdd gnd cell_6t
Xbit_r247_c76 bl[76] br[76] wl[247] vdd gnd cell_6t
Xbit_r248_c76 bl[76] br[76] wl[248] vdd gnd cell_6t
Xbit_r249_c76 bl[76] br[76] wl[249] vdd gnd cell_6t
Xbit_r250_c76 bl[76] br[76] wl[250] vdd gnd cell_6t
Xbit_r251_c76 bl[76] br[76] wl[251] vdd gnd cell_6t
Xbit_r252_c76 bl[76] br[76] wl[252] vdd gnd cell_6t
Xbit_r253_c76 bl[76] br[76] wl[253] vdd gnd cell_6t
Xbit_r254_c76 bl[76] br[76] wl[254] vdd gnd cell_6t
Xbit_r255_c76 bl[76] br[76] wl[255] vdd gnd cell_6t
Xbit_r0_c77 bl[77] br[77] wl[0] vdd gnd cell_6t
Xbit_r1_c77 bl[77] br[77] wl[1] vdd gnd cell_6t
Xbit_r2_c77 bl[77] br[77] wl[2] vdd gnd cell_6t
Xbit_r3_c77 bl[77] br[77] wl[3] vdd gnd cell_6t
Xbit_r4_c77 bl[77] br[77] wl[4] vdd gnd cell_6t
Xbit_r5_c77 bl[77] br[77] wl[5] vdd gnd cell_6t
Xbit_r6_c77 bl[77] br[77] wl[6] vdd gnd cell_6t
Xbit_r7_c77 bl[77] br[77] wl[7] vdd gnd cell_6t
Xbit_r8_c77 bl[77] br[77] wl[8] vdd gnd cell_6t
Xbit_r9_c77 bl[77] br[77] wl[9] vdd gnd cell_6t
Xbit_r10_c77 bl[77] br[77] wl[10] vdd gnd cell_6t
Xbit_r11_c77 bl[77] br[77] wl[11] vdd gnd cell_6t
Xbit_r12_c77 bl[77] br[77] wl[12] vdd gnd cell_6t
Xbit_r13_c77 bl[77] br[77] wl[13] vdd gnd cell_6t
Xbit_r14_c77 bl[77] br[77] wl[14] vdd gnd cell_6t
Xbit_r15_c77 bl[77] br[77] wl[15] vdd gnd cell_6t
Xbit_r16_c77 bl[77] br[77] wl[16] vdd gnd cell_6t
Xbit_r17_c77 bl[77] br[77] wl[17] vdd gnd cell_6t
Xbit_r18_c77 bl[77] br[77] wl[18] vdd gnd cell_6t
Xbit_r19_c77 bl[77] br[77] wl[19] vdd gnd cell_6t
Xbit_r20_c77 bl[77] br[77] wl[20] vdd gnd cell_6t
Xbit_r21_c77 bl[77] br[77] wl[21] vdd gnd cell_6t
Xbit_r22_c77 bl[77] br[77] wl[22] vdd gnd cell_6t
Xbit_r23_c77 bl[77] br[77] wl[23] vdd gnd cell_6t
Xbit_r24_c77 bl[77] br[77] wl[24] vdd gnd cell_6t
Xbit_r25_c77 bl[77] br[77] wl[25] vdd gnd cell_6t
Xbit_r26_c77 bl[77] br[77] wl[26] vdd gnd cell_6t
Xbit_r27_c77 bl[77] br[77] wl[27] vdd gnd cell_6t
Xbit_r28_c77 bl[77] br[77] wl[28] vdd gnd cell_6t
Xbit_r29_c77 bl[77] br[77] wl[29] vdd gnd cell_6t
Xbit_r30_c77 bl[77] br[77] wl[30] vdd gnd cell_6t
Xbit_r31_c77 bl[77] br[77] wl[31] vdd gnd cell_6t
Xbit_r32_c77 bl[77] br[77] wl[32] vdd gnd cell_6t
Xbit_r33_c77 bl[77] br[77] wl[33] vdd gnd cell_6t
Xbit_r34_c77 bl[77] br[77] wl[34] vdd gnd cell_6t
Xbit_r35_c77 bl[77] br[77] wl[35] vdd gnd cell_6t
Xbit_r36_c77 bl[77] br[77] wl[36] vdd gnd cell_6t
Xbit_r37_c77 bl[77] br[77] wl[37] vdd gnd cell_6t
Xbit_r38_c77 bl[77] br[77] wl[38] vdd gnd cell_6t
Xbit_r39_c77 bl[77] br[77] wl[39] vdd gnd cell_6t
Xbit_r40_c77 bl[77] br[77] wl[40] vdd gnd cell_6t
Xbit_r41_c77 bl[77] br[77] wl[41] vdd gnd cell_6t
Xbit_r42_c77 bl[77] br[77] wl[42] vdd gnd cell_6t
Xbit_r43_c77 bl[77] br[77] wl[43] vdd gnd cell_6t
Xbit_r44_c77 bl[77] br[77] wl[44] vdd gnd cell_6t
Xbit_r45_c77 bl[77] br[77] wl[45] vdd gnd cell_6t
Xbit_r46_c77 bl[77] br[77] wl[46] vdd gnd cell_6t
Xbit_r47_c77 bl[77] br[77] wl[47] vdd gnd cell_6t
Xbit_r48_c77 bl[77] br[77] wl[48] vdd gnd cell_6t
Xbit_r49_c77 bl[77] br[77] wl[49] vdd gnd cell_6t
Xbit_r50_c77 bl[77] br[77] wl[50] vdd gnd cell_6t
Xbit_r51_c77 bl[77] br[77] wl[51] vdd gnd cell_6t
Xbit_r52_c77 bl[77] br[77] wl[52] vdd gnd cell_6t
Xbit_r53_c77 bl[77] br[77] wl[53] vdd gnd cell_6t
Xbit_r54_c77 bl[77] br[77] wl[54] vdd gnd cell_6t
Xbit_r55_c77 bl[77] br[77] wl[55] vdd gnd cell_6t
Xbit_r56_c77 bl[77] br[77] wl[56] vdd gnd cell_6t
Xbit_r57_c77 bl[77] br[77] wl[57] vdd gnd cell_6t
Xbit_r58_c77 bl[77] br[77] wl[58] vdd gnd cell_6t
Xbit_r59_c77 bl[77] br[77] wl[59] vdd gnd cell_6t
Xbit_r60_c77 bl[77] br[77] wl[60] vdd gnd cell_6t
Xbit_r61_c77 bl[77] br[77] wl[61] vdd gnd cell_6t
Xbit_r62_c77 bl[77] br[77] wl[62] vdd gnd cell_6t
Xbit_r63_c77 bl[77] br[77] wl[63] vdd gnd cell_6t
Xbit_r64_c77 bl[77] br[77] wl[64] vdd gnd cell_6t
Xbit_r65_c77 bl[77] br[77] wl[65] vdd gnd cell_6t
Xbit_r66_c77 bl[77] br[77] wl[66] vdd gnd cell_6t
Xbit_r67_c77 bl[77] br[77] wl[67] vdd gnd cell_6t
Xbit_r68_c77 bl[77] br[77] wl[68] vdd gnd cell_6t
Xbit_r69_c77 bl[77] br[77] wl[69] vdd gnd cell_6t
Xbit_r70_c77 bl[77] br[77] wl[70] vdd gnd cell_6t
Xbit_r71_c77 bl[77] br[77] wl[71] vdd gnd cell_6t
Xbit_r72_c77 bl[77] br[77] wl[72] vdd gnd cell_6t
Xbit_r73_c77 bl[77] br[77] wl[73] vdd gnd cell_6t
Xbit_r74_c77 bl[77] br[77] wl[74] vdd gnd cell_6t
Xbit_r75_c77 bl[77] br[77] wl[75] vdd gnd cell_6t
Xbit_r76_c77 bl[77] br[77] wl[76] vdd gnd cell_6t
Xbit_r77_c77 bl[77] br[77] wl[77] vdd gnd cell_6t
Xbit_r78_c77 bl[77] br[77] wl[78] vdd gnd cell_6t
Xbit_r79_c77 bl[77] br[77] wl[79] vdd gnd cell_6t
Xbit_r80_c77 bl[77] br[77] wl[80] vdd gnd cell_6t
Xbit_r81_c77 bl[77] br[77] wl[81] vdd gnd cell_6t
Xbit_r82_c77 bl[77] br[77] wl[82] vdd gnd cell_6t
Xbit_r83_c77 bl[77] br[77] wl[83] vdd gnd cell_6t
Xbit_r84_c77 bl[77] br[77] wl[84] vdd gnd cell_6t
Xbit_r85_c77 bl[77] br[77] wl[85] vdd gnd cell_6t
Xbit_r86_c77 bl[77] br[77] wl[86] vdd gnd cell_6t
Xbit_r87_c77 bl[77] br[77] wl[87] vdd gnd cell_6t
Xbit_r88_c77 bl[77] br[77] wl[88] vdd gnd cell_6t
Xbit_r89_c77 bl[77] br[77] wl[89] vdd gnd cell_6t
Xbit_r90_c77 bl[77] br[77] wl[90] vdd gnd cell_6t
Xbit_r91_c77 bl[77] br[77] wl[91] vdd gnd cell_6t
Xbit_r92_c77 bl[77] br[77] wl[92] vdd gnd cell_6t
Xbit_r93_c77 bl[77] br[77] wl[93] vdd gnd cell_6t
Xbit_r94_c77 bl[77] br[77] wl[94] vdd gnd cell_6t
Xbit_r95_c77 bl[77] br[77] wl[95] vdd gnd cell_6t
Xbit_r96_c77 bl[77] br[77] wl[96] vdd gnd cell_6t
Xbit_r97_c77 bl[77] br[77] wl[97] vdd gnd cell_6t
Xbit_r98_c77 bl[77] br[77] wl[98] vdd gnd cell_6t
Xbit_r99_c77 bl[77] br[77] wl[99] vdd gnd cell_6t
Xbit_r100_c77 bl[77] br[77] wl[100] vdd gnd cell_6t
Xbit_r101_c77 bl[77] br[77] wl[101] vdd gnd cell_6t
Xbit_r102_c77 bl[77] br[77] wl[102] vdd gnd cell_6t
Xbit_r103_c77 bl[77] br[77] wl[103] vdd gnd cell_6t
Xbit_r104_c77 bl[77] br[77] wl[104] vdd gnd cell_6t
Xbit_r105_c77 bl[77] br[77] wl[105] vdd gnd cell_6t
Xbit_r106_c77 bl[77] br[77] wl[106] vdd gnd cell_6t
Xbit_r107_c77 bl[77] br[77] wl[107] vdd gnd cell_6t
Xbit_r108_c77 bl[77] br[77] wl[108] vdd gnd cell_6t
Xbit_r109_c77 bl[77] br[77] wl[109] vdd gnd cell_6t
Xbit_r110_c77 bl[77] br[77] wl[110] vdd gnd cell_6t
Xbit_r111_c77 bl[77] br[77] wl[111] vdd gnd cell_6t
Xbit_r112_c77 bl[77] br[77] wl[112] vdd gnd cell_6t
Xbit_r113_c77 bl[77] br[77] wl[113] vdd gnd cell_6t
Xbit_r114_c77 bl[77] br[77] wl[114] vdd gnd cell_6t
Xbit_r115_c77 bl[77] br[77] wl[115] vdd gnd cell_6t
Xbit_r116_c77 bl[77] br[77] wl[116] vdd gnd cell_6t
Xbit_r117_c77 bl[77] br[77] wl[117] vdd gnd cell_6t
Xbit_r118_c77 bl[77] br[77] wl[118] vdd gnd cell_6t
Xbit_r119_c77 bl[77] br[77] wl[119] vdd gnd cell_6t
Xbit_r120_c77 bl[77] br[77] wl[120] vdd gnd cell_6t
Xbit_r121_c77 bl[77] br[77] wl[121] vdd gnd cell_6t
Xbit_r122_c77 bl[77] br[77] wl[122] vdd gnd cell_6t
Xbit_r123_c77 bl[77] br[77] wl[123] vdd gnd cell_6t
Xbit_r124_c77 bl[77] br[77] wl[124] vdd gnd cell_6t
Xbit_r125_c77 bl[77] br[77] wl[125] vdd gnd cell_6t
Xbit_r126_c77 bl[77] br[77] wl[126] vdd gnd cell_6t
Xbit_r127_c77 bl[77] br[77] wl[127] vdd gnd cell_6t
Xbit_r128_c77 bl[77] br[77] wl[128] vdd gnd cell_6t
Xbit_r129_c77 bl[77] br[77] wl[129] vdd gnd cell_6t
Xbit_r130_c77 bl[77] br[77] wl[130] vdd gnd cell_6t
Xbit_r131_c77 bl[77] br[77] wl[131] vdd gnd cell_6t
Xbit_r132_c77 bl[77] br[77] wl[132] vdd gnd cell_6t
Xbit_r133_c77 bl[77] br[77] wl[133] vdd gnd cell_6t
Xbit_r134_c77 bl[77] br[77] wl[134] vdd gnd cell_6t
Xbit_r135_c77 bl[77] br[77] wl[135] vdd gnd cell_6t
Xbit_r136_c77 bl[77] br[77] wl[136] vdd gnd cell_6t
Xbit_r137_c77 bl[77] br[77] wl[137] vdd gnd cell_6t
Xbit_r138_c77 bl[77] br[77] wl[138] vdd gnd cell_6t
Xbit_r139_c77 bl[77] br[77] wl[139] vdd gnd cell_6t
Xbit_r140_c77 bl[77] br[77] wl[140] vdd gnd cell_6t
Xbit_r141_c77 bl[77] br[77] wl[141] vdd gnd cell_6t
Xbit_r142_c77 bl[77] br[77] wl[142] vdd gnd cell_6t
Xbit_r143_c77 bl[77] br[77] wl[143] vdd gnd cell_6t
Xbit_r144_c77 bl[77] br[77] wl[144] vdd gnd cell_6t
Xbit_r145_c77 bl[77] br[77] wl[145] vdd gnd cell_6t
Xbit_r146_c77 bl[77] br[77] wl[146] vdd gnd cell_6t
Xbit_r147_c77 bl[77] br[77] wl[147] vdd gnd cell_6t
Xbit_r148_c77 bl[77] br[77] wl[148] vdd gnd cell_6t
Xbit_r149_c77 bl[77] br[77] wl[149] vdd gnd cell_6t
Xbit_r150_c77 bl[77] br[77] wl[150] vdd gnd cell_6t
Xbit_r151_c77 bl[77] br[77] wl[151] vdd gnd cell_6t
Xbit_r152_c77 bl[77] br[77] wl[152] vdd gnd cell_6t
Xbit_r153_c77 bl[77] br[77] wl[153] vdd gnd cell_6t
Xbit_r154_c77 bl[77] br[77] wl[154] vdd gnd cell_6t
Xbit_r155_c77 bl[77] br[77] wl[155] vdd gnd cell_6t
Xbit_r156_c77 bl[77] br[77] wl[156] vdd gnd cell_6t
Xbit_r157_c77 bl[77] br[77] wl[157] vdd gnd cell_6t
Xbit_r158_c77 bl[77] br[77] wl[158] vdd gnd cell_6t
Xbit_r159_c77 bl[77] br[77] wl[159] vdd gnd cell_6t
Xbit_r160_c77 bl[77] br[77] wl[160] vdd gnd cell_6t
Xbit_r161_c77 bl[77] br[77] wl[161] vdd gnd cell_6t
Xbit_r162_c77 bl[77] br[77] wl[162] vdd gnd cell_6t
Xbit_r163_c77 bl[77] br[77] wl[163] vdd gnd cell_6t
Xbit_r164_c77 bl[77] br[77] wl[164] vdd gnd cell_6t
Xbit_r165_c77 bl[77] br[77] wl[165] vdd gnd cell_6t
Xbit_r166_c77 bl[77] br[77] wl[166] vdd gnd cell_6t
Xbit_r167_c77 bl[77] br[77] wl[167] vdd gnd cell_6t
Xbit_r168_c77 bl[77] br[77] wl[168] vdd gnd cell_6t
Xbit_r169_c77 bl[77] br[77] wl[169] vdd gnd cell_6t
Xbit_r170_c77 bl[77] br[77] wl[170] vdd gnd cell_6t
Xbit_r171_c77 bl[77] br[77] wl[171] vdd gnd cell_6t
Xbit_r172_c77 bl[77] br[77] wl[172] vdd gnd cell_6t
Xbit_r173_c77 bl[77] br[77] wl[173] vdd gnd cell_6t
Xbit_r174_c77 bl[77] br[77] wl[174] vdd gnd cell_6t
Xbit_r175_c77 bl[77] br[77] wl[175] vdd gnd cell_6t
Xbit_r176_c77 bl[77] br[77] wl[176] vdd gnd cell_6t
Xbit_r177_c77 bl[77] br[77] wl[177] vdd gnd cell_6t
Xbit_r178_c77 bl[77] br[77] wl[178] vdd gnd cell_6t
Xbit_r179_c77 bl[77] br[77] wl[179] vdd gnd cell_6t
Xbit_r180_c77 bl[77] br[77] wl[180] vdd gnd cell_6t
Xbit_r181_c77 bl[77] br[77] wl[181] vdd gnd cell_6t
Xbit_r182_c77 bl[77] br[77] wl[182] vdd gnd cell_6t
Xbit_r183_c77 bl[77] br[77] wl[183] vdd gnd cell_6t
Xbit_r184_c77 bl[77] br[77] wl[184] vdd gnd cell_6t
Xbit_r185_c77 bl[77] br[77] wl[185] vdd gnd cell_6t
Xbit_r186_c77 bl[77] br[77] wl[186] vdd gnd cell_6t
Xbit_r187_c77 bl[77] br[77] wl[187] vdd gnd cell_6t
Xbit_r188_c77 bl[77] br[77] wl[188] vdd gnd cell_6t
Xbit_r189_c77 bl[77] br[77] wl[189] vdd gnd cell_6t
Xbit_r190_c77 bl[77] br[77] wl[190] vdd gnd cell_6t
Xbit_r191_c77 bl[77] br[77] wl[191] vdd gnd cell_6t
Xbit_r192_c77 bl[77] br[77] wl[192] vdd gnd cell_6t
Xbit_r193_c77 bl[77] br[77] wl[193] vdd gnd cell_6t
Xbit_r194_c77 bl[77] br[77] wl[194] vdd gnd cell_6t
Xbit_r195_c77 bl[77] br[77] wl[195] vdd gnd cell_6t
Xbit_r196_c77 bl[77] br[77] wl[196] vdd gnd cell_6t
Xbit_r197_c77 bl[77] br[77] wl[197] vdd gnd cell_6t
Xbit_r198_c77 bl[77] br[77] wl[198] vdd gnd cell_6t
Xbit_r199_c77 bl[77] br[77] wl[199] vdd gnd cell_6t
Xbit_r200_c77 bl[77] br[77] wl[200] vdd gnd cell_6t
Xbit_r201_c77 bl[77] br[77] wl[201] vdd gnd cell_6t
Xbit_r202_c77 bl[77] br[77] wl[202] vdd gnd cell_6t
Xbit_r203_c77 bl[77] br[77] wl[203] vdd gnd cell_6t
Xbit_r204_c77 bl[77] br[77] wl[204] vdd gnd cell_6t
Xbit_r205_c77 bl[77] br[77] wl[205] vdd gnd cell_6t
Xbit_r206_c77 bl[77] br[77] wl[206] vdd gnd cell_6t
Xbit_r207_c77 bl[77] br[77] wl[207] vdd gnd cell_6t
Xbit_r208_c77 bl[77] br[77] wl[208] vdd gnd cell_6t
Xbit_r209_c77 bl[77] br[77] wl[209] vdd gnd cell_6t
Xbit_r210_c77 bl[77] br[77] wl[210] vdd gnd cell_6t
Xbit_r211_c77 bl[77] br[77] wl[211] vdd gnd cell_6t
Xbit_r212_c77 bl[77] br[77] wl[212] vdd gnd cell_6t
Xbit_r213_c77 bl[77] br[77] wl[213] vdd gnd cell_6t
Xbit_r214_c77 bl[77] br[77] wl[214] vdd gnd cell_6t
Xbit_r215_c77 bl[77] br[77] wl[215] vdd gnd cell_6t
Xbit_r216_c77 bl[77] br[77] wl[216] vdd gnd cell_6t
Xbit_r217_c77 bl[77] br[77] wl[217] vdd gnd cell_6t
Xbit_r218_c77 bl[77] br[77] wl[218] vdd gnd cell_6t
Xbit_r219_c77 bl[77] br[77] wl[219] vdd gnd cell_6t
Xbit_r220_c77 bl[77] br[77] wl[220] vdd gnd cell_6t
Xbit_r221_c77 bl[77] br[77] wl[221] vdd gnd cell_6t
Xbit_r222_c77 bl[77] br[77] wl[222] vdd gnd cell_6t
Xbit_r223_c77 bl[77] br[77] wl[223] vdd gnd cell_6t
Xbit_r224_c77 bl[77] br[77] wl[224] vdd gnd cell_6t
Xbit_r225_c77 bl[77] br[77] wl[225] vdd gnd cell_6t
Xbit_r226_c77 bl[77] br[77] wl[226] vdd gnd cell_6t
Xbit_r227_c77 bl[77] br[77] wl[227] vdd gnd cell_6t
Xbit_r228_c77 bl[77] br[77] wl[228] vdd gnd cell_6t
Xbit_r229_c77 bl[77] br[77] wl[229] vdd gnd cell_6t
Xbit_r230_c77 bl[77] br[77] wl[230] vdd gnd cell_6t
Xbit_r231_c77 bl[77] br[77] wl[231] vdd gnd cell_6t
Xbit_r232_c77 bl[77] br[77] wl[232] vdd gnd cell_6t
Xbit_r233_c77 bl[77] br[77] wl[233] vdd gnd cell_6t
Xbit_r234_c77 bl[77] br[77] wl[234] vdd gnd cell_6t
Xbit_r235_c77 bl[77] br[77] wl[235] vdd gnd cell_6t
Xbit_r236_c77 bl[77] br[77] wl[236] vdd gnd cell_6t
Xbit_r237_c77 bl[77] br[77] wl[237] vdd gnd cell_6t
Xbit_r238_c77 bl[77] br[77] wl[238] vdd gnd cell_6t
Xbit_r239_c77 bl[77] br[77] wl[239] vdd gnd cell_6t
Xbit_r240_c77 bl[77] br[77] wl[240] vdd gnd cell_6t
Xbit_r241_c77 bl[77] br[77] wl[241] vdd gnd cell_6t
Xbit_r242_c77 bl[77] br[77] wl[242] vdd gnd cell_6t
Xbit_r243_c77 bl[77] br[77] wl[243] vdd gnd cell_6t
Xbit_r244_c77 bl[77] br[77] wl[244] vdd gnd cell_6t
Xbit_r245_c77 bl[77] br[77] wl[245] vdd gnd cell_6t
Xbit_r246_c77 bl[77] br[77] wl[246] vdd gnd cell_6t
Xbit_r247_c77 bl[77] br[77] wl[247] vdd gnd cell_6t
Xbit_r248_c77 bl[77] br[77] wl[248] vdd gnd cell_6t
Xbit_r249_c77 bl[77] br[77] wl[249] vdd gnd cell_6t
Xbit_r250_c77 bl[77] br[77] wl[250] vdd gnd cell_6t
Xbit_r251_c77 bl[77] br[77] wl[251] vdd gnd cell_6t
Xbit_r252_c77 bl[77] br[77] wl[252] vdd gnd cell_6t
Xbit_r253_c77 bl[77] br[77] wl[253] vdd gnd cell_6t
Xbit_r254_c77 bl[77] br[77] wl[254] vdd gnd cell_6t
Xbit_r255_c77 bl[77] br[77] wl[255] vdd gnd cell_6t
Xbit_r0_c78 bl[78] br[78] wl[0] vdd gnd cell_6t
Xbit_r1_c78 bl[78] br[78] wl[1] vdd gnd cell_6t
Xbit_r2_c78 bl[78] br[78] wl[2] vdd gnd cell_6t
Xbit_r3_c78 bl[78] br[78] wl[3] vdd gnd cell_6t
Xbit_r4_c78 bl[78] br[78] wl[4] vdd gnd cell_6t
Xbit_r5_c78 bl[78] br[78] wl[5] vdd gnd cell_6t
Xbit_r6_c78 bl[78] br[78] wl[6] vdd gnd cell_6t
Xbit_r7_c78 bl[78] br[78] wl[7] vdd gnd cell_6t
Xbit_r8_c78 bl[78] br[78] wl[8] vdd gnd cell_6t
Xbit_r9_c78 bl[78] br[78] wl[9] vdd gnd cell_6t
Xbit_r10_c78 bl[78] br[78] wl[10] vdd gnd cell_6t
Xbit_r11_c78 bl[78] br[78] wl[11] vdd gnd cell_6t
Xbit_r12_c78 bl[78] br[78] wl[12] vdd gnd cell_6t
Xbit_r13_c78 bl[78] br[78] wl[13] vdd gnd cell_6t
Xbit_r14_c78 bl[78] br[78] wl[14] vdd gnd cell_6t
Xbit_r15_c78 bl[78] br[78] wl[15] vdd gnd cell_6t
Xbit_r16_c78 bl[78] br[78] wl[16] vdd gnd cell_6t
Xbit_r17_c78 bl[78] br[78] wl[17] vdd gnd cell_6t
Xbit_r18_c78 bl[78] br[78] wl[18] vdd gnd cell_6t
Xbit_r19_c78 bl[78] br[78] wl[19] vdd gnd cell_6t
Xbit_r20_c78 bl[78] br[78] wl[20] vdd gnd cell_6t
Xbit_r21_c78 bl[78] br[78] wl[21] vdd gnd cell_6t
Xbit_r22_c78 bl[78] br[78] wl[22] vdd gnd cell_6t
Xbit_r23_c78 bl[78] br[78] wl[23] vdd gnd cell_6t
Xbit_r24_c78 bl[78] br[78] wl[24] vdd gnd cell_6t
Xbit_r25_c78 bl[78] br[78] wl[25] vdd gnd cell_6t
Xbit_r26_c78 bl[78] br[78] wl[26] vdd gnd cell_6t
Xbit_r27_c78 bl[78] br[78] wl[27] vdd gnd cell_6t
Xbit_r28_c78 bl[78] br[78] wl[28] vdd gnd cell_6t
Xbit_r29_c78 bl[78] br[78] wl[29] vdd gnd cell_6t
Xbit_r30_c78 bl[78] br[78] wl[30] vdd gnd cell_6t
Xbit_r31_c78 bl[78] br[78] wl[31] vdd gnd cell_6t
Xbit_r32_c78 bl[78] br[78] wl[32] vdd gnd cell_6t
Xbit_r33_c78 bl[78] br[78] wl[33] vdd gnd cell_6t
Xbit_r34_c78 bl[78] br[78] wl[34] vdd gnd cell_6t
Xbit_r35_c78 bl[78] br[78] wl[35] vdd gnd cell_6t
Xbit_r36_c78 bl[78] br[78] wl[36] vdd gnd cell_6t
Xbit_r37_c78 bl[78] br[78] wl[37] vdd gnd cell_6t
Xbit_r38_c78 bl[78] br[78] wl[38] vdd gnd cell_6t
Xbit_r39_c78 bl[78] br[78] wl[39] vdd gnd cell_6t
Xbit_r40_c78 bl[78] br[78] wl[40] vdd gnd cell_6t
Xbit_r41_c78 bl[78] br[78] wl[41] vdd gnd cell_6t
Xbit_r42_c78 bl[78] br[78] wl[42] vdd gnd cell_6t
Xbit_r43_c78 bl[78] br[78] wl[43] vdd gnd cell_6t
Xbit_r44_c78 bl[78] br[78] wl[44] vdd gnd cell_6t
Xbit_r45_c78 bl[78] br[78] wl[45] vdd gnd cell_6t
Xbit_r46_c78 bl[78] br[78] wl[46] vdd gnd cell_6t
Xbit_r47_c78 bl[78] br[78] wl[47] vdd gnd cell_6t
Xbit_r48_c78 bl[78] br[78] wl[48] vdd gnd cell_6t
Xbit_r49_c78 bl[78] br[78] wl[49] vdd gnd cell_6t
Xbit_r50_c78 bl[78] br[78] wl[50] vdd gnd cell_6t
Xbit_r51_c78 bl[78] br[78] wl[51] vdd gnd cell_6t
Xbit_r52_c78 bl[78] br[78] wl[52] vdd gnd cell_6t
Xbit_r53_c78 bl[78] br[78] wl[53] vdd gnd cell_6t
Xbit_r54_c78 bl[78] br[78] wl[54] vdd gnd cell_6t
Xbit_r55_c78 bl[78] br[78] wl[55] vdd gnd cell_6t
Xbit_r56_c78 bl[78] br[78] wl[56] vdd gnd cell_6t
Xbit_r57_c78 bl[78] br[78] wl[57] vdd gnd cell_6t
Xbit_r58_c78 bl[78] br[78] wl[58] vdd gnd cell_6t
Xbit_r59_c78 bl[78] br[78] wl[59] vdd gnd cell_6t
Xbit_r60_c78 bl[78] br[78] wl[60] vdd gnd cell_6t
Xbit_r61_c78 bl[78] br[78] wl[61] vdd gnd cell_6t
Xbit_r62_c78 bl[78] br[78] wl[62] vdd gnd cell_6t
Xbit_r63_c78 bl[78] br[78] wl[63] vdd gnd cell_6t
Xbit_r64_c78 bl[78] br[78] wl[64] vdd gnd cell_6t
Xbit_r65_c78 bl[78] br[78] wl[65] vdd gnd cell_6t
Xbit_r66_c78 bl[78] br[78] wl[66] vdd gnd cell_6t
Xbit_r67_c78 bl[78] br[78] wl[67] vdd gnd cell_6t
Xbit_r68_c78 bl[78] br[78] wl[68] vdd gnd cell_6t
Xbit_r69_c78 bl[78] br[78] wl[69] vdd gnd cell_6t
Xbit_r70_c78 bl[78] br[78] wl[70] vdd gnd cell_6t
Xbit_r71_c78 bl[78] br[78] wl[71] vdd gnd cell_6t
Xbit_r72_c78 bl[78] br[78] wl[72] vdd gnd cell_6t
Xbit_r73_c78 bl[78] br[78] wl[73] vdd gnd cell_6t
Xbit_r74_c78 bl[78] br[78] wl[74] vdd gnd cell_6t
Xbit_r75_c78 bl[78] br[78] wl[75] vdd gnd cell_6t
Xbit_r76_c78 bl[78] br[78] wl[76] vdd gnd cell_6t
Xbit_r77_c78 bl[78] br[78] wl[77] vdd gnd cell_6t
Xbit_r78_c78 bl[78] br[78] wl[78] vdd gnd cell_6t
Xbit_r79_c78 bl[78] br[78] wl[79] vdd gnd cell_6t
Xbit_r80_c78 bl[78] br[78] wl[80] vdd gnd cell_6t
Xbit_r81_c78 bl[78] br[78] wl[81] vdd gnd cell_6t
Xbit_r82_c78 bl[78] br[78] wl[82] vdd gnd cell_6t
Xbit_r83_c78 bl[78] br[78] wl[83] vdd gnd cell_6t
Xbit_r84_c78 bl[78] br[78] wl[84] vdd gnd cell_6t
Xbit_r85_c78 bl[78] br[78] wl[85] vdd gnd cell_6t
Xbit_r86_c78 bl[78] br[78] wl[86] vdd gnd cell_6t
Xbit_r87_c78 bl[78] br[78] wl[87] vdd gnd cell_6t
Xbit_r88_c78 bl[78] br[78] wl[88] vdd gnd cell_6t
Xbit_r89_c78 bl[78] br[78] wl[89] vdd gnd cell_6t
Xbit_r90_c78 bl[78] br[78] wl[90] vdd gnd cell_6t
Xbit_r91_c78 bl[78] br[78] wl[91] vdd gnd cell_6t
Xbit_r92_c78 bl[78] br[78] wl[92] vdd gnd cell_6t
Xbit_r93_c78 bl[78] br[78] wl[93] vdd gnd cell_6t
Xbit_r94_c78 bl[78] br[78] wl[94] vdd gnd cell_6t
Xbit_r95_c78 bl[78] br[78] wl[95] vdd gnd cell_6t
Xbit_r96_c78 bl[78] br[78] wl[96] vdd gnd cell_6t
Xbit_r97_c78 bl[78] br[78] wl[97] vdd gnd cell_6t
Xbit_r98_c78 bl[78] br[78] wl[98] vdd gnd cell_6t
Xbit_r99_c78 bl[78] br[78] wl[99] vdd gnd cell_6t
Xbit_r100_c78 bl[78] br[78] wl[100] vdd gnd cell_6t
Xbit_r101_c78 bl[78] br[78] wl[101] vdd gnd cell_6t
Xbit_r102_c78 bl[78] br[78] wl[102] vdd gnd cell_6t
Xbit_r103_c78 bl[78] br[78] wl[103] vdd gnd cell_6t
Xbit_r104_c78 bl[78] br[78] wl[104] vdd gnd cell_6t
Xbit_r105_c78 bl[78] br[78] wl[105] vdd gnd cell_6t
Xbit_r106_c78 bl[78] br[78] wl[106] vdd gnd cell_6t
Xbit_r107_c78 bl[78] br[78] wl[107] vdd gnd cell_6t
Xbit_r108_c78 bl[78] br[78] wl[108] vdd gnd cell_6t
Xbit_r109_c78 bl[78] br[78] wl[109] vdd gnd cell_6t
Xbit_r110_c78 bl[78] br[78] wl[110] vdd gnd cell_6t
Xbit_r111_c78 bl[78] br[78] wl[111] vdd gnd cell_6t
Xbit_r112_c78 bl[78] br[78] wl[112] vdd gnd cell_6t
Xbit_r113_c78 bl[78] br[78] wl[113] vdd gnd cell_6t
Xbit_r114_c78 bl[78] br[78] wl[114] vdd gnd cell_6t
Xbit_r115_c78 bl[78] br[78] wl[115] vdd gnd cell_6t
Xbit_r116_c78 bl[78] br[78] wl[116] vdd gnd cell_6t
Xbit_r117_c78 bl[78] br[78] wl[117] vdd gnd cell_6t
Xbit_r118_c78 bl[78] br[78] wl[118] vdd gnd cell_6t
Xbit_r119_c78 bl[78] br[78] wl[119] vdd gnd cell_6t
Xbit_r120_c78 bl[78] br[78] wl[120] vdd gnd cell_6t
Xbit_r121_c78 bl[78] br[78] wl[121] vdd gnd cell_6t
Xbit_r122_c78 bl[78] br[78] wl[122] vdd gnd cell_6t
Xbit_r123_c78 bl[78] br[78] wl[123] vdd gnd cell_6t
Xbit_r124_c78 bl[78] br[78] wl[124] vdd gnd cell_6t
Xbit_r125_c78 bl[78] br[78] wl[125] vdd gnd cell_6t
Xbit_r126_c78 bl[78] br[78] wl[126] vdd gnd cell_6t
Xbit_r127_c78 bl[78] br[78] wl[127] vdd gnd cell_6t
Xbit_r128_c78 bl[78] br[78] wl[128] vdd gnd cell_6t
Xbit_r129_c78 bl[78] br[78] wl[129] vdd gnd cell_6t
Xbit_r130_c78 bl[78] br[78] wl[130] vdd gnd cell_6t
Xbit_r131_c78 bl[78] br[78] wl[131] vdd gnd cell_6t
Xbit_r132_c78 bl[78] br[78] wl[132] vdd gnd cell_6t
Xbit_r133_c78 bl[78] br[78] wl[133] vdd gnd cell_6t
Xbit_r134_c78 bl[78] br[78] wl[134] vdd gnd cell_6t
Xbit_r135_c78 bl[78] br[78] wl[135] vdd gnd cell_6t
Xbit_r136_c78 bl[78] br[78] wl[136] vdd gnd cell_6t
Xbit_r137_c78 bl[78] br[78] wl[137] vdd gnd cell_6t
Xbit_r138_c78 bl[78] br[78] wl[138] vdd gnd cell_6t
Xbit_r139_c78 bl[78] br[78] wl[139] vdd gnd cell_6t
Xbit_r140_c78 bl[78] br[78] wl[140] vdd gnd cell_6t
Xbit_r141_c78 bl[78] br[78] wl[141] vdd gnd cell_6t
Xbit_r142_c78 bl[78] br[78] wl[142] vdd gnd cell_6t
Xbit_r143_c78 bl[78] br[78] wl[143] vdd gnd cell_6t
Xbit_r144_c78 bl[78] br[78] wl[144] vdd gnd cell_6t
Xbit_r145_c78 bl[78] br[78] wl[145] vdd gnd cell_6t
Xbit_r146_c78 bl[78] br[78] wl[146] vdd gnd cell_6t
Xbit_r147_c78 bl[78] br[78] wl[147] vdd gnd cell_6t
Xbit_r148_c78 bl[78] br[78] wl[148] vdd gnd cell_6t
Xbit_r149_c78 bl[78] br[78] wl[149] vdd gnd cell_6t
Xbit_r150_c78 bl[78] br[78] wl[150] vdd gnd cell_6t
Xbit_r151_c78 bl[78] br[78] wl[151] vdd gnd cell_6t
Xbit_r152_c78 bl[78] br[78] wl[152] vdd gnd cell_6t
Xbit_r153_c78 bl[78] br[78] wl[153] vdd gnd cell_6t
Xbit_r154_c78 bl[78] br[78] wl[154] vdd gnd cell_6t
Xbit_r155_c78 bl[78] br[78] wl[155] vdd gnd cell_6t
Xbit_r156_c78 bl[78] br[78] wl[156] vdd gnd cell_6t
Xbit_r157_c78 bl[78] br[78] wl[157] vdd gnd cell_6t
Xbit_r158_c78 bl[78] br[78] wl[158] vdd gnd cell_6t
Xbit_r159_c78 bl[78] br[78] wl[159] vdd gnd cell_6t
Xbit_r160_c78 bl[78] br[78] wl[160] vdd gnd cell_6t
Xbit_r161_c78 bl[78] br[78] wl[161] vdd gnd cell_6t
Xbit_r162_c78 bl[78] br[78] wl[162] vdd gnd cell_6t
Xbit_r163_c78 bl[78] br[78] wl[163] vdd gnd cell_6t
Xbit_r164_c78 bl[78] br[78] wl[164] vdd gnd cell_6t
Xbit_r165_c78 bl[78] br[78] wl[165] vdd gnd cell_6t
Xbit_r166_c78 bl[78] br[78] wl[166] vdd gnd cell_6t
Xbit_r167_c78 bl[78] br[78] wl[167] vdd gnd cell_6t
Xbit_r168_c78 bl[78] br[78] wl[168] vdd gnd cell_6t
Xbit_r169_c78 bl[78] br[78] wl[169] vdd gnd cell_6t
Xbit_r170_c78 bl[78] br[78] wl[170] vdd gnd cell_6t
Xbit_r171_c78 bl[78] br[78] wl[171] vdd gnd cell_6t
Xbit_r172_c78 bl[78] br[78] wl[172] vdd gnd cell_6t
Xbit_r173_c78 bl[78] br[78] wl[173] vdd gnd cell_6t
Xbit_r174_c78 bl[78] br[78] wl[174] vdd gnd cell_6t
Xbit_r175_c78 bl[78] br[78] wl[175] vdd gnd cell_6t
Xbit_r176_c78 bl[78] br[78] wl[176] vdd gnd cell_6t
Xbit_r177_c78 bl[78] br[78] wl[177] vdd gnd cell_6t
Xbit_r178_c78 bl[78] br[78] wl[178] vdd gnd cell_6t
Xbit_r179_c78 bl[78] br[78] wl[179] vdd gnd cell_6t
Xbit_r180_c78 bl[78] br[78] wl[180] vdd gnd cell_6t
Xbit_r181_c78 bl[78] br[78] wl[181] vdd gnd cell_6t
Xbit_r182_c78 bl[78] br[78] wl[182] vdd gnd cell_6t
Xbit_r183_c78 bl[78] br[78] wl[183] vdd gnd cell_6t
Xbit_r184_c78 bl[78] br[78] wl[184] vdd gnd cell_6t
Xbit_r185_c78 bl[78] br[78] wl[185] vdd gnd cell_6t
Xbit_r186_c78 bl[78] br[78] wl[186] vdd gnd cell_6t
Xbit_r187_c78 bl[78] br[78] wl[187] vdd gnd cell_6t
Xbit_r188_c78 bl[78] br[78] wl[188] vdd gnd cell_6t
Xbit_r189_c78 bl[78] br[78] wl[189] vdd gnd cell_6t
Xbit_r190_c78 bl[78] br[78] wl[190] vdd gnd cell_6t
Xbit_r191_c78 bl[78] br[78] wl[191] vdd gnd cell_6t
Xbit_r192_c78 bl[78] br[78] wl[192] vdd gnd cell_6t
Xbit_r193_c78 bl[78] br[78] wl[193] vdd gnd cell_6t
Xbit_r194_c78 bl[78] br[78] wl[194] vdd gnd cell_6t
Xbit_r195_c78 bl[78] br[78] wl[195] vdd gnd cell_6t
Xbit_r196_c78 bl[78] br[78] wl[196] vdd gnd cell_6t
Xbit_r197_c78 bl[78] br[78] wl[197] vdd gnd cell_6t
Xbit_r198_c78 bl[78] br[78] wl[198] vdd gnd cell_6t
Xbit_r199_c78 bl[78] br[78] wl[199] vdd gnd cell_6t
Xbit_r200_c78 bl[78] br[78] wl[200] vdd gnd cell_6t
Xbit_r201_c78 bl[78] br[78] wl[201] vdd gnd cell_6t
Xbit_r202_c78 bl[78] br[78] wl[202] vdd gnd cell_6t
Xbit_r203_c78 bl[78] br[78] wl[203] vdd gnd cell_6t
Xbit_r204_c78 bl[78] br[78] wl[204] vdd gnd cell_6t
Xbit_r205_c78 bl[78] br[78] wl[205] vdd gnd cell_6t
Xbit_r206_c78 bl[78] br[78] wl[206] vdd gnd cell_6t
Xbit_r207_c78 bl[78] br[78] wl[207] vdd gnd cell_6t
Xbit_r208_c78 bl[78] br[78] wl[208] vdd gnd cell_6t
Xbit_r209_c78 bl[78] br[78] wl[209] vdd gnd cell_6t
Xbit_r210_c78 bl[78] br[78] wl[210] vdd gnd cell_6t
Xbit_r211_c78 bl[78] br[78] wl[211] vdd gnd cell_6t
Xbit_r212_c78 bl[78] br[78] wl[212] vdd gnd cell_6t
Xbit_r213_c78 bl[78] br[78] wl[213] vdd gnd cell_6t
Xbit_r214_c78 bl[78] br[78] wl[214] vdd gnd cell_6t
Xbit_r215_c78 bl[78] br[78] wl[215] vdd gnd cell_6t
Xbit_r216_c78 bl[78] br[78] wl[216] vdd gnd cell_6t
Xbit_r217_c78 bl[78] br[78] wl[217] vdd gnd cell_6t
Xbit_r218_c78 bl[78] br[78] wl[218] vdd gnd cell_6t
Xbit_r219_c78 bl[78] br[78] wl[219] vdd gnd cell_6t
Xbit_r220_c78 bl[78] br[78] wl[220] vdd gnd cell_6t
Xbit_r221_c78 bl[78] br[78] wl[221] vdd gnd cell_6t
Xbit_r222_c78 bl[78] br[78] wl[222] vdd gnd cell_6t
Xbit_r223_c78 bl[78] br[78] wl[223] vdd gnd cell_6t
Xbit_r224_c78 bl[78] br[78] wl[224] vdd gnd cell_6t
Xbit_r225_c78 bl[78] br[78] wl[225] vdd gnd cell_6t
Xbit_r226_c78 bl[78] br[78] wl[226] vdd gnd cell_6t
Xbit_r227_c78 bl[78] br[78] wl[227] vdd gnd cell_6t
Xbit_r228_c78 bl[78] br[78] wl[228] vdd gnd cell_6t
Xbit_r229_c78 bl[78] br[78] wl[229] vdd gnd cell_6t
Xbit_r230_c78 bl[78] br[78] wl[230] vdd gnd cell_6t
Xbit_r231_c78 bl[78] br[78] wl[231] vdd gnd cell_6t
Xbit_r232_c78 bl[78] br[78] wl[232] vdd gnd cell_6t
Xbit_r233_c78 bl[78] br[78] wl[233] vdd gnd cell_6t
Xbit_r234_c78 bl[78] br[78] wl[234] vdd gnd cell_6t
Xbit_r235_c78 bl[78] br[78] wl[235] vdd gnd cell_6t
Xbit_r236_c78 bl[78] br[78] wl[236] vdd gnd cell_6t
Xbit_r237_c78 bl[78] br[78] wl[237] vdd gnd cell_6t
Xbit_r238_c78 bl[78] br[78] wl[238] vdd gnd cell_6t
Xbit_r239_c78 bl[78] br[78] wl[239] vdd gnd cell_6t
Xbit_r240_c78 bl[78] br[78] wl[240] vdd gnd cell_6t
Xbit_r241_c78 bl[78] br[78] wl[241] vdd gnd cell_6t
Xbit_r242_c78 bl[78] br[78] wl[242] vdd gnd cell_6t
Xbit_r243_c78 bl[78] br[78] wl[243] vdd gnd cell_6t
Xbit_r244_c78 bl[78] br[78] wl[244] vdd gnd cell_6t
Xbit_r245_c78 bl[78] br[78] wl[245] vdd gnd cell_6t
Xbit_r246_c78 bl[78] br[78] wl[246] vdd gnd cell_6t
Xbit_r247_c78 bl[78] br[78] wl[247] vdd gnd cell_6t
Xbit_r248_c78 bl[78] br[78] wl[248] vdd gnd cell_6t
Xbit_r249_c78 bl[78] br[78] wl[249] vdd gnd cell_6t
Xbit_r250_c78 bl[78] br[78] wl[250] vdd gnd cell_6t
Xbit_r251_c78 bl[78] br[78] wl[251] vdd gnd cell_6t
Xbit_r252_c78 bl[78] br[78] wl[252] vdd gnd cell_6t
Xbit_r253_c78 bl[78] br[78] wl[253] vdd gnd cell_6t
Xbit_r254_c78 bl[78] br[78] wl[254] vdd gnd cell_6t
Xbit_r255_c78 bl[78] br[78] wl[255] vdd gnd cell_6t
Xbit_r0_c79 bl[79] br[79] wl[0] vdd gnd cell_6t
Xbit_r1_c79 bl[79] br[79] wl[1] vdd gnd cell_6t
Xbit_r2_c79 bl[79] br[79] wl[2] vdd gnd cell_6t
Xbit_r3_c79 bl[79] br[79] wl[3] vdd gnd cell_6t
Xbit_r4_c79 bl[79] br[79] wl[4] vdd gnd cell_6t
Xbit_r5_c79 bl[79] br[79] wl[5] vdd gnd cell_6t
Xbit_r6_c79 bl[79] br[79] wl[6] vdd gnd cell_6t
Xbit_r7_c79 bl[79] br[79] wl[7] vdd gnd cell_6t
Xbit_r8_c79 bl[79] br[79] wl[8] vdd gnd cell_6t
Xbit_r9_c79 bl[79] br[79] wl[9] vdd gnd cell_6t
Xbit_r10_c79 bl[79] br[79] wl[10] vdd gnd cell_6t
Xbit_r11_c79 bl[79] br[79] wl[11] vdd gnd cell_6t
Xbit_r12_c79 bl[79] br[79] wl[12] vdd gnd cell_6t
Xbit_r13_c79 bl[79] br[79] wl[13] vdd gnd cell_6t
Xbit_r14_c79 bl[79] br[79] wl[14] vdd gnd cell_6t
Xbit_r15_c79 bl[79] br[79] wl[15] vdd gnd cell_6t
Xbit_r16_c79 bl[79] br[79] wl[16] vdd gnd cell_6t
Xbit_r17_c79 bl[79] br[79] wl[17] vdd gnd cell_6t
Xbit_r18_c79 bl[79] br[79] wl[18] vdd gnd cell_6t
Xbit_r19_c79 bl[79] br[79] wl[19] vdd gnd cell_6t
Xbit_r20_c79 bl[79] br[79] wl[20] vdd gnd cell_6t
Xbit_r21_c79 bl[79] br[79] wl[21] vdd gnd cell_6t
Xbit_r22_c79 bl[79] br[79] wl[22] vdd gnd cell_6t
Xbit_r23_c79 bl[79] br[79] wl[23] vdd gnd cell_6t
Xbit_r24_c79 bl[79] br[79] wl[24] vdd gnd cell_6t
Xbit_r25_c79 bl[79] br[79] wl[25] vdd gnd cell_6t
Xbit_r26_c79 bl[79] br[79] wl[26] vdd gnd cell_6t
Xbit_r27_c79 bl[79] br[79] wl[27] vdd gnd cell_6t
Xbit_r28_c79 bl[79] br[79] wl[28] vdd gnd cell_6t
Xbit_r29_c79 bl[79] br[79] wl[29] vdd gnd cell_6t
Xbit_r30_c79 bl[79] br[79] wl[30] vdd gnd cell_6t
Xbit_r31_c79 bl[79] br[79] wl[31] vdd gnd cell_6t
Xbit_r32_c79 bl[79] br[79] wl[32] vdd gnd cell_6t
Xbit_r33_c79 bl[79] br[79] wl[33] vdd gnd cell_6t
Xbit_r34_c79 bl[79] br[79] wl[34] vdd gnd cell_6t
Xbit_r35_c79 bl[79] br[79] wl[35] vdd gnd cell_6t
Xbit_r36_c79 bl[79] br[79] wl[36] vdd gnd cell_6t
Xbit_r37_c79 bl[79] br[79] wl[37] vdd gnd cell_6t
Xbit_r38_c79 bl[79] br[79] wl[38] vdd gnd cell_6t
Xbit_r39_c79 bl[79] br[79] wl[39] vdd gnd cell_6t
Xbit_r40_c79 bl[79] br[79] wl[40] vdd gnd cell_6t
Xbit_r41_c79 bl[79] br[79] wl[41] vdd gnd cell_6t
Xbit_r42_c79 bl[79] br[79] wl[42] vdd gnd cell_6t
Xbit_r43_c79 bl[79] br[79] wl[43] vdd gnd cell_6t
Xbit_r44_c79 bl[79] br[79] wl[44] vdd gnd cell_6t
Xbit_r45_c79 bl[79] br[79] wl[45] vdd gnd cell_6t
Xbit_r46_c79 bl[79] br[79] wl[46] vdd gnd cell_6t
Xbit_r47_c79 bl[79] br[79] wl[47] vdd gnd cell_6t
Xbit_r48_c79 bl[79] br[79] wl[48] vdd gnd cell_6t
Xbit_r49_c79 bl[79] br[79] wl[49] vdd gnd cell_6t
Xbit_r50_c79 bl[79] br[79] wl[50] vdd gnd cell_6t
Xbit_r51_c79 bl[79] br[79] wl[51] vdd gnd cell_6t
Xbit_r52_c79 bl[79] br[79] wl[52] vdd gnd cell_6t
Xbit_r53_c79 bl[79] br[79] wl[53] vdd gnd cell_6t
Xbit_r54_c79 bl[79] br[79] wl[54] vdd gnd cell_6t
Xbit_r55_c79 bl[79] br[79] wl[55] vdd gnd cell_6t
Xbit_r56_c79 bl[79] br[79] wl[56] vdd gnd cell_6t
Xbit_r57_c79 bl[79] br[79] wl[57] vdd gnd cell_6t
Xbit_r58_c79 bl[79] br[79] wl[58] vdd gnd cell_6t
Xbit_r59_c79 bl[79] br[79] wl[59] vdd gnd cell_6t
Xbit_r60_c79 bl[79] br[79] wl[60] vdd gnd cell_6t
Xbit_r61_c79 bl[79] br[79] wl[61] vdd gnd cell_6t
Xbit_r62_c79 bl[79] br[79] wl[62] vdd gnd cell_6t
Xbit_r63_c79 bl[79] br[79] wl[63] vdd gnd cell_6t
Xbit_r64_c79 bl[79] br[79] wl[64] vdd gnd cell_6t
Xbit_r65_c79 bl[79] br[79] wl[65] vdd gnd cell_6t
Xbit_r66_c79 bl[79] br[79] wl[66] vdd gnd cell_6t
Xbit_r67_c79 bl[79] br[79] wl[67] vdd gnd cell_6t
Xbit_r68_c79 bl[79] br[79] wl[68] vdd gnd cell_6t
Xbit_r69_c79 bl[79] br[79] wl[69] vdd gnd cell_6t
Xbit_r70_c79 bl[79] br[79] wl[70] vdd gnd cell_6t
Xbit_r71_c79 bl[79] br[79] wl[71] vdd gnd cell_6t
Xbit_r72_c79 bl[79] br[79] wl[72] vdd gnd cell_6t
Xbit_r73_c79 bl[79] br[79] wl[73] vdd gnd cell_6t
Xbit_r74_c79 bl[79] br[79] wl[74] vdd gnd cell_6t
Xbit_r75_c79 bl[79] br[79] wl[75] vdd gnd cell_6t
Xbit_r76_c79 bl[79] br[79] wl[76] vdd gnd cell_6t
Xbit_r77_c79 bl[79] br[79] wl[77] vdd gnd cell_6t
Xbit_r78_c79 bl[79] br[79] wl[78] vdd gnd cell_6t
Xbit_r79_c79 bl[79] br[79] wl[79] vdd gnd cell_6t
Xbit_r80_c79 bl[79] br[79] wl[80] vdd gnd cell_6t
Xbit_r81_c79 bl[79] br[79] wl[81] vdd gnd cell_6t
Xbit_r82_c79 bl[79] br[79] wl[82] vdd gnd cell_6t
Xbit_r83_c79 bl[79] br[79] wl[83] vdd gnd cell_6t
Xbit_r84_c79 bl[79] br[79] wl[84] vdd gnd cell_6t
Xbit_r85_c79 bl[79] br[79] wl[85] vdd gnd cell_6t
Xbit_r86_c79 bl[79] br[79] wl[86] vdd gnd cell_6t
Xbit_r87_c79 bl[79] br[79] wl[87] vdd gnd cell_6t
Xbit_r88_c79 bl[79] br[79] wl[88] vdd gnd cell_6t
Xbit_r89_c79 bl[79] br[79] wl[89] vdd gnd cell_6t
Xbit_r90_c79 bl[79] br[79] wl[90] vdd gnd cell_6t
Xbit_r91_c79 bl[79] br[79] wl[91] vdd gnd cell_6t
Xbit_r92_c79 bl[79] br[79] wl[92] vdd gnd cell_6t
Xbit_r93_c79 bl[79] br[79] wl[93] vdd gnd cell_6t
Xbit_r94_c79 bl[79] br[79] wl[94] vdd gnd cell_6t
Xbit_r95_c79 bl[79] br[79] wl[95] vdd gnd cell_6t
Xbit_r96_c79 bl[79] br[79] wl[96] vdd gnd cell_6t
Xbit_r97_c79 bl[79] br[79] wl[97] vdd gnd cell_6t
Xbit_r98_c79 bl[79] br[79] wl[98] vdd gnd cell_6t
Xbit_r99_c79 bl[79] br[79] wl[99] vdd gnd cell_6t
Xbit_r100_c79 bl[79] br[79] wl[100] vdd gnd cell_6t
Xbit_r101_c79 bl[79] br[79] wl[101] vdd gnd cell_6t
Xbit_r102_c79 bl[79] br[79] wl[102] vdd gnd cell_6t
Xbit_r103_c79 bl[79] br[79] wl[103] vdd gnd cell_6t
Xbit_r104_c79 bl[79] br[79] wl[104] vdd gnd cell_6t
Xbit_r105_c79 bl[79] br[79] wl[105] vdd gnd cell_6t
Xbit_r106_c79 bl[79] br[79] wl[106] vdd gnd cell_6t
Xbit_r107_c79 bl[79] br[79] wl[107] vdd gnd cell_6t
Xbit_r108_c79 bl[79] br[79] wl[108] vdd gnd cell_6t
Xbit_r109_c79 bl[79] br[79] wl[109] vdd gnd cell_6t
Xbit_r110_c79 bl[79] br[79] wl[110] vdd gnd cell_6t
Xbit_r111_c79 bl[79] br[79] wl[111] vdd gnd cell_6t
Xbit_r112_c79 bl[79] br[79] wl[112] vdd gnd cell_6t
Xbit_r113_c79 bl[79] br[79] wl[113] vdd gnd cell_6t
Xbit_r114_c79 bl[79] br[79] wl[114] vdd gnd cell_6t
Xbit_r115_c79 bl[79] br[79] wl[115] vdd gnd cell_6t
Xbit_r116_c79 bl[79] br[79] wl[116] vdd gnd cell_6t
Xbit_r117_c79 bl[79] br[79] wl[117] vdd gnd cell_6t
Xbit_r118_c79 bl[79] br[79] wl[118] vdd gnd cell_6t
Xbit_r119_c79 bl[79] br[79] wl[119] vdd gnd cell_6t
Xbit_r120_c79 bl[79] br[79] wl[120] vdd gnd cell_6t
Xbit_r121_c79 bl[79] br[79] wl[121] vdd gnd cell_6t
Xbit_r122_c79 bl[79] br[79] wl[122] vdd gnd cell_6t
Xbit_r123_c79 bl[79] br[79] wl[123] vdd gnd cell_6t
Xbit_r124_c79 bl[79] br[79] wl[124] vdd gnd cell_6t
Xbit_r125_c79 bl[79] br[79] wl[125] vdd gnd cell_6t
Xbit_r126_c79 bl[79] br[79] wl[126] vdd gnd cell_6t
Xbit_r127_c79 bl[79] br[79] wl[127] vdd gnd cell_6t
Xbit_r128_c79 bl[79] br[79] wl[128] vdd gnd cell_6t
Xbit_r129_c79 bl[79] br[79] wl[129] vdd gnd cell_6t
Xbit_r130_c79 bl[79] br[79] wl[130] vdd gnd cell_6t
Xbit_r131_c79 bl[79] br[79] wl[131] vdd gnd cell_6t
Xbit_r132_c79 bl[79] br[79] wl[132] vdd gnd cell_6t
Xbit_r133_c79 bl[79] br[79] wl[133] vdd gnd cell_6t
Xbit_r134_c79 bl[79] br[79] wl[134] vdd gnd cell_6t
Xbit_r135_c79 bl[79] br[79] wl[135] vdd gnd cell_6t
Xbit_r136_c79 bl[79] br[79] wl[136] vdd gnd cell_6t
Xbit_r137_c79 bl[79] br[79] wl[137] vdd gnd cell_6t
Xbit_r138_c79 bl[79] br[79] wl[138] vdd gnd cell_6t
Xbit_r139_c79 bl[79] br[79] wl[139] vdd gnd cell_6t
Xbit_r140_c79 bl[79] br[79] wl[140] vdd gnd cell_6t
Xbit_r141_c79 bl[79] br[79] wl[141] vdd gnd cell_6t
Xbit_r142_c79 bl[79] br[79] wl[142] vdd gnd cell_6t
Xbit_r143_c79 bl[79] br[79] wl[143] vdd gnd cell_6t
Xbit_r144_c79 bl[79] br[79] wl[144] vdd gnd cell_6t
Xbit_r145_c79 bl[79] br[79] wl[145] vdd gnd cell_6t
Xbit_r146_c79 bl[79] br[79] wl[146] vdd gnd cell_6t
Xbit_r147_c79 bl[79] br[79] wl[147] vdd gnd cell_6t
Xbit_r148_c79 bl[79] br[79] wl[148] vdd gnd cell_6t
Xbit_r149_c79 bl[79] br[79] wl[149] vdd gnd cell_6t
Xbit_r150_c79 bl[79] br[79] wl[150] vdd gnd cell_6t
Xbit_r151_c79 bl[79] br[79] wl[151] vdd gnd cell_6t
Xbit_r152_c79 bl[79] br[79] wl[152] vdd gnd cell_6t
Xbit_r153_c79 bl[79] br[79] wl[153] vdd gnd cell_6t
Xbit_r154_c79 bl[79] br[79] wl[154] vdd gnd cell_6t
Xbit_r155_c79 bl[79] br[79] wl[155] vdd gnd cell_6t
Xbit_r156_c79 bl[79] br[79] wl[156] vdd gnd cell_6t
Xbit_r157_c79 bl[79] br[79] wl[157] vdd gnd cell_6t
Xbit_r158_c79 bl[79] br[79] wl[158] vdd gnd cell_6t
Xbit_r159_c79 bl[79] br[79] wl[159] vdd gnd cell_6t
Xbit_r160_c79 bl[79] br[79] wl[160] vdd gnd cell_6t
Xbit_r161_c79 bl[79] br[79] wl[161] vdd gnd cell_6t
Xbit_r162_c79 bl[79] br[79] wl[162] vdd gnd cell_6t
Xbit_r163_c79 bl[79] br[79] wl[163] vdd gnd cell_6t
Xbit_r164_c79 bl[79] br[79] wl[164] vdd gnd cell_6t
Xbit_r165_c79 bl[79] br[79] wl[165] vdd gnd cell_6t
Xbit_r166_c79 bl[79] br[79] wl[166] vdd gnd cell_6t
Xbit_r167_c79 bl[79] br[79] wl[167] vdd gnd cell_6t
Xbit_r168_c79 bl[79] br[79] wl[168] vdd gnd cell_6t
Xbit_r169_c79 bl[79] br[79] wl[169] vdd gnd cell_6t
Xbit_r170_c79 bl[79] br[79] wl[170] vdd gnd cell_6t
Xbit_r171_c79 bl[79] br[79] wl[171] vdd gnd cell_6t
Xbit_r172_c79 bl[79] br[79] wl[172] vdd gnd cell_6t
Xbit_r173_c79 bl[79] br[79] wl[173] vdd gnd cell_6t
Xbit_r174_c79 bl[79] br[79] wl[174] vdd gnd cell_6t
Xbit_r175_c79 bl[79] br[79] wl[175] vdd gnd cell_6t
Xbit_r176_c79 bl[79] br[79] wl[176] vdd gnd cell_6t
Xbit_r177_c79 bl[79] br[79] wl[177] vdd gnd cell_6t
Xbit_r178_c79 bl[79] br[79] wl[178] vdd gnd cell_6t
Xbit_r179_c79 bl[79] br[79] wl[179] vdd gnd cell_6t
Xbit_r180_c79 bl[79] br[79] wl[180] vdd gnd cell_6t
Xbit_r181_c79 bl[79] br[79] wl[181] vdd gnd cell_6t
Xbit_r182_c79 bl[79] br[79] wl[182] vdd gnd cell_6t
Xbit_r183_c79 bl[79] br[79] wl[183] vdd gnd cell_6t
Xbit_r184_c79 bl[79] br[79] wl[184] vdd gnd cell_6t
Xbit_r185_c79 bl[79] br[79] wl[185] vdd gnd cell_6t
Xbit_r186_c79 bl[79] br[79] wl[186] vdd gnd cell_6t
Xbit_r187_c79 bl[79] br[79] wl[187] vdd gnd cell_6t
Xbit_r188_c79 bl[79] br[79] wl[188] vdd gnd cell_6t
Xbit_r189_c79 bl[79] br[79] wl[189] vdd gnd cell_6t
Xbit_r190_c79 bl[79] br[79] wl[190] vdd gnd cell_6t
Xbit_r191_c79 bl[79] br[79] wl[191] vdd gnd cell_6t
Xbit_r192_c79 bl[79] br[79] wl[192] vdd gnd cell_6t
Xbit_r193_c79 bl[79] br[79] wl[193] vdd gnd cell_6t
Xbit_r194_c79 bl[79] br[79] wl[194] vdd gnd cell_6t
Xbit_r195_c79 bl[79] br[79] wl[195] vdd gnd cell_6t
Xbit_r196_c79 bl[79] br[79] wl[196] vdd gnd cell_6t
Xbit_r197_c79 bl[79] br[79] wl[197] vdd gnd cell_6t
Xbit_r198_c79 bl[79] br[79] wl[198] vdd gnd cell_6t
Xbit_r199_c79 bl[79] br[79] wl[199] vdd gnd cell_6t
Xbit_r200_c79 bl[79] br[79] wl[200] vdd gnd cell_6t
Xbit_r201_c79 bl[79] br[79] wl[201] vdd gnd cell_6t
Xbit_r202_c79 bl[79] br[79] wl[202] vdd gnd cell_6t
Xbit_r203_c79 bl[79] br[79] wl[203] vdd gnd cell_6t
Xbit_r204_c79 bl[79] br[79] wl[204] vdd gnd cell_6t
Xbit_r205_c79 bl[79] br[79] wl[205] vdd gnd cell_6t
Xbit_r206_c79 bl[79] br[79] wl[206] vdd gnd cell_6t
Xbit_r207_c79 bl[79] br[79] wl[207] vdd gnd cell_6t
Xbit_r208_c79 bl[79] br[79] wl[208] vdd gnd cell_6t
Xbit_r209_c79 bl[79] br[79] wl[209] vdd gnd cell_6t
Xbit_r210_c79 bl[79] br[79] wl[210] vdd gnd cell_6t
Xbit_r211_c79 bl[79] br[79] wl[211] vdd gnd cell_6t
Xbit_r212_c79 bl[79] br[79] wl[212] vdd gnd cell_6t
Xbit_r213_c79 bl[79] br[79] wl[213] vdd gnd cell_6t
Xbit_r214_c79 bl[79] br[79] wl[214] vdd gnd cell_6t
Xbit_r215_c79 bl[79] br[79] wl[215] vdd gnd cell_6t
Xbit_r216_c79 bl[79] br[79] wl[216] vdd gnd cell_6t
Xbit_r217_c79 bl[79] br[79] wl[217] vdd gnd cell_6t
Xbit_r218_c79 bl[79] br[79] wl[218] vdd gnd cell_6t
Xbit_r219_c79 bl[79] br[79] wl[219] vdd gnd cell_6t
Xbit_r220_c79 bl[79] br[79] wl[220] vdd gnd cell_6t
Xbit_r221_c79 bl[79] br[79] wl[221] vdd gnd cell_6t
Xbit_r222_c79 bl[79] br[79] wl[222] vdd gnd cell_6t
Xbit_r223_c79 bl[79] br[79] wl[223] vdd gnd cell_6t
Xbit_r224_c79 bl[79] br[79] wl[224] vdd gnd cell_6t
Xbit_r225_c79 bl[79] br[79] wl[225] vdd gnd cell_6t
Xbit_r226_c79 bl[79] br[79] wl[226] vdd gnd cell_6t
Xbit_r227_c79 bl[79] br[79] wl[227] vdd gnd cell_6t
Xbit_r228_c79 bl[79] br[79] wl[228] vdd gnd cell_6t
Xbit_r229_c79 bl[79] br[79] wl[229] vdd gnd cell_6t
Xbit_r230_c79 bl[79] br[79] wl[230] vdd gnd cell_6t
Xbit_r231_c79 bl[79] br[79] wl[231] vdd gnd cell_6t
Xbit_r232_c79 bl[79] br[79] wl[232] vdd gnd cell_6t
Xbit_r233_c79 bl[79] br[79] wl[233] vdd gnd cell_6t
Xbit_r234_c79 bl[79] br[79] wl[234] vdd gnd cell_6t
Xbit_r235_c79 bl[79] br[79] wl[235] vdd gnd cell_6t
Xbit_r236_c79 bl[79] br[79] wl[236] vdd gnd cell_6t
Xbit_r237_c79 bl[79] br[79] wl[237] vdd gnd cell_6t
Xbit_r238_c79 bl[79] br[79] wl[238] vdd gnd cell_6t
Xbit_r239_c79 bl[79] br[79] wl[239] vdd gnd cell_6t
Xbit_r240_c79 bl[79] br[79] wl[240] vdd gnd cell_6t
Xbit_r241_c79 bl[79] br[79] wl[241] vdd gnd cell_6t
Xbit_r242_c79 bl[79] br[79] wl[242] vdd gnd cell_6t
Xbit_r243_c79 bl[79] br[79] wl[243] vdd gnd cell_6t
Xbit_r244_c79 bl[79] br[79] wl[244] vdd gnd cell_6t
Xbit_r245_c79 bl[79] br[79] wl[245] vdd gnd cell_6t
Xbit_r246_c79 bl[79] br[79] wl[246] vdd gnd cell_6t
Xbit_r247_c79 bl[79] br[79] wl[247] vdd gnd cell_6t
Xbit_r248_c79 bl[79] br[79] wl[248] vdd gnd cell_6t
Xbit_r249_c79 bl[79] br[79] wl[249] vdd gnd cell_6t
Xbit_r250_c79 bl[79] br[79] wl[250] vdd gnd cell_6t
Xbit_r251_c79 bl[79] br[79] wl[251] vdd gnd cell_6t
Xbit_r252_c79 bl[79] br[79] wl[252] vdd gnd cell_6t
Xbit_r253_c79 bl[79] br[79] wl[253] vdd gnd cell_6t
Xbit_r254_c79 bl[79] br[79] wl[254] vdd gnd cell_6t
Xbit_r255_c79 bl[79] br[79] wl[255] vdd gnd cell_6t
Xbit_r0_c80 bl[80] br[80] wl[0] vdd gnd cell_6t
Xbit_r1_c80 bl[80] br[80] wl[1] vdd gnd cell_6t
Xbit_r2_c80 bl[80] br[80] wl[2] vdd gnd cell_6t
Xbit_r3_c80 bl[80] br[80] wl[3] vdd gnd cell_6t
Xbit_r4_c80 bl[80] br[80] wl[4] vdd gnd cell_6t
Xbit_r5_c80 bl[80] br[80] wl[5] vdd gnd cell_6t
Xbit_r6_c80 bl[80] br[80] wl[6] vdd gnd cell_6t
Xbit_r7_c80 bl[80] br[80] wl[7] vdd gnd cell_6t
Xbit_r8_c80 bl[80] br[80] wl[8] vdd gnd cell_6t
Xbit_r9_c80 bl[80] br[80] wl[9] vdd gnd cell_6t
Xbit_r10_c80 bl[80] br[80] wl[10] vdd gnd cell_6t
Xbit_r11_c80 bl[80] br[80] wl[11] vdd gnd cell_6t
Xbit_r12_c80 bl[80] br[80] wl[12] vdd gnd cell_6t
Xbit_r13_c80 bl[80] br[80] wl[13] vdd gnd cell_6t
Xbit_r14_c80 bl[80] br[80] wl[14] vdd gnd cell_6t
Xbit_r15_c80 bl[80] br[80] wl[15] vdd gnd cell_6t
Xbit_r16_c80 bl[80] br[80] wl[16] vdd gnd cell_6t
Xbit_r17_c80 bl[80] br[80] wl[17] vdd gnd cell_6t
Xbit_r18_c80 bl[80] br[80] wl[18] vdd gnd cell_6t
Xbit_r19_c80 bl[80] br[80] wl[19] vdd gnd cell_6t
Xbit_r20_c80 bl[80] br[80] wl[20] vdd gnd cell_6t
Xbit_r21_c80 bl[80] br[80] wl[21] vdd gnd cell_6t
Xbit_r22_c80 bl[80] br[80] wl[22] vdd gnd cell_6t
Xbit_r23_c80 bl[80] br[80] wl[23] vdd gnd cell_6t
Xbit_r24_c80 bl[80] br[80] wl[24] vdd gnd cell_6t
Xbit_r25_c80 bl[80] br[80] wl[25] vdd gnd cell_6t
Xbit_r26_c80 bl[80] br[80] wl[26] vdd gnd cell_6t
Xbit_r27_c80 bl[80] br[80] wl[27] vdd gnd cell_6t
Xbit_r28_c80 bl[80] br[80] wl[28] vdd gnd cell_6t
Xbit_r29_c80 bl[80] br[80] wl[29] vdd gnd cell_6t
Xbit_r30_c80 bl[80] br[80] wl[30] vdd gnd cell_6t
Xbit_r31_c80 bl[80] br[80] wl[31] vdd gnd cell_6t
Xbit_r32_c80 bl[80] br[80] wl[32] vdd gnd cell_6t
Xbit_r33_c80 bl[80] br[80] wl[33] vdd gnd cell_6t
Xbit_r34_c80 bl[80] br[80] wl[34] vdd gnd cell_6t
Xbit_r35_c80 bl[80] br[80] wl[35] vdd gnd cell_6t
Xbit_r36_c80 bl[80] br[80] wl[36] vdd gnd cell_6t
Xbit_r37_c80 bl[80] br[80] wl[37] vdd gnd cell_6t
Xbit_r38_c80 bl[80] br[80] wl[38] vdd gnd cell_6t
Xbit_r39_c80 bl[80] br[80] wl[39] vdd gnd cell_6t
Xbit_r40_c80 bl[80] br[80] wl[40] vdd gnd cell_6t
Xbit_r41_c80 bl[80] br[80] wl[41] vdd gnd cell_6t
Xbit_r42_c80 bl[80] br[80] wl[42] vdd gnd cell_6t
Xbit_r43_c80 bl[80] br[80] wl[43] vdd gnd cell_6t
Xbit_r44_c80 bl[80] br[80] wl[44] vdd gnd cell_6t
Xbit_r45_c80 bl[80] br[80] wl[45] vdd gnd cell_6t
Xbit_r46_c80 bl[80] br[80] wl[46] vdd gnd cell_6t
Xbit_r47_c80 bl[80] br[80] wl[47] vdd gnd cell_6t
Xbit_r48_c80 bl[80] br[80] wl[48] vdd gnd cell_6t
Xbit_r49_c80 bl[80] br[80] wl[49] vdd gnd cell_6t
Xbit_r50_c80 bl[80] br[80] wl[50] vdd gnd cell_6t
Xbit_r51_c80 bl[80] br[80] wl[51] vdd gnd cell_6t
Xbit_r52_c80 bl[80] br[80] wl[52] vdd gnd cell_6t
Xbit_r53_c80 bl[80] br[80] wl[53] vdd gnd cell_6t
Xbit_r54_c80 bl[80] br[80] wl[54] vdd gnd cell_6t
Xbit_r55_c80 bl[80] br[80] wl[55] vdd gnd cell_6t
Xbit_r56_c80 bl[80] br[80] wl[56] vdd gnd cell_6t
Xbit_r57_c80 bl[80] br[80] wl[57] vdd gnd cell_6t
Xbit_r58_c80 bl[80] br[80] wl[58] vdd gnd cell_6t
Xbit_r59_c80 bl[80] br[80] wl[59] vdd gnd cell_6t
Xbit_r60_c80 bl[80] br[80] wl[60] vdd gnd cell_6t
Xbit_r61_c80 bl[80] br[80] wl[61] vdd gnd cell_6t
Xbit_r62_c80 bl[80] br[80] wl[62] vdd gnd cell_6t
Xbit_r63_c80 bl[80] br[80] wl[63] vdd gnd cell_6t
Xbit_r64_c80 bl[80] br[80] wl[64] vdd gnd cell_6t
Xbit_r65_c80 bl[80] br[80] wl[65] vdd gnd cell_6t
Xbit_r66_c80 bl[80] br[80] wl[66] vdd gnd cell_6t
Xbit_r67_c80 bl[80] br[80] wl[67] vdd gnd cell_6t
Xbit_r68_c80 bl[80] br[80] wl[68] vdd gnd cell_6t
Xbit_r69_c80 bl[80] br[80] wl[69] vdd gnd cell_6t
Xbit_r70_c80 bl[80] br[80] wl[70] vdd gnd cell_6t
Xbit_r71_c80 bl[80] br[80] wl[71] vdd gnd cell_6t
Xbit_r72_c80 bl[80] br[80] wl[72] vdd gnd cell_6t
Xbit_r73_c80 bl[80] br[80] wl[73] vdd gnd cell_6t
Xbit_r74_c80 bl[80] br[80] wl[74] vdd gnd cell_6t
Xbit_r75_c80 bl[80] br[80] wl[75] vdd gnd cell_6t
Xbit_r76_c80 bl[80] br[80] wl[76] vdd gnd cell_6t
Xbit_r77_c80 bl[80] br[80] wl[77] vdd gnd cell_6t
Xbit_r78_c80 bl[80] br[80] wl[78] vdd gnd cell_6t
Xbit_r79_c80 bl[80] br[80] wl[79] vdd gnd cell_6t
Xbit_r80_c80 bl[80] br[80] wl[80] vdd gnd cell_6t
Xbit_r81_c80 bl[80] br[80] wl[81] vdd gnd cell_6t
Xbit_r82_c80 bl[80] br[80] wl[82] vdd gnd cell_6t
Xbit_r83_c80 bl[80] br[80] wl[83] vdd gnd cell_6t
Xbit_r84_c80 bl[80] br[80] wl[84] vdd gnd cell_6t
Xbit_r85_c80 bl[80] br[80] wl[85] vdd gnd cell_6t
Xbit_r86_c80 bl[80] br[80] wl[86] vdd gnd cell_6t
Xbit_r87_c80 bl[80] br[80] wl[87] vdd gnd cell_6t
Xbit_r88_c80 bl[80] br[80] wl[88] vdd gnd cell_6t
Xbit_r89_c80 bl[80] br[80] wl[89] vdd gnd cell_6t
Xbit_r90_c80 bl[80] br[80] wl[90] vdd gnd cell_6t
Xbit_r91_c80 bl[80] br[80] wl[91] vdd gnd cell_6t
Xbit_r92_c80 bl[80] br[80] wl[92] vdd gnd cell_6t
Xbit_r93_c80 bl[80] br[80] wl[93] vdd gnd cell_6t
Xbit_r94_c80 bl[80] br[80] wl[94] vdd gnd cell_6t
Xbit_r95_c80 bl[80] br[80] wl[95] vdd gnd cell_6t
Xbit_r96_c80 bl[80] br[80] wl[96] vdd gnd cell_6t
Xbit_r97_c80 bl[80] br[80] wl[97] vdd gnd cell_6t
Xbit_r98_c80 bl[80] br[80] wl[98] vdd gnd cell_6t
Xbit_r99_c80 bl[80] br[80] wl[99] vdd gnd cell_6t
Xbit_r100_c80 bl[80] br[80] wl[100] vdd gnd cell_6t
Xbit_r101_c80 bl[80] br[80] wl[101] vdd gnd cell_6t
Xbit_r102_c80 bl[80] br[80] wl[102] vdd gnd cell_6t
Xbit_r103_c80 bl[80] br[80] wl[103] vdd gnd cell_6t
Xbit_r104_c80 bl[80] br[80] wl[104] vdd gnd cell_6t
Xbit_r105_c80 bl[80] br[80] wl[105] vdd gnd cell_6t
Xbit_r106_c80 bl[80] br[80] wl[106] vdd gnd cell_6t
Xbit_r107_c80 bl[80] br[80] wl[107] vdd gnd cell_6t
Xbit_r108_c80 bl[80] br[80] wl[108] vdd gnd cell_6t
Xbit_r109_c80 bl[80] br[80] wl[109] vdd gnd cell_6t
Xbit_r110_c80 bl[80] br[80] wl[110] vdd gnd cell_6t
Xbit_r111_c80 bl[80] br[80] wl[111] vdd gnd cell_6t
Xbit_r112_c80 bl[80] br[80] wl[112] vdd gnd cell_6t
Xbit_r113_c80 bl[80] br[80] wl[113] vdd gnd cell_6t
Xbit_r114_c80 bl[80] br[80] wl[114] vdd gnd cell_6t
Xbit_r115_c80 bl[80] br[80] wl[115] vdd gnd cell_6t
Xbit_r116_c80 bl[80] br[80] wl[116] vdd gnd cell_6t
Xbit_r117_c80 bl[80] br[80] wl[117] vdd gnd cell_6t
Xbit_r118_c80 bl[80] br[80] wl[118] vdd gnd cell_6t
Xbit_r119_c80 bl[80] br[80] wl[119] vdd gnd cell_6t
Xbit_r120_c80 bl[80] br[80] wl[120] vdd gnd cell_6t
Xbit_r121_c80 bl[80] br[80] wl[121] vdd gnd cell_6t
Xbit_r122_c80 bl[80] br[80] wl[122] vdd gnd cell_6t
Xbit_r123_c80 bl[80] br[80] wl[123] vdd gnd cell_6t
Xbit_r124_c80 bl[80] br[80] wl[124] vdd gnd cell_6t
Xbit_r125_c80 bl[80] br[80] wl[125] vdd gnd cell_6t
Xbit_r126_c80 bl[80] br[80] wl[126] vdd gnd cell_6t
Xbit_r127_c80 bl[80] br[80] wl[127] vdd gnd cell_6t
Xbit_r128_c80 bl[80] br[80] wl[128] vdd gnd cell_6t
Xbit_r129_c80 bl[80] br[80] wl[129] vdd gnd cell_6t
Xbit_r130_c80 bl[80] br[80] wl[130] vdd gnd cell_6t
Xbit_r131_c80 bl[80] br[80] wl[131] vdd gnd cell_6t
Xbit_r132_c80 bl[80] br[80] wl[132] vdd gnd cell_6t
Xbit_r133_c80 bl[80] br[80] wl[133] vdd gnd cell_6t
Xbit_r134_c80 bl[80] br[80] wl[134] vdd gnd cell_6t
Xbit_r135_c80 bl[80] br[80] wl[135] vdd gnd cell_6t
Xbit_r136_c80 bl[80] br[80] wl[136] vdd gnd cell_6t
Xbit_r137_c80 bl[80] br[80] wl[137] vdd gnd cell_6t
Xbit_r138_c80 bl[80] br[80] wl[138] vdd gnd cell_6t
Xbit_r139_c80 bl[80] br[80] wl[139] vdd gnd cell_6t
Xbit_r140_c80 bl[80] br[80] wl[140] vdd gnd cell_6t
Xbit_r141_c80 bl[80] br[80] wl[141] vdd gnd cell_6t
Xbit_r142_c80 bl[80] br[80] wl[142] vdd gnd cell_6t
Xbit_r143_c80 bl[80] br[80] wl[143] vdd gnd cell_6t
Xbit_r144_c80 bl[80] br[80] wl[144] vdd gnd cell_6t
Xbit_r145_c80 bl[80] br[80] wl[145] vdd gnd cell_6t
Xbit_r146_c80 bl[80] br[80] wl[146] vdd gnd cell_6t
Xbit_r147_c80 bl[80] br[80] wl[147] vdd gnd cell_6t
Xbit_r148_c80 bl[80] br[80] wl[148] vdd gnd cell_6t
Xbit_r149_c80 bl[80] br[80] wl[149] vdd gnd cell_6t
Xbit_r150_c80 bl[80] br[80] wl[150] vdd gnd cell_6t
Xbit_r151_c80 bl[80] br[80] wl[151] vdd gnd cell_6t
Xbit_r152_c80 bl[80] br[80] wl[152] vdd gnd cell_6t
Xbit_r153_c80 bl[80] br[80] wl[153] vdd gnd cell_6t
Xbit_r154_c80 bl[80] br[80] wl[154] vdd gnd cell_6t
Xbit_r155_c80 bl[80] br[80] wl[155] vdd gnd cell_6t
Xbit_r156_c80 bl[80] br[80] wl[156] vdd gnd cell_6t
Xbit_r157_c80 bl[80] br[80] wl[157] vdd gnd cell_6t
Xbit_r158_c80 bl[80] br[80] wl[158] vdd gnd cell_6t
Xbit_r159_c80 bl[80] br[80] wl[159] vdd gnd cell_6t
Xbit_r160_c80 bl[80] br[80] wl[160] vdd gnd cell_6t
Xbit_r161_c80 bl[80] br[80] wl[161] vdd gnd cell_6t
Xbit_r162_c80 bl[80] br[80] wl[162] vdd gnd cell_6t
Xbit_r163_c80 bl[80] br[80] wl[163] vdd gnd cell_6t
Xbit_r164_c80 bl[80] br[80] wl[164] vdd gnd cell_6t
Xbit_r165_c80 bl[80] br[80] wl[165] vdd gnd cell_6t
Xbit_r166_c80 bl[80] br[80] wl[166] vdd gnd cell_6t
Xbit_r167_c80 bl[80] br[80] wl[167] vdd gnd cell_6t
Xbit_r168_c80 bl[80] br[80] wl[168] vdd gnd cell_6t
Xbit_r169_c80 bl[80] br[80] wl[169] vdd gnd cell_6t
Xbit_r170_c80 bl[80] br[80] wl[170] vdd gnd cell_6t
Xbit_r171_c80 bl[80] br[80] wl[171] vdd gnd cell_6t
Xbit_r172_c80 bl[80] br[80] wl[172] vdd gnd cell_6t
Xbit_r173_c80 bl[80] br[80] wl[173] vdd gnd cell_6t
Xbit_r174_c80 bl[80] br[80] wl[174] vdd gnd cell_6t
Xbit_r175_c80 bl[80] br[80] wl[175] vdd gnd cell_6t
Xbit_r176_c80 bl[80] br[80] wl[176] vdd gnd cell_6t
Xbit_r177_c80 bl[80] br[80] wl[177] vdd gnd cell_6t
Xbit_r178_c80 bl[80] br[80] wl[178] vdd gnd cell_6t
Xbit_r179_c80 bl[80] br[80] wl[179] vdd gnd cell_6t
Xbit_r180_c80 bl[80] br[80] wl[180] vdd gnd cell_6t
Xbit_r181_c80 bl[80] br[80] wl[181] vdd gnd cell_6t
Xbit_r182_c80 bl[80] br[80] wl[182] vdd gnd cell_6t
Xbit_r183_c80 bl[80] br[80] wl[183] vdd gnd cell_6t
Xbit_r184_c80 bl[80] br[80] wl[184] vdd gnd cell_6t
Xbit_r185_c80 bl[80] br[80] wl[185] vdd gnd cell_6t
Xbit_r186_c80 bl[80] br[80] wl[186] vdd gnd cell_6t
Xbit_r187_c80 bl[80] br[80] wl[187] vdd gnd cell_6t
Xbit_r188_c80 bl[80] br[80] wl[188] vdd gnd cell_6t
Xbit_r189_c80 bl[80] br[80] wl[189] vdd gnd cell_6t
Xbit_r190_c80 bl[80] br[80] wl[190] vdd gnd cell_6t
Xbit_r191_c80 bl[80] br[80] wl[191] vdd gnd cell_6t
Xbit_r192_c80 bl[80] br[80] wl[192] vdd gnd cell_6t
Xbit_r193_c80 bl[80] br[80] wl[193] vdd gnd cell_6t
Xbit_r194_c80 bl[80] br[80] wl[194] vdd gnd cell_6t
Xbit_r195_c80 bl[80] br[80] wl[195] vdd gnd cell_6t
Xbit_r196_c80 bl[80] br[80] wl[196] vdd gnd cell_6t
Xbit_r197_c80 bl[80] br[80] wl[197] vdd gnd cell_6t
Xbit_r198_c80 bl[80] br[80] wl[198] vdd gnd cell_6t
Xbit_r199_c80 bl[80] br[80] wl[199] vdd gnd cell_6t
Xbit_r200_c80 bl[80] br[80] wl[200] vdd gnd cell_6t
Xbit_r201_c80 bl[80] br[80] wl[201] vdd gnd cell_6t
Xbit_r202_c80 bl[80] br[80] wl[202] vdd gnd cell_6t
Xbit_r203_c80 bl[80] br[80] wl[203] vdd gnd cell_6t
Xbit_r204_c80 bl[80] br[80] wl[204] vdd gnd cell_6t
Xbit_r205_c80 bl[80] br[80] wl[205] vdd gnd cell_6t
Xbit_r206_c80 bl[80] br[80] wl[206] vdd gnd cell_6t
Xbit_r207_c80 bl[80] br[80] wl[207] vdd gnd cell_6t
Xbit_r208_c80 bl[80] br[80] wl[208] vdd gnd cell_6t
Xbit_r209_c80 bl[80] br[80] wl[209] vdd gnd cell_6t
Xbit_r210_c80 bl[80] br[80] wl[210] vdd gnd cell_6t
Xbit_r211_c80 bl[80] br[80] wl[211] vdd gnd cell_6t
Xbit_r212_c80 bl[80] br[80] wl[212] vdd gnd cell_6t
Xbit_r213_c80 bl[80] br[80] wl[213] vdd gnd cell_6t
Xbit_r214_c80 bl[80] br[80] wl[214] vdd gnd cell_6t
Xbit_r215_c80 bl[80] br[80] wl[215] vdd gnd cell_6t
Xbit_r216_c80 bl[80] br[80] wl[216] vdd gnd cell_6t
Xbit_r217_c80 bl[80] br[80] wl[217] vdd gnd cell_6t
Xbit_r218_c80 bl[80] br[80] wl[218] vdd gnd cell_6t
Xbit_r219_c80 bl[80] br[80] wl[219] vdd gnd cell_6t
Xbit_r220_c80 bl[80] br[80] wl[220] vdd gnd cell_6t
Xbit_r221_c80 bl[80] br[80] wl[221] vdd gnd cell_6t
Xbit_r222_c80 bl[80] br[80] wl[222] vdd gnd cell_6t
Xbit_r223_c80 bl[80] br[80] wl[223] vdd gnd cell_6t
Xbit_r224_c80 bl[80] br[80] wl[224] vdd gnd cell_6t
Xbit_r225_c80 bl[80] br[80] wl[225] vdd gnd cell_6t
Xbit_r226_c80 bl[80] br[80] wl[226] vdd gnd cell_6t
Xbit_r227_c80 bl[80] br[80] wl[227] vdd gnd cell_6t
Xbit_r228_c80 bl[80] br[80] wl[228] vdd gnd cell_6t
Xbit_r229_c80 bl[80] br[80] wl[229] vdd gnd cell_6t
Xbit_r230_c80 bl[80] br[80] wl[230] vdd gnd cell_6t
Xbit_r231_c80 bl[80] br[80] wl[231] vdd gnd cell_6t
Xbit_r232_c80 bl[80] br[80] wl[232] vdd gnd cell_6t
Xbit_r233_c80 bl[80] br[80] wl[233] vdd gnd cell_6t
Xbit_r234_c80 bl[80] br[80] wl[234] vdd gnd cell_6t
Xbit_r235_c80 bl[80] br[80] wl[235] vdd gnd cell_6t
Xbit_r236_c80 bl[80] br[80] wl[236] vdd gnd cell_6t
Xbit_r237_c80 bl[80] br[80] wl[237] vdd gnd cell_6t
Xbit_r238_c80 bl[80] br[80] wl[238] vdd gnd cell_6t
Xbit_r239_c80 bl[80] br[80] wl[239] vdd gnd cell_6t
Xbit_r240_c80 bl[80] br[80] wl[240] vdd gnd cell_6t
Xbit_r241_c80 bl[80] br[80] wl[241] vdd gnd cell_6t
Xbit_r242_c80 bl[80] br[80] wl[242] vdd gnd cell_6t
Xbit_r243_c80 bl[80] br[80] wl[243] vdd gnd cell_6t
Xbit_r244_c80 bl[80] br[80] wl[244] vdd gnd cell_6t
Xbit_r245_c80 bl[80] br[80] wl[245] vdd gnd cell_6t
Xbit_r246_c80 bl[80] br[80] wl[246] vdd gnd cell_6t
Xbit_r247_c80 bl[80] br[80] wl[247] vdd gnd cell_6t
Xbit_r248_c80 bl[80] br[80] wl[248] vdd gnd cell_6t
Xbit_r249_c80 bl[80] br[80] wl[249] vdd gnd cell_6t
Xbit_r250_c80 bl[80] br[80] wl[250] vdd gnd cell_6t
Xbit_r251_c80 bl[80] br[80] wl[251] vdd gnd cell_6t
Xbit_r252_c80 bl[80] br[80] wl[252] vdd gnd cell_6t
Xbit_r253_c80 bl[80] br[80] wl[253] vdd gnd cell_6t
Xbit_r254_c80 bl[80] br[80] wl[254] vdd gnd cell_6t
Xbit_r255_c80 bl[80] br[80] wl[255] vdd gnd cell_6t
Xbit_r0_c81 bl[81] br[81] wl[0] vdd gnd cell_6t
Xbit_r1_c81 bl[81] br[81] wl[1] vdd gnd cell_6t
Xbit_r2_c81 bl[81] br[81] wl[2] vdd gnd cell_6t
Xbit_r3_c81 bl[81] br[81] wl[3] vdd gnd cell_6t
Xbit_r4_c81 bl[81] br[81] wl[4] vdd gnd cell_6t
Xbit_r5_c81 bl[81] br[81] wl[5] vdd gnd cell_6t
Xbit_r6_c81 bl[81] br[81] wl[6] vdd gnd cell_6t
Xbit_r7_c81 bl[81] br[81] wl[7] vdd gnd cell_6t
Xbit_r8_c81 bl[81] br[81] wl[8] vdd gnd cell_6t
Xbit_r9_c81 bl[81] br[81] wl[9] vdd gnd cell_6t
Xbit_r10_c81 bl[81] br[81] wl[10] vdd gnd cell_6t
Xbit_r11_c81 bl[81] br[81] wl[11] vdd gnd cell_6t
Xbit_r12_c81 bl[81] br[81] wl[12] vdd gnd cell_6t
Xbit_r13_c81 bl[81] br[81] wl[13] vdd gnd cell_6t
Xbit_r14_c81 bl[81] br[81] wl[14] vdd gnd cell_6t
Xbit_r15_c81 bl[81] br[81] wl[15] vdd gnd cell_6t
Xbit_r16_c81 bl[81] br[81] wl[16] vdd gnd cell_6t
Xbit_r17_c81 bl[81] br[81] wl[17] vdd gnd cell_6t
Xbit_r18_c81 bl[81] br[81] wl[18] vdd gnd cell_6t
Xbit_r19_c81 bl[81] br[81] wl[19] vdd gnd cell_6t
Xbit_r20_c81 bl[81] br[81] wl[20] vdd gnd cell_6t
Xbit_r21_c81 bl[81] br[81] wl[21] vdd gnd cell_6t
Xbit_r22_c81 bl[81] br[81] wl[22] vdd gnd cell_6t
Xbit_r23_c81 bl[81] br[81] wl[23] vdd gnd cell_6t
Xbit_r24_c81 bl[81] br[81] wl[24] vdd gnd cell_6t
Xbit_r25_c81 bl[81] br[81] wl[25] vdd gnd cell_6t
Xbit_r26_c81 bl[81] br[81] wl[26] vdd gnd cell_6t
Xbit_r27_c81 bl[81] br[81] wl[27] vdd gnd cell_6t
Xbit_r28_c81 bl[81] br[81] wl[28] vdd gnd cell_6t
Xbit_r29_c81 bl[81] br[81] wl[29] vdd gnd cell_6t
Xbit_r30_c81 bl[81] br[81] wl[30] vdd gnd cell_6t
Xbit_r31_c81 bl[81] br[81] wl[31] vdd gnd cell_6t
Xbit_r32_c81 bl[81] br[81] wl[32] vdd gnd cell_6t
Xbit_r33_c81 bl[81] br[81] wl[33] vdd gnd cell_6t
Xbit_r34_c81 bl[81] br[81] wl[34] vdd gnd cell_6t
Xbit_r35_c81 bl[81] br[81] wl[35] vdd gnd cell_6t
Xbit_r36_c81 bl[81] br[81] wl[36] vdd gnd cell_6t
Xbit_r37_c81 bl[81] br[81] wl[37] vdd gnd cell_6t
Xbit_r38_c81 bl[81] br[81] wl[38] vdd gnd cell_6t
Xbit_r39_c81 bl[81] br[81] wl[39] vdd gnd cell_6t
Xbit_r40_c81 bl[81] br[81] wl[40] vdd gnd cell_6t
Xbit_r41_c81 bl[81] br[81] wl[41] vdd gnd cell_6t
Xbit_r42_c81 bl[81] br[81] wl[42] vdd gnd cell_6t
Xbit_r43_c81 bl[81] br[81] wl[43] vdd gnd cell_6t
Xbit_r44_c81 bl[81] br[81] wl[44] vdd gnd cell_6t
Xbit_r45_c81 bl[81] br[81] wl[45] vdd gnd cell_6t
Xbit_r46_c81 bl[81] br[81] wl[46] vdd gnd cell_6t
Xbit_r47_c81 bl[81] br[81] wl[47] vdd gnd cell_6t
Xbit_r48_c81 bl[81] br[81] wl[48] vdd gnd cell_6t
Xbit_r49_c81 bl[81] br[81] wl[49] vdd gnd cell_6t
Xbit_r50_c81 bl[81] br[81] wl[50] vdd gnd cell_6t
Xbit_r51_c81 bl[81] br[81] wl[51] vdd gnd cell_6t
Xbit_r52_c81 bl[81] br[81] wl[52] vdd gnd cell_6t
Xbit_r53_c81 bl[81] br[81] wl[53] vdd gnd cell_6t
Xbit_r54_c81 bl[81] br[81] wl[54] vdd gnd cell_6t
Xbit_r55_c81 bl[81] br[81] wl[55] vdd gnd cell_6t
Xbit_r56_c81 bl[81] br[81] wl[56] vdd gnd cell_6t
Xbit_r57_c81 bl[81] br[81] wl[57] vdd gnd cell_6t
Xbit_r58_c81 bl[81] br[81] wl[58] vdd gnd cell_6t
Xbit_r59_c81 bl[81] br[81] wl[59] vdd gnd cell_6t
Xbit_r60_c81 bl[81] br[81] wl[60] vdd gnd cell_6t
Xbit_r61_c81 bl[81] br[81] wl[61] vdd gnd cell_6t
Xbit_r62_c81 bl[81] br[81] wl[62] vdd gnd cell_6t
Xbit_r63_c81 bl[81] br[81] wl[63] vdd gnd cell_6t
Xbit_r64_c81 bl[81] br[81] wl[64] vdd gnd cell_6t
Xbit_r65_c81 bl[81] br[81] wl[65] vdd gnd cell_6t
Xbit_r66_c81 bl[81] br[81] wl[66] vdd gnd cell_6t
Xbit_r67_c81 bl[81] br[81] wl[67] vdd gnd cell_6t
Xbit_r68_c81 bl[81] br[81] wl[68] vdd gnd cell_6t
Xbit_r69_c81 bl[81] br[81] wl[69] vdd gnd cell_6t
Xbit_r70_c81 bl[81] br[81] wl[70] vdd gnd cell_6t
Xbit_r71_c81 bl[81] br[81] wl[71] vdd gnd cell_6t
Xbit_r72_c81 bl[81] br[81] wl[72] vdd gnd cell_6t
Xbit_r73_c81 bl[81] br[81] wl[73] vdd gnd cell_6t
Xbit_r74_c81 bl[81] br[81] wl[74] vdd gnd cell_6t
Xbit_r75_c81 bl[81] br[81] wl[75] vdd gnd cell_6t
Xbit_r76_c81 bl[81] br[81] wl[76] vdd gnd cell_6t
Xbit_r77_c81 bl[81] br[81] wl[77] vdd gnd cell_6t
Xbit_r78_c81 bl[81] br[81] wl[78] vdd gnd cell_6t
Xbit_r79_c81 bl[81] br[81] wl[79] vdd gnd cell_6t
Xbit_r80_c81 bl[81] br[81] wl[80] vdd gnd cell_6t
Xbit_r81_c81 bl[81] br[81] wl[81] vdd gnd cell_6t
Xbit_r82_c81 bl[81] br[81] wl[82] vdd gnd cell_6t
Xbit_r83_c81 bl[81] br[81] wl[83] vdd gnd cell_6t
Xbit_r84_c81 bl[81] br[81] wl[84] vdd gnd cell_6t
Xbit_r85_c81 bl[81] br[81] wl[85] vdd gnd cell_6t
Xbit_r86_c81 bl[81] br[81] wl[86] vdd gnd cell_6t
Xbit_r87_c81 bl[81] br[81] wl[87] vdd gnd cell_6t
Xbit_r88_c81 bl[81] br[81] wl[88] vdd gnd cell_6t
Xbit_r89_c81 bl[81] br[81] wl[89] vdd gnd cell_6t
Xbit_r90_c81 bl[81] br[81] wl[90] vdd gnd cell_6t
Xbit_r91_c81 bl[81] br[81] wl[91] vdd gnd cell_6t
Xbit_r92_c81 bl[81] br[81] wl[92] vdd gnd cell_6t
Xbit_r93_c81 bl[81] br[81] wl[93] vdd gnd cell_6t
Xbit_r94_c81 bl[81] br[81] wl[94] vdd gnd cell_6t
Xbit_r95_c81 bl[81] br[81] wl[95] vdd gnd cell_6t
Xbit_r96_c81 bl[81] br[81] wl[96] vdd gnd cell_6t
Xbit_r97_c81 bl[81] br[81] wl[97] vdd gnd cell_6t
Xbit_r98_c81 bl[81] br[81] wl[98] vdd gnd cell_6t
Xbit_r99_c81 bl[81] br[81] wl[99] vdd gnd cell_6t
Xbit_r100_c81 bl[81] br[81] wl[100] vdd gnd cell_6t
Xbit_r101_c81 bl[81] br[81] wl[101] vdd gnd cell_6t
Xbit_r102_c81 bl[81] br[81] wl[102] vdd gnd cell_6t
Xbit_r103_c81 bl[81] br[81] wl[103] vdd gnd cell_6t
Xbit_r104_c81 bl[81] br[81] wl[104] vdd gnd cell_6t
Xbit_r105_c81 bl[81] br[81] wl[105] vdd gnd cell_6t
Xbit_r106_c81 bl[81] br[81] wl[106] vdd gnd cell_6t
Xbit_r107_c81 bl[81] br[81] wl[107] vdd gnd cell_6t
Xbit_r108_c81 bl[81] br[81] wl[108] vdd gnd cell_6t
Xbit_r109_c81 bl[81] br[81] wl[109] vdd gnd cell_6t
Xbit_r110_c81 bl[81] br[81] wl[110] vdd gnd cell_6t
Xbit_r111_c81 bl[81] br[81] wl[111] vdd gnd cell_6t
Xbit_r112_c81 bl[81] br[81] wl[112] vdd gnd cell_6t
Xbit_r113_c81 bl[81] br[81] wl[113] vdd gnd cell_6t
Xbit_r114_c81 bl[81] br[81] wl[114] vdd gnd cell_6t
Xbit_r115_c81 bl[81] br[81] wl[115] vdd gnd cell_6t
Xbit_r116_c81 bl[81] br[81] wl[116] vdd gnd cell_6t
Xbit_r117_c81 bl[81] br[81] wl[117] vdd gnd cell_6t
Xbit_r118_c81 bl[81] br[81] wl[118] vdd gnd cell_6t
Xbit_r119_c81 bl[81] br[81] wl[119] vdd gnd cell_6t
Xbit_r120_c81 bl[81] br[81] wl[120] vdd gnd cell_6t
Xbit_r121_c81 bl[81] br[81] wl[121] vdd gnd cell_6t
Xbit_r122_c81 bl[81] br[81] wl[122] vdd gnd cell_6t
Xbit_r123_c81 bl[81] br[81] wl[123] vdd gnd cell_6t
Xbit_r124_c81 bl[81] br[81] wl[124] vdd gnd cell_6t
Xbit_r125_c81 bl[81] br[81] wl[125] vdd gnd cell_6t
Xbit_r126_c81 bl[81] br[81] wl[126] vdd gnd cell_6t
Xbit_r127_c81 bl[81] br[81] wl[127] vdd gnd cell_6t
Xbit_r128_c81 bl[81] br[81] wl[128] vdd gnd cell_6t
Xbit_r129_c81 bl[81] br[81] wl[129] vdd gnd cell_6t
Xbit_r130_c81 bl[81] br[81] wl[130] vdd gnd cell_6t
Xbit_r131_c81 bl[81] br[81] wl[131] vdd gnd cell_6t
Xbit_r132_c81 bl[81] br[81] wl[132] vdd gnd cell_6t
Xbit_r133_c81 bl[81] br[81] wl[133] vdd gnd cell_6t
Xbit_r134_c81 bl[81] br[81] wl[134] vdd gnd cell_6t
Xbit_r135_c81 bl[81] br[81] wl[135] vdd gnd cell_6t
Xbit_r136_c81 bl[81] br[81] wl[136] vdd gnd cell_6t
Xbit_r137_c81 bl[81] br[81] wl[137] vdd gnd cell_6t
Xbit_r138_c81 bl[81] br[81] wl[138] vdd gnd cell_6t
Xbit_r139_c81 bl[81] br[81] wl[139] vdd gnd cell_6t
Xbit_r140_c81 bl[81] br[81] wl[140] vdd gnd cell_6t
Xbit_r141_c81 bl[81] br[81] wl[141] vdd gnd cell_6t
Xbit_r142_c81 bl[81] br[81] wl[142] vdd gnd cell_6t
Xbit_r143_c81 bl[81] br[81] wl[143] vdd gnd cell_6t
Xbit_r144_c81 bl[81] br[81] wl[144] vdd gnd cell_6t
Xbit_r145_c81 bl[81] br[81] wl[145] vdd gnd cell_6t
Xbit_r146_c81 bl[81] br[81] wl[146] vdd gnd cell_6t
Xbit_r147_c81 bl[81] br[81] wl[147] vdd gnd cell_6t
Xbit_r148_c81 bl[81] br[81] wl[148] vdd gnd cell_6t
Xbit_r149_c81 bl[81] br[81] wl[149] vdd gnd cell_6t
Xbit_r150_c81 bl[81] br[81] wl[150] vdd gnd cell_6t
Xbit_r151_c81 bl[81] br[81] wl[151] vdd gnd cell_6t
Xbit_r152_c81 bl[81] br[81] wl[152] vdd gnd cell_6t
Xbit_r153_c81 bl[81] br[81] wl[153] vdd gnd cell_6t
Xbit_r154_c81 bl[81] br[81] wl[154] vdd gnd cell_6t
Xbit_r155_c81 bl[81] br[81] wl[155] vdd gnd cell_6t
Xbit_r156_c81 bl[81] br[81] wl[156] vdd gnd cell_6t
Xbit_r157_c81 bl[81] br[81] wl[157] vdd gnd cell_6t
Xbit_r158_c81 bl[81] br[81] wl[158] vdd gnd cell_6t
Xbit_r159_c81 bl[81] br[81] wl[159] vdd gnd cell_6t
Xbit_r160_c81 bl[81] br[81] wl[160] vdd gnd cell_6t
Xbit_r161_c81 bl[81] br[81] wl[161] vdd gnd cell_6t
Xbit_r162_c81 bl[81] br[81] wl[162] vdd gnd cell_6t
Xbit_r163_c81 bl[81] br[81] wl[163] vdd gnd cell_6t
Xbit_r164_c81 bl[81] br[81] wl[164] vdd gnd cell_6t
Xbit_r165_c81 bl[81] br[81] wl[165] vdd gnd cell_6t
Xbit_r166_c81 bl[81] br[81] wl[166] vdd gnd cell_6t
Xbit_r167_c81 bl[81] br[81] wl[167] vdd gnd cell_6t
Xbit_r168_c81 bl[81] br[81] wl[168] vdd gnd cell_6t
Xbit_r169_c81 bl[81] br[81] wl[169] vdd gnd cell_6t
Xbit_r170_c81 bl[81] br[81] wl[170] vdd gnd cell_6t
Xbit_r171_c81 bl[81] br[81] wl[171] vdd gnd cell_6t
Xbit_r172_c81 bl[81] br[81] wl[172] vdd gnd cell_6t
Xbit_r173_c81 bl[81] br[81] wl[173] vdd gnd cell_6t
Xbit_r174_c81 bl[81] br[81] wl[174] vdd gnd cell_6t
Xbit_r175_c81 bl[81] br[81] wl[175] vdd gnd cell_6t
Xbit_r176_c81 bl[81] br[81] wl[176] vdd gnd cell_6t
Xbit_r177_c81 bl[81] br[81] wl[177] vdd gnd cell_6t
Xbit_r178_c81 bl[81] br[81] wl[178] vdd gnd cell_6t
Xbit_r179_c81 bl[81] br[81] wl[179] vdd gnd cell_6t
Xbit_r180_c81 bl[81] br[81] wl[180] vdd gnd cell_6t
Xbit_r181_c81 bl[81] br[81] wl[181] vdd gnd cell_6t
Xbit_r182_c81 bl[81] br[81] wl[182] vdd gnd cell_6t
Xbit_r183_c81 bl[81] br[81] wl[183] vdd gnd cell_6t
Xbit_r184_c81 bl[81] br[81] wl[184] vdd gnd cell_6t
Xbit_r185_c81 bl[81] br[81] wl[185] vdd gnd cell_6t
Xbit_r186_c81 bl[81] br[81] wl[186] vdd gnd cell_6t
Xbit_r187_c81 bl[81] br[81] wl[187] vdd gnd cell_6t
Xbit_r188_c81 bl[81] br[81] wl[188] vdd gnd cell_6t
Xbit_r189_c81 bl[81] br[81] wl[189] vdd gnd cell_6t
Xbit_r190_c81 bl[81] br[81] wl[190] vdd gnd cell_6t
Xbit_r191_c81 bl[81] br[81] wl[191] vdd gnd cell_6t
Xbit_r192_c81 bl[81] br[81] wl[192] vdd gnd cell_6t
Xbit_r193_c81 bl[81] br[81] wl[193] vdd gnd cell_6t
Xbit_r194_c81 bl[81] br[81] wl[194] vdd gnd cell_6t
Xbit_r195_c81 bl[81] br[81] wl[195] vdd gnd cell_6t
Xbit_r196_c81 bl[81] br[81] wl[196] vdd gnd cell_6t
Xbit_r197_c81 bl[81] br[81] wl[197] vdd gnd cell_6t
Xbit_r198_c81 bl[81] br[81] wl[198] vdd gnd cell_6t
Xbit_r199_c81 bl[81] br[81] wl[199] vdd gnd cell_6t
Xbit_r200_c81 bl[81] br[81] wl[200] vdd gnd cell_6t
Xbit_r201_c81 bl[81] br[81] wl[201] vdd gnd cell_6t
Xbit_r202_c81 bl[81] br[81] wl[202] vdd gnd cell_6t
Xbit_r203_c81 bl[81] br[81] wl[203] vdd gnd cell_6t
Xbit_r204_c81 bl[81] br[81] wl[204] vdd gnd cell_6t
Xbit_r205_c81 bl[81] br[81] wl[205] vdd gnd cell_6t
Xbit_r206_c81 bl[81] br[81] wl[206] vdd gnd cell_6t
Xbit_r207_c81 bl[81] br[81] wl[207] vdd gnd cell_6t
Xbit_r208_c81 bl[81] br[81] wl[208] vdd gnd cell_6t
Xbit_r209_c81 bl[81] br[81] wl[209] vdd gnd cell_6t
Xbit_r210_c81 bl[81] br[81] wl[210] vdd gnd cell_6t
Xbit_r211_c81 bl[81] br[81] wl[211] vdd gnd cell_6t
Xbit_r212_c81 bl[81] br[81] wl[212] vdd gnd cell_6t
Xbit_r213_c81 bl[81] br[81] wl[213] vdd gnd cell_6t
Xbit_r214_c81 bl[81] br[81] wl[214] vdd gnd cell_6t
Xbit_r215_c81 bl[81] br[81] wl[215] vdd gnd cell_6t
Xbit_r216_c81 bl[81] br[81] wl[216] vdd gnd cell_6t
Xbit_r217_c81 bl[81] br[81] wl[217] vdd gnd cell_6t
Xbit_r218_c81 bl[81] br[81] wl[218] vdd gnd cell_6t
Xbit_r219_c81 bl[81] br[81] wl[219] vdd gnd cell_6t
Xbit_r220_c81 bl[81] br[81] wl[220] vdd gnd cell_6t
Xbit_r221_c81 bl[81] br[81] wl[221] vdd gnd cell_6t
Xbit_r222_c81 bl[81] br[81] wl[222] vdd gnd cell_6t
Xbit_r223_c81 bl[81] br[81] wl[223] vdd gnd cell_6t
Xbit_r224_c81 bl[81] br[81] wl[224] vdd gnd cell_6t
Xbit_r225_c81 bl[81] br[81] wl[225] vdd gnd cell_6t
Xbit_r226_c81 bl[81] br[81] wl[226] vdd gnd cell_6t
Xbit_r227_c81 bl[81] br[81] wl[227] vdd gnd cell_6t
Xbit_r228_c81 bl[81] br[81] wl[228] vdd gnd cell_6t
Xbit_r229_c81 bl[81] br[81] wl[229] vdd gnd cell_6t
Xbit_r230_c81 bl[81] br[81] wl[230] vdd gnd cell_6t
Xbit_r231_c81 bl[81] br[81] wl[231] vdd gnd cell_6t
Xbit_r232_c81 bl[81] br[81] wl[232] vdd gnd cell_6t
Xbit_r233_c81 bl[81] br[81] wl[233] vdd gnd cell_6t
Xbit_r234_c81 bl[81] br[81] wl[234] vdd gnd cell_6t
Xbit_r235_c81 bl[81] br[81] wl[235] vdd gnd cell_6t
Xbit_r236_c81 bl[81] br[81] wl[236] vdd gnd cell_6t
Xbit_r237_c81 bl[81] br[81] wl[237] vdd gnd cell_6t
Xbit_r238_c81 bl[81] br[81] wl[238] vdd gnd cell_6t
Xbit_r239_c81 bl[81] br[81] wl[239] vdd gnd cell_6t
Xbit_r240_c81 bl[81] br[81] wl[240] vdd gnd cell_6t
Xbit_r241_c81 bl[81] br[81] wl[241] vdd gnd cell_6t
Xbit_r242_c81 bl[81] br[81] wl[242] vdd gnd cell_6t
Xbit_r243_c81 bl[81] br[81] wl[243] vdd gnd cell_6t
Xbit_r244_c81 bl[81] br[81] wl[244] vdd gnd cell_6t
Xbit_r245_c81 bl[81] br[81] wl[245] vdd gnd cell_6t
Xbit_r246_c81 bl[81] br[81] wl[246] vdd gnd cell_6t
Xbit_r247_c81 bl[81] br[81] wl[247] vdd gnd cell_6t
Xbit_r248_c81 bl[81] br[81] wl[248] vdd gnd cell_6t
Xbit_r249_c81 bl[81] br[81] wl[249] vdd gnd cell_6t
Xbit_r250_c81 bl[81] br[81] wl[250] vdd gnd cell_6t
Xbit_r251_c81 bl[81] br[81] wl[251] vdd gnd cell_6t
Xbit_r252_c81 bl[81] br[81] wl[252] vdd gnd cell_6t
Xbit_r253_c81 bl[81] br[81] wl[253] vdd gnd cell_6t
Xbit_r254_c81 bl[81] br[81] wl[254] vdd gnd cell_6t
Xbit_r255_c81 bl[81] br[81] wl[255] vdd gnd cell_6t
Xbit_r0_c82 bl[82] br[82] wl[0] vdd gnd cell_6t
Xbit_r1_c82 bl[82] br[82] wl[1] vdd gnd cell_6t
Xbit_r2_c82 bl[82] br[82] wl[2] vdd gnd cell_6t
Xbit_r3_c82 bl[82] br[82] wl[3] vdd gnd cell_6t
Xbit_r4_c82 bl[82] br[82] wl[4] vdd gnd cell_6t
Xbit_r5_c82 bl[82] br[82] wl[5] vdd gnd cell_6t
Xbit_r6_c82 bl[82] br[82] wl[6] vdd gnd cell_6t
Xbit_r7_c82 bl[82] br[82] wl[7] vdd gnd cell_6t
Xbit_r8_c82 bl[82] br[82] wl[8] vdd gnd cell_6t
Xbit_r9_c82 bl[82] br[82] wl[9] vdd gnd cell_6t
Xbit_r10_c82 bl[82] br[82] wl[10] vdd gnd cell_6t
Xbit_r11_c82 bl[82] br[82] wl[11] vdd gnd cell_6t
Xbit_r12_c82 bl[82] br[82] wl[12] vdd gnd cell_6t
Xbit_r13_c82 bl[82] br[82] wl[13] vdd gnd cell_6t
Xbit_r14_c82 bl[82] br[82] wl[14] vdd gnd cell_6t
Xbit_r15_c82 bl[82] br[82] wl[15] vdd gnd cell_6t
Xbit_r16_c82 bl[82] br[82] wl[16] vdd gnd cell_6t
Xbit_r17_c82 bl[82] br[82] wl[17] vdd gnd cell_6t
Xbit_r18_c82 bl[82] br[82] wl[18] vdd gnd cell_6t
Xbit_r19_c82 bl[82] br[82] wl[19] vdd gnd cell_6t
Xbit_r20_c82 bl[82] br[82] wl[20] vdd gnd cell_6t
Xbit_r21_c82 bl[82] br[82] wl[21] vdd gnd cell_6t
Xbit_r22_c82 bl[82] br[82] wl[22] vdd gnd cell_6t
Xbit_r23_c82 bl[82] br[82] wl[23] vdd gnd cell_6t
Xbit_r24_c82 bl[82] br[82] wl[24] vdd gnd cell_6t
Xbit_r25_c82 bl[82] br[82] wl[25] vdd gnd cell_6t
Xbit_r26_c82 bl[82] br[82] wl[26] vdd gnd cell_6t
Xbit_r27_c82 bl[82] br[82] wl[27] vdd gnd cell_6t
Xbit_r28_c82 bl[82] br[82] wl[28] vdd gnd cell_6t
Xbit_r29_c82 bl[82] br[82] wl[29] vdd gnd cell_6t
Xbit_r30_c82 bl[82] br[82] wl[30] vdd gnd cell_6t
Xbit_r31_c82 bl[82] br[82] wl[31] vdd gnd cell_6t
Xbit_r32_c82 bl[82] br[82] wl[32] vdd gnd cell_6t
Xbit_r33_c82 bl[82] br[82] wl[33] vdd gnd cell_6t
Xbit_r34_c82 bl[82] br[82] wl[34] vdd gnd cell_6t
Xbit_r35_c82 bl[82] br[82] wl[35] vdd gnd cell_6t
Xbit_r36_c82 bl[82] br[82] wl[36] vdd gnd cell_6t
Xbit_r37_c82 bl[82] br[82] wl[37] vdd gnd cell_6t
Xbit_r38_c82 bl[82] br[82] wl[38] vdd gnd cell_6t
Xbit_r39_c82 bl[82] br[82] wl[39] vdd gnd cell_6t
Xbit_r40_c82 bl[82] br[82] wl[40] vdd gnd cell_6t
Xbit_r41_c82 bl[82] br[82] wl[41] vdd gnd cell_6t
Xbit_r42_c82 bl[82] br[82] wl[42] vdd gnd cell_6t
Xbit_r43_c82 bl[82] br[82] wl[43] vdd gnd cell_6t
Xbit_r44_c82 bl[82] br[82] wl[44] vdd gnd cell_6t
Xbit_r45_c82 bl[82] br[82] wl[45] vdd gnd cell_6t
Xbit_r46_c82 bl[82] br[82] wl[46] vdd gnd cell_6t
Xbit_r47_c82 bl[82] br[82] wl[47] vdd gnd cell_6t
Xbit_r48_c82 bl[82] br[82] wl[48] vdd gnd cell_6t
Xbit_r49_c82 bl[82] br[82] wl[49] vdd gnd cell_6t
Xbit_r50_c82 bl[82] br[82] wl[50] vdd gnd cell_6t
Xbit_r51_c82 bl[82] br[82] wl[51] vdd gnd cell_6t
Xbit_r52_c82 bl[82] br[82] wl[52] vdd gnd cell_6t
Xbit_r53_c82 bl[82] br[82] wl[53] vdd gnd cell_6t
Xbit_r54_c82 bl[82] br[82] wl[54] vdd gnd cell_6t
Xbit_r55_c82 bl[82] br[82] wl[55] vdd gnd cell_6t
Xbit_r56_c82 bl[82] br[82] wl[56] vdd gnd cell_6t
Xbit_r57_c82 bl[82] br[82] wl[57] vdd gnd cell_6t
Xbit_r58_c82 bl[82] br[82] wl[58] vdd gnd cell_6t
Xbit_r59_c82 bl[82] br[82] wl[59] vdd gnd cell_6t
Xbit_r60_c82 bl[82] br[82] wl[60] vdd gnd cell_6t
Xbit_r61_c82 bl[82] br[82] wl[61] vdd gnd cell_6t
Xbit_r62_c82 bl[82] br[82] wl[62] vdd gnd cell_6t
Xbit_r63_c82 bl[82] br[82] wl[63] vdd gnd cell_6t
Xbit_r64_c82 bl[82] br[82] wl[64] vdd gnd cell_6t
Xbit_r65_c82 bl[82] br[82] wl[65] vdd gnd cell_6t
Xbit_r66_c82 bl[82] br[82] wl[66] vdd gnd cell_6t
Xbit_r67_c82 bl[82] br[82] wl[67] vdd gnd cell_6t
Xbit_r68_c82 bl[82] br[82] wl[68] vdd gnd cell_6t
Xbit_r69_c82 bl[82] br[82] wl[69] vdd gnd cell_6t
Xbit_r70_c82 bl[82] br[82] wl[70] vdd gnd cell_6t
Xbit_r71_c82 bl[82] br[82] wl[71] vdd gnd cell_6t
Xbit_r72_c82 bl[82] br[82] wl[72] vdd gnd cell_6t
Xbit_r73_c82 bl[82] br[82] wl[73] vdd gnd cell_6t
Xbit_r74_c82 bl[82] br[82] wl[74] vdd gnd cell_6t
Xbit_r75_c82 bl[82] br[82] wl[75] vdd gnd cell_6t
Xbit_r76_c82 bl[82] br[82] wl[76] vdd gnd cell_6t
Xbit_r77_c82 bl[82] br[82] wl[77] vdd gnd cell_6t
Xbit_r78_c82 bl[82] br[82] wl[78] vdd gnd cell_6t
Xbit_r79_c82 bl[82] br[82] wl[79] vdd gnd cell_6t
Xbit_r80_c82 bl[82] br[82] wl[80] vdd gnd cell_6t
Xbit_r81_c82 bl[82] br[82] wl[81] vdd gnd cell_6t
Xbit_r82_c82 bl[82] br[82] wl[82] vdd gnd cell_6t
Xbit_r83_c82 bl[82] br[82] wl[83] vdd gnd cell_6t
Xbit_r84_c82 bl[82] br[82] wl[84] vdd gnd cell_6t
Xbit_r85_c82 bl[82] br[82] wl[85] vdd gnd cell_6t
Xbit_r86_c82 bl[82] br[82] wl[86] vdd gnd cell_6t
Xbit_r87_c82 bl[82] br[82] wl[87] vdd gnd cell_6t
Xbit_r88_c82 bl[82] br[82] wl[88] vdd gnd cell_6t
Xbit_r89_c82 bl[82] br[82] wl[89] vdd gnd cell_6t
Xbit_r90_c82 bl[82] br[82] wl[90] vdd gnd cell_6t
Xbit_r91_c82 bl[82] br[82] wl[91] vdd gnd cell_6t
Xbit_r92_c82 bl[82] br[82] wl[92] vdd gnd cell_6t
Xbit_r93_c82 bl[82] br[82] wl[93] vdd gnd cell_6t
Xbit_r94_c82 bl[82] br[82] wl[94] vdd gnd cell_6t
Xbit_r95_c82 bl[82] br[82] wl[95] vdd gnd cell_6t
Xbit_r96_c82 bl[82] br[82] wl[96] vdd gnd cell_6t
Xbit_r97_c82 bl[82] br[82] wl[97] vdd gnd cell_6t
Xbit_r98_c82 bl[82] br[82] wl[98] vdd gnd cell_6t
Xbit_r99_c82 bl[82] br[82] wl[99] vdd gnd cell_6t
Xbit_r100_c82 bl[82] br[82] wl[100] vdd gnd cell_6t
Xbit_r101_c82 bl[82] br[82] wl[101] vdd gnd cell_6t
Xbit_r102_c82 bl[82] br[82] wl[102] vdd gnd cell_6t
Xbit_r103_c82 bl[82] br[82] wl[103] vdd gnd cell_6t
Xbit_r104_c82 bl[82] br[82] wl[104] vdd gnd cell_6t
Xbit_r105_c82 bl[82] br[82] wl[105] vdd gnd cell_6t
Xbit_r106_c82 bl[82] br[82] wl[106] vdd gnd cell_6t
Xbit_r107_c82 bl[82] br[82] wl[107] vdd gnd cell_6t
Xbit_r108_c82 bl[82] br[82] wl[108] vdd gnd cell_6t
Xbit_r109_c82 bl[82] br[82] wl[109] vdd gnd cell_6t
Xbit_r110_c82 bl[82] br[82] wl[110] vdd gnd cell_6t
Xbit_r111_c82 bl[82] br[82] wl[111] vdd gnd cell_6t
Xbit_r112_c82 bl[82] br[82] wl[112] vdd gnd cell_6t
Xbit_r113_c82 bl[82] br[82] wl[113] vdd gnd cell_6t
Xbit_r114_c82 bl[82] br[82] wl[114] vdd gnd cell_6t
Xbit_r115_c82 bl[82] br[82] wl[115] vdd gnd cell_6t
Xbit_r116_c82 bl[82] br[82] wl[116] vdd gnd cell_6t
Xbit_r117_c82 bl[82] br[82] wl[117] vdd gnd cell_6t
Xbit_r118_c82 bl[82] br[82] wl[118] vdd gnd cell_6t
Xbit_r119_c82 bl[82] br[82] wl[119] vdd gnd cell_6t
Xbit_r120_c82 bl[82] br[82] wl[120] vdd gnd cell_6t
Xbit_r121_c82 bl[82] br[82] wl[121] vdd gnd cell_6t
Xbit_r122_c82 bl[82] br[82] wl[122] vdd gnd cell_6t
Xbit_r123_c82 bl[82] br[82] wl[123] vdd gnd cell_6t
Xbit_r124_c82 bl[82] br[82] wl[124] vdd gnd cell_6t
Xbit_r125_c82 bl[82] br[82] wl[125] vdd gnd cell_6t
Xbit_r126_c82 bl[82] br[82] wl[126] vdd gnd cell_6t
Xbit_r127_c82 bl[82] br[82] wl[127] vdd gnd cell_6t
Xbit_r128_c82 bl[82] br[82] wl[128] vdd gnd cell_6t
Xbit_r129_c82 bl[82] br[82] wl[129] vdd gnd cell_6t
Xbit_r130_c82 bl[82] br[82] wl[130] vdd gnd cell_6t
Xbit_r131_c82 bl[82] br[82] wl[131] vdd gnd cell_6t
Xbit_r132_c82 bl[82] br[82] wl[132] vdd gnd cell_6t
Xbit_r133_c82 bl[82] br[82] wl[133] vdd gnd cell_6t
Xbit_r134_c82 bl[82] br[82] wl[134] vdd gnd cell_6t
Xbit_r135_c82 bl[82] br[82] wl[135] vdd gnd cell_6t
Xbit_r136_c82 bl[82] br[82] wl[136] vdd gnd cell_6t
Xbit_r137_c82 bl[82] br[82] wl[137] vdd gnd cell_6t
Xbit_r138_c82 bl[82] br[82] wl[138] vdd gnd cell_6t
Xbit_r139_c82 bl[82] br[82] wl[139] vdd gnd cell_6t
Xbit_r140_c82 bl[82] br[82] wl[140] vdd gnd cell_6t
Xbit_r141_c82 bl[82] br[82] wl[141] vdd gnd cell_6t
Xbit_r142_c82 bl[82] br[82] wl[142] vdd gnd cell_6t
Xbit_r143_c82 bl[82] br[82] wl[143] vdd gnd cell_6t
Xbit_r144_c82 bl[82] br[82] wl[144] vdd gnd cell_6t
Xbit_r145_c82 bl[82] br[82] wl[145] vdd gnd cell_6t
Xbit_r146_c82 bl[82] br[82] wl[146] vdd gnd cell_6t
Xbit_r147_c82 bl[82] br[82] wl[147] vdd gnd cell_6t
Xbit_r148_c82 bl[82] br[82] wl[148] vdd gnd cell_6t
Xbit_r149_c82 bl[82] br[82] wl[149] vdd gnd cell_6t
Xbit_r150_c82 bl[82] br[82] wl[150] vdd gnd cell_6t
Xbit_r151_c82 bl[82] br[82] wl[151] vdd gnd cell_6t
Xbit_r152_c82 bl[82] br[82] wl[152] vdd gnd cell_6t
Xbit_r153_c82 bl[82] br[82] wl[153] vdd gnd cell_6t
Xbit_r154_c82 bl[82] br[82] wl[154] vdd gnd cell_6t
Xbit_r155_c82 bl[82] br[82] wl[155] vdd gnd cell_6t
Xbit_r156_c82 bl[82] br[82] wl[156] vdd gnd cell_6t
Xbit_r157_c82 bl[82] br[82] wl[157] vdd gnd cell_6t
Xbit_r158_c82 bl[82] br[82] wl[158] vdd gnd cell_6t
Xbit_r159_c82 bl[82] br[82] wl[159] vdd gnd cell_6t
Xbit_r160_c82 bl[82] br[82] wl[160] vdd gnd cell_6t
Xbit_r161_c82 bl[82] br[82] wl[161] vdd gnd cell_6t
Xbit_r162_c82 bl[82] br[82] wl[162] vdd gnd cell_6t
Xbit_r163_c82 bl[82] br[82] wl[163] vdd gnd cell_6t
Xbit_r164_c82 bl[82] br[82] wl[164] vdd gnd cell_6t
Xbit_r165_c82 bl[82] br[82] wl[165] vdd gnd cell_6t
Xbit_r166_c82 bl[82] br[82] wl[166] vdd gnd cell_6t
Xbit_r167_c82 bl[82] br[82] wl[167] vdd gnd cell_6t
Xbit_r168_c82 bl[82] br[82] wl[168] vdd gnd cell_6t
Xbit_r169_c82 bl[82] br[82] wl[169] vdd gnd cell_6t
Xbit_r170_c82 bl[82] br[82] wl[170] vdd gnd cell_6t
Xbit_r171_c82 bl[82] br[82] wl[171] vdd gnd cell_6t
Xbit_r172_c82 bl[82] br[82] wl[172] vdd gnd cell_6t
Xbit_r173_c82 bl[82] br[82] wl[173] vdd gnd cell_6t
Xbit_r174_c82 bl[82] br[82] wl[174] vdd gnd cell_6t
Xbit_r175_c82 bl[82] br[82] wl[175] vdd gnd cell_6t
Xbit_r176_c82 bl[82] br[82] wl[176] vdd gnd cell_6t
Xbit_r177_c82 bl[82] br[82] wl[177] vdd gnd cell_6t
Xbit_r178_c82 bl[82] br[82] wl[178] vdd gnd cell_6t
Xbit_r179_c82 bl[82] br[82] wl[179] vdd gnd cell_6t
Xbit_r180_c82 bl[82] br[82] wl[180] vdd gnd cell_6t
Xbit_r181_c82 bl[82] br[82] wl[181] vdd gnd cell_6t
Xbit_r182_c82 bl[82] br[82] wl[182] vdd gnd cell_6t
Xbit_r183_c82 bl[82] br[82] wl[183] vdd gnd cell_6t
Xbit_r184_c82 bl[82] br[82] wl[184] vdd gnd cell_6t
Xbit_r185_c82 bl[82] br[82] wl[185] vdd gnd cell_6t
Xbit_r186_c82 bl[82] br[82] wl[186] vdd gnd cell_6t
Xbit_r187_c82 bl[82] br[82] wl[187] vdd gnd cell_6t
Xbit_r188_c82 bl[82] br[82] wl[188] vdd gnd cell_6t
Xbit_r189_c82 bl[82] br[82] wl[189] vdd gnd cell_6t
Xbit_r190_c82 bl[82] br[82] wl[190] vdd gnd cell_6t
Xbit_r191_c82 bl[82] br[82] wl[191] vdd gnd cell_6t
Xbit_r192_c82 bl[82] br[82] wl[192] vdd gnd cell_6t
Xbit_r193_c82 bl[82] br[82] wl[193] vdd gnd cell_6t
Xbit_r194_c82 bl[82] br[82] wl[194] vdd gnd cell_6t
Xbit_r195_c82 bl[82] br[82] wl[195] vdd gnd cell_6t
Xbit_r196_c82 bl[82] br[82] wl[196] vdd gnd cell_6t
Xbit_r197_c82 bl[82] br[82] wl[197] vdd gnd cell_6t
Xbit_r198_c82 bl[82] br[82] wl[198] vdd gnd cell_6t
Xbit_r199_c82 bl[82] br[82] wl[199] vdd gnd cell_6t
Xbit_r200_c82 bl[82] br[82] wl[200] vdd gnd cell_6t
Xbit_r201_c82 bl[82] br[82] wl[201] vdd gnd cell_6t
Xbit_r202_c82 bl[82] br[82] wl[202] vdd gnd cell_6t
Xbit_r203_c82 bl[82] br[82] wl[203] vdd gnd cell_6t
Xbit_r204_c82 bl[82] br[82] wl[204] vdd gnd cell_6t
Xbit_r205_c82 bl[82] br[82] wl[205] vdd gnd cell_6t
Xbit_r206_c82 bl[82] br[82] wl[206] vdd gnd cell_6t
Xbit_r207_c82 bl[82] br[82] wl[207] vdd gnd cell_6t
Xbit_r208_c82 bl[82] br[82] wl[208] vdd gnd cell_6t
Xbit_r209_c82 bl[82] br[82] wl[209] vdd gnd cell_6t
Xbit_r210_c82 bl[82] br[82] wl[210] vdd gnd cell_6t
Xbit_r211_c82 bl[82] br[82] wl[211] vdd gnd cell_6t
Xbit_r212_c82 bl[82] br[82] wl[212] vdd gnd cell_6t
Xbit_r213_c82 bl[82] br[82] wl[213] vdd gnd cell_6t
Xbit_r214_c82 bl[82] br[82] wl[214] vdd gnd cell_6t
Xbit_r215_c82 bl[82] br[82] wl[215] vdd gnd cell_6t
Xbit_r216_c82 bl[82] br[82] wl[216] vdd gnd cell_6t
Xbit_r217_c82 bl[82] br[82] wl[217] vdd gnd cell_6t
Xbit_r218_c82 bl[82] br[82] wl[218] vdd gnd cell_6t
Xbit_r219_c82 bl[82] br[82] wl[219] vdd gnd cell_6t
Xbit_r220_c82 bl[82] br[82] wl[220] vdd gnd cell_6t
Xbit_r221_c82 bl[82] br[82] wl[221] vdd gnd cell_6t
Xbit_r222_c82 bl[82] br[82] wl[222] vdd gnd cell_6t
Xbit_r223_c82 bl[82] br[82] wl[223] vdd gnd cell_6t
Xbit_r224_c82 bl[82] br[82] wl[224] vdd gnd cell_6t
Xbit_r225_c82 bl[82] br[82] wl[225] vdd gnd cell_6t
Xbit_r226_c82 bl[82] br[82] wl[226] vdd gnd cell_6t
Xbit_r227_c82 bl[82] br[82] wl[227] vdd gnd cell_6t
Xbit_r228_c82 bl[82] br[82] wl[228] vdd gnd cell_6t
Xbit_r229_c82 bl[82] br[82] wl[229] vdd gnd cell_6t
Xbit_r230_c82 bl[82] br[82] wl[230] vdd gnd cell_6t
Xbit_r231_c82 bl[82] br[82] wl[231] vdd gnd cell_6t
Xbit_r232_c82 bl[82] br[82] wl[232] vdd gnd cell_6t
Xbit_r233_c82 bl[82] br[82] wl[233] vdd gnd cell_6t
Xbit_r234_c82 bl[82] br[82] wl[234] vdd gnd cell_6t
Xbit_r235_c82 bl[82] br[82] wl[235] vdd gnd cell_6t
Xbit_r236_c82 bl[82] br[82] wl[236] vdd gnd cell_6t
Xbit_r237_c82 bl[82] br[82] wl[237] vdd gnd cell_6t
Xbit_r238_c82 bl[82] br[82] wl[238] vdd gnd cell_6t
Xbit_r239_c82 bl[82] br[82] wl[239] vdd gnd cell_6t
Xbit_r240_c82 bl[82] br[82] wl[240] vdd gnd cell_6t
Xbit_r241_c82 bl[82] br[82] wl[241] vdd gnd cell_6t
Xbit_r242_c82 bl[82] br[82] wl[242] vdd gnd cell_6t
Xbit_r243_c82 bl[82] br[82] wl[243] vdd gnd cell_6t
Xbit_r244_c82 bl[82] br[82] wl[244] vdd gnd cell_6t
Xbit_r245_c82 bl[82] br[82] wl[245] vdd gnd cell_6t
Xbit_r246_c82 bl[82] br[82] wl[246] vdd gnd cell_6t
Xbit_r247_c82 bl[82] br[82] wl[247] vdd gnd cell_6t
Xbit_r248_c82 bl[82] br[82] wl[248] vdd gnd cell_6t
Xbit_r249_c82 bl[82] br[82] wl[249] vdd gnd cell_6t
Xbit_r250_c82 bl[82] br[82] wl[250] vdd gnd cell_6t
Xbit_r251_c82 bl[82] br[82] wl[251] vdd gnd cell_6t
Xbit_r252_c82 bl[82] br[82] wl[252] vdd gnd cell_6t
Xbit_r253_c82 bl[82] br[82] wl[253] vdd gnd cell_6t
Xbit_r254_c82 bl[82] br[82] wl[254] vdd gnd cell_6t
Xbit_r255_c82 bl[82] br[82] wl[255] vdd gnd cell_6t
Xbit_r0_c83 bl[83] br[83] wl[0] vdd gnd cell_6t
Xbit_r1_c83 bl[83] br[83] wl[1] vdd gnd cell_6t
Xbit_r2_c83 bl[83] br[83] wl[2] vdd gnd cell_6t
Xbit_r3_c83 bl[83] br[83] wl[3] vdd gnd cell_6t
Xbit_r4_c83 bl[83] br[83] wl[4] vdd gnd cell_6t
Xbit_r5_c83 bl[83] br[83] wl[5] vdd gnd cell_6t
Xbit_r6_c83 bl[83] br[83] wl[6] vdd gnd cell_6t
Xbit_r7_c83 bl[83] br[83] wl[7] vdd gnd cell_6t
Xbit_r8_c83 bl[83] br[83] wl[8] vdd gnd cell_6t
Xbit_r9_c83 bl[83] br[83] wl[9] vdd gnd cell_6t
Xbit_r10_c83 bl[83] br[83] wl[10] vdd gnd cell_6t
Xbit_r11_c83 bl[83] br[83] wl[11] vdd gnd cell_6t
Xbit_r12_c83 bl[83] br[83] wl[12] vdd gnd cell_6t
Xbit_r13_c83 bl[83] br[83] wl[13] vdd gnd cell_6t
Xbit_r14_c83 bl[83] br[83] wl[14] vdd gnd cell_6t
Xbit_r15_c83 bl[83] br[83] wl[15] vdd gnd cell_6t
Xbit_r16_c83 bl[83] br[83] wl[16] vdd gnd cell_6t
Xbit_r17_c83 bl[83] br[83] wl[17] vdd gnd cell_6t
Xbit_r18_c83 bl[83] br[83] wl[18] vdd gnd cell_6t
Xbit_r19_c83 bl[83] br[83] wl[19] vdd gnd cell_6t
Xbit_r20_c83 bl[83] br[83] wl[20] vdd gnd cell_6t
Xbit_r21_c83 bl[83] br[83] wl[21] vdd gnd cell_6t
Xbit_r22_c83 bl[83] br[83] wl[22] vdd gnd cell_6t
Xbit_r23_c83 bl[83] br[83] wl[23] vdd gnd cell_6t
Xbit_r24_c83 bl[83] br[83] wl[24] vdd gnd cell_6t
Xbit_r25_c83 bl[83] br[83] wl[25] vdd gnd cell_6t
Xbit_r26_c83 bl[83] br[83] wl[26] vdd gnd cell_6t
Xbit_r27_c83 bl[83] br[83] wl[27] vdd gnd cell_6t
Xbit_r28_c83 bl[83] br[83] wl[28] vdd gnd cell_6t
Xbit_r29_c83 bl[83] br[83] wl[29] vdd gnd cell_6t
Xbit_r30_c83 bl[83] br[83] wl[30] vdd gnd cell_6t
Xbit_r31_c83 bl[83] br[83] wl[31] vdd gnd cell_6t
Xbit_r32_c83 bl[83] br[83] wl[32] vdd gnd cell_6t
Xbit_r33_c83 bl[83] br[83] wl[33] vdd gnd cell_6t
Xbit_r34_c83 bl[83] br[83] wl[34] vdd gnd cell_6t
Xbit_r35_c83 bl[83] br[83] wl[35] vdd gnd cell_6t
Xbit_r36_c83 bl[83] br[83] wl[36] vdd gnd cell_6t
Xbit_r37_c83 bl[83] br[83] wl[37] vdd gnd cell_6t
Xbit_r38_c83 bl[83] br[83] wl[38] vdd gnd cell_6t
Xbit_r39_c83 bl[83] br[83] wl[39] vdd gnd cell_6t
Xbit_r40_c83 bl[83] br[83] wl[40] vdd gnd cell_6t
Xbit_r41_c83 bl[83] br[83] wl[41] vdd gnd cell_6t
Xbit_r42_c83 bl[83] br[83] wl[42] vdd gnd cell_6t
Xbit_r43_c83 bl[83] br[83] wl[43] vdd gnd cell_6t
Xbit_r44_c83 bl[83] br[83] wl[44] vdd gnd cell_6t
Xbit_r45_c83 bl[83] br[83] wl[45] vdd gnd cell_6t
Xbit_r46_c83 bl[83] br[83] wl[46] vdd gnd cell_6t
Xbit_r47_c83 bl[83] br[83] wl[47] vdd gnd cell_6t
Xbit_r48_c83 bl[83] br[83] wl[48] vdd gnd cell_6t
Xbit_r49_c83 bl[83] br[83] wl[49] vdd gnd cell_6t
Xbit_r50_c83 bl[83] br[83] wl[50] vdd gnd cell_6t
Xbit_r51_c83 bl[83] br[83] wl[51] vdd gnd cell_6t
Xbit_r52_c83 bl[83] br[83] wl[52] vdd gnd cell_6t
Xbit_r53_c83 bl[83] br[83] wl[53] vdd gnd cell_6t
Xbit_r54_c83 bl[83] br[83] wl[54] vdd gnd cell_6t
Xbit_r55_c83 bl[83] br[83] wl[55] vdd gnd cell_6t
Xbit_r56_c83 bl[83] br[83] wl[56] vdd gnd cell_6t
Xbit_r57_c83 bl[83] br[83] wl[57] vdd gnd cell_6t
Xbit_r58_c83 bl[83] br[83] wl[58] vdd gnd cell_6t
Xbit_r59_c83 bl[83] br[83] wl[59] vdd gnd cell_6t
Xbit_r60_c83 bl[83] br[83] wl[60] vdd gnd cell_6t
Xbit_r61_c83 bl[83] br[83] wl[61] vdd gnd cell_6t
Xbit_r62_c83 bl[83] br[83] wl[62] vdd gnd cell_6t
Xbit_r63_c83 bl[83] br[83] wl[63] vdd gnd cell_6t
Xbit_r64_c83 bl[83] br[83] wl[64] vdd gnd cell_6t
Xbit_r65_c83 bl[83] br[83] wl[65] vdd gnd cell_6t
Xbit_r66_c83 bl[83] br[83] wl[66] vdd gnd cell_6t
Xbit_r67_c83 bl[83] br[83] wl[67] vdd gnd cell_6t
Xbit_r68_c83 bl[83] br[83] wl[68] vdd gnd cell_6t
Xbit_r69_c83 bl[83] br[83] wl[69] vdd gnd cell_6t
Xbit_r70_c83 bl[83] br[83] wl[70] vdd gnd cell_6t
Xbit_r71_c83 bl[83] br[83] wl[71] vdd gnd cell_6t
Xbit_r72_c83 bl[83] br[83] wl[72] vdd gnd cell_6t
Xbit_r73_c83 bl[83] br[83] wl[73] vdd gnd cell_6t
Xbit_r74_c83 bl[83] br[83] wl[74] vdd gnd cell_6t
Xbit_r75_c83 bl[83] br[83] wl[75] vdd gnd cell_6t
Xbit_r76_c83 bl[83] br[83] wl[76] vdd gnd cell_6t
Xbit_r77_c83 bl[83] br[83] wl[77] vdd gnd cell_6t
Xbit_r78_c83 bl[83] br[83] wl[78] vdd gnd cell_6t
Xbit_r79_c83 bl[83] br[83] wl[79] vdd gnd cell_6t
Xbit_r80_c83 bl[83] br[83] wl[80] vdd gnd cell_6t
Xbit_r81_c83 bl[83] br[83] wl[81] vdd gnd cell_6t
Xbit_r82_c83 bl[83] br[83] wl[82] vdd gnd cell_6t
Xbit_r83_c83 bl[83] br[83] wl[83] vdd gnd cell_6t
Xbit_r84_c83 bl[83] br[83] wl[84] vdd gnd cell_6t
Xbit_r85_c83 bl[83] br[83] wl[85] vdd gnd cell_6t
Xbit_r86_c83 bl[83] br[83] wl[86] vdd gnd cell_6t
Xbit_r87_c83 bl[83] br[83] wl[87] vdd gnd cell_6t
Xbit_r88_c83 bl[83] br[83] wl[88] vdd gnd cell_6t
Xbit_r89_c83 bl[83] br[83] wl[89] vdd gnd cell_6t
Xbit_r90_c83 bl[83] br[83] wl[90] vdd gnd cell_6t
Xbit_r91_c83 bl[83] br[83] wl[91] vdd gnd cell_6t
Xbit_r92_c83 bl[83] br[83] wl[92] vdd gnd cell_6t
Xbit_r93_c83 bl[83] br[83] wl[93] vdd gnd cell_6t
Xbit_r94_c83 bl[83] br[83] wl[94] vdd gnd cell_6t
Xbit_r95_c83 bl[83] br[83] wl[95] vdd gnd cell_6t
Xbit_r96_c83 bl[83] br[83] wl[96] vdd gnd cell_6t
Xbit_r97_c83 bl[83] br[83] wl[97] vdd gnd cell_6t
Xbit_r98_c83 bl[83] br[83] wl[98] vdd gnd cell_6t
Xbit_r99_c83 bl[83] br[83] wl[99] vdd gnd cell_6t
Xbit_r100_c83 bl[83] br[83] wl[100] vdd gnd cell_6t
Xbit_r101_c83 bl[83] br[83] wl[101] vdd gnd cell_6t
Xbit_r102_c83 bl[83] br[83] wl[102] vdd gnd cell_6t
Xbit_r103_c83 bl[83] br[83] wl[103] vdd gnd cell_6t
Xbit_r104_c83 bl[83] br[83] wl[104] vdd gnd cell_6t
Xbit_r105_c83 bl[83] br[83] wl[105] vdd gnd cell_6t
Xbit_r106_c83 bl[83] br[83] wl[106] vdd gnd cell_6t
Xbit_r107_c83 bl[83] br[83] wl[107] vdd gnd cell_6t
Xbit_r108_c83 bl[83] br[83] wl[108] vdd gnd cell_6t
Xbit_r109_c83 bl[83] br[83] wl[109] vdd gnd cell_6t
Xbit_r110_c83 bl[83] br[83] wl[110] vdd gnd cell_6t
Xbit_r111_c83 bl[83] br[83] wl[111] vdd gnd cell_6t
Xbit_r112_c83 bl[83] br[83] wl[112] vdd gnd cell_6t
Xbit_r113_c83 bl[83] br[83] wl[113] vdd gnd cell_6t
Xbit_r114_c83 bl[83] br[83] wl[114] vdd gnd cell_6t
Xbit_r115_c83 bl[83] br[83] wl[115] vdd gnd cell_6t
Xbit_r116_c83 bl[83] br[83] wl[116] vdd gnd cell_6t
Xbit_r117_c83 bl[83] br[83] wl[117] vdd gnd cell_6t
Xbit_r118_c83 bl[83] br[83] wl[118] vdd gnd cell_6t
Xbit_r119_c83 bl[83] br[83] wl[119] vdd gnd cell_6t
Xbit_r120_c83 bl[83] br[83] wl[120] vdd gnd cell_6t
Xbit_r121_c83 bl[83] br[83] wl[121] vdd gnd cell_6t
Xbit_r122_c83 bl[83] br[83] wl[122] vdd gnd cell_6t
Xbit_r123_c83 bl[83] br[83] wl[123] vdd gnd cell_6t
Xbit_r124_c83 bl[83] br[83] wl[124] vdd gnd cell_6t
Xbit_r125_c83 bl[83] br[83] wl[125] vdd gnd cell_6t
Xbit_r126_c83 bl[83] br[83] wl[126] vdd gnd cell_6t
Xbit_r127_c83 bl[83] br[83] wl[127] vdd gnd cell_6t
Xbit_r128_c83 bl[83] br[83] wl[128] vdd gnd cell_6t
Xbit_r129_c83 bl[83] br[83] wl[129] vdd gnd cell_6t
Xbit_r130_c83 bl[83] br[83] wl[130] vdd gnd cell_6t
Xbit_r131_c83 bl[83] br[83] wl[131] vdd gnd cell_6t
Xbit_r132_c83 bl[83] br[83] wl[132] vdd gnd cell_6t
Xbit_r133_c83 bl[83] br[83] wl[133] vdd gnd cell_6t
Xbit_r134_c83 bl[83] br[83] wl[134] vdd gnd cell_6t
Xbit_r135_c83 bl[83] br[83] wl[135] vdd gnd cell_6t
Xbit_r136_c83 bl[83] br[83] wl[136] vdd gnd cell_6t
Xbit_r137_c83 bl[83] br[83] wl[137] vdd gnd cell_6t
Xbit_r138_c83 bl[83] br[83] wl[138] vdd gnd cell_6t
Xbit_r139_c83 bl[83] br[83] wl[139] vdd gnd cell_6t
Xbit_r140_c83 bl[83] br[83] wl[140] vdd gnd cell_6t
Xbit_r141_c83 bl[83] br[83] wl[141] vdd gnd cell_6t
Xbit_r142_c83 bl[83] br[83] wl[142] vdd gnd cell_6t
Xbit_r143_c83 bl[83] br[83] wl[143] vdd gnd cell_6t
Xbit_r144_c83 bl[83] br[83] wl[144] vdd gnd cell_6t
Xbit_r145_c83 bl[83] br[83] wl[145] vdd gnd cell_6t
Xbit_r146_c83 bl[83] br[83] wl[146] vdd gnd cell_6t
Xbit_r147_c83 bl[83] br[83] wl[147] vdd gnd cell_6t
Xbit_r148_c83 bl[83] br[83] wl[148] vdd gnd cell_6t
Xbit_r149_c83 bl[83] br[83] wl[149] vdd gnd cell_6t
Xbit_r150_c83 bl[83] br[83] wl[150] vdd gnd cell_6t
Xbit_r151_c83 bl[83] br[83] wl[151] vdd gnd cell_6t
Xbit_r152_c83 bl[83] br[83] wl[152] vdd gnd cell_6t
Xbit_r153_c83 bl[83] br[83] wl[153] vdd gnd cell_6t
Xbit_r154_c83 bl[83] br[83] wl[154] vdd gnd cell_6t
Xbit_r155_c83 bl[83] br[83] wl[155] vdd gnd cell_6t
Xbit_r156_c83 bl[83] br[83] wl[156] vdd gnd cell_6t
Xbit_r157_c83 bl[83] br[83] wl[157] vdd gnd cell_6t
Xbit_r158_c83 bl[83] br[83] wl[158] vdd gnd cell_6t
Xbit_r159_c83 bl[83] br[83] wl[159] vdd gnd cell_6t
Xbit_r160_c83 bl[83] br[83] wl[160] vdd gnd cell_6t
Xbit_r161_c83 bl[83] br[83] wl[161] vdd gnd cell_6t
Xbit_r162_c83 bl[83] br[83] wl[162] vdd gnd cell_6t
Xbit_r163_c83 bl[83] br[83] wl[163] vdd gnd cell_6t
Xbit_r164_c83 bl[83] br[83] wl[164] vdd gnd cell_6t
Xbit_r165_c83 bl[83] br[83] wl[165] vdd gnd cell_6t
Xbit_r166_c83 bl[83] br[83] wl[166] vdd gnd cell_6t
Xbit_r167_c83 bl[83] br[83] wl[167] vdd gnd cell_6t
Xbit_r168_c83 bl[83] br[83] wl[168] vdd gnd cell_6t
Xbit_r169_c83 bl[83] br[83] wl[169] vdd gnd cell_6t
Xbit_r170_c83 bl[83] br[83] wl[170] vdd gnd cell_6t
Xbit_r171_c83 bl[83] br[83] wl[171] vdd gnd cell_6t
Xbit_r172_c83 bl[83] br[83] wl[172] vdd gnd cell_6t
Xbit_r173_c83 bl[83] br[83] wl[173] vdd gnd cell_6t
Xbit_r174_c83 bl[83] br[83] wl[174] vdd gnd cell_6t
Xbit_r175_c83 bl[83] br[83] wl[175] vdd gnd cell_6t
Xbit_r176_c83 bl[83] br[83] wl[176] vdd gnd cell_6t
Xbit_r177_c83 bl[83] br[83] wl[177] vdd gnd cell_6t
Xbit_r178_c83 bl[83] br[83] wl[178] vdd gnd cell_6t
Xbit_r179_c83 bl[83] br[83] wl[179] vdd gnd cell_6t
Xbit_r180_c83 bl[83] br[83] wl[180] vdd gnd cell_6t
Xbit_r181_c83 bl[83] br[83] wl[181] vdd gnd cell_6t
Xbit_r182_c83 bl[83] br[83] wl[182] vdd gnd cell_6t
Xbit_r183_c83 bl[83] br[83] wl[183] vdd gnd cell_6t
Xbit_r184_c83 bl[83] br[83] wl[184] vdd gnd cell_6t
Xbit_r185_c83 bl[83] br[83] wl[185] vdd gnd cell_6t
Xbit_r186_c83 bl[83] br[83] wl[186] vdd gnd cell_6t
Xbit_r187_c83 bl[83] br[83] wl[187] vdd gnd cell_6t
Xbit_r188_c83 bl[83] br[83] wl[188] vdd gnd cell_6t
Xbit_r189_c83 bl[83] br[83] wl[189] vdd gnd cell_6t
Xbit_r190_c83 bl[83] br[83] wl[190] vdd gnd cell_6t
Xbit_r191_c83 bl[83] br[83] wl[191] vdd gnd cell_6t
Xbit_r192_c83 bl[83] br[83] wl[192] vdd gnd cell_6t
Xbit_r193_c83 bl[83] br[83] wl[193] vdd gnd cell_6t
Xbit_r194_c83 bl[83] br[83] wl[194] vdd gnd cell_6t
Xbit_r195_c83 bl[83] br[83] wl[195] vdd gnd cell_6t
Xbit_r196_c83 bl[83] br[83] wl[196] vdd gnd cell_6t
Xbit_r197_c83 bl[83] br[83] wl[197] vdd gnd cell_6t
Xbit_r198_c83 bl[83] br[83] wl[198] vdd gnd cell_6t
Xbit_r199_c83 bl[83] br[83] wl[199] vdd gnd cell_6t
Xbit_r200_c83 bl[83] br[83] wl[200] vdd gnd cell_6t
Xbit_r201_c83 bl[83] br[83] wl[201] vdd gnd cell_6t
Xbit_r202_c83 bl[83] br[83] wl[202] vdd gnd cell_6t
Xbit_r203_c83 bl[83] br[83] wl[203] vdd gnd cell_6t
Xbit_r204_c83 bl[83] br[83] wl[204] vdd gnd cell_6t
Xbit_r205_c83 bl[83] br[83] wl[205] vdd gnd cell_6t
Xbit_r206_c83 bl[83] br[83] wl[206] vdd gnd cell_6t
Xbit_r207_c83 bl[83] br[83] wl[207] vdd gnd cell_6t
Xbit_r208_c83 bl[83] br[83] wl[208] vdd gnd cell_6t
Xbit_r209_c83 bl[83] br[83] wl[209] vdd gnd cell_6t
Xbit_r210_c83 bl[83] br[83] wl[210] vdd gnd cell_6t
Xbit_r211_c83 bl[83] br[83] wl[211] vdd gnd cell_6t
Xbit_r212_c83 bl[83] br[83] wl[212] vdd gnd cell_6t
Xbit_r213_c83 bl[83] br[83] wl[213] vdd gnd cell_6t
Xbit_r214_c83 bl[83] br[83] wl[214] vdd gnd cell_6t
Xbit_r215_c83 bl[83] br[83] wl[215] vdd gnd cell_6t
Xbit_r216_c83 bl[83] br[83] wl[216] vdd gnd cell_6t
Xbit_r217_c83 bl[83] br[83] wl[217] vdd gnd cell_6t
Xbit_r218_c83 bl[83] br[83] wl[218] vdd gnd cell_6t
Xbit_r219_c83 bl[83] br[83] wl[219] vdd gnd cell_6t
Xbit_r220_c83 bl[83] br[83] wl[220] vdd gnd cell_6t
Xbit_r221_c83 bl[83] br[83] wl[221] vdd gnd cell_6t
Xbit_r222_c83 bl[83] br[83] wl[222] vdd gnd cell_6t
Xbit_r223_c83 bl[83] br[83] wl[223] vdd gnd cell_6t
Xbit_r224_c83 bl[83] br[83] wl[224] vdd gnd cell_6t
Xbit_r225_c83 bl[83] br[83] wl[225] vdd gnd cell_6t
Xbit_r226_c83 bl[83] br[83] wl[226] vdd gnd cell_6t
Xbit_r227_c83 bl[83] br[83] wl[227] vdd gnd cell_6t
Xbit_r228_c83 bl[83] br[83] wl[228] vdd gnd cell_6t
Xbit_r229_c83 bl[83] br[83] wl[229] vdd gnd cell_6t
Xbit_r230_c83 bl[83] br[83] wl[230] vdd gnd cell_6t
Xbit_r231_c83 bl[83] br[83] wl[231] vdd gnd cell_6t
Xbit_r232_c83 bl[83] br[83] wl[232] vdd gnd cell_6t
Xbit_r233_c83 bl[83] br[83] wl[233] vdd gnd cell_6t
Xbit_r234_c83 bl[83] br[83] wl[234] vdd gnd cell_6t
Xbit_r235_c83 bl[83] br[83] wl[235] vdd gnd cell_6t
Xbit_r236_c83 bl[83] br[83] wl[236] vdd gnd cell_6t
Xbit_r237_c83 bl[83] br[83] wl[237] vdd gnd cell_6t
Xbit_r238_c83 bl[83] br[83] wl[238] vdd gnd cell_6t
Xbit_r239_c83 bl[83] br[83] wl[239] vdd gnd cell_6t
Xbit_r240_c83 bl[83] br[83] wl[240] vdd gnd cell_6t
Xbit_r241_c83 bl[83] br[83] wl[241] vdd gnd cell_6t
Xbit_r242_c83 bl[83] br[83] wl[242] vdd gnd cell_6t
Xbit_r243_c83 bl[83] br[83] wl[243] vdd gnd cell_6t
Xbit_r244_c83 bl[83] br[83] wl[244] vdd gnd cell_6t
Xbit_r245_c83 bl[83] br[83] wl[245] vdd gnd cell_6t
Xbit_r246_c83 bl[83] br[83] wl[246] vdd gnd cell_6t
Xbit_r247_c83 bl[83] br[83] wl[247] vdd gnd cell_6t
Xbit_r248_c83 bl[83] br[83] wl[248] vdd gnd cell_6t
Xbit_r249_c83 bl[83] br[83] wl[249] vdd gnd cell_6t
Xbit_r250_c83 bl[83] br[83] wl[250] vdd gnd cell_6t
Xbit_r251_c83 bl[83] br[83] wl[251] vdd gnd cell_6t
Xbit_r252_c83 bl[83] br[83] wl[252] vdd gnd cell_6t
Xbit_r253_c83 bl[83] br[83] wl[253] vdd gnd cell_6t
Xbit_r254_c83 bl[83] br[83] wl[254] vdd gnd cell_6t
Xbit_r255_c83 bl[83] br[83] wl[255] vdd gnd cell_6t
Xbit_r0_c84 bl[84] br[84] wl[0] vdd gnd cell_6t
Xbit_r1_c84 bl[84] br[84] wl[1] vdd gnd cell_6t
Xbit_r2_c84 bl[84] br[84] wl[2] vdd gnd cell_6t
Xbit_r3_c84 bl[84] br[84] wl[3] vdd gnd cell_6t
Xbit_r4_c84 bl[84] br[84] wl[4] vdd gnd cell_6t
Xbit_r5_c84 bl[84] br[84] wl[5] vdd gnd cell_6t
Xbit_r6_c84 bl[84] br[84] wl[6] vdd gnd cell_6t
Xbit_r7_c84 bl[84] br[84] wl[7] vdd gnd cell_6t
Xbit_r8_c84 bl[84] br[84] wl[8] vdd gnd cell_6t
Xbit_r9_c84 bl[84] br[84] wl[9] vdd gnd cell_6t
Xbit_r10_c84 bl[84] br[84] wl[10] vdd gnd cell_6t
Xbit_r11_c84 bl[84] br[84] wl[11] vdd gnd cell_6t
Xbit_r12_c84 bl[84] br[84] wl[12] vdd gnd cell_6t
Xbit_r13_c84 bl[84] br[84] wl[13] vdd gnd cell_6t
Xbit_r14_c84 bl[84] br[84] wl[14] vdd gnd cell_6t
Xbit_r15_c84 bl[84] br[84] wl[15] vdd gnd cell_6t
Xbit_r16_c84 bl[84] br[84] wl[16] vdd gnd cell_6t
Xbit_r17_c84 bl[84] br[84] wl[17] vdd gnd cell_6t
Xbit_r18_c84 bl[84] br[84] wl[18] vdd gnd cell_6t
Xbit_r19_c84 bl[84] br[84] wl[19] vdd gnd cell_6t
Xbit_r20_c84 bl[84] br[84] wl[20] vdd gnd cell_6t
Xbit_r21_c84 bl[84] br[84] wl[21] vdd gnd cell_6t
Xbit_r22_c84 bl[84] br[84] wl[22] vdd gnd cell_6t
Xbit_r23_c84 bl[84] br[84] wl[23] vdd gnd cell_6t
Xbit_r24_c84 bl[84] br[84] wl[24] vdd gnd cell_6t
Xbit_r25_c84 bl[84] br[84] wl[25] vdd gnd cell_6t
Xbit_r26_c84 bl[84] br[84] wl[26] vdd gnd cell_6t
Xbit_r27_c84 bl[84] br[84] wl[27] vdd gnd cell_6t
Xbit_r28_c84 bl[84] br[84] wl[28] vdd gnd cell_6t
Xbit_r29_c84 bl[84] br[84] wl[29] vdd gnd cell_6t
Xbit_r30_c84 bl[84] br[84] wl[30] vdd gnd cell_6t
Xbit_r31_c84 bl[84] br[84] wl[31] vdd gnd cell_6t
Xbit_r32_c84 bl[84] br[84] wl[32] vdd gnd cell_6t
Xbit_r33_c84 bl[84] br[84] wl[33] vdd gnd cell_6t
Xbit_r34_c84 bl[84] br[84] wl[34] vdd gnd cell_6t
Xbit_r35_c84 bl[84] br[84] wl[35] vdd gnd cell_6t
Xbit_r36_c84 bl[84] br[84] wl[36] vdd gnd cell_6t
Xbit_r37_c84 bl[84] br[84] wl[37] vdd gnd cell_6t
Xbit_r38_c84 bl[84] br[84] wl[38] vdd gnd cell_6t
Xbit_r39_c84 bl[84] br[84] wl[39] vdd gnd cell_6t
Xbit_r40_c84 bl[84] br[84] wl[40] vdd gnd cell_6t
Xbit_r41_c84 bl[84] br[84] wl[41] vdd gnd cell_6t
Xbit_r42_c84 bl[84] br[84] wl[42] vdd gnd cell_6t
Xbit_r43_c84 bl[84] br[84] wl[43] vdd gnd cell_6t
Xbit_r44_c84 bl[84] br[84] wl[44] vdd gnd cell_6t
Xbit_r45_c84 bl[84] br[84] wl[45] vdd gnd cell_6t
Xbit_r46_c84 bl[84] br[84] wl[46] vdd gnd cell_6t
Xbit_r47_c84 bl[84] br[84] wl[47] vdd gnd cell_6t
Xbit_r48_c84 bl[84] br[84] wl[48] vdd gnd cell_6t
Xbit_r49_c84 bl[84] br[84] wl[49] vdd gnd cell_6t
Xbit_r50_c84 bl[84] br[84] wl[50] vdd gnd cell_6t
Xbit_r51_c84 bl[84] br[84] wl[51] vdd gnd cell_6t
Xbit_r52_c84 bl[84] br[84] wl[52] vdd gnd cell_6t
Xbit_r53_c84 bl[84] br[84] wl[53] vdd gnd cell_6t
Xbit_r54_c84 bl[84] br[84] wl[54] vdd gnd cell_6t
Xbit_r55_c84 bl[84] br[84] wl[55] vdd gnd cell_6t
Xbit_r56_c84 bl[84] br[84] wl[56] vdd gnd cell_6t
Xbit_r57_c84 bl[84] br[84] wl[57] vdd gnd cell_6t
Xbit_r58_c84 bl[84] br[84] wl[58] vdd gnd cell_6t
Xbit_r59_c84 bl[84] br[84] wl[59] vdd gnd cell_6t
Xbit_r60_c84 bl[84] br[84] wl[60] vdd gnd cell_6t
Xbit_r61_c84 bl[84] br[84] wl[61] vdd gnd cell_6t
Xbit_r62_c84 bl[84] br[84] wl[62] vdd gnd cell_6t
Xbit_r63_c84 bl[84] br[84] wl[63] vdd gnd cell_6t
Xbit_r64_c84 bl[84] br[84] wl[64] vdd gnd cell_6t
Xbit_r65_c84 bl[84] br[84] wl[65] vdd gnd cell_6t
Xbit_r66_c84 bl[84] br[84] wl[66] vdd gnd cell_6t
Xbit_r67_c84 bl[84] br[84] wl[67] vdd gnd cell_6t
Xbit_r68_c84 bl[84] br[84] wl[68] vdd gnd cell_6t
Xbit_r69_c84 bl[84] br[84] wl[69] vdd gnd cell_6t
Xbit_r70_c84 bl[84] br[84] wl[70] vdd gnd cell_6t
Xbit_r71_c84 bl[84] br[84] wl[71] vdd gnd cell_6t
Xbit_r72_c84 bl[84] br[84] wl[72] vdd gnd cell_6t
Xbit_r73_c84 bl[84] br[84] wl[73] vdd gnd cell_6t
Xbit_r74_c84 bl[84] br[84] wl[74] vdd gnd cell_6t
Xbit_r75_c84 bl[84] br[84] wl[75] vdd gnd cell_6t
Xbit_r76_c84 bl[84] br[84] wl[76] vdd gnd cell_6t
Xbit_r77_c84 bl[84] br[84] wl[77] vdd gnd cell_6t
Xbit_r78_c84 bl[84] br[84] wl[78] vdd gnd cell_6t
Xbit_r79_c84 bl[84] br[84] wl[79] vdd gnd cell_6t
Xbit_r80_c84 bl[84] br[84] wl[80] vdd gnd cell_6t
Xbit_r81_c84 bl[84] br[84] wl[81] vdd gnd cell_6t
Xbit_r82_c84 bl[84] br[84] wl[82] vdd gnd cell_6t
Xbit_r83_c84 bl[84] br[84] wl[83] vdd gnd cell_6t
Xbit_r84_c84 bl[84] br[84] wl[84] vdd gnd cell_6t
Xbit_r85_c84 bl[84] br[84] wl[85] vdd gnd cell_6t
Xbit_r86_c84 bl[84] br[84] wl[86] vdd gnd cell_6t
Xbit_r87_c84 bl[84] br[84] wl[87] vdd gnd cell_6t
Xbit_r88_c84 bl[84] br[84] wl[88] vdd gnd cell_6t
Xbit_r89_c84 bl[84] br[84] wl[89] vdd gnd cell_6t
Xbit_r90_c84 bl[84] br[84] wl[90] vdd gnd cell_6t
Xbit_r91_c84 bl[84] br[84] wl[91] vdd gnd cell_6t
Xbit_r92_c84 bl[84] br[84] wl[92] vdd gnd cell_6t
Xbit_r93_c84 bl[84] br[84] wl[93] vdd gnd cell_6t
Xbit_r94_c84 bl[84] br[84] wl[94] vdd gnd cell_6t
Xbit_r95_c84 bl[84] br[84] wl[95] vdd gnd cell_6t
Xbit_r96_c84 bl[84] br[84] wl[96] vdd gnd cell_6t
Xbit_r97_c84 bl[84] br[84] wl[97] vdd gnd cell_6t
Xbit_r98_c84 bl[84] br[84] wl[98] vdd gnd cell_6t
Xbit_r99_c84 bl[84] br[84] wl[99] vdd gnd cell_6t
Xbit_r100_c84 bl[84] br[84] wl[100] vdd gnd cell_6t
Xbit_r101_c84 bl[84] br[84] wl[101] vdd gnd cell_6t
Xbit_r102_c84 bl[84] br[84] wl[102] vdd gnd cell_6t
Xbit_r103_c84 bl[84] br[84] wl[103] vdd gnd cell_6t
Xbit_r104_c84 bl[84] br[84] wl[104] vdd gnd cell_6t
Xbit_r105_c84 bl[84] br[84] wl[105] vdd gnd cell_6t
Xbit_r106_c84 bl[84] br[84] wl[106] vdd gnd cell_6t
Xbit_r107_c84 bl[84] br[84] wl[107] vdd gnd cell_6t
Xbit_r108_c84 bl[84] br[84] wl[108] vdd gnd cell_6t
Xbit_r109_c84 bl[84] br[84] wl[109] vdd gnd cell_6t
Xbit_r110_c84 bl[84] br[84] wl[110] vdd gnd cell_6t
Xbit_r111_c84 bl[84] br[84] wl[111] vdd gnd cell_6t
Xbit_r112_c84 bl[84] br[84] wl[112] vdd gnd cell_6t
Xbit_r113_c84 bl[84] br[84] wl[113] vdd gnd cell_6t
Xbit_r114_c84 bl[84] br[84] wl[114] vdd gnd cell_6t
Xbit_r115_c84 bl[84] br[84] wl[115] vdd gnd cell_6t
Xbit_r116_c84 bl[84] br[84] wl[116] vdd gnd cell_6t
Xbit_r117_c84 bl[84] br[84] wl[117] vdd gnd cell_6t
Xbit_r118_c84 bl[84] br[84] wl[118] vdd gnd cell_6t
Xbit_r119_c84 bl[84] br[84] wl[119] vdd gnd cell_6t
Xbit_r120_c84 bl[84] br[84] wl[120] vdd gnd cell_6t
Xbit_r121_c84 bl[84] br[84] wl[121] vdd gnd cell_6t
Xbit_r122_c84 bl[84] br[84] wl[122] vdd gnd cell_6t
Xbit_r123_c84 bl[84] br[84] wl[123] vdd gnd cell_6t
Xbit_r124_c84 bl[84] br[84] wl[124] vdd gnd cell_6t
Xbit_r125_c84 bl[84] br[84] wl[125] vdd gnd cell_6t
Xbit_r126_c84 bl[84] br[84] wl[126] vdd gnd cell_6t
Xbit_r127_c84 bl[84] br[84] wl[127] vdd gnd cell_6t
Xbit_r128_c84 bl[84] br[84] wl[128] vdd gnd cell_6t
Xbit_r129_c84 bl[84] br[84] wl[129] vdd gnd cell_6t
Xbit_r130_c84 bl[84] br[84] wl[130] vdd gnd cell_6t
Xbit_r131_c84 bl[84] br[84] wl[131] vdd gnd cell_6t
Xbit_r132_c84 bl[84] br[84] wl[132] vdd gnd cell_6t
Xbit_r133_c84 bl[84] br[84] wl[133] vdd gnd cell_6t
Xbit_r134_c84 bl[84] br[84] wl[134] vdd gnd cell_6t
Xbit_r135_c84 bl[84] br[84] wl[135] vdd gnd cell_6t
Xbit_r136_c84 bl[84] br[84] wl[136] vdd gnd cell_6t
Xbit_r137_c84 bl[84] br[84] wl[137] vdd gnd cell_6t
Xbit_r138_c84 bl[84] br[84] wl[138] vdd gnd cell_6t
Xbit_r139_c84 bl[84] br[84] wl[139] vdd gnd cell_6t
Xbit_r140_c84 bl[84] br[84] wl[140] vdd gnd cell_6t
Xbit_r141_c84 bl[84] br[84] wl[141] vdd gnd cell_6t
Xbit_r142_c84 bl[84] br[84] wl[142] vdd gnd cell_6t
Xbit_r143_c84 bl[84] br[84] wl[143] vdd gnd cell_6t
Xbit_r144_c84 bl[84] br[84] wl[144] vdd gnd cell_6t
Xbit_r145_c84 bl[84] br[84] wl[145] vdd gnd cell_6t
Xbit_r146_c84 bl[84] br[84] wl[146] vdd gnd cell_6t
Xbit_r147_c84 bl[84] br[84] wl[147] vdd gnd cell_6t
Xbit_r148_c84 bl[84] br[84] wl[148] vdd gnd cell_6t
Xbit_r149_c84 bl[84] br[84] wl[149] vdd gnd cell_6t
Xbit_r150_c84 bl[84] br[84] wl[150] vdd gnd cell_6t
Xbit_r151_c84 bl[84] br[84] wl[151] vdd gnd cell_6t
Xbit_r152_c84 bl[84] br[84] wl[152] vdd gnd cell_6t
Xbit_r153_c84 bl[84] br[84] wl[153] vdd gnd cell_6t
Xbit_r154_c84 bl[84] br[84] wl[154] vdd gnd cell_6t
Xbit_r155_c84 bl[84] br[84] wl[155] vdd gnd cell_6t
Xbit_r156_c84 bl[84] br[84] wl[156] vdd gnd cell_6t
Xbit_r157_c84 bl[84] br[84] wl[157] vdd gnd cell_6t
Xbit_r158_c84 bl[84] br[84] wl[158] vdd gnd cell_6t
Xbit_r159_c84 bl[84] br[84] wl[159] vdd gnd cell_6t
Xbit_r160_c84 bl[84] br[84] wl[160] vdd gnd cell_6t
Xbit_r161_c84 bl[84] br[84] wl[161] vdd gnd cell_6t
Xbit_r162_c84 bl[84] br[84] wl[162] vdd gnd cell_6t
Xbit_r163_c84 bl[84] br[84] wl[163] vdd gnd cell_6t
Xbit_r164_c84 bl[84] br[84] wl[164] vdd gnd cell_6t
Xbit_r165_c84 bl[84] br[84] wl[165] vdd gnd cell_6t
Xbit_r166_c84 bl[84] br[84] wl[166] vdd gnd cell_6t
Xbit_r167_c84 bl[84] br[84] wl[167] vdd gnd cell_6t
Xbit_r168_c84 bl[84] br[84] wl[168] vdd gnd cell_6t
Xbit_r169_c84 bl[84] br[84] wl[169] vdd gnd cell_6t
Xbit_r170_c84 bl[84] br[84] wl[170] vdd gnd cell_6t
Xbit_r171_c84 bl[84] br[84] wl[171] vdd gnd cell_6t
Xbit_r172_c84 bl[84] br[84] wl[172] vdd gnd cell_6t
Xbit_r173_c84 bl[84] br[84] wl[173] vdd gnd cell_6t
Xbit_r174_c84 bl[84] br[84] wl[174] vdd gnd cell_6t
Xbit_r175_c84 bl[84] br[84] wl[175] vdd gnd cell_6t
Xbit_r176_c84 bl[84] br[84] wl[176] vdd gnd cell_6t
Xbit_r177_c84 bl[84] br[84] wl[177] vdd gnd cell_6t
Xbit_r178_c84 bl[84] br[84] wl[178] vdd gnd cell_6t
Xbit_r179_c84 bl[84] br[84] wl[179] vdd gnd cell_6t
Xbit_r180_c84 bl[84] br[84] wl[180] vdd gnd cell_6t
Xbit_r181_c84 bl[84] br[84] wl[181] vdd gnd cell_6t
Xbit_r182_c84 bl[84] br[84] wl[182] vdd gnd cell_6t
Xbit_r183_c84 bl[84] br[84] wl[183] vdd gnd cell_6t
Xbit_r184_c84 bl[84] br[84] wl[184] vdd gnd cell_6t
Xbit_r185_c84 bl[84] br[84] wl[185] vdd gnd cell_6t
Xbit_r186_c84 bl[84] br[84] wl[186] vdd gnd cell_6t
Xbit_r187_c84 bl[84] br[84] wl[187] vdd gnd cell_6t
Xbit_r188_c84 bl[84] br[84] wl[188] vdd gnd cell_6t
Xbit_r189_c84 bl[84] br[84] wl[189] vdd gnd cell_6t
Xbit_r190_c84 bl[84] br[84] wl[190] vdd gnd cell_6t
Xbit_r191_c84 bl[84] br[84] wl[191] vdd gnd cell_6t
Xbit_r192_c84 bl[84] br[84] wl[192] vdd gnd cell_6t
Xbit_r193_c84 bl[84] br[84] wl[193] vdd gnd cell_6t
Xbit_r194_c84 bl[84] br[84] wl[194] vdd gnd cell_6t
Xbit_r195_c84 bl[84] br[84] wl[195] vdd gnd cell_6t
Xbit_r196_c84 bl[84] br[84] wl[196] vdd gnd cell_6t
Xbit_r197_c84 bl[84] br[84] wl[197] vdd gnd cell_6t
Xbit_r198_c84 bl[84] br[84] wl[198] vdd gnd cell_6t
Xbit_r199_c84 bl[84] br[84] wl[199] vdd gnd cell_6t
Xbit_r200_c84 bl[84] br[84] wl[200] vdd gnd cell_6t
Xbit_r201_c84 bl[84] br[84] wl[201] vdd gnd cell_6t
Xbit_r202_c84 bl[84] br[84] wl[202] vdd gnd cell_6t
Xbit_r203_c84 bl[84] br[84] wl[203] vdd gnd cell_6t
Xbit_r204_c84 bl[84] br[84] wl[204] vdd gnd cell_6t
Xbit_r205_c84 bl[84] br[84] wl[205] vdd gnd cell_6t
Xbit_r206_c84 bl[84] br[84] wl[206] vdd gnd cell_6t
Xbit_r207_c84 bl[84] br[84] wl[207] vdd gnd cell_6t
Xbit_r208_c84 bl[84] br[84] wl[208] vdd gnd cell_6t
Xbit_r209_c84 bl[84] br[84] wl[209] vdd gnd cell_6t
Xbit_r210_c84 bl[84] br[84] wl[210] vdd gnd cell_6t
Xbit_r211_c84 bl[84] br[84] wl[211] vdd gnd cell_6t
Xbit_r212_c84 bl[84] br[84] wl[212] vdd gnd cell_6t
Xbit_r213_c84 bl[84] br[84] wl[213] vdd gnd cell_6t
Xbit_r214_c84 bl[84] br[84] wl[214] vdd gnd cell_6t
Xbit_r215_c84 bl[84] br[84] wl[215] vdd gnd cell_6t
Xbit_r216_c84 bl[84] br[84] wl[216] vdd gnd cell_6t
Xbit_r217_c84 bl[84] br[84] wl[217] vdd gnd cell_6t
Xbit_r218_c84 bl[84] br[84] wl[218] vdd gnd cell_6t
Xbit_r219_c84 bl[84] br[84] wl[219] vdd gnd cell_6t
Xbit_r220_c84 bl[84] br[84] wl[220] vdd gnd cell_6t
Xbit_r221_c84 bl[84] br[84] wl[221] vdd gnd cell_6t
Xbit_r222_c84 bl[84] br[84] wl[222] vdd gnd cell_6t
Xbit_r223_c84 bl[84] br[84] wl[223] vdd gnd cell_6t
Xbit_r224_c84 bl[84] br[84] wl[224] vdd gnd cell_6t
Xbit_r225_c84 bl[84] br[84] wl[225] vdd gnd cell_6t
Xbit_r226_c84 bl[84] br[84] wl[226] vdd gnd cell_6t
Xbit_r227_c84 bl[84] br[84] wl[227] vdd gnd cell_6t
Xbit_r228_c84 bl[84] br[84] wl[228] vdd gnd cell_6t
Xbit_r229_c84 bl[84] br[84] wl[229] vdd gnd cell_6t
Xbit_r230_c84 bl[84] br[84] wl[230] vdd gnd cell_6t
Xbit_r231_c84 bl[84] br[84] wl[231] vdd gnd cell_6t
Xbit_r232_c84 bl[84] br[84] wl[232] vdd gnd cell_6t
Xbit_r233_c84 bl[84] br[84] wl[233] vdd gnd cell_6t
Xbit_r234_c84 bl[84] br[84] wl[234] vdd gnd cell_6t
Xbit_r235_c84 bl[84] br[84] wl[235] vdd gnd cell_6t
Xbit_r236_c84 bl[84] br[84] wl[236] vdd gnd cell_6t
Xbit_r237_c84 bl[84] br[84] wl[237] vdd gnd cell_6t
Xbit_r238_c84 bl[84] br[84] wl[238] vdd gnd cell_6t
Xbit_r239_c84 bl[84] br[84] wl[239] vdd gnd cell_6t
Xbit_r240_c84 bl[84] br[84] wl[240] vdd gnd cell_6t
Xbit_r241_c84 bl[84] br[84] wl[241] vdd gnd cell_6t
Xbit_r242_c84 bl[84] br[84] wl[242] vdd gnd cell_6t
Xbit_r243_c84 bl[84] br[84] wl[243] vdd gnd cell_6t
Xbit_r244_c84 bl[84] br[84] wl[244] vdd gnd cell_6t
Xbit_r245_c84 bl[84] br[84] wl[245] vdd gnd cell_6t
Xbit_r246_c84 bl[84] br[84] wl[246] vdd gnd cell_6t
Xbit_r247_c84 bl[84] br[84] wl[247] vdd gnd cell_6t
Xbit_r248_c84 bl[84] br[84] wl[248] vdd gnd cell_6t
Xbit_r249_c84 bl[84] br[84] wl[249] vdd gnd cell_6t
Xbit_r250_c84 bl[84] br[84] wl[250] vdd gnd cell_6t
Xbit_r251_c84 bl[84] br[84] wl[251] vdd gnd cell_6t
Xbit_r252_c84 bl[84] br[84] wl[252] vdd gnd cell_6t
Xbit_r253_c84 bl[84] br[84] wl[253] vdd gnd cell_6t
Xbit_r254_c84 bl[84] br[84] wl[254] vdd gnd cell_6t
Xbit_r255_c84 bl[84] br[84] wl[255] vdd gnd cell_6t
Xbit_r0_c85 bl[85] br[85] wl[0] vdd gnd cell_6t
Xbit_r1_c85 bl[85] br[85] wl[1] vdd gnd cell_6t
Xbit_r2_c85 bl[85] br[85] wl[2] vdd gnd cell_6t
Xbit_r3_c85 bl[85] br[85] wl[3] vdd gnd cell_6t
Xbit_r4_c85 bl[85] br[85] wl[4] vdd gnd cell_6t
Xbit_r5_c85 bl[85] br[85] wl[5] vdd gnd cell_6t
Xbit_r6_c85 bl[85] br[85] wl[6] vdd gnd cell_6t
Xbit_r7_c85 bl[85] br[85] wl[7] vdd gnd cell_6t
Xbit_r8_c85 bl[85] br[85] wl[8] vdd gnd cell_6t
Xbit_r9_c85 bl[85] br[85] wl[9] vdd gnd cell_6t
Xbit_r10_c85 bl[85] br[85] wl[10] vdd gnd cell_6t
Xbit_r11_c85 bl[85] br[85] wl[11] vdd gnd cell_6t
Xbit_r12_c85 bl[85] br[85] wl[12] vdd gnd cell_6t
Xbit_r13_c85 bl[85] br[85] wl[13] vdd gnd cell_6t
Xbit_r14_c85 bl[85] br[85] wl[14] vdd gnd cell_6t
Xbit_r15_c85 bl[85] br[85] wl[15] vdd gnd cell_6t
Xbit_r16_c85 bl[85] br[85] wl[16] vdd gnd cell_6t
Xbit_r17_c85 bl[85] br[85] wl[17] vdd gnd cell_6t
Xbit_r18_c85 bl[85] br[85] wl[18] vdd gnd cell_6t
Xbit_r19_c85 bl[85] br[85] wl[19] vdd gnd cell_6t
Xbit_r20_c85 bl[85] br[85] wl[20] vdd gnd cell_6t
Xbit_r21_c85 bl[85] br[85] wl[21] vdd gnd cell_6t
Xbit_r22_c85 bl[85] br[85] wl[22] vdd gnd cell_6t
Xbit_r23_c85 bl[85] br[85] wl[23] vdd gnd cell_6t
Xbit_r24_c85 bl[85] br[85] wl[24] vdd gnd cell_6t
Xbit_r25_c85 bl[85] br[85] wl[25] vdd gnd cell_6t
Xbit_r26_c85 bl[85] br[85] wl[26] vdd gnd cell_6t
Xbit_r27_c85 bl[85] br[85] wl[27] vdd gnd cell_6t
Xbit_r28_c85 bl[85] br[85] wl[28] vdd gnd cell_6t
Xbit_r29_c85 bl[85] br[85] wl[29] vdd gnd cell_6t
Xbit_r30_c85 bl[85] br[85] wl[30] vdd gnd cell_6t
Xbit_r31_c85 bl[85] br[85] wl[31] vdd gnd cell_6t
Xbit_r32_c85 bl[85] br[85] wl[32] vdd gnd cell_6t
Xbit_r33_c85 bl[85] br[85] wl[33] vdd gnd cell_6t
Xbit_r34_c85 bl[85] br[85] wl[34] vdd gnd cell_6t
Xbit_r35_c85 bl[85] br[85] wl[35] vdd gnd cell_6t
Xbit_r36_c85 bl[85] br[85] wl[36] vdd gnd cell_6t
Xbit_r37_c85 bl[85] br[85] wl[37] vdd gnd cell_6t
Xbit_r38_c85 bl[85] br[85] wl[38] vdd gnd cell_6t
Xbit_r39_c85 bl[85] br[85] wl[39] vdd gnd cell_6t
Xbit_r40_c85 bl[85] br[85] wl[40] vdd gnd cell_6t
Xbit_r41_c85 bl[85] br[85] wl[41] vdd gnd cell_6t
Xbit_r42_c85 bl[85] br[85] wl[42] vdd gnd cell_6t
Xbit_r43_c85 bl[85] br[85] wl[43] vdd gnd cell_6t
Xbit_r44_c85 bl[85] br[85] wl[44] vdd gnd cell_6t
Xbit_r45_c85 bl[85] br[85] wl[45] vdd gnd cell_6t
Xbit_r46_c85 bl[85] br[85] wl[46] vdd gnd cell_6t
Xbit_r47_c85 bl[85] br[85] wl[47] vdd gnd cell_6t
Xbit_r48_c85 bl[85] br[85] wl[48] vdd gnd cell_6t
Xbit_r49_c85 bl[85] br[85] wl[49] vdd gnd cell_6t
Xbit_r50_c85 bl[85] br[85] wl[50] vdd gnd cell_6t
Xbit_r51_c85 bl[85] br[85] wl[51] vdd gnd cell_6t
Xbit_r52_c85 bl[85] br[85] wl[52] vdd gnd cell_6t
Xbit_r53_c85 bl[85] br[85] wl[53] vdd gnd cell_6t
Xbit_r54_c85 bl[85] br[85] wl[54] vdd gnd cell_6t
Xbit_r55_c85 bl[85] br[85] wl[55] vdd gnd cell_6t
Xbit_r56_c85 bl[85] br[85] wl[56] vdd gnd cell_6t
Xbit_r57_c85 bl[85] br[85] wl[57] vdd gnd cell_6t
Xbit_r58_c85 bl[85] br[85] wl[58] vdd gnd cell_6t
Xbit_r59_c85 bl[85] br[85] wl[59] vdd gnd cell_6t
Xbit_r60_c85 bl[85] br[85] wl[60] vdd gnd cell_6t
Xbit_r61_c85 bl[85] br[85] wl[61] vdd gnd cell_6t
Xbit_r62_c85 bl[85] br[85] wl[62] vdd gnd cell_6t
Xbit_r63_c85 bl[85] br[85] wl[63] vdd gnd cell_6t
Xbit_r64_c85 bl[85] br[85] wl[64] vdd gnd cell_6t
Xbit_r65_c85 bl[85] br[85] wl[65] vdd gnd cell_6t
Xbit_r66_c85 bl[85] br[85] wl[66] vdd gnd cell_6t
Xbit_r67_c85 bl[85] br[85] wl[67] vdd gnd cell_6t
Xbit_r68_c85 bl[85] br[85] wl[68] vdd gnd cell_6t
Xbit_r69_c85 bl[85] br[85] wl[69] vdd gnd cell_6t
Xbit_r70_c85 bl[85] br[85] wl[70] vdd gnd cell_6t
Xbit_r71_c85 bl[85] br[85] wl[71] vdd gnd cell_6t
Xbit_r72_c85 bl[85] br[85] wl[72] vdd gnd cell_6t
Xbit_r73_c85 bl[85] br[85] wl[73] vdd gnd cell_6t
Xbit_r74_c85 bl[85] br[85] wl[74] vdd gnd cell_6t
Xbit_r75_c85 bl[85] br[85] wl[75] vdd gnd cell_6t
Xbit_r76_c85 bl[85] br[85] wl[76] vdd gnd cell_6t
Xbit_r77_c85 bl[85] br[85] wl[77] vdd gnd cell_6t
Xbit_r78_c85 bl[85] br[85] wl[78] vdd gnd cell_6t
Xbit_r79_c85 bl[85] br[85] wl[79] vdd gnd cell_6t
Xbit_r80_c85 bl[85] br[85] wl[80] vdd gnd cell_6t
Xbit_r81_c85 bl[85] br[85] wl[81] vdd gnd cell_6t
Xbit_r82_c85 bl[85] br[85] wl[82] vdd gnd cell_6t
Xbit_r83_c85 bl[85] br[85] wl[83] vdd gnd cell_6t
Xbit_r84_c85 bl[85] br[85] wl[84] vdd gnd cell_6t
Xbit_r85_c85 bl[85] br[85] wl[85] vdd gnd cell_6t
Xbit_r86_c85 bl[85] br[85] wl[86] vdd gnd cell_6t
Xbit_r87_c85 bl[85] br[85] wl[87] vdd gnd cell_6t
Xbit_r88_c85 bl[85] br[85] wl[88] vdd gnd cell_6t
Xbit_r89_c85 bl[85] br[85] wl[89] vdd gnd cell_6t
Xbit_r90_c85 bl[85] br[85] wl[90] vdd gnd cell_6t
Xbit_r91_c85 bl[85] br[85] wl[91] vdd gnd cell_6t
Xbit_r92_c85 bl[85] br[85] wl[92] vdd gnd cell_6t
Xbit_r93_c85 bl[85] br[85] wl[93] vdd gnd cell_6t
Xbit_r94_c85 bl[85] br[85] wl[94] vdd gnd cell_6t
Xbit_r95_c85 bl[85] br[85] wl[95] vdd gnd cell_6t
Xbit_r96_c85 bl[85] br[85] wl[96] vdd gnd cell_6t
Xbit_r97_c85 bl[85] br[85] wl[97] vdd gnd cell_6t
Xbit_r98_c85 bl[85] br[85] wl[98] vdd gnd cell_6t
Xbit_r99_c85 bl[85] br[85] wl[99] vdd gnd cell_6t
Xbit_r100_c85 bl[85] br[85] wl[100] vdd gnd cell_6t
Xbit_r101_c85 bl[85] br[85] wl[101] vdd gnd cell_6t
Xbit_r102_c85 bl[85] br[85] wl[102] vdd gnd cell_6t
Xbit_r103_c85 bl[85] br[85] wl[103] vdd gnd cell_6t
Xbit_r104_c85 bl[85] br[85] wl[104] vdd gnd cell_6t
Xbit_r105_c85 bl[85] br[85] wl[105] vdd gnd cell_6t
Xbit_r106_c85 bl[85] br[85] wl[106] vdd gnd cell_6t
Xbit_r107_c85 bl[85] br[85] wl[107] vdd gnd cell_6t
Xbit_r108_c85 bl[85] br[85] wl[108] vdd gnd cell_6t
Xbit_r109_c85 bl[85] br[85] wl[109] vdd gnd cell_6t
Xbit_r110_c85 bl[85] br[85] wl[110] vdd gnd cell_6t
Xbit_r111_c85 bl[85] br[85] wl[111] vdd gnd cell_6t
Xbit_r112_c85 bl[85] br[85] wl[112] vdd gnd cell_6t
Xbit_r113_c85 bl[85] br[85] wl[113] vdd gnd cell_6t
Xbit_r114_c85 bl[85] br[85] wl[114] vdd gnd cell_6t
Xbit_r115_c85 bl[85] br[85] wl[115] vdd gnd cell_6t
Xbit_r116_c85 bl[85] br[85] wl[116] vdd gnd cell_6t
Xbit_r117_c85 bl[85] br[85] wl[117] vdd gnd cell_6t
Xbit_r118_c85 bl[85] br[85] wl[118] vdd gnd cell_6t
Xbit_r119_c85 bl[85] br[85] wl[119] vdd gnd cell_6t
Xbit_r120_c85 bl[85] br[85] wl[120] vdd gnd cell_6t
Xbit_r121_c85 bl[85] br[85] wl[121] vdd gnd cell_6t
Xbit_r122_c85 bl[85] br[85] wl[122] vdd gnd cell_6t
Xbit_r123_c85 bl[85] br[85] wl[123] vdd gnd cell_6t
Xbit_r124_c85 bl[85] br[85] wl[124] vdd gnd cell_6t
Xbit_r125_c85 bl[85] br[85] wl[125] vdd gnd cell_6t
Xbit_r126_c85 bl[85] br[85] wl[126] vdd gnd cell_6t
Xbit_r127_c85 bl[85] br[85] wl[127] vdd gnd cell_6t
Xbit_r128_c85 bl[85] br[85] wl[128] vdd gnd cell_6t
Xbit_r129_c85 bl[85] br[85] wl[129] vdd gnd cell_6t
Xbit_r130_c85 bl[85] br[85] wl[130] vdd gnd cell_6t
Xbit_r131_c85 bl[85] br[85] wl[131] vdd gnd cell_6t
Xbit_r132_c85 bl[85] br[85] wl[132] vdd gnd cell_6t
Xbit_r133_c85 bl[85] br[85] wl[133] vdd gnd cell_6t
Xbit_r134_c85 bl[85] br[85] wl[134] vdd gnd cell_6t
Xbit_r135_c85 bl[85] br[85] wl[135] vdd gnd cell_6t
Xbit_r136_c85 bl[85] br[85] wl[136] vdd gnd cell_6t
Xbit_r137_c85 bl[85] br[85] wl[137] vdd gnd cell_6t
Xbit_r138_c85 bl[85] br[85] wl[138] vdd gnd cell_6t
Xbit_r139_c85 bl[85] br[85] wl[139] vdd gnd cell_6t
Xbit_r140_c85 bl[85] br[85] wl[140] vdd gnd cell_6t
Xbit_r141_c85 bl[85] br[85] wl[141] vdd gnd cell_6t
Xbit_r142_c85 bl[85] br[85] wl[142] vdd gnd cell_6t
Xbit_r143_c85 bl[85] br[85] wl[143] vdd gnd cell_6t
Xbit_r144_c85 bl[85] br[85] wl[144] vdd gnd cell_6t
Xbit_r145_c85 bl[85] br[85] wl[145] vdd gnd cell_6t
Xbit_r146_c85 bl[85] br[85] wl[146] vdd gnd cell_6t
Xbit_r147_c85 bl[85] br[85] wl[147] vdd gnd cell_6t
Xbit_r148_c85 bl[85] br[85] wl[148] vdd gnd cell_6t
Xbit_r149_c85 bl[85] br[85] wl[149] vdd gnd cell_6t
Xbit_r150_c85 bl[85] br[85] wl[150] vdd gnd cell_6t
Xbit_r151_c85 bl[85] br[85] wl[151] vdd gnd cell_6t
Xbit_r152_c85 bl[85] br[85] wl[152] vdd gnd cell_6t
Xbit_r153_c85 bl[85] br[85] wl[153] vdd gnd cell_6t
Xbit_r154_c85 bl[85] br[85] wl[154] vdd gnd cell_6t
Xbit_r155_c85 bl[85] br[85] wl[155] vdd gnd cell_6t
Xbit_r156_c85 bl[85] br[85] wl[156] vdd gnd cell_6t
Xbit_r157_c85 bl[85] br[85] wl[157] vdd gnd cell_6t
Xbit_r158_c85 bl[85] br[85] wl[158] vdd gnd cell_6t
Xbit_r159_c85 bl[85] br[85] wl[159] vdd gnd cell_6t
Xbit_r160_c85 bl[85] br[85] wl[160] vdd gnd cell_6t
Xbit_r161_c85 bl[85] br[85] wl[161] vdd gnd cell_6t
Xbit_r162_c85 bl[85] br[85] wl[162] vdd gnd cell_6t
Xbit_r163_c85 bl[85] br[85] wl[163] vdd gnd cell_6t
Xbit_r164_c85 bl[85] br[85] wl[164] vdd gnd cell_6t
Xbit_r165_c85 bl[85] br[85] wl[165] vdd gnd cell_6t
Xbit_r166_c85 bl[85] br[85] wl[166] vdd gnd cell_6t
Xbit_r167_c85 bl[85] br[85] wl[167] vdd gnd cell_6t
Xbit_r168_c85 bl[85] br[85] wl[168] vdd gnd cell_6t
Xbit_r169_c85 bl[85] br[85] wl[169] vdd gnd cell_6t
Xbit_r170_c85 bl[85] br[85] wl[170] vdd gnd cell_6t
Xbit_r171_c85 bl[85] br[85] wl[171] vdd gnd cell_6t
Xbit_r172_c85 bl[85] br[85] wl[172] vdd gnd cell_6t
Xbit_r173_c85 bl[85] br[85] wl[173] vdd gnd cell_6t
Xbit_r174_c85 bl[85] br[85] wl[174] vdd gnd cell_6t
Xbit_r175_c85 bl[85] br[85] wl[175] vdd gnd cell_6t
Xbit_r176_c85 bl[85] br[85] wl[176] vdd gnd cell_6t
Xbit_r177_c85 bl[85] br[85] wl[177] vdd gnd cell_6t
Xbit_r178_c85 bl[85] br[85] wl[178] vdd gnd cell_6t
Xbit_r179_c85 bl[85] br[85] wl[179] vdd gnd cell_6t
Xbit_r180_c85 bl[85] br[85] wl[180] vdd gnd cell_6t
Xbit_r181_c85 bl[85] br[85] wl[181] vdd gnd cell_6t
Xbit_r182_c85 bl[85] br[85] wl[182] vdd gnd cell_6t
Xbit_r183_c85 bl[85] br[85] wl[183] vdd gnd cell_6t
Xbit_r184_c85 bl[85] br[85] wl[184] vdd gnd cell_6t
Xbit_r185_c85 bl[85] br[85] wl[185] vdd gnd cell_6t
Xbit_r186_c85 bl[85] br[85] wl[186] vdd gnd cell_6t
Xbit_r187_c85 bl[85] br[85] wl[187] vdd gnd cell_6t
Xbit_r188_c85 bl[85] br[85] wl[188] vdd gnd cell_6t
Xbit_r189_c85 bl[85] br[85] wl[189] vdd gnd cell_6t
Xbit_r190_c85 bl[85] br[85] wl[190] vdd gnd cell_6t
Xbit_r191_c85 bl[85] br[85] wl[191] vdd gnd cell_6t
Xbit_r192_c85 bl[85] br[85] wl[192] vdd gnd cell_6t
Xbit_r193_c85 bl[85] br[85] wl[193] vdd gnd cell_6t
Xbit_r194_c85 bl[85] br[85] wl[194] vdd gnd cell_6t
Xbit_r195_c85 bl[85] br[85] wl[195] vdd gnd cell_6t
Xbit_r196_c85 bl[85] br[85] wl[196] vdd gnd cell_6t
Xbit_r197_c85 bl[85] br[85] wl[197] vdd gnd cell_6t
Xbit_r198_c85 bl[85] br[85] wl[198] vdd gnd cell_6t
Xbit_r199_c85 bl[85] br[85] wl[199] vdd gnd cell_6t
Xbit_r200_c85 bl[85] br[85] wl[200] vdd gnd cell_6t
Xbit_r201_c85 bl[85] br[85] wl[201] vdd gnd cell_6t
Xbit_r202_c85 bl[85] br[85] wl[202] vdd gnd cell_6t
Xbit_r203_c85 bl[85] br[85] wl[203] vdd gnd cell_6t
Xbit_r204_c85 bl[85] br[85] wl[204] vdd gnd cell_6t
Xbit_r205_c85 bl[85] br[85] wl[205] vdd gnd cell_6t
Xbit_r206_c85 bl[85] br[85] wl[206] vdd gnd cell_6t
Xbit_r207_c85 bl[85] br[85] wl[207] vdd gnd cell_6t
Xbit_r208_c85 bl[85] br[85] wl[208] vdd gnd cell_6t
Xbit_r209_c85 bl[85] br[85] wl[209] vdd gnd cell_6t
Xbit_r210_c85 bl[85] br[85] wl[210] vdd gnd cell_6t
Xbit_r211_c85 bl[85] br[85] wl[211] vdd gnd cell_6t
Xbit_r212_c85 bl[85] br[85] wl[212] vdd gnd cell_6t
Xbit_r213_c85 bl[85] br[85] wl[213] vdd gnd cell_6t
Xbit_r214_c85 bl[85] br[85] wl[214] vdd gnd cell_6t
Xbit_r215_c85 bl[85] br[85] wl[215] vdd gnd cell_6t
Xbit_r216_c85 bl[85] br[85] wl[216] vdd gnd cell_6t
Xbit_r217_c85 bl[85] br[85] wl[217] vdd gnd cell_6t
Xbit_r218_c85 bl[85] br[85] wl[218] vdd gnd cell_6t
Xbit_r219_c85 bl[85] br[85] wl[219] vdd gnd cell_6t
Xbit_r220_c85 bl[85] br[85] wl[220] vdd gnd cell_6t
Xbit_r221_c85 bl[85] br[85] wl[221] vdd gnd cell_6t
Xbit_r222_c85 bl[85] br[85] wl[222] vdd gnd cell_6t
Xbit_r223_c85 bl[85] br[85] wl[223] vdd gnd cell_6t
Xbit_r224_c85 bl[85] br[85] wl[224] vdd gnd cell_6t
Xbit_r225_c85 bl[85] br[85] wl[225] vdd gnd cell_6t
Xbit_r226_c85 bl[85] br[85] wl[226] vdd gnd cell_6t
Xbit_r227_c85 bl[85] br[85] wl[227] vdd gnd cell_6t
Xbit_r228_c85 bl[85] br[85] wl[228] vdd gnd cell_6t
Xbit_r229_c85 bl[85] br[85] wl[229] vdd gnd cell_6t
Xbit_r230_c85 bl[85] br[85] wl[230] vdd gnd cell_6t
Xbit_r231_c85 bl[85] br[85] wl[231] vdd gnd cell_6t
Xbit_r232_c85 bl[85] br[85] wl[232] vdd gnd cell_6t
Xbit_r233_c85 bl[85] br[85] wl[233] vdd gnd cell_6t
Xbit_r234_c85 bl[85] br[85] wl[234] vdd gnd cell_6t
Xbit_r235_c85 bl[85] br[85] wl[235] vdd gnd cell_6t
Xbit_r236_c85 bl[85] br[85] wl[236] vdd gnd cell_6t
Xbit_r237_c85 bl[85] br[85] wl[237] vdd gnd cell_6t
Xbit_r238_c85 bl[85] br[85] wl[238] vdd gnd cell_6t
Xbit_r239_c85 bl[85] br[85] wl[239] vdd gnd cell_6t
Xbit_r240_c85 bl[85] br[85] wl[240] vdd gnd cell_6t
Xbit_r241_c85 bl[85] br[85] wl[241] vdd gnd cell_6t
Xbit_r242_c85 bl[85] br[85] wl[242] vdd gnd cell_6t
Xbit_r243_c85 bl[85] br[85] wl[243] vdd gnd cell_6t
Xbit_r244_c85 bl[85] br[85] wl[244] vdd gnd cell_6t
Xbit_r245_c85 bl[85] br[85] wl[245] vdd gnd cell_6t
Xbit_r246_c85 bl[85] br[85] wl[246] vdd gnd cell_6t
Xbit_r247_c85 bl[85] br[85] wl[247] vdd gnd cell_6t
Xbit_r248_c85 bl[85] br[85] wl[248] vdd gnd cell_6t
Xbit_r249_c85 bl[85] br[85] wl[249] vdd gnd cell_6t
Xbit_r250_c85 bl[85] br[85] wl[250] vdd gnd cell_6t
Xbit_r251_c85 bl[85] br[85] wl[251] vdd gnd cell_6t
Xbit_r252_c85 bl[85] br[85] wl[252] vdd gnd cell_6t
Xbit_r253_c85 bl[85] br[85] wl[253] vdd gnd cell_6t
Xbit_r254_c85 bl[85] br[85] wl[254] vdd gnd cell_6t
Xbit_r255_c85 bl[85] br[85] wl[255] vdd gnd cell_6t
Xbit_r0_c86 bl[86] br[86] wl[0] vdd gnd cell_6t
Xbit_r1_c86 bl[86] br[86] wl[1] vdd gnd cell_6t
Xbit_r2_c86 bl[86] br[86] wl[2] vdd gnd cell_6t
Xbit_r3_c86 bl[86] br[86] wl[3] vdd gnd cell_6t
Xbit_r4_c86 bl[86] br[86] wl[4] vdd gnd cell_6t
Xbit_r5_c86 bl[86] br[86] wl[5] vdd gnd cell_6t
Xbit_r6_c86 bl[86] br[86] wl[6] vdd gnd cell_6t
Xbit_r7_c86 bl[86] br[86] wl[7] vdd gnd cell_6t
Xbit_r8_c86 bl[86] br[86] wl[8] vdd gnd cell_6t
Xbit_r9_c86 bl[86] br[86] wl[9] vdd gnd cell_6t
Xbit_r10_c86 bl[86] br[86] wl[10] vdd gnd cell_6t
Xbit_r11_c86 bl[86] br[86] wl[11] vdd gnd cell_6t
Xbit_r12_c86 bl[86] br[86] wl[12] vdd gnd cell_6t
Xbit_r13_c86 bl[86] br[86] wl[13] vdd gnd cell_6t
Xbit_r14_c86 bl[86] br[86] wl[14] vdd gnd cell_6t
Xbit_r15_c86 bl[86] br[86] wl[15] vdd gnd cell_6t
Xbit_r16_c86 bl[86] br[86] wl[16] vdd gnd cell_6t
Xbit_r17_c86 bl[86] br[86] wl[17] vdd gnd cell_6t
Xbit_r18_c86 bl[86] br[86] wl[18] vdd gnd cell_6t
Xbit_r19_c86 bl[86] br[86] wl[19] vdd gnd cell_6t
Xbit_r20_c86 bl[86] br[86] wl[20] vdd gnd cell_6t
Xbit_r21_c86 bl[86] br[86] wl[21] vdd gnd cell_6t
Xbit_r22_c86 bl[86] br[86] wl[22] vdd gnd cell_6t
Xbit_r23_c86 bl[86] br[86] wl[23] vdd gnd cell_6t
Xbit_r24_c86 bl[86] br[86] wl[24] vdd gnd cell_6t
Xbit_r25_c86 bl[86] br[86] wl[25] vdd gnd cell_6t
Xbit_r26_c86 bl[86] br[86] wl[26] vdd gnd cell_6t
Xbit_r27_c86 bl[86] br[86] wl[27] vdd gnd cell_6t
Xbit_r28_c86 bl[86] br[86] wl[28] vdd gnd cell_6t
Xbit_r29_c86 bl[86] br[86] wl[29] vdd gnd cell_6t
Xbit_r30_c86 bl[86] br[86] wl[30] vdd gnd cell_6t
Xbit_r31_c86 bl[86] br[86] wl[31] vdd gnd cell_6t
Xbit_r32_c86 bl[86] br[86] wl[32] vdd gnd cell_6t
Xbit_r33_c86 bl[86] br[86] wl[33] vdd gnd cell_6t
Xbit_r34_c86 bl[86] br[86] wl[34] vdd gnd cell_6t
Xbit_r35_c86 bl[86] br[86] wl[35] vdd gnd cell_6t
Xbit_r36_c86 bl[86] br[86] wl[36] vdd gnd cell_6t
Xbit_r37_c86 bl[86] br[86] wl[37] vdd gnd cell_6t
Xbit_r38_c86 bl[86] br[86] wl[38] vdd gnd cell_6t
Xbit_r39_c86 bl[86] br[86] wl[39] vdd gnd cell_6t
Xbit_r40_c86 bl[86] br[86] wl[40] vdd gnd cell_6t
Xbit_r41_c86 bl[86] br[86] wl[41] vdd gnd cell_6t
Xbit_r42_c86 bl[86] br[86] wl[42] vdd gnd cell_6t
Xbit_r43_c86 bl[86] br[86] wl[43] vdd gnd cell_6t
Xbit_r44_c86 bl[86] br[86] wl[44] vdd gnd cell_6t
Xbit_r45_c86 bl[86] br[86] wl[45] vdd gnd cell_6t
Xbit_r46_c86 bl[86] br[86] wl[46] vdd gnd cell_6t
Xbit_r47_c86 bl[86] br[86] wl[47] vdd gnd cell_6t
Xbit_r48_c86 bl[86] br[86] wl[48] vdd gnd cell_6t
Xbit_r49_c86 bl[86] br[86] wl[49] vdd gnd cell_6t
Xbit_r50_c86 bl[86] br[86] wl[50] vdd gnd cell_6t
Xbit_r51_c86 bl[86] br[86] wl[51] vdd gnd cell_6t
Xbit_r52_c86 bl[86] br[86] wl[52] vdd gnd cell_6t
Xbit_r53_c86 bl[86] br[86] wl[53] vdd gnd cell_6t
Xbit_r54_c86 bl[86] br[86] wl[54] vdd gnd cell_6t
Xbit_r55_c86 bl[86] br[86] wl[55] vdd gnd cell_6t
Xbit_r56_c86 bl[86] br[86] wl[56] vdd gnd cell_6t
Xbit_r57_c86 bl[86] br[86] wl[57] vdd gnd cell_6t
Xbit_r58_c86 bl[86] br[86] wl[58] vdd gnd cell_6t
Xbit_r59_c86 bl[86] br[86] wl[59] vdd gnd cell_6t
Xbit_r60_c86 bl[86] br[86] wl[60] vdd gnd cell_6t
Xbit_r61_c86 bl[86] br[86] wl[61] vdd gnd cell_6t
Xbit_r62_c86 bl[86] br[86] wl[62] vdd gnd cell_6t
Xbit_r63_c86 bl[86] br[86] wl[63] vdd gnd cell_6t
Xbit_r64_c86 bl[86] br[86] wl[64] vdd gnd cell_6t
Xbit_r65_c86 bl[86] br[86] wl[65] vdd gnd cell_6t
Xbit_r66_c86 bl[86] br[86] wl[66] vdd gnd cell_6t
Xbit_r67_c86 bl[86] br[86] wl[67] vdd gnd cell_6t
Xbit_r68_c86 bl[86] br[86] wl[68] vdd gnd cell_6t
Xbit_r69_c86 bl[86] br[86] wl[69] vdd gnd cell_6t
Xbit_r70_c86 bl[86] br[86] wl[70] vdd gnd cell_6t
Xbit_r71_c86 bl[86] br[86] wl[71] vdd gnd cell_6t
Xbit_r72_c86 bl[86] br[86] wl[72] vdd gnd cell_6t
Xbit_r73_c86 bl[86] br[86] wl[73] vdd gnd cell_6t
Xbit_r74_c86 bl[86] br[86] wl[74] vdd gnd cell_6t
Xbit_r75_c86 bl[86] br[86] wl[75] vdd gnd cell_6t
Xbit_r76_c86 bl[86] br[86] wl[76] vdd gnd cell_6t
Xbit_r77_c86 bl[86] br[86] wl[77] vdd gnd cell_6t
Xbit_r78_c86 bl[86] br[86] wl[78] vdd gnd cell_6t
Xbit_r79_c86 bl[86] br[86] wl[79] vdd gnd cell_6t
Xbit_r80_c86 bl[86] br[86] wl[80] vdd gnd cell_6t
Xbit_r81_c86 bl[86] br[86] wl[81] vdd gnd cell_6t
Xbit_r82_c86 bl[86] br[86] wl[82] vdd gnd cell_6t
Xbit_r83_c86 bl[86] br[86] wl[83] vdd gnd cell_6t
Xbit_r84_c86 bl[86] br[86] wl[84] vdd gnd cell_6t
Xbit_r85_c86 bl[86] br[86] wl[85] vdd gnd cell_6t
Xbit_r86_c86 bl[86] br[86] wl[86] vdd gnd cell_6t
Xbit_r87_c86 bl[86] br[86] wl[87] vdd gnd cell_6t
Xbit_r88_c86 bl[86] br[86] wl[88] vdd gnd cell_6t
Xbit_r89_c86 bl[86] br[86] wl[89] vdd gnd cell_6t
Xbit_r90_c86 bl[86] br[86] wl[90] vdd gnd cell_6t
Xbit_r91_c86 bl[86] br[86] wl[91] vdd gnd cell_6t
Xbit_r92_c86 bl[86] br[86] wl[92] vdd gnd cell_6t
Xbit_r93_c86 bl[86] br[86] wl[93] vdd gnd cell_6t
Xbit_r94_c86 bl[86] br[86] wl[94] vdd gnd cell_6t
Xbit_r95_c86 bl[86] br[86] wl[95] vdd gnd cell_6t
Xbit_r96_c86 bl[86] br[86] wl[96] vdd gnd cell_6t
Xbit_r97_c86 bl[86] br[86] wl[97] vdd gnd cell_6t
Xbit_r98_c86 bl[86] br[86] wl[98] vdd gnd cell_6t
Xbit_r99_c86 bl[86] br[86] wl[99] vdd gnd cell_6t
Xbit_r100_c86 bl[86] br[86] wl[100] vdd gnd cell_6t
Xbit_r101_c86 bl[86] br[86] wl[101] vdd gnd cell_6t
Xbit_r102_c86 bl[86] br[86] wl[102] vdd gnd cell_6t
Xbit_r103_c86 bl[86] br[86] wl[103] vdd gnd cell_6t
Xbit_r104_c86 bl[86] br[86] wl[104] vdd gnd cell_6t
Xbit_r105_c86 bl[86] br[86] wl[105] vdd gnd cell_6t
Xbit_r106_c86 bl[86] br[86] wl[106] vdd gnd cell_6t
Xbit_r107_c86 bl[86] br[86] wl[107] vdd gnd cell_6t
Xbit_r108_c86 bl[86] br[86] wl[108] vdd gnd cell_6t
Xbit_r109_c86 bl[86] br[86] wl[109] vdd gnd cell_6t
Xbit_r110_c86 bl[86] br[86] wl[110] vdd gnd cell_6t
Xbit_r111_c86 bl[86] br[86] wl[111] vdd gnd cell_6t
Xbit_r112_c86 bl[86] br[86] wl[112] vdd gnd cell_6t
Xbit_r113_c86 bl[86] br[86] wl[113] vdd gnd cell_6t
Xbit_r114_c86 bl[86] br[86] wl[114] vdd gnd cell_6t
Xbit_r115_c86 bl[86] br[86] wl[115] vdd gnd cell_6t
Xbit_r116_c86 bl[86] br[86] wl[116] vdd gnd cell_6t
Xbit_r117_c86 bl[86] br[86] wl[117] vdd gnd cell_6t
Xbit_r118_c86 bl[86] br[86] wl[118] vdd gnd cell_6t
Xbit_r119_c86 bl[86] br[86] wl[119] vdd gnd cell_6t
Xbit_r120_c86 bl[86] br[86] wl[120] vdd gnd cell_6t
Xbit_r121_c86 bl[86] br[86] wl[121] vdd gnd cell_6t
Xbit_r122_c86 bl[86] br[86] wl[122] vdd gnd cell_6t
Xbit_r123_c86 bl[86] br[86] wl[123] vdd gnd cell_6t
Xbit_r124_c86 bl[86] br[86] wl[124] vdd gnd cell_6t
Xbit_r125_c86 bl[86] br[86] wl[125] vdd gnd cell_6t
Xbit_r126_c86 bl[86] br[86] wl[126] vdd gnd cell_6t
Xbit_r127_c86 bl[86] br[86] wl[127] vdd gnd cell_6t
Xbit_r128_c86 bl[86] br[86] wl[128] vdd gnd cell_6t
Xbit_r129_c86 bl[86] br[86] wl[129] vdd gnd cell_6t
Xbit_r130_c86 bl[86] br[86] wl[130] vdd gnd cell_6t
Xbit_r131_c86 bl[86] br[86] wl[131] vdd gnd cell_6t
Xbit_r132_c86 bl[86] br[86] wl[132] vdd gnd cell_6t
Xbit_r133_c86 bl[86] br[86] wl[133] vdd gnd cell_6t
Xbit_r134_c86 bl[86] br[86] wl[134] vdd gnd cell_6t
Xbit_r135_c86 bl[86] br[86] wl[135] vdd gnd cell_6t
Xbit_r136_c86 bl[86] br[86] wl[136] vdd gnd cell_6t
Xbit_r137_c86 bl[86] br[86] wl[137] vdd gnd cell_6t
Xbit_r138_c86 bl[86] br[86] wl[138] vdd gnd cell_6t
Xbit_r139_c86 bl[86] br[86] wl[139] vdd gnd cell_6t
Xbit_r140_c86 bl[86] br[86] wl[140] vdd gnd cell_6t
Xbit_r141_c86 bl[86] br[86] wl[141] vdd gnd cell_6t
Xbit_r142_c86 bl[86] br[86] wl[142] vdd gnd cell_6t
Xbit_r143_c86 bl[86] br[86] wl[143] vdd gnd cell_6t
Xbit_r144_c86 bl[86] br[86] wl[144] vdd gnd cell_6t
Xbit_r145_c86 bl[86] br[86] wl[145] vdd gnd cell_6t
Xbit_r146_c86 bl[86] br[86] wl[146] vdd gnd cell_6t
Xbit_r147_c86 bl[86] br[86] wl[147] vdd gnd cell_6t
Xbit_r148_c86 bl[86] br[86] wl[148] vdd gnd cell_6t
Xbit_r149_c86 bl[86] br[86] wl[149] vdd gnd cell_6t
Xbit_r150_c86 bl[86] br[86] wl[150] vdd gnd cell_6t
Xbit_r151_c86 bl[86] br[86] wl[151] vdd gnd cell_6t
Xbit_r152_c86 bl[86] br[86] wl[152] vdd gnd cell_6t
Xbit_r153_c86 bl[86] br[86] wl[153] vdd gnd cell_6t
Xbit_r154_c86 bl[86] br[86] wl[154] vdd gnd cell_6t
Xbit_r155_c86 bl[86] br[86] wl[155] vdd gnd cell_6t
Xbit_r156_c86 bl[86] br[86] wl[156] vdd gnd cell_6t
Xbit_r157_c86 bl[86] br[86] wl[157] vdd gnd cell_6t
Xbit_r158_c86 bl[86] br[86] wl[158] vdd gnd cell_6t
Xbit_r159_c86 bl[86] br[86] wl[159] vdd gnd cell_6t
Xbit_r160_c86 bl[86] br[86] wl[160] vdd gnd cell_6t
Xbit_r161_c86 bl[86] br[86] wl[161] vdd gnd cell_6t
Xbit_r162_c86 bl[86] br[86] wl[162] vdd gnd cell_6t
Xbit_r163_c86 bl[86] br[86] wl[163] vdd gnd cell_6t
Xbit_r164_c86 bl[86] br[86] wl[164] vdd gnd cell_6t
Xbit_r165_c86 bl[86] br[86] wl[165] vdd gnd cell_6t
Xbit_r166_c86 bl[86] br[86] wl[166] vdd gnd cell_6t
Xbit_r167_c86 bl[86] br[86] wl[167] vdd gnd cell_6t
Xbit_r168_c86 bl[86] br[86] wl[168] vdd gnd cell_6t
Xbit_r169_c86 bl[86] br[86] wl[169] vdd gnd cell_6t
Xbit_r170_c86 bl[86] br[86] wl[170] vdd gnd cell_6t
Xbit_r171_c86 bl[86] br[86] wl[171] vdd gnd cell_6t
Xbit_r172_c86 bl[86] br[86] wl[172] vdd gnd cell_6t
Xbit_r173_c86 bl[86] br[86] wl[173] vdd gnd cell_6t
Xbit_r174_c86 bl[86] br[86] wl[174] vdd gnd cell_6t
Xbit_r175_c86 bl[86] br[86] wl[175] vdd gnd cell_6t
Xbit_r176_c86 bl[86] br[86] wl[176] vdd gnd cell_6t
Xbit_r177_c86 bl[86] br[86] wl[177] vdd gnd cell_6t
Xbit_r178_c86 bl[86] br[86] wl[178] vdd gnd cell_6t
Xbit_r179_c86 bl[86] br[86] wl[179] vdd gnd cell_6t
Xbit_r180_c86 bl[86] br[86] wl[180] vdd gnd cell_6t
Xbit_r181_c86 bl[86] br[86] wl[181] vdd gnd cell_6t
Xbit_r182_c86 bl[86] br[86] wl[182] vdd gnd cell_6t
Xbit_r183_c86 bl[86] br[86] wl[183] vdd gnd cell_6t
Xbit_r184_c86 bl[86] br[86] wl[184] vdd gnd cell_6t
Xbit_r185_c86 bl[86] br[86] wl[185] vdd gnd cell_6t
Xbit_r186_c86 bl[86] br[86] wl[186] vdd gnd cell_6t
Xbit_r187_c86 bl[86] br[86] wl[187] vdd gnd cell_6t
Xbit_r188_c86 bl[86] br[86] wl[188] vdd gnd cell_6t
Xbit_r189_c86 bl[86] br[86] wl[189] vdd gnd cell_6t
Xbit_r190_c86 bl[86] br[86] wl[190] vdd gnd cell_6t
Xbit_r191_c86 bl[86] br[86] wl[191] vdd gnd cell_6t
Xbit_r192_c86 bl[86] br[86] wl[192] vdd gnd cell_6t
Xbit_r193_c86 bl[86] br[86] wl[193] vdd gnd cell_6t
Xbit_r194_c86 bl[86] br[86] wl[194] vdd gnd cell_6t
Xbit_r195_c86 bl[86] br[86] wl[195] vdd gnd cell_6t
Xbit_r196_c86 bl[86] br[86] wl[196] vdd gnd cell_6t
Xbit_r197_c86 bl[86] br[86] wl[197] vdd gnd cell_6t
Xbit_r198_c86 bl[86] br[86] wl[198] vdd gnd cell_6t
Xbit_r199_c86 bl[86] br[86] wl[199] vdd gnd cell_6t
Xbit_r200_c86 bl[86] br[86] wl[200] vdd gnd cell_6t
Xbit_r201_c86 bl[86] br[86] wl[201] vdd gnd cell_6t
Xbit_r202_c86 bl[86] br[86] wl[202] vdd gnd cell_6t
Xbit_r203_c86 bl[86] br[86] wl[203] vdd gnd cell_6t
Xbit_r204_c86 bl[86] br[86] wl[204] vdd gnd cell_6t
Xbit_r205_c86 bl[86] br[86] wl[205] vdd gnd cell_6t
Xbit_r206_c86 bl[86] br[86] wl[206] vdd gnd cell_6t
Xbit_r207_c86 bl[86] br[86] wl[207] vdd gnd cell_6t
Xbit_r208_c86 bl[86] br[86] wl[208] vdd gnd cell_6t
Xbit_r209_c86 bl[86] br[86] wl[209] vdd gnd cell_6t
Xbit_r210_c86 bl[86] br[86] wl[210] vdd gnd cell_6t
Xbit_r211_c86 bl[86] br[86] wl[211] vdd gnd cell_6t
Xbit_r212_c86 bl[86] br[86] wl[212] vdd gnd cell_6t
Xbit_r213_c86 bl[86] br[86] wl[213] vdd gnd cell_6t
Xbit_r214_c86 bl[86] br[86] wl[214] vdd gnd cell_6t
Xbit_r215_c86 bl[86] br[86] wl[215] vdd gnd cell_6t
Xbit_r216_c86 bl[86] br[86] wl[216] vdd gnd cell_6t
Xbit_r217_c86 bl[86] br[86] wl[217] vdd gnd cell_6t
Xbit_r218_c86 bl[86] br[86] wl[218] vdd gnd cell_6t
Xbit_r219_c86 bl[86] br[86] wl[219] vdd gnd cell_6t
Xbit_r220_c86 bl[86] br[86] wl[220] vdd gnd cell_6t
Xbit_r221_c86 bl[86] br[86] wl[221] vdd gnd cell_6t
Xbit_r222_c86 bl[86] br[86] wl[222] vdd gnd cell_6t
Xbit_r223_c86 bl[86] br[86] wl[223] vdd gnd cell_6t
Xbit_r224_c86 bl[86] br[86] wl[224] vdd gnd cell_6t
Xbit_r225_c86 bl[86] br[86] wl[225] vdd gnd cell_6t
Xbit_r226_c86 bl[86] br[86] wl[226] vdd gnd cell_6t
Xbit_r227_c86 bl[86] br[86] wl[227] vdd gnd cell_6t
Xbit_r228_c86 bl[86] br[86] wl[228] vdd gnd cell_6t
Xbit_r229_c86 bl[86] br[86] wl[229] vdd gnd cell_6t
Xbit_r230_c86 bl[86] br[86] wl[230] vdd gnd cell_6t
Xbit_r231_c86 bl[86] br[86] wl[231] vdd gnd cell_6t
Xbit_r232_c86 bl[86] br[86] wl[232] vdd gnd cell_6t
Xbit_r233_c86 bl[86] br[86] wl[233] vdd gnd cell_6t
Xbit_r234_c86 bl[86] br[86] wl[234] vdd gnd cell_6t
Xbit_r235_c86 bl[86] br[86] wl[235] vdd gnd cell_6t
Xbit_r236_c86 bl[86] br[86] wl[236] vdd gnd cell_6t
Xbit_r237_c86 bl[86] br[86] wl[237] vdd gnd cell_6t
Xbit_r238_c86 bl[86] br[86] wl[238] vdd gnd cell_6t
Xbit_r239_c86 bl[86] br[86] wl[239] vdd gnd cell_6t
Xbit_r240_c86 bl[86] br[86] wl[240] vdd gnd cell_6t
Xbit_r241_c86 bl[86] br[86] wl[241] vdd gnd cell_6t
Xbit_r242_c86 bl[86] br[86] wl[242] vdd gnd cell_6t
Xbit_r243_c86 bl[86] br[86] wl[243] vdd gnd cell_6t
Xbit_r244_c86 bl[86] br[86] wl[244] vdd gnd cell_6t
Xbit_r245_c86 bl[86] br[86] wl[245] vdd gnd cell_6t
Xbit_r246_c86 bl[86] br[86] wl[246] vdd gnd cell_6t
Xbit_r247_c86 bl[86] br[86] wl[247] vdd gnd cell_6t
Xbit_r248_c86 bl[86] br[86] wl[248] vdd gnd cell_6t
Xbit_r249_c86 bl[86] br[86] wl[249] vdd gnd cell_6t
Xbit_r250_c86 bl[86] br[86] wl[250] vdd gnd cell_6t
Xbit_r251_c86 bl[86] br[86] wl[251] vdd gnd cell_6t
Xbit_r252_c86 bl[86] br[86] wl[252] vdd gnd cell_6t
Xbit_r253_c86 bl[86] br[86] wl[253] vdd gnd cell_6t
Xbit_r254_c86 bl[86] br[86] wl[254] vdd gnd cell_6t
Xbit_r255_c86 bl[86] br[86] wl[255] vdd gnd cell_6t
Xbit_r0_c87 bl[87] br[87] wl[0] vdd gnd cell_6t
Xbit_r1_c87 bl[87] br[87] wl[1] vdd gnd cell_6t
Xbit_r2_c87 bl[87] br[87] wl[2] vdd gnd cell_6t
Xbit_r3_c87 bl[87] br[87] wl[3] vdd gnd cell_6t
Xbit_r4_c87 bl[87] br[87] wl[4] vdd gnd cell_6t
Xbit_r5_c87 bl[87] br[87] wl[5] vdd gnd cell_6t
Xbit_r6_c87 bl[87] br[87] wl[6] vdd gnd cell_6t
Xbit_r7_c87 bl[87] br[87] wl[7] vdd gnd cell_6t
Xbit_r8_c87 bl[87] br[87] wl[8] vdd gnd cell_6t
Xbit_r9_c87 bl[87] br[87] wl[9] vdd gnd cell_6t
Xbit_r10_c87 bl[87] br[87] wl[10] vdd gnd cell_6t
Xbit_r11_c87 bl[87] br[87] wl[11] vdd gnd cell_6t
Xbit_r12_c87 bl[87] br[87] wl[12] vdd gnd cell_6t
Xbit_r13_c87 bl[87] br[87] wl[13] vdd gnd cell_6t
Xbit_r14_c87 bl[87] br[87] wl[14] vdd gnd cell_6t
Xbit_r15_c87 bl[87] br[87] wl[15] vdd gnd cell_6t
Xbit_r16_c87 bl[87] br[87] wl[16] vdd gnd cell_6t
Xbit_r17_c87 bl[87] br[87] wl[17] vdd gnd cell_6t
Xbit_r18_c87 bl[87] br[87] wl[18] vdd gnd cell_6t
Xbit_r19_c87 bl[87] br[87] wl[19] vdd gnd cell_6t
Xbit_r20_c87 bl[87] br[87] wl[20] vdd gnd cell_6t
Xbit_r21_c87 bl[87] br[87] wl[21] vdd gnd cell_6t
Xbit_r22_c87 bl[87] br[87] wl[22] vdd gnd cell_6t
Xbit_r23_c87 bl[87] br[87] wl[23] vdd gnd cell_6t
Xbit_r24_c87 bl[87] br[87] wl[24] vdd gnd cell_6t
Xbit_r25_c87 bl[87] br[87] wl[25] vdd gnd cell_6t
Xbit_r26_c87 bl[87] br[87] wl[26] vdd gnd cell_6t
Xbit_r27_c87 bl[87] br[87] wl[27] vdd gnd cell_6t
Xbit_r28_c87 bl[87] br[87] wl[28] vdd gnd cell_6t
Xbit_r29_c87 bl[87] br[87] wl[29] vdd gnd cell_6t
Xbit_r30_c87 bl[87] br[87] wl[30] vdd gnd cell_6t
Xbit_r31_c87 bl[87] br[87] wl[31] vdd gnd cell_6t
Xbit_r32_c87 bl[87] br[87] wl[32] vdd gnd cell_6t
Xbit_r33_c87 bl[87] br[87] wl[33] vdd gnd cell_6t
Xbit_r34_c87 bl[87] br[87] wl[34] vdd gnd cell_6t
Xbit_r35_c87 bl[87] br[87] wl[35] vdd gnd cell_6t
Xbit_r36_c87 bl[87] br[87] wl[36] vdd gnd cell_6t
Xbit_r37_c87 bl[87] br[87] wl[37] vdd gnd cell_6t
Xbit_r38_c87 bl[87] br[87] wl[38] vdd gnd cell_6t
Xbit_r39_c87 bl[87] br[87] wl[39] vdd gnd cell_6t
Xbit_r40_c87 bl[87] br[87] wl[40] vdd gnd cell_6t
Xbit_r41_c87 bl[87] br[87] wl[41] vdd gnd cell_6t
Xbit_r42_c87 bl[87] br[87] wl[42] vdd gnd cell_6t
Xbit_r43_c87 bl[87] br[87] wl[43] vdd gnd cell_6t
Xbit_r44_c87 bl[87] br[87] wl[44] vdd gnd cell_6t
Xbit_r45_c87 bl[87] br[87] wl[45] vdd gnd cell_6t
Xbit_r46_c87 bl[87] br[87] wl[46] vdd gnd cell_6t
Xbit_r47_c87 bl[87] br[87] wl[47] vdd gnd cell_6t
Xbit_r48_c87 bl[87] br[87] wl[48] vdd gnd cell_6t
Xbit_r49_c87 bl[87] br[87] wl[49] vdd gnd cell_6t
Xbit_r50_c87 bl[87] br[87] wl[50] vdd gnd cell_6t
Xbit_r51_c87 bl[87] br[87] wl[51] vdd gnd cell_6t
Xbit_r52_c87 bl[87] br[87] wl[52] vdd gnd cell_6t
Xbit_r53_c87 bl[87] br[87] wl[53] vdd gnd cell_6t
Xbit_r54_c87 bl[87] br[87] wl[54] vdd gnd cell_6t
Xbit_r55_c87 bl[87] br[87] wl[55] vdd gnd cell_6t
Xbit_r56_c87 bl[87] br[87] wl[56] vdd gnd cell_6t
Xbit_r57_c87 bl[87] br[87] wl[57] vdd gnd cell_6t
Xbit_r58_c87 bl[87] br[87] wl[58] vdd gnd cell_6t
Xbit_r59_c87 bl[87] br[87] wl[59] vdd gnd cell_6t
Xbit_r60_c87 bl[87] br[87] wl[60] vdd gnd cell_6t
Xbit_r61_c87 bl[87] br[87] wl[61] vdd gnd cell_6t
Xbit_r62_c87 bl[87] br[87] wl[62] vdd gnd cell_6t
Xbit_r63_c87 bl[87] br[87] wl[63] vdd gnd cell_6t
Xbit_r64_c87 bl[87] br[87] wl[64] vdd gnd cell_6t
Xbit_r65_c87 bl[87] br[87] wl[65] vdd gnd cell_6t
Xbit_r66_c87 bl[87] br[87] wl[66] vdd gnd cell_6t
Xbit_r67_c87 bl[87] br[87] wl[67] vdd gnd cell_6t
Xbit_r68_c87 bl[87] br[87] wl[68] vdd gnd cell_6t
Xbit_r69_c87 bl[87] br[87] wl[69] vdd gnd cell_6t
Xbit_r70_c87 bl[87] br[87] wl[70] vdd gnd cell_6t
Xbit_r71_c87 bl[87] br[87] wl[71] vdd gnd cell_6t
Xbit_r72_c87 bl[87] br[87] wl[72] vdd gnd cell_6t
Xbit_r73_c87 bl[87] br[87] wl[73] vdd gnd cell_6t
Xbit_r74_c87 bl[87] br[87] wl[74] vdd gnd cell_6t
Xbit_r75_c87 bl[87] br[87] wl[75] vdd gnd cell_6t
Xbit_r76_c87 bl[87] br[87] wl[76] vdd gnd cell_6t
Xbit_r77_c87 bl[87] br[87] wl[77] vdd gnd cell_6t
Xbit_r78_c87 bl[87] br[87] wl[78] vdd gnd cell_6t
Xbit_r79_c87 bl[87] br[87] wl[79] vdd gnd cell_6t
Xbit_r80_c87 bl[87] br[87] wl[80] vdd gnd cell_6t
Xbit_r81_c87 bl[87] br[87] wl[81] vdd gnd cell_6t
Xbit_r82_c87 bl[87] br[87] wl[82] vdd gnd cell_6t
Xbit_r83_c87 bl[87] br[87] wl[83] vdd gnd cell_6t
Xbit_r84_c87 bl[87] br[87] wl[84] vdd gnd cell_6t
Xbit_r85_c87 bl[87] br[87] wl[85] vdd gnd cell_6t
Xbit_r86_c87 bl[87] br[87] wl[86] vdd gnd cell_6t
Xbit_r87_c87 bl[87] br[87] wl[87] vdd gnd cell_6t
Xbit_r88_c87 bl[87] br[87] wl[88] vdd gnd cell_6t
Xbit_r89_c87 bl[87] br[87] wl[89] vdd gnd cell_6t
Xbit_r90_c87 bl[87] br[87] wl[90] vdd gnd cell_6t
Xbit_r91_c87 bl[87] br[87] wl[91] vdd gnd cell_6t
Xbit_r92_c87 bl[87] br[87] wl[92] vdd gnd cell_6t
Xbit_r93_c87 bl[87] br[87] wl[93] vdd gnd cell_6t
Xbit_r94_c87 bl[87] br[87] wl[94] vdd gnd cell_6t
Xbit_r95_c87 bl[87] br[87] wl[95] vdd gnd cell_6t
Xbit_r96_c87 bl[87] br[87] wl[96] vdd gnd cell_6t
Xbit_r97_c87 bl[87] br[87] wl[97] vdd gnd cell_6t
Xbit_r98_c87 bl[87] br[87] wl[98] vdd gnd cell_6t
Xbit_r99_c87 bl[87] br[87] wl[99] vdd gnd cell_6t
Xbit_r100_c87 bl[87] br[87] wl[100] vdd gnd cell_6t
Xbit_r101_c87 bl[87] br[87] wl[101] vdd gnd cell_6t
Xbit_r102_c87 bl[87] br[87] wl[102] vdd gnd cell_6t
Xbit_r103_c87 bl[87] br[87] wl[103] vdd gnd cell_6t
Xbit_r104_c87 bl[87] br[87] wl[104] vdd gnd cell_6t
Xbit_r105_c87 bl[87] br[87] wl[105] vdd gnd cell_6t
Xbit_r106_c87 bl[87] br[87] wl[106] vdd gnd cell_6t
Xbit_r107_c87 bl[87] br[87] wl[107] vdd gnd cell_6t
Xbit_r108_c87 bl[87] br[87] wl[108] vdd gnd cell_6t
Xbit_r109_c87 bl[87] br[87] wl[109] vdd gnd cell_6t
Xbit_r110_c87 bl[87] br[87] wl[110] vdd gnd cell_6t
Xbit_r111_c87 bl[87] br[87] wl[111] vdd gnd cell_6t
Xbit_r112_c87 bl[87] br[87] wl[112] vdd gnd cell_6t
Xbit_r113_c87 bl[87] br[87] wl[113] vdd gnd cell_6t
Xbit_r114_c87 bl[87] br[87] wl[114] vdd gnd cell_6t
Xbit_r115_c87 bl[87] br[87] wl[115] vdd gnd cell_6t
Xbit_r116_c87 bl[87] br[87] wl[116] vdd gnd cell_6t
Xbit_r117_c87 bl[87] br[87] wl[117] vdd gnd cell_6t
Xbit_r118_c87 bl[87] br[87] wl[118] vdd gnd cell_6t
Xbit_r119_c87 bl[87] br[87] wl[119] vdd gnd cell_6t
Xbit_r120_c87 bl[87] br[87] wl[120] vdd gnd cell_6t
Xbit_r121_c87 bl[87] br[87] wl[121] vdd gnd cell_6t
Xbit_r122_c87 bl[87] br[87] wl[122] vdd gnd cell_6t
Xbit_r123_c87 bl[87] br[87] wl[123] vdd gnd cell_6t
Xbit_r124_c87 bl[87] br[87] wl[124] vdd gnd cell_6t
Xbit_r125_c87 bl[87] br[87] wl[125] vdd gnd cell_6t
Xbit_r126_c87 bl[87] br[87] wl[126] vdd gnd cell_6t
Xbit_r127_c87 bl[87] br[87] wl[127] vdd gnd cell_6t
Xbit_r128_c87 bl[87] br[87] wl[128] vdd gnd cell_6t
Xbit_r129_c87 bl[87] br[87] wl[129] vdd gnd cell_6t
Xbit_r130_c87 bl[87] br[87] wl[130] vdd gnd cell_6t
Xbit_r131_c87 bl[87] br[87] wl[131] vdd gnd cell_6t
Xbit_r132_c87 bl[87] br[87] wl[132] vdd gnd cell_6t
Xbit_r133_c87 bl[87] br[87] wl[133] vdd gnd cell_6t
Xbit_r134_c87 bl[87] br[87] wl[134] vdd gnd cell_6t
Xbit_r135_c87 bl[87] br[87] wl[135] vdd gnd cell_6t
Xbit_r136_c87 bl[87] br[87] wl[136] vdd gnd cell_6t
Xbit_r137_c87 bl[87] br[87] wl[137] vdd gnd cell_6t
Xbit_r138_c87 bl[87] br[87] wl[138] vdd gnd cell_6t
Xbit_r139_c87 bl[87] br[87] wl[139] vdd gnd cell_6t
Xbit_r140_c87 bl[87] br[87] wl[140] vdd gnd cell_6t
Xbit_r141_c87 bl[87] br[87] wl[141] vdd gnd cell_6t
Xbit_r142_c87 bl[87] br[87] wl[142] vdd gnd cell_6t
Xbit_r143_c87 bl[87] br[87] wl[143] vdd gnd cell_6t
Xbit_r144_c87 bl[87] br[87] wl[144] vdd gnd cell_6t
Xbit_r145_c87 bl[87] br[87] wl[145] vdd gnd cell_6t
Xbit_r146_c87 bl[87] br[87] wl[146] vdd gnd cell_6t
Xbit_r147_c87 bl[87] br[87] wl[147] vdd gnd cell_6t
Xbit_r148_c87 bl[87] br[87] wl[148] vdd gnd cell_6t
Xbit_r149_c87 bl[87] br[87] wl[149] vdd gnd cell_6t
Xbit_r150_c87 bl[87] br[87] wl[150] vdd gnd cell_6t
Xbit_r151_c87 bl[87] br[87] wl[151] vdd gnd cell_6t
Xbit_r152_c87 bl[87] br[87] wl[152] vdd gnd cell_6t
Xbit_r153_c87 bl[87] br[87] wl[153] vdd gnd cell_6t
Xbit_r154_c87 bl[87] br[87] wl[154] vdd gnd cell_6t
Xbit_r155_c87 bl[87] br[87] wl[155] vdd gnd cell_6t
Xbit_r156_c87 bl[87] br[87] wl[156] vdd gnd cell_6t
Xbit_r157_c87 bl[87] br[87] wl[157] vdd gnd cell_6t
Xbit_r158_c87 bl[87] br[87] wl[158] vdd gnd cell_6t
Xbit_r159_c87 bl[87] br[87] wl[159] vdd gnd cell_6t
Xbit_r160_c87 bl[87] br[87] wl[160] vdd gnd cell_6t
Xbit_r161_c87 bl[87] br[87] wl[161] vdd gnd cell_6t
Xbit_r162_c87 bl[87] br[87] wl[162] vdd gnd cell_6t
Xbit_r163_c87 bl[87] br[87] wl[163] vdd gnd cell_6t
Xbit_r164_c87 bl[87] br[87] wl[164] vdd gnd cell_6t
Xbit_r165_c87 bl[87] br[87] wl[165] vdd gnd cell_6t
Xbit_r166_c87 bl[87] br[87] wl[166] vdd gnd cell_6t
Xbit_r167_c87 bl[87] br[87] wl[167] vdd gnd cell_6t
Xbit_r168_c87 bl[87] br[87] wl[168] vdd gnd cell_6t
Xbit_r169_c87 bl[87] br[87] wl[169] vdd gnd cell_6t
Xbit_r170_c87 bl[87] br[87] wl[170] vdd gnd cell_6t
Xbit_r171_c87 bl[87] br[87] wl[171] vdd gnd cell_6t
Xbit_r172_c87 bl[87] br[87] wl[172] vdd gnd cell_6t
Xbit_r173_c87 bl[87] br[87] wl[173] vdd gnd cell_6t
Xbit_r174_c87 bl[87] br[87] wl[174] vdd gnd cell_6t
Xbit_r175_c87 bl[87] br[87] wl[175] vdd gnd cell_6t
Xbit_r176_c87 bl[87] br[87] wl[176] vdd gnd cell_6t
Xbit_r177_c87 bl[87] br[87] wl[177] vdd gnd cell_6t
Xbit_r178_c87 bl[87] br[87] wl[178] vdd gnd cell_6t
Xbit_r179_c87 bl[87] br[87] wl[179] vdd gnd cell_6t
Xbit_r180_c87 bl[87] br[87] wl[180] vdd gnd cell_6t
Xbit_r181_c87 bl[87] br[87] wl[181] vdd gnd cell_6t
Xbit_r182_c87 bl[87] br[87] wl[182] vdd gnd cell_6t
Xbit_r183_c87 bl[87] br[87] wl[183] vdd gnd cell_6t
Xbit_r184_c87 bl[87] br[87] wl[184] vdd gnd cell_6t
Xbit_r185_c87 bl[87] br[87] wl[185] vdd gnd cell_6t
Xbit_r186_c87 bl[87] br[87] wl[186] vdd gnd cell_6t
Xbit_r187_c87 bl[87] br[87] wl[187] vdd gnd cell_6t
Xbit_r188_c87 bl[87] br[87] wl[188] vdd gnd cell_6t
Xbit_r189_c87 bl[87] br[87] wl[189] vdd gnd cell_6t
Xbit_r190_c87 bl[87] br[87] wl[190] vdd gnd cell_6t
Xbit_r191_c87 bl[87] br[87] wl[191] vdd gnd cell_6t
Xbit_r192_c87 bl[87] br[87] wl[192] vdd gnd cell_6t
Xbit_r193_c87 bl[87] br[87] wl[193] vdd gnd cell_6t
Xbit_r194_c87 bl[87] br[87] wl[194] vdd gnd cell_6t
Xbit_r195_c87 bl[87] br[87] wl[195] vdd gnd cell_6t
Xbit_r196_c87 bl[87] br[87] wl[196] vdd gnd cell_6t
Xbit_r197_c87 bl[87] br[87] wl[197] vdd gnd cell_6t
Xbit_r198_c87 bl[87] br[87] wl[198] vdd gnd cell_6t
Xbit_r199_c87 bl[87] br[87] wl[199] vdd gnd cell_6t
Xbit_r200_c87 bl[87] br[87] wl[200] vdd gnd cell_6t
Xbit_r201_c87 bl[87] br[87] wl[201] vdd gnd cell_6t
Xbit_r202_c87 bl[87] br[87] wl[202] vdd gnd cell_6t
Xbit_r203_c87 bl[87] br[87] wl[203] vdd gnd cell_6t
Xbit_r204_c87 bl[87] br[87] wl[204] vdd gnd cell_6t
Xbit_r205_c87 bl[87] br[87] wl[205] vdd gnd cell_6t
Xbit_r206_c87 bl[87] br[87] wl[206] vdd gnd cell_6t
Xbit_r207_c87 bl[87] br[87] wl[207] vdd gnd cell_6t
Xbit_r208_c87 bl[87] br[87] wl[208] vdd gnd cell_6t
Xbit_r209_c87 bl[87] br[87] wl[209] vdd gnd cell_6t
Xbit_r210_c87 bl[87] br[87] wl[210] vdd gnd cell_6t
Xbit_r211_c87 bl[87] br[87] wl[211] vdd gnd cell_6t
Xbit_r212_c87 bl[87] br[87] wl[212] vdd gnd cell_6t
Xbit_r213_c87 bl[87] br[87] wl[213] vdd gnd cell_6t
Xbit_r214_c87 bl[87] br[87] wl[214] vdd gnd cell_6t
Xbit_r215_c87 bl[87] br[87] wl[215] vdd gnd cell_6t
Xbit_r216_c87 bl[87] br[87] wl[216] vdd gnd cell_6t
Xbit_r217_c87 bl[87] br[87] wl[217] vdd gnd cell_6t
Xbit_r218_c87 bl[87] br[87] wl[218] vdd gnd cell_6t
Xbit_r219_c87 bl[87] br[87] wl[219] vdd gnd cell_6t
Xbit_r220_c87 bl[87] br[87] wl[220] vdd gnd cell_6t
Xbit_r221_c87 bl[87] br[87] wl[221] vdd gnd cell_6t
Xbit_r222_c87 bl[87] br[87] wl[222] vdd gnd cell_6t
Xbit_r223_c87 bl[87] br[87] wl[223] vdd gnd cell_6t
Xbit_r224_c87 bl[87] br[87] wl[224] vdd gnd cell_6t
Xbit_r225_c87 bl[87] br[87] wl[225] vdd gnd cell_6t
Xbit_r226_c87 bl[87] br[87] wl[226] vdd gnd cell_6t
Xbit_r227_c87 bl[87] br[87] wl[227] vdd gnd cell_6t
Xbit_r228_c87 bl[87] br[87] wl[228] vdd gnd cell_6t
Xbit_r229_c87 bl[87] br[87] wl[229] vdd gnd cell_6t
Xbit_r230_c87 bl[87] br[87] wl[230] vdd gnd cell_6t
Xbit_r231_c87 bl[87] br[87] wl[231] vdd gnd cell_6t
Xbit_r232_c87 bl[87] br[87] wl[232] vdd gnd cell_6t
Xbit_r233_c87 bl[87] br[87] wl[233] vdd gnd cell_6t
Xbit_r234_c87 bl[87] br[87] wl[234] vdd gnd cell_6t
Xbit_r235_c87 bl[87] br[87] wl[235] vdd gnd cell_6t
Xbit_r236_c87 bl[87] br[87] wl[236] vdd gnd cell_6t
Xbit_r237_c87 bl[87] br[87] wl[237] vdd gnd cell_6t
Xbit_r238_c87 bl[87] br[87] wl[238] vdd gnd cell_6t
Xbit_r239_c87 bl[87] br[87] wl[239] vdd gnd cell_6t
Xbit_r240_c87 bl[87] br[87] wl[240] vdd gnd cell_6t
Xbit_r241_c87 bl[87] br[87] wl[241] vdd gnd cell_6t
Xbit_r242_c87 bl[87] br[87] wl[242] vdd gnd cell_6t
Xbit_r243_c87 bl[87] br[87] wl[243] vdd gnd cell_6t
Xbit_r244_c87 bl[87] br[87] wl[244] vdd gnd cell_6t
Xbit_r245_c87 bl[87] br[87] wl[245] vdd gnd cell_6t
Xbit_r246_c87 bl[87] br[87] wl[246] vdd gnd cell_6t
Xbit_r247_c87 bl[87] br[87] wl[247] vdd gnd cell_6t
Xbit_r248_c87 bl[87] br[87] wl[248] vdd gnd cell_6t
Xbit_r249_c87 bl[87] br[87] wl[249] vdd gnd cell_6t
Xbit_r250_c87 bl[87] br[87] wl[250] vdd gnd cell_6t
Xbit_r251_c87 bl[87] br[87] wl[251] vdd gnd cell_6t
Xbit_r252_c87 bl[87] br[87] wl[252] vdd gnd cell_6t
Xbit_r253_c87 bl[87] br[87] wl[253] vdd gnd cell_6t
Xbit_r254_c87 bl[87] br[87] wl[254] vdd gnd cell_6t
Xbit_r255_c87 bl[87] br[87] wl[255] vdd gnd cell_6t
Xbit_r0_c88 bl[88] br[88] wl[0] vdd gnd cell_6t
Xbit_r1_c88 bl[88] br[88] wl[1] vdd gnd cell_6t
Xbit_r2_c88 bl[88] br[88] wl[2] vdd gnd cell_6t
Xbit_r3_c88 bl[88] br[88] wl[3] vdd gnd cell_6t
Xbit_r4_c88 bl[88] br[88] wl[4] vdd gnd cell_6t
Xbit_r5_c88 bl[88] br[88] wl[5] vdd gnd cell_6t
Xbit_r6_c88 bl[88] br[88] wl[6] vdd gnd cell_6t
Xbit_r7_c88 bl[88] br[88] wl[7] vdd gnd cell_6t
Xbit_r8_c88 bl[88] br[88] wl[8] vdd gnd cell_6t
Xbit_r9_c88 bl[88] br[88] wl[9] vdd gnd cell_6t
Xbit_r10_c88 bl[88] br[88] wl[10] vdd gnd cell_6t
Xbit_r11_c88 bl[88] br[88] wl[11] vdd gnd cell_6t
Xbit_r12_c88 bl[88] br[88] wl[12] vdd gnd cell_6t
Xbit_r13_c88 bl[88] br[88] wl[13] vdd gnd cell_6t
Xbit_r14_c88 bl[88] br[88] wl[14] vdd gnd cell_6t
Xbit_r15_c88 bl[88] br[88] wl[15] vdd gnd cell_6t
Xbit_r16_c88 bl[88] br[88] wl[16] vdd gnd cell_6t
Xbit_r17_c88 bl[88] br[88] wl[17] vdd gnd cell_6t
Xbit_r18_c88 bl[88] br[88] wl[18] vdd gnd cell_6t
Xbit_r19_c88 bl[88] br[88] wl[19] vdd gnd cell_6t
Xbit_r20_c88 bl[88] br[88] wl[20] vdd gnd cell_6t
Xbit_r21_c88 bl[88] br[88] wl[21] vdd gnd cell_6t
Xbit_r22_c88 bl[88] br[88] wl[22] vdd gnd cell_6t
Xbit_r23_c88 bl[88] br[88] wl[23] vdd gnd cell_6t
Xbit_r24_c88 bl[88] br[88] wl[24] vdd gnd cell_6t
Xbit_r25_c88 bl[88] br[88] wl[25] vdd gnd cell_6t
Xbit_r26_c88 bl[88] br[88] wl[26] vdd gnd cell_6t
Xbit_r27_c88 bl[88] br[88] wl[27] vdd gnd cell_6t
Xbit_r28_c88 bl[88] br[88] wl[28] vdd gnd cell_6t
Xbit_r29_c88 bl[88] br[88] wl[29] vdd gnd cell_6t
Xbit_r30_c88 bl[88] br[88] wl[30] vdd gnd cell_6t
Xbit_r31_c88 bl[88] br[88] wl[31] vdd gnd cell_6t
Xbit_r32_c88 bl[88] br[88] wl[32] vdd gnd cell_6t
Xbit_r33_c88 bl[88] br[88] wl[33] vdd gnd cell_6t
Xbit_r34_c88 bl[88] br[88] wl[34] vdd gnd cell_6t
Xbit_r35_c88 bl[88] br[88] wl[35] vdd gnd cell_6t
Xbit_r36_c88 bl[88] br[88] wl[36] vdd gnd cell_6t
Xbit_r37_c88 bl[88] br[88] wl[37] vdd gnd cell_6t
Xbit_r38_c88 bl[88] br[88] wl[38] vdd gnd cell_6t
Xbit_r39_c88 bl[88] br[88] wl[39] vdd gnd cell_6t
Xbit_r40_c88 bl[88] br[88] wl[40] vdd gnd cell_6t
Xbit_r41_c88 bl[88] br[88] wl[41] vdd gnd cell_6t
Xbit_r42_c88 bl[88] br[88] wl[42] vdd gnd cell_6t
Xbit_r43_c88 bl[88] br[88] wl[43] vdd gnd cell_6t
Xbit_r44_c88 bl[88] br[88] wl[44] vdd gnd cell_6t
Xbit_r45_c88 bl[88] br[88] wl[45] vdd gnd cell_6t
Xbit_r46_c88 bl[88] br[88] wl[46] vdd gnd cell_6t
Xbit_r47_c88 bl[88] br[88] wl[47] vdd gnd cell_6t
Xbit_r48_c88 bl[88] br[88] wl[48] vdd gnd cell_6t
Xbit_r49_c88 bl[88] br[88] wl[49] vdd gnd cell_6t
Xbit_r50_c88 bl[88] br[88] wl[50] vdd gnd cell_6t
Xbit_r51_c88 bl[88] br[88] wl[51] vdd gnd cell_6t
Xbit_r52_c88 bl[88] br[88] wl[52] vdd gnd cell_6t
Xbit_r53_c88 bl[88] br[88] wl[53] vdd gnd cell_6t
Xbit_r54_c88 bl[88] br[88] wl[54] vdd gnd cell_6t
Xbit_r55_c88 bl[88] br[88] wl[55] vdd gnd cell_6t
Xbit_r56_c88 bl[88] br[88] wl[56] vdd gnd cell_6t
Xbit_r57_c88 bl[88] br[88] wl[57] vdd gnd cell_6t
Xbit_r58_c88 bl[88] br[88] wl[58] vdd gnd cell_6t
Xbit_r59_c88 bl[88] br[88] wl[59] vdd gnd cell_6t
Xbit_r60_c88 bl[88] br[88] wl[60] vdd gnd cell_6t
Xbit_r61_c88 bl[88] br[88] wl[61] vdd gnd cell_6t
Xbit_r62_c88 bl[88] br[88] wl[62] vdd gnd cell_6t
Xbit_r63_c88 bl[88] br[88] wl[63] vdd gnd cell_6t
Xbit_r64_c88 bl[88] br[88] wl[64] vdd gnd cell_6t
Xbit_r65_c88 bl[88] br[88] wl[65] vdd gnd cell_6t
Xbit_r66_c88 bl[88] br[88] wl[66] vdd gnd cell_6t
Xbit_r67_c88 bl[88] br[88] wl[67] vdd gnd cell_6t
Xbit_r68_c88 bl[88] br[88] wl[68] vdd gnd cell_6t
Xbit_r69_c88 bl[88] br[88] wl[69] vdd gnd cell_6t
Xbit_r70_c88 bl[88] br[88] wl[70] vdd gnd cell_6t
Xbit_r71_c88 bl[88] br[88] wl[71] vdd gnd cell_6t
Xbit_r72_c88 bl[88] br[88] wl[72] vdd gnd cell_6t
Xbit_r73_c88 bl[88] br[88] wl[73] vdd gnd cell_6t
Xbit_r74_c88 bl[88] br[88] wl[74] vdd gnd cell_6t
Xbit_r75_c88 bl[88] br[88] wl[75] vdd gnd cell_6t
Xbit_r76_c88 bl[88] br[88] wl[76] vdd gnd cell_6t
Xbit_r77_c88 bl[88] br[88] wl[77] vdd gnd cell_6t
Xbit_r78_c88 bl[88] br[88] wl[78] vdd gnd cell_6t
Xbit_r79_c88 bl[88] br[88] wl[79] vdd gnd cell_6t
Xbit_r80_c88 bl[88] br[88] wl[80] vdd gnd cell_6t
Xbit_r81_c88 bl[88] br[88] wl[81] vdd gnd cell_6t
Xbit_r82_c88 bl[88] br[88] wl[82] vdd gnd cell_6t
Xbit_r83_c88 bl[88] br[88] wl[83] vdd gnd cell_6t
Xbit_r84_c88 bl[88] br[88] wl[84] vdd gnd cell_6t
Xbit_r85_c88 bl[88] br[88] wl[85] vdd gnd cell_6t
Xbit_r86_c88 bl[88] br[88] wl[86] vdd gnd cell_6t
Xbit_r87_c88 bl[88] br[88] wl[87] vdd gnd cell_6t
Xbit_r88_c88 bl[88] br[88] wl[88] vdd gnd cell_6t
Xbit_r89_c88 bl[88] br[88] wl[89] vdd gnd cell_6t
Xbit_r90_c88 bl[88] br[88] wl[90] vdd gnd cell_6t
Xbit_r91_c88 bl[88] br[88] wl[91] vdd gnd cell_6t
Xbit_r92_c88 bl[88] br[88] wl[92] vdd gnd cell_6t
Xbit_r93_c88 bl[88] br[88] wl[93] vdd gnd cell_6t
Xbit_r94_c88 bl[88] br[88] wl[94] vdd gnd cell_6t
Xbit_r95_c88 bl[88] br[88] wl[95] vdd gnd cell_6t
Xbit_r96_c88 bl[88] br[88] wl[96] vdd gnd cell_6t
Xbit_r97_c88 bl[88] br[88] wl[97] vdd gnd cell_6t
Xbit_r98_c88 bl[88] br[88] wl[98] vdd gnd cell_6t
Xbit_r99_c88 bl[88] br[88] wl[99] vdd gnd cell_6t
Xbit_r100_c88 bl[88] br[88] wl[100] vdd gnd cell_6t
Xbit_r101_c88 bl[88] br[88] wl[101] vdd gnd cell_6t
Xbit_r102_c88 bl[88] br[88] wl[102] vdd gnd cell_6t
Xbit_r103_c88 bl[88] br[88] wl[103] vdd gnd cell_6t
Xbit_r104_c88 bl[88] br[88] wl[104] vdd gnd cell_6t
Xbit_r105_c88 bl[88] br[88] wl[105] vdd gnd cell_6t
Xbit_r106_c88 bl[88] br[88] wl[106] vdd gnd cell_6t
Xbit_r107_c88 bl[88] br[88] wl[107] vdd gnd cell_6t
Xbit_r108_c88 bl[88] br[88] wl[108] vdd gnd cell_6t
Xbit_r109_c88 bl[88] br[88] wl[109] vdd gnd cell_6t
Xbit_r110_c88 bl[88] br[88] wl[110] vdd gnd cell_6t
Xbit_r111_c88 bl[88] br[88] wl[111] vdd gnd cell_6t
Xbit_r112_c88 bl[88] br[88] wl[112] vdd gnd cell_6t
Xbit_r113_c88 bl[88] br[88] wl[113] vdd gnd cell_6t
Xbit_r114_c88 bl[88] br[88] wl[114] vdd gnd cell_6t
Xbit_r115_c88 bl[88] br[88] wl[115] vdd gnd cell_6t
Xbit_r116_c88 bl[88] br[88] wl[116] vdd gnd cell_6t
Xbit_r117_c88 bl[88] br[88] wl[117] vdd gnd cell_6t
Xbit_r118_c88 bl[88] br[88] wl[118] vdd gnd cell_6t
Xbit_r119_c88 bl[88] br[88] wl[119] vdd gnd cell_6t
Xbit_r120_c88 bl[88] br[88] wl[120] vdd gnd cell_6t
Xbit_r121_c88 bl[88] br[88] wl[121] vdd gnd cell_6t
Xbit_r122_c88 bl[88] br[88] wl[122] vdd gnd cell_6t
Xbit_r123_c88 bl[88] br[88] wl[123] vdd gnd cell_6t
Xbit_r124_c88 bl[88] br[88] wl[124] vdd gnd cell_6t
Xbit_r125_c88 bl[88] br[88] wl[125] vdd gnd cell_6t
Xbit_r126_c88 bl[88] br[88] wl[126] vdd gnd cell_6t
Xbit_r127_c88 bl[88] br[88] wl[127] vdd gnd cell_6t
Xbit_r128_c88 bl[88] br[88] wl[128] vdd gnd cell_6t
Xbit_r129_c88 bl[88] br[88] wl[129] vdd gnd cell_6t
Xbit_r130_c88 bl[88] br[88] wl[130] vdd gnd cell_6t
Xbit_r131_c88 bl[88] br[88] wl[131] vdd gnd cell_6t
Xbit_r132_c88 bl[88] br[88] wl[132] vdd gnd cell_6t
Xbit_r133_c88 bl[88] br[88] wl[133] vdd gnd cell_6t
Xbit_r134_c88 bl[88] br[88] wl[134] vdd gnd cell_6t
Xbit_r135_c88 bl[88] br[88] wl[135] vdd gnd cell_6t
Xbit_r136_c88 bl[88] br[88] wl[136] vdd gnd cell_6t
Xbit_r137_c88 bl[88] br[88] wl[137] vdd gnd cell_6t
Xbit_r138_c88 bl[88] br[88] wl[138] vdd gnd cell_6t
Xbit_r139_c88 bl[88] br[88] wl[139] vdd gnd cell_6t
Xbit_r140_c88 bl[88] br[88] wl[140] vdd gnd cell_6t
Xbit_r141_c88 bl[88] br[88] wl[141] vdd gnd cell_6t
Xbit_r142_c88 bl[88] br[88] wl[142] vdd gnd cell_6t
Xbit_r143_c88 bl[88] br[88] wl[143] vdd gnd cell_6t
Xbit_r144_c88 bl[88] br[88] wl[144] vdd gnd cell_6t
Xbit_r145_c88 bl[88] br[88] wl[145] vdd gnd cell_6t
Xbit_r146_c88 bl[88] br[88] wl[146] vdd gnd cell_6t
Xbit_r147_c88 bl[88] br[88] wl[147] vdd gnd cell_6t
Xbit_r148_c88 bl[88] br[88] wl[148] vdd gnd cell_6t
Xbit_r149_c88 bl[88] br[88] wl[149] vdd gnd cell_6t
Xbit_r150_c88 bl[88] br[88] wl[150] vdd gnd cell_6t
Xbit_r151_c88 bl[88] br[88] wl[151] vdd gnd cell_6t
Xbit_r152_c88 bl[88] br[88] wl[152] vdd gnd cell_6t
Xbit_r153_c88 bl[88] br[88] wl[153] vdd gnd cell_6t
Xbit_r154_c88 bl[88] br[88] wl[154] vdd gnd cell_6t
Xbit_r155_c88 bl[88] br[88] wl[155] vdd gnd cell_6t
Xbit_r156_c88 bl[88] br[88] wl[156] vdd gnd cell_6t
Xbit_r157_c88 bl[88] br[88] wl[157] vdd gnd cell_6t
Xbit_r158_c88 bl[88] br[88] wl[158] vdd gnd cell_6t
Xbit_r159_c88 bl[88] br[88] wl[159] vdd gnd cell_6t
Xbit_r160_c88 bl[88] br[88] wl[160] vdd gnd cell_6t
Xbit_r161_c88 bl[88] br[88] wl[161] vdd gnd cell_6t
Xbit_r162_c88 bl[88] br[88] wl[162] vdd gnd cell_6t
Xbit_r163_c88 bl[88] br[88] wl[163] vdd gnd cell_6t
Xbit_r164_c88 bl[88] br[88] wl[164] vdd gnd cell_6t
Xbit_r165_c88 bl[88] br[88] wl[165] vdd gnd cell_6t
Xbit_r166_c88 bl[88] br[88] wl[166] vdd gnd cell_6t
Xbit_r167_c88 bl[88] br[88] wl[167] vdd gnd cell_6t
Xbit_r168_c88 bl[88] br[88] wl[168] vdd gnd cell_6t
Xbit_r169_c88 bl[88] br[88] wl[169] vdd gnd cell_6t
Xbit_r170_c88 bl[88] br[88] wl[170] vdd gnd cell_6t
Xbit_r171_c88 bl[88] br[88] wl[171] vdd gnd cell_6t
Xbit_r172_c88 bl[88] br[88] wl[172] vdd gnd cell_6t
Xbit_r173_c88 bl[88] br[88] wl[173] vdd gnd cell_6t
Xbit_r174_c88 bl[88] br[88] wl[174] vdd gnd cell_6t
Xbit_r175_c88 bl[88] br[88] wl[175] vdd gnd cell_6t
Xbit_r176_c88 bl[88] br[88] wl[176] vdd gnd cell_6t
Xbit_r177_c88 bl[88] br[88] wl[177] vdd gnd cell_6t
Xbit_r178_c88 bl[88] br[88] wl[178] vdd gnd cell_6t
Xbit_r179_c88 bl[88] br[88] wl[179] vdd gnd cell_6t
Xbit_r180_c88 bl[88] br[88] wl[180] vdd gnd cell_6t
Xbit_r181_c88 bl[88] br[88] wl[181] vdd gnd cell_6t
Xbit_r182_c88 bl[88] br[88] wl[182] vdd gnd cell_6t
Xbit_r183_c88 bl[88] br[88] wl[183] vdd gnd cell_6t
Xbit_r184_c88 bl[88] br[88] wl[184] vdd gnd cell_6t
Xbit_r185_c88 bl[88] br[88] wl[185] vdd gnd cell_6t
Xbit_r186_c88 bl[88] br[88] wl[186] vdd gnd cell_6t
Xbit_r187_c88 bl[88] br[88] wl[187] vdd gnd cell_6t
Xbit_r188_c88 bl[88] br[88] wl[188] vdd gnd cell_6t
Xbit_r189_c88 bl[88] br[88] wl[189] vdd gnd cell_6t
Xbit_r190_c88 bl[88] br[88] wl[190] vdd gnd cell_6t
Xbit_r191_c88 bl[88] br[88] wl[191] vdd gnd cell_6t
Xbit_r192_c88 bl[88] br[88] wl[192] vdd gnd cell_6t
Xbit_r193_c88 bl[88] br[88] wl[193] vdd gnd cell_6t
Xbit_r194_c88 bl[88] br[88] wl[194] vdd gnd cell_6t
Xbit_r195_c88 bl[88] br[88] wl[195] vdd gnd cell_6t
Xbit_r196_c88 bl[88] br[88] wl[196] vdd gnd cell_6t
Xbit_r197_c88 bl[88] br[88] wl[197] vdd gnd cell_6t
Xbit_r198_c88 bl[88] br[88] wl[198] vdd gnd cell_6t
Xbit_r199_c88 bl[88] br[88] wl[199] vdd gnd cell_6t
Xbit_r200_c88 bl[88] br[88] wl[200] vdd gnd cell_6t
Xbit_r201_c88 bl[88] br[88] wl[201] vdd gnd cell_6t
Xbit_r202_c88 bl[88] br[88] wl[202] vdd gnd cell_6t
Xbit_r203_c88 bl[88] br[88] wl[203] vdd gnd cell_6t
Xbit_r204_c88 bl[88] br[88] wl[204] vdd gnd cell_6t
Xbit_r205_c88 bl[88] br[88] wl[205] vdd gnd cell_6t
Xbit_r206_c88 bl[88] br[88] wl[206] vdd gnd cell_6t
Xbit_r207_c88 bl[88] br[88] wl[207] vdd gnd cell_6t
Xbit_r208_c88 bl[88] br[88] wl[208] vdd gnd cell_6t
Xbit_r209_c88 bl[88] br[88] wl[209] vdd gnd cell_6t
Xbit_r210_c88 bl[88] br[88] wl[210] vdd gnd cell_6t
Xbit_r211_c88 bl[88] br[88] wl[211] vdd gnd cell_6t
Xbit_r212_c88 bl[88] br[88] wl[212] vdd gnd cell_6t
Xbit_r213_c88 bl[88] br[88] wl[213] vdd gnd cell_6t
Xbit_r214_c88 bl[88] br[88] wl[214] vdd gnd cell_6t
Xbit_r215_c88 bl[88] br[88] wl[215] vdd gnd cell_6t
Xbit_r216_c88 bl[88] br[88] wl[216] vdd gnd cell_6t
Xbit_r217_c88 bl[88] br[88] wl[217] vdd gnd cell_6t
Xbit_r218_c88 bl[88] br[88] wl[218] vdd gnd cell_6t
Xbit_r219_c88 bl[88] br[88] wl[219] vdd gnd cell_6t
Xbit_r220_c88 bl[88] br[88] wl[220] vdd gnd cell_6t
Xbit_r221_c88 bl[88] br[88] wl[221] vdd gnd cell_6t
Xbit_r222_c88 bl[88] br[88] wl[222] vdd gnd cell_6t
Xbit_r223_c88 bl[88] br[88] wl[223] vdd gnd cell_6t
Xbit_r224_c88 bl[88] br[88] wl[224] vdd gnd cell_6t
Xbit_r225_c88 bl[88] br[88] wl[225] vdd gnd cell_6t
Xbit_r226_c88 bl[88] br[88] wl[226] vdd gnd cell_6t
Xbit_r227_c88 bl[88] br[88] wl[227] vdd gnd cell_6t
Xbit_r228_c88 bl[88] br[88] wl[228] vdd gnd cell_6t
Xbit_r229_c88 bl[88] br[88] wl[229] vdd gnd cell_6t
Xbit_r230_c88 bl[88] br[88] wl[230] vdd gnd cell_6t
Xbit_r231_c88 bl[88] br[88] wl[231] vdd gnd cell_6t
Xbit_r232_c88 bl[88] br[88] wl[232] vdd gnd cell_6t
Xbit_r233_c88 bl[88] br[88] wl[233] vdd gnd cell_6t
Xbit_r234_c88 bl[88] br[88] wl[234] vdd gnd cell_6t
Xbit_r235_c88 bl[88] br[88] wl[235] vdd gnd cell_6t
Xbit_r236_c88 bl[88] br[88] wl[236] vdd gnd cell_6t
Xbit_r237_c88 bl[88] br[88] wl[237] vdd gnd cell_6t
Xbit_r238_c88 bl[88] br[88] wl[238] vdd gnd cell_6t
Xbit_r239_c88 bl[88] br[88] wl[239] vdd gnd cell_6t
Xbit_r240_c88 bl[88] br[88] wl[240] vdd gnd cell_6t
Xbit_r241_c88 bl[88] br[88] wl[241] vdd gnd cell_6t
Xbit_r242_c88 bl[88] br[88] wl[242] vdd gnd cell_6t
Xbit_r243_c88 bl[88] br[88] wl[243] vdd gnd cell_6t
Xbit_r244_c88 bl[88] br[88] wl[244] vdd gnd cell_6t
Xbit_r245_c88 bl[88] br[88] wl[245] vdd gnd cell_6t
Xbit_r246_c88 bl[88] br[88] wl[246] vdd gnd cell_6t
Xbit_r247_c88 bl[88] br[88] wl[247] vdd gnd cell_6t
Xbit_r248_c88 bl[88] br[88] wl[248] vdd gnd cell_6t
Xbit_r249_c88 bl[88] br[88] wl[249] vdd gnd cell_6t
Xbit_r250_c88 bl[88] br[88] wl[250] vdd gnd cell_6t
Xbit_r251_c88 bl[88] br[88] wl[251] vdd gnd cell_6t
Xbit_r252_c88 bl[88] br[88] wl[252] vdd gnd cell_6t
Xbit_r253_c88 bl[88] br[88] wl[253] vdd gnd cell_6t
Xbit_r254_c88 bl[88] br[88] wl[254] vdd gnd cell_6t
Xbit_r255_c88 bl[88] br[88] wl[255] vdd gnd cell_6t
Xbit_r0_c89 bl[89] br[89] wl[0] vdd gnd cell_6t
Xbit_r1_c89 bl[89] br[89] wl[1] vdd gnd cell_6t
Xbit_r2_c89 bl[89] br[89] wl[2] vdd gnd cell_6t
Xbit_r3_c89 bl[89] br[89] wl[3] vdd gnd cell_6t
Xbit_r4_c89 bl[89] br[89] wl[4] vdd gnd cell_6t
Xbit_r5_c89 bl[89] br[89] wl[5] vdd gnd cell_6t
Xbit_r6_c89 bl[89] br[89] wl[6] vdd gnd cell_6t
Xbit_r7_c89 bl[89] br[89] wl[7] vdd gnd cell_6t
Xbit_r8_c89 bl[89] br[89] wl[8] vdd gnd cell_6t
Xbit_r9_c89 bl[89] br[89] wl[9] vdd gnd cell_6t
Xbit_r10_c89 bl[89] br[89] wl[10] vdd gnd cell_6t
Xbit_r11_c89 bl[89] br[89] wl[11] vdd gnd cell_6t
Xbit_r12_c89 bl[89] br[89] wl[12] vdd gnd cell_6t
Xbit_r13_c89 bl[89] br[89] wl[13] vdd gnd cell_6t
Xbit_r14_c89 bl[89] br[89] wl[14] vdd gnd cell_6t
Xbit_r15_c89 bl[89] br[89] wl[15] vdd gnd cell_6t
Xbit_r16_c89 bl[89] br[89] wl[16] vdd gnd cell_6t
Xbit_r17_c89 bl[89] br[89] wl[17] vdd gnd cell_6t
Xbit_r18_c89 bl[89] br[89] wl[18] vdd gnd cell_6t
Xbit_r19_c89 bl[89] br[89] wl[19] vdd gnd cell_6t
Xbit_r20_c89 bl[89] br[89] wl[20] vdd gnd cell_6t
Xbit_r21_c89 bl[89] br[89] wl[21] vdd gnd cell_6t
Xbit_r22_c89 bl[89] br[89] wl[22] vdd gnd cell_6t
Xbit_r23_c89 bl[89] br[89] wl[23] vdd gnd cell_6t
Xbit_r24_c89 bl[89] br[89] wl[24] vdd gnd cell_6t
Xbit_r25_c89 bl[89] br[89] wl[25] vdd gnd cell_6t
Xbit_r26_c89 bl[89] br[89] wl[26] vdd gnd cell_6t
Xbit_r27_c89 bl[89] br[89] wl[27] vdd gnd cell_6t
Xbit_r28_c89 bl[89] br[89] wl[28] vdd gnd cell_6t
Xbit_r29_c89 bl[89] br[89] wl[29] vdd gnd cell_6t
Xbit_r30_c89 bl[89] br[89] wl[30] vdd gnd cell_6t
Xbit_r31_c89 bl[89] br[89] wl[31] vdd gnd cell_6t
Xbit_r32_c89 bl[89] br[89] wl[32] vdd gnd cell_6t
Xbit_r33_c89 bl[89] br[89] wl[33] vdd gnd cell_6t
Xbit_r34_c89 bl[89] br[89] wl[34] vdd gnd cell_6t
Xbit_r35_c89 bl[89] br[89] wl[35] vdd gnd cell_6t
Xbit_r36_c89 bl[89] br[89] wl[36] vdd gnd cell_6t
Xbit_r37_c89 bl[89] br[89] wl[37] vdd gnd cell_6t
Xbit_r38_c89 bl[89] br[89] wl[38] vdd gnd cell_6t
Xbit_r39_c89 bl[89] br[89] wl[39] vdd gnd cell_6t
Xbit_r40_c89 bl[89] br[89] wl[40] vdd gnd cell_6t
Xbit_r41_c89 bl[89] br[89] wl[41] vdd gnd cell_6t
Xbit_r42_c89 bl[89] br[89] wl[42] vdd gnd cell_6t
Xbit_r43_c89 bl[89] br[89] wl[43] vdd gnd cell_6t
Xbit_r44_c89 bl[89] br[89] wl[44] vdd gnd cell_6t
Xbit_r45_c89 bl[89] br[89] wl[45] vdd gnd cell_6t
Xbit_r46_c89 bl[89] br[89] wl[46] vdd gnd cell_6t
Xbit_r47_c89 bl[89] br[89] wl[47] vdd gnd cell_6t
Xbit_r48_c89 bl[89] br[89] wl[48] vdd gnd cell_6t
Xbit_r49_c89 bl[89] br[89] wl[49] vdd gnd cell_6t
Xbit_r50_c89 bl[89] br[89] wl[50] vdd gnd cell_6t
Xbit_r51_c89 bl[89] br[89] wl[51] vdd gnd cell_6t
Xbit_r52_c89 bl[89] br[89] wl[52] vdd gnd cell_6t
Xbit_r53_c89 bl[89] br[89] wl[53] vdd gnd cell_6t
Xbit_r54_c89 bl[89] br[89] wl[54] vdd gnd cell_6t
Xbit_r55_c89 bl[89] br[89] wl[55] vdd gnd cell_6t
Xbit_r56_c89 bl[89] br[89] wl[56] vdd gnd cell_6t
Xbit_r57_c89 bl[89] br[89] wl[57] vdd gnd cell_6t
Xbit_r58_c89 bl[89] br[89] wl[58] vdd gnd cell_6t
Xbit_r59_c89 bl[89] br[89] wl[59] vdd gnd cell_6t
Xbit_r60_c89 bl[89] br[89] wl[60] vdd gnd cell_6t
Xbit_r61_c89 bl[89] br[89] wl[61] vdd gnd cell_6t
Xbit_r62_c89 bl[89] br[89] wl[62] vdd gnd cell_6t
Xbit_r63_c89 bl[89] br[89] wl[63] vdd gnd cell_6t
Xbit_r64_c89 bl[89] br[89] wl[64] vdd gnd cell_6t
Xbit_r65_c89 bl[89] br[89] wl[65] vdd gnd cell_6t
Xbit_r66_c89 bl[89] br[89] wl[66] vdd gnd cell_6t
Xbit_r67_c89 bl[89] br[89] wl[67] vdd gnd cell_6t
Xbit_r68_c89 bl[89] br[89] wl[68] vdd gnd cell_6t
Xbit_r69_c89 bl[89] br[89] wl[69] vdd gnd cell_6t
Xbit_r70_c89 bl[89] br[89] wl[70] vdd gnd cell_6t
Xbit_r71_c89 bl[89] br[89] wl[71] vdd gnd cell_6t
Xbit_r72_c89 bl[89] br[89] wl[72] vdd gnd cell_6t
Xbit_r73_c89 bl[89] br[89] wl[73] vdd gnd cell_6t
Xbit_r74_c89 bl[89] br[89] wl[74] vdd gnd cell_6t
Xbit_r75_c89 bl[89] br[89] wl[75] vdd gnd cell_6t
Xbit_r76_c89 bl[89] br[89] wl[76] vdd gnd cell_6t
Xbit_r77_c89 bl[89] br[89] wl[77] vdd gnd cell_6t
Xbit_r78_c89 bl[89] br[89] wl[78] vdd gnd cell_6t
Xbit_r79_c89 bl[89] br[89] wl[79] vdd gnd cell_6t
Xbit_r80_c89 bl[89] br[89] wl[80] vdd gnd cell_6t
Xbit_r81_c89 bl[89] br[89] wl[81] vdd gnd cell_6t
Xbit_r82_c89 bl[89] br[89] wl[82] vdd gnd cell_6t
Xbit_r83_c89 bl[89] br[89] wl[83] vdd gnd cell_6t
Xbit_r84_c89 bl[89] br[89] wl[84] vdd gnd cell_6t
Xbit_r85_c89 bl[89] br[89] wl[85] vdd gnd cell_6t
Xbit_r86_c89 bl[89] br[89] wl[86] vdd gnd cell_6t
Xbit_r87_c89 bl[89] br[89] wl[87] vdd gnd cell_6t
Xbit_r88_c89 bl[89] br[89] wl[88] vdd gnd cell_6t
Xbit_r89_c89 bl[89] br[89] wl[89] vdd gnd cell_6t
Xbit_r90_c89 bl[89] br[89] wl[90] vdd gnd cell_6t
Xbit_r91_c89 bl[89] br[89] wl[91] vdd gnd cell_6t
Xbit_r92_c89 bl[89] br[89] wl[92] vdd gnd cell_6t
Xbit_r93_c89 bl[89] br[89] wl[93] vdd gnd cell_6t
Xbit_r94_c89 bl[89] br[89] wl[94] vdd gnd cell_6t
Xbit_r95_c89 bl[89] br[89] wl[95] vdd gnd cell_6t
Xbit_r96_c89 bl[89] br[89] wl[96] vdd gnd cell_6t
Xbit_r97_c89 bl[89] br[89] wl[97] vdd gnd cell_6t
Xbit_r98_c89 bl[89] br[89] wl[98] vdd gnd cell_6t
Xbit_r99_c89 bl[89] br[89] wl[99] vdd gnd cell_6t
Xbit_r100_c89 bl[89] br[89] wl[100] vdd gnd cell_6t
Xbit_r101_c89 bl[89] br[89] wl[101] vdd gnd cell_6t
Xbit_r102_c89 bl[89] br[89] wl[102] vdd gnd cell_6t
Xbit_r103_c89 bl[89] br[89] wl[103] vdd gnd cell_6t
Xbit_r104_c89 bl[89] br[89] wl[104] vdd gnd cell_6t
Xbit_r105_c89 bl[89] br[89] wl[105] vdd gnd cell_6t
Xbit_r106_c89 bl[89] br[89] wl[106] vdd gnd cell_6t
Xbit_r107_c89 bl[89] br[89] wl[107] vdd gnd cell_6t
Xbit_r108_c89 bl[89] br[89] wl[108] vdd gnd cell_6t
Xbit_r109_c89 bl[89] br[89] wl[109] vdd gnd cell_6t
Xbit_r110_c89 bl[89] br[89] wl[110] vdd gnd cell_6t
Xbit_r111_c89 bl[89] br[89] wl[111] vdd gnd cell_6t
Xbit_r112_c89 bl[89] br[89] wl[112] vdd gnd cell_6t
Xbit_r113_c89 bl[89] br[89] wl[113] vdd gnd cell_6t
Xbit_r114_c89 bl[89] br[89] wl[114] vdd gnd cell_6t
Xbit_r115_c89 bl[89] br[89] wl[115] vdd gnd cell_6t
Xbit_r116_c89 bl[89] br[89] wl[116] vdd gnd cell_6t
Xbit_r117_c89 bl[89] br[89] wl[117] vdd gnd cell_6t
Xbit_r118_c89 bl[89] br[89] wl[118] vdd gnd cell_6t
Xbit_r119_c89 bl[89] br[89] wl[119] vdd gnd cell_6t
Xbit_r120_c89 bl[89] br[89] wl[120] vdd gnd cell_6t
Xbit_r121_c89 bl[89] br[89] wl[121] vdd gnd cell_6t
Xbit_r122_c89 bl[89] br[89] wl[122] vdd gnd cell_6t
Xbit_r123_c89 bl[89] br[89] wl[123] vdd gnd cell_6t
Xbit_r124_c89 bl[89] br[89] wl[124] vdd gnd cell_6t
Xbit_r125_c89 bl[89] br[89] wl[125] vdd gnd cell_6t
Xbit_r126_c89 bl[89] br[89] wl[126] vdd gnd cell_6t
Xbit_r127_c89 bl[89] br[89] wl[127] vdd gnd cell_6t
Xbit_r128_c89 bl[89] br[89] wl[128] vdd gnd cell_6t
Xbit_r129_c89 bl[89] br[89] wl[129] vdd gnd cell_6t
Xbit_r130_c89 bl[89] br[89] wl[130] vdd gnd cell_6t
Xbit_r131_c89 bl[89] br[89] wl[131] vdd gnd cell_6t
Xbit_r132_c89 bl[89] br[89] wl[132] vdd gnd cell_6t
Xbit_r133_c89 bl[89] br[89] wl[133] vdd gnd cell_6t
Xbit_r134_c89 bl[89] br[89] wl[134] vdd gnd cell_6t
Xbit_r135_c89 bl[89] br[89] wl[135] vdd gnd cell_6t
Xbit_r136_c89 bl[89] br[89] wl[136] vdd gnd cell_6t
Xbit_r137_c89 bl[89] br[89] wl[137] vdd gnd cell_6t
Xbit_r138_c89 bl[89] br[89] wl[138] vdd gnd cell_6t
Xbit_r139_c89 bl[89] br[89] wl[139] vdd gnd cell_6t
Xbit_r140_c89 bl[89] br[89] wl[140] vdd gnd cell_6t
Xbit_r141_c89 bl[89] br[89] wl[141] vdd gnd cell_6t
Xbit_r142_c89 bl[89] br[89] wl[142] vdd gnd cell_6t
Xbit_r143_c89 bl[89] br[89] wl[143] vdd gnd cell_6t
Xbit_r144_c89 bl[89] br[89] wl[144] vdd gnd cell_6t
Xbit_r145_c89 bl[89] br[89] wl[145] vdd gnd cell_6t
Xbit_r146_c89 bl[89] br[89] wl[146] vdd gnd cell_6t
Xbit_r147_c89 bl[89] br[89] wl[147] vdd gnd cell_6t
Xbit_r148_c89 bl[89] br[89] wl[148] vdd gnd cell_6t
Xbit_r149_c89 bl[89] br[89] wl[149] vdd gnd cell_6t
Xbit_r150_c89 bl[89] br[89] wl[150] vdd gnd cell_6t
Xbit_r151_c89 bl[89] br[89] wl[151] vdd gnd cell_6t
Xbit_r152_c89 bl[89] br[89] wl[152] vdd gnd cell_6t
Xbit_r153_c89 bl[89] br[89] wl[153] vdd gnd cell_6t
Xbit_r154_c89 bl[89] br[89] wl[154] vdd gnd cell_6t
Xbit_r155_c89 bl[89] br[89] wl[155] vdd gnd cell_6t
Xbit_r156_c89 bl[89] br[89] wl[156] vdd gnd cell_6t
Xbit_r157_c89 bl[89] br[89] wl[157] vdd gnd cell_6t
Xbit_r158_c89 bl[89] br[89] wl[158] vdd gnd cell_6t
Xbit_r159_c89 bl[89] br[89] wl[159] vdd gnd cell_6t
Xbit_r160_c89 bl[89] br[89] wl[160] vdd gnd cell_6t
Xbit_r161_c89 bl[89] br[89] wl[161] vdd gnd cell_6t
Xbit_r162_c89 bl[89] br[89] wl[162] vdd gnd cell_6t
Xbit_r163_c89 bl[89] br[89] wl[163] vdd gnd cell_6t
Xbit_r164_c89 bl[89] br[89] wl[164] vdd gnd cell_6t
Xbit_r165_c89 bl[89] br[89] wl[165] vdd gnd cell_6t
Xbit_r166_c89 bl[89] br[89] wl[166] vdd gnd cell_6t
Xbit_r167_c89 bl[89] br[89] wl[167] vdd gnd cell_6t
Xbit_r168_c89 bl[89] br[89] wl[168] vdd gnd cell_6t
Xbit_r169_c89 bl[89] br[89] wl[169] vdd gnd cell_6t
Xbit_r170_c89 bl[89] br[89] wl[170] vdd gnd cell_6t
Xbit_r171_c89 bl[89] br[89] wl[171] vdd gnd cell_6t
Xbit_r172_c89 bl[89] br[89] wl[172] vdd gnd cell_6t
Xbit_r173_c89 bl[89] br[89] wl[173] vdd gnd cell_6t
Xbit_r174_c89 bl[89] br[89] wl[174] vdd gnd cell_6t
Xbit_r175_c89 bl[89] br[89] wl[175] vdd gnd cell_6t
Xbit_r176_c89 bl[89] br[89] wl[176] vdd gnd cell_6t
Xbit_r177_c89 bl[89] br[89] wl[177] vdd gnd cell_6t
Xbit_r178_c89 bl[89] br[89] wl[178] vdd gnd cell_6t
Xbit_r179_c89 bl[89] br[89] wl[179] vdd gnd cell_6t
Xbit_r180_c89 bl[89] br[89] wl[180] vdd gnd cell_6t
Xbit_r181_c89 bl[89] br[89] wl[181] vdd gnd cell_6t
Xbit_r182_c89 bl[89] br[89] wl[182] vdd gnd cell_6t
Xbit_r183_c89 bl[89] br[89] wl[183] vdd gnd cell_6t
Xbit_r184_c89 bl[89] br[89] wl[184] vdd gnd cell_6t
Xbit_r185_c89 bl[89] br[89] wl[185] vdd gnd cell_6t
Xbit_r186_c89 bl[89] br[89] wl[186] vdd gnd cell_6t
Xbit_r187_c89 bl[89] br[89] wl[187] vdd gnd cell_6t
Xbit_r188_c89 bl[89] br[89] wl[188] vdd gnd cell_6t
Xbit_r189_c89 bl[89] br[89] wl[189] vdd gnd cell_6t
Xbit_r190_c89 bl[89] br[89] wl[190] vdd gnd cell_6t
Xbit_r191_c89 bl[89] br[89] wl[191] vdd gnd cell_6t
Xbit_r192_c89 bl[89] br[89] wl[192] vdd gnd cell_6t
Xbit_r193_c89 bl[89] br[89] wl[193] vdd gnd cell_6t
Xbit_r194_c89 bl[89] br[89] wl[194] vdd gnd cell_6t
Xbit_r195_c89 bl[89] br[89] wl[195] vdd gnd cell_6t
Xbit_r196_c89 bl[89] br[89] wl[196] vdd gnd cell_6t
Xbit_r197_c89 bl[89] br[89] wl[197] vdd gnd cell_6t
Xbit_r198_c89 bl[89] br[89] wl[198] vdd gnd cell_6t
Xbit_r199_c89 bl[89] br[89] wl[199] vdd gnd cell_6t
Xbit_r200_c89 bl[89] br[89] wl[200] vdd gnd cell_6t
Xbit_r201_c89 bl[89] br[89] wl[201] vdd gnd cell_6t
Xbit_r202_c89 bl[89] br[89] wl[202] vdd gnd cell_6t
Xbit_r203_c89 bl[89] br[89] wl[203] vdd gnd cell_6t
Xbit_r204_c89 bl[89] br[89] wl[204] vdd gnd cell_6t
Xbit_r205_c89 bl[89] br[89] wl[205] vdd gnd cell_6t
Xbit_r206_c89 bl[89] br[89] wl[206] vdd gnd cell_6t
Xbit_r207_c89 bl[89] br[89] wl[207] vdd gnd cell_6t
Xbit_r208_c89 bl[89] br[89] wl[208] vdd gnd cell_6t
Xbit_r209_c89 bl[89] br[89] wl[209] vdd gnd cell_6t
Xbit_r210_c89 bl[89] br[89] wl[210] vdd gnd cell_6t
Xbit_r211_c89 bl[89] br[89] wl[211] vdd gnd cell_6t
Xbit_r212_c89 bl[89] br[89] wl[212] vdd gnd cell_6t
Xbit_r213_c89 bl[89] br[89] wl[213] vdd gnd cell_6t
Xbit_r214_c89 bl[89] br[89] wl[214] vdd gnd cell_6t
Xbit_r215_c89 bl[89] br[89] wl[215] vdd gnd cell_6t
Xbit_r216_c89 bl[89] br[89] wl[216] vdd gnd cell_6t
Xbit_r217_c89 bl[89] br[89] wl[217] vdd gnd cell_6t
Xbit_r218_c89 bl[89] br[89] wl[218] vdd gnd cell_6t
Xbit_r219_c89 bl[89] br[89] wl[219] vdd gnd cell_6t
Xbit_r220_c89 bl[89] br[89] wl[220] vdd gnd cell_6t
Xbit_r221_c89 bl[89] br[89] wl[221] vdd gnd cell_6t
Xbit_r222_c89 bl[89] br[89] wl[222] vdd gnd cell_6t
Xbit_r223_c89 bl[89] br[89] wl[223] vdd gnd cell_6t
Xbit_r224_c89 bl[89] br[89] wl[224] vdd gnd cell_6t
Xbit_r225_c89 bl[89] br[89] wl[225] vdd gnd cell_6t
Xbit_r226_c89 bl[89] br[89] wl[226] vdd gnd cell_6t
Xbit_r227_c89 bl[89] br[89] wl[227] vdd gnd cell_6t
Xbit_r228_c89 bl[89] br[89] wl[228] vdd gnd cell_6t
Xbit_r229_c89 bl[89] br[89] wl[229] vdd gnd cell_6t
Xbit_r230_c89 bl[89] br[89] wl[230] vdd gnd cell_6t
Xbit_r231_c89 bl[89] br[89] wl[231] vdd gnd cell_6t
Xbit_r232_c89 bl[89] br[89] wl[232] vdd gnd cell_6t
Xbit_r233_c89 bl[89] br[89] wl[233] vdd gnd cell_6t
Xbit_r234_c89 bl[89] br[89] wl[234] vdd gnd cell_6t
Xbit_r235_c89 bl[89] br[89] wl[235] vdd gnd cell_6t
Xbit_r236_c89 bl[89] br[89] wl[236] vdd gnd cell_6t
Xbit_r237_c89 bl[89] br[89] wl[237] vdd gnd cell_6t
Xbit_r238_c89 bl[89] br[89] wl[238] vdd gnd cell_6t
Xbit_r239_c89 bl[89] br[89] wl[239] vdd gnd cell_6t
Xbit_r240_c89 bl[89] br[89] wl[240] vdd gnd cell_6t
Xbit_r241_c89 bl[89] br[89] wl[241] vdd gnd cell_6t
Xbit_r242_c89 bl[89] br[89] wl[242] vdd gnd cell_6t
Xbit_r243_c89 bl[89] br[89] wl[243] vdd gnd cell_6t
Xbit_r244_c89 bl[89] br[89] wl[244] vdd gnd cell_6t
Xbit_r245_c89 bl[89] br[89] wl[245] vdd gnd cell_6t
Xbit_r246_c89 bl[89] br[89] wl[246] vdd gnd cell_6t
Xbit_r247_c89 bl[89] br[89] wl[247] vdd gnd cell_6t
Xbit_r248_c89 bl[89] br[89] wl[248] vdd gnd cell_6t
Xbit_r249_c89 bl[89] br[89] wl[249] vdd gnd cell_6t
Xbit_r250_c89 bl[89] br[89] wl[250] vdd gnd cell_6t
Xbit_r251_c89 bl[89] br[89] wl[251] vdd gnd cell_6t
Xbit_r252_c89 bl[89] br[89] wl[252] vdd gnd cell_6t
Xbit_r253_c89 bl[89] br[89] wl[253] vdd gnd cell_6t
Xbit_r254_c89 bl[89] br[89] wl[254] vdd gnd cell_6t
Xbit_r255_c89 bl[89] br[89] wl[255] vdd gnd cell_6t
Xbit_r0_c90 bl[90] br[90] wl[0] vdd gnd cell_6t
Xbit_r1_c90 bl[90] br[90] wl[1] vdd gnd cell_6t
Xbit_r2_c90 bl[90] br[90] wl[2] vdd gnd cell_6t
Xbit_r3_c90 bl[90] br[90] wl[3] vdd gnd cell_6t
Xbit_r4_c90 bl[90] br[90] wl[4] vdd gnd cell_6t
Xbit_r5_c90 bl[90] br[90] wl[5] vdd gnd cell_6t
Xbit_r6_c90 bl[90] br[90] wl[6] vdd gnd cell_6t
Xbit_r7_c90 bl[90] br[90] wl[7] vdd gnd cell_6t
Xbit_r8_c90 bl[90] br[90] wl[8] vdd gnd cell_6t
Xbit_r9_c90 bl[90] br[90] wl[9] vdd gnd cell_6t
Xbit_r10_c90 bl[90] br[90] wl[10] vdd gnd cell_6t
Xbit_r11_c90 bl[90] br[90] wl[11] vdd gnd cell_6t
Xbit_r12_c90 bl[90] br[90] wl[12] vdd gnd cell_6t
Xbit_r13_c90 bl[90] br[90] wl[13] vdd gnd cell_6t
Xbit_r14_c90 bl[90] br[90] wl[14] vdd gnd cell_6t
Xbit_r15_c90 bl[90] br[90] wl[15] vdd gnd cell_6t
Xbit_r16_c90 bl[90] br[90] wl[16] vdd gnd cell_6t
Xbit_r17_c90 bl[90] br[90] wl[17] vdd gnd cell_6t
Xbit_r18_c90 bl[90] br[90] wl[18] vdd gnd cell_6t
Xbit_r19_c90 bl[90] br[90] wl[19] vdd gnd cell_6t
Xbit_r20_c90 bl[90] br[90] wl[20] vdd gnd cell_6t
Xbit_r21_c90 bl[90] br[90] wl[21] vdd gnd cell_6t
Xbit_r22_c90 bl[90] br[90] wl[22] vdd gnd cell_6t
Xbit_r23_c90 bl[90] br[90] wl[23] vdd gnd cell_6t
Xbit_r24_c90 bl[90] br[90] wl[24] vdd gnd cell_6t
Xbit_r25_c90 bl[90] br[90] wl[25] vdd gnd cell_6t
Xbit_r26_c90 bl[90] br[90] wl[26] vdd gnd cell_6t
Xbit_r27_c90 bl[90] br[90] wl[27] vdd gnd cell_6t
Xbit_r28_c90 bl[90] br[90] wl[28] vdd gnd cell_6t
Xbit_r29_c90 bl[90] br[90] wl[29] vdd gnd cell_6t
Xbit_r30_c90 bl[90] br[90] wl[30] vdd gnd cell_6t
Xbit_r31_c90 bl[90] br[90] wl[31] vdd gnd cell_6t
Xbit_r32_c90 bl[90] br[90] wl[32] vdd gnd cell_6t
Xbit_r33_c90 bl[90] br[90] wl[33] vdd gnd cell_6t
Xbit_r34_c90 bl[90] br[90] wl[34] vdd gnd cell_6t
Xbit_r35_c90 bl[90] br[90] wl[35] vdd gnd cell_6t
Xbit_r36_c90 bl[90] br[90] wl[36] vdd gnd cell_6t
Xbit_r37_c90 bl[90] br[90] wl[37] vdd gnd cell_6t
Xbit_r38_c90 bl[90] br[90] wl[38] vdd gnd cell_6t
Xbit_r39_c90 bl[90] br[90] wl[39] vdd gnd cell_6t
Xbit_r40_c90 bl[90] br[90] wl[40] vdd gnd cell_6t
Xbit_r41_c90 bl[90] br[90] wl[41] vdd gnd cell_6t
Xbit_r42_c90 bl[90] br[90] wl[42] vdd gnd cell_6t
Xbit_r43_c90 bl[90] br[90] wl[43] vdd gnd cell_6t
Xbit_r44_c90 bl[90] br[90] wl[44] vdd gnd cell_6t
Xbit_r45_c90 bl[90] br[90] wl[45] vdd gnd cell_6t
Xbit_r46_c90 bl[90] br[90] wl[46] vdd gnd cell_6t
Xbit_r47_c90 bl[90] br[90] wl[47] vdd gnd cell_6t
Xbit_r48_c90 bl[90] br[90] wl[48] vdd gnd cell_6t
Xbit_r49_c90 bl[90] br[90] wl[49] vdd gnd cell_6t
Xbit_r50_c90 bl[90] br[90] wl[50] vdd gnd cell_6t
Xbit_r51_c90 bl[90] br[90] wl[51] vdd gnd cell_6t
Xbit_r52_c90 bl[90] br[90] wl[52] vdd gnd cell_6t
Xbit_r53_c90 bl[90] br[90] wl[53] vdd gnd cell_6t
Xbit_r54_c90 bl[90] br[90] wl[54] vdd gnd cell_6t
Xbit_r55_c90 bl[90] br[90] wl[55] vdd gnd cell_6t
Xbit_r56_c90 bl[90] br[90] wl[56] vdd gnd cell_6t
Xbit_r57_c90 bl[90] br[90] wl[57] vdd gnd cell_6t
Xbit_r58_c90 bl[90] br[90] wl[58] vdd gnd cell_6t
Xbit_r59_c90 bl[90] br[90] wl[59] vdd gnd cell_6t
Xbit_r60_c90 bl[90] br[90] wl[60] vdd gnd cell_6t
Xbit_r61_c90 bl[90] br[90] wl[61] vdd gnd cell_6t
Xbit_r62_c90 bl[90] br[90] wl[62] vdd gnd cell_6t
Xbit_r63_c90 bl[90] br[90] wl[63] vdd gnd cell_6t
Xbit_r64_c90 bl[90] br[90] wl[64] vdd gnd cell_6t
Xbit_r65_c90 bl[90] br[90] wl[65] vdd gnd cell_6t
Xbit_r66_c90 bl[90] br[90] wl[66] vdd gnd cell_6t
Xbit_r67_c90 bl[90] br[90] wl[67] vdd gnd cell_6t
Xbit_r68_c90 bl[90] br[90] wl[68] vdd gnd cell_6t
Xbit_r69_c90 bl[90] br[90] wl[69] vdd gnd cell_6t
Xbit_r70_c90 bl[90] br[90] wl[70] vdd gnd cell_6t
Xbit_r71_c90 bl[90] br[90] wl[71] vdd gnd cell_6t
Xbit_r72_c90 bl[90] br[90] wl[72] vdd gnd cell_6t
Xbit_r73_c90 bl[90] br[90] wl[73] vdd gnd cell_6t
Xbit_r74_c90 bl[90] br[90] wl[74] vdd gnd cell_6t
Xbit_r75_c90 bl[90] br[90] wl[75] vdd gnd cell_6t
Xbit_r76_c90 bl[90] br[90] wl[76] vdd gnd cell_6t
Xbit_r77_c90 bl[90] br[90] wl[77] vdd gnd cell_6t
Xbit_r78_c90 bl[90] br[90] wl[78] vdd gnd cell_6t
Xbit_r79_c90 bl[90] br[90] wl[79] vdd gnd cell_6t
Xbit_r80_c90 bl[90] br[90] wl[80] vdd gnd cell_6t
Xbit_r81_c90 bl[90] br[90] wl[81] vdd gnd cell_6t
Xbit_r82_c90 bl[90] br[90] wl[82] vdd gnd cell_6t
Xbit_r83_c90 bl[90] br[90] wl[83] vdd gnd cell_6t
Xbit_r84_c90 bl[90] br[90] wl[84] vdd gnd cell_6t
Xbit_r85_c90 bl[90] br[90] wl[85] vdd gnd cell_6t
Xbit_r86_c90 bl[90] br[90] wl[86] vdd gnd cell_6t
Xbit_r87_c90 bl[90] br[90] wl[87] vdd gnd cell_6t
Xbit_r88_c90 bl[90] br[90] wl[88] vdd gnd cell_6t
Xbit_r89_c90 bl[90] br[90] wl[89] vdd gnd cell_6t
Xbit_r90_c90 bl[90] br[90] wl[90] vdd gnd cell_6t
Xbit_r91_c90 bl[90] br[90] wl[91] vdd gnd cell_6t
Xbit_r92_c90 bl[90] br[90] wl[92] vdd gnd cell_6t
Xbit_r93_c90 bl[90] br[90] wl[93] vdd gnd cell_6t
Xbit_r94_c90 bl[90] br[90] wl[94] vdd gnd cell_6t
Xbit_r95_c90 bl[90] br[90] wl[95] vdd gnd cell_6t
Xbit_r96_c90 bl[90] br[90] wl[96] vdd gnd cell_6t
Xbit_r97_c90 bl[90] br[90] wl[97] vdd gnd cell_6t
Xbit_r98_c90 bl[90] br[90] wl[98] vdd gnd cell_6t
Xbit_r99_c90 bl[90] br[90] wl[99] vdd gnd cell_6t
Xbit_r100_c90 bl[90] br[90] wl[100] vdd gnd cell_6t
Xbit_r101_c90 bl[90] br[90] wl[101] vdd gnd cell_6t
Xbit_r102_c90 bl[90] br[90] wl[102] vdd gnd cell_6t
Xbit_r103_c90 bl[90] br[90] wl[103] vdd gnd cell_6t
Xbit_r104_c90 bl[90] br[90] wl[104] vdd gnd cell_6t
Xbit_r105_c90 bl[90] br[90] wl[105] vdd gnd cell_6t
Xbit_r106_c90 bl[90] br[90] wl[106] vdd gnd cell_6t
Xbit_r107_c90 bl[90] br[90] wl[107] vdd gnd cell_6t
Xbit_r108_c90 bl[90] br[90] wl[108] vdd gnd cell_6t
Xbit_r109_c90 bl[90] br[90] wl[109] vdd gnd cell_6t
Xbit_r110_c90 bl[90] br[90] wl[110] vdd gnd cell_6t
Xbit_r111_c90 bl[90] br[90] wl[111] vdd gnd cell_6t
Xbit_r112_c90 bl[90] br[90] wl[112] vdd gnd cell_6t
Xbit_r113_c90 bl[90] br[90] wl[113] vdd gnd cell_6t
Xbit_r114_c90 bl[90] br[90] wl[114] vdd gnd cell_6t
Xbit_r115_c90 bl[90] br[90] wl[115] vdd gnd cell_6t
Xbit_r116_c90 bl[90] br[90] wl[116] vdd gnd cell_6t
Xbit_r117_c90 bl[90] br[90] wl[117] vdd gnd cell_6t
Xbit_r118_c90 bl[90] br[90] wl[118] vdd gnd cell_6t
Xbit_r119_c90 bl[90] br[90] wl[119] vdd gnd cell_6t
Xbit_r120_c90 bl[90] br[90] wl[120] vdd gnd cell_6t
Xbit_r121_c90 bl[90] br[90] wl[121] vdd gnd cell_6t
Xbit_r122_c90 bl[90] br[90] wl[122] vdd gnd cell_6t
Xbit_r123_c90 bl[90] br[90] wl[123] vdd gnd cell_6t
Xbit_r124_c90 bl[90] br[90] wl[124] vdd gnd cell_6t
Xbit_r125_c90 bl[90] br[90] wl[125] vdd gnd cell_6t
Xbit_r126_c90 bl[90] br[90] wl[126] vdd gnd cell_6t
Xbit_r127_c90 bl[90] br[90] wl[127] vdd gnd cell_6t
Xbit_r128_c90 bl[90] br[90] wl[128] vdd gnd cell_6t
Xbit_r129_c90 bl[90] br[90] wl[129] vdd gnd cell_6t
Xbit_r130_c90 bl[90] br[90] wl[130] vdd gnd cell_6t
Xbit_r131_c90 bl[90] br[90] wl[131] vdd gnd cell_6t
Xbit_r132_c90 bl[90] br[90] wl[132] vdd gnd cell_6t
Xbit_r133_c90 bl[90] br[90] wl[133] vdd gnd cell_6t
Xbit_r134_c90 bl[90] br[90] wl[134] vdd gnd cell_6t
Xbit_r135_c90 bl[90] br[90] wl[135] vdd gnd cell_6t
Xbit_r136_c90 bl[90] br[90] wl[136] vdd gnd cell_6t
Xbit_r137_c90 bl[90] br[90] wl[137] vdd gnd cell_6t
Xbit_r138_c90 bl[90] br[90] wl[138] vdd gnd cell_6t
Xbit_r139_c90 bl[90] br[90] wl[139] vdd gnd cell_6t
Xbit_r140_c90 bl[90] br[90] wl[140] vdd gnd cell_6t
Xbit_r141_c90 bl[90] br[90] wl[141] vdd gnd cell_6t
Xbit_r142_c90 bl[90] br[90] wl[142] vdd gnd cell_6t
Xbit_r143_c90 bl[90] br[90] wl[143] vdd gnd cell_6t
Xbit_r144_c90 bl[90] br[90] wl[144] vdd gnd cell_6t
Xbit_r145_c90 bl[90] br[90] wl[145] vdd gnd cell_6t
Xbit_r146_c90 bl[90] br[90] wl[146] vdd gnd cell_6t
Xbit_r147_c90 bl[90] br[90] wl[147] vdd gnd cell_6t
Xbit_r148_c90 bl[90] br[90] wl[148] vdd gnd cell_6t
Xbit_r149_c90 bl[90] br[90] wl[149] vdd gnd cell_6t
Xbit_r150_c90 bl[90] br[90] wl[150] vdd gnd cell_6t
Xbit_r151_c90 bl[90] br[90] wl[151] vdd gnd cell_6t
Xbit_r152_c90 bl[90] br[90] wl[152] vdd gnd cell_6t
Xbit_r153_c90 bl[90] br[90] wl[153] vdd gnd cell_6t
Xbit_r154_c90 bl[90] br[90] wl[154] vdd gnd cell_6t
Xbit_r155_c90 bl[90] br[90] wl[155] vdd gnd cell_6t
Xbit_r156_c90 bl[90] br[90] wl[156] vdd gnd cell_6t
Xbit_r157_c90 bl[90] br[90] wl[157] vdd gnd cell_6t
Xbit_r158_c90 bl[90] br[90] wl[158] vdd gnd cell_6t
Xbit_r159_c90 bl[90] br[90] wl[159] vdd gnd cell_6t
Xbit_r160_c90 bl[90] br[90] wl[160] vdd gnd cell_6t
Xbit_r161_c90 bl[90] br[90] wl[161] vdd gnd cell_6t
Xbit_r162_c90 bl[90] br[90] wl[162] vdd gnd cell_6t
Xbit_r163_c90 bl[90] br[90] wl[163] vdd gnd cell_6t
Xbit_r164_c90 bl[90] br[90] wl[164] vdd gnd cell_6t
Xbit_r165_c90 bl[90] br[90] wl[165] vdd gnd cell_6t
Xbit_r166_c90 bl[90] br[90] wl[166] vdd gnd cell_6t
Xbit_r167_c90 bl[90] br[90] wl[167] vdd gnd cell_6t
Xbit_r168_c90 bl[90] br[90] wl[168] vdd gnd cell_6t
Xbit_r169_c90 bl[90] br[90] wl[169] vdd gnd cell_6t
Xbit_r170_c90 bl[90] br[90] wl[170] vdd gnd cell_6t
Xbit_r171_c90 bl[90] br[90] wl[171] vdd gnd cell_6t
Xbit_r172_c90 bl[90] br[90] wl[172] vdd gnd cell_6t
Xbit_r173_c90 bl[90] br[90] wl[173] vdd gnd cell_6t
Xbit_r174_c90 bl[90] br[90] wl[174] vdd gnd cell_6t
Xbit_r175_c90 bl[90] br[90] wl[175] vdd gnd cell_6t
Xbit_r176_c90 bl[90] br[90] wl[176] vdd gnd cell_6t
Xbit_r177_c90 bl[90] br[90] wl[177] vdd gnd cell_6t
Xbit_r178_c90 bl[90] br[90] wl[178] vdd gnd cell_6t
Xbit_r179_c90 bl[90] br[90] wl[179] vdd gnd cell_6t
Xbit_r180_c90 bl[90] br[90] wl[180] vdd gnd cell_6t
Xbit_r181_c90 bl[90] br[90] wl[181] vdd gnd cell_6t
Xbit_r182_c90 bl[90] br[90] wl[182] vdd gnd cell_6t
Xbit_r183_c90 bl[90] br[90] wl[183] vdd gnd cell_6t
Xbit_r184_c90 bl[90] br[90] wl[184] vdd gnd cell_6t
Xbit_r185_c90 bl[90] br[90] wl[185] vdd gnd cell_6t
Xbit_r186_c90 bl[90] br[90] wl[186] vdd gnd cell_6t
Xbit_r187_c90 bl[90] br[90] wl[187] vdd gnd cell_6t
Xbit_r188_c90 bl[90] br[90] wl[188] vdd gnd cell_6t
Xbit_r189_c90 bl[90] br[90] wl[189] vdd gnd cell_6t
Xbit_r190_c90 bl[90] br[90] wl[190] vdd gnd cell_6t
Xbit_r191_c90 bl[90] br[90] wl[191] vdd gnd cell_6t
Xbit_r192_c90 bl[90] br[90] wl[192] vdd gnd cell_6t
Xbit_r193_c90 bl[90] br[90] wl[193] vdd gnd cell_6t
Xbit_r194_c90 bl[90] br[90] wl[194] vdd gnd cell_6t
Xbit_r195_c90 bl[90] br[90] wl[195] vdd gnd cell_6t
Xbit_r196_c90 bl[90] br[90] wl[196] vdd gnd cell_6t
Xbit_r197_c90 bl[90] br[90] wl[197] vdd gnd cell_6t
Xbit_r198_c90 bl[90] br[90] wl[198] vdd gnd cell_6t
Xbit_r199_c90 bl[90] br[90] wl[199] vdd gnd cell_6t
Xbit_r200_c90 bl[90] br[90] wl[200] vdd gnd cell_6t
Xbit_r201_c90 bl[90] br[90] wl[201] vdd gnd cell_6t
Xbit_r202_c90 bl[90] br[90] wl[202] vdd gnd cell_6t
Xbit_r203_c90 bl[90] br[90] wl[203] vdd gnd cell_6t
Xbit_r204_c90 bl[90] br[90] wl[204] vdd gnd cell_6t
Xbit_r205_c90 bl[90] br[90] wl[205] vdd gnd cell_6t
Xbit_r206_c90 bl[90] br[90] wl[206] vdd gnd cell_6t
Xbit_r207_c90 bl[90] br[90] wl[207] vdd gnd cell_6t
Xbit_r208_c90 bl[90] br[90] wl[208] vdd gnd cell_6t
Xbit_r209_c90 bl[90] br[90] wl[209] vdd gnd cell_6t
Xbit_r210_c90 bl[90] br[90] wl[210] vdd gnd cell_6t
Xbit_r211_c90 bl[90] br[90] wl[211] vdd gnd cell_6t
Xbit_r212_c90 bl[90] br[90] wl[212] vdd gnd cell_6t
Xbit_r213_c90 bl[90] br[90] wl[213] vdd gnd cell_6t
Xbit_r214_c90 bl[90] br[90] wl[214] vdd gnd cell_6t
Xbit_r215_c90 bl[90] br[90] wl[215] vdd gnd cell_6t
Xbit_r216_c90 bl[90] br[90] wl[216] vdd gnd cell_6t
Xbit_r217_c90 bl[90] br[90] wl[217] vdd gnd cell_6t
Xbit_r218_c90 bl[90] br[90] wl[218] vdd gnd cell_6t
Xbit_r219_c90 bl[90] br[90] wl[219] vdd gnd cell_6t
Xbit_r220_c90 bl[90] br[90] wl[220] vdd gnd cell_6t
Xbit_r221_c90 bl[90] br[90] wl[221] vdd gnd cell_6t
Xbit_r222_c90 bl[90] br[90] wl[222] vdd gnd cell_6t
Xbit_r223_c90 bl[90] br[90] wl[223] vdd gnd cell_6t
Xbit_r224_c90 bl[90] br[90] wl[224] vdd gnd cell_6t
Xbit_r225_c90 bl[90] br[90] wl[225] vdd gnd cell_6t
Xbit_r226_c90 bl[90] br[90] wl[226] vdd gnd cell_6t
Xbit_r227_c90 bl[90] br[90] wl[227] vdd gnd cell_6t
Xbit_r228_c90 bl[90] br[90] wl[228] vdd gnd cell_6t
Xbit_r229_c90 bl[90] br[90] wl[229] vdd gnd cell_6t
Xbit_r230_c90 bl[90] br[90] wl[230] vdd gnd cell_6t
Xbit_r231_c90 bl[90] br[90] wl[231] vdd gnd cell_6t
Xbit_r232_c90 bl[90] br[90] wl[232] vdd gnd cell_6t
Xbit_r233_c90 bl[90] br[90] wl[233] vdd gnd cell_6t
Xbit_r234_c90 bl[90] br[90] wl[234] vdd gnd cell_6t
Xbit_r235_c90 bl[90] br[90] wl[235] vdd gnd cell_6t
Xbit_r236_c90 bl[90] br[90] wl[236] vdd gnd cell_6t
Xbit_r237_c90 bl[90] br[90] wl[237] vdd gnd cell_6t
Xbit_r238_c90 bl[90] br[90] wl[238] vdd gnd cell_6t
Xbit_r239_c90 bl[90] br[90] wl[239] vdd gnd cell_6t
Xbit_r240_c90 bl[90] br[90] wl[240] vdd gnd cell_6t
Xbit_r241_c90 bl[90] br[90] wl[241] vdd gnd cell_6t
Xbit_r242_c90 bl[90] br[90] wl[242] vdd gnd cell_6t
Xbit_r243_c90 bl[90] br[90] wl[243] vdd gnd cell_6t
Xbit_r244_c90 bl[90] br[90] wl[244] vdd gnd cell_6t
Xbit_r245_c90 bl[90] br[90] wl[245] vdd gnd cell_6t
Xbit_r246_c90 bl[90] br[90] wl[246] vdd gnd cell_6t
Xbit_r247_c90 bl[90] br[90] wl[247] vdd gnd cell_6t
Xbit_r248_c90 bl[90] br[90] wl[248] vdd gnd cell_6t
Xbit_r249_c90 bl[90] br[90] wl[249] vdd gnd cell_6t
Xbit_r250_c90 bl[90] br[90] wl[250] vdd gnd cell_6t
Xbit_r251_c90 bl[90] br[90] wl[251] vdd gnd cell_6t
Xbit_r252_c90 bl[90] br[90] wl[252] vdd gnd cell_6t
Xbit_r253_c90 bl[90] br[90] wl[253] vdd gnd cell_6t
Xbit_r254_c90 bl[90] br[90] wl[254] vdd gnd cell_6t
Xbit_r255_c90 bl[90] br[90] wl[255] vdd gnd cell_6t
Xbit_r0_c91 bl[91] br[91] wl[0] vdd gnd cell_6t
Xbit_r1_c91 bl[91] br[91] wl[1] vdd gnd cell_6t
Xbit_r2_c91 bl[91] br[91] wl[2] vdd gnd cell_6t
Xbit_r3_c91 bl[91] br[91] wl[3] vdd gnd cell_6t
Xbit_r4_c91 bl[91] br[91] wl[4] vdd gnd cell_6t
Xbit_r5_c91 bl[91] br[91] wl[5] vdd gnd cell_6t
Xbit_r6_c91 bl[91] br[91] wl[6] vdd gnd cell_6t
Xbit_r7_c91 bl[91] br[91] wl[7] vdd gnd cell_6t
Xbit_r8_c91 bl[91] br[91] wl[8] vdd gnd cell_6t
Xbit_r9_c91 bl[91] br[91] wl[9] vdd gnd cell_6t
Xbit_r10_c91 bl[91] br[91] wl[10] vdd gnd cell_6t
Xbit_r11_c91 bl[91] br[91] wl[11] vdd gnd cell_6t
Xbit_r12_c91 bl[91] br[91] wl[12] vdd gnd cell_6t
Xbit_r13_c91 bl[91] br[91] wl[13] vdd gnd cell_6t
Xbit_r14_c91 bl[91] br[91] wl[14] vdd gnd cell_6t
Xbit_r15_c91 bl[91] br[91] wl[15] vdd gnd cell_6t
Xbit_r16_c91 bl[91] br[91] wl[16] vdd gnd cell_6t
Xbit_r17_c91 bl[91] br[91] wl[17] vdd gnd cell_6t
Xbit_r18_c91 bl[91] br[91] wl[18] vdd gnd cell_6t
Xbit_r19_c91 bl[91] br[91] wl[19] vdd gnd cell_6t
Xbit_r20_c91 bl[91] br[91] wl[20] vdd gnd cell_6t
Xbit_r21_c91 bl[91] br[91] wl[21] vdd gnd cell_6t
Xbit_r22_c91 bl[91] br[91] wl[22] vdd gnd cell_6t
Xbit_r23_c91 bl[91] br[91] wl[23] vdd gnd cell_6t
Xbit_r24_c91 bl[91] br[91] wl[24] vdd gnd cell_6t
Xbit_r25_c91 bl[91] br[91] wl[25] vdd gnd cell_6t
Xbit_r26_c91 bl[91] br[91] wl[26] vdd gnd cell_6t
Xbit_r27_c91 bl[91] br[91] wl[27] vdd gnd cell_6t
Xbit_r28_c91 bl[91] br[91] wl[28] vdd gnd cell_6t
Xbit_r29_c91 bl[91] br[91] wl[29] vdd gnd cell_6t
Xbit_r30_c91 bl[91] br[91] wl[30] vdd gnd cell_6t
Xbit_r31_c91 bl[91] br[91] wl[31] vdd gnd cell_6t
Xbit_r32_c91 bl[91] br[91] wl[32] vdd gnd cell_6t
Xbit_r33_c91 bl[91] br[91] wl[33] vdd gnd cell_6t
Xbit_r34_c91 bl[91] br[91] wl[34] vdd gnd cell_6t
Xbit_r35_c91 bl[91] br[91] wl[35] vdd gnd cell_6t
Xbit_r36_c91 bl[91] br[91] wl[36] vdd gnd cell_6t
Xbit_r37_c91 bl[91] br[91] wl[37] vdd gnd cell_6t
Xbit_r38_c91 bl[91] br[91] wl[38] vdd gnd cell_6t
Xbit_r39_c91 bl[91] br[91] wl[39] vdd gnd cell_6t
Xbit_r40_c91 bl[91] br[91] wl[40] vdd gnd cell_6t
Xbit_r41_c91 bl[91] br[91] wl[41] vdd gnd cell_6t
Xbit_r42_c91 bl[91] br[91] wl[42] vdd gnd cell_6t
Xbit_r43_c91 bl[91] br[91] wl[43] vdd gnd cell_6t
Xbit_r44_c91 bl[91] br[91] wl[44] vdd gnd cell_6t
Xbit_r45_c91 bl[91] br[91] wl[45] vdd gnd cell_6t
Xbit_r46_c91 bl[91] br[91] wl[46] vdd gnd cell_6t
Xbit_r47_c91 bl[91] br[91] wl[47] vdd gnd cell_6t
Xbit_r48_c91 bl[91] br[91] wl[48] vdd gnd cell_6t
Xbit_r49_c91 bl[91] br[91] wl[49] vdd gnd cell_6t
Xbit_r50_c91 bl[91] br[91] wl[50] vdd gnd cell_6t
Xbit_r51_c91 bl[91] br[91] wl[51] vdd gnd cell_6t
Xbit_r52_c91 bl[91] br[91] wl[52] vdd gnd cell_6t
Xbit_r53_c91 bl[91] br[91] wl[53] vdd gnd cell_6t
Xbit_r54_c91 bl[91] br[91] wl[54] vdd gnd cell_6t
Xbit_r55_c91 bl[91] br[91] wl[55] vdd gnd cell_6t
Xbit_r56_c91 bl[91] br[91] wl[56] vdd gnd cell_6t
Xbit_r57_c91 bl[91] br[91] wl[57] vdd gnd cell_6t
Xbit_r58_c91 bl[91] br[91] wl[58] vdd gnd cell_6t
Xbit_r59_c91 bl[91] br[91] wl[59] vdd gnd cell_6t
Xbit_r60_c91 bl[91] br[91] wl[60] vdd gnd cell_6t
Xbit_r61_c91 bl[91] br[91] wl[61] vdd gnd cell_6t
Xbit_r62_c91 bl[91] br[91] wl[62] vdd gnd cell_6t
Xbit_r63_c91 bl[91] br[91] wl[63] vdd gnd cell_6t
Xbit_r64_c91 bl[91] br[91] wl[64] vdd gnd cell_6t
Xbit_r65_c91 bl[91] br[91] wl[65] vdd gnd cell_6t
Xbit_r66_c91 bl[91] br[91] wl[66] vdd gnd cell_6t
Xbit_r67_c91 bl[91] br[91] wl[67] vdd gnd cell_6t
Xbit_r68_c91 bl[91] br[91] wl[68] vdd gnd cell_6t
Xbit_r69_c91 bl[91] br[91] wl[69] vdd gnd cell_6t
Xbit_r70_c91 bl[91] br[91] wl[70] vdd gnd cell_6t
Xbit_r71_c91 bl[91] br[91] wl[71] vdd gnd cell_6t
Xbit_r72_c91 bl[91] br[91] wl[72] vdd gnd cell_6t
Xbit_r73_c91 bl[91] br[91] wl[73] vdd gnd cell_6t
Xbit_r74_c91 bl[91] br[91] wl[74] vdd gnd cell_6t
Xbit_r75_c91 bl[91] br[91] wl[75] vdd gnd cell_6t
Xbit_r76_c91 bl[91] br[91] wl[76] vdd gnd cell_6t
Xbit_r77_c91 bl[91] br[91] wl[77] vdd gnd cell_6t
Xbit_r78_c91 bl[91] br[91] wl[78] vdd gnd cell_6t
Xbit_r79_c91 bl[91] br[91] wl[79] vdd gnd cell_6t
Xbit_r80_c91 bl[91] br[91] wl[80] vdd gnd cell_6t
Xbit_r81_c91 bl[91] br[91] wl[81] vdd gnd cell_6t
Xbit_r82_c91 bl[91] br[91] wl[82] vdd gnd cell_6t
Xbit_r83_c91 bl[91] br[91] wl[83] vdd gnd cell_6t
Xbit_r84_c91 bl[91] br[91] wl[84] vdd gnd cell_6t
Xbit_r85_c91 bl[91] br[91] wl[85] vdd gnd cell_6t
Xbit_r86_c91 bl[91] br[91] wl[86] vdd gnd cell_6t
Xbit_r87_c91 bl[91] br[91] wl[87] vdd gnd cell_6t
Xbit_r88_c91 bl[91] br[91] wl[88] vdd gnd cell_6t
Xbit_r89_c91 bl[91] br[91] wl[89] vdd gnd cell_6t
Xbit_r90_c91 bl[91] br[91] wl[90] vdd gnd cell_6t
Xbit_r91_c91 bl[91] br[91] wl[91] vdd gnd cell_6t
Xbit_r92_c91 bl[91] br[91] wl[92] vdd gnd cell_6t
Xbit_r93_c91 bl[91] br[91] wl[93] vdd gnd cell_6t
Xbit_r94_c91 bl[91] br[91] wl[94] vdd gnd cell_6t
Xbit_r95_c91 bl[91] br[91] wl[95] vdd gnd cell_6t
Xbit_r96_c91 bl[91] br[91] wl[96] vdd gnd cell_6t
Xbit_r97_c91 bl[91] br[91] wl[97] vdd gnd cell_6t
Xbit_r98_c91 bl[91] br[91] wl[98] vdd gnd cell_6t
Xbit_r99_c91 bl[91] br[91] wl[99] vdd gnd cell_6t
Xbit_r100_c91 bl[91] br[91] wl[100] vdd gnd cell_6t
Xbit_r101_c91 bl[91] br[91] wl[101] vdd gnd cell_6t
Xbit_r102_c91 bl[91] br[91] wl[102] vdd gnd cell_6t
Xbit_r103_c91 bl[91] br[91] wl[103] vdd gnd cell_6t
Xbit_r104_c91 bl[91] br[91] wl[104] vdd gnd cell_6t
Xbit_r105_c91 bl[91] br[91] wl[105] vdd gnd cell_6t
Xbit_r106_c91 bl[91] br[91] wl[106] vdd gnd cell_6t
Xbit_r107_c91 bl[91] br[91] wl[107] vdd gnd cell_6t
Xbit_r108_c91 bl[91] br[91] wl[108] vdd gnd cell_6t
Xbit_r109_c91 bl[91] br[91] wl[109] vdd gnd cell_6t
Xbit_r110_c91 bl[91] br[91] wl[110] vdd gnd cell_6t
Xbit_r111_c91 bl[91] br[91] wl[111] vdd gnd cell_6t
Xbit_r112_c91 bl[91] br[91] wl[112] vdd gnd cell_6t
Xbit_r113_c91 bl[91] br[91] wl[113] vdd gnd cell_6t
Xbit_r114_c91 bl[91] br[91] wl[114] vdd gnd cell_6t
Xbit_r115_c91 bl[91] br[91] wl[115] vdd gnd cell_6t
Xbit_r116_c91 bl[91] br[91] wl[116] vdd gnd cell_6t
Xbit_r117_c91 bl[91] br[91] wl[117] vdd gnd cell_6t
Xbit_r118_c91 bl[91] br[91] wl[118] vdd gnd cell_6t
Xbit_r119_c91 bl[91] br[91] wl[119] vdd gnd cell_6t
Xbit_r120_c91 bl[91] br[91] wl[120] vdd gnd cell_6t
Xbit_r121_c91 bl[91] br[91] wl[121] vdd gnd cell_6t
Xbit_r122_c91 bl[91] br[91] wl[122] vdd gnd cell_6t
Xbit_r123_c91 bl[91] br[91] wl[123] vdd gnd cell_6t
Xbit_r124_c91 bl[91] br[91] wl[124] vdd gnd cell_6t
Xbit_r125_c91 bl[91] br[91] wl[125] vdd gnd cell_6t
Xbit_r126_c91 bl[91] br[91] wl[126] vdd gnd cell_6t
Xbit_r127_c91 bl[91] br[91] wl[127] vdd gnd cell_6t
Xbit_r128_c91 bl[91] br[91] wl[128] vdd gnd cell_6t
Xbit_r129_c91 bl[91] br[91] wl[129] vdd gnd cell_6t
Xbit_r130_c91 bl[91] br[91] wl[130] vdd gnd cell_6t
Xbit_r131_c91 bl[91] br[91] wl[131] vdd gnd cell_6t
Xbit_r132_c91 bl[91] br[91] wl[132] vdd gnd cell_6t
Xbit_r133_c91 bl[91] br[91] wl[133] vdd gnd cell_6t
Xbit_r134_c91 bl[91] br[91] wl[134] vdd gnd cell_6t
Xbit_r135_c91 bl[91] br[91] wl[135] vdd gnd cell_6t
Xbit_r136_c91 bl[91] br[91] wl[136] vdd gnd cell_6t
Xbit_r137_c91 bl[91] br[91] wl[137] vdd gnd cell_6t
Xbit_r138_c91 bl[91] br[91] wl[138] vdd gnd cell_6t
Xbit_r139_c91 bl[91] br[91] wl[139] vdd gnd cell_6t
Xbit_r140_c91 bl[91] br[91] wl[140] vdd gnd cell_6t
Xbit_r141_c91 bl[91] br[91] wl[141] vdd gnd cell_6t
Xbit_r142_c91 bl[91] br[91] wl[142] vdd gnd cell_6t
Xbit_r143_c91 bl[91] br[91] wl[143] vdd gnd cell_6t
Xbit_r144_c91 bl[91] br[91] wl[144] vdd gnd cell_6t
Xbit_r145_c91 bl[91] br[91] wl[145] vdd gnd cell_6t
Xbit_r146_c91 bl[91] br[91] wl[146] vdd gnd cell_6t
Xbit_r147_c91 bl[91] br[91] wl[147] vdd gnd cell_6t
Xbit_r148_c91 bl[91] br[91] wl[148] vdd gnd cell_6t
Xbit_r149_c91 bl[91] br[91] wl[149] vdd gnd cell_6t
Xbit_r150_c91 bl[91] br[91] wl[150] vdd gnd cell_6t
Xbit_r151_c91 bl[91] br[91] wl[151] vdd gnd cell_6t
Xbit_r152_c91 bl[91] br[91] wl[152] vdd gnd cell_6t
Xbit_r153_c91 bl[91] br[91] wl[153] vdd gnd cell_6t
Xbit_r154_c91 bl[91] br[91] wl[154] vdd gnd cell_6t
Xbit_r155_c91 bl[91] br[91] wl[155] vdd gnd cell_6t
Xbit_r156_c91 bl[91] br[91] wl[156] vdd gnd cell_6t
Xbit_r157_c91 bl[91] br[91] wl[157] vdd gnd cell_6t
Xbit_r158_c91 bl[91] br[91] wl[158] vdd gnd cell_6t
Xbit_r159_c91 bl[91] br[91] wl[159] vdd gnd cell_6t
Xbit_r160_c91 bl[91] br[91] wl[160] vdd gnd cell_6t
Xbit_r161_c91 bl[91] br[91] wl[161] vdd gnd cell_6t
Xbit_r162_c91 bl[91] br[91] wl[162] vdd gnd cell_6t
Xbit_r163_c91 bl[91] br[91] wl[163] vdd gnd cell_6t
Xbit_r164_c91 bl[91] br[91] wl[164] vdd gnd cell_6t
Xbit_r165_c91 bl[91] br[91] wl[165] vdd gnd cell_6t
Xbit_r166_c91 bl[91] br[91] wl[166] vdd gnd cell_6t
Xbit_r167_c91 bl[91] br[91] wl[167] vdd gnd cell_6t
Xbit_r168_c91 bl[91] br[91] wl[168] vdd gnd cell_6t
Xbit_r169_c91 bl[91] br[91] wl[169] vdd gnd cell_6t
Xbit_r170_c91 bl[91] br[91] wl[170] vdd gnd cell_6t
Xbit_r171_c91 bl[91] br[91] wl[171] vdd gnd cell_6t
Xbit_r172_c91 bl[91] br[91] wl[172] vdd gnd cell_6t
Xbit_r173_c91 bl[91] br[91] wl[173] vdd gnd cell_6t
Xbit_r174_c91 bl[91] br[91] wl[174] vdd gnd cell_6t
Xbit_r175_c91 bl[91] br[91] wl[175] vdd gnd cell_6t
Xbit_r176_c91 bl[91] br[91] wl[176] vdd gnd cell_6t
Xbit_r177_c91 bl[91] br[91] wl[177] vdd gnd cell_6t
Xbit_r178_c91 bl[91] br[91] wl[178] vdd gnd cell_6t
Xbit_r179_c91 bl[91] br[91] wl[179] vdd gnd cell_6t
Xbit_r180_c91 bl[91] br[91] wl[180] vdd gnd cell_6t
Xbit_r181_c91 bl[91] br[91] wl[181] vdd gnd cell_6t
Xbit_r182_c91 bl[91] br[91] wl[182] vdd gnd cell_6t
Xbit_r183_c91 bl[91] br[91] wl[183] vdd gnd cell_6t
Xbit_r184_c91 bl[91] br[91] wl[184] vdd gnd cell_6t
Xbit_r185_c91 bl[91] br[91] wl[185] vdd gnd cell_6t
Xbit_r186_c91 bl[91] br[91] wl[186] vdd gnd cell_6t
Xbit_r187_c91 bl[91] br[91] wl[187] vdd gnd cell_6t
Xbit_r188_c91 bl[91] br[91] wl[188] vdd gnd cell_6t
Xbit_r189_c91 bl[91] br[91] wl[189] vdd gnd cell_6t
Xbit_r190_c91 bl[91] br[91] wl[190] vdd gnd cell_6t
Xbit_r191_c91 bl[91] br[91] wl[191] vdd gnd cell_6t
Xbit_r192_c91 bl[91] br[91] wl[192] vdd gnd cell_6t
Xbit_r193_c91 bl[91] br[91] wl[193] vdd gnd cell_6t
Xbit_r194_c91 bl[91] br[91] wl[194] vdd gnd cell_6t
Xbit_r195_c91 bl[91] br[91] wl[195] vdd gnd cell_6t
Xbit_r196_c91 bl[91] br[91] wl[196] vdd gnd cell_6t
Xbit_r197_c91 bl[91] br[91] wl[197] vdd gnd cell_6t
Xbit_r198_c91 bl[91] br[91] wl[198] vdd gnd cell_6t
Xbit_r199_c91 bl[91] br[91] wl[199] vdd gnd cell_6t
Xbit_r200_c91 bl[91] br[91] wl[200] vdd gnd cell_6t
Xbit_r201_c91 bl[91] br[91] wl[201] vdd gnd cell_6t
Xbit_r202_c91 bl[91] br[91] wl[202] vdd gnd cell_6t
Xbit_r203_c91 bl[91] br[91] wl[203] vdd gnd cell_6t
Xbit_r204_c91 bl[91] br[91] wl[204] vdd gnd cell_6t
Xbit_r205_c91 bl[91] br[91] wl[205] vdd gnd cell_6t
Xbit_r206_c91 bl[91] br[91] wl[206] vdd gnd cell_6t
Xbit_r207_c91 bl[91] br[91] wl[207] vdd gnd cell_6t
Xbit_r208_c91 bl[91] br[91] wl[208] vdd gnd cell_6t
Xbit_r209_c91 bl[91] br[91] wl[209] vdd gnd cell_6t
Xbit_r210_c91 bl[91] br[91] wl[210] vdd gnd cell_6t
Xbit_r211_c91 bl[91] br[91] wl[211] vdd gnd cell_6t
Xbit_r212_c91 bl[91] br[91] wl[212] vdd gnd cell_6t
Xbit_r213_c91 bl[91] br[91] wl[213] vdd gnd cell_6t
Xbit_r214_c91 bl[91] br[91] wl[214] vdd gnd cell_6t
Xbit_r215_c91 bl[91] br[91] wl[215] vdd gnd cell_6t
Xbit_r216_c91 bl[91] br[91] wl[216] vdd gnd cell_6t
Xbit_r217_c91 bl[91] br[91] wl[217] vdd gnd cell_6t
Xbit_r218_c91 bl[91] br[91] wl[218] vdd gnd cell_6t
Xbit_r219_c91 bl[91] br[91] wl[219] vdd gnd cell_6t
Xbit_r220_c91 bl[91] br[91] wl[220] vdd gnd cell_6t
Xbit_r221_c91 bl[91] br[91] wl[221] vdd gnd cell_6t
Xbit_r222_c91 bl[91] br[91] wl[222] vdd gnd cell_6t
Xbit_r223_c91 bl[91] br[91] wl[223] vdd gnd cell_6t
Xbit_r224_c91 bl[91] br[91] wl[224] vdd gnd cell_6t
Xbit_r225_c91 bl[91] br[91] wl[225] vdd gnd cell_6t
Xbit_r226_c91 bl[91] br[91] wl[226] vdd gnd cell_6t
Xbit_r227_c91 bl[91] br[91] wl[227] vdd gnd cell_6t
Xbit_r228_c91 bl[91] br[91] wl[228] vdd gnd cell_6t
Xbit_r229_c91 bl[91] br[91] wl[229] vdd gnd cell_6t
Xbit_r230_c91 bl[91] br[91] wl[230] vdd gnd cell_6t
Xbit_r231_c91 bl[91] br[91] wl[231] vdd gnd cell_6t
Xbit_r232_c91 bl[91] br[91] wl[232] vdd gnd cell_6t
Xbit_r233_c91 bl[91] br[91] wl[233] vdd gnd cell_6t
Xbit_r234_c91 bl[91] br[91] wl[234] vdd gnd cell_6t
Xbit_r235_c91 bl[91] br[91] wl[235] vdd gnd cell_6t
Xbit_r236_c91 bl[91] br[91] wl[236] vdd gnd cell_6t
Xbit_r237_c91 bl[91] br[91] wl[237] vdd gnd cell_6t
Xbit_r238_c91 bl[91] br[91] wl[238] vdd gnd cell_6t
Xbit_r239_c91 bl[91] br[91] wl[239] vdd gnd cell_6t
Xbit_r240_c91 bl[91] br[91] wl[240] vdd gnd cell_6t
Xbit_r241_c91 bl[91] br[91] wl[241] vdd gnd cell_6t
Xbit_r242_c91 bl[91] br[91] wl[242] vdd gnd cell_6t
Xbit_r243_c91 bl[91] br[91] wl[243] vdd gnd cell_6t
Xbit_r244_c91 bl[91] br[91] wl[244] vdd gnd cell_6t
Xbit_r245_c91 bl[91] br[91] wl[245] vdd gnd cell_6t
Xbit_r246_c91 bl[91] br[91] wl[246] vdd gnd cell_6t
Xbit_r247_c91 bl[91] br[91] wl[247] vdd gnd cell_6t
Xbit_r248_c91 bl[91] br[91] wl[248] vdd gnd cell_6t
Xbit_r249_c91 bl[91] br[91] wl[249] vdd gnd cell_6t
Xbit_r250_c91 bl[91] br[91] wl[250] vdd gnd cell_6t
Xbit_r251_c91 bl[91] br[91] wl[251] vdd gnd cell_6t
Xbit_r252_c91 bl[91] br[91] wl[252] vdd gnd cell_6t
Xbit_r253_c91 bl[91] br[91] wl[253] vdd gnd cell_6t
Xbit_r254_c91 bl[91] br[91] wl[254] vdd gnd cell_6t
Xbit_r255_c91 bl[91] br[91] wl[255] vdd gnd cell_6t
Xbit_r0_c92 bl[92] br[92] wl[0] vdd gnd cell_6t
Xbit_r1_c92 bl[92] br[92] wl[1] vdd gnd cell_6t
Xbit_r2_c92 bl[92] br[92] wl[2] vdd gnd cell_6t
Xbit_r3_c92 bl[92] br[92] wl[3] vdd gnd cell_6t
Xbit_r4_c92 bl[92] br[92] wl[4] vdd gnd cell_6t
Xbit_r5_c92 bl[92] br[92] wl[5] vdd gnd cell_6t
Xbit_r6_c92 bl[92] br[92] wl[6] vdd gnd cell_6t
Xbit_r7_c92 bl[92] br[92] wl[7] vdd gnd cell_6t
Xbit_r8_c92 bl[92] br[92] wl[8] vdd gnd cell_6t
Xbit_r9_c92 bl[92] br[92] wl[9] vdd gnd cell_6t
Xbit_r10_c92 bl[92] br[92] wl[10] vdd gnd cell_6t
Xbit_r11_c92 bl[92] br[92] wl[11] vdd gnd cell_6t
Xbit_r12_c92 bl[92] br[92] wl[12] vdd gnd cell_6t
Xbit_r13_c92 bl[92] br[92] wl[13] vdd gnd cell_6t
Xbit_r14_c92 bl[92] br[92] wl[14] vdd gnd cell_6t
Xbit_r15_c92 bl[92] br[92] wl[15] vdd gnd cell_6t
Xbit_r16_c92 bl[92] br[92] wl[16] vdd gnd cell_6t
Xbit_r17_c92 bl[92] br[92] wl[17] vdd gnd cell_6t
Xbit_r18_c92 bl[92] br[92] wl[18] vdd gnd cell_6t
Xbit_r19_c92 bl[92] br[92] wl[19] vdd gnd cell_6t
Xbit_r20_c92 bl[92] br[92] wl[20] vdd gnd cell_6t
Xbit_r21_c92 bl[92] br[92] wl[21] vdd gnd cell_6t
Xbit_r22_c92 bl[92] br[92] wl[22] vdd gnd cell_6t
Xbit_r23_c92 bl[92] br[92] wl[23] vdd gnd cell_6t
Xbit_r24_c92 bl[92] br[92] wl[24] vdd gnd cell_6t
Xbit_r25_c92 bl[92] br[92] wl[25] vdd gnd cell_6t
Xbit_r26_c92 bl[92] br[92] wl[26] vdd gnd cell_6t
Xbit_r27_c92 bl[92] br[92] wl[27] vdd gnd cell_6t
Xbit_r28_c92 bl[92] br[92] wl[28] vdd gnd cell_6t
Xbit_r29_c92 bl[92] br[92] wl[29] vdd gnd cell_6t
Xbit_r30_c92 bl[92] br[92] wl[30] vdd gnd cell_6t
Xbit_r31_c92 bl[92] br[92] wl[31] vdd gnd cell_6t
Xbit_r32_c92 bl[92] br[92] wl[32] vdd gnd cell_6t
Xbit_r33_c92 bl[92] br[92] wl[33] vdd gnd cell_6t
Xbit_r34_c92 bl[92] br[92] wl[34] vdd gnd cell_6t
Xbit_r35_c92 bl[92] br[92] wl[35] vdd gnd cell_6t
Xbit_r36_c92 bl[92] br[92] wl[36] vdd gnd cell_6t
Xbit_r37_c92 bl[92] br[92] wl[37] vdd gnd cell_6t
Xbit_r38_c92 bl[92] br[92] wl[38] vdd gnd cell_6t
Xbit_r39_c92 bl[92] br[92] wl[39] vdd gnd cell_6t
Xbit_r40_c92 bl[92] br[92] wl[40] vdd gnd cell_6t
Xbit_r41_c92 bl[92] br[92] wl[41] vdd gnd cell_6t
Xbit_r42_c92 bl[92] br[92] wl[42] vdd gnd cell_6t
Xbit_r43_c92 bl[92] br[92] wl[43] vdd gnd cell_6t
Xbit_r44_c92 bl[92] br[92] wl[44] vdd gnd cell_6t
Xbit_r45_c92 bl[92] br[92] wl[45] vdd gnd cell_6t
Xbit_r46_c92 bl[92] br[92] wl[46] vdd gnd cell_6t
Xbit_r47_c92 bl[92] br[92] wl[47] vdd gnd cell_6t
Xbit_r48_c92 bl[92] br[92] wl[48] vdd gnd cell_6t
Xbit_r49_c92 bl[92] br[92] wl[49] vdd gnd cell_6t
Xbit_r50_c92 bl[92] br[92] wl[50] vdd gnd cell_6t
Xbit_r51_c92 bl[92] br[92] wl[51] vdd gnd cell_6t
Xbit_r52_c92 bl[92] br[92] wl[52] vdd gnd cell_6t
Xbit_r53_c92 bl[92] br[92] wl[53] vdd gnd cell_6t
Xbit_r54_c92 bl[92] br[92] wl[54] vdd gnd cell_6t
Xbit_r55_c92 bl[92] br[92] wl[55] vdd gnd cell_6t
Xbit_r56_c92 bl[92] br[92] wl[56] vdd gnd cell_6t
Xbit_r57_c92 bl[92] br[92] wl[57] vdd gnd cell_6t
Xbit_r58_c92 bl[92] br[92] wl[58] vdd gnd cell_6t
Xbit_r59_c92 bl[92] br[92] wl[59] vdd gnd cell_6t
Xbit_r60_c92 bl[92] br[92] wl[60] vdd gnd cell_6t
Xbit_r61_c92 bl[92] br[92] wl[61] vdd gnd cell_6t
Xbit_r62_c92 bl[92] br[92] wl[62] vdd gnd cell_6t
Xbit_r63_c92 bl[92] br[92] wl[63] vdd gnd cell_6t
Xbit_r64_c92 bl[92] br[92] wl[64] vdd gnd cell_6t
Xbit_r65_c92 bl[92] br[92] wl[65] vdd gnd cell_6t
Xbit_r66_c92 bl[92] br[92] wl[66] vdd gnd cell_6t
Xbit_r67_c92 bl[92] br[92] wl[67] vdd gnd cell_6t
Xbit_r68_c92 bl[92] br[92] wl[68] vdd gnd cell_6t
Xbit_r69_c92 bl[92] br[92] wl[69] vdd gnd cell_6t
Xbit_r70_c92 bl[92] br[92] wl[70] vdd gnd cell_6t
Xbit_r71_c92 bl[92] br[92] wl[71] vdd gnd cell_6t
Xbit_r72_c92 bl[92] br[92] wl[72] vdd gnd cell_6t
Xbit_r73_c92 bl[92] br[92] wl[73] vdd gnd cell_6t
Xbit_r74_c92 bl[92] br[92] wl[74] vdd gnd cell_6t
Xbit_r75_c92 bl[92] br[92] wl[75] vdd gnd cell_6t
Xbit_r76_c92 bl[92] br[92] wl[76] vdd gnd cell_6t
Xbit_r77_c92 bl[92] br[92] wl[77] vdd gnd cell_6t
Xbit_r78_c92 bl[92] br[92] wl[78] vdd gnd cell_6t
Xbit_r79_c92 bl[92] br[92] wl[79] vdd gnd cell_6t
Xbit_r80_c92 bl[92] br[92] wl[80] vdd gnd cell_6t
Xbit_r81_c92 bl[92] br[92] wl[81] vdd gnd cell_6t
Xbit_r82_c92 bl[92] br[92] wl[82] vdd gnd cell_6t
Xbit_r83_c92 bl[92] br[92] wl[83] vdd gnd cell_6t
Xbit_r84_c92 bl[92] br[92] wl[84] vdd gnd cell_6t
Xbit_r85_c92 bl[92] br[92] wl[85] vdd gnd cell_6t
Xbit_r86_c92 bl[92] br[92] wl[86] vdd gnd cell_6t
Xbit_r87_c92 bl[92] br[92] wl[87] vdd gnd cell_6t
Xbit_r88_c92 bl[92] br[92] wl[88] vdd gnd cell_6t
Xbit_r89_c92 bl[92] br[92] wl[89] vdd gnd cell_6t
Xbit_r90_c92 bl[92] br[92] wl[90] vdd gnd cell_6t
Xbit_r91_c92 bl[92] br[92] wl[91] vdd gnd cell_6t
Xbit_r92_c92 bl[92] br[92] wl[92] vdd gnd cell_6t
Xbit_r93_c92 bl[92] br[92] wl[93] vdd gnd cell_6t
Xbit_r94_c92 bl[92] br[92] wl[94] vdd gnd cell_6t
Xbit_r95_c92 bl[92] br[92] wl[95] vdd gnd cell_6t
Xbit_r96_c92 bl[92] br[92] wl[96] vdd gnd cell_6t
Xbit_r97_c92 bl[92] br[92] wl[97] vdd gnd cell_6t
Xbit_r98_c92 bl[92] br[92] wl[98] vdd gnd cell_6t
Xbit_r99_c92 bl[92] br[92] wl[99] vdd gnd cell_6t
Xbit_r100_c92 bl[92] br[92] wl[100] vdd gnd cell_6t
Xbit_r101_c92 bl[92] br[92] wl[101] vdd gnd cell_6t
Xbit_r102_c92 bl[92] br[92] wl[102] vdd gnd cell_6t
Xbit_r103_c92 bl[92] br[92] wl[103] vdd gnd cell_6t
Xbit_r104_c92 bl[92] br[92] wl[104] vdd gnd cell_6t
Xbit_r105_c92 bl[92] br[92] wl[105] vdd gnd cell_6t
Xbit_r106_c92 bl[92] br[92] wl[106] vdd gnd cell_6t
Xbit_r107_c92 bl[92] br[92] wl[107] vdd gnd cell_6t
Xbit_r108_c92 bl[92] br[92] wl[108] vdd gnd cell_6t
Xbit_r109_c92 bl[92] br[92] wl[109] vdd gnd cell_6t
Xbit_r110_c92 bl[92] br[92] wl[110] vdd gnd cell_6t
Xbit_r111_c92 bl[92] br[92] wl[111] vdd gnd cell_6t
Xbit_r112_c92 bl[92] br[92] wl[112] vdd gnd cell_6t
Xbit_r113_c92 bl[92] br[92] wl[113] vdd gnd cell_6t
Xbit_r114_c92 bl[92] br[92] wl[114] vdd gnd cell_6t
Xbit_r115_c92 bl[92] br[92] wl[115] vdd gnd cell_6t
Xbit_r116_c92 bl[92] br[92] wl[116] vdd gnd cell_6t
Xbit_r117_c92 bl[92] br[92] wl[117] vdd gnd cell_6t
Xbit_r118_c92 bl[92] br[92] wl[118] vdd gnd cell_6t
Xbit_r119_c92 bl[92] br[92] wl[119] vdd gnd cell_6t
Xbit_r120_c92 bl[92] br[92] wl[120] vdd gnd cell_6t
Xbit_r121_c92 bl[92] br[92] wl[121] vdd gnd cell_6t
Xbit_r122_c92 bl[92] br[92] wl[122] vdd gnd cell_6t
Xbit_r123_c92 bl[92] br[92] wl[123] vdd gnd cell_6t
Xbit_r124_c92 bl[92] br[92] wl[124] vdd gnd cell_6t
Xbit_r125_c92 bl[92] br[92] wl[125] vdd gnd cell_6t
Xbit_r126_c92 bl[92] br[92] wl[126] vdd gnd cell_6t
Xbit_r127_c92 bl[92] br[92] wl[127] vdd gnd cell_6t
Xbit_r128_c92 bl[92] br[92] wl[128] vdd gnd cell_6t
Xbit_r129_c92 bl[92] br[92] wl[129] vdd gnd cell_6t
Xbit_r130_c92 bl[92] br[92] wl[130] vdd gnd cell_6t
Xbit_r131_c92 bl[92] br[92] wl[131] vdd gnd cell_6t
Xbit_r132_c92 bl[92] br[92] wl[132] vdd gnd cell_6t
Xbit_r133_c92 bl[92] br[92] wl[133] vdd gnd cell_6t
Xbit_r134_c92 bl[92] br[92] wl[134] vdd gnd cell_6t
Xbit_r135_c92 bl[92] br[92] wl[135] vdd gnd cell_6t
Xbit_r136_c92 bl[92] br[92] wl[136] vdd gnd cell_6t
Xbit_r137_c92 bl[92] br[92] wl[137] vdd gnd cell_6t
Xbit_r138_c92 bl[92] br[92] wl[138] vdd gnd cell_6t
Xbit_r139_c92 bl[92] br[92] wl[139] vdd gnd cell_6t
Xbit_r140_c92 bl[92] br[92] wl[140] vdd gnd cell_6t
Xbit_r141_c92 bl[92] br[92] wl[141] vdd gnd cell_6t
Xbit_r142_c92 bl[92] br[92] wl[142] vdd gnd cell_6t
Xbit_r143_c92 bl[92] br[92] wl[143] vdd gnd cell_6t
Xbit_r144_c92 bl[92] br[92] wl[144] vdd gnd cell_6t
Xbit_r145_c92 bl[92] br[92] wl[145] vdd gnd cell_6t
Xbit_r146_c92 bl[92] br[92] wl[146] vdd gnd cell_6t
Xbit_r147_c92 bl[92] br[92] wl[147] vdd gnd cell_6t
Xbit_r148_c92 bl[92] br[92] wl[148] vdd gnd cell_6t
Xbit_r149_c92 bl[92] br[92] wl[149] vdd gnd cell_6t
Xbit_r150_c92 bl[92] br[92] wl[150] vdd gnd cell_6t
Xbit_r151_c92 bl[92] br[92] wl[151] vdd gnd cell_6t
Xbit_r152_c92 bl[92] br[92] wl[152] vdd gnd cell_6t
Xbit_r153_c92 bl[92] br[92] wl[153] vdd gnd cell_6t
Xbit_r154_c92 bl[92] br[92] wl[154] vdd gnd cell_6t
Xbit_r155_c92 bl[92] br[92] wl[155] vdd gnd cell_6t
Xbit_r156_c92 bl[92] br[92] wl[156] vdd gnd cell_6t
Xbit_r157_c92 bl[92] br[92] wl[157] vdd gnd cell_6t
Xbit_r158_c92 bl[92] br[92] wl[158] vdd gnd cell_6t
Xbit_r159_c92 bl[92] br[92] wl[159] vdd gnd cell_6t
Xbit_r160_c92 bl[92] br[92] wl[160] vdd gnd cell_6t
Xbit_r161_c92 bl[92] br[92] wl[161] vdd gnd cell_6t
Xbit_r162_c92 bl[92] br[92] wl[162] vdd gnd cell_6t
Xbit_r163_c92 bl[92] br[92] wl[163] vdd gnd cell_6t
Xbit_r164_c92 bl[92] br[92] wl[164] vdd gnd cell_6t
Xbit_r165_c92 bl[92] br[92] wl[165] vdd gnd cell_6t
Xbit_r166_c92 bl[92] br[92] wl[166] vdd gnd cell_6t
Xbit_r167_c92 bl[92] br[92] wl[167] vdd gnd cell_6t
Xbit_r168_c92 bl[92] br[92] wl[168] vdd gnd cell_6t
Xbit_r169_c92 bl[92] br[92] wl[169] vdd gnd cell_6t
Xbit_r170_c92 bl[92] br[92] wl[170] vdd gnd cell_6t
Xbit_r171_c92 bl[92] br[92] wl[171] vdd gnd cell_6t
Xbit_r172_c92 bl[92] br[92] wl[172] vdd gnd cell_6t
Xbit_r173_c92 bl[92] br[92] wl[173] vdd gnd cell_6t
Xbit_r174_c92 bl[92] br[92] wl[174] vdd gnd cell_6t
Xbit_r175_c92 bl[92] br[92] wl[175] vdd gnd cell_6t
Xbit_r176_c92 bl[92] br[92] wl[176] vdd gnd cell_6t
Xbit_r177_c92 bl[92] br[92] wl[177] vdd gnd cell_6t
Xbit_r178_c92 bl[92] br[92] wl[178] vdd gnd cell_6t
Xbit_r179_c92 bl[92] br[92] wl[179] vdd gnd cell_6t
Xbit_r180_c92 bl[92] br[92] wl[180] vdd gnd cell_6t
Xbit_r181_c92 bl[92] br[92] wl[181] vdd gnd cell_6t
Xbit_r182_c92 bl[92] br[92] wl[182] vdd gnd cell_6t
Xbit_r183_c92 bl[92] br[92] wl[183] vdd gnd cell_6t
Xbit_r184_c92 bl[92] br[92] wl[184] vdd gnd cell_6t
Xbit_r185_c92 bl[92] br[92] wl[185] vdd gnd cell_6t
Xbit_r186_c92 bl[92] br[92] wl[186] vdd gnd cell_6t
Xbit_r187_c92 bl[92] br[92] wl[187] vdd gnd cell_6t
Xbit_r188_c92 bl[92] br[92] wl[188] vdd gnd cell_6t
Xbit_r189_c92 bl[92] br[92] wl[189] vdd gnd cell_6t
Xbit_r190_c92 bl[92] br[92] wl[190] vdd gnd cell_6t
Xbit_r191_c92 bl[92] br[92] wl[191] vdd gnd cell_6t
Xbit_r192_c92 bl[92] br[92] wl[192] vdd gnd cell_6t
Xbit_r193_c92 bl[92] br[92] wl[193] vdd gnd cell_6t
Xbit_r194_c92 bl[92] br[92] wl[194] vdd gnd cell_6t
Xbit_r195_c92 bl[92] br[92] wl[195] vdd gnd cell_6t
Xbit_r196_c92 bl[92] br[92] wl[196] vdd gnd cell_6t
Xbit_r197_c92 bl[92] br[92] wl[197] vdd gnd cell_6t
Xbit_r198_c92 bl[92] br[92] wl[198] vdd gnd cell_6t
Xbit_r199_c92 bl[92] br[92] wl[199] vdd gnd cell_6t
Xbit_r200_c92 bl[92] br[92] wl[200] vdd gnd cell_6t
Xbit_r201_c92 bl[92] br[92] wl[201] vdd gnd cell_6t
Xbit_r202_c92 bl[92] br[92] wl[202] vdd gnd cell_6t
Xbit_r203_c92 bl[92] br[92] wl[203] vdd gnd cell_6t
Xbit_r204_c92 bl[92] br[92] wl[204] vdd gnd cell_6t
Xbit_r205_c92 bl[92] br[92] wl[205] vdd gnd cell_6t
Xbit_r206_c92 bl[92] br[92] wl[206] vdd gnd cell_6t
Xbit_r207_c92 bl[92] br[92] wl[207] vdd gnd cell_6t
Xbit_r208_c92 bl[92] br[92] wl[208] vdd gnd cell_6t
Xbit_r209_c92 bl[92] br[92] wl[209] vdd gnd cell_6t
Xbit_r210_c92 bl[92] br[92] wl[210] vdd gnd cell_6t
Xbit_r211_c92 bl[92] br[92] wl[211] vdd gnd cell_6t
Xbit_r212_c92 bl[92] br[92] wl[212] vdd gnd cell_6t
Xbit_r213_c92 bl[92] br[92] wl[213] vdd gnd cell_6t
Xbit_r214_c92 bl[92] br[92] wl[214] vdd gnd cell_6t
Xbit_r215_c92 bl[92] br[92] wl[215] vdd gnd cell_6t
Xbit_r216_c92 bl[92] br[92] wl[216] vdd gnd cell_6t
Xbit_r217_c92 bl[92] br[92] wl[217] vdd gnd cell_6t
Xbit_r218_c92 bl[92] br[92] wl[218] vdd gnd cell_6t
Xbit_r219_c92 bl[92] br[92] wl[219] vdd gnd cell_6t
Xbit_r220_c92 bl[92] br[92] wl[220] vdd gnd cell_6t
Xbit_r221_c92 bl[92] br[92] wl[221] vdd gnd cell_6t
Xbit_r222_c92 bl[92] br[92] wl[222] vdd gnd cell_6t
Xbit_r223_c92 bl[92] br[92] wl[223] vdd gnd cell_6t
Xbit_r224_c92 bl[92] br[92] wl[224] vdd gnd cell_6t
Xbit_r225_c92 bl[92] br[92] wl[225] vdd gnd cell_6t
Xbit_r226_c92 bl[92] br[92] wl[226] vdd gnd cell_6t
Xbit_r227_c92 bl[92] br[92] wl[227] vdd gnd cell_6t
Xbit_r228_c92 bl[92] br[92] wl[228] vdd gnd cell_6t
Xbit_r229_c92 bl[92] br[92] wl[229] vdd gnd cell_6t
Xbit_r230_c92 bl[92] br[92] wl[230] vdd gnd cell_6t
Xbit_r231_c92 bl[92] br[92] wl[231] vdd gnd cell_6t
Xbit_r232_c92 bl[92] br[92] wl[232] vdd gnd cell_6t
Xbit_r233_c92 bl[92] br[92] wl[233] vdd gnd cell_6t
Xbit_r234_c92 bl[92] br[92] wl[234] vdd gnd cell_6t
Xbit_r235_c92 bl[92] br[92] wl[235] vdd gnd cell_6t
Xbit_r236_c92 bl[92] br[92] wl[236] vdd gnd cell_6t
Xbit_r237_c92 bl[92] br[92] wl[237] vdd gnd cell_6t
Xbit_r238_c92 bl[92] br[92] wl[238] vdd gnd cell_6t
Xbit_r239_c92 bl[92] br[92] wl[239] vdd gnd cell_6t
Xbit_r240_c92 bl[92] br[92] wl[240] vdd gnd cell_6t
Xbit_r241_c92 bl[92] br[92] wl[241] vdd gnd cell_6t
Xbit_r242_c92 bl[92] br[92] wl[242] vdd gnd cell_6t
Xbit_r243_c92 bl[92] br[92] wl[243] vdd gnd cell_6t
Xbit_r244_c92 bl[92] br[92] wl[244] vdd gnd cell_6t
Xbit_r245_c92 bl[92] br[92] wl[245] vdd gnd cell_6t
Xbit_r246_c92 bl[92] br[92] wl[246] vdd gnd cell_6t
Xbit_r247_c92 bl[92] br[92] wl[247] vdd gnd cell_6t
Xbit_r248_c92 bl[92] br[92] wl[248] vdd gnd cell_6t
Xbit_r249_c92 bl[92] br[92] wl[249] vdd gnd cell_6t
Xbit_r250_c92 bl[92] br[92] wl[250] vdd gnd cell_6t
Xbit_r251_c92 bl[92] br[92] wl[251] vdd gnd cell_6t
Xbit_r252_c92 bl[92] br[92] wl[252] vdd gnd cell_6t
Xbit_r253_c92 bl[92] br[92] wl[253] vdd gnd cell_6t
Xbit_r254_c92 bl[92] br[92] wl[254] vdd gnd cell_6t
Xbit_r255_c92 bl[92] br[92] wl[255] vdd gnd cell_6t
Xbit_r0_c93 bl[93] br[93] wl[0] vdd gnd cell_6t
Xbit_r1_c93 bl[93] br[93] wl[1] vdd gnd cell_6t
Xbit_r2_c93 bl[93] br[93] wl[2] vdd gnd cell_6t
Xbit_r3_c93 bl[93] br[93] wl[3] vdd gnd cell_6t
Xbit_r4_c93 bl[93] br[93] wl[4] vdd gnd cell_6t
Xbit_r5_c93 bl[93] br[93] wl[5] vdd gnd cell_6t
Xbit_r6_c93 bl[93] br[93] wl[6] vdd gnd cell_6t
Xbit_r7_c93 bl[93] br[93] wl[7] vdd gnd cell_6t
Xbit_r8_c93 bl[93] br[93] wl[8] vdd gnd cell_6t
Xbit_r9_c93 bl[93] br[93] wl[9] vdd gnd cell_6t
Xbit_r10_c93 bl[93] br[93] wl[10] vdd gnd cell_6t
Xbit_r11_c93 bl[93] br[93] wl[11] vdd gnd cell_6t
Xbit_r12_c93 bl[93] br[93] wl[12] vdd gnd cell_6t
Xbit_r13_c93 bl[93] br[93] wl[13] vdd gnd cell_6t
Xbit_r14_c93 bl[93] br[93] wl[14] vdd gnd cell_6t
Xbit_r15_c93 bl[93] br[93] wl[15] vdd gnd cell_6t
Xbit_r16_c93 bl[93] br[93] wl[16] vdd gnd cell_6t
Xbit_r17_c93 bl[93] br[93] wl[17] vdd gnd cell_6t
Xbit_r18_c93 bl[93] br[93] wl[18] vdd gnd cell_6t
Xbit_r19_c93 bl[93] br[93] wl[19] vdd gnd cell_6t
Xbit_r20_c93 bl[93] br[93] wl[20] vdd gnd cell_6t
Xbit_r21_c93 bl[93] br[93] wl[21] vdd gnd cell_6t
Xbit_r22_c93 bl[93] br[93] wl[22] vdd gnd cell_6t
Xbit_r23_c93 bl[93] br[93] wl[23] vdd gnd cell_6t
Xbit_r24_c93 bl[93] br[93] wl[24] vdd gnd cell_6t
Xbit_r25_c93 bl[93] br[93] wl[25] vdd gnd cell_6t
Xbit_r26_c93 bl[93] br[93] wl[26] vdd gnd cell_6t
Xbit_r27_c93 bl[93] br[93] wl[27] vdd gnd cell_6t
Xbit_r28_c93 bl[93] br[93] wl[28] vdd gnd cell_6t
Xbit_r29_c93 bl[93] br[93] wl[29] vdd gnd cell_6t
Xbit_r30_c93 bl[93] br[93] wl[30] vdd gnd cell_6t
Xbit_r31_c93 bl[93] br[93] wl[31] vdd gnd cell_6t
Xbit_r32_c93 bl[93] br[93] wl[32] vdd gnd cell_6t
Xbit_r33_c93 bl[93] br[93] wl[33] vdd gnd cell_6t
Xbit_r34_c93 bl[93] br[93] wl[34] vdd gnd cell_6t
Xbit_r35_c93 bl[93] br[93] wl[35] vdd gnd cell_6t
Xbit_r36_c93 bl[93] br[93] wl[36] vdd gnd cell_6t
Xbit_r37_c93 bl[93] br[93] wl[37] vdd gnd cell_6t
Xbit_r38_c93 bl[93] br[93] wl[38] vdd gnd cell_6t
Xbit_r39_c93 bl[93] br[93] wl[39] vdd gnd cell_6t
Xbit_r40_c93 bl[93] br[93] wl[40] vdd gnd cell_6t
Xbit_r41_c93 bl[93] br[93] wl[41] vdd gnd cell_6t
Xbit_r42_c93 bl[93] br[93] wl[42] vdd gnd cell_6t
Xbit_r43_c93 bl[93] br[93] wl[43] vdd gnd cell_6t
Xbit_r44_c93 bl[93] br[93] wl[44] vdd gnd cell_6t
Xbit_r45_c93 bl[93] br[93] wl[45] vdd gnd cell_6t
Xbit_r46_c93 bl[93] br[93] wl[46] vdd gnd cell_6t
Xbit_r47_c93 bl[93] br[93] wl[47] vdd gnd cell_6t
Xbit_r48_c93 bl[93] br[93] wl[48] vdd gnd cell_6t
Xbit_r49_c93 bl[93] br[93] wl[49] vdd gnd cell_6t
Xbit_r50_c93 bl[93] br[93] wl[50] vdd gnd cell_6t
Xbit_r51_c93 bl[93] br[93] wl[51] vdd gnd cell_6t
Xbit_r52_c93 bl[93] br[93] wl[52] vdd gnd cell_6t
Xbit_r53_c93 bl[93] br[93] wl[53] vdd gnd cell_6t
Xbit_r54_c93 bl[93] br[93] wl[54] vdd gnd cell_6t
Xbit_r55_c93 bl[93] br[93] wl[55] vdd gnd cell_6t
Xbit_r56_c93 bl[93] br[93] wl[56] vdd gnd cell_6t
Xbit_r57_c93 bl[93] br[93] wl[57] vdd gnd cell_6t
Xbit_r58_c93 bl[93] br[93] wl[58] vdd gnd cell_6t
Xbit_r59_c93 bl[93] br[93] wl[59] vdd gnd cell_6t
Xbit_r60_c93 bl[93] br[93] wl[60] vdd gnd cell_6t
Xbit_r61_c93 bl[93] br[93] wl[61] vdd gnd cell_6t
Xbit_r62_c93 bl[93] br[93] wl[62] vdd gnd cell_6t
Xbit_r63_c93 bl[93] br[93] wl[63] vdd gnd cell_6t
Xbit_r64_c93 bl[93] br[93] wl[64] vdd gnd cell_6t
Xbit_r65_c93 bl[93] br[93] wl[65] vdd gnd cell_6t
Xbit_r66_c93 bl[93] br[93] wl[66] vdd gnd cell_6t
Xbit_r67_c93 bl[93] br[93] wl[67] vdd gnd cell_6t
Xbit_r68_c93 bl[93] br[93] wl[68] vdd gnd cell_6t
Xbit_r69_c93 bl[93] br[93] wl[69] vdd gnd cell_6t
Xbit_r70_c93 bl[93] br[93] wl[70] vdd gnd cell_6t
Xbit_r71_c93 bl[93] br[93] wl[71] vdd gnd cell_6t
Xbit_r72_c93 bl[93] br[93] wl[72] vdd gnd cell_6t
Xbit_r73_c93 bl[93] br[93] wl[73] vdd gnd cell_6t
Xbit_r74_c93 bl[93] br[93] wl[74] vdd gnd cell_6t
Xbit_r75_c93 bl[93] br[93] wl[75] vdd gnd cell_6t
Xbit_r76_c93 bl[93] br[93] wl[76] vdd gnd cell_6t
Xbit_r77_c93 bl[93] br[93] wl[77] vdd gnd cell_6t
Xbit_r78_c93 bl[93] br[93] wl[78] vdd gnd cell_6t
Xbit_r79_c93 bl[93] br[93] wl[79] vdd gnd cell_6t
Xbit_r80_c93 bl[93] br[93] wl[80] vdd gnd cell_6t
Xbit_r81_c93 bl[93] br[93] wl[81] vdd gnd cell_6t
Xbit_r82_c93 bl[93] br[93] wl[82] vdd gnd cell_6t
Xbit_r83_c93 bl[93] br[93] wl[83] vdd gnd cell_6t
Xbit_r84_c93 bl[93] br[93] wl[84] vdd gnd cell_6t
Xbit_r85_c93 bl[93] br[93] wl[85] vdd gnd cell_6t
Xbit_r86_c93 bl[93] br[93] wl[86] vdd gnd cell_6t
Xbit_r87_c93 bl[93] br[93] wl[87] vdd gnd cell_6t
Xbit_r88_c93 bl[93] br[93] wl[88] vdd gnd cell_6t
Xbit_r89_c93 bl[93] br[93] wl[89] vdd gnd cell_6t
Xbit_r90_c93 bl[93] br[93] wl[90] vdd gnd cell_6t
Xbit_r91_c93 bl[93] br[93] wl[91] vdd gnd cell_6t
Xbit_r92_c93 bl[93] br[93] wl[92] vdd gnd cell_6t
Xbit_r93_c93 bl[93] br[93] wl[93] vdd gnd cell_6t
Xbit_r94_c93 bl[93] br[93] wl[94] vdd gnd cell_6t
Xbit_r95_c93 bl[93] br[93] wl[95] vdd gnd cell_6t
Xbit_r96_c93 bl[93] br[93] wl[96] vdd gnd cell_6t
Xbit_r97_c93 bl[93] br[93] wl[97] vdd gnd cell_6t
Xbit_r98_c93 bl[93] br[93] wl[98] vdd gnd cell_6t
Xbit_r99_c93 bl[93] br[93] wl[99] vdd gnd cell_6t
Xbit_r100_c93 bl[93] br[93] wl[100] vdd gnd cell_6t
Xbit_r101_c93 bl[93] br[93] wl[101] vdd gnd cell_6t
Xbit_r102_c93 bl[93] br[93] wl[102] vdd gnd cell_6t
Xbit_r103_c93 bl[93] br[93] wl[103] vdd gnd cell_6t
Xbit_r104_c93 bl[93] br[93] wl[104] vdd gnd cell_6t
Xbit_r105_c93 bl[93] br[93] wl[105] vdd gnd cell_6t
Xbit_r106_c93 bl[93] br[93] wl[106] vdd gnd cell_6t
Xbit_r107_c93 bl[93] br[93] wl[107] vdd gnd cell_6t
Xbit_r108_c93 bl[93] br[93] wl[108] vdd gnd cell_6t
Xbit_r109_c93 bl[93] br[93] wl[109] vdd gnd cell_6t
Xbit_r110_c93 bl[93] br[93] wl[110] vdd gnd cell_6t
Xbit_r111_c93 bl[93] br[93] wl[111] vdd gnd cell_6t
Xbit_r112_c93 bl[93] br[93] wl[112] vdd gnd cell_6t
Xbit_r113_c93 bl[93] br[93] wl[113] vdd gnd cell_6t
Xbit_r114_c93 bl[93] br[93] wl[114] vdd gnd cell_6t
Xbit_r115_c93 bl[93] br[93] wl[115] vdd gnd cell_6t
Xbit_r116_c93 bl[93] br[93] wl[116] vdd gnd cell_6t
Xbit_r117_c93 bl[93] br[93] wl[117] vdd gnd cell_6t
Xbit_r118_c93 bl[93] br[93] wl[118] vdd gnd cell_6t
Xbit_r119_c93 bl[93] br[93] wl[119] vdd gnd cell_6t
Xbit_r120_c93 bl[93] br[93] wl[120] vdd gnd cell_6t
Xbit_r121_c93 bl[93] br[93] wl[121] vdd gnd cell_6t
Xbit_r122_c93 bl[93] br[93] wl[122] vdd gnd cell_6t
Xbit_r123_c93 bl[93] br[93] wl[123] vdd gnd cell_6t
Xbit_r124_c93 bl[93] br[93] wl[124] vdd gnd cell_6t
Xbit_r125_c93 bl[93] br[93] wl[125] vdd gnd cell_6t
Xbit_r126_c93 bl[93] br[93] wl[126] vdd gnd cell_6t
Xbit_r127_c93 bl[93] br[93] wl[127] vdd gnd cell_6t
Xbit_r128_c93 bl[93] br[93] wl[128] vdd gnd cell_6t
Xbit_r129_c93 bl[93] br[93] wl[129] vdd gnd cell_6t
Xbit_r130_c93 bl[93] br[93] wl[130] vdd gnd cell_6t
Xbit_r131_c93 bl[93] br[93] wl[131] vdd gnd cell_6t
Xbit_r132_c93 bl[93] br[93] wl[132] vdd gnd cell_6t
Xbit_r133_c93 bl[93] br[93] wl[133] vdd gnd cell_6t
Xbit_r134_c93 bl[93] br[93] wl[134] vdd gnd cell_6t
Xbit_r135_c93 bl[93] br[93] wl[135] vdd gnd cell_6t
Xbit_r136_c93 bl[93] br[93] wl[136] vdd gnd cell_6t
Xbit_r137_c93 bl[93] br[93] wl[137] vdd gnd cell_6t
Xbit_r138_c93 bl[93] br[93] wl[138] vdd gnd cell_6t
Xbit_r139_c93 bl[93] br[93] wl[139] vdd gnd cell_6t
Xbit_r140_c93 bl[93] br[93] wl[140] vdd gnd cell_6t
Xbit_r141_c93 bl[93] br[93] wl[141] vdd gnd cell_6t
Xbit_r142_c93 bl[93] br[93] wl[142] vdd gnd cell_6t
Xbit_r143_c93 bl[93] br[93] wl[143] vdd gnd cell_6t
Xbit_r144_c93 bl[93] br[93] wl[144] vdd gnd cell_6t
Xbit_r145_c93 bl[93] br[93] wl[145] vdd gnd cell_6t
Xbit_r146_c93 bl[93] br[93] wl[146] vdd gnd cell_6t
Xbit_r147_c93 bl[93] br[93] wl[147] vdd gnd cell_6t
Xbit_r148_c93 bl[93] br[93] wl[148] vdd gnd cell_6t
Xbit_r149_c93 bl[93] br[93] wl[149] vdd gnd cell_6t
Xbit_r150_c93 bl[93] br[93] wl[150] vdd gnd cell_6t
Xbit_r151_c93 bl[93] br[93] wl[151] vdd gnd cell_6t
Xbit_r152_c93 bl[93] br[93] wl[152] vdd gnd cell_6t
Xbit_r153_c93 bl[93] br[93] wl[153] vdd gnd cell_6t
Xbit_r154_c93 bl[93] br[93] wl[154] vdd gnd cell_6t
Xbit_r155_c93 bl[93] br[93] wl[155] vdd gnd cell_6t
Xbit_r156_c93 bl[93] br[93] wl[156] vdd gnd cell_6t
Xbit_r157_c93 bl[93] br[93] wl[157] vdd gnd cell_6t
Xbit_r158_c93 bl[93] br[93] wl[158] vdd gnd cell_6t
Xbit_r159_c93 bl[93] br[93] wl[159] vdd gnd cell_6t
Xbit_r160_c93 bl[93] br[93] wl[160] vdd gnd cell_6t
Xbit_r161_c93 bl[93] br[93] wl[161] vdd gnd cell_6t
Xbit_r162_c93 bl[93] br[93] wl[162] vdd gnd cell_6t
Xbit_r163_c93 bl[93] br[93] wl[163] vdd gnd cell_6t
Xbit_r164_c93 bl[93] br[93] wl[164] vdd gnd cell_6t
Xbit_r165_c93 bl[93] br[93] wl[165] vdd gnd cell_6t
Xbit_r166_c93 bl[93] br[93] wl[166] vdd gnd cell_6t
Xbit_r167_c93 bl[93] br[93] wl[167] vdd gnd cell_6t
Xbit_r168_c93 bl[93] br[93] wl[168] vdd gnd cell_6t
Xbit_r169_c93 bl[93] br[93] wl[169] vdd gnd cell_6t
Xbit_r170_c93 bl[93] br[93] wl[170] vdd gnd cell_6t
Xbit_r171_c93 bl[93] br[93] wl[171] vdd gnd cell_6t
Xbit_r172_c93 bl[93] br[93] wl[172] vdd gnd cell_6t
Xbit_r173_c93 bl[93] br[93] wl[173] vdd gnd cell_6t
Xbit_r174_c93 bl[93] br[93] wl[174] vdd gnd cell_6t
Xbit_r175_c93 bl[93] br[93] wl[175] vdd gnd cell_6t
Xbit_r176_c93 bl[93] br[93] wl[176] vdd gnd cell_6t
Xbit_r177_c93 bl[93] br[93] wl[177] vdd gnd cell_6t
Xbit_r178_c93 bl[93] br[93] wl[178] vdd gnd cell_6t
Xbit_r179_c93 bl[93] br[93] wl[179] vdd gnd cell_6t
Xbit_r180_c93 bl[93] br[93] wl[180] vdd gnd cell_6t
Xbit_r181_c93 bl[93] br[93] wl[181] vdd gnd cell_6t
Xbit_r182_c93 bl[93] br[93] wl[182] vdd gnd cell_6t
Xbit_r183_c93 bl[93] br[93] wl[183] vdd gnd cell_6t
Xbit_r184_c93 bl[93] br[93] wl[184] vdd gnd cell_6t
Xbit_r185_c93 bl[93] br[93] wl[185] vdd gnd cell_6t
Xbit_r186_c93 bl[93] br[93] wl[186] vdd gnd cell_6t
Xbit_r187_c93 bl[93] br[93] wl[187] vdd gnd cell_6t
Xbit_r188_c93 bl[93] br[93] wl[188] vdd gnd cell_6t
Xbit_r189_c93 bl[93] br[93] wl[189] vdd gnd cell_6t
Xbit_r190_c93 bl[93] br[93] wl[190] vdd gnd cell_6t
Xbit_r191_c93 bl[93] br[93] wl[191] vdd gnd cell_6t
Xbit_r192_c93 bl[93] br[93] wl[192] vdd gnd cell_6t
Xbit_r193_c93 bl[93] br[93] wl[193] vdd gnd cell_6t
Xbit_r194_c93 bl[93] br[93] wl[194] vdd gnd cell_6t
Xbit_r195_c93 bl[93] br[93] wl[195] vdd gnd cell_6t
Xbit_r196_c93 bl[93] br[93] wl[196] vdd gnd cell_6t
Xbit_r197_c93 bl[93] br[93] wl[197] vdd gnd cell_6t
Xbit_r198_c93 bl[93] br[93] wl[198] vdd gnd cell_6t
Xbit_r199_c93 bl[93] br[93] wl[199] vdd gnd cell_6t
Xbit_r200_c93 bl[93] br[93] wl[200] vdd gnd cell_6t
Xbit_r201_c93 bl[93] br[93] wl[201] vdd gnd cell_6t
Xbit_r202_c93 bl[93] br[93] wl[202] vdd gnd cell_6t
Xbit_r203_c93 bl[93] br[93] wl[203] vdd gnd cell_6t
Xbit_r204_c93 bl[93] br[93] wl[204] vdd gnd cell_6t
Xbit_r205_c93 bl[93] br[93] wl[205] vdd gnd cell_6t
Xbit_r206_c93 bl[93] br[93] wl[206] vdd gnd cell_6t
Xbit_r207_c93 bl[93] br[93] wl[207] vdd gnd cell_6t
Xbit_r208_c93 bl[93] br[93] wl[208] vdd gnd cell_6t
Xbit_r209_c93 bl[93] br[93] wl[209] vdd gnd cell_6t
Xbit_r210_c93 bl[93] br[93] wl[210] vdd gnd cell_6t
Xbit_r211_c93 bl[93] br[93] wl[211] vdd gnd cell_6t
Xbit_r212_c93 bl[93] br[93] wl[212] vdd gnd cell_6t
Xbit_r213_c93 bl[93] br[93] wl[213] vdd gnd cell_6t
Xbit_r214_c93 bl[93] br[93] wl[214] vdd gnd cell_6t
Xbit_r215_c93 bl[93] br[93] wl[215] vdd gnd cell_6t
Xbit_r216_c93 bl[93] br[93] wl[216] vdd gnd cell_6t
Xbit_r217_c93 bl[93] br[93] wl[217] vdd gnd cell_6t
Xbit_r218_c93 bl[93] br[93] wl[218] vdd gnd cell_6t
Xbit_r219_c93 bl[93] br[93] wl[219] vdd gnd cell_6t
Xbit_r220_c93 bl[93] br[93] wl[220] vdd gnd cell_6t
Xbit_r221_c93 bl[93] br[93] wl[221] vdd gnd cell_6t
Xbit_r222_c93 bl[93] br[93] wl[222] vdd gnd cell_6t
Xbit_r223_c93 bl[93] br[93] wl[223] vdd gnd cell_6t
Xbit_r224_c93 bl[93] br[93] wl[224] vdd gnd cell_6t
Xbit_r225_c93 bl[93] br[93] wl[225] vdd gnd cell_6t
Xbit_r226_c93 bl[93] br[93] wl[226] vdd gnd cell_6t
Xbit_r227_c93 bl[93] br[93] wl[227] vdd gnd cell_6t
Xbit_r228_c93 bl[93] br[93] wl[228] vdd gnd cell_6t
Xbit_r229_c93 bl[93] br[93] wl[229] vdd gnd cell_6t
Xbit_r230_c93 bl[93] br[93] wl[230] vdd gnd cell_6t
Xbit_r231_c93 bl[93] br[93] wl[231] vdd gnd cell_6t
Xbit_r232_c93 bl[93] br[93] wl[232] vdd gnd cell_6t
Xbit_r233_c93 bl[93] br[93] wl[233] vdd gnd cell_6t
Xbit_r234_c93 bl[93] br[93] wl[234] vdd gnd cell_6t
Xbit_r235_c93 bl[93] br[93] wl[235] vdd gnd cell_6t
Xbit_r236_c93 bl[93] br[93] wl[236] vdd gnd cell_6t
Xbit_r237_c93 bl[93] br[93] wl[237] vdd gnd cell_6t
Xbit_r238_c93 bl[93] br[93] wl[238] vdd gnd cell_6t
Xbit_r239_c93 bl[93] br[93] wl[239] vdd gnd cell_6t
Xbit_r240_c93 bl[93] br[93] wl[240] vdd gnd cell_6t
Xbit_r241_c93 bl[93] br[93] wl[241] vdd gnd cell_6t
Xbit_r242_c93 bl[93] br[93] wl[242] vdd gnd cell_6t
Xbit_r243_c93 bl[93] br[93] wl[243] vdd gnd cell_6t
Xbit_r244_c93 bl[93] br[93] wl[244] vdd gnd cell_6t
Xbit_r245_c93 bl[93] br[93] wl[245] vdd gnd cell_6t
Xbit_r246_c93 bl[93] br[93] wl[246] vdd gnd cell_6t
Xbit_r247_c93 bl[93] br[93] wl[247] vdd gnd cell_6t
Xbit_r248_c93 bl[93] br[93] wl[248] vdd gnd cell_6t
Xbit_r249_c93 bl[93] br[93] wl[249] vdd gnd cell_6t
Xbit_r250_c93 bl[93] br[93] wl[250] vdd gnd cell_6t
Xbit_r251_c93 bl[93] br[93] wl[251] vdd gnd cell_6t
Xbit_r252_c93 bl[93] br[93] wl[252] vdd gnd cell_6t
Xbit_r253_c93 bl[93] br[93] wl[253] vdd gnd cell_6t
Xbit_r254_c93 bl[93] br[93] wl[254] vdd gnd cell_6t
Xbit_r255_c93 bl[93] br[93] wl[255] vdd gnd cell_6t
Xbit_r0_c94 bl[94] br[94] wl[0] vdd gnd cell_6t
Xbit_r1_c94 bl[94] br[94] wl[1] vdd gnd cell_6t
Xbit_r2_c94 bl[94] br[94] wl[2] vdd gnd cell_6t
Xbit_r3_c94 bl[94] br[94] wl[3] vdd gnd cell_6t
Xbit_r4_c94 bl[94] br[94] wl[4] vdd gnd cell_6t
Xbit_r5_c94 bl[94] br[94] wl[5] vdd gnd cell_6t
Xbit_r6_c94 bl[94] br[94] wl[6] vdd gnd cell_6t
Xbit_r7_c94 bl[94] br[94] wl[7] vdd gnd cell_6t
Xbit_r8_c94 bl[94] br[94] wl[8] vdd gnd cell_6t
Xbit_r9_c94 bl[94] br[94] wl[9] vdd gnd cell_6t
Xbit_r10_c94 bl[94] br[94] wl[10] vdd gnd cell_6t
Xbit_r11_c94 bl[94] br[94] wl[11] vdd gnd cell_6t
Xbit_r12_c94 bl[94] br[94] wl[12] vdd gnd cell_6t
Xbit_r13_c94 bl[94] br[94] wl[13] vdd gnd cell_6t
Xbit_r14_c94 bl[94] br[94] wl[14] vdd gnd cell_6t
Xbit_r15_c94 bl[94] br[94] wl[15] vdd gnd cell_6t
Xbit_r16_c94 bl[94] br[94] wl[16] vdd gnd cell_6t
Xbit_r17_c94 bl[94] br[94] wl[17] vdd gnd cell_6t
Xbit_r18_c94 bl[94] br[94] wl[18] vdd gnd cell_6t
Xbit_r19_c94 bl[94] br[94] wl[19] vdd gnd cell_6t
Xbit_r20_c94 bl[94] br[94] wl[20] vdd gnd cell_6t
Xbit_r21_c94 bl[94] br[94] wl[21] vdd gnd cell_6t
Xbit_r22_c94 bl[94] br[94] wl[22] vdd gnd cell_6t
Xbit_r23_c94 bl[94] br[94] wl[23] vdd gnd cell_6t
Xbit_r24_c94 bl[94] br[94] wl[24] vdd gnd cell_6t
Xbit_r25_c94 bl[94] br[94] wl[25] vdd gnd cell_6t
Xbit_r26_c94 bl[94] br[94] wl[26] vdd gnd cell_6t
Xbit_r27_c94 bl[94] br[94] wl[27] vdd gnd cell_6t
Xbit_r28_c94 bl[94] br[94] wl[28] vdd gnd cell_6t
Xbit_r29_c94 bl[94] br[94] wl[29] vdd gnd cell_6t
Xbit_r30_c94 bl[94] br[94] wl[30] vdd gnd cell_6t
Xbit_r31_c94 bl[94] br[94] wl[31] vdd gnd cell_6t
Xbit_r32_c94 bl[94] br[94] wl[32] vdd gnd cell_6t
Xbit_r33_c94 bl[94] br[94] wl[33] vdd gnd cell_6t
Xbit_r34_c94 bl[94] br[94] wl[34] vdd gnd cell_6t
Xbit_r35_c94 bl[94] br[94] wl[35] vdd gnd cell_6t
Xbit_r36_c94 bl[94] br[94] wl[36] vdd gnd cell_6t
Xbit_r37_c94 bl[94] br[94] wl[37] vdd gnd cell_6t
Xbit_r38_c94 bl[94] br[94] wl[38] vdd gnd cell_6t
Xbit_r39_c94 bl[94] br[94] wl[39] vdd gnd cell_6t
Xbit_r40_c94 bl[94] br[94] wl[40] vdd gnd cell_6t
Xbit_r41_c94 bl[94] br[94] wl[41] vdd gnd cell_6t
Xbit_r42_c94 bl[94] br[94] wl[42] vdd gnd cell_6t
Xbit_r43_c94 bl[94] br[94] wl[43] vdd gnd cell_6t
Xbit_r44_c94 bl[94] br[94] wl[44] vdd gnd cell_6t
Xbit_r45_c94 bl[94] br[94] wl[45] vdd gnd cell_6t
Xbit_r46_c94 bl[94] br[94] wl[46] vdd gnd cell_6t
Xbit_r47_c94 bl[94] br[94] wl[47] vdd gnd cell_6t
Xbit_r48_c94 bl[94] br[94] wl[48] vdd gnd cell_6t
Xbit_r49_c94 bl[94] br[94] wl[49] vdd gnd cell_6t
Xbit_r50_c94 bl[94] br[94] wl[50] vdd gnd cell_6t
Xbit_r51_c94 bl[94] br[94] wl[51] vdd gnd cell_6t
Xbit_r52_c94 bl[94] br[94] wl[52] vdd gnd cell_6t
Xbit_r53_c94 bl[94] br[94] wl[53] vdd gnd cell_6t
Xbit_r54_c94 bl[94] br[94] wl[54] vdd gnd cell_6t
Xbit_r55_c94 bl[94] br[94] wl[55] vdd gnd cell_6t
Xbit_r56_c94 bl[94] br[94] wl[56] vdd gnd cell_6t
Xbit_r57_c94 bl[94] br[94] wl[57] vdd gnd cell_6t
Xbit_r58_c94 bl[94] br[94] wl[58] vdd gnd cell_6t
Xbit_r59_c94 bl[94] br[94] wl[59] vdd gnd cell_6t
Xbit_r60_c94 bl[94] br[94] wl[60] vdd gnd cell_6t
Xbit_r61_c94 bl[94] br[94] wl[61] vdd gnd cell_6t
Xbit_r62_c94 bl[94] br[94] wl[62] vdd gnd cell_6t
Xbit_r63_c94 bl[94] br[94] wl[63] vdd gnd cell_6t
Xbit_r64_c94 bl[94] br[94] wl[64] vdd gnd cell_6t
Xbit_r65_c94 bl[94] br[94] wl[65] vdd gnd cell_6t
Xbit_r66_c94 bl[94] br[94] wl[66] vdd gnd cell_6t
Xbit_r67_c94 bl[94] br[94] wl[67] vdd gnd cell_6t
Xbit_r68_c94 bl[94] br[94] wl[68] vdd gnd cell_6t
Xbit_r69_c94 bl[94] br[94] wl[69] vdd gnd cell_6t
Xbit_r70_c94 bl[94] br[94] wl[70] vdd gnd cell_6t
Xbit_r71_c94 bl[94] br[94] wl[71] vdd gnd cell_6t
Xbit_r72_c94 bl[94] br[94] wl[72] vdd gnd cell_6t
Xbit_r73_c94 bl[94] br[94] wl[73] vdd gnd cell_6t
Xbit_r74_c94 bl[94] br[94] wl[74] vdd gnd cell_6t
Xbit_r75_c94 bl[94] br[94] wl[75] vdd gnd cell_6t
Xbit_r76_c94 bl[94] br[94] wl[76] vdd gnd cell_6t
Xbit_r77_c94 bl[94] br[94] wl[77] vdd gnd cell_6t
Xbit_r78_c94 bl[94] br[94] wl[78] vdd gnd cell_6t
Xbit_r79_c94 bl[94] br[94] wl[79] vdd gnd cell_6t
Xbit_r80_c94 bl[94] br[94] wl[80] vdd gnd cell_6t
Xbit_r81_c94 bl[94] br[94] wl[81] vdd gnd cell_6t
Xbit_r82_c94 bl[94] br[94] wl[82] vdd gnd cell_6t
Xbit_r83_c94 bl[94] br[94] wl[83] vdd gnd cell_6t
Xbit_r84_c94 bl[94] br[94] wl[84] vdd gnd cell_6t
Xbit_r85_c94 bl[94] br[94] wl[85] vdd gnd cell_6t
Xbit_r86_c94 bl[94] br[94] wl[86] vdd gnd cell_6t
Xbit_r87_c94 bl[94] br[94] wl[87] vdd gnd cell_6t
Xbit_r88_c94 bl[94] br[94] wl[88] vdd gnd cell_6t
Xbit_r89_c94 bl[94] br[94] wl[89] vdd gnd cell_6t
Xbit_r90_c94 bl[94] br[94] wl[90] vdd gnd cell_6t
Xbit_r91_c94 bl[94] br[94] wl[91] vdd gnd cell_6t
Xbit_r92_c94 bl[94] br[94] wl[92] vdd gnd cell_6t
Xbit_r93_c94 bl[94] br[94] wl[93] vdd gnd cell_6t
Xbit_r94_c94 bl[94] br[94] wl[94] vdd gnd cell_6t
Xbit_r95_c94 bl[94] br[94] wl[95] vdd gnd cell_6t
Xbit_r96_c94 bl[94] br[94] wl[96] vdd gnd cell_6t
Xbit_r97_c94 bl[94] br[94] wl[97] vdd gnd cell_6t
Xbit_r98_c94 bl[94] br[94] wl[98] vdd gnd cell_6t
Xbit_r99_c94 bl[94] br[94] wl[99] vdd gnd cell_6t
Xbit_r100_c94 bl[94] br[94] wl[100] vdd gnd cell_6t
Xbit_r101_c94 bl[94] br[94] wl[101] vdd gnd cell_6t
Xbit_r102_c94 bl[94] br[94] wl[102] vdd gnd cell_6t
Xbit_r103_c94 bl[94] br[94] wl[103] vdd gnd cell_6t
Xbit_r104_c94 bl[94] br[94] wl[104] vdd gnd cell_6t
Xbit_r105_c94 bl[94] br[94] wl[105] vdd gnd cell_6t
Xbit_r106_c94 bl[94] br[94] wl[106] vdd gnd cell_6t
Xbit_r107_c94 bl[94] br[94] wl[107] vdd gnd cell_6t
Xbit_r108_c94 bl[94] br[94] wl[108] vdd gnd cell_6t
Xbit_r109_c94 bl[94] br[94] wl[109] vdd gnd cell_6t
Xbit_r110_c94 bl[94] br[94] wl[110] vdd gnd cell_6t
Xbit_r111_c94 bl[94] br[94] wl[111] vdd gnd cell_6t
Xbit_r112_c94 bl[94] br[94] wl[112] vdd gnd cell_6t
Xbit_r113_c94 bl[94] br[94] wl[113] vdd gnd cell_6t
Xbit_r114_c94 bl[94] br[94] wl[114] vdd gnd cell_6t
Xbit_r115_c94 bl[94] br[94] wl[115] vdd gnd cell_6t
Xbit_r116_c94 bl[94] br[94] wl[116] vdd gnd cell_6t
Xbit_r117_c94 bl[94] br[94] wl[117] vdd gnd cell_6t
Xbit_r118_c94 bl[94] br[94] wl[118] vdd gnd cell_6t
Xbit_r119_c94 bl[94] br[94] wl[119] vdd gnd cell_6t
Xbit_r120_c94 bl[94] br[94] wl[120] vdd gnd cell_6t
Xbit_r121_c94 bl[94] br[94] wl[121] vdd gnd cell_6t
Xbit_r122_c94 bl[94] br[94] wl[122] vdd gnd cell_6t
Xbit_r123_c94 bl[94] br[94] wl[123] vdd gnd cell_6t
Xbit_r124_c94 bl[94] br[94] wl[124] vdd gnd cell_6t
Xbit_r125_c94 bl[94] br[94] wl[125] vdd gnd cell_6t
Xbit_r126_c94 bl[94] br[94] wl[126] vdd gnd cell_6t
Xbit_r127_c94 bl[94] br[94] wl[127] vdd gnd cell_6t
Xbit_r128_c94 bl[94] br[94] wl[128] vdd gnd cell_6t
Xbit_r129_c94 bl[94] br[94] wl[129] vdd gnd cell_6t
Xbit_r130_c94 bl[94] br[94] wl[130] vdd gnd cell_6t
Xbit_r131_c94 bl[94] br[94] wl[131] vdd gnd cell_6t
Xbit_r132_c94 bl[94] br[94] wl[132] vdd gnd cell_6t
Xbit_r133_c94 bl[94] br[94] wl[133] vdd gnd cell_6t
Xbit_r134_c94 bl[94] br[94] wl[134] vdd gnd cell_6t
Xbit_r135_c94 bl[94] br[94] wl[135] vdd gnd cell_6t
Xbit_r136_c94 bl[94] br[94] wl[136] vdd gnd cell_6t
Xbit_r137_c94 bl[94] br[94] wl[137] vdd gnd cell_6t
Xbit_r138_c94 bl[94] br[94] wl[138] vdd gnd cell_6t
Xbit_r139_c94 bl[94] br[94] wl[139] vdd gnd cell_6t
Xbit_r140_c94 bl[94] br[94] wl[140] vdd gnd cell_6t
Xbit_r141_c94 bl[94] br[94] wl[141] vdd gnd cell_6t
Xbit_r142_c94 bl[94] br[94] wl[142] vdd gnd cell_6t
Xbit_r143_c94 bl[94] br[94] wl[143] vdd gnd cell_6t
Xbit_r144_c94 bl[94] br[94] wl[144] vdd gnd cell_6t
Xbit_r145_c94 bl[94] br[94] wl[145] vdd gnd cell_6t
Xbit_r146_c94 bl[94] br[94] wl[146] vdd gnd cell_6t
Xbit_r147_c94 bl[94] br[94] wl[147] vdd gnd cell_6t
Xbit_r148_c94 bl[94] br[94] wl[148] vdd gnd cell_6t
Xbit_r149_c94 bl[94] br[94] wl[149] vdd gnd cell_6t
Xbit_r150_c94 bl[94] br[94] wl[150] vdd gnd cell_6t
Xbit_r151_c94 bl[94] br[94] wl[151] vdd gnd cell_6t
Xbit_r152_c94 bl[94] br[94] wl[152] vdd gnd cell_6t
Xbit_r153_c94 bl[94] br[94] wl[153] vdd gnd cell_6t
Xbit_r154_c94 bl[94] br[94] wl[154] vdd gnd cell_6t
Xbit_r155_c94 bl[94] br[94] wl[155] vdd gnd cell_6t
Xbit_r156_c94 bl[94] br[94] wl[156] vdd gnd cell_6t
Xbit_r157_c94 bl[94] br[94] wl[157] vdd gnd cell_6t
Xbit_r158_c94 bl[94] br[94] wl[158] vdd gnd cell_6t
Xbit_r159_c94 bl[94] br[94] wl[159] vdd gnd cell_6t
Xbit_r160_c94 bl[94] br[94] wl[160] vdd gnd cell_6t
Xbit_r161_c94 bl[94] br[94] wl[161] vdd gnd cell_6t
Xbit_r162_c94 bl[94] br[94] wl[162] vdd gnd cell_6t
Xbit_r163_c94 bl[94] br[94] wl[163] vdd gnd cell_6t
Xbit_r164_c94 bl[94] br[94] wl[164] vdd gnd cell_6t
Xbit_r165_c94 bl[94] br[94] wl[165] vdd gnd cell_6t
Xbit_r166_c94 bl[94] br[94] wl[166] vdd gnd cell_6t
Xbit_r167_c94 bl[94] br[94] wl[167] vdd gnd cell_6t
Xbit_r168_c94 bl[94] br[94] wl[168] vdd gnd cell_6t
Xbit_r169_c94 bl[94] br[94] wl[169] vdd gnd cell_6t
Xbit_r170_c94 bl[94] br[94] wl[170] vdd gnd cell_6t
Xbit_r171_c94 bl[94] br[94] wl[171] vdd gnd cell_6t
Xbit_r172_c94 bl[94] br[94] wl[172] vdd gnd cell_6t
Xbit_r173_c94 bl[94] br[94] wl[173] vdd gnd cell_6t
Xbit_r174_c94 bl[94] br[94] wl[174] vdd gnd cell_6t
Xbit_r175_c94 bl[94] br[94] wl[175] vdd gnd cell_6t
Xbit_r176_c94 bl[94] br[94] wl[176] vdd gnd cell_6t
Xbit_r177_c94 bl[94] br[94] wl[177] vdd gnd cell_6t
Xbit_r178_c94 bl[94] br[94] wl[178] vdd gnd cell_6t
Xbit_r179_c94 bl[94] br[94] wl[179] vdd gnd cell_6t
Xbit_r180_c94 bl[94] br[94] wl[180] vdd gnd cell_6t
Xbit_r181_c94 bl[94] br[94] wl[181] vdd gnd cell_6t
Xbit_r182_c94 bl[94] br[94] wl[182] vdd gnd cell_6t
Xbit_r183_c94 bl[94] br[94] wl[183] vdd gnd cell_6t
Xbit_r184_c94 bl[94] br[94] wl[184] vdd gnd cell_6t
Xbit_r185_c94 bl[94] br[94] wl[185] vdd gnd cell_6t
Xbit_r186_c94 bl[94] br[94] wl[186] vdd gnd cell_6t
Xbit_r187_c94 bl[94] br[94] wl[187] vdd gnd cell_6t
Xbit_r188_c94 bl[94] br[94] wl[188] vdd gnd cell_6t
Xbit_r189_c94 bl[94] br[94] wl[189] vdd gnd cell_6t
Xbit_r190_c94 bl[94] br[94] wl[190] vdd gnd cell_6t
Xbit_r191_c94 bl[94] br[94] wl[191] vdd gnd cell_6t
Xbit_r192_c94 bl[94] br[94] wl[192] vdd gnd cell_6t
Xbit_r193_c94 bl[94] br[94] wl[193] vdd gnd cell_6t
Xbit_r194_c94 bl[94] br[94] wl[194] vdd gnd cell_6t
Xbit_r195_c94 bl[94] br[94] wl[195] vdd gnd cell_6t
Xbit_r196_c94 bl[94] br[94] wl[196] vdd gnd cell_6t
Xbit_r197_c94 bl[94] br[94] wl[197] vdd gnd cell_6t
Xbit_r198_c94 bl[94] br[94] wl[198] vdd gnd cell_6t
Xbit_r199_c94 bl[94] br[94] wl[199] vdd gnd cell_6t
Xbit_r200_c94 bl[94] br[94] wl[200] vdd gnd cell_6t
Xbit_r201_c94 bl[94] br[94] wl[201] vdd gnd cell_6t
Xbit_r202_c94 bl[94] br[94] wl[202] vdd gnd cell_6t
Xbit_r203_c94 bl[94] br[94] wl[203] vdd gnd cell_6t
Xbit_r204_c94 bl[94] br[94] wl[204] vdd gnd cell_6t
Xbit_r205_c94 bl[94] br[94] wl[205] vdd gnd cell_6t
Xbit_r206_c94 bl[94] br[94] wl[206] vdd gnd cell_6t
Xbit_r207_c94 bl[94] br[94] wl[207] vdd gnd cell_6t
Xbit_r208_c94 bl[94] br[94] wl[208] vdd gnd cell_6t
Xbit_r209_c94 bl[94] br[94] wl[209] vdd gnd cell_6t
Xbit_r210_c94 bl[94] br[94] wl[210] vdd gnd cell_6t
Xbit_r211_c94 bl[94] br[94] wl[211] vdd gnd cell_6t
Xbit_r212_c94 bl[94] br[94] wl[212] vdd gnd cell_6t
Xbit_r213_c94 bl[94] br[94] wl[213] vdd gnd cell_6t
Xbit_r214_c94 bl[94] br[94] wl[214] vdd gnd cell_6t
Xbit_r215_c94 bl[94] br[94] wl[215] vdd gnd cell_6t
Xbit_r216_c94 bl[94] br[94] wl[216] vdd gnd cell_6t
Xbit_r217_c94 bl[94] br[94] wl[217] vdd gnd cell_6t
Xbit_r218_c94 bl[94] br[94] wl[218] vdd gnd cell_6t
Xbit_r219_c94 bl[94] br[94] wl[219] vdd gnd cell_6t
Xbit_r220_c94 bl[94] br[94] wl[220] vdd gnd cell_6t
Xbit_r221_c94 bl[94] br[94] wl[221] vdd gnd cell_6t
Xbit_r222_c94 bl[94] br[94] wl[222] vdd gnd cell_6t
Xbit_r223_c94 bl[94] br[94] wl[223] vdd gnd cell_6t
Xbit_r224_c94 bl[94] br[94] wl[224] vdd gnd cell_6t
Xbit_r225_c94 bl[94] br[94] wl[225] vdd gnd cell_6t
Xbit_r226_c94 bl[94] br[94] wl[226] vdd gnd cell_6t
Xbit_r227_c94 bl[94] br[94] wl[227] vdd gnd cell_6t
Xbit_r228_c94 bl[94] br[94] wl[228] vdd gnd cell_6t
Xbit_r229_c94 bl[94] br[94] wl[229] vdd gnd cell_6t
Xbit_r230_c94 bl[94] br[94] wl[230] vdd gnd cell_6t
Xbit_r231_c94 bl[94] br[94] wl[231] vdd gnd cell_6t
Xbit_r232_c94 bl[94] br[94] wl[232] vdd gnd cell_6t
Xbit_r233_c94 bl[94] br[94] wl[233] vdd gnd cell_6t
Xbit_r234_c94 bl[94] br[94] wl[234] vdd gnd cell_6t
Xbit_r235_c94 bl[94] br[94] wl[235] vdd gnd cell_6t
Xbit_r236_c94 bl[94] br[94] wl[236] vdd gnd cell_6t
Xbit_r237_c94 bl[94] br[94] wl[237] vdd gnd cell_6t
Xbit_r238_c94 bl[94] br[94] wl[238] vdd gnd cell_6t
Xbit_r239_c94 bl[94] br[94] wl[239] vdd gnd cell_6t
Xbit_r240_c94 bl[94] br[94] wl[240] vdd gnd cell_6t
Xbit_r241_c94 bl[94] br[94] wl[241] vdd gnd cell_6t
Xbit_r242_c94 bl[94] br[94] wl[242] vdd gnd cell_6t
Xbit_r243_c94 bl[94] br[94] wl[243] vdd gnd cell_6t
Xbit_r244_c94 bl[94] br[94] wl[244] vdd gnd cell_6t
Xbit_r245_c94 bl[94] br[94] wl[245] vdd gnd cell_6t
Xbit_r246_c94 bl[94] br[94] wl[246] vdd gnd cell_6t
Xbit_r247_c94 bl[94] br[94] wl[247] vdd gnd cell_6t
Xbit_r248_c94 bl[94] br[94] wl[248] vdd gnd cell_6t
Xbit_r249_c94 bl[94] br[94] wl[249] vdd gnd cell_6t
Xbit_r250_c94 bl[94] br[94] wl[250] vdd gnd cell_6t
Xbit_r251_c94 bl[94] br[94] wl[251] vdd gnd cell_6t
Xbit_r252_c94 bl[94] br[94] wl[252] vdd gnd cell_6t
Xbit_r253_c94 bl[94] br[94] wl[253] vdd gnd cell_6t
Xbit_r254_c94 bl[94] br[94] wl[254] vdd gnd cell_6t
Xbit_r255_c94 bl[94] br[94] wl[255] vdd gnd cell_6t
Xbit_r0_c95 bl[95] br[95] wl[0] vdd gnd cell_6t
Xbit_r1_c95 bl[95] br[95] wl[1] vdd gnd cell_6t
Xbit_r2_c95 bl[95] br[95] wl[2] vdd gnd cell_6t
Xbit_r3_c95 bl[95] br[95] wl[3] vdd gnd cell_6t
Xbit_r4_c95 bl[95] br[95] wl[4] vdd gnd cell_6t
Xbit_r5_c95 bl[95] br[95] wl[5] vdd gnd cell_6t
Xbit_r6_c95 bl[95] br[95] wl[6] vdd gnd cell_6t
Xbit_r7_c95 bl[95] br[95] wl[7] vdd gnd cell_6t
Xbit_r8_c95 bl[95] br[95] wl[8] vdd gnd cell_6t
Xbit_r9_c95 bl[95] br[95] wl[9] vdd gnd cell_6t
Xbit_r10_c95 bl[95] br[95] wl[10] vdd gnd cell_6t
Xbit_r11_c95 bl[95] br[95] wl[11] vdd gnd cell_6t
Xbit_r12_c95 bl[95] br[95] wl[12] vdd gnd cell_6t
Xbit_r13_c95 bl[95] br[95] wl[13] vdd gnd cell_6t
Xbit_r14_c95 bl[95] br[95] wl[14] vdd gnd cell_6t
Xbit_r15_c95 bl[95] br[95] wl[15] vdd gnd cell_6t
Xbit_r16_c95 bl[95] br[95] wl[16] vdd gnd cell_6t
Xbit_r17_c95 bl[95] br[95] wl[17] vdd gnd cell_6t
Xbit_r18_c95 bl[95] br[95] wl[18] vdd gnd cell_6t
Xbit_r19_c95 bl[95] br[95] wl[19] vdd gnd cell_6t
Xbit_r20_c95 bl[95] br[95] wl[20] vdd gnd cell_6t
Xbit_r21_c95 bl[95] br[95] wl[21] vdd gnd cell_6t
Xbit_r22_c95 bl[95] br[95] wl[22] vdd gnd cell_6t
Xbit_r23_c95 bl[95] br[95] wl[23] vdd gnd cell_6t
Xbit_r24_c95 bl[95] br[95] wl[24] vdd gnd cell_6t
Xbit_r25_c95 bl[95] br[95] wl[25] vdd gnd cell_6t
Xbit_r26_c95 bl[95] br[95] wl[26] vdd gnd cell_6t
Xbit_r27_c95 bl[95] br[95] wl[27] vdd gnd cell_6t
Xbit_r28_c95 bl[95] br[95] wl[28] vdd gnd cell_6t
Xbit_r29_c95 bl[95] br[95] wl[29] vdd gnd cell_6t
Xbit_r30_c95 bl[95] br[95] wl[30] vdd gnd cell_6t
Xbit_r31_c95 bl[95] br[95] wl[31] vdd gnd cell_6t
Xbit_r32_c95 bl[95] br[95] wl[32] vdd gnd cell_6t
Xbit_r33_c95 bl[95] br[95] wl[33] vdd gnd cell_6t
Xbit_r34_c95 bl[95] br[95] wl[34] vdd gnd cell_6t
Xbit_r35_c95 bl[95] br[95] wl[35] vdd gnd cell_6t
Xbit_r36_c95 bl[95] br[95] wl[36] vdd gnd cell_6t
Xbit_r37_c95 bl[95] br[95] wl[37] vdd gnd cell_6t
Xbit_r38_c95 bl[95] br[95] wl[38] vdd gnd cell_6t
Xbit_r39_c95 bl[95] br[95] wl[39] vdd gnd cell_6t
Xbit_r40_c95 bl[95] br[95] wl[40] vdd gnd cell_6t
Xbit_r41_c95 bl[95] br[95] wl[41] vdd gnd cell_6t
Xbit_r42_c95 bl[95] br[95] wl[42] vdd gnd cell_6t
Xbit_r43_c95 bl[95] br[95] wl[43] vdd gnd cell_6t
Xbit_r44_c95 bl[95] br[95] wl[44] vdd gnd cell_6t
Xbit_r45_c95 bl[95] br[95] wl[45] vdd gnd cell_6t
Xbit_r46_c95 bl[95] br[95] wl[46] vdd gnd cell_6t
Xbit_r47_c95 bl[95] br[95] wl[47] vdd gnd cell_6t
Xbit_r48_c95 bl[95] br[95] wl[48] vdd gnd cell_6t
Xbit_r49_c95 bl[95] br[95] wl[49] vdd gnd cell_6t
Xbit_r50_c95 bl[95] br[95] wl[50] vdd gnd cell_6t
Xbit_r51_c95 bl[95] br[95] wl[51] vdd gnd cell_6t
Xbit_r52_c95 bl[95] br[95] wl[52] vdd gnd cell_6t
Xbit_r53_c95 bl[95] br[95] wl[53] vdd gnd cell_6t
Xbit_r54_c95 bl[95] br[95] wl[54] vdd gnd cell_6t
Xbit_r55_c95 bl[95] br[95] wl[55] vdd gnd cell_6t
Xbit_r56_c95 bl[95] br[95] wl[56] vdd gnd cell_6t
Xbit_r57_c95 bl[95] br[95] wl[57] vdd gnd cell_6t
Xbit_r58_c95 bl[95] br[95] wl[58] vdd gnd cell_6t
Xbit_r59_c95 bl[95] br[95] wl[59] vdd gnd cell_6t
Xbit_r60_c95 bl[95] br[95] wl[60] vdd gnd cell_6t
Xbit_r61_c95 bl[95] br[95] wl[61] vdd gnd cell_6t
Xbit_r62_c95 bl[95] br[95] wl[62] vdd gnd cell_6t
Xbit_r63_c95 bl[95] br[95] wl[63] vdd gnd cell_6t
Xbit_r64_c95 bl[95] br[95] wl[64] vdd gnd cell_6t
Xbit_r65_c95 bl[95] br[95] wl[65] vdd gnd cell_6t
Xbit_r66_c95 bl[95] br[95] wl[66] vdd gnd cell_6t
Xbit_r67_c95 bl[95] br[95] wl[67] vdd gnd cell_6t
Xbit_r68_c95 bl[95] br[95] wl[68] vdd gnd cell_6t
Xbit_r69_c95 bl[95] br[95] wl[69] vdd gnd cell_6t
Xbit_r70_c95 bl[95] br[95] wl[70] vdd gnd cell_6t
Xbit_r71_c95 bl[95] br[95] wl[71] vdd gnd cell_6t
Xbit_r72_c95 bl[95] br[95] wl[72] vdd gnd cell_6t
Xbit_r73_c95 bl[95] br[95] wl[73] vdd gnd cell_6t
Xbit_r74_c95 bl[95] br[95] wl[74] vdd gnd cell_6t
Xbit_r75_c95 bl[95] br[95] wl[75] vdd gnd cell_6t
Xbit_r76_c95 bl[95] br[95] wl[76] vdd gnd cell_6t
Xbit_r77_c95 bl[95] br[95] wl[77] vdd gnd cell_6t
Xbit_r78_c95 bl[95] br[95] wl[78] vdd gnd cell_6t
Xbit_r79_c95 bl[95] br[95] wl[79] vdd gnd cell_6t
Xbit_r80_c95 bl[95] br[95] wl[80] vdd gnd cell_6t
Xbit_r81_c95 bl[95] br[95] wl[81] vdd gnd cell_6t
Xbit_r82_c95 bl[95] br[95] wl[82] vdd gnd cell_6t
Xbit_r83_c95 bl[95] br[95] wl[83] vdd gnd cell_6t
Xbit_r84_c95 bl[95] br[95] wl[84] vdd gnd cell_6t
Xbit_r85_c95 bl[95] br[95] wl[85] vdd gnd cell_6t
Xbit_r86_c95 bl[95] br[95] wl[86] vdd gnd cell_6t
Xbit_r87_c95 bl[95] br[95] wl[87] vdd gnd cell_6t
Xbit_r88_c95 bl[95] br[95] wl[88] vdd gnd cell_6t
Xbit_r89_c95 bl[95] br[95] wl[89] vdd gnd cell_6t
Xbit_r90_c95 bl[95] br[95] wl[90] vdd gnd cell_6t
Xbit_r91_c95 bl[95] br[95] wl[91] vdd gnd cell_6t
Xbit_r92_c95 bl[95] br[95] wl[92] vdd gnd cell_6t
Xbit_r93_c95 bl[95] br[95] wl[93] vdd gnd cell_6t
Xbit_r94_c95 bl[95] br[95] wl[94] vdd gnd cell_6t
Xbit_r95_c95 bl[95] br[95] wl[95] vdd gnd cell_6t
Xbit_r96_c95 bl[95] br[95] wl[96] vdd gnd cell_6t
Xbit_r97_c95 bl[95] br[95] wl[97] vdd gnd cell_6t
Xbit_r98_c95 bl[95] br[95] wl[98] vdd gnd cell_6t
Xbit_r99_c95 bl[95] br[95] wl[99] vdd gnd cell_6t
Xbit_r100_c95 bl[95] br[95] wl[100] vdd gnd cell_6t
Xbit_r101_c95 bl[95] br[95] wl[101] vdd gnd cell_6t
Xbit_r102_c95 bl[95] br[95] wl[102] vdd gnd cell_6t
Xbit_r103_c95 bl[95] br[95] wl[103] vdd gnd cell_6t
Xbit_r104_c95 bl[95] br[95] wl[104] vdd gnd cell_6t
Xbit_r105_c95 bl[95] br[95] wl[105] vdd gnd cell_6t
Xbit_r106_c95 bl[95] br[95] wl[106] vdd gnd cell_6t
Xbit_r107_c95 bl[95] br[95] wl[107] vdd gnd cell_6t
Xbit_r108_c95 bl[95] br[95] wl[108] vdd gnd cell_6t
Xbit_r109_c95 bl[95] br[95] wl[109] vdd gnd cell_6t
Xbit_r110_c95 bl[95] br[95] wl[110] vdd gnd cell_6t
Xbit_r111_c95 bl[95] br[95] wl[111] vdd gnd cell_6t
Xbit_r112_c95 bl[95] br[95] wl[112] vdd gnd cell_6t
Xbit_r113_c95 bl[95] br[95] wl[113] vdd gnd cell_6t
Xbit_r114_c95 bl[95] br[95] wl[114] vdd gnd cell_6t
Xbit_r115_c95 bl[95] br[95] wl[115] vdd gnd cell_6t
Xbit_r116_c95 bl[95] br[95] wl[116] vdd gnd cell_6t
Xbit_r117_c95 bl[95] br[95] wl[117] vdd gnd cell_6t
Xbit_r118_c95 bl[95] br[95] wl[118] vdd gnd cell_6t
Xbit_r119_c95 bl[95] br[95] wl[119] vdd gnd cell_6t
Xbit_r120_c95 bl[95] br[95] wl[120] vdd gnd cell_6t
Xbit_r121_c95 bl[95] br[95] wl[121] vdd gnd cell_6t
Xbit_r122_c95 bl[95] br[95] wl[122] vdd gnd cell_6t
Xbit_r123_c95 bl[95] br[95] wl[123] vdd gnd cell_6t
Xbit_r124_c95 bl[95] br[95] wl[124] vdd gnd cell_6t
Xbit_r125_c95 bl[95] br[95] wl[125] vdd gnd cell_6t
Xbit_r126_c95 bl[95] br[95] wl[126] vdd gnd cell_6t
Xbit_r127_c95 bl[95] br[95] wl[127] vdd gnd cell_6t
Xbit_r128_c95 bl[95] br[95] wl[128] vdd gnd cell_6t
Xbit_r129_c95 bl[95] br[95] wl[129] vdd gnd cell_6t
Xbit_r130_c95 bl[95] br[95] wl[130] vdd gnd cell_6t
Xbit_r131_c95 bl[95] br[95] wl[131] vdd gnd cell_6t
Xbit_r132_c95 bl[95] br[95] wl[132] vdd gnd cell_6t
Xbit_r133_c95 bl[95] br[95] wl[133] vdd gnd cell_6t
Xbit_r134_c95 bl[95] br[95] wl[134] vdd gnd cell_6t
Xbit_r135_c95 bl[95] br[95] wl[135] vdd gnd cell_6t
Xbit_r136_c95 bl[95] br[95] wl[136] vdd gnd cell_6t
Xbit_r137_c95 bl[95] br[95] wl[137] vdd gnd cell_6t
Xbit_r138_c95 bl[95] br[95] wl[138] vdd gnd cell_6t
Xbit_r139_c95 bl[95] br[95] wl[139] vdd gnd cell_6t
Xbit_r140_c95 bl[95] br[95] wl[140] vdd gnd cell_6t
Xbit_r141_c95 bl[95] br[95] wl[141] vdd gnd cell_6t
Xbit_r142_c95 bl[95] br[95] wl[142] vdd gnd cell_6t
Xbit_r143_c95 bl[95] br[95] wl[143] vdd gnd cell_6t
Xbit_r144_c95 bl[95] br[95] wl[144] vdd gnd cell_6t
Xbit_r145_c95 bl[95] br[95] wl[145] vdd gnd cell_6t
Xbit_r146_c95 bl[95] br[95] wl[146] vdd gnd cell_6t
Xbit_r147_c95 bl[95] br[95] wl[147] vdd gnd cell_6t
Xbit_r148_c95 bl[95] br[95] wl[148] vdd gnd cell_6t
Xbit_r149_c95 bl[95] br[95] wl[149] vdd gnd cell_6t
Xbit_r150_c95 bl[95] br[95] wl[150] vdd gnd cell_6t
Xbit_r151_c95 bl[95] br[95] wl[151] vdd gnd cell_6t
Xbit_r152_c95 bl[95] br[95] wl[152] vdd gnd cell_6t
Xbit_r153_c95 bl[95] br[95] wl[153] vdd gnd cell_6t
Xbit_r154_c95 bl[95] br[95] wl[154] vdd gnd cell_6t
Xbit_r155_c95 bl[95] br[95] wl[155] vdd gnd cell_6t
Xbit_r156_c95 bl[95] br[95] wl[156] vdd gnd cell_6t
Xbit_r157_c95 bl[95] br[95] wl[157] vdd gnd cell_6t
Xbit_r158_c95 bl[95] br[95] wl[158] vdd gnd cell_6t
Xbit_r159_c95 bl[95] br[95] wl[159] vdd gnd cell_6t
Xbit_r160_c95 bl[95] br[95] wl[160] vdd gnd cell_6t
Xbit_r161_c95 bl[95] br[95] wl[161] vdd gnd cell_6t
Xbit_r162_c95 bl[95] br[95] wl[162] vdd gnd cell_6t
Xbit_r163_c95 bl[95] br[95] wl[163] vdd gnd cell_6t
Xbit_r164_c95 bl[95] br[95] wl[164] vdd gnd cell_6t
Xbit_r165_c95 bl[95] br[95] wl[165] vdd gnd cell_6t
Xbit_r166_c95 bl[95] br[95] wl[166] vdd gnd cell_6t
Xbit_r167_c95 bl[95] br[95] wl[167] vdd gnd cell_6t
Xbit_r168_c95 bl[95] br[95] wl[168] vdd gnd cell_6t
Xbit_r169_c95 bl[95] br[95] wl[169] vdd gnd cell_6t
Xbit_r170_c95 bl[95] br[95] wl[170] vdd gnd cell_6t
Xbit_r171_c95 bl[95] br[95] wl[171] vdd gnd cell_6t
Xbit_r172_c95 bl[95] br[95] wl[172] vdd gnd cell_6t
Xbit_r173_c95 bl[95] br[95] wl[173] vdd gnd cell_6t
Xbit_r174_c95 bl[95] br[95] wl[174] vdd gnd cell_6t
Xbit_r175_c95 bl[95] br[95] wl[175] vdd gnd cell_6t
Xbit_r176_c95 bl[95] br[95] wl[176] vdd gnd cell_6t
Xbit_r177_c95 bl[95] br[95] wl[177] vdd gnd cell_6t
Xbit_r178_c95 bl[95] br[95] wl[178] vdd gnd cell_6t
Xbit_r179_c95 bl[95] br[95] wl[179] vdd gnd cell_6t
Xbit_r180_c95 bl[95] br[95] wl[180] vdd gnd cell_6t
Xbit_r181_c95 bl[95] br[95] wl[181] vdd gnd cell_6t
Xbit_r182_c95 bl[95] br[95] wl[182] vdd gnd cell_6t
Xbit_r183_c95 bl[95] br[95] wl[183] vdd gnd cell_6t
Xbit_r184_c95 bl[95] br[95] wl[184] vdd gnd cell_6t
Xbit_r185_c95 bl[95] br[95] wl[185] vdd gnd cell_6t
Xbit_r186_c95 bl[95] br[95] wl[186] vdd gnd cell_6t
Xbit_r187_c95 bl[95] br[95] wl[187] vdd gnd cell_6t
Xbit_r188_c95 bl[95] br[95] wl[188] vdd gnd cell_6t
Xbit_r189_c95 bl[95] br[95] wl[189] vdd gnd cell_6t
Xbit_r190_c95 bl[95] br[95] wl[190] vdd gnd cell_6t
Xbit_r191_c95 bl[95] br[95] wl[191] vdd gnd cell_6t
Xbit_r192_c95 bl[95] br[95] wl[192] vdd gnd cell_6t
Xbit_r193_c95 bl[95] br[95] wl[193] vdd gnd cell_6t
Xbit_r194_c95 bl[95] br[95] wl[194] vdd gnd cell_6t
Xbit_r195_c95 bl[95] br[95] wl[195] vdd gnd cell_6t
Xbit_r196_c95 bl[95] br[95] wl[196] vdd gnd cell_6t
Xbit_r197_c95 bl[95] br[95] wl[197] vdd gnd cell_6t
Xbit_r198_c95 bl[95] br[95] wl[198] vdd gnd cell_6t
Xbit_r199_c95 bl[95] br[95] wl[199] vdd gnd cell_6t
Xbit_r200_c95 bl[95] br[95] wl[200] vdd gnd cell_6t
Xbit_r201_c95 bl[95] br[95] wl[201] vdd gnd cell_6t
Xbit_r202_c95 bl[95] br[95] wl[202] vdd gnd cell_6t
Xbit_r203_c95 bl[95] br[95] wl[203] vdd gnd cell_6t
Xbit_r204_c95 bl[95] br[95] wl[204] vdd gnd cell_6t
Xbit_r205_c95 bl[95] br[95] wl[205] vdd gnd cell_6t
Xbit_r206_c95 bl[95] br[95] wl[206] vdd gnd cell_6t
Xbit_r207_c95 bl[95] br[95] wl[207] vdd gnd cell_6t
Xbit_r208_c95 bl[95] br[95] wl[208] vdd gnd cell_6t
Xbit_r209_c95 bl[95] br[95] wl[209] vdd gnd cell_6t
Xbit_r210_c95 bl[95] br[95] wl[210] vdd gnd cell_6t
Xbit_r211_c95 bl[95] br[95] wl[211] vdd gnd cell_6t
Xbit_r212_c95 bl[95] br[95] wl[212] vdd gnd cell_6t
Xbit_r213_c95 bl[95] br[95] wl[213] vdd gnd cell_6t
Xbit_r214_c95 bl[95] br[95] wl[214] vdd gnd cell_6t
Xbit_r215_c95 bl[95] br[95] wl[215] vdd gnd cell_6t
Xbit_r216_c95 bl[95] br[95] wl[216] vdd gnd cell_6t
Xbit_r217_c95 bl[95] br[95] wl[217] vdd gnd cell_6t
Xbit_r218_c95 bl[95] br[95] wl[218] vdd gnd cell_6t
Xbit_r219_c95 bl[95] br[95] wl[219] vdd gnd cell_6t
Xbit_r220_c95 bl[95] br[95] wl[220] vdd gnd cell_6t
Xbit_r221_c95 bl[95] br[95] wl[221] vdd gnd cell_6t
Xbit_r222_c95 bl[95] br[95] wl[222] vdd gnd cell_6t
Xbit_r223_c95 bl[95] br[95] wl[223] vdd gnd cell_6t
Xbit_r224_c95 bl[95] br[95] wl[224] vdd gnd cell_6t
Xbit_r225_c95 bl[95] br[95] wl[225] vdd gnd cell_6t
Xbit_r226_c95 bl[95] br[95] wl[226] vdd gnd cell_6t
Xbit_r227_c95 bl[95] br[95] wl[227] vdd gnd cell_6t
Xbit_r228_c95 bl[95] br[95] wl[228] vdd gnd cell_6t
Xbit_r229_c95 bl[95] br[95] wl[229] vdd gnd cell_6t
Xbit_r230_c95 bl[95] br[95] wl[230] vdd gnd cell_6t
Xbit_r231_c95 bl[95] br[95] wl[231] vdd gnd cell_6t
Xbit_r232_c95 bl[95] br[95] wl[232] vdd gnd cell_6t
Xbit_r233_c95 bl[95] br[95] wl[233] vdd gnd cell_6t
Xbit_r234_c95 bl[95] br[95] wl[234] vdd gnd cell_6t
Xbit_r235_c95 bl[95] br[95] wl[235] vdd gnd cell_6t
Xbit_r236_c95 bl[95] br[95] wl[236] vdd gnd cell_6t
Xbit_r237_c95 bl[95] br[95] wl[237] vdd gnd cell_6t
Xbit_r238_c95 bl[95] br[95] wl[238] vdd gnd cell_6t
Xbit_r239_c95 bl[95] br[95] wl[239] vdd gnd cell_6t
Xbit_r240_c95 bl[95] br[95] wl[240] vdd gnd cell_6t
Xbit_r241_c95 bl[95] br[95] wl[241] vdd gnd cell_6t
Xbit_r242_c95 bl[95] br[95] wl[242] vdd gnd cell_6t
Xbit_r243_c95 bl[95] br[95] wl[243] vdd gnd cell_6t
Xbit_r244_c95 bl[95] br[95] wl[244] vdd gnd cell_6t
Xbit_r245_c95 bl[95] br[95] wl[245] vdd gnd cell_6t
Xbit_r246_c95 bl[95] br[95] wl[246] vdd gnd cell_6t
Xbit_r247_c95 bl[95] br[95] wl[247] vdd gnd cell_6t
Xbit_r248_c95 bl[95] br[95] wl[248] vdd gnd cell_6t
Xbit_r249_c95 bl[95] br[95] wl[249] vdd gnd cell_6t
Xbit_r250_c95 bl[95] br[95] wl[250] vdd gnd cell_6t
Xbit_r251_c95 bl[95] br[95] wl[251] vdd gnd cell_6t
Xbit_r252_c95 bl[95] br[95] wl[252] vdd gnd cell_6t
Xbit_r253_c95 bl[95] br[95] wl[253] vdd gnd cell_6t
Xbit_r254_c95 bl[95] br[95] wl[254] vdd gnd cell_6t
Xbit_r255_c95 bl[95] br[95] wl[255] vdd gnd cell_6t
Xbit_r0_c96 bl[96] br[96] wl[0] vdd gnd cell_6t
Xbit_r1_c96 bl[96] br[96] wl[1] vdd gnd cell_6t
Xbit_r2_c96 bl[96] br[96] wl[2] vdd gnd cell_6t
Xbit_r3_c96 bl[96] br[96] wl[3] vdd gnd cell_6t
Xbit_r4_c96 bl[96] br[96] wl[4] vdd gnd cell_6t
Xbit_r5_c96 bl[96] br[96] wl[5] vdd gnd cell_6t
Xbit_r6_c96 bl[96] br[96] wl[6] vdd gnd cell_6t
Xbit_r7_c96 bl[96] br[96] wl[7] vdd gnd cell_6t
Xbit_r8_c96 bl[96] br[96] wl[8] vdd gnd cell_6t
Xbit_r9_c96 bl[96] br[96] wl[9] vdd gnd cell_6t
Xbit_r10_c96 bl[96] br[96] wl[10] vdd gnd cell_6t
Xbit_r11_c96 bl[96] br[96] wl[11] vdd gnd cell_6t
Xbit_r12_c96 bl[96] br[96] wl[12] vdd gnd cell_6t
Xbit_r13_c96 bl[96] br[96] wl[13] vdd gnd cell_6t
Xbit_r14_c96 bl[96] br[96] wl[14] vdd gnd cell_6t
Xbit_r15_c96 bl[96] br[96] wl[15] vdd gnd cell_6t
Xbit_r16_c96 bl[96] br[96] wl[16] vdd gnd cell_6t
Xbit_r17_c96 bl[96] br[96] wl[17] vdd gnd cell_6t
Xbit_r18_c96 bl[96] br[96] wl[18] vdd gnd cell_6t
Xbit_r19_c96 bl[96] br[96] wl[19] vdd gnd cell_6t
Xbit_r20_c96 bl[96] br[96] wl[20] vdd gnd cell_6t
Xbit_r21_c96 bl[96] br[96] wl[21] vdd gnd cell_6t
Xbit_r22_c96 bl[96] br[96] wl[22] vdd gnd cell_6t
Xbit_r23_c96 bl[96] br[96] wl[23] vdd gnd cell_6t
Xbit_r24_c96 bl[96] br[96] wl[24] vdd gnd cell_6t
Xbit_r25_c96 bl[96] br[96] wl[25] vdd gnd cell_6t
Xbit_r26_c96 bl[96] br[96] wl[26] vdd gnd cell_6t
Xbit_r27_c96 bl[96] br[96] wl[27] vdd gnd cell_6t
Xbit_r28_c96 bl[96] br[96] wl[28] vdd gnd cell_6t
Xbit_r29_c96 bl[96] br[96] wl[29] vdd gnd cell_6t
Xbit_r30_c96 bl[96] br[96] wl[30] vdd gnd cell_6t
Xbit_r31_c96 bl[96] br[96] wl[31] vdd gnd cell_6t
Xbit_r32_c96 bl[96] br[96] wl[32] vdd gnd cell_6t
Xbit_r33_c96 bl[96] br[96] wl[33] vdd gnd cell_6t
Xbit_r34_c96 bl[96] br[96] wl[34] vdd gnd cell_6t
Xbit_r35_c96 bl[96] br[96] wl[35] vdd gnd cell_6t
Xbit_r36_c96 bl[96] br[96] wl[36] vdd gnd cell_6t
Xbit_r37_c96 bl[96] br[96] wl[37] vdd gnd cell_6t
Xbit_r38_c96 bl[96] br[96] wl[38] vdd gnd cell_6t
Xbit_r39_c96 bl[96] br[96] wl[39] vdd gnd cell_6t
Xbit_r40_c96 bl[96] br[96] wl[40] vdd gnd cell_6t
Xbit_r41_c96 bl[96] br[96] wl[41] vdd gnd cell_6t
Xbit_r42_c96 bl[96] br[96] wl[42] vdd gnd cell_6t
Xbit_r43_c96 bl[96] br[96] wl[43] vdd gnd cell_6t
Xbit_r44_c96 bl[96] br[96] wl[44] vdd gnd cell_6t
Xbit_r45_c96 bl[96] br[96] wl[45] vdd gnd cell_6t
Xbit_r46_c96 bl[96] br[96] wl[46] vdd gnd cell_6t
Xbit_r47_c96 bl[96] br[96] wl[47] vdd gnd cell_6t
Xbit_r48_c96 bl[96] br[96] wl[48] vdd gnd cell_6t
Xbit_r49_c96 bl[96] br[96] wl[49] vdd gnd cell_6t
Xbit_r50_c96 bl[96] br[96] wl[50] vdd gnd cell_6t
Xbit_r51_c96 bl[96] br[96] wl[51] vdd gnd cell_6t
Xbit_r52_c96 bl[96] br[96] wl[52] vdd gnd cell_6t
Xbit_r53_c96 bl[96] br[96] wl[53] vdd gnd cell_6t
Xbit_r54_c96 bl[96] br[96] wl[54] vdd gnd cell_6t
Xbit_r55_c96 bl[96] br[96] wl[55] vdd gnd cell_6t
Xbit_r56_c96 bl[96] br[96] wl[56] vdd gnd cell_6t
Xbit_r57_c96 bl[96] br[96] wl[57] vdd gnd cell_6t
Xbit_r58_c96 bl[96] br[96] wl[58] vdd gnd cell_6t
Xbit_r59_c96 bl[96] br[96] wl[59] vdd gnd cell_6t
Xbit_r60_c96 bl[96] br[96] wl[60] vdd gnd cell_6t
Xbit_r61_c96 bl[96] br[96] wl[61] vdd gnd cell_6t
Xbit_r62_c96 bl[96] br[96] wl[62] vdd gnd cell_6t
Xbit_r63_c96 bl[96] br[96] wl[63] vdd gnd cell_6t
Xbit_r64_c96 bl[96] br[96] wl[64] vdd gnd cell_6t
Xbit_r65_c96 bl[96] br[96] wl[65] vdd gnd cell_6t
Xbit_r66_c96 bl[96] br[96] wl[66] vdd gnd cell_6t
Xbit_r67_c96 bl[96] br[96] wl[67] vdd gnd cell_6t
Xbit_r68_c96 bl[96] br[96] wl[68] vdd gnd cell_6t
Xbit_r69_c96 bl[96] br[96] wl[69] vdd gnd cell_6t
Xbit_r70_c96 bl[96] br[96] wl[70] vdd gnd cell_6t
Xbit_r71_c96 bl[96] br[96] wl[71] vdd gnd cell_6t
Xbit_r72_c96 bl[96] br[96] wl[72] vdd gnd cell_6t
Xbit_r73_c96 bl[96] br[96] wl[73] vdd gnd cell_6t
Xbit_r74_c96 bl[96] br[96] wl[74] vdd gnd cell_6t
Xbit_r75_c96 bl[96] br[96] wl[75] vdd gnd cell_6t
Xbit_r76_c96 bl[96] br[96] wl[76] vdd gnd cell_6t
Xbit_r77_c96 bl[96] br[96] wl[77] vdd gnd cell_6t
Xbit_r78_c96 bl[96] br[96] wl[78] vdd gnd cell_6t
Xbit_r79_c96 bl[96] br[96] wl[79] vdd gnd cell_6t
Xbit_r80_c96 bl[96] br[96] wl[80] vdd gnd cell_6t
Xbit_r81_c96 bl[96] br[96] wl[81] vdd gnd cell_6t
Xbit_r82_c96 bl[96] br[96] wl[82] vdd gnd cell_6t
Xbit_r83_c96 bl[96] br[96] wl[83] vdd gnd cell_6t
Xbit_r84_c96 bl[96] br[96] wl[84] vdd gnd cell_6t
Xbit_r85_c96 bl[96] br[96] wl[85] vdd gnd cell_6t
Xbit_r86_c96 bl[96] br[96] wl[86] vdd gnd cell_6t
Xbit_r87_c96 bl[96] br[96] wl[87] vdd gnd cell_6t
Xbit_r88_c96 bl[96] br[96] wl[88] vdd gnd cell_6t
Xbit_r89_c96 bl[96] br[96] wl[89] vdd gnd cell_6t
Xbit_r90_c96 bl[96] br[96] wl[90] vdd gnd cell_6t
Xbit_r91_c96 bl[96] br[96] wl[91] vdd gnd cell_6t
Xbit_r92_c96 bl[96] br[96] wl[92] vdd gnd cell_6t
Xbit_r93_c96 bl[96] br[96] wl[93] vdd gnd cell_6t
Xbit_r94_c96 bl[96] br[96] wl[94] vdd gnd cell_6t
Xbit_r95_c96 bl[96] br[96] wl[95] vdd gnd cell_6t
Xbit_r96_c96 bl[96] br[96] wl[96] vdd gnd cell_6t
Xbit_r97_c96 bl[96] br[96] wl[97] vdd gnd cell_6t
Xbit_r98_c96 bl[96] br[96] wl[98] vdd gnd cell_6t
Xbit_r99_c96 bl[96] br[96] wl[99] vdd gnd cell_6t
Xbit_r100_c96 bl[96] br[96] wl[100] vdd gnd cell_6t
Xbit_r101_c96 bl[96] br[96] wl[101] vdd gnd cell_6t
Xbit_r102_c96 bl[96] br[96] wl[102] vdd gnd cell_6t
Xbit_r103_c96 bl[96] br[96] wl[103] vdd gnd cell_6t
Xbit_r104_c96 bl[96] br[96] wl[104] vdd gnd cell_6t
Xbit_r105_c96 bl[96] br[96] wl[105] vdd gnd cell_6t
Xbit_r106_c96 bl[96] br[96] wl[106] vdd gnd cell_6t
Xbit_r107_c96 bl[96] br[96] wl[107] vdd gnd cell_6t
Xbit_r108_c96 bl[96] br[96] wl[108] vdd gnd cell_6t
Xbit_r109_c96 bl[96] br[96] wl[109] vdd gnd cell_6t
Xbit_r110_c96 bl[96] br[96] wl[110] vdd gnd cell_6t
Xbit_r111_c96 bl[96] br[96] wl[111] vdd gnd cell_6t
Xbit_r112_c96 bl[96] br[96] wl[112] vdd gnd cell_6t
Xbit_r113_c96 bl[96] br[96] wl[113] vdd gnd cell_6t
Xbit_r114_c96 bl[96] br[96] wl[114] vdd gnd cell_6t
Xbit_r115_c96 bl[96] br[96] wl[115] vdd gnd cell_6t
Xbit_r116_c96 bl[96] br[96] wl[116] vdd gnd cell_6t
Xbit_r117_c96 bl[96] br[96] wl[117] vdd gnd cell_6t
Xbit_r118_c96 bl[96] br[96] wl[118] vdd gnd cell_6t
Xbit_r119_c96 bl[96] br[96] wl[119] vdd gnd cell_6t
Xbit_r120_c96 bl[96] br[96] wl[120] vdd gnd cell_6t
Xbit_r121_c96 bl[96] br[96] wl[121] vdd gnd cell_6t
Xbit_r122_c96 bl[96] br[96] wl[122] vdd gnd cell_6t
Xbit_r123_c96 bl[96] br[96] wl[123] vdd gnd cell_6t
Xbit_r124_c96 bl[96] br[96] wl[124] vdd gnd cell_6t
Xbit_r125_c96 bl[96] br[96] wl[125] vdd gnd cell_6t
Xbit_r126_c96 bl[96] br[96] wl[126] vdd gnd cell_6t
Xbit_r127_c96 bl[96] br[96] wl[127] vdd gnd cell_6t
Xbit_r128_c96 bl[96] br[96] wl[128] vdd gnd cell_6t
Xbit_r129_c96 bl[96] br[96] wl[129] vdd gnd cell_6t
Xbit_r130_c96 bl[96] br[96] wl[130] vdd gnd cell_6t
Xbit_r131_c96 bl[96] br[96] wl[131] vdd gnd cell_6t
Xbit_r132_c96 bl[96] br[96] wl[132] vdd gnd cell_6t
Xbit_r133_c96 bl[96] br[96] wl[133] vdd gnd cell_6t
Xbit_r134_c96 bl[96] br[96] wl[134] vdd gnd cell_6t
Xbit_r135_c96 bl[96] br[96] wl[135] vdd gnd cell_6t
Xbit_r136_c96 bl[96] br[96] wl[136] vdd gnd cell_6t
Xbit_r137_c96 bl[96] br[96] wl[137] vdd gnd cell_6t
Xbit_r138_c96 bl[96] br[96] wl[138] vdd gnd cell_6t
Xbit_r139_c96 bl[96] br[96] wl[139] vdd gnd cell_6t
Xbit_r140_c96 bl[96] br[96] wl[140] vdd gnd cell_6t
Xbit_r141_c96 bl[96] br[96] wl[141] vdd gnd cell_6t
Xbit_r142_c96 bl[96] br[96] wl[142] vdd gnd cell_6t
Xbit_r143_c96 bl[96] br[96] wl[143] vdd gnd cell_6t
Xbit_r144_c96 bl[96] br[96] wl[144] vdd gnd cell_6t
Xbit_r145_c96 bl[96] br[96] wl[145] vdd gnd cell_6t
Xbit_r146_c96 bl[96] br[96] wl[146] vdd gnd cell_6t
Xbit_r147_c96 bl[96] br[96] wl[147] vdd gnd cell_6t
Xbit_r148_c96 bl[96] br[96] wl[148] vdd gnd cell_6t
Xbit_r149_c96 bl[96] br[96] wl[149] vdd gnd cell_6t
Xbit_r150_c96 bl[96] br[96] wl[150] vdd gnd cell_6t
Xbit_r151_c96 bl[96] br[96] wl[151] vdd gnd cell_6t
Xbit_r152_c96 bl[96] br[96] wl[152] vdd gnd cell_6t
Xbit_r153_c96 bl[96] br[96] wl[153] vdd gnd cell_6t
Xbit_r154_c96 bl[96] br[96] wl[154] vdd gnd cell_6t
Xbit_r155_c96 bl[96] br[96] wl[155] vdd gnd cell_6t
Xbit_r156_c96 bl[96] br[96] wl[156] vdd gnd cell_6t
Xbit_r157_c96 bl[96] br[96] wl[157] vdd gnd cell_6t
Xbit_r158_c96 bl[96] br[96] wl[158] vdd gnd cell_6t
Xbit_r159_c96 bl[96] br[96] wl[159] vdd gnd cell_6t
Xbit_r160_c96 bl[96] br[96] wl[160] vdd gnd cell_6t
Xbit_r161_c96 bl[96] br[96] wl[161] vdd gnd cell_6t
Xbit_r162_c96 bl[96] br[96] wl[162] vdd gnd cell_6t
Xbit_r163_c96 bl[96] br[96] wl[163] vdd gnd cell_6t
Xbit_r164_c96 bl[96] br[96] wl[164] vdd gnd cell_6t
Xbit_r165_c96 bl[96] br[96] wl[165] vdd gnd cell_6t
Xbit_r166_c96 bl[96] br[96] wl[166] vdd gnd cell_6t
Xbit_r167_c96 bl[96] br[96] wl[167] vdd gnd cell_6t
Xbit_r168_c96 bl[96] br[96] wl[168] vdd gnd cell_6t
Xbit_r169_c96 bl[96] br[96] wl[169] vdd gnd cell_6t
Xbit_r170_c96 bl[96] br[96] wl[170] vdd gnd cell_6t
Xbit_r171_c96 bl[96] br[96] wl[171] vdd gnd cell_6t
Xbit_r172_c96 bl[96] br[96] wl[172] vdd gnd cell_6t
Xbit_r173_c96 bl[96] br[96] wl[173] vdd gnd cell_6t
Xbit_r174_c96 bl[96] br[96] wl[174] vdd gnd cell_6t
Xbit_r175_c96 bl[96] br[96] wl[175] vdd gnd cell_6t
Xbit_r176_c96 bl[96] br[96] wl[176] vdd gnd cell_6t
Xbit_r177_c96 bl[96] br[96] wl[177] vdd gnd cell_6t
Xbit_r178_c96 bl[96] br[96] wl[178] vdd gnd cell_6t
Xbit_r179_c96 bl[96] br[96] wl[179] vdd gnd cell_6t
Xbit_r180_c96 bl[96] br[96] wl[180] vdd gnd cell_6t
Xbit_r181_c96 bl[96] br[96] wl[181] vdd gnd cell_6t
Xbit_r182_c96 bl[96] br[96] wl[182] vdd gnd cell_6t
Xbit_r183_c96 bl[96] br[96] wl[183] vdd gnd cell_6t
Xbit_r184_c96 bl[96] br[96] wl[184] vdd gnd cell_6t
Xbit_r185_c96 bl[96] br[96] wl[185] vdd gnd cell_6t
Xbit_r186_c96 bl[96] br[96] wl[186] vdd gnd cell_6t
Xbit_r187_c96 bl[96] br[96] wl[187] vdd gnd cell_6t
Xbit_r188_c96 bl[96] br[96] wl[188] vdd gnd cell_6t
Xbit_r189_c96 bl[96] br[96] wl[189] vdd gnd cell_6t
Xbit_r190_c96 bl[96] br[96] wl[190] vdd gnd cell_6t
Xbit_r191_c96 bl[96] br[96] wl[191] vdd gnd cell_6t
Xbit_r192_c96 bl[96] br[96] wl[192] vdd gnd cell_6t
Xbit_r193_c96 bl[96] br[96] wl[193] vdd gnd cell_6t
Xbit_r194_c96 bl[96] br[96] wl[194] vdd gnd cell_6t
Xbit_r195_c96 bl[96] br[96] wl[195] vdd gnd cell_6t
Xbit_r196_c96 bl[96] br[96] wl[196] vdd gnd cell_6t
Xbit_r197_c96 bl[96] br[96] wl[197] vdd gnd cell_6t
Xbit_r198_c96 bl[96] br[96] wl[198] vdd gnd cell_6t
Xbit_r199_c96 bl[96] br[96] wl[199] vdd gnd cell_6t
Xbit_r200_c96 bl[96] br[96] wl[200] vdd gnd cell_6t
Xbit_r201_c96 bl[96] br[96] wl[201] vdd gnd cell_6t
Xbit_r202_c96 bl[96] br[96] wl[202] vdd gnd cell_6t
Xbit_r203_c96 bl[96] br[96] wl[203] vdd gnd cell_6t
Xbit_r204_c96 bl[96] br[96] wl[204] vdd gnd cell_6t
Xbit_r205_c96 bl[96] br[96] wl[205] vdd gnd cell_6t
Xbit_r206_c96 bl[96] br[96] wl[206] vdd gnd cell_6t
Xbit_r207_c96 bl[96] br[96] wl[207] vdd gnd cell_6t
Xbit_r208_c96 bl[96] br[96] wl[208] vdd gnd cell_6t
Xbit_r209_c96 bl[96] br[96] wl[209] vdd gnd cell_6t
Xbit_r210_c96 bl[96] br[96] wl[210] vdd gnd cell_6t
Xbit_r211_c96 bl[96] br[96] wl[211] vdd gnd cell_6t
Xbit_r212_c96 bl[96] br[96] wl[212] vdd gnd cell_6t
Xbit_r213_c96 bl[96] br[96] wl[213] vdd gnd cell_6t
Xbit_r214_c96 bl[96] br[96] wl[214] vdd gnd cell_6t
Xbit_r215_c96 bl[96] br[96] wl[215] vdd gnd cell_6t
Xbit_r216_c96 bl[96] br[96] wl[216] vdd gnd cell_6t
Xbit_r217_c96 bl[96] br[96] wl[217] vdd gnd cell_6t
Xbit_r218_c96 bl[96] br[96] wl[218] vdd gnd cell_6t
Xbit_r219_c96 bl[96] br[96] wl[219] vdd gnd cell_6t
Xbit_r220_c96 bl[96] br[96] wl[220] vdd gnd cell_6t
Xbit_r221_c96 bl[96] br[96] wl[221] vdd gnd cell_6t
Xbit_r222_c96 bl[96] br[96] wl[222] vdd gnd cell_6t
Xbit_r223_c96 bl[96] br[96] wl[223] vdd gnd cell_6t
Xbit_r224_c96 bl[96] br[96] wl[224] vdd gnd cell_6t
Xbit_r225_c96 bl[96] br[96] wl[225] vdd gnd cell_6t
Xbit_r226_c96 bl[96] br[96] wl[226] vdd gnd cell_6t
Xbit_r227_c96 bl[96] br[96] wl[227] vdd gnd cell_6t
Xbit_r228_c96 bl[96] br[96] wl[228] vdd gnd cell_6t
Xbit_r229_c96 bl[96] br[96] wl[229] vdd gnd cell_6t
Xbit_r230_c96 bl[96] br[96] wl[230] vdd gnd cell_6t
Xbit_r231_c96 bl[96] br[96] wl[231] vdd gnd cell_6t
Xbit_r232_c96 bl[96] br[96] wl[232] vdd gnd cell_6t
Xbit_r233_c96 bl[96] br[96] wl[233] vdd gnd cell_6t
Xbit_r234_c96 bl[96] br[96] wl[234] vdd gnd cell_6t
Xbit_r235_c96 bl[96] br[96] wl[235] vdd gnd cell_6t
Xbit_r236_c96 bl[96] br[96] wl[236] vdd gnd cell_6t
Xbit_r237_c96 bl[96] br[96] wl[237] vdd gnd cell_6t
Xbit_r238_c96 bl[96] br[96] wl[238] vdd gnd cell_6t
Xbit_r239_c96 bl[96] br[96] wl[239] vdd gnd cell_6t
Xbit_r240_c96 bl[96] br[96] wl[240] vdd gnd cell_6t
Xbit_r241_c96 bl[96] br[96] wl[241] vdd gnd cell_6t
Xbit_r242_c96 bl[96] br[96] wl[242] vdd gnd cell_6t
Xbit_r243_c96 bl[96] br[96] wl[243] vdd gnd cell_6t
Xbit_r244_c96 bl[96] br[96] wl[244] vdd gnd cell_6t
Xbit_r245_c96 bl[96] br[96] wl[245] vdd gnd cell_6t
Xbit_r246_c96 bl[96] br[96] wl[246] vdd gnd cell_6t
Xbit_r247_c96 bl[96] br[96] wl[247] vdd gnd cell_6t
Xbit_r248_c96 bl[96] br[96] wl[248] vdd gnd cell_6t
Xbit_r249_c96 bl[96] br[96] wl[249] vdd gnd cell_6t
Xbit_r250_c96 bl[96] br[96] wl[250] vdd gnd cell_6t
Xbit_r251_c96 bl[96] br[96] wl[251] vdd gnd cell_6t
Xbit_r252_c96 bl[96] br[96] wl[252] vdd gnd cell_6t
Xbit_r253_c96 bl[96] br[96] wl[253] vdd gnd cell_6t
Xbit_r254_c96 bl[96] br[96] wl[254] vdd gnd cell_6t
Xbit_r255_c96 bl[96] br[96] wl[255] vdd gnd cell_6t
Xbit_r0_c97 bl[97] br[97] wl[0] vdd gnd cell_6t
Xbit_r1_c97 bl[97] br[97] wl[1] vdd gnd cell_6t
Xbit_r2_c97 bl[97] br[97] wl[2] vdd gnd cell_6t
Xbit_r3_c97 bl[97] br[97] wl[3] vdd gnd cell_6t
Xbit_r4_c97 bl[97] br[97] wl[4] vdd gnd cell_6t
Xbit_r5_c97 bl[97] br[97] wl[5] vdd gnd cell_6t
Xbit_r6_c97 bl[97] br[97] wl[6] vdd gnd cell_6t
Xbit_r7_c97 bl[97] br[97] wl[7] vdd gnd cell_6t
Xbit_r8_c97 bl[97] br[97] wl[8] vdd gnd cell_6t
Xbit_r9_c97 bl[97] br[97] wl[9] vdd gnd cell_6t
Xbit_r10_c97 bl[97] br[97] wl[10] vdd gnd cell_6t
Xbit_r11_c97 bl[97] br[97] wl[11] vdd gnd cell_6t
Xbit_r12_c97 bl[97] br[97] wl[12] vdd gnd cell_6t
Xbit_r13_c97 bl[97] br[97] wl[13] vdd gnd cell_6t
Xbit_r14_c97 bl[97] br[97] wl[14] vdd gnd cell_6t
Xbit_r15_c97 bl[97] br[97] wl[15] vdd gnd cell_6t
Xbit_r16_c97 bl[97] br[97] wl[16] vdd gnd cell_6t
Xbit_r17_c97 bl[97] br[97] wl[17] vdd gnd cell_6t
Xbit_r18_c97 bl[97] br[97] wl[18] vdd gnd cell_6t
Xbit_r19_c97 bl[97] br[97] wl[19] vdd gnd cell_6t
Xbit_r20_c97 bl[97] br[97] wl[20] vdd gnd cell_6t
Xbit_r21_c97 bl[97] br[97] wl[21] vdd gnd cell_6t
Xbit_r22_c97 bl[97] br[97] wl[22] vdd gnd cell_6t
Xbit_r23_c97 bl[97] br[97] wl[23] vdd gnd cell_6t
Xbit_r24_c97 bl[97] br[97] wl[24] vdd gnd cell_6t
Xbit_r25_c97 bl[97] br[97] wl[25] vdd gnd cell_6t
Xbit_r26_c97 bl[97] br[97] wl[26] vdd gnd cell_6t
Xbit_r27_c97 bl[97] br[97] wl[27] vdd gnd cell_6t
Xbit_r28_c97 bl[97] br[97] wl[28] vdd gnd cell_6t
Xbit_r29_c97 bl[97] br[97] wl[29] vdd gnd cell_6t
Xbit_r30_c97 bl[97] br[97] wl[30] vdd gnd cell_6t
Xbit_r31_c97 bl[97] br[97] wl[31] vdd gnd cell_6t
Xbit_r32_c97 bl[97] br[97] wl[32] vdd gnd cell_6t
Xbit_r33_c97 bl[97] br[97] wl[33] vdd gnd cell_6t
Xbit_r34_c97 bl[97] br[97] wl[34] vdd gnd cell_6t
Xbit_r35_c97 bl[97] br[97] wl[35] vdd gnd cell_6t
Xbit_r36_c97 bl[97] br[97] wl[36] vdd gnd cell_6t
Xbit_r37_c97 bl[97] br[97] wl[37] vdd gnd cell_6t
Xbit_r38_c97 bl[97] br[97] wl[38] vdd gnd cell_6t
Xbit_r39_c97 bl[97] br[97] wl[39] vdd gnd cell_6t
Xbit_r40_c97 bl[97] br[97] wl[40] vdd gnd cell_6t
Xbit_r41_c97 bl[97] br[97] wl[41] vdd gnd cell_6t
Xbit_r42_c97 bl[97] br[97] wl[42] vdd gnd cell_6t
Xbit_r43_c97 bl[97] br[97] wl[43] vdd gnd cell_6t
Xbit_r44_c97 bl[97] br[97] wl[44] vdd gnd cell_6t
Xbit_r45_c97 bl[97] br[97] wl[45] vdd gnd cell_6t
Xbit_r46_c97 bl[97] br[97] wl[46] vdd gnd cell_6t
Xbit_r47_c97 bl[97] br[97] wl[47] vdd gnd cell_6t
Xbit_r48_c97 bl[97] br[97] wl[48] vdd gnd cell_6t
Xbit_r49_c97 bl[97] br[97] wl[49] vdd gnd cell_6t
Xbit_r50_c97 bl[97] br[97] wl[50] vdd gnd cell_6t
Xbit_r51_c97 bl[97] br[97] wl[51] vdd gnd cell_6t
Xbit_r52_c97 bl[97] br[97] wl[52] vdd gnd cell_6t
Xbit_r53_c97 bl[97] br[97] wl[53] vdd gnd cell_6t
Xbit_r54_c97 bl[97] br[97] wl[54] vdd gnd cell_6t
Xbit_r55_c97 bl[97] br[97] wl[55] vdd gnd cell_6t
Xbit_r56_c97 bl[97] br[97] wl[56] vdd gnd cell_6t
Xbit_r57_c97 bl[97] br[97] wl[57] vdd gnd cell_6t
Xbit_r58_c97 bl[97] br[97] wl[58] vdd gnd cell_6t
Xbit_r59_c97 bl[97] br[97] wl[59] vdd gnd cell_6t
Xbit_r60_c97 bl[97] br[97] wl[60] vdd gnd cell_6t
Xbit_r61_c97 bl[97] br[97] wl[61] vdd gnd cell_6t
Xbit_r62_c97 bl[97] br[97] wl[62] vdd gnd cell_6t
Xbit_r63_c97 bl[97] br[97] wl[63] vdd gnd cell_6t
Xbit_r64_c97 bl[97] br[97] wl[64] vdd gnd cell_6t
Xbit_r65_c97 bl[97] br[97] wl[65] vdd gnd cell_6t
Xbit_r66_c97 bl[97] br[97] wl[66] vdd gnd cell_6t
Xbit_r67_c97 bl[97] br[97] wl[67] vdd gnd cell_6t
Xbit_r68_c97 bl[97] br[97] wl[68] vdd gnd cell_6t
Xbit_r69_c97 bl[97] br[97] wl[69] vdd gnd cell_6t
Xbit_r70_c97 bl[97] br[97] wl[70] vdd gnd cell_6t
Xbit_r71_c97 bl[97] br[97] wl[71] vdd gnd cell_6t
Xbit_r72_c97 bl[97] br[97] wl[72] vdd gnd cell_6t
Xbit_r73_c97 bl[97] br[97] wl[73] vdd gnd cell_6t
Xbit_r74_c97 bl[97] br[97] wl[74] vdd gnd cell_6t
Xbit_r75_c97 bl[97] br[97] wl[75] vdd gnd cell_6t
Xbit_r76_c97 bl[97] br[97] wl[76] vdd gnd cell_6t
Xbit_r77_c97 bl[97] br[97] wl[77] vdd gnd cell_6t
Xbit_r78_c97 bl[97] br[97] wl[78] vdd gnd cell_6t
Xbit_r79_c97 bl[97] br[97] wl[79] vdd gnd cell_6t
Xbit_r80_c97 bl[97] br[97] wl[80] vdd gnd cell_6t
Xbit_r81_c97 bl[97] br[97] wl[81] vdd gnd cell_6t
Xbit_r82_c97 bl[97] br[97] wl[82] vdd gnd cell_6t
Xbit_r83_c97 bl[97] br[97] wl[83] vdd gnd cell_6t
Xbit_r84_c97 bl[97] br[97] wl[84] vdd gnd cell_6t
Xbit_r85_c97 bl[97] br[97] wl[85] vdd gnd cell_6t
Xbit_r86_c97 bl[97] br[97] wl[86] vdd gnd cell_6t
Xbit_r87_c97 bl[97] br[97] wl[87] vdd gnd cell_6t
Xbit_r88_c97 bl[97] br[97] wl[88] vdd gnd cell_6t
Xbit_r89_c97 bl[97] br[97] wl[89] vdd gnd cell_6t
Xbit_r90_c97 bl[97] br[97] wl[90] vdd gnd cell_6t
Xbit_r91_c97 bl[97] br[97] wl[91] vdd gnd cell_6t
Xbit_r92_c97 bl[97] br[97] wl[92] vdd gnd cell_6t
Xbit_r93_c97 bl[97] br[97] wl[93] vdd gnd cell_6t
Xbit_r94_c97 bl[97] br[97] wl[94] vdd gnd cell_6t
Xbit_r95_c97 bl[97] br[97] wl[95] vdd gnd cell_6t
Xbit_r96_c97 bl[97] br[97] wl[96] vdd gnd cell_6t
Xbit_r97_c97 bl[97] br[97] wl[97] vdd gnd cell_6t
Xbit_r98_c97 bl[97] br[97] wl[98] vdd gnd cell_6t
Xbit_r99_c97 bl[97] br[97] wl[99] vdd gnd cell_6t
Xbit_r100_c97 bl[97] br[97] wl[100] vdd gnd cell_6t
Xbit_r101_c97 bl[97] br[97] wl[101] vdd gnd cell_6t
Xbit_r102_c97 bl[97] br[97] wl[102] vdd gnd cell_6t
Xbit_r103_c97 bl[97] br[97] wl[103] vdd gnd cell_6t
Xbit_r104_c97 bl[97] br[97] wl[104] vdd gnd cell_6t
Xbit_r105_c97 bl[97] br[97] wl[105] vdd gnd cell_6t
Xbit_r106_c97 bl[97] br[97] wl[106] vdd gnd cell_6t
Xbit_r107_c97 bl[97] br[97] wl[107] vdd gnd cell_6t
Xbit_r108_c97 bl[97] br[97] wl[108] vdd gnd cell_6t
Xbit_r109_c97 bl[97] br[97] wl[109] vdd gnd cell_6t
Xbit_r110_c97 bl[97] br[97] wl[110] vdd gnd cell_6t
Xbit_r111_c97 bl[97] br[97] wl[111] vdd gnd cell_6t
Xbit_r112_c97 bl[97] br[97] wl[112] vdd gnd cell_6t
Xbit_r113_c97 bl[97] br[97] wl[113] vdd gnd cell_6t
Xbit_r114_c97 bl[97] br[97] wl[114] vdd gnd cell_6t
Xbit_r115_c97 bl[97] br[97] wl[115] vdd gnd cell_6t
Xbit_r116_c97 bl[97] br[97] wl[116] vdd gnd cell_6t
Xbit_r117_c97 bl[97] br[97] wl[117] vdd gnd cell_6t
Xbit_r118_c97 bl[97] br[97] wl[118] vdd gnd cell_6t
Xbit_r119_c97 bl[97] br[97] wl[119] vdd gnd cell_6t
Xbit_r120_c97 bl[97] br[97] wl[120] vdd gnd cell_6t
Xbit_r121_c97 bl[97] br[97] wl[121] vdd gnd cell_6t
Xbit_r122_c97 bl[97] br[97] wl[122] vdd gnd cell_6t
Xbit_r123_c97 bl[97] br[97] wl[123] vdd gnd cell_6t
Xbit_r124_c97 bl[97] br[97] wl[124] vdd gnd cell_6t
Xbit_r125_c97 bl[97] br[97] wl[125] vdd gnd cell_6t
Xbit_r126_c97 bl[97] br[97] wl[126] vdd gnd cell_6t
Xbit_r127_c97 bl[97] br[97] wl[127] vdd gnd cell_6t
Xbit_r128_c97 bl[97] br[97] wl[128] vdd gnd cell_6t
Xbit_r129_c97 bl[97] br[97] wl[129] vdd gnd cell_6t
Xbit_r130_c97 bl[97] br[97] wl[130] vdd gnd cell_6t
Xbit_r131_c97 bl[97] br[97] wl[131] vdd gnd cell_6t
Xbit_r132_c97 bl[97] br[97] wl[132] vdd gnd cell_6t
Xbit_r133_c97 bl[97] br[97] wl[133] vdd gnd cell_6t
Xbit_r134_c97 bl[97] br[97] wl[134] vdd gnd cell_6t
Xbit_r135_c97 bl[97] br[97] wl[135] vdd gnd cell_6t
Xbit_r136_c97 bl[97] br[97] wl[136] vdd gnd cell_6t
Xbit_r137_c97 bl[97] br[97] wl[137] vdd gnd cell_6t
Xbit_r138_c97 bl[97] br[97] wl[138] vdd gnd cell_6t
Xbit_r139_c97 bl[97] br[97] wl[139] vdd gnd cell_6t
Xbit_r140_c97 bl[97] br[97] wl[140] vdd gnd cell_6t
Xbit_r141_c97 bl[97] br[97] wl[141] vdd gnd cell_6t
Xbit_r142_c97 bl[97] br[97] wl[142] vdd gnd cell_6t
Xbit_r143_c97 bl[97] br[97] wl[143] vdd gnd cell_6t
Xbit_r144_c97 bl[97] br[97] wl[144] vdd gnd cell_6t
Xbit_r145_c97 bl[97] br[97] wl[145] vdd gnd cell_6t
Xbit_r146_c97 bl[97] br[97] wl[146] vdd gnd cell_6t
Xbit_r147_c97 bl[97] br[97] wl[147] vdd gnd cell_6t
Xbit_r148_c97 bl[97] br[97] wl[148] vdd gnd cell_6t
Xbit_r149_c97 bl[97] br[97] wl[149] vdd gnd cell_6t
Xbit_r150_c97 bl[97] br[97] wl[150] vdd gnd cell_6t
Xbit_r151_c97 bl[97] br[97] wl[151] vdd gnd cell_6t
Xbit_r152_c97 bl[97] br[97] wl[152] vdd gnd cell_6t
Xbit_r153_c97 bl[97] br[97] wl[153] vdd gnd cell_6t
Xbit_r154_c97 bl[97] br[97] wl[154] vdd gnd cell_6t
Xbit_r155_c97 bl[97] br[97] wl[155] vdd gnd cell_6t
Xbit_r156_c97 bl[97] br[97] wl[156] vdd gnd cell_6t
Xbit_r157_c97 bl[97] br[97] wl[157] vdd gnd cell_6t
Xbit_r158_c97 bl[97] br[97] wl[158] vdd gnd cell_6t
Xbit_r159_c97 bl[97] br[97] wl[159] vdd gnd cell_6t
Xbit_r160_c97 bl[97] br[97] wl[160] vdd gnd cell_6t
Xbit_r161_c97 bl[97] br[97] wl[161] vdd gnd cell_6t
Xbit_r162_c97 bl[97] br[97] wl[162] vdd gnd cell_6t
Xbit_r163_c97 bl[97] br[97] wl[163] vdd gnd cell_6t
Xbit_r164_c97 bl[97] br[97] wl[164] vdd gnd cell_6t
Xbit_r165_c97 bl[97] br[97] wl[165] vdd gnd cell_6t
Xbit_r166_c97 bl[97] br[97] wl[166] vdd gnd cell_6t
Xbit_r167_c97 bl[97] br[97] wl[167] vdd gnd cell_6t
Xbit_r168_c97 bl[97] br[97] wl[168] vdd gnd cell_6t
Xbit_r169_c97 bl[97] br[97] wl[169] vdd gnd cell_6t
Xbit_r170_c97 bl[97] br[97] wl[170] vdd gnd cell_6t
Xbit_r171_c97 bl[97] br[97] wl[171] vdd gnd cell_6t
Xbit_r172_c97 bl[97] br[97] wl[172] vdd gnd cell_6t
Xbit_r173_c97 bl[97] br[97] wl[173] vdd gnd cell_6t
Xbit_r174_c97 bl[97] br[97] wl[174] vdd gnd cell_6t
Xbit_r175_c97 bl[97] br[97] wl[175] vdd gnd cell_6t
Xbit_r176_c97 bl[97] br[97] wl[176] vdd gnd cell_6t
Xbit_r177_c97 bl[97] br[97] wl[177] vdd gnd cell_6t
Xbit_r178_c97 bl[97] br[97] wl[178] vdd gnd cell_6t
Xbit_r179_c97 bl[97] br[97] wl[179] vdd gnd cell_6t
Xbit_r180_c97 bl[97] br[97] wl[180] vdd gnd cell_6t
Xbit_r181_c97 bl[97] br[97] wl[181] vdd gnd cell_6t
Xbit_r182_c97 bl[97] br[97] wl[182] vdd gnd cell_6t
Xbit_r183_c97 bl[97] br[97] wl[183] vdd gnd cell_6t
Xbit_r184_c97 bl[97] br[97] wl[184] vdd gnd cell_6t
Xbit_r185_c97 bl[97] br[97] wl[185] vdd gnd cell_6t
Xbit_r186_c97 bl[97] br[97] wl[186] vdd gnd cell_6t
Xbit_r187_c97 bl[97] br[97] wl[187] vdd gnd cell_6t
Xbit_r188_c97 bl[97] br[97] wl[188] vdd gnd cell_6t
Xbit_r189_c97 bl[97] br[97] wl[189] vdd gnd cell_6t
Xbit_r190_c97 bl[97] br[97] wl[190] vdd gnd cell_6t
Xbit_r191_c97 bl[97] br[97] wl[191] vdd gnd cell_6t
Xbit_r192_c97 bl[97] br[97] wl[192] vdd gnd cell_6t
Xbit_r193_c97 bl[97] br[97] wl[193] vdd gnd cell_6t
Xbit_r194_c97 bl[97] br[97] wl[194] vdd gnd cell_6t
Xbit_r195_c97 bl[97] br[97] wl[195] vdd gnd cell_6t
Xbit_r196_c97 bl[97] br[97] wl[196] vdd gnd cell_6t
Xbit_r197_c97 bl[97] br[97] wl[197] vdd gnd cell_6t
Xbit_r198_c97 bl[97] br[97] wl[198] vdd gnd cell_6t
Xbit_r199_c97 bl[97] br[97] wl[199] vdd gnd cell_6t
Xbit_r200_c97 bl[97] br[97] wl[200] vdd gnd cell_6t
Xbit_r201_c97 bl[97] br[97] wl[201] vdd gnd cell_6t
Xbit_r202_c97 bl[97] br[97] wl[202] vdd gnd cell_6t
Xbit_r203_c97 bl[97] br[97] wl[203] vdd gnd cell_6t
Xbit_r204_c97 bl[97] br[97] wl[204] vdd gnd cell_6t
Xbit_r205_c97 bl[97] br[97] wl[205] vdd gnd cell_6t
Xbit_r206_c97 bl[97] br[97] wl[206] vdd gnd cell_6t
Xbit_r207_c97 bl[97] br[97] wl[207] vdd gnd cell_6t
Xbit_r208_c97 bl[97] br[97] wl[208] vdd gnd cell_6t
Xbit_r209_c97 bl[97] br[97] wl[209] vdd gnd cell_6t
Xbit_r210_c97 bl[97] br[97] wl[210] vdd gnd cell_6t
Xbit_r211_c97 bl[97] br[97] wl[211] vdd gnd cell_6t
Xbit_r212_c97 bl[97] br[97] wl[212] vdd gnd cell_6t
Xbit_r213_c97 bl[97] br[97] wl[213] vdd gnd cell_6t
Xbit_r214_c97 bl[97] br[97] wl[214] vdd gnd cell_6t
Xbit_r215_c97 bl[97] br[97] wl[215] vdd gnd cell_6t
Xbit_r216_c97 bl[97] br[97] wl[216] vdd gnd cell_6t
Xbit_r217_c97 bl[97] br[97] wl[217] vdd gnd cell_6t
Xbit_r218_c97 bl[97] br[97] wl[218] vdd gnd cell_6t
Xbit_r219_c97 bl[97] br[97] wl[219] vdd gnd cell_6t
Xbit_r220_c97 bl[97] br[97] wl[220] vdd gnd cell_6t
Xbit_r221_c97 bl[97] br[97] wl[221] vdd gnd cell_6t
Xbit_r222_c97 bl[97] br[97] wl[222] vdd gnd cell_6t
Xbit_r223_c97 bl[97] br[97] wl[223] vdd gnd cell_6t
Xbit_r224_c97 bl[97] br[97] wl[224] vdd gnd cell_6t
Xbit_r225_c97 bl[97] br[97] wl[225] vdd gnd cell_6t
Xbit_r226_c97 bl[97] br[97] wl[226] vdd gnd cell_6t
Xbit_r227_c97 bl[97] br[97] wl[227] vdd gnd cell_6t
Xbit_r228_c97 bl[97] br[97] wl[228] vdd gnd cell_6t
Xbit_r229_c97 bl[97] br[97] wl[229] vdd gnd cell_6t
Xbit_r230_c97 bl[97] br[97] wl[230] vdd gnd cell_6t
Xbit_r231_c97 bl[97] br[97] wl[231] vdd gnd cell_6t
Xbit_r232_c97 bl[97] br[97] wl[232] vdd gnd cell_6t
Xbit_r233_c97 bl[97] br[97] wl[233] vdd gnd cell_6t
Xbit_r234_c97 bl[97] br[97] wl[234] vdd gnd cell_6t
Xbit_r235_c97 bl[97] br[97] wl[235] vdd gnd cell_6t
Xbit_r236_c97 bl[97] br[97] wl[236] vdd gnd cell_6t
Xbit_r237_c97 bl[97] br[97] wl[237] vdd gnd cell_6t
Xbit_r238_c97 bl[97] br[97] wl[238] vdd gnd cell_6t
Xbit_r239_c97 bl[97] br[97] wl[239] vdd gnd cell_6t
Xbit_r240_c97 bl[97] br[97] wl[240] vdd gnd cell_6t
Xbit_r241_c97 bl[97] br[97] wl[241] vdd gnd cell_6t
Xbit_r242_c97 bl[97] br[97] wl[242] vdd gnd cell_6t
Xbit_r243_c97 bl[97] br[97] wl[243] vdd gnd cell_6t
Xbit_r244_c97 bl[97] br[97] wl[244] vdd gnd cell_6t
Xbit_r245_c97 bl[97] br[97] wl[245] vdd gnd cell_6t
Xbit_r246_c97 bl[97] br[97] wl[246] vdd gnd cell_6t
Xbit_r247_c97 bl[97] br[97] wl[247] vdd gnd cell_6t
Xbit_r248_c97 bl[97] br[97] wl[248] vdd gnd cell_6t
Xbit_r249_c97 bl[97] br[97] wl[249] vdd gnd cell_6t
Xbit_r250_c97 bl[97] br[97] wl[250] vdd gnd cell_6t
Xbit_r251_c97 bl[97] br[97] wl[251] vdd gnd cell_6t
Xbit_r252_c97 bl[97] br[97] wl[252] vdd gnd cell_6t
Xbit_r253_c97 bl[97] br[97] wl[253] vdd gnd cell_6t
Xbit_r254_c97 bl[97] br[97] wl[254] vdd gnd cell_6t
Xbit_r255_c97 bl[97] br[97] wl[255] vdd gnd cell_6t
Xbit_r0_c98 bl[98] br[98] wl[0] vdd gnd cell_6t
Xbit_r1_c98 bl[98] br[98] wl[1] vdd gnd cell_6t
Xbit_r2_c98 bl[98] br[98] wl[2] vdd gnd cell_6t
Xbit_r3_c98 bl[98] br[98] wl[3] vdd gnd cell_6t
Xbit_r4_c98 bl[98] br[98] wl[4] vdd gnd cell_6t
Xbit_r5_c98 bl[98] br[98] wl[5] vdd gnd cell_6t
Xbit_r6_c98 bl[98] br[98] wl[6] vdd gnd cell_6t
Xbit_r7_c98 bl[98] br[98] wl[7] vdd gnd cell_6t
Xbit_r8_c98 bl[98] br[98] wl[8] vdd gnd cell_6t
Xbit_r9_c98 bl[98] br[98] wl[9] vdd gnd cell_6t
Xbit_r10_c98 bl[98] br[98] wl[10] vdd gnd cell_6t
Xbit_r11_c98 bl[98] br[98] wl[11] vdd gnd cell_6t
Xbit_r12_c98 bl[98] br[98] wl[12] vdd gnd cell_6t
Xbit_r13_c98 bl[98] br[98] wl[13] vdd gnd cell_6t
Xbit_r14_c98 bl[98] br[98] wl[14] vdd gnd cell_6t
Xbit_r15_c98 bl[98] br[98] wl[15] vdd gnd cell_6t
Xbit_r16_c98 bl[98] br[98] wl[16] vdd gnd cell_6t
Xbit_r17_c98 bl[98] br[98] wl[17] vdd gnd cell_6t
Xbit_r18_c98 bl[98] br[98] wl[18] vdd gnd cell_6t
Xbit_r19_c98 bl[98] br[98] wl[19] vdd gnd cell_6t
Xbit_r20_c98 bl[98] br[98] wl[20] vdd gnd cell_6t
Xbit_r21_c98 bl[98] br[98] wl[21] vdd gnd cell_6t
Xbit_r22_c98 bl[98] br[98] wl[22] vdd gnd cell_6t
Xbit_r23_c98 bl[98] br[98] wl[23] vdd gnd cell_6t
Xbit_r24_c98 bl[98] br[98] wl[24] vdd gnd cell_6t
Xbit_r25_c98 bl[98] br[98] wl[25] vdd gnd cell_6t
Xbit_r26_c98 bl[98] br[98] wl[26] vdd gnd cell_6t
Xbit_r27_c98 bl[98] br[98] wl[27] vdd gnd cell_6t
Xbit_r28_c98 bl[98] br[98] wl[28] vdd gnd cell_6t
Xbit_r29_c98 bl[98] br[98] wl[29] vdd gnd cell_6t
Xbit_r30_c98 bl[98] br[98] wl[30] vdd gnd cell_6t
Xbit_r31_c98 bl[98] br[98] wl[31] vdd gnd cell_6t
Xbit_r32_c98 bl[98] br[98] wl[32] vdd gnd cell_6t
Xbit_r33_c98 bl[98] br[98] wl[33] vdd gnd cell_6t
Xbit_r34_c98 bl[98] br[98] wl[34] vdd gnd cell_6t
Xbit_r35_c98 bl[98] br[98] wl[35] vdd gnd cell_6t
Xbit_r36_c98 bl[98] br[98] wl[36] vdd gnd cell_6t
Xbit_r37_c98 bl[98] br[98] wl[37] vdd gnd cell_6t
Xbit_r38_c98 bl[98] br[98] wl[38] vdd gnd cell_6t
Xbit_r39_c98 bl[98] br[98] wl[39] vdd gnd cell_6t
Xbit_r40_c98 bl[98] br[98] wl[40] vdd gnd cell_6t
Xbit_r41_c98 bl[98] br[98] wl[41] vdd gnd cell_6t
Xbit_r42_c98 bl[98] br[98] wl[42] vdd gnd cell_6t
Xbit_r43_c98 bl[98] br[98] wl[43] vdd gnd cell_6t
Xbit_r44_c98 bl[98] br[98] wl[44] vdd gnd cell_6t
Xbit_r45_c98 bl[98] br[98] wl[45] vdd gnd cell_6t
Xbit_r46_c98 bl[98] br[98] wl[46] vdd gnd cell_6t
Xbit_r47_c98 bl[98] br[98] wl[47] vdd gnd cell_6t
Xbit_r48_c98 bl[98] br[98] wl[48] vdd gnd cell_6t
Xbit_r49_c98 bl[98] br[98] wl[49] vdd gnd cell_6t
Xbit_r50_c98 bl[98] br[98] wl[50] vdd gnd cell_6t
Xbit_r51_c98 bl[98] br[98] wl[51] vdd gnd cell_6t
Xbit_r52_c98 bl[98] br[98] wl[52] vdd gnd cell_6t
Xbit_r53_c98 bl[98] br[98] wl[53] vdd gnd cell_6t
Xbit_r54_c98 bl[98] br[98] wl[54] vdd gnd cell_6t
Xbit_r55_c98 bl[98] br[98] wl[55] vdd gnd cell_6t
Xbit_r56_c98 bl[98] br[98] wl[56] vdd gnd cell_6t
Xbit_r57_c98 bl[98] br[98] wl[57] vdd gnd cell_6t
Xbit_r58_c98 bl[98] br[98] wl[58] vdd gnd cell_6t
Xbit_r59_c98 bl[98] br[98] wl[59] vdd gnd cell_6t
Xbit_r60_c98 bl[98] br[98] wl[60] vdd gnd cell_6t
Xbit_r61_c98 bl[98] br[98] wl[61] vdd gnd cell_6t
Xbit_r62_c98 bl[98] br[98] wl[62] vdd gnd cell_6t
Xbit_r63_c98 bl[98] br[98] wl[63] vdd gnd cell_6t
Xbit_r64_c98 bl[98] br[98] wl[64] vdd gnd cell_6t
Xbit_r65_c98 bl[98] br[98] wl[65] vdd gnd cell_6t
Xbit_r66_c98 bl[98] br[98] wl[66] vdd gnd cell_6t
Xbit_r67_c98 bl[98] br[98] wl[67] vdd gnd cell_6t
Xbit_r68_c98 bl[98] br[98] wl[68] vdd gnd cell_6t
Xbit_r69_c98 bl[98] br[98] wl[69] vdd gnd cell_6t
Xbit_r70_c98 bl[98] br[98] wl[70] vdd gnd cell_6t
Xbit_r71_c98 bl[98] br[98] wl[71] vdd gnd cell_6t
Xbit_r72_c98 bl[98] br[98] wl[72] vdd gnd cell_6t
Xbit_r73_c98 bl[98] br[98] wl[73] vdd gnd cell_6t
Xbit_r74_c98 bl[98] br[98] wl[74] vdd gnd cell_6t
Xbit_r75_c98 bl[98] br[98] wl[75] vdd gnd cell_6t
Xbit_r76_c98 bl[98] br[98] wl[76] vdd gnd cell_6t
Xbit_r77_c98 bl[98] br[98] wl[77] vdd gnd cell_6t
Xbit_r78_c98 bl[98] br[98] wl[78] vdd gnd cell_6t
Xbit_r79_c98 bl[98] br[98] wl[79] vdd gnd cell_6t
Xbit_r80_c98 bl[98] br[98] wl[80] vdd gnd cell_6t
Xbit_r81_c98 bl[98] br[98] wl[81] vdd gnd cell_6t
Xbit_r82_c98 bl[98] br[98] wl[82] vdd gnd cell_6t
Xbit_r83_c98 bl[98] br[98] wl[83] vdd gnd cell_6t
Xbit_r84_c98 bl[98] br[98] wl[84] vdd gnd cell_6t
Xbit_r85_c98 bl[98] br[98] wl[85] vdd gnd cell_6t
Xbit_r86_c98 bl[98] br[98] wl[86] vdd gnd cell_6t
Xbit_r87_c98 bl[98] br[98] wl[87] vdd gnd cell_6t
Xbit_r88_c98 bl[98] br[98] wl[88] vdd gnd cell_6t
Xbit_r89_c98 bl[98] br[98] wl[89] vdd gnd cell_6t
Xbit_r90_c98 bl[98] br[98] wl[90] vdd gnd cell_6t
Xbit_r91_c98 bl[98] br[98] wl[91] vdd gnd cell_6t
Xbit_r92_c98 bl[98] br[98] wl[92] vdd gnd cell_6t
Xbit_r93_c98 bl[98] br[98] wl[93] vdd gnd cell_6t
Xbit_r94_c98 bl[98] br[98] wl[94] vdd gnd cell_6t
Xbit_r95_c98 bl[98] br[98] wl[95] vdd gnd cell_6t
Xbit_r96_c98 bl[98] br[98] wl[96] vdd gnd cell_6t
Xbit_r97_c98 bl[98] br[98] wl[97] vdd gnd cell_6t
Xbit_r98_c98 bl[98] br[98] wl[98] vdd gnd cell_6t
Xbit_r99_c98 bl[98] br[98] wl[99] vdd gnd cell_6t
Xbit_r100_c98 bl[98] br[98] wl[100] vdd gnd cell_6t
Xbit_r101_c98 bl[98] br[98] wl[101] vdd gnd cell_6t
Xbit_r102_c98 bl[98] br[98] wl[102] vdd gnd cell_6t
Xbit_r103_c98 bl[98] br[98] wl[103] vdd gnd cell_6t
Xbit_r104_c98 bl[98] br[98] wl[104] vdd gnd cell_6t
Xbit_r105_c98 bl[98] br[98] wl[105] vdd gnd cell_6t
Xbit_r106_c98 bl[98] br[98] wl[106] vdd gnd cell_6t
Xbit_r107_c98 bl[98] br[98] wl[107] vdd gnd cell_6t
Xbit_r108_c98 bl[98] br[98] wl[108] vdd gnd cell_6t
Xbit_r109_c98 bl[98] br[98] wl[109] vdd gnd cell_6t
Xbit_r110_c98 bl[98] br[98] wl[110] vdd gnd cell_6t
Xbit_r111_c98 bl[98] br[98] wl[111] vdd gnd cell_6t
Xbit_r112_c98 bl[98] br[98] wl[112] vdd gnd cell_6t
Xbit_r113_c98 bl[98] br[98] wl[113] vdd gnd cell_6t
Xbit_r114_c98 bl[98] br[98] wl[114] vdd gnd cell_6t
Xbit_r115_c98 bl[98] br[98] wl[115] vdd gnd cell_6t
Xbit_r116_c98 bl[98] br[98] wl[116] vdd gnd cell_6t
Xbit_r117_c98 bl[98] br[98] wl[117] vdd gnd cell_6t
Xbit_r118_c98 bl[98] br[98] wl[118] vdd gnd cell_6t
Xbit_r119_c98 bl[98] br[98] wl[119] vdd gnd cell_6t
Xbit_r120_c98 bl[98] br[98] wl[120] vdd gnd cell_6t
Xbit_r121_c98 bl[98] br[98] wl[121] vdd gnd cell_6t
Xbit_r122_c98 bl[98] br[98] wl[122] vdd gnd cell_6t
Xbit_r123_c98 bl[98] br[98] wl[123] vdd gnd cell_6t
Xbit_r124_c98 bl[98] br[98] wl[124] vdd gnd cell_6t
Xbit_r125_c98 bl[98] br[98] wl[125] vdd gnd cell_6t
Xbit_r126_c98 bl[98] br[98] wl[126] vdd gnd cell_6t
Xbit_r127_c98 bl[98] br[98] wl[127] vdd gnd cell_6t
Xbit_r128_c98 bl[98] br[98] wl[128] vdd gnd cell_6t
Xbit_r129_c98 bl[98] br[98] wl[129] vdd gnd cell_6t
Xbit_r130_c98 bl[98] br[98] wl[130] vdd gnd cell_6t
Xbit_r131_c98 bl[98] br[98] wl[131] vdd gnd cell_6t
Xbit_r132_c98 bl[98] br[98] wl[132] vdd gnd cell_6t
Xbit_r133_c98 bl[98] br[98] wl[133] vdd gnd cell_6t
Xbit_r134_c98 bl[98] br[98] wl[134] vdd gnd cell_6t
Xbit_r135_c98 bl[98] br[98] wl[135] vdd gnd cell_6t
Xbit_r136_c98 bl[98] br[98] wl[136] vdd gnd cell_6t
Xbit_r137_c98 bl[98] br[98] wl[137] vdd gnd cell_6t
Xbit_r138_c98 bl[98] br[98] wl[138] vdd gnd cell_6t
Xbit_r139_c98 bl[98] br[98] wl[139] vdd gnd cell_6t
Xbit_r140_c98 bl[98] br[98] wl[140] vdd gnd cell_6t
Xbit_r141_c98 bl[98] br[98] wl[141] vdd gnd cell_6t
Xbit_r142_c98 bl[98] br[98] wl[142] vdd gnd cell_6t
Xbit_r143_c98 bl[98] br[98] wl[143] vdd gnd cell_6t
Xbit_r144_c98 bl[98] br[98] wl[144] vdd gnd cell_6t
Xbit_r145_c98 bl[98] br[98] wl[145] vdd gnd cell_6t
Xbit_r146_c98 bl[98] br[98] wl[146] vdd gnd cell_6t
Xbit_r147_c98 bl[98] br[98] wl[147] vdd gnd cell_6t
Xbit_r148_c98 bl[98] br[98] wl[148] vdd gnd cell_6t
Xbit_r149_c98 bl[98] br[98] wl[149] vdd gnd cell_6t
Xbit_r150_c98 bl[98] br[98] wl[150] vdd gnd cell_6t
Xbit_r151_c98 bl[98] br[98] wl[151] vdd gnd cell_6t
Xbit_r152_c98 bl[98] br[98] wl[152] vdd gnd cell_6t
Xbit_r153_c98 bl[98] br[98] wl[153] vdd gnd cell_6t
Xbit_r154_c98 bl[98] br[98] wl[154] vdd gnd cell_6t
Xbit_r155_c98 bl[98] br[98] wl[155] vdd gnd cell_6t
Xbit_r156_c98 bl[98] br[98] wl[156] vdd gnd cell_6t
Xbit_r157_c98 bl[98] br[98] wl[157] vdd gnd cell_6t
Xbit_r158_c98 bl[98] br[98] wl[158] vdd gnd cell_6t
Xbit_r159_c98 bl[98] br[98] wl[159] vdd gnd cell_6t
Xbit_r160_c98 bl[98] br[98] wl[160] vdd gnd cell_6t
Xbit_r161_c98 bl[98] br[98] wl[161] vdd gnd cell_6t
Xbit_r162_c98 bl[98] br[98] wl[162] vdd gnd cell_6t
Xbit_r163_c98 bl[98] br[98] wl[163] vdd gnd cell_6t
Xbit_r164_c98 bl[98] br[98] wl[164] vdd gnd cell_6t
Xbit_r165_c98 bl[98] br[98] wl[165] vdd gnd cell_6t
Xbit_r166_c98 bl[98] br[98] wl[166] vdd gnd cell_6t
Xbit_r167_c98 bl[98] br[98] wl[167] vdd gnd cell_6t
Xbit_r168_c98 bl[98] br[98] wl[168] vdd gnd cell_6t
Xbit_r169_c98 bl[98] br[98] wl[169] vdd gnd cell_6t
Xbit_r170_c98 bl[98] br[98] wl[170] vdd gnd cell_6t
Xbit_r171_c98 bl[98] br[98] wl[171] vdd gnd cell_6t
Xbit_r172_c98 bl[98] br[98] wl[172] vdd gnd cell_6t
Xbit_r173_c98 bl[98] br[98] wl[173] vdd gnd cell_6t
Xbit_r174_c98 bl[98] br[98] wl[174] vdd gnd cell_6t
Xbit_r175_c98 bl[98] br[98] wl[175] vdd gnd cell_6t
Xbit_r176_c98 bl[98] br[98] wl[176] vdd gnd cell_6t
Xbit_r177_c98 bl[98] br[98] wl[177] vdd gnd cell_6t
Xbit_r178_c98 bl[98] br[98] wl[178] vdd gnd cell_6t
Xbit_r179_c98 bl[98] br[98] wl[179] vdd gnd cell_6t
Xbit_r180_c98 bl[98] br[98] wl[180] vdd gnd cell_6t
Xbit_r181_c98 bl[98] br[98] wl[181] vdd gnd cell_6t
Xbit_r182_c98 bl[98] br[98] wl[182] vdd gnd cell_6t
Xbit_r183_c98 bl[98] br[98] wl[183] vdd gnd cell_6t
Xbit_r184_c98 bl[98] br[98] wl[184] vdd gnd cell_6t
Xbit_r185_c98 bl[98] br[98] wl[185] vdd gnd cell_6t
Xbit_r186_c98 bl[98] br[98] wl[186] vdd gnd cell_6t
Xbit_r187_c98 bl[98] br[98] wl[187] vdd gnd cell_6t
Xbit_r188_c98 bl[98] br[98] wl[188] vdd gnd cell_6t
Xbit_r189_c98 bl[98] br[98] wl[189] vdd gnd cell_6t
Xbit_r190_c98 bl[98] br[98] wl[190] vdd gnd cell_6t
Xbit_r191_c98 bl[98] br[98] wl[191] vdd gnd cell_6t
Xbit_r192_c98 bl[98] br[98] wl[192] vdd gnd cell_6t
Xbit_r193_c98 bl[98] br[98] wl[193] vdd gnd cell_6t
Xbit_r194_c98 bl[98] br[98] wl[194] vdd gnd cell_6t
Xbit_r195_c98 bl[98] br[98] wl[195] vdd gnd cell_6t
Xbit_r196_c98 bl[98] br[98] wl[196] vdd gnd cell_6t
Xbit_r197_c98 bl[98] br[98] wl[197] vdd gnd cell_6t
Xbit_r198_c98 bl[98] br[98] wl[198] vdd gnd cell_6t
Xbit_r199_c98 bl[98] br[98] wl[199] vdd gnd cell_6t
Xbit_r200_c98 bl[98] br[98] wl[200] vdd gnd cell_6t
Xbit_r201_c98 bl[98] br[98] wl[201] vdd gnd cell_6t
Xbit_r202_c98 bl[98] br[98] wl[202] vdd gnd cell_6t
Xbit_r203_c98 bl[98] br[98] wl[203] vdd gnd cell_6t
Xbit_r204_c98 bl[98] br[98] wl[204] vdd gnd cell_6t
Xbit_r205_c98 bl[98] br[98] wl[205] vdd gnd cell_6t
Xbit_r206_c98 bl[98] br[98] wl[206] vdd gnd cell_6t
Xbit_r207_c98 bl[98] br[98] wl[207] vdd gnd cell_6t
Xbit_r208_c98 bl[98] br[98] wl[208] vdd gnd cell_6t
Xbit_r209_c98 bl[98] br[98] wl[209] vdd gnd cell_6t
Xbit_r210_c98 bl[98] br[98] wl[210] vdd gnd cell_6t
Xbit_r211_c98 bl[98] br[98] wl[211] vdd gnd cell_6t
Xbit_r212_c98 bl[98] br[98] wl[212] vdd gnd cell_6t
Xbit_r213_c98 bl[98] br[98] wl[213] vdd gnd cell_6t
Xbit_r214_c98 bl[98] br[98] wl[214] vdd gnd cell_6t
Xbit_r215_c98 bl[98] br[98] wl[215] vdd gnd cell_6t
Xbit_r216_c98 bl[98] br[98] wl[216] vdd gnd cell_6t
Xbit_r217_c98 bl[98] br[98] wl[217] vdd gnd cell_6t
Xbit_r218_c98 bl[98] br[98] wl[218] vdd gnd cell_6t
Xbit_r219_c98 bl[98] br[98] wl[219] vdd gnd cell_6t
Xbit_r220_c98 bl[98] br[98] wl[220] vdd gnd cell_6t
Xbit_r221_c98 bl[98] br[98] wl[221] vdd gnd cell_6t
Xbit_r222_c98 bl[98] br[98] wl[222] vdd gnd cell_6t
Xbit_r223_c98 bl[98] br[98] wl[223] vdd gnd cell_6t
Xbit_r224_c98 bl[98] br[98] wl[224] vdd gnd cell_6t
Xbit_r225_c98 bl[98] br[98] wl[225] vdd gnd cell_6t
Xbit_r226_c98 bl[98] br[98] wl[226] vdd gnd cell_6t
Xbit_r227_c98 bl[98] br[98] wl[227] vdd gnd cell_6t
Xbit_r228_c98 bl[98] br[98] wl[228] vdd gnd cell_6t
Xbit_r229_c98 bl[98] br[98] wl[229] vdd gnd cell_6t
Xbit_r230_c98 bl[98] br[98] wl[230] vdd gnd cell_6t
Xbit_r231_c98 bl[98] br[98] wl[231] vdd gnd cell_6t
Xbit_r232_c98 bl[98] br[98] wl[232] vdd gnd cell_6t
Xbit_r233_c98 bl[98] br[98] wl[233] vdd gnd cell_6t
Xbit_r234_c98 bl[98] br[98] wl[234] vdd gnd cell_6t
Xbit_r235_c98 bl[98] br[98] wl[235] vdd gnd cell_6t
Xbit_r236_c98 bl[98] br[98] wl[236] vdd gnd cell_6t
Xbit_r237_c98 bl[98] br[98] wl[237] vdd gnd cell_6t
Xbit_r238_c98 bl[98] br[98] wl[238] vdd gnd cell_6t
Xbit_r239_c98 bl[98] br[98] wl[239] vdd gnd cell_6t
Xbit_r240_c98 bl[98] br[98] wl[240] vdd gnd cell_6t
Xbit_r241_c98 bl[98] br[98] wl[241] vdd gnd cell_6t
Xbit_r242_c98 bl[98] br[98] wl[242] vdd gnd cell_6t
Xbit_r243_c98 bl[98] br[98] wl[243] vdd gnd cell_6t
Xbit_r244_c98 bl[98] br[98] wl[244] vdd gnd cell_6t
Xbit_r245_c98 bl[98] br[98] wl[245] vdd gnd cell_6t
Xbit_r246_c98 bl[98] br[98] wl[246] vdd gnd cell_6t
Xbit_r247_c98 bl[98] br[98] wl[247] vdd gnd cell_6t
Xbit_r248_c98 bl[98] br[98] wl[248] vdd gnd cell_6t
Xbit_r249_c98 bl[98] br[98] wl[249] vdd gnd cell_6t
Xbit_r250_c98 bl[98] br[98] wl[250] vdd gnd cell_6t
Xbit_r251_c98 bl[98] br[98] wl[251] vdd gnd cell_6t
Xbit_r252_c98 bl[98] br[98] wl[252] vdd gnd cell_6t
Xbit_r253_c98 bl[98] br[98] wl[253] vdd gnd cell_6t
Xbit_r254_c98 bl[98] br[98] wl[254] vdd gnd cell_6t
Xbit_r255_c98 bl[98] br[98] wl[255] vdd gnd cell_6t
Xbit_r0_c99 bl[99] br[99] wl[0] vdd gnd cell_6t
Xbit_r1_c99 bl[99] br[99] wl[1] vdd gnd cell_6t
Xbit_r2_c99 bl[99] br[99] wl[2] vdd gnd cell_6t
Xbit_r3_c99 bl[99] br[99] wl[3] vdd gnd cell_6t
Xbit_r4_c99 bl[99] br[99] wl[4] vdd gnd cell_6t
Xbit_r5_c99 bl[99] br[99] wl[5] vdd gnd cell_6t
Xbit_r6_c99 bl[99] br[99] wl[6] vdd gnd cell_6t
Xbit_r7_c99 bl[99] br[99] wl[7] vdd gnd cell_6t
Xbit_r8_c99 bl[99] br[99] wl[8] vdd gnd cell_6t
Xbit_r9_c99 bl[99] br[99] wl[9] vdd gnd cell_6t
Xbit_r10_c99 bl[99] br[99] wl[10] vdd gnd cell_6t
Xbit_r11_c99 bl[99] br[99] wl[11] vdd gnd cell_6t
Xbit_r12_c99 bl[99] br[99] wl[12] vdd gnd cell_6t
Xbit_r13_c99 bl[99] br[99] wl[13] vdd gnd cell_6t
Xbit_r14_c99 bl[99] br[99] wl[14] vdd gnd cell_6t
Xbit_r15_c99 bl[99] br[99] wl[15] vdd gnd cell_6t
Xbit_r16_c99 bl[99] br[99] wl[16] vdd gnd cell_6t
Xbit_r17_c99 bl[99] br[99] wl[17] vdd gnd cell_6t
Xbit_r18_c99 bl[99] br[99] wl[18] vdd gnd cell_6t
Xbit_r19_c99 bl[99] br[99] wl[19] vdd gnd cell_6t
Xbit_r20_c99 bl[99] br[99] wl[20] vdd gnd cell_6t
Xbit_r21_c99 bl[99] br[99] wl[21] vdd gnd cell_6t
Xbit_r22_c99 bl[99] br[99] wl[22] vdd gnd cell_6t
Xbit_r23_c99 bl[99] br[99] wl[23] vdd gnd cell_6t
Xbit_r24_c99 bl[99] br[99] wl[24] vdd gnd cell_6t
Xbit_r25_c99 bl[99] br[99] wl[25] vdd gnd cell_6t
Xbit_r26_c99 bl[99] br[99] wl[26] vdd gnd cell_6t
Xbit_r27_c99 bl[99] br[99] wl[27] vdd gnd cell_6t
Xbit_r28_c99 bl[99] br[99] wl[28] vdd gnd cell_6t
Xbit_r29_c99 bl[99] br[99] wl[29] vdd gnd cell_6t
Xbit_r30_c99 bl[99] br[99] wl[30] vdd gnd cell_6t
Xbit_r31_c99 bl[99] br[99] wl[31] vdd gnd cell_6t
Xbit_r32_c99 bl[99] br[99] wl[32] vdd gnd cell_6t
Xbit_r33_c99 bl[99] br[99] wl[33] vdd gnd cell_6t
Xbit_r34_c99 bl[99] br[99] wl[34] vdd gnd cell_6t
Xbit_r35_c99 bl[99] br[99] wl[35] vdd gnd cell_6t
Xbit_r36_c99 bl[99] br[99] wl[36] vdd gnd cell_6t
Xbit_r37_c99 bl[99] br[99] wl[37] vdd gnd cell_6t
Xbit_r38_c99 bl[99] br[99] wl[38] vdd gnd cell_6t
Xbit_r39_c99 bl[99] br[99] wl[39] vdd gnd cell_6t
Xbit_r40_c99 bl[99] br[99] wl[40] vdd gnd cell_6t
Xbit_r41_c99 bl[99] br[99] wl[41] vdd gnd cell_6t
Xbit_r42_c99 bl[99] br[99] wl[42] vdd gnd cell_6t
Xbit_r43_c99 bl[99] br[99] wl[43] vdd gnd cell_6t
Xbit_r44_c99 bl[99] br[99] wl[44] vdd gnd cell_6t
Xbit_r45_c99 bl[99] br[99] wl[45] vdd gnd cell_6t
Xbit_r46_c99 bl[99] br[99] wl[46] vdd gnd cell_6t
Xbit_r47_c99 bl[99] br[99] wl[47] vdd gnd cell_6t
Xbit_r48_c99 bl[99] br[99] wl[48] vdd gnd cell_6t
Xbit_r49_c99 bl[99] br[99] wl[49] vdd gnd cell_6t
Xbit_r50_c99 bl[99] br[99] wl[50] vdd gnd cell_6t
Xbit_r51_c99 bl[99] br[99] wl[51] vdd gnd cell_6t
Xbit_r52_c99 bl[99] br[99] wl[52] vdd gnd cell_6t
Xbit_r53_c99 bl[99] br[99] wl[53] vdd gnd cell_6t
Xbit_r54_c99 bl[99] br[99] wl[54] vdd gnd cell_6t
Xbit_r55_c99 bl[99] br[99] wl[55] vdd gnd cell_6t
Xbit_r56_c99 bl[99] br[99] wl[56] vdd gnd cell_6t
Xbit_r57_c99 bl[99] br[99] wl[57] vdd gnd cell_6t
Xbit_r58_c99 bl[99] br[99] wl[58] vdd gnd cell_6t
Xbit_r59_c99 bl[99] br[99] wl[59] vdd gnd cell_6t
Xbit_r60_c99 bl[99] br[99] wl[60] vdd gnd cell_6t
Xbit_r61_c99 bl[99] br[99] wl[61] vdd gnd cell_6t
Xbit_r62_c99 bl[99] br[99] wl[62] vdd gnd cell_6t
Xbit_r63_c99 bl[99] br[99] wl[63] vdd gnd cell_6t
Xbit_r64_c99 bl[99] br[99] wl[64] vdd gnd cell_6t
Xbit_r65_c99 bl[99] br[99] wl[65] vdd gnd cell_6t
Xbit_r66_c99 bl[99] br[99] wl[66] vdd gnd cell_6t
Xbit_r67_c99 bl[99] br[99] wl[67] vdd gnd cell_6t
Xbit_r68_c99 bl[99] br[99] wl[68] vdd gnd cell_6t
Xbit_r69_c99 bl[99] br[99] wl[69] vdd gnd cell_6t
Xbit_r70_c99 bl[99] br[99] wl[70] vdd gnd cell_6t
Xbit_r71_c99 bl[99] br[99] wl[71] vdd gnd cell_6t
Xbit_r72_c99 bl[99] br[99] wl[72] vdd gnd cell_6t
Xbit_r73_c99 bl[99] br[99] wl[73] vdd gnd cell_6t
Xbit_r74_c99 bl[99] br[99] wl[74] vdd gnd cell_6t
Xbit_r75_c99 bl[99] br[99] wl[75] vdd gnd cell_6t
Xbit_r76_c99 bl[99] br[99] wl[76] vdd gnd cell_6t
Xbit_r77_c99 bl[99] br[99] wl[77] vdd gnd cell_6t
Xbit_r78_c99 bl[99] br[99] wl[78] vdd gnd cell_6t
Xbit_r79_c99 bl[99] br[99] wl[79] vdd gnd cell_6t
Xbit_r80_c99 bl[99] br[99] wl[80] vdd gnd cell_6t
Xbit_r81_c99 bl[99] br[99] wl[81] vdd gnd cell_6t
Xbit_r82_c99 bl[99] br[99] wl[82] vdd gnd cell_6t
Xbit_r83_c99 bl[99] br[99] wl[83] vdd gnd cell_6t
Xbit_r84_c99 bl[99] br[99] wl[84] vdd gnd cell_6t
Xbit_r85_c99 bl[99] br[99] wl[85] vdd gnd cell_6t
Xbit_r86_c99 bl[99] br[99] wl[86] vdd gnd cell_6t
Xbit_r87_c99 bl[99] br[99] wl[87] vdd gnd cell_6t
Xbit_r88_c99 bl[99] br[99] wl[88] vdd gnd cell_6t
Xbit_r89_c99 bl[99] br[99] wl[89] vdd gnd cell_6t
Xbit_r90_c99 bl[99] br[99] wl[90] vdd gnd cell_6t
Xbit_r91_c99 bl[99] br[99] wl[91] vdd gnd cell_6t
Xbit_r92_c99 bl[99] br[99] wl[92] vdd gnd cell_6t
Xbit_r93_c99 bl[99] br[99] wl[93] vdd gnd cell_6t
Xbit_r94_c99 bl[99] br[99] wl[94] vdd gnd cell_6t
Xbit_r95_c99 bl[99] br[99] wl[95] vdd gnd cell_6t
Xbit_r96_c99 bl[99] br[99] wl[96] vdd gnd cell_6t
Xbit_r97_c99 bl[99] br[99] wl[97] vdd gnd cell_6t
Xbit_r98_c99 bl[99] br[99] wl[98] vdd gnd cell_6t
Xbit_r99_c99 bl[99] br[99] wl[99] vdd gnd cell_6t
Xbit_r100_c99 bl[99] br[99] wl[100] vdd gnd cell_6t
Xbit_r101_c99 bl[99] br[99] wl[101] vdd gnd cell_6t
Xbit_r102_c99 bl[99] br[99] wl[102] vdd gnd cell_6t
Xbit_r103_c99 bl[99] br[99] wl[103] vdd gnd cell_6t
Xbit_r104_c99 bl[99] br[99] wl[104] vdd gnd cell_6t
Xbit_r105_c99 bl[99] br[99] wl[105] vdd gnd cell_6t
Xbit_r106_c99 bl[99] br[99] wl[106] vdd gnd cell_6t
Xbit_r107_c99 bl[99] br[99] wl[107] vdd gnd cell_6t
Xbit_r108_c99 bl[99] br[99] wl[108] vdd gnd cell_6t
Xbit_r109_c99 bl[99] br[99] wl[109] vdd gnd cell_6t
Xbit_r110_c99 bl[99] br[99] wl[110] vdd gnd cell_6t
Xbit_r111_c99 bl[99] br[99] wl[111] vdd gnd cell_6t
Xbit_r112_c99 bl[99] br[99] wl[112] vdd gnd cell_6t
Xbit_r113_c99 bl[99] br[99] wl[113] vdd gnd cell_6t
Xbit_r114_c99 bl[99] br[99] wl[114] vdd gnd cell_6t
Xbit_r115_c99 bl[99] br[99] wl[115] vdd gnd cell_6t
Xbit_r116_c99 bl[99] br[99] wl[116] vdd gnd cell_6t
Xbit_r117_c99 bl[99] br[99] wl[117] vdd gnd cell_6t
Xbit_r118_c99 bl[99] br[99] wl[118] vdd gnd cell_6t
Xbit_r119_c99 bl[99] br[99] wl[119] vdd gnd cell_6t
Xbit_r120_c99 bl[99] br[99] wl[120] vdd gnd cell_6t
Xbit_r121_c99 bl[99] br[99] wl[121] vdd gnd cell_6t
Xbit_r122_c99 bl[99] br[99] wl[122] vdd gnd cell_6t
Xbit_r123_c99 bl[99] br[99] wl[123] vdd gnd cell_6t
Xbit_r124_c99 bl[99] br[99] wl[124] vdd gnd cell_6t
Xbit_r125_c99 bl[99] br[99] wl[125] vdd gnd cell_6t
Xbit_r126_c99 bl[99] br[99] wl[126] vdd gnd cell_6t
Xbit_r127_c99 bl[99] br[99] wl[127] vdd gnd cell_6t
Xbit_r128_c99 bl[99] br[99] wl[128] vdd gnd cell_6t
Xbit_r129_c99 bl[99] br[99] wl[129] vdd gnd cell_6t
Xbit_r130_c99 bl[99] br[99] wl[130] vdd gnd cell_6t
Xbit_r131_c99 bl[99] br[99] wl[131] vdd gnd cell_6t
Xbit_r132_c99 bl[99] br[99] wl[132] vdd gnd cell_6t
Xbit_r133_c99 bl[99] br[99] wl[133] vdd gnd cell_6t
Xbit_r134_c99 bl[99] br[99] wl[134] vdd gnd cell_6t
Xbit_r135_c99 bl[99] br[99] wl[135] vdd gnd cell_6t
Xbit_r136_c99 bl[99] br[99] wl[136] vdd gnd cell_6t
Xbit_r137_c99 bl[99] br[99] wl[137] vdd gnd cell_6t
Xbit_r138_c99 bl[99] br[99] wl[138] vdd gnd cell_6t
Xbit_r139_c99 bl[99] br[99] wl[139] vdd gnd cell_6t
Xbit_r140_c99 bl[99] br[99] wl[140] vdd gnd cell_6t
Xbit_r141_c99 bl[99] br[99] wl[141] vdd gnd cell_6t
Xbit_r142_c99 bl[99] br[99] wl[142] vdd gnd cell_6t
Xbit_r143_c99 bl[99] br[99] wl[143] vdd gnd cell_6t
Xbit_r144_c99 bl[99] br[99] wl[144] vdd gnd cell_6t
Xbit_r145_c99 bl[99] br[99] wl[145] vdd gnd cell_6t
Xbit_r146_c99 bl[99] br[99] wl[146] vdd gnd cell_6t
Xbit_r147_c99 bl[99] br[99] wl[147] vdd gnd cell_6t
Xbit_r148_c99 bl[99] br[99] wl[148] vdd gnd cell_6t
Xbit_r149_c99 bl[99] br[99] wl[149] vdd gnd cell_6t
Xbit_r150_c99 bl[99] br[99] wl[150] vdd gnd cell_6t
Xbit_r151_c99 bl[99] br[99] wl[151] vdd gnd cell_6t
Xbit_r152_c99 bl[99] br[99] wl[152] vdd gnd cell_6t
Xbit_r153_c99 bl[99] br[99] wl[153] vdd gnd cell_6t
Xbit_r154_c99 bl[99] br[99] wl[154] vdd gnd cell_6t
Xbit_r155_c99 bl[99] br[99] wl[155] vdd gnd cell_6t
Xbit_r156_c99 bl[99] br[99] wl[156] vdd gnd cell_6t
Xbit_r157_c99 bl[99] br[99] wl[157] vdd gnd cell_6t
Xbit_r158_c99 bl[99] br[99] wl[158] vdd gnd cell_6t
Xbit_r159_c99 bl[99] br[99] wl[159] vdd gnd cell_6t
Xbit_r160_c99 bl[99] br[99] wl[160] vdd gnd cell_6t
Xbit_r161_c99 bl[99] br[99] wl[161] vdd gnd cell_6t
Xbit_r162_c99 bl[99] br[99] wl[162] vdd gnd cell_6t
Xbit_r163_c99 bl[99] br[99] wl[163] vdd gnd cell_6t
Xbit_r164_c99 bl[99] br[99] wl[164] vdd gnd cell_6t
Xbit_r165_c99 bl[99] br[99] wl[165] vdd gnd cell_6t
Xbit_r166_c99 bl[99] br[99] wl[166] vdd gnd cell_6t
Xbit_r167_c99 bl[99] br[99] wl[167] vdd gnd cell_6t
Xbit_r168_c99 bl[99] br[99] wl[168] vdd gnd cell_6t
Xbit_r169_c99 bl[99] br[99] wl[169] vdd gnd cell_6t
Xbit_r170_c99 bl[99] br[99] wl[170] vdd gnd cell_6t
Xbit_r171_c99 bl[99] br[99] wl[171] vdd gnd cell_6t
Xbit_r172_c99 bl[99] br[99] wl[172] vdd gnd cell_6t
Xbit_r173_c99 bl[99] br[99] wl[173] vdd gnd cell_6t
Xbit_r174_c99 bl[99] br[99] wl[174] vdd gnd cell_6t
Xbit_r175_c99 bl[99] br[99] wl[175] vdd gnd cell_6t
Xbit_r176_c99 bl[99] br[99] wl[176] vdd gnd cell_6t
Xbit_r177_c99 bl[99] br[99] wl[177] vdd gnd cell_6t
Xbit_r178_c99 bl[99] br[99] wl[178] vdd gnd cell_6t
Xbit_r179_c99 bl[99] br[99] wl[179] vdd gnd cell_6t
Xbit_r180_c99 bl[99] br[99] wl[180] vdd gnd cell_6t
Xbit_r181_c99 bl[99] br[99] wl[181] vdd gnd cell_6t
Xbit_r182_c99 bl[99] br[99] wl[182] vdd gnd cell_6t
Xbit_r183_c99 bl[99] br[99] wl[183] vdd gnd cell_6t
Xbit_r184_c99 bl[99] br[99] wl[184] vdd gnd cell_6t
Xbit_r185_c99 bl[99] br[99] wl[185] vdd gnd cell_6t
Xbit_r186_c99 bl[99] br[99] wl[186] vdd gnd cell_6t
Xbit_r187_c99 bl[99] br[99] wl[187] vdd gnd cell_6t
Xbit_r188_c99 bl[99] br[99] wl[188] vdd gnd cell_6t
Xbit_r189_c99 bl[99] br[99] wl[189] vdd gnd cell_6t
Xbit_r190_c99 bl[99] br[99] wl[190] vdd gnd cell_6t
Xbit_r191_c99 bl[99] br[99] wl[191] vdd gnd cell_6t
Xbit_r192_c99 bl[99] br[99] wl[192] vdd gnd cell_6t
Xbit_r193_c99 bl[99] br[99] wl[193] vdd gnd cell_6t
Xbit_r194_c99 bl[99] br[99] wl[194] vdd gnd cell_6t
Xbit_r195_c99 bl[99] br[99] wl[195] vdd gnd cell_6t
Xbit_r196_c99 bl[99] br[99] wl[196] vdd gnd cell_6t
Xbit_r197_c99 bl[99] br[99] wl[197] vdd gnd cell_6t
Xbit_r198_c99 bl[99] br[99] wl[198] vdd gnd cell_6t
Xbit_r199_c99 bl[99] br[99] wl[199] vdd gnd cell_6t
Xbit_r200_c99 bl[99] br[99] wl[200] vdd gnd cell_6t
Xbit_r201_c99 bl[99] br[99] wl[201] vdd gnd cell_6t
Xbit_r202_c99 bl[99] br[99] wl[202] vdd gnd cell_6t
Xbit_r203_c99 bl[99] br[99] wl[203] vdd gnd cell_6t
Xbit_r204_c99 bl[99] br[99] wl[204] vdd gnd cell_6t
Xbit_r205_c99 bl[99] br[99] wl[205] vdd gnd cell_6t
Xbit_r206_c99 bl[99] br[99] wl[206] vdd gnd cell_6t
Xbit_r207_c99 bl[99] br[99] wl[207] vdd gnd cell_6t
Xbit_r208_c99 bl[99] br[99] wl[208] vdd gnd cell_6t
Xbit_r209_c99 bl[99] br[99] wl[209] vdd gnd cell_6t
Xbit_r210_c99 bl[99] br[99] wl[210] vdd gnd cell_6t
Xbit_r211_c99 bl[99] br[99] wl[211] vdd gnd cell_6t
Xbit_r212_c99 bl[99] br[99] wl[212] vdd gnd cell_6t
Xbit_r213_c99 bl[99] br[99] wl[213] vdd gnd cell_6t
Xbit_r214_c99 bl[99] br[99] wl[214] vdd gnd cell_6t
Xbit_r215_c99 bl[99] br[99] wl[215] vdd gnd cell_6t
Xbit_r216_c99 bl[99] br[99] wl[216] vdd gnd cell_6t
Xbit_r217_c99 bl[99] br[99] wl[217] vdd gnd cell_6t
Xbit_r218_c99 bl[99] br[99] wl[218] vdd gnd cell_6t
Xbit_r219_c99 bl[99] br[99] wl[219] vdd gnd cell_6t
Xbit_r220_c99 bl[99] br[99] wl[220] vdd gnd cell_6t
Xbit_r221_c99 bl[99] br[99] wl[221] vdd gnd cell_6t
Xbit_r222_c99 bl[99] br[99] wl[222] vdd gnd cell_6t
Xbit_r223_c99 bl[99] br[99] wl[223] vdd gnd cell_6t
Xbit_r224_c99 bl[99] br[99] wl[224] vdd gnd cell_6t
Xbit_r225_c99 bl[99] br[99] wl[225] vdd gnd cell_6t
Xbit_r226_c99 bl[99] br[99] wl[226] vdd gnd cell_6t
Xbit_r227_c99 bl[99] br[99] wl[227] vdd gnd cell_6t
Xbit_r228_c99 bl[99] br[99] wl[228] vdd gnd cell_6t
Xbit_r229_c99 bl[99] br[99] wl[229] vdd gnd cell_6t
Xbit_r230_c99 bl[99] br[99] wl[230] vdd gnd cell_6t
Xbit_r231_c99 bl[99] br[99] wl[231] vdd gnd cell_6t
Xbit_r232_c99 bl[99] br[99] wl[232] vdd gnd cell_6t
Xbit_r233_c99 bl[99] br[99] wl[233] vdd gnd cell_6t
Xbit_r234_c99 bl[99] br[99] wl[234] vdd gnd cell_6t
Xbit_r235_c99 bl[99] br[99] wl[235] vdd gnd cell_6t
Xbit_r236_c99 bl[99] br[99] wl[236] vdd gnd cell_6t
Xbit_r237_c99 bl[99] br[99] wl[237] vdd gnd cell_6t
Xbit_r238_c99 bl[99] br[99] wl[238] vdd gnd cell_6t
Xbit_r239_c99 bl[99] br[99] wl[239] vdd gnd cell_6t
Xbit_r240_c99 bl[99] br[99] wl[240] vdd gnd cell_6t
Xbit_r241_c99 bl[99] br[99] wl[241] vdd gnd cell_6t
Xbit_r242_c99 bl[99] br[99] wl[242] vdd gnd cell_6t
Xbit_r243_c99 bl[99] br[99] wl[243] vdd gnd cell_6t
Xbit_r244_c99 bl[99] br[99] wl[244] vdd gnd cell_6t
Xbit_r245_c99 bl[99] br[99] wl[245] vdd gnd cell_6t
Xbit_r246_c99 bl[99] br[99] wl[246] vdd gnd cell_6t
Xbit_r247_c99 bl[99] br[99] wl[247] vdd gnd cell_6t
Xbit_r248_c99 bl[99] br[99] wl[248] vdd gnd cell_6t
Xbit_r249_c99 bl[99] br[99] wl[249] vdd gnd cell_6t
Xbit_r250_c99 bl[99] br[99] wl[250] vdd gnd cell_6t
Xbit_r251_c99 bl[99] br[99] wl[251] vdd gnd cell_6t
Xbit_r252_c99 bl[99] br[99] wl[252] vdd gnd cell_6t
Xbit_r253_c99 bl[99] br[99] wl[253] vdd gnd cell_6t
Xbit_r254_c99 bl[99] br[99] wl[254] vdd gnd cell_6t
Xbit_r255_c99 bl[99] br[99] wl[255] vdd gnd cell_6t
Xbit_r0_c100 bl[100] br[100] wl[0] vdd gnd cell_6t
Xbit_r1_c100 bl[100] br[100] wl[1] vdd gnd cell_6t
Xbit_r2_c100 bl[100] br[100] wl[2] vdd gnd cell_6t
Xbit_r3_c100 bl[100] br[100] wl[3] vdd gnd cell_6t
Xbit_r4_c100 bl[100] br[100] wl[4] vdd gnd cell_6t
Xbit_r5_c100 bl[100] br[100] wl[5] vdd gnd cell_6t
Xbit_r6_c100 bl[100] br[100] wl[6] vdd gnd cell_6t
Xbit_r7_c100 bl[100] br[100] wl[7] vdd gnd cell_6t
Xbit_r8_c100 bl[100] br[100] wl[8] vdd gnd cell_6t
Xbit_r9_c100 bl[100] br[100] wl[9] vdd gnd cell_6t
Xbit_r10_c100 bl[100] br[100] wl[10] vdd gnd cell_6t
Xbit_r11_c100 bl[100] br[100] wl[11] vdd gnd cell_6t
Xbit_r12_c100 bl[100] br[100] wl[12] vdd gnd cell_6t
Xbit_r13_c100 bl[100] br[100] wl[13] vdd gnd cell_6t
Xbit_r14_c100 bl[100] br[100] wl[14] vdd gnd cell_6t
Xbit_r15_c100 bl[100] br[100] wl[15] vdd gnd cell_6t
Xbit_r16_c100 bl[100] br[100] wl[16] vdd gnd cell_6t
Xbit_r17_c100 bl[100] br[100] wl[17] vdd gnd cell_6t
Xbit_r18_c100 bl[100] br[100] wl[18] vdd gnd cell_6t
Xbit_r19_c100 bl[100] br[100] wl[19] vdd gnd cell_6t
Xbit_r20_c100 bl[100] br[100] wl[20] vdd gnd cell_6t
Xbit_r21_c100 bl[100] br[100] wl[21] vdd gnd cell_6t
Xbit_r22_c100 bl[100] br[100] wl[22] vdd gnd cell_6t
Xbit_r23_c100 bl[100] br[100] wl[23] vdd gnd cell_6t
Xbit_r24_c100 bl[100] br[100] wl[24] vdd gnd cell_6t
Xbit_r25_c100 bl[100] br[100] wl[25] vdd gnd cell_6t
Xbit_r26_c100 bl[100] br[100] wl[26] vdd gnd cell_6t
Xbit_r27_c100 bl[100] br[100] wl[27] vdd gnd cell_6t
Xbit_r28_c100 bl[100] br[100] wl[28] vdd gnd cell_6t
Xbit_r29_c100 bl[100] br[100] wl[29] vdd gnd cell_6t
Xbit_r30_c100 bl[100] br[100] wl[30] vdd gnd cell_6t
Xbit_r31_c100 bl[100] br[100] wl[31] vdd gnd cell_6t
Xbit_r32_c100 bl[100] br[100] wl[32] vdd gnd cell_6t
Xbit_r33_c100 bl[100] br[100] wl[33] vdd gnd cell_6t
Xbit_r34_c100 bl[100] br[100] wl[34] vdd gnd cell_6t
Xbit_r35_c100 bl[100] br[100] wl[35] vdd gnd cell_6t
Xbit_r36_c100 bl[100] br[100] wl[36] vdd gnd cell_6t
Xbit_r37_c100 bl[100] br[100] wl[37] vdd gnd cell_6t
Xbit_r38_c100 bl[100] br[100] wl[38] vdd gnd cell_6t
Xbit_r39_c100 bl[100] br[100] wl[39] vdd gnd cell_6t
Xbit_r40_c100 bl[100] br[100] wl[40] vdd gnd cell_6t
Xbit_r41_c100 bl[100] br[100] wl[41] vdd gnd cell_6t
Xbit_r42_c100 bl[100] br[100] wl[42] vdd gnd cell_6t
Xbit_r43_c100 bl[100] br[100] wl[43] vdd gnd cell_6t
Xbit_r44_c100 bl[100] br[100] wl[44] vdd gnd cell_6t
Xbit_r45_c100 bl[100] br[100] wl[45] vdd gnd cell_6t
Xbit_r46_c100 bl[100] br[100] wl[46] vdd gnd cell_6t
Xbit_r47_c100 bl[100] br[100] wl[47] vdd gnd cell_6t
Xbit_r48_c100 bl[100] br[100] wl[48] vdd gnd cell_6t
Xbit_r49_c100 bl[100] br[100] wl[49] vdd gnd cell_6t
Xbit_r50_c100 bl[100] br[100] wl[50] vdd gnd cell_6t
Xbit_r51_c100 bl[100] br[100] wl[51] vdd gnd cell_6t
Xbit_r52_c100 bl[100] br[100] wl[52] vdd gnd cell_6t
Xbit_r53_c100 bl[100] br[100] wl[53] vdd gnd cell_6t
Xbit_r54_c100 bl[100] br[100] wl[54] vdd gnd cell_6t
Xbit_r55_c100 bl[100] br[100] wl[55] vdd gnd cell_6t
Xbit_r56_c100 bl[100] br[100] wl[56] vdd gnd cell_6t
Xbit_r57_c100 bl[100] br[100] wl[57] vdd gnd cell_6t
Xbit_r58_c100 bl[100] br[100] wl[58] vdd gnd cell_6t
Xbit_r59_c100 bl[100] br[100] wl[59] vdd gnd cell_6t
Xbit_r60_c100 bl[100] br[100] wl[60] vdd gnd cell_6t
Xbit_r61_c100 bl[100] br[100] wl[61] vdd gnd cell_6t
Xbit_r62_c100 bl[100] br[100] wl[62] vdd gnd cell_6t
Xbit_r63_c100 bl[100] br[100] wl[63] vdd gnd cell_6t
Xbit_r64_c100 bl[100] br[100] wl[64] vdd gnd cell_6t
Xbit_r65_c100 bl[100] br[100] wl[65] vdd gnd cell_6t
Xbit_r66_c100 bl[100] br[100] wl[66] vdd gnd cell_6t
Xbit_r67_c100 bl[100] br[100] wl[67] vdd gnd cell_6t
Xbit_r68_c100 bl[100] br[100] wl[68] vdd gnd cell_6t
Xbit_r69_c100 bl[100] br[100] wl[69] vdd gnd cell_6t
Xbit_r70_c100 bl[100] br[100] wl[70] vdd gnd cell_6t
Xbit_r71_c100 bl[100] br[100] wl[71] vdd gnd cell_6t
Xbit_r72_c100 bl[100] br[100] wl[72] vdd gnd cell_6t
Xbit_r73_c100 bl[100] br[100] wl[73] vdd gnd cell_6t
Xbit_r74_c100 bl[100] br[100] wl[74] vdd gnd cell_6t
Xbit_r75_c100 bl[100] br[100] wl[75] vdd gnd cell_6t
Xbit_r76_c100 bl[100] br[100] wl[76] vdd gnd cell_6t
Xbit_r77_c100 bl[100] br[100] wl[77] vdd gnd cell_6t
Xbit_r78_c100 bl[100] br[100] wl[78] vdd gnd cell_6t
Xbit_r79_c100 bl[100] br[100] wl[79] vdd gnd cell_6t
Xbit_r80_c100 bl[100] br[100] wl[80] vdd gnd cell_6t
Xbit_r81_c100 bl[100] br[100] wl[81] vdd gnd cell_6t
Xbit_r82_c100 bl[100] br[100] wl[82] vdd gnd cell_6t
Xbit_r83_c100 bl[100] br[100] wl[83] vdd gnd cell_6t
Xbit_r84_c100 bl[100] br[100] wl[84] vdd gnd cell_6t
Xbit_r85_c100 bl[100] br[100] wl[85] vdd gnd cell_6t
Xbit_r86_c100 bl[100] br[100] wl[86] vdd gnd cell_6t
Xbit_r87_c100 bl[100] br[100] wl[87] vdd gnd cell_6t
Xbit_r88_c100 bl[100] br[100] wl[88] vdd gnd cell_6t
Xbit_r89_c100 bl[100] br[100] wl[89] vdd gnd cell_6t
Xbit_r90_c100 bl[100] br[100] wl[90] vdd gnd cell_6t
Xbit_r91_c100 bl[100] br[100] wl[91] vdd gnd cell_6t
Xbit_r92_c100 bl[100] br[100] wl[92] vdd gnd cell_6t
Xbit_r93_c100 bl[100] br[100] wl[93] vdd gnd cell_6t
Xbit_r94_c100 bl[100] br[100] wl[94] vdd gnd cell_6t
Xbit_r95_c100 bl[100] br[100] wl[95] vdd gnd cell_6t
Xbit_r96_c100 bl[100] br[100] wl[96] vdd gnd cell_6t
Xbit_r97_c100 bl[100] br[100] wl[97] vdd gnd cell_6t
Xbit_r98_c100 bl[100] br[100] wl[98] vdd gnd cell_6t
Xbit_r99_c100 bl[100] br[100] wl[99] vdd gnd cell_6t
Xbit_r100_c100 bl[100] br[100] wl[100] vdd gnd cell_6t
Xbit_r101_c100 bl[100] br[100] wl[101] vdd gnd cell_6t
Xbit_r102_c100 bl[100] br[100] wl[102] vdd gnd cell_6t
Xbit_r103_c100 bl[100] br[100] wl[103] vdd gnd cell_6t
Xbit_r104_c100 bl[100] br[100] wl[104] vdd gnd cell_6t
Xbit_r105_c100 bl[100] br[100] wl[105] vdd gnd cell_6t
Xbit_r106_c100 bl[100] br[100] wl[106] vdd gnd cell_6t
Xbit_r107_c100 bl[100] br[100] wl[107] vdd gnd cell_6t
Xbit_r108_c100 bl[100] br[100] wl[108] vdd gnd cell_6t
Xbit_r109_c100 bl[100] br[100] wl[109] vdd gnd cell_6t
Xbit_r110_c100 bl[100] br[100] wl[110] vdd gnd cell_6t
Xbit_r111_c100 bl[100] br[100] wl[111] vdd gnd cell_6t
Xbit_r112_c100 bl[100] br[100] wl[112] vdd gnd cell_6t
Xbit_r113_c100 bl[100] br[100] wl[113] vdd gnd cell_6t
Xbit_r114_c100 bl[100] br[100] wl[114] vdd gnd cell_6t
Xbit_r115_c100 bl[100] br[100] wl[115] vdd gnd cell_6t
Xbit_r116_c100 bl[100] br[100] wl[116] vdd gnd cell_6t
Xbit_r117_c100 bl[100] br[100] wl[117] vdd gnd cell_6t
Xbit_r118_c100 bl[100] br[100] wl[118] vdd gnd cell_6t
Xbit_r119_c100 bl[100] br[100] wl[119] vdd gnd cell_6t
Xbit_r120_c100 bl[100] br[100] wl[120] vdd gnd cell_6t
Xbit_r121_c100 bl[100] br[100] wl[121] vdd gnd cell_6t
Xbit_r122_c100 bl[100] br[100] wl[122] vdd gnd cell_6t
Xbit_r123_c100 bl[100] br[100] wl[123] vdd gnd cell_6t
Xbit_r124_c100 bl[100] br[100] wl[124] vdd gnd cell_6t
Xbit_r125_c100 bl[100] br[100] wl[125] vdd gnd cell_6t
Xbit_r126_c100 bl[100] br[100] wl[126] vdd gnd cell_6t
Xbit_r127_c100 bl[100] br[100] wl[127] vdd gnd cell_6t
Xbit_r128_c100 bl[100] br[100] wl[128] vdd gnd cell_6t
Xbit_r129_c100 bl[100] br[100] wl[129] vdd gnd cell_6t
Xbit_r130_c100 bl[100] br[100] wl[130] vdd gnd cell_6t
Xbit_r131_c100 bl[100] br[100] wl[131] vdd gnd cell_6t
Xbit_r132_c100 bl[100] br[100] wl[132] vdd gnd cell_6t
Xbit_r133_c100 bl[100] br[100] wl[133] vdd gnd cell_6t
Xbit_r134_c100 bl[100] br[100] wl[134] vdd gnd cell_6t
Xbit_r135_c100 bl[100] br[100] wl[135] vdd gnd cell_6t
Xbit_r136_c100 bl[100] br[100] wl[136] vdd gnd cell_6t
Xbit_r137_c100 bl[100] br[100] wl[137] vdd gnd cell_6t
Xbit_r138_c100 bl[100] br[100] wl[138] vdd gnd cell_6t
Xbit_r139_c100 bl[100] br[100] wl[139] vdd gnd cell_6t
Xbit_r140_c100 bl[100] br[100] wl[140] vdd gnd cell_6t
Xbit_r141_c100 bl[100] br[100] wl[141] vdd gnd cell_6t
Xbit_r142_c100 bl[100] br[100] wl[142] vdd gnd cell_6t
Xbit_r143_c100 bl[100] br[100] wl[143] vdd gnd cell_6t
Xbit_r144_c100 bl[100] br[100] wl[144] vdd gnd cell_6t
Xbit_r145_c100 bl[100] br[100] wl[145] vdd gnd cell_6t
Xbit_r146_c100 bl[100] br[100] wl[146] vdd gnd cell_6t
Xbit_r147_c100 bl[100] br[100] wl[147] vdd gnd cell_6t
Xbit_r148_c100 bl[100] br[100] wl[148] vdd gnd cell_6t
Xbit_r149_c100 bl[100] br[100] wl[149] vdd gnd cell_6t
Xbit_r150_c100 bl[100] br[100] wl[150] vdd gnd cell_6t
Xbit_r151_c100 bl[100] br[100] wl[151] vdd gnd cell_6t
Xbit_r152_c100 bl[100] br[100] wl[152] vdd gnd cell_6t
Xbit_r153_c100 bl[100] br[100] wl[153] vdd gnd cell_6t
Xbit_r154_c100 bl[100] br[100] wl[154] vdd gnd cell_6t
Xbit_r155_c100 bl[100] br[100] wl[155] vdd gnd cell_6t
Xbit_r156_c100 bl[100] br[100] wl[156] vdd gnd cell_6t
Xbit_r157_c100 bl[100] br[100] wl[157] vdd gnd cell_6t
Xbit_r158_c100 bl[100] br[100] wl[158] vdd gnd cell_6t
Xbit_r159_c100 bl[100] br[100] wl[159] vdd gnd cell_6t
Xbit_r160_c100 bl[100] br[100] wl[160] vdd gnd cell_6t
Xbit_r161_c100 bl[100] br[100] wl[161] vdd gnd cell_6t
Xbit_r162_c100 bl[100] br[100] wl[162] vdd gnd cell_6t
Xbit_r163_c100 bl[100] br[100] wl[163] vdd gnd cell_6t
Xbit_r164_c100 bl[100] br[100] wl[164] vdd gnd cell_6t
Xbit_r165_c100 bl[100] br[100] wl[165] vdd gnd cell_6t
Xbit_r166_c100 bl[100] br[100] wl[166] vdd gnd cell_6t
Xbit_r167_c100 bl[100] br[100] wl[167] vdd gnd cell_6t
Xbit_r168_c100 bl[100] br[100] wl[168] vdd gnd cell_6t
Xbit_r169_c100 bl[100] br[100] wl[169] vdd gnd cell_6t
Xbit_r170_c100 bl[100] br[100] wl[170] vdd gnd cell_6t
Xbit_r171_c100 bl[100] br[100] wl[171] vdd gnd cell_6t
Xbit_r172_c100 bl[100] br[100] wl[172] vdd gnd cell_6t
Xbit_r173_c100 bl[100] br[100] wl[173] vdd gnd cell_6t
Xbit_r174_c100 bl[100] br[100] wl[174] vdd gnd cell_6t
Xbit_r175_c100 bl[100] br[100] wl[175] vdd gnd cell_6t
Xbit_r176_c100 bl[100] br[100] wl[176] vdd gnd cell_6t
Xbit_r177_c100 bl[100] br[100] wl[177] vdd gnd cell_6t
Xbit_r178_c100 bl[100] br[100] wl[178] vdd gnd cell_6t
Xbit_r179_c100 bl[100] br[100] wl[179] vdd gnd cell_6t
Xbit_r180_c100 bl[100] br[100] wl[180] vdd gnd cell_6t
Xbit_r181_c100 bl[100] br[100] wl[181] vdd gnd cell_6t
Xbit_r182_c100 bl[100] br[100] wl[182] vdd gnd cell_6t
Xbit_r183_c100 bl[100] br[100] wl[183] vdd gnd cell_6t
Xbit_r184_c100 bl[100] br[100] wl[184] vdd gnd cell_6t
Xbit_r185_c100 bl[100] br[100] wl[185] vdd gnd cell_6t
Xbit_r186_c100 bl[100] br[100] wl[186] vdd gnd cell_6t
Xbit_r187_c100 bl[100] br[100] wl[187] vdd gnd cell_6t
Xbit_r188_c100 bl[100] br[100] wl[188] vdd gnd cell_6t
Xbit_r189_c100 bl[100] br[100] wl[189] vdd gnd cell_6t
Xbit_r190_c100 bl[100] br[100] wl[190] vdd gnd cell_6t
Xbit_r191_c100 bl[100] br[100] wl[191] vdd gnd cell_6t
Xbit_r192_c100 bl[100] br[100] wl[192] vdd gnd cell_6t
Xbit_r193_c100 bl[100] br[100] wl[193] vdd gnd cell_6t
Xbit_r194_c100 bl[100] br[100] wl[194] vdd gnd cell_6t
Xbit_r195_c100 bl[100] br[100] wl[195] vdd gnd cell_6t
Xbit_r196_c100 bl[100] br[100] wl[196] vdd gnd cell_6t
Xbit_r197_c100 bl[100] br[100] wl[197] vdd gnd cell_6t
Xbit_r198_c100 bl[100] br[100] wl[198] vdd gnd cell_6t
Xbit_r199_c100 bl[100] br[100] wl[199] vdd gnd cell_6t
Xbit_r200_c100 bl[100] br[100] wl[200] vdd gnd cell_6t
Xbit_r201_c100 bl[100] br[100] wl[201] vdd gnd cell_6t
Xbit_r202_c100 bl[100] br[100] wl[202] vdd gnd cell_6t
Xbit_r203_c100 bl[100] br[100] wl[203] vdd gnd cell_6t
Xbit_r204_c100 bl[100] br[100] wl[204] vdd gnd cell_6t
Xbit_r205_c100 bl[100] br[100] wl[205] vdd gnd cell_6t
Xbit_r206_c100 bl[100] br[100] wl[206] vdd gnd cell_6t
Xbit_r207_c100 bl[100] br[100] wl[207] vdd gnd cell_6t
Xbit_r208_c100 bl[100] br[100] wl[208] vdd gnd cell_6t
Xbit_r209_c100 bl[100] br[100] wl[209] vdd gnd cell_6t
Xbit_r210_c100 bl[100] br[100] wl[210] vdd gnd cell_6t
Xbit_r211_c100 bl[100] br[100] wl[211] vdd gnd cell_6t
Xbit_r212_c100 bl[100] br[100] wl[212] vdd gnd cell_6t
Xbit_r213_c100 bl[100] br[100] wl[213] vdd gnd cell_6t
Xbit_r214_c100 bl[100] br[100] wl[214] vdd gnd cell_6t
Xbit_r215_c100 bl[100] br[100] wl[215] vdd gnd cell_6t
Xbit_r216_c100 bl[100] br[100] wl[216] vdd gnd cell_6t
Xbit_r217_c100 bl[100] br[100] wl[217] vdd gnd cell_6t
Xbit_r218_c100 bl[100] br[100] wl[218] vdd gnd cell_6t
Xbit_r219_c100 bl[100] br[100] wl[219] vdd gnd cell_6t
Xbit_r220_c100 bl[100] br[100] wl[220] vdd gnd cell_6t
Xbit_r221_c100 bl[100] br[100] wl[221] vdd gnd cell_6t
Xbit_r222_c100 bl[100] br[100] wl[222] vdd gnd cell_6t
Xbit_r223_c100 bl[100] br[100] wl[223] vdd gnd cell_6t
Xbit_r224_c100 bl[100] br[100] wl[224] vdd gnd cell_6t
Xbit_r225_c100 bl[100] br[100] wl[225] vdd gnd cell_6t
Xbit_r226_c100 bl[100] br[100] wl[226] vdd gnd cell_6t
Xbit_r227_c100 bl[100] br[100] wl[227] vdd gnd cell_6t
Xbit_r228_c100 bl[100] br[100] wl[228] vdd gnd cell_6t
Xbit_r229_c100 bl[100] br[100] wl[229] vdd gnd cell_6t
Xbit_r230_c100 bl[100] br[100] wl[230] vdd gnd cell_6t
Xbit_r231_c100 bl[100] br[100] wl[231] vdd gnd cell_6t
Xbit_r232_c100 bl[100] br[100] wl[232] vdd gnd cell_6t
Xbit_r233_c100 bl[100] br[100] wl[233] vdd gnd cell_6t
Xbit_r234_c100 bl[100] br[100] wl[234] vdd gnd cell_6t
Xbit_r235_c100 bl[100] br[100] wl[235] vdd gnd cell_6t
Xbit_r236_c100 bl[100] br[100] wl[236] vdd gnd cell_6t
Xbit_r237_c100 bl[100] br[100] wl[237] vdd gnd cell_6t
Xbit_r238_c100 bl[100] br[100] wl[238] vdd gnd cell_6t
Xbit_r239_c100 bl[100] br[100] wl[239] vdd gnd cell_6t
Xbit_r240_c100 bl[100] br[100] wl[240] vdd gnd cell_6t
Xbit_r241_c100 bl[100] br[100] wl[241] vdd gnd cell_6t
Xbit_r242_c100 bl[100] br[100] wl[242] vdd gnd cell_6t
Xbit_r243_c100 bl[100] br[100] wl[243] vdd gnd cell_6t
Xbit_r244_c100 bl[100] br[100] wl[244] vdd gnd cell_6t
Xbit_r245_c100 bl[100] br[100] wl[245] vdd gnd cell_6t
Xbit_r246_c100 bl[100] br[100] wl[246] vdd gnd cell_6t
Xbit_r247_c100 bl[100] br[100] wl[247] vdd gnd cell_6t
Xbit_r248_c100 bl[100] br[100] wl[248] vdd gnd cell_6t
Xbit_r249_c100 bl[100] br[100] wl[249] vdd gnd cell_6t
Xbit_r250_c100 bl[100] br[100] wl[250] vdd gnd cell_6t
Xbit_r251_c100 bl[100] br[100] wl[251] vdd gnd cell_6t
Xbit_r252_c100 bl[100] br[100] wl[252] vdd gnd cell_6t
Xbit_r253_c100 bl[100] br[100] wl[253] vdd gnd cell_6t
Xbit_r254_c100 bl[100] br[100] wl[254] vdd gnd cell_6t
Xbit_r255_c100 bl[100] br[100] wl[255] vdd gnd cell_6t
Xbit_r0_c101 bl[101] br[101] wl[0] vdd gnd cell_6t
Xbit_r1_c101 bl[101] br[101] wl[1] vdd gnd cell_6t
Xbit_r2_c101 bl[101] br[101] wl[2] vdd gnd cell_6t
Xbit_r3_c101 bl[101] br[101] wl[3] vdd gnd cell_6t
Xbit_r4_c101 bl[101] br[101] wl[4] vdd gnd cell_6t
Xbit_r5_c101 bl[101] br[101] wl[5] vdd gnd cell_6t
Xbit_r6_c101 bl[101] br[101] wl[6] vdd gnd cell_6t
Xbit_r7_c101 bl[101] br[101] wl[7] vdd gnd cell_6t
Xbit_r8_c101 bl[101] br[101] wl[8] vdd gnd cell_6t
Xbit_r9_c101 bl[101] br[101] wl[9] vdd gnd cell_6t
Xbit_r10_c101 bl[101] br[101] wl[10] vdd gnd cell_6t
Xbit_r11_c101 bl[101] br[101] wl[11] vdd gnd cell_6t
Xbit_r12_c101 bl[101] br[101] wl[12] vdd gnd cell_6t
Xbit_r13_c101 bl[101] br[101] wl[13] vdd gnd cell_6t
Xbit_r14_c101 bl[101] br[101] wl[14] vdd gnd cell_6t
Xbit_r15_c101 bl[101] br[101] wl[15] vdd gnd cell_6t
Xbit_r16_c101 bl[101] br[101] wl[16] vdd gnd cell_6t
Xbit_r17_c101 bl[101] br[101] wl[17] vdd gnd cell_6t
Xbit_r18_c101 bl[101] br[101] wl[18] vdd gnd cell_6t
Xbit_r19_c101 bl[101] br[101] wl[19] vdd gnd cell_6t
Xbit_r20_c101 bl[101] br[101] wl[20] vdd gnd cell_6t
Xbit_r21_c101 bl[101] br[101] wl[21] vdd gnd cell_6t
Xbit_r22_c101 bl[101] br[101] wl[22] vdd gnd cell_6t
Xbit_r23_c101 bl[101] br[101] wl[23] vdd gnd cell_6t
Xbit_r24_c101 bl[101] br[101] wl[24] vdd gnd cell_6t
Xbit_r25_c101 bl[101] br[101] wl[25] vdd gnd cell_6t
Xbit_r26_c101 bl[101] br[101] wl[26] vdd gnd cell_6t
Xbit_r27_c101 bl[101] br[101] wl[27] vdd gnd cell_6t
Xbit_r28_c101 bl[101] br[101] wl[28] vdd gnd cell_6t
Xbit_r29_c101 bl[101] br[101] wl[29] vdd gnd cell_6t
Xbit_r30_c101 bl[101] br[101] wl[30] vdd gnd cell_6t
Xbit_r31_c101 bl[101] br[101] wl[31] vdd gnd cell_6t
Xbit_r32_c101 bl[101] br[101] wl[32] vdd gnd cell_6t
Xbit_r33_c101 bl[101] br[101] wl[33] vdd gnd cell_6t
Xbit_r34_c101 bl[101] br[101] wl[34] vdd gnd cell_6t
Xbit_r35_c101 bl[101] br[101] wl[35] vdd gnd cell_6t
Xbit_r36_c101 bl[101] br[101] wl[36] vdd gnd cell_6t
Xbit_r37_c101 bl[101] br[101] wl[37] vdd gnd cell_6t
Xbit_r38_c101 bl[101] br[101] wl[38] vdd gnd cell_6t
Xbit_r39_c101 bl[101] br[101] wl[39] vdd gnd cell_6t
Xbit_r40_c101 bl[101] br[101] wl[40] vdd gnd cell_6t
Xbit_r41_c101 bl[101] br[101] wl[41] vdd gnd cell_6t
Xbit_r42_c101 bl[101] br[101] wl[42] vdd gnd cell_6t
Xbit_r43_c101 bl[101] br[101] wl[43] vdd gnd cell_6t
Xbit_r44_c101 bl[101] br[101] wl[44] vdd gnd cell_6t
Xbit_r45_c101 bl[101] br[101] wl[45] vdd gnd cell_6t
Xbit_r46_c101 bl[101] br[101] wl[46] vdd gnd cell_6t
Xbit_r47_c101 bl[101] br[101] wl[47] vdd gnd cell_6t
Xbit_r48_c101 bl[101] br[101] wl[48] vdd gnd cell_6t
Xbit_r49_c101 bl[101] br[101] wl[49] vdd gnd cell_6t
Xbit_r50_c101 bl[101] br[101] wl[50] vdd gnd cell_6t
Xbit_r51_c101 bl[101] br[101] wl[51] vdd gnd cell_6t
Xbit_r52_c101 bl[101] br[101] wl[52] vdd gnd cell_6t
Xbit_r53_c101 bl[101] br[101] wl[53] vdd gnd cell_6t
Xbit_r54_c101 bl[101] br[101] wl[54] vdd gnd cell_6t
Xbit_r55_c101 bl[101] br[101] wl[55] vdd gnd cell_6t
Xbit_r56_c101 bl[101] br[101] wl[56] vdd gnd cell_6t
Xbit_r57_c101 bl[101] br[101] wl[57] vdd gnd cell_6t
Xbit_r58_c101 bl[101] br[101] wl[58] vdd gnd cell_6t
Xbit_r59_c101 bl[101] br[101] wl[59] vdd gnd cell_6t
Xbit_r60_c101 bl[101] br[101] wl[60] vdd gnd cell_6t
Xbit_r61_c101 bl[101] br[101] wl[61] vdd gnd cell_6t
Xbit_r62_c101 bl[101] br[101] wl[62] vdd gnd cell_6t
Xbit_r63_c101 bl[101] br[101] wl[63] vdd gnd cell_6t
Xbit_r64_c101 bl[101] br[101] wl[64] vdd gnd cell_6t
Xbit_r65_c101 bl[101] br[101] wl[65] vdd gnd cell_6t
Xbit_r66_c101 bl[101] br[101] wl[66] vdd gnd cell_6t
Xbit_r67_c101 bl[101] br[101] wl[67] vdd gnd cell_6t
Xbit_r68_c101 bl[101] br[101] wl[68] vdd gnd cell_6t
Xbit_r69_c101 bl[101] br[101] wl[69] vdd gnd cell_6t
Xbit_r70_c101 bl[101] br[101] wl[70] vdd gnd cell_6t
Xbit_r71_c101 bl[101] br[101] wl[71] vdd gnd cell_6t
Xbit_r72_c101 bl[101] br[101] wl[72] vdd gnd cell_6t
Xbit_r73_c101 bl[101] br[101] wl[73] vdd gnd cell_6t
Xbit_r74_c101 bl[101] br[101] wl[74] vdd gnd cell_6t
Xbit_r75_c101 bl[101] br[101] wl[75] vdd gnd cell_6t
Xbit_r76_c101 bl[101] br[101] wl[76] vdd gnd cell_6t
Xbit_r77_c101 bl[101] br[101] wl[77] vdd gnd cell_6t
Xbit_r78_c101 bl[101] br[101] wl[78] vdd gnd cell_6t
Xbit_r79_c101 bl[101] br[101] wl[79] vdd gnd cell_6t
Xbit_r80_c101 bl[101] br[101] wl[80] vdd gnd cell_6t
Xbit_r81_c101 bl[101] br[101] wl[81] vdd gnd cell_6t
Xbit_r82_c101 bl[101] br[101] wl[82] vdd gnd cell_6t
Xbit_r83_c101 bl[101] br[101] wl[83] vdd gnd cell_6t
Xbit_r84_c101 bl[101] br[101] wl[84] vdd gnd cell_6t
Xbit_r85_c101 bl[101] br[101] wl[85] vdd gnd cell_6t
Xbit_r86_c101 bl[101] br[101] wl[86] vdd gnd cell_6t
Xbit_r87_c101 bl[101] br[101] wl[87] vdd gnd cell_6t
Xbit_r88_c101 bl[101] br[101] wl[88] vdd gnd cell_6t
Xbit_r89_c101 bl[101] br[101] wl[89] vdd gnd cell_6t
Xbit_r90_c101 bl[101] br[101] wl[90] vdd gnd cell_6t
Xbit_r91_c101 bl[101] br[101] wl[91] vdd gnd cell_6t
Xbit_r92_c101 bl[101] br[101] wl[92] vdd gnd cell_6t
Xbit_r93_c101 bl[101] br[101] wl[93] vdd gnd cell_6t
Xbit_r94_c101 bl[101] br[101] wl[94] vdd gnd cell_6t
Xbit_r95_c101 bl[101] br[101] wl[95] vdd gnd cell_6t
Xbit_r96_c101 bl[101] br[101] wl[96] vdd gnd cell_6t
Xbit_r97_c101 bl[101] br[101] wl[97] vdd gnd cell_6t
Xbit_r98_c101 bl[101] br[101] wl[98] vdd gnd cell_6t
Xbit_r99_c101 bl[101] br[101] wl[99] vdd gnd cell_6t
Xbit_r100_c101 bl[101] br[101] wl[100] vdd gnd cell_6t
Xbit_r101_c101 bl[101] br[101] wl[101] vdd gnd cell_6t
Xbit_r102_c101 bl[101] br[101] wl[102] vdd gnd cell_6t
Xbit_r103_c101 bl[101] br[101] wl[103] vdd gnd cell_6t
Xbit_r104_c101 bl[101] br[101] wl[104] vdd gnd cell_6t
Xbit_r105_c101 bl[101] br[101] wl[105] vdd gnd cell_6t
Xbit_r106_c101 bl[101] br[101] wl[106] vdd gnd cell_6t
Xbit_r107_c101 bl[101] br[101] wl[107] vdd gnd cell_6t
Xbit_r108_c101 bl[101] br[101] wl[108] vdd gnd cell_6t
Xbit_r109_c101 bl[101] br[101] wl[109] vdd gnd cell_6t
Xbit_r110_c101 bl[101] br[101] wl[110] vdd gnd cell_6t
Xbit_r111_c101 bl[101] br[101] wl[111] vdd gnd cell_6t
Xbit_r112_c101 bl[101] br[101] wl[112] vdd gnd cell_6t
Xbit_r113_c101 bl[101] br[101] wl[113] vdd gnd cell_6t
Xbit_r114_c101 bl[101] br[101] wl[114] vdd gnd cell_6t
Xbit_r115_c101 bl[101] br[101] wl[115] vdd gnd cell_6t
Xbit_r116_c101 bl[101] br[101] wl[116] vdd gnd cell_6t
Xbit_r117_c101 bl[101] br[101] wl[117] vdd gnd cell_6t
Xbit_r118_c101 bl[101] br[101] wl[118] vdd gnd cell_6t
Xbit_r119_c101 bl[101] br[101] wl[119] vdd gnd cell_6t
Xbit_r120_c101 bl[101] br[101] wl[120] vdd gnd cell_6t
Xbit_r121_c101 bl[101] br[101] wl[121] vdd gnd cell_6t
Xbit_r122_c101 bl[101] br[101] wl[122] vdd gnd cell_6t
Xbit_r123_c101 bl[101] br[101] wl[123] vdd gnd cell_6t
Xbit_r124_c101 bl[101] br[101] wl[124] vdd gnd cell_6t
Xbit_r125_c101 bl[101] br[101] wl[125] vdd gnd cell_6t
Xbit_r126_c101 bl[101] br[101] wl[126] vdd gnd cell_6t
Xbit_r127_c101 bl[101] br[101] wl[127] vdd gnd cell_6t
Xbit_r128_c101 bl[101] br[101] wl[128] vdd gnd cell_6t
Xbit_r129_c101 bl[101] br[101] wl[129] vdd gnd cell_6t
Xbit_r130_c101 bl[101] br[101] wl[130] vdd gnd cell_6t
Xbit_r131_c101 bl[101] br[101] wl[131] vdd gnd cell_6t
Xbit_r132_c101 bl[101] br[101] wl[132] vdd gnd cell_6t
Xbit_r133_c101 bl[101] br[101] wl[133] vdd gnd cell_6t
Xbit_r134_c101 bl[101] br[101] wl[134] vdd gnd cell_6t
Xbit_r135_c101 bl[101] br[101] wl[135] vdd gnd cell_6t
Xbit_r136_c101 bl[101] br[101] wl[136] vdd gnd cell_6t
Xbit_r137_c101 bl[101] br[101] wl[137] vdd gnd cell_6t
Xbit_r138_c101 bl[101] br[101] wl[138] vdd gnd cell_6t
Xbit_r139_c101 bl[101] br[101] wl[139] vdd gnd cell_6t
Xbit_r140_c101 bl[101] br[101] wl[140] vdd gnd cell_6t
Xbit_r141_c101 bl[101] br[101] wl[141] vdd gnd cell_6t
Xbit_r142_c101 bl[101] br[101] wl[142] vdd gnd cell_6t
Xbit_r143_c101 bl[101] br[101] wl[143] vdd gnd cell_6t
Xbit_r144_c101 bl[101] br[101] wl[144] vdd gnd cell_6t
Xbit_r145_c101 bl[101] br[101] wl[145] vdd gnd cell_6t
Xbit_r146_c101 bl[101] br[101] wl[146] vdd gnd cell_6t
Xbit_r147_c101 bl[101] br[101] wl[147] vdd gnd cell_6t
Xbit_r148_c101 bl[101] br[101] wl[148] vdd gnd cell_6t
Xbit_r149_c101 bl[101] br[101] wl[149] vdd gnd cell_6t
Xbit_r150_c101 bl[101] br[101] wl[150] vdd gnd cell_6t
Xbit_r151_c101 bl[101] br[101] wl[151] vdd gnd cell_6t
Xbit_r152_c101 bl[101] br[101] wl[152] vdd gnd cell_6t
Xbit_r153_c101 bl[101] br[101] wl[153] vdd gnd cell_6t
Xbit_r154_c101 bl[101] br[101] wl[154] vdd gnd cell_6t
Xbit_r155_c101 bl[101] br[101] wl[155] vdd gnd cell_6t
Xbit_r156_c101 bl[101] br[101] wl[156] vdd gnd cell_6t
Xbit_r157_c101 bl[101] br[101] wl[157] vdd gnd cell_6t
Xbit_r158_c101 bl[101] br[101] wl[158] vdd gnd cell_6t
Xbit_r159_c101 bl[101] br[101] wl[159] vdd gnd cell_6t
Xbit_r160_c101 bl[101] br[101] wl[160] vdd gnd cell_6t
Xbit_r161_c101 bl[101] br[101] wl[161] vdd gnd cell_6t
Xbit_r162_c101 bl[101] br[101] wl[162] vdd gnd cell_6t
Xbit_r163_c101 bl[101] br[101] wl[163] vdd gnd cell_6t
Xbit_r164_c101 bl[101] br[101] wl[164] vdd gnd cell_6t
Xbit_r165_c101 bl[101] br[101] wl[165] vdd gnd cell_6t
Xbit_r166_c101 bl[101] br[101] wl[166] vdd gnd cell_6t
Xbit_r167_c101 bl[101] br[101] wl[167] vdd gnd cell_6t
Xbit_r168_c101 bl[101] br[101] wl[168] vdd gnd cell_6t
Xbit_r169_c101 bl[101] br[101] wl[169] vdd gnd cell_6t
Xbit_r170_c101 bl[101] br[101] wl[170] vdd gnd cell_6t
Xbit_r171_c101 bl[101] br[101] wl[171] vdd gnd cell_6t
Xbit_r172_c101 bl[101] br[101] wl[172] vdd gnd cell_6t
Xbit_r173_c101 bl[101] br[101] wl[173] vdd gnd cell_6t
Xbit_r174_c101 bl[101] br[101] wl[174] vdd gnd cell_6t
Xbit_r175_c101 bl[101] br[101] wl[175] vdd gnd cell_6t
Xbit_r176_c101 bl[101] br[101] wl[176] vdd gnd cell_6t
Xbit_r177_c101 bl[101] br[101] wl[177] vdd gnd cell_6t
Xbit_r178_c101 bl[101] br[101] wl[178] vdd gnd cell_6t
Xbit_r179_c101 bl[101] br[101] wl[179] vdd gnd cell_6t
Xbit_r180_c101 bl[101] br[101] wl[180] vdd gnd cell_6t
Xbit_r181_c101 bl[101] br[101] wl[181] vdd gnd cell_6t
Xbit_r182_c101 bl[101] br[101] wl[182] vdd gnd cell_6t
Xbit_r183_c101 bl[101] br[101] wl[183] vdd gnd cell_6t
Xbit_r184_c101 bl[101] br[101] wl[184] vdd gnd cell_6t
Xbit_r185_c101 bl[101] br[101] wl[185] vdd gnd cell_6t
Xbit_r186_c101 bl[101] br[101] wl[186] vdd gnd cell_6t
Xbit_r187_c101 bl[101] br[101] wl[187] vdd gnd cell_6t
Xbit_r188_c101 bl[101] br[101] wl[188] vdd gnd cell_6t
Xbit_r189_c101 bl[101] br[101] wl[189] vdd gnd cell_6t
Xbit_r190_c101 bl[101] br[101] wl[190] vdd gnd cell_6t
Xbit_r191_c101 bl[101] br[101] wl[191] vdd gnd cell_6t
Xbit_r192_c101 bl[101] br[101] wl[192] vdd gnd cell_6t
Xbit_r193_c101 bl[101] br[101] wl[193] vdd gnd cell_6t
Xbit_r194_c101 bl[101] br[101] wl[194] vdd gnd cell_6t
Xbit_r195_c101 bl[101] br[101] wl[195] vdd gnd cell_6t
Xbit_r196_c101 bl[101] br[101] wl[196] vdd gnd cell_6t
Xbit_r197_c101 bl[101] br[101] wl[197] vdd gnd cell_6t
Xbit_r198_c101 bl[101] br[101] wl[198] vdd gnd cell_6t
Xbit_r199_c101 bl[101] br[101] wl[199] vdd gnd cell_6t
Xbit_r200_c101 bl[101] br[101] wl[200] vdd gnd cell_6t
Xbit_r201_c101 bl[101] br[101] wl[201] vdd gnd cell_6t
Xbit_r202_c101 bl[101] br[101] wl[202] vdd gnd cell_6t
Xbit_r203_c101 bl[101] br[101] wl[203] vdd gnd cell_6t
Xbit_r204_c101 bl[101] br[101] wl[204] vdd gnd cell_6t
Xbit_r205_c101 bl[101] br[101] wl[205] vdd gnd cell_6t
Xbit_r206_c101 bl[101] br[101] wl[206] vdd gnd cell_6t
Xbit_r207_c101 bl[101] br[101] wl[207] vdd gnd cell_6t
Xbit_r208_c101 bl[101] br[101] wl[208] vdd gnd cell_6t
Xbit_r209_c101 bl[101] br[101] wl[209] vdd gnd cell_6t
Xbit_r210_c101 bl[101] br[101] wl[210] vdd gnd cell_6t
Xbit_r211_c101 bl[101] br[101] wl[211] vdd gnd cell_6t
Xbit_r212_c101 bl[101] br[101] wl[212] vdd gnd cell_6t
Xbit_r213_c101 bl[101] br[101] wl[213] vdd gnd cell_6t
Xbit_r214_c101 bl[101] br[101] wl[214] vdd gnd cell_6t
Xbit_r215_c101 bl[101] br[101] wl[215] vdd gnd cell_6t
Xbit_r216_c101 bl[101] br[101] wl[216] vdd gnd cell_6t
Xbit_r217_c101 bl[101] br[101] wl[217] vdd gnd cell_6t
Xbit_r218_c101 bl[101] br[101] wl[218] vdd gnd cell_6t
Xbit_r219_c101 bl[101] br[101] wl[219] vdd gnd cell_6t
Xbit_r220_c101 bl[101] br[101] wl[220] vdd gnd cell_6t
Xbit_r221_c101 bl[101] br[101] wl[221] vdd gnd cell_6t
Xbit_r222_c101 bl[101] br[101] wl[222] vdd gnd cell_6t
Xbit_r223_c101 bl[101] br[101] wl[223] vdd gnd cell_6t
Xbit_r224_c101 bl[101] br[101] wl[224] vdd gnd cell_6t
Xbit_r225_c101 bl[101] br[101] wl[225] vdd gnd cell_6t
Xbit_r226_c101 bl[101] br[101] wl[226] vdd gnd cell_6t
Xbit_r227_c101 bl[101] br[101] wl[227] vdd gnd cell_6t
Xbit_r228_c101 bl[101] br[101] wl[228] vdd gnd cell_6t
Xbit_r229_c101 bl[101] br[101] wl[229] vdd gnd cell_6t
Xbit_r230_c101 bl[101] br[101] wl[230] vdd gnd cell_6t
Xbit_r231_c101 bl[101] br[101] wl[231] vdd gnd cell_6t
Xbit_r232_c101 bl[101] br[101] wl[232] vdd gnd cell_6t
Xbit_r233_c101 bl[101] br[101] wl[233] vdd gnd cell_6t
Xbit_r234_c101 bl[101] br[101] wl[234] vdd gnd cell_6t
Xbit_r235_c101 bl[101] br[101] wl[235] vdd gnd cell_6t
Xbit_r236_c101 bl[101] br[101] wl[236] vdd gnd cell_6t
Xbit_r237_c101 bl[101] br[101] wl[237] vdd gnd cell_6t
Xbit_r238_c101 bl[101] br[101] wl[238] vdd gnd cell_6t
Xbit_r239_c101 bl[101] br[101] wl[239] vdd gnd cell_6t
Xbit_r240_c101 bl[101] br[101] wl[240] vdd gnd cell_6t
Xbit_r241_c101 bl[101] br[101] wl[241] vdd gnd cell_6t
Xbit_r242_c101 bl[101] br[101] wl[242] vdd gnd cell_6t
Xbit_r243_c101 bl[101] br[101] wl[243] vdd gnd cell_6t
Xbit_r244_c101 bl[101] br[101] wl[244] vdd gnd cell_6t
Xbit_r245_c101 bl[101] br[101] wl[245] vdd gnd cell_6t
Xbit_r246_c101 bl[101] br[101] wl[246] vdd gnd cell_6t
Xbit_r247_c101 bl[101] br[101] wl[247] vdd gnd cell_6t
Xbit_r248_c101 bl[101] br[101] wl[248] vdd gnd cell_6t
Xbit_r249_c101 bl[101] br[101] wl[249] vdd gnd cell_6t
Xbit_r250_c101 bl[101] br[101] wl[250] vdd gnd cell_6t
Xbit_r251_c101 bl[101] br[101] wl[251] vdd gnd cell_6t
Xbit_r252_c101 bl[101] br[101] wl[252] vdd gnd cell_6t
Xbit_r253_c101 bl[101] br[101] wl[253] vdd gnd cell_6t
Xbit_r254_c101 bl[101] br[101] wl[254] vdd gnd cell_6t
Xbit_r255_c101 bl[101] br[101] wl[255] vdd gnd cell_6t
Xbit_r0_c102 bl[102] br[102] wl[0] vdd gnd cell_6t
Xbit_r1_c102 bl[102] br[102] wl[1] vdd gnd cell_6t
Xbit_r2_c102 bl[102] br[102] wl[2] vdd gnd cell_6t
Xbit_r3_c102 bl[102] br[102] wl[3] vdd gnd cell_6t
Xbit_r4_c102 bl[102] br[102] wl[4] vdd gnd cell_6t
Xbit_r5_c102 bl[102] br[102] wl[5] vdd gnd cell_6t
Xbit_r6_c102 bl[102] br[102] wl[6] vdd gnd cell_6t
Xbit_r7_c102 bl[102] br[102] wl[7] vdd gnd cell_6t
Xbit_r8_c102 bl[102] br[102] wl[8] vdd gnd cell_6t
Xbit_r9_c102 bl[102] br[102] wl[9] vdd gnd cell_6t
Xbit_r10_c102 bl[102] br[102] wl[10] vdd gnd cell_6t
Xbit_r11_c102 bl[102] br[102] wl[11] vdd gnd cell_6t
Xbit_r12_c102 bl[102] br[102] wl[12] vdd gnd cell_6t
Xbit_r13_c102 bl[102] br[102] wl[13] vdd gnd cell_6t
Xbit_r14_c102 bl[102] br[102] wl[14] vdd gnd cell_6t
Xbit_r15_c102 bl[102] br[102] wl[15] vdd gnd cell_6t
Xbit_r16_c102 bl[102] br[102] wl[16] vdd gnd cell_6t
Xbit_r17_c102 bl[102] br[102] wl[17] vdd gnd cell_6t
Xbit_r18_c102 bl[102] br[102] wl[18] vdd gnd cell_6t
Xbit_r19_c102 bl[102] br[102] wl[19] vdd gnd cell_6t
Xbit_r20_c102 bl[102] br[102] wl[20] vdd gnd cell_6t
Xbit_r21_c102 bl[102] br[102] wl[21] vdd gnd cell_6t
Xbit_r22_c102 bl[102] br[102] wl[22] vdd gnd cell_6t
Xbit_r23_c102 bl[102] br[102] wl[23] vdd gnd cell_6t
Xbit_r24_c102 bl[102] br[102] wl[24] vdd gnd cell_6t
Xbit_r25_c102 bl[102] br[102] wl[25] vdd gnd cell_6t
Xbit_r26_c102 bl[102] br[102] wl[26] vdd gnd cell_6t
Xbit_r27_c102 bl[102] br[102] wl[27] vdd gnd cell_6t
Xbit_r28_c102 bl[102] br[102] wl[28] vdd gnd cell_6t
Xbit_r29_c102 bl[102] br[102] wl[29] vdd gnd cell_6t
Xbit_r30_c102 bl[102] br[102] wl[30] vdd gnd cell_6t
Xbit_r31_c102 bl[102] br[102] wl[31] vdd gnd cell_6t
Xbit_r32_c102 bl[102] br[102] wl[32] vdd gnd cell_6t
Xbit_r33_c102 bl[102] br[102] wl[33] vdd gnd cell_6t
Xbit_r34_c102 bl[102] br[102] wl[34] vdd gnd cell_6t
Xbit_r35_c102 bl[102] br[102] wl[35] vdd gnd cell_6t
Xbit_r36_c102 bl[102] br[102] wl[36] vdd gnd cell_6t
Xbit_r37_c102 bl[102] br[102] wl[37] vdd gnd cell_6t
Xbit_r38_c102 bl[102] br[102] wl[38] vdd gnd cell_6t
Xbit_r39_c102 bl[102] br[102] wl[39] vdd gnd cell_6t
Xbit_r40_c102 bl[102] br[102] wl[40] vdd gnd cell_6t
Xbit_r41_c102 bl[102] br[102] wl[41] vdd gnd cell_6t
Xbit_r42_c102 bl[102] br[102] wl[42] vdd gnd cell_6t
Xbit_r43_c102 bl[102] br[102] wl[43] vdd gnd cell_6t
Xbit_r44_c102 bl[102] br[102] wl[44] vdd gnd cell_6t
Xbit_r45_c102 bl[102] br[102] wl[45] vdd gnd cell_6t
Xbit_r46_c102 bl[102] br[102] wl[46] vdd gnd cell_6t
Xbit_r47_c102 bl[102] br[102] wl[47] vdd gnd cell_6t
Xbit_r48_c102 bl[102] br[102] wl[48] vdd gnd cell_6t
Xbit_r49_c102 bl[102] br[102] wl[49] vdd gnd cell_6t
Xbit_r50_c102 bl[102] br[102] wl[50] vdd gnd cell_6t
Xbit_r51_c102 bl[102] br[102] wl[51] vdd gnd cell_6t
Xbit_r52_c102 bl[102] br[102] wl[52] vdd gnd cell_6t
Xbit_r53_c102 bl[102] br[102] wl[53] vdd gnd cell_6t
Xbit_r54_c102 bl[102] br[102] wl[54] vdd gnd cell_6t
Xbit_r55_c102 bl[102] br[102] wl[55] vdd gnd cell_6t
Xbit_r56_c102 bl[102] br[102] wl[56] vdd gnd cell_6t
Xbit_r57_c102 bl[102] br[102] wl[57] vdd gnd cell_6t
Xbit_r58_c102 bl[102] br[102] wl[58] vdd gnd cell_6t
Xbit_r59_c102 bl[102] br[102] wl[59] vdd gnd cell_6t
Xbit_r60_c102 bl[102] br[102] wl[60] vdd gnd cell_6t
Xbit_r61_c102 bl[102] br[102] wl[61] vdd gnd cell_6t
Xbit_r62_c102 bl[102] br[102] wl[62] vdd gnd cell_6t
Xbit_r63_c102 bl[102] br[102] wl[63] vdd gnd cell_6t
Xbit_r64_c102 bl[102] br[102] wl[64] vdd gnd cell_6t
Xbit_r65_c102 bl[102] br[102] wl[65] vdd gnd cell_6t
Xbit_r66_c102 bl[102] br[102] wl[66] vdd gnd cell_6t
Xbit_r67_c102 bl[102] br[102] wl[67] vdd gnd cell_6t
Xbit_r68_c102 bl[102] br[102] wl[68] vdd gnd cell_6t
Xbit_r69_c102 bl[102] br[102] wl[69] vdd gnd cell_6t
Xbit_r70_c102 bl[102] br[102] wl[70] vdd gnd cell_6t
Xbit_r71_c102 bl[102] br[102] wl[71] vdd gnd cell_6t
Xbit_r72_c102 bl[102] br[102] wl[72] vdd gnd cell_6t
Xbit_r73_c102 bl[102] br[102] wl[73] vdd gnd cell_6t
Xbit_r74_c102 bl[102] br[102] wl[74] vdd gnd cell_6t
Xbit_r75_c102 bl[102] br[102] wl[75] vdd gnd cell_6t
Xbit_r76_c102 bl[102] br[102] wl[76] vdd gnd cell_6t
Xbit_r77_c102 bl[102] br[102] wl[77] vdd gnd cell_6t
Xbit_r78_c102 bl[102] br[102] wl[78] vdd gnd cell_6t
Xbit_r79_c102 bl[102] br[102] wl[79] vdd gnd cell_6t
Xbit_r80_c102 bl[102] br[102] wl[80] vdd gnd cell_6t
Xbit_r81_c102 bl[102] br[102] wl[81] vdd gnd cell_6t
Xbit_r82_c102 bl[102] br[102] wl[82] vdd gnd cell_6t
Xbit_r83_c102 bl[102] br[102] wl[83] vdd gnd cell_6t
Xbit_r84_c102 bl[102] br[102] wl[84] vdd gnd cell_6t
Xbit_r85_c102 bl[102] br[102] wl[85] vdd gnd cell_6t
Xbit_r86_c102 bl[102] br[102] wl[86] vdd gnd cell_6t
Xbit_r87_c102 bl[102] br[102] wl[87] vdd gnd cell_6t
Xbit_r88_c102 bl[102] br[102] wl[88] vdd gnd cell_6t
Xbit_r89_c102 bl[102] br[102] wl[89] vdd gnd cell_6t
Xbit_r90_c102 bl[102] br[102] wl[90] vdd gnd cell_6t
Xbit_r91_c102 bl[102] br[102] wl[91] vdd gnd cell_6t
Xbit_r92_c102 bl[102] br[102] wl[92] vdd gnd cell_6t
Xbit_r93_c102 bl[102] br[102] wl[93] vdd gnd cell_6t
Xbit_r94_c102 bl[102] br[102] wl[94] vdd gnd cell_6t
Xbit_r95_c102 bl[102] br[102] wl[95] vdd gnd cell_6t
Xbit_r96_c102 bl[102] br[102] wl[96] vdd gnd cell_6t
Xbit_r97_c102 bl[102] br[102] wl[97] vdd gnd cell_6t
Xbit_r98_c102 bl[102] br[102] wl[98] vdd gnd cell_6t
Xbit_r99_c102 bl[102] br[102] wl[99] vdd gnd cell_6t
Xbit_r100_c102 bl[102] br[102] wl[100] vdd gnd cell_6t
Xbit_r101_c102 bl[102] br[102] wl[101] vdd gnd cell_6t
Xbit_r102_c102 bl[102] br[102] wl[102] vdd gnd cell_6t
Xbit_r103_c102 bl[102] br[102] wl[103] vdd gnd cell_6t
Xbit_r104_c102 bl[102] br[102] wl[104] vdd gnd cell_6t
Xbit_r105_c102 bl[102] br[102] wl[105] vdd gnd cell_6t
Xbit_r106_c102 bl[102] br[102] wl[106] vdd gnd cell_6t
Xbit_r107_c102 bl[102] br[102] wl[107] vdd gnd cell_6t
Xbit_r108_c102 bl[102] br[102] wl[108] vdd gnd cell_6t
Xbit_r109_c102 bl[102] br[102] wl[109] vdd gnd cell_6t
Xbit_r110_c102 bl[102] br[102] wl[110] vdd gnd cell_6t
Xbit_r111_c102 bl[102] br[102] wl[111] vdd gnd cell_6t
Xbit_r112_c102 bl[102] br[102] wl[112] vdd gnd cell_6t
Xbit_r113_c102 bl[102] br[102] wl[113] vdd gnd cell_6t
Xbit_r114_c102 bl[102] br[102] wl[114] vdd gnd cell_6t
Xbit_r115_c102 bl[102] br[102] wl[115] vdd gnd cell_6t
Xbit_r116_c102 bl[102] br[102] wl[116] vdd gnd cell_6t
Xbit_r117_c102 bl[102] br[102] wl[117] vdd gnd cell_6t
Xbit_r118_c102 bl[102] br[102] wl[118] vdd gnd cell_6t
Xbit_r119_c102 bl[102] br[102] wl[119] vdd gnd cell_6t
Xbit_r120_c102 bl[102] br[102] wl[120] vdd gnd cell_6t
Xbit_r121_c102 bl[102] br[102] wl[121] vdd gnd cell_6t
Xbit_r122_c102 bl[102] br[102] wl[122] vdd gnd cell_6t
Xbit_r123_c102 bl[102] br[102] wl[123] vdd gnd cell_6t
Xbit_r124_c102 bl[102] br[102] wl[124] vdd gnd cell_6t
Xbit_r125_c102 bl[102] br[102] wl[125] vdd gnd cell_6t
Xbit_r126_c102 bl[102] br[102] wl[126] vdd gnd cell_6t
Xbit_r127_c102 bl[102] br[102] wl[127] vdd gnd cell_6t
Xbit_r128_c102 bl[102] br[102] wl[128] vdd gnd cell_6t
Xbit_r129_c102 bl[102] br[102] wl[129] vdd gnd cell_6t
Xbit_r130_c102 bl[102] br[102] wl[130] vdd gnd cell_6t
Xbit_r131_c102 bl[102] br[102] wl[131] vdd gnd cell_6t
Xbit_r132_c102 bl[102] br[102] wl[132] vdd gnd cell_6t
Xbit_r133_c102 bl[102] br[102] wl[133] vdd gnd cell_6t
Xbit_r134_c102 bl[102] br[102] wl[134] vdd gnd cell_6t
Xbit_r135_c102 bl[102] br[102] wl[135] vdd gnd cell_6t
Xbit_r136_c102 bl[102] br[102] wl[136] vdd gnd cell_6t
Xbit_r137_c102 bl[102] br[102] wl[137] vdd gnd cell_6t
Xbit_r138_c102 bl[102] br[102] wl[138] vdd gnd cell_6t
Xbit_r139_c102 bl[102] br[102] wl[139] vdd gnd cell_6t
Xbit_r140_c102 bl[102] br[102] wl[140] vdd gnd cell_6t
Xbit_r141_c102 bl[102] br[102] wl[141] vdd gnd cell_6t
Xbit_r142_c102 bl[102] br[102] wl[142] vdd gnd cell_6t
Xbit_r143_c102 bl[102] br[102] wl[143] vdd gnd cell_6t
Xbit_r144_c102 bl[102] br[102] wl[144] vdd gnd cell_6t
Xbit_r145_c102 bl[102] br[102] wl[145] vdd gnd cell_6t
Xbit_r146_c102 bl[102] br[102] wl[146] vdd gnd cell_6t
Xbit_r147_c102 bl[102] br[102] wl[147] vdd gnd cell_6t
Xbit_r148_c102 bl[102] br[102] wl[148] vdd gnd cell_6t
Xbit_r149_c102 bl[102] br[102] wl[149] vdd gnd cell_6t
Xbit_r150_c102 bl[102] br[102] wl[150] vdd gnd cell_6t
Xbit_r151_c102 bl[102] br[102] wl[151] vdd gnd cell_6t
Xbit_r152_c102 bl[102] br[102] wl[152] vdd gnd cell_6t
Xbit_r153_c102 bl[102] br[102] wl[153] vdd gnd cell_6t
Xbit_r154_c102 bl[102] br[102] wl[154] vdd gnd cell_6t
Xbit_r155_c102 bl[102] br[102] wl[155] vdd gnd cell_6t
Xbit_r156_c102 bl[102] br[102] wl[156] vdd gnd cell_6t
Xbit_r157_c102 bl[102] br[102] wl[157] vdd gnd cell_6t
Xbit_r158_c102 bl[102] br[102] wl[158] vdd gnd cell_6t
Xbit_r159_c102 bl[102] br[102] wl[159] vdd gnd cell_6t
Xbit_r160_c102 bl[102] br[102] wl[160] vdd gnd cell_6t
Xbit_r161_c102 bl[102] br[102] wl[161] vdd gnd cell_6t
Xbit_r162_c102 bl[102] br[102] wl[162] vdd gnd cell_6t
Xbit_r163_c102 bl[102] br[102] wl[163] vdd gnd cell_6t
Xbit_r164_c102 bl[102] br[102] wl[164] vdd gnd cell_6t
Xbit_r165_c102 bl[102] br[102] wl[165] vdd gnd cell_6t
Xbit_r166_c102 bl[102] br[102] wl[166] vdd gnd cell_6t
Xbit_r167_c102 bl[102] br[102] wl[167] vdd gnd cell_6t
Xbit_r168_c102 bl[102] br[102] wl[168] vdd gnd cell_6t
Xbit_r169_c102 bl[102] br[102] wl[169] vdd gnd cell_6t
Xbit_r170_c102 bl[102] br[102] wl[170] vdd gnd cell_6t
Xbit_r171_c102 bl[102] br[102] wl[171] vdd gnd cell_6t
Xbit_r172_c102 bl[102] br[102] wl[172] vdd gnd cell_6t
Xbit_r173_c102 bl[102] br[102] wl[173] vdd gnd cell_6t
Xbit_r174_c102 bl[102] br[102] wl[174] vdd gnd cell_6t
Xbit_r175_c102 bl[102] br[102] wl[175] vdd gnd cell_6t
Xbit_r176_c102 bl[102] br[102] wl[176] vdd gnd cell_6t
Xbit_r177_c102 bl[102] br[102] wl[177] vdd gnd cell_6t
Xbit_r178_c102 bl[102] br[102] wl[178] vdd gnd cell_6t
Xbit_r179_c102 bl[102] br[102] wl[179] vdd gnd cell_6t
Xbit_r180_c102 bl[102] br[102] wl[180] vdd gnd cell_6t
Xbit_r181_c102 bl[102] br[102] wl[181] vdd gnd cell_6t
Xbit_r182_c102 bl[102] br[102] wl[182] vdd gnd cell_6t
Xbit_r183_c102 bl[102] br[102] wl[183] vdd gnd cell_6t
Xbit_r184_c102 bl[102] br[102] wl[184] vdd gnd cell_6t
Xbit_r185_c102 bl[102] br[102] wl[185] vdd gnd cell_6t
Xbit_r186_c102 bl[102] br[102] wl[186] vdd gnd cell_6t
Xbit_r187_c102 bl[102] br[102] wl[187] vdd gnd cell_6t
Xbit_r188_c102 bl[102] br[102] wl[188] vdd gnd cell_6t
Xbit_r189_c102 bl[102] br[102] wl[189] vdd gnd cell_6t
Xbit_r190_c102 bl[102] br[102] wl[190] vdd gnd cell_6t
Xbit_r191_c102 bl[102] br[102] wl[191] vdd gnd cell_6t
Xbit_r192_c102 bl[102] br[102] wl[192] vdd gnd cell_6t
Xbit_r193_c102 bl[102] br[102] wl[193] vdd gnd cell_6t
Xbit_r194_c102 bl[102] br[102] wl[194] vdd gnd cell_6t
Xbit_r195_c102 bl[102] br[102] wl[195] vdd gnd cell_6t
Xbit_r196_c102 bl[102] br[102] wl[196] vdd gnd cell_6t
Xbit_r197_c102 bl[102] br[102] wl[197] vdd gnd cell_6t
Xbit_r198_c102 bl[102] br[102] wl[198] vdd gnd cell_6t
Xbit_r199_c102 bl[102] br[102] wl[199] vdd gnd cell_6t
Xbit_r200_c102 bl[102] br[102] wl[200] vdd gnd cell_6t
Xbit_r201_c102 bl[102] br[102] wl[201] vdd gnd cell_6t
Xbit_r202_c102 bl[102] br[102] wl[202] vdd gnd cell_6t
Xbit_r203_c102 bl[102] br[102] wl[203] vdd gnd cell_6t
Xbit_r204_c102 bl[102] br[102] wl[204] vdd gnd cell_6t
Xbit_r205_c102 bl[102] br[102] wl[205] vdd gnd cell_6t
Xbit_r206_c102 bl[102] br[102] wl[206] vdd gnd cell_6t
Xbit_r207_c102 bl[102] br[102] wl[207] vdd gnd cell_6t
Xbit_r208_c102 bl[102] br[102] wl[208] vdd gnd cell_6t
Xbit_r209_c102 bl[102] br[102] wl[209] vdd gnd cell_6t
Xbit_r210_c102 bl[102] br[102] wl[210] vdd gnd cell_6t
Xbit_r211_c102 bl[102] br[102] wl[211] vdd gnd cell_6t
Xbit_r212_c102 bl[102] br[102] wl[212] vdd gnd cell_6t
Xbit_r213_c102 bl[102] br[102] wl[213] vdd gnd cell_6t
Xbit_r214_c102 bl[102] br[102] wl[214] vdd gnd cell_6t
Xbit_r215_c102 bl[102] br[102] wl[215] vdd gnd cell_6t
Xbit_r216_c102 bl[102] br[102] wl[216] vdd gnd cell_6t
Xbit_r217_c102 bl[102] br[102] wl[217] vdd gnd cell_6t
Xbit_r218_c102 bl[102] br[102] wl[218] vdd gnd cell_6t
Xbit_r219_c102 bl[102] br[102] wl[219] vdd gnd cell_6t
Xbit_r220_c102 bl[102] br[102] wl[220] vdd gnd cell_6t
Xbit_r221_c102 bl[102] br[102] wl[221] vdd gnd cell_6t
Xbit_r222_c102 bl[102] br[102] wl[222] vdd gnd cell_6t
Xbit_r223_c102 bl[102] br[102] wl[223] vdd gnd cell_6t
Xbit_r224_c102 bl[102] br[102] wl[224] vdd gnd cell_6t
Xbit_r225_c102 bl[102] br[102] wl[225] vdd gnd cell_6t
Xbit_r226_c102 bl[102] br[102] wl[226] vdd gnd cell_6t
Xbit_r227_c102 bl[102] br[102] wl[227] vdd gnd cell_6t
Xbit_r228_c102 bl[102] br[102] wl[228] vdd gnd cell_6t
Xbit_r229_c102 bl[102] br[102] wl[229] vdd gnd cell_6t
Xbit_r230_c102 bl[102] br[102] wl[230] vdd gnd cell_6t
Xbit_r231_c102 bl[102] br[102] wl[231] vdd gnd cell_6t
Xbit_r232_c102 bl[102] br[102] wl[232] vdd gnd cell_6t
Xbit_r233_c102 bl[102] br[102] wl[233] vdd gnd cell_6t
Xbit_r234_c102 bl[102] br[102] wl[234] vdd gnd cell_6t
Xbit_r235_c102 bl[102] br[102] wl[235] vdd gnd cell_6t
Xbit_r236_c102 bl[102] br[102] wl[236] vdd gnd cell_6t
Xbit_r237_c102 bl[102] br[102] wl[237] vdd gnd cell_6t
Xbit_r238_c102 bl[102] br[102] wl[238] vdd gnd cell_6t
Xbit_r239_c102 bl[102] br[102] wl[239] vdd gnd cell_6t
Xbit_r240_c102 bl[102] br[102] wl[240] vdd gnd cell_6t
Xbit_r241_c102 bl[102] br[102] wl[241] vdd gnd cell_6t
Xbit_r242_c102 bl[102] br[102] wl[242] vdd gnd cell_6t
Xbit_r243_c102 bl[102] br[102] wl[243] vdd gnd cell_6t
Xbit_r244_c102 bl[102] br[102] wl[244] vdd gnd cell_6t
Xbit_r245_c102 bl[102] br[102] wl[245] vdd gnd cell_6t
Xbit_r246_c102 bl[102] br[102] wl[246] vdd gnd cell_6t
Xbit_r247_c102 bl[102] br[102] wl[247] vdd gnd cell_6t
Xbit_r248_c102 bl[102] br[102] wl[248] vdd gnd cell_6t
Xbit_r249_c102 bl[102] br[102] wl[249] vdd gnd cell_6t
Xbit_r250_c102 bl[102] br[102] wl[250] vdd gnd cell_6t
Xbit_r251_c102 bl[102] br[102] wl[251] vdd gnd cell_6t
Xbit_r252_c102 bl[102] br[102] wl[252] vdd gnd cell_6t
Xbit_r253_c102 bl[102] br[102] wl[253] vdd gnd cell_6t
Xbit_r254_c102 bl[102] br[102] wl[254] vdd gnd cell_6t
Xbit_r255_c102 bl[102] br[102] wl[255] vdd gnd cell_6t
Xbit_r0_c103 bl[103] br[103] wl[0] vdd gnd cell_6t
Xbit_r1_c103 bl[103] br[103] wl[1] vdd gnd cell_6t
Xbit_r2_c103 bl[103] br[103] wl[2] vdd gnd cell_6t
Xbit_r3_c103 bl[103] br[103] wl[3] vdd gnd cell_6t
Xbit_r4_c103 bl[103] br[103] wl[4] vdd gnd cell_6t
Xbit_r5_c103 bl[103] br[103] wl[5] vdd gnd cell_6t
Xbit_r6_c103 bl[103] br[103] wl[6] vdd gnd cell_6t
Xbit_r7_c103 bl[103] br[103] wl[7] vdd gnd cell_6t
Xbit_r8_c103 bl[103] br[103] wl[8] vdd gnd cell_6t
Xbit_r9_c103 bl[103] br[103] wl[9] vdd gnd cell_6t
Xbit_r10_c103 bl[103] br[103] wl[10] vdd gnd cell_6t
Xbit_r11_c103 bl[103] br[103] wl[11] vdd gnd cell_6t
Xbit_r12_c103 bl[103] br[103] wl[12] vdd gnd cell_6t
Xbit_r13_c103 bl[103] br[103] wl[13] vdd gnd cell_6t
Xbit_r14_c103 bl[103] br[103] wl[14] vdd gnd cell_6t
Xbit_r15_c103 bl[103] br[103] wl[15] vdd gnd cell_6t
Xbit_r16_c103 bl[103] br[103] wl[16] vdd gnd cell_6t
Xbit_r17_c103 bl[103] br[103] wl[17] vdd gnd cell_6t
Xbit_r18_c103 bl[103] br[103] wl[18] vdd gnd cell_6t
Xbit_r19_c103 bl[103] br[103] wl[19] vdd gnd cell_6t
Xbit_r20_c103 bl[103] br[103] wl[20] vdd gnd cell_6t
Xbit_r21_c103 bl[103] br[103] wl[21] vdd gnd cell_6t
Xbit_r22_c103 bl[103] br[103] wl[22] vdd gnd cell_6t
Xbit_r23_c103 bl[103] br[103] wl[23] vdd gnd cell_6t
Xbit_r24_c103 bl[103] br[103] wl[24] vdd gnd cell_6t
Xbit_r25_c103 bl[103] br[103] wl[25] vdd gnd cell_6t
Xbit_r26_c103 bl[103] br[103] wl[26] vdd gnd cell_6t
Xbit_r27_c103 bl[103] br[103] wl[27] vdd gnd cell_6t
Xbit_r28_c103 bl[103] br[103] wl[28] vdd gnd cell_6t
Xbit_r29_c103 bl[103] br[103] wl[29] vdd gnd cell_6t
Xbit_r30_c103 bl[103] br[103] wl[30] vdd gnd cell_6t
Xbit_r31_c103 bl[103] br[103] wl[31] vdd gnd cell_6t
Xbit_r32_c103 bl[103] br[103] wl[32] vdd gnd cell_6t
Xbit_r33_c103 bl[103] br[103] wl[33] vdd gnd cell_6t
Xbit_r34_c103 bl[103] br[103] wl[34] vdd gnd cell_6t
Xbit_r35_c103 bl[103] br[103] wl[35] vdd gnd cell_6t
Xbit_r36_c103 bl[103] br[103] wl[36] vdd gnd cell_6t
Xbit_r37_c103 bl[103] br[103] wl[37] vdd gnd cell_6t
Xbit_r38_c103 bl[103] br[103] wl[38] vdd gnd cell_6t
Xbit_r39_c103 bl[103] br[103] wl[39] vdd gnd cell_6t
Xbit_r40_c103 bl[103] br[103] wl[40] vdd gnd cell_6t
Xbit_r41_c103 bl[103] br[103] wl[41] vdd gnd cell_6t
Xbit_r42_c103 bl[103] br[103] wl[42] vdd gnd cell_6t
Xbit_r43_c103 bl[103] br[103] wl[43] vdd gnd cell_6t
Xbit_r44_c103 bl[103] br[103] wl[44] vdd gnd cell_6t
Xbit_r45_c103 bl[103] br[103] wl[45] vdd gnd cell_6t
Xbit_r46_c103 bl[103] br[103] wl[46] vdd gnd cell_6t
Xbit_r47_c103 bl[103] br[103] wl[47] vdd gnd cell_6t
Xbit_r48_c103 bl[103] br[103] wl[48] vdd gnd cell_6t
Xbit_r49_c103 bl[103] br[103] wl[49] vdd gnd cell_6t
Xbit_r50_c103 bl[103] br[103] wl[50] vdd gnd cell_6t
Xbit_r51_c103 bl[103] br[103] wl[51] vdd gnd cell_6t
Xbit_r52_c103 bl[103] br[103] wl[52] vdd gnd cell_6t
Xbit_r53_c103 bl[103] br[103] wl[53] vdd gnd cell_6t
Xbit_r54_c103 bl[103] br[103] wl[54] vdd gnd cell_6t
Xbit_r55_c103 bl[103] br[103] wl[55] vdd gnd cell_6t
Xbit_r56_c103 bl[103] br[103] wl[56] vdd gnd cell_6t
Xbit_r57_c103 bl[103] br[103] wl[57] vdd gnd cell_6t
Xbit_r58_c103 bl[103] br[103] wl[58] vdd gnd cell_6t
Xbit_r59_c103 bl[103] br[103] wl[59] vdd gnd cell_6t
Xbit_r60_c103 bl[103] br[103] wl[60] vdd gnd cell_6t
Xbit_r61_c103 bl[103] br[103] wl[61] vdd gnd cell_6t
Xbit_r62_c103 bl[103] br[103] wl[62] vdd gnd cell_6t
Xbit_r63_c103 bl[103] br[103] wl[63] vdd gnd cell_6t
Xbit_r64_c103 bl[103] br[103] wl[64] vdd gnd cell_6t
Xbit_r65_c103 bl[103] br[103] wl[65] vdd gnd cell_6t
Xbit_r66_c103 bl[103] br[103] wl[66] vdd gnd cell_6t
Xbit_r67_c103 bl[103] br[103] wl[67] vdd gnd cell_6t
Xbit_r68_c103 bl[103] br[103] wl[68] vdd gnd cell_6t
Xbit_r69_c103 bl[103] br[103] wl[69] vdd gnd cell_6t
Xbit_r70_c103 bl[103] br[103] wl[70] vdd gnd cell_6t
Xbit_r71_c103 bl[103] br[103] wl[71] vdd gnd cell_6t
Xbit_r72_c103 bl[103] br[103] wl[72] vdd gnd cell_6t
Xbit_r73_c103 bl[103] br[103] wl[73] vdd gnd cell_6t
Xbit_r74_c103 bl[103] br[103] wl[74] vdd gnd cell_6t
Xbit_r75_c103 bl[103] br[103] wl[75] vdd gnd cell_6t
Xbit_r76_c103 bl[103] br[103] wl[76] vdd gnd cell_6t
Xbit_r77_c103 bl[103] br[103] wl[77] vdd gnd cell_6t
Xbit_r78_c103 bl[103] br[103] wl[78] vdd gnd cell_6t
Xbit_r79_c103 bl[103] br[103] wl[79] vdd gnd cell_6t
Xbit_r80_c103 bl[103] br[103] wl[80] vdd gnd cell_6t
Xbit_r81_c103 bl[103] br[103] wl[81] vdd gnd cell_6t
Xbit_r82_c103 bl[103] br[103] wl[82] vdd gnd cell_6t
Xbit_r83_c103 bl[103] br[103] wl[83] vdd gnd cell_6t
Xbit_r84_c103 bl[103] br[103] wl[84] vdd gnd cell_6t
Xbit_r85_c103 bl[103] br[103] wl[85] vdd gnd cell_6t
Xbit_r86_c103 bl[103] br[103] wl[86] vdd gnd cell_6t
Xbit_r87_c103 bl[103] br[103] wl[87] vdd gnd cell_6t
Xbit_r88_c103 bl[103] br[103] wl[88] vdd gnd cell_6t
Xbit_r89_c103 bl[103] br[103] wl[89] vdd gnd cell_6t
Xbit_r90_c103 bl[103] br[103] wl[90] vdd gnd cell_6t
Xbit_r91_c103 bl[103] br[103] wl[91] vdd gnd cell_6t
Xbit_r92_c103 bl[103] br[103] wl[92] vdd gnd cell_6t
Xbit_r93_c103 bl[103] br[103] wl[93] vdd gnd cell_6t
Xbit_r94_c103 bl[103] br[103] wl[94] vdd gnd cell_6t
Xbit_r95_c103 bl[103] br[103] wl[95] vdd gnd cell_6t
Xbit_r96_c103 bl[103] br[103] wl[96] vdd gnd cell_6t
Xbit_r97_c103 bl[103] br[103] wl[97] vdd gnd cell_6t
Xbit_r98_c103 bl[103] br[103] wl[98] vdd gnd cell_6t
Xbit_r99_c103 bl[103] br[103] wl[99] vdd gnd cell_6t
Xbit_r100_c103 bl[103] br[103] wl[100] vdd gnd cell_6t
Xbit_r101_c103 bl[103] br[103] wl[101] vdd gnd cell_6t
Xbit_r102_c103 bl[103] br[103] wl[102] vdd gnd cell_6t
Xbit_r103_c103 bl[103] br[103] wl[103] vdd gnd cell_6t
Xbit_r104_c103 bl[103] br[103] wl[104] vdd gnd cell_6t
Xbit_r105_c103 bl[103] br[103] wl[105] vdd gnd cell_6t
Xbit_r106_c103 bl[103] br[103] wl[106] vdd gnd cell_6t
Xbit_r107_c103 bl[103] br[103] wl[107] vdd gnd cell_6t
Xbit_r108_c103 bl[103] br[103] wl[108] vdd gnd cell_6t
Xbit_r109_c103 bl[103] br[103] wl[109] vdd gnd cell_6t
Xbit_r110_c103 bl[103] br[103] wl[110] vdd gnd cell_6t
Xbit_r111_c103 bl[103] br[103] wl[111] vdd gnd cell_6t
Xbit_r112_c103 bl[103] br[103] wl[112] vdd gnd cell_6t
Xbit_r113_c103 bl[103] br[103] wl[113] vdd gnd cell_6t
Xbit_r114_c103 bl[103] br[103] wl[114] vdd gnd cell_6t
Xbit_r115_c103 bl[103] br[103] wl[115] vdd gnd cell_6t
Xbit_r116_c103 bl[103] br[103] wl[116] vdd gnd cell_6t
Xbit_r117_c103 bl[103] br[103] wl[117] vdd gnd cell_6t
Xbit_r118_c103 bl[103] br[103] wl[118] vdd gnd cell_6t
Xbit_r119_c103 bl[103] br[103] wl[119] vdd gnd cell_6t
Xbit_r120_c103 bl[103] br[103] wl[120] vdd gnd cell_6t
Xbit_r121_c103 bl[103] br[103] wl[121] vdd gnd cell_6t
Xbit_r122_c103 bl[103] br[103] wl[122] vdd gnd cell_6t
Xbit_r123_c103 bl[103] br[103] wl[123] vdd gnd cell_6t
Xbit_r124_c103 bl[103] br[103] wl[124] vdd gnd cell_6t
Xbit_r125_c103 bl[103] br[103] wl[125] vdd gnd cell_6t
Xbit_r126_c103 bl[103] br[103] wl[126] vdd gnd cell_6t
Xbit_r127_c103 bl[103] br[103] wl[127] vdd gnd cell_6t
Xbit_r128_c103 bl[103] br[103] wl[128] vdd gnd cell_6t
Xbit_r129_c103 bl[103] br[103] wl[129] vdd gnd cell_6t
Xbit_r130_c103 bl[103] br[103] wl[130] vdd gnd cell_6t
Xbit_r131_c103 bl[103] br[103] wl[131] vdd gnd cell_6t
Xbit_r132_c103 bl[103] br[103] wl[132] vdd gnd cell_6t
Xbit_r133_c103 bl[103] br[103] wl[133] vdd gnd cell_6t
Xbit_r134_c103 bl[103] br[103] wl[134] vdd gnd cell_6t
Xbit_r135_c103 bl[103] br[103] wl[135] vdd gnd cell_6t
Xbit_r136_c103 bl[103] br[103] wl[136] vdd gnd cell_6t
Xbit_r137_c103 bl[103] br[103] wl[137] vdd gnd cell_6t
Xbit_r138_c103 bl[103] br[103] wl[138] vdd gnd cell_6t
Xbit_r139_c103 bl[103] br[103] wl[139] vdd gnd cell_6t
Xbit_r140_c103 bl[103] br[103] wl[140] vdd gnd cell_6t
Xbit_r141_c103 bl[103] br[103] wl[141] vdd gnd cell_6t
Xbit_r142_c103 bl[103] br[103] wl[142] vdd gnd cell_6t
Xbit_r143_c103 bl[103] br[103] wl[143] vdd gnd cell_6t
Xbit_r144_c103 bl[103] br[103] wl[144] vdd gnd cell_6t
Xbit_r145_c103 bl[103] br[103] wl[145] vdd gnd cell_6t
Xbit_r146_c103 bl[103] br[103] wl[146] vdd gnd cell_6t
Xbit_r147_c103 bl[103] br[103] wl[147] vdd gnd cell_6t
Xbit_r148_c103 bl[103] br[103] wl[148] vdd gnd cell_6t
Xbit_r149_c103 bl[103] br[103] wl[149] vdd gnd cell_6t
Xbit_r150_c103 bl[103] br[103] wl[150] vdd gnd cell_6t
Xbit_r151_c103 bl[103] br[103] wl[151] vdd gnd cell_6t
Xbit_r152_c103 bl[103] br[103] wl[152] vdd gnd cell_6t
Xbit_r153_c103 bl[103] br[103] wl[153] vdd gnd cell_6t
Xbit_r154_c103 bl[103] br[103] wl[154] vdd gnd cell_6t
Xbit_r155_c103 bl[103] br[103] wl[155] vdd gnd cell_6t
Xbit_r156_c103 bl[103] br[103] wl[156] vdd gnd cell_6t
Xbit_r157_c103 bl[103] br[103] wl[157] vdd gnd cell_6t
Xbit_r158_c103 bl[103] br[103] wl[158] vdd gnd cell_6t
Xbit_r159_c103 bl[103] br[103] wl[159] vdd gnd cell_6t
Xbit_r160_c103 bl[103] br[103] wl[160] vdd gnd cell_6t
Xbit_r161_c103 bl[103] br[103] wl[161] vdd gnd cell_6t
Xbit_r162_c103 bl[103] br[103] wl[162] vdd gnd cell_6t
Xbit_r163_c103 bl[103] br[103] wl[163] vdd gnd cell_6t
Xbit_r164_c103 bl[103] br[103] wl[164] vdd gnd cell_6t
Xbit_r165_c103 bl[103] br[103] wl[165] vdd gnd cell_6t
Xbit_r166_c103 bl[103] br[103] wl[166] vdd gnd cell_6t
Xbit_r167_c103 bl[103] br[103] wl[167] vdd gnd cell_6t
Xbit_r168_c103 bl[103] br[103] wl[168] vdd gnd cell_6t
Xbit_r169_c103 bl[103] br[103] wl[169] vdd gnd cell_6t
Xbit_r170_c103 bl[103] br[103] wl[170] vdd gnd cell_6t
Xbit_r171_c103 bl[103] br[103] wl[171] vdd gnd cell_6t
Xbit_r172_c103 bl[103] br[103] wl[172] vdd gnd cell_6t
Xbit_r173_c103 bl[103] br[103] wl[173] vdd gnd cell_6t
Xbit_r174_c103 bl[103] br[103] wl[174] vdd gnd cell_6t
Xbit_r175_c103 bl[103] br[103] wl[175] vdd gnd cell_6t
Xbit_r176_c103 bl[103] br[103] wl[176] vdd gnd cell_6t
Xbit_r177_c103 bl[103] br[103] wl[177] vdd gnd cell_6t
Xbit_r178_c103 bl[103] br[103] wl[178] vdd gnd cell_6t
Xbit_r179_c103 bl[103] br[103] wl[179] vdd gnd cell_6t
Xbit_r180_c103 bl[103] br[103] wl[180] vdd gnd cell_6t
Xbit_r181_c103 bl[103] br[103] wl[181] vdd gnd cell_6t
Xbit_r182_c103 bl[103] br[103] wl[182] vdd gnd cell_6t
Xbit_r183_c103 bl[103] br[103] wl[183] vdd gnd cell_6t
Xbit_r184_c103 bl[103] br[103] wl[184] vdd gnd cell_6t
Xbit_r185_c103 bl[103] br[103] wl[185] vdd gnd cell_6t
Xbit_r186_c103 bl[103] br[103] wl[186] vdd gnd cell_6t
Xbit_r187_c103 bl[103] br[103] wl[187] vdd gnd cell_6t
Xbit_r188_c103 bl[103] br[103] wl[188] vdd gnd cell_6t
Xbit_r189_c103 bl[103] br[103] wl[189] vdd gnd cell_6t
Xbit_r190_c103 bl[103] br[103] wl[190] vdd gnd cell_6t
Xbit_r191_c103 bl[103] br[103] wl[191] vdd gnd cell_6t
Xbit_r192_c103 bl[103] br[103] wl[192] vdd gnd cell_6t
Xbit_r193_c103 bl[103] br[103] wl[193] vdd gnd cell_6t
Xbit_r194_c103 bl[103] br[103] wl[194] vdd gnd cell_6t
Xbit_r195_c103 bl[103] br[103] wl[195] vdd gnd cell_6t
Xbit_r196_c103 bl[103] br[103] wl[196] vdd gnd cell_6t
Xbit_r197_c103 bl[103] br[103] wl[197] vdd gnd cell_6t
Xbit_r198_c103 bl[103] br[103] wl[198] vdd gnd cell_6t
Xbit_r199_c103 bl[103] br[103] wl[199] vdd gnd cell_6t
Xbit_r200_c103 bl[103] br[103] wl[200] vdd gnd cell_6t
Xbit_r201_c103 bl[103] br[103] wl[201] vdd gnd cell_6t
Xbit_r202_c103 bl[103] br[103] wl[202] vdd gnd cell_6t
Xbit_r203_c103 bl[103] br[103] wl[203] vdd gnd cell_6t
Xbit_r204_c103 bl[103] br[103] wl[204] vdd gnd cell_6t
Xbit_r205_c103 bl[103] br[103] wl[205] vdd gnd cell_6t
Xbit_r206_c103 bl[103] br[103] wl[206] vdd gnd cell_6t
Xbit_r207_c103 bl[103] br[103] wl[207] vdd gnd cell_6t
Xbit_r208_c103 bl[103] br[103] wl[208] vdd gnd cell_6t
Xbit_r209_c103 bl[103] br[103] wl[209] vdd gnd cell_6t
Xbit_r210_c103 bl[103] br[103] wl[210] vdd gnd cell_6t
Xbit_r211_c103 bl[103] br[103] wl[211] vdd gnd cell_6t
Xbit_r212_c103 bl[103] br[103] wl[212] vdd gnd cell_6t
Xbit_r213_c103 bl[103] br[103] wl[213] vdd gnd cell_6t
Xbit_r214_c103 bl[103] br[103] wl[214] vdd gnd cell_6t
Xbit_r215_c103 bl[103] br[103] wl[215] vdd gnd cell_6t
Xbit_r216_c103 bl[103] br[103] wl[216] vdd gnd cell_6t
Xbit_r217_c103 bl[103] br[103] wl[217] vdd gnd cell_6t
Xbit_r218_c103 bl[103] br[103] wl[218] vdd gnd cell_6t
Xbit_r219_c103 bl[103] br[103] wl[219] vdd gnd cell_6t
Xbit_r220_c103 bl[103] br[103] wl[220] vdd gnd cell_6t
Xbit_r221_c103 bl[103] br[103] wl[221] vdd gnd cell_6t
Xbit_r222_c103 bl[103] br[103] wl[222] vdd gnd cell_6t
Xbit_r223_c103 bl[103] br[103] wl[223] vdd gnd cell_6t
Xbit_r224_c103 bl[103] br[103] wl[224] vdd gnd cell_6t
Xbit_r225_c103 bl[103] br[103] wl[225] vdd gnd cell_6t
Xbit_r226_c103 bl[103] br[103] wl[226] vdd gnd cell_6t
Xbit_r227_c103 bl[103] br[103] wl[227] vdd gnd cell_6t
Xbit_r228_c103 bl[103] br[103] wl[228] vdd gnd cell_6t
Xbit_r229_c103 bl[103] br[103] wl[229] vdd gnd cell_6t
Xbit_r230_c103 bl[103] br[103] wl[230] vdd gnd cell_6t
Xbit_r231_c103 bl[103] br[103] wl[231] vdd gnd cell_6t
Xbit_r232_c103 bl[103] br[103] wl[232] vdd gnd cell_6t
Xbit_r233_c103 bl[103] br[103] wl[233] vdd gnd cell_6t
Xbit_r234_c103 bl[103] br[103] wl[234] vdd gnd cell_6t
Xbit_r235_c103 bl[103] br[103] wl[235] vdd gnd cell_6t
Xbit_r236_c103 bl[103] br[103] wl[236] vdd gnd cell_6t
Xbit_r237_c103 bl[103] br[103] wl[237] vdd gnd cell_6t
Xbit_r238_c103 bl[103] br[103] wl[238] vdd gnd cell_6t
Xbit_r239_c103 bl[103] br[103] wl[239] vdd gnd cell_6t
Xbit_r240_c103 bl[103] br[103] wl[240] vdd gnd cell_6t
Xbit_r241_c103 bl[103] br[103] wl[241] vdd gnd cell_6t
Xbit_r242_c103 bl[103] br[103] wl[242] vdd gnd cell_6t
Xbit_r243_c103 bl[103] br[103] wl[243] vdd gnd cell_6t
Xbit_r244_c103 bl[103] br[103] wl[244] vdd gnd cell_6t
Xbit_r245_c103 bl[103] br[103] wl[245] vdd gnd cell_6t
Xbit_r246_c103 bl[103] br[103] wl[246] vdd gnd cell_6t
Xbit_r247_c103 bl[103] br[103] wl[247] vdd gnd cell_6t
Xbit_r248_c103 bl[103] br[103] wl[248] vdd gnd cell_6t
Xbit_r249_c103 bl[103] br[103] wl[249] vdd gnd cell_6t
Xbit_r250_c103 bl[103] br[103] wl[250] vdd gnd cell_6t
Xbit_r251_c103 bl[103] br[103] wl[251] vdd gnd cell_6t
Xbit_r252_c103 bl[103] br[103] wl[252] vdd gnd cell_6t
Xbit_r253_c103 bl[103] br[103] wl[253] vdd gnd cell_6t
Xbit_r254_c103 bl[103] br[103] wl[254] vdd gnd cell_6t
Xbit_r255_c103 bl[103] br[103] wl[255] vdd gnd cell_6t
Xbit_r0_c104 bl[104] br[104] wl[0] vdd gnd cell_6t
Xbit_r1_c104 bl[104] br[104] wl[1] vdd gnd cell_6t
Xbit_r2_c104 bl[104] br[104] wl[2] vdd gnd cell_6t
Xbit_r3_c104 bl[104] br[104] wl[3] vdd gnd cell_6t
Xbit_r4_c104 bl[104] br[104] wl[4] vdd gnd cell_6t
Xbit_r5_c104 bl[104] br[104] wl[5] vdd gnd cell_6t
Xbit_r6_c104 bl[104] br[104] wl[6] vdd gnd cell_6t
Xbit_r7_c104 bl[104] br[104] wl[7] vdd gnd cell_6t
Xbit_r8_c104 bl[104] br[104] wl[8] vdd gnd cell_6t
Xbit_r9_c104 bl[104] br[104] wl[9] vdd gnd cell_6t
Xbit_r10_c104 bl[104] br[104] wl[10] vdd gnd cell_6t
Xbit_r11_c104 bl[104] br[104] wl[11] vdd gnd cell_6t
Xbit_r12_c104 bl[104] br[104] wl[12] vdd gnd cell_6t
Xbit_r13_c104 bl[104] br[104] wl[13] vdd gnd cell_6t
Xbit_r14_c104 bl[104] br[104] wl[14] vdd gnd cell_6t
Xbit_r15_c104 bl[104] br[104] wl[15] vdd gnd cell_6t
Xbit_r16_c104 bl[104] br[104] wl[16] vdd gnd cell_6t
Xbit_r17_c104 bl[104] br[104] wl[17] vdd gnd cell_6t
Xbit_r18_c104 bl[104] br[104] wl[18] vdd gnd cell_6t
Xbit_r19_c104 bl[104] br[104] wl[19] vdd gnd cell_6t
Xbit_r20_c104 bl[104] br[104] wl[20] vdd gnd cell_6t
Xbit_r21_c104 bl[104] br[104] wl[21] vdd gnd cell_6t
Xbit_r22_c104 bl[104] br[104] wl[22] vdd gnd cell_6t
Xbit_r23_c104 bl[104] br[104] wl[23] vdd gnd cell_6t
Xbit_r24_c104 bl[104] br[104] wl[24] vdd gnd cell_6t
Xbit_r25_c104 bl[104] br[104] wl[25] vdd gnd cell_6t
Xbit_r26_c104 bl[104] br[104] wl[26] vdd gnd cell_6t
Xbit_r27_c104 bl[104] br[104] wl[27] vdd gnd cell_6t
Xbit_r28_c104 bl[104] br[104] wl[28] vdd gnd cell_6t
Xbit_r29_c104 bl[104] br[104] wl[29] vdd gnd cell_6t
Xbit_r30_c104 bl[104] br[104] wl[30] vdd gnd cell_6t
Xbit_r31_c104 bl[104] br[104] wl[31] vdd gnd cell_6t
Xbit_r32_c104 bl[104] br[104] wl[32] vdd gnd cell_6t
Xbit_r33_c104 bl[104] br[104] wl[33] vdd gnd cell_6t
Xbit_r34_c104 bl[104] br[104] wl[34] vdd gnd cell_6t
Xbit_r35_c104 bl[104] br[104] wl[35] vdd gnd cell_6t
Xbit_r36_c104 bl[104] br[104] wl[36] vdd gnd cell_6t
Xbit_r37_c104 bl[104] br[104] wl[37] vdd gnd cell_6t
Xbit_r38_c104 bl[104] br[104] wl[38] vdd gnd cell_6t
Xbit_r39_c104 bl[104] br[104] wl[39] vdd gnd cell_6t
Xbit_r40_c104 bl[104] br[104] wl[40] vdd gnd cell_6t
Xbit_r41_c104 bl[104] br[104] wl[41] vdd gnd cell_6t
Xbit_r42_c104 bl[104] br[104] wl[42] vdd gnd cell_6t
Xbit_r43_c104 bl[104] br[104] wl[43] vdd gnd cell_6t
Xbit_r44_c104 bl[104] br[104] wl[44] vdd gnd cell_6t
Xbit_r45_c104 bl[104] br[104] wl[45] vdd gnd cell_6t
Xbit_r46_c104 bl[104] br[104] wl[46] vdd gnd cell_6t
Xbit_r47_c104 bl[104] br[104] wl[47] vdd gnd cell_6t
Xbit_r48_c104 bl[104] br[104] wl[48] vdd gnd cell_6t
Xbit_r49_c104 bl[104] br[104] wl[49] vdd gnd cell_6t
Xbit_r50_c104 bl[104] br[104] wl[50] vdd gnd cell_6t
Xbit_r51_c104 bl[104] br[104] wl[51] vdd gnd cell_6t
Xbit_r52_c104 bl[104] br[104] wl[52] vdd gnd cell_6t
Xbit_r53_c104 bl[104] br[104] wl[53] vdd gnd cell_6t
Xbit_r54_c104 bl[104] br[104] wl[54] vdd gnd cell_6t
Xbit_r55_c104 bl[104] br[104] wl[55] vdd gnd cell_6t
Xbit_r56_c104 bl[104] br[104] wl[56] vdd gnd cell_6t
Xbit_r57_c104 bl[104] br[104] wl[57] vdd gnd cell_6t
Xbit_r58_c104 bl[104] br[104] wl[58] vdd gnd cell_6t
Xbit_r59_c104 bl[104] br[104] wl[59] vdd gnd cell_6t
Xbit_r60_c104 bl[104] br[104] wl[60] vdd gnd cell_6t
Xbit_r61_c104 bl[104] br[104] wl[61] vdd gnd cell_6t
Xbit_r62_c104 bl[104] br[104] wl[62] vdd gnd cell_6t
Xbit_r63_c104 bl[104] br[104] wl[63] vdd gnd cell_6t
Xbit_r64_c104 bl[104] br[104] wl[64] vdd gnd cell_6t
Xbit_r65_c104 bl[104] br[104] wl[65] vdd gnd cell_6t
Xbit_r66_c104 bl[104] br[104] wl[66] vdd gnd cell_6t
Xbit_r67_c104 bl[104] br[104] wl[67] vdd gnd cell_6t
Xbit_r68_c104 bl[104] br[104] wl[68] vdd gnd cell_6t
Xbit_r69_c104 bl[104] br[104] wl[69] vdd gnd cell_6t
Xbit_r70_c104 bl[104] br[104] wl[70] vdd gnd cell_6t
Xbit_r71_c104 bl[104] br[104] wl[71] vdd gnd cell_6t
Xbit_r72_c104 bl[104] br[104] wl[72] vdd gnd cell_6t
Xbit_r73_c104 bl[104] br[104] wl[73] vdd gnd cell_6t
Xbit_r74_c104 bl[104] br[104] wl[74] vdd gnd cell_6t
Xbit_r75_c104 bl[104] br[104] wl[75] vdd gnd cell_6t
Xbit_r76_c104 bl[104] br[104] wl[76] vdd gnd cell_6t
Xbit_r77_c104 bl[104] br[104] wl[77] vdd gnd cell_6t
Xbit_r78_c104 bl[104] br[104] wl[78] vdd gnd cell_6t
Xbit_r79_c104 bl[104] br[104] wl[79] vdd gnd cell_6t
Xbit_r80_c104 bl[104] br[104] wl[80] vdd gnd cell_6t
Xbit_r81_c104 bl[104] br[104] wl[81] vdd gnd cell_6t
Xbit_r82_c104 bl[104] br[104] wl[82] vdd gnd cell_6t
Xbit_r83_c104 bl[104] br[104] wl[83] vdd gnd cell_6t
Xbit_r84_c104 bl[104] br[104] wl[84] vdd gnd cell_6t
Xbit_r85_c104 bl[104] br[104] wl[85] vdd gnd cell_6t
Xbit_r86_c104 bl[104] br[104] wl[86] vdd gnd cell_6t
Xbit_r87_c104 bl[104] br[104] wl[87] vdd gnd cell_6t
Xbit_r88_c104 bl[104] br[104] wl[88] vdd gnd cell_6t
Xbit_r89_c104 bl[104] br[104] wl[89] vdd gnd cell_6t
Xbit_r90_c104 bl[104] br[104] wl[90] vdd gnd cell_6t
Xbit_r91_c104 bl[104] br[104] wl[91] vdd gnd cell_6t
Xbit_r92_c104 bl[104] br[104] wl[92] vdd gnd cell_6t
Xbit_r93_c104 bl[104] br[104] wl[93] vdd gnd cell_6t
Xbit_r94_c104 bl[104] br[104] wl[94] vdd gnd cell_6t
Xbit_r95_c104 bl[104] br[104] wl[95] vdd gnd cell_6t
Xbit_r96_c104 bl[104] br[104] wl[96] vdd gnd cell_6t
Xbit_r97_c104 bl[104] br[104] wl[97] vdd gnd cell_6t
Xbit_r98_c104 bl[104] br[104] wl[98] vdd gnd cell_6t
Xbit_r99_c104 bl[104] br[104] wl[99] vdd gnd cell_6t
Xbit_r100_c104 bl[104] br[104] wl[100] vdd gnd cell_6t
Xbit_r101_c104 bl[104] br[104] wl[101] vdd gnd cell_6t
Xbit_r102_c104 bl[104] br[104] wl[102] vdd gnd cell_6t
Xbit_r103_c104 bl[104] br[104] wl[103] vdd gnd cell_6t
Xbit_r104_c104 bl[104] br[104] wl[104] vdd gnd cell_6t
Xbit_r105_c104 bl[104] br[104] wl[105] vdd gnd cell_6t
Xbit_r106_c104 bl[104] br[104] wl[106] vdd gnd cell_6t
Xbit_r107_c104 bl[104] br[104] wl[107] vdd gnd cell_6t
Xbit_r108_c104 bl[104] br[104] wl[108] vdd gnd cell_6t
Xbit_r109_c104 bl[104] br[104] wl[109] vdd gnd cell_6t
Xbit_r110_c104 bl[104] br[104] wl[110] vdd gnd cell_6t
Xbit_r111_c104 bl[104] br[104] wl[111] vdd gnd cell_6t
Xbit_r112_c104 bl[104] br[104] wl[112] vdd gnd cell_6t
Xbit_r113_c104 bl[104] br[104] wl[113] vdd gnd cell_6t
Xbit_r114_c104 bl[104] br[104] wl[114] vdd gnd cell_6t
Xbit_r115_c104 bl[104] br[104] wl[115] vdd gnd cell_6t
Xbit_r116_c104 bl[104] br[104] wl[116] vdd gnd cell_6t
Xbit_r117_c104 bl[104] br[104] wl[117] vdd gnd cell_6t
Xbit_r118_c104 bl[104] br[104] wl[118] vdd gnd cell_6t
Xbit_r119_c104 bl[104] br[104] wl[119] vdd gnd cell_6t
Xbit_r120_c104 bl[104] br[104] wl[120] vdd gnd cell_6t
Xbit_r121_c104 bl[104] br[104] wl[121] vdd gnd cell_6t
Xbit_r122_c104 bl[104] br[104] wl[122] vdd gnd cell_6t
Xbit_r123_c104 bl[104] br[104] wl[123] vdd gnd cell_6t
Xbit_r124_c104 bl[104] br[104] wl[124] vdd gnd cell_6t
Xbit_r125_c104 bl[104] br[104] wl[125] vdd gnd cell_6t
Xbit_r126_c104 bl[104] br[104] wl[126] vdd gnd cell_6t
Xbit_r127_c104 bl[104] br[104] wl[127] vdd gnd cell_6t
Xbit_r128_c104 bl[104] br[104] wl[128] vdd gnd cell_6t
Xbit_r129_c104 bl[104] br[104] wl[129] vdd gnd cell_6t
Xbit_r130_c104 bl[104] br[104] wl[130] vdd gnd cell_6t
Xbit_r131_c104 bl[104] br[104] wl[131] vdd gnd cell_6t
Xbit_r132_c104 bl[104] br[104] wl[132] vdd gnd cell_6t
Xbit_r133_c104 bl[104] br[104] wl[133] vdd gnd cell_6t
Xbit_r134_c104 bl[104] br[104] wl[134] vdd gnd cell_6t
Xbit_r135_c104 bl[104] br[104] wl[135] vdd gnd cell_6t
Xbit_r136_c104 bl[104] br[104] wl[136] vdd gnd cell_6t
Xbit_r137_c104 bl[104] br[104] wl[137] vdd gnd cell_6t
Xbit_r138_c104 bl[104] br[104] wl[138] vdd gnd cell_6t
Xbit_r139_c104 bl[104] br[104] wl[139] vdd gnd cell_6t
Xbit_r140_c104 bl[104] br[104] wl[140] vdd gnd cell_6t
Xbit_r141_c104 bl[104] br[104] wl[141] vdd gnd cell_6t
Xbit_r142_c104 bl[104] br[104] wl[142] vdd gnd cell_6t
Xbit_r143_c104 bl[104] br[104] wl[143] vdd gnd cell_6t
Xbit_r144_c104 bl[104] br[104] wl[144] vdd gnd cell_6t
Xbit_r145_c104 bl[104] br[104] wl[145] vdd gnd cell_6t
Xbit_r146_c104 bl[104] br[104] wl[146] vdd gnd cell_6t
Xbit_r147_c104 bl[104] br[104] wl[147] vdd gnd cell_6t
Xbit_r148_c104 bl[104] br[104] wl[148] vdd gnd cell_6t
Xbit_r149_c104 bl[104] br[104] wl[149] vdd gnd cell_6t
Xbit_r150_c104 bl[104] br[104] wl[150] vdd gnd cell_6t
Xbit_r151_c104 bl[104] br[104] wl[151] vdd gnd cell_6t
Xbit_r152_c104 bl[104] br[104] wl[152] vdd gnd cell_6t
Xbit_r153_c104 bl[104] br[104] wl[153] vdd gnd cell_6t
Xbit_r154_c104 bl[104] br[104] wl[154] vdd gnd cell_6t
Xbit_r155_c104 bl[104] br[104] wl[155] vdd gnd cell_6t
Xbit_r156_c104 bl[104] br[104] wl[156] vdd gnd cell_6t
Xbit_r157_c104 bl[104] br[104] wl[157] vdd gnd cell_6t
Xbit_r158_c104 bl[104] br[104] wl[158] vdd gnd cell_6t
Xbit_r159_c104 bl[104] br[104] wl[159] vdd gnd cell_6t
Xbit_r160_c104 bl[104] br[104] wl[160] vdd gnd cell_6t
Xbit_r161_c104 bl[104] br[104] wl[161] vdd gnd cell_6t
Xbit_r162_c104 bl[104] br[104] wl[162] vdd gnd cell_6t
Xbit_r163_c104 bl[104] br[104] wl[163] vdd gnd cell_6t
Xbit_r164_c104 bl[104] br[104] wl[164] vdd gnd cell_6t
Xbit_r165_c104 bl[104] br[104] wl[165] vdd gnd cell_6t
Xbit_r166_c104 bl[104] br[104] wl[166] vdd gnd cell_6t
Xbit_r167_c104 bl[104] br[104] wl[167] vdd gnd cell_6t
Xbit_r168_c104 bl[104] br[104] wl[168] vdd gnd cell_6t
Xbit_r169_c104 bl[104] br[104] wl[169] vdd gnd cell_6t
Xbit_r170_c104 bl[104] br[104] wl[170] vdd gnd cell_6t
Xbit_r171_c104 bl[104] br[104] wl[171] vdd gnd cell_6t
Xbit_r172_c104 bl[104] br[104] wl[172] vdd gnd cell_6t
Xbit_r173_c104 bl[104] br[104] wl[173] vdd gnd cell_6t
Xbit_r174_c104 bl[104] br[104] wl[174] vdd gnd cell_6t
Xbit_r175_c104 bl[104] br[104] wl[175] vdd gnd cell_6t
Xbit_r176_c104 bl[104] br[104] wl[176] vdd gnd cell_6t
Xbit_r177_c104 bl[104] br[104] wl[177] vdd gnd cell_6t
Xbit_r178_c104 bl[104] br[104] wl[178] vdd gnd cell_6t
Xbit_r179_c104 bl[104] br[104] wl[179] vdd gnd cell_6t
Xbit_r180_c104 bl[104] br[104] wl[180] vdd gnd cell_6t
Xbit_r181_c104 bl[104] br[104] wl[181] vdd gnd cell_6t
Xbit_r182_c104 bl[104] br[104] wl[182] vdd gnd cell_6t
Xbit_r183_c104 bl[104] br[104] wl[183] vdd gnd cell_6t
Xbit_r184_c104 bl[104] br[104] wl[184] vdd gnd cell_6t
Xbit_r185_c104 bl[104] br[104] wl[185] vdd gnd cell_6t
Xbit_r186_c104 bl[104] br[104] wl[186] vdd gnd cell_6t
Xbit_r187_c104 bl[104] br[104] wl[187] vdd gnd cell_6t
Xbit_r188_c104 bl[104] br[104] wl[188] vdd gnd cell_6t
Xbit_r189_c104 bl[104] br[104] wl[189] vdd gnd cell_6t
Xbit_r190_c104 bl[104] br[104] wl[190] vdd gnd cell_6t
Xbit_r191_c104 bl[104] br[104] wl[191] vdd gnd cell_6t
Xbit_r192_c104 bl[104] br[104] wl[192] vdd gnd cell_6t
Xbit_r193_c104 bl[104] br[104] wl[193] vdd gnd cell_6t
Xbit_r194_c104 bl[104] br[104] wl[194] vdd gnd cell_6t
Xbit_r195_c104 bl[104] br[104] wl[195] vdd gnd cell_6t
Xbit_r196_c104 bl[104] br[104] wl[196] vdd gnd cell_6t
Xbit_r197_c104 bl[104] br[104] wl[197] vdd gnd cell_6t
Xbit_r198_c104 bl[104] br[104] wl[198] vdd gnd cell_6t
Xbit_r199_c104 bl[104] br[104] wl[199] vdd gnd cell_6t
Xbit_r200_c104 bl[104] br[104] wl[200] vdd gnd cell_6t
Xbit_r201_c104 bl[104] br[104] wl[201] vdd gnd cell_6t
Xbit_r202_c104 bl[104] br[104] wl[202] vdd gnd cell_6t
Xbit_r203_c104 bl[104] br[104] wl[203] vdd gnd cell_6t
Xbit_r204_c104 bl[104] br[104] wl[204] vdd gnd cell_6t
Xbit_r205_c104 bl[104] br[104] wl[205] vdd gnd cell_6t
Xbit_r206_c104 bl[104] br[104] wl[206] vdd gnd cell_6t
Xbit_r207_c104 bl[104] br[104] wl[207] vdd gnd cell_6t
Xbit_r208_c104 bl[104] br[104] wl[208] vdd gnd cell_6t
Xbit_r209_c104 bl[104] br[104] wl[209] vdd gnd cell_6t
Xbit_r210_c104 bl[104] br[104] wl[210] vdd gnd cell_6t
Xbit_r211_c104 bl[104] br[104] wl[211] vdd gnd cell_6t
Xbit_r212_c104 bl[104] br[104] wl[212] vdd gnd cell_6t
Xbit_r213_c104 bl[104] br[104] wl[213] vdd gnd cell_6t
Xbit_r214_c104 bl[104] br[104] wl[214] vdd gnd cell_6t
Xbit_r215_c104 bl[104] br[104] wl[215] vdd gnd cell_6t
Xbit_r216_c104 bl[104] br[104] wl[216] vdd gnd cell_6t
Xbit_r217_c104 bl[104] br[104] wl[217] vdd gnd cell_6t
Xbit_r218_c104 bl[104] br[104] wl[218] vdd gnd cell_6t
Xbit_r219_c104 bl[104] br[104] wl[219] vdd gnd cell_6t
Xbit_r220_c104 bl[104] br[104] wl[220] vdd gnd cell_6t
Xbit_r221_c104 bl[104] br[104] wl[221] vdd gnd cell_6t
Xbit_r222_c104 bl[104] br[104] wl[222] vdd gnd cell_6t
Xbit_r223_c104 bl[104] br[104] wl[223] vdd gnd cell_6t
Xbit_r224_c104 bl[104] br[104] wl[224] vdd gnd cell_6t
Xbit_r225_c104 bl[104] br[104] wl[225] vdd gnd cell_6t
Xbit_r226_c104 bl[104] br[104] wl[226] vdd gnd cell_6t
Xbit_r227_c104 bl[104] br[104] wl[227] vdd gnd cell_6t
Xbit_r228_c104 bl[104] br[104] wl[228] vdd gnd cell_6t
Xbit_r229_c104 bl[104] br[104] wl[229] vdd gnd cell_6t
Xbit_r230_c104 bl[104] br[104] wl[230] vdd gnd cell_6t
Xbit_r231_c104 bl[104] br[104] wl[231] vdd gnd cell_6t
Xbit_r232_c104 bl[104] br[104] wl[232] vdd gnd cell_6t
Xbit_r233_c104 bl[104] br[104] wl[233] vdd gnd cell_6t
Xbit_r234_c104 bl[104] br[104] wl[234] vdd gnd cell_6t
Xbit_r235_c104 bl[104] br[104] wl[235] vdd gnd cell_6t
Xbit_r236_c104 bl[104] br[104] wl[236] vdd gnd cell_6t
Xbit_r237_c104 bl[104] br[104] wl[237] vdd gnd cell_6t
Xbit_r238_c104 bl[104] br[104] wl[238] vdd gnd cell_6t
Xbit_r239_c104 bl[104] br[104] wl[239] vdd gnd cell_6t
Xbit_r240_c104 bl[104] br[104] wl[240] vdd gnd cell_6t
Xbit_r241_c104 bl[104] br[104] wl[241] vdd gnd cell_6t
Xbit_r242_c104 bl[104] br[104] wl[242] vdd gnd cell_6t
Xbit_r243_c104 bl[104] br[104] wl[243] vdd gnd cell_6t
Xbit_r244_c104 bl[104] br[104] wl[244] vdd gnd cell_6t
Xbit_r245_c104 bl[104] br[104] wl[245] vdd gnd cell_6t
Xbit_r246_c104 bl[104] br[104] wl[246] vdd gnd cell_6t
Xbit_r247_c104 bl[104] br[104] wl[247] vdd gnd cell_6t
Xbit_r248_c104 bl[104] br[104] wl[248] vdd gnd cell_6t
Xbit_r249_c104 bl[104] br[104] wl[249] vdd gnd cell_6t
Xbit_r250_c104 bl[104] br[104] wl[250] vdd gnd cell_6t
Xbit_r251_c104 bl[104] br[104] wl[251] vdd gnd cell_6t
Xbit_r252_c104 bl[104] br[104] wl[252] vdd gnd cell_6t
Xbit_r253_c104 bl[104] br[104] wl[253] vdd gnd cell_6t
Xbit_r254_c104 bl[104] br[104] wl[254] vdd gnd cell_6t
Xbit_r255_c104 bl[104] br[104] wl[255] vdd gnd cell_6t
Xbit_r0_c105 bl[105] br[105] wl[0] vdd gnd cell_6t
Xbit_r1_c105 bl[105] br[105] wl[1] vdd gnd cell_6t
Xbit_r2_c105 bl[105] br[105] wl[2] vdd gnd cell_6t
Xbit_r3_c105 bl[105] br[105] wl[3] vdd gnd cell_6t
Xbit_r4_c105 bl[105] br[105] wl[4] vdd gnd cell_6t
Xbit_r5_c105 bl[105] br[105] wl[5] vdd gnd cell_6t
Xbit_r6_c105 bl[105] br[105] wl[6] vdd gnd cell_6t
Xbit_r7_c105 bl[105] br[105] wl[7] vdd gnd cell_6t
Xbit_r8_c105 bl[105] br[105] wl[8] vdd gnd cell_6t
Xbit_r9_c105 bl[105] br[105] wl[9] vdd gnd cell_6t
Xbit_r10_c105 bl[105] br[105] wl[10] vdd gnd cell_6t
Xbit_r11_c105 bl[105] br[105] wl[11] vdd gnd cell_6t
Xbit_r12_c105 bl[105] br[105] wl[12] vdd gnd cell_6t
Xbit_r13_c105 bl[105] br[105] wl[13] vdd gnd cell_6t
Xbit_r14_c105 bl[105] br[105] wl[14] vdd gnd cell_6t
Xbit_r15_c105 bl[105] br[105] wl[15] vdd gnd cell_6t
Xbit_r16_c105 bl[105] br[105] wl[16] vdd gnd cell_6t
Xbit_r17_c105 bl[105] br[105] wl[17] vdd gnd cell_6t
Xbit_r18_c105 bl[105] br[105] wl[18] vdd gnd cell_6t
Xbit_r19_c105 bl[105] br[105] wl[19] vdd gnd cell_6t
Xbit_r20_c105 bl[105] br[105] wl[20] vdd gnd cell_6t
Xbit_r21_c105 bl[105] br[105] wl[21] vdd gnd cell_6t
Xbit_r22_c105 bl[105] br[105] wl[22] vdd gnd cell_6t
Xbit_r23_c105 bl[105] br[105] wl[23] vdd gnd cell_6t
Xbit_r24_c105 bl[105] br[105] wl[24] vdd gnd cell_6t
Xbit_r25_c105 bl[105] br[105] wl[25] vdd gnd cell_6t
Xbit_r26_c105 bl[105] br[105] wl[26] vdd gnd cell_6t
Xbit_r27_c105 bl[105] br[105] wl[27] vdd gnd cell_6t
Xbit_r28_c105 bl[105] br[105] wl[28] vdd gnd cell_6t
Xbit_r29_c105 bl[105] br[105] wl[29] vdd gnd cell_6t
Xbit_r30_c105 bl[105] br[105] wl[30] vdd gnd cell_6t
Xbit_r31_c105 bl[105] br[105] wl[31] vdd gnd cell_6t
Xbit_r32_c105 bl[105] br[105] wl[32] vdd gnd cell_6t
Xbit_r33_c105 bl[105] br[105] wl[33] vdd gnd cell_6t
Xbit_r34_c105 bl[105] br[105] wl[34] vdd gnd cell_6t
Xbit_r35_c105 bl[105] br[105] wl[35] vdd gnd cell_6t
Xbit_r36_c105 bl[105] br[105] wl[36] vdd gnd cell_6t
Xbit_r37_c105 bl[105] br[105] wl[37] vdd gnd cell_6t
Xbit_r38_c105 bl[105] br[105] wl[38] vdd gnd cell_6t
Xbit_r39_c105 bl[105] br[105] wl[39] vdd gnd cell_6t
Xbit_r40_c105 bl[105] br[105] wl[40] vdd gnd cell_6t
Xbit_r41_c105 bl[105] br[105] wl[41] vdd gnd cell_6t
Xbit_r42_c105 bl[105] br[105] wl[42] vdd gnd cell_6t
Xbit_r43_c105 bl[105] br[105] wl[43] vdd gnd cell_6t
Xbit_r44_c105 bl[105] br[105] wl[44] vdd gnd cell_6t
Xbit_r45_c105 bl[105] br[105] wl[45] vdd gnd cell_6t
Xbit_r46_c105 bl[105] br[105] wl[46] vdd gnd cell_6t
Xbit_r47_c105 bl[105] br[105] wl[47] vdd gnd cell_6t
Xbit_r48_c105 bl[105] br[105] wl[48] vdd gnd cell_6t
Xbit_r49_c105 bl[105] br[105] wl[49] vdd gnd cell_6t
Xbit_r50_c105 bl[105] br[105] wl[50] vdd gnd cell_6t
Xbit_r51_c105 bl[105] br[105] wl[51] vdd gnd cell_6t
Xbit_r52_c105 bl[105] br[105] wl[52] vdd gnd cell_6t
Xbit_r53_c105 bl[105] br[105] wl[53] vdd gnd cell_6t
Xbit_r54_c105 bl[105] br[105] wl[54] vdd gnd cell_6t
Xbit_r55_c105 bl[105] br[105] wl[55] vdd gnd cell_6t
Xbit_r56_c105 bl[105] br[105] wl[56] vdd gnd cell_6t
Xbit_r57_c105 bl[105] br[105] wl[57] vdd gnd cell_6t
Xbit_r58_c105 bl[105] br[105] wl[58] vdd gnd cell_6t
Xbit_r59_c105 bl[105] br[105] wl[59] vdd gnd cell_6t
Xbit_r60_c105 bl[105] br[105] wl[60] vdd gnd cell_6t
Xbit_r61_c105 bl[105] br[105] wl[61] vdd gnd cell_6t
Xbit_r62_c105 bl[105] br[105] wl[62] vdd gnd cell_6t
Xbit_r63_c105 bl[105] br[105] wl[63] vdd gnd cell_6t
Xbit_r64_c105 bl[105] br[105] wl[64] vdd gnd cell_6t
Xbit_r65_c105 bl[105] br[105] wl[65] vdd gnd cell_6t
Xbit_r66_c105 bl[105] br[105] wl[66] vdd gnd cell_6t
Xbit_r67_c105 bl[105] br[105] wl[67] vdd gnd cell_6t
Xbit_r68_c105 bl[105] br[105] wl[68] vdd gnd cell_6t
Xbit_r69_c105 bl[105] br[105] wl[69] vdd gnd cell_6t
Xbit_r70_c105 bl[105] br[105] wl[70] vdd gnd cell_6t
Xbit_r71_c105 bl[105] br[105] wl[71] vdd gnd cell_6t
Xbit_r72_c105 bl[105] br[105] wl[72] vdd gnd cell_6t
Xbit_r73_c105 bl[105] br[105] wl[73] vdd gnd cell_6t
Xbit_r74_c105 bl[105] br[105] wl[74] vdd gnd cell_6t
Xbit_r75_c105 bl[105] br[105] wl[75] vdd gnd cell_6t
Xbit_r76_c105 bl[105] br[105] wl[76] vdd gnd cell_6t
Xbit_r77_c105 bl[105] br[105] wl[77] vdd gnd cell_6t
Xbit_r78_c105 bl[105] br[105] wl[78] vdd gnd cell_6t
Xbit_r79_c105 bl[105] br[105] wl[79] vdd gnd cell_6t
Xbit_r80_c105 bl[105] br[105] wl[80] vdd gnd cell_6t
Xbit_r81_c105 bl[105] br[105] wl[81] vdd gnd cell_6t
Xbit_r82_c105 bl[105] br[105] wl[82] vdd gnd cell_6t
Xbit_r83_c105 bl[105] br[105] wl[83] vdd gnd cell_6t
Xbit_r84_c105 bl[105] br[105] wl[84] vdd gnd cell_6t
Xbit_r85_c105 bl[105] br[105] wl[85] vdd gnd cell_6t
Xbit_r86_c105 bl[105] br[105] wl[86] vdd gnd cell_6t
Xbit_r87_c105 bl[105] br[105] wl[87] vdd gnd cell_6t
Xbit_r88_c105 bl[105] br[105] wl[88] vdd gnd cell_6t
Xbit_r89_c105 bl[105] br[105] wl[89] vdd gnd cell_6t
Xbit_r90_c105 bl[105] br[105] wl[90] vdd gnd cell_6t
Xbit_r91_c105 bl[105] br[105] wl[91] vdd gnd cell_6t
Xbit_r92_c105 bl[105] br[105] wl[92] vdd gnd cell_6t
Xbit_r93_c105 bl[105] br[105] wl[93] vdd gnd cell_6t
Xbit_r94_c105 bl[105] br[105] wl[94] vdd gnd cell_6t
Xbit_r95_c105 bl[105] br[105] wl[95] vdd gnd cell_6t
Xbit_r96_c105 bl[105] br[105] wl[96] vdd gnd cell_6t
Xbit_r97_c105 bl[105] br[105] wl[97] vdd gnd cell_6t
Xbit_r98_c105 bl[105] br[105] wl[98] vdd gnd cell_6t
Xbit_r99_c105 bl[105] br[105] wl[99] vdd gnd cell_6t
Xbit_r100_c105 bl[105] br[105] wl[100] vdd gnd cell_6t
Xbit_r101_c105 bl[105] br[105] wl[101] vdd gnd cell_6t
Xbit_r102_c105 bl[105] br[105] wl[102] vdd gnd cell_6t
Xbit_r103_c105 bl[105] br[105] wl[103] vdd gnd cell_6t
Xbit_r104_c105 bl[105] br[105] wl[104] vdd gnd cell_6t
Xbit_r105_c105 bl[105] br[105] wl[105] vdd gnd cell_6t
Xbit_r106_c105 bl[105] br[105] wl[106] vdd gnd cell_6t
Xbit_r107_c105 bl[105] br[105] wl[107] vdd gnd cell_6t
Xbit_r108_c105 bl[105] br[105] wl[108] vdd gnd cell_6t
Xbit_r109_c105 bl[105] br[105] wl[109] vdd gnd cell_6t
Xbit_r110_c105 bl[105] br[105] wl[110] vdd gnd cell_6t
Xbit_r111_c105 bl[105] br[105] wl[111] vdd gnd cell_6t
Xbit_r112_c105 bl[105] br[105] wl[112] vdd gnd cell_6t
Xbit_r113_c105 bl[105] br[105] wl[113] vdd gnd cell_6t
Xbit_r114_c105 bl[105] br[105] wl[114] vdd gnd cell_6t
Xbit_r115_c105 bl[105] br[105] wl[115] vdd gnd cell_6t
Xbit_r116_c105 bl[105] br[105] wl[116] vdd gnd cell_6t
Xbit_r117_c105 bl[105] br[105] wl[117] vdd gnd cell_6t
Xbit_r118_c105 bl[105] br[105] wl[118] vdd gnd cell_6t
Xbit_r119_c105 bl[105] br[105] wl[119] vdd gnd cell_6t
Xbit_r120_c105 bl[105] br[105] wl[120] vdd gnd cell_6t
Xbit_r121_c105 bl[105] br[105] wl[121] vdd gnd cell_6t
Xbit_r122_c105 bl[105] br[105] wl[122] vdd gnd cell_6t
Xbit_r123_c105 bl[105] br[105] wl[123] vdd gnd cell_6t
Xbit_r124_c105 bl[105] br[105] wl[124] vdd gnd cell_6t
Xbit_r125_c105 bl[105] br[105] wl[125] vdd gnd cell_6t
Xbit_r126_c105 bl[105] br[105] wl[126] vdd gnd cell_6t
Xbit_r127_c105 bl[105] br[105] wl[127] vdd gnd cell_6t
Xbit_r128_c105 bl[105] br[105] wl[128] vdd gnd cell_6t
Xbit_r129_c105 bl[105] br[105] wl[129] vdd gnd cell_6t
Xbit_r130_c105 bl[105] br[105] wl[130] vdd gnd cell_6t
Xbit_r131_c105 bl[105] br[105] wl[131] vdd gnd cell_6t
Xbit_r132_c105 bl[105] br[105] wl[132] vdd gnd cell_6t
Xbit_r133_c105 bl[105] br[105] wl[133] vdd gnd cell_6t
Xbit_r134_c105 bl[105] br[105] wl[134] vdd gnd cell_6t
Xbit_r135_c105 bl[105] br[105] wl[135] vdd gnd cell_6t
Xbit_r136_c105 bl[105] br[105] wl[136] vdd gnd cell_6t
Xbit_r137_c105 bl[105] br[105] wl[137] vdd gnd cell_6t
Xbit_r138_c105 bl[105] br[105] wl[138] vdd gnd cell_6t
Xbit_r139_c105 bl[105] br[105] wl[139] vdd gnd cell_6t
Xbit_r140_c105 bl[105] br[105] wl[140] vdd gnd cell_6t
Xbit_r141_c105 bl[105] br[105] wl[141] vdd gnd cell_6t
Xbit_r142_c105 bl[105] br[105] wl[142] vdd gnd cell_6t
Xbit_r143_c105 bl[105] br[105] wl[143] vdd gnd cell_6t
Xbit_r144_c105 bl[105] br[105] wl[144] vdd gnd cell_6t
Xbit_r145_c105 bl[105] br[105] wl[145] vdd gnd cell_6t
Xbit_r146_c105 bl[105] br[105] wl[146] vdd gnd cell_6t
Xbit_r147_c105 bl[105] br[105] wl[147] vdd gnd cell_6t
Xbit_r148_c105 bl[105] br[105] wl[148] vdd gnd cell_6t
Xbit_r149_c105 bl[105] br[105] wl[149] vdd gnd cell_6t
Xbit_r150_c105 bl[105] br[105] wl[150] vdd gnd cell_6t
Xbit_r151_c105 bl[105] br[105] wl[151] vdd gnd cell_6t
Xbit_r152_c105 bl[105] br[105] wl[152] vdd gnd cell_6t
Xbit_r153_c105 bl[105] br[105] wl[153] vdd gnd cell_6t
Xbit_r154_c105 bl[105] br[105] wl[154] vdd gnd cell_6t
Xbit_r155_c105 bl[105] br[105] wl[155] vdd gnd cell_6t
Xbit_r156_c105 bl[105] br[105] wl[156] vdd gnd cell_6t
Xbit_r157_c105 bl[105] br[105] wl[157] vdd gnd cell_6t
Xbit_r158_c105 bl[105] br[105] wl[158] vdd gnd cell_6t
Xbit_r159_c105 bl[105] br[105] wl[159] vdd gnd cell_6t
Xbit_r160_c105 bl[105] br[105] wl[160] vdd gnd cell_6t
Xbit_r161_c105 bl[105] br[105] wl[161] vdd gnd cell_6t
Xbit_r162_c105 bl[105] br[105] wl[162] vdd gnd cell_6t
Xbit_r163_c105 bl[105] br[105] wl[163] vdd gnd cell_6t
Xbit_r164_c105 bl[105] br[105] wl[164] vdd gnd cell_6t
Xbit_r165_c105 bl[105] br[105] wl[165] vdd gnd cell_6t
Xbit_r166_c105 bl[105] br[105] wl[166] vdd gnd cell_6t
Xbit_r167_c105 bl[105] br[105] wl[167] vdd gnd cell_6t
Xbit_r168_c105 bl[105] br[105] wl[168] vdd gnd cell_6t
Xbit_r169_c105 bl[105] br[105] wl[169] vdd gnd cell_6t
Xbit_r170_c105 bl[105] br[105] wl[170] vdd gnd cell_6t
Xbit_r171_c105 bl[105] br[105] wl[171] vdd gnd cell_6t
Xbit_r172_c105 bl[105] br[105] wl[172] vdd gnd cell_6t
Xbit_r173_c105 bl[105] br[105] wl[173] vdd gnd cell_6t
Xbit_r174_c105 bl[105] br[105] wl[174] vdd gnd cell_6t
Xbit_r175_c105 bl[105] br[105] wl[175] vdd gnd cell_6t
Xbit_r176_c105 bl[105] br[105] wl[176] vdd gnd cell_6t
Xbit_r177_c105 bl[105] br[105] wl[177] vdd gnd cell_6t
Xbit_r178_c105 bl[105] br[105] wl[178] vdd gnd cell_6t
Xbit_r179_c105 bl[105] br[105] wl[179] vdd gnd cell_6t
Xbit_r180_c105 bl[105] br[105] wl[180] vdd gnd cell_6t
Xbit_r181_c105 bl[105] br[105] wl[181] vdd gnd cell_6t
Xbit_r182_c105 bl[105] br[105] wl[182] vdd gnd cell_6t
Xbit_r183_c105 bl[105] br[105] wl[183] vdd gnd cell_6t
Xbit_r184_c105 bl[105] br[105] wl[184] vdd gnd cell_6t
Xbit_r185_c105 bl[105] br[105] wl[185] vdd gnd cell_6t
Xbit_r186_c105 bl[105] br[105] wl[186] vdd gnd cell_6t
Xbit_r187_c105 bl[105] br[105] wl[187] vdd gnd cell_6t
Xbit_r188_c105 bl[105] br[105] wl[188] vdd gnd cell_6t
Xbit_r189_c105 bl[105] br[105] wl[189] vdd gnd cell_6t
Xbit_r190_c105 bl[105] br[105] wl[190] vdd gnd cell_6t
Xbit_r191_c105 bl[105] br[105] wl[191] vdd gnd cell_6t
Xbit_r192_c105 bl[105] br[105] wl[192] vdd gnd cell_6t
Xbit_r193_c105 bl[105] br[105] wl[193] vdd gnd cell_6t
Xbit_r194_c105 bl[105] br[105] wl[194] vdd gnd cell_6t
Xbit_r195_c105 bl[105] br[105] wl[195] vdd gnd cell_6t
Xbit_r196_c105 bl[105] br[105] wl[196] vdd gnd cell_6t
Xbit_r197_c105 bl[105] br[105] wl[197] vdd gnd cell_6t
Xbit_r198_c105 bl[105] br[105] wl[198] vdd gnd cell_6t
Xbit_r199_c105 bl[105] br[105] wl[199] vdd gnd cell_6t
Xbit_r200_c105 bl[105] br[105] wl[200] vdd gnd cell_6t
Xbit_r201_c105 bl[105] br[105] wl[201] vdd gnd cell_6t
Xbit_r202_c105 bl[105] br[105] wl[202] vdd gnd cell_6t
Xbit_r203_c105 bl[105] br[105] wl[203] vdd gnd cell_6t
Xbit_r204_c105 bl[105] br[105] wl[204] vdd gnd cell_6t
Xbit_r205_c105 bl[105] br[105] wl[205] vdd gnd cell_6t
Xbit_r206_c105 bl[105] br[105] wl[206] vdd gnd cell_6t
Xbit_r207_c105 bl[105] br[105] wl[207] vdd gnd cell_6t
Xbit_r208_c105 bl[105] br[105] wl[208] vdd gnd cell_6t
Xbit_r209_c105 bl[105] br[105] wl[209] vdd gnd cell_6t
Xbit_r210_c105 bl[105] br[105] wl[210] vdd gnd cell_6t
Xbit_r211_c105 bl[105] br[105] wl[211] vdd gnd cell_6t
Xbit_r212_c105 bl[105] br[105] wl[212] vdd gnd cell_6t
Xbit_r213_c105 bl[105] br[105] wl[213] vdd gnd cell_6t
Xbit_r214_c105 bl[105] br[105] wl[214] vdd gnd cell_6t
Xbit_r215_c105 bl[105] br[105] wl[215] vdd gnd cell_6t
Xbit_r216_c105 bl[105] br[105] wl[216] vdd gnd cell_6t
Xbit_r217_c105 bl[105] br[105] wl[217] vdd gnd cell_6t
Xbit_r218_c105 bl[105] br[105] wl[218] vdd gnd cell_6t
Xbit_r219_c105 bl[105] br[105] wl[219] vdd gnd cell_6t
Xbit_r220_c105 bl[105] br[105] wl[220] vdd gnd cell_6t
Xbit_r221_c105 bl[105] br[105] wl[221] vdd gnd cell_6t
Xbit_r222_c105 bl[105] br[105] wl[222] vdd gnd cell_6t
Xbit_r223_c105 bl[105] br[105] wl[223] vdd gnd cell_6t
Xbit_r224_c105 bl[105] br[105] wl[224] vdd gnd cell_6t
Xbit_r225_c105 bl[105] br[105] wl[225] vdd gnd cell_6t
Xbit_r226_c105 bl[105] br[105] wl[226] vdd gnd cell_6t
Xbit_r227_c105 bl[105] br[105] wl[227] vdd gnd cell_6t
Xbit_r228_c105 bl[105] br[105] wl[228] vdd gnd cell_6t
Xbit_r229_c105 bl[105] br[105] wl[229] vdd gnd cell_6t
Xbit_r230_c105 bl[105] br[105] wl[230] vdd gnd cell_6t
Xbit_r231_c105 bl[105] br[105] wl[231] vdd gnd cell_6t
Xbit_r232_c105 bl[105] br[105] wl[232] vdd gnd cell_6t
Xbit_r233_c105 bl[105] br[105] wl[233] vdd gnd cell_6t
Xbit_r234_c105 bl[105] br[105] wl[234] vdd gnd cell_6t
Xbit_r235_c105 bl[105] br[105] wl[235] vdd gnd cell_6t
Xbit_r236_c105 bl[105] br[105] wl[236] vdd gnd cell_6t
Xbit_r237_c105 bl[105] br[105] wl[237] vdd gnd cell_6t
Xbit_r238_c105 bl[105] br[105] wl[238] vdd gnd cell_6t
Xbit_r239_c105 bl[105] br[105] wl[239] vdd gnd cell_6t
Xbit_r240_c105 bl[105] br[105] wl[240] vdd gnd cell_6t
Xbit_r241_c105 bl[105] br[105] wl[241] vdd gnd cell_6t
Xbit_r242_c105 bl[105] br[105] wl[242] vdd gnd cell_6t
Xbit_r243_c105 bl[105] br[105] wl[243] vdd gnd cell_6t
Xbit_r244_c105 bl[105] br[105] wl[244] vdd gnd cell_6t
Xbit_r245_c105 bl[105] br[105] wl[245] vdd gnd cell_6t
Xbit_r246_c105 bl[105] br[105] wl[246] vdd gnd cell_6t
Xbit_r247_c105 bl[105] br[105] wl[247] vdd gnd cell_6t
Xbit_r248_c105 bl[105] br[105] wl[248] vdd gnd cell_6t
Xbit_r249_c105 bl[105] br[105] wl[249] vdd gnd cell_6t
Xbit_r250_c105 bl[105] br[105] wl[250] vdd gnd cell_6t
Xbit_r251_c105 bl[105] br[105] wl[251] vdd gnd cell_6t
Xbit_r252_c105 bl[105] br[105] wl[252] vdd gnd cell_6t
Xbit_r253_c105 bl[105] br[105] wl[253] vdd gnd cell_6t
Xbit_r254_c105 bl[105] br[105] wl[254] vdd gnd cell_6t
Xbit_r255_c105 bl[105] br[105] wl[255] vdd gnd cell_6t
Xbit_r0_c106 bl[106] br[106] wl[0] vdd gnd cell_6t
Xbit_r1_c106 bl[106] br[106] wl[1] vdd gnd cell_6t
Xbit_r2_c106 bl[106] br[106] wl[2] vdd gnd cell_6t
Xbit_r3_c106 bl[106] br[106] wl[3] vdd gnd cell_6t
Xbit_r4_c106 bl[106] br[106] wl[4] vdd gnd cell_6t
Xbit_r5_c106 bl[106] br[106] wl[5] vdd gnd cell_6t
Xbit_r6_c106 bl[106] br[106] wl[6] vdd gnd cell_6t
Xbit_r7_c106 bl[106] br[106] wl[7] vdd gnd cell_6t
Xbit_r8_c106 bl[106] br[106] wl[8] vdd gnd cell_6t
Xbit_r9_c106 bl[106] br[106] wl[9] vdd gnd cell_6t
Xbit_r10_c106 bl[106] br[106] wl[10] vdd gnd cell_6t
Xbit_r11_c106 bl[106] br[106] wl[11] vdd gnd cell_6t
Xbit_r12_c106 bl[106] br[106] wl[12] vdd gnd cell_6t
Xbit_r13_c106 bl[106] br[106] wl[13] vdd gnd cell_6t
Xbit_r14_c106 bl[106] br[106] wl[14] vdd gnd cell_6t
Xbit_r15_c106 bl[106] br[106] wl[15] vdd gnd cell_6t
Xbit_r16_c106 bl[106] br[106] wl[16] vdd gnd cell_6t
Xbit_r17_c106 bl[106] br[106] wl[17] vdd gnd cell_6t
Xbit_r18_c106 bl[106] br[106] wl[18] vdd gnd cell_6t
Xbit_r19_c106 bl[106] br[106] wl[19] vdd gnd cell_6t
Xbit_r20_c106 bl[106] br[106] wl[20] vdd gnd cell_6t
Xbit_r21_c106 bl[106] br[106] wl[21] vdd gnd cell_6t
Xbit_r22_c106 bl[106] br[106] wl[22] vdd gnd cell_6t
Xbit_r23_c106 bl[106] br[106] wl[23] vdd gnd cell_6t
Xbit_r24_c106 bl[106] br[106] wl[24] vdd gnd cell_6t
Xbit_r25_c106 bl[106] br[106] wl[25] vdd gnd cell_6t
Xbit_r26_c106 bl[106] br[106] wl[26] vdd gnd cell_6t
Xbit_r27_c106 bl[106] br[106] wl[27] vdd gnd cell_6t
Xbit_r28_c106 bl[106] br[106] wl[28] vdd gnd cell_6t
Xbit_r29_c106 bl[106] br[106] wl[29] vdd gnd cell_6t
Xbit_r30_c106 bl[106] br[106] wl[30] vdd gnd cell_6t
Xbit_r31_c106 bl[106] br[106] wl[31] vdd gnd cell_6t
Xbit_r32_c106 bl[106] br[106] wl[32] vdd gnd cell_6t
Xbit_r33_c106 bl[106] br[106] wl[33] vdd gnd cell_6t
Xbit_r34_c106 bl[106] br[106] wl[34] vdd gnd cell_6t
Xbit_r35_c106 bl[106] br[106] wl[35] vdd gnd cell_6t
Xbit_r36_c106 bl[106] br[106] wl[36] vdd gnd cell_6t
Xbit_r37_c106 bl[106] br[106] wl[37] vdd gnd cell_6t
Xbit_r38_c106 bl[106] br[106] wl[38] vdd gnd cell_6t
Xbit_r39_c106 bl[106] br[106] wl[39] vdd gnd cell_6t
Xbit_r40_c106 bl[106] br[106] wl[40] vdd gnd cell_6t
Xbit_r41_c106 bl[106] br[106] wl[41] vdd gnd cell_6t
Xbit_r42_c106 bl[106] br[106] wl[42] vdd gnd cell_6t
Xbit_r43_c106 bl[106] br[106] wl[43] vdd gnd cell_6t
Xbit_r44_c106 bl[106] br[106] wl[44] vdd gnd cell_6t
Xbit_r45_c106 bl[106] br[106] wl[45] vdd gnd cell_6t
Xbit_r46_c106 bl[106] br[106] wl[46] vdd gnd cell_6t
Xbit_r47_c106 bl[106] br[106] wl[47] vdd gnd cell_6t
Xbit_r48_c106 bl[106] br[106] wl[48] vdd gnd cell_6t
Xbit_r49_c106 bl[106] br[106] wl[49] vdd gnd cell_6t
Xbit_r50_c106 bl[106] br[106] wl[50] vdd gnd cell_6t
Xbit_r51_c106 bl[106] br[106] wl[51] vdd gnd cell_6t
Xbit_r52_c106 bl[106] br[106] wl[52] vdd gnd cell_6t
Xbit_r53_c106 bl[106] br[106] wl[53] vdd gnd cell_6t
Xbit_r54_c106 bl[106] br[106] wl[54] vdd gnd cell_6t
Xbit_r55_c106 bl[106] br[106] wl[55] vdd gnd cell_6t
Xbit_r56_c106 bl[106] br[106] wl[56] vdd gnd cell_6t
Xbit_r57_c106 bl[106] br[106] wl[57] vdd gnd cell_6t
Xbit_r58_c106 bl[106] br[106] wl[58] vdd gnd cell_6t
Xbit_r59_c106 bl[106] br[106] wl[59] vdd gnd cell_6t
Xbit_r60_c106 bl[106] br[106] wl[60] vdd gnd cell_6t
Xbit_r61_c106 bl[106] br[106] wl[61] vdd gnd cell_6t
Xbit_r62_c106 bl[106] br[106] wl[62] vdd gnd cell_6t
Xbit_r63_c106 bl[106] br[106] wl[63] vdd gnd cell_6t
Xbit_r64_c106 bl[106] br[106] wl[64] vdd gnd cell_6t
Xbit_r65_c106 bl[106] br[106] wl[65] vdd gnd cell_6t
Xbit_r66_c106 bl[106] br[106] wl[66] vdd gnd cell_6t
Xbit_r67_c106 bl[106] br[106] wl[67] vdd gnd cell_6t
Xbit_r68_c106 bl[106] br[106] wl[68] vdd gnd cell_6t
Xbit_r69_c106 bl[106] br[106] wl[69] vdd gnd cell_6t
Xbit_r70_c106 bl[106] br[106] wl[70] vdd gnd cell_6t
Xbit_r71_c106 bl[106] br[106] wl[71] vdd gnd cell_6t
Xbit_r72_c106 bl[106] br[106] wl[72] vdd gnd cell_6t
Xbit_r73_c106 bl[106] br[106] wl[73] vdd gnd cell_6t
Xbit_r74_c106 bl[106] br[106] wl[74] vdd gnd cell_6t
Xbit_r75_c106 bl[106] br[106] wl[75] vdd gnd cell_6t
Xbit_r76_c106 bl[106] br[106] wl[76] vdd gnd cell_6t
Xbit_r77_c106 bl[106] br[106] wl[77] vdd gnd cell_6t
Xbit_r78_c106 bl[106] br[106] wl[78] vdd gnd cell_6t
Xbit_r79_c106 bl[106] br[106] wl[79] vdd gnd cell_6t
Xbit_r80_c106 bl[106] br[106] wl[80] vdd gnd cell_6t
Xbit_r81_c106 bl[106] br[106] wl[81] vdd gnd cell_6t
Xbit_r82_c106 bl[106] br[106] wl[82] vdd gnd cell_6t
Xbit_r83_c106 bl[106] br[106] wl[83] vdd gnd cell_6t
Xbit_r84_c106 bl[106] br[106] wl[84] vdd gnd cell_6t
Xbit_r85_c106 bl[106] br[106] wl[85] vdd gnd cell_6t
Xbit_r86_c106 bl[106] br[106] wl[86] vdd gnd cell_6t
Xbit_r87_c106 bl[106] br[106] wl[87] vdd gnd cell_6t
Xbit_r88_c106 bl[106] br[106] wl[88] vdd gnd cell_6t
Xbit_r89_c106 bl[106] br[106] wl[89] vdd gnd cell_6t
Xbit_r90_c106 bl[106] br[106] wl[90] vdd gnd cell_6t
Xbit_r91_c106 bl[106] br[106] wl[91] vdd gnd cell_6t
Xbit_r92_c106 bl[106] br[106] wl[92] vdd gnd cell_6t
Xbit_r93_c106 bl[106] br[106] wl[93] vdd gnd cell_6t
Xbit_r94_c106 bl[106] br[106] wl[94] vdd gnd cell_6t
Xbit_r95_c106 bl[106] br[106] wl[95] vdd gnd cell_6t
Xbit_r96_c106 bl[106] br[106] wl[96] vdd gnd cell_6t
Xbit_r97_c106 bl[106] br[106] wl[97] vdd gnd cell_6t
Xbit_r98_c106 bl[106] br[106] wl[98] vdd gnd cell_6t
Xbit_r99_c106 bl[106] br[106] wl[99] vdd gnd cell_6t
Xbit_r100_c106 bl[106] br[106] wl[100] vdd gnd cell_6t
Xbit_r101_c106 bl[106] br[106] wl[101] vdd gnd cell_6t
Xbit_r102_c106 bl[106] br[106] wl[102] vdd gnd cell_6t
Xbit_r103_c106 bl[106] br[106] wl[103] vdd gnd cell_6t
Xbit_r104_c106 bl[106] br[106] wl[104] vdd gnd cell_6t
Xbit_r105_c106 bl[106] br[106] wl[105] vdd gnd cell_6t
Xbit_r106_c106 bl[106] br[106] wl[106] vdd gnd cell_6t
Xbit_r107_c106 bl[106] br[106] wl[107] vdd gnd cell_6t
Xbit_r108_c106 bl[106] br[106] wl[108] vdd gnd cell_6t
Xbit_r109_c106 bl[106] br[106] wl[109] vdd gnd cell_6t
Xbit_r110_c106 bl[106] br[106] wl[110] vdd gnd cell_6t
Xbit_r111_c106 bl[106] br[106] wl[111] vdd gnd cell_6t
Xbit_r112_c106 bl[106] br[106] wl[112] vdd gnd cell_6t
Xbit_r113_c106 bl[106] br[106] wl[113] vdd gnd cell_6t
Xbit_r114_c106 bl[106] br[106] wl[114] vdd gnd cell_6t
Xbit_r115_c106 bl[106] br[106] wl[115] vdd gnd cell_6t
Xbit_r116_c106 bl[106] br[106] wl[116] vdd gnd cell_6t
Xbit_r117_c106 bl[106] br[106] wl[117] vdd gnd cell_6t
Xbit_r118_c106 bl[106] br[106] wl[118] vdd gnd cell_6t
Xbit_r119_c106 bl[106] br[106] wl[119] vdd gnd cell_6t
Xbit_r120_c106 bl[106] br[106] wl[120] vdd gnd cell_6t
Xbit_r121_c106 bl[106] br[106] wl[121] vdd gnd cell_6t
Xbit_r122_c106 bl[106] br[106] wl[122] vdd gnd cell_6t
Xbit_r123_c106 bl[106] br[106] wl[123] vdd gnd cell_6t
Xbit_r124_c106 bl[106] br[106] wl[124] vdd gnd cell_6t
Xbit_r125_c106 bl[106] br[106] wl[125] vdd gnd cell_6t
Xbit_r126_c106 bl[106] br[106] wl[126] vdd gnd cell_6t
Xbit_r127_c106 bl[106] br[106] wl[127] vdd gnd cell_6t
Xbit_r128_c106 bl[106] br[106] wl[128] vdd gnd cell_6t
Xbit_r129_c106 bl[106] br[106] wl[129] vdd gnd cell_6t
Xbit_r130_c106 bl[106] br[106] wl[130] vdd gnd cell_6t
Xbit_r131_c106 bl[106] br[106] wl[131] vdd gnd cell_6t
Xbit_r132_c106 bl[106] br[106] wl[132] vdd gnd cell_6t
Xbit_r133_c106 bl[106] br[106] wl[133] vdd gnd cell_6t
Xbit_r134_c106 bl[106] br[106] wl[134] vdd gnd cell_6t
Xbit_r135_c106 bl[106] br[106] wl[135] vdd gnd cell_6t
Xbit_r136_c106 bl[106] br[106] wl[136] vdd gnd cell_6t
Xbit_r137_c106 bl[106] br[106] wl[137] vdd gnd cell_6t
Xbit_r138_c106 bl[106] br[106] wl[138] vdd gnd cell_6t
Xbit_r139_c106 bl[106] br[106] wl[139] vdd gnd cell_6t
Xbit_r140_c106 bl[106] br[106] wl[140] vdd gnd cell_6t
Xbit_r141_c106 bl[106] br[106] wl[141] vdd gnd cell_6t
Xbit_r142_c106 bl[106] br[106] wl[142] vdd gnd cell_6t
Xbit_r143_c106 bl[106] br[106] wl[143] vdd gnd cell_6t
Xbit_r144_c106 bl[106] br[106] wl[144] vdd gnd cell_6t
Xbit_r145_c106 bl[106] br[106] wl[145] vdd gnd cell_6t
Xbit_r146_c106 bl[106] br[106] wl[146] vdd gnd cell_6t
Xbit_r147_c106 bl[106] br[106] wl[147] vdd gnd cell_6t
Xbit_r148_c106 bl[106] br[106] wl[148] vdd gnd cell_6t
Xbit_r149_c106 bl[106] br[106] wl[149] vdd gnd cell_6t
Xbit_r150_c106 bl[106] br[106] wl[150] vdd gnd cell_6t
Xbit_r151_c106 bl[106] br[106] wl[151] vdd gnd cell_6t
Xbit_r152_c106 bl[106] br[106] wl[152] vdd gnd cell_6t
Xbit_r153_c106 bl[106] br[106] wl[153] vdd gnd cell_6t
Xbit_r154_c106 bl[106] br[106] wl[154] vdd gnd cell_6t
Xbit_r155_c106 bl[106] br[106] wl[155] vdd gnd cell_6t
Xbit_r156_c106 bl[106] br[106] wl[156] vdd gnd cell_6t
Xbit_r157_c106 bl[106] br[106] wl[157] vdd gnd cell_6t
Xbit_r158_c106 bl[106] br[106] wl[158] vdd gnd cell_6t
Xbit_r159_c106 bl[106] br[106] wl[159] vdd gnd cell_6t
Xbit_r160_c106 bl[106] br[106] wl[160] vdd gnd cell_6t
Xbit_r161_c106 bl[106] br[106] wl[161] vdd gnd cell_6t
Xbit_r162_c106 bl[106] br[106] wl[162] vdd gnd cell_6t
Xbit_r163_c106 bl[106] br[106] wl[163] vdd gnd cell_6t
Xbit_r164_c106 bl[106] br[106] wl[164] vdd gnd cell_6t
Xbit_r165_c106 bl[106] br[106] wl[165] vdd gnd cell_6t
Xbit_r166_c106 bl[106] br[106] wl[166] vdd gnd cell_6t
Xbit_r167_c106 bl[106] br[106] wl[167] vdd gnd cell_6t
Xbit_r168_c106 bl[106] br[106] wl[168] vdd gnd cell_6t
Xbit_r169_c106 bl[106] br[106] wl[169] vdd gnd cell_6t
Xbit_r170_c106 bl[106] br[106] wl[170] vdd gnd cell_6t
Xbit_r171_c106 bl[106] br[106] wl[171] vdd gnd cell_6t
Xbit_r172_c106 bl[106] br[106] wl[172] vdd gnd cell_6t
Xbit_r173_c106 bl[106] br[106] wl[173] vdd gnd cell_6t
Xbit_r174_c106 bl[106] br[106] wl[174] vdd gnd cell_6t
Xbit_r175_c106 bl[106] br[106] wl[175] vdd gnd cell_6t
Xbit_r176_c106 bl[106] br[106] wl[176] vdd gnd cell_6t
Xbit_r177_c106 bl[106] br[106] wl[177] vdd gnd cell_6t
Xbit_r178_c106 bl[106] br[106] wl[178] vdd gnd cell_6t
Xbit_r179_c106 bl[106] br[106] wl[179] vdd gnd cell_6t
Xbit_r180_c106 bl[106] br[106] wl[180] vdd gnd cell_6t
Xbit_r181_c106 bl[106] br[106] wl[181] vdd gnd cell_6t
Xbit_r182_c106 bl[106] br[106] wl[182] vdd gnd cell_6t
Xbit_r183_c106 bl[106] br[106] wl[183] vdd gnd cell_6t
Xbit_r184_c106 bl[106] br[106] wl[184] vdd gnd cell_6t
Xbit_r185_c106 bl[106] br[106] wl[185] vdd gnd cell_6t
Xbit_r186_c106 bl[106] br[106] wl[186] vdd gnd cell_6t
Xbit_r187_c106 bl[106] br[106] wl[187] vdd gnd cell_6t
Xbit_r188_c106 bl[106] br[106] wl[188] vdd gnd cell_6t
Xbit_r189_c106 bl[106] br[106] wl[189] vdd gnd cell_6t
Xbit_r190_c106 bl[106] br[106] wl[190] vdd gnd cell_6t
Xbit_r191_c106 bl[106] br[106] wl[191] vdd gnd cell_6t
Xbit_r192_c106 bl[106] br[106] wl[192] vdd gnd cell_6t
Xbit_r193_c106 bl[106] br[106] wl[193] vdd gnd cell_6t
Xbit_r194_c106 bl[106] br[106] wl[194] vdd gnd cell_6t
Xbit_r195_c106 bl[106] br[106] wl[195] vdd gnd cell_6t
Xbit_r196_c106 bl[106] br[106] wl[196] vdd gnd cell_6t
Xbit_r197_c106 bl[106] br[106] wl[197] vdd gnd cell_6t
Xbit_r198_c106 bl[106] br[106] wl[198] vdd gnd cell_6t
Xbit_r199_c106 bl[106] br[106] wl[199] vdd gnd cell_6t
Xbit_r200_c106 bl[106] br[106] wl[200] vdd gnd cell_6t
Xbit_r201_c106 bl[106] br[106] wl[201] vdd gnd cell_6t
Xbit_r202_c106 bl[106] br[106] wl[202] vdd gnd cell_6t
Xbit_r203_c106 bl[106] br[106] wl[203] vdd gnd cell_6t
Xbit_r204_c106 bl[106] br[106] wl[204] vdd gnd cell_6t
Xbit_r205_c106 bl[106] br[106] wl[205] vdd gnd cell_6t
Xbit_r206_c106 bl[106] br[106] wl[206] vdd gnd cell_6t
Xbit_r207_c106 bl[106] br[106] wl[207] vdd gnd cell_6t
Xbit_r208_c106 bl[106] br[106] wl[208] vdd gnd cell_6t
Xbit_r209_c106 bl[106] br[106] wl[209] vdd gnd cell_6t
Xbit_r210_c106 bl[106] br[106] wl[210] vdd gnd cell_6t
Xbit_r211_c106 bl[106] br[106] wl[211] vdd gnd cell_6t
Xbit_r212_c106 bl[106] br[106] wl[212] vdd gnd cell_6t
Xbit_r213_c106 bl[106] br[106] wl[213] vdd gnd cell_6t
Xbit_r214_c106 bl[106] br[106] wl[214] vdd gnd cell_6t
Xbit_r215_c106 bl[106] br[106] wl[215] vdd gnd cell_6t
Xbit_r216_c106 bl[106] br[106] wl[216] vdd gnd cell_6t
Xbit_r217_c106 bl[106] br[106] wl[217] vdd gnd cell_6t
Xbit_r218_c106 bl[106] br[106] wl[218] vdd gnd cell_6t
Xbit_r219_c106 bl[106] br[106] wl[219] vdd gnd cell_6t
Xbit_r220_c106 bl[106] br[106] wl[220] vdd gnd cell_6t
Xbit_r221_c106 bl[106] br[106] wl[221] vdd gnd cell_6t
Xbit_r222_c106 bl[106] br[106] wl[222] vdd gnd cell_6t
Xbit_r223_c106 bl[106] br[106] wl[223] vdd gnd cell_6t
Xbit_r224_c106 bl[106] br[106] wl[224] vdd gnd cell_6t
Xbit_r225_c106 bl[106] br[106] wl[225] vdd gnd cell_6t
Xbit_r226_c106 bl[106] br[106] wl[226] vdd gnd cell_6t
Xbit_r227_c106 bl[106] br[106] wl[227] vdd gnd cell_6t
Xbit_r228_c106 bl[106] br[106] wl[228] vdd gnd cell_6t
Xbit_r229_c106 bl[106] br[106] wl[229] vdd gnd cell_6t
Xbit_r230_c106 bl[106] br[106] wl[230] vdd gnd cell_6t
Xbit_r231_c106 bl[106] br[106] wl[231] vdd gnd cell_6t
Xbit_r232_c106 bl[106] br[106] wl[232] vdd gnd cell_6t
Xbit_r233_c106 bl[106] br[106] wl[233] vdd gnd cell_6t
Xbit_r234_c106 bl[106] br[106] wl[234] vdd gnd cell_6t
Xbit_r235_c106 bl[106] br[106] wl[235] vdd gnd cell_6t
Xbit_r236_c106 bl[106] br[106] wl[236] vdd gnd cell_6t
Xbit_r237_c106 bl[106] br[106] wl[237] vdd gnd cell_6t
Xbit_r238_c106 bl[106] br[106] wl[238] vdd gnd cell_6t
Xbit_r239_c106 bl[106] br[106] wl[239] vdd gnd cell_6t
Xbit_r240_c106 bl[106] br[106] wl[240] vdd gnd cell_6t
Xbit_r241_c106 bl[106] br[106] wl[241] vdd gnd cell_6t
Xbit_r242_c106 bl[106] br[106] wl[242] vdd gnd cell_6t
Xbit_r243_c106 bl[106] br[106] wl[243] vdd gnd cell_6t
Xbit_r244_c106 bl[106] br[106] wl[244] vdd gnd cell_6t
Xbit_r245_c106 bl[106] br[106] wl[245] vdd gnd cell_6t
Xbit_r246_c106 bl[106] br[106] wl[246] vdd gnd cell_6t
Xbit_r247_c106 bl[106] br[106] wl[247] vdd gnd cell_6t
Xbit_r248_c106 bl[106] br[106] wl[248] vdd gnd cell_6t
Xbit_r249_c106 bl[106] br[106] wl[249] vdd gnd cell_6t
Xbit_r250_c106 bl[106] br[106] wl[250] vdd gnd cell_6t
Xbit_r251_c106 bl[106] br[106] wl[251] vdd gnd cell_6t
Xbit_r252_c106 bl[106] br[106] wl[252] vdd gnd cell_6t
Xbit_r253_c106 bl[106] br[106] wl[253] vdd gnd cell_6t
Xbit_r254_c106 bl[106] br[106] wl[254] vdd gnd cell_6t
Xbit_r255_c106 bl[106] br[106] wl[255] vdd gnd cell_6t
Xbit_r0_c107 bl[107] br[107] wl[0] vdd gnd cell_6t
Xbit_r1_c107 bl[107] br[107] wl[1] vdd gnd cell_6t
Xbit_r2_c107 bl[107] br[107] wl[2] vdd gnd cell_6t
Xbit_r3_c107 bl[107] br[107] wl[3] vdd gnd cell_6t
Xbit_r4_c107 bl[107] br[107] wl[4] vdd gnd cell_6t
Xbit_r5_c107 bl[107] br[107] wl[5] vdd gnd cell_6t
Xbit_r6_c107 bl[107] br[107] wl[6] vdd gnd cell_6t
Xbit_r7_c107 bl[107] br[107] wl[7] vdd gnd cell_6t
Xbit_r8_c107 bl[107] br[107] wl[8] vdd gnd cell_6t
Xbit_r9_c107 bl[107] br[107] wl[9] vdd gnd cell_6t
Xbit_r10_c107 bl[107] br[107] wl[10] vdd gnd cell_6t
Xbit_r11_c107 bl[107] br[107] wl[11] vdd gnd cell_6t
Xbit_r12_c107 bl[107] br[107] wl[12] vdd gnd cell_6t
Xbit_r13_c107 bl[107] br[107] wl[13] vdd gnd cell_6t
Xbit_r14_c107 bl[107] br[107] wl[14] vdd gnd cell_6t
Xbit_r15_c107 bl[107] br[107] wl[15] vdd gnd cell_6t
Xbit_r16_c107 bl[107] br[107] wl[16] vdd gnd cell_6t
Xbit_r17_c107 bl[107] br[107] wl[17] vdd gnd cell_6t
Xbit_r18_c107 bl[107] br[107] wl[18] vdd gnd cell_6t
Xbit_r19_c107 bl[107] br[107] wl[19] vdd gnd cell_6t
Xbit_r20_c107 bl[107] br[107] wl[20] vdd gnd cell_6t
Xbit_r21_c107 bl[107] br[107] wl[21] vdd gnd cell_6t
Xbit_r22_c107 bl[107] br[107] wl[22] vdd gnd cell_6t
Xbit_r23_c107 bl[107] br[107] wl[23] vdd gnd cell_6t
Xbit_r24_c107 bl[107] br[107] wl[24] vdd gnd cell_6t
Xbit_r25_c107 bl[107] br[107] wl[25] vdd gnd cell_6t
Xbit_r26_c107 bl[107] br[107] wl[26] vdd gnd cell_6t
Xbit_r27_c107 bl[107] br[107] wl[27] vdd gnd cell_6t
Xbit_r28_c107 bl[107] br[107] wl[28] vdd gnd cell_6t
Xbit_r29_c107 bl[107] br[107] wl[29] vdd gnd cell_6t
Xbit_r30_c107 bl[107] br[107] wl[30] vdd gnd cell_6t
Xbit_r31_c107 bl[107] br[107] wl[31] vdd gnd cell_6t
Xbit_r32_c107 bl[107] br[107] wl[32] vdd gnd cell_6t
Xbit_r33_c107 bl[107] br[107] wl[33] vdd gnd cell_6t
Xbit_r34_c107 bl[107] br[107] wl[34] vdd gnd cell_6t
Xbit_r35_c107 bl[107] br[107] wl[35] vdd gnd cell_6t
Xbit_r36_c107 bl[107] br[107] wl[36] vdd gnd cell_6t
Xbit_r37_c107 bl[107] br[107] wl[37] vdd gnd cell_6t
Xbit_r38_c107 bl[107] br[107] wl[38] vdd gnd cell_6t
Xbit_r39_c107 bl[107] br[107] wl[39] vdd gnd cell_6t
Xbit_r40_c107 bl[107] br[107] wl[40] vdd gnd cell_6t
Xbit_r41_c107 bl[107] br[107] wl[41] vdd gnd cell_6t
Xbit_r42_c107 bl[107] br[107] wl[42] vdd gnd cell_6t
Xbit_r43_c107 bl[107] br[107] wl[43] vdd gnd cell_6t
Xbit_r44_c107 bl[107] br[107] wl[44] vdd gnd cell_6t
Xbit_r45_c107 bl[107] br[107] wl[45] vdd gnd cell_6t
Xbit_r46_c107 bl[107] br[107] wl[46] vdd gnd cell_6t
Xbit_r47_c107 bl[107] br[107] wl[47] vdd gnd cell_6t
Xbit_r48_c107 bl[107] br[107] wl[48] vdd gnd cell_6t
Xbit_r49_c107 bl[107] br[107] wl[49] vdd gnd cell_6t
Xbit_r50_c107 bl[107] br[107] wl[50] vdd gnd cell_6t
Xbit_r51_c107 bl[107] br[107] wl[51] vdd gnd cell_6t
Xbit_r52_c107 bl[107] br[107] wl[52] vdd gnd cell_6t
Xbit_r53_c107 bl[107] br[107] wl[53] vdd gnd cell_6t
Xbit_r54_c107 bl[107] br[107] wl[54] vdd gnd cell_6t
Xbit_r55_c107 bl[107] br[107] wl[55] vdd gnd cell_6t
Xbit_r56_c107 bl[107] br[107] wl[56] vdd gnd cell_6t
Xbit_r57_c107 bl[107] br[107] wl[57] vdd gnd cell_6t
Xbit_r58_c107 bl[107] br[107] wl[58] vdd gnd cell_6t
Xbit_r59_c107 bl[107] br[107] wl[59] vdd gnd cell_6t
Xbit_r60_c107 bl[107] br[107] wl[60] vdd gnd cell_6t
Xbit_r61_c107 bl[107] br[107] wl[61] vdd gnd cell_6t
Xbit_r62_c107 bl[107] br[107] wl[62] vdd gnd cell_6t
Xbit_r63_c107 bl[107] br[107] wl[63] vdd gnd cell_6t
Xbit_r64_c107 bl[107] br[107] wl[64] vdd gnd cell_6t
Xbit_r65_c107 bl[107] br[107] wl[65] vdd gnd cell_6t
Xbit_r66_c107 bl[107] br[107] wl[66] vdd gnd cell_6t
Xbit_r67_c107 bl[107] br[107] wl[67] vdd gnd cell_6t
Xbit_r68_c107 bl[107] br[107] wl[68] vdd gnd cell_6t
Xbit_r69_c107 bl[107] br[107] wl[69] vdd gnd cell_6t
Xbit_r70_c107 bl[107] br[107] wl[70] vdd gnd cell_6t
Xbit_r71_c107 bl[107] br[107] wl[71] vdd gnd cell_6t
Xbit_r72_c107 bl[107] br[107] wl[72] vdd gnd cell_6t
Xbit_r73_c107 bl[107] br[107] wl[73] vdd gnd cell_6t
Xbit_r74_c107 bl[107] br[107] wl[74] vdd gnd cell_6t
Xbit_r75_c107 bl[107] br[107] wl[75] vdd gnd cell_6t
Xbit_r76_c107 bl[107] br[107] wl[76] vdd gnd cell_6t
Xbit_r77_c107 bl[107] br[107] wl[77] vdd gnd cell_6t
Xbit_r78_c107 bl[107] br[107] wl[78] vdd gnd cell_6t
Xbit_r79_c107 bl[107] br[107] wl[79] vdd gnd cell_6t
Xbit_r80_c107 bl[107] br[107] wl[80] vdd gnd cell_6t
Xbit_r81_c107 bl[107] br[107] wl[81] vdd gnd cell_6t
Xbit_r82_c107 bl[107] br[107] wl[82] vdd gnd cell_6t
Xbit_r83_c107 bl[107] br[107] wl[83] vdd gnd cell_6t
Xbit_r84_c107 bl[107] br[107] wl[84] vdd gnd cell_6t
Xbit_r85_c107 bl[107] br[107] wl[85] vdd gnd cell_6t
Xbit_r86_c107 bl[107] br[107] wl[86] vdd gnd cell_6t
Xbit_r87_c107 bl[107] br[107] wl[87] vdd gnd cell_6t
Xbit_r88_c107 bl[107] br[107] wl[88] vdd gnd cell_6t
Xbit_r89_c107 bl[107] br[107] wl[89] vdd gnd cell_6t
Xbit_r90_c107 bl[107] br[107] wl[90] vdd gnd cell_6t
Xbit_r91_c107 bl[107] br[107] wl[91] vdd gnd cell_6t
Xbit_r92_c107 bl[107] br[107] wl[92] vdd gnd cell_6t
Xbit_r93_c107 bl[107] br[107] wl[93] vdd gnd cell_6t
Xbit_r94_c107 bl[107] br[107] wl[94] vdd gnd cell_6t
Xbit_r95_c107 bl[107] br[107] wl[95] vdd gnd cell_6t
Xbit_r96_c107 bl[107] br[107] wl[96] vdd gnd cell_6t
Xbit_r97_c107 bl[107] br[107] wl[97] vdd gnd cell_6t
Xbit_r98_c107 bl[107] br[107] wl[98] vdd gnd cell_6t
Xbit_r99_c107 bl[107] br[107] wl[99] vdd gnd cell_6t
Xbit_r100_c107 bl[107] br[107] wl[100] vdd gnd cell_6t
Xbit_r101_c107 bl[107] br[107] wl[101] vdd gnd cell_6t
Xbit_r102_c107 bl[107] br[107] wl[102] vdd gnd cell_6t
Xbit_r103_c107 bl[107] br[107] wl[103] vdd gnd cell_6t
Xbit_r104_c107 bl[107] br[107] wl[104] vdd gnd cell_6t
Xbit_r105_c107 bl[107] br[107] wl[105] vdd gnd cell_6t
Xbit_r106_c107 bl[107] br[107] wl[106] vdd gnd cell_6t
Xbit_r107_c107 bl[107] br[107] wl[107] vdd gnd cell_6t
Xbit_r108_c107 bl[107] br[107] wl[108] vdd gnd cell_6t
Xbit_r109_c107 bl[107] br[107] wl[109] vdd gnd cell_6t
Xbit_r110_c107 bl[107] br[107] wl[110] vdd gnd cell_6t
Xbit_r111_c107 bl[107] br[107] wl[111] vdd gnd cell_6t
Xbit_r112_c107 bl[107] br[107] wl[112] vdd gnd cell_6t
Xbit_r113_c107 bl[107] br[107] wl[113] vdd gnd cell_6t
Xbit_r114_c107 bl[107] br[107] wl[114] vdd gnd cell_6t
Xbit_r115_c107 bl[107] br[107] wl[115] vdd gnd cell_6t
Xbit_r116_c107 bl[107] br[107] wl[116] vdd gnd cell_6t
Xbit_r117_c107 bl[107] br[107] wl[117] vdd gnd cell_6t
Xbit_r118_c107 bl[107] br[107] wl[118] vdd gnd cell_6t
Xbit_r119_c107 bl[107] br[107] wl[119] vdd gnd cell_6t
Xbit_r120_c107 bl[107] br[107] wl[120] vdd gnd cell_6t
Xbit_r121_c107 bl[107] br[107] wl[121] vdd gnd cell_6t
Xbit_r122_c107 bl[107] br[107] wl[122] vdd gnd cell_6t
Xbit_r123_c107 bl[107] br[107] wl[123] vdd gnd cell_6t
Xbit_r124_c107 bl[107] br[107] wl[124] vdd gnd cell_6t
Xbit_r125_c107 bl[107] br[107] wl[125] vdd gnd cell_6t
Xbit_r126_c107 bl[107] br[107] wl[126] vdd gnd cell_6t
Xbit_r127_c107 bl[107] br[107] wl[127] vdd gnd cell_6t
Xbit_r128_c107 bl[107] br[107] wl[128] vdd gnd cell_6t
Xbit_r129_c107 bl[107] br[107] wl[129] vdd gnd cell_6t
Xbit_r130_c107 bl[107] br[107] wl[130] vdd gnd cell_6t
Xbit_r131_c107 bl[107] br[107] wl[131] vdd gnd cell_6t
Xbit_r132_c107 bl[107] br[107] wl[132] vdd gnd cell_6t
Xbit_r133_c107 bl[107] br[107] wl[133] vdd gnd cell_6t
Xbit_r134_c107 bl[107] br[107] wl[134] vdd gnd cell_6t
Xbit_r135_c107 bl[107] br[107] wl[135] vdd gnd cell_6t
Xbit_r136_c107 bl[107] br[107] wl[136] vdd gnd cell_6t
Xbit_r137_c107 bl[107] br[107] wl[137] vdd gnd cell_6t
Xbit_r138_c107 bl[107] br[107] wl[138] vdd gnd cell_6t
Xbit_r139_c107 bl[107] br[107] wl[139] vdd gnd cell_6t
Xbit_r140_c107 bl[107] br[107] wl[140] vdd gnd cell_6t
Xbit_r141_c107 bl[107] br[107] wl[141] vdd gnd cell_6t
Xbit_r142_c107 bl[107] br[107] wl[142] vdd gnd cell_6t
Xbit_r143_c107 bl[107] br[107] wl[143] vdd gnd cell_6t
Xbit_r144_c107 bl[107] br[107] wl[144] vdd gnd cell_6t
Xbit_r145_c107 bl[107] br[107] wl[145] vdd gnd cell_6t
Xbit_r146_c107 bl[107] br[107] wl[146] vdd gnd cell_6t
Xbit_r147_c107 bl[107] br[107] wl[147] vdd gnd cell_6t
Xbit_r148_c107 bl[107] br[107] wl[148] vdd gnd cell_6t
Xbit_r149_c107 bl[107] br[107] wl[149] vdd gnd cell_6t
Xbit_r150_c107 bl[107] br[107] wl[150] vdd gnd cell_6t
Xbit_r151_c107 bl[107] br[107] wl[151] vdd gnd cell_6t
Xbit_r152_c107 bl[107] br[107] wl[152] vdd gnd cell_6t
Xbit_r153_c107 bl[107] br[107] wl[153] vdd gnd cell_6t
Xbit_r154_c107 bl[107] br[107] wl[154] vdd gnd cell_6t
Xbit_r155_c107 bl[107] br[107] wl[155] vdd gnd cell_6t
Xbit_r156_c107 bl[107] br[107] wl[156] vdd gnd cell_6t
Xbit_r157_c107 bl[107] br[107] wl[157] vdd gnd cell_6t
Xbit_r158_c107 bl[107] br[107] wl[158] vdd gnd cell_6t
Xbit_r159_c107 bl[107] br[107] wl[159] vdd gnd cell_6t
Xbit_r160_c107 bl[107] br[107] wl[160] vdd gnd cell_6t
Xbit_r161_c107 bl[107] br[107] wl[161] vdd gnd cell_6t
Xbit_r162_c107 bl[107] br[107] wl[162] vdd gnd cell_6t
Xbit_r163_c107 bl[107] br[107] wl[163] vdd gnd cell_6t
Xbit_r164_c107 bl[107] br[107] wl[164] vdd gnd cell_6t
Xbit_r165_c107 bl[107] br[107] wl[165] vdd gnd cell_6t
Xbit_r166_c107 bl[107] br[107] wl[166] vdd gnd cell_6t
Xbit_r167_c107 bl[107] br[107] wl[167] vdd gnd cell_6t
Xbit_r168_c107 bl[107] br[107] wl[168] vdd gnd cell_6t
Xbit_r169_c107 bl[107] br[107] wl[169] vdd gnd cell_6t
Xbit_r170_c107 bl[107] br[107] wl[170] vdd gnd cell_6t
Xbit_r171_c107 bl[107] br[107] wl[171] vdd gnd cell_6t
Xbit_r172_c107 bl[107] br[107] wl[172] vdd gnd cell_6t
Xbit_r173_c107 bl[107] br[107] wl[173] vdd gnd cell_6t
Xbit_r174_c107 bl[107] br[107] wl[174] vdd gnd cell_6t
Xbit_r175_c107 bl[107] br[107] wl[175] vdd gnd cell_6t
Xbit_r176_c107 bl[107] br[107] wl[176] vdd gnd cell_6t
Xbit_r177_c107 bl[107] br[107] wl[177] vdd gnd cell_6t
Xbit_r178_c107 bl[107] br[107] wl[178] vdd gnd cell_6t
Xbit_r179_c107 bl[107] br[107] wl[179] vdd gnd cell_6t
Xbit_r180_c107 bl[107] br[107] wl[180] vdd gnd cell_6t
Xbit_r181_c107 bl[107] br[107] wl[181] vdd gnd cell_6t
Xbit_r182_c107 bl[107] br[107] wl[182] vdd gnd cell_6t
Xbit_r183_c107 bl[107] br[107] wl[183] vdd gnd cell_6t
Xbit_r184_c107 bl[107] br[107] wl[184] vdd gnd cell_6t
Xbit_r185_c107 bl[107] br[107] wl[185] vdd gnd cell_6t
Xbit_r186_c107 bl[107] br[107] wl[186] vdd gnd cell_6t
Xbit_r187_c107 bl[107] br[107] wl[187] vdd gnd cell_6t
Xbit_r188_c107 bl[107] br[107] wl[188] vdd gnd cell_6t
Xbit_r189_c107 bl[107] br[107] wl[189] vdd gnd cell_6t
Xbit_r190_c107 bl[107] br[107] wl[190] vdd gnd cell_6t
Xbit_r191_c107 bl[107] br[107] wl[191] vdd gnd cell_6t
Xbit_r192_c107 bl[107] br[107] wl[192] vdd gnd cell_6t
Xbit_r193_c107 bl[107] br[107] wl[193] vdd gnd cell_6t
Xbit_r194_c107 bl[107] br[107] wl[194] vdd gnd cell_6t
Xbit_r195_c107 bl[107] br[107] wl[195] vdd gnd cell_6t
Xbit_r196_c107 bl[107] br[107] wl[196] vdd gnd cell_6t
Xbit_r197_c107 bl[107] br[107] wl[197] vdd gnd cell_6t
Xbit_r198_c107 bl[107] br[107] wl[198] vdd gnd cell_6t
Xbit_r199_c107 bl[107] br[107] wl[199] vdd gnd cell_6t
Xbit_r200_c107 bl[107] br[107] wl[200] vdd gnd cell_6t
Xbit_r201_c107 bl[107] br[107] wl[201] vdd gnd cell_6t
Xbit_r202_c107 bl[107] br[107] wl[202] vdd gnd cell_6t
Xbit_r203_c107 bl[107] br[107] wl[203] vdd gnd cell_6t
Xbit_r204_c107 bl[107] br[107] wl[204] vdd gnd cell_6t
Xbit_r205_c107 bl[107] br[107] wl[205] vdd gnd cell_6t
Xbit_r206_c107 bl[107] br[107] wl[206] vdd gnd cell_6t
Xbit_r207_c107 bl[107] br[107] wl[207] vdd gnd cell_6t
Xbit_r208_c107 bl[107] br[107] wl[208] vdd gnd cell_6t
Xbit_r209_c107 bl[107] br[107] wl[209] vdd gnd cell_6t
Xbit_r210_c107 bl[107] br[107] wl[210] vdd gnd cell_6t
Xbit_r211_c107 bl[107] br[107] wl[211] vdd gnd cell_6t
Xbit_r212_c107 bl[107] br[107] wl[212] vdd gnd cell_6t
Xbit_r213_c107 bl[107] br[107] wl[213] vdd gnd cell_6t
Xbit_r214_c107 bl[107] br[107] wl[214] vdd gnd cell_6t
Xbit_r215_c107 bl[107] br[107] wl[215] vdd gnd cell_6t
Xbit_r216_c107 bl[107] br[107] wl[216] vdd gnd cell_6t
Xbit_r217_c107 bl[107] br[107] wl[217] vdd gnd cell_6t
Xbit_r218_c107 bl[107] br[107] wl[218] vdd gnd cell_6t
Xbit_r219_c107 bl[107] br[107] wl[219] vdd gnd cell_6t
Xbit_r220_c107 bl[107] br[107] wl[220] vdd gnd cell_6t
Xbit_r221_c107 bl[107] br[107] wl[221] vdd gnd cell_6t
Xbit_r222_c107 bl[107] br[107] wl[222] vdd gnd cell_6t
Xbit_r223_c107 bl[107] br[107] wl[223] vdd gnd cell_6t
Xbit_r224_c107 bl[107] br[107] wl[224] vdd gnd cell_6t
Xbit_r225_c107 bl[107] br[107] wl[225] vdd gnd cell_6t
Xbit_r226_c107 bl[107] br[107] wl[226] vdd gnd cell_6t
Xbit_r227_c107 bl[107] br[107] wl[227] vdd gnd cell_6t
Xbit_r228_c107 bl[107] br[107] wl[228] vdd gnd cell_6t
Xbit_r229_c107 bl[107] br[107] wl[229] vdd gnd cell_6t
Xbit_r230_c107 bl[107] br[107] wl[230] vdd gnd cell_6t
Xbit_r231_c107 bl[107] br[107] wl[231] vdd gnd cell_6t
Xbit_r232_c107 bl[107] br[107] wl[232] vdd gnd cell_6t
Xbit_r233_c107 bl[107] br[107] wl[233] vdd gnd cell_6t
Xbit_r234_c107 bl[107] br[107] wl[234] vdd gnd cell_6t
Xbit_r235_c107 bl[107] br[107] wl[235] vdd gnd cell_6t
Xbit_r236_c107 bl[107] br[107] wl[236] vdd gnd cell_6t
Xbit_r237_c107 bl[107] br[107] wl[237] vdd gnd cell_6t
Xbit_r238_c107 bl[107] br[107] wl[238] vdd gnd cell_6t
Xbit_r239_c107 bl[107] br[107] wl[239] vdd gnd cell_6t
Xbit_r240_c107 bl[107] br[107] wl[240] vdd gnd cell_6t
Xbit_r241_c107 bl[107] br[107] wl[241] vdd gnd cell_6t
Xbit_r242_c107 bl[107] br[107] wl[242] vdd gnd cell_6t
Xbit_r243_c107 bl[107] br[107] wl[243] vdd gnd cell_6t
Xbit_r244_c107 bl[107] br[107] wl[244] vdd gnd cell_6t
Xbit_r245_c107 bl[107] br[107] wl[245] vdd gnd cell_6t
Xbit_r246_c107 bl[107] br[107] wl[246] vdd gnd cell_6t
Xbit_r247_c107 bl[107] br[107] wl[247] vdd gnd cell_6t
Xbit_r248_c107 bl[107] br[107] wl[248] vdd gnd cell_6t
Xbit_r249_c107 bl[107] br[107] wl[249] vdd gnd cell_6t
Xbit_r250_c107 bl[107] br[107] wl[250] vdd gnd cell_6t
Xbit_r251_c107 bl[107] br[107] wl[251] vdd gnd cell_6t
Xbit_r252_c107 bl[107] br[107] wl[252] vdd gnd cell_6t
Xbit_r253_c107 bl[107] br[107] wl[253] vdd gnd cell_6t
Xbit_r254_c107 bl[107] br[107] wl[254] vdd gnd cell_6t
Xbit_r255_c107 bl[107] br[107] wl[255] vdd gnd cell_6t
Xbit_r0_c108 bl[108] br[108] wl[0] vdd gnd cell_6t
Xbit_r1_c108 bl[108] br[108] wl[1] vdd gnd cell_6t
Xbit_r2_c108 bl[108] br[108] wl[2] vdd gnd cell_6t
Xbit_r3_c108 bl[108] br[108] wl[3] vdd gnd cell_6t
Xbit_r4_c108 bl[108] br[108] wl[4] vdd gnd cell_6t
Xbit_r5_c108 bl[108] br[108] wl[5] vdd gnd cell_6t
Xbit_r6_c108 bl[108] br[108] wl[6] vdd gnd cell_6t
Xbit_r7_c108 bl[108] br[108] wl[7] vdd gnd cell_6t
Xbit_r8_c108 bl[108] br[108] wl[8] vdd gnd cell_6t
Xbit_r9_c108 bl[108] br[108] wl[9] vdd gnd cell_6t
Xbit_r10_c108 bl[108] br[108] wl[10] vdd gnd cell_6t
Xbit_r11_c108 bl[108] br[108] wl[11] vdd gnd cell_6t
Xbit_r12_c108 bl[108] br[108] wl[12] vdd gnd cell_6t
Xbit_r13_c108 bl[108] br[108] wl[13] vdd gnd cell_6t
Xbit_r14_c108 bl[108] br[108] wl[14] vdd gnd cell_6t
Xbit_r15_c108 bl[108] br[108] wl[15] vdd gnd cell_6t
Xbit_r16_c108 bl[108] br[108] wl[16] vdd gnd cell_6t
Xbit_r17_c108 bl[108] br[108] wl[17] vdd gnd cell_6t
Xbit_r18_c108 bl[108] br[108] wl[18] vdd gnd cell_6t
Xbit_r19_c108 bl[108] br[108] wl[19] vdd gnd cell_6t
Xbit_r20_c108 bl[108] br[108] wl[20] vdd gnd cell_6t
Xbit_r21_c108 bl[108] br[108] wl[21] vdd gnd cell_6t
Xbit_r22_c108 bl[108] br[108] wl[22] vdd gnd cell_6t
Xbit_r23_c108 bl[108] br[108] wl[23] vdd gnd cell_6t
Xbit_r24_c108 bl[108] br[108] wl[24] vdd gnd cell_6t
Xbit_r25_c108 bl[108] br[108] wl[25] vdd gnd cell_6t
Xbit_r26_c108 bl[108] br[108] wl[26] vdd gnd cell_6t
Xbit_r27_c108 bl[108] br[108] wl[27] vdd gnd cell_6t
Xbit_r28_c108 bl[108] br[108] wl[28] vdd gnd cell_6t
Xbit_r29_c108 bl[108] br[108] wl[29] vdd gnd cell_6t
Xbit_r30_c108 bl[108] br[108] wl[30] vdd gnd cell_6t
Xbit_r31_c108 bl[108] br[108] wl[31] vdd gnd cell_6t
Xbit_r32_c108 bl[108] br[108] wl[32] vdd gnd cell_6t
Xbit_r33_c108 bl[108] br[108] wl[33] vdd gnd cell_6t
Xbit_r34_c108 bl[108] br[108] wl[34] vdd gnd cell_6t
Xbit_r35_c108 bl[108] br[108] wl[35] vdd gnd cell_6t
Xbit_r36_c108 bl[108] br[108] wl[36] vdd gnd cell_6t
Xbit_r37_c108 bl[108] br[108] wl[37] vdd gnd cell_6t
Xbit_r38_c108 bl[108] br[108] wl[38] vdd gnd cell_6t
Xbit_r39_c108 bl[108] br[108] wl[39] vdd gnd cell_6t
Xbit_r40_c108 bl[108] br[108] wl[40] vdd gnd cell_6t
Xbit_r41_c108 bl[108] br[108] wl[41] vdd gnd cell_6t
Xbit_r42_c108 bl[108] br[108] wl[42] vdd gnd cell_6t
Xbit_r43_c108 bl[108] br[108] wl[43] vdd gnd cell_6t
Xbit_r44_c108 bl[108] br[108] wl[44] vdd gnd cell_6t
Xbit_r45_c108 bl[108] br[108] wl[45] vdd gnd cell_6t
Xbit_r46_c108 bl[108] br[108] wl[46] vdd gnd cell_6t
Xbit_r47_c108 bl[108] br[108] wl[47] vdd gnd cell_6t
Xbit_r48_c108 bl[108] br[108] wl[48] vdd gnd cell_6t
Xbit_r49_c108 bl[108] br[108] wl[49] vdd gnd cell_6t
Xbit_r50_c108 bl[108] br[108] wl[50] vdd gnd cell_6t
Xbit_r51_c108 bl[108] br[108] wl[51] vdd gnd cell_6t
Xbit_r52_c108 bl[108] br[108] wl[52] vdd gnd cell_6t
Xbit_r53_c108 bl[108] br[108] wl[53] vdd gnd cell_6t
Xbit_r54_c108 bl[108] br[108] wl[54] vdd gnd cell_6t
Xbit_r55_c108 bl[108] br[108] wl[55] vdd gnd cell_6t
Xbit_r56_c108 bl[108] br[108] wl[56] vdd gnd cell_6t
Xbit_r57_c108 bl[108] br[108] wl[57] vdd gnd cell_6t
Xbit_r58_c108 bl[108] br[108] wl[58] vdd gnd cell_6t
Xbit_r59_c108 bl[108] br[108] wl[59] vdd gnd cell_6t
Xbit_r60_c108 bl[108] br[108] wl[60] vdd gnd cell_6t
Xbit_r61_c108 bl[108] br[108] wl[61] vdd gnd cell_6t
Xbit_r62_c108 bl[108] br[108] wl[62] vdd gnd cell_6t
Xbit_r63_c108 bl[108] br[108] wl[63] vdd gnd cell_6t
Xbit_r64_c108 bl[108] br[108] wl[64] vdd gnd cell_6t
Xbit_r65_c108 bl[108] br[108] wl[65] vdd gnd cell_6t
Xbit_r66_c108 bl[108] br[108] wl[66] vdd gnd cell_6t
Xbit_r67_c108 bl[108] br[108] wl[67] vdd gnd cell_6t
Xbit_r68_c108 bl[108] br[108] wl[68] vdd gnd cell_6t
Xbit_r69_c108 bl[108] br[108] wl[69] vdd gnd cell_6t
Xbit_r70_c108 bl[108] br[108] wl[70] vdd gnd cell_6t
Xbit_r71_c108 bl[108] br[108] wl[71] vdd gnd cell_6t
Xbit_r72_c108 bl[108] br[108] wl[72] vdd gnd cell_6t
Xbit_r73_c108 bl[108] br[108] wl[73] vdd gnd cell_6t
Xbit_r74_c108 bl[108] br[108] wl[74] vdd gnd cell_6t
Xbit_r75_c108 bl[108] br[108] wl[75] vdd gnd cell_6t
Xbit_r76_c108 bl[108] br[108] wl[76] vdd gnd cell_6t
Xbit_r77_c108 bl[108] br[108] wl[77] vdd gnd cell_6t
Xbit_r78_c108 bl[108] br[108] wl[78] vdd gnd cell_6t
Xbit_r79_c108 bl[108] br[108] wl[79] vdd gnd cell_6t
Xbit_r80_c108 bl[108] br[108] wl[80] vdd gnd cell_6t
Xbit_r81_c108 bl[108] br[108] wl[81] vdd gnd cell_6t
Xbit_r82_c108 bl[108] br[108] wl[82] vdd gnd cell_6t
Xbit_r83_c108 bl[108] br[108] wl[83] vdd gnd cell_6t
Xbit_r84_c108 bl[108] br[108] wl[84] vdd gnd cell_6t
Xbit_r85_c108 bl[108] br[108] wl[85] vdd gnd cell_6t
Xbit_r86_c108 bl[108] br[108] wl[86] vdd gnd cell_6t
Xbit_r87_c108 bl[108] br[108] wl[87] vdd gnd cell_6t
Xbit_r88_c108 bl[108] br[108] wl[88] vdd gnd cell_6t
Xbit_r89_c108 bl[108] br[108] wl[89] vdd gnd cell_6t
Xbit_r90_c108 bl[108] br[108] wl[90] vdd gnd cell_6t
Xbit_r91_c108 bl[108] br[108] wl[91] vdd gnd cell_6t
Xbit_r92_c108 bl[108] br[108] wl[92] vdd gnd cell_6t
Xbit_r93_c108 bl[108] br[108] wl[93] vdd gnd cell_6t
Xbit_r94_c108 bl[108] br[108] wl[94] vdd gnd cell_6t
Xbit_r95_c108 bl[108] br[108] wl[95] vdd gnd cell_6t
Xbit_r96_c108 bl[108] br[108] wl[96] vdd gnd cell_6t
Xbit_r97_c108 bl[108] br[108] wl[97] vdd gnd cell_6t
Xbit_r98_c108 bl[108] br[108] wl[98] vdd gnd cell_6t
Xbit_r99_c108 bl[108] br[108] wl[99] vdd gnd cell_6t
Xbit_r100_c108 bl[108] br[108] wl[100] vdd gnd cell_6t
Xbit_r101_c108 bl[108] br[108] wl[101] vdd gnd cell_6t
Xbit_r102_c108 bl[108] br[108] wl[102] vdd gnd cell_6t
Xbit_r103_c108 bl[108] br[108] wl[103] vdd gnd cell_6t
Xbit_r104_c108 bl[108] br[108] wl[104] vdd gnd cell_6t
Xbit_r105_c108 bl[108] br[108] wl[105] vdd gnd cell_6t
Xbit_r106_c108 bl[108] br[108] wl[106] vdd gnd cell_6t
Xbit_r107_c108 bl[108] br[108] wl[107] vdd gnd cell_6t
Xbit_r108_c108 bl[108] br[108] wl[108] vdd gnd cell_6t
Xbit_r109_c108 bl[108] br[108] wl[109] vdd gnd cell_6t
Xbit_r110_c108 bl[108] br[108] wl[110] vdd gnd cell_6t
Xbit_r111_c108 bl[108] br[108] wl[111] vdd gnd cell_6t
Xbit_r112_c108 bl[108] br[108] wl[112] vdd gnd cell_6t
Xbit_r113_c108 bl[108] br[108] wl[113] vdd gnd cell_6t
Xbit_r114_c108 bl[108] br[108] wl[114] vdd gnd cell_6t
Xbit_r115_c108 bl[108] br[108] wl[115] vdd gnd cell_6t
Xbit_r116_c108 bl[108] br[108] wl[116] vdd gnd cell_6t
Xbit_r117_c108 bl[108] br[108] wl[117] vdd gnd cell_6t
Xbit_r118_c108 bl[108] br[108] wl[118] vdd gnd cell_6t
Xbit_r119_c108 bl[108] br[108] wl[119] vdd gnd cell_6t
Xbit_r120_c108 bl[108] br[108] wl[120] vdd gnd cell_6t
Xbit_r121_c108 bl[108] br[108] wl[121] vdd gnd cell_6t
Xbit_r122_c108 bl[108] br[108] wl[122] vdd gnd cell_6t
Xbit_r123_c108 bl[108] br[108] wl[123] vdd gnd cell_6t
Xbit_r124_c108 bl[108] br[108] wl[124] vdd gnd cell_6t
Xbit_r125_c108 bl[108] br[108] wl[125] vdd gnd cell_6t
Xbit_r126_c108 bl[108] br[108] wl[126] vdd gnd cell_6t
Xbit_r127_c108 bl[108] br[108] wl[127] vdd gnd cell_6t
Xbit_r128_c108 bl[108] br[108] wl[128] vdd gnd cell_6t
Xbit_r129_c108 bl[108] br[108] wl[129] vdd gnd cell_6t
Xbit_r130_c108 bl[108] br[108] wl[130] vdd gnd cell_6t
Xbit_r131_c108 bl[108] br[108] wl[131] vdd gnd cell_6t
Xbit_r132_c108 bl[108] br[108] wl[132] vdd gnd cell_6t
Xbit_r133_c108 bl[108] br[108] wl[133] vdd gnd cell_6t
Xbit_r134_c108 bl[108] br[108] wl[134] vdd gnd cell_6t
Xbit_r135_c108 bl[108] br[108] wl[135] vdd gnd cell_6t
Xbit_r136_c108 bl[108] br[108] wl[136] vdd gnd cell_6t
Xbit_r137_c108 bl[108] br[108] wl[137] vdd gnd cell_6t
Xbit_r138_c108 bl[108] br[108] wl[138] vdd gnd cell_6t
Xbit_r139_c108 bl[108] br[108] wl[139] vdd gnd cell_6t
Xbit_r140_c108 bl[108] br[108] wl[140] vdd gnd cell_6t
Xbit_r141_c108 bl[108] br[108] wl[141] vdd gnd cell_6t
Xbit_r142_c108 bl[108] br[108] wl[142] vdd gnd cell_6t
Xbit_r143_c108 bl[108] br[108] wl[143] vdd gnd cell_6t
Xbit_r144_c108 bl[108] br[108] wl[144] vdd gnd cell_6t
Xbit_r145_c108 bl[108] br[108] wl[145] vdd gnd cell_6t
Xbit_r146_c108 bl[108] br[108] wl[146] vdd gnd cell_6t
Xbit_r147_c108 bl[108] br[108] wl[147] vdd gnd cell_6t
Xbit_r148_c108 bl[108] br[108] wl[148] vdd gnd cell_6t
Xbit_r149_c108 bl[108] br[108] wl[149] vdd gnd cell_6t
Xbit_r150_c108 bl[108] br[108] wl[150] vdd gnd cell_6t
Xbit_r151_c108 bl[108] br[108] wl[151] vdd gnd cell_6t
Xbit_r152_c108 bl[108] br[108] wl[152] vdd gnd cell_6t
Xbit_r153_c108 bl[108] br[108] wl[153] vdd gnd cell_6t
Xbit_r154_c108 bl[108] br[108] wl[154] vdd gnd cell_6t
Xbit_r155_c108 bl[108] br[108] wl[155] vdd gnd cell_6t
Xbit_r156_c108 bl[108] br[108] wl[156] vdd gnd cell_6t
Xbit_r157_c108 bl[108] br[108] wl[157] vdd gnd cell_6t
Xbit_r158_c108 bl[108] br[108] wl[158] vdd gnd cell_6t
Xbit_r159_c108 bl[108] br[108] wl[159] vdd gnd cell_6t
Xbit_r160_c108 bl[108] br[108] wl[160] vdd gnd cell_6t
Xbit_r161_c108 bl[108] br[108] wl[161] vdd gnd cell_6t
Xbit_r162_c108 bl[108] br[108] wl[162] vdd gnd cell_6t
Xbit_r163_c108 bl[108] br[108] wl[163] vdd gnd cell_6t
Xbit_r164_c108 bl[108] br[108] wl[164] vdd gnd cell_6t
Xbit_r165_c108 bl[108] br[108] wl[165] vdd gnd cell_6t
Xbit_r166_c108 bl[108] br[108] wl[166] vdd gnd cell_6t
Xbit_r167_c108 bl[108] br[108] wl[167] vdd gnd cell_6t
Xbit_r168_c108 bl[108] br[108] wl[168] vdd gnd cell_6t
Xbit_r169_c108 bl[108] br[108] wl[169] vdd gnd cell_6t
Xbit_r170_c108 bl[108] br[108] wl[170] vdd gnd cell_6t
Xbit_r171_c108 bl[108] br[108] wl[171] vdd gnd cell_6t
Xbit_r172_c108 bl[108] br[108] wl[172] vdd gnd cell_6t
Xbit_r173_c108 bl[108] br[108] wl[173] vdd gnd cell_6t
Xbit_r174_c108 bl[108] br[108] wl[174] vdd gnd cell_6t
Xbit_r175_c108 bl[108] br[108] wl[175] vdd gnd cell_6t
Xbit_r176_c108 bl[108] br[108] wl[176] vdd gnd cell_6t
Xbit_r177_c108 bl[108] br[108] wl[177] vdd gnd cell_6t
Xbit_r178_c108 bl[108] br[108] wl[178] vdd gnd cell_6t
Xbit_r179_c108 bl[108] br[108] wl[179] vdd gnd cell_6t
Xbit_r180_c108 bl[108] br[108] wl[180] vdd gnd cell_6t
Xbit_r181_c108 bl[108] br[108] wl[181] vdd gnd cell_6t
Xbit_r182_c108 bl[108] br[108] wl[182] vdd gnd cell_6t
Xbit_r183_c108 bl[108] br[108] wl[183] vdd gnd cell_6t
Xbit_r184_c108 bl[108] br[108] wl[184] vdd gnd cell_6t
Xbit_r185_c108 bl[108] br[108] wl[185] vdd gnd cell_6t
Xbit_r186_c108 bl[108] br[108] wl[186] vdd gnd cell_6t
Xbit_r187_c108 bl[108] br[108] wl[187] vdd gnd cell_6t
Xbit_r188_c108 bl[108] br[108] wl[188] vdd gnd cell_6t
Xbit_r189_c108 bl[108] br[108] wl[189] vdd gnd cell_6t
Xbit_r190_c108 bl[108] br[108] wl[190] vdd gnd cell_6t
Xbit_r191_c108 bl[108] br[108] wl[191] vdd gnd cell_6t
Xbit_r192_c108 bl[108] br[108] wl[192] vdd gnd cell_6t
Xbit_r193_c108 bl[108] br[108] wl[193] vdd gnd cell_6t
Xbit_r194_c108 bl[108] br[108] wl[194] vdd gnd cell_6t
Xbit_r195_c108 bl[108] br[108] wl[195] vdd gnd cell_6t
Xbit_r196_c108 bl[108] br[108] wl[196] vdd gnd cell_6t
Xbit_r197_c108 bl[108] br[108] wl[197] vdd gnd cell_6t
Xbit_r198_c108 bl[108] br[108] wl[198] vdd gnd cell_6t
Xbit_r199_c108 bl[108] br[108] wl[199] vdd gnd cell_6t
Xbit_r200_c108 bl[108] br[108] wl[200] vdd gnd cell_6t
Xbit_r201_c108 bl[108] br[108] wl[201] vdd gnd cell_6t
Xbit_r202_c108 bl[108] br[108] wl[202] vdd gnd cell_6t
Xbit_r203_c108 bl[108] br[108] wl[203] vdd gnd cell_6t
Xbit_r204_c108 bl[108] br[108] wl[204] vdd gnd cell_6t
Xbit_r205_c108 bl[108] br[108] wl[205] vdd gnd cell_6t
Xbit_r206_c108 bl[108] br[108] wl[206] vdd gnd cell_6t
Xbit_r207_c108 bl[108] br[108] wl[207] vdd gnd cell_6t
Xbit_r208_c108 bl[108] br[108] wl[208] vdd gnd cell_6t
Xbit_r209_c108 bl[108] br[108] wl[209] vdd gnd cell_6t
Xbit_r210_c108 bl[108] br[108] wl[210] vdd gnd cell_6t
Xbit_r211_c108 bl[108] br[108] wl[211] vdd gnd cell_6t
Xbit_r212_c108 bl[108] br[108] wl[212] vdd gnd cell_6t
Xbit_r213_c108 bl[108] br[108] wl[213] vdd gnd cell_6t
Xbit_r214_c108 bl[108] br[108] wl[214] vdd gnd cell_6t
Xbit_r215_c108 bl[108] br[108] wl[215] vdd gnd cell_6t
Xbit_r216_c108 bl[108] br[108] wl[216] vdd gnd cell_6t
Xbit_r217_c108 bl[108] br[108] wl[217] vdd gnd cell_6t
Xbit_r218_c108 bl[108] br[108] wl[218] vdd gnd cell_6t
Xbit_r219_c108 bl[108] br[108] wl[219] vdd gnd cell_6t
Xbit_r220_c108 bl[108] br[108] wl[220] vdd gnd cell_6t
Xbit_r221_c108 bl[108] br[108] wl[221] vdd gnd cell_6t
Xbit_r222_c108 bl[108] br[108] wl[222] vdd gnd cell_6t
Xbit_r223_c108 bl[108] br[108] wl[223] vdd gnd cell_6t
Xbit_r224_c108 bl[108] br[108] wl[224] vdd gnd cell_6t
Xbit_r225_c108 bl[108] br[108] wl[225] vdd gnd cell_6t
Xbit_r226_c108 bl[108] br[108] wl[226] vdd gnd cell_6t
Xbit_r227_c108 bl[108] br[108] wl[227] vdd gnd cell_6t
Xbit_r228_c108 bl[108] br[108] wl[228] vdd gnd cell_6t
Xbit_r229_c108 bl[108] br[108] wl[229] vdd gnd cell_6t
Xbit_r230_c108 bl[108] br[108] wl[230] vdd gnd cell_6t
Xbit_r231_c108 bl[108] br[108] wl[231] vdd gnd cell_6t
Xbit_r232_c108 bl[108] br[108] wl[232] vdd gnd cell_6t
Xbit_r233_c108 bl[108] br[108] wl[233] vdd gnd cell_6t
Xbit_r234_c108 bl[108] br[108] wl[234] vdd gnd cell_6t
Xbit_r235_c108 bl[108] br[108] wl[235] vdd gnd cell_6t
Xbit_r236_c108 bl[108] br[108] wl[236] vdd gnd cell_6t
Xbit_r237_c108 bl[108] br[108] wl[237] vdd gnd cell_6t
Xbit_r238_c108 bl[108] br[108] wl[238] vdd gnd cell_6t
Xbit_r239_c108 bl[108] br[108] wl[239] vdd gnd cell_6t
Xbit_r240_c108 bl[108] br[108] wl[240] vdd gnd cell_6t
Xbit_r241_c108 bl[108] br[108] wl[241] vdd gnd cell_6t
Xbit_r242_c108 bl[108] br[108] wl[242] vdd gnd cell_6t
Xbit_r243_c108 bl[108] br[108] wl[243] vdd gnd cell_6t
Xbit_r244_c108 bl[108] br[108] wl[244] vdd gnd cell_6t
Xbit_r245_c108 bl[108] br[108] wl[245] vdd gnd cell_6t
Xbit_r246_c108 bl[108] br[108] wl[246] vdd gnd cell_6t
Xbit_r247_c108 bl[108] br[108] wl[247] vdd gnd cell_6t
Xbit_r248_c108 bl[108] br[108] wl[248] vdd gnd cell_6t
Xbit_r249_c108 bl[108] br[108] wl[249] vdd gnd cell_6t
Xbit_r250_c108 bl[108] br[108] wl[250] vdd gnd cell_6t
Xbit_r251_c108 bl[108] br[108] wl[251] vdd gnd cell_6t
Xbit_r252_c108 bl[108] br[108] wl[252] vdd gnd cell_6t
Xbit_r253_c108 bl[108] br[108] wl[253] vdd gnd cell_6t
Xbit_r254_c108 bl[108] br[108] wl[254] vdd gnd cell_6t
Xbit_r255_c108 bl[108] br[108] wl[255] vdd gnd cell_6t
Xbit_r0_c109 bl[109] br[109] wl[0] vdd gnd cell_6t
Xbit_r1_c109 bl[109] br[109] wl[1] vdd gnd cell_6t
Xbit_r2_c109 bl[109] br[109] wl[2] vdd gnd cell_6t
Xbit_r3_c109 bl[109] br[109] wl[3] vdd gnd cell_6t
Xbit_r4_c109 bl[109] br[109] wl[4] vdd gnd cell_6t
Xbit_r5_c109 bl[109] br[109] wl[5] vdd gnd cell_6t
Xbit_r6_c109 bl[109] br[109] wl[6] vdd gnd cell_6t
Xbit_r7_c109 bl[109] br[109] wl[7] vdd gnd cell_6t
Xbit_r8_c109 bl[109] br[109] wl[8] vdd gnd cell_6t
Xbit_r9_c109 bl[109] br[109] wl[9] vdd gnd cell_6t
Xbit_r10_c109 bl[109] br[109] wl[10] vdd gnd cell_6t
Xbit_r11_c109 bl[109] br[109] wl[11] vdd gnd cell_6t
Xbit_r12_c109 bl[109] br[109] wl[12] vdd gnd cell_6t
Xbit_r13_c109 bl[109] br[109] wl[13] vdd gnd cell_6t
Xbit_r14_c109 bl[109] br[109] wl[14] vdd gnd cell_6t
Xbit_r15_c109 bl[109] br[109] wl[15] vdd gnd cell_6t
Xbit_r16_c109 bl[109] br[109] wl[16] vdd gnd cell_6t
Xbit_r17_c109 bl[109] br[109] wl[17] vdd gnd cell_6t
Xbit_r18_c109 bl[109] br[109] wl[18] vdd gnd cell_6t
Xbit_r19_c109 bl[109] br[109] wl[19] vdd gnd cell_6t
Xbit_r20_c109 bl[109] br[109] wl[20] vdd gnd cell_6t
Xbit_r21_c109 bl[109] br[109] wl[21] vdd gnd cell_6t
Xbit_r22_c109 bl[109] br[109] wl[22] vdd gnd cell_6t
Xbit_r23_c109 bl[109] br[109] wl[23] vdd gnd cell_6t
Xbit_r24_c109 bl[109] br[109] wl[24] vdd gnd cell_6t
Xbit_r25_c109 bl[109] br[109] wl[25] vdd gnd cell_6t
Xbit_r26_c109 bl[109] br[109] wl[26] vdd gnd cell_6t
Xbit_r27_c109 bl[109] br[109] wl[27] vdd gnd cell_6t
Xbit_r28_c109 bl[109] br[109] wl[28] vdd gnd cell_6t
Xbit_r29_c109 bl[109] br[109] wl[29] vdd gnd cell_6t
Xbit_r30_c109 bl[109] br[109] wl[30] vdd gnd cell_6t
Xbit_r31_c109 bl[109] br[109] wl[31] vdd gnd cell_6t
Xbit_r32_c109 bl[109] br[109] wl[32] vdd gnd cell_6t
Xbit_r33_c109 bl[109] br[109] wl[33] vdd gnd cell_6t
Xbit_r34_c109 bl[109] br[109] wl[34] vdd gnd cell_6t
Xbit_r35_c109 bl[109] br[109] wl[35] vdd gnd cell_6t
Xbit_r36_c109 bl[109] br[109] wl[36] vdd gnd cell_6t
Xbit_r37_c109 bl[109] br[109] wl[37] vdd gnd cell_6t
Xbit_r38_c109 bl[109] br[109] wl[38] vdd gnd cell_6t
Xbit_r39_c109 bl[109] br[109] wl[39] vdd gnd cell_6t
Xbit_r40_c109 bl[109] br[109] wl[40] vdd gnd cell_6t
Xbit_r41_c109 bl[109] br[109] wl[41] vdd gnd cell_6t
Xbit_r42_c109 bl[109] br[109] wl[42] vdd gnd cell_6t
Xbit_r43_c109 bl[109] br[109] wl[43] vdd gnd cell_6t
Xbit_r44_c109 bl[109] br[109] wl[44] vdd gnd cell_6t
Xbit_r45_c109 bl[109] br[109] wl[45] vdd gnd cell_6t
Xbit_r46_c109 bl[109] br[109] wl[46] vdd gnd cell_6t
Xbit_r47_c109 bl[109] br[109] wl[47] vdd gnd cell_6t
Xbit_r48_c109 bl[109] br[109] wl[48] vdd gnd cell_6t
Xbit_r49_c109 bl[109] br[109] wl[49] vdd gnd cell_6t
Xbit_r50_c109 bl[109] br[109] wl[50] vdd gnd cell_6t
Xbit_r51_c109 bl[109] br[109] wl[51] vdd gnd cell_6t
Xbit_r52_c109 bl[109] br[109] wl[52] vdd gnd cell_6t
Xbit_r53_c109 bl[109] br[109] wl[53] vdd gnd cell_6t
Xbit_r54_c109 bl[109] br[109] wl[54] vdd gnd cell_6t
Xbit_r55_c109 bl[109] br[109] wl[55] vdd gnd cell_6t
Xbit_r56_c109 bl[109] br[109] wl[56] vdd gnd cell_6t
Xbit_r57_c109 bl[109] br[109] wl[57] vdd gnd cell_6t
Xbit_r58_c109 bl[109] br[109] wl[58] vdd gnd cell_6t
Xbit_r59_c109 bl[109] br[109] wl[59] vdd gnd cell_6t
Xbit_r60_c109 bl[109] br[109] wl[60] vdd gnd cell_6t
Xbit_r61_c109 bl[109] br[109] wl[61] vdd gnd cell_6t
Xbit_r62_c109 bl[109] br[109] wl[62] vdd gnd cell_6t
Xbit_r63_c109 bl[109] br[109] wl[63] vdd gnd cell_6t
Xbit_r64_c109 bl[109] br[109] wl[64] vdd gnd cell_6t
Xbit_r65_c109 bl[109] br[109] wl[65] vdd gnd cell_6t
Xbit_r66_c109 bl[109] br[109] wl[66] vdd gnd cell_6t
Xbit_r67_c109 bl[109] br[109] wl[67] vdd gnd cell_6t
Xbit_r68_c109 bl[109] br[109] wl[68] vdd gnd cell_6t
Xbit_r69_c109 bl[109] br[109] wl[69] vdd gnd cell_6t
Xbit_r70_c109 bl[109] br[109] wl[70] vdd gnd cell_6t
Xbit_r71_c109 bl[109] br[109] wl[71] vdd gnd cell_6t
Xbit_r72_c109 bl[109] br[109] wl[72] vdd gnd cell_6t
Xbit_r73_c109 bl[109] br[109] wl[73] vdd gnd cell_6t
Xbit_r74_c109 bl[109] br[109] wl[74] vdd gnd cell_6t
Xbit_r75_c109 bl[109] br[109] wl[75] vdd gnd cell_6t
Xbit_r76_c109 bl[109] br[109] wl[76] vdd gnd cell_6t
Xbit_r77_c109 bl[109] br[109] wl[77] vdd gnd cell_6t
Xbit_r78_c109 bl[109] br[109] wl[78] vdd gnd cell_6t
Xbit_r79_c109 bl[109] br[109] wl[79] vdd gnd cell_6t
Xbit_r80_c109 bl[109] br[109] wl[80] vdd gnd cell_6t
Xbit_r81_c109 bl[109] br[109] wl[81] vdd gnd cell_6t
Xbit_r82_c109 bl[109] br[109] wl[82] vdd gnd cell_6t
Xbit_r83_c109 bl[109] br[109] wl[83] vdd gnd cell_6t
Xbit_r84_c109 bl[109] br[109] wl[84] vdd gnd cell_6t
Xbit_r85_c109 bl[109] br[109] wl[85] vdd gnd cell_6t
Xbit_r86_c109 bl[109] br[109] wl[86] vdd gnd cell_6t
Xbit_r87_c109 bl[109] br[109] wl[87] vdd gnd cell_6t
Xbit_r88_c109 bl[109] br[109] wl[88] vdd gnd cell_6t
Xbit_r89_c109 bl[109] br[109] wl[89] vdd gnd cell_6t
Xbit_r90_c109 bl[109] br[109] wl[90] vdd gnd cell_6t
Xbit_r91_c109 bl[109] br[109] wl[91] vdd gnd cell_6t
Xbit_r92_c109 bl[109] br[109] wl[92] vdd gnd cell_6t
Xbit_r93_c109 bl[109] br[109] wl[93] vdd gnd cell_6t
Xbit_r94_c109 bl[109] br[109] wl[94] vdd gnd cell_6t
Xbit_r95_c109 bl[109] br[109] wl[95] vdd gnd cell_6t
Xbit_r96_c109 bl[109] br[109] wl[96] vdd gnd cell_6t
Xbit_r97_c109 bl[109] br[109] wl[97] vdd gnd cell_6t
Xbit_r98_c109 bl[109] br[109] wl[98] vdd gnd cell_6t
Xbit_r99_c109 bl[109] br[109] wl[99] vdd gnd cell_6t
Xbit_r100_c109 bl[109] br[109] wl[100] vdd gnd cell_6t
Xbit_r101_c109 bl[109] br[109] wl[101] vdd gnd cell_6t
Xbit_r102_c109 bl[109] br[109] wl[102] vdd gnd cell_6t
Xbit_r103_c109 bl[109] br[109] wl[103] vdd gnd cell_6t
Xbit_r104_c109 bl[109] br[109] wl[104] vdd gnd cell_6t
Xbit_r105_c109 bl[109] br[109] wl[105] vdd gnd cell_6t
Xbit_r106_c109 bl[109] br[109] wl[106] vdd gnd cell_6t
Xbit_r107_c109 bl[109] br[109] wl[107] vdd gnd cell_6t
Xbit_r108_c109 bl[109] br[109] wl[108] vdd gnd cell_6t
Xbit_r109_c109 bl[109] br[109] wl[109] vdd gnd cell_6t
Xbit_r110_c109 bl[109] br[109] wl[110] vdd gnd cell_6t
Xbit_r111_c109 bl[109] br[109] wl[111] vdd gnd cell_6t
Xbit_r112_c109 bl[109] br[109] wl[112] vdd gnd cell_6t
Xbit_r113_c109 bl[109] br[109] wl[113] vdd gnd cell_6t
Xbit_r114_c109 bl[109] br[109] wl[114] vdd gnd cell_6t
Xbit_r115_c109 bl[109] br[109] wl[115] vdd gnd cell_6t
Xbit_r116_c109 bl[109] br[109] wl[116] vdd gnd cell_6t
Xbit_r117_c109 bl[109] br[109] wl[117] vdd gnd cell_6t
Xbit_r118_c109 bl[109] br[109] wl[118] vdd gnd cell_6t
Xbit_r119_c109 bl[109] br[109] wl[119] vdd gnd cell_6t
Xbit_r120_c109 bl[109] br[109] wl[120] vdd gnd cell_6t
Xbit_r121_c109 bl[109] br[109] wl[121] vdd gnd cell_6t
Xbit_r122_c109 bl[109] br[109] wl[122] vdd gnd cell_6t
Xbit_r123_c109 bl[109] br[109] wl[123] vdd gnd cell_6t
Xbit_r124_c109 bl[109] br[109] wl[124] vdd gnd cell_6t
Xbit_r125_c109 bl[109] br[109] wl[125] vdd gnd cell_6t
Xbit_r126_c109 bl[109] br[109] wl[126] vdd gnd cell_6t
Xbit_r127_c109 bl[109] br[109] wl[127] vdd gnd cell_6t
Xbit_r128_c109 bl[109] br[109] wl[128] vdd gnd cell_6t
Xbit_r129_c109 bl[109] br[109] wl[129] vdd gnd cell_6t
Xbit_r130_c109 bl[109] br[109] wl[130] vdd gnd cell_6t
Xbit_r131_c109 bl[109] br[109] wl[131] vdd gnd cell_6t
Xbit_r132_c109 bl[109] br[109] wl[132] vdd gnd cell_6t
Xbit_r133_c109 bl[109] br[109] wl[133] vdd gnd cell_6t
Xbit_r134_c109 bl[109] br[109] wl[134] vdd gnd cell_6t
Xbit_r135_c109 bl[109] br[109] wl[135] vdd gnd cell_6t
Xbit_r136_c109 bl[109] br[109] wl[136] vdd gnd cell_6t
Xbit_r137_c109 bl[109] br[109] wl[137] vdd gnd cell_6t
Xbit_r138_c109 bl[109] br[109] wl[138] vdd gnd cell_6t
Xbit_r139_c109 bl[109] br[109] wl[139] vdd gnd cell_6t
Xbit_r140_c109 bl[109] br[109] wl[140] vdd gnd cell_6t
Xbit_r141_c109 bl[109] br[109] wl[141] vdd gnd cell_6t
Xbit_r142_c109 bl[109] br[109] wl[142] vdd gnd cell_6t
Xbit_r143_c109 bl[109] br[109] wl[143] vdd gnd cell_6t
Xbit_r144_c109 bl[109] br[109] wl[144] vdd gnd cell_6t
Xbit_r145_c109 bl[109] br[109] wl[145] vdd gnd cell_6t
Xbit_r146_c109 bl[109] br[109] wl[146] vdd gnd cell_6t
Xbit_r147_c109 bl[109] br[109] wl[147] vdd gnd cell_6t
Xbit_r148_c109 bl[109] br[109] wl[148] vdd gnd cell_6t
Xbit_r149_c109 bl[109] br[109] wl[149] vdd gnd cell_6t
Xbit_r150_c109 bl[109] br[109] wl[150] vdd gnd cell_6t
Xbit_r151_c109 bl[109] br[109] wl[151] vdd gnd cell_6t
Xbit_r152_c109 bl[109] br[109] wl[152] vdd gnd cell_6t
Xbit_r153_c109 bl[109] br[109] wl[153] vdd gnd cell_6t
Xbit_r154_c109 bl[109] br[109] wl[154] vdd gnd cell_6t
Xbit_r155_c109 bl[109] br[109] wl[155] vdd gnd cell_6t
Xbit_r156_c109 bl[109] br[109] wl[156] vdd gnd cell_6t
Xbit_r157_c109 bl[109] br[109] wl[157] vdd gnd cell_6t
Xbit_r158_c109 bl[109] br[109] wl[158] vdd gnd cell_6t
Xbit_r159_c109 bl[109] br[109] wl[159] vdd gnd cell_6t
Xbit_r160_c109 bl[109] br[109] wl[160] vdd gnd cell_6t
Xbit_r161_c109 bl[109] br[109] wl[161] vdd gnd cell_6t
Xbit_r162_c109 bl[109] br[109] wl[162] vdd gnd cell_6t
Xbit_r163_c109 bl[109] br[109] wl[163] vdd gnd cell_6t
Xbit_r164_c109 bl[109] br[109] wl[164] vdd gnd cell_6t
Xbit_r165_c109 bl[109] br[109] wl[165] vdd gnd cell_6t
Xbit_r166_c109 bl[109] br[109] wl[166] vdd gnd cell_6t
Xbit_r167_c109 bl[109] br[109] wl[167] vdd gnd cell_6t
Xbit_r168_c109 bl[109] br[109] wl[168] vdd gnd cell_6t
Xbit_r169_c109 bl[109] br[109] wl[169] vdd gnd cell_6t
Xbit_r170_c109 bl[109] br[109] wl[170] vdd gnd cell_6t
Xbit_r171_c109 bl[109] br[109] wl[171] vdd gnd cell_6t
Xbit_r172_c109 bl[109] br[109] wl[172] vdd gnd cell_6t
Xbit_r173_c109 bl[109] br[109] wl[173] vdd gnd cell_6t
Xbit_r174_c109 bl[109] br[109] wl[174] vdd gnd cell_6t
Xbit_r175_c109 bl[109] br[109] wl[175] vdd gnd cell_6t
Xbit_r176_c109 bl[109] br[109] wl[176] vdd gnd cell_6t
Xbit_r177_c109 bl[109] br[109] wl[177] vdd gnd cell_6t
Xbit_r178_c109 bl[109] br[109] wl[178] vdd gnd cell_6t
Xbit_r179_c109 bl[109] br[109] wl[179] vdd gnd cell_6t
Xbit_r180_c109 bl[109] br[109] wl[180] vdd gnd cell_6t
Xbit_r181_c109 bl[109] br[109] wl[181] vdd gnd cell_6t
Xbit_r182_c109 bl[109] br[109] wl[182] vdd gnd cell_6t
Xbit_r183_c109 bl[109] br[109] wl[183] vdd gnd cell_6t
Xbit_r184_c109 bl[109] br[109] wl[184] vdd gnd cell_6t
Xbit_r185_c109 bl[109] br[109] wl[185] vdd gnd cell_6t
Xbit_r186_c109 bl[109] br[109] wl[186] vdd gnd cell_6t
Xbit_r187_c109 bl[109] br[109] wl[187] vdd gnd cell_6t
Xbit_r188_c109 bl[109] br[109] wl[188] vdd gnd cell_6t
Xbit_r189_c109 bl[109] br[109] wl[189] vdd gnd cell_6t
Xbit_r190_c109 bl[109] br[109] wl[190] vdd gnd cell_6t
Xbit_r191_c109 bl[109] br[109] wl[191] vdd gnd cell_6t
Xbit_r192_c109 bl[109] br[109] wl[192] vdd gnd cell_6t
Xbit_r193_c109 bl[109] br[109] wl[193] vdd gnd cell_6t
Xbit_r194_c109 bl[109] br[109] wl[194] vdd gnd cell_6t
Xbit_r195_c109 bl[109] br[109] wl[195] vdd gnd cell_6t
Xbit_r196_c109 bl[109] br[109] wl[196] vdd gnd cell_6t
Xbit_r197_c109 bl[109] br[109] wl[197] vdd gnd cell_6t
Xbit_r198_c109 bl[109] br[109] wl[198] vdd gnd cell_6t
Xbit_r199_c109 bl[109] br[109] wl[199] vdd gnd cell_6t
Xbit_r200_c109 bl[109] br[109] wl[200] vdd gnd cell_6t
Xbit_r201_c109 bl[109] br[109] wl[201] vdd gnd cell_6t
Xbit_r202_c109 bl[109] br[109] wl[202] vdd gnd cell_6t
Xbit_r203_c109 bl[109] br[109] wl[203] vdd gnd cell_6t
Xbit_r204_c109 bl[109] br[109] wl[204] vdd gnd cell_6t
Xbit_r205_c109 bl[109] br[109] wl[205] vdd gnd cell_6t
Xbit_r206_c109 bl[109] br[109] wl[206] vdd gnd cell_6t
Xbit_r207_c109 bl[109] br[109] wl[207] vdd gnd cell_6t
Xbit_r208_c109 bl[109] br[109] wl[208] vdd gnd cell_6t
Xbit_r209_c109 bl[109] br[109] wl[209] vdd gnd cell_6t
Xbit_r210_c109 bl[109] br[109] wl[210] vdd gnd cell_6t
Xbit_r211_c109 bl[109] br[109] wl[211] vdd gnd cell_6t
Xbit_r212_c109 bl[109] br[109] wl[212] vdd gnd cell_6t
Xbit_r213_c109 bl[109] br[109] wl[213] vdd gnd cell_6t
Xbit_r214_c109 bl[109] br[109] wl[214] vdd gnd cell_6t
Xbit_r215_c109 bl[109] br[109] wl[215] vdd gnd cell_6t
Xbit_r216_c109 bl[109] br[109] wl[216] vdd gnd cell_6t
Xbit_r217_c109 bl[109] br[109] wl[217] vdd gnd cell_6t
Xbit_r218_c109 bl[109] br[109] wl[218] vdd gnd cell_6t
Xbit_r219_c109 bl[109] br[109] wl[219] vdd gnd cell_6t
Xbit_r220_c109 bl[109] br[109] wl[220] vdd gnd cell_6t
Xbit_r221_c109 bl[109] br[109] wl[221] vdd gnd cell_6t
Xbit_r222_c109 bl[109] br[109] wl[222] vdd gnd cell_6t
Xbit_r223_c109 bl[109] br[109] wl[223] vdd gnd cell_6t
Xbit_r224_c109 bl[109] br[109] wl[224] vdd gnd cell_6t
Xbit_r225_c109 bl[109] br[109] wl[225] vdd gnd cell_6t
Xbit_r226_c109 bl[109] br[109] wl[226] vdd gnd cell_6t
Xbit_r227_c109 bl[109] br[109] wl[227] vdd gnd cell_6t
Xbit_r228_c109 bl[109] br[109] wl[228] vdd gnd cell_6t
Xbit_r229_c109 bl[109] br[109] wl[229] vdd gnd cell_6t
Xbit_r230_c109 bl[109] br[109] wl[230] vdd gnd cell_6t
Xbit_r231_c109 bl[109] br[109] wl[231] vdd gnd cell_6t
Xbit_r232_c109 bl[109] br[109] wl[232] vdd gnd cell_6t
Xbit_r233_c109 bl[109] br[109] wl[233] vdd gnd cell_6t
Xbit_r234_c109 bl[109] br[109] wl[234] vdd gnd cell_6t
Xbit_r235_c109 bl[109] br[109] wl[235] vdd gnd cell_6t
Xbit_r236_c109 bl[109] br[109] wl[236] vdd gnd cell_6t
Xbit_r237_c109 bl[109] br[109] wl[237] vdd gnd cell_6t
Xbit_r238_c109 bl[109] br[109] wl[238] vdd gnd cell_6t
Xbit_r239_c109 bl[109] br[109] wl[239] vdd gnd cell_6t
Xbit_r240_c109 bl[109] br[109] wl[240] vdd gnd cell_6t
Xbit_r241_c109 bl[109] br[109] wl[241] vdd gnd cell_6t
Xbit_r242_c109 bl[109] br[109] wl[242] vdd gnd cell_6t
Xbit_r243_c109 bl[109] br[109] wl[243] vdd gnd cell_6t
Xbit_r244_c109 bl[109] br[109] wl[244] vdd gnd cell_6t
Xbit_r245_c109 bl[109] br[109] wl[245] vdd gnd cell_6t
Xbit_r246_c109 bl[109] br[109] wl[246] vdd gnd cell_6t
Xbit_r247_c109 bl[109] br[109] wl[247] vdd gnd cell_6t
Xbit_r248_c109 bl[109] br[109] wl[248] vdd gnd cell_6t
Xbit_r249_c109 bl[109] br[109] wl[249] vdd gnd cell_6t
Xbit_r250_c109 bl[109] br[109] wl[250] vdd gnd cell_6t
Xbit_r251_c109 bl[109] br[109] wl[251] vdd gnd cell_6t
Xbit_r252_c109 bl[109] br[109] wl[252] vdd gnd cell_6t
Xbit_r253_c109 bl[109] br[109] wl[253] vdd gnd cell_6t
Xbit_r254_c109 bl[109] br[109] wl[254] vdd gnd cell_6t
Xbit_r255_c109 bl[109] br[109] wl[255] vdd gnd cell_6t
Xbit_r0_c110 bl[110] br[110] wl[0] vdd gnd cell_6t
Xbit_r1_c110 bl[110] br[110] wl[1] vdd gnd cell_6t
Xbit_r2_c110 bl[110] br[110] wl[2] vdd gnd cell_6t
Xbit_r3_c110 bl[110] br[110] wl[3] vdd gnd cell_6t
Xbit_r4_c110 bl[110] br[110] wl[4] vdd gnd cell_6t
Xbit_r5_c110 bl[110] br[110] wl[5] vdd gnd cell_6t
Xbit_r6_c110 bl[110] br[110] wl[6] vdd gnd cell_6t
Xbit_r7_c110 bl[110] br[110] wl[7] vdd gnd cell_6t
Xbit_r8_c110 bl[110] br[110] wl[8] vdd gnd cell_6t
Xbit_r9_c110 bl[110] br[110] wl[9] vdd gnd cell_6t
Xbit_r10_c110 bl[110] br[110] wl[10] vdd gnd cell_6t
Xbit_r11_c110 bl[110] br[110] wl[11] vdd gnd cell_6t
Xbit_r12_c110 bl[110] br[110] wl[12] vdd gnd cell_6t
Xbit_r13_c110 bl[110] br[110] wl[13] vdd gnd cell_6t
Xbit_r14_c110 bl[110] br[110] wl[14] vdd gnd cell_6t
Xbit_r15_c110 bl[110] br[110] wl[15] vdd gnd cell_6t
Xbit_r16_c110 bl[110] br[110] wl[16] vdd gnd cell_6t
Xbit_r17_c110 bl[110] br[110] wl[17] vdd gnd cell_6t
Xbit_r18_c110 bl[110] br[110] wl[18] vdd gnd cell_6t
Xbit_r19_c110 bl[110] br[110] wl[19] vdd gnd cell_6t
Xbit_r20_c110 bl[110] br[110] wl[20] vdd gnd cell_6t
Xbit_r21_c110 bl[110] br[110] wl[21] vdd gnd cell_6t
Xbit_r22_c110 bl[110] br[110] wl[22] vdd gnd cell_6t
Xbit_r23_c110 bl[110] br[110] wl[23] vdd gnd cell_6t
Xbit_r24_c110 bl[110] br[110] wl[24] vdd gnd cell_6t
Xbit_r25_c110 bl[110] br[110] wl[25] vdd gnd cell_6t
Xbit_r26_c110 bl[110] br[110] wl[26] vdd gnd cell_6t
Xbit_r27_c110 bl[110] br[110] wl[27] vdd gnd cell_6t
Xbit_r28_c110 bl[110] br[110] wl[28] vdd gnd cell_6t
Xbit_r29_c110 bl[110] br[110] wl[29] vdd gnd cell_6t
Xbit_r30_c110 bl[110] br[110] wl[30] vdd gnd cell_6t
Xbit_r31_c110 bl[110] br[110] wl[31] vdd gnd cell_6t
Xbit_r32_c110 bl[110] br[110] wl[32] vdd gnd cell_6t
Xbit_r33_c110 bl[110] br[110] wl[33] vdd gnd cell_6t
Xbit_r34_c110 bl[110] br[110] wl[34] vdd gnd cell_6t
Xbit_r35_c110 bl[110] br[110] wl[35] vdd gnd cell_6t
Xbit_r36_c110 bl[110] br[110] wl[36] vdd gnd cell_6t
Xbit_r37_c110 bl[110] br[110] wl[37] vdd gnd cell_6t
Xbit_r38_c110 bl[110] br[110] wl[38] vdd gnd cell_6t
Xbit_r39_c110 bl[110] br[110] wl[39] vdd gnd cell_6t
Xbit_r40_c110 bl[110] br[110] wl[40] vdd gnd cell_6t
Xbit_r41_c110 bl[110] br[110] wl[41] vdd gnd cell_6t
Xbit_r42_c110 bl[110] br[110] wl[42] vdd gnd cell_6t
Xbit_r43_c110 bl[110] br[110] wl[43] vdd gnd cell_6t
Xbit_r44_c110 bl[110] br[110] wl[44] vdd gnd cell_6t
Xbit_r45_c110 bl[110] br[110] wl[45] vdd gnd cell_6t
Xbit_r46_c110 bl[110] br[110] wl[46] vdd gnd cell_6t
Xbit_r47_c110 bl[110] br[110] wl[47] vdd gnd cell_6t
Xbit_r48_c110 bl[110] br[110] wl[48] vdd gnd cell_6t
Xbit_r49_c110 bl[110] br[110] wl[49] vdd gnd cell_6t
Xbit_r50_c110 bl[110] br[110] wl[50] vdd gnd cell_6t
Xbit_r51_c110 bl[110] br[110] wl[51] vdd gnd cell_6t
Xbit_r52_c110 bl[110] br[110] wl[52] vdd gnd cell_6t
Xbit_r53_c110 bl[110] br[110] wl[53] vdd gnd cell_6t
Xbit_r54_c110 bl[110] br[110] wl[54] vdd gnd cell_6t
Xbit_r55_c110 bl[110] br[110] wl[55] vdd gnd cell_6t
Xbit_r56_c110 bl[110] br[110] wl[56] vdd gnd cell_6t
Xbit_r57_c110 bl[110] br[110] wl[57] vdd gnd cell_6t
Xbit_r58_c110 bl[110] br[110] wl[58] vdd gnd cell_6t
Xbit_r59_c110 bl[110] br[110] wl[59] vdd gnd cell_6t
Xbit_r60_c110 bl[110] br[110] wl[60] vdd gnd cell_6t
Xbit_r61_c110 bl[110] br[110] wl[61] vdd gnd cell_6t
Xbit_r62_c110 bl[110] br[110] wl[62] vdd gnd cell_6t
Xbit_r63_c110 bl[110] br[110] wl[63] vdd gnd cell_6t
Xbit_r64_c110 bl[110] br[110] wl[64] vdd gnd cell_6t
Xbit_r65_c110 bl[110] br[110] wl[65] vdd gnd cell_6t
Xbit_r66_c110 bl[110] br[110] wl[66] vdd gnd cell_6t
Xbit_r67_c110 bl[110] br[110] wl[67] vdd gnd cell_6t
Xbit_r68_c110 bl[110] br[110] wl[68] vdd gnd cell_6t
Xbit_r69_c110 bl[110] br[110] wl[69] vdd gnd cell_6t
Xbit_r70_c110 bl[110] br[110] wl[70] vdd gnd cell_6t
Xbit_r71_c110 bl[110] br[110] wl[71] vdd gnd cell_6t
Xbit_r72_c110 bl[110] br[110] wl[72] vdd gnd cell_6t
Xbit_r73_c110 bl[110] br[110] wl[73] vdd gnd cell_6t
Xbit_r74_c110 bl[110] br[110] wl[74] vdd gnd cell_6t
Xbit_r75_c110 bl[110] br[110] wl[75] vdd gnd cell_6t
Xbit_r76_c110 bl[110] br[110] wl[76] vdd gnd cell_6t
Xbit_r77_c110 bl[110] br[110] wl[77] vdd gnd cell_6t
Xbit_r78_c110 bl[110] br[110] wl[78] vdd gnd cell_6t
Xbit_r79_c110 bl[110] br[110] wl[79] vdd gnd cell_6t
Xbit_r80_c110 bl[110] br[110] wl[80] vdd gnd cell_6t
Xbit_r81_c110 bl[110] br[110] wl[81] vdd gnd cell_6t
Xbit_r82_c110 bl[110] br[110] wl[82] vdd gnd cell_6t
Xbit_r83_c110 bl[110] br[110] wl[83] vdd gnd cell_6t
Xbit_r84_c110 bl[110] br[110] wl[84] vdd gnd cell_6t
Xbit_r85_c110 bl[110] br[110] wl[85] vdd gnd cell_6t
Xbit_r86_c110 bl[110] br[110] wl[86] vdd gnd cell_6t
Xbit_r87_c110 bl[110] br[110] wl[87] vdd gnd cell_6t
Xbit_r88_c110 bl[110] br[110] wl[88] vdd gnd cell_6t
Xbit_r89_c110 bl[110] br[110] wl[89] vdd gnd cell_6t
Xbit_r90_c110 bl[110] br[110] wl[90] vdd gnd cell_6t
Xbit_r91_c110 bl[110] br[110] wl[91] vdd gnd cell_6t
Xbit_r92_c110 bl[110] br[110] wl[92] vdd gnd cell_6t
Xbit_r93_c110 bl[110] br[110] wl[93] vdd gnd cell_6t
Xbit_r94_c110 bl[110] br[110] wl[94] vdd gnd cell_6t
Xbit_r95_c110 bl[110] br[110] wl[95] vdd gnd cell_6t
Xbit_r96_c110 bl[110] br[110] wl[96] vdd gnd cell_6t
Xbit_r97_c110 bl[110] br[110] wl[97] vdd gnd cell_6t
Xbit_r98_c110 bl[110] br[110] wl[98] vdd gnd cell_6t
Xbit_r99_c110 bl[110] br[110] wl[99] vdd gnd cell_6t
Xbit_r100_c110 bl[110] br[110] wl[100] vdd gnd cell_6t
Xbit_r101_c110 bl[110] br[110] wl[101] vdd gnd cell_6t
Xbit_r102_c110 bl[110] br[110] wl[102] vdd gnd cell_6t
Xbit_r103_c110 bl[110] br[110] wl[103] vdd gnd cell_6t
Xbit_r104_c110 bl[110] br[110] wl[104] vdd gnd cell_6t
Xbit_r105_c110 bl[110] br[110] wl[105] vdd gnd cell_6t
Xbit_r106_c110 bl[110] br[110] wl[106] vdd gnd cell_6t
Xbit_r107_c110 bl[110] br[110] wl[107] vdd gnd cell_6t
Xbit_r108_c110 bl[110] br[110] wl[108] vdd gnd cell_6t
Xbit_r109_c110 bl[110] br[110] wl[109] vdd gnd cell_6t
Xbit_r110_c110 bl[110] br[110] wl[110] vdd gnd cell_6t
Xbit_r111_c110 bl[110] br[110] wl[111] vdd gnd cell_6t
Xbit_r112_c110 bl[110] br[110] wl[112] vdd gnd cell_6t
Xbit_r113_c110 bl[110] br[110] wl[113] vdd gnd cell_6t
Xbit_r114_c110 bl[110] br[110] wl[114] vdd gnd cell_6t
Xbit_r115_c110 bl[110] br[110] wl[115] vdd gnd cell_6t
Xbit_r116_c110 bl[110] br[110] wl[116] vdd gnd cell_6t
Xbit_r117_c110 bl[110] br[110] wl[117] vdd gnd cell_6t
Xbit_r118_c110 bl[110] br[110] wl[118] vdd gnd cell_6t
Xbit_r119_c110 bl[110] br[110] wl[119] vdd gnd cell_6t
Xbit_r120_c110 bl[110] br[110] wl[120] vdd gnd cell_6t
Xbit_r121_c110 bl[110] br[110] wl[121] vdd gnd cell_6t
Xbit_r122_c110 bl[110] br[110] wl[122] vdd gnd cell_6t
Xbit_r123_c110 bl[110] br[110] wl[123] vdd gnd cell_6t
Xbit_r124_c110 bl[110] br[110] wl[124] vdd gnd cell_6t
Xbit_r125_c110 bl[110] br[110] wl[125] vdd gnd cell_6t
Xbit_r126_c110 bl[110] br[110] wl[126] vdd gnd cell_6t
Xbit_r127_c110 bl[110] br[110] wl[127] vdd gnd cell_6t
Xbit_r128_c110 bl[110] br[110] wl[128] vdd gnd cell_6t
Xbit_r129_c110 bl[110] br[110] wl[129] vdd gnd cell_6t
Xbit_r130_c110 bl[110] br[110] wl[130] vdd gnd cell_6t
Xbit_r131_c110 bl[110] br[110] wl[131] vdd gnd cell_6t
Xbit_r132_c110 bl[110] br[110] wl[132] vdd gnd cell_6t
Xbit_r133_c110 bl[110] br[110] wl[133] vdd gnd cell_6t
Xbit_r134_c110 bl[110] br[110] wl[134] vdd gnd cell_6t
Xbit_r135_c110 bl[110] br[110] wl[135] vdd gnd cell_6t
Xbit_r136_c110 bl[110] br[110] wl[136] vdd gnd cell_6t
Xbit_r137_c110 bl[110] br[110] wl[137] vdd gnd cell_6t
Xbit_r138_c110 bl[110] br[110] wl[138] vdd gnd cell_6t
Xbit_r139_c110 bl[110] br[110] wl[139] vdd gnd cell_6t
Xbit_r140_c110 bl[110] br[110] wl[140] vdd gnd cell_6t
Xbit_r141_c110 bl[110] br[110] wl[141] vdd gnd cell_6t
Xbit_r142_c110 bl[110] br[110] wl[142] vdd gnd cell_6t
Xbit_r143_c110 bl[110] br[110] wl[143] vdd gnd cell_6t
Xbit_r144_c110 bl[110] br[110] wl[144] vdd gnd cell_6t
Xbit_r145_c110 bl[110] br[110] wl[145] vdd gnd cell_6t
Xbit_r146_c110 bl[110] br[110] wl[146] vdd gnd cell_6t
Xbit_r147_c110 bl[110] br[110] wl[147] vdd gnd cell_6t
Xbit_r148_c110 bl[110] br[110] wl[148] vdd gnd cell_6t
Xbit_r149_c110 bl[110] br[110] wl[149] vdd gnd cell_6t
Xbit_r150_c110 bl[110] br[110] wl[150] vdd gnd cell_6t
Xbit_r151_c110 bl[110] br[110] wl[151] vdd gnd cell_6t
Xbit_r152_c110 bl[110] br[110] wl[152] vdd gnd cell_6t
Xbit_r153_c110 bl[110] br[110] wl[153] vdd gnd cell_6t
Xbit_r154_c110 bl[110] br[110] wl[154] vdd gnd cell_6t
Xbit_r155_c110 bl[110] br[110] wl[155] vdd gnd cell_6t
Xbit_r156_c110 bl[110] br[110] wl[156] vdd gnd cell_6t
Xbit_r157_c110 bl[110] br[110] wl[157] vdd gnd cell_6t
Xbit_r158_c110 bl[110] br[110] wl[158] vdd gnd cell_6t
Xbit_r159_c110 bl[110] br[110] wl[159] vdd gnd cell_6t
Xbit_r160_c110 bl[110] br[110] wl[160] vdd gnd cell_6t
Xbit_r161_c110 bl[110] br[110] wl[161] vdd gnd cell_6t
Xbit_r162_c110 bl[110] br[110] wl[162] vdd gnd cell_6t
Xbit_r163_c110 bl[110] br[110] wl[163] vdd gnd cell_6t
Xbit_r164_c110 bl[110] br[110] wl[164] vdd gnd cell_6t
Xbit_r165_c110 bl[110] br[110] wl[165] vdd gnd cell_6t
Xbit_r166_c110 bl[110] br[110] wl[166] vdd gnd cell_6t
Xbit_r167_c110 bl[110] br[110] wl[167] vdd gnd cell_6t
Xbit_r168_c110 bl[110] br[110] wl[168] vdd gnd cell_6t
Xbit_r169_c110 bl[110] br[110] wl[169] vdd gnd cell_6t
Xbit_r170_c110 bl[110] br[110] wl[170] vdd gnd cell_6t
Xbit_r171_c110 bl[110] br[110] wl[171] vdd gnd cell_6t
Xbit_r172_c110 bl[110] br[110] wl[172] vdd gnd cell_6t
Xbit_r173_c110 bl[110] br[110] wl[173] vdd gnd cell_6t
Xbit_r174_c110 bl[110] br[110] wl[174] vdd gnd cell_6t
Xbit_r175_c110 bl[110] br[110] wl[175] vdd gnd cell_6t
Xbit_r176_c110 bl[110] br[110] wl[176] vdd gnd cell_6t
Xbit_r177_c110 bl[110] br[110] wl[177] vdd gnd cell_6t
Xbit_r178_c110 bl[110] br[110] wl[178] vdd gnd cell_6t
Xbit_r179_c110 bl[110] br[110] wl[179] vdd gnd cell_6t
Xbit_r180_c110 bl[110] br[110] wl[180] vdd gnd cell_6t
Xbit_r181_c110 bl[110] br[110] wl[181] vdd gnd cell_6t
Xbit_r182_c110 bl[110] br[110] wl[182] vdd gnd cell_6t
Xbit_r183_c110 bl[110] br[110] wl[183] vdd gnd cell_6t
Xbit_r184_c110 bl[110] br[110] wl[184] vdd gnd cell_6t
Xbit_r185_c110 bl[110] br[110] wl[185] vdd gnd cell_6t
Xbit_r186_c110 bl[110] br[110] wl[186] vdd gnd cell_6t
Xbit_r187_c110 bl[110] br[110] wl[187] vdd gnd cell_6t
Xbit_r188_c110 bl[110] br[110] wl[188] vdd gnd cell_6t
Xbit_r189_c110 bl[110] br[110] wl[189] vdd gnd cell_6t
Xbit_r190_c110 bl[110] br[110] wl[190] vdd gnd cell_6t
Xbit_r191_c110 bl[110] br[110] wl[191] vdd gnd cell_6t
Xbit_r192_c110 bl[110] br[110] wl[192] vdd gnd cell_6t
Xbit_r193_c110 bl[110] br[110] wl[193] vdd gnd cell_6t
Xbit_r194_c110 bl[110] br[110] wl[194] vdd gnd cell_6t
Xbit_r195_c110 bl[110] br[110] wl[195] vdd gnd cell_6t
Xbit_r196_c110 bl[110] br[110] wl[196] vdd gnd cell_6t
Xbit_r197_c110 bl[110] br[110] wl[197] vdd gnd cell_6t
Xbit_r198_c110 bl[110] br[110] wl[198] vdd gnd cell_6t
Xbit_r199_c110 bl[110] br[110] wl[199] vdd gnd cell_6t
Xbit_r200_c110 bl[110] br[110] wl[200] vdd gnd cell_6t
Xbit_r201_c110 bl[110] br[110] wl[201] vdd gnd cell_6t
Xbit_r202_c110 bl[110] br[110] wl[202] vdd gnd cell_6t
Xbit_r203_c110 bl[110] br[110] wl[203] vdd gnd cell_6t
Xbit_r204_c110 bl[110] br[110] wl[204] vdd gnd cell_6t
Xbit_r205_c110 bl[110] br[110] wl[205] vdd gnd cell_6t
Xbit_r206_c110 bl[110] br[110] wl[206] vdd gnd cell_6t
Xbit_r207_c110 bl[110] br[110] wl[207] vdd gnd cell_6t
Xbit_r208_c110 bl[110] br[110] wl[208] vdd gnd cell_6t
Xbit_r209_c110 bl[110] br[110] wl[209] vdd gnd cell_6t
Xbit_r210_c110 bl[110] br[110] wl[210] vdd gnd cell_6t
Xbit_r211_c110 bl[110] br[110] wl[211] vdd gnd cell_6t
Xbit_r212_c110 bl[110] br[110] wl[212] vdd gnd cell_6t
Xbit_r213_c110 bl[110] br[110] wl[213] vdd gnd cell_6t
Xbit_r214_c110 bl[110] br[110] wl[214] vdd gnd cell_6t
Xbit_r215_c110 bl[110] br[110] wl[215] vdd gnd cell_6t
Xbit_r216_c110 bl[110] br[110] wl[216] vdd gnd cell_6t
Xbit_r217_c110 bl[110] br[110] wl[217] vdd gnd cell_6t
Xbit_r218_c110 bl[110] br[110] wl[218] vdd gnd cell_6t
Xbit_r219_c110 bl[110] br[110] wl[219] vdd gnd cell_6t
Xbit_r220_c110 bl[110] br[110] wl[220] vdd gnd cell_6t
Xbit_r221_c110 bl[110] br[110] wl[221] vdd gnd cell_6t
Xbit_r222_c110 bl[110] br[110] wl[222] vdd gnd cell_6t
Xbit_r223_c110 bl[110] br[110] wl[223] vdd gnd cell_6t
Xbit_r224_c110 bl[110] br[110] wl[224] vdd gnd cell_6t
Xbit_r225_c110 bl[110] br[110] wl[225] vdd gnd cell_6t
Xbit_r226_c110 bl[110] br[110] wl[226] vdd gnd cell_6t
Xbit_r227_c110 bl[110] br[110] wl[227] vdd gnd cell_6t
Xbit_r228_c110 bl[110] br[110] wl[228] vdd gnd cell_6t
Xbit_r229_c110 bl[110] br[110] wl[229] vdd gnd cell_6t
Xbit_r230_c110 bl[110] br[110] wl[230] vdd gnd cell_6t
Xbit_r231_c110 bl[110] br[110] wl[231] vdd gnd cell_6t
Xbit_r232_c110 bl[110] br[110] wl[232] vdd gnd cell_6t
Xbit_r233_c110 bl[110] br[110] wl[233] vdd gnd cell_6t
Xbit_r234_c110 bl[110] br[110] wl[234] vdd gnd cell_6t
Xbit_r235_c110 bl[110] br[110] wl[235] vdd gnd cell_6t
Xbit_r236_c110 bl[110] br[110] wl[236] vdd gnd cell_6t
Xbit_r237_c110 bl[110] br[110] wl[237] vdd gnd cell_6t
Xbit_r238_c110 bl[110] br[110] wl[238] vdd gnd cell_6t
Xbit_r239_c110 bl[110] br[110] wl[239] vdd gnd cell_6t
Xbit_r240_c110 bl[110] br[110] wl[240] vdd gnd cell_6t
Xbit_r241_c110 bl[110] br[110] wl[241] vdd gnd cell_6t
Xbit_r242_c110 bl[110] br[110] wl[242] vdd gnd cell_6t
Xbit_r243_c110 bl[110] br[110] wl[243] vdd gnd cell_6t
Xbit_r244_c110 bl[110] br[110] wl[244] vdd gnd cell_6t
Xbit_r245_c110 bl[110] br[110] wl[245] vdd gnd cell_6t
Xbit_r246_c110 bl[110] br[110] wl[246] vdd gnd cell_6t
Xbit_r247_c110 bl[110] br[110] wl[247] vdd gnd cell_6t
Xbit_r248_c110 bl[110] br[110] wl[248] vdd gnd cell_6t
Xbit_r249_c110 bl[110] br[110] wl[249] vdd gnd cell_6t
Xbit_r250_c110 bl[110] br[110] wl[250] vdd gnd cell_6t
Xbit_r251_c110 bl[110] br[110] wl[251] vdd gnd cell_6t
Xbit_r252_c110 bl[110] br[110] wl[252] vdd gnd cell_6t
Xbit_r253_c110 bl[110] br[110] wl[253] vdd gnd cell_6t
Xbit_r254_c110 bl[110] br[110] wl[254] vdd gnd cell_6t
Xbit_r255_c110 bl[110] br[110] wl[255] vdd gnd cell_6t
Xbit_r0_c111 bl[111] br[111] wl[0] vdd gnd cell_6t
Xbit_r1_c111 bl[111] br[111] wl[1] vdd gnd cell_6t
Xbit_r2_c111 bl[111] br[111] wl[2] vdd gnd cell_6t
Xbit_r3_c111 bl[111] br[111] wl[3] vdd gnd cell_6t
Xbit_r4_c111 bl[111] br[111] wl[4] vdd gnd cell_6t
Xbit_r5_c111 bl[111] br[111] wl[5] vdd gnd cell_6t
Xbit_r6_c111 bl[111] br[111] wl[6] vdd gnd cell_6t
Xbit_r7_c111 bl[111] br[111] wl[7] vdd gnd cell_6t
Xbit_r8_c111 bl[111] br[111] wl[8] vdd gnd cell_6t
Xbit_r9_c111 bl[111] br[111] wl[9] vdd gnd cell_6t
Xbit_r10_c111 bl[111] br[111] wl[10] vdd gnd cell_6t
Xbit_r11_c111 bl[111] br[111] wl[11] vdd gnd cell_6t
Xbit_r12_c111 bl[111] br[111] wl[12] vdd gnd cell_6t
Xbit_r13_c111 bl[111] br[111] wl[13] vdd gnd cell_6t
Xbit_r14_c111 bl[111] br[111] wl[14] vdd gnd cell_6t
Xbit_r15_c111 bl[111] br[111] wl[15] vdd gnd cell_6t
Xbit_r16_c111 bl[111] br[111] wl[16] vdd gnd cell_6t
Xbit_r17_c111 bl[111] br[111] wl[17] vdd gnd cell_6t
Xbit_r18_c111 bl[111] br[111] wl[18] vdd gnd cell_6t
Xbit_r19_c111 bl[111] br[111] wl[19] vdd gnd cell_6t
Xbit_r20_c111 bl[111] br[111] wl[20] vdd gnd cell_6t
Xbit_r21_c111 bl[111] br[111] wl[21] vdd gnd cell_6t
Xbit_r22_c111 bl[111] br[111] wl[22] vdd gnd cell_6t
Xbit_r23_c111 bl[111] br[111] wl[23] vdd gnd cell_6t
Xbit_r24_c111 bl[111] br[111] wl[24] vdd gnd cell_6t
Xbit_r25_c111 bl[111] br[111] wl[25] vdd gnd cell_6t
Xbit_r26_c111 bl[111] br[111] wl[26] vdd gnd cell_6t
Xbit_r27_c111 bl[111] br[111] wl[27] vdd gnd cell_6t
Xbit_r28_c111 bl[111] br[111] wl[28] vdd gnd cell_6t
Xbit_r29_c111 bl[111] br[111] wl[29] vdd gnd cell_6t
Xbit_r30_c111 bl[111] br[111] wl[30] vdd gnd cell_6t
Xbit_r31_c111 bl[111] br[111] wl[31] vdd gnd cell_6t
Xbit_r32_c111 bl[111] br[111] wl[32] vdd gnd cell_6t
Xbit_r33_c111 bl[111] br[111] wl[33] vdd gnd cell_6t
Xbit_r34_c111 bl[111] br[111] wl[34] vdd gnd cell_6t
Xbit_r35_c111 bl[111] br[111] wl[35] vdd gnd cell_6t
Xbit_r36_c111 bl[111] br[111] wl[36] vdd gnd cell_6t
Xbit_r37_c111 bl[111] br[111] wl[37] vdd gnd cell_6t
Xbit_r38_c111 bl[111] br[111] wl[38] vdd gnd cell_6t
Xbit_r39_c111 bl[111] br[111] wl[39] vdd gnd cell_6t
Xbit_r40_c111 bl[111] br[111] wl[40] vdd gnd cell_6t
Xbit_r41_c111 bl[111] br[111] wl[41] vdd gnd cell_6t
Xbit_r42_c111 bl[111] br[111] wl[42] vdd gnd cell_6t
Xbit_r43_c111 bl[111] br[111] wl[43] vdd gnd cell_6t
Xbit_r44_c111 bl[111] br[111] wl[44] vdd gnd cell_6t
Xbit_r45_c111 bl[111] br[111] wl[45] vdd gnd cell_6t
Xbit_r46_c111 bl[111] br[111] wl[46] vdd gnd cell_6t
Xbit_r47_c111 bl[111] br[111] wl[47] vdd gnd cell_6t
Xbit_r48_c111 bl[111] br[111] wl[48] vdd gnd cell_6t
Xbit_r49_c111 bl[111] br[111] wl[49] vdd gnd cell_6t
Xbit_r50_c111 bl[111] br[111] wl[50] vdd gnd cell_6t
Xbit_r51_c111 bl[111] br[111] wl[51] vdd gnd cell_6t
Xbit_r52_c111 bl[111] br[111] wl[52] vdd gnd cell_6t
Xbit_r53_c111 bl[111] br[111] wl[53] vdd gnd cell_6t
Xbit_r54_c111 bl[111] br[111] wl[54] vdd gnd cell_6t
Xbit_r55_c111 bl[111] br[111] wl[55] vdd gnd cell_6t
Xbit_r56_c111 bl[111] br[111] wl[56] vdd gnd cell_6t
Xbit_r57_c111 bl[111] br[111] wl[57] vdd gnd cell_6t
Xbit_r58_c111 bl[111] br[111] wl[58] vdd gnd cell_6t
Xbit_r59_c111 bl[111] br[111] wl[59] vdd gnd cell_6t
Xbit_r60_c111 bl[111] br[111] wl[60] vdd gnd cell_6t
Xbit_r61_c111 bl[111] br[111] wl[61] vdd gnd cell_6t
Xbit_r62_c111 bl[111] br[111] wl[62] vdd gnd cell_6t
Xbit_r63_c111 bl[111] br[111] wl[63] vdd gnd cell_6t
Xbit_r64_c111 bl[111] br[111] wl[64] vdd gnd cell_6t
Xbit_r65_c111 bl[111] br[111] wl[65] vdd gnd cell_6t
Xbit_r66_c111 bl[111] br[111] wl[66] vdd gnd cell_6t
Xbit_r67_c111 bl[111] br[111] wl[67] vdd gnd cell_6t
Xbit_r68_c111 bl[111] br[111] wl[68] vdd gnd cell_6t
Xbit_r69_c111 bl[111] br[111] wl[69] vdd gnd cell_6t
Xbit_r70_c111 bl[111] br[111] wl[70] vdd gnd cell_6t
Xbit_r71_c111 bl[111] br[111] wl[71] vdd gnd cell_6t
Xbit_r72_c111 bl[111] br[111] wl[72] vdd gnd cell_6t
Xbit_r73_c111 bl[111] br[111] wl[73] vdd gnd cell_6t
Xbit_r74_c111 bl[111] br[111] wl[74] vdd gnd cell_6t
Xbit_r75_c111 bl[111] br[111] wl[75] vdd gnd cell_6t
Xbit_r76_c111 bl[111] br[111] wl[76] vdd gnd cell_6t
Xbit_r77_c111 bl[111] br[111] wl[77] vdd gnd cell_6t
Xbit_r78_c111 bl[111] br[111] wl[78] vdd gnd cell_6t
Xbit_r79_c111 bl[111] br[111] wl[79] vdd gnd cell_6t
Xbit_r80_c111 bl[111] br[111] wl[80] vdd gnd cell_6t
Xbit_r81_c111 bl[111] br[111] wl[81] vdd gnd cell_6t
Xbit_r82_c111 bl[111] br[111] wl[82] vdd gnd cell_6t
Xbit_r83_c111 bl[111] br[111] wl[83] vdd gnd cell_6t
Xbit_r84_c111 bl[111] br[111] wl[84] vdd gnd cell_6t
Xbit_r85_c111 bl[111] br[111] wl[85] vdd gnd cell_6t
Xbit_r86_c111 bl[111] br[111] wl[86] vdd gnd cell_6t
Xbit_r87_c111 bl[111] br[111] wl[87] vdd gnd cell_6t
Xbit_r88_c111 bl[111] br[111] wl[88] vdd gnd cell_6t
Xbit_r89_c111 bl[111] br[111] wl[89] vdd gnd cell_6t
Xbit_r90_c111 bl[111] br[111] wl[90] vdd gnd cell_6t
Xbit_r91_c111 bl[111] br[111] wl[91] vdd gnd cell_6t
Xbit_r92_c111 bl[111] br[111] wl[92] vdd gnd cell_6t
Xbit_r93_c111 bl[111] br[111] wl[93] vdd gnd cell_6t
Xbit_r94_c111 bl[111] br[111] wl[94] vdd gnd cell_6t
Xbit_r95_c111 bl[111] br[111] wl[95] vdd gnd cell_6t
Xbit_r96_c111 bl[111] br[111] wl[96] vdd gnd cell_6t
Xbit_r97_c111 bl[111] br[111] wl[97] vdd gnd cell_6t
Xbit_r98_c111 bl[111] br[111] wl[98] vdd gnd cell_6t
Xbit_r99_c111 bl[111] br[111] wl[99] vdd gnd cell_6t
Xbit_r100_c111 bl[111] br[111] wl[100] vdd gnd cell_6t
Xbit_r101_c111 bl[111] br[111] wl[101] vdd gnd cell_6t
Xbit_r102_c111 bl[111] br[111] wl[102] vdd gnd cell_6t
Xbit_r103_c111 bl[111] br[111] wl[103] vdd gnd cell_6t
Xbit_r104_c111 bl[111] br[111] wl[104] vdd gnd cell_6t
Xbit_r105_c111 bl[111] br[111] wl[105] vdd gnd cell_6t
Xbit_r106_c111 bl[111] br[111] wl[106] vdd gnd cell_6t
Xbit_r107_c111 bl[111] br[111] wl[107] vdd gnd cell_6t
Xbit_r108_c111 bl[111] br[111] wl[108] vdd gnd cell_6t
Xbit_r109_c111 bl[111] br[111] wl[109] vdd gnd cell_6t
Xbit_r110_c111 bl[111] br[111] wl[110] vdd gnd cell_6t
Xbit_r111_c111 bl[111] br[111] wl[111] vdd gnd cell_6t
Xbit_r112_c111 bl[111] br[111] wl[112] vdd gnd cell_6t
Xbit_r113_c111 bl[111] br[111] wl[113] vdd gnd cell_6t
Xbit_r114_c111 bl[111] br[111] wl[114] vdd gnd cell_6t
Xbit_r115_c111 bl[111] br[111] wl[115] vdd gnd cell_6t
Xbit_r116_c111 bl[111] br[111] wl[116] vdd gnd cell_6t
Xbit_r117_c111 bl[111] br[111] wl[117] vdd gnd cell_6t
Xbit_r118_c111 bl[111] br[111] wl[118] vdd gnd cell_6t
Xbit_r119_c111 bl[111] br[111] wl[119] vdd gnd cell_6t
Xbit_r120_c111 bl[111] br[111] wl[120] vdd gnd cell_6t
Xbit_r121_c111 bl[111] br[111] wl[121] vdd gnd cell_6t
Xbit_r122_c111 bl[111] br[111] wl[122] vdd gnd cell_6t
Xbit_r123_c111 bl[111] br[111] wl[123] vdd gnd cell_6t
Xbit_r124_c111 bl[111] br[111] wl[124] vdd gnd cell_6t
Xbit_r125_c111 bl[111] br[111] wl[125] vdd gnd cell_6t
Xbit_r126_c111 bl[111] br[111] wl[126] vdd gnd cell_6t
Xbit_r127_c111 bl[111] br[111] wl[127] vdd gnd cell_6t
Xbit_r128_c111 bl[111] br[111] wl[128] vdd gnd cell_6t
Xbit_r129_c111 bl[111] br[111] wl[129] vdd gnd cell_6t
Xbit_r130_c111 bl[111] br[111] wl[130] vdd gnd cell_6t
Xbit_r131_c111 bl[111] br[111] wl[131] vdd gnd cell_6t
Xbit_r132_c111 bl[111] br[111] wl[132] vdd gnd cell_6t
Xbit_r133_c111 bl[111] br[111] wl[133] vdd gnd cell_6t
Xbit_r134_c111 bl[111] br[111] wl[134] vdd gnd cell_6t
Xbit_r135_c111 bl[111] br[111] wl[135] vdd gnd cell_6t
Xbit_r136_c111 bl[111] br[111] wl[136] vdd gnd cell_6t
Xbit_r137_c111 bl[111] br[111] wl[137] vdd gnd cell_6t
Xbit_r138_c111 bl[111] br[111] wl[138] vdd gnd cell_6t
Xbit_r139_c111 bl[111] br[111] wl[139] vdd gnd cell_6t
Xbit_r140_c111 bl[111] br[111] wl[140] vdd gnd cell_6t
Xbit_r141_c111 bl[111] br[111] wl[141] vdd gnd cell_6t
Xbit_r142_c111 bl[111] br[111] wl[142] vdd gnd cell_6t
Xbit_r143_c111 bl[111] br[111] wl[143] vdd gnd cell_6t
Xbit_r144_c111 bl[111] br[111] wl[144] vdd gnd cell_6t
Xbit_r145_c111 bl[111] br[111] wl[145] vdd gnd cell_6t
Xbit_r146_c111 bl[111] br[111] wl[146] vdd gnd cell_6t
Xbit_r147_c111 bl[111] br[111] wl[147] vdd gnd cell_6t
Xbit_r148_c111 bl[111] br[111] wl[148] vdd gnd cell_6t
Xbit_r149_c111 bl[111] br[111] wl[149] vdd gnd cell_6t
Xbit_r150_c111 bl[111] br[111] wl[150] vdd gnd cell_6t
Xbit_r151_c111 bl[111] br[111] wl[151] vdd gnd cell_6t
Xbit_r152_c111 bl[111] br[111] wl[152] vdd gnd cell_6t
Xbit_r153_c111 bl[111] br[111] wl[153] vdd gnd cell_6t
Xbit_r154_c111 bl[111] br[111] wl[154] vdd gnd cell_6t
Xbit_r155_c111 bl[111] br[111] wl[155] vdd gnd cell_6t
Xbit_r156_c111 bl[111] br[111] wl[156] vdd gnd cell_6t
Xbit_r157_c111 bl[111] br[111] wl[157] vdd gnd cell_6t
Xbit_r158_c111 bl[111] br[111] wl[158] vdd gnd cell_6t
Xbit_r159_c111 bl[111] br[111] wl[159] vdd gnd cell_6t
Xbit_r160_c111 bl[111] br[111] wl[160] vdd gnd cell_6t
Xbit_r161_c111 bl[111] br[111] wl[161] vdd gnd cell_6t
Xbit_r162_c111 bl[111] br[111] wl[162] vdd gnd cell_6t
Xbit_r163_c111 bl[111] br[111] wl[163] vdd gnd cell_6t
Xbit_r164_c111 bl[111] br[111] wl[164] vdd gnd cell_6t
Xbit_r165_c111 bl[111] br[111] wl[165] vdd gnd cell_6t
Xbit_r166_c111 bl[111] br[111] wl[166] vdd gnd cell_6t
Xbit_r167_c111 bl[111] br[111] wl[167] vdd gnd cell_6t
Xbit_r168_c111 bl[111] br[111] wl[168] vdd gnd cell_6t
Xbit_r169_c111 bl[111] br[111] wl[169] vdd gnd cell_6t
Xbit_r170_c111 bl[111] br[111] wl[170] vdd gnd cell_6t
Xbit_r171_c111 bl[111] br[111] wl[171] vdd gnd cell_6t
Xbit_r172_c111 bl[111] br[111] wl[172] vdd gnd cell_6t
Xbit_r173_c111 bl[111] br[111] wl[173] vdd gnd cell_6t
Xbit_r174_c111 bl[111] br[111] wl[174] vdd gnd cell_6t
Xbit_r175_c111 bl[111] br[111] wl[175] vdd gnd cell_6t
Xbit_r176_c111 bl[111] br[111] wl[176] vdd gnd cell_6t
Xbit_r177_c111 bl[111] br[111] wl[177] vdd gnd cell_6t
Xbit_r178_c111 bl[111] br[111] wl[178] vdd gnd cell_6t
Xbit_r179_c111 bl[111] br[111] wl[179] vdd gnd cell_6t
Xbit_r180_c111 bl[111] br[111] wl[180] vdd gnd cell_6t
Xbit_r181_c111 bl[111] br[111] wl[181] vdd gnd cell_6t
Xbit_r182_c111 bl[111] br[111] wl[182] vdd gnd cell_6t
Xbit_r183_c111 bl[111] br[111] wl[183] vdd gnd cell_6t
Xbit_r184_c111 bl[111] br[111] wl[184] vdd gnd cell_6t
Xbit_r185_c111 bl[111] br[111] wl[185] vdd gnd cell_6t
Xbit_r186_c111 bl[111] br[111] wl[186] vdd gnd cell_6t
Xbit_r187_c111 bl[111] br[111] wl[187] vdd gnd cell_6t
Xbit_r188_c111 bl[111] br[111] wl[188] vdd gnd cell_6t
Xbit_r189_c111 bl[111] br[111] wl[189] vdd gnd cell_6t
Xbit_r190_c111 bl[111] br[111] wl[190] vdd gnd cell_6t
Xbit_r191_c111 bl[111] br[111] wl[191] vdd gnd cell_6t
Xbit_r192_c111 bl[111] br[111] wl[192] vdd gnd cell_6t
Xbit_r193_c111 bl[111] br[111] wl[193] vdd gnd cell_6t
Xbit_r194_c111 bl[111] br[111] wl[194] vdd gnd cell_6t
Xbit_r195_c111 bl[111] br[111] wl[195] vdd gnd cell_6t
Xbit_r196_c111 bl[111] br[111] wl[196] vdd gnd cell_6t
Xbit_r197_c111 bl[111] br[111] wl[197] vdd gnd cell_6t
Xbit_r198_c111 bl[111] br[111] wl[198] vdd gnd cell_6t
Xbit_r199_c111 bl[111] br[111] wl[199] vdd gnd cell_6t
Xbit_r200_c111 bl[111] br[111] wl[200] vdd gnd cell_6t
Xbit_r201_c111 bl[111] br[111] wl[201] vdd gnd cell_6t
Xbit_r202_c111 bl[111] br[111] wl[202] vdd gnd cell_6t
Xbit_r203_c111 bl[111] br[111] wl[203] vdd gnd cell_6t
Xbit_r204_c111 bl[111] br[111] wl[204] vdd gnd cell_6t
Xbit_r205_c111 bl[111] br[111] wl[205] vdd gnd cell_6t
Xbit_r206_c111 bl[111] br[111] wl[206] vdd gnd cell_6t
Xbit_r207_c111 bl[111] br[111] wl[207] vdd gnd cell_6t
Xbit_r208_c111 bl[111] br[111] wl[208] vdd gnd cell_6t
Xbit_r209_c111 bl[111] br[111] wl[209] vdd gnd cell_6t
Xbit_r210_c111 bl[111] br[111] wl[210] vdd gnd cell_6t
Xbit_r211_c111 bl[111] br[111] wl[211] vdd gnd cell_6t
Xbit_r212_c111 bl[111] br[111] wl[212] vdd gnd cell_6t
Xbit_r213_c111 bl[111] br[111] wl[213] vdd gnd cell_6t
Xbit_r214_c111 bl[111] br[111] wl[214] vdd gnd cell_6t
Xbit_r215_c111 bl[111] br[111] wl[215] vdd gnd cell_6t
Xbit_r216_c111 bl[111] br[111] wl[216] vdd gnd cell_6t
Xbit_r217_c111 bl[111] br[111] wl[217] vdd gnd cell_6t
Xbit_r218_c111 bl[111] br[111] wl[218] vdd gnd cell_6t
Xbit_r219_c111 bl[111] br[111] wl[219] vdd gnd cell_6t
Xbit_r220_c111 bl[111] br[111] wl[220] vdd gnd cell_6t
Xbit_r221_c111 bl[111] br[111] wl[221] vdd gnd cell_6t
Xbit_r222_c111 bl[111] br[111] wl[222] vdd gnd cell_6t
Xbit_r223_c111 bl[111] br[111] wl[223] vdd gnd cell_6t
Xbit_r224_c111 bl[111] br[111] wl[224] vdd gnd cell_6t
Xbit_r225_c111 bl[111] br[111] wl[225] vdd gnd cell_6t
Xbit_r226_c111 bl[111] br[111] wl[226] vdd gnd cell_6t
Xbit_r227_c111 bl[111] br[111] wl[227] vdd gnd cell_6t
Xbit_r228_c111 bl[111] br[111] wl[228] vdd gnd cell_6t
Xbit_r229_c111 bl[111] br[111] wl[229] vdd gnd cell_6t
Xbit_r230_c111 bl[111] br[111] wl[230] vdd gnd cell_6t
Xbit_r231_c111 bl[111] br[111] wl[231] vdd gnd cell_6t
Xbit_r232_c111 bl[111] br[111] wl[232] vdd gnd cell_6t
Xbit_r233_c111 bl[111] br[111] wl[233] vdd gnd cell_6t
Xbit_r234_c111 bl[111] br[111] wl[234] vdd gnd cell_6t
Xbit_r235_c111 bl[111] br[111] wl[235] vdd gnd cell_6t
Xbit_r236_c111 bl[111] br[111] wl[236] vdd gnd cell_6t
Xbit_r237_c111 bl[111] br[111] wl[237] vdd gnd cell_6t
Xbit_r238_c111 bl[111] br[111] wl[238] vdd gnd cell_6t
Xbit_r239_c111 bl[111] br[111] wl[239] vdd gnd cell_6t
Xbit_r240_c111 bl[111] br[111] wl[240] vdd gnd cell_6t
Xbit_r241_c111 bl[111] br[111] wl[241] vdd gnd cell_6t
Xbit_r242_c111 bl[111] br[111] wl[242] vdd gnd cell_6t
Xbit_r243_c111 bl[111] br[111] wl[243] vdd gnd cell_6t
Xbit_r244_c111 bl[111] br[111] wl[244] vdd gnd cell_6t
Xbit_r245_c111 bl[111] br[111] wl[245] vdd gnd cell_6t
Xbit_r246_c111 bl[111] br[111] wl[246] vdd gnd cell_6t
Xbit_r247_c111 bl[111] br[111] wl[247] vdd gnd cell_6t
Xbit_r248_c111 bl[111] br[111] wl[248] vdd gnd cell_6t
Xbit_r249_c111 bl[111] br[111] wl[249] vdd gnd cell_6t
Xbit_r250_c111 bl[111] br[111] wl[250] vdd gnd cell_6t
Xbit_r251_c111 bl[111] br[111] wl[251] vdd gnd cell_6t
Xbit_r252_c111 bl[111] br[111] wl[252] vdd gnd cell_6t
Xbit_r253_c111 bl[111] br[111] wl[253] vdd gnd cell_6t
Xbit_r254_c111 bl[111] br[111] wl[254] vdd gnd cell_6t
Xbit_r255_c111 bl[111] br[111] wl[255] vdd gnd cell_6t
Xbit_r0_c112 bl[112] br[112] wl[0] vdd gnd cell_6t
Xbit_r1_c112 bl[112] br[112] wl[1] vdd gnd cell_6t
Xbit_r2_c112 bl[112] br[112] wl[2] vdd gnd cell_6t
Xbit_r3_c112 bl[112] br[112] wl[3] vdd gnd cell_6t
Xbit_r4_c112 bl[112] br[112] wl[4] vdd gnd cell_6t
Xbit_r5_c112 bl[112] br[112] wl[5] vdd gnd cell_6t
Xbit_r6_c112 bl[112] br[112] wl[6] vdd gnd cell_6t
Xbit_r7_c112 bl[112] br[112] wl[7] vdd gnd cell_6t
Xbit_r8_c112 bl[112] br[112] wl[8] vdd gnd cell_6t
Xbit_r9_c112 bl[112] br[112] wl[9] vdd gnd cell_6t
Xbit_r10_c112 bl[112] br[112] wl[10] vdd gnd cell_6t
Xbit_r11_c112 bl[112] br[112] wl[11] vdd gnd cell_6t
Xbit_r12_c112 bl[112] br[112] wl[12] vdd gnd cell_6t
Xbit_r13_c112 bl[112] br[112] wl[13] vdd gnd cell_6t
Xbit_r14_c112 bl[112] br[112] wl[14] vdd gnd cell_6t
Xbit_r15_c112 bl[112] br[112] wl[15] vdd gnd cell_6t
Xbit_r16_c112 bl[112] br[112] wl[16] vdd gnd cell_6t
Xbit_r17_c112 bl[112] br[112] wl[17] vdd gnd cell_6t
Xbit_r18_c112 bl[112] br[112] wl[18] vdd gnd cell_6t
Xbit_r19_c112 bl[112] br[112] wl[19] vdd gnd cell_6t
Xbit_r20_c112 bl[112] br[112] wl[20] vdd gnd cell_6t
Xbit_r21_c112 bl[112] br[112] wl[21] vdd gnd cell_6t
Xbit_r22_c112 bl[112] br[112] wl[22] vdd gnd cell_6t
Xbit_r23_c112 bl[112] br[112] wl[23] vdd gnd cell_6t
Xbit_r24_c112 bl[112] br[112] wl[24] vdd gnd cell_6t
Xbit_r25_c112 bl[112] br[112] wl[25] vdd gnd cell_6t
Xbit_r26_c112 bl[112] br[112] wl[26] vdd gnd cell_6t
Xbit_r27_c112 bl[112] br[112] wl[27] vdd gnd cell_6t
Xbit_r28_c112 bl[112] br[112] wl[28] vdd gnd cell_6t
Xbit_r29_c112 bl[112] br[112] wl[29] vdd gnd cell_6t
Xbit_r30_c112 bl[112] br[112] wl[30] vdd gnd cell_6t
Xbit_r31_c112 bl[112] br[112] wl[31] vdd gnd cell_6t
Xbit_r32_c112 bl[112] br[112] wl[32] vdd gnd cell_6t
Xbit_r33_c112 bl[112] br[112] wl[33] vdd gnd cell_6t
Xbit_r34_c112 bl[112] br[112] wl[34] vdd gnd cell_6t
Xbit_r35_c112 bl[112] br[112] wl[35] vdd gnd cell_6t
Xbit_r36_c112 bl[112] br[112] wl[36] vdd gnd cell_6t
Xbit_r37_c112 bl[112] br[112] wl[37] vdd gnd cell_6t
Xbit_r38_c112 bl[112] br[112] wl[38] vdd gnd cell_6t
Xbit_r39_c112 bl[112] br[112] wl[39] vdd gnd cell_6t
Xbit_r40_c112 bl[112] br[112] wl[40] vdd gnd cell_6t
Xbit_r41_c112 bl[112] br[112] wl[41] vdd gnd cell_6t
Xbit_r42_c112 bl[112] br[112] wl[42] vdd gnd cell_6t
Xbit_r43_c112 bl[112] br[112] wl[43] vdd gnd cell_6t
Xbit_r44_c112 bl[112] br[112] wl[44] vdd gnd cell_6t
Xbit_r45_c112 bl[112] br[112] wl[45] vdd gnd cell_6t
Xbit_r46_c112 bl[112] br[112] wl[46] vdd gnd cell_6t
Xbit_r47_c112 bl[112] br[112] wl[47] vdd gnd cell_6t
Xbit_r48_c112 bl[112] br[112] wl[48] vdd gnd cell_6t
Xbit_r49_c112 bl[112] br[112] wl[49] vdd gnd cell_6t
Xbit_r50_c112 bl[112] br[112] wl[50] vdd gnd cell_6t
Xbit_r51_c112 bl[112] br[112] wl[51] vdd gnd cell_6t
Xbit_r52_c112 bl[112] br[112] wl[52] vdd gnd cell_6t
Xbit_r53_c112 bl[112] br[112] wl[53] vdd gnd cell_6t
Xbit_r54_c112 bl[112] br[112] wl[54] vdd gnd cell_6t
Xbit_r55_c112 bl[112] br[112] wl[55] vdd gnd cell_6t
Xbit_r56_c112 bl[112] br[112] wl[56] vdd gnd cell_6t
Xbit_r57_c112 bl[112] br[112] wl[57] vdd gnd cell_6t
Xbit_r58_c112 bl[112] br[112] wl[58] vdd gnd cell_6t
Xbit_r59_c112 bl[112] br[112] wl[59] vdd gnd cell_6t
Xbit_r60_c112 bl[112] br[112] wl[60] vdd gnd cell_6t
Xbit_r61_c112 bl[112] br[112] wl[61] vdd gnd cell_6t
Xbit_r62_c112 bl[112] br[112] wl[62] vdd gnd cell_6t
Xbit_r63_c112 bl[112] br[112] wl[63] vdd gnd cell_6t
Xbit_r64_c112 bl[112] br[112] wl[64] vdd gnd cell_6t
Xbit_r65_c112 bl[112] br[112] wl[65] vdd gnd cell_6t
Xbit_r66_c112 bl[112] br[112] wl[66] vdd gnd cell_6t
Xbit_r67_c112 bl[112] br[112] wl[67] vdd gnd cell_6t
Xbit_r68_c112 bl[112] br[112] wl[68] vdd gnd cell_6t
Xbit_r69_c112 bl[112] br[112] wl[69] vdd gnd cell_6t
Xbit_r70_c112 bl[112] br[112] wl[70] vdd gnd cell_6t
Xbit_r71_c112 bl[112] br[112] wl[71] vdd gnd cell_6t
Xbit_r72_c112 bl[112] br[112] wl[72] vdd gnd cell_6t
Xbit_r73_c112 bl[112] br[112] wl[73] vdd gnd cell_6t
Xbit_r74_c112 bl[112] br[112] wl[74] vdd gnd cell_6t
Xbit_r75_c112 bl[112] br[112] wl[75] vdd gnd cell_6t
Xbit_r76_c112 bl[112] br[112] wl[76] vdd gnd cell_6t
Xbit_r77_c112 bl[112] br[112] wl[77] vdd gnd cell_6t
Xbit_r78_c112 bl[112] br[112] wl[78] vdd gnd cell_6t
Xbit_r79_c112 bl[112] br[112] wl[79] vdd gnd cell_6t
Xbit_r80_c112 bl[112] br[112] wl[80] vdd gnd cell_6t
Xbit_r81_c112 bl[112] br[112] wl[81] vdd gnd cell_6t
Xbit_r82_c112 bl[112] br[112] wl[82] vdd gnd cell_6t
Xbit_r83_c112 bl[112] br[112] wl[83] vdd gnd cell_6t
Xbit_r84_c112 bl[112] br[112] wl[84] vdd gnd cell_6t
Xbit_r85_c112 bl[112] br[112] wl[85] vdd gnd cell_6t
Xbit_r86_c112 bl[112] br[112] wl[86] vdd gnd cell_6t
Xbit_r87_c112 bl[112] br[112] wl[87] vdd gnd cell_6t
Xbit_r88_c112 bl[112] br[112] wl[88] vdd gnd cell_6t
Xbit_r89_c112 bl[112] br[112] wl[89] vdd gnd cell_6t
Xbit_r90_c112 bl[112] br[112] wl[90] vdd gnd cell_6t
Xbit_r91_c112 bl[112] br[112] wl[91] vdd gnd cell_6t
Xbit_r92_c112 bl[112] br[112] wl[92] vdd gnd cell_6t
Xbit_r93_c112 bl[112] br[112] wl[93] vdd gnd cell_6t
Xbit_r94_c112 bl[112] br[112] wl[94] vdd gnd cell_6t
Xbit_r95_c112 bl[112] br[112] wl[95] vdd gnd cell_6t
Xbit_r96_c112 bl[112] br[112] wl[96] vdd gnd cell_6t
Xbit_r97_c112 bl[112] br[112] wl[97] vdd gnd cell_6t
Xbit_r98_c112 bl[112] br[112] wl[98] vdd gnd cell_6t
Xbit_r99_c112 bl[112] br[112] wl[99] vdd gnd cell_6t
Xbit_r100_c112 bl[112] br[112] wl[100] vdd gnd cell_6t
Xbit_r101_c112 bl[112] br[112] wl[101] vdd gnd cell_6t
Xbit_r102_c112 bl[112] br[112] wl[102] vdd gnd cell_6t
Xbit_r103_c112 bl[112] br[112] wl[103] vdd gnd cell_6t
Xbit_r104_c112 bl[112] br[112] wl[104] vdd gnd cell_6t
Xbit_r105_c112 bl[112] br[112] wl[105] vdd gnd cell_6t
Xbit_r106_c112 bl[112] br[112] wl[106] vdd gnd cell_6t
Xbit_r107_c112 bl[112] br[112] wl[107] vdd gnd cell_6t
Xbit_r108_c112 bl[112] br[112] wl[108] vdd gnd cell_6t
Xbit_r109_c112 bl[112] br[112] wl[109] vdd gnd cell_6t
Xbit_r110_c112 bl[112] br[112] wl[110] vdd gnd cell_6t
Xbit_r111_c112 bl[112] br[112] wl[111] vdd gnd cell_6t
Xbit_r112_c112 bl[112] br[112] wl[112] vdd gnd cell_6t
Xbit_r113_c112 bl[112] br[112] wl[113] vdd gnd cell_6t
Xbit_r114_c112 bl[112] br[112] wl[114] vdd gnd cell_6t
Xbit_r115_c112 bl[112] br[112] wl[115] vdd gnd cell_6t
Xbit_r116_c112 bl[112] br[112] wl[116] vdd gnd cell_6t
Xbit_r117_c112 bl[112] br[112] wl[117] vdd gnd cell_6t
Xbit_r118_c112 bl[112] br[112] wl[118] vdd gnd cell_6t
Xbit_r119_c112 bl[112] br[112] wl[119] vdd gnd cell_6t
Xbit_r120_c112 bl[112] br[112] wl[120] vdd gnd cell_6t
Xbit_r121_c112 bl[112] br[112] wl[121] vdd gnd cell_6t
Xbit_r122_c112 bl[112] br[112] wl[122] vdd gnd cell_6t
Xbit_r123_c112 bl[112] br[112] wl[123] vdd gnd cell_6t
Xbit_r124_c112 bl[112] br[112] wl[124] vdd gnd cell_6t
Xbit_r125_c112 bl[112] br[112] wl[125] vdd gnd cell_6t
Xbit_r126_c112 bl[112] br[112] wl[126] vdd gnd cell_6t
Xbit_r127_c112 bl[112] br[112] wl[127] vdd gnd cell_6t
Xbit_r128_c112 bl[112] br[112] wl[128] vdd gnd cell_6t
Xbit_r129_c112 bl[112] br[112] wl[129] vdd gnd cell_6t
Xbit_r130_c112 bl[112] br[112] wl[130] vdd gnd cell_6t
Xbit_r131_c112 bl[112] br[112] wl[131] vdd gnd cell_6t
Xbit_r132_c112 bl[112] br[112] wl[132] vdd gnd cell_6t
Xbit_r133_c112 bl[112] br[112] wl[133] vdd gnd cell_6t
Xbit_r134_c112 bl[112] br[112] wl[134] vdd gnd cell_6t
Xbit_r135_c112 bl[112] br[112] wl[135] vdd gnd cell_6t
Xbit_r136_c112 bl[112] br[112] wl[136] vdd gnd cell_6t
Xbit_r137_c112 bl[112] br[112] wl[137] vdd gnd cell_6t
Xbit_r138_c112 bl[112] br[112] wl[138] vdd gnd cell_6t
Xbit_r139_c112 bl[112] br[112] wl[139] vdd gnd cell_6t
Xbit_r140_c112 bl[112] br[112] wl[140] vdd gnd cell_6t
Xbit_r141_c112 bl[112] br[112] wl[141] vdd gnd cell_6t
Xbit_r142_c112 bl[112] br[112] wl[142] vdd gnd cell_6t
Xbit_r143_c112 bl[112] br[112] wl[143] vdd gnd cell_6t
Xbit_r144_c112 bl[112] br[112] wl[144] vdd gnd cell_6t
Xbit_r145_c112 bl[112] br[112] wl[145] vdd gnd cell_6t
Xbit_r146_c112 bl[112] br[112] wl[146] vdd gnd cell_6t
Xbit_r147_c112 bl[112] br[112] wl[147] vdd gnd cell_6t
Xbit_r148_c112 bl[112] br[112] wl[148] vdd gnd cell_6t
Xbit_r149_c112 bl[112] br[112] wl[149] vdd gnd cell_6t
Xbit_r150_c112 bl[112] br[112] wl[150] vdd gnd cell_6t
Xbit_r151_c112 bl[112] br[112] wl[151] vdd gnd cell_6t
Xbit_r152_c112 bl[112] br[112] wl[152] vdd gnd cell_6t
Xbit_r153_c112 bl[112] br[112] wl[153] vdd gnd cell_6t
Xbit_r154_c112 bl[112] br[112] wl[154] vdd gnd cell_6t
Xbit_r155_c112 bl[112] br[112] wl[155] vdd gnd cell_6t
Xbit_r156_c112 bl[112] br[112] wl[156] vdd gnd cell_6t
Xbit_r157_c112 bl[112] br[112] wl[157] vdd gnd cell_6t
Xbit_r158_c112 bl[112] br[112] wl[158] vdd gnd cell_6t
Xbit_r159_c112 bl[112] br[112] wl[159] vdd gnd cell_6t
Xbit_r160_c112 bl[112] br[112] wl[160] vdd gnd cell_6t
Xbit_r161_c112 bl[112] br[112] wl[161] vdd gnd cell_6t
Xbit_r162_c112 bl[112] br[112] wl[162] vdd gnd cell_6t
Xbit_r163_c112 bl[112] br[112] wl[163] vdd gnd cell_6t
Xbit_r164_c112 bl[112] br[112] wl[164] vdd gnd cell_6t
Xbit_r165_c112 bl[112] br[112] wl[165] vdd gnd cell_6t
Xbit_r166_c112 bl[112] br[112] wl[166] vdd gnd cell_6t
Xbit_r167_c112 bl[112] br[112] wl[167] vdd gnd cell_6t
Xbit_r168_c112 bl[112] br[112] wl[168] vdd gnd cell_6t
Xbit_r169_c112 bl[112] br[112] wl[169] vdd gnd cell_6t
Xbit_r170_c112 bl[112] br[112] wl[170] vdd gnd cell_6t
Xbit_r171_c112 bl[112] br[112] wl[171] vdd gnd cell_6t
Xbit_r172_c112 bl[112] br[112] wl[172] vdd gnd cell_6t
Xbit_r173_c112 bl[112] br[112] wl[173] vdd gnd cell_6t
Xbit_r174_c112 bl[112] br[112] wl[174] vdd gnd cell_6t
Xbit_r175_c112 bl[112] br[112] wl[175] vdd gnd cell_6t
Xbit_r176_c112 bl[112] br[112] wl[176] vdd gnd cell_6t
Xbit_r177_c112 bl[112] br[112] wl[177] vdd gnd cell_6t
Xbit_r178_c112 bl[112] br[112] wl[178] vdd gnd cell_6t
Xbit_r179_c112 bl[112] br[112] wl[179] vdd gnd cell_6t
Xbit_r180_c112 bl[112] br[112] wl[180] vdd gnd cell_6t
Xbit_r181_c112 bl[112] br[112] wl[181] vdd gnd cell_6t
Xbit_r182_c112 bl[112] br[112] wl[182] vdd gnd cell_6t
Xbit_r183_c112 bl[112] br[112] wl[183] vdd gnd cell_6t
Xbit_r184_c112 bl[112] br[112] wl[184] vdd gnd cell_6t
Xbit_r185_c112 bl[112] br[112] wl[185] vdd gnd cell_6t
Xbit_r186_c112 bl[112] br[112] wl[186] vdd gnd cell_6t
Xbit_r187_c112 bl[112] br[112] wl[187] vdd gnd cell_6t
Xbit_r188_c112 bl[112] br[112] wl[188] vdd gnd cell_6t
Xbit_r189_c112 bl[112] br[112] wl[189] vdd gnd cell_6t
Xbit_r190_c112 bl[112] br[112] wl[190] vdd gnd cell_6t
Xbit_r191_c112 bl[112] br[112] wl[191] vdd gnd cell_6t
Xbit_r192_c112 bl[112] br[112] wl[192] vdd gnd cell_6t
Xbit_r193_c112 bl[112] br[112] wl[193] vdd gnd cell_6t
Xbit_r194_c112 bl[112] br[112] wl[194] vdd gnd cell_6t
Xbit_r195_c112 bl[112] br[112] wl[195] vdd gnd cell_6t
Xbit_r196_c112 bl[112] br[112] wl[196] vdd gnd cell_6t
Xbit_r197_c112 bl[112] br[112] wl[197] vdd gnd cell_6t
Xbit_r198_c112 bl[112] br[112] wl[198] vdd gnd cell_6t
Xbit_r199_c112 bl[112] br[112] wl[199] vdd gnd cell_6t
Xbit_r200_c112 bl[112] br[112] wl[200] vdd gnd cell_6t
Xbit_r201_c112 bl[112] br[112] wl[201] vdd gnd cell_6t
Xbit_r202_c112 bl[112] br[112] wl[202] vdd gnd cell_6t
Xbit_r203_c112 bl[112] br[112] wl[203] vdd gnd cell_6t
Xbit_r204_c112 bl[112] br[112] wl[204] vdd gnd cell_6t
Xbit_r205_c112 bl[112] br[112] wl[205] vdd gnd cell_6t
Xbit_r206_c112 bl[112] br[112] wl[206] vdd gnd cell_6t
Xbit_r207_c112 bl[112] br[112] wl[207] vdd gnd cell_6t
Xbit_r208_c112 bl[112] br[112] wl[208] vdd gnd cell_6t
Xbit_r209_c112 bl[112] br[112] wl[209] vdd gnd cell_6t
Xbit_r210_c112 bl[112] br[112] wl[210] vdd gnd cell_6t
Xbit_r211_c112 bl[112] br[112] wl[211] vdd gnd cell_6t
Xbit_r212_c112 bl[112] br[112] wl[212] vdd gnd cell_6t
Xbit_r213_c112 bl[112] br[112] wl[213] vdd gnd cell_6t
Xbit_r214_c112 bl[112] br[112] wl[214] vdd gnd cell_6t
Xbit_r215_c112 bl[112] br[112] wl[215] vdd gnd cell_6t
Xbit_r216_c112 bl[112] br[112] wl[216] vdd gnd cell_6t
Xbit_r217_c112 bl[112] br[112] wl[217] vdd gnd cell_6t
Xbit_r218_c112 bl[112] br[112] wl[218] vdd gnd cell_6t
Xbit_r219_c112 bl[112] br[112] wl[219] vdd gnd cell_6t
Xbit_r220_c112 bl[112] br[112] wl[220] vdd gnd cell_6t
Xbit_r221_c112 bl[112] br[112] wl[221] vdd gnd cell_6t
Xbit_r222_c112 bl[112] br[112] wl[222] vdd gnd cell_6t
Xbit_r223_c112 bl[112] br[112] wl[223] vdd gnd cell_6t
Xbit_r224_c112 bl[112] br[112] wl[224] vdd gnd cell_6t
Xbit_r225_c112 bl[112] br[112] wl[225] vdd gnd cell_6t
Xbit_r226_c112 bl[112] br[112] wl[226] vdd gnd cell_6t
Xbit_r227_c112 bl[112] br[112] wl[227] vdd gnd cell_6t
Xbit_r228_c112 bl[112] br[112] wl[228] vdd gnd cell_6t
Xbit_r229_c112 bl[112] br[112] wl[229] vdd gnd cell_6t
Xbit_r230_c112 bl[112] br[112] wl[230] vdd gnd cell_6t
Xbit_r231_c112 bl[112] br[112] wl[231] vdd gnd cell_6t
Xbit_r232_c112 bl[112] br[112] wl[232] vdd gnd cell_6t
Xbit_r233_c112 bl[112] br[112] wl[233] vdd gnd cell_6t
Xbit_r234_c112 bl[112] br[112] wl[234] vdd gnd cell_6t
Xbit_r235_c112 bl[112] br[112] wl[235] vdd gnd cell_6t
Xbit_r236_c112 bl[112] br[112] wl[236] vdd gnd cell_6t
Xbit_r237_c112 bl[112] br[112] wl[237] vdd gnd cell_6t
Xbit_r238_c112 bl[112] br[112] wl[238] vdd gnd cell_6t
Xbit_r239_c112 bl[112] br[112] wl[239] vdd gnd cell_6t
Xbit_r240_c112 bl[112] br[112] wl[240] vdd gnd cell_6t
Xbit_r241_c112 bl[112] br[112] wl[241] vdd gnd cell_6t
Xbit_r242_c112 bl[112] br[112] wl[242] vdd gnd cell_6t
Xbit_r243_c112 bl[112] br[112] wl[243] vdd gnd cell_6t
Xbit_r244_c112 bl[112] br[112] wl[244] vdd gnd cell_6t
Xbit_r245_c112 bl[112] br[112] wl[245] vdd gnd cell_6t
Xbit_r246_c112 bl[112] br[112] wl[246] vdd gnd cell_6t
Xbit_r247_c112 bl[112] br[112] wl[247] vdd gnd cell_6t
Xbit_r248_c112 bl[112] br[112] wl[248] vdd gnd cell_6t
Xbit_r249_c112 bl[112] br[112] wl[249] vdd gnd cell_6t
Xbit_r250_c112 bl[112] br[112] wl[250] vdd gnd cell_6t
Xbit_r251_c112 bl[112] br[112] wl[251] vdd gnd cell_6t
Xbit_r252_c112 bl[112] br[112] wl[252] vdd gnd cell_6t
Xbit_r253_c112 bl[112] br[112] wl[253] vdd gnd cell_6t
Xbit_r254_c112 bl[112] br[112] wl[254] vdd gnd cell_6t
Xbit_r255_c112 bl[112] br[112] wl[255] vdd gnd cell_6t
Xbit_r0_c113 bl[113] br[113] wl[0] vdd gnd cell_6t
Xbit_r1_c113 bl[113] br[113] wl[1] vdd gnd cell_6t
Xbit_r2_c113 bl[113] br[113] wl[2] vdd gnd cell_6t
Xbit_r3_c113 bl[113] br[113] wl[3] vdd gnd cell_6t
Xbit_r4_c113 bl[113] br[113] wl[4] vdd gnd cell_6t
Xbit_r5_c113 bl[113] br[113] wl[5] vdd gnd cell_6t
Xbit_r6_c113 bl[113] br[113] wl[6] vdd gnd cell_6t
Xbit_r7_c113 bl[113] br[113] wl[7] vdd gnd cell_6t
Xbit_r8_c113 bl[113] br[113] wl[8] vdd gnd cell_6t
Xbit_r9_c113 bl[113] br[113] wl[9] vdd gnd cell_6t
Xbit_r10_c113 bl[113] br[113] wl[10] vdd gnd cell_6t
Xbit_r11_c113 bl[113] br[113] wl[11] vdd gnd cell_6t
Xbit_r12_c113 bl[113] br[113] wl[12] vdd gnd cell_6t
Xbit_r13_c113 bl[113] br[113] wl[13] vdd gnd cell_6t
Xbit_r14_c113 bl[113] br[113] wl[14] vdd gnd cell_6t
Xbit_r15_c113 bl[113] br[113] wl[15] vdd gnd cell_6t
Xbit_r16_c113 bl[113] br[113] wl[16] vdd gnd cell_6t
Xbit_r17_c113 bl[113] br[113] wl[17] vdd gnd cell_6t
Xbit_r18_c113 bl[113] br[113] wl[18] vdd gnd cell_6t
Xbit_r19_c113 bl[113] br[113] wl[19] vdd gnd cell_6t
Xbit_r20_c113 bl[113] br[113] wl[20] vdd gnd cell_6t
Xbit_r21_c113 bl[113] br[113] wl[21] vdd gnd cell_6t
Xbit_r22_c113 bl[113] br[113] wl[22] vdd gnd cell_6t
Xbit_r23_c113 bl[113] br[113] wl[23] vdd gnd cell_6t
Xbit_r24_c113 bl[113] br[113] wl[24] vdd gnd cell_6t
Xbit_r25_c113 bl[113] br[113] wl[25] vdd gnd cell_6t
Xbit_r26_c113 bl[113] br[113] wl[26] vdd gnd cell_6t
Xbit_r27_c113 bl[113] br[113] wl[27] vdd gnd cell_6t
Xbit_r28_c113 bl[113] br[113] wl[28] vdd gnd cell_6t
Xbit_r29_c113 bl[113] br[113] wl[29] vdd gnd cell_6t
Xbit_r30_c113 bl[113] br[113] wl[30] vdd gnd cell_6t
Xbit_r31_c113 bl[113] br[113] wl[31] vdd gnd cell_6t
Xbit_r32_c113 bl[113] br[113] wl[32] vdd gnd cell_6t
Xbit_r33_c113 bl[113] br[113] wl[33] vdd gnd cell_6t
Xbit_r34_c113 bl[113] br[113] wl[34] vdd gnd cell_6t
Xbit_r35_c113 bl[113] br[113] wl[35] vdd gnd cell_6t
Xbit_r36_c113 bl[113] br[113] wl[36] vdd gnd cell_6t
Xbit_r37_c113 bl[113] br[113] wl[37] vdd gnd cell_6t
Xbit_r38_c113 bl[113] br[113] wl[38] vdd gnd cell_6t
Xbit_r39_c113 bl[113] br[113] wl[39] vdd gnd cell_6t
Xbit_r40_c113 bl[113] br[113] wl[40] vdd gnd cell_6t
Xbit_r41_c113 bl[113] br[113] wl[41] vdd gnd cell_6t
Xbit_r42_c113 bl[113] br[113] wl[42] vdd gnd cell_6t
Xbit_r43_c113 bl[113] br[113] wl[43] vdd gnd cell_6t
Xbit_r44_c113 bl[113] br[113] wl[44] vdd gnd cell_6t
Xbit_r45_c113 bl[113] br[113] wl[45] vdd gnd cell_6t
Xbit_r46_c113 bl[113] br[113] wl[46] vdd gnd cell_6t
Xbit_r47_c113 bl[113] br[113] wl[47] vdd gnd cell_6t
Xbit_r48_c113 bl[113] br[113] wl[48] vdd gnd cell_6t
Xbit_r49_c113 bl[113] br[113] wl[49] vdd gnd cell_6t
Xbit_r50_c113 bl[113] br[113] wl[50] vdd gnd cell_6t
Xbit_r51_c113 bl[113] br[113] wl[51] vdd gnd cell_6t
Xbit_r52_c113 bl[113] br[113] wl[52] vdd gnd cell_6t
Xbit_r53_c113 bl[113] br[113] wl[53] vdd gnd cell_6t
Xbit_r54_c113 bl[113] br[113] wl[54] vdd gnd cell_6t
Xbit_r55_c113 bl[113] br[113] wl[55] vdd gnd cell_6t
Xbit_r56_c113 bl[113] br[113] wl[56] vdd gnd cell_6t
Xbit_r57_c113 bl[113] br[113] wl[57] vdd gnd cell_6t
Xbit_r58_c113 bl[113] br[113] wl[58] vdd gnd cell_6t
Xbit_r59_c113 bl[113] br[113] wl[59] vdd gnd cell_6t
Xbit_r60_c113 bl[113] br[113] wl[60] vdd gnd cell_6t
Xbit_r61_c113 bl[113] br[113] wl[61] vdd gnd cell_6t
Xbit_r62_c113 bl[113] br[113] wl[62] vdd gnd cell_6t
Xbit_r63_c113 bl[113] br[113] wl[63] vdd gnd cell_6t
Xbit_r64_c113 bl[113] br[113] wl[64] vdd gnd cell_6t
Xbit_r65_c113 bl[113] br[113] wl[65] vdd gnd cell_6t
Xbit_r66_c113 bl[113] br[113] wl[66] vdd gnd cell_6t
Xbit_r67_c113 bl[113] br[113] wl[67] vdd gnd cell_6t
Xbit_r68_c113 bl[113] br[113] wl[68] vdd gnd cell_6t
Xbit_r69_c113 bl[113] br[113] wl[69] vdd gnd cell_6t
Xbit_r70_c113 bl[113] br[113] wl[70] vdd gnd cell_6t
Xbit_r71_c113 bl[113] br[113] wl[71] vdd gnd cell_6t
Xbit_r72_c113 bl[113] br[113] wl[72] vdd gnd cell_6t
Xbit_r73_c113 bl[113] br[113] wl[73] vdd gnd cell_6t
Xbit_r74_c113 bl[113] br[113] wl[74] vdd gnd cell_6t
Xbit_r75_c113 bl[113] br[113] wl[75] vdd gnd cell_6t
Xbit_r76_c113 bl[113] br[113] wl[76] vdd gnd cell_6t
Xbit_r77_c113 bl[113] br[113] wl[77] vdd gnd cell_6t
Xbit_r78_c113 bl[113] br[113] wl[78] vdd gnd cell_6t
Xbit_r79_c113 bl[113] br[113] wl[79] vdd gnd cell_6t
Xbit_r80_c113 bl[113] br[113] wl[80] vdd gnd cell_6t
Xbit_r81_c113 bl[113] br[113] wl[81] vdd gnd cell_6t
Xbit_r82_c113 bl[113] br[113] wl[82] vdd gnd cell_6t
Xbit_r83_c113 bl[113] br[113] wl[83] vdd gnd cell_6t
Xbit_r84_c113 bl[113] br[113] wl[84] vdd gnd cell_6t
Xbit_r85_c113 bl[113] br[113] wl[85] vdd gnd cell_6t
Xbit_r86_c113 bl[113] br[113] wl[86] vdd gnd cell_6t
Xbit_r87_c113 bl[113] br[113] wl[87] vdd gnd cell_6t
Xbit_r88_c113 bl[113] br[113] wl[88] vdd gnd cell_6t
Xbit_r89_c113 bl[113] br[113] wl[89] vdd gnd cell_6t
Xbit_r90_c113 bl[113] br[113] wl[90] vdd gnd cell_6t
Xbit_r91_c113 bl[113] br[113] wl[91] vdd gnd cell_6t
Xbit_r92_c113 bl[113] br[113] wl[92] vdd gnd cell_6t
Xbit_r93_c113 bl[113] br[113] wl[93] vdd gnd cell_6t
Xbit_r94_c113 bl[113] br[113] wl[94] vdd gnd cell_6t
Xbit_r95_c113 bl[113] br[113] wl[95] vdd gnd cell_6t
Xbit_r96_c113 bl[113] br[113] wl[96] vdd gnd cell_6t
Xbit_r97_c113 bl[113] br[113] wl[97] vdd gnd cell_6t
Xbit_r98_c113 bl[113] br[113] wl[98] vdd gnd cell_6t
Xbit_r99_c113 bl[113] br[113] wl[99] vdd gnd cell_6t
Xbit_r100_c113 bl[113] br[113] wl[100] vdd gnd cell_6t
Xbit_r101_c113 bl[113] br[113] wl[101] vdd gnd cell_6t
Xbit_r102_c113 bl[113] br[113] wl[102] vdd gnd cell_6t
Xbit_r103_c113 bl[113] br[113] wl[103] vdd gnd cell_6t
Xbit_r104_c113 bl[113] br[113] wl[104] vdd gnd cell_6t
Xbit_r105_c113 bl[113] br[113] wl[105] vdd gnd cell_6t
Xbit_r106_c113 bl[113] br[113] wl[106] vdd gnd cell_6t
Xbit_r107_c113 bl[113] br[113] wl[107] vdd gnd cell_6t
Xbit_r108_c113 bl[113] br[113] wl[108] vdd gnd cell_6t
Xbit_r109_c113 bl[113] br[113] wl[109] vdd gnd cell_6t
Xbit_r110_c113 bl[113] br[113] wl[110] vdd gnd cell_6t
Xbit_r111_c113 bl[113] br[113] wl[111] vdd gnd cell_6t
Xbit_r112_c113 bl[113] br[113] wl[112] vdd gnd cell_6t
Xbit_r113_c113 bl[113] br[113] wl[113] vdd gnd cell_6t
Xbit_r114_c113 bl[113] br[113] wl[114] vdd gnd cell_6t
Xbit_r115_c113 bl[113] br[113] wl[115] vdd gnd cell_6t
Xbit_r116_c113 bl[113] br[113] wl[116] vdd gnd cell_6t
Xbit_r117_c113 bl[113] br[113] wl[117] vdd gnd cell_6t
Xbit_r118_c113 bl[113] br[113] wl[118] vdd gnd cell_6t
Xbit_r119_c113 bl[113] br[113] wl[119] vdd gnd cell_6t
Xbit_r120_c113 bl[113] br[113] wl[120] vdd gnd cell_6t
Xbit_r121_c113 bl[113] br[113] wl[121] vdd gnd cell_6t
Xbit_r122_c113 bl[113] br[113] wl[122] vdd gnd cell_6t
Xbit_r123_c113 bl[113] br[113] wl[123] vdd gnd cell_6t
Xbit_r124_c113 bl[113] br[113] wl[124] vdd gnd cell_6t
Xbit_r125_c113 bl[113] br[113] wl[125] vdd gnd cell_6t
Xbit_r126_c113 bl[113] br[113] wl[126] vdd gnd cell_6t
Xbit_r127_c113 bl[113] br[113] wl[127] vdd gnd cell_6t
Xbit_r128_c113 bl[113] br[113] wl[128] vdd gnd cell_6t
Xbit_r129_c113 bl[113] br[113] wl[129] vdd gnd cell_6t
Xbit_r130_c113 bl[113] br[113] wl[130] vdd gnd cell_6t
Xbit_r131_c113 bl[113] br[113] wl[131] vdd gnd cell_6t
Xbit_r132_c113 bl[113] br[113] wl[132] vdd gnd cell_6t
Xbit_r133_c113 bl[113] br[113] wl[133] vdd gnd cell_6t
Xbit_r134_c113 bl[113] br[113] wl[134] vdd gnd cell_6t
Xbit_r135_c113 bl[113] br[113] wl[135] vdd gnd cell_6t
Xbit_r136_c113 bl[113] br[113] wl[136] vdd gnd cell_6t
Xbit_r137_c113 bl[113] br[113] wl[137] vdd gnd cell_6t
Xbit_r138_c113 bl[113] br[113] wl[138] vdd gnd cell_6t
Xbit_r139_c113 bl[113] br[113] wl[139] vdd gnd cell_6t
Xbit_r140_c113 bl[113] br[113] wl[140] vdd gnd cell_6t
Xbit_r141_c113 bl[113] br[113] wl[141] vdd gnd cell_6t
Xbit_r142_c113 bl[113] br[113] wl[142] vdd gnd cell_6t
Xbit_r143_c113 bl[113] br[113] wl[143] vdd gnd cell_6t
Xbit_r144_c113 bl[113] br[113] wl[144] vdd gnd cell_6t
Xbit_r145_c113 bl[113] br[113] wl[145] vdd gnd cell_6t
Xbit_r146_c113 bl[113] br[113] wl[146] vdd gnd cell_6t
Xbit_r147_c113 bl[113] br[113] wl[147] vdd gnd cell_6t
Xbit_r148_c113 bl[113] br[113] wl[148] vdd gnd cell_6t
Xbit_r149_c113 bl[113] br[113] wl[149] vdd gnd cell_6t
Xbit_r150_c113 bl[113] br[113] wl[150] vdd gnd cell_6t
Xbit_r151_c113 bl[113] br[113] wl[151] vdd gnd cell_6t
Xbit_r152_c113 bl[113] br[113] wl[152] vdd gnd cell_6t
Xbit_r153_c113 bl[113] br[113] wl[153] vdd gnd cell_6t
Xbit_r154_c113 bl[113] br[113] wl[154] vdd gnd cell_6t
Xbit_r155_c113 bl[113] br[113] wl[155] vdd gnd cell_6t
Xbit_r156_c113 bl[113] br[113] wl[156] vdd gnd cell_6t
Xbit_r157_c113 bl[113] br[113] wl[157] vdd gnd cell_6t
Xbit_r158_c113 bl[113] br[113] wl[158] vdd gnd cell_6t
Xbit_r159_c113 bl[113] br[113] wl[159] vdd gnd cell_6t
Xbit_r160_c113 bl[113] br[113] wl[160] vdd gnd cell_6t
Xbit_r161_c113 bl[113] br[113] wl[161] vdd gnd cell_6t
Xbit_r162_c113 bl[113] br[113] wl[162] vdd gnd cell_6t
Xbit_r163_c113 bl[113] br[113] wl[163] vdd gnd cell_6t
Xbit_r164_c113 bl[113] br[113] wl[164] vdd gnd cell_6t
Xbit_r165_c113 bl[113] br[113] wl[165] vdd gnd cell_6t
Xbit_r166_c113 bl[113] br[113] wl[166] vdd gnd cell_6t
Xbit_r167_c113 bl[113] br[113] wl[167] vdd gnd cell_6t
Xbit_r168_c113 bl[113] br[113] wl[168] vdd gnd cell_6t
Xbit_r169_c113 bl[113] br[113] wl[169] vdd gnd cell_6t
Xbit_r170_c113 bl[113] br[113] wl[170] vdd gnd cell_6t
Xbit_r171_c113 bl[113] br[113] wl[171] vdd gnd cell_6t
Xbit_r172_c113 bl[113] br[113] wl[172] vdd gnd cell_6t
Xbit_r173_c113 bl[113] br[113] wl[173] vdd gnd cell_6t
Xbit_r174_c113 bl[113] br[113] wl[174] vdd gnd cell_6t
Xbit_r175_c113 bl[113] br[113] wl[175] vdd gnd cell_6t
Xbit_r176_c113 bl[113] br[113] wl[176] vdd gnd cell_6t
Xbit_r177_c113 bl[113] br[113] wl[177] vdd gnd cell_6t
Xbit_r178_c113 bl[113] br[113] wl[178] vdd gnd cell_6t
Xbit_r179_c113 bl[113] br[113] wl[179] vdd gnd cell_6t
Xbit_r180_c113 bl[113] br[113] wl[180] vdd gnd cell_6t
Xbit_r181_c113 bl[113] br[113] wl[181] vdd gnd cell_6t
Xbit_r182_c113 bl[113] br[113] wl[182] vdd gnd cell_6t
Xbit_r183_c113 bl[113] br[113] wl[183] vdd gnd cell_6t
Xbit_r184_c113 bl[113] br[113] wl[184] vdd gnd cell_6t
Xbit_r185_c113 bl[113] br[113] wl[185] vdd gnd cell_6t
Xbit_r186_c113 bl[113] br[113] wl[186] vdd gnd cell_6t
Xbit_r187_c113 bl[113] br[113] wl[187] vdd gnd cell_6t
Xbit_r188_c113 bl[113] br[113] wl[188] vdd gnd cell_6t
Xbit_r189_c113 bl[113] br[113] wl[189] vdd gnd cell_6t
Xbit_r190_c113 bl[113] br[113] wl[190] vdd gnd cell_6t
Xbit_r191_c113 bl[113] br[113] wl[191] vdd gnd cell_6t
Xbit_r192_c113 bl[113] br[113] wl[192] vdd gnd cell_6t
Xbit_r193_c113 bl[113] br[113] wl[193] vdd gnd cell_6t
Xbit_r194_c113 bl[113] br[113] wl[194] vdd gnd cell_6t
Xbit_r195_c113 bl[113] br[113] wl[195] vdd gnd cell_6t
Xbit_r196_c113 bl[113] br[113] wl[196] vdd gnd cell_6t
Xbit_r197_c113 bl[113] br[113] wl[197] vdd gnd cell_6t
Xbit_r198_c113 bl[113] br[113] wl[198] vdd gnd cell_6t
Xbit_r199_c113 bl[113] br[113] wl[199] vdd gnd cell_6t
Xbit_r200_c113 bl[113] br[113] wl[200] vdd gnd cell_6t
Xbit_r201_c113 bl[113] br[113] wl[201] vdd gnd cell_6t
Xbit_r202_c113 bl[113] br[113] wl[202] vdd gnd cell_6t
Xbit_r203_c113 bl[113] br[113] wl[203] vdd gnd cell_6t
Xbit_r204_c113 bl[113] br[113] wl[204] vdd gnd cell_6t
Xbit_r205_c113 bl[113] br[113] wl[205] vdd gnd cell_6t
Xbit_r206_c113 bl[113] br[113] wl[206] vdd gnd cell_6t
Xbit_r207_c113 bl[113] br[113] wl[207] vdd gnd cell_6t
Xbit_r208_c113 bl[113] br[113] wl[208] vdd gnd cell_6t
Xbit_r209_c113 bl[113] br[113] wl[209] vdd gnd cell_6t
Xbit_r210_c113 bl[113] br[113] wl[210] vdd gnd cell_6t
Xbit_r211_c113 bl[113] br[113] wl[211] vdd gnd cell_6t
Xbit_r212_c113 bl[113] br[113] wl[212] vdd gnd cell_6t
Xbit_r213_c113 bl[113] br[113] wl[213] vdd gnd cell_6t
Xbit_r214_c113 bl[113] br[113] wl[214] vdd gnd cell_6t
Xbit_r215_c113 bl[113] br[113] wl[215] vdd gnd cell_6t
Xbit_r216_c113 bl[113] br[113] wl[216] vdd gnd cell_6t
Xbit_r217_c113 bl[113] br[113] wl[217] vdd gnd cell_6t
Xbit_r218_c113 bl[113] br[113] wl[218] vdd gnd cell_6t
Xbit_r219_c113 bl[113] br[113] wl[219] vdd gnd cell_6t
Xbit_r220_c113 bl[113] br[113] wl[220] vdd gnd cell_6t
Xbit_r221_c113 bl[113] br[113] wl[221] vdd gnd cell_6t
Xbit_r222_c113 bl[113] br[113] wl[222] vdd gnd cell_6t
Xbit_r223_c113 bl[113] br[113] wl[223] vdd gnd cell_6t
Xbit_r224_c113 bl[113] br[113] wl[224] vdd gnd cell_6t
Xbit_r225_c113 bl[113] br[113] wl[225] vdd gnd cell_6t
Xbit_r226_c113 bl[113] br[113] wl[226] vdd gnd cell_6t
Xbit_r227_c113 bl[113] br[113] wl[227] vdd gnd cell_6t
Xbit_r228_c113 bl[113] br[113] wl[228] vdd gnd cell_6t
Xbit_r229_c113 bl[113] br[113] wl[229] vdd gnd cell_6t
Xbit_r230_c113 bl[113] br[113] wl[230] vdd gnd cell_6t
Xbit_r231_c113 bl[113] br[113] wl[231] vdd gnd cell_6t
Xbit_r232_c113 bl[113] br[113] wl[232] vdd gnd cell_6t
Xbit_r233_c113 bl[113] br[113] wl[233] vdd gnd cell_6t
Xbit_r234_c113 bl[113] br[113] wl[234] vdd gnd cell_6t
Xbit_r235_c113 bl[113] br[113] wl[235] vdd gnd cell_6t
Xbit_r236_c113 bl[113] br[113] wl[236] vdd gnd cell_6t
Xbit_r237_c113 bl[113] br[113] wl[237] vdd gnd cell_6t
Xbit_r238_c113 bl[113] br[113] wl[238] vdd gnd cell_6t
Xbit_r239_c113 bl[113] br[113] wl[239] vdd gnd cell_6t
Xbit_r240_c113 bl[113] br[113] wl[240] vdd gnd cell_6t
Xbit_r241_c113 bl[113] br[113] wl[241] vdd gnd cell_6t
Xbit_r242_c113 bl[113] br[113] wl[242] vdd gnd cell_6t
Xbit_r243_c113 bl[113] br[113] wl[243] vdd gnd cell_6t
Xbit_r244_c113 bl[113] br[113] wl[244] vdd gnd cell_6t
Xbit_r245_c113 bl[113] br[113] wl[245] vdd gnd cell_6t
Xbit_r246_c113 bl[113] br[113] wl[246] vdd gnd cell_6t
Xbit_r247_c113 bl[113] br[113] wl[247] vdd gnd cell_6t
Xbit_r248_c113 bl[113] br[113] wl[248] vdd gnd cell_6t
Xbit_r249_c113 bl[113] br[113] wl[249] vdd gnd cell_6t
Xbit_r250_c113 bl[113] br[113] wl[250] vdd gnd cell_6t
Xbit_r251_c113 bl[113] br[113] wl[251] vdd gnd cell_6t
Xbit_r252_c113 bl[113] br[113] wl[252] vdd gnd cell_6t
Xbit_r253_c113 bl[113] br[113] wl[253] vdd gnd cell_6t
Xbit_r254_c113 bl[113] br[113] wl[254] vdd gnd cell_6t
Xbit_r255_c113 bl[113] br[113] wl[255] vdd gnd cell_6t
Xbit_r0_c114 bl[114] br[114] wl[0] vdd gnd cell_6t
Xbit_r1_c114 bl[114] br[114] wl[1] vdd gnd cell_6t
Xbit_r2_c114 bl[114] br[114] wl[2] vdd gnd cell_6t
Xbit_r3_c114 bl[114] br[114] wl[3] vdd gnd cell_6t
Xbit_r4_c114 bl[114] br[114] wl[4] vdd gnd cell_6t
Xbit_r5_c114 bl[114] br[114] wl[5] vdd gnd cell_6t
Xbit_r6_c114 bl[114] br[114] wl[6] vdd gnd cell_6t
Xbit_r7_c114 bl[114] br[114] wl[7] vdd gnd cell_6t
Xbit_r8_c114 bl[114] br[114] wl[8] vdd gnd cell_6t
Xbit_r9_c114 bl[114] br[114] wl[9] vdd gnd cell_6t
Xbit_r10_c114 bl[114] br[114] wl[10] vdd gnd cell_6t
Xbit_r11_c114 bl[114] br[114] wl[11] vdd gnd cell_6t
Xbit_r12_c114 bl[114] br[114] wl[12] vdd gnd cell_6t
Xbit_r13_c114 bl[114] br[114] wl[13] vdd gnd cell_6t
Xbit_r14_c114 bl[114] br[114] wl[14] vdd gnd cell_6t
Xbit_r15_c114 bl[114] br[114] wl[15] vdd gnd cell_6t
Xbit_r16_c114 bl[114] br[114] wl[16] vdd gnd cell_6t
Xbit_r17_c114 bl[114] br[114] wl[17] vdd gnd cell_6t
Xbit_r18_c114 bl[114] br[114] wl[18] vdd gnd cell_6t
Xbit_r19_c114 bl[114] br[114] wl[19] vdd gnd cell_6t
Xbit_r20_c114 bl[114] br[114] wl[20] vdd gnd cell_6t
Xbit_r21_c114 bl[114] br[114] wl[21] vdd gnd cell_6t
Xbit_r22_c114 bl[114] br[114] wl[22] vdd gnd cell_6t
Xbit_r23_c114 bl[114] br[114] wl[23] vdd gnd cell_6t
Xbit_r24_c114 bl[114] br[114] wl[24] vdd gnd cell_6t
Xbit_r25_c114 bl[114] br[114] wl[25] vdd gnd cell_6t
Xbit_r26_c114 bl[114] br[114] wl[26] vdd gnd cell_6t
Xbit_r27_c114 bl[114] br[114] wl[27] vdd gnd cell_6t
Xbit_r28_c114 bl[114] br[114] wl[28] vdd gnd cell_6t
Xbit_r29_c114 bl[114] br[114] wl[29] vdd gnd cell_6t
Xbit_r30_c114 bl[114] br[114] wl[30] vdd gnd cell_6t
Xbit_r31_c114 bl[114] br[114] wl[31] vdd gnd cell_6t
Xbit_r32_c114 bl[114] br[114] wl[32] vdd gnd cell_6t
Xbit_r33_c114 bl[114] br[114] wl[33] vdd gnd cell_6t
Xbit_r34_c114 bl[114] br[114] wl[34] vdd gnd cell_6t
Xbit_r35_c114 bl[114] br[114] wl[35] vdd gnd cell_6t
Xbit_r36_c114 bl[114] br[114] wl[36] vdd gnd cell_6t
Xbit_r37_c114 bl[114] br[114] wl[37] vdd gnd cell_6t
Xbit_r38_c114 bl[114] br[114] wl[38] vdd gnd cell_6t
Xbit_r39_c114 bl[114] br[114] wl[39] vdd gnd cell_6t
Xbit_r40_c114 bl[114] br[114] wl[40] vdd gnd cell_6t
Xbit_r41_c114 bl[114] br[114] wl[41] vdd gnd cell_6t
Xbit_r42_c114 bl[114] br[114] wl[42] vdd gnd cell_6t
Xbit_r43_c114 bl[114] br[114] wl[43] vdd gnd cell_6t
Xbit_r44_c114 bl[114] br[114] wl[44] vdd gnd cell_6t
Xbit_r45_c114 bl[114] br[114] wl[45] vdd gnd cell_6t
Xbit_r46_c114 bl[114] br[114] wl[46] vdd gnd cell_6t
Xbit_r47_c114 bl[114] br[114] wl[47] vdd gnd cell_6t
Xbit_r48_c114 bl[114] br[114] wl[48] vdd gnd cell_6t
Xbit_r49_c114 bl[114] br[114] wl[49] vdd gnd cell_6t
Xbit_r50_c114 bl[114] br[114] wl[50] vdd gnd cell_6t
Xbit_r51_c114 bl[114] br[114] wl[51] vdd gnd cell_6t
Xbit_r52_c114 bl[114] br[114] wl[52] vdd gnd cell_6t
Xbit_r53_c114 bl[114] br[114] wl[53] vdd gnd cell_6t
Xbit_r54_c114 bl[114] br[114] wl[54] vdd gnd cell_6t
Xbit_r55_c114 bl[114] br[114] wl[55] vdd gnd cell_6t
Xbit_r56_c114 bl[114] br[114] wl[56] vdd gnd cell_6t
Xbit_r57_c114 bl[114] br[114] wl[57] vdd gnd cell_6t
Xbit_r58_c114 bl[114] br[114] wl[58] vdd gnd cell_6t
Xbit_r59_c114 bl[114] br[114] wl[59] vdd gnd cell_6t
Xbit_r60_c114 bl[114] br[114] wl[60] vdd gnd cell_6t
Xbit_r61_c114 bl[114] br[114] wl[61] vdd gnd cell_6t
Xbit_r62_c114 bl[114] br[114] wl[62] vdd gnd cell_6t
Xbit_r63_c114 bl[114] br[114] wl[63] vdd gnd cell_6t
Xbit_r64_c114 bl[114] br[114] wl[64] vdd gnd cell_6t
Xbit_r65_c114 bl[114] br[114] wl[65] vdd gnd cell_6t
Xbit_r66_c114 bl[114] br[114] wl[66] vdd gnd cell_6t
Xbit_r67_c114 bl[114] br[114] wl[67] vdd gnd cell_6t
Xbit_r68_c114 bl[114] br[114] wl[68] vdd gnd cell_6t
Xbit_r69_c114 bl[114] br[114] wl[69] vdd gnd cell_6t
Xbit_r70_c114 bl[114] br[114] wl[70] vdd gnd cell_6t
Xbit_r71_c114 bl[114] br[114] wl[71] vdd gnd cell_6t
Xbit_r72_c114 bl[114] br[114] wl[72] vdd gnd cell_6t
Xbit_r73_c114 bl[114] br[114] wl[73] vdd gnd cell_6t
Xbit_r74_c114 bl[114] br[114] wl[74] vdd gnd cell_6t
Xbit_r75_c114 bl[114] br[114] wl[75] vdd gnd cell_6t
Xbit_r76_c114 bl[114] br[114] wl[76] vdd gnd cell_6t
Xbit_r77_c114 bl[114] br[114] wl[77] vdd gnd cell_6t
Xbit_r78_c114 bl[114] br[114] wl[78] vdd gnd cell_6t
Xbit_r79_c114 bl[114] br[114] wl[79] vdd gnd cell_6t
Xbit_r80_c114 bl[114] br[114] wl[80] vdd gnd cell_6t
Xbit_r81_c114 bl[114] br[114] wl[81] vdd gnd cell_6t
Xbit_r82_c114 bl[114] br[114] wl[82] vdd gnd cell_6t
Xbit_r83_c114 bl[114] br[114] wl[83] vdd gnd cell_6t
Xbit_r84_c114 bl[114] br[114] wl[84] vdd gnd cell_6t
Xbit_r85_c114 bl[114] br[114] wl[85] vdd gnd cell_6t
Xbit_r86_c114 bl[114] br[114] wl[86] vdd gnd cell_6t
Xbit_r87_c114 bl[114] br[114] wl[87] vdd gnd cell_6t
Xbit_r88_c114 bl[114] br[114] wl[88] vdd gnd cell_6t
Xbit_r89_c114 bl[114] br[114] wl[89] vdd gnd cell_6t
Xbit_r90_c114 bl[114] br[114] wl[90] vdd gnd cell_6t
Xbit_r91_c114 bl[114] br[114] wl[91] vdd gnd cell_6t
Xbit_r92_c114 bl[114] br[114] wl[92] vdd gnd cell_6t
Xbit_r93_c114 bl[114] br[114] wl[93] vdd gnd cell_6t
Xbit_r94_c114 bl[114] br[114] wl[94] vdd gnd cell_6t
Xbit_r95_c114 bl[114] br[114] wl[95] vdd gnd cell_6t
Xbit_r96_c114 bl[114] br[114] wl[96] vdd gnd cell_6t
Xbit_r97_c114 bl[114] br[114] wl[97] vdd gnd cell_6t
Xbit_r98_c114 bl[114] br[114] wl[98] vdd gnd cell_6t
Xbit_r99_c114 bl[114] br[114] wl[99] vdd gnd cell_6t
Xbit_r100_c114 bl[114] br[114] wl[100] vdd gnd cell_6t
Xbit_r101_c114 bl[114] br[114] wl[101] vdd gnd cell_6t
Xbit_r102_c114 bl[114] br[114] wl[102] vdd gnd cell_6t
Xbit_r103_c114 bl[114] br[114] wl[103] vdd gnd cell_6t
Xbit_r104_c114 bl[114] br[114] wl[104] vdd gnd cell_6t
Xbit_r105_c114 bl[114] br[114] wl[105] vdd gnd cell_6t
Xbit_r106_c114 bl[114] br[114] wl[106] vdd gnd cell_6t
Xbit_r107_c114 bl[114] br[114] wl[107] vdd gnd cell_6t
Xbit_r108_c114 bl[114] br[114] wl[108] vdd gnd cell_6t
Xbit_r109_c114 bl[114] br[114] wl[109] vdd gnd cell_6t
Xbit_r110_c114 bl[114] br[114] wl[110] vdd gnd cell_6t
Xbit_r111_c114 bl[114] br[114] wl[111] vdd gnd cell_6t
Xbit_r112_c114 bl[114] br[114] wl[112] vdd gnd cell_6t
Xbit_r113_c114 bl[114] br[114] wl[113] vdd gnd cell_6t
Xbit_r114_c114 bl[114] br[114] wl[114] vdd gnd cell_6t
Xbit_r115_c114 bl[114] br[114] wl[115] vdd gnd cell_6t
Xbit_r116_c114 bl[114] br[114] wl[116] vdd gnd cell_6t
Xbit_r117_c114 bl[114] br[114] wl[117] vdd gnd cell_6t
Xbit_r118_c114 bl[114] br[114] wl[118] vdd gnd cell_6t
Xbit_r119_c114 bl[114] br[114] wl[119] vdd gnd cell_6t
Xbit_r120_c114 bl[114] br[114] wl[120] vdd gnd cell_6t
Xbit_r121_c114 bl[114] br[114] wl[121] vdd gnd cell_6t
Xbit_r122_c114 bl[114] br[114] wl[122] vdd gnd cell_6t
Xbit_r123_c114 bl[114] br[114] wl[123] vdd gnd cell_6t
Xbit_r124_c114 bl[114] br[114] wl[124] vdd gnd cell_6t
Xbit_r125_c114 bl[114] br[114] wl[125] vdd gnd cell_6t
Xbit_r126_c114 bl[114] br[114] wl[126] vdd gnd cell_6t
Xbit_r127_c114 bl[114] br[114] wl[127] vdd gnd cell_6t
Xbit_r128_c114 bl[114] br[114] wl[128] vdd gnd cell_6t
Xbit_r129_c114 bl[114] br[114] wl[129] vdd gnd cell_6t
Xbit_r130_c114 bl[114] br[114] wl[130] vdd gnd cell_6t
Xbit_r131_c114 bl[114] br[114] wl[131] vdd gnd cell_6t
Xbit_r132_c114 bl[114] br[114] wl[132] vdd gnd cell_6t
Xbit_r133_c114 bl[114] br[114] wl[133] vdd gnd cell_6t
Xbit_r134_c114 bl[114] br[114] wl[134] vdd gnd cell_6t
Xbit_r135_c114 bl[114] br[114] wl[135] vdd gnd cell_6t
Xbit_r136_c114 bl[114] br[114] wl[136] vdd gnd cell_6t
Xbit_r137_c114 bl[114] br[114] wl[137] vdd gnd cell_6t
Xbit_r138_c114 bl[114] br[114] wl[138] vdd gnd cell_6t
Xbit_r139_c114 bl[114] br[114] wl[139] vdd gnd cell_6t
Xbit_r140_c114 bl[114] br[114] wl[140] vdd gnd cell_6t
Xbit_r141_c114 bl[114] br[114] wl[141] vdd gnd cell_6t
Xbit_r142_c114 bl[114] br[114] wl[142] vdd gnd cell_6t
Xbit_r143_c114 bl[114] br[114] wl[143] vdd gnd cell_6t
Xbit_r144_c114 bl[114] br[114] wl[144] vdd gnd cell_6t
Xbit_r145_c114 bl[114] br[114] wl[145] vdd gnd cell_6t
Xbit_r146_c114 bl[114] br[114] wl[146] vdd gnd cell_6t
Xbit_r147_c114 bl[114] br[114] wl[147] vdd gnd cell_6t
Xbit_r148_c114 bl[114] br[114] wl[148] vdd gnd cell_6t
Xbit_r149_c114 bl[114] br[114] wl[149] vdd gnd cell_6t
Xbit_r150_c114 bl[114] br[114] wl[150] vdd gnd cell_6t
Xbit_r151_c114 bl[114] br[114] wl[151] vdd gnd cell_6t
Xbit_r152_c114 bl[114] br[114] wl[152] vdd gnd cell_6t
Xbit_r153_c114 bl[114] br[114] wl[153] vdd gnd cell_6t
Xbit_r154_c114 bl[114] br[114] wl[154] vdd gnd cell_6t
Xbit_r155_c114 bl[114] br[114] wl[155] vdd gnd cell_6t
Xbit_r156_c114 bl[114] br[114] wl[156] vdd gnd cell_6t
Xbit_r157_c114 bl[114] br[114] wl[157] vdd gnd cell_6t
Xbit_r158_c114 bl[114] br[114] wl[158] vdd gnd cell_6t
Xbit_r159_c114 bl[114] br[114] wl[159] vdd gnd cell_6t
Xbit_r160_c114 bl[114] br[114] wl[160] vdd gnd cell_6t
Xbit_r161_c114 bl[114] br[114] wl[161] vdd gnd cell_6t
Xbit_r162_c114 bl[114] br[114] wl[162] vdd gnd cell_6t
Xbit_r163_c114 bl[114] br[114] wl[163] vdd gnd cell_6t
Xbit_r164_c114 bl[114] br[114] wl[164] vdd gnd cell_6t
Xbit_r165_c114 bl[114] br[114] wl[165] vdd gnd cell_6t
Xbit_r166_c114 bl[114] br[114] wl[166] vdd gnd cell_6t
Xbit_r167_c114 bl[114] br[114] wl[167] vdd gnd cell_6t
Xbit_r168_c114 bl[114] br[114] wl[168] vdd gnd cell_6t
Xbit_r169_c114 bl[114] br[114] wl[169] vdd gnd cell_6t
Xbit_r170_c114 bl[114] br[114] wl[170] vdd gnd cell_6t
Xbit_r171_c114 bl[114] br[114] wl[171] vdd gnd cell_6t
Xbit_r172_c114 bl[114] br[114] wl[172] vdd gnd cell_6t
Xbit_r173_c114 bl[114] br[114] wl[173] vdd gnd cell_6t
Xbit_r174_c114 bl[114] br[114] wl[174] vdd gnd cell_6t
Xbit_r175_c114 bl[114] br[114] wl[175] vdd gnd cell_6t
Xbit_r176_c114 bl[114] br[114] wl[176] vdd gnd cell_6t
Xbit_r177_c114 bl[114] br[114] wl[177] vdd gnd cell_6t
Xbit_r178_c114 bl[114] br[114] wl[178] vdd gnd cell_6t
Xbit_r179_c114 bl[114] br[114] wl[179] vdd gnd cell_6t
Xbit_r180_c114 bl[114] br[114] wl[180] vdd gnd cell_6t
Xbit_r181_c114 bl[114] br[114] wl[181] vdd gnd cell_6t
Xbit_r182_c114 bl[114] br[114] wl[182] vdd gnd cell_6t
Xbit_r183_c114 bl[114] br[114] wl[183] vdd gnd cell_6t
Xbit_r184_c114 bl[114] br[114] wl[184] vdd gnd cell_6t
Xbit_r185_c114 bl[114] br[114] wl[185] vdd gnd cell_6t
Xbit_r186_c114 bl[114] br[114] wl[186] vdd gnd cell_6t
Xbit_r187_c114 bl[114] br[114] wl[187] vdd gnd cell_6t
Xbit_r188_c114 bl[114] br[114] wl[188] vdd gnd cell_6t
Xbit_r189_c114 bl[114] br[114] wl[189] vdd gnd cell_6t
Xbit_r190_c114 bl[114] br[114] wl[190] vdd gnd cell_6t
Xbit_r191_c114 bl[114] br[114] wl[191] vdd gnd cell_6t
Xbit_r192_c114 bl[114] br[114] wl[192] vdd gnd cell_6t
Xbit_r193_c114 bl[114] br[114] wl[193] vdd gnd cell_6t
Xbit_r194_c114 bl[114] br[114] wl[194] vdd gnd cell_6t
Xbit_r195_c114 bl[114] br[114] wl[195] vdd gnd cell_6t
Xbit_r196_c114 bl[114] br[114] wl[196] vdd gnd cell_6t
Xbit_r197_c114 bl[114] br[114] wl[197] vdd gnd cell_6t
Xbit_r198_c114 bl[114] br[114] wl[198] vdd gnd cell_6t
Xbit_r199_c114 bl[114] br[114] wl[199] vdd gnd cell_6t
Xbit_r200_c114 bl[114] br[114] wl[200] vdd gnd cell_6t
Xbit_r201_c114 bl[114] br[114] wl[201] vdd gnd cell_6t
Xbit_r202_c114 bl[114] br[114] wl[202] vdd gnd cell_6t
Xbit_r203_c114 bl[114] br[114] wl[203] vdd gnd cell_6t
Xbit_r204_c114 bl[114] br[114] wl[204] vdd gnd cell_6t
Xbit_r205_c114 bl[114] br[114] wl[205] vdd gnd cell_6t
Xbit_r206_c114 bl[114] br[114] wl[206] vdd gnd cell_6t
Xbit_r207_c114 bl[114] br[114] wl[207] vdd gnd cell_6t
Xbit_r208_c114 bl[114] br[114] wl[208] vdd gnd cell_6t
Xbit_r209_c114 bl[114] br[114] wl[209] vdd gnd cell_6t
Xbit_r210_c114 bl[114] br[114] wl[210] vdd gnd cell_6t
Xbit_r211_c114 bl[114] br[114] wl[211] vdd gnd cell_6t
Xbit_r212_c114 bl[114] br[114] wl[212] vdd gnd cell_6t
Xbit_r213_c114 bl[114] br[114] wl[213] vdd gnd cell_6t
Xbit_r214_c114 bl[114] br[114] wl[214] vdd gnd cell_6t
Xbit_r215_c114 bl[114] br[114] wl[215] vdd gnd cell_6t
Xbit_r216_c114 bl[114] br[114] wl[216] vdd gnd cell_6t
Xbit_r217_c114 bl[114] br[114] wl[217] vdd gnd cell_6t
Xbit_r218_c114 bl[114] br[114] wl[218] vdd gnd cell_6t
Xbit_r219_c114 bl[114] br[114] wl[219] vdd gnd cell_6t
Xbit_r220_c114 bl[114] br[114] wl[220] vdd gnd cell_6t
Xbit_r221_c114 bl[114] br[114] wl[221] vdd gnd cell_6t
Xbit_r222_c114 bl[114] br[114] wl[222] vdd gnd cell_6t
Xbit_r223_c114 bl[114] br[114] wl[223] vdd gnd cell_6t
Xbit_r224_c114 bl[114] br[114] wl[224] vdd gnd cell_6t
Xbit_r225_c114 bl[114] br[114] wl[225] vdd gnd cell_6t
Xbit_r226_c114 bl[114] br[114] wl[226] vdd gnd cell_6t
Xbit_r227_c114 bl[114] br[114] wl[227] vdd gnd cell_6t
Xbit_r228_c114 bl[114] br[114] wl[228] vdd gnd cell_6t
Xbit_r229_c114 bl[114] br[114] wl[229] vdd gnd cell_6t
Xbit_r230_c114 bl[114] br[114] wl[230] vdd gnd cell_6t
Xbit_r231_c114 bl[114] br[114] wl[231] vdd gnd cell_6t
Xbit_r232_c114 bl[114] br[114] wl[232] vdd gnd cell_6t
Xbit_r233_c114 bl[114] br[114] wl[233] vdd gnd cell_6t
Xbit_r234_c114 bl[114] br[114] wl[234] vdd gnd cell_6t
Xbit_r235_c114 bl[114] br[114] wl[235] vdd gnd cell_6t
Xbit_r236_c114 bl[114] br[114] wl[236] vdd gnd cell_6t
Xbit_r237_c114 bl[114] br[114] wl[237] vdd gnd cell_6t
Xbit_r238_c114 bl[114] br[114] wl[238] vdd gnd cell_6t
Xbit_r239_c114 bl[114] br[114] wl[239] vdd gnd cell_6t
Xbit_r240_c114 bl[114] br[114] wl[240] vdd gnd cell_6t
Xbit_r241_c114 bl[114] br[114] wl[241] vdd gnd cell_6t
Xbit_r242_c114 bl[114] br[114] wl[242] vdd gnd cell_6t
Xbit_r243_c114 bl[114] br[114] wl[243] vdd gnd cell_6t
Xbit_r244_c114 bl[114] br[114] wl[244] vdd gnd cell_6t
Xbit_r245_c114 bl[114] br[114] wl[245] vdd gnd cell_6t
Xbit_r246_c114 bl[114] br[114] wl[246] vdd gnd cell_6t
Xbit_r247_c114 bl[114] br[114] wl[247] vdd gnd cell_6t
Xbit_r248_c114 bl[114] br[114] wl[248] vdd gnd cell_6t
Xbit_r249_c114 bl[114] br[114] wl[249] vdd gnd cell_6t
Xbit_r250_c114 bl[114] br[114] wl[250] vdd gnd cell_6t
Xbit_r251_c114 bl[114] br[114] wl[251] vdd gnd cell_6t
Xbit_r252_c114 bl[114] br[114] wl[252] vdd gnd cell_6t
Xbit_r253_c114 bl[114] br[114] wl[253] vdd gnd cell_6t
Xbit_r254_c114 bl[114] br[114] wl[254] vdd gnd cell_6t
Xbit_r255_c114 bl[114] br[114] wl[255] vdd gnd cell_6t
Xbit_r0_c115 bl[115] br[115] wl[0] vdd gnd cell_6t
Xbit_r1_c115 bl[115] br[115] wl[1] vdd gnd cell_6t
Xbit_r2_c115 bl[115] br[115] wl[2] vdd gnd cell_6t
Xbit_r3_c115 bl[115] br[115] wl[3] vdd gnd cell_6t
Xbit_r4_c115 bl[115] br[115] wl[4] vdd gnd cell_6t
Xbit_r5_c115 bl[115] br[115] wl[5] vdd gnd cell_6t
Xbit_r6_c115 bl[115] br[115] wl[6] vdd gnd cell_6t
Xbit_r7_c115 bl[115] br[115] wl[7] vdd gnd cell_6t
Xbit_r8_c115 bl[115] br[115] wl[8] vdd gnd cell_6t
Xbit_r9_c115 bl[115] br[115] wl[9] vdd gnd cell_6t
Xbit_r10_c115 bl[115] br[115] wl[10] vdd gnd cell_6t
Xbit_r11_c115 bl[115] br[115] wl[11] vdd gnd cell_6t
Xbit_r12_c115 bl[115] br[115] wl[12] vdd gnd cell_6t
Xbit_r13_c115 bl[115] br[115] wl[13] vdd gnd cell_6t
Xbit_r14_c115 bl[115] br[115] wl[14] vdd gnd cell_6t
Xbit_r15_c115 bl[115] br[115] wl[15] vdd gnd cell_6t
Xbit_r16_c115 bl[115] br[115] wl[16] vdd gnd cell_6t
Xbit_r17_c115 bl[115] br[115] wl[17] vdd gnd cell_6t
Xbit_r18_c115 bl[115] br[115] wl[18] vdd gnd cell_6t
Xbit_r19_c115 bl[115] br[115] wl[19] vdd gnd cell_6t
Xbit_r20_c115 bl[115] br[115] wl[20] vdd gnd cell_6t
Xbit_r21_c115 bl[115] br[115] wl[21] vdd gnd cell_6t
Xbit_r22_c115 bl[115] br[115] wl[22] vdd gnd cell_6t
Xbit_r23_c115 bl[115] br[115] wl[23] vdd gnd cell_6t
Xbit_r24_c115 bl[115] br[115] wl[24] vdd gnd cell_6t
Xbit_r25_c115 bl[115] br[115] wl[25] vdd gnd cell_6t
Xbit_r26_c115 bl[115] br[115] wl[26] vdd gnd cell_6t
Xbit_r27_c115 bl[115] br[115] wl[27] vdd gnd cell_6t
Xbit_r28_c115 bl[115] br[115] wl[28] vdd gnd cell_6t
Xbit_r29_c115 bl[115] br[115] wl[29] vdd gnd cell_6t
Xbit_r30_c115 bl[115] br[115] wl[30] vdd gnd cell_6t
Xbit_r31_c115 bl[115] br[115] wl[31] vdd gnd cell_6t
Xbit_r32_c115 bl[115] br[115] wl[32] vdd gnd cell_6t
Xbit_r33_c115 bl[115] br[115] wl[33] vdd gnd cell_6t
Xbit_r34_c115 bl[115] br[115] wl[34] vdd gnd cell_6t
Xbit_r35_c115 bl[115] br[115] wl[35] vdd gnd cell_6t
Xbit_r36_c115 bl[115] br[115] wl[36] vdd gnd cell_6t
Xbit_r37_c115 bl[115] br[115] wl[37] vdd gnd cell_6t
Xbit_r38_c115 bl[115] br[115] wl[38] vdd gnd cell_6t
Xbit_r39_c115 bl[115] br[115] wl[39] vdd gnd cell_6t
Xbit_r40_c115 bl[115] br[115] wl[40] vdd gnd cell_6t
Xbit_r41_c115 bl[115] br[115] wl[41] vdd gnd cell_6t
Xbit_r42_c115 bl[115] br[115] wl[42] vdd gnd cell_6t
Xbit_r43_c115 bl[115] br[115] wl[43] vdd gnd cell_6t
Xbit_r44_c115 bl[115] br[115] wl[44] vdd gnd cell_6t
Xbit_r45_c115 bl[115] br[115] wl[45] vdd gnd cell_6t
Xbit_r46_c115 bl[115] br[115] wl[46] vdd gnd cell_6t
Xbit_r47_c115 bl[115] br[115] wl[47] vdd gnd cell_6t
Xbit_r48_c115 bl[115] br[115] wl[48] vdd gnd cell_6t
Xbit_r49_c115 bl[115] br[115] wl[49] vdd gnd cell_6t
Xbit_r50_c115 bl[115] br[115] wl[50] vdd gnd cell_6t
Xbit_r51_c115 bl[115] br[115] wl[51] vdd gnd cell_6t
Xbit_r52_c115 bl[115] br[115] wl[52] vdd gnd cell_6t
Xbit_r53_c115 bl[115] br[115] wl[53] vdd gnd cell_6t
Xbit_r54_c115 bl[115] br[115] wl[54] vdd gnd cell_6t
Xbit_r55_c115 bl[115] br[115] wl[55] vdd gnd cell_6t
Xbit_r56_c115 bl[115] br[115] wl[56] vdd gnd cell_6t
Xbit_r57_c115 bl[115] br[115] wl[57] vdd gnd cell_6t
Xbit_r58_c115 bl[115] br[115] wl[58] vdd gnd cell_6t
Xbit_r59_c115 bl[115] br[115] wl[59] vdd gnd cell_6t
Xbit_r60_c115 bl[115] br[115] wl[60] vdd gnd cell_6t
Xbit_r61_c115 bl[115] br[115] wl[61] vdd gnd cell_6t
Xbit_r62_c115 bl[115] br[115] wl[62] vdd gnd cell_6t
Xbit_r63_c115 bl[115] br[115] wl[63] vdd gnd cell_6t
Xbit_r64_c115 bl[115] br[115] wl[64] vdd gnd cell_6t
Xbit_r65_c115 bl[115] br[115] wl[65] vdd gnd cell_6t
Xbit_r66_c115 bl[115] br[115] wl[66] vdd gnd cell_6t
Xbit_r67_c115 bl[115] br[115] wl[67] vdd gnd cell_6t
Xbit_r68_c115 bl[115] br[115] wl[68] vdd gnd cell_6t
Xbit_r69_c115 bl[115] br[115] wl[69] vdd gnd cell_6t
Xbit_r70_c115 bl[115] br[115] wl[70] vdd gnd cell_6t
Xbit_r71_c115 bl[115] br[115] wl[71] vdd gnd cell_6t
Xbit_r72_c115 bl[115] br[115] wl[72] vdd gnd cell_6t
Xbit_r73_c115 bl[115] br[115] wl[73] vdd gnd cell_6t
Xbit_r74_c115 bl[115] br[115] wl[74] vdd gnd cell_6t
Xbit_r75_c115 bl[115] br[115] wl[75] vdd gnd cell_6t
Xbit_r76_c115 bl[115] br[115] wl[76] vdd gnd cell_6t
Xbit_r77_c115 bl[115] br[115] wl[77] vdd gnd cell_6t
Xbit_r78_c115 bl[115] br[115] wl[78] vdd gnd cell_6t
Xbit_r79_c115 bl[115] br[115] wl[79] vdd gnd cell_6t
Xbit_r80_c115 bl[115] br[115] wl[80] vdd gnd cell_6t
Xbit_r81_c115 bl[115] br[115] wl[81] vdd gnd cell_6t
Xbit_r82_c115 bl[115] br[115] wl[82] vdd gnd cell_6t
Xbit_r83_c115 bl[115] br[115] wl[83] vdd gnd cell_6t
Xbit_r84_c115 bl[115] br[115] wl[84] vdd gnd cell_6t
Xbit_r85_c115 bl[115] br[115] wl[85] vdd gnd cell_6t
Xbit_r86_c115 bl[115] br[115] wl[86] vdd gnd cell_6t
Xbit_r87_c115 bl[115] br[115] wl[87] vdd gnd cell_6t
Xbit_r88_c115 bl[115] br[115] wl[88] vdd gnd cell_6t
Xbit_r89_c115 bl[115] br[115] wl[89] vdd gnd cell_6t
Xbit_r90_c115 bl[115] br[115] wl[90] vdd gnd cell_6t
Xbit_r91_c115 bl[115] br[115] wl[91] vdd gnd cell_6t
Xbit_r92_c115 bl[115] br[115] wl[92] vdd gnd cell_6t
Xbit_r93_c115 bl[115] br[115] wl[93] vdd gnd cell_6t
Xbit_r94_c115 bl[115] br[115] wl[94] vdd gnd cell_6t
Xbit_r95_c115 bl[115] br[115] wl[95] vdd gnd cell_6t
Xbit_r96_c115 bl[115] br[115] wl[96] vdd gnd cell_6t
Xbit_r97_c115 bl[115] br[115] wl[97] vdd gnd cell_6t
Xbit_r98_c115 bl[115] br[115] wl[98] vdd gnd cell_6t
Xbit_r99_c115 bl[115] br[115] wl[99] vdd gnd cell_6t
Xbit_r100_c115 bl[115] br[115] wl[100] vdd gnd cell_6t
Xbit_r101_c115 bl[115] br[115] wl[101] vdd gnd cell_6t
Xbit_r102_c115 bl[115] br[115] wl[102] vdd gnd cell_6t
Xbit_r103_c115 bl[115] br[115] wl[103] vdd gnd cell_6t
Xbit_r104_c115 bl[115] br[115] wl[104] vdd gnd cell_6t
Xbit_r105_c115 bl[115] br[115] wl[105] vdd gnd cell_6t
Xbit_r106_c115 bl[115] br[115] wl[106] vdd gnd cell_6t
Xbit_r107_c115 bl[115] br[115] wl[107] vdd gnd cell_6t
Xbit_r108_c115 bl[115] br[115] wl[108] vdd gnd cell_6t
Xbit_r109_c115 bl[115] br[115] wl[109] vdd gnd cell_6t
Xbit_r110_c115 bl[115] br[115] wl[110] vdd gnd cell_6t
Xbit_r111_c115 bl[115] br[115] wl[111] vdd gnd cell_6t
Xbit_r112_c115 bl[115] br[115] wl[112] vdd gnd cell_6t
Xbit_r113_c115 bl[115] br[115] wl[113] vdd gnd cell_6t
Xbit_r114_c115 bl[115] br[115] wl[114] vdd gnd cell_6t
Xbit_r115_c115 bl[115] br[115] wl[115] vdd gnd cell_6t
Xbit_r116_c115 bl[115] br[115] wl[116] vdd gnd cell_6t
Xbit_r117_c115 bl[115] br[115] wl[117] vdd gnd cell_6t
Xbit_r118_c115 bl[115] br[115] wl[118] vdd gnd cell_6t
Xbit_r119_c115 bl[115] br[115] wl[119] vdd gnd cell_6t
Xbit_r120_c115 bl[115] br[115] wl[120] vdd gnd cell_6t
Xbit_r121_c115 bl[115] br[115] wl[121] vdd gnd cell_6t
Xbit_r122_c115 bl[115] br[115] wl[122] vdd gnd cell_6t
Xbit_r123_c115 bl[115] br[115] wl[123] vdd gnd cell_6t
Xbit_r124_c115 bl[115] br[115] wl[124] vdd gnd cell_6t
Xbit_r125_c115 bl[115] br[115] wl[125] vdd gnd cell_6t
Xbit_r126_c115 bl[115] br[115] wl[126] vdd gnd cell_6t
Xbit_r127_c115 bl[115] br[115] wl[127] vdd gnd cell_6t
Xbit_r128_c115 bl[115] br[115] wl[128] vdd gnd cell_6t
Xbit_r129_c115 bl[115] br[115] wl[129] vdd gnd cell_6t
Xbit_r130_c115 bl[115] br[115] wl[130] vdd gnd cell_6t
Xbit_r131_c115 bl[115] br[115] wl[131] vdd gnd cell_6t
Xbit_r132_c115 bl[115] br[115] wl[132] vdd gnd cell_6t
Xbit_r133_c115 bl[115] br[115] wl[133] vdd gnd cell_6t
Xbit_r134_c115 bl[115] br[115] wl[134] vdd gnd cell_6t
Xbit_r135_c115 bl[115] br[115] wl[135] vdd gnd cell_6t
Xbit_r136_c115 bl[115] br[115] wl[136] vdd gnd cell_6t
Xbit_r137_c115 bl[115] br[115] wl[137] vdd gnd cell_6t
Xbit_r138_c115 bl[115] br[115] wl[138] vdd gnd cell_6t
Xbit_r139_c115 bl[115] br[115] wl[139] vdd gnd cell_6t
Xbit_r140_c115 bl[115] br[115] wl[140] vdd gnd cell_6t
Xbit_r141_c115 bl[115] br[115] wl[141] vdd gnd cell_6t
Xbit_r142_c115 bl[115] br[115] wl[142] vdd gnd cell_6t
Xbit_r143_c115 bl[115] br[115] wl[143] vdd gnd cell_6t
Xbit_r144_c115 bl[115] br[115] wl[144] vdd gnd cell_6t
Xbit_r145_c115 bl[115] br[115] wl[145] vdd gnd cell_6t
Xbit_r146_c115 bl[115] br[115] wl[146] vdd gnd cell_6t
Xbit_r147_c115 bl[115] br[115] wl[147] vdd gnd cell_6t
Xbit_r148_c115 bl[115] br[115] wl[148] vdd gnd cell_6t
Xbit_r149_c115 bl[115] br[115] wl[149] vdd gnd cell_6t
Xbit_r150_c115 bl[115] br[115] wl[150] vdd gnd cell_6t
Xbit_r151_c115 bl[115] br[115] wl[151] vdd gnd cell_6t
Xbit_r152_c115 bl[115] br[115] wl[152] vdd gnd cell_6t
Xbit_r153_c115 bl[115] br[115] wl[153] vdd gnd cell_6t
Xbit_r154_c115 bl[115] br[115] wl[154] vdd gnd cell_6t
Xbit_r155_c115 bl[115] br[115] wl[155] vdd gnd cell_6t
Xbit_r156_c115 bl[115] br[115] wl[156] vdd gnd cell_6t
Xbit_r157_c115 bl[115] br[115] wl[157] vdd gnd cell_6t
Xbit_r158_c115 bl[115] br[115] wl[158] vdd gnd cell_6t
Xbit_r159_c115 bl[115] br[115] wl[159] vdd gnd cell_6t
Xbit_r160_c115 bl[115] br[115] wl[160] vdd gnd cell_6t
Xbit_r161_c115 bl[115] br[115] wl[161] vdd gnd cell_6t
Xbit_r162_c115 bl[115] br[115] wl[162] vdd gnd cell_6t
Xbit_r163_c115 bl[115] br[115] wl[163] vdd gnd cell_6t
Xbit_r164_c115 bl[115] br[115] wl[164] vdd gnd cell_6t
Xbit_r165_c115 bl[115] br[115] wl[165] vdd gnd cell_6t
Xbit_r166_c115 bl[115] br[115] wl[166] vdd gnd cell_6t
Xbit_r167_c115 bl[115] br[115] wl[167] vdd gnd cell_6t
Xbit_r168_c115 bl[115] br[115] wl[168] vdd gnd cell_6t
Xbit_r169_c115 bl[115] br[115] wl[169] vdd gnd cell_6t
Xbit_r170_c115 bl[115] br[115] wl[170] vdd gnd cell_6t
Xbit_r171_c115 bl[115] br[115] wl[171] vdd gnd cell_6t
Xbit_r172_c115 bl[115] br[115] wl[172] vdd gnd cell_6t
Xbit_r173_c115 bl[115] br[115] wl[173] vdd gnd cell_6t
Xbit_r174_c115 bl[115] br[115] wl[174] vdd gnd cell_6t
Xbit_r175_c115 bl[115] br[115] wl[175] vdd gnd cell_6t
Xbit_r176_c115 bl[115] br[115] wl[176] vdd gnd cell_6t
Xbit_r177_c115 bl[115] br[115] wl[177] vdd gnd cell_6t
Xbit_r178_c115 bl[115] br[115] wl[178] vdd gnd cell_6t
Xbit_r179_c115 bl[115] br[115] wl[179] vdd gnd cell_6t
Xbit_r180_c115 bl[115] br[115] wl[180] vdd gnd cell_6t
Xbit_r181_c115 bl[115] br[115] wl[181] vdd gnd cell_6t
Xbit_r182_c115 bl[115] br[115] wl[182] vdd gnd cell_6t
Xbit_r183_c115 bl[115] br[115] wl[183] vdd gnd cell_6t
Xbit_r184_c115 bl[115] br[115] wl[184] vdd gnd cell_6t
Xbit_r185_c115 bl[115] br[115] wl[185] vdd gnd cell_6t
Xbit_r186_c115 bl[115] br[115] wl[186] vdd gnd cell_6t
Xbit_r187_c115 bl[115] br[115] wl[187] vdd gnd cell_6t
Xbit_r188_c115 bl[115] br[115] wl[188] vdd gnd cell_6t
Xbit_r189_c115 bl[115] br[115] wl[189] vdd gnd cell_6t
Xbit_r190_c115 bl[115] br[115] wl[190] vdd gnd cell_6t
Xbit_r191_c115 bl[115] br[115] wl[191] vdd gnd cell_6t
Xbit_r192_c115 bl[115] br[115] wl[192] vdd gnd cell_6t
Xbit_r193_c115 bl[115] br[115] wl[193] vdd gnd cell_6t
Xbit_r194_c115 bl[115] br[115] wl[194] vdd gnd cell_6t
Xbit_r195_c115 bl[115] br[115] wl[195] vdd gnd cell_6t
Xbit_r196_c115 bl[115] br[115] wl[196] vdd gnd cell_6t
Xbit_r197_c115 bl[115] br[115] wl[197] vdd gnd cell_6t
Xbit_r198_c115 bl[115] br[115] wl[198] vdd gnd cell_6t
Xbit_r199_c115 bl[115] br[115] wl[199] vdd gnd cell_6t
Xbit_r200_c115 bl[115] br[115] wl[200] vdd gnd cell_6t
Xbit_r201_c115 bl[115] br[115] wl[201] vdd gnd cell_6t
Xbit_r202_c115 bl[115] br[115] wl[202] vdd gnd cell_6t
Xbit_r203_c115 bl[115] br[115] wl[203] vdd gnd cell_6t
Xbit_r204_c115 bl[115] br[115] wl[204] vdd gnd cell_6t
Xbit_r205_c115 bl[115] br[115] wl[205] vdd gnd cell_6t
Xbit_r206_c115 bl[115] br[115] wl[206] vdd gnd cell_6t
Xbit_r207_c115 bl[115] br[115] wl[207] vdd gnd cell_6t
Xbit_r208_c115 bl[115] br[115] wl[208] vdd gnd cell_6t
Xbit_r209_c115 bl[115] br[115] wl[209] vdd gnd cell_6t
Xbit_r210_c115 bl[115] br[115] wl[210] vdd gnd cell_6t
Xbit_r211_c115 bl[115] br[115] wl[211] vdd gnd cell_6t
Xbit_r212_c115 bl[115] br[115] wl[212] vdd gnd cell_6t
Xbit_r213_c115 bl[115] br[115] wl[213] vdd gnd cell_6t
Xbit_r214_c115 bl[115] br[115] wl[214] vdd gnd cell_6t
Xbit_r215_c115 bl[115] br[115] wl[215] vdd gnd cell_6t
Xbit_r216_c115 bl[115] br[115] wl[216] vdd gnd cell_6t
Xbit_r217_c115 bl[115] br[115] wl[217] vdd gnd cell_6t
Xbit_r218_c115 bl[115] br[115] wl[218] vdd gnd cell_6t
Xbit_r219_c115 bl[115] br[115] wl[219] vdd gnd cell_6t
Xbit_r220_c115 bl[115] br[115] wl[220] vdd gnd cell_6t
Xbit_r221_c115 bl[115] br[115] wl[221] vdd gnd cell_6t
Xbit_r222_c115 bl[115] br[115] wl[222] vdd gnd cell_6t
Xbit_r223_c115 bl[115] br[115] wl[223] vdd gnd cell_6t
Xbit_r224_c115 bl[115] br[115] wl[224] vdd gnd cell_6t
Xbit_r225_c115 bl[115] br[115] wl[225] vdd gnd cell_6t
Xbit_r226_c115 bl[115] br[115] wl[226] vdd gnd cell_6t
Xbit_r227_c115 bl[115] br[115] wl[227] vdd gnd cell_6t
Xbit_r228_c115 bl[115] br[115] wl[228] vdd gnd cell_6t
Xbit_r229_c115 bl[115] br[115] wl[229] vdd gnd cell_6t
Xbit_r230_c115 bl[115] br[115] wl[230] vdd gnd cell_6t
Xbit_r231_c115 bl[115] br[115] wl[231] vdd gnd cell_6t
Xbit_r232_c115 bl[115] br[115] wl[232] vdd gnd cell_6t
Xbit_r233_c115 bl[115] br[115] wl[233] vdd gnd cell_6t
Xbit_r234_c115 bl[115] br[115] wl[234] vdd gnd cell_6t
Xbit_r235_c115 bl[115] br[115] wl[235] vdd gnd cell_6t
Xbit_r236_c115 bl[115] br[115] wl[236] vdd gnd cell_6t
Xbit_r237_c115 bl[115] br[115] wl[237] vdd gnd cell_6t
Xbit_r238_c115 bl[115] br[115] wl[238] vdd gnd cell_6t
Xbit_r239_c115 bl[115] br[115] wl[239] vdd gnd cell_6t
Xbit_r240_c115 bl[115] br[115] wl[240] vdd gnd cell_6t
Xbit_r241_c115 bl[115] br[115] wl[241] vdd gnd cell_6t
Xbit_r242_c115 bl[115] br[115] wl[242] vdd gnd cell_6t
Xbit_r243_c115 bl[115] br[115] wl[243] vdd gnd cell_6t
Xbit_r244_c115 bl[115] br[115] wl[244] vdd gnd cell_6t
Xbit_r245_c115 bl[115] br[115] wl[245] vdd gnd cell_6t
Xbit_r246_c115 bl[115] br[115] wl[246] vdd gnd cell_6t
Xbit_r247_c115 bl[115] br[115] wl[247] vdd gnd cell_6t
Xbit_r248_c115 bl[115] br[115] wl[248] vdd gnd cell_6t
Xbit_r249_c115 bl[115] br[115] wl[249] vdd gnd cell_6t
Xbit_r250_c115 bl[115] br[115] wl[250] vdd gnd cell_6t
Xbit_r251_c115 bl[115] br[115] wl[251] vdd gnd cell_6t
Xbit_r252_c115 bl[115] br[115] wl[252] vdd gnd cell_6t
Xbit_r253_c115 bl[115] br[115] wl[253] vdd gnd cell_6t
Xbit_r254_c115 bl[115] br[115] wl[254] vdd gnd cell_6t
Xbit_r255_c115 bl[115] br[115] wl[255] vdd gnd cell_6t
Xbit_r0_c116 bl[116] br[116] wl[0] vdd gnd cell_6t
Xbit_r1_c116 bl[116] br[116] wl[1] vdd gnd cell_6t
Xbit_r2_c116 bl[116] br[116] wl[2] vdd gnd cell_6t
Xbit_r3_c116 bl[116] br[116] wl[3] vdd gnd cell_6t
Xbit_r4_c116 bl[116] br[116] wl[4] vdd gnd cell_6t
Xbit_r5_c116 bl[116] br[116] wl[5] vdd gnd cell_6t
Xbit_r6_c116 bl[116] br[116] wl[6] vdd gnd cell_6t
Xbit_r7_c116 bl[116] br[116] wl[7] vdd gnd cell_6t
Xbit_r8_c116 bl[116] br[116] wl[8] vdd gnd cell_6t
Xbit_r9_c116 bl[116] br[116] wl[9] vdd gnd cell_6t
Xbit_r10_c116 bl[116] br[116] wl[10] vdd gnd cell_6t
Xbit_r11_c116 bl[116] br[116] wl[11] vdd gnd cell_6t
Xbit_r12_c116 bl[116] br[116] wl[12] vdd gnd cell_6t
Xbit_r13_c116 bl[116] br[116] wl[13] vdd gnd cell_6t
Xbit_r14_c116 bl[116] br[116] wl[14] vdd gnd cell_6t
Xbit_r15_c116 bl[116] br[116] wl[15] vdd gnd cell_6t
Xbit_r16_c116 bl[116] br[116] wl[16] vdd gnd cell_6t
Xbit_r17_c116 bl[116] br[116] wl[17] vdd gnd cell_6t
Xbit_r18_c116 bl[116] br[116] wl[18] vdd gnd cell_6t
Xbit_r19_c116 bl[116] br[116] wl[19] vdd gnd cell_6t
Xbit_r20_c116 bl[116] br[116] wl[20] vdd gnd cell_6t
Xbit_r21_c116 bl[116] br[116] wl[21] vdd gnd cell_6t
Xbit_r22_c116 bl[116] br[116] wl[22] vdd gnd cell_6t
Xbit_r23_c116 bl[116] br[116] wl[23] vdd gnd cell_6t
Xbit_r24_c116 bl[116] br[116] wl[24] vdd gnd cell_6t
Xbit_r25_c116 bl[116] br[116] wl[25] vdd gnd cell_6t
Xbit_r26_c116 bl[116] br[116] wl[26] vdd gnd cell_6t
Xbit_r27_c116 bl[116] br[116] wl[27] vdd gnd cell_6t
Xbit_r28_c116 bl[116] br[116] wl[28] vdd gnd cell_6t
Xbit_r29_c116 bl[116] br[116] wl[29] vdd gnd cell_6t
Xbit_r30_c116 bl[116] br[116] wl[30] vdd gnd cell_6t
Xbit_r31_c116 bl[116] br[116] wl[31] vdd gnd cell_6t
Xbit_r32_c116 bl[116] br[116] wl[32] vdd gnd cell_6t
Xbit_r33_c116 bl[116] br[116] wl[33] vdd gnd cell_6t
Xbit_r34_c116 bl[116] br[116] wl[34] vdd gnd cell_6t
Xbit_r35_c116 bl[116] br[116] wl[35] vdd gnd cell_6t
Xbit_r36_c116 bl[116] br[116] wl[36] vdd gnd cell_6t
Xbit_r37_c116 bl[116] br[116] wl[37] vdd gnd cell_6t
Xbit_r38_c116 bl[116] br[116] wl[38] vdd gnd cell_6t
Xbit_r39_c116 bl[116] br[116] wl[39] vdd gnd cell_6t
Xbit_r40_c116 bl[116] br[116] wl[40] vdd gnd cell_6t
Xbit_r41_c116 bl[116] br[116] wl[41] vdd gnd cell_6t
Xbit_r42_c116 bl[116] br[116] wl[42] vdd gnd cell_6t
Xbit_r43_c116 bl[116] br[116] wl[43] vdd gnd cell_6t
Xbit_r44_c116 bl[116] br[116] wl[44] vdd gnd cell_6t
Xbit_r45_c116 bl[116] br[116] wl[45] vdd gnd cell_6t
Xbit_r46_c116 bl[116] br[116] wl[46] vdd gnd cell_6t
Xbit_r47_c116 bl[116] br[116] wl[47] vdd gnd cell_6t
Xbit_r48_c116 bl[116] br[116] wl[48] vdd gnd cell_6t
Xbit_r49_c116 bl[116] br[116] wl[49] vdd gnd cell_6t
Xbit_r50_c116 bl[116] br[116] wl[50] vdd gnd cell_6t
Xbit_r51_c116 bl[116] br[116] wl[51] vdd gnd cell_6t
Xbit_r52_c116 bl[116] br[116] wl[52] vdd gnd cell_6t
Xbit_r53_c116 bl[116] br[116] wl[53] vdd gnd cell_6t
Xbit_r54_c116 bl[116] br[116] wl[54] vdd gnd cell_6t
Xbit_r55_c116 bl[116] br[116] wl[55] vdd gnd cell_6t
Xbit_r56_c116 bl[116] br[116] wl[56] vdd gnd cell_6t
Xbit_r57_c116 bl[116] br[116] wl[57] vdd gnd cell_6t
Xbit_r58_c116 bl[116] br[116] wl[58] vdd gnd cell_6t
Xbit_r59_c116 bl[116] br[116] wl[59] vdd gnd cell_6t
Xbit_r60_c116 bl[116] br[116] wl[60] vdd gnd cell_6t
Xbit_r61_c116 bl[116] br[116] wl[61] vdd gnd cell_6t
Xbit_r62_c116 bl[116] br[116] wl[62] vdd gnd cell_6t
Xbit_r63_c116 bl[116] br[116] wl[63] vdd gnd cell_6t
Xbit_r64_c116 bl[116] br[116] wl[64] vdd gnd cell_6t
Xbit_r65_c116 bl[116] br[116] wl[65] vdd gnd cell_6t
Xbit_r66_c116 bl[116] br[116] wl[66] vdd gnd cell_6t
Xbit_r67_c116 bl[116] br[116] wl[67] vdd gnd cell_6t
Xbit_r68_c116 bl[116] br[116] wl[68] vdd gnd cell_6t
Xbit_r69_c116 bl[116] br[116] wl[69] vdd gnd cell_6t
Xbit_r70_c116 bl[116] br[116] wl[70] vdd gnd cell_6t
Xbit_r71_c116 bl[116] br[116] wl[71] vdd gnd cell_6t
Xbit_r72_c116 bl[116] br[116] wl[72] vdd gnd cell_6t
Xbit_r73_c116 bl[116] br[116] wl[73] vdd gnd cell_6t
Xbit_r74_c116 bl[116] br[116] wl[74] vdd gnd cell_6t
Xbit_r75_c116 bl[116] br[116] wl[75] vdd gnd cell_6t
Xbit_r76_c116 bl[116] br[116] wl[76] vdd gnd cell_6t
Xbit_r77_c116 bl[116] br[116] wl[77] vdd gnd cell_6t
Xbit_r78_c116 bl[116] br[116] wl[78] vdd gnd cell_6t
Xbit_r79_c116 bl[116] br[116] wl[79] vdd gnd cell_6t
Xbit_r80_c116 bl[116] br[116] wl[80] vdd gnd cell_6t
Xbit_r81_c116 bl[116] br[116] wl[81] vdd gnd cell_6t
Xbit_r82_c116 bl[116] br[116] wl[82] vdd gnd cell_6t
Xbit_r83_c116 bl[116] br[116] wl[83] vdd gnd cell_6t
Xbit_r84_c116 bl[116] br[116] wl[84] vdd gnd cell_6t
Xbit_r85_c116 bl[116] br[116] wl[85] vdd gnd cell_6t
Xbit_r86_c116 bl[116] br[116] wl[86] vdd gnd cell_6t
Xbit_r87_c116 bl[116] br[116] wl[87] vdd gnd cell_6t
Xbit_r88_c116 bl[116] br[116] wl[88] vdd gnd cell_6t
Xbit_r89_c116 bl[116] br[116] wl[89] vdd gnd cell_6t
Xbit_r90_c116 bl[116] br[116] wl[90] vdd gnd cell_6t
Xbit_r91_c116 bl[116] br[116] wl[91] vdd gnd cell_6t
Xbit_r92_c116 bl[116] br[116] wl[92] vdd gnd cell_6t
Xbit_r93_c116 bl[116] br[116] wl[93] vdd gnd cell_6t
Xbit_r94_c116 bl[116] br[116] wl[94] vdd gnd cell_6t
Xbit_r95_c116 bl[116] br[116] wl[95] vdd gnd cell_6t
Xbit_r96_c116 bl[116] br[116] wl[96] vdd gnd cell_6t
Xbit_r97_c116 bl[116] br[116] wl[97] vdd gnd cell_6t
Xbit_r98_c116 bl[116] br[116] wl[98] vdd gnd cell_6t
Xbit_r99_c116 bl[116] br[116] wl[99] vdd gnd cell_6t
Xbit_r100_c116 bl[116] br[116] wl[100] vdd gnd cell_6t
Xbit_r101_c116 bl[116] br[116] wl[101] vdd gnd cell_6t
Xbit_r102_c116 bl[116] br[116] wl[102] vdd gnd cell_6t
Xbit_r103_c116 bl[116] br[116] wl[103] vdd gnd cell_6t
Xbit_r104_c116 bl[116] br[116] wl[104] vdd gnd cell_6t
Xbit_r105_c116 bl[116] br[116] wl[105] vdd gnd cell_6t
Xbit_r106_c116 bl[116] br[116] wl[106] vdd gnd cell_6t
Xbit_r107_c116 bl[116] br[116] wl[107] vdd gnd cell_6t
Xbit_r108_c116 bl[116] br[116] wl[108] vdd gnd cell_6t
Xbit_r109_c116 bl[116] br[116] wl[109] vdd gnd cell_6t
Xbit_r110_c116 bl[116] br[116] wl[110] vdd gnd cell_6t
Xbit_r111_c116 bl[116] br[116] wl[111] vdd gnd cell_6t
Xbit_r112_c116 bl[116] br[116] wl[112] vdd gnd cell_6t
Xbit_r113_c116 bl[116] br[116] wl[113] vdd gnd cell_6t
Xbit_r114_c116 bl[116] br[116] wl[114] vdd gnd cell_6t
Xbit_r115_c116 bl[116] br[116] wl[115] vdd gnd cell_6t
Xbit_r116_c116 bl[116] br[116] wl[116] vdd gnd cell_6t
Xbit_r117_c116 bl[116] br[116] wl[117] vdd gnd cell_6t
Xbit_r118_c116 bl[116] br[116] wl[118] vdd gnd cell_6t
Xbit_r119_c116 bl[116] br[116] wl[119] vdd gnd cell_6t
Xbit_r120_c116 bl[116] br[116] wl[120] vdd gnd cell_6t
Xbit_r121_c116 bl[116] br[116] wl[121] vdd gnd cell_6t
Xbit_r122_c116 bl[116] br[116] wl[122] vdd gnd cell_6t
Xbit_r123_c116 bl[116] br[116] wl[123] vdd gnd cell_6t
Xbit_r124_c116 bl[116] br[116] wl[124] vdd gnd cell_6t
Xbit_r125_c116 bl[116] br[116] wl[125] vdd gnd cell_6t
Xbit_r126_c116 bl[116] br[116] wl[126] vdd gnd cell_6t
Xbit_r127_c116 bl[116] br[116] wl[127] vdd gnd cell_6t
Xbit_r128_c116 bl[116] br[116] wl[128] vdd gnd cell_6t
Xbit_r129_c116 bl[116] br[116] wl[129] vdd gnd cell_6t
Xbit_r130_c116 bl[116] br[116] wl[130] vdd gnd cell_6t
Xbit_r131_c116 bl[116] br[116] wl[131] vdd gnd cell_6t
Xbit_r132_c116 bl[116] br[116] wl[132] vdd gnd cell_6t
Xbit_r133_c116 bl[116] br[116] wl[133] vdd gnd cell_6t
Xbit_r134_c116 bl[116] br[116] wl[134] vdd gnd cell_6t
Xbit_r135_c116 bl[116] br[116] wl[135] vdd gnd cell_6t
Xbit_r136_c116 bl[116] br[116] wl[136] vdd gnd cell_6t
Xbit_r137_c116 bl[116] br[116] wl[137] vdd gnd cell_6t
Xbit_r138_c116 bl[116] br[116] wl[138] vdd gnd cell_6t
Xbit_r139_c116 bl[116] br[116] wl[139] vdd gnd cell_6t
Xbit_r140_c116 bl[116] br[116] wl[140] vdd gnd cell_6t
Xbit_r141_c116 bl[116] br[116] wl[141] vdd gnd cell_6t
Xbit_r142_c116 bl[116] br[116] wl[142] vdd gnd cell_6t
Xbit_r143_c116 bl[116] br[116] wl[143] vdd gnd cell_6t
Xbit_r144_c116 bl[116] br[116] wl[144] vdd gnd cell_6t
Xbit_r145_c116 bl[116] br[116] wl[145] vdd gnd cell_6t
Xbit_r146_c116 bl[116] br[116] wl[146] vdd gnd cell_6t
Xbit_r147_c116 bl[116] br[116] wl[147] vdd gnd cell_6t
Xbit_r148_c116 bl[116] br[116] wl[148] vdd gnd cell_6t
Xbit_r149_c116 bl[116] br[116] wl[149] vdd gnd cell_6t
Xbit_r150_c116 bl[116] br[116] wl[150] vdd gnd cell_6t
Xbit_r151_c116 bl[116] br[116] wl[151] vdd gnd cell_6t
Xbit_r152_c116 bl[116] br[116] wl[152] vdd gnd cell_6t
Xbit_r153_c116 bl[116] br[116] wl[153] vdd gnd cell_6t
Xbit_r154_c116 bl[116] br[116] wl[154] vdd gnd cell_6t
Xbit_r155_c116 bl[116] br[116] wl[155] vdd gnd cell_6t
Xbit_r156_c116 bl[116] br[116] wl[156] vdd gnd cell_6t
Xbit_r157_c116 bl[116] br[116] wl[157] vdd gnd cell_6t
Xbit_r158_c116 bl[116] br[116] wl[158] vdd gnd cell_6t
Xbit_r159_c116 bl[116] br[116] wl[159] vdd gnd cell_6t
Xbit_r160_c116 bl[116] br[116] wl[160] vdd gnd cell_6t
Xbit_r161_c116 bl[116] br[116] wl[161] vdd gnd cell_6t
Xbit_r162_c116 bl[116] br[116] wl[162] vdd gnd cell_6t
Xbit_r163_c116 bl[116] br[116] wl[163] vdd gnd cell_6t
Xbit_r164_c116 bl[116] br[116] wl[164] vdd gnd cell_6t
Xbit_r165_c116 bl[116] br[116] wl[165] vdd gnd cell_6t
Xbit_r166_c116 bl[116] br[116] wl[166] vdd gnd cell_6t
Xbit_r167_c116 bl[116] br[116] wl[167] vdd gnd cell_6t
Xbit_r168_c116 bl[116] br[116] wl[168] vdd gnd cell_6t
Xbit_r169_c116 bl[116] br[116] wl[169] vdd gnd cell_6t
Xbit_r170_c116 bl[116] br[116] wl[170] vdd gnd cell_6t
Xbit_r171_c116 bl[116] br[116] wl[171] vdd gnd cell_6t
Xbit_r172_c116 bl[116] br[116] wl[172] vdd gnd cell_6t
Xbit_r173_c116 bl[116] br[116] wl[173] vdd gnd cell_6t
Xbit_r174_c116 bl[116] br[116] wl[174] vdd gnd cell_6t
Xbit_r175_c116 bl[116] br[116] wl[175] vdd gnd cell_6t
Xbit_r176_c116 bl[116] br[116] wl[176] vdd gnd cell_6t
Xbit_r177_c116 bl[116] br[116] wl[177] vdd gnd cell_6t
Xbit_r178_c116 bl[116] br[116] wl[178] vdd gnd cell_6t
Xbit_r179_c116 bl[116] br[116] wl[179] vdd gnd cell_6t
Xbit_r180_c116 bl[116] br[116] wl[180] vdd gnd cell_6t
Xbit_r181_c116 bl[116] br[116] wl[181] vdd gnd cell_6t
Xbit_r182_c116 bl[116] br[116] wl[182] vdd gnd cell_6t
Xbit_r183_c116 bl[116] br[116] wl[183] vdd gnd cell_6t
Xbit_r184_c116 bl[116] br[116] wl[184] vdd gnd cell_6t
Xbit_r185_c116 bl[116] br[116] wl[185] vdd gnd cell_6t
Xbit_r186_c116 bl[116] br[116] wl[186] vdd gnd cell_6t
Xbit_r187_c116 bl[116] br[116] wl[187] vdd gnd cell_6t
Xbit_r188_c116 bl[116] br[116] wl[188] vdd gnd cell_6t
Xbit_r189_c116 bl[116] br[116] wl[189] vdd gnd cell_6t
Xbit_r190_c116 bl[116] br[116] wl[190] vdd gnd cell_6t
Xbit_r191_c116 bl[116] br[116] wl[191] vdd gnd cell_6t
Xbit_r192_c116 bl[116] br[116] wl[192] vdd gnd cell_6t
Xbit_r193_c116 bl[116] br[116] wl[193] vdd gnd cell_6t
Xbit_r194_c116 bl[116] br[116] wl[194] vdd gnd cell_6t
Xbit_r195_c116 bl[116] br[116] wl[195] vdd gnd cell_6t
Xbit_r196_c116 bl[116] br[116] wl[196] vdd gnd cell_6t
Xbit_r197_c116 bl[116] br[116] wl[197] vdd gnd cell_6t
Xbit_r198_c116 bl[116] br[116] wl[198] vdd gnd cell_6t
Xbit_r199_c116 bl[116] br[116] wl[199] vdd gnd cell_6t
Xbit_r200_c116 bl[116] br[116] wl[200] vdd gnd cell_6t
Xbit_r201_c116 bl[116] br[116] wl[201] vdd gnd cell_6t
Xbit_r202_c116 bl[116] br[116] wl[202] vdd gnd cell_6t
Xbit_r203_c116 bl[116] br[116] wl[203] vdd gnd cell_6t
Xbit_r204_c116 bl[116] br[116] wl[204] vdd gnd cell_6t
Xbit_r205_c116 bl[116] br[116] wl[205] vdd gnd cell_6t
Xbit_r206_c116 bl[116] br[116] wl[206] vdd gnd cell_6t
Xbit_r207_c116 bl[116] br[116] wl[207] vdd gnd cell_6t
Xbit_r208_c116 bl[116] br[116] wl[208] vdd gnd cell_6t
Xbit_r209_c116 bl[116] br[116] wl[209] vdd gnd cell_6t
Xbit_r210_c116 bl[116] br[116] wl[210] vdd gnd cell_6t
Xbit_r211_c116 bl[116] br[116] wl[211] vdd gnd cell_6t
Xbit_r212_c116 bl[116] br[116] wl[212] vdd gnd cell_6t
Xbit_r213_c116 bl[116] br[116] wl[213] vdd gnd cell_6t
Xbit_r214_c116 bl[116] br[116] wl[214] vdd gnd cell_6t
Xbit_r215_c116 bl[116] br[116] wl[215] vdd gnd cell_6t
Xbit_r216_c116 bl[116] br[116] wl[216] vdd gnd cell_6t
Xbit_r217_c116 bl[116] br[116] wl[217] vdd gnd cell_6t
Xbit_r218_c116 bl[116] br[116] wl[218] vdd gnd cell_6t
Xbit_r219_c116 bl[116] br[116] wl[219] vdd gnd cell_6t
Xbit_r220_c116 bl[116] br[116] wl[220] vdd gnd cell_6t
Xbit_r221_c116 bl[116] br[116] wl[221] vdd gnd cell_6t
Xbit_r222_c116 bl[116] br[116] wl[222] vdd gnd cell_6t
Xbit_r223_c116 bl[116] br[116] wl[223] vdd gnd cell_6t
Xbit_r224_c116 bl[116] br[116] wl[224] vdd gnd cell_6t
Xbit_r225_c116 bl[116] br[116] wl[225] vdd gnd cell_6t
Xbit_r226_c116 bl[116] br[116] wl[226] vdd gnd cell_6t
Xbit_r227_c116 bl[116] br[116] wl[227] vdd gnd cell_6t
Xbit_r228_c116 bl[116] br[116] wl[228] vdd gnd cell_6t
Xbit_r229_c116 bl[116] br[116] wl[229] vdd gnd cell_6t
Xbit_r230_c116 bl[116] br[116] wl[230] vdd gnd cell_6t
Xbit_r231_c116 bl[116] br[116] wl[231] vdd gnd cell_6t
Xbit_r232_c116 bl[116] br[116] wl[232] vdd gnd cell_6t
Xbit_r233_c116 bl[116] br[116] wl[233] vdd gnd cell_6t
Xbit_r234_c116 bl[116] br[116] wl[234] vdd gnd cell_6t
Xbit_r235_c116 bl[116] br[116] wl[235] vdd gnd cell_6t
Xbit_r236_c116 bl[116] br[116] wl[236] vdd gnd cell_6t
Xbit_r237_c116 bl[116] br[116] wl[237] vdd gnd cell_6t
Xbit_r238_c116 bl[116] br[116] wl[238] vdd gnd cell_6t
Xbit_r239_c116 bl[116] br[116] wl[239] vdd gnd cell_6t
Xbit_r240_c116 bl[116] br[116] wl[240] vdd gnd cell_6t
Xbit_r241_c116 bl[116] br[116] wl[241] vdd gnd cell_6t
Xbit_r242_c116 bl[116] br[116] wl[242] vdd gnd cell_6t
Xbit_r243_c116 bl[116] br[116] wl[243] vdd gnd cell_6t
Xbit_r244_c116 bl[116] br[116] wl[244] vdd gnd cell_6t
Xbit_r245_c116 bl[116] br[116] wl[245] vdd gnd cell_6t
Xbit_r246_c116 bl[116] br[116] wl[246] vdd gnd cell_6t
Xbit_r247_c116 bl[116] br[116] wl[247] vdd gnd cell_6t
Xbit_r248_c116 bl[116] br[116] wl[248] vdd gnd cell_6t
Xbit_r249_c116 bl[116] br[116] wl[249] vdd gnd cell_6t
Xbit_r250_c116 bl[116] br[116] wl[250] vdd gnd cell_6t
Xbit_r251_c116 bl[116] br[116] wl[251] vdd gnd cell_6t
Xbit_r252_c116 bl[116] br[116] wl[252] vdd gnd cell_6t
Xbit_r253_c116 bl[116] br[116] wl[253] vdd gnd cell_6t
Xbit_r254_c116 bl[116] br[116] wl[254] vdd gnd cell_6t
Xbit_r255_c116 bl[116] br[116] wl[255] vdd gnd cell_6t
Xbit_r0_c117 bl[117] br[117] wl[0] vdd gnd cell_6t
Xbit_r1_c117 bl[117] br[117] wl[1] vdd gnd cell_6t
Xbit_r2_c117 bl[117] br[117] wl[2] vdd gnd cell_6t
Xbit_r3_c117 bl[117] br[117] wl[3] vdd gnd cell_6t
Xbit_r4_c117 bl[117] br[117] wl[4] vdd gnd cell_6t
Xbit_r5_c117 bl[117] br[117] wl[5] vdd gnd cell_6t
Xbit_r6_c117 bl[117] br[117] wl[6] vdd gnd cell_6t
Xbit_r7_c117 bl[117] br[117] wl[7] vdd gnd cell_6t
Xbit_r8_c117 bl[117] br[117] wl[8] vdd gnd cell_6t
Xbit_r9_c117 bl[117] br[117] wl[9] vdd gnd cell_6t
Xbit_r10_c117 bl[117] br[117] wl[10] vdd gnd cell_6t
Xbit_r11_c117 bl[117] br[117] wl[11] vdd gnd cell_6t
Xbit_r12_c117 bl[117] br[117] wl[12] vdd gnd cell_6t
Xbit_r13_c117 bl[117] br[117] wl[13] vdd gnd cell_6t
Xbit_r14_c117 bl[117] br[117] wl[14] vdd gnd cell_6t
Xbit_r15_c117 bl[117] br[117] wl[15] vdd gnd cell_6t
Xbit_r16_c117 bl[117] br[117] wl[16] vdd gnd cell_6t
Xbit_r17_c117 bl[117] br[117] wl[17] vdd gnd cell_6t
Xbit_r18_c117 bl[117] br[117] wl[18] vdd gnd cell_6t
Xbit_r19_c117 bl[117] br[117] wl[19] vdd gnd cell_6t
Xbit_r20_c117 bl[117] br[117] wl[20] vdd gnd cell_6t
Xbit_r21_c117 bl[117] br[117] wl[21] vdd gnd cell_6t
Xbit_r22_c117 bl[117] br[117] wl[22] vdd gnd cell_6t
Xbit_r23_c117 bl[117] br[117] wl[23] vdd gnd cell_6t
Xbit_r24_c117 bl[117] br[117] wl[24] vdd gnd cell_6t
Xbit_r25_c117 bl[117] br[117] wl[25] vdd gnd cell_6t
Xbit_r26_c117 bl[117] br[117] wl[26] vdd gnd cell_6t
Xbit_r27_c117 bl[117] br[117] wl[27] vdd gnd cell_6t
Xbit_r28_c117 bl[117] br[117] wl[28] vdd gnd cell_6t
Xbit_r29_c117 bl[117] br[117] wl[29] vdd gnd cell_6t
Xbit_r30_c117 bl[117] br[117] wl[30] vdd gnd cell_6t
Xbit_r31_c117 bl[117] br[117] wl[31] vdd gnd cell_6t
Xbit_r32_c117 bl[117] br[117] wl[32] vdd gnd cell_6t
Xbit_r33_c117 bl[117] br[117] wl[33] vdd gnd cell_6t
Xbit_r34_c117 bl[117] br[117] wl[34] vdd gnd cell_6t
Xbit_r35_c117 bl[117] br[117] wl[35] vdd gnd cell_6t
Xbit_r36_c117 bl[117] br[117] wl[36] vdd gnd cell_6t
Xbit_r37_c117 bl[117] br[117] wl[37] vdd gnd cell_6t
Xbit_r38_c117 bl[117] br[117] wl[38] vdd gnd cell_6t
Xbit_r39_c117 bl[117] br[117] wl[39] vdd gnd cell_6t
Xbit_r40_c117 bl[117] br[117] wl[40] vdd gnd cell_6t
Xbit_r41_c117 bl[117] br[117] wl[41] vdd gnd cell_6t
Xbit_r42_c117 bl[117] br[117] wl[42] vdd gnd cell_6t
Xbit_r43_c117 bl[117] br[117] wl[43] vdd gnd cell_6t
Xbit_r44_c117 bl[117] br[117] wl[44] vdd gnd cell_6t
Xbit_r45_c117 bl[117] br[117] wl[45] vdd gnd cell_6t
Xbit_r46_c117 bl[117] br[117] wl[46] vdd gnd cell_6t
Xbit_r47_c117 bl[117] br[117] wl[47] vdd gnd cell_6t
Xbit_r48_c117 bl[117] br[117] wl[48] vdd gnd cell_6t
Xbit_r49_c117 bl[117] br[117] wl[49] vdd gnd cell_6t
Xbit_r50_c117 bl[117] br[117] wl[50] vdd gnd cell_6t
Xbit_r51_c117 bl[117] br[117] wl[51] vdd gnd cell_6t
Xbit_r52_c117 bl[117] br[117] wl[52] vdd gnd cell_6t
Xbit_r53_c117 bl[117] br[117] wl[53] vdd gnd cell_6t
Xbit_r54_c117 bl[117] br[117] wl[54] vdd gnd cell_6t
Xbit_r55_c117 bl[117] br[117] wl[55] vdd gnd cell_6t
Xbit_r56_c117 bl[117] br[117] wl[56] vdd gnd cell_6t
Xbit_r57_c117 bl[117] br[117] wl[57] vdd gnd cell_6t
Xbit_r58_c117 bl[117] br[117] wl[58] vdd gnd cell_6t
Xbit_r59_c117 bl[117] br[117] wl[59] vdd gnd cell_6t
Xbit_r60_c117 bl[117] br[117] wl[60] vdd gnd cell_6t
Xbit_r61_c117 bl[117] br[117] wl[61] vdd gnd cell_6t
Xbit_r62_c117 bl[117] br[117] wl[62] vdd gnd cell_6t
Xbit_r63_c117 bl[117] br[117] wl[63] vdd gnd cell_6t
Xbit_r64_c117 bl[117] br[117] wl[64] vdd gnd cell_6t
Xbit_r65_c117 bl[117] br[117] wl[65] vdd gnd cell_6t
Xbit_r66_c117 bl[117] br[117] wl[66] vdd gnd cell_6t
Xbit_r67_c117 bl[117] br[117] wl[67] vdd gnd cell_6t
Xbit_r68_c117 bl[117] br[117] wl[68] vdd gnd cell_6t
Xbit_r69_c117 bl[117] br[117] wl[69] vdd gnd cell_6t
Xbit_r70_c117 bl[117] br[117] wl[70] vdd gnd cell_6t
Xbit_r71_c117 bl[117] br[117] wl[71] vdd gnd cell_6t
Xbit_r72_c117 bl[117] br[117] wl[72] vdd gnd cell_6t
Xbit_r73_c117 bl[117] br[117] wl[73] vdd gnd cell_6t
Xbit_r74_c117 bl[117] br[117] wl[74] vdd gnd cell_6t
Xbit_r75_c117 bl[117] br[117] wl[75] vdd gnd cell_6t
Xbit_r76_c117 bl[117] br[117] wl[76] vdd gnd cell_6t
Xbit_r77_c117 bl[117] br[117] wl[77] vdd gnd cell_6t
Xbit_r78_c117 bl[117] br[117] wl[78] vdd gnd cell_6t
Xbit_r79_c117 bl[117] br[117] wl[79] vdd gnd cell_6t
Xbit_r80_c117 bl[117] br[117] wl[80] vdd gnd cell_6t
Xbit_r81_c117 bl[117] br[117] wl[81] vdd gnd cell_6t
Xbit_r82_c117 bl[117] br[117] wl[82] vdd gnd cell_6t
Xbit_r83_c117 bl[117] br[117] wl[83] vdd gnd cell_6t
Xbit_r84_c117 bl[117] br[117] wl[84] vdd gnd cell_6t
Xbit_r85_c117 bl[117] br[117] wl[85] vdd gnd cell_6t
Xbit_r86_c117 bl[117] br[117] wl[86] vdd gnd cell_6t
Xbit_r87_c117 bl[117] br[117] wl[87] vdd gnd cell_6t
Xbit_r88_c117 bl[117] br[117] wl[88] vdd gnd cell_6t
Xbit_r89_c117 bl[117] br[117] wl[89] vdd gnd cell_6t
Xbit_r90_c117 bl[117] br[117] wl[90] vdd gnd cell_6t
Xbit_r91_c117 bl[117] br[117] wl[91] vdd gnd cell_6t
Xbit_r92_c117 bl[117] br[117] wl[92] vdd gnd cell_6t
Xbit_r93_c117 bl[117] br[117] wl[93] vdd gnd cell_6t
Xbit_r94_c117 bl[117] br[117] wl[94] vdd gnd cell_6t
Xbit_r95_c117 bl[117] br[117] wl[95] vdd gnd cell_6t
Xbit_r96_c117 bl[117] br[117] wl[96] vdd gnd cell_6t
Xbit_r97_c117 bl[117] br[117] wl[97] vdd gnd cell_6t
Xbit_r98_c117 bl[117] br[117] wl[98] vdd gnd cell_6t
Xbit_r99_c117 bl[117] br[117] wl[99] vdd gnd cell_6t
Xbit_r100_c117 bl[117] br[117] wl[100] vdd gnd cell_6t
Xbit_r101_c117 bl[117] br[117] wl[101] vdd gnd cell_6t
Xbit_r102_c117 bl[117] br[117] wl[102] vdd gnd cell_6t
Xbit_r103_c117 bl[117] br[117] wl[103] vdd gnd cell_6t
Xbit_r104_c117 bl[117] br[117] wl[104] vdd gnd cell_6t
Xbit_r105_c117 bl[117] br[117] wl[105] vdd gnd cell_6t
Xbit_r106_c117 bl[117] br[117] wl[106] vdd gnd cell_6t
Xbit_r107_c117 bl[117] br[117] wl[107] vdd gnd cell_6t
Xbit_r108_c117 bl[117] br[117] wl[108] vdd gnd cell_6t
Xbit_r109_c117 bl[117] br[117] wl[109] vdd gnd cell_6t
Xbit_r110_c117 bl[117] br[117] wl[110] vdd gnd cell_6t
Xbit_r111_c117 bl[117] br[117] wl[111] vdd gnd cell_6t
Xbit_r112_c117 bl[117] br[117] wl[112] vdd gnd cell_6t
Xbit_r113_c117 bl[117] br[117] wl[113] vdd gnd cell_6t
Xbit_r114_c117 bl[117] br[117] wl[114] vdd gnd cell_6t
Xbit_r115_c117 bl[117] br[117] wl[115] vdd gnd cell_6t
Xbit_r116_c117 bl[117] br[117] wl[116] vdd gnd cell_6t
Xbit_r117_c117 bl[117] br[117] wl[117] vdd gnd cell_6t
Xbit_r118_c117 bl[117] br[117] wl[118] vdd gnd cell_6t
Xbit_r119_c117 bl[117] br[117] wl[119] vdd gnd cell_6t
Xbit_r120_c117 bl[117] br[117] wl[120] vdd gnd cell_6t
Xbit_r121_c117 bl[117] br[117] wl[121] vdd gnd cell_6t
Xbit_r122_c117 bl[117] br[117] wl[122] vdd gnd cell_6t
Xbit_r123_c117 bl[117] br[117] wl[123] vdd gnd cell_6t
Xbit_r124_c117 bl[117] br[117] wl[124] vdd gnd cell_6t
Xbit_r125_c117 bl[117] br[117] wl[125] vdd gnd cell_6t
Xbit_r126_c117 bl[117] br[117] wl[126] vdd gnd cell_6t
Xbit_r127_c117 bl[117] br[117] wl[127] vdd gnd cell_6t
Xbit_r128_c117 bl[117] br[117] wl[128] vdd gnd cell_6t
Xbit_r129_c117 bl[117] br[117] wl[129] vdd gnd cell_6t
Xbit_r130_c117 bl[117] br[117] wl[130] vdd gnd cell_6t
Xbit_r131_c117 bl[117] br[117] wl[131] vdd gnd cell_6t
Xbit_r132_c117 bl[117] br[117] wl[132] vdd gnd cell_6t
Xbit_r133_c117 bl[117] br[117] wl[133] vdd gnd cell_6t
Xbit_r134_c117 bl[117] br[117] wl[134] vdd gnd cell_6t
Xbit_r135_c117 bl[117] br[117] wl[135] vdd gnd cell_6t
Xbit_r136_c117 bl[117] br[117] wl[136] vdd gnd cell_6t
Xbit_r137_c117 bl[117] br[117] wl[137] vdd gnd cell_6t
Xbit_r138_c117 bl[117] br[117] wl[138] vdd gnd cell_6t
Xbit_r139_c117 bl[117] br[117] wl[139] vdd gnd cell_6t
Xbit_r140_c117 bl[117] br[117] wl[140] vdd gnd cell_6t
Xbit_r141_c117 bl[117] br[117] wl[141] vdd gnd cell_6t
Xbit_r142_c117 bl[117] br[117] wl[142] vdd gnd cell_6t
Xbit_r143_c117 bl[117] br[117] wl[143] vdd gnd cell_6t
Xbit_r144_c117 bl[117] br[117] wl[144] vdd gnd cell_6t
Xbit_r145_c117 bl[117] br[117] wl[145] vdd gnd cell_6t
Xbit_r146_c117 bl[117] br[117] wl[146] vdd gnd cell_6t
Xbit_r147_c117 bl[117] br[117] wl[147] vdd gnd cell_6t
Xbit_r148_c117 bl[117] br[117] wl[148] vdd gnd cell_6t
Xbit_r149_c117 bl[117] br[117] wl[149] vdd gnd cell_6t
Xbit_r150_c117 bl[117] br[117] wl[150] vdd gnd cell_6t
Xbit_r151_c117 bl[117] br[117] wl[151] vdd gnd cell_6t
Xbit_r152_c117 bl[117] br[117] wl[152] vdd gnd cell_6t
Xbit_r153_c117 bl[117] br[117] wl[153] vdd gnd cell_6t
Xbit_r154_c117 bl[117] br[117] wl[154] vdd gnd cell_6t
Xbit_r155_c117 bl[117] br[117] wl[155] vdd gnd cell_6t
Xbit_r156_c117 bl[117] br[117] wl[156] vdd gnd cell_6t
Xbit_r157_c117 bl[117] br[117] wl[157] vdd gnd cell_6t
Xbit_r158_c117 bl[117] br[117] wl[158] vdd gnd cell_6t
Xbit_r159_c117 bl[117] br[117] wl[159] vdd gnd cell_6t
Xbit_r160_c117 bl[117] br[117] wl[160] vdd gnd cell_6t
Xbit_r161_c117 bl[117] br[117] wl[161] vdd gnd cell_6t
Xbit_r162_c117 bl[117] br[117] wl[162] vdd gnd cell_6t
Xbit_r163_c117 bl[117] br[117] wl[163] vdd gnd cell_6t
Xbit_r164_c117 bl[117] br[117] wl[164] vdd gnd cell_6t
Xbit_r165_c117 bl[117] br[117] wl[165] vdd gnd cell_6t
Xbit_r166_c117 bl[117] br[117] wl[166] vdd gnd cell_6t
Xbit_r167_c117 bl[117] br[117] wl[167] vdd gnd cell_6t
Xbit_r168_c117 bl[117] br[117] wl[168] vdd gnd cell_6t
Xbit_r169_c117 bl[117] br[117] wl[169] vdd gnd cell_6t
Xbit_r170_c117 bl[117] br[117] wl[170] vdd gnd cell_6t
Xbit_r171_c117 bl[117] br[117] wl[171] vdd gnd cell_6t
Xbit_r172_c117 bl[117] br[117] wl[172] vdd gnd cell_6t
Xbit_r173_c117 bl[117] br[117] wl[173] vdd gnd cell_6t
Xbit_r174_c117 bl[117] br[117] wl[174] vdd gnd cell_6t
Xbit_r175_c117 bl[117] br[117] wl[175] vdd gnd cell_6t
Xbit_r176_c117 bl[117] br[117] wl[176] vdd gnd cell_6t
Xbit_r177_c117 bl[117] br[117] wl[177] vdd gnd cell_6t
Xbit_r178_c117 bl[117] br[117] wl[178] vdd gnd cell_6t
Xbit_r179_c117 bl[117] br[117] wl[179] vdd gnd cell_6t
Xbit_r180_c117 bl[117] br[117] wl[180] vdd gnd cell_6t
Xbit_r181_c117 bl[117] br[117] wl[181] vdd gnd cell_6t
Xbit_r182_c117 bl[117] br[117] wl[182] vdd gnd cell_6t
Xbit_r183_c117 bl[117] br[117] wl[183] vdd gnd cell_6t
Xbit_r184_c117 bl[117] br[117] wl[184] vdd gnd cell_6t
Xbit_r185_c117 bl[117] br[117] wl[185] vdd gnd cell_6t
Xbit_r186_c117 bl[117] br[117] wl[186] vdd gnd cell_6t
Xbit_r187_c117 bl[117] br[117] wl[187] vdd gnd cell_6t
Xbit_r188_c117 bl[117] br[117] wl[188] vdd gnd cell_6t
Xbit_r189_c117 bl[117] br[117] wl[189] vdd gnd cell_6t
Xbit_r190_c117 bl[117] br[117] wl[190] vdd gnd cell_6t
Xbit_r191_c117 bl[117] br[117] wl[191] vdd gnd cell_6t
Xbit_r192_c117 bl[117] br[117] wl[192] vdd gnd cell_6t
Xbit_r193_c117 bl[117] br[117] wl[193] vdd gnd cell_6t
Xbit_r194_c117 bl[117] br[117] wl[194] vdd gnd cell_6t
Xbit_r195_c117 bl[117] br[117] wl[195] vdd gnd cell_6t
Xbit_r196_c117 bl[117] br[117] wl[196] vdd gnd cell_6t
Xbit_r197_c117 bl[117] br[117] wl[197] vdd gnd cell_6t
Xbit_r198_c117 bl[117] br[117] wl[198] vdd gnd cell_6t
Xbit_r199_c117 bl[117] br[117] wl[199] vdd gnd cell_6t
Xbit_r200_c117 bl[117] br[117] wl[200] vdd gnd cell_6t
Xbit_r201_c117 bl[117] br[117] wl[201] vdd gnd cell_6t
Xbit_r202_c117 bl[117] br[117] wl[202] vdd gnd cell_6t
Xbit_r203_c117 bl[117] br[117] wl[203] vdd gnd cell_6t
Xbit_r204_c117 bl[117] br[117] wl[204] vdd gnd cell_6t
Xbit_r205_c117 bl[117] br[117] wl[205] vdd gnd cell_6t
Xbit_r206_c117 bl[117] br[117] wl[206] vdd gnd cell_6t
Xbit_r207_c117 bl[117] br[117] wl[207] vdd gnd cell_6t
Xbit_r208_c117 bl[117] br[117] wl[208] vdd gnd cell_6t
Xbit_r209_c117 bl[117] br[117] wl[209] vdd gnd cell_6t
Xbit_r210_c117 bl[117] br[117] wl[210] vdd gnd cell_6t
Xbit_r211_c117 bl[117] br[117] wl[211] vdd gnd cell_6t
Xbit_r212_c117 bl[117] br[117] wl[212] vdd gnd cell_6t
Xbit_r213_c117 bl[117] br[117] wl[213] vdd gnd cell_6t
Xbit_r214_c117 bl[117] br[117] wl[214] vdd gnd cell_6t
Xbit_r215_c117 bl[117] br[117] wl[215] vdd gnd cell_6t
Xbit_r216_c117 bl[117] br[117] wl[216] vdd gnd cell_6t
Xbit_r217_c117 bl[117] br[117] wl[217] vdd gnd cell_6t
Xbit_r218_c117 bl[117] br[117] wl[218] vdd gnd cell_6t
Xbit_r219_c117 bl[117] br[117] wl[219] vdd gnd cell_6t
Xbit_r220_c117 bl[117] br[117] wl[220] vdd gnd cell_6t
Xbit_r221_c117 bl[117] br[117] wl[221] vdd gnd cell_6t
Xbit_r222_c117 bl[117] br[117] wl[222] vdd gnd cell_6t
Xbit_r223_c117 bl[117] br[117] wl[223] vdd gnd cell_6t
Xbit_r224_c117 bl[117] br[117] wl[224] vdd gnd cell_6t
Xbit_r225_c117 bl[117] br[117] wl[225] vdd gnd cell_6t
Xbit_r226_c117 bl[117] br[117] wl[226] vdd gnd cell_6t
Xbit_r227_c117 bl[117] br[117] wl[227] vdd gnd cell_6t
Xbit_r228_c117 bl[117] br[117] wl[228] vdd gnd cell_6t
Xbit_r229_c117 bl[117] br[117] wl[229] vdd gnd cell_6t
Xbit_r230_c117 bl[117] br[117] wl[230] vdd gnd cell_6t
Xbit_r231_c117 bl[117] br[117] wl[231] vdd gnd cell_6t
Xbit_r232_c117 bl[117] br[117] wl[232] vdd gnd cell_6t
Xbit_r233_c117 bl[117] br[117] wl[233] vdd gnd cell_6t
Xbit_r234_c117 bl[117] br[117] wl[234] vdd gnd cell_6t
Xbit_r235_c117 bl[117] br[117] wl[235] vdd gnd cell_6t
Xbit_r236_c117 bl[117] br[117] wl[236] vdd gnd cell_6t
Xbit_r237_c117 bl[117] br[117] wl[237] vdd gnd cell_6t
Xbit_r238_c117 bl[117] br[117] wl[238] vdd gnd cell_6t
Xbit_r239_c117 bl[117] br[117] wl[239] vdd gnd cell_6t
Xbit_r240_c117 bl[117] br[117] wl[240] vdd gnd cell_6t
Xbit_r241_c117 bl[117] br[117] wl[241] vdd gnd cell_6t
Xbit_r242_c117 bl[117] br[117] wl[242] vdd gnd cell_6t
Xbit_r243_c117 bl[117] br[117] wl[243] vdd gnd cell_6t
Xbit_r244_c117 bl[117] br[117] wl[244] vdd gnd cell_6t
Xbit_r245_c117 bl[117] br[117] wl[245] vdd gnd cell_6t
Xbit_r246_c117 bl[117] br[117] wl[246] vdd gnd cell_6t
Xbit_r247_c117 bl[117] br[117] wl[247] vdd gnd cell_6t
Xbit_r248_c117 bl[117] br[117] wl[248] vdd gnd cell_6t
Xbit_r249_c117 bl[117] br[117] wl[249] vdd gnd cell_6t
Xbit_r250_c117 bl[117] br[117] wl[250] vdd gnd cell_6t
Xbit_r251_c117 bl[117] br[117] wl[251] vdd gnd cell_6t
Xbit_r252_c117 bl[117] br[117] wl[252] vdd gnd cell_6t
Xbit_r253_c117 bl[117] br[117] wl[253] vdd gnd cell_6t
Xbit_r254_c117 bl[117] br[117] wl[254] vdd gnd cell_6t
Xbit_r255_c117 bl[117] br[117] wl[255] vdd gnd cell_6t
Xbit_r0_c118 bl[118] br[118] wl[0] vdd gnd cell_6t
Xbit_r1_c118 bl[118] br[118] wl[1] vdd gnd cell_6t
Xbit_r2_c118 bl[118] br[118] wl[2] vdd gnd cell_6t
Xbit_r3_c118 bl[118] br[118] wl[3] vdd gnd cell_6t
Xbit_r4_c118 bl[118] br[118] wl[4] vdd gnd cell_6t
Xbit_r5_c118 bl[118] br[118] wl[5] vdd gnd cell_6t
Xbit_r6_c118 bl[118] br[118] wl[6] vdd gnd cell_6t
Xbit_r7_c118 bl[118] br[118] wl[7] vdd gnd cell_6t
Xbit_r8_c118 bl[118] br[118] wl[8] vdd gnd cell_6t
Xbit_r9_c118 bl[118] br[118] wl[9] vdd gnd cell_6t
Xbit_r10_c118 bl[118] br[118] wl[10] vdd gnd cell_6t
Xbit_r11_c118 bl[118] br[118] wl[11] vdd gnd cell_6t
Xbit_r12_c118 bl[118] br[118] wl[12] vdd gnd cell_6t
Xbit_r13_c118 bl[118] br[118] wl[13] vdd gnd cell_6t
Xbit_r14_c118 bl[118] br[118] wl[14] vdd gnd cell_6t
Xbit_r15_c118 bl[118] br[118] wl[15] vdd gnd cell_6t
Xbit_r16_c118 bl[118] br[118] wl[16] vdd gnd cell_6t
Xbit_r17_c118 bl[118] br[118] wl[17] vdd gnd cell_6t
Xbit_r18_c118 bl[118] br[118] wl[18] vdd gnd cell_6t
Xbit_r19_c118 bl[118] br[118] wl[19] vdd gnd cell_6t
Xbit_r20_c118 bl[118] br[118] wl[20] vdd gnd cell_6t
Xbit_r21_c118 bl[118] br[118] wl[21] vdd gnd cell_6t
Xbit_r22_c118 bl[118] br[118] wl[22] vdd gnd cell_6t
Xbit_r23_c118 bl[118] br[118] wl[23] vdd gnd cell_6t
Xbit_r24_c118 bl[118] br[118] wl[24] vdd gnd cell_6t
Xbit_r25_c118 bl[118] br[118] wl[25] vdd gnd cell_6t
Xbit_r26_c118 bl[118] br[118] wl[26] vdd gnd cell_6t
Xbit_r27_c118 bl[118] br[118] wl[27] vdd gnd cell_6t
Xbit_r28_c118 bl[118] br[118] wl[28] vdd gnd cell_6t
Xbit_r29_c118 bl[118] br[118] wl[29] vdd gnd cell_6t
Xbit_r30_c118 bl[118] br[118] wl[30] vdd gnd cell_6t
Xbit_r31_c118 bl[118] br[118] wl[31] vdd gnd cell_6t
Xbit_r32_c118 bl[118] br[118] wl[32] vdd gnd cell_6t
Xbit_r33_c118 bl[118] br[118] wl[33] vdd gnd cell_6t
Xbit_r34_c118 bl[118] br[118] wl[34] vdd gnd cell_6t
Xbit_r35_c118 bl[118] br[118] wl[35] vdd gnd cell_6t
Xbit_r36_c118 bl[118] br[118] wl[36] vdd gnd cell_6t
Xbit_r37_c118 bl[118] br[118] wl[37] vdd gnd cell_6t
Xbit_r38_c118 bl[118] br[118] wl[38] vdd gnd cell_6t
Xbit_r39_c118 bl[118] br[118] wl[39] vdd gnd cell_6t
Xbit_r40_c118 bl[118] br[118] wl[40] vdd gnd cell_6t
Xbit_r41_c118 bl[118] br[118] wl[41] vdd gnd cell_6t
Xbit_r42_c118 bl[118] br[118] wl[42] vdd gnd cell_6t
Xbit_r43_c118 bl[118] br[118] wl[43] vdd gnd cell_6t
Xbit_r44_c118 bl[118] br[118] wl[44] vdd gnd cell_6t
Xbit_r45_c118 bl[118] br[118] wl[45] vdd gnd cell_6t
Xbit_r46_c118 bl[118] br[118] wl[46] vdd gnd cell_6t
Xbit_r47_c118 bl[118] br[118] wl[47] vdd gnd cell_6t
Xbit_r48_c118 bl[118] br[118] wl[48] vdd gnd cell_6t
Xbit_r49_c118 bl[118] br[118] wl[49] vdd gnd cell_6t
Xbit_r50_c118 bl[118] br[118] wl[50] vdd gnd cell_6t
Xbit_r51_c118 bl[118] br[118] wl[51] vdd gnd cell_6t
Xbit_r52_c118 bl[118] br[118] wl[52] vdd gnd cell_6t
Xbit_r53_c118 bl[118] br[118] wl[53] vdd gnd cell_6t
Xbit_r54_c118 bl[118] br[118] wl[54] vdd gnd cell_6t
Xbit_r55_c118 bl[118] br[118] wl[55] vdd gnd cell_6t
Xbit_r56_c118 bl[118] br[118] wl[56] vdd gnd cell_6t
Xbit_r57_c118 bl[118] br[118] wl[57] vdd gnd cell_6t
Xbit_r58_c118 bl[118] br[118] wl[58] vdd gnd cell_6t
Xbit_r59_c118 bl[118] br[118] wl[59] vdd gnd cell_6t
Xbit_r60_c118 bl[118] br[118] wl[60] vdd gnd cell_6t
Xbit_r61_c118 bl[118] br[118] wl[61] vdd gnd cell_6t
Xbit_r62_c118 bl[118] br[118] wl[62] vdd gnd cell_6t
Xbit_r63_c118 bl[118] br[118] wl[63] vdd gnd cell_6t
Xbit_r64_c118 bl[118] br[118] wl[64] vdd gnd cell_6t
Xbit_r65_c118 bl[118] br[118] wl[65] vdd gnd cell_6t
Xbit_r66_c118 bl[118] br[118] wl[66] vdd gnd cell_6t
Xbit_r67_c118 bl[118] br[118] wl[67] vdd gnd cell_6t
Xbit_r68_c118 bl[118] br[118] wl[68] vdd gnd cell_6t
Xbit_r69_c118 bl[118] br[118] wl[69] vdd gnd cell_6t
Xbit_r70_c118 bl[118] br[118] wl[70] vdd gnd cell_6t
Xbit_r71_c118 bl[118] br[118] wl[71] vdd gnd cell_6t
Xbit_r72_c118 bl[118] br[118] wl[72] vdd gnd cell_6t
Xbit_r73_c118 bl[118] br[118] wl[73] vdd gnd cell_6t
Xbit_r74_c118 bl[118] br[118] wl[74] vdd gnd cell_6t
Xbit_r75_c118 bl[118] br[118] wl[75] vdd gnd cell_6t
Xbit_r76_c118 bl[118] br[118] wl[76] vdd gnd cell_6t
Xbit_r77_c118 bl[118] br[118] wl[77] vdd gnd cell_6t
Xbit_r78_c118 bl[118] br[118] wl[78] vdd gnd cell_6t
Xbit_r79_c118 bl[118] br[118] wl[79] vdd gnd cell_6t
Xbit_r80_c118 bl[118] br[118] wl[80] vdd gnd cell_6t
Xbit_r81_c118 bl[118] br[118] wl[81] vdd gnd cell_6t
Xbit_r82_c118 bl[118] br[118] wl[82] vdd gnd cell_6t
Xbit_r83_c118 bl[118] br[118] wl[83] vdd gnd cell_6t
Xbit_r84_c118 bl[118] br[118] wl[84] vdd gnd cell_6t
Xbit_r85_c118 bl[118] br[118] wl[85] vdd gnd cell_6t
Xbit_r86_c118 bl[118] br[118] wl[86] vdd gnd cell_6t
Xbit_r87_c118 bl[118] br[118] wl[87] vdd gnd cell_6t
Xbit_r88_c118 bl[118] br[118] wl[88] vdd gnd cell_6t
Xbit_r89_c118 bl[118] br[118] wl[89] vdd gnd cell_6t
Xbit_r90_c118 bl[118] br[118] wl[90] vdd gnd cell_6t
Xbit_r91_c118 bl[118] br[118] wl[91] vdd gnd cell_6t
Xbit_r92_c118 bl[118] br[118] wl[92] vdd gnd cell_6t
Xbit_r93_c118 bl[118] br[118] wl[93] vdd gnd cell_6t
Xbit_r94_c118 bl[118] br[118] wl[94] vdd gnd cell_6t
Xbit_r95_c118 bl[118] br[118] wl[95] vdd gnd cell_6t
Xbit_r96_c118 bl[118] br[118] wl[96] vdd gnd cell_6t
Xbit_r97_c118 bl[118] br[118] wl[97] vdd gnd cell_6t
Xbit_r98_c118 bl[118] br[118] wl[98] vdd gnd cell_6t
Xbit_r99_c118 bl[118] br[118] wl[99] vdd gnd cell_6t
Xbit_r100_c118 bl[118] br[118] wl[100] vdd gnd cell_6t
Xbit_r101_c118 bl[118] br[118] wl[101] vdd gnd cell_6t
Xbit_r102_c118 bl[118] br[118] wl[102] vdd gnd cell_6t
Xbit_r103_c118 bl[118] br[118] wl[103] vdd gnd cell_6t
Xbit_r104_c118 bl[118] br[118] wl[104] vdd gnd cell_6t
Xbit_r105_c118 bl[118] br[118] wl[105] vdd gnd cell_6t
Xbit_r106_c118 bl[118] br[118] wl[106] vdd gnd cell_6t
Xbit_r107_c118 bl[118] br[118] wl[107] vdd gnd cell_6t
Xbit_r108_c118 bl[118] br[118] wl[108] vdd gnd cell_6t
Xbit_r109_c118 bl[118] br[118] wl[109] vdd gnd cell_6t
Xbit_r110_c118 bl[118] br[118] wl[110] vdd gnd cell_6t
Xbit_r111_c118 bl[118] br[118] wl[111] vdd gnd cell_6t
Xbit_r112_c118 bl[118] br[118] wl[112] vdd gnd cell_6t
Xbit_r113_c118 bl[118] br[118] wl[113] vdd gnd cell_6t
Xbit_r114_c118 bl[118] br[118] wl[114] vdd gnd cell_6t
Xbit_r115_c118 bl[118] br[118] wl[115] vdd gnd cell_6t
Xbit_r116_c118 bl[118] br[118] wl[116] vdd gnd cell_6t
Xbit_r117_c118 bl[118] br[118] wl[117] vdd gnd cell_6t
Xbit_r118_c118 bl[118] br[118] wl[118] vdd gnd cell_6t
Xbit_r119_c118 bl[118] br[118] wl[119] vdd gnd cell_6t
Xbit_r120_c118 bl[118] br[118] wl[120] vdd gnd cell_6t
Xbit_r121_c118 bl[118] br[118] wl[121] vdd gnd cell_6t
Xbit_r122_c118 bl[118] br[118] wl[122] vdd gnd cell_6t
Xbit_r123_c118 bl[118] br[118] wl[123] vdd gnd cell_6t
Xbit_r124_c118 bl[118] br[118] wl[124] vdd gnd cell_6t
Xbit_r125_c118 bl[118] br[118] wl[125] vdd gnd cell_6t
Xbit_r126_c118 bl[118] br[118] wl[126] vdd gnd cell_6t
Xbit_r127_c118 bl[118] br[118] wl[127] vdd gnd cell_6t
Xbit_r128_c118 bl[118] br[118] wl[128] vdd gnd cell_6t
Xbit_r129_c118 bl[118] br[118] wl[129] vdd gnd cell_6t
Xbit_r130_c118 bl[118] br[118] wl[130] vdd gnd cell_6t
Xbit_r131_c118 bl[118] br[118] wl[131] vdd gnd cell_6t
Xbit_r132_c118 bl[118] br[118] wl[132] vdd gnd cell_6t
Xbit_r133_c118 bl[118] br[118] wl[133] vdd gnd cell_6t
Xbit_r134_c118 bl[118] br[118] wl[134] vdd gnd cell_6t
Xbit_r135_c118 bl[118] br[118] wl[135] vdd gnd cell_6t
Xbit_r136_c118 bl[118] br[118] wl[136] vdd gnd cell_6t
Xbit_r137_c118 bl[118] br[118] wl[137] vdd gnd cell_6t
Xbit_r138_c118 bl[118] br[118] wl[138] vdd gnd cell_6t
Xbit_r139_c118 bl[118] br[118] wl[139] vdd gnd cell_6t
Xbit_r140_c118 bl[118] br[118] wl[140] vdd gnd cell_6t
Xbit_r141_c118 bl[118] br[118] wl[141] vdd gnd cell_6t
Xbit_r142_c118 bl[118] br[118] wl[142] vdd gnd cell_6t
Xbit_r143_c118 bl[118] br[118] wl[143] vdd gnd cell_6t
Xbit_r144_c118 bl[118] br[118] wl[144] vdd gnd cell_6t
Xbit_r145_c118 bl[118] br[118] wl[145] vdd gnd cell_6t
Xbit_r146_c118 bl[118] br[118] wl[146] vdd gnd cell_6t
Xbit_r147_c118 bl[118] br[118] wl[147] vdd gnd cell_6t
Xbit_r148_c118 bl[118] br[118] wl[148] vdd gnd cell_6t
Xbit_r149_c118 bl[118] br[118] wl[149] vdd gnd cell_6t
Xbit_r150_c118 bl[118] br[118] wl[150] vdd gnd cell_6t
Xbit_r151_c118 bl[118] br[118] wl[151] vdd gnd cell_6t
Xbit_r152_c118 bl[118] br[118] wl[152] vdd gnd cell_6t
Xbit_r153_c118 bl[118] br[118] wl[153] vdd gnd cell_6t
Xbit_r154_c118 bl[118] br[118] wl[154] vdd gnd cell_6t
Xbit_r155_c118 bl[118] br[118] wl[155] vdd gnd cell_6t
Xbit_r156_c118 bl[118] br[118] wl[156] vdd gnd cell_6t
Xbit_r157_c118 bl[118] br[118] wl[157] vdd gnd cell_6t
Xbit_r158_c118 bl[118] br[118] wl[158] vdd gnd cell_6t
Xbit_r159_c118 bl[118] br[118] wl[159] vdd gnd cell_6t
Xbit_r160_c118 bl[118] br[118] wl[160] vdd gnd cell_6t
Xbit_r161_c118 bl[118] br[118] wl[161] vdd gnd cell_6t
Xbit_r162_c118 bl[118] br[118] wl[162] vdd gnd cell_6t
Xbit_r163_c118 bl[118] br[118] wl[163] vdd gnd cell_6t
Xbit_r164_c118 bl[118] br[118] wl[164] vdd gnd cell_6t
Xbit_r165_c118 bl[118] br[118] wl[165] vdd gnd cell_6t
Xbit_r166_c118 bl[118] br[118] wl[166] vdd gnd cell_6t
Xbit_r167_c118 bl[118] br[118] wl[167] vdd gnd cell_6t
Xbit_r168_c118 bl[118] br[118] wl[168] vdd gnd cell_6t
Xbit_r169_c118 bl[118] br[118] wl[169] vdd gnd cell_6t
Xbit_r170_c118 bl[118] br[118] wl[170] vdd gnd cell_6t
Xbit_r171_c118 bl[118] br[118] wl[171] vdd gnd cell_6t
Xbit_r172_c118 bl[118] br[118] wl[172] vdd gnd cell_6t
Xbit_r173_c118 bl[118] br[118] wl[173] vdd gnd cell_6t
Xbit_r174_c118 bl[118] br[118] wl[174] vdd gnd cell_6t
Xbit_r175_c118 bl[118] br[118] wl[175] vdd gnd cell_6t
Xbit_r176_c118 bl[118] br[118] wl[176] vdd gnd cell_6t
Xbit_r177_c118 bl[118] br[118] wl[177] vdd gnd cell_6t
Xbit_r178_c118 bl[118] br[118] wl[178] vdd gnd cell_6t
Xbit_r179_c118 bl[118] br[118] wl[179] vdd gnd cell_6t
Xbit_r180_c118 bl[118] br[118] wl[180] vdd gnd cell_6t
Xbit_r181_c118 bl[118] br[118] wl[181] vdd gnd cell_6t
Xbit_r182_c118 bl[118] br[118] wl[182] vdd gnd cell_6t
Xbit_r183_c118 bl[118] br[118] wl[183] vdd gnd cell_6t
Xbit_r184_c118 bl[118] br[118] wl[184] vdd gnd cell_6t
Xbit_r185_c118 bl[118] br[118] wl[185] vdd gnd cell_6t
Xbit_r186_c118 bl[118] br[118] wl[186] vdd gnd cell_6t
Xbit_r187_c118 bl[118] br[118] wl[187] vdd gnd cell_6t
Xbit_r188_c118 bl[118] br[118] wl[188] vdd gnd cell_6t
Xbit_r189_c118 bl[118] br[118] wl[189] vdd gnd cell_6t
Xbit_r190_c118 bl[118] br[118] wl[190] vdd gnd cell_6t
Xbit_r191_c118 bl[118] br[118] wl[191] vdd gnd cell_6t
Xbit_r192_c118 bl[118] br[118] wl[192] vdd gnd cell_6t
Xbit_r193_c118 bl[118] br[118] wl[193] vdd gnd cell_6t
Xbit_r194_c118 bl[118] br[118] wl[194] vdd gnd cell_6t
Xbit_r195_c118 bl[118] br[118] wl[195] vdd gnd cell_6t
Xbit_r196_c118 bl[118] br[118] wl[196] vdd gnd cell_6t
Xbit_r197_c118 bl[118] br[118] wl[197] vdd gnd cell_6t
Xbit_r198_c118 bl[118] br[118] wl[198] vdd gnd cell_6t
Xbit_r199_c118 bl[118] br[118] wl[199] vdd gnd cell_6t
Xbit_r200_c118 bl[118] br[118] wl[200] vdd gnd cell_6t
Xbit_r201_c118 bl[118] br[118] wl[201] vdd gnd cell_6t
Xbit_r202_c118 bl[118] br[118] wl[202] vdd gnd cell_6t
Xbit_r203_c118 bl[118] br[118] wl[203] vdd gnd cell_6t
Xbit_r204_c118 bl[118] br[118] wl[204] vdd gnd cell_6t
Xbit_r205_c118 bl[118] br[118] wl[205] vdd gnd cell_6t
Xbit_r206_c118 bl[118] br[118] wl[206] vdd gnd cell_6t
Xbit_r207_c118 bl[118] br[118] wl[207] vdd gnd cell_6t
Xbit_r208_c118 bl[118] br[118] wl[208] vdd gnd cell_6t
Xbit_r209_c118 bl[118] br[118] wl[209] vdd gnd cell_6t
Xbit_r210_c118 bl[118] br[118] wl[210] vdd gnd cell_6t
Xbit_r211_c118 bl[118] br[118] wl[211] vdd gnd cell_6t
Xbit_r212_c118 bl[118] br[118] wl[212] vdd gnd cell_6t
Xbit_r213_c118 bl[118] br[118] wl[213] vdd gnd cell_6t
Xbit_r214_c118 bl[118] br[118] wl[214] vdd gnd cell_6t
Xbit_r215_c118 bl[118] br[118] wl[215] vdd gnd cell_6t
Xbit_r216_c118 bl[118] br[118] wl[216] vdd gnd cell_6t
Xbit_r217_c118 bl[118] br[118] wl[217] vdd gnd cell_6t
Xbit_r218_c118 bl[118] br[118] wl[218] vdd gnd cell_6t
Xbit_r219_c118 bl[118] br[118] wl[219] vdd gnd cell_6t
Xbit_r220_c118 bl[118] br[118] wl[220] vdd gnd cell_6t
Xbit_r221_c118 bl[118] br[118] wl[221] vdd gnd cell_6t
Xbit_r222_c118 bl[118] br[118] wl[222] vdd gnd cell_6t
Xbit_r223_c118 bl[118] br[118] wl[223] vdd gnd cell_6t
Xbit_r224_c118 bl[118] br[118] wl[224] vdd gnd cell_6t
Xbit_r225_c118 bl[118] br[118] wl[225] vdd gnd cell_6t
Xbit_r226_c118 bl[118] br[118] wl[226] vdd gnd cell_6t
Xbit_r227_c118 bl[118] br[118] wl[227] vdd gnd cell_6t
Xbit_r228_c118 bl[118] br[118] wl[228] vdd gnd cell_6t
Xbit_r229_c118 bl[118] br[118] wl[229] vdd gnd cell_6t
Xbit_r230_c118 bl[118] br[118] wl[230] vdd gnd cell_6t
Xbit_r231_c118 bl[118] br[118] wl[231] vdd gnd cell_6t
Xbit_r232_c118 bl[118] br[118] wl[232] vdd gnd cell_6t
Xbit_r233_c118 bl[118] br[118] wl[233] vdd gnd cell_6t
Xbit_r234_c118 bl[118] br[118] wl[234] vdd gnd cell_6t
Xbit_r235_c118 bl[118] br[118] wl[235] vdd gnd cell_6t
Xbit_r236_c118 bl[118] br[118] wl[236] vdd gnd cell_6t
Xbit_r237_c118 bl[118] br[118] wl[237] vdd gnd cell_6t
Xbit_r238_c118 bl[118] br[118] wl[238] vdd gnd cell_6t
Xbit_r239_c118 bl[118] br[118] wl[239] vdd gnd cell_6t
Xbit_r240_c118 bl[118] br[118] wl[240] vdd gnd cell_6t
Xbit_r241_c118 bl[118] br[118] wl[241] vdd gnd cell_6t
Xbit_r242_c118 bl[118] br[118] wl[242] vdd gnd cell_6t
Xbit_r243_c118 bl[118] br[118] wl[243] vdd gnd cell_6t
Xbit_r244_c118 bl[118] br[118] wl[244] vdd gnd cell_6t
Xbit_r245_c118 bl[118] br[118] wl[245] vdd gnd cell_6t
Xbit_r246_c118 bl[118] br[118] wl[246] vdd gnd cell_6t
Xbit_r247_c118 bl[118] br[118] wl[247] vdd gnd cell_6t
Xbit_r248_c118 bl[118] br[118] wl[248] vdd gnd cell_6t
Xbit_r249_c118 bl[118] br[118] wl[249] vdd gnd cell_6t
Xbit_r250_c118 bl[118] br[118] wl[250] vdd gnd cell_6t
Xbit_r251_c118 bl[118] br[118] wl[251] vdd gnd cell_6t
Xbit_r252_c118 bl[118] br[118] wl[252] vdd gnd cell_6t
Xbit_r253_c118 bl[118] br[118] wl[253] vdd gnd cell_6t
Xbit_r254_c118 bl[118] br[118] wl[254] vdd gnd cell_6t
Xbit_r255_c118 bl[118] br[118] wl[255] vdd gnd cell_6t
Xbit_r0_c119 bl[119] br[119] wl[0] vdd gnd cell_6t
Xbit_r1_c119 bl[119] br[119] wl[1] vdd gnd cell_6t
Xbit_r2_c119 bl[119] br[119] wl[2] vdd gnd cell_6t
Xbit_r3_c119 bl[119] br[119] wl[3] vdd gnd cell_6t
Xbit_r4_c119 bl[119] br[119] wl[4] vdd gnd cell_6t
Xbit_r5_c119 bl[119] br[119] wl[5] vdd gnd cell_6t
Xbit_r6_c119 bl[119] br[119] wl[6] vdd gnd cell_6t
Xbit_r7_c119 bl[119] br[119] wl[7] vdd gnd cell_6t
Xbit_r8_c119 bl[119] br[119] wl[8] vdd gnd cell_6t
Xbit_r9_c119 bl[119] br[119] wl[9] vdd gnd cell_6t
Xbit_r10_c119 bl[119] br[119] wl[10] vdd gnd cell_6t
Xbit_r11_c119 bl[119] br[119] wl[11] vdd gnd cell_6t
Xbit_r12_c119 bl[119] br[119] wl[12] vdd gnd cell_6t
Xbit_r13_c119 bl[119] br[119] wl[13] vdd gnd cell_6t
Xbit_r14_c119 bl[119] br[119] wl[14] vdd gnd cell_6t
Xbit_r15_c119 bl[119] br[119] wl[15] vdd gnd cell_6t
Xbit_r16_c119 bl[119] br[119] wl[16] vdd gnd cell_6t
Xbit_r17_c119 bl[119] br[119] wl[17] vdd gnd cell_6t
Xbit_r18_c119 bl[119] br[119] wl[18] vdd gnd cell_6t
Xbit_r19_c119 bl[119] br[119] wl[19] vdd gnd cell_6t
Xbit_r20_c119 bl[119] br[119] wl[20] vdd gnd cell_6t
Xbit_r21_c119 bl[119] br[119] wl[21] vdd gnd cell_6t
Xbit_r22_c119 bl[119] br[119] wl[22] vdd gnd cell_6t
Xbit_r23_c119 bl[119] br[119] wl[23] vdd gnd cell_6t
Xbit_r24_c119 bl[119] br[119] wl[24] vdd gnd cell_6t
Xbit_r25_c119 bl[119] br[119] wl[25] vdd gnd cell_6t
Xbit_r26_c119 bl[119] br[119] wl[26] vdd gnd cell_6t
Xbit_r27_c119 bl[119] br[119] wl[27] vdd gnd cell_6t
Xbit_r28_c119 bl[119] br[119] wl[28] vdd gnd cell_6t
Xbit_r29_c119 bl[119] br[119] wl[29] vdd gnd cell_6t
Xbit_r30_c119 bl[119] br[119] wl[30] vdd gnd cell_6t
Xbit_r31_c119 bl[119] br[119] wl[31] vdd gnd cell_6t
Xbit_r32_c119 bl[119] br[119] wl[32] vdd gnd cell_6t
Xbit_r33_c119 bl[119] br[119] wl[33] vdd gnd cell_6t
Xbit_r34_c119 bl[119] br[119] wl[34] vdd gnd cell_6t
Xbit_r35_c119 bl[119] br[119] wl[35] vdd gnd cell_6t
Xbit_r36_c119 bl[119] br[119] wl[36] vdd gnd cell_6t
Xbit_r37_c119 bl[119] br[119] wl[37] vdd gnd cell_6t
Xbit_r38_c119 bl[119] br[119] wl[38] vdd gnd cell_6t
Xbit_r39_c119 bl[119] br[119] wl[39] vdd gnd cell_6t
Xbit_r40_c119 bl[119] br[119] wl[40] vdd gnd cell_6t
Xbit_r41_c119 bl[119] br[119] wl[41] vdd gnd cell_6t
Xbit_r42_c119 bl[119] br[119] wl[42] vdd gnd cell_6t
Xbit_r43_c119 bl[119] br[119] wl[43] vdd gnd cell_6t
Xbit_r44_c119 bl[119] br[119] wl[44] vdd gnd cell_6t
Xbit_r45_c119 bl[119] br[119] wl[45] vdd gnd cell_6t
Xbit_r46_c119 bl[119] br[119] wl[46] vdd gnd cell_6t
Xbit_r47_c119 bl[119] br[119] wl[47] vdd gnd cell_6t
Xbit_r48_c119 bl[119] br[119] wl[48] vdd gnd cell_6t
Xbit_r49_c119 bl[119] br[119] wl[49] vdd gnd cell_6t
Xbit_r50_c119 bl[119] br[119] wl[50] vdd gnd cell_6t
Xbit_r51_c119 bl[119] br[119] wl[51] vdd gnd cell_6t
Xbit_r52_c119 bl[119] br[119] wl[52] vdd gnd cell_6t
Xbit_r53_c119 bl[119] br[119] wl[53] vdd gnd cell_6t
Xbit_r54_c119 bl[119] br[119] wl[54] vdd gnd cell_6t
Xbit_r55_c119 bl[119] br[119] wl[55] vdd gnd cell_6t
Xbit_r56_c119 bl[119] br[119] wl[56] vdd gnd cell_6t
Xbit_r57_c119 bl[119] br[119] wl[57] vdd gnd cell_6t
Xbit_r58_c119 bl[119] br[119] wl[58] vdd gnd cell_6t
Xbit_r59_c119 bl[119] br[119] wl[59] vdd gnd cell_6t
Xbit_r60_c119 bl[119] br[119] wl[60] vdd gnd cell_6t
Xbit_r61_c119 bl[119] br[119] wl[61] vdd gnd cell_6t
Xbit_r62_c119 bl[119] br[119] wl[62] vdd gnd cell_6t
Xbit_r63_c119 bl[119] br[119] wl[63] vdd gnd cell_6t
Xbit_r64_c119 bl[119] br[119] wl[64] vdd gnd cell_6t
Xbit_r65_c119 bl[119] br[119] wl[65] vdd gnd cell_6t
Xbit_r66_c119 bl[119] br[119] wl[66] vdd gnd cell_6t
Xbit_r67_c119 bl[119] br[119] wl[67] vdd gnd cell_6t
Xbit_r68_c119 bl[119] br[119] wl[68] vdd gnd cell_6t
Xbit_r69_c119 bl[119] br[119] wl[69] vdd gnd cell_6t
Xbit_r70_c119 bl[119] br[119] wl[70] vdd gnd cell_6t
Xbit_r71_c119 bl[119] br[119] wl[71] vdd gnd cell_6t
Xbit_r72_c119 bl[119] br[119] wl[72] vdd gnd cell_6t
Xbit_r73_c119 bl[119] br[119] wl[73] vdd gnd cell_6t
Xbit_r74_c119 bl[119] br[119] wl[74] vdd gnd cell_6t
Xbit_r75_c119 bl[119] br[119] wl[75] vdd gnd cell_6t
Xbit_r76_c119 bl[119] br[119] wl[76] vdd gnd cell_6t
Xbit_r77_c119 bl[119] br[119] wl[77] vdd gnd cell_6t
Xbit_r78_c119 bl[119] br[119] wl[78] vdd gnd cell_6t
Xbit_r79_c119 bl[119] br[119] wl[79] vdd gnd cell_6t
Xbit_r80_c119 bl[119] br[119] wl[80] vdd gnd cell_6t
Xbit_r81_c119 bl[119] br[119] wl[81] vdd gnd cell_6t
Xbit_r82_c119 bl[119] br[119] wl[82] vdd gnd cell_6t
Xbit_r83_c119 bl[119] br[119] wl[83] vdd gnd cell_6t
Xbit_r84_c119 bl[119] br[119] wl[84] vdd gnd cell_6t
Xbit_r85_c119 bl[119] br[119] wl[85] vdd gnd cell_6t
Xbit_r86_c119 bl[119] br[119] wl[86] vdd gnd cell_6t
Xbit_r87_c119 bl[119] br[119] wl[87] vdd gnd cell_6t
Xbit_r88_c119 bl[119] br[119] wl[88] vdd gnd cell_6t
Xbit_r89_c119 bl[119] br[119] wl[89] vdd gnd cell_6t
Xbit_r90_c119 bl[119] br[119] wl[90] vdd gnd cell_6t
Xbit_r91_c119 bl[119] br[119] wl[91] vdd gnd cell_6t
Xbit_r92_c119 bl[119] br[119] wl[92] vdd gnd cell_6t
Xbit_r93_c119 bl[119] br[119] wl[93] vdd gnd cell_6t
Xbit_r94_c119 bl[119] br[119] wl[94] vdd gnd cell_6t
Xbit_r95_c119 bl[119] br[119] wl[95] vdd gnd cell_6t
Xbit_r96_c119 bl[119] br[119] wl[96] vdd gnd cell_6t
Xbit_r97_c119 bl[119] br[119] wl[97] vdd gnd cell_6t
Xbit_r98_c119 bl[119] br[119] wl[98] vdd gnd cell_6t
Xbit_r99_c119 bl[119] br[119] wl[99] vdd gnd cell_6t
Xbit_r100_c119 bl[119] br[119] wl[100] vdd gnd cell_6t
Xbit_r101_c119 bl[119] br[119] wl[101] vdd gnd cell_6t
Xbit_r102_c119 bl[119] br[119] wl[102] vdd gnd cell_6t
Xbit_r103_c119 bl[119] br[119] wl[103] vdd gnd cell_6t
Xbit_r104_c119 bl[119] br[119] wl[104] vdd gnd cell_6t
Xbit_r105_c119 bl[119] br[119] wl[105] vdd gnd cell_6t
Xbit_r106_c119 bl[119] br[119] wl[106] vdd gnd cell_6t
Xbit_r107_c119 bl[119] br[119] wl[107] vdd gnd cell_6t
Xbit_r108_c119 bl[119] br[119] wl[108] vdd gnd cell_6t
Xbit_r109_c119 bl[119] br[119] wl[109] vdd gnd cell_6t
Xbit_r110_c119 bl[119] br[119] wl[110] vdd gnd cell_6t
Xbit_r111_c119 bl[119] br[119] wl[111] vdd gnd cell_6t
Xbit_r112_c119 bl[119] br[119] wl[112] vdd gnd cell_6t
Xbit_r113_c119 bl[119] br[119] wl[113] vdd gnd cell_6t
Xbit_r114_c119 bl[119] br[119] wl[114] vdd gnd cell_6t
Xbit_r115_c119 bl[119] br[119] wl[115] vdd gnd cell_6t
Xbit_r116_c119 bl[119] br[119] wl[116] vdd gnd cell_6t
Xbit_r117_c119 bl[119] br[119] wl[117] vdd gnd cell_6t
Xbit_r118_c119 bl[119] br[119] wl[118] vdd gnd cell_6t
Xbit_r119_c119 bl[119] br[119] wl[119] vdd gnd cell_6t
Xbit_r120_c119 bl[119] br[119] wl[120] vdd gnd cell_6t
Xbit_r121_c119 bl[119] br[119] wl[121] vdd gnd cell_6t
Xbit_r122_c119 bl[119] br[119] wl[122] vdd gnd cell_6t
Xbit_r123_c119 bl[119] br[119] wl[123] vdd gnd cell_6t
Xbit_r124_c119 bl[119] br[119] wl[124] vdd gnd cell_6t
Xbit_r125_c119 bl[119] br[119] wl[125] vdd gnd cell_6t
Xbit_r126_c119 bl[119] br[119] wl[126] vdd gnd cell_6t
Xbit_r127_c119 bl[119] br[119] wl[127] vdd gnd cell_6t
Xbit_r128_c119 bl[119] br[119] wl[128] vdd gnd cell_6t
Xbit_r129_c119 bl[119] br[119] wl[129] vdd gnd cell_6t
Xbit_r130_c119 bl[119] br[119] wl[130] vdd gnd cell_6t
Xbit_r131_c119 bl[119] br[119] wl[131] vdd gnd cell_6t
Xbit_r132_c119 bl[119] br[119] wl[132] vdd gnd cell_6t
Xbit_r133_c119 bl[119] br[119] wl[133] vdd gnd cell_6t
Xbit_r134_c119 bl[119] br[119] wl[134] vdd gnd cell_6t
Xbit_r135_c119 bl[119] br[119] wl[135] vdd gnd cell_6t
Xbit_r136_c119 bl[119] br[119] wl[136] vdd gnd cell_6t
Xbit_r137_c119 bl[119] br[119] wl[137] vdd gnd cell_6t
Xbit_r138_c119 bl[119] br[119] wl[138] vdd gnd cell_6t
Xbit_r139_c119 bl[119] br[119] wl[139] vdd gnd cell_6t
Xbit_r140_c119 bl[119] br[119] wl[140] vdd gnd cell_6t
Xbit_r141_c119 bl[119] br[119] wl[141] vdd gnd cell_6t
Xbit_r142_c119 bl[119] br[119] wl[142] vdd gnd cell_6t
Xbit_r143_c119 bl[119] br[119] wl[143] vdd gnd cell_6t
Xbit_r144_c119 bl[119] br[119] wl[144] vdd gnd cell_6t
Xbit_r145_c119 bl[119] br[119] wl[145] vdd gnd cell_6t
Xbit_r146_c119 bl[119] br[119] wl[146] vdd gnd cell_6t
Xbit_r147_c119 bl[119] br[119] wl[147] vdd gnd cell_6t
Xbit_r148_c119 bl[119] br[119] wl[148] vdd gnd cell_6t
Xbit_r149_c119 bl[119] br[119] wl[149] vdd gnd cell_6t
Xbit_r150_c119 bl[119] br[119] wl[150] vdd gnd cell_6t
Xbit_r151_c119 bl[119] br[119] wl[151] vdd gnd cell_6t
Xbit_r152_c119 bl[119] br[119] wl[152] vdd gnd cell_6t
Xbit_r153_c119 bl[119] br[119] wl[153] vdd gnd cell_6t
Xbit_r154_c119 bl[119] br[119] wl[154] vdd gnd cell_6t
Xbit_r155_c119 bl[119] br[119] wl[155] vdd gnd cell_6t
Xbit_r156_c119 bl[119] br[119] wl[156] vdd gnd cell_6t
Xbit_r157_c119 bl[119] br[119] wl[157] vdd gnd cell_6t
Xbit_r158_c119 bl[119] br[119] wl[158] vdd gnd cell_6t
Xbit_r159_c119 bl[119] br[119] wl[159] vdd gnd cell_6t
Xbit_r160_c119 bl[119] br[119] wl[160] vdd gnd cell_6t
Xbit_r161_c119 bl[119] br[119] wl[161] vdd gnd cell_6t
Xbit_r162_c119 bl[119] br[119] wl[162] vdd gnd cell_6t
Xbit_r163_c119 bl[119] br[119] wl[163] vdd gnd cell_6t
Xbit_r164_c119 bl[119] br[119] wl[164] vdd gnd cell_6t
Xbit_r165_c119 bl[119] br[119] wl[165] vdd gnd cell_6t
Xbit_r166_c119 bl[119] br[119] wl[166] vdd gnd cell_6t
Xbit_r167_c119 bl[119] br[119] wl[167] vdd gnd cell_6t
Xbit_r168_c119 bl[119] br[119] wl[168] vdd gnd cell_6t
Xbit_r169_c119 bl[119] br[119] wl[169] vdd gnd cell_6t
Xbit_r170_c119 bl[119] br[119] wl[170] vdd gnd cell_6t
Xbit_r171_c119 bl[119] br[119] wl[171] vdd gnd cell_6t
Xbit_r172_c119 bl[119] br[119] wl[172] vdd gnd cell_6t
Xbit_r173_c119 bl[119] br[119] wl[173] vdd gnd cell_6t
Xbit_r174_c119 bl[119] br[119] wl[174] vdd gnd cell_6t
Xbit_r175_c119 bl[119] br[119] wl[175] vdd gnd cell_6t
Xbit_r176_c119 bl[119] br[119] wl[176] vdd gnd cell_6t
Xbit_r177_c119 bl[119] br[119] wl[177] vdd gnd cell_6t
Xbit_r178_c119 bl[119] br[119] wl[178] vdd gnd cell_6t
Xbit_r179_c119 bl[119] br[119] wl[179] vdd gnd cell_6t
Xbit_r180_c119 bl[119] br[119] wl[180] vdd gnd cell_6t
Xbit_r181_c119 bl[119] br[119] wl[181] vdd gnd cell_6t
Xbit_r182_c119 bl[119] br[119] wl[182] vdd gnd cell_6t
Xbit_r183_c119 bl[119] br[119] wl[183] vdd gnd cell_6t
Xbit_r184_c119 bl[119] br[119] wl[184] vdd gnd cell_6t
Xbit_r185_c119 bl[119] br[119] wl[185] vdd gnd cell_6t
Xbit_r186_c119 bl[119] br[119] wl[186] vdd gnd cell_6t
Xbit_r187_c119 bl[119] br[119] wl[187] vdd gnd cell_6t
Xbit_r188_c119 bl[119] br[119] wl[188] vdd gnd cell_6t
Xbit_r189_c119 bl[119] br[119] wl[189] vdd gnd cell_6t
Xbit_r190_c119 bl[119] br[119] wl[190] vdd gnd cell_6t
Xbit_r191_c119 bl[119] br[119] wl[191] vdd gnd cell_6t
Xbit_r192_c119 bl[119] br[119] wl[192] vdd gnd cell_6t
Xbit_r193_c119 bl[119] br[119] wl[193] vdd gnd cell_6t
Xbit_r194_c119 bl[119] br[119] wl[194] vdd gnd cell_6t
Xbit_r195_c119 bl[119] br[119] wl[195] vdd gnd cell_6t
Xbit_r196_c119 bl[119] br[119] wl[196] vdd gnd cell_6t
Xbit_r197_c119 bl[119] br[119] wl[197] vdd gnd cell_6t
Xbit_r198_c119 bl[119] br[119] wl[198] vdd gnd cell_6t
Xbit_r199_c119 bl[119] br[119] wl[199] vdd gnd cell_6t
Xbit_r200_c119 bl[119] br[119] wl[200] vdd gnd cell_6t
Xbit_r201_c119 bl[119] br[119] wl[201] vdd gnd cell_6t
Xbit_r202_c119 bl[119] br[119] wl[202] vdd gnd cell_6t
Xbit_r203_c119 bl[119] br[119] wl[203] vdd gnd cell_6t
Xbit_r204_c119 bl[119] br[119] wl[204] vdd gnd cell_6t
Xbit_r205_c119 bl[119] br[119] wl[205] vdd gnd cell_6t
Xbit_r206_c119 bl[119] br[119] wl[206] vdd gnd cell_6t
Xbit_r207_c119 bl[119] br[119] wl[207] vdd gnd cell_6t
Xbit_r208_c119 bl[119] br[119] wl[208] vdd gnd cell_6t
Xbit_r209_c119 bl[119] br[119] wl[209] vdd gnd cell_6t
Xbit_r210_c119 bl[119] br[119] wl[210] vdd gnd cell_6t
Xbit_r211_c119 bl[119] br[119] wl[211] vdd gnd cell_6t
Xbit_r212_c119 bl[119] br[119] wl[212] vdd gnd cell_6t
Xbit_r213_c119 bl[119] br[119] wl[213] vdd gnd cell_6t
Xbit_r214_c119 bl[119] br[119] wl[214] vdd gnd cell_6t
Xbit_r215_c119 bl[119] br[119] wl[215] vdd gnd cell_6t
Xbit_r216_c119 bl[119] br[119] wl[216] vdd gnd cell_6t
Xbit_r217_c119 bl[119] br[119] wl[217] vdd gnd cell_6t
Xbit_r218_c119 bl[119] br[119] wl[218] vdd gnd cell_6t
Xbit_r219_c119 bl[119] br[119] wl[219] vdd gnd cell_6t
Xbit_r220_c119 bl[119] br[119] wl[220] vdd gnd cell_6t
Xbit_r221_c119 bl[119] br[119] wl[221] vdd gnd cell_6t
Xbit_r222_c119 bl[119] br[119] wl[222] vdd gnd cell_6t
Xbit_r223_c119 bl[119] br[119] wl[223] vdd gnd cell_6t
Xbit_r224_c119 bl[119] br[119] wl[224] vdd gnd cell_6t
Xbit_r225_c119 bl[119] br[119] wl[225] vdd gnd cell_6t
Xbit_r226_c119 bl[119] br[119] wl[226] vdd gnd cell_6t
Xbit_r227_c119 bl[119] br[119] wl[227] vdd gnd cell_6t
Xbit_r228_c119 bl[119] br[119] wl[228] vdd gnd cell_6t
Xbit_r229_c119 bl[119] br[119] wl[229] vdd gnd cell_6t
Xbit_r230_c119 bl[119] br[119] wl[230] vdd gnd cell_6t
Xbit_r231_c119 bl[119] br[119] wl[231] vdd gnd cell_6t
Xbit_r232_c119 bl[119] br[119] wl[232] vdd gnd cell_6t
Xbit_r233_c119 bl[119] br[119] wl[233] vdd gnd cell_6t
Xbit_r234_c119 bl[119] br[119] wl[234] vdd gnd cell_6t
Xbit_r235_c119 bl[119] br[119] wl[235] vdd gnd cell_6t
Xbit_r236_c119 bl[119] br[119] wl[236] vdd gnd cell_6t
Xbit_r237_c119 bl[119] br[119] wl[237] vdd gnd cell_6t
Xbit_r238_c119 bl[119] br[119] wl[238] vdd gnd cell_6t
Xbit_r239_c119 bl[119] br[119] wl[239] vdd gnd cell_6t
Xbit_r240_c119 bl[119] br[119] wl[240] vdd gnd cell_6t
Xbit_r241_c119 bl[119] br[119] wl[241] vdd gnd cell_6t
Xbit_r242_c119 bl[119] br[119] wl[242] vdd gnd cell_6t
Xbit_r243_c119 bl[119] br[119] wl[243] vdd gnd cell_6t
Xbit_r244_c119 bl[119] br[119] wl[244] vdd gnd cell_6t
Xbit_r245_c119 bl[119] br[119] wl[245] vdd gnd cell_6t
Xbit_r246_c119 bl[119] br[119] wl[246] vdd gnd cell_6t
Xbit_r247_c119 bl[119] br[119] wl[247] vdd gnd cell_6t
Xbit_r248_c119 bl[119] br[119] wl[248] vdd gnd cell_6t
Xbit_r249_c119 bl[119] br[119] wl[249] vdd gnd cell_6t
Xbit_r250_c119 bl[119] br[119] wl[250] vdd gnd cell_6t
Xbit_r251_c119 bl[119] br[119] wl[251] vdd gnd cell_6t
Xbit_r252_c119 bl[119] br[119] wl[252] vdd gnd cell_6t
Xbit_r253_c119 bl[119] br[119] wl[253] vdd gnd cell_6t
Xbit_r254_c119 bl[119] br[119] wl[254] vdd gnd cell_6t
Xbit_r255_c119 bl[119] br[119] wl[255] vdd gnd cell_6t
Xbit_r0_c120 bl[120] br[120] wl[0] vdd gnd cell_6t
Xbit_r1_c120 bl[120] br[120] wl[1] vdd gnd cell_6t
Xbit_r2_c120 bl[120] br[120] wl[2] vdd gnd cell_6t
Xbit_r3_c120 bl[120] br[120] wl[3] vdd gnd cell_6t
Xbit_r4_c120 bl[120] br[120] wl[4] vdd gnd cell_6t
Xbit_r5_c120 bl[120] br[120] wl[5] vdd gnd cell_6t
Xbit_r6_c120 bl[120] br[120] wl[6] vdd gnd cell_6t
Xbit_r7_c120 bl[120] br[120] wl[7] vdd gnd cell_6t
Xbit_r8_c120 bl[120] br[120] wl[8] vdd gnd cell_6t
Xbit_r9_c120 bl[120] br[120] wl[9] vdd gnd cell_6t
Xbit_r10_c120 bl[120] br[120] wl[10] vdd gnd cell_6t
Xbit_r11_c120 bl[120] br[120] wl[11] vdd gnd cell_6t
Xbit_r12_c120 bl[120] br[120] wl[12] vdd gnd cell_6t
Xbit_r13_c120 bl[120] br[120] wl[13] vdd gnd cell_6t
Xbit_r14_c120 bl[120] br[120] wl[14] vdd gnd cell_6t
Xbit_r15_c120 bl[120] br[120] wl[15] vdd gnd cell_6t
Xbit_r16_c120 bl[120] br[120] wl[16] vdd gnd cell_6t
Xbit_r17_c120 bl[120] br[120] wl[17] vdd gnd cell_6t
Xbit_r18_c120 bl[120] br[120] wl[18] vdd gnd cell_6t
Xbit_r19_c120 bl[120] br[120] wl[19] vdd gnd cell_6t
Xbit_r20_c120 bl[120] br[120] wl[20] vdd gnd cell_6t
Xbit_r21_c120 bl[120] br[120] wl[21] vdd gnd cell_6t
Xbit_r22_c120 bl[120] br[120] wl[22] vdd gnd cell_6t
Xbit_r23_c120 bl[120] br[120] wl[23] vdd gnd cell_6t
Xbit_r24_c120 bl[120] br[120] wl[24] vdd gnd cell_6t
Xbit_r25_c120 bl[120] br[120] wl[25] vdd gnd cell_6t
Xbit_r26_c120 bl[120] br[120] wl[26] vdd gnd cell_6t
Xbit_r27_c120 bl[120] br[120] wl[27] vdd gnd cell_6t
Xbit_r28_c120 bl[120] br[120] wl[28] vdd gnd cell_6t
Xbit_r29_c120 bl[120] br[120] wl[29] vdd gnd cell_6t
Xbit_r30_c120 bl[120] br[120] wl[30] vdd gnd cell_6t
Xbit_r31_c120 bl[120] br[120] wl[31] vdd gnd cell_6t
Xbit_r32_c120 bl[120] br[120] wl[32] vdd gnd cell_6t
Xbit_r33_c120 bl[120] br[120] wl[33] vdd gnd cell_6t
Xbit_r34_c120 bl[120] br[120] wl[34] vdd gnd cell_6t
Xbit_r35_c120 bl[120] br[120] wl[35] vdd gnd cell_6t
Xbit_r36_c120 bl[120] br[120] wl[36] vdd gnd cell_6t
Xbit_r37_c120 bl[120] br[120] wl[37] vdd gnd cell_6t
Xbit_r38_c120 bl[120] br[120] wl[38] vdd gnd cell_6t
Xbit_r39_c120 bl[120] br[120] wl[39] vdd gnd cell_6t
Xbit_r40_c120 bl[120] br[120] wl[40] vdd gnd cell_6t
Xbit_r41_c120 bl[120] br[120] wl[41] vdd gnd cell_6t
Xbit_r42_c120 bl[120] br[120] wl[42] vdd gnd cell_6t
Xbit_r43_c120 bl[120] br[120] wl[43] vdd gnd cell_6t
Xbit_r44_c120 bl[120] br[120] wl[44] vdd gnd cell_6t
Xbit_r45_c120 bl[120] br[120] wl[45] vdd gnd cell_6t
Xbit_r46_c120 bl[120] br[120] wl[46] vdd gnd cell_6t
Xbit_r47_c120 bl[120] br[120] wl[47] vdd gnd cell_6t
Xbit_r48_c120 bl[120] br[120] wl[48] vdd gnd cell_6t
Xbit_r49_c120 bl[120] br[120] wl[49] vdd gnd cell_6t
Xbit_r50_c120 bl[120] br[120] wl[50] vdd gnd cell_6t
Xbit_r51_c120 bl[120] br[120] wl[51] vdd gnd cell_6t
Xbit_r52_c120 bl[120] br[120] wl[52] vdd gnd cell_6t
Xbit_r53_c120 bl[120] br[120] wl[53] vdd gnd cell_6t
Xbit_r54_c120 bl[120] br[120] wl[54] vdd gnd cell_6t
Xbit_r55_c120 bl[120] br[120] wl[55] vdd gnd cell_6t
Xbit_r56_c120 bl[120] br[120] wl[56] vdd gnd cell_6t
Xbit_r57_c120 bl[120] br[120] wl[57] vdd gnd cell_6t
Xbit_r58_c120 bl[120] br[120] wl[58] vdd gnd cell_6t
Xbit_r59_c120 bl[120] br[120] wl[59] vdd gnd cell_6t
Xbit_r60_c120 bl[120] br[120] wl[60] vdd gnd cell_6t
Xbit_r61_c120 bl[120] br[120] wl[61] vdd gnd cell_6t
Xbit_r62_c120 bl[120] br[120] wl[62] vdd gnd cell_6t
Xbit_r63_c120 bl[120] br[120] wl[63] vdd gnd cell_6t
Xbit_r64_c120 bl[120] br[120] wl[64] vdd gnd cell_6t
Xbit_r65_c120 bl[120] br[120] wl[65] vdd gnd cell_6t
Xbit_r66_c120 bl[120] br[120] wl[66] vdd gnd cell_6t
Xbit_r67_c120 bl[120] br[120] wl[67] vdd gnd cell_6t
Xbit_r68_c120 bl[120] br[120] wl[68] vdd gnd cell_6t
Xbit_r69_c120 bl[120] br[120] wl[69] vdd gnd cell_6t
Xbit_r70_c120 bl[120] br[120] wl[70] vdd gnd cell_6t
Xbit_r71_c120 bl[120] br[120] wl[71] vdd gnd cell_6t
Xbit_r72_c120 bl[120] br[120] wl[72] vdd gnd cell_6t
Xbit_r73_c120 bl[120] br[120] wl[73] vdd gnd cell_6t
Xbit_r74_c120 bl[120] br[120] wl[74] vdd gnd cell_6t
Xbit_r75_c120 bl[120] br[120] wl[75] vdd gnd cell_6t
Xbit_r76_c120 bl[120] br[120] wl[76] vdd gnd cell_6t
Xbit_r77_c120 bl[120] br[120] wl[77] vdd gnd cell_6t
Xbit_r78_c120 bl[120] br[120] wl[78] vdd gnd cell_6t
Xbit_r79_c120 bl[120] br[120] wl[79] vdd gnd cell_6t
Xbit_r80_c120 bl[120] br[120] wl[80] vdd gnd cell_6t
Xbit_r81_c120 bl[120] br[120] wl[81] vdd gnd cell_6t
Xbit_r82_c120 bl[120] br[120] wl[82] vdd gnd cell_6t
Xbit_r83_c120 bl[120] br[120] wl[83] vdd gnd cell_6t
Xbit_r84_c120 bl[120] br[120] wl[84] vdd gnd cell_6t
Xbit_r85_c120 bl[120] br[120] wl[85] vdd gnd cell_6t
Xbit_r86_c120 bl[120] br[120] wl[86] vdd gnd cell_6t
Xbit_r87_c120 bl[120] br[120] wl[87] vdd gnd cell_6t
Xbit_r88_c120 bl[120] br[120] wl[88] vdd gnd cell_6t
Xbit_r89_c120 bl[120] br[120] wl[89] vdd gnd cell_6t
Xbit_r90_c120 bl[120] br[120] wl[90] vdd gnd cell_6t
Xbit_r91_c120 bl[120] br[120] wl[91] vdd gnd cell_6t
Xbit_r92_c120 bl[120] br[120] wl[92] vdd gnd cell_6t
Xbit_r93_c120 bl[120] br[120] wl[93] vdd gnd cell_6t
Xbit_r94_c120 bl[120] br[120] wl[94] vdd gnd cell_6t
Xbit_r95_c120 bl[120] br[120] wl[95] vdd gnd cell_6t
Xbit_r96_c120 bl[120] br[120] wl[96] vdd gnd cell_6t
Xbit_r97_c120 bl[120] br[120] wl[97] vdd gnd cell_6t
Xbit_r98_c120 bl[120] br[120] wl[98] vdd gnd cell_6t
Xbit_r99_c120 bl[120] br[120] wl[99] vdd gnd cell_6t
Xbit_r100_c120 bl[120] br[120] wl[100] vdd gnd cell_6t
Xbit_r101_c120 bl[120] br[120] wl[101] vdd gnd cell_6t
Xbit_r102_c120 bl[120] br[120] wl[102] vdd gnd cell_6t
Xbit_r103_c120 bl[120] br[120] wl[103] vdd gnd cell_6t
Xbit_r104_c120 bl[120] br[120] wl[104] vdd gnd cell_6t
Xbit_r105_c120 bl[120] br[120] wl[105] vdd gnd cell_6t
Xbit_r106_c120 bl[120] br[120] wl[106] vdd gnd cell_6t
Xbit_r107_c120 bl[120] br[120] wl[107] vdd gnd cell_6t
Xbit_r108_c120 bl[120] br[120] wl[108] vdd gnd cell_6t
Xbit_r109_c120 bl[120] br[120] wl[109] vdd gnd cell_6t
Xbit_r110_c120 bl[120] br[120] wl[110] vdd gnd cell_6t
Xbit_r111_c120 bl[120] br[120] wl[111] vdd gnd cell_6t
Xbit_r112_c120 bl[120] br[120] wl[112] vdd gnd cell_6t
Xbit_r113_c120 bl[120] br[120] wl[113] vdd gnd cell_6t
Xbit_r114_c120 bl[120] br[120] wl[114] vdd gnd cell_6t
Xbit_r115_c120 bl[120] br[120] wl[115] vdd gnd cell_6t
Xbit_r116_c120 bl[120] br[120] wl[116] vdd gnd cell_6t
Xbit_r117_c120 bl[120] br[120] wl[117] vdd gnd cell_6t
Xbit_r118_c120 bl[120] br[120] wl[118] vdd gnd cell_6t
Xbit_r119_c120 bl[120] br[120] wl[119] vdd gnd cell_6t
Xbit_r120_c120 bl[120] br[120] wl[120] vdd gnd cell_6t
Xbit_r121_c120 bl[120] br[120] wl[121] vdd gnd cell_6t
Xbit_r122_c120 bl[120] br[120] wl[122] vdd gnd cell_6t
Xbit_r123_c120 bl[120] br[120] wl[123] vdd gnd cell_6t
Xbit_r124_c120 bl[120] br[120] wl[124] vdd gnd cell_6t
Xbit_r125_c120 bl[120] br[120] wl[125] vdd gnd cell_6t
Xbit_r126_c120 bl[120] br[120] wl[126] vdd gnd cell_6t
Xbit_r127_c120 bl[120] br[120] wl[127] vdd gnd cell_6t
Xbit_r128_c120 bl[120] br[120] wl[128] vdd gnd cell_6t
Xbit_r129_c120 bl[120] br[120] wl[129] vdd gnd cell_6t
Xbit_r130_c120 bl[120] br[120] wl[130] vdd gnd cell_6t
Xbit_r131_c120 bl[120] br[120] wl[131] vdd gnd cell_6t
Xbit_r132_c120 bl[120] br[120] wl[132] vdd gnd cell_6t
Xbit_r133_c120 bl[120] br[120] wl[133] vdd gnd cell_6t
Xbit_r134_c120 bl[120] br[120] wl[134] vdd gnd cell_6t
Xbit_r135_c120 bl[120] br[120] wl[135] vdd gnd cell_6t
Xbit_r136_c120 bl[120] br[120] wl[136] vdd gnd cell_6t
Xbit_r137_c120 bl[120] br[120] wl[137] vdd gnd cell_6t
Xbit_r138_c120 bl[120] br[120] wl[138] vdd gnd cell_6t
Xbit_r139_c120 bl[120] br[120] wl[139] vdd gnd cell_6t
Xbit_r140_c120 bl[120] br[120] wl[140] vdd gnd cell_6t
Xbit_r141_c120 bl[120] br[120] wl[141] vdd gnd cell_6t
Xbit_r142_c120 bl[120] br[120] wl[142] vdd gnd cell_6t
Xbit_r143_c120 bl[120] br[120] wl[143] vdd gnd cell_6t
Xbit_r144_c120 bl[120] br[120] wl[144] vdd gnd cell_6t
Xbit_r145_c120 bl[120] br[120] wl[145] vdd gnd cell_6t
Xbit_r146_c120 bl[120] br[120] wl[146] vdd gnd cell_6t
Xbit_r147_c120 bl[120] br[120] wl[147] vdd gnd cell_6t
Xbit_r148_c120 bl[120] br[120] wl[148] vdd gnd cell_6t
Xbit_r149_c120 bl[120] br[120] wl[149] vdd gnd cell_6t
Xbit_r150_c120 bl[120] br[120] wl[150] vdd gnd cell_6t
Xbit_r151_c120 bl[120] br[120] wl[151] vdd gnd cell_6t
Xbit_r152_c120 bl[120] br[120] wl[152] vdd gnd cell_6t
Xbit_r153_c120 bl[120] br[120] wl[153] vdd gnd cell_6t
Xbit_r154_c120 bl[120] br[120] wl[154] vdd gnd cell_6t
Xbit_r155_c120 bl[120] br[120] wl[155] vdd gnd cell_6t
Xbit_r156_c120 bl[120] br[120] wl[156] vdd gnd cell_6t
Xbit_r157_c120 bl[120] br[120] wl[157] vdd gnd cell_6t
Xbit_r158_c120 bl[120] br[120] wl[158] vdd gnd cell_6t
Xbit_r159_c120 bl[120] br[120] wl[159] vdd gnd cell_6t
Xbit_r160_c120 bl[120] br[120] wl[160] vdd gnd cell_6t
Xbit_r161_c120 bl[120] br[120] wl[161] vdd gnd cell_6t
Xbit_r162_c120 bl[120] br[120] wl[162] vdd gnd cell_6t
Xbit_r163_c120 bl[120] br[120] wl[163] vdd gnd cell_6t
Xbit_r164_c120 bl[120] br[120] wl[164] vdd gnd cell_6t
Xbit_r165_c120 bl[120] br[120] wl[165] vdd gnd cell_6t
Xbit_r166_c120 bl[120] br[120] wl[166] vdd gnd cell_6t
Xbit_r167_c120 bl[120] br[120] wl[167] vdd gnd cell_6t
Xbit_r168_c120 bl[120] br[120] wl[168] vdd gnd cell_6t
Xbit_r169_c120 bl[120] br[120] wl[169] vdd gnd cell_6t
Xbit_r170_c120 bl[120] br[120] wl[170] vdd gnd cell_6t
Xbit_r171_c120 bl[120] br[120] wl[171] vdd gnd cell_6t
Xbit_r172_c120 bl[120] br[120] wl[172] vdd gnd cell_6t
Xbit_r173_c120 bl[120] br[120] wl[173] vdd gnd cell_6t
Xbit_r174_c120 bl[120] br[120] wl[174] vdd gnd cell_6t
Xbit_r175_c120 bl[120] br[120] wl[175] vdd gnd cell_6t
Xbit_r176_c120 bl[120] br[120] wl[176] vdd gnd cell_6t
Xbit_r177_c120 bl[120] br[120] wl[177] vdd gnd cell_6t
Xbit_r178_c120 bl[120] br[120] wl[178] vdd gnd cell_6t
Xbit_r179_c120 bl[120] br[120] wl[179] vdd gnd cell_6t
Xbit_r180_c120 bl[120] br[120] wl[180] vdd gnd cell_6t
Xbit_r181_c120 bl[120] br[120] wl[181] vdd gnd cell_6t
Xbit_r182_c120 bl[120] br[120] wl[182] vdd gnd cell_6t
Xbit_r183_c120 bl[120] br[120] wl[183] vdd gnd cell_6t
Xbit_r184_c120 bl[120] br[120] wl[184] vdd gnd cell_6t
Xbit_r185_c120 bl[120] br[120] wl[185] vdd gnd cell_6t
Xbit_r186_c120 bl[120] br[120] wl[186] vdd gnd cell_6t
Xbit_r187_c120 bl[120] br[120] wl[187] vdd gnd cell_6t
Xbit_r188_c120 bl[120] br[120] wl[188] vdd gnd cell_6t
Xbit_r189_c120 bl[120] br[120] wl[189] vdd gnd cell_6t
Xbit_r190_c120 bl[120] br[120] wl[190] vdd gnd cell_6t
Xbit_r191_c120 bl[120] br[120] wl[191] vdd gnd cell_6t
Xbit_r192_c120 bl[120] br[120] wl[192] vdd gnd cell_6t
Xbit_r193_c120 bl[120] br[120] wl[193] vdd gnd cell_6t
Xbit_r194_c120 bl[120] br[120] wl[194] vdd gnd cell_6t
Xbit_r195_c120 bl[120] br[120] wl[195] vdd gnd cell_6t
Xbit_r196_c120 bl[120] br[120] wl[196] vdd gnd cell_6t
Xbit_r197_c120 bl[120] br[120] wl[197] vdd gnd cell_6t
Xbit_r198_c120 bl[120] br[120] wl[198] vdd gnd cell_6t
Xbit_r199_c120 bl[120] br[120] wl[199] vdd gnd cell_6t
Xbit_r200_c120 bl[120] br[120] wl[200] vdd gnd cell_6t
Xbit_r201_c120 bl[120] br[120] wl[201] vdd gnd cell_6t
Xbit_r202_c120 bl[120] br[120] wl[202] vdd gnd cell_6t
Xbit_r203_c120 bl[120] br[120] wl[203] vdd gnd cell_6t
Xbit_r204_c120 bl[120] br[120] wl[204] vdd gnd cell_6t
Xbit_r205_c120 bl[120] br[120] wl[205] vdd gnd cell_6t
Xbit_r206_c120 bl[120] br[120] wl[206] vdd gnd cell_6t
Xbit_r207_c120 bl[120] br[120] wl[207] vdd gnd cell_6t
Xbit_r208_c120 bl[120] br[120] wl[208] vdd gnd cell_6t
Xbit_r209_c120 bl[120] br[120] wl[209] vdd gnd cell_6t
Xbit_r210_c120 bl[120] br[120] wl[210] vdd gnd cell_6t
Xbit_r211_c120 bl[120] br[120] wl[211] vdd gnd cell_6t
Xbit_r212_c120 bl[120] br[120] wl[212] vdd gnd cell_6t
Xbit_r213_c120 bl[120] br[120] wl[213] vdd gnd cell_6t
Xbit_r214_c120 bl[120] br[120] wl[214] vdd gnd cell_6t
Xbit_r215_c120 bl[120] br[120] wl[215] vdd gnd cell_6t
Xbit_r216_c120 bl[120] br[120] wl[216] vdd gnd cell_6t
Xbit_r217_c120 bl[120] br[120] wl[217] vdd gnd cell_6t
Xbit_r218_c120 bl[120] br[120] wl[218] vdd gnd cell_6t
Xbit_r219_c120 bl[120] br[120] wl[219] vdd gnd cell_6t
Xbit_r220_c120 bl[120] br[120] wl[220] vdd gnd cell_6t
Xbit_r221_c120 bl[120] br[120] wl[221] vdd gnd cell_6t
Xbit_r222_c120 bl[120] br[120] wl[222] vdd gnd cell_6t
Xbit_r223_c120 bl[120] br[120] wl[223] vdd gnd cell_6t
Xbit_r224_c120 bl[120] br[120] wl[224] vdd gnd cell_6t
Xbit_r225_c120 bl[120] br[120] wl[225] vdd gnd cell_6t
Xbit_r226_c120 bl[120] br[120] wl[226] vdd gnd cell_6t
Xbit_r227_c120 bl[120] br[120] wl[227] vdd gnd cell_6t
Xbit_r228_c120 bl[120] br[120] wl[228] vdd gnd cell_6t
Xbit_r229_c120 bl[120] br[120] wl[229] vdd gnd cell_6t
Xbit_r230_c120 bl[120] br[120] wl[230] vdd gnd cell_6t
Xbit_r231_c120 bl[120] br[120] wl[231] vdd gnd cell_6t
Xbit_r232_c120 bl[120] br[120] wl[232] vdd gnd cell_6t
Xbit_r233_c120 bl[120] br[120] wl[233] vdd gnd cell_6t
Xbit_r234_c120 bl[120] br[120] wl[234] vdd gnd cell_6t
Xbit_r235_c120 bl[120] br[120] wl[235] vdd gnd cell_6t
Xbit_r236_c120 bl[120] br[120] wl[236] vdd gnd cell_6t
Xbit_r237_c120 bl[120] br[120] wl[237] vdd gnd cell_6t
Xbit_r238_c120 bl[120] br[120] wl[238] vdd gnd cell_6t
Xbit_r239_c120 bl[120] br[120] wl[239] vdd gnd cell_6t
Xbit_r240_c120 bl[120] br[120] wl[240] vdd gnd cell_6t
Xbit_r241_c120 bl[120] br[120] wl[241] vdd gnd cell_6t
Xbit_r242_c120 bl[120] br[120] wl[242] vdd gnd cell_6t
Xbit_r243_c120 bl[120] br[120] wl[243] vdd gnd cell_6t
Xbit_r244_c120 bl[120] br[120] wl[244] vdd gnd cell_6t
Xbit_r245_c120 bl[120] br[120] wl[245] vdd gnd cell_6t
Xbit_r246_c120 bl[120] br[120] wl[246] vdd gnd cell_6t
Xbit_r247_c120 bl[120] br[120] wl[247] vdd gnd cell_6t
Xbit_r248_c120 bl[120] br[120] wl[248] vdd gnd cell_6t
Xbit_r249_c120 bl[120] br[120] wl[249] vdd gnd cell_6t
Xbit_r250_c120 bl[120] br[120] wl[250] vdd gnd cell_6t
Xbit_r251_c120 bl[120] br[120] wl[251] vdd gnd cell_6t
Xbit_r252_c120 bl[120] br[120] wl[252] vdd gnd cell_6t
Xbit_r253_c120 bl[120] br[120] wl[253] vdd gnd cell_6t
Xbit_r254_c120 bl[120] br[120] wl[254] vdd gnd cell_6t
Xbit_r255_c120 bl[120] br[120] wl[255] vdd gnd cell_6t
Xbit_r0_c121 bl[121] br[121] wl[0] vdd gnd cell_6t
Xbit_r1_c121 bl[121] br[121] wl[1] vdd gnd cell_6t
Xbit_r2_c121 bl[121] br[121] wl[2] vdd gnd cell_6t
Xbit_r3_c121 bl[121] br[121] wl[3] vdd gnd cell_6t
Xbit_r4_c121 bl[121] br[121] wl[4] vdd gnd cell_6t
Xbit_r5_c121 bl[121] br[121] wl[5] vdd gnd cell_6t
Xbit_r6_c121 bl[121] br[121] wl[6] vdd gnd cell_6t
Xbit_r7_c121 bl[121] br[121] wl[7] vdd gnd cell_6t
Xbit_r8_c121 bl[121] br[121] wl[8] vdd gnd cell_6t
Xbit_r9_c121 bl[121] br[121] wl[9] vdd gnd cell_6t
Xbit_r10_c121 bl[121] br[121] wl[10] vdd gnd cell_6t
Xbit_r11_c121 bl[121] br[121] wl[11] vdd gnd cell_6t
Xbit_r12_c121 bl[121] br[121] wl[12] vdd gnd cell_6t
Xbit_r13_c121 bl[121] br[121] wl[13] vdd gnd cell_6t
Xbit_r14_c121 bl[121] br[121] wl[14] vdd gnd cell_6t
Xbit_r15_c121 bl[121] br[121] wl[15] vdd gnd cell_6t
Xbit_r16_c121 bl[121] br[121] wl[16] vdd gnd cell_6t
Xbit_r17_c121 bl[121] br[121] wl[17] vdd gnd cell_6t
Xbit_r18_c121 bl[121] br[121] wl[18] vdd gnd cell_6t
Xbit_r19_c121 bl[121] br[121] wl[19] vdd gnd cell_6t
Xbit_r20_c121 bl[121] br[121] wl[20] vdd gnd cell_6t
Xbit_r21_c121 bl[121] br[121] wl[21] vdd gnd cell_6t
Xbit_r22_c121 bl[121] br[121] wl[22] vdd gnd cell_6t
Xbit_r23_c121 bl[121] br[121] wl[23] vdd gnd cell_6t
Xbit_r24_c121 bl[121] br[121] wl[24] vdd gnd cell_6t
Xbit_r25_c121 bl[121] br[121] wl[25] vdd gnd cell_6t
Xbit_r26_c121 bl[121] br[121] wl[26] vdd gnd cell_6t
Xbit_r27_c121 bl[121] br[121] wl[27] vdd gnd cell_6t
Xbit_r28_c121 bl[121] br[121] wl[28] vdd gnd cell_6t
Xbit_r29_c121 bl[121] br[121] wl[29] vdd gnd cell_6t
Xbit_r30_c121 bl[121] br[121] wl[30] vdd gnd cell_6t
Xbit_r31_c121 bl[121] br[121] wl[31] vdd gnd cell_6t
Xbit_r32_c121 bl[121] br[121] wl[32] vdd gnd cell_6t
Xbit_r33_c121 bl[121] br[121] wl[33] vdd gnd cell_6t
Xbit_r34_c121 bl[121] br[121] wl[34] vdd gnd cell_6t
Xbit_r35_c121 bl[121] br[121] wl[35] vdd gnd cell_6t
Xbit_r36_c121 bl[121] br[121] wl[36] vdd gnd cell_6t
Xbit_r37_c121 bl[121] br[121] wl[37] vdd gnd cell_6t
Xbit_r38_c121 bl[121] br[121] wl[38] vdd gnd cell_6t
Xbit_r39_c121 bl[121] br[121] wl[39] vdd gnd cell_6t
Xbit_r40_c121 bl[121] br[121] wl[40] vdd gnd cell_6t
Xbit_r41_c121 bl[121] br[121] wl[41] vdd gnd cell_6t
Xbit_r42_c121 bl[121] br[121] wl[42] vdd gnd cell_6t
Xbit_r43_c121 bl[121] br[121] wl[43] vdd gnd cell_6t
Xbit_r44_c121 bl[121] br[121] wl[44] vdd gnd cell_6t
Xbit_r45_c121 bl[121] br[121] wl[45] vdd gnd cell_6t
Xbit_r46_c121 bl[121] br[121] wl[46] vdd gnd cell_6t
Xbit_r47_c121 bl[121] br[121] wl[47] vdd gnd cell_6t
Xbit_r48_c121 bl[121] br[121] wl[48] vdd gnd cell_6t
Xbit_r49_c121 bl[121] br[121] wl[49] vdd gnd cell_6t
Xbit_r50_c121 bl[121] br[121] wl[50] vdd gnd cell_6t
Xbit_r51_c121 bl[121] br[121] wl[51] vdd gnd cell_6t
Xbit_r52_c121 bl[121] br[121] wl[52] vdd gnd cell_6t
Xbit_r53_c121 bl[121] br[121] wl[53] vdd gnd cell_6t
Xbit_r54_c121 bl[121] br[121] wl[54] vdd gnd cell_6t
Xbit_r55_c121 bl[121] br[121] wl[55] vdd gnd cell_6t
Xbit_r56_c121 bl[121] br[121] wl[56] vdd gnd cell_6t
Xbit_r57_c121 bl[121] br[121] wl[57] vdd gnd cell_6t
Xbit_r58_c121 bl[121] br[121] wl[58] vdd gnd cell_6t
Xbit_r59_c121 bl[121] br[121] wl[59] vdd gnd cell_6t
Xbit_r60_c121 bl[121] br[121] wl[60] vdd gnd cell_6t
Xbit_r61_c121 bl[121] br[121] wl[61] vdd gnd cell_6t
Xbit_r62_c121 bl[121] br[121] wl[62] vdd gnd cell_6t
Xbit_r63_c121 bl[121] br[121] wl[63] vdd gnd cell_6t
Xbit_r64_c121 bl[121] br[121] wl[64] vdd gnd cell_6t
Xbit_r65_c121 bl[121] br[121] wl[65] vdd gnd cell_6t
Xbit_r66_c121 bl[121] br[121] wl[66] vdd gnd cell_6t
Xbit_r67_c121 bl[121] br[121] wl[67] vdd gnd cell_6t
Xbit_r68_c121 bl[121] br[121] wl[68] vdd gnd cell_6t
Xbit_r69_c121 bl[121] br[121] wl[69] vdd gnd cell_6t
Xbit_r70_c121 bl[121] br[121] wl[70] vdd gnd cell_6t
Xbit_r71_c121 bl[121] br[121] wl[71] vdd gnd cell_6t
Xbit_r72_c121 bl[121] br[121] wl[72] vdd gnd cell_6t
Xbit_r73_c121 bl[121] br[121] wl[73] vdd gnd cell_6t
Xbit_r74_c121 bl[121] br[121] wl[74] vdd gnd cell_6t
Xbit_r75_c121 bl[121] br[121] wl[75] vdd gnd cell_6t
Xbit_r76_c121 bl[121] br[121] wl[76] vdd gnd cell_6t
Xbit_r77_c121 bl[121] br[121] wl[77] vdd gnd cell_6t
Xbit_r78_c121 bl[121] br[121] wl[78] vdd gnd cell_6t
Xbit_r79_c121 bl[121] br[121] wl[79] vdd gnd cell_6t
Xbit_r80_c121 bl[121] br[121] wl[80] vdd gnd cell_6t
Xbit_r81_c121 bl[121] br[121] wl[81] vdd gnd cell_6t
Xbit_r82_c121 bl[121] br[121] wl[82] vdd gnd cell_6t
Xbit_r83_c121 bl[121] br[121] wl[83] vdd gnd cell_6t
Xbit_r84_c121 bl[121] br[121] wl[84] vdd gnd cell_6t
Xbit_r85_c121 bl[121] br[121] wl[85] vdd gnd cell_6t
Xbit_r86_c121 bl[121] br[121] wl[86] vdd gnd cell_6t
Xbit_r87_c121 bl[121] br[121] wl[87] vdd gnd cell_6t
Xbit_r88_c121 bl[121] br[121] wl[88] vdd gnd cell_6t
Xbit_r89_c121 bl[121] br[121] wl[89] vdd gnd cell_6t
Xbit_r90_c121 bl[121] br[121] wl[90] vdd gnd cell_6t
Xbit_r91_c121 bl[121] br[121] wl[91] vdd gnd cell_6t
Xbit_r92_c121 bl[121] br[121] wl[92] vdd gnd cell_6t
Xbit_r93_c121 bl[121] br[121] wl[93] vdd gnd cell_6t
Xbit_r94_c121 bl[121] br[121] wl[94] vdd gnd cell_6t
Xbit_r95_c121 bl[121] br[121] wl[95] vdd gnd cell_6t
Xbit_r96_c121 bl[121] br[121] wl[96] vdd gnd cell_6t
Xbit_r97_c121 bl[121] br[121] wl[97] vdd gnd cell_6t
Xbit_r98_c121 bl[121] br[121] wl[98] vdd gnd cell_6t
Xbit_r99_c121 bl[121] br[121] wl[99] vdd gnd cell_6t
Xbit_r100_c121 bl[121] br[121] wl[100] vdd gnd cell_6t
Xbit_r101_c121 bl[121] br[121] wl[101] vdd gnd cell_6t
Xbit_r102_c121 bl[121] br[121] wl[102] vdd gnd cell_6t
Xbit_r103_c121 bl[121] br[121] wl[103] vdd gnd cell_6t
Xbit_r104_c121 bl[121] br[121] wl[104] vdd gnd cell_6t
Xbit_r105_c121 bl[121] br[121] wl[105] vdd gnd cell_6t
Xbit_r106_c121 bl[121] br[121] wl[106] vdd gnd cell_6t
Xbit_r107_c121 bl[121] br[121] wl[107] vdd gnd cell_6t
Xbit_r108_c121 bl[121] br[121] wl[108] vdd gnd cell_6t
Xbit_r109_c121 bl[121] br[121] wl[109] vdd gnd cell_6t
Xbit_r110_c121 bl[121] br[121] wl[110] vdd gnd cell_6t
Xbit_r111_c121 bl[121] br[121] wl[111] vdd gnd cell_6t
Xbit_r112_c121 bl[121] br[121] wl[112] vdd gnd cell_6t
Xbit_r113_c121 bl[121] br[121] wl[113] vdd gnd cell_6t
Xbit_r114_c121 bl[121] br[121] wl[114] vdd gnd cell_6t
Xbit_r115_c121 bl[121] br[121] wl[115] vdd gnd cell_6t
Xbit_r116_c121 bl[121] br[121] wl[116] vdd gnd cell_6t
Xbit_r117_c121 bl[121] br[121] wl[117] vdd gnd cell_6t
Xbit_r118_c121 bl[121] br[121] wl[118] vdd gnd cell_6t
Xbit_r119_c121 bl[121] br[121] wl[119] vdd gnd cell_6t
Xbit_r120_c121 bl[121] br[121] wl[120] vdd gnd cell_6t
Xbit_r121_c121 bl[121] br[121] wl[121] vdd gnd cell_6t
Xbit_r122_c121 bl[121] br[121] wl[122] vdd gnd cell_6t
Xbit_r123_c121 bl[121] br[121] wl[123] vdd gnd cell_6t
Xbit_r124_c121 bl[121] br[121] wl[124] vdd gnd cell_6t
Xbit_r125_c121 bl[121] br[121] wl[125] vdd gnd cell_6t
Xbit_r126_c121 bl[121] br[121] wl[126] vdd gnd cell_6t
Xbit_r127_c121 bl[121] br[121] wl[127] vdd gnd cell_6t
Xbit_r128_c121 bl[121] br[121] wl[128] vdd gnd cell_6t
Xbit_r129_c121 bl[121] br[121] wl[129] vdd gnd cell_6t
Xbit_r130_c121 bl[121] br[121] wl[130] vdd gnd cell_6t
Xbit_r131_c121 bl[121] br[121] wl[131] vdd gnd cell_6t
Xbit_r132_c121 bl[121] br[121] wl[132] vdd gnd cell_6t
Xbit_r133_c121 bl[121] br[121] wl[133] vdd gnd cell_6t
Xbit_r134_c121 bl[121] br[121] wl[134] vdd gnd cell_6t
Xbit_r135_c121 bl[121] br[121] wl[135] vdd gnd cell_6t
Xbit_r136_c121 bl[121] br[121] wl[136] vdd gnd cell_6t
Xbit_r137_c121 bl[121] br[121] wl[137] vdd gnd cell_6t
Xbit_r138_c121 bl[121] br[121] wl[138] vdd gnd cell_6t
Xbit_r139_c121 bl[121] br[121] wl[139] vdd gnd cell_6t
Xbit_r140_c121 bl[121] br[121] wl[140] vdd gnd cell_6t
Xbit_r141_c121 bl[121] br[121] wl[141] vdd gnd cell_6t
Xbit_r142_c121 bl[121] br[121] wl[142] vdd gnd cell_6t
Xbit_r143_c121 bl[121] br[121] wl[143] vdd gnd cell_6t
Xbit_r144_c121 bl[121] br[121] wl[144] vdd gnd cell_6t
Xbit_r145_c121 bl[121] br[121] wl[145] vdd gnd cell_6t
Xbit_r146_c121 bl[121] br[121] wl[146] vdd gnd cell_6t
Xbit_r147_c121 bl[121] br[121] wl[147] vdd gnd cell_6t
Xbit_r148_c121 bl[121] br[121] wl[148] vdd gnd cell_6t
Xbit_r149_c121 bl[121] br[121] wl[149] vdd gnd cell_6t
Xbit_r150_c121 bl[121] br[121] wl[150] vdd gnd cell_6t
Xbit_r151_c121 bl[121] br[121] wl[151] vdd gnd cell_6t
Xbit_r152_c121 bl[121] br[121] wl[152] vdd gnd cell_6t
Xbit_r153_c121 bl[121] br[121] wl[153] vdd gnd cell_6t
Xbit_r154_c121 bl[121] br[121] wl[154] vdd gnd cell_6t
Xbit_r155_c121 bl[121] br[121] wl[155] vdd gnd cell_6t
Xbit_r156_c121 bl[121] br[121] wl[156] vdd gnd cell_6t
Xbit_r157_c121 bl[121] br[121] wl[157] vdd gnd cell_6t
Xbit_r158_c121 bl[121] br[121] wl[158] vdd gnd cell_6t
Xbit_r159_c121 bl[121] br[121] wl[159] vdd gnd cell_6t
Xbit_r160_c121 bl[121] br[121] wl[160] vdd gnd cell_6t
Xbit_r161_c121 bl[121] br[121] wl[161] vdd gnd cell_6t
Xbit_r162_c121 bl[121] br[121] wl[162] vdd gnd cell_6t
Xbit_r163_c121 bl[121] br[121] wl[163] vdd gnd cell_6t
Xbit_r164_c121 bl[121] br[121] wl[164] vdd gnd cell_6t
Xbit_r165_c121 bl[121] br[121] wl[165] vdd gnd cell_6t
Xbit_r166_c121 bl[121] br[121] wl[166] vdd gnd cell_6t
Xbit_r167_c121 bl[121] br[121] wl[167] vdd gnd cell_6t
Xbit_r168_c121 bl[121] br[121] wl[168] vdd gnd cell_6t
Xbit_r169_c121 bl[121] br[121] wl[169] vdd gnd cell_6t
Xbit_r170_c121 bl[121] br[121] wl[170] vdd gnd cell_6t
Xbit_r171_c121 bl[121] br[121] wl[171] vdd gnd cell_6t
Xbit_r172_c121 bl[121] br[121] wl[172] vdd gnd cell_6t
Xbit_r173_c121 bl[121] br[121] wl[173] vdd gnd cell_6t
Xbit_r174_c121 bl[121] br[121] wl[174] vdd gnd cell_6t
Xbit_r175_c121 bl[121] br[121] wl[175] vdd gnd cell_6t
Xbit_r176_c121 bl[121] br[121] wl[176] vdd gnd cell_6t
Xbit_r177_c121 bl[121] br[121] wl[177] vdd gnd cell_6t
Xbit_r178_c121 bl[121] br[121] wl[178] vdd gnd cell_6t
Xbit_r179_c121 bl[121] br[121] wl[179] vdd gnd cell_6t
Xbit_r180_c121 bl[121] br[121] wl[180] vdd gnd cell_6t
Xbit_r181_c121 bl[121] br[121] wl[181] vdd gnd cell_6t
Xbit_r182_c121 bl[121] br[121] wl[182] vdd gnd cell_6t
Xbit_r183_c121 bl[121] br[121] wl[183] vdd gnd cell_6t
Xbit_r184_c121 bl[121] br[121] wl[184] vdd gnd cell_6t
Xbit_r185_c121 bl[121] br[121] wl[185] vdd gnd cell_6t
Xbit_r186_c121 bl[121] br[121] wl[186] vdd gnd cell_6t
Xbit_r187_c121 bl[121] br[121] wl[187] vdd gnd cell_6t
Xbit_r188_c121 bl[121] br[121] wl[188] vdd gnd cell_6t
Xbit_r189_c121 bl[121] br[121] wl[189] vdd gnd cell_6t
Xbit_r190_c121 bl[121] br[121] wl[190] vdd gnd cell_6t
Xbit_r191_c121 bl[121] br[121] wl[191] vdd gnd cell_6t
Xbit_r192_c121 bl[121] br[121] wl[192] vdd gnd cell_6t
Xbit_r193_c121 bl[121] br[121] wl[193] vdd gnd cell_6t
Xbit_r194_c121 bl[121] br[121] wl[194] vdd gnd cell_6t
Xbit_r195_c121 bl[121] br[121] wl[195] vdd gnd cell_6t
Xbit_r196_c121 bl[121] br[121] wl[196] vdd gnd cell_6t
Xbit_r197_c121 bl[121] br[121] wl[197] vdd gnd cell_6t
Xbit_r198_c121 bl[121] br[121] wl[198] vdd gnd cell_6t
Xbit_r199_c121 bl[121] br[121] wl[199] vdd gnd cell_6t
Xbit_r200_c121 bl[121] br[121] wl[200] vdd gnd cell_6t
Xbit_r201_c121 bl[121] br[121] wl[201] vdd gnd cell_6t
Xbit_r202_c121 bl[121] br[121] wl[202] vdd gnd cell_6t
Xbit_r203_c121 bl[121] br[121] wl[203] vdd gnd cell_6t
Xbit_r204_c121 bl[121] br[121] wl[204] vdd gnd cell_6t
Xbit_r205_c121 bl[121] br[121] wl[205] vdd gnd cell_6t
Xbit_r206_c121 bl[121] br[121] wl[206] vdd gnd cell_6t
Xbit_r207_c121 bl[121] br[121] wl[207] vdd gnd cell_6t
Xbit_r208_c121 bl[121] br[121] wl[208] vdd gnd cell_6t
Xbit_r209_c121 bl[121] br[121] wl[209] vdd gnd cell_6t
Xbit_r210_c121 bl[121] br[121] wl[210] vdd gnd cell_6t
Xbit_r211_c121 bl[121] br[121] wl[211] vdd gnd cell_6t
Xbit_r212_c121 bl[121] br[121] wl[212] vdd gnd cell_6t
Xbit_r213_c121 bl[121] br[121] wl[213] vdd gnd cell_6t
Xbit_r214_c121 bl[121] br[121] wl[214] vdd gnd cell_6t
Xbit_r215_c121 bl[121] br[121] wl[215] vdd gnd cell_6t
Xbit_r216_c121 bl[121] br[121] wl[216] vdd gnd cell_6t
Xbit_r217_c121 bl[121] br[121] wl[217] vdd gnd cell_6t
Xbit_r218_c121 bl[121] br[121] wl[218] vdd gnd cell_6t
Xbit_r219_c121 bl[121] br[121] wl[219] vdd gnd cell_6t
Xbit_r220_c121 bl[121] br[121] wl[220] vdd gnd cell_6t
Xbit_r221_c121 bl[121] br[121] wl[221] vdd gnd cell_6t
Xbit_r222_c121 bl[121] br[121] wl[222] vdd gnd cell_6t
Xbit_r223_c121 bl[121] br[121] wl[223] vdd gnd cell_6t
Xbit_r224_c121 bl[121] br[121] wl[224] vdd gnd cell_6t
Xbit_r225_c121 bl[121] br[121] wl[225] vdd gnd cell_6t
Xbit_r226_c121 bl[121] br[121] wl[226] vdd gnd cell_6t
Xbit_r227_c121 bl[121] br[121] wl[227] vdd gnd cell_6t
Xbit_r228_c121 bl[121] br[121] wl[228] vdd gnd cell_6t
Xbit_r229_c121 bl[121] br[121] wl[229] vdd gnd cell_6t
Xbit_r230_c121 bl[121] br[121] wl[230] vdd gnd cell_6t
Xbit_r231_c121 bl[121] br[121] wl[231] vdd gnd cell_6t
Xbit_r232_c121 bl[121] br[121] wl[232] vdd gnd cell_6t
Xbit_r233_c121 bl[121] br[121] wl[233] vdd gnd cell_6t
Xbit_r234_c121 bl[121] br[121] wl[234] vdd gnd cell_6t
Xbit_r235_c121 bl[121] br[121] wl[235] vdd gnd cell_6t
Xbit_r236_c121 bl[121] br[121] wl[236] vdd gnd cell_6t
Xbit_r237_c121 bl[121] br[121] wl[237] vdd gnd cell_6t
Xbit_r238_c121 bl[121] br[121] wl[238] vdd gnd cell_6t
Xbit_r239_c121 bl[121] br[121] wl[239] vdd gnd cell_6t
Xbit_r240_c121 bl[121] br[121] wl[240] vdd gnd cell_6t
Xbit_r241_c121 bl[121] br[121] wl[241] vdd gnd cell_6t
Xbit_r242_c121 bl[121] br[121] wl[242] vdd gnd cell_6t
Xbit_r243_c121 bl[121] br[121] wl[243] vdd gnd cell_6t
Xbit_r244_c121 bl[121] br[121] wl[244] vdd gnd cell_6t
Xbit_r245_c121 bl[121] br[121] wl[245] vdd gnd cell_6t
Xbit_r246_c121 bl[121] br[121] wl[246] vdd gnd cell_6t
Xbit_r247_c121 bl[121] br[121] wl[247] vdd gnd cell_6t
Xbit_r248_c121 bl[121] br[121] wl[248] vdd gnd cell_6t
Xbit_r249_c121 bl[121] br[121] wl[249] vdd gnd cell_6t
Xbit_r250_c121 bl[121] br[121] wl[250] vdd gnd cell_6t
Xbit_r251_c121 bl[121] br[121] wl[251] vdd gnd cell_6t
Xbit_r252_c121 bl[121] br[121] wl[252] vdd gnd cell_6t
Xbit_r253_c121 bl[121] br[121] wl[253] vdd gnd cell_6t
Xbit_r254_c121 bl[121] br[121] wl[254] vdd gnd cell_6t
Xbit_r255_c121 bl[121] br[121] wl[255] vdd gnd cell_6t
Xbit_r0_c122 bl[122] br[122] wl[0] vdd gnd cell_6t
Xbit_r1_c122 bl[122] br[122] wl[1] vdd gnd cell_6t
Xbit_r2_c122 bl[122] br[122] wl[2] vdd gnd cell_6t
Xbit_r3_c122 bl[122] br[122] wl[3] vdd gnd cell_6t
Xbit_r4_c122 bl[122] br[122] wl[4] vdd gnd cell_6t
Xbit_r5_c122 bl[122] br[122] wl[5] vdd gnd cell_6t
Xbit_r6_c122 bl[122] br[122] wl[6] vdd gnd cell_6t
Xbit_r7_c122 bl[122] br[122] wl[7] vdd gnd cell_6t
Xbit_r8_c122 bl[122] br[122] wl[8] vdd gnd cell_6t
Xbit_r9_c122 bl[122] br[122] wl[9] vdd gnd cell_6t
Xbit_r10_c122 bl[122] br[122] wl[10] vdd gnd cell_6t
Xbit_r11_c122 bl[122] br[122] wl[11] vdd gnd cell_6t
Xbit_r12_c122 bl[122] br[122] wl[12] vdd gnd cell_6t
Xbit_r13_c122 bl[122] br[122] wl[13] vdd gnd cell_6t
Xbit_r14_c122 bl[122] br[122] wl[14] vdd gnd cell_6t
Xbit_r15_c122 bl[122] br[122] wl[15] vdd gnd cell_6t
Xbit_r16_c122 bl[122] br[122] wl[16] vdd gnd cell_6t
Xbit_r17_c122 bl[122] br[122] wl[17] vdd gnd cell_6t
Xbit_r18_c122 bl[122] br[122] wl[18] vdd gnd cell_6t
Xbit_r19_c122 bl[122] br[122] wl[19] vdd gnd cell_6t
Xbit_r20_c122 bl[122] br[122] wl[20] vdd gnd cell_6t
Xbit_r21_c122 bl[122] br[122] wl[21] vdd gnd cell_6t
Xbit_r22_c122 bl[122] br[122] wl[22] vdd gnd cell_6t
Xbit_r23_c122 bl[122] br[122] wl[23] vdd gnd cell_6t
Xbit_r24_c122 bl[122] br[122] wl[24] vdd gnd cell_6t
Xbit_r25_c122 bl[122] br[122] wl[25] vdd gnd cell_6t
Xbit_r26_c122 bl[122] br[122] wl[26] vdd gnd cell_6t
Xbit_r27_c122 bl[122] br[122] wl[27] vdd gnd cell_6t
Xbit_r28_c122 bl[122] br[122] wl[28] vdd gnd cell_6t
Xbit_r29_c122 bl[122] br[122] wl[29] vdd gnd cell_6t
Xbit_r30_c122 bl[122] br[122] wl[30] vdd gnd cell_6t
Xbit_r31_c122 bl[122] br[122] wl[31] vdd gnd cell_6t
Xbit_r32_c122 bl[122] br[122] wl[32] vdd gnd cell_6t
Xbit_r33_c122 bl[122] br[122] wl[33] vdd gnd cell_6t
Xbit_r34_c122 bl[122] br[122] wl[34] vdd gnd cell_6t
Xbit_r35_c122 bl[122] br[122] wl[35] vdd gnd cell_6t
Xbit_r36_c122 bl[122] br[122] wl[36] vdd gnd cell_6t
Xbit_r37_c122 bl[122] br[122] wl[37] vdd gnd cell_6t
Xbit_r38_c122 bl[122] br[122] wl[38] vdd gnd cell_6t
Xbit_r39_c122 bl[122] br[122] wl[39] vdd gnd cell_6t
Xbit_r40_c122 bl[122] br[122] wl[40] vdd gnd cell_6t
Xbit_r41_c122 bl[122] br[122] wl[41] vdd gnd cell_6t
Xbit_r42_c122 bl[122] br[122] wl[42] vdd gnd cell_6t
Xbit_r43_c122 bl[122] br[122] wl[43] vdd gnd cell_6t
Xbit_r44_c122 bl[122] br[122] wl[44] vdd gnd cell_6t
Xbit_r45_c122 bl[122] br[122] wl[45] vdd gnd cell_6t
Xbit_r46_c122 bl[122] br[122] wl[46] vdd gnd cell_6t
Xbit_r47_c122 bl[122] br[122] wl[47] vdd gnd cell_6t
Xbit_r48_c122 bl[122] br[122] wl[48] vdd gnd cell_6t
Xbit_r49_c122 bl[122] br[122] wl[49] vdd gnd cell_6t
Xbit_r50_c122 bl[122] br[122] wl[50] vdd gnd cell_6t
Xbit_r51_c122 bl[122] br[122] wl[51] vdd gnd cell_6t
Xbit_r52_c122 bl[122] br[122] wl[52] vdd gnd cell_6t
Xbit_r53_c122 bl[122] br[122] wl[53] vdd gnd cell_6t
Xbit_r54_c122 bl[122] br[122] wl[54] vdd gnd cell_6t
Xbit_r55_c122 bl[122] br[122] wl[55] vdd gnd cell_6t
Xbit_r56_c122 bl[122] br[122] wl[56] vdd gnd cell_6t
Xbit_r57_c122 bl[122] br[122] wl[57] vdd gnd cell_6t
Xbit_r58_c122 bl[122] br[122] wl[58] vdd gnd cell_6t
Xbit_r59_c122 bl[122] br[122] wl[59] vdd gnd cell_6t
Xbit_r60_c122 bl[122] br[122] wl[60] vdd gnd cell_6t
Xbit_r61_c122 bl[122] br[122] wl[61] vdd gnd cell_6t
Xbit_r62_c122 bl[122] br[122] wl[62] vdd gnd cell_6t
Xbit_r63_c122 bl[122] br[122] wl[63] vdd gnd cell_6t
Xbit_r64_c122 bl[122] br[122] wl[64] vdd gnd cell_6t
Xbit_r65_c122 bl[122] br[122] wl[65] vdd gnd cell_6t
Xbit_r66_c122 bl[122] br[122] wl[66] vdd gnd cell_6t
Xbit_r67_c122 bl[122] br[122] wl[67] vdd gnd cell_6t
Xbit_r68_c122 bl[122] br[122] wl[68] vdd gnd cell_6t
Xbit_r69_c122 bl[122] br[122] wl[69] vdd gnd cell_6t
Xbit_r70_c122 bl[122] br[122] wl[70] vdd gnd cell_6t
Xbit_r71_c122 bl[122] br[122] wl[71] vdd gnd cell_6t
Xbit_r72_c122 bl[122] br[122] wl[72] vdd gnd cell_6t
Xbit_r73_c122 bl[122] br[122] wl[73] vdd gnd cell_6t
Xbit_r74_c122 bl[122] br[122] wl[74] vdd gnd cell_6t
Xbit_r75_c122 bl[122] br[122] wl[75] vdd gnd cell_6t
Xbit_r76_c122 bl[122] br[122] wl[76] vdd gnd cell_6t
Xbit_r77_c122 bl[122] br[122] wl[77] vdd gnd cell_6t
Xbit_r78_c122 bl[122] br[122] wl[78] vdd gnd cell_6t
Xbit_r79_c122 bl[122] br[122] wl[79] vdd gnd cell_6t
Xbit_r80_c122 bl[122] br[122] wl[80] vdd gnd cell_6t
Xbit_r81_c122 bl[122] br[122] wl[81] vdd gnd cell_6t
Xbit_r82_c122 bl[122] br[122] wl[82] vdd gnd cell_6t
Xbit_r83_c122 bl[122] br[122] wl[83] vdd gnd cell_6t
Xbit_r84_c122 bl[122] br[122] wl[84] vdd gnd cell_6t
Xbit_r85_c122 bl[122] br[122] wl[85] vdd gnd cell_6t
Xbit_r86_c122 bl[122] br[122] wl[86] vdd gnd cell_6t
Xbit_r87_c122 bl[122] br[122] wl[87] vdd gnd cell_6t
Xbit_r88_c122 bl[122] br[122] wl[88] vdd gnd cell_6t
Xbit_r89_c122 bl[122] br[122] wl[89] vdd gnd cell_6t
Xbit_r90_c122 bl[122] br[122] wl[90] vdd gnd cell_6t
Xbit_r91_c122 bl[122] br[122] wl[91] vdd gnd cell_6t
Xbit_r92_c122 bl[122] br[122] wl[92] vdd gnd cell_6t
Xbit_r93_c122 bl[122] br[122] wl[93] vdd gnd cell_6t
Xbit_r94_c122 bl[122] br[122] wl[94] vdd gnd cell_6t
Xbit_r95_c122 bl[122] br[122] wl[95] vdd gnd cell_6t
Xbit_r96_c122 bl[122] br[122] wl[96] vdd gnd cell_6t
Xbit_r97_c122 bl[122] br[122] wl[97] vdd gnd cell_6t
Xbit_r98_c122 bl[122] br[122] wl[98] vdd gnd cell_6t
Xbit_r99_c122 bl[122] br[122] wl[99] vdd gnd cell_6t
Xbit_r100_c122 bl[122] br[122] wl[100] vdd gnd cell_6t
Xbit_r101_c122 bl[122] br[122] wl[101] vdd gnd cell_6t
Xbit_r102_c122 bl[122] br[122] wl[102] vdd gnd cell_6t
Xbit_r103_c122 bl[122] br[122] wl[103] vdd gnd cell_6t
Xbit_r104_c122 bl[122] br[122] wl[104] vdd gnd cell_6t
Xbit_r105_c122 bl[122] br[122] wl[105] vdd gnd cell_6t
Xbit_r106_c122 bl[122] br[122] wl[106] vdd gnd cell_6t
Xbit_r107_c122 bl[122] br[122] wl[107] vdd gnd cell_6t
Xbit_r108_c122 bl[122] br[122] wl[108] vdd gnd cell_6t
Xbit_r109_c122 bl[122] br[122] wl[109] vdd gnd cell_6t
Xbit_r110_c122 bl[122] br[122] wl[110] vdd gnd cell_6t
Xbit_r111_c122 bl[122] br[122] wl[111] vdd gnd cell_6t
Xbit_r112_c122 bl[122] br[122] wl[112] vdd gnd cell_6t
Xbit_r113_c122 bl[122] br[122] wl[113] vdd gnd cell_6t
Xbit_r114_c122 bl[122] br[122] wl[114] vdd gnd cell_6t
Xbit_r115_c122 bl[122] br[122] wl[115] vdd gnd cell_6t
Xbit_r116_c122 bl[122] br[122] wl[116] vdd gnd cell_6t
Xbit_r117_c122 bl[122] br[122] wl[117] vdd gnd cell_6t
Xbit_r118_c122 bl[122] br[122] wl[118] vdd gnd cell_6t
Xbit_r119_c122 bl[122] br[122] wl[119] vdd gnd cell_6t
Xbit_r120_c122 bl[122] br[122] wl[120] vdd gnd cell_6t
Xbit_r121_c122 bl[122] br[122] wl[121] vdd gnd cell_6t
Xbit_r122_c122 bl[122] br[122] wl[122] vdd gnd cell_6t
Xbit_r123_c122 bl[122] br[122] wl[123] vdd gnd cell_6t
Xbit_r124_c122 bl[122] br[122] wl[124] vdd gnd cell_6t
Xbit_r125_c122 bl[122] br[122] wl[125] vdd gnd cell_6t
Xbit_r126_c122 bl[122] br[122] wl[126] vdd gnd cell_6t
Xbit_r127_c122 bl[122] br[122] wl[127] vdd gnd cell_6t
Xbit_r128_c122 bl[122] br[122] wl[128] vdd gnd cell_6t
Xbit_r129_c122 bl[122] br[122] wl[129] vdd gnd cell_6t
Xbit_r130_c122 bl[122] br[122] wl[130] vdd gnd cell_6t
Xbit_r131_c122 bl[122] br[122] wl[131] vdd gnd cell_6t
Xbit_r132_c122 bl[122] br[122] wl[132] vdd gnd cell_6t
Xbit_r133_c122 bl[122] br[122] wl[133] vdd gnd cell_6t
Xbit_r134_c122 bl[122] br[122] wl[134] vdd gnd cell_6t
Xbit_r135_c122 bl[122] br[122] wl[135] vdd gnd cell_6t
Xbit_r136_c122 bl[122] br[122] wl[136] vdd gnd cell_6t
Xbit_r137_c122 bl[122] br[122] wl[137] vdd gnd cell_6t
Xbit_r138_c122 bl[122] br[122] wl[138] vdd gnd cell_6t
Xbit_r139_c122 bl[122] br[122] wl[139] vdd gnd cell_6t
Xbit_r140_c122 bl[122] br[122] wl[140] vdd gnd cell_6t
Xbit_r141_c122 bl[122] br[122] wl[141] vdd gnd cell_6t
Xbit_r142_c122 bl[122] br[122] wl[142] vdd gnd cell_6t
Xbit_r143_c122 bl[122] br[122] wl[143] vdd gnd cell_6t
Xbit_r144_c122 bl[122] br[122] wl[144] vdd gnd cell_6t
Xbit_r145_c122 bl[122] br[122] wl[145] vdd gnd cell_6t
Xbit_r146_c122 bl[122] br[122] wl[146] vdd gnd cell_6t
Xbit_r147_c122 bl[122] br[122] wl[147] vdd gnd cell_6t
Xbit_r148_c122 bl[122] br[122] wl[148] vdd gnd cell_6t
Xbit_r149_c122 bl[122] br[122] wl[149] vdd gnd cell_6t
Xbit_r150_c122 bl[122] br[122] wl[150] vdd gnd cell_6t
Xbit_r151_c122 bl[122] br[122] wl[151] vdd gnd cell_6t
Xbit_r152_c122 bl[122] br[122] wl[152] vdd gnd cell_6t
Xbit_r153_c122 bl[122] br[122] wl[153] vdd gnd cell_6t
Xbit_r154_c122 bl[122] br[122] wl[154] vdd gnd cell_6t
Xbit_r155_c122 bl[122] br[122] wl[155] vdd gnd cell_6t
Xbit_r156_c122 bl[122] br[122] wl[156] vdd gnd cell_6t
Xbit_r157_c122 bl[122] br[122] wl[157] vdd gnd cell_6t
Xbit_r158_c122 bl[122] br[122] wl[158] vdd gnd cell_6t
Xbit_r159_c122 bl[122] br[122] wl[159] vdd gnd cell_6t
Xbit_r160_c122 bl[122] br[122] wl[160] vdd gnd cell_6t
Xbit_r161_c122 bl[122] br[122] wl[161] vdd gnd cell_6t
Xbit_r162_c122 bl[122] br[122] wl[162] vdd gnd cell_6t
Xbit_r163_c122 bl[122] br[122] wl[163] vdd gnd cell_6t
Xbit_r164_c122 bl[122] br[122] wl[164] vdd gnd cell_6t
Xbit_r165_c122 bl[122] br[122] wl[165] vdd gnd cell_6t
Xbit_r166_c122 bl[122] br[122] wl[166] vdd gnd cell_6t
Xbit_r167_c122 bl[122] br[122] wl[167] vdd gnd cell_6t
Xbit_r168_c122 bl[122] br[122] wl[168] vdd gnd cell_6t
Xbit_r169_c122 bl[122] br[122] wl[169] vdd gnd cell_6t
Xbit_r170_c122 bl[122] br[122] wl[170] vdd gnd cell_6t
Xbit_r171_c122 bl[122] br[122] wl[171] vdd gnd cell_6t
Xbit_r172_c122 bl[122] br[122] wl[172] vdd gnd cell_6t
Xbit_r173_c122 bl[122] br[122] wl[173] vdd gnd cell_6t
Xbit_r174_c122 bl[122] br[122] wl[174] vdd gnd cell_6t
Xbit_r175_c122 bl[122] br[122] wl[175] vdd gnd cell_6t
Xbit_r176_c122 bl[122] br[122] wl[176] vdd gnd cell_6t
Xbit_r177_c122 bl[122] br[122] wl[177] vdd gnd cell_6t
Xbit_r178_c122 bl[122] br[122] wl[178] vdd gnd cell_6t
Xbit_r179_c122 bl[122] br[122] wl[179] vdd gnd cell_6t
Xbit_r180_c122 bl[122] br[122] wl[180] vdd gnd cell_6t
Xbit_r181_c122 bl[122] br[122] wl[181] vdd gnd cell_6t
Xbit_r182_c122 bl[122] br[122] wl[182] vdd gnd cell_6t
Xbit_r183_c122 bl[122] br[122] wl[183] vdd gnd cell_6t
Xbit_r184_c122 bl[122] br[122] wl[184] vdd gnd cell_6t
Xbit_r185_c122 bl[122] br[122] wl[185] vdd gnd cell_6t
Xbit_r186_c122 bl[122] br[122] wl[186] vdd gnd cell_6t
Xbit_r187_c122 bl[122] br[122] wl[187] vdd gnd cell_6t
Xbit_r188_c122 bl[122] br[122] wl[188] vdd gnd cell_6t
Xbit_r189_c122 bl[122] br[122] wl[189] vdd gnd cell_6t
Xbit_r190_c122 bl[122] br[122] wl[190] vdd gnd cell_6t
Xbit_r191_c122 bl[122] br[122] wl[191] vdd gnd cell_6t
Xbit_r192_c122 bl[122] br[122] wl[192] vdd gnd cell_6t
Xbit_r193_c122 bl[122] br[122] wl[193] vdd gnd cell_6t
Xbit_r194_c122 bl[122] br[122] wl[194] vdd gnd cell_6t
Xbit_r195_c122 bl[122] br[122] wl[195] vdd gnd cell_6t
Xbit_r196_c122 bl[122] br[122] wl[196] vdd gnd cell_6t
Xbit_r197_c122 bl[122] br[122] wl[197] vdd gnd cell_6t
Xbit_r198_c122 bl[122] br[122] wl[198] vdd gnd cell_6t
Xbit_r199_c122 bl[122] br[122] wl[199] vdd gnd cell_6t
Xbit_r200_c122 bl[122] br[122] wl[200] vdd gnd cell_6t
Xbit_r201_c122 bl[122] br[122] wl[201] vdd gnd cell_6t
Xbit_r202_c122 bl[122] br[122] wl[202] vdd gnd cell_6t
Xbit_r203_c122 bl[122] br[122] wl[203] vdd gnd cell_6t
Xbit_r204_c122 bl[122] br[122] wl[204] vdd gnd cell_6t
Xbit_r205_c122 bl[122] br[122] wl[205] vdd gnd cell_6t
Xbit_r206_c122 bl[122] br[122] wl[206] vdd gnd cell_6t
Xbit_r207_c122 bl[122] br[122] wl[207] vdd gnd cell_6t
Xbit_r208_c122 bl[122] br[122] wl[208] vdd gnd cell_6t
Xbit_r209_c122 bl[122] br[122] wl[209] vdd gnd cell_6t
Xbit_r210_c122 bl[122] br[122] wl[210] vdd gnd cell_6t
Xbit_r211_c122 bl[122] br[122] wl[211] vdd gnd cell_6t
Xbit_r212_c122 bl[122] br[122] wl[212] vdd gnd cell_6t
Xbit_r213_c122 bl[122] br[122] wl[213] vdd gnd cell_6t
Xbit_r214_c122 bl[122] br[122] wl[214] vdd gnd cell_6t
Xbit_r215_c122 bl[122] br[122] wl[215] vdd gnd cell_6t
Xbit_r216_c122 bl[122] br[122] wl[216] vdd gnd cell_6t
Xbit_r217_c122 bl[122] br[122] wl[217] vdd gnd cell_6t
Xbit_r218_c122 bl[122] br[122] wl[218] vdd gnd cell_6t
Xbit_r219_c122 bl[122] br[122] wl[219] vdd gnd cell_6t
Xbit_r220_c122 bl[122] br[122] wl[220] vdd gnd cell_6t
Xbit_r221_c122 bl[122] br[122] wl[221] vdd gnd cell_6t
Xbit_r222_c122 bl[122] br[122] wl[222] vdd gnd cell_6t
Xbit_r223_c122 bl[122] br[122] wl[223] vdd gnd cell_6t
Xbit_r224_c122 bl[122] br[122] wl[224] vdd gnd cell_6t
Xbit_r225_c122 bl[122] br[122] wl[225] vdd gnd cell_6t
Xbit_r226_c122 bl[122] br[122] wl[226] vdd gnd cell_6t
Xbit_r227_c122 bl[122] br[122] wl[227] vdd gnd cell_6t
Xbit_r228_c122 bl[122] br[122] wl[228] vdd gnd cell_6t
Xbit_r229_c122 bl[122] br[122] wl[229] vdd gnd cell_6t
Xbit_r230_c122 bl[122] br[122] wl[230] vdd gnd cell_6t
Xbit_r231_c122 bl[122] br[122] wl[231] vdd gnd cell_6t
Xbit_r232_c122 bl[122] br[122] wl[232] vdd gnd cell_6t
Xbit_r233_c122 bl[122] br[122] wl[233] vdd gnd cell_6t
Xbit_r234_c122 bl[122] br[122] wl[234] vdd gnd cell_6t
Xbit_r235_c122 bl[122] br[122] wl[235] vdd gnd cell_6t
Xbit_r236_c122 bl[122] br[122] wl[236] vdd gnd cell_6t
Xbit_r237_c122 bl[122] br[122] wl[237] vdd gnd cell_6t
Xbit_r238_c122 bl[122] br[122] wl[238] vdd gnd cell_6t
Xbit_r239_c122 bl[122] br[122] wl[239] vdd gnd cell_6t
Xbit_r240_c122 bl[122] br[122] wl[240] vdd gnd cell_6t
Xbit_r241_c122 bl[122] br[122] wl[241] vdd gnd cell_6t
Xbit_r242_c122 bl[122] br[122] wl[242] vdd gnd cell_6t
Xbit_r243_c122 bl[122] br[122] wl[243] vdd gnd cell_6t
Xbit_r244_c122 bl[122] br[122] wl[244] vdd gnd cell_6t
Xbit_r245_c122 bl[122] br[122] wl[245] vdd gnd cell_6t
Xbit_r246_c122 bl[122] br[122] wl[246] vdd gnd cell_6t
Xbit_r247_c122 bl[122] br[122] wl[247] vdd gnd cell_6t
Xbit_r248_c122 bl[122] br[122] wl[248] vdd gnd cell_6t
Xbit_r249_c122 bl[122] br[122] wl[249] vdd gnd cell_6t
Xbit_r250_c122 bl[122] br[122] wl[250] vdd gnd cell_6t
Xbit_r251_c122 bl[122] br[122] wl[251] vdd gnd cell_6t
Xbit_r252_c122 bl[122] br[122] wl[252] vdd gnd cell_6t
Xbit_r253_c122 bl[122] br[122] wl[253] vdd gnd cell_6t
Xbit_r254_c122 bl[122] br[122] wl[254] vdd gnd cell_6t
Xbit_r255_c122 bl[122] br[122] wl[255] vdd gnd cell_6t
Xbit_r0_c123 bl[123] br[123] wl[0] vdd gnd cell_6t
Xbit_r1_c123 bl[123] br[123] wl[1] vdd gnd cell_6t
Xbit_r2_c123 bl[123] br[123] wl[2] vdd gnd cell_6t
Xbit_r3_c123 bl[123] br[123] wl[3] vdd gnd cell_6t
Xbit_r4_c123 bl[123] br[123] wl[4] vdd gnd cell_6t
Xbit_r5_c123 bl[123] br[123] wl[5] vdd gnd cell_6t
Xbit_r6_c123 bl[123] br[123] wl[6] vdd gnd cell_6t
Xbit_r7_c123 bl[123] br[123] wl[7] vdd gnd cell_6t
Xbit_r8_c123 bl[123] br[123] wl[8] vdd gnd cell_6t
Xbit_r9_c123 bl[123] br[123] wl[9] vdd gnd cell_6t
Xbit_r10_c123 bl[123] br[123] wl[10] vdd gnd cell_6t
Xbit_r11_c123 bl[123] br[123] wl[11] vdd gnd cell_6t
Xbit_r12_c123 bl[123] br[123] wl[12] vdd gnd cell_6t
Xbit_r13_c123 bl[123] br[123] wl[13] vdd gnd cell_6t
Xbit_r14_c123 bl[123] br[123] wl[14] vdd gnd cell_6t
Xbit_r15_c123 bl[123] br[123] wl[15] vdd gnd cell_6t
Xbit_r16_c123 bl[123] br[123] wl[16] vdd gnd cell_6t
Xbit_r17_c123 bl[123] br[123] wl[17] vdd gnd cell_6t
Xbit_r18_c123 bl[123] br[123] wl[18] vdd gnd cell_6t
Xbit_r19_c123 bl[123] br[123] wl[19] vdd gnd cell_6t
Xbit_r20_c123 bl[123] br[123] wl[20] vdd gnd cell_6t
Xbit_r21_c123 bl[123] br[123] wl[21] vdd gnd cell_6t
Xbit_r22_c123 bl[123] br[123] wl[22] vdd gnd cell_6t
Xbit_r23_c123 bl[123] br[123] wl[23] vdd gnd cell_6t
Xbit_r24_c123 bl[123] br[123] wl[24] vdd gnd cell_6t
Xbit_r25_c123 bl[123] br[123] wl[25] vdd gnd cell_6t
Xbit_r26_c123 bl[123] br[123] wl[26] vdd gnd cell_6t
Xbit_r27_c123 bl[123] br[123] wl[27] vdd gnd cell_6t
Xbit_r28_c123 bl[123] br[123] wl[28] vdd gnd cell_6t
Xbit_r29_c123 bl[123] br[123] wl[29] vdd gnd cell_6t
Xbit_r30_c123 bl[123] br[123] wl[30] vdd gnd cell_6t
Xbit_r31_c123 bl[123] br[123] wl[31] vdd gnd cell_6t
Xbit_r32_c123 bl[123] br[123] wl[32] vdd gnd cell_6t
Xbit_r33_c123 bl[123] br[123] wl[33] vdd gnd cell_6t
Xbit_r34_c123 bl[123] br[123] wl[34] vdd gnd cell_6t
Xbit_r35_c123 bl[123] br[123] wl[35] vdd gnd cell_6t
Xbit_r36_c123 bl[123] br[123] wl[36] vdd gnd cell_6t
Xbit_r37_c123 bl[123] br[123] wl[37] vdd gnd cell_6t
Xbit_r38_c123 bl[123] br[123] wl[38] vdd gnd cell_6t
Xbit_r39_c123 bl[123] br[123] wl[39] vdd gnd cell_6t
Xbit_r40_c123 bl[123] br[123] wl[40] vdd gnd cell_6t
Xbit_r41_c123 bl[123] br[123] wl[41] vdd gnd cell_6t
Xbit_r42_c123 bl[123] br[123] wl[42] vdd gnd cell_6t
Xbit_r43_c123 bl[123] br[123] wl[43] vdd gnd cell_6t
Xbit_r44_c123 bl[123] br[123] wl[44] vdd gnd cell_6t
Xbit_r45_c123 bl[123] br[123] wl[45] vdd gnd cell_6t
Xbit_r46_c123 bl[123] br[123] wl[46] vdd gnd cell_6t
Xbit_r47_c123 bl[123] br[123] wl[47] vdd gnd cell_6t
Xbit_r48_c123 bl[123] br[123] wl[48] vdd gnd cell_6t
Xbit_r49_c123 bl[123] br[123] wl[49] vdd gnd cell_6t
Xbit_r50_c123 bl[123] br[123] wl[50] vdd gnd cell_6t
Xbit_r51_c123 bl[123] br[123] wl[51] vdd gnd cell_6t
Xbit_r52_c123 bl[123] br[123] wl[52] vdd gnd cell_6t
Xbit_r53_c123 bl[123] br[123] wl[53] vdd gnd cell_6t
Xbit_r54_c123 bl[123] br[123] wl[54] vdd gnd cell_6t
Xbit_r55_c123 bl[123] br[123] wl[55] vdd gnd cell_6t
Xbit_r56_c123 bl[123] br[123] wl[56] vdd gnd cell_6t
Xbit_r57_c123 bl[123] br[123] wl[57] vdd gnd cell_6t
Xbit_r58_c123 bl[123] br[123] wl[58] vdd gnd cell_6t
Xbit_r59_c123 bl[123] br[123] wl[59] vdd gnd cell_6t
Xbit_r60_c123 bl[123] br[123] wl[60] vdd gnd cell_6t
Xbit_r61_c123 bl[123] br[123] wl[61] vdd gnd cell_6t
Xbit_r62_c123 bl[123] br[123] wl[62] vdd gnd cell_6t
Xbit_r63_c123 bl[123] br[123] wl[63] vdd gnd cell_6t
Xbit_r64_c123 bl[123] br[123] wl[64] vdd gnd cell_6t
Xbit_r65_c123 bl[123] br[123] wl[65] vdd gnd cell_6t
Xbit_r66_c123 bl[123] br[123] wl[66] vdd gnd cell_6t
Xbit_r67_c123 bl[123] br[123] wl[67] vdd gnd cell_6t
Xbit_r68_c123 bl[123] br[123] wl[68] vdd gnd cell_6t
Xbit_r69_c123 bl[123] br[123] wl[69] vdd gnd cell_6t
Xbit_r70_c123 bl[123] br[123] wl[70] vdd gnd cell_6t
Xbit_r71_c123 bl[123] br[123] wl[71] vdd gnd cell_6t
Xbit_r72_c123 bl[123] br[123] wl[72] vdd gnd cell_6t
Xbit_r73_c123 bl[123] br[123] wl[73] vdd gnd cell_6t
Xbit_r74_c123 bl[123] br[123] wl[74] vdd gnd cell_6t
Xbit_r75_c123 bl[123] br[123] wl[75] vdd gnd cell_6t
Xbit_r76_c123 bl[123] br[123] wl[76] vdd gnd cell_6t
Xbit_r77_c123 bl[123] br[123] wl[77] vdd gnd cell_6t
Xbit_r78_c123 bl[123] br[123] wl[78] vdd gnd cell_6t
Xbit_r79_c123 bl[123] br[123] wl[79] vdd gnd cell_6t
Xbit_r80_c123 bl[123] br[123] wl[80] vdd gnd cell_6t
Xbit_r81_c123 bl[123] br[123] wl[81] vdd gnd cell_6t
Xbit_r82_c123 bl[123] br[123] wl[82] vdd gnd cell_6t
Xbit_r83_c123 bl[123] br[123] wl[83] vdd gnd cell_6t
Xbit_r84_c123 bl[123] br[123] wl[84] vdd gnd cell_6t
Xbit_r85_c123 bl[123] br[123] wl[85] vdd gnd cell_6t
Xbit_r86_c123 bl[123] br[123] wl[86] vdd gnd cell_6t
Xbit_r87_c123 bl[123] br[123] wl[87] vdd gnd cell_6t
Xbit_r88_c123 bl[123] br[123] wl[88] vdd gnd cell_6t
Xbit_r89_c123 bl[123] br[123] wl[89] vdd gnd cell_6t
Xbit_r90_c123 bl[123] br[123] wl[90] vdd gnd cell_6t
Xbit_r91_c123 bl[123] br[123] wl[91] vdd gnd cell_6t
Xbit_r92_c123 bl[123] br[123] wl[92] vdd gnd cell_6t
Xbit_r93_c123 bl[123] br[123] wl[93] vdd gnd cell_6t
Xbit_r94_c123 bl[123] br[123] wl[94] vdd gnd cell_6t
Xbit_r95_c123 bl[123] br[123] wl[95] vdd gnd cell_6t
Xbit_r96_c123 bl[123] br[123] wl[96] vdd gnd cell_6t
Xbit_r97_c123 bl[123] br[123] wl[97] vdd gnd cell_6t
Xbit_r98_c123 bl[123] br[123] wl[98] vdd gnd cell_6t
Xbit_r99_c123 bl[123] br[123] wl[99] vdd gnd cell_6t
Xbit_r100_c123 bl[123] br[123] wl[100] vdd gnd cell_6t
Xbit_r101_c123 bl[123] br[123] wl[101] vdd gnd cell_6t
Xbit_r102_c123 bl[123] br[123] wl[102] vdd gnd cell_6t
Xbit_r103_c123 bl[123] br[123] wl[103] vdd gnd cell_6t
Xbit_r104_c123 bl[123] br[123] wl[104] vdd gnd cell_6t
Xbit_r105_c123 bl[123] br[123] wl[105] vdd gnd cell_6t
Xbit_r106_c123 bl[123] br[123] wl[106] vdd gnd cell_6t
Xbit_r107_c123 bl[123] br[123] wl[107] vdd gnd cell_6t
Xbit_r108_c123 bl[123] br[123] wl[108] vdd gnd cell_6t
Xbit_r109_c123 bl[123] br[123] wl[109] vdd gnd cell_6t
Xbit_r110_c123 bl[123] br[123] wl[110] vdd gnd cell_6t
Xbit_r111_c123 bl[123] br[123] wl[111] vdd gnd cell_6t
Xbit_r112_c123 bl[123] br[123] wl[112] vdd gnd cell_6t
Xbit_r113_c123 bl[123] br[123] wl[113] vdd gnd cell_6t
Xbit_r114_c123 bl[123] br[123] wl[114] vdd gnd cell_6t
Xbit_r115_c123 bl[123] br[123] wl[115] vdd gnd cell_6t
Xbit_r116_c123 bl[123] br[123] wl[116] vdd gnd cell_6t
Xbit_r117_c123 bl[123] br[123] wl[117] vdd gnd cell_6t
Xbit_r118_c123 bl[123] br[123] wl[118] vdd gnd cell_6t
Xbit_r119_c123 bl[123] br[123] wl[119] vdd gnd cell_6t
Xbit_r120_c123 bl[123] br[123] wl[120] vdd gnd cell_6t
Xbit_r121_c123 bl[123] br[123] wl[121] vdd gnd cell_6t
Xbit_r122_c123 bl[123] br[123] wl[122] vdd gnd cell_6t
Xbit_r123_c123 bl[123] br[123] wl[123] vdd gnd cell_6t
Xbit_r124_c123 bl[123] br[123] wl[124] vdd gnd cell_6t
Xbit_r125_c123 bl[123] br[123] wl[125] vdd gnd cell_6t
Xbit_r126_c123 bl[123] br[123] wl[126] vdd gnd cell_6t
Xbit_r127_c123 bl[123] br[123] wl[127] vdd gnd cell_6t
Xbit_r128_c123 bl[123] br[123] wl[128] vdd gnd cell_6t
Xbit_r129_c123 bl[123] br[123] wl[129] vdd gnd cell_6t
Xbit_r130_c123 bl[123] br[123] wl[130] vdd gnd cell_6t
Xbit_r131_c123 bl[123] br[123] wl[131] vdd gnd cell_6t
Xbit_r132_c123 bl[123] br[123] wl[132] vdd gnd cell_6t
Xbit_r133_c123 bl[123] br[123] wl[133] vdd gnd cell_6t
Xbit_r134_c123 bl[123] br[123] wl[134] vdd gnd cell_6t
Xbit_r135_c123 bl[123] br[123] wl[135] vdd gnd cell_6t
Xbit_r136_c123 bl[123] br[123] wl[136] vdd gnd cell_6t
Xbit_r137_c123 bl[123] br[123] wl[137] vdd gnd cell_6t
Xbit_r138_c123 bl[123] br[123] wl[138] vdd gnd cell_6t
Xbit_r139_c123 bl[123] br[123] wl[139] vdd gnd cell_6t
Xbit_r140_c123 bl[123] br[123] wl[140] vdd gnd cell_6t
Xbit_r141_c123 bl[123] br[123] wl[141] vdd gnd cell_6t
Xbit_r142_c123 bl[123] br[123] wl[142] vdd gnd cell_6t
Xbit_r143_c123 bl[123] br[123] wl[143] vdd gnd cell_6t
Xbit_r144_c123 bl[123] br[123] wl[144] vdd gnd cell_6t
Xbit_r145_c123 bl[123] br[123] wl[145] vdd gnd cell_6t
Xbit_r146_c123 bl[123] br[123] wl[146] vdd gnd cell_6t
Xbit_r147_c123 bl[123] br[123] wl[147] vdd gnd cell_6t
Xbit_r148_c123 bl[123] br[123] wl[148] vdd gnd cell_6t
Xbit_r149_c123 bl[123] br[123] wl[149] vdd gnd cell_6t
Xbit_r150_c123 bl[123] br[123] wl[150] vdd gnd cell_6t
Xbit_r151_c123 bl[123] br[123] wl[151] vdd gnd cell_6t
Xbit_r152_c123 bl[123] br[123] wl[152] vdd gnd cell_6t
Xbit_r153_c123 bl[123] br[123] wl[153] vdd gnd cell_6t
Xbit_r154_c123 bl[123] br[123] wl[154] vdd gnd cell_6t
Xbit_r155_c123 bl[123] br[123] wl[155] vdd gnd cell_6t
Xbit_r156_c123 bl[123] br[123] wl[156] vdd gnd cell_6t
Xbit_r157_c123 bl[123] br[123] wl[157] vdd gnd cell_6t
Xbit_r158_c123 bl[123] br[123] wl[158] vdd gnd cell_6t
Xbit_r159_c123 bl[123] br[123] wl[159] vdd gnd cell_6t
Xbit_r160_c123 bl[123] br[123] wl[160] vdd gnd cell_6t
Xbit_r161_c123 bl[123] br[123] wl[161] vdd gnd cell_6t
Xbit_r162_c123 bl[123] br[123] wl[162] vdd gnd cell_6t
Xbit_r163_c123 bl[123] br[123] wl[163] vdd gnd cell_6t
Xbit_r164_c123 bl[123] br[123] wl[164] vdd gnd cell_6t
Xbit_r165_c123 bl[123] br[123] wl[165] vdd gnd cell_6t
Xbit_r166_c123 bl[123] br[123] wl[166] vdd gnd cell_6t
Xbit_r167_c123 bl[123] br[123] wl[167] vdd gnd cell_6t
Xbit_r168_c123 bl[123] br[123] wl[168] vdd gnd cell_6t
Xbit_r169_c123 bl[123] br[123] wl[169] vdd gnd cell_6t
Xbit_r170_c123 bl[123] br[123] wl[170] vdd gnd cell_6t
Xbit_r171_c123 bl[123] br[123] wl[171] vdd gnd cell_6t
Xbit_r172_c123 bl[123] br[123] wl[172] vdd gnd cell_6t
Xbit_r173_c123 bl[123] br[123] wl[173] vdd gnd cell_6t
Xbit_r174_c123 bl[123] br[123] wl[174] vdd gnd cell_6t
Xbit_r175_c123 bl[123] br[123] wl[175] vdd gnd cell_6t
Xbit_r176_c123 bl[123] br[123] wl[176] vdd gnd cell_6t
Xbit_r177_c123 bl[123] br[123] wl[177] vdd gnd cell_6t
Xbit_r178_c123 bl[123] br[123] wl[178] vdd gnd cell_6t
Xbit_r179_c123 bl[123] br[123] wl[179] vdd gnd cell_6t
Xbit_r180_c123 bl[123] br[123] wl[180] vdd gnd cell_6t
Xbit_r181_c123 bl[123] br[123] wl[181] vdd gnd cell_6t
Xbit_r182_c123 bl[123] br[123] wl[182] vdd gnd cell_6t
Xbit_r183_c123 bl[123] br[123] wl[183] vdd gnd cell_6t
Xbit_r184_c123 bl[123] br[123] wl[184] vdd gnd cell_6t
Xbit_r185_c123 bl[123] br[123] wl[185] vdd gnd cell_6t
Xbit_r186_c123 bl[123] br[123] wl[186] vdd gnd cell_6t
Xbit_r187_c123 bl[123] br[123] wl[187] vdd gnd cell_6t
Xbit_r188_c123 bl[123] br[123] wl[188] vdd gnd cell_6t
Xbit_r189_c123 bl[123] br[123] wl[189] vdd gnd cell_6t
Xbit_r190_c123 bl[123] br[123] wl[190] vdd gnd cell_6t
Xbit_r191_c123 bl[123] br[123] wl[191] vdd gnd cell_6t
Xbit_r192_c123 bl[123] br[123] wl[192] vdd gnd cell_6t
Xbit_r193_c123 bl[123] br[123] wl[193] vdd gnd cell_6t
Xbit_r194_c123 bl[123] br[123] wl[194] vdd gnd cell_6t
Xbit_r195_c123 bl[123] br[123] wl[195] vdd gnd cell_6t
Xbit_r196_c123 bl[123] br[123] wl[196] vdd gnd cell_6t
Xbit_r197_c123 bl[123] br[123] wl[197] vdd gnd cell_6t
Xbit_r198_c123 bl[123] br[123] wl[198] vdd gnd cell_6t
Xbit_r199_c123 bl[123] br[123] wl[199] vdd gnd cell_6t
Xbit_r200_c123 bl[123] br[123] wl[200] vdd gnd cell_6t
Xbit_r201_c123 bl[123] br[123] wl[201] vdd gnd cell_6t
Xbit_r202_c123 bl[123] br[123] wl[202] vdd gnd cell_6t
Xbit_r203_c123 bl[123] br[123] wl[203] vdd gnd cell_6t
Xbit_r204_c123 bl[123] br[123] wl[204] vdd gnd cell_6t
Xbit_r205_c123 bl[123] br[123] wl[205] vdd gnd cell_6t
Xbit_r206_c123 bl[123] br[123] wl[206] vdd gnd cell_6t
Xbit_r207_c123 bl[123] br[123] wl[207] vdd gnd cell_6t
Xbit_r208_c123 bl[123] br[123] wl[208] vdd gnd cell_6t
Xbit_r209_c123 bl[123] br[123] wl[209] vdd gnd cell_6t
Xbit_r210_c123 bl[123] br[123] wl[210] vdd gnd cell_6t
Xbit_r211_c123 bl[123] br[123] wl[211] vdd gnd cell_6t
Xbit_r212_c123 bl[123] br[123] wl[212] vdd gnd cell_6t
Xbit_r213_c123 bl[123] br[123] wl[213] vdd gnd cell_6t
Xbit_r214_c123 bl[123] br[123] wl[214] vdd gnd cell_6t
Xbit_r215_c123 bl[123] br[123] wl[215] vdd gnd cell_6t
Xbit_r216_c123 bl[123] br[123] wl[216] vdd gnd cell_6t
Xbit_r217_c123 bl[123] br[123] wl[217] vdd gnd cell_6t
Xbit_r218_c123 bl[123] br[123] wl[218] vdd gnd cell_6t
Xbit_r219_c123 bl[123] br[123] wl[219] vdd gnd cell_6t
Xbit_r220_c123 bl[123] br[123] wl[220] vdd gnd cell_6t
Xbit_r221_c123 bl[123] br[123] wl[221] vdd gnd cell_6t
Xbit_r222_c123 bl[123] br[123] wl[222] vdd gnd cell_6t
Xbit_r223_c123 bl[123] br[123] wl[223] vdd gnd cell_6t
Xbit_r224_c123 bl[123] br[123] wl[224] vdd gnd cell_6t
Xbit_r225_c123 bl[123] br[123] wl[225] vdd gnd cell_6t
Xbit_r226_c123 bl[123] br[123] wl[226] vdd gnd cell_6t
Xbit_r227_c123 bl[123] br[123] wl[227] vdd gnd cell_6t
Xbit_r228_c123 bl[123] br[123] wl[228] vdd gnd cell_6t
Xbit_r229_c123 bl[123] br[123] wl[229] vdd gnd cell_6t
Xbit_r230_c123 bl[123] br[123] wl[230] vdd gnd cell_6t
Xbit_r231_c123 bl[123] br[123] wl[231] vdd gnd cell_6t
Xbit_r232_c123 bl[123] br[123] wl[232] vdd gnd cell_6t
Xbit_r233_c123 bl[123] br[123] wl[233] vdd gnd cell_6t
Xbit_r234_c123 bl[123] br[123] wl[234] vdd gnd cell_6t
Xbit_r235_c123 bl[123] br[123] wl[235] vdd gnd cell_6t
Xbit_r236_c123 bl[123] br[123] wl[236] vdd gnd cell_6t
Xbit_r237_c123 bl[123] br[123] wl[237] vdd gnd cell_6t
Xbit_r238_c123 bl[123] br[123] wl[238] vdd gnd cell_6t
Xbit_r239_c123 bl[123] br[123] wl[239] vdd gnd cell_6t
Xbit_r240_c123 bl[123] br[123] wl[240] vdd gnd cell_6t
Xbit_r241_c123 bl[123] br[123] wl[241] vdd gnd cell_6t
Xbit_r242_c123 bl[123] br[123] wl[242] vdd gnd cell_6t
Xbit_r243_c123 bl[123] br[123] wl[243] vdd gnd cell_6t
Xbit_r244_c123 bl[123] br[123] wl[244] vdd gnd cell_6t
Xbit_r245_c123 bl[123] br[123] wl[245] vdd gnd cell_6t
Xbit_r246_c123 bl[123] br[123] wl[246] vdd gnd cell_6t
Xbit_r247_c123 bl[123] br[123] wl[247] vdd gnd cell_6t
Xbit_r248_c123 bl[123] br[123] wl[248] vdd gnd cell_6t
Xbit_r249_c123 bl[123] br[123] wl[249] vdd gnd cell_6t
Xbit_r250_c123 bl[123] br[123] wl[250] vdd gnd cell_6t
Xbit_r251_c123 bl[123] br[123] wl[251] vdd gnd cell_6t
Xbit_r252_c123 bl[123] br[123] wl[252] vdd gnd cell_6t
Xbit_r253_c123 bl[123] br[123] wl[253] vdd gnd cell_6t
Xbit_r254_c123 bl[123] br[123] wl[254] vdd gnd cell_6t
Xbit_r255_c123 bl[123] br[123] wl[255] vdd gnd cell_6t
Xbit_r0_c124 bl[124] br[124] wl[0] vdd gnd cell_6t
Xbit_r1_c124 bl[124] br[124] wl[1] vdd gnd cell_6t
Xbit_r2_c124 bl[124] br[124] wl[2] vdd gnd cell_6t
Xbit_r3_c124 bl[124] br[124] wl[3] vdd gnd cell_6t
Xbit_r4_c124 bl[124] br[124] wl[4] vdd gnd cell_6t
Xbit_r5_c124 bl[124] br[124] wl[5] vdd gnd cell_6t
Xbit_r6_c124 bl[124] br[124] wl[6] vdd gnd cell_6t
Xbit_r7_c124 bl[124] br[124] wl[7] vdd gnd cell_6t
Xbit_r8_c124 bl[124] br[124] wl[8] vdd gnd cell_6t
Xbit_r9_c124 bl[124] br[124] wl[9] vdd gnd cell_6t
Xbit_r10_c124 bl[124] br[124] wl[10] vdd gnd cell_6t
Xbit_r11_c124 bl[124] br[124] wl[11] vdd gnd cell_6t
Xbit_r12_c124 bl[124] br[124] wl[12] vdd gnd cell_6t
Xbit_r13_c124 bl[124] br[124] wl[13] vdd gnd cell_6t
Xbit_r14_c124 bl[124] br[124] wl[14] vdd gnd cell_6t
Xbit_r15_c124 bl[124] br[124] wl[15] vdd gnd cell_6t
Xbit_r16_c124 bl[124] br[124] wl[16] vdd gnd cell_6t
Xbit_r17_c124 bl[124] br[124] wl[17] vdd gnd cell_6t
Xbit_r18_c124 bl[124] br[124] wl[18] vdd gnd cell_6t
Xbit_r19_c124 bl[124] br[124] wl[19] vdd gnd cell_6t
Xbit_r20_c124 bl[124] br[124] wl[20] vdd gnd cell_6t
Xbit_r21_c124 bl[124] br[124] wl[21] vdd gnd cell_6t
Xbit_r22_c124 bl[124] br[124] wl[22] vdd gnd cell_6t
Xbit_r23_c124 bl[124] br[124] wl[23] vdd gnd cell_6t
Xbit_r24_c124 bl[124] br[124] wl[24] vdd gnd cell_6t
Xbit_r25_c124 bl[124] br[124] wl[25] vdd gnd cell_6t
Xbit_r26_c124 bl[124] br[124] wl[26] vdd gnd cell_6t
Xbit_r27_c124 bl[124] br[124] wl[27] vdd gnd cell_6t
Xbit_r28_c124 bl[124] br[124] wl[28] vdd gnd cell_6t
Xbit_r29_c124 bl[124] br[124] wl[29] vdd gnd cell_6t
Xbit_r30_c124 bl[124] br[124] wl[30] vdd gnd cell_6t
Xbit_r31_c124 bl[124] br[124] wl[31] vdd gnd cell_6t
Xbit_r32_c124 bl[124] br[124] wl[32] vdd gnd cell_6t
Xbit_r33_c124 bl[124] br[124] wl[33] vdd gnd cell_6t
Xbit_r34_c124 bl[124] br[124] wl[34] vdd gnd cell_6t
Xbit_r35_c124 bl[124] br[124] wl[35] vdd gnd cell_6t
Xbit_r36_c124 bl[124] br[124] wl[36] vdd gnd cell_6t
Xbit_r37_c124 bl[124] br[124] wl[37] vdd gnd cell_6t
Xbit_r38_c124 bl[124] br[124] wl[38] vdd gnd cell_6t
Xbit_r39_c124 bl[124] br[124] wl[39] vdd gnd cell_6t
Xbit_r40_c124 bl[124] br[124] wl[40] vdd gnd cell_6t
Xbit_r41_c124 bl[124] br[124] wl[41] vdd gnd cell_6t
Xbit_r42_c124 bl[124] br[124] wl[42] vdd gnd cell_6t
Xbit_r43_c124 bl[124] br[124] wl[43] vdd gnd cell_6t
Xbit_r44_c124 bl[124] br[124] wl[44] vdd gnd cell_6t
Xbit_r45_c124 bl[124] br[124] wl[45] vdd gnd cell_6t
Xbit_r46_c124 bl[124] br[124] wl[46] vdd gnd cell_6t
Xbit_r47_c124 bl[124] br[124] wl[47] vdd gnd cell_6t
Xbit_r48_c124 bl[124] br[124] wl[48] vdd gnd cell_6t
Xbit_r49_c124 bl[124] br[124] wl[49] vdd gnd cell_6t
Xbit_r50_c124 bl[124] br[124] wl[50] vdd gnd cell_6t
Xbit_r51_c124 bl[124] br[124] wl[51] vdd gnd cell_6t
Xbit_r52_c124 bl[124] br[124] wl[52] vdd gnd cell_6t
Xbit_r53_c124 bl[124] br[124] wl[53] vdd gnd cell_6t
Xbit_r54_c124 bl[124] br[124] wl[54] vdd gnd cell_6t
Xbit_r55_c124 bl[124] br[124] wl[55] vdd gnd cell_6t
Xbit_r56_c124 bl[124] br[124] wl[56] vdd gnd cell_6t
Xbit_r57_c124 bl[124] br[124] wl[57] vdd gnd cell_6t
Xbit_r58_c124 bl[124] br[124] wl[58] vdd gnd cell_6t
Xbit_r59_c124 bl[124] br[124] wl[59] vdd gnd cell_6t
Xbit_r60_c124 bl[124] br[124] wl[60] vdd gnd cell_6t
Xbit_r61_c124 bl[124] br[124] wl[61] vdd gnd cell_6t
Xbit_r62_c124 bl[124] br[124] wl[62] vdd gnd cell_6t
Xbit_r63_c124 bl[124] br[124] wl[63] vdd gnd cell_6t
Xbit_r64_c124 bl[124] br[124] wl[64] vdd gnd cell_6t
Xbit_r65_c124 bl[124] br[124] wl[65] vdd gnd cell_6t
Xbit_r66_c124 bl[124] br[124] wl[66] vdd gnd cell_6t
Xbit_r67_c124 bl[124] br[124] wl[67] vdd gnd cell_6t
Xbit_r68_c124 bl[124] br[124] wl[68] vdd gnd cell_6t
Xbit_r69_c124 bl[124] br[124] wl[69] vdd gnd cell_6t
Xbit_r70_c124 bl[124] br[124] wl[70] vdd gnd cell_6t
Xbit_r71_c124 bl[124] br[124] wl[71] vdd gnd cell_6t
Xbit_r72_c124 bl[124] br[124] wl[72] vdd gnd cell_6t
Xbit_r73_c124 bl[124] br[124] wl[73] vdd gnd cell_6t
Xbit_r74_c124 bl[124] br[124] wl[74] vdd gnd cell_6t
Xbit_r75_c124 bl[124] br[124] wl[75] vdd gnd cell_6t
Xbit_r76_c124 bl[124] br[124] wl[76] vdd gnd cell_6t
Xbit_r77_c124 bl[124] br[124] wl[77] vdd gnd cell_6t
Xbit_r78_c124 bl[124] br[124] wl[78] vdd gnd cell_6t
Xbit_r79_c124 bl[124] br[124] wl[79] vdd gnd cell_6t
Xbit_r80_c124 bl[124] br[124] wl[80] vdd gnd cell_6t
Xbit_r81_c124 bl[124] br[124] wl[81] vdd gnd cell_6t
Xbit_r82_c124 bl[124] br[124] wl[82] vdd gnd cell_6t
Xbit_r83_c124 bl[124] br[124] wl[83] vdd gnd cell_6t
Xbit_r84_c124 bl[124] br[124] wl[84] vdd gnd cell_6t
Xbit_r85_c124 bl[124] br[124] wl[85] vdd gnd cell_6t
Xbit_r86_c124 bl[124] br[124] wl[86] vdd gnd cell_6t
Xbit_r87_c124 bl[124] br[124] wl[87] vdd gnd cell_6t
Xbit_r88_c124 bl[124] br[124] wl[88] vdd gnd cell_6t
Xbit_r89_c124 bl[124] br[124] wl[89] vdd gnd cell_6t
Xbit_r90_c124 bl[124] br[124] wl[90] vdd gnd cell_6t
Xbit_r91_c124 bl[124] br[124] wl[91] vdd gnd cell_6t
Xbit_r92_c124 bl[124] br[124] wl[92] vdd gnd cell_6t
Xbit_r93_c124 bl[124] br[124] wl[93] vdd gnd cell_6t
Xbit_r94_c124 bl[124] br[124] wl[94] vdd gnd cell_6t
Xbit_r95_c124 bl[124] br[124] wl[95] vdd gnd cell_6t
Xbit_r96_c124 bl[124] br[124] wl[96] vdd gnd cell_6t
Xbit_r97_c124 bl[124] br[124] wl[97] vdd gnd cell_6t
Xbit_r98_c124 bl[124] br[124] wl[98] vdd gnd cell_6t
Xbit_r99_c124 bl[124] br[124] wl[99] vdd gnd cell_6t
Xbit_r100_c124 bl[124] br[124] wl[100] vdd gnd cell_6t
Xbit_r101_c124 bl[124] br[124] wl[101] vdd gnd cell_6t
Xbit_r102_c124 bl[124] br[124] wl[102] vdd gnd cell_6t
Xbit_r103_c124 bl[124] br[124] wl[103] vdd gnd cell_6t
Xbit_r104_c124 bl[124] br[124] wl[104] vdd gnd cell_6t
Xbit_r105_c124 bl[124] br[124] wl[105] vdd gnd cell_6t
Xbit_r106_c124 bl[124] br[124] wl[106] vdd gnd cell_6t
Xbit_r107_c124 bl[124] br[124] wl[107] vdd gnd cell_6t
Xbit_r108_c124 bl[124] br[124] wl[108] vdd gnd cell_6t
Xbit_r109_c124 bl[124] br[124] wl[109] vdd gnd cell_6t
Xbit_r110_c124 bl[124] br[124] wl[110] vdd gnd cell_6t
Xbit_r111_c124 bl[124] br[124] wl[111] vdd gnd cell_6t
Xbit_r112_c124 bl[124] br[124] wl[112] vdd gnd cell_6t
Xbit_r113_c124 bl[124] br[124] wl[113] vdd gnd cell_6t
Xbit_r114_c124 bl[124] br[124] wl[114] vdd gnd cell_6t
Xbit_r115_c124 bl[124] br[124] wl[115] vdd gnd cell_6t
Xbit_r116_c124 bl[124] br[124] wl[116] vdd gnd cell_6t
Xbit_r117_c124 bl[124] br[124] wl[117] vdd gnd cell_6t
Xbit_r118_c124 bl[124] br[124] wl[118] vdd gnd cell_6t
Xbit_r119_c124 bl[124] br[124] wl[119] vdd gnd cell_6t
Xbit_r120_c124 bl[124] br[124] wl[120] vdd gnd cell_6t
Xbit_r121_c124 bl[124] br[124] wl[121] vdd gnd cell_6t
Xbit_r122_c124 bl[124] br[124] wl[122] vdd gnd cell_6t
Xbit_r123_c124 bl[124] br[124] wl[123] vdd gnd cell_6t
Xbit_r124_c124 bl[124] br[124] wl[124] vdd gnd cell_6t
Xbit_r125_c124 bl[124] br[124] wl[125] vdd gnd cell_6t
Xbit_r126_c124 bl[124] br[124] wl[126] vdd gnd cell_6t
Xbit_r127_c124 bl[124] br[124] wl[127] vdd gnd cell_6t
Xbit_r128_c124 bl[124] br[124] wl[128] vdd gnd cell_6t
Xbit_r129_c124 bl[124] br[124] wl[129] vdd gnd cell_6t
Xbit_r130_c124 bl[124] br[124] wl[130] vdd gnd cell_6t
Xbit_r131_c124 bl[124] br[124] wl[131] vdd gnd cell_6t
Xbit_r132_c124 bl[124] br[124] wl[132] vdd gnd cell_6t
Xbit_r133_c124 bl[124] br[124] wl[133] vdd gnd cell_6t
Xbit_r134_c124 bl[124] br[124] wl[134] vdd gnd cell_6t
Xbit_r135_c124 bl[124] br[124] wl[135] vdd gnd cell_6t
Xbit_r136_c124 bl[124] br[124] wl[136] vdd gnd cell_6t
Xbit_r137_c124 bl[124] br[124] wl[137] vdd gnd cell_6t
Xbit_r138_c124 bl[124] br[124] wl[138] vdd gnd cell_6t
Xbit_r139_c124 bl[124] br[124] wl[139] vdd gnd cell_6t
Xbit_r140_c124 bl[124] br[124] wl[140] vdd gnd cell_6t
Xbit_r141_c124 bl[124] br[124] wl[141] vdd gnd cell_6t
Xbit_r142_c124 bl[124] br[124] wl[142] vdd gnd cell_6t
Xbit_r143_c124 bl[124] br[124] wl[143] vdd gnd cell_6t
Xbit_r144_c124 bl[124] br[124] wl[144] vdd gnd cell_6t
Xbit_r145_c124 bl[124] br[124] wl[145] vdd gnd cell_6t
Xbit_r146_c124 bl[124] br[124] wl[146] vdd gnd cell_6t
Xbit_r147_c124 bl[124] br[124] wl[147] vdd gnd cell_6t
Xbit_r148_c124 bl[124] br[124] wl[148] vdd gnd cell_6t
Xbit_r149_c124 bl[124] br[124] wl[149] vdd gnd cell_6t
Xbit_r150_c124 bl[124] br[124] wl[150] vdd gnd cell_6t
Xbit_r151_c124 bl[124] br[124] wl[151] vdd gnd cell_6t
Xbit_r152_c124 bl[124] br[124] wl[152] vdd gnd cell_6t
Xbit_r153_c124 bl[124] br[124] wl[153] vdd gnd cell_6t
Xbit_r154_c124 bl[124] br[124] wl[154] vdd gnd cell_6t
Xbit_r155_c124 bl[124] br[124] wl[155] vdd gnd cell_6t
Xbit_r156_c124 bl[124] br[124] wl[156] vdd gnd cell_6t
Xbit_r157_c124 bl[124] br[124] wl[157] vdd gnd cell_6t
Xbit_r158_c124 bl[124] br[124] wl[158] vdd gnd cell_6t
Xbit_r159_c124 bl[124] br[124] wl[159] vdd gnd cell_6t
Xbit_r160_c124 bl[124] br[124] wl[160] vdd gnd cell_6t
Xbit_r161_c124 bl[124] br[124] wl[161] vdd gnd cell_6t
Xbit_r162_c124 bl[124] br[124] wl[162] vdd gnd cell_6t
Xbit_r163_c124 bl[124] br[124] wl[163] vdd gnd cell_6t
Xbit_r164_c124 bl[124] br[124] wl[164] vdd gnd cell_6t
Xbit_r165_c124 bl[124] br[124] wl[165] vdd gnd cell_6t
Xbit_r166_c124 bl[124] br[124] wl[166] vdd gnd cell_6t
Xbit_r167_c124 bl[124] br[124] wl[167] vdd gnd cell_6t
Xbit_r168_c124 bl[124] br[124] wl[168] vdd gnd cell_6t
Xbit_r169_c124 bl[124] br[124] wl[169] vdd gnd cell_6t
Xbit_r170_c124 bl[124] br[124] wl[170] vdd gnd cell_6t
Xbit_r171_c124 bl[124] br[124] wl[171] vdd gnd cell_6t
Xbit_r172_c124 bl[124] br[124] wl[172] vdd gnd cell_6t
Xbit_r173_c124 bl[124] br[124] wl[173] vdd gnd cell_6t
Xbit_r174_c124 bl[124] br[124] wl[174] vdd gnd cell_6t
Xbit_r175_c124 bl[124] br[124] wl[175] vdd gnd cell_6t
Xbit_r176_c124 bl[124] br[124] wl[176] vdd gnd cell_6t
Xbit_r177_c124 bl[124] br[124] wl[177] vdd gnd cell_6t
Xbit_r178_c124 bl[124] br[124] wl[178] vdd gnd cell_6t
Xbit_r179_c124 bl[124] br[124] wl[179] vdd gnd cell_6t
Xbit_r180_c124 bl[124] br[124] wl[180] vdd gnd cell_6t
Xbit_r181_c124 bl[124] br[124] wl[181] vdd gnd cell_6t
Xbit_r182_c124 bl[124] br[124] wl[182] vdd gnd cell_6t
Xbit_r183_c124 bl[124] br[124] wl[183] vdd gnd cell_6t
Xbit_r184_c124 bl[124] br[124] wl[184] vdd gnd cell_6t
Xbit_r185_c124 bl[124] br[124] wl[185] vdd gnd cell_6t
Xbit_r186_c124 bl[124] br[124] wl[186] vdd gnd cell_6t
Xbit_r187_c124 bl[124] br[124] wl[187] vdd gnd cell_6t
Xbit_r188_c124 bl[124] br[124] wl[188] vdd gnd cell_6t
Xbit_r189_c124 bl[124] br[124] wl[189] vdd gnd cell_6t
Xbit_r190_c124 bl[124] br[124] wl[190] vdd gnd cell_6t
Xbit_r191_c124 bl[124] br[124] wl[191] vdd gnd cell_6t
Xbit_r192_c124 bl[124] br[124] wl[192] vdd gnd cell_6t
Xbit_r193_c124 bl[124] br[124] wl[193] vdd gnd cell_6t
Xbit_r194_c124 bl[124] br[124] wl[194] vdd gnd cell_6t
Xbit_r195_c124 bl[124] br[124] wl[195] vdd gnd cell_6t
Xbit_r196_c124 bl[124] br[124] wl[196] vdd gnd cell_6t
Xbit_r197_c124 bl[124] br[124] wl[197] vdd gnd cell_6t
Xbit_r198_c124 bl[124] br[124] wl[198] vdd gnd cell_6t
Xbit_r199_c124 bl[124] br[124] wl[199] vdd gnd cell_6t
Xbit_r200_c124 bl[124] br[124] wl[200] vdd gnd cell_6t
Xbit_r201_c124 bl[124] br[124] wl[201] vdd gnd cell_6t
Xbit_r202_c124 bl[124] br[124] wl[202] vdd gnd cell_6t
Xbit_r203_c124 bl[124] br[124] wl[203] vdd gnd cell_6t
Xbit_r204_c124 bl[124] br[124] wl[204] vdd gnd cell_6t
Xbit_r205_c124 bl[124] br[124] wl[205] vdd gnd cell_6t
Xbit_r206_c124 bl[124] br[124] wl[206] vdd gnd cell_6t
Xbit_r207_c124 bl[124] br[124] wl[207] vdd gnd cell_6t
Xbit_r208_c124 bl[124] br[124] wl[208] vdd gnd cell_6t
Xbit_r209_c124 bl[124] br[124] wl[209] vdd gnd cell_6t
Xbit_r210_c124 bl[124] br[124] wl[210] vdd gnd cell_6t
Xbit_r211_c124 bl[124] br[124] wl[211] vdd gnd cell_6t
Xbit_r212_c124 bl[124] br[124] wl[212] vdd gnd cell_6t
Xbit_r213_c124 bl[124] br[124] wl[213] vdd gnd cell_6t
Xbit_r214_c124 bl[124] br[124] wl[214] vdd gnd cell_6t
Xbit_r215_c124 bl[124] br[124] wl[215] vdd gnd cell_6t
Xbit_r216_c124 bl[124] br[124] wl[216] vdd gnd cell_6t
Xbit_r217_c124 bl[124] br[124] wl[217] vdd gnd cell_6t
Xbit_r218_c124 bl[124] br[124] wl[218] vdd gnd cell_6t
Xbit_r219_c124 bl[124] br[124] wl[219] vdd gnd cell_6t
Xbit_r220_c124 bl[124] br[124] wl[220] vdd gnd cell_6t
Xbit_r221_c124 bl[124] br[124] wl[221] vdd gnd cell_6t
Xbit_r222_c124 bl[124] br[124] wl[222] vdd gnd cell_6t
Xbit_r223_c124 bl[124] br[124] wl[223] vdd gnd cell_6t
Xbit_r224_c124 bl[124] br[124] wl[224] vdd gnd cell_6t
Xbit_r225_c124 bl[124] br[124] wl[225] vdd gnd cell_6t
Xbit_r226_c124 bl[124] br[124] wl[226] vdd gnd cell_6t
Xbit_r227_c124 bl[124] br[124] wl[227] vdd gnd cell_6t
Xbit_r228_c124 bl[124] br[124] wl[228] vdd gnd cell_6t
Xbit_r229_c124 bl[124] br[124] wl[229] vdd gnd cell_6t
Xbit_r230_c124 bl[124] br[124] wl[230] vdd gnd cell_6t
Xbit_r231_c124 bl[124] br[124] wl[231] vdd gnd cell_6t
Xbit_r232_c124 bl[124] br[124] wl[232] vdd gnd cell_6t
Xbit_r233_c124 bl[124] br[124] wl[233] vdd gnd cell_6t
Xbit_r234_c124 bl[124] br[124] wl[234] vdd gnd cell_6t
Xbit_r235_c124 bl[124] br[124] wl[235] vdd gnd cell_6t
Xbit_r236_c124 bl[124] br[124] wl[236] vdd gnd cell_6t
Xbit_r237_c124 bl[124] br[124] wl[237] vdd gnd cell_6t
Xbit_r238_c124 bl[124] br[124] wl[238] vdd gnd cell_6t
Xbit_r239_c124 bl[124] br[124] wl[239] vdd gnd cell_6t
Xbit_r240_c124 bl[124] br[124] wl[240] vdd gnd cell_6t
Xbit_r241_c124 bl[124] br[124] wl[241] vdd gnd cell_6t
Xbit_r242_c124 bl[124] br[124] wl[242] vdd gnd cell_6t
Xbit_r243_c124 bl[124] br[124] wl[243] vdd gnd cell_6t
Xbit_r244_c124 bl[124] br[124] wl[244] vdd gnd cell_6t
Xbit_r245_c124 bl[124] br[124] wl[245] vdd gnd cell_6t
Xbit_r246_c124 bl[124] br[124] wl[246] vdd gnd cell_6t
Xbit_r247_c124 bl[124] br[124] wl[247] vdd gnd cell_6t
Xbit_r248_c124 bl[124] br[124] wl[248] vdd gnd cell_6t
Xbit_r249_c124 bl[124] br[124] wl[249] vdd gnd cell_6t
Xbit_r250_c124 bl[124] br[124] wl[250] vdd gnd cell_6t
Xbit_r251_c124 bl[124] br[124] wl[251] vdd gnd cell_6t
Xbit_r252_c124 bl[124] br[124] wl[252] vdd gnd cell_6t
Xbit_r253_c124 bl[124] br[124] wl[253] vdd gnd cell_6t
Xbit_r254_c124 bl[124] br[124] wl[254] vdd gnd cell_6t
Xbit_r255_c124 bl[124] br[124] wl[255] vdd gnd cell_6t
Xbit_r0_c125 bl[125] br[125] wl[0] vdd gnd cell_6t
Xbit_r1_c125 bl[125] br[125] wl[1] vdd gnd cell_6t
Xbit_r2_c125 bl[125] br[125] wl[2] vdd gnd cell_6t
Xbit_r3_c125 bl[125] br[125] wl[3] vdd gnd cell_6t
Xbit_r4_c125 bl[125] br[125] wl[4] vdd gnd cell_6t
Xbit_r5_c125 bl[125] br[125] wl[5] vdd gnd cell_6t
Xbit_r6_c125 bl[125] br[125] wl[6] vdd gnd cell_6t
Xbit_r7_c125 bl[125] br[125] wl[7] vdd gnd cell_6t
Xbit_r8_c125 bl[125] br[125] wl[8] vdd gnd cell_6t
Xbit_r9_c125 bl[125] br[125] wl[9] vdd gnd cell_6t
Xbit_r10_c125 bl[125] br[125] wl[10] vdd gnd cell_6t
Xbit_r11_c125 bl[125] br[125] wl[11] vdd gnd cell_6t
Xbit_r12_c125 bl[125] br[125] wl[12] vdd gnd cell_6t
Xbit_r13_c125 bl[125] br[125] wl[13] vdd gnd cell_6t
Xbit_r14_c125 bl[125] br[125] wl[14] vdd gnd cell_6t
Xbit_r15_c125 bl[125] br[125] wl[15] vdd gnd cell_6t
Xbit_r16_c125 bl[125] br[125] wl[16] vdd gnd cell_6t
Xbit_r17_c125 bl[125] br[125] wl[17] vdd gnd cell_6t
Xbit_r18_c125 bl[125] br[125] wl[18] vdd gnd cell_6t
Xbit_r19_c125 bl[125] br[125] wl[19] vdd gnd cell_6t
Xbit_r20_c125 bl[125] br[125] wl[20] vdd gnd cell_6t
Xbit_r21_c125 bl[125] br[125] wl[21] vdd gnd cell_6t
Xbit_r22_c125 bl[125] br[125] wl[22] vdd gnd cell_6t
Xbit_r23_c125 bl[125] br[125] wl[23] vdd gnd cell_6t
Xbit_r24_c125 bl[125] br[125] wl[24] vdd gnd cell_6t
Xbit_r25_c125 bl[125] br[125] wl[25] vdd gnd cell_6t
Xbit_r26_c125 bl[125] br[125] wl[26] vdd gnd cell_6t
Xbit_r27_c125 bl[125] br[125] wl[27] vdd gnd cell_6t
Xbit_r28_c125 bl[125] br[125] wl[28] vdd gnd cell_6t
Xbit_r29_c125 bl[125] br[125] wl[29] vdd gnd cell_6t
Xbit_r30_c125 bl[125] br[125] wl[30] vdd gnd cell_6t
Xbit_r31_c125 bl[125] br[125] wl[31] vdd gnd cell_6t
Xbit_r32_c125 bl[125] br[125] wl[32] vdd gnd cell_6t
Xbit_r33_c125 bl[125] br[125] wl[33] vdd gnd cell_6t
Xbit_r34_c125 bl[125] br[125] wl[34] vdd gnd cell_6t
Xbit_r35_c125 bl[125] br[125] wl[35] vdd gnd cell_6t
Xbit_r36_c125 bl[125] br[125] wl[36] vdd gnd cell_6t
Xbit_r37_c125 bl[125] br[125] wl[37] vdd gnd cell_6t
Xbit_r38_c125 bl[125] br[125] wl[38] vdd gnd cell_6t
Xbit_r39_c125 bl[125] br[125] wl[39] vdd gnd cell_6t
Xbit_r40_c125 bl[125] br[125] wl[40] vdd gnd cell_6t
Xbit_r41_c125 bl[125] br[125] wl[41] vdd gnd cell_6t
Xbit_r42_c125 bl[125] br[125] wl[42] vdd gnd cell_6t
Xbit_r43_c125 bl[125] br[125] wl[43] vdd gnd cell_6t
Xbit_r44_c125 bl[125] br[125] wl[44] vdd gnd cell_6t
Xbit_r45_c125 bl[125] br[125] wl[45] vdd gnd cell_6t
Xbit_r46_c125 bl[125] br[125] wl[46] vdd gnd cell_6t
Xbit_r47_c125 bl[125] br[125] wl[47] vdd gnd cell_6t
Xbit_r48_c125 bl[125] br[125] wl[48] vdd gnd cell_6t
Xbit_r49_c125 bl[125] br[125] wl[49] vdd gnd cell_6t
Xbit_r50_c125 bl[125] br[125] wl[50] vdd gnd cell_6t
Xbit_r51_c125 bl[125] br[125] wl[51] vdd gnd cell_6t
Xbit_r52_c125 bl[125] br[125] wl[52] vdd gnd cell_6t
Xbit_r53_c125 bl[125] br[125] wl[53] vdd gnd cell_6t
Xbit_r54_c125 bl[125] br[125] wl[54] vdd gnd cell_6t
Xbit_r55_c125 bl[125] br[125] wl[55] vdd gnd cell_6t
Xbit_r56_c125 bl[125] br[125] wl[56] vdd gnd cell_6t
Xbit_r57_c125 bl[125] br[125] wl[57] vdd gnd cell_6t
Xbit_r58_c125 bl[125] br[125] wl[58] vdd gnd cell_6t
Xbit_r59_c125 bl[125] br[125] wl[59] vdd gnd cell_6t
Xbit_r60_c125 bl[125] br[125] wl[60] vdd gnd cell_6t
Xbit_r61_c125 bl[125] br[125] wl[61] vdd gnd cell_6t
Xbit_r62_c125 bl[125] br[125] wl[62] vdd gnd cell_6t
Xbit_r63_c125 bl[125] br[125] wl[63] vdd gnd cell_6t
Xbit_r64_c125 bl[125] br[125] wl[64] vdd gnd cell_6t
Xbit_r65_c125 bl[125] br[125] wl[65] vdd gnd cell_6t
Xbit_r66_c125 bl[125] br[125] wl[66] vdd gnd cell_6t
Xbit_r67_c125 bl[125] br[125] wl[67] vdd gnd cell_6t
Xbit_r68_c125 bl[125] br[125] wl[68] vdd gnd cell_6t
Xbit_r69_c125 bl[125] br[125] wl[69] vdd gnd cell_6t
Xbit_r70_c125 bl[125] br[125] wl[70] vdd gnd cell_6t
Xbit_r71_c125 bl[125] br[125] wl[71] vdd gnd cell_6t
Xbit_r72_c125 bl[125] br[125] wl[72] vdd gnd cell_6t
Xbit_r73_c125 bl[125] br[125] wl[73] vdd gnd cell_6t
Xbit_r74_c125 bl[125] br[125] wl[74] vdd gnd cell_6t
Xbit_r75_c125 bl[125] br[125] wl[75] vdd gnd cell_6t
Xbit_r76_c125 bl[125] br[125] wl[76] vdd gnd cell_6t
Xbit_r77_c125 bl[125] br[125] wl[77] vdd gnd cell_6t
Xbit_r78_c125 bl[125] br[125] wl[78] vdd gnd cell_6t
Xbit_r79_c125 bl[125] br[125] wl[79] vdd gnd cell_6t
Xbit_r80_c125 bl[125] br[125] wl[80] vdd gnd cell_6t
Xbit_r81_c125 bl[125] br[125] wl[81] vdd gnd cell_6t
Xbit_r82_c125 bl[125] br[125] wl[82] vdd gnd cell_6t
Xbit_r83_c125 bl[125] br[125] wl[83] vdd gnd cell_6t
Xbit_r84_c125 bl[125] br[125] wl[84] vdd gnd cell_6t
Xbit_r85_c125 bl[125] br[125] wl[85] vdd gnd cell_6t
Xbit_r86_c125 bl[125] br[125] wl[86] vdd gnd cell_6t
Xbit_r87_c125 bl[125] br[125] wl[87] vdd gnd cell_6t
Xbit_r88_c125 bl[125] br[125] wl[88] vdd gnd cell_6t
Xbit_r89_c125 bl[125] br[125] wl[89] vdd gnd cell_6t
Xbit_r90_c125 bl[125] br[125] wl[90] vdd gnd cell_6t
Xbit_r91_c125 bl[125] br[125] wl[91] vdd gnd cell_6t
Xbit_r92_c125 bl[125] br[125] wl[92] vdd gnd cell_6t
Xbit_r93_c125 bl[125] br[125] wl[93] vdd gnd cell_6t
Xbit_r94_c125 bl[125] br[125] wl[94] vdd gnd cell_6t
Xbit_r95_c125 bl[125] br[125] wl[95] vdd gnd cell_6t
Xbit_r96_c125 bl[125] br[125] wl[96] vdd gnd cell_6t
Xbit_r97_c125 bl[125] br[125] wl[97] vdd gnd cell_6t
Xbit_r98_c125 bl[125] br[125] wl[98] vdd gnd cell_6t
Xbit_r99_c125 bl[125] br[125] wl[99] vdd gnd cell_6t
Xbit_r100_c125 bl[125] br[125] wl[100] vdd gnd cell_6t
Xbit_r101_c125 bl[125] br[125] wl[101] vdd gnd cell_6t
Xbit_r102_c125 bl[125] br[125] wl[102] vdd gnd cell_6t
Xbit_r103_c125 bl[125] br[125] wl[103] vdd gnd cell_6t
Xbit_r104_c125 bl[125] br[125] wl[104] vdd gnd cell_6t
Xbit_r105_c125 bl[125] br[125] wl[105] vdd gnd cell_6t
Xbit_r106_c125 bl[125] br[125] wl[106] vdd gnd cell_6t
Xbit_r107_c125 bl[125] br[125] wl[107] vdd gnd cell_6t
Xbit_r108_c125 bl[125] br[125] wl[108] vdd gnd cell_6t
Xbit_r109_c125 bl[125] br[125] wl[109] vdd gnd cell_6t
Xbit_r110_c125 bl[125] br[125] wl[110] vdd gnd cell_6t
Xbit_r111_c125 bl[125] br[125] wl[111] vdd gnd cell_6t
Xbit_r112_c125 bl[125] br[125] wl[112] vdd gnd cell_6t
Xbit_r113_c125 bl[125] br[125] wl[113] vdd gnd cell_6t
Xbit_r114_c125 bl[125] br[125] wl[114] vdd gnd cell_6t
Xbit_r115_c125 bl[125] br[125] wl[115] vdd gnd cell_6t
Xbit_r116_c125 bl[125] br[125] wl[116] vdd gnd cell_6t
Xbit_r117_c125 bl[125] br[125] wl[117] vdd gnd cell_6t
Xbit_r118_c125 bl[125] br[125] wl[118] vdd gnd cell_6t
Xbit_r119_c125 bl[125] br[125] wl[119] vdd gnd cell_6t
Xbit_r120_c125 bl[125] br[125] wl[120] vdd gnd cell_6t
Xbit_r121_c125 bl[125] br[125] wl[121] vdd gnd cell_6t
Xbit_r122_c125 bl[125] br[125] wl[122] vdd gnd cell_6t
Xbit_r123_c125 bl[125] br[125] wl[123] vdd gnd cell_6t
Xbit_r124_c125 bl[125] br[125] wl[124] vdd gnd cell_6t
Xbit_r125_c125 bl[125] br[125] wl[125] vdd gnd cell_6t
Xbit_r126_c125 bl[125] br[125] wl[126] vdd gnd cell_6t
Xbit_r127_c125 bl[125] br[125] wl[127] vdd gnd cell_6t
Xbit_r128_c125 bl[125] br[125] wl[128] vdd gnd cell_6t
Xbit_r129_c125 bl[125] br[125] wl[129] vdd gnd cell_6t
Xbit_r130_c125 bl[125] br[125] wl[130] vdd gnd cell_6t
Xbit_r131_c125 bl[125] br[125] wl[131] vdd gnd cell_6t
Xbit_r132_c125 bl[125] br[125] wl[132] vdd gnd cell_6t
Xbit_r133_c125 bl[125] br[125] wl[133] vdd gnd cell_6t
Xbit_r134_c125 bl[125] br[125] wl[134] vdd gnd cell_6t
Xbit_r135_c125 bl[125] br[125] wl[135] vdd gnd cell_6t
Xbit_r136_c125 bl[125] br[125] wl[136] vdd gnd cell_6t
Xbit_r137_c125 bl[125] br[125] wl[137] vdd gnd cell_6t
Xbit_r138_c125 bl[125] br[125] wl[138] vdd gnd cell_6t
Xbit_r139_c125 bl[125] br[125] wl[139] vdd gnd cell_6t
Xbit_r140_c125 bl[125] br[125] wl[140] vdd gnd cell_6t
Xbit_r141_c125 bl[125] br[125] wl[141] vdd gnd cell_6t
Xbit_r142_c125 bl[125] br[125] wl[142] vdd gnd cell_6t
Xbit_r143_c125 bl[125] br[125] wl[143] vdd gnd cell_6t
Xbit_r144_c125 bl[125] br[125] wl[144] vdd gnd cell_6t
Xbit_r145_c125 bl[125] br[125] wl[145] vdd gnd cell_6t
Xbit_r146_c125 bl[125] br[125] wl[146] vdd gnd cell_6t
Xbit_r147_c125 bl[125] br[125] wl[147] vdd gnd cell_6t
Xbit_r148_c125 bl[125] br[125] wl[148] vdd gnd cell_6t
Xbit_r149_c125 bl[125] br[125] wl[149] vdd gnd cell_6t
Xbit_r150_c125 bl[125] br[125] wl[150] vdd gnd cell_6t
Xbit_r151_c125 bl[125] br[125] wl[151] vdd gnd cell_6t
Xbit_r152_c125 bl[125] br[125] wl[152] vdd gnd cell_6t
Xbit_r153_c125 bl[125] br[125] wl[153] vdd gnd cell_6t
Xbit_r154_c125 bl[125] br[125] wl[154] vdd gnd cell_6t
Xbit_r155_c125 bl[125] br[125] wl[155] vdd gnd cell_6t
Xbit_r156_c125 bl[125] br[125] wl[156] vdd gnd cell_6t
Xbit_r157_c125 bl[125] br[125] wl[157] vdd gnd cell_6t
Xbit_r158_c125 bl[125] br[125] wl[158] vdd gnd cell_6t
Xbit_r159_c125 bl[125] br[125] wl[159] vdd gnd cell_6t
Xbit_r160_c125 bl[125] br[125] wl[160] vdd gnd cell_6t
Xbit_r161_c125 bl[125] br[125] wl[161] vdd gnd cell_6t
Xbit_r162_c125 bl[125] br[125] wl[162] vdd gnd cell_6t
Xbit_r163_c125 bl[125] br[125] wl[163] vdd gnd cell_6t
Xbit_r164_c125 bl[125] br[125] wl[164] vdd gnd cell_6t
Xbit_r165_c125 bl[125] br[125] wl[165] vdd gnd cell_6t
Xbit_r166_c125 bl[125] br[125] wl[166] vdd gnd cell_6t
Xbit_r167_c125 bl[125] br[125] wl[167] vdd gnd cell_6t
Xbit_r168_c125 bl[125] br[125] wl[168] vdd gnd cell_6t
Xbit_r169_c125 bl[125] br[125] wl[169] vdd gnd cell_6t
Xbit_r170_c125 bl[125] br[125] wl[170] vdd gnd cell_6t
Xbit_r171_c125 bl[125] br[125] wl[171] vdd gnd cell_6t
Xbit_r172_c125 bl[125] br[125] wl[172] vdd gnd cell_6t
Xbit_r173_c125 bl[125] br[125] wl[173] vdd gnd cell_6t
Xbit_r174_c125 bl[125] br[125] wl[174] vdd gnd cell_6t
Xbit_r175_c125 bl[125] br[125] wl[175] vdd gnd cell_6t
Xbit_r176_c125 bl[125] br[125] wl[176] vdd gnd cell_6t
Xbit_r177_c125 bl[125] br[125] wl[177] vdd gnd cell_6t
Xbit_r178_c125 bl[125] br[125] wl[178] vdd gnd cell_6t
Xbit_r179_c125 bl[125] br[125] wl[179] vdd gnd cell_6t
Xbit_r180_c125 bl[125] br[125] wl[180] vdd gnd cell_6t
Xbit_r181_c125 bl[125] br[125] wl[181] vdd gnd cell_6t
Xbit_r182_c125 bl[125] br[125] wl[182] vdd gnd cell_6t
Xbit_r183_c125 bl[125] br[125] wl[183] vdd gnd cell_6t
Xbit_r184_c125 bl[125] br[125] wl[184] vdd gnd cell_6t
Xbit_r185_c125 bl[125] br[125] wl[185] vdd gnd cell_6t
Xbit_r186_c125 bl[125] br[125] wl[186] vdd gnd cell_6t
Xbit_r187_c125 bl[125] br[125] wl[187] vdd gnd cell_6t
Xbit_r188_c125 bl[125] br[125] wl[188] vdd gnd cell_6t
Xbit_r189_c125 bl[125] br[125] wl[189] vdd gnd cell_6t
Xbit_r190_c125 bl[125] br[125] wl[190] vdd gnd cell_6t
Xbit_r191_c125 bl[125] br[125] wl[191] vdd gnd cell_6t
Xbit_r192_c125 bl[125] br[125] wl[192] vdd gnd cell_6t
Xbit_r193_c125 bl[125] br[125] wl[193] vdd gnd cell_6t
Xbit_r194_c125 bl[125] br[125] wl[194] vdd gnd cell_6t
Xbit_r195_c125 bl[125] br[125] wl[195] vdd gnd cell_6t
Xbit_r196_c125 bl[125] br[125] wl[196] vdd gnd cell_6t
Xbit_r197_c125 bl[125] br[125] wl[197] vdd gnd cell_6t
Xbit_r198_c125 bl[125] br[125] wl[198] vdd gnd cell_6t
Xbit_r199_c125 bl[125] br[125] wl[199] vdd gnd cell_6t
Xbit_r200_c125 bl[125] br[125] wl[200] vdd gnd cell_6t
Xbit_r201_c125 bl[125] br[125] wl[201] vdd gnd cell_6t
Xbit_r202_c125 bl[125] br[125] wl[202] vdd gnd cell_6t
Xbit_r203_c125 bl[125] br[125] wl[203] vdd gnd cell_6t
Xbit_r204_c125 bl[125] br[125] wl[204] vdd gnd cell_6t
Xbit_r205_c125 bl[125] br[125] wl[205] vdd gnd cell_6t
Xbit_r206_c125 bl[125] br[125] wl[206] vdd gnd cell_6t
Xbit_r207_c125 bl[125] br[125] wl[207] vdd gnd cell_6t
Xbit_r208_c125 bl[125] br[125] wl[208] vdd gnd cell_6t
Xbit_r209_c125 bl[125] br[125] wl[209] vdd gnd cell_6t
Xbit_r210_c125 bl[125] br[125] wl[210] vdd gnd cell_6t
Xbit_r211_c125 bl[125] br[125] wl[211] vdd gnd cell_6t
Xbit_r212_c125 bl[125] br[125] wl[212] vdd gnd cell_6t
Xbit_r213_c125 bl[125] br[125] wl[213] vdd gnd cell_6t
Xbit_r214_c125 bl[125] br[125] wl[214] vdd gnd cell_6t
Xbit_r215_c125 bl[125] br[125] wl[215] vdd gnd cell_6t
Xbit_r216_c125 bl[125] br[125] wl[216] vdd gnd cell_6t
Xbit_r217_c125 bl[125] br[125] wl[217] vdd gnd cell_6t
Xbit_r218_c125 bl[125] br[125] wl[218] vdd gnd cell_6t
Xbit_r219_c125 bl[125] br[125] wl[219] vdd gnd cell_6t
Xbit_r220_c125 bl[125] br[125] wl[220] vdd gnd cell_6t
Xbit_r221_c125 bl[125] br[125] wl[221] vdd gnd cell_6t
Xbit_r222_c125 bl[125] br[125] wl[222] vdd gnd cell_6t
Xbit_r223_c125 bl[125] br[125] wl[223] vdd gnd cell_6t
Xbit_r224_c125 bl[125] br[125] wl[224] vdd gnd cell_6t
Xbit_r225_c125 bl[125] br[125] wl[225] vdd gnd cell_6t
Xbit_r226_c125 bl[125] br[125] wl[226] vdd gnd cell_6t
Xbit_r227_c125 bl[125] br[125] wl[227] vdd gnd cell_6t
Xbit_r228_c125 bl[125] br[125] wl[228] vdd gnd cell_6t
Xbit_r229_c125 bl[125] br[125] wl[229] vdd gnd cell_6t
Xbit_r230_c125 bl[125] br[125] wl[230] vdd gnd cell_6t
Xbit_r231_c125 bl[125] br[125] wl[231] vdd gnd cell_6t
Xbit_r232_c125 bl[125] br[125] wl[232] vdd gnd cell_6t
Xbit_r233_c125 bl[125] br[125] wl[233] vdd gnd cell_6t
Xbit_r234_c125 bl[125] br[125] wl[234] vdd gnd cell_6t
Xbit_r235_c125 bl[125] br[125] wl[235] vdd gnd cell_6t
Xbit_r236_c125 bl[125] br[125] wl[236] vdd gnd cell_6t
Xbit_r237_c125 bl[125] br[125] wl[237] vdd gnd cell_6t
Xbit_r238_c125 bl[125] br[125] wl[238] vdd gnd cell_6t
Xbit_r239_c125 bl[125] br[125] wl[239] vdd gnd cell_6t
Xbit_r240_c125 bl[125] br[125] wl[240] vdd gnd cell_6t
Xbit_r241_c125 bl[125] br[125] wl[241] vdd gnd cell_6t
Xbit_r242_c125 bl[125] br[125] wl[242] vdd gnd cell_6t
Xbit_r243_c125 bl[125] br[125] wl[243] vdd gnd cell_6t
Xbit_r244_c125 bl[125] br[125] wl[244] vdd gnd cell_6t
Xbit_r245_c125 bl[125] br[125] wl[245] vdd gnd cell_6t
Xbit_r246_c125 bl[125] br[125] wl[246] vdd gnd cell_6t
Xbit_r247_c125 bl[125] br[125] wl[247] vdd gnd cell_6t
Xbit_r248_c125 bl[125] br[125] wl[248] vdd gnd cell_6t
Xbit_r249_c125 bl[125] br[125] wl[249] vdd gnd cell_6t
Xbit_r250_c125 bl[125] br[125] wl[250] vdd gnd cell_6t
Xbit_r251_c125 bl[125] br[125] wl[251] vdd gnd cell_6t
Xbit_r252_c125 bl[125] br[125] wl[252] vdd gnd cell_6t
Xbit_r253_c125 bl[125] br[125] wl[253] vdd gnd cell_6t
Xbit_r254_c125 bl[125] br[125] wl[254] vdd gnd cell_6t
Xbit_r255_c125 bl[125] br[125] wl[255] vdd gnd cell_6t
Xbit_r0_c126 bl[126] br[126] wl[0] vdd gnd cell_6t
Xbit_r1_c126 bl[126] br[126] wl[1] vdd gnd cell_6t
Xbit_r2_c126 bl[126] br[126] wl[2] vdd gnd cell_6t
Xbit_r3_c126 bl[126] br[126] wl[3] vdd gnd cell_6t
Xbit_r4_c126 bl[126] br[126] wl[4] vdd gnd cell_6t
Xbit_r5_c126 bl[126] br[126] wl[5] vdd gnd cell_6t
Xbit_r6_c126 bl[126] br[126] wl[6] vdd gnd cell_6t
Xbit_r7_c126 bl[126] br[126] wl[7] vdd gnd cell_6t
Xbit_r8_c126 bl[126] br[126] wl[8] vdd gnd cell_6t
Xbit_r9_c126 bl[126] br[126] wl[9] vdd gnd cell_6t
Xbit_r10_c126 bl[126] br[126] wl[10] vdd gnd cell_6t
Xbit_r11_c126 bl[126] br[126] wl[11] vdd gnd cell_6t
Xbit_r12_c126 bl[126] br[126] wl[12] vdd gnd cell_6t
Xbit_r13_c126 bl[126] br[126] wl[13] vdd gnd cell_6t
Xbit_r14_c126 bl[126] br[126] wl[14] vdd gnd cell_6t
Xbit_r15_c126 bl[126] br[126] wl[15] vdd gnd cell_6t
Xbit_r16_c126 bl[126] br[126] wl[16] vdd gnd cell_6t
Xbit_r17_c126 bl[126] br[126] wl[17] vdd gnd cell_6t
Xbit_r18_c126 bl[126] br[126] wl[18] vdd gnd cell_6t
Xbit_r19_c126 bl[126] br[126] wl[19] vdd gnd cell_6t
Xbit_r20_c126 bl[126] br[126] wl[20] vdd gnd cell_6t
Xbit_r21_c126 bl[126] br[126] wl[21] vdd gnd cell_6t
Xbit_r22_c126 bl[126] br[126] wl[22] vdd gnd cell_6t
Xbit_r23_c126 bl[126] br[126] wl[23] vdd gnd cell_6t
Xbit_r24_c126 bl[126] br[126] wl[24] vdd gnd cell_6t
Xbit_r25_c126 bl[126] br[126] wl[25] vdd gnd cell_6t
Xbit_r26_c126 bl[126] br[126] wl[26] vdd gnd cell_6t
Xbit_r27_c126 bl[126] br[126] wl[27] vdd gnd cell_6t
Xbit_r28_c126 bl[126] br[126] wl[28] vdd gnd cell_6t
Xbit_r29_c126 bl[126] br[126] wl[29] vdd gnd cell_6t
Xbit_r30_c126 bl[126] br[126] wl[30] vdd gnd cell_6t
Xbit_r31_c126 bl[126] br[126] wl[31] vdd gnd cell_6t
Xbit_r32_c126 bl[126] br[126] wl[32] vdd gnd cell_6t
Xbit_r33_c126 bl[126] br[126] wl[33] vdd gnd cell_6t
Xbit_r34_c126 bl[126] br[126] wl[34] vdd gnd cell_6t
Xbit_r35_c126 bl[126] br[126] wl[35] vdd gnd cell_6t
Xbit_r36_c126 bl[126] br[126] wl[36] vdd gnd cell_6t
Xbit_r37_c126 bl[126] br[126] wl[37] vdd gnd cell_6t
Xbit_r38_c126 bl[126] br[126] wl[38] vdd gnd cell_6t
Xbit_r39_c126 bl[126] br[126] wl[39] vdd gnd cell_6t
Xbit_r40_c126 bl[126] br[126] wl[40] vdd gnd cell_6t
Xbit_r41_c126 bl[126] br[126] wl[41] vdd gnd cell_6t
Xbit_r42_c126 bl[126] br[126] wl[42] vdd gnd cell_6t
Xbit_r43_c126 bl[126] br[126] wl[43] vdd gnd cell_6t
Xbit_r44_c126 bl[126] br[126] wl[44] vdd gnd cell_6t
Xbit_r45_c126 bl[126] br[126] wl[45] vdd gnd cell_6t
Xbit_r46_c126 bl[126] br[126] wl[46] vdd gnd cell_6t
Xbit_r47_c126 bl[126] br[126] wl[47] vdd gnd cell_6t
Xbit_r48_c126 bl[126] br[126] wl[48] vdd gnd cell_6t
Xbit_r49_c126 bl[126] br[126] wl[49] vdd gnd cell_6t
Xbit_r50_c126 bl[126] br[126] wl[50] vdd gnd cell_6t
Xbit_r51_c126 bl[126] br[126] wl[51] vdd gnd cell_6t
Xbit_r52_c126 bl[126] br[126] wl[52] vdd gnd cell_6t
Xbit_r53_c126 bl[126] br[126] wl[53] vdd gnd cell_6t
Xbit_r54_c126 bl[126] br[126] wl[54] vdd gnd cell_6t
Xbit_r55_c126 bl[126] br[126] wl[55] vdd gnd cell_6t
Xbit_r56_c126 bl[126] br[126] wl[56] vdd gnd cell_6t
Xbit_r57_c126 bl[126] br[126] wl[57] vdd gnd cell_6t
Xbit_r58_c126 bl[126] br[126] wl[58] vdd gnd cell_6t
Xbit_r59_c126 bl[126] br[126] wl[59] vdd gnd cell_6t
Xbit_r60_c126 bl[126] br[126] wl[60] vdd gnd cell_6t
Xbit_r61_c126 bl[126] br[126] wl[61] vdd gnd cell_6t
Xbit_r62_c126 bl[126] br[126] wl[62] vdd gnd cell_6t
Xbit_r63_c126 bl[126] br[126] wl[63] vdd gnd cell_6t
Xbit_r64_c126 bl[126] br[126] wl[64] vdd gnd cell_6t
Xbit_r65_c126 bl[126] br[126] wl[65] vdd gnd cell_6t
Xbit_r66_c126 bl[126] br[126] wl[66] vdd gnd cell_6t
Xbit_r67_c126 bl[126] br[126] wl[67] vdd gnd cell_6t
Xbit_r68_c126 bl[126] br[126] wl[68] vdd gnd cell_6t
Xbit_r69_c126 bl[126] br[126] wl[69] vdd gnd cell_6t
Xbit_r70_c126 bl[126] br[126] wl[70] vdd gnd cell_6t
Xbit_r71_c126 bl[126] br[126] wl[71] vdd gnd cell_6t
Xbit_r72_c126 bl[126] br[126] wl[72] vdd gnd cell_6t
Xbit_r73_c126 bl[126] br[126] wl[73] vdd gnd cell_6t
Xbit_r74_c126 bl[126] br[126] wl[74] vdd gnd cell_6t
Xbit_r75_c126 bl[126] br[126] wl[75] vdd gnd cell_6t
Xbit_r76_c126 bl[126] br[126] wl[76] vdd gnd cell_6t
Xbit_r77_c126 bl[126] br[126] wl[77] vdd gnd cell_6t
Xbit_r78_c126 bl[126] br[126] wl[78] vdd gnd cell_6t
Xbit_r79_c126 bl[126] br[126] wl[79] vdd gnd cell_6t
Xbit_r80_c126 bl[126] br[126] wl[80] vdd gnd cell_6t
Xbit_r81_c126 bl[126] br[126] wl[81] vdd gnd cell_6t
Xbit_r82_c126 bl[126] br[126] wl[82] vdd gnd cell_6t
Xbit_r83_c126 bl[126] br[126] wl[83] vdd gnd cell_6t
Xbit_r84_c126 bl[126] br[126] wl[84] vdd gnd cell_6t
Xbit_r85_c126 bl[126] br[126] wl[85] vdd gnd cell_6t
Xbit_r86_c126 bl[126] br[126] wl[86] vdd gnd cell_6t
Xbit_r87_c126 bl[126] br[126] wl[87] vdd gnd cell_6t
Xbit_r88_c126 bl[126] br[126] wl[88] vdd gnd cell_6t
Xbit_r89_c126 bl[126] br[126] wl[89] vdd gnd cell_6t
Xbit_r90_c126 bl[126] br[126] wl[90] vdd gnd cell_6t
Xbit_r91_c126 bl[126] br[126] wl[91] vdd gnd cell_6t
Xbit_r92_c126 bl[126] br[126] wl[92] vdd gnd cell_6t
Xbit_r93_c126 bl[126] br[126] wl[93] vdd gnd cell_6t
Xbit_r94_c126 bl[126] br[126] wl[94] vdd gnd cell_6t
Xbit_r95_c126 bl[126] br[126] wl[95] vdd gnd cell_6t
Xbit_r96_c126 bl[126] br[126] wl[96] vdd gnd cell_6t
Xbit_r97_c126 bl[126] br[126] wl[97] vdd gnd cell_6t
Xbit_r98_c126 bl[126] br[126] wl[98] vdd gnd cell_6t
Xbit_r99_c126 bl[126] br[126] wl[99] vdd gnd cell_6t
Xbit_r100_c126 bl[126] br[126] wl[100] vdd gnd cell_6t
Xbit_r101_c126 bl[126] br[126] wl[101] vdd gnd cell_6t
Xbit_r102_c126 bl[126] br[126] wl[102] vdd gnd cell_6t
Xbit_r103_c126 bl[126] br[126] wl[103] vdd gnd cell_6t
Xbit_r104_c126 bl[126] br[126] wl[104] vdd gnd cell_6t
Xbit_r105_c126 bl[126] br[126] wl[105] vdd gnd cell_6t
Xbit_r106_c126 bl[126] br[126] wl[106] vdd gnd cell_6t
Xbit_r107_c126 bl[126] br[126] wl[107] vdd gnd cell_6t
Xbit_r108_c126 bl[126] br[126] wl[108] vdd gnd cell_6t
Xbit_r109_c126 bl[126] br[126] wl[109] vdd gnd cell_6t
Xbit_r110_c126 bl[126] br[126] wl[110] vdd gnd cell_6t
Xbit_r111_c126 bl[126] br[126] wl[111] vdd gnd cell_6t
Xbit_r112_c126 bl[126] br[126] wl[112] vdd gnd cell_6t
Xbit_r113_c126 bl[126] br[126] wl[113] vdd gnd cell_6t
Xbit_r114_c126 bl[126] br[126] wl[114] vdd gnd cell_6t
Xbit_r115_c126 bl[126] br[126] wl[115] vdd gnd cell_6t
Xbit_r116_c126 bl[126] br[126] wl[116] vdd gnd cell_6t
Xbit_r117_c126 bl[126] br[126] wl[117] vdd gnd cell_6t
Xbit_r118_c126 bl[126] br[126] wl[118] vdd gnd cell_6t
Xbit_r119_c126 bl[126] br[126] wl[119] vdd gnd cell_6t
Xbit_r120_c126 bl[126] br[126] wl[120] vdd gnd cell_6t
Xbit_r121_c126 bl[126] br[126] wl[121] vdd gnd cell_6t
Xbit_r122_c126 bl[126] br[126] wl[122] vdd gnd cell_6t
Xbit_r123_c126 bl[126] br[126] wl[123] vdd gnd cell_6t
Xbit_r124_c126 bl[126] br[126] wl[124] vdd gnd cell_6t
Xbit_r125_c126 bl[126] br[126] wl[125] vdd gnd cell_6t
Xbit_r126_c126 bl[126] br[126] wl[126] vdd gnd cell_6t
Xbit_r127_c126 bl[126] br[126] wl[127] vdd gnd cell_6t
Xbit_r128_c126 bl[126] br[126] wl[128] vdd gnd cell_6t
Xbit_r129_c126 bl[126] br[126] wl[129] vdd gnd cell_6t
Xbit_r130_c126 bl[126] br[126] wl[130] vdd gnd cell_6t
Xbit_r131_c126 bl[126] br[126] wl[131] vdd gnd cell_6t
Xbit_r132_c126 bl[126] br[126] wl[132] vdd gnd cell_6t
Xbit_r133_c126 bl[126] br[126] wl[133] vdd gnd cell_6t
Xbit_r134_c126 bl[126] br[126] wl[134] vdd gnd cell_6t
Xbit_r135_c126 bl[126] br[126] wl[135] vdd gnd cell_6t
Xbit_r136_c126 bl[126] br[126] wl[136] vdd gnd cell_6t
Xbit_r137_c126 bl[126] br[126] wl[137] vdd gnd cell_6t
Xbit_r138_c126 bl[126] br[126] wl[138] vdd gnd cell_6t
Xbit_r139_c126 bl[126] br[126] wl[139] vdd gnd cell_6t
Xbit_r140_c126 bl[126] br[126] wl[140] vdd gnd cell_6t
Xbit_r141_c126 bl[126] br[126] wl[141] vdd gnd cell_6t
Xbit_r142_c126 bl[126] br[126] wl[142] vdd gnd cell_6t
Xbit_r143_c126 bl[126] br[126] wl[143] vdd gnd cell_6t
Xbit_r144_c126 bl[126] br[126] wl[144] vdd gnd cell_6t
Xbit_r145_c126 bl[126] br[126] wl[145] vdd gnd cell_6t
Xbit_r146_c126 bl[126] br[126] wl[146] vdd gnd cell_6t
Xbit_r147_c126 bl[126] br[126] wl[147] vdd gnd cell_6t
Xbit_r148_c126 bl[126] br[126] wl[148] vdd gnd cell_6t
Xbit_r149_c126 bl[126] br[126] wl[149] vdd gnd cell_6t
Xbit_r150_c126 bl[126] br[126] wl[150] vdd gnd cell_6t
Xbit_r151_c126 bl[126] br[126] wl[151] vdd gnd cell_6t
Xbit_r152_c126 bl[126] br[126] wl[152] vdd gnd cell_6t
Xbit_r153_c126 bl[126] br[126] wl[153] vdd gnd cell_6t
Xbit_r154_c126 bl[126] br[126] wl[154] vdd gnd cell_6t
Xbit_r155_c126 bl[126] br[126] wl[155] vdd gnd cell_6t
Xbit_r156_c126 bl[126] br[126] wl[156] vdd gnd cell_6t
Xbit_r157_c126 bl[126] br[126] wl[157] vdd gnd cell_6t
Xbit_r158_c126 bl[126] br[126] wl[158] vdd gnd cell_6t
Xbit_r159_c126 bl[126] br[126] wl[159] vdd gnd cell_6t
Xbit_r160_c126 bl[126] br[126] wl[160] vdd gnd cell_6t
Xbit_r161_c126 bl[126] br[126] wl[161] vdd gnd cell_6t
Xbit_r162_c126 bl[126] br[126] wl[162] vdd gnd cell_6t
Xbit_r163_c126 bl[126] br[126] wl[163] vdd gnd cell_6t
Xbit_r164_c126 bl[126] br[126] wl[164] vdd gnd cell_6t
Xbit_r165_c126 bl[126] br[126] wl[165] vdd gnd cell_6t
Xbit_r166_c126 bl[126] br[126] wl[166] vdd gnd cell_6t
Xbit_r167_c126 bl[126] br[126] wl[167] vdd gnd cell_6t
Xbit_r168_c126 bl[126] br[126] wl[168] vdd gnd cell_6t
Xbit_r169_c126 bl[126] br[126] wl[169] vdd gnd cell_6t
Xbit_r170_c126 bl[126] br[126] wl[170] vdd gnd cell_6t
Xbit_r171_c126 bl[126] br[126] wl[171] vdd gnd cell_6t
Xbit_r172_c126 bl[126] br[126] wl[172] vdd gnd cell_6t
Xbit_r173_c126 bl[126] br[126] wl[173] vdd gnd cell_6t
Xbit_r174_c126 bl[126] br[126] wl[174] vdd gnd cell_6t
Xbit_r175_c126 bl[126] br[126] wl[175] vdd gnd cell_6t
Xbit_r176_c126 bl[126] br[126] wl[176] vdd gnd cell_6t
Xbit_r177_c126 bl[126] br[126] wl[177] vdd gnd cell_6t
Xbit_r178_c126 bl[126] br[126] wl[178] vdd gnd cell_6t
Xbit_r179_c126 bl[126] br[126] wl[179] vdd gnd cell_6t
Xbit_r180_c126 bl[126] br[126] wl[180] vdd gnd cell_6t
Xbit_r181_c126 bl[126] br[126] wl[181] vdd gnd cell_6t
Xbit_r182_c126 bl[126] br[126] wl[182] vdd gnd cell_6t
Xbit_r183_c126 bl[126] br[126] wl[183] vdd gnd cell_6t
Xbit_r184_c126 bl[126] br[126] wl[184] vdd gnd cell_6t
Xbit_r185_c126 bl[126] br[126] wl[185] vdd gnd cell_6t
Xbit_r186_c126 bl[126] br[126] wl[186] vdd gnd cell_6t
Xbit_r187_c126 bl[126] br[126] wl[187] vdd gnd cell_6t
Xbit_r188_c126 bl[126] br[126] wl[188] vdd gnd cell_6t
Xbit_r189_c126 bl[126] br[126] wl[189] vdd gnd cell_6t
Xbit_r190_c126 bl[126] br[126] wl[190] vdd gnd cell_6t
Xbit_r191_c126 bl[126] br[126] wl[191] vdd gnd cell_6t
Xbit_r192_c126 bl[126] br[126] wl[192] vdd gnd cell_6t
Xbit_r193_c126 bl[126] br[126] wl[193] vdd gnd cell_6t
Xbit_r194_c126 bl[126] br[126] wl[194] vdd gnd cell_6t
Xbit_r195_c126 bl[126] br[126] wl[195] vdd gnd cell_6t
Xbit_r196_c126 bl[126] br[126] wl[196] vdd gnd cell_6t
Xbit_r197_c126 bl[126] br[126] wl[197] vdd gnd cell_6t
Xbit_r198_c126 bl[126] br[126] wl[198] vdd gnd cell_6t
Xbit_r199_c126 bl[126] br[126] wl[199] vdd gnd cell_6t
Xbit_r200_c126 bl[126] br[126] wl[200] vdd gnd cell_6t
Xbit_r201_c126 bl[126] br[126] wl[201] vdd gnd cell_6t
Xbit_r202_c126 bl[126] br[126] wl[202] vdd gnd cell_6t
Xbit_r203_c126 bl[126] br[126] wl[203] vdd gnd cell_6t
Xbit_r204_c126 bl[126] br[126] wl[204] vdd gnd cell_6t
Xbit_r205_c126 bl[126] br[126] wl[205] vdd gnd cell_6t
Xbit_r206_c126 bl[126] br[126] wl[206] vdd gnd cell_6t
Xbit_r207_c126 bl[126] br[126] wl[207] vdd gnd cell_6t
Xbit_r208_c126 bl[126] br[126] wl[208] vdd gnd cell_6t
Xbit_r209_c126 bl[126] br[126] wl[209] vdd gnd cell_6t
Xbit_r210_c126 bl[126] br[126] wl[210] vdd gnd cell_6t
Xbit_r211_c126 bl[126] br[126] wl[211] vdd gnd cell_6t
Xbit_r212_c126 bl[126] br[126] wl[212] vdd gnd cell_6t
Xbit_r213_c126 bl[126] br[126] wl[213] vdd gnd cell_6t
Xbit_r214_c126 bl[126] br[126] wl[214] vdd gnd cell_6t
Xbit_r215_c126 bl[126] br[126] wl[215] vdd gnd cell_6t
Xbit_r216_c126 bl[126] br[126] wl[216] vdd gnd cell_6t
Xbit_r217_c126 bl[126] br[126] wl[217] vdd gnd cell_6t
Xbit_r218_c126 bl[126] br[126] wl[218] vdd gnd cell_6t
Xbit_r219_c126 bl[126] br[126] wl[219] vdd gnd cell_6t
Xbit_r220_c126 bl[126] br[126] wl[220] vdd gnd cell_6t
Xbit_r221_c126 bl[126] br[126] wl[221] vdd gnd cell_6t
Xbit_r222_c126 bl[126] br[126] wl[222] vdd gnd cell_6t
Xbit_r223_c126 bl[126] br[126] wl[223] vdd gnd cell_6t
Xbit_r224_c126 bl[126] br[126] wl[224] vdd gnd cell_6t
Xbit_r225_c126 bl[126] br[126] wl[225] vdd gnd cell_6t
Xbit_r226_c126 bl[126] br[126] wl[226] vdd gnd cell_6t
Xbit_r227_c126 bl[126] br[126] wl[227] vdd gnd cell_6t
Xbit_r228_c126 bl[126] br[126] wl[228] vdd gnd cell_6t
Xbit_r229_c126 bl[126] br[126] wl[229] vdd gnd cell_6t
Xbit_r230_c126 bl[126] br[126] wl[230] vdd gnd cell_6t
Xbit_r231_c126 bl[126] br[126] wl[231] vdd gnd cell_6t
Xbit_r232_c126 bl[126] br[126] wl[232] vdd gnd cell_6t
Xbit_r233_c126 bl[126] br[126] wl[233] vdd gnd cell_6t
Xbit_r234_c126 bl[126] br[126] wl[234] vdd gnd cell_6t
Xbit_r235_c126 bl[126] br[126] wl[235] vdd gnd cell_6t
Xbit_r236_c126 bl[126] br[126] wl[236] vdd gnd cell_6t
Xbit_r237_c126 bl[126] br[126] wl[237] vdd gnd cell_6t
Xbit_r238_c126 bl[126] br[126] wl[238] vdd gnd cell_6t
Xbit_r239_c126 bl[126] br[126] wl[239] vdd gnd cell_6t
Xbit_r240_c126 bl[126] br[126] wl[240] vdd gnd cell_6t
Xbit_r241_c126 bl[126] br[126] wl[241] vdd gnd cell_6t
Xbit_r242_c126 bl[126] br[126] wl[242] vdd gnd cell_6t
Xbit_r243_c126 bl[126] br[126] wl[243] vdd gnd cell_6t
Xbit_r244_c126 bl[126] br[126] wl[244] vdd gnd cell_6t
Xbit_r245_c126 bl[126] br[126] wl[245] vdd gnd cell_6t
Xbit_r246_c126 bl[126] br[126] wl[246] vdd gnd cell_6t
Xbit_r247_c126 bl[126] br[126] wl[247] vdd gnd cell_6t
Xbit_r248_c126 bl[126] br[126] wl[248] vdd gnd cell_6t
Xbit_r249_c126 bl[126] br[126] wl[249] vdd gnd cell_6t
Xbit_r250_c126 bl[126] br[126] wl[250] vdd gnd cell_6t
Xbit_r251_c126 bl[126] br[126] wl[251] vdd gnd cell_6t
Xbit_r252_c126 bl[126] br[126] wl[252] vdd gnd cell_6t
Xbit_r253_c126 bl[126] br[126] wl[253] vdd gnd cell_6t
Xbit_r254_c126 bl[126] br[126] wl[254] vdd gnd cell_6t
Xbit_r255_c126 bl[126] br[126] wl[255] vdd gnd cell_6t
Xbit_r0_c127 bl[127] br[127] wl[0] vdd gnd cell_6t
Xbit_r1_c127 bl[127] br[127] wl[1] vdd gnd cell_6t
Xbit_r2_c127 bl[127] br[127] wl[2] vdd gnd cell_6t
Xbit_r3_c127 bl[127] br[127] wl[3] vdd gnd cell_6t
Xbit_r4_c127 bl[127] br[127] wl[4] vdd gnd cell_6t
Xbit_r5_c127 bl[127] br[127] wl[5] vdd gnd cell_6t
Xbit_r6_c127 bl[127] br[127] wl[6] vdd gnd cell_6t
Xbit_r7_c127 bl[127] br[127] wl[7] vdd gnd cell_6t
Xbit_r8_c127 bl[127] br[127] wl[8] vdd gnd cell_6t
Xbit_r9_c127 bl[127] br[127] wl[9] vdd gnd cell_6t
Xbit_r10_c127 bl[127] br[127] wl[10] vdd gnd cell_6t
Xbit_r11_c127 bl[127] br[127] wl[11] vdd gnd cell_6t
Xbit_r12_c127 bl[127] br[127] wl[12] vdd gnd cell_6t
Xbit_r13_c127 bl[127] br[127] wl[13] vdd gnd cell_6t
Xbit_r14_c127 bl[127] br[127] wl[14] vdd gnd cell_6t
Xbit_r15_c127 bl[127] br[127] wl[15] vdd gnd cell_6t
Xbit_r16_c127 bl[127] br[127] wl[16] vdd gnd cell_6t
Xbit_r17_c127 bl[127] br[127] wl[17] vdd gnd cell_6t
Xbit_r18_c127 bl[127] br[127] wl[18] vdd gnd cell_6t
Xbit_r19_c127 bl[127] br[127] wl[19] vdd gnd cell_6t
Xbit_r20_c127 bl[127] br[127] wl[20] vdd gnd cell_6t
Xbit_r21_c127 bl[127] br[127] wl[21] vdd gnd cell_6t
Xbit_r22_c127 bl[127] br[127] wl[22] vdd gnd cell_6t
Xbit_r23_c127 bl[127] br[127] wl[23] vdd gnd cell_6t
Xbit_r24_c127 bl[127] br[127] wl[24] vdd gnd cell_6t
Xbit_r25_c127 bl[127] br[127] wl[25] vdd gnd cell_6t
Xbit_r26_c127 bl[127] br[127] wl[26] vdd gnd cell_6t
Xbit_r27_c127 bl[127] br[127] wl[27] vdd gnd cell_6t
Xbit_r28_c127 bl[127] br[127] wl[28] vdd gnd cell_6t
Xbit_r29_c127 bl[127] br[127] wl[29] vdd gnd cell_6t
Xbit_r30_c127 bl[127] br[127] wl[30] vdd gnd cell_6t
Xbit_r31_c127 bl[127] br[127] wl[31] vdd gnd cell_6t
Xbit_r32_c127 bl[127] br[127] wl[32] vdd gnd cell_6t
Xbit_r33_c127 bl[127] br[127] wl[33] vdd gnd cell_6t
Xbit_r34_c127 bl[127] br[127] wl[34] vdd gnd cell_6t
Xbit_r35_c127 bl[127] br[127] wl[35] vdd gnd cell_6t
Xbit_r36_c127 bl[127] br[127] wl[36] vdd gnd cell_6t
Xbit_r37_c127 bl[127] br[127] wl[37] vdd gnd cell_6t
Xbit_r38_c127 bl[127] br[127] wl[38] vdd gnd cell_6t
Xbit_r39_c127 bl[127] br[127] wl[39] vdd gnd cell_6t
Xbit_r40_c127 bl[127] br[127] wl[40] vdd gnd cell_6t
Xbit_r41_c127 bl[127] br[127] wl[41] vdd gnd cell_6t
Xbit_r42_c127 bl[127] br[127] wl[42] vdd gnd cell_6t
Xbit_r43_c127 bl[127] br[127] wl[43] vdd gnd cell_6t
Xbit_r44_c127 bl[127] br[127] wl[44] vdd gnd cell_6t
Xbit_r45_c127 bl[127] br[127] wl[45] vdd gnd cell_6t
Xbit_r46_c127 bl[127] br[127] wl[46] vdd gnd cell_6t
Xbit_r47_c127 bl[127] br[127] wl[47] vdd gnd cell_6t
Xbit_r48_c127 bl[127] br[127] wl[48] vdd gnd cell_6t
Xbit_r49_c127 bl[127] br[127] wl[49] vdd gnd cell_6t
Xbit_r50_c127 bl[127] br[127] wl[50] vdd gnd cell_6t
Xbit_r51_c127 bl[127] br[127] wl[51] vdd gnd cell_6t
Xbit_r52_c127 bl[127] br[127] wl[52] vdd gnd cell_6t
Xbit_r53_c127 bl[127] br[127] wl[53] vdd gnd cell_6t
Xbit_r54_c127 bl[127] br[127] wl[54] vdd gnd cell_6t
Xbit_r55_c127 bl[127] br[127] wl[55] vdd gnd cell_6t
Xbit_r56_c127 bl[127] br[127] wl[56] vdd gnd cell_6t
Xbit_r57_c127 bl[127] br[127] wl[57] vdd gnd cell_6t
Xbit_r58_c127 bl[127] br[127] wl[58] vdd gnd cell_6t
Xbit_r59_c127 bl[127] br[127] wl[59] vdd gnd cell_6t
Xbit_r60_c127 bl[127] br[127] wl[60] vdd gnd cell_6t
Xbit_r61_c127 bl[127] br[127] wl[61] vdd gnd cell_6t
Xbit_r62_c127 bl[127] br[127] wl[62] vdd gnd cell_6t
Xbit_r63_c127 bl[127] br[127] wl[63] vdd gnd cell_6t
Xbit_r64_c127 bl[127] br[127] wl[64] vdd gnd cell_6t
Xbit_r65_c127 bl[127] br[127] wl[65] vdd gnd cell_6t
Xbit_r66_c127 bl[127] br[127] wl[66] vdd gnd cell_6t
Xbit_r67_c127 bl[127] br[127] wl[67] vdd gnd cell_6t
Xbit_r68_c127 bl[127] br[127] wl[68] vdd gnd cell_6t
Xbit_r69_c127 bl[127] br[127] wl[69] vdd gnd cell_6t
Xbit_r70_c127 bl[127] br[127] wl[70] vdd gnd cell_6t
Xbit_r71_c127 bl[127] br[127] wl[71] vdd gnd cell_6t
Xbit_r72_c127 bl[127] br[127] wl[72] vdd gnd cell_6t
Xbit_r73_c127 bl[127] br[127] wl[73] vdd gnd cell_6t
Xbit_r74_c127 bl[127] br[127] wl[74] vdd gnd cell_6t
Xbit_r75_c127 bl[127] br[127] wl[75] vdd gnd cell_6t
Xbit_r76_c127 bl[127] br[127] wl[76] vdd gnd cell_6t
Xbit_r77_c127 bl[127] br[127] wl[77] vdd gnd cell_6t
Xbit_r78_c127 bl[127] br[127] wl[78] vdd gnd cell_6t
Xbit_r79_c127 bl[127] br[127] wl[79] vdd gnd cell_6t
Xbit_r80_c127 bl[127] br[127] wl[80] vdd gnd cell_6t
Xbit_r81_c127 bl[127] br[127] wl[81] vdd gnd cell_6t
Xbit_r82_c127 bl[127] br[127] wl[82] vdd gnd cell_6t
Xbit_r83_c127 bl[127] br[127] wl[83] vdd gnd cell_6t
Xbit_r84_c127 bl[127] br[127] wl[84] vdd gnd cell_6t
Xbit_r85_c127 bl[127] br[127] wl[85] vdd gnd cell_6t
Xbit_r86_c127 bl[127] br[127] wl[86] vdd gnd cell_6t
Xbit_r87_c127 bl[127] br[127] wl[87] vdd gnd cell_6t
Xbit_r88_c127 bl[127] br[127] wl[88] vdd gnd cell_6t
Xbit_r89_c127 bl[127] br[127] wl[89] vdd gnd cell_6t
Xbit_r90_c127 bl[127] br[127] wl[90] vdd gnd cell_6t
Xbit_r91_c127 bl[127] br[127] wl[91] vdd gnd cell_6t
Xbit_r92_c127 bl[127] br[127] wl[92] vdd gnd cell_6t
Xbit_r93_c127 bl[127] br[127] wl[93] vdd gnd cell_6t
Xbit_r94_c127 bl[127] br[127] wl[94] vdd gnd cell_6t
Xbit_r95_c127 bl[127] br[127] wl[95] vdd gnd cell_6t
Xbit_r96_c127 bl[127] br[127] wl[96] vdd gnd cell_6t
Xbit_r97_c127 bl[127] br[127] wl[97] vdd gnd cell_6t
Xbit_r98_c127 bl[127] br[127] wl[98] vdd gnd cell_6t
Xbit_r99_c127 bl[127] br[127] wl[99] vdd gnd cell_6t
Xbit_r100_c127 bl[127] br[127] wl[100] vdd gnd cell_6t
Xbit_r101_c127 bl[127] br[127] wl[101] vdd gnd cell_6t
Xbit_r102_c127 bl[127] br[127] wl[102] vdd gnd cell_6t
Xbit_r103_c127 bl[127] br[127] wl[103] vdd gnd cell_6t
Xbit_r104_c127 bl[127] br[127] wl[104] vdd gnd cell_6t
Xbit_r105_c127 bl[127] br[127] wl[105] vdd gnd cell_6t
Xbit_r106_c127 bl[127] br[127] wl[106] vdd gnd cell_6t
Xbit_r107_c127 bl[127] br[127] wl[107] vdd gnd cell_6t
Xbit_r108_c127 bl[127] br[127] wl[108] vdd gnd cell_6t
Xbit_r109_c127 bl[127] br[127] wl[109] vdd gnd cell_6t
Xbit_r110_c127 bl[127] br[127] wl[110] vdd gnd cell_6t
Xbit_r111_c127 bl[127] br[127] wl[111] vdd gnd cell_6t
Xbit_r112_c127 bl[127] br[127] wl[112] vdd gnd cell_6t
Xbit_r113_c127 bl[127] br[127] wl[113] vdd gnd cell_6t
Xbit_r114_c127 bl[127] br[127] wl[114] vdd gnd cell_6t
Xbit_r115_c127 bl[127] br[127] wl[115] vdd gnd cell_6t
Xbit_r116_c127 bl[127] br[127] wl[116] vdd gnd cell_6t
Xbit_r117_c127 bl[127] br[127] wl[117] vdd gnd cell_6t
Xbit_r118_c127 bl[127] br[127] wl[118] vdd gnd cell_6t
Xbit_r119_c127 bl[127] br[127] wl[119] vdd gnd cell_6t
Xbit_r120_c127 bl[127] br[127] wl[120] vdd gnd cell_6t
Xbit_r121_c127 bl[127] br[127] wl[121] vdd gnd cell_6t
Xbit_r122_c127 bl[127] br[127] wl[122] vdd gnd cell_6t
Xbit_r123_c127 bl[127] br[127] wl[123] vdd gnd cell_6t
Xbit_r124_c127 bl[127] br[127] wl[124] vdd gnd cell_6t
Xbit_r125_c127 bl[127] br[127] wl[125] vdd gnd cell_6t
Xbit_r126_c127 bl[127] br[127] wl[126] vdd gnd cell_6t
Xbit_r127_c127 bl[127] br[127] wl[127] vdd gnd cell_6t
Xbit_r128_c127 bl[127] br[127] wl[128] vdd gnd cell_6t
Xbit_r129_c127 bl[127] br[127] wl[129] vdd gnd cell_6t
Xbit_r130_c127 bl[127] br[127] wl[130] vdd gnd cell_6t
Xbit_r131_c127 bl[127] br[127] wl[131] vdd gnd cell_6t
Xbit_r132_c127 bl[127] br[127] wl[132] vdd gnd cell_6t
Xbit_r133_c127 bl[127] br[127] wl[133] vdd gnd cell_6t
Xbit_r134_c127 bl[127] br[127] wl[134] vdd gnd cell_6t
Xbit_r135_c127 bl[127] br[127] wl[135] vdd gnd cell_6t
Xbit_r136_c127 bl[127] br[127] wl[136] vdd gnd cell_6t
Xbit_r137_c127 bl[127] br[127] wl[137] vdd gnd cell_6t
Xbit_r138_c127 bl[127] br[127] wl[138] vdd gnd cell_6t
Xbit_r139_c127 bl[127] br[127] wl[139] vdd gnd cell_6t
Xbit_r140_c127 bl[127] br[127] wl[140] vdd gnd cell_6t
Xbit_r141_c127 bl[127] br[127] wl[141] vdd gnd cell_6t
Xbit_r142_c127 bl[127] br[127] wl[142] vdd gnd cell_6t
Xbit_r143_c127 bl[127] br[127] wl[143] vdd gnd cell_6t
Xbit_r144_c127 bl[127] br[127] wl[144] vdd gnd cell_6t
Xbit_r145_c127 bl[127] br[127] wl[145] vdd gnd cell_6t
Xbit_r146_c127 bl[127] br[127] wl[146] vdd gnd cell_6t
Xbit_r147_c127 bl[127] br[127] wl[147] vdd gnd cell_6t
Xbit_r148_c127 bl[127] br[127] wl[148] vdd gnd cell_6t
Xbit_r149_c127 bl[127] br[127] wl[149] vdd gnd cell_6t
Xbit_r150_c127 bl[127] br[127] wl[150] vdd gnd cell_6t
Xbit_r151_c127 bl[127] br[127] wl[151] vdd gnd cell_6t
Xbit_r152_c127 bl[127] br[127] wl[152] vdd gnd cell_6t
Xbit_r153_c127 bl[127] br[127] wl[153] vdd gnd cell_6t
Xbit_r154_c127 bl[127] br[127] wl[154] vdd gnd cell_6t
Xbit_r155_c127 bl[127] br[127] wl[155] vdd gnd cell_6t
Xbit_r156_c127 bl[127] br[127] wl[156] vdd gnd cell_6t
Xbit_r157_c127 bl[127] br[127] wl[157] vdd gnd cell_6t
Xbit_r158_c127 bl[127] br[127] wl[158] vdd gnd cell_6t
Xbit_r159_c127 bl[127] br[127] wl[159] vdd gnd cell_6t
Xbit_r160_c127 bl[127] br[127] wl[160] vdd gnd cell_6t
Xbit_r161_c127 bl[127] br[127] wl[161] vdd gnd cell_6t
Xbit_r162_c127 bl[127] br[127] wl[162] vdd gnd cell_6t
Xbit_r163_c127 bl[127] br[127] wl[163] vdd gnd cell_6t
Xbit_r164_c127 bl[127] br[127] wl[164] vdd gnd cell_6t
Xbit_r165_c127 bl[127] br[127] wl[165] vdd gnd cell_6t
Xbit_r166_c127 bl[127] br[127] wl[166] vdd gnd cell_6t
Xbit_r167_c127 bl[127] br[127] wl[167] vdd gnd cell_6t
Xbit_r168_c127 bl[127] br[127] wl[168] vdd gnd cell_6t
Xbit_r169_c127 bl[127] br[127] wl[169] vdd gnd cell_6t
Xbit_r170_c127 bl[127] br[127] wl[170] vdd gnd cell_6t
Xbit_r171_c127 bl[127] br[127] wl[171] vdd gnd cell_6t
Xbit_r172_c127 bl[127] br[127] wl[172] vdd gnd cell_6t
Xbit_r173_c127 bl[127] br[127] wl[173] vdd gnd cell_6t
Xbit_r174_c127 bl[127] br[127] wl[174] vdd gnd cell_6t
Xbit_r175_c127 bl[127] br[127] wl[175] vdd gnd cell_6t
Xbit_r176_c127 bl[127] br[127] wl[176] vdd gnd cell_6t
Xbit_r177_c127 bl[127] br[127] wl[177] vdd gnd cell_6t
Xbit_r178_c127 bl[127] br[127] wl[178] vdd gnd cell_6t
Xbit_r179_c127 bl[127] br[127] wl[179] vdd gnd cell_6t
Xbit_r180_c127 bl[127] br[127] wl[180] vdd gnd cell_6t
Xbit_r181_c127 bl[127] br[127] wl[181] vdd gnd cell_6t
Xbit_r182_c127 bl[127] br[127] wl[182] vdd gnd cell_6t
Xbit_r183_c127 bl[127] br[127] wl[183] vdd gnd cell_6t
Xbit_r184_c127 bl[127] br[127] wl[184] vdd gnd cell_6t
Xbit_r185_c127 bl[127] br[127] wl[185] vdd gnd cell_6t
Xbit_r186_c127 bl[127] br[127] wl[186] vdd gnd cell_6t
Xbit_r187_c127 bl[127] br[127] wl[187] vdd gnd cell_6t
Xbit_r188_c127 bl[127] br[127] wl[188] vdd gnd cell_6t
Xbit_r189_c127 bl[127] br[127] wl[189] vdd gnd cell_6t
Xbit_r190_c127 bl[127] br[127] wl[190] vdd gnd cell_6t
Xbit_r191_c127 bl[127] br[127] wl[191] vdd gnd cell_6t
Xbit_r192_c127 bl[127] br[127] wl[192] vdd gnd cell_6t
Xbit_r193_c127 bl[127] br[127] wl[193] vdd gnd cell_6t
Xbit_r194_c127 bl[127] br[127] wl[194] vdd gnd cell_6t
Xbit_r195_c127 bl[127] br[127] wl[195] vdd gnd cell_6t
Xbit_r196_c127 bl[127] br[127] wl[196] vdd gnd cell_6t
Xbit_r197_c127 bl[127] br[127] wl[197] vdd gnd cell_6t
Xbit_r198_c127 bl[127] br[127] wl[198] vdd gnd cell_6t
Xbit_r199_c127 bl[127] br[127] wl[199] vdd gnd cell_6t
Xbit_r200_c127 bl[127] br[127] wl[200] vdd gnd cell_6t
Xbit_r201_c127 bl[127] br[127] wl[201] vdd gnd cell_6t
Xbit_r202_c127 bl[127] br[127] wl[202] vdd gnd cell_6t
Xbit_r203_c127 bl[127] br[127] wl[203] vdd gnd cell_6t
Xbit_r204_c127 bl[127] br[127] wl[204] vdd gnd cell_6t
Xbit_r205_c127 bl[127] br[127] wl[205] vdd gnd cell_6t
Xbit_r206_c127 bl[127] br[127] wl[206] vdd gnd cell_6t
Xbit_r207_c127 bl[127] br[127] wl[207] vdd gnd cell_6t
Xbit_r208_c127 bl[127] br[127] wl[208] vdd gnd cell_6t
Xbit_r209_c127 bl[127] br[127] wl[209] vdd gnd cell_6t
Xbit_r210_c127 bl[127] br[127] wl[210] vdd gnd cell_6t
Xbit_r211_c127 bl[127] br[127] wl[211] vdd gnd cell_6t
Xbit_r212_c127 bl[127] br[127] wl[212] vdd gnd cell_6t
Xbit_r213_c127 bl[127] br[127] wl[213] vdd gnd cell_6t
Xbit_r214_c127 bl[127] br[127] wl[214] vdd gnd cell_6t
Xbit_r215_c127 bl[127] br[127] wl[215] vdd gnd cell_6t
Xbit_r216_c127 bl[127] br[127] wl[216] vdd gnd cell_6t
Xbit_r217_c127 bl[127] br[127] wl[217] vdd gnd cell_6t
Xbit_r218_c127 bl[127] br[127] wl[218] vdd gnd cell_6t
Xbit_r219_c127 bl[127] br[127] wl[219] vdd gnd cell_6t
Xbit_r220_c127 bl[127] br[127] wl[220] vdd gnd cell_6t
Xbit_r221_c127 bl[127] br[127] wl[221] vdd gnd cell_6t
Xbit_r222_c127 bl[127] br[127] wl[222] vdd gnd cell_6t
Xbit_r223_c127 bl[127] br[127] wl[223] vdd gnd cell_6t
Xbit_r224_c127 bl[127] br[127] wl[224] vdd gnd cell_6t
Xbit_r225_c127 bl[127] br[127] wl[225] vdd gnd cell_6t
Xbit_r226_c127 bl[127] br[127] wl[226] vdd gnd cell_6t
Xbit_r227_c127 bl[127] br[127] wl[227] vdd gnd cell_6t
Xbit_r228_c127 bl[127] br[127] wl[228] vdd gnd cell_6t
Xbit_r229_c127 bl[127] br[127] wl[229] vdd gnd cell_6t
Xbit_r230_c127 bl[127] br[127] wl[230] vdd gnd cell_6t
Xbit_r231_c127 bl[127] br[127] wl[231] vdd gnd cell_6t
Xbit_r232_c127 bl[127] br[127] wl[232] vdd gnd cell_6t
Xbit_r233_c127 bl[127] br[127] wl[233] vdd gnd cell_6t
Xbit_r234_c127 bl[127] br[127] wl[234] vdd gnd cell_6t
Xbit_r235_c127 bl[127] br[127] wl[235] vdd gnd cell_6t
Xbit_r236_c127 bl[127] br[127] wl[236] vdd gnd cell_6t
Xbit_r237_c127 bl[127] br[127] wl[237] vdd gnd cell_6t
Xbit_r238_c127 bl[127] br[127] wl[238] vdd gnd cell_6t
Xbit_r239_c127 bl[127] br[127] wl[239] vdd gnd cell_6t
Xbit_r240_c127 bl[127] br[127] wl[240] vdd gnd cell_6t
Xbit_r241_c127 bl[127] br[127] wl[241] vdd gnd cell_6t
Xbit_r242_c127 bl[127] br[127] wl[242] vdd gnd cell_6t
Xbit_r243_c127 bl[127] br[127] wl[243] vdd gnd cell_6t
Xbit_r244_c127 bl[127] br[127] wl[244] vdd gnd cell_6t
Xbit_r245_c127 bl[127] br[127] wl[245] vdd gnd cell_6t
Xbit_r246_c127 bl[127] br[127] wl[246] vdd gnd cell_6t
Xbit_r247_c127 bl[127] br[127] wl[247] vdd gnd cell_6t
Xbit_r248_c127 bl[127] br[127] wl[248] vdd gnd cell_6t
Xbit_r249_c127 bl[127] br[127] wl[249] vdd gnd cell_6t
Xbit_r250_c127 bl[127] br[127] wl[250] vdd gnd cell_6t
Xbit_r251_c127 bl[127] br[127] wl[251] vdd gnd cell_6t
Xbit_r252_c127 bl[127] br[127] wl[252] vdd gnd cell_6t
Xbit_r253_c127 bl[127] br[127] wl[253] vdd gnd cell_6t
Xbit_r254_c127 bl[127] br[127] wl[254] vdd gnd cell_6t
Xbit_r255_c127 bl[127] br[127] wl[255] vdd gnd cell_6t
Xbit_r0_c128 bl[128] br[128] wl[0] vdd gnd cell_6t
Xbit_r1_c128 bl[128] br[128] wl[1] vdd gnd cell_6t
Xbit_r2_c128 bl[128] br[128] wl[2] vdd gnd cell_6t
Xbit_r3_c128 bl[128] br[128] wl[3] vdd gnd cell_6t
Xbit_r4_c128 bl[128] br[128] wl[4] vdd gnd cell_6t
Xbit_r5_c128 bl[128] br[128] wl[5] vdd gnd cell_6t
Xbit_r6_c128 bl[128] br[128] wl[6] vdd gnd cell_6t
Xbit_r7_c128 bl[128] br[128] wl[7] vdd gnd cell_6t
Xbit_r8_c128 bl[128] br[128] wl[8] vdd gnd cell_6t
Xbit_r9_c128 bl[128] br[128] wl[9] vdd gnd cell_6t
Xbit_r10_c128 bl[128] br[128] wl[10] vdd gnd cell_6t
Xbit_r11_c128 bl[128] br[128] wl[11] vdd gnd cell_6t
Xbit_r12_c128 bl[128] br[128] wl[12] vdd gnd cell_6t
Xbit_r13_c128 bl[128] br[128] wl[13] vdd gnd cell_6t
Xbit_r14_c128 bl[128] br[128] wl[14] vdd gnd cell_6t
Xbit_r15_c128 bl[128] br[128] wl[15] vdd gnd cell_6t
Xbit_r16_c128 bl[128] br[128] wl[16] vdd gnd cell_6t
Xbit_r17_c128 bl[128] br[128] wl[17] vdd gnd cell_6t
Xbit_r18_c128 bl[128] br[128] wl[18] vdd gnd cell_6t
Xbit_r19_c128 bl[128] br[128] wl[19] vdd gnd cell_6t
Xbit_r20_c128 bl[128] br[128] wl[20] vdd gnd cell_6t
Xbit_r21_c128 bl[128] br[128] wl[21] vdd gnd cell_6t
Xbit_r22_c128 bl[128] br[128] wl[22] vdd gnd cell_6t
Xbit_r23_c128 bl[128] br[128] wl[23] vdd gnd cell_6t
Xbit_r24_c128 bl[128] br[128] wl[24] vdd gnd cell_6t
Xbit_r25_c128 bl[128] br[128] wl[25] vdd gnd cell_6t
Xbit_r26_c128 bl[128] br[128] wl[26] vdd gnd cell_6t
Xbit_r27_c128 bl[128] br[128] wl[27] vdd gnd cell_6t
Xbit_r28_c128 bl[128] br[128] wl[28] vdd gnd cell_6t
Xbit_r29_c128 bl[128] br[128] wl[29] vdd gnd cell_6t
Xbit_r30_c128 bl[128] br[128] wl[30] vdd gnd cell_6t
Xbit_r31_c128 bl[128] br[128] wl[31] vdd gnd cell_6t
Xbit_r32_c128 bl[128] br[128] wl[32] vdd gnd cell_6t
Xbit_r33_c128 bl[128] br[128] wl[33] vdd gnd cell_6t
Xbit_r34_c128 bl[128] br[128] wl[34] vdd gnd cell_6t
Xbit_r35_c128 bl[128] br[128] wl[35] vdd gnd cell_6t
Xbit_r36_c128 bl[128] br[128] wl[36] vdd gnd cell_6t
Xbit_r37_c128 bl[128] br[128] wl[37] vdd gnd cell_6t
Xbit_r38_c128 bl[128] br[128] wl[38] vdd gnd cell_6t
Xbit_r39_c128 bl[128] br[128] wl[39] vdd gnd cell_6t
Xbit_r40_c128 bl[128] br[128] wl[40] vdd gnd cell_6t
Xbit_r41_c128 bl[128] br[128] wl[41] vdd gnd cell_6t
Xbit_r42_c128 bl[128] br[128] wl[42] vdd gnd cell_6t
Xbit_r43_c128 bl[128] br[128] wl[43] vdd gnd cell_6t
Xbit_r44_c128 bl[128] br[128] wl[44] vdd gnd cell_6t
Xbit_r45_c128 bl[128] br[128] wl[45] vdd gnd cell_6t
Xbit_r46_c128 bl[128] br[128] wl[46] vdd gnd cell_6t
Xbit_r47_c128 bl[128] br[128] wl[47] vdd gnd cell_6t
Xbit_r48_c128 bl[128] br[128] wl[48] vdd gnd cell_6t
Xbit_r49_c128 bl[128] br[128] wl[49] vdd gnd cell_6t
Xbit_r50_c128 bl[128] br[128] wl[50] vdd gnd cell_6t
Xbit_r51_c128 bl[128] br[128] wl[51] vdd gnd cell_6t
Xbit_r52_c128 bl[128] br[128] wl[52] vdd gnd cell_6t
Xbit_r53_c128 bl[128] br[128] wl[53] vdd gnd cell_6t
Xbit_r54_c128 bl[128] br[128] wl[54] vdd gnd cell_6t
Xbit_r55_c128 bl[128] br[128] wl[55] vdd gnd cell_6t
Xbit_r56_c128 bl[128] br[128] wl[56] vdd gnd cell_6t
Xbit_r57_c128 bl[128] br[128] wl[57] vdd gnd cell_6t
Xbit_r58_c128 bl[128] br[128] wl[58] vdd gnd cell_6t
Xbit_r59_c128 bl[128] br[128] wl[59] vdd gnd cell_6t
Xbit_r60_c128 bl[128] br[128] wl[60] vdd gnd cell_6t
Xbit_r61_c128 bl[128] br[128] wl[61] vdd gnd cell_6t
Xbit_r62_c128 bl[128] br[128] wl[62] vdd gnd cell_6t
Xbit_r63_c128 bl[128] br[128] wl[63] vdd gnd cell_6t
Xbit_r64_c128 bl[128] br[128] wl[64] vdd gnd cell_6t
Xbit_r65_c128 bl[128] br[128] wl[65] vdd gnd cell_6t
Xbit_r66_c128 bl[128] br[128] wl[66] vdd gnd cell_6t
Xbit_r67_c128 bl[128] br[128] wl[67] vdd gnd cell_6t
Xbit_r68_c128 bl[128] br[128] wl[68] vdd gnd cell_6t
Xbit_r69_c128 bl[128] br[128] wl[69] vdd gnd cell_6t
Xbit_r70_c128 bl[128] br[128] wl[70] vdd gnd cell_6t
Xbit_r71_c128 bl[128] br[128] wl[71] vdd gnd cell_6t
Xbit_r72_c128 bl[128] br[128] wl[72] vdd gnd cell_6t
Xbit_r73_c128 bl[128] br[128] wl[73] vdd gnd cell_6t
Xbit_r74_c128 bl[128] br[128] wl[74] vdd gnd cell_6t
Xbit_r75_c128 bl[128] br[128] wl[75] vdd gnd cell_6t
Xbit_r76_c128 bl[128] br[128] wl[76] vdd gnd cell_6t
Xbit_r77_c128 bl[128] br[128] wl[77] vdd gnd cell_6t
Xbit_r78_c128 bl[128] br[128] wl[78] vdd gnd cell_6t
Xbit_r79_c128 bl[128] br[128] wl[79] vdd gnd cell_6t
Xbit_r80_c128 bl[128] br[128] wl[80] vdd gnd cell_6t
Xbit_r81_c128 bl[128] br[128] wl[81] vdd gnd cell_6t
Xbit_r82_c128 bl[128] br[128] wl[82] vdd gnd cell_6t
Xbit_r83_c128 bl[128] br[128] wl[83] vdd gnd cell_6t
Xbit_r84_c128 bl[128] br[128] wl[84] vdd gnd cell_6t
Xbit_r85_c128 bl[128] br[128] wl[85] vdd gnd cell_6t
Xbit_r86_c128 bl[128] br[128] wl[86] vdd gnd cell_6t
Xbit_r87_c128 bl[128] br[128] wl[87] vdd gnd cell_6t
Xbit_r88_c128 bl[128] br[128] wl[88] vdd gnd cell_6t
Xbit_r89_c128 bl[128] br[128] wl[89] vdd gnd cell_6t
Xbit_r90_c128 bl[128] br[128] wl[90] vdd gnd cell_6t
Xbit_r91_c128 bl[128] br[128] wl[91] vdd gnd cell_6t
Xbit_r92_c128 bl[128] br[128] wl[92] vdd gnd cell_6t
Xbit_r93_c128 bl[128] br[128] wl[93] vdd gnd cell_6t
Xbit_r94_c128 bl[128] br[128] wl[94] vdd gnd cell_6t
Xbit_r95_c128 bl[128] br[128] wl[95] vdd gnd cell_6t
Xbit_r96_c128 bl[128] br[128] wl[96] vdd gnd cell_6t
Xbit_r97_c128 bl[128] br[128] wl[97] vdd gnd cell_6t
Xbit_r98_c128 bl[128] br[128] wl[98] vdd gnd cell_6t
Xbit_r99_c128 bl[128] br[128] wl[99] vdd gnd cell_6t
Xbit_r100_c128 bl[128] br[128] wl[100] vdd gnd cell_6t
Xbit_r101_c128 bl[128] br[128] wl[101] vdd gnd cell_6t
Xbit_r102_c128 bl[128] br[128] wl[102] vdd gnd cell_6t
Xbit_r103_c128 bl[128] br[128] wl[103] vdd gnd cell_6t
Xbit_r104_c128 bl[128] br[128] wl[104] vdd gnd cell_6t
Xbit_r105_c128 bl[128] br[128] wl[105] vdd gnd cell_6t
Xbit_r106_c128 bl[128] br[128] wl[106] vdd gnd cell_6t
Xbit_r107_c128 bl[128] br[128] wl[107] vdd gnd cell_6t
Xbit_r108_c128 bl[128] br[128] wl[108] vdd gnd cell_6t
Xbit_r109_c128 bl[128] br[128] wl[109] vdd gnd cell_6t
Xbit_r110_c128 bl[128] br[128] wl[110] vdd gnd cell_6t
Xbit_r111_c128 bl[128] br[128] wl[111] vdd gnd cell_6t
Xbit_r112_c128 bl[128] br[128] wl[112] vdd gnd cell_6t
Xbit_r113_c128 bl[128] br[128] wl[113] vdd gnd cell_6t
Xbit_r114_c128 bl[128] br[128] wl[114] vdd gnd cell_6t
Xbit_r115_c128 bl[128] br[128] wl[115] vdd gnd cell_6t
Xbit_r116_c128 bl[128] br[128] wl[116] vdd gnd cell_6t
Xbit_r117_c128 bl[128] br[128] wl[117] vdd gnd cell_6t
Xbit_r118_c128 bl[128] br[128] wl[118] vdd gnd cell_6t
Xbit_r119_c128 bl[128] br[128] wl[119] vdd gnd cell_6t
Xbit_r120_c128 bl[128] br[128] wl[120] vdd gnd cell_6t
Xbit_r121_c128 bl[128] br[128] wl[121] vdd gnd cell_6t
Xbit_r122_c128 bl[128] br[128] wl[122] vdd gnd cell_6t
Xbit_r123_c128 bl[128] br[128] wl[123] vdd gnd cell_6t
Xbit_r124_c128 bl[128] br[128] wl[124] vdd gnd cell_6t
Xbit_r125_c128 bl[128] br[128] wl[125] vdd gnd cell_6t
Xbit_r126_c128 bl[128] br[128] wl[126] vdd gnd cell_6t
Xbit_r127_c128 bl[128] br[128] wl[127] vdd gnd cell_6t
Xbit_r128_c128 bl[128] br[128] wl[128] vdd gnd cell_6t
Xbit_r129_c128 bl[128] br[128] wl[129] vdd gnd cell_6t
Xbit_r130_c128 bl[128] br[128] wl[130] vdd gnd cell_6t
Xbit_r131_c128 bl[128] br[128] wl[131] vdd gnd cell_6t
Xbit_r132_c128 bl[128] br[128] wl[132] vdd gnd cell_6t
Xbit_r133_c128 bl[128] br[128] wl[133] vdd gnd cell_6t
Xbit_r134_c128 bl[128] br[128] wl[134] vdd gnd cell_6t
Xbit_r135_c128 bl[128] br[128] wl[135] vdd gnd cell_6t
Xbit_r136_c128 bl[128] br[128] wl[136] vdd gnd cell_6t
Xbit_r137_c128 bl[128] br[128] wl[137] vdd gnd cell_6t
Xbit_r138_c128 bl[128] br[128] wl[138] vdd gnd cell_6t
Xbit_r139_c128 bl[128] br[128] wl[139] vdd gnd cell_6t
Xbit_r140_c128 bl[128] br[128] wl[140] vdd gnd cell_6t
Xbit_r141_c128 bl[128] br[128] wl[141] vdd gnd cell_6t
Xbit_r142_c128 bl[128] br[128] wl[142] vdd gnd cell_6t
Xbit_r143_c128 bl[128] br[128] wl[143] vdd gnd cell_6t
Xbit_r144_c128 bl[128] br[128] wl[144] vdd gnd cell_6t
Xbit_r145_c128 bl[128] br[128] wl[145] vdd gnd cell_6t
Xbit_r146_c128 bl[128] br[128] wl[146] vdd gnd cell_6t
Xbit_r147_c128 bl[128] br[128] wl[147] vdd gnd cell_6t
Xbit_r148_c128 bl[128] br[128] wl[148] vdd gnd cell_6t
Xbit_r149_c128 bl[128] br[128] wl[149] vdd gnd cell_6t
Xbit_r150_c128 bl[128] br[128] wl[150] vdd gnd cell_6t
Xbit_r151_c128 bl[128] br[128] wl[151] vdd gnd cell_6t
Xbit_r152_c128 bl[128] br[128] wl[152] vdd gnd cell_6t
Xbit_r153_c128 bl[128] br[128] wl[153] vdd gnd cell_6t
Xbit_r154_c128 bl[128] br[128] wl[154] vdd gnd cell_6t
Xbit_r155_c128 bl[128] br[128] wl[155] vdd gnd cell_6t
Xbit_r156_c128 bl[128] br[128] wl[156] vdd gnd cell_6t
Xbit_r157_c128 bl[128] br[128] wl[157] vdd gnd cell_6t
Xbit_r158_c128 bl[128] br[128] wl[158] vdd gnd cell_6t
Xbit_r159_c128 bl[128] br[128] wl[159] vdd gnd cell_6t
Xbit_r160_c128 bl[128] br[128] wl[160] vdd gnd cell_6t
Xbit_r161_c128 bl[128] br[128] wl[161] vdd gnd cell_6t
Xbit_r162_c128 bl[128] br[128] wl[162] vdd gnd cell_6t
Xbit_r163_c128 bl[128] br[128] wl[163] vdd gnd cell_6t
Xbit_r164_c128 bl[128] br[128] wl[164] vdd gnd cell_6t
Xbit_r165_c128 bl[128] br[128] wl[165] vdd gnd cell_6t
Xbit_r166_c128 bl[128] br[128] wl[166] vdd gnd cell_6t
Xbit_r167_c128 bl[128] br[128] wl[167] vdd gnd cell_6t
Xbit_r168_c128 bl[128] br[128] wl[168] vdd gnd cell_6t
Xbit_r169_c128 bl[128] br[128] wl[169] vdd gnd cell_6t
Xbit_r170_c128 bl[128] br[128] wl[170] vdd gnd cell_6t
Xbit_r171_c128 bl[128] br[128] wl[171] vdd gnd cell_6t
Xbit_r172_c128 bl[128] br[128] wl[172] vdd gnd cell_6t
Xbit_r173_c128 bl[128] br[128] wl[173] vdd gnd cell_6t
Xbit_r174_c128 bl[128] br[128] wl[174] vdd gnd cell_6t
Xbit_r175_c128 bl[128] br[128] wl[175] vdd gnd cell_6t
Xbit_r176_c128 bl[128] br[128] wl[176] vdd gnd cell_6t
Xbit_r177_c128 bl[128] br[128] wl[177] vdd gnd cell_6t
Xbit_r178_c128 bl[128] br[128] wl[178] vdd gnd cell_6t
Xbit_r179_c128 bl[128] br[128] wl[179] vdd gnd cell_6t
Xbit_r180_c128 bl[128] br[128] wl[180] vdd gnd cell_6t
Xbit_r181_c128 bl[128] br[128] wl[181] vdd gnd cell_6t
Xbit_r182_c128 bl[128] br[128] wl[182] vdd gnd cell_6t
Xbit_r183_c128 bl[128] br[128] wl[183] vdd gnd cell_6t
Xbit_r184_c128 bl[128] br[128] wl[184] vdd gnd cell_6t
Xbit_r185_c128 bl[128] br[128] wl[185] vdd gnd cell_6t
Xbit_r186_c128 bl[128] br[128] wl[186] vdd gnd cell_6t
Xbit_r187_c128 bl[128] br[128] wl[187] vdd gnd cell_6t
Xbit_r188_c128 bl[128] br[128] wl[188] vdd gnd cell_6t
Xbit_r189_c128 bl[128] br[128] wl[189] vdd gnd cell_6t
Xbit_r190_c128 bl[128] br[128] wl[190] vdd gnd cell_6t
Xbit_r191_c128 bl[128] br[128] wl[191] vdd gnd cell_6t
Xbit_r192_c128 bl[128] br[128] wl[192] vdd gnd cell_6t
Xbit_r193_c128 bl[128] br[128] wl[193] vdd gnd cell_6t
Xbit_r194_c128 bl[128] br[128] wl[194] vdd gnd cell_6t
Xbit_r195_c128 bl[128] br[128] wl[195] vdd gnd cell_6t
Xbit_r196_c128 bl[128] br[128] wl[196] vdd gnd cell_6t
Xbit_r197_c128 bl[128] br[128] wl[197] vdd gnd cell_6t
Xbit_r198_c128 bl[128] br[128] wl[198] vdd gnd cell_6t
Xbit_r199_c128 bl[128] br[128] wl[199] vdd gnd cell_6t
Xbit_r200_c128 bl[128] br[128] wl[200] vdd gnd cell_6t
Xbit_r201_c128 bl[128] br[128] wl[201] vdd gnd cell_6t
Xbit_r202_c128 bl[128] br[128] wl[202] vdd gnd cell_6t
Xbit_r203_c128 bl[128] br[128] wl[203] vdd gnd cell_6t
Xbit_r204_c128 bl[128] br[128] wl[204] vdd gnd cell_6t
Xbit_r205_c128 bl[128] br[128] wl[205] vdd gnd cell_6t
Xbit_r206_c128 bl[128] br[128] wl[206] vdd gnd cell_6t
Xbit_r207_c128 bl[128] br[128] wl[207] vdd gnd cell_6t
Xbit_r208_c128 bl[128] br[128] wl[208] vdd gnd cell_6t
Xbit_r209_c128 bl[128] br[128] wl[209] vdd gnd cell_6t
Xbit_r210_c128 bl[128] br[128] wl[210] vdd gnd cell_6t
Xbit_r211_c128 bl[128] br[128] wl[211] vdd gnd cell_6t
Xbit_r212_c128 bl[128] br[128] wl[212] vdd gnd cell_6t
Xbit_r213_c128 bl[128] br[128] wl[213] vdd gnd cell_6t
Xbit_r214_c128 bl[128] br[128] wl[214] vdd gnd cell_6t
Xbit_r215_c128 bl[128] br[128] wl[215] vdd gnd cell_6t
Xbit_r216_c128 bl[128] br[128] wl[216] vdd gnd cell_6t
Xbit_r217_c128 bl[128] br[128] wl[217] vdd gnd cell_6t
Xbit_r218_c128 bl[128] br[128] wl[218] vdd gnd cell_6t
Xbit_r219_c128 bl[128] br[128] wl[219] vdd gnd cell_6t
Xbit_r220_c128 bl[128] br[128] wl[220] vdd gnd cell_6t
Xbit_r221_c128 bl[128] br[128] wl[221] vdd gnd cell_6t
Xbit_r222_c128 bl[128] br[128] wl[222] vdd gnd cell_6t
Xbit_r223_c128 bl[128] br[128] wl[223] vdd gnd cell_6t
Xbit_r224_c128 bl[128] br[128] wl[224] vdd gnd cell_6t
Xbit_r225_c128 bl[128] br[128] wl[225] vdd gnd cell_6t
Xbit_r226_c128 bl[128] br[128] wl[226] vdd gnd cell_6t
Xbit_r227_c128 bl[128] br[128] wl[227] vdd gnd cell_6t
Xbit_r228_c128 bl[128] br[128] wl[228] vdd gnd cell_6t
Xbit_r229_c128 bl[128] br[128] wl[229] vdd gnd cell_6t
Xbit_r230_c128 bl[128] br[128] wl[230] vdd gnd cell_6t
Xbit_r231_c128 bl[128] br[128] wl[231] vdd gnd cell_6t
Xbit_r232_c128 bl[128] br[128] wl[232] vdd gnd cell_6t
Xbit_r233_c128 bl[128] br[128] wl[233] vdd gnd cell_6t
Xbit_r234_c128 bl[128] br[128] wl[234] vdd gnd cell_6t
Xbit_r235_c128 bl[128] br[128] wl[235] vdd gnd cell_6t
Xbit_r236_c128 bl[128] br[128] wl[236] vdd gnd cell_6t
Xbit_r237_c128 bl[128] br[128] wl[237] vdd gnd cell_6t
Xbit_r238_c128 bl[128] br[128] wl[238] vdd gnd cell_6t
Xbit_r239_c128 bl[128] br[128] wl[239] vdd gnd cell_6t
Xbit_r240_c128 bl[128] br[128] wl[240] vdd gnd cell_6t
Xbit_r241_c128 bl[128] br[128] wl[241] vdd gnd cell_6t
Xbit_r242_c128 bl[128] br[128] wl[242] vdd gnd cell_6t
Xbit_r243_c128 bl[128] br[128] wl[243] vdd gnd cell_6t
Xbit_r244_c128 bl[128] br[128] wl[244] vdd gnd cell_6t
Xbit_r245_c128 bl[128] br[128] wl[245] vdd gnd cell_6t
Xbit_r246_c128 bl[128] br[128] wl[246] vdd gnd cell_6t
Xbit_r247_c128 bl[128] br[128] wl[247] vdd gnd cell_6t
Xbit_r248_c128 bl[128] br[128] wl[248] vdd gnd cell_6t
Xbit_r249_c128 bl[128] br[128] wl[249] vdd gnd cell_6t
Xbit_r250_c128 bl[128] br[128] wl[250] vdd gnd cell_6t
Xbit_r251_c128 bl[128] br[128] wl[251] vdd gnd cell_6t
Xbit_r252_c128 bl[128] br[128] wl[252] vdd gnd cell_6t
Xbit_r253_c128 bl[128] br[128] wl[253] vdd gnd cell_6t
Xbit_r254_c128 bl[128] br[128] wl[254] vdd gnd cell_6t
Xbit_r255_c128 bl[128] br[128] wl[255] vdd gnd cell_6t
Xbit_r0_c129 bl[129] br[129] wl[0] vdd gnd cell_6t
Xbit_r1_c129 bl[129] br[129] wl[1] vdd gnd cell_6t
Xbit_r2_c129 bl[129] br[129] wl[2] vdd gnd cell_6t
Xbit_r3_c129 bl[129] br[129] wl[3] vdd gnd cell_6t
Xbit_r4_c129 bl[129] br[129] wl[4] vdd gnd cell_6t
Xbit_r5_c129 bl[129] br[129] wl[5] vdd gnd cell_6t
Xbit_r6_c129 bl[129] br[129] wl[6] vdd gnd cell_6t
Xbit_r7_c129 bl[129] br[129] wl[7] vdd gnd cell_6t
Xbit_r8_c129 bl[129] br[129] wl[8] vdd gnd cell_6t
Xbit_r9_c129 bl[129] br[129] wl[9] vdd gnd cell_6t
Xbit_r10_c129 bl[129] br[129] wl[10] vdd gnd cell_6t
Xbit_r11_c129 bl[129] br[129] wl[11] vdd gnd cell_6t
Xbit_r12_c129 bl[129] br[129] wl[12] vdd gnd cell_6t
Xbit_r13_c129 bl[129] br[129] wl[13] vdd gnd cell_6t
Xbit_r14_c129 bl[129] br[129] wl[14] vdd gnd cell_6t
Xbit_r15_c129 bl[129] br[129] wl[15] vdd gnd cell_6t
Xbit_r16_c129 bl[129] br[129] wl[16] vdd gnd cell_6t
Xbit_r17_c129 bl[129] br[129] wl[17] vdd gnd cell_6t
Xbit_r18_c129 bl[129] br[129] wl[18] vdd gnd cell_6t
Xbit_r19_c129 bl[129] br[129] wl[19] vdd gnd cell_6t
Xbit_r20_c129 bl[129] br[129] wl[20] vdd gnd cell_6t
Xbit_r21_c129 bl[129] br[129] wl[21] vdd gnd cell_6t
Xbit_r22_c129 bl[129] br[129] wl[22] vdd gnd cell_6t
Xbit_r23_c129 bl[129] br[129] wl[23] vdd gnd cell_6t
Xbit_r24_c129 bl[129] br[129] wl[24] vdd gnd cell_6t
Xbit_r25_c129 bl[129] br[129] wl[25] vdd gnd cell_6t
Xbit_r26_c129 bl[129] br[129] wl[26] vdd gnd cell_6t
Xbit_r27_c129 bl[129] br[129] wl[27] vdd gnd cell_6t
Xbit_r28_c129 bl[129] br[129] wl[28] vdd gnd cell_6t
Xbit_r29_c129 bl[129] br[129] wl[29] vdd gnd cell_6t
Xbit_r30_c129 bl[129] br[129] wl[30] vdd gnd cell_6t
Xbit_r31_c129 bl[129] br[129] wl[31] vdd gnd cell_6t
Xbit_r32_c129 bl[129] br[129] wl[32] vdd gnd cell_6t
Xbit_r33_c129 bl[129] br[129] wl[33] vdd gnd cell_6t
Xbit_r34_c129 bl[129] br[129] wl[34] vdd gnd cell_6t
Xbit_r35_c129 bl[129] br[129] wl[35] vdd gnd cell_6t
Xbit_r36_c129 bl[129] br[129] wl[36] vdd gnd cell_6t
Xbit_r37_c129 bl[129] br[129] wl[37] vdd gnd cell_6t
Xbit_r38_c129 bl[129] br[129] wl[38] vdd gnd cell_6t
Xbit_r39_c129 bl[129] br[129] wl[39] vdd gnd cell_6t
Xbit_r40_c129 bl[129] br[129] wl[40] vdd gnd cell_6t
Xbit_r41_c129 bl[129] br[129] wl[41] vdd gnd cell_6t
Xbit_r42_c129 bl[129] br[129] wl[42] vdd gnd cell_6t
Xbit_r43_c129 bl[129] br[129] wl[43] vdd gnd cell_6t
Xbit_r44_c129 bl[129] br[129] wl[44] vdd gnd cell_6t
Xbit_r45_c129 bl[129] br[129] wl[45] vdd gnd cell_6t
Xbit_r46_c129 bl[129] br[129] wl[46] vdd gnd cell_6t
Xbit_r47_c129 bl[129] br[129] wl[47] vdd gnd cell_6t
Xbit_r48_c129 bl[129] br[129] wl[48] vdd gnd cell_6t
Xbit_r49_c129 bl[129] br[129] wl[49] vdd gnd cell_6t
Xbit_r50_c129 bl[129] br[129] wl[50] vdd gnd cell_6t
Xbit_r51_c129 bl[129] br[129] wl[51] vdd gnd cell_6t
Xbit_r52_c129 bl[129] br[129] wl[52] vdd gnd cell_6t
Xbit_r53_c129 bl[129] br[129] wl[53] vdd gnd cell_6t
Xbit_r54_c129 bl[129] br[129] wl[54] vdd gnd cell_6t
Xbit_r55_c129 bl[129] br[129] wl[55] vdd gnd cell_6t
Xbit_r56_c129 bl[129] br[129] wl[56] vdd gnd cell_6t
Xbit_r57_c129 bl[129] br[129] wl[57] vdd gnd cell_6t
Xbit_r58_c129 bl[129] br[129] wl[58] vdd gnd cell_6t
Xbit_r59_c129 bl[129] br[129] wl[59] vdd gnd cell_6t
Xbit_r60_c129 bl[129] br[129] wl[60] vdd gnd cell_6t
Xbit_r61_c129 bl[129] br[129] wl[61] vdd gnd cell_6t
Xbit_r62_c129 bl[129] br[129] wl[62] vdd gnd cell_6t
Xbit_r63_c129 bl[129] br[129] wl[63] vdd gnd cell_6t
Xbit_r64_c129 bl[129] br[129] wl[64] vdd gnd cell_6t
Xbit_r65_c129 bl[129] br[129] wl[65] vdd gnd cell_6t
Xbit_r66_c129 bl[129] br[129] wl[66] vdd gnd cell_6t
Xbit_r67_c129 bl[129] br[129] wl[67] vdd gnd cell_6t
Xbit_r68_c129 bl[129] br[129] wl[68] vdd gnd cell_6t
Xbit_r69_c129 bl[129] br[129] wl[69] vdd gnd cell_6t
Xbit_r70_c129 bl[129] br[129] wl[70] vdd gnd cell_6t
Xbit_r71_c129 bl[129] br[129] wl[71] vdd gnd cell_6t
Xbit_r72_c129 bl[129] br[129] wl[72] vdd gnd cell_6t
Xbit_r73_c129 bl[129] br[129] wl[73] vdd gnd cell_6t
Xbit_r74_c129 bl[129] br[129] wl[74] vdd gnd cell_6t
Xbit_r75_c129 bl[129] br[129] wl[75] vdd gnd cell_6t
Xbit_r76_c129 bl[129] br[129] wl[76] vdd gnd cell_6t
Xbit_r77_c129 bl[129] br[129] wl[77] vdd gnd cell_6t
Xbit_r78_c129 bl[129] br[129] wl[78] vdd gnd cell_6t
Xbit_r79_c129 bl[129] br[129] wl[79] vdd gnd cell_6t
Xbit_r80_c129 bl[129] br[129] wl[80] vdd gnd cell_6t
Xbit_r81_c129 bl[129] br[129] wl[81] vdd gnd cell_6t
Xbit_r82_c129 bl[129] br[129] wl[82] vdd gnd cell_6t
Xbit_r83_c129 bl[129] br[129] wl[83] vdd gnd cell_6t
Xbit_r84_c129 bl[129] br[129] wl[84] vdd gnd cell_6t
Xbit_r85_c129 bl[129] br[129] wl[85] vdd gnd cell_6t
Xbit_r86_c129 bl[129] br[129] wl[86] vdd gnd cell_6t
Xbit_r87_c129 bl[129] br[129] wl[87] vdd gnd cell_6t
Xbit_r88_c129 bl[129] br[129] wl[88] vdd gnd cell_6t
Xbit_r89_c129 bl[129] br[129] wl[89] vdd gnd cell_6t
Xbit_r90_c129 bl[129] br[129] wl[90] vdd gnd cell_6t
Xbit_r91_c129 bl[129] br[129] wl[91] vdd gnd cell_6t
Xbit_r92_c129 bl[129] br[129] wl[92] vdd gnd cell_6t
Xbit_r93_c129 bl[129] br[129] wl[93] vdd gnd cell_6t
Xbit_r94_c129 bl[129] br[129] wl[94] vdd gnd cell_6t
Xbit_r95_c129 bl[129] br[129] wl[95] vdd gnd cell_6t
Xbit_r96_c129 bl[129] br[129] wl[96] vdd gnd cell_6t
Xbit_r97_c129 bl[129] br[129] wl[97] vdd gnd cell_6t
Xbit_r98_c129 bl[129] br[129] wl[98] vdd gnd cell_6t
Xbit_r99_c129 bl[129] br[129] wl[99] vdd gnd cell_6t
Xbit_r100_c129 bl[129] br[129] wl[100] vdd gnd cell_6t
Xbit_r101_c129 bl[129] br[129] wl[101] vdd gnd cell_6t
Xbit_r102_c129 bl[129] br[129] wl[102] vdd gnd cell_6t
Xbit_r103_c129 bl[129] br[129] wl[103] vdd gnd cell_6t
Xbit_r104_c129 bl[129] br[129] wl[104] vdd gnd cell_6t
Xbit_r105_c129 bl[129] br[129] wl[105] vdd gnd cell_6t
Xbit_r106_c129 bl[129] br[129] wl[106] vdd gnd cell_6t
Xbit_r107_c129 bl[129] br[129] wl[107] vdd gnd cell_6t
Xbit_r108_c129 bl[129] br[129] wl[108] vdd gnd cell_6t
Xbit_r109_c129 bl[129] br[129] wl[109] vdd gnd cell_6t
Xbit_r110_c129 bl[129] br[129] wl[110] vdd gnd cell_6t
Xbit_r111_c129 bl[129] br[129] wl[111] vdd gnd cell_6t
Xbit_r112_c129 bl[129] br[129] wl[112] vdd gnd cell_6t
Xbit_r113_c129 bl[129] br[129] wl[113] vdd gnd cell_6t
Xbit_r114_c129 bl[129] br[129] wl[114] vdd gnd cell_6t
Xbit_r115_c129 bl[129] br[129] wl[115] vdd gnd cell_6t
Xbit_r116_c129 bl[129] br[129] wl[116] vdd gnd cell_6t
Xbit_r117_c129 bl[129] br[129] wl[117] vdd gnd cell_6t
Xbit_r118_c129 bl[129] br[129] wl[118] vdd gnd cell_6t
Xbit_r119_c129 bl[129] br[129] wl[119] vdd gnd cell_6t
Xbit_r120_c129 bl[129] br[129] wl[120] vdd gnd cell_6t
Xbit_r121_c129 bl[129] br[129] wl[121] vdd gnd cell_6t
Xbit_r122_c129 bl[129] br[129] wl[122] vdd gnd cell_6t
Xbit_r123_c129 bl[129] br[129] wl[123] vdd gnd cell_6t
Xbit_r124_c129 bl[129] br[129] wl[124] vdd gnd cell_6t
Xbit_r125_c129 bl[129] br[129] wl[125] vdd gnd cell_6t
Xbit_r126_c129 bl[129] br[129] wl[126] vdd gnd cell_6t
Xbit_r127_c129 bl[129] br[129] wl[127] vdd gnd cell_6t
Xbit_r128_c129 bl[129] br[129] wl[128] vdd gnd cell_6t
Xbit_r129_c129 bl[129] br[129] wl[129] vdd gnd cell_6t
Xbit_r130_c129 bl[129] br[129] wl[130] vdd gnd cell_6t
Xbit_r131_c129 bl[129] br[129] wl[131] vdd gnd cell_6t
Xbit_r132_c129 bl[129] br[129] wl[132] vdd gnd cell_6t
Xbit_r133_c129 bl[129] br[129] wl[133] vdd gnd cell_6t
Xbit_r134_c129 bl[129] br[129] wl[134] vdd gnd cell_6t
Xbit_r135_c129 bl[129] br[129] wl[135] vdd gnd cell_6t
Xbit_r136_c129 bl[129] br[129] wl[136] vdd gnd cell_6t
Xbit_r137_c129 bl[129] br[129] wl[137] vdd gnd cell_6t
Xbit_r138_c129 bl[129] br[129] wl[138] vdd gnd cell_6t
Xbit_r139_c129 bl[129] br[129] wl[139] vdd gnd cell_6t
Xbit_r140_c129 bl[129] br[129] wl[140] vdd gnd cell_6t
Xbit_r141_c129 bl[129] br[129] wl[141] vdd gnd cell_6t
Xbit_r142_c129 bl[129] br[129] wl[142] vdd gnd cell_6t
Xbit_r143_c129 bl[129] br[129] wl[143] vdd gnd cell_6t
Xbit_r144_c129 bl[129] br[129] wl[144] vdd gnd cell_6t
Xbit_r145_c129 bl[129] br[129] wl[145] vdd gnd cell_6t
Xbit_r146_c129 bl[129] br[129] wl[146] vdd gnd cell_6t
Xbit_r147_c129 bl[129] br[129] wl[147] vdd gnd cell_6t
Xbit_r148_c129 bl[129] br[129] wl[148] vdd gnd cell_6t
Xbit_r149_c129 bl[129] br[129] wl[149] vdd gnd cell_6t
Xbit_r150_c129 bl[129] br[129] wl[150] vdd gnd cell_6t
Xbit_r151_c129 bl[129] br[129] wl[151] vdd gnd cell_6t
Xbit_r152_c129 bl[129] br[129] wl[152] vdd gnd cell_6t
Xbit_r153_c129 bl[129] br[129] wl[153] vdd gnd cell_6t
Xbit_r154_c129 bl[129] br[129] wl[154] vdd gnd cell_6t
Xbit_r155_c129 bl[129] br[129] wl[155] vdd gnd cell_6t
Xbit_r156_c129 bl[129] br[129] wl[156] vdd gnd cell_6t
Xbit_r157_c129 bl[129] br[129] wl[157] vdd gnd cell_6t
Xbit_r158_c129 bl[129] br[129] wl[158] vdd gnd cell_6t
Xbit_r159_c129 bl[129] br[129] wl[159] vdd gnd cell_6t
Xbit_r160_c129 bl[129] br[129] wl[160] vdd gnd cell_6t
Xbit_r161_c129 bl[129] br[129] wl[161] vdd gnd cell_6t
Xbit_r162_c129 bl[129] br[129] wl[162] vdd gnd cell_6t
Xbit_r163_c129 bl[129] br[129] wl[163] vdd gnd cell_6t
Xbit_r164_c129 bl[129] br[129] wl[164] vdd gnd cell_6t
Xbit_r165_c129 bl[129] br[129] wl[165] vdd gnd cell_6t
Xbit_r166_c129 bl[129] br[129] wl[166] vdd gnd cell_6t
Xbit_r167_c129 bl[129] br[129] wl[167] vdd gnd cell_6t
Xbit_r168_c129 bl[129] br[129] wl[168] vdd gnd cell_6t
Xbit_r169_c129 bl[129] br[129] wl[169] vdd gnd cell_6t
Xbit_r170_c129 bl[129] br[129] wl[170] vdd gnd cell_6t
Xbit_r171_c129 bl[129] br[129] wl[171] vdd gnd cell_6t
Xbit_r172_c129 bl[129] br[129] wl[172] vdd gnd cell_6t
Xbit_r173_c129 bl[129] br[129] wl[173] vdd gnd cell_6t
Xbit_r174_c129 bl[129] br[129] wl[174] vdd gnd cell_6t
Xbit_r175_c129 bl[129] br[129] wl[175] vdd gnd cell_6t
Xbit_r176_c129 bl[129] br[129] wl[176] vdd gnd cell_6t
Xbit_r177_c129 bl[129] br[129] wl[177] vdd gnd cell_6t
Xbit_r178_c129 bl[129] br[129] wl[178] vdd gnd cell_6t
Xbit_r179_c129 bl[129] br[129] wl[179] vdd gnd cell_6t
Xbit_r180_c129 bl[129] br[129] wl[180] vdd gnd cell_6t
Xbit_r181_c129 bl[129] br[129] wl[181] vdd gnd cell_6t
Xbit_r182_c129 bl[129] br[129] wl[182] vdd gnd cell_6t
Xbit_r183_c129 bl[129] br[129] wl[183] vdd gnd cell_6t
Xbit_r184_c129 bl[129] br[129] wl[184] vdd gnd cell_6t
Xbit_r185_c129 bl[129] br[129] wl[185] vdd gnd cell_6t
Xbit_r186_c129 bl[129] br[129] wl[186] vdd gnd cell_6t
Xbit_r187_c129 bl[129] br[129] wl[187] vdd gnd cell_6t
Xbit_r188_c129 bl[129] br[129] wl[188] vdd gnd cell_6t
Xbit_r189_c129 bl[129] br[129] wl[189] vdd gnd cell_6t
Xbit_r190_c129 bl[129] br[129] wl[190] vdd gnd cell_6t
Xbit_r191_c129 bl[129] br[129] wl[191] vdd gnd cell_6t
Xbit_r192_c129 bl[129] br[129] wl[192] vdd gnd cell_6t
Xbit_r193_c129 bl[129] br[129] wl[193] vdd gnd cell_6t
Xbit_r194_c129 bl[129] br[129] wl[194] vdd gnd cell_6t
Xbit_r195_c129 bl[129] br[129] wl[195] vdd gnd cell_6t
Xbit_r196_c129 bl[129] br[129] wl[196] vdd gnd cell_6t
Xbit_r197_c129 bl[129] br[129] wl[197] vdd gnd cell_6t
Xbit_r198_c129 bl[129] br[129] wl[198] vdd gnd cell_6t
Xbit_r199_c129 bl[129] br[129] wl[199] vdd gnd cell_6t
Xbit_r200_c129 bl[129] br[129] wl[200] vdd gnd cell_6t
Xbit_r201_c129 bl[129] br[129] wl[201] vdd gnd cell_6t
Xbit_r202_c129 bl[129] br[129] wl[202] vdd gnd cell_6t
Xbit_r203_c129 bl[129] br[129] wl[203] vdd gnd cell_6t
Xbit_r204_c129 bl[129] br[129] wl[204] vdd gnd cell_6t
Xbit_r205_c129 bl[129] br[129] wl[205] vdd gnd cell_6t
Xbit_r206_c129 bl[129] br[129] wl[206] vdd gnd cell_6t
Xbit_r207_c129 bl[129] br[129] wl[207] vdd gnd cell_6t
Xbit_r208_c129 bl[129] br[129] wl[208] vdd gnd cell_6t
Xbit_r209_c129 bl[129] br[129] wl[209] vdd gnd cell_6t
Xbit_r210_c129 bl[129] br[129] wl[210] vdd gnd cell_6t
Xbit_r211_c129 bl[129] br[129] wl[211] vdd gnd cell_6t
Xbit_r212_c129 bl[129] br[129] wl[212] vdd gnd cell_6t
Xbit_r213_c129 bl[129] br[129] wl[213] vdd gnd cell_6t
Xbit_r214_c129 bl[129] br[129] wl[214] vdd gnd cell_6t
Xbit_r215_c129 bl[129] br[129] wl[215] vdd gnd cell_6t
Xbit_r216_c129 bl[129] br[129] wl[216] vdd gnd cell_6t
Xbit_r217_c129 bl[129] br[129] wl[217] vdd gnd cell_6t
Xbit_r218_c129 bl[129] br[129] wl[218] vdd gnd cell_6t
Xbit_r219_c129 bl[129] br[129] wl[219] vdd gnd cell_6t
Xbit_r220_c129 bl[129] br[129] wl[220] vdd gnd cell_6t
Xbit_r221_c129 bl[129] br[129] wl[221] vdd gnd cell_6t
Xbit_r222_c129 bl[129] br[129] wl[222] vdd gnd cell_6t
Xbit_r223_c129 bl[129] br[129] wl[223] vdd gnd cell_6t
Xbit_r224_c129 bl[129] br[129] wl[224] vdd gnd cell_6t
Xbit_r225_c129 bl[129] br[129] wl[225] vdd gnd cell_6t
Xbit_r226_c129 bl[129] br[129] wl[226] vdd gnd cell_6t
Xbit_r227_c129 bl[129] br[129] wl[227] vdd gnd cell_6t
Xbit_r228_c129 bl[129] br[129] wl[228] vdd gnd cell_6t
Xbit_r229_c129 bl[129] br[129] wl[229] vdd gnd cell_6t
Xbit_r230_c129 bl[129] br[129] wl[230] vdd gnd cell_6t
Xbit_r231_c129 bl[129] br[129] wl[231] vdd gnd cell_6t
Xbit_r232_c129 bl[129] br[129] wl[232] vdd gnd cell_6t
Xbit_r233_c129 bl[129] br[129] wl[233] vdd gnd cell_6t
Xbit_r234_c129 bl[129] br[129] wl[234] vdd gnd cell_6t
Xbit_r235_c129 bl[129] br[129] wl[235] vdd gnd cell_6t
Xbit_r236_c129 bl[129] br[129] wl[236] vdd gnd cell_6t
Xbit_r237_c129 bl[129] br[129] wl[237] vdd gnd cell_6t
Xbit_r238_c129 bl[129] br[129] wl[238] vdd gnd cell_6t
Xbit_r239_c129 bl[129] br[129] wl[239] vdd gnd cell_6t
Xbit_r240_c129 bl[129] br[129] wl[240] vdd gnd cell_6t
Xbit_r241_c129 bl[129] br[129] wl[241] vdd gnd cell_6t
Xbit_r242_c129 bl[129] br[129] wl[242] vdd gnd cell_6t
Xbit_r243_c129 bl[129] br[129] wl[243] vdd gnd cell_6t
Xbit_r244_c129 bl[129] br[129] wl[244] vdd gnd cell_6t
Xbit_r245_c129 bl[129] br[129] wl[245] vdd gnd cell_6t
Xbit_r246_c129 bl[129] br[129] wl[246] vdd gnd cell_6t
Xbit_r247_c129 bl[129] br[129] wl[247] vdd gnd cell_6t
Xbit_r248_c129 bl[129] br[129] wl[248] vdd gnd cell_6t
Xbit_r249_c129 bl[129] br[129] wl[249] vdd gnd cell_6t
Xbit_r250_c129 bl[129] br[129] wl[250] vdd gnd cell_6t
Xbit_r251_c129 bl[129] br[129] wl[251] vdd gnd cell_6t
Xbit_r252_c129 bl[129] br[129] wl[252] vdd gnd cell_6t
Xbit_r253_c129 bl[129] br[129] wl[253] vdd gnd cell_6t
Xbit_r254_c129 bl[129] br[129] wl[254] vdd gnd cell_6t
Xbit_r255_c129 bl[129] br[129] wl[255] vdd gnd cell_6t
Xbit_r0_c130 bl[130] br[130] wl[0] vdd gnd cell_6t
Xbit_r1_c130 bl[130] br[130] wl[1] vdd gnd cell_6t
Xbit_r2_c130 bl[130] br[130] wl[2] vdd gnd cell_6t
Xbit_r3_c130 bl[130] br[130] wl[3] vdd gnd cell_6t
Xbit_r4_c130 bl[130] br[130] wl[4] vdd gnd cell_6t
Xbit_r5_c130 bl[130] br[130] wl[5] vdd gnd cell_6t
Xbit_r6_c130 bl[130] br[130] wl[6] vdd gnd cell_6t
Xbit_r7_c130 bl[130] br[130] wl[7] vdd gnd cell_6t
Xbit_r8_c130 bl[130] br[130] wl[8] vdd gnd cell_6t
Xbit_r9_c130 bl[130] br[130] wl[9] vdd gnd cell_6t
Xbit_r10_c130 bl[130] br[130] wl[10] vdd gnd cell_6t
Xbit_r11_c130 bl[130] br[130] wl[11] vdd gnd cell_6t
Xbit_r12_c130 bl[130] br[130] wl[12] vdd gnd cell_6t
Xbit_r13_c130 bl[130] br[130] wl[13] vdd gnd cell_6t
Xbit_r14_c130 bl[130] br[130] wl[14] vdd gnd cell_6t
Xbit_r15_c130 bl[130] br[130] wl[15] vdd gnd cell_6t
Xbit_r16_c130 bl[130] br[130] wl[16] vdd gnd cell_6t
Xbit_r17_c130 bl[130] br[130] wl[17] vdd gnd cell_6t
Xbit_r18_c130 bl[130] br[130] wl[18] vdd gnd cell_6t
Xbit_r19_c130 bl[130] br[130] wl[19] vdd gnd cell_6t
Xbit_r20_c130 bl[130] br[130] wl[20] vdd gnd cell_6t
Xbit_r21_c130 bl[130] br[130] wl[21] vdd gnd cell_6t
Xbit_r22_c130 bl[130] br[130] wl[22] vdd gnd cell_6t
Xbit_r23_c130 bl[130] br[130] wl[23] vdd gnd cell_6t
Xbit_r24_c130 bl[130] br[130] wl[24] vdd gnd cell_6t
Xbit_r25_c130 bl[130] br[130] wl[25] vdd gnd cell_6t
Xbit_r26_c130 bl[130] br[130] wl[26] vdd gnd cell_6t
Xbit_r27_c130 bl[130] br[130] wl[27] vdd gnd cell_6t
Xbit_r28_c130 bl[130] br[130] wl[28] vdd gnd cell_6t
Xbit_r29_c130 bl[130] br[130] wl[29] vdd gnd cell_6t
Xbit_r30_c130 bl[130] br[130] wl[30] vdd gnd cell_6t
Xbit_r31_c130 bl[130] br[130] wl[31] vdd gnd cell_6t
Xbit_r32_c130 bl[130] br[130] wl[32] vdd gnd cell_6t
Xbit_r33_c130 bl[130] br[130] wl[33] vdd gnd cell_6t
Xbit_r34_c130 bl[130] br[130] wl[34] vdd gnd cell_6t
Xbit_r35_c130 bl[130] br[130] wl[35] vdd gnd cell_6t
Xbit_r36_c130 bl[130] br[130] wl[36] vdd gnd cell_6t
Xbit_r37_c130 bl[130] br[130] wl[37] vdd gnd cell_6t
Xbit_r38_c130 bl[130] br[130] wl[38] vdd gnd cell_6t
Xbit_r39_c130 bl[130] br[130] wl[39] vdd gnd cell_6t
Xbit_r40_c130 bl[130] br[130] wl[40] vdd gnd cell_6t
Xbit_r41_c130 bl[130] br[130] wl[41] vdd gnd cell_6t
Xbit_r42_c130 bl[130] br[130] wl[42] vdd gnd cell_6t
Xbit_r43_c130 bl[130] br[130] wl[43] vdd gnd cell_6t
Xbit_r44_c130 bl[130] br[130] wl[44] vdd gnd cell_6t
Xbit_r45_c130 bl[130] br[130] wl[45] vdd gnd cell_6t
Xbit_r46_c130 bl[130] br[130] wl[46] vdd gnd cell_6t
Xbit_r47_c130 bl[130] br[130] wl[47] vdd gnd cell_6t
Xbit_r48_c130 bl[130] br[130] wl[48] vdd gnd cell_6t
Xbit_r49_c130 bl[130] br[130] wl[49] vdd gnd cell_6t
Xbit_r50_c130 bl[130] br[130] wl[50] vdd gnd cell_6t
Xbit_r51_c130 bl[130] br[130] wl[51] vdd gnd cell_6t
Xbit_r52_c130 bl[130] br[130] wl[52] vdd gnd cell_6t
Xbit_r53_c130 bl[130] br[130] wl[53] vdd gnd cell_6t
Xbit_r54_c130 bl[130] br[130] wl[54] vdd gnd cell_6t
Xbit_r55_c130 bl[130] br[130] wl[55] vdd gnd cell_6t
Xbit_r56_c130 bl[130] br[130] wl[56] vdd gnd cell_6t
Xbit_r57_c130 bl[130] br[130] wl[57] vdd gnd cell_6t
Xbit_r58_c130 bl[130] br[130] wl[58] vdd gnd cell_6t
Xbit_r59_c130 bl[130] br[130] wl[59] vdd gnd cell_6t
Xbit_r60_c130 bl[130] br[130] wl[60] vdd gnd cell_6t
Xbit_r61_c130 bl[130] br[130] wl[61] vdd gnd cell_6t
Xbit_r62_c130 bl[130] br[130] wl[62] vdd gnd cell_6t
Xbit_r63_c130 bl[130] br[130] wl[63] vdd gnd cell_6t
Xbit_r64_c130 bl[130] br[130] wl[64] vdd gnd cell_6t
Xbit_r65_c130 bl[130] br[130] wl[65] vdd gnd cell_6t
Xbit_r66_c130 bl[130] br[130] wl[66] vdd gnd cell_6t
Xbit_r67_c130 bl[130] br[130] wl[67] vdd gnd cell_6t
Xbit_r68_c130 bl[130] br[130] wl[68] vdd gnd cell_6t
Xbit_r69_c130 bl[130] br[130] wl[69] vdd gnd cell_6t
Xbit_r70_c130 bl[130] br[130] wl[70] vdd gnd cell_6t
Xbit_r71_c130 bl[130] br[130] wl[71] vdd gnd cell_6t
Xbit_r72_c130 bl[130] br[130] wl[72] vdd gnd cell_6t
Xbit_r73_c130 bl[130] br[130] wl[73] vdd gnd cell_6t
Xbit_r74_c130 bl[130] br[130] wl[74] vdd gnd cell_6t
Xbit_r75_c130 bl[130] br[130] wl[75] vdd gnd cell_6t
Xbit_r76_c130 bl[130] br[130] wl[76] vdd gnd cell_6t
Xbit_r77_c130 bl[130] br[130] wl[77] vdd gnd cell_6t
Xbit_r78_c130 bl[130] br[130] wl[78] vdd gnd cell_6t
Xbit_r79_c130 bl[130] br[130] wl[79] vdd gnd cell_6t
Xbit_r80_c130 bl[130] br[130] wl[80] vdd gnd cell_6t
Xbit_r81_c130 bl[130] br[130] wl[81] vdd gnd cell_6t
Xbit_r82_c130 bl[130] br[130] wl[82] vdd gnd cell_6t
Xbit_r83_c130 bl[130] br[130] wl[83] vdd gnd cell_6t
Xbit_r84_c130 bl[130] br[130] wl[84] vdd gnd cell_6t
Xbit_r85_c130 bl[130] br[130] wl[85] vdd gnd cell_6t
Xbit_r86_c130 bl[130] br[130] wl[86] vdd gnd cell_6t
Xbit_r87_c130 bl[130] br[130] wl[87] vdd gnd cell_6t
Xbit_r88_c130 bl[130] br[130] wl[88] vdd gnd cell_6t
Xbit_r89_c130 bl[130] br[130] wl[89] vdd gnd cell_6t
Xbit_r90_c130 bl[130] br[130] wl[90] vdd gnd cell_6t
Xbit_r91_c130 bl[130] br[130] wl[91] vdd gnd cell_6t
Xbit_r92_c130 bl[130] br[130] wl[92] vdd gnd cell_6t
Xbit_r93_c130 bl[130] br[130] wl[93] vdd gnd cell_6t
Xbit_r94_c130 bl[130] br[130] wl[94] vdd gnd cell_6t
Xbit_r95_c130 bl[130] br[130] wl[95] vdd gnd cell_6t
Xbit_r96_c130 bl[130] br[130] wl[96] vdd gnd cell_6t
Xbit_r97_c130 bl[130] br[130] wl[97] vdd gnd cell_6t
Xbit_r98_c130 bl[130] br[130] wl[98] vdd gnd cell_6t
Xbit_r99_c130 bl[130] br[130] wl[99] vdd gnd cell_6t
Xbit_r100_c130 bl[130] br[130] wl[100] vdd gnd cell_6t
Xbit_r101_c130 bl[130] br[130] wl[101] vdd gnd cell_6t
Xbit_r102_c130 bl[130] br[130] wl[102] vdd gnd cell_6t
Xbit_r103_c130 bl[130] br[130] wl[103] vdd gnd cell_6t
Xbit_r104_c130 bl[130] br[130] wl[104] vdd gnd cell_6t
Xbit_r105_c130 bl[130] br[130] wl[105] vdd gnd cell_6t
Xbit_r106_c130 bl[130] br[130] wl[106] vdd gnd cell_6t
Xbit_r107_c130 bl[130] br[130] wl[107] vdd gnd cell_6t
Xbit_r108_c130 bl[130] br[130] wl[108] vdd gnd cell_6t
Xbit_r109_c130 bl[130] br[130] wl[109] vdd gnd cell_6t
Xbit_r110_c130 bl[130] br[130] wl[110] vdd gnd cell_6t
Xbit_r111_c130 bl[130] br[130] wl[111] vdd gnd cell_6t
Xbit_r112_c130 bl[130] br[130] wl[112] vdd gnd cell_6t
Xbit_r113_c130 bl[130] br[130] wl[113] vdd gnd cell_6t
Xbit_r114_c130 bl[130] br[130] wl[114] vdd gnd cell_6t
Xbit_r115_c130 bl[130] br[130] wl[115] vdd gnd cell_6t
Xbit_r116_c130 bl[130] br[130] wl[116] vdd gnd cell_6t
Xbit_r117_c130 bl[130] br[130] wl[117] vdd gnd cell_6t
Xbit_r118_c130 bl[130] br[130] wl[118] vdd gnd cell_6t
Xbit_r119_c130 bl[130] br[130] wl[119] vdd gnd cell_6t
Xbit_r120_c130 bl[130] br[130] wl[120] vdd gnd cell_6t
Xbit_r121_c130 bl[130] br[130] wl[121] vdd gnd cell_6t
Xbit_r122_c130 bl[130] br[130] wl[122] vdd gnd cell_6t
Xbit_r123_c130 bl[130] br[130] wl[123] vdd gnd cell_6t
Xbit_r124_c130 bl[130] br[130] wl[124] vdd gnd cell_6t
Xbit_r125_c130 bl[130] br[130] wl[125] vdd gnd cell_6t
Xbit_r126_c130 bl[130] br[130] wl[126] vdd gnd cell_6t
Xbit_r127_c130 bl[130] br[130] wl[127] vdd gnd cell_6t
Xbit_r128_c130 bl[130] br[130] wl[128] vdd gnd cell_6t
Xbit_r129_c130 bl[130] br[130] wl[129] vdd gnd cell_6t
Xbit_r130_c130 bl[130] br[130] wl[130] vdd gnd cell_6t
Xbit_r131_c130 bl[130] br[130] wl[131] vdd gnd cell_6t
Xbit_r132_c130 bl[130] br[130] wl[132] vdd gnd cell_6t
Xbit_r133_c130 bl[130] br[130] wl[133] vdd gnd cell_6t
Xbit_r134_c130 bl[130] br[130] wl[134] vdd gnd cell_6t
Xbit_r135_c130 bl[130] br[130] wl[135] vdd gnd cell_6t
Xbit_r136_c130 bl[130] br[130] wl[136] vdd gnd cell_6t
Xbit_r137_c130 bl[130] br[130] wl[137] vdd gnd cell_6t
Xbit_r138_c130 bl[130] br[130] wl[138] vdd gnd cell_6t
Xbit_r139_c130 bl[130] br[130] wl[139] vdd gnd cell_6t
Xbit_r140_c130 bl[130] br[130] wl[140] vdd gnd cell_6t
Xbit_r141_c130 bl[130] br[130] wl[141] vdd gnd cell_6t
Xbit_r142_c130 bl[130] br[130] wl[142] vdd gnd cell_6t
Xbit_r143_c130 bl[130] br[130] wl[143] vdd gnd cell_6t
Xbit_r144_c130 bl[130] br[130] wl[144] vdd gnd cell_6t
Xbit_r145_c130 bl[130] br[130] wl[145] vdd gnd cell_6t
Xbit_r146_c130 bl[130] br[130] wl[146] vdd gnd cell_6t
Xbit_r147_c130 bl[130] br[130] wl[147] vdd gnd cell_6t
Xbit_r148_c130 bl[130] br[130] wl[148] vdd gnd cell_6t
Xbit_r149_c130 bl[130] br[130] wl[149] vdd gnd cell_6t
Xbit_r150_c130 bl[130] br[130] wl[150] vdd gnd cell_6t
Xbit_r151_c130 bl[130] br[130] wl[151] vdd gnd cell_6t
Xbit_r152_c130 bl[130] br[130] wl[152] vdd gnd cell_6t
Xbit_r153_c130 bl[130] br[130] wl[153] vdd gnd cell_6t
Xbit_r154_c130 bl[130] br[130] wl[154] vdd gnd cell_6t
Xbit_r155_c130 bl[130] br[130] wl[155] vdd gnd cell_6t
Xbit_r156_c130 bl[130] br[130] wl[156] vdd gnd cell_6t
Xbit_r157_c130 bl[130] br[130] wl[157] vdd gnd cell_6t
Xbit_r158_c130 bl[130] br[130] wl[158] vdd gnd cell_6t
Xbit_r159_c130 bl[130] br[130] wl[159] vdd gnd cell_6t
Xbit_r160_c130 bl[130] br[130] wl[160] vdd gnd cell_6t
Xbit_r161_c130 bl[130] br[130] wl[161] vdd gnd cell_6t
Xbit_r162_c130 bl[130] br[130] wl[162] vdd gnd cell_6t
Xbit_r163_c130 bl[130] br[130] wl[163] vdd gnd cell_6t
Xbit_r164_c130 bl[130] br[130] wl[164] vdd gnd cell_6t
Xbit_r165_c130 bl[130] br[130] wl[165] vdd gnd cell_6t
Xbit_r166_c130 bl[130] br[130] wl[166] vdd gnd cell_6t
Xbit_r167_c130 bl[130] br[130] wl[167] vdd gnd cell_6t
Xbit_r168_c130 bl[130] br[130] wl[168] vdd gnd cell_6t
Xbit_r169_c130 bl[130] br[130] wl[169] vdd gnd cell_6t
Xbit_r170_c130 bl[130] br[130] wl[170] vdd gnd cell_6t
Xbit_r171_c130 bl[130] br[130] wl[171] vdd gnd cell_6t
Xbit_r172_c130 bl[130] br[130] wl[172] vdd gnd cell_6t
Xbit_r173_c130 bl[130] br[130] wl[173] vdd gnd cell_6t
Xbit_r174_c130 bl[130] br[130] wl[174] vdd gnd cell_6t
Xbit_r175_c130 bl[130] br[130] wl[175] vdd gnd cell_6t
Xbit_r176_c130 bl[130] br[130] wl[176] vdd gnd cell_6t
Xbit_r177_c130 bl[130] br[130] wl[177] vdd gnd cell_6t
Xbit_r178_c130 bl[130] br[130] wl[178] vdd gnd cell_6t
Xbit_r179_c130 bl[130] br[130] wl[179] vdd gnd cell_6t
Xbit_r180_c130 bl[130] br[130] wl[180] vdd gnd cell_6t
Xbit_r181_c130 bl[130] br[130] wl[181] vdd gnd cell_6t
Xbit_r182_c130 bl[130] br[130] wl[182] vdd gnd cell_6t
Xbit_r183_c130 bl[130] br[130] wl[183] vdd gnd cell_6t
Xbit_r184_c130 bl[130] br[130] wl[184] vdd gnd cell_6t
Xbit_r185_c130 bl[130] br[130] wl[185] vdd gnd cell_6t
Xbit_r186_c130 bl[130] br[130] wl[186] vdd gnd cell_6t
Xbit_r187_c130 bl[130] br[130] wl[187] vdd gnd cell_6t
Xbit_r188_c130 bl[130] br[130] wl[188] vdd gnd cell_6t
Xbit_r189_c130 bl[130] br[130] wl[189] vdd gnd cell_6t
Xbit_r190_c130 bl[130] br[130] wl[190] vdd gnd cell_6t
Xbit_r191_c130 bl[130] br[130] wl[191] vdd gnd cell_6t
Xbit_r192_c130 bl[130] br[130] wl[192] vdd gnd cell_6t
Xbit_r193_c130 bl[130] br[130] wl[193] vdd gnd cell_6t
Xbit_r194_c130 bl[130] br[130] wl[194] vdd gnd cell_6t
Xbit_r195_c130 bl[130] br[130] wl[195] vdd gnd cell_6t
Xbit_r196_c130 bl[130] br[130] wl[196] vdd gnd cell_6t
Xbit_r197_c130 bl[130] br[130] wl[197] vdd gnd cell_6t
Xbit_r198_c130 bl[130] br[130] wl[198] vdd gnd cell_6t
Xbit_r199_c130 bl[130] br[130] wl[199] vdd gnd cell_6t
Xbit_r200_c130 bl[130] br[130] wl[200] vdd gnd cell_6t
Xbit_r201_c130 bl[130] br[130] wl[201] vdd gnd cell_6t
Xbit_r202_c130 bl[130] br[130] wl[202] vdd gnd cell_6t
Xbit_r203_c130 bl[130] br[130] wl[203] vdd gnd cell_6t
Xbit_r204_c130 bl[130] br[130] wl[204] vdd gnd cell_6t
Xbit_r205_c130 bl[130] br[130] wl[205] vdd gnd cell_6t
Xbit_r206_c130 bl[130] br[130] wl[206] vdd gnd cell_6t
Xbit_r207_c130 bl[130] br[130] wl[207] vdd gnd cell_6t
Xbit_r208_c130 bl[130] br[130] wl[208] vdd gnd cell_6t
Xbit_r209_c130 bl[130] br[130] wl[209] vdd gnd cell_6t
Xbit_r210_c130 bl[130] br[130] wl[210] vdd gnd cell_6t
Xbit_r211_c130 bl[130] br[130] wl[211] vdd gnd cell_6t
Xbit_r212_c130 bl[130] br[130] wl[212] vdd gnd cell_6t
Xbit_r213_c130 bl[130] br[130] wl[213] vdd gnd cell_6t
Xbit_r214_c130 bl[130] br[130] wl[214] vdd gnd cell_6t
Xbit_r215_c130 bl[130] br[130] wl[215] vdd gnd cell_6t
Xbit_r216_c130 bl[130] br[130] wl[216] vdd gnd cell_6t
Xbit_r217_c130 bl[130] br[130] wl[217] vdd gnd cell_6t
Xbit_r218_c130 bl[130] br[130] wl[218] vdd gnd cell_6t
Xbit_r219_c130 bl[130] br[130] wl[219] vdd gnd cell_6t
Xbit_r220_c130 bl[130] br[130] wl[220] vdd gnd cell_6t
Xbit_r221_c130 bl[130] br[130] wl[221] vdd gnd cell_6t
Xbit_r222_c130 bl[130] br[130] wl[222] vdd gnd cell_6t
Xbit_r223_c130 bl[130] br[130] wl[223] vdd gnd cell_6t
Xbit_r224_c130 bl[130] br[130] wl[224] vdd gnd cell_6t
Xbit_r225_c130 bl[130] br[130] wl[225] vdd gnd cell_6t
Xbit_r226_c130 bl[130] br[130] wl[226] vdd gnd cell_6t
Xbit_r227_c130 bl[130] br[130] wl[227] vdd gnd cell_6t
Xbit_r228_c130 bl[130] br[130] wl[228] vdd gnd cell_6t
Xbit_r229_c130 bl[130] br[130] wl[229] vdd gnd cell_6t
Xbit_r230_c130 bl[130] br[130] wl[230] vdd gnd cell_6t
Xbit_r231_c130 bl[130] br[130] wl[231] vdd gnd cell_6t
Xbit_r232_c130 bl[130] br[130] wl[232] vdd gnd cell_6t
Xbit_r233_c130 bl[130] br[130] wl[233] vdd gnd cell_6t
Xbit_r234_c130 bl[130] br[130] wl[234] vdd gnd cell_6t
Xbit_r235_c130 bl[130] br[130] wl[235] vdd gnd cell_6t
Xbit_r236_c130 bl[130] br[130] wl[236] vdd gnd cell_6t
Xbit_r237_c130 bl[130] br[130] wl[237] vdd gnd cell_6t
Xbit_r238_c130 bl[130] br[130] wl[238] vdd gnd cell_6t
Xbit_r239_c130 bl[130] br[130] wl[239] vdd gnd cell_6t
Xbit_r240_c130 bl[130] br[130] wl[240] vdd gnd cell_6t
Xbit_r241_c130 bl[130] br[130] wl[241] vdd gnd cell_6t
Xbit_r242_c130 bl[130] br[130] wl[242] vdd gnd cell_6t
Xbit_r243_c130 bl[130] br[130] wl[243] vdd gnd cell_6t
Xbit_r244_c130 bl[130] br[130] wl[244] vdd gnd cell_6t
Xbit_r245_c130 bl[130] br[130] wl[245] vdd gnd cell_6t
Xbit_r246_c130 bl[130] br[130] wl[246] vdd gnd cell_6t
Xbit_r247_c130 bl[130] br[130] wl[247] vdd gnd cell_6t
Xbit_r248_c130 bl[130] br[130] wl[248] vdd gnd cell_6t
Xbit_r249_c130 bl[130] br[130] wl[249] vdd gnd cell_6t
Xbit_r250_c130 bl[130] br[130] wl[250] vdd gnd cell_6t
Xbit_r251_c130 bl[130] br[130] wl[251] vdd gnd cell_6t
Xbit_r252_c130 bl[130] br[130] wl[252] vdd gnd cell_6t
Xbit_r253_c130 bl[130] br[130] wl[253] vdd gnd cell_6t
Xbit_r254_c130 bl[130] br[130] wl[254] vdd gnd cell_6t
Xbit_r255_c130 bl[130] br[130] wl[255] vdd gnd cell_6t
Xbit_r0_c131 bl[131] br[131] wl[0] vdd gnd cell_6t
Xbit_r1_c131 bl[131] br[131] wl[1] vdd gnd cell_6t
Xbit_r2_c131 bl[131] br[131] wl[2] vdd gnd cell_6t
Xbit_r3_c131 bl[131] br[131] wl[3] vdd gnd cell_6t
Xbit_r4_c131 bl[131] br[131] wl[4] vdd gnd cell_6t
Xbit_r5_c131 bl[131] br[131] wl[5] vdd gnd cell_6t
Xbit_r6_c131 bl[131] br[131] wl[6] vdd gnd cell_6t
Xbit_r7_c131 bl[131] br[131] wl[7] vdd gnd cell_6t
Xbit_r8_c131 bl[131] br[131] wl[8] vdd gnd cell_6t
Xbit_r9_c131 bl[131] br[131] wl[9] vdd gnd cell_6t
Xbit_r10_c131 bl[131] br[131] wl[10] vdd gnd cell_6t
Xbit_r11_c131 bl[131] br[131] wl[11] vdd gnd cell_6t
Xbit_r12_c131 bl[131] br[131] wl[12] vdd gnd cell_6t
Xbit_r13_c131 bl[131] br[131] wl[13] vdd gnd cell_6t
Xbit_r14_c131 bl[131] br[131] wl[14] vdd gnd cell_6t
Xbit_r15_c131 bl[131] br[131] wl[15] vdd gnd cell_6t
Xbit_r16_c131 bl[131] br[131] wl[16] vdd gnd cell_6t
Xbit_r17_c131 bl[131] br[131] wl[17] vdd gnd cell_6t
Xbit_r18_c131 bl[131] br[131] wl[18] vdd gnd cell_6t
Xbit_r19_c131 bl[131] br[131] wl[19] vdd gnd cell_6t
Xbit_r20_c131 bl[131] br[131] wl[20] vdd gnd cell_6t
Xbit_r21_c131 bl[131] br[131] wl[21] vdd gnd cell_6t
Xbit_r22_c131 bl[131] br[131] wl[22] vdd gnd cell_6t
Xbit_r23_c131 bl[131] br[131] wl[23] vdd gnd cell_6t
Xbit_r24_c131 bl[131] br[131] wl[24] vdd gnd cell_6t
Xbit_r25_c131 bl[131] br[131] wl[25] vdd gnd cell_6t
Xbit_r26_c131 bl[131] br[131] wl[26] vdd gnd cell_6t
Xbit_r27_c131 bl[131] br[131] wl[27] vdd gnd cell_6t
Xbit_r28_c131 bl[131] br[131] wl[28] vdd gnd cell_6t
Xbit_r29_c131 bl[131] br[131] wl[29] vdd gnd cell_6t
Xbit_r30_c131 bl[131] br[131] wl[30] vdd gnd cell_6t
Xbit_r31_c131 bl[131] br[131] wl[31] vdd gnd cell_6t
Xbit_r32_c131 bl[131] br[131] wl[32] vdd gnd cell_6t
Xbit_r33_c131 bl[131] br[131] wl[33] vdd gnd cell_6t
Xbit_r34_c131 bl[131] br[131] wl[34] vdd gnd cell_6t
Xbit_r35_c131 bl[131] br[131] wl[35] vdd gnd cell_6t
Xbit_r36_c131 bl[131] br[131] wl[36] vdd gnd cell_6t
Xbit_r37_c131 bl[131] br[131] wl[37] vdd gnd cell_6t
Xbit_r38_c131 bl[131] br[131] wl[38] vdd gnd cell_6t
Xbit_r39_c131 bl[131] br[131] wl[39] vdd gnd cell_6t
Xbit_r40_c131 bl[131] br[131] wl[40] vdd gnd cell_6t
Xbit_r41_c131 bl[131] br[131] wl[41] vdd gnd cell_6t
Xbit_r42_c131 bl[131] br[131] wl[42] vdd gnd cell_6t
Xbit_r43_c131 bl[131] br[131] wl[43] vdd gnd cell_6t
Xbit_r44_c131 bl[131] br[131] wl[44] vdd gnd cell_6t
Xbit_r45_c131 bl[131] br[131] wl[45] vdd gnd cell_6t
Xbit_r46_c131 bl[131] br[131] wl[46] vdd gnd cell_6t
Xbit_r47_c131 bl[131] br[131] wl[47] vdd gnd cell_6t
Xbit_r48_c131 bl[131] br[131] wl[48] vdd gnd cell_6t
Xbit_r49_c131 bl[131] br[131] wl[49] vdd gnd cell_6t
Xbit_r50_c131 bl[131] br[131] wl[50] vdd gnd cell_6t
Xbit_r51_c131 bl[131] br[131] wl[51] vdd gnd cell_6t
Xbit_r52_c131 bl[131] br[131] wl[52] vdd gnd cell_6t
Xbit_r53_c131 bl[131] br[131] wl[53] vdd gnd cell_6t
Xbit_r54_c131 bl[131] br[131] wl[54] vdd gnd cell_6t
Xbit_r55_c131 bl[131] br[131] wl[55] vdd gnd cell_6t
Xbit_r56_c131 bl[131] br[131] wl[56] vdd gnd cell_6t
Xbit_r57_c131 bl[131] br[131] wl[57] vdd gnd cell_6t
Xbit_r58_c131 bl[131] br[131] wl[58] vdd gnd cell_6t
Xbit_r59_c131 bl[131] br[131] wl[59] vdd gnd cell_6t
Xbit_r60_c131 bl[131] br[131] wl[60] vdd gnd cell_6t
Xbit_r61_c131 bl[131] br[131] wl[61] vdd gnd cell_6t
Xbit_r62_c131 bl[131] br[131] wl[62] vdd gnd cell_6t
Xbit_r63_c131 bl[131] br[131] wl[63] vdd gnd cell_6t
Xbit_r64_c131 bl[131] br[131] wl[64] vdd gnd cell_6t
Xbit_r65_c131 bl[131] br[131] wl[65] vdd gnd cell_6t
Xbit_r66_c131 bl[131] br[131] wl[66] vdd gnd cell_6t
Xbit_r67_c131 bl[131] br[131] wl[67] vdd gnd cell_6t
Xbit_r68_c131 bl[131] br[131] wl[68] vdd gnd cell_6t
Xbit_r69_c131 bl[131] br[131] wl[69] vdd gnd cell_6t
Xbit_r70_c131 bl[131] br[131] wl[70] vdd gnd cell_6t
Xbit_r71_c131 bl[131] br[131] wl[71] vdd gnd cell_6t
Xbit_r72_c131 bl[131] br[131] wl[72] vdd gnd cell_6t
Xbit_r73_c131 bl[131] br[131] wl[73] vdd gnd cell_6t
Xbit_r74_c131 bl[131] br[131] wl[74] vdd gnd cell_6t
Xbit_r75_c131 bl[131] br[131] wl[75] vdd gnd cell_6t
Xbit_r76_c131 bl[131] br[131] wl[76] vdd gnd cell_6t
Xbit_r77_c131 bl[131] br[131] wl[77] vdd gnd cell_6t
Xbit_r78_c131 bl[131] br[131] wl[78] vdd gnd cell_6t
Xbit_r79_c131 bl[131] br[131] wl[79] vdd gnd cell_6t
Xbit_r80_c131 bl[131] br[131] wl[80] vdd gnd cell_6t
Xbit_r81_c131 bl[131] br[131] wl[81] vdd gnd cell_6t
Xbit_r82_c131 bl[131] br[131] wl[82] vdd gnd cell_6t
Xbit_r83_c131 bl[131] br[131] wl[83] vdd gnd cell_6t
Xbit_r84_c131 bl[131] br[131] wl[84] vdd gnd cell_6t
Xbit_r85_c131 bl[131] br[131] wl[85] vdd gnd cell_6t
Xbit_r86_c131 bl[131] br[131] wl[86] vdd gnd cell_6t
Xbit_r87_c131 bl[131] br[131] wl[87] vdd gnd cell_6t
Xbit_r88_c131 bl[131] br[131] wl[88] vdd gnd cell_6t
Xbit_r89_c131 bl[131] br[131] wl[89] vdd gnd cell_6t
Xbit_r90_c131 bl[131] br[131] wl[90] vdd gnd cell_6t
Xbit_r91_c131 bl[131] br[131] wl[91] vdd gnd cell_6t
Xbit_r92_c131 bl[131] br[131] wl[92] vdd gnd cell_6t
Xbit_r93_c131 bl[131] br[131] wl[93] vdd gnd cell_6t
Xbit_r94_c131 bl[131] br[131] wl[94] vdd gnd cell_6t
Xbit_r95_c131 bl[131] br[131] wl[95] vdd gnd cell_6t
Xbit_r96_c131 bl[131] br[131] wl[96] vdd gnd cell_6t
Xbit_r97_c131 bl[131] br[131] wl[97] vdd gnd cell_6t
Xbit_r98_c131 bl[131] br[131] wl[98] vdd gnd cell_6t
Xbit_r99_c131 bl[131] br[131] wl[99] vdd gnd cell_6t
Xbit_r100_c131 bl[131] br[131] wl[100] vdd gnd cell_6t
Xbit_r101_c131 bl[131] br[131] wl[101] vdd gnd cell_6t
Xbit_r102_c131 bl[131] br[131] wl[102] vdd gnd cell_6t
Xbit_r103_c131 bl[131] br[131] wl[103] vdd gnd cell_6t
Xbit_r104_c131 bl[131] br[131] wl[104] vdd gnd cell_6t
Xbit_r105_c131 bl[131] br[131] wl[105] vdd gnd cell_6t
Xbit_r106_c131 bl[131] br[131] wl[106] vdd gnd cell_6t
Xbit_r107_c131 bl[131] br[131] wl[107] vdd gnd cell_6t
Xbit_r108_c131 bl[131] br[131] wl[108] vdd gnd cell_6t
Xbit_r109_c131 bl[131] br[131] wl[109] vdd gnd cell_6t
Xbit_r110_c131 bl[131] br[131] wl[110] vdd gnd cell_6t
Xbit_r111_c131 bl[131] br[131] wl[111] vdd gnd cell_6t
Xbit_r112_c131 bl[131] br[131] wl[112] vdd gnd cell_6t
Xbit_r113_c131 bl[131] br[131] wl[113] vdd gnd cell_6t
Xbit_r114_c131 bl[131] br[131] wl[114] vdd gnd cell_6t
Xbit_r115_c131 bl[131] br[131] wl[115] vdd gnd cell_6t
Xbit_r116_c131 bl[131] br[131] wl[116] vdd gnd cell_6t
Xbit_r117_c131 bl[131] br[131] wl[117] vdd gnd cell_6t
Xbit_r118_c131 bl[131] br[131] wl[118] vdd gnd cell_6t
Xbit_r119_c131 bl[131] br[131] wl[119] vdd gnd cell_6t
Xbit_r120_c131 bl[131] br[131] wl[120] vdd gnd cell_6t
Xbit_r121_c131 bl[131] br[131] wl[121] vdd gnd cell_6t
Xbit_r122_c131 bl[131] br[131] wl[122] vdd gnd cell_6t
Xbit_r123_c131 bl[131] br[131] wl[123] vdd gnd cell_6t
Xbit_r124_c131 bl[131] br[131] wl[124] vdd gnd cell_6t
Xbit_r125_c131 bl[131] br[131] wl[125] vdd gnd cell_6t
Xbit_r126_c131 bl[131] br[131] wl[126] vdd gnd cell_6t
Xbit_r127_c131 bl[131] br[131] wl[127] vdd gnd cell_6t
Xbit_r128_c131 bl[131] br[131] wl[128] vdd gnd cell_6t
Xbit_r129_c131 bl[131] br[131] wl[129] vdd gnd cell_6t
Xbit_r130_c131 bl[131] br[131] wl[130] vdd gnd cell_6t
Xbit_r131_c131 bl[131] br[131] wl[131] vdd gnd cell_6t
Xbit_r132_c131 bl[131] br[131] wl[132] vdd gnd cell_6t
Xbit_r133_c131 bl[131] br[131] wl[133] vdd gnd cell_6t
Xbit_r134_c131 bl[131] br[131] wl[134] vdd gnd cell_6t
Xbit_r135_c131 bl[131] br[131] wl[135] vdd gnd cell_6t
Xbit_r136_c131 bl[131] br[131] wl[136] vdd gnd cell_6t
Xbit_r137_c131 bl[131] br[131] wl[137] vdd gnd cell_6t
Xbit_r138_c131 bl[131] br[131] wl[138] vdd gnd cell_6t
Xbit_r139_c131 bl[131] br[131] wl[139] vdd gnd cell_6t
Xbit_r140_c131 bl[131] br[131] wl[140] vdd gnd cell_6t
Xbit_r141_c131 bl[131] br[131] wl[141] vdd gnd cell_6t
Xbit_r142_c131 bl[131] br[131] wl[142] vdd gnd cell_6t
Xbit_r143_c131 bl[131] br[131] wl[143] vdd gnd cell_6t
Xbit_r144_c131 bl[131] br[131] wl[144] vdd gnd cell_6t
Xbit_r145_c131 bl[131] br[131] wl[145] vdd gnd cell_6t
Xbit_r146_c131 bl[131] br[131] wl[146] vdd gnd cell_6t
Xbit_r147_c131 bl[131] br[131] wl[147] vdd gnd cell_6t
Xbit_r148_c131 bl[131] br[131] wl[148] vdd gnd cell_6t
Xbit_r149_c131 bl[131] br[131] wl[149] vdd gnd cell_6t
Xbit_r150_c131 bl[131] br[131] wl[150] vdd gnd cell_6t
Xbit_r151_c131 bl[131] br[131] wl[151] vdd gnd cell_6t
Xbit_r152_c131 bl[131] br[131] wl[152] vdd gnd cell_6t
Xbit_r153_c131 bl[131] br[131] wl[153] vdd gnd cell_6t
Xbit_r154_c131 bl[131] br[131] wl[154] vdd gnd cell_6t
Xbit_r155_c131 bl[131] br[131] wl[155] vdd gnd cell_6t
Xbit_r156_c131 bl[131] br[131] wl[156] vdd gnd cell_6t
Xbit_r157_c131 bl[131] br[131] wl[157] vdd gnd cell_6t
Xbit_r158_c131 bl[131] br[131] wl[158] vdd gnd cell_6t
Xbit_r159_c131 bl[131] br[131] wl[159] vdd gnd cell_6t
Xbit_r160_c131 bl[131] br[131] wl[160] vdd gnd cell_6t
Xbit_r161_c131 bl[131] br[131] wl[161] vdd gnd cell_6t
Xbit_r162_c131 bl[131] br[131] wl[162] vdd gnd cell_6t
Xbit_r163_c131 bl[131] br[131] wl[163] vdd gnd cell_6t
Xbit_r164_c131 bl[131] br[131] wl[164] vdd gnd cell_6t
Xbit_r165_c131 bl[131] br[131] wl[165] vdd gnd cell_6t
Xbit_r166_c131 bl[131] br[131] wl[166] vdd gnd cell_6t
Xbit_r167_c131 bl[131] br[131] wl[167] vdd gnd cell_6t
Xbit_r168_c131 bl[131] br[131] wl[168] vdd gnd cell_6t
Xbit_r169_c131 bl[131] br[131] wl[169] vdd gnd cell_6t
Xbit_r170_c131 bl[131] br[131] wl[170] vdd gnd cell_6t
Xbit_r171_c131 bl[131] br[131] wl[171] vdd gnd cell_6t
Xbit_r172_c131 bl[131] br[131] wl[172] vdd gnd cell_6t
Xbit_r173_c131 bl[131] br[131] wl[173] vdd gnd cell_6t
Xbit_r174_c131 bl[131] br[131] wl[174] vdd gnd cell_6t
Xbit_r175_c131 bl[131] br[131] wl[175] vdd gnd cell_6t
Xbit_r176_c131 bl[131] br[131] wl[176] vdd gnd cell_6t
Xbit_r177_c131 bl[131] br[131] wl[177] vdd gnd cell_6t
Xbit_r178_c131 bl[131] br[131] wl[178] vdd gnd cell_6t
Xbit_r179_c131 bl[131] br[131] wl[179] vdd gnd cell_6t
Xbit_r180_c131 bl[131] br[131] wl[180] vdd gnd cell_6t
Xbit_r181_c131 bl[131] br[131] wl[181] vdd gnd cell_6t
Xbit_r182_c131 bl[131] br[131] wl[182] vdd gnd cell_6t
Xbit_r183_c131 bl[131] br[131] wl[183] vdd gnd cell_6t
Xbit_r184_c131 bl[131] br[131] wl[184] vdd gnd cell_6t
Xbit_r185_c131 bl[131] br[131] wl[185] vdd gnd cell_6t
Xbit_r186_c131 bl[131] br[131] wl[186] vdd gnd cell_6t
Xbit_r187_c131 bl[131] br[131] wl[187] vdd gnd cell_6t
Xbit_r188_c131 bl[131] br[131] wl[188] vdd gnd cell_6t
Xbit_r189_c131 bl[131] br[131] wl[189] vdd gnd cell_6t
Xbit_r190_c131 bl[131] br[131] wl[190] vdd gnd cell_6t
Xbit_r191_c131 bl[131] br[131] wl[191] vdd gnd cell_6t
Xbit_r192_c131 bl[131] br[131] wl[192] vdd gnd cell_6t
Xbit_r193_c131 bl[131] br[131] wl[193] vdd gnd cell_6t
Xbit_r194_c131 bl[131] br[131] wl[194] vdd gnd cell_6t
Xbit_r195_c131 bl[131] br[131] wl[195] vdd gnd cell_6t
Xbit_r196_c131 bl[131] br[131] wl[196] vdd gnd cell_6t
Xbit_r197_c131 bl[131] br[131] wl[197] vdd gnd cell_6t
Xbit_r198_c131 bl[131] br[131] wl[198] vdd gnd cell_6t
Xbit_r199_c131 bl[131] br[131] wl[199] vdd gnd cell_6t
Xbit_r200_c131 bl[131] br[131] wl[200] vdd gnd cell_6t
Xbit_r201_c131 bl[131] br[131] wl[201] vdd gnd cell_6t
Xbit_r202_c131 bl[131] br[131] wl[202] vdd gnd cell_6t
Xbit_r203_c131 bl[131] br[131] wl[203] vdd gnd cell_6t
Xbit_r204_c131 bl[131] br[131] wl[204] vdd gnd cell_6t
Xbit_r205_c131 bl[131] br[131] wl[205] vdd gnd cell_6t
Xbit_r206_c131 bl[131] br[131] wl[206] vdd gnd cell_6t
Xbit_r207_c131 bl[131] br[131] wl[207] vdd gnd cell_6t
Xbit_r208_c131 bl[131] br[131] wl[208] vdd gnd cell_6t
Xbit_r209_c131 bl[131] br[131] wl[209] vdd gnd cell_6t
Xbit_r210_c131 bl[131] br[131] wl[210] vdd gnd cell_6t
Xbit_r211_c131 bl[131] br[131] wl[211] vdd gnd cell_6t
Xbit_r212_c131 bl[131] br[131] wl[212] vdd gnd cell_6t
Xbit_r213_c131 bl[131] br[131] wl[213] vdd gnd cell_6t
Xbit_r214_c131 bl[131] br[131] wl[214] vdd gnd cell_6t
Xbit_r215_c131 bl[131] br[131] wl[215] vdd gnd cell_6t
Xbit_r216_c131 bl[131] br[131] wl[216] vdd gnd cell_6t
Xbit_r217_c131 bl[131] br[131] wl[217] vdd gnd cell_6t
Xbit_r218_c131 bl[131] br[131] wl[218] vdd gnd cell_6t
Xbit_r219_c131 bl[131] br[131] wl[219] vdd gnd cell_6t
Xbit_r220_c131 bl[131] br[131] wl[220] vdd gnd cell_6t
Xbit_r221_c131 bl[131] br[131] wl[221] vdd gnd cell_6t
Xbit_r222_c131 bl[131] br[131] wl[222] vdd gnd cell_6t
Xbit_r223_c131 bl[131] br[131] wl[223] vdd gnd cell_6t
Xbit_r224_c131 bl[131] br[131] wl[224] vdd gnd cell_6t
Xbit_r225_c131 bl[131] br[131] wl[225] vdd gnd cell_6t
Xbit_r226_c131 bl[131] br[131] wl[226] vdd gnd cell_6t
Xbit_r227_c131 bl[131] br[131] wl[227] vdd gnd cell_6t
Xbit_r228_c131 bl[131] br[131] wl[228] vdd gnd cell_6t
Xbit_r229_c131 bl[131] br[131] wl[229] vdd gnd cell_6t
Xbit_r230_c131 bl[131] br[131] wl[230] vdd gnd cell_6t
Xbit_r231_c131 bl[131] br[131] wl[231] vdd gnd cell_6t
Xbit_r232_c131 bl[131] br[131] wl[232] vdd gnd cell_6t
Xbit_r233_c131 bl[131] br[131] wl[233] vdd gnd cell_6t
Xbit_r234_c131 bl[131] br[131] wl[234] vdd gnd cell_6t
Xbit_r235_c131 bl[131] br[131] wl[235] vdd gnd cell_6t
Xbit_r236_c131 bl[131] br[131] wl[236] vdd gnd cell_6t
Xbit_r237_c131 bl[131] br[131] wl[237] vdd gnd cell_6t
Xbit_r238_c131 bl[131] br[131] wl[238] vdd gnd cell_6t
Xbit_r239_c131 bl[131] br[131] wl[239] vdd gnd cell_6t
Xbit_r240_c131 bl[131] br[131] wl[240] vdd gnd cell_6t
Xbit_r241_c131 bl[131] br[131] wl[241] vdd gnd cell_6t
Xbit_r242_c131 bl[131] br[131] wl[242] vdd gnd cell_6t
Xbit_r243_c131 bl[131] br[131] wl[243] vdd gnd cell_6t
Xbit_r244_c131 bl[131] br[131] wl[244] vdd gnd cell_6t
Xbit_r245_c131 bl[131] br[131] wl[245] vdd gnd cell_6t
Xbit_r246_c131 bl[131] br[131] wl[246] vdd gnd cell_6t
Xbit_r247_c131 bl[131] br[131] wl[247] vdd gnd cell_6t
Xbit_r248_c131 bl[131] br[131] wl[248] vdd gnd cell_6t
Xbit_r249_c131 bl[131] br[131] wl[249] vdd gnd cell_6t
Xbit_r250_c131 bl[131] br[131] wl[250] vdd gnd cell_6t
Xbit_r251_c131 bl[131] br[131] wl[251] vdd gnd cell_6t
Xbit_r252_c131 bl[131] br[131] wl[252] vdd gnd cell_6t
Xbit_r253_c131 bl[131] br[131] wl[253] vdd gnd cell_6t
Xbit_r254_c131 bl[131] br[131] wl[254] vdd gnd cell_6t
Xbit_r255_c131 bl[131] br[131] wl[255] vdd gnd cell_6t
Xbit_r0_c132 bl[132] br[132] wl[0] vdd gnd cell_6t
Xbit_r1_c132 bl[132] br[132] wl[1] vdd gnd cell_6t
Xbit_r2_c132 bl[132] br[132] wl[2] vdd gnd cell_6t
Xbit_r3_c132 bl[132] br[132] wl[3] vdd gnd cell_6t
Xbit_r4_c132 bl[132] br[132] wl[4] vdd gnd cell_6t
Xbit_r5_c132 bl[132] br[132] wl[5] vdd gnd cell_6t
Xbit_r6_c132 bl[132] br[132] wl[6] vdd gnd cell_6t
Xbit_r7_c132 bl[132] br[132] wl[7] vdd gnd cell_6t
Xbit_r8_c132 bl[132] br[132] wl[8] vdd gnd cell_6t
Xbit_r9_c132 bl[132] br[132] wl[9] vdd gnd cell_6t
Xbit_r10_c132 bl[132] br[132] wl[10] vdd gnd cell_6t
Xbit_r11_c132 bl[132] br[132] wl[11] vdd gnd cell_6t
Xbit_r12_c132 bl[132] br[132] wl[12] vdd gnd cell_6t
Xbit_r13_c132 bl[132] br[132] wl[13] vdd gnd cell_6t
Xbit_r14_c132 bl[132] br[132] wl[14] vdd gnd cell_6t
Xbit_r15_c132 bl[132] br[132] wl[15] vdd gnd cell_6t
Xbit_r16_c132 bl[132] br[132] wl[16] vdd gnd cell_6t
Xbit_r17_c132 bl[132] br[132] wl[17] vdd gnd cell_6t
Xbit_r18_c132 bl[132] br[132] wl[18] vdd gnd cell_6t
Xbit_r19_c132 bl[132] br[132] wl[19] vdd gnd cell_6t
Xbit_r20_c132 bl[132] br[132] wl[20] vdd gnd cell_6t
Xbit_r21_c132 bl[132] br[132] wl[21] vdd gnd cell_6t
Xbit_r22_c132 bl[132] br[132] wl[22] vdd gnd cell_6t
Xbit_r23_c132 bl[132] br[132] wl[23] vdd gnd cell_6t
Xbit_r24_c132 bl[132] br[132] wl[24] vdd gnd cell_6t
Xbit_r25_c132 bl[132] br[132] wl[25] vdd gnd cell_6t
Xbit_r26_c132 bl[132] br[132] wl[26] vdd gnd cell_6t
Xbit_r27_c132 bl[132] br[132] wl[27] vdd gnd cell_6t
Xbit_r28_c132 bl[132] br[132] wl[28] vdd gnd cell_6t
Xbit_r29_c132 bl[132] br[132] wl[29] vdd gnd cell_6t
Xbit_r30_c132 bl[132] br[132] wl[30] vdd gnd cell_6t
Xbit_r31_c132 bl[132] br[132] wl[31] vdd gnd cell_6t
Xbit_r32_c132 bl[132] br[132] wl[32] vdd gnd cell_6t
Xbit_r33_c132 bl[132] br[132] wl[33] vdd gnd cell_6t
Xbit_r34_c132 bl[132] br[132] wl[34] vdd gnd cell_6t
Xbit_r35_c132 bl[132] br[132] wl[35] vdd gnd cell_6t
Xbit_r36_c132 bl[132] br[132] wl[36] vdd gnd cell_6t
Xbit_r37_c132 bl[132] br[132] wl[37] vdd gnd cell_6t
Xbit_r38_c132 bl[132] br[132] wl[38] vdd gnd cell_6t
Xbit_r39_c132 bl[132] br[132] wl[39] vdd gnd cell_6t
Xbit_r40_c132 bl[132] br[132] wl[40] vdd gnd cell_6t
Xbit_r41_c132 bl[132] br[132] wl[41] vdd gnd cell_6t
Xbit_r42_c132 bl[132] br[132] wl[42] vdd gnd cell_6t
Xbit_r43_c132 bl[132] br[132] wl[43] vdd gnd cell_6t
Xbit_r44_c132 bl[132] br[132] wl[44] vdd gnd cell_6t
Xbit_r45_c132 bl[132] br[132] wl[45] vdd gnd cell_6t
Xbit_r46_c132 bl[132] br[132] wl[46] vdd gnd cell_6t
Xbit_r47_c132 bl[132] br[132] wl[47] vdd gnd cell_6t
Xbit_r48_c132 bl[132] br[132] wl[48] vdd gnd cell_6t
Xbit_r49_c132 bl[132] br[132] wl[49] vdd gnd cell_6t
Xbit_r50_c132 bl[132] br[132] wl[50] vdd gnd cell_6t
Xbit_r51_c132 bl[132] br[132] wl[51] vdd gnd cell_6t
Xbit_r52_c132 bl[132] br[132] wl[52] vdd gnd cell_6t
Xbit_r53_c132 bl[132] br[132] wl[53] vdd gnd cell_6t
Xbit_r54_c132 bl[132] br[132] wl[54] vdd gnd cell_6t
Xbit_r55_c132 bl[132] br[132] wl[55] vdd gnd cell_6t
Xbit_r56_c132 bl[132] br[132] wl[56] vdd gnd cell_6t
Xbit_r57_c132 bl[132] br[132] wl[57] vdd gnd cell_6t
Xbit_r58_c132 bl[132] br[132] wl[58] vdd gnd cell_6t
Xbit_r59_c132 bl[132] br[132] wl[59] vdd gnd cell_6t
Xbit_r60_c132 bl[132] br[132] wl[60] vdd gnd cell_6t
Xbit_r61_c132 bl[132] br[132] wl[61] vdd gnd cell_6t
Xbit_r62_c132 bl[132] br[132] wl[62] vdd gnd cell_6t
Xbit_r63_c132 bl[132] br[132] wl[63] vdd gnd cell_6t
Xbit_r64_c132 bl[132] br[132] wl[64] vdd gnd cell_6t
Xbit_r65_c132 bl[132] br[132] wl[65] vdd gnd cell_6t
Xbit_r66_c132 bl[132] br[132] wl[66] vdd gnd cell_6t
Xbit_r67_c132 bl[132] br[132] wl[67] vdd gnd cell_6t
Xbit_r68_c132 bl[132] br[132] wl[68] vdd gnd cell_6t
Xbit_r69_c132 bl[132] br[132] wl[69] vdd gnd cell_6t
Xbit_r70_c132 bl[132] br[132] wl[70] vdd gnd cell_6t
Xbit_r71_c132 bl[132] br[132] wl[71] vdd gnd cell_6t
Xbit_r72_c132 bl[132] br[132] wl[72] vdd gnd cell_6t
Xbit_r73_c132 bl[132] br[132] wl[73] vdd gnd cell_6t
Xbit_r74_c132 bl[132] br[132] wl[74] vdd gnd cell_6t
Xbit_r75_c132 bl[132] br[132] wl[75] vdd gnd cell_6t
Xbit_r76_c132 bl[132] br[132] wl[76] vdd gnd cell_6t
Xbit_r77_c132 bl[132] br[132] wl[77] vdd gnd cell_6t
Xbit_r78_c132 bl[132] br[132] wl[78] vdd gnd cell_6t
Xbit_r79_c132 bl[132] br[132] wl[79] vdd gnd cell_6t
Xbit_r80_c132 bl[132] br[132] wl[80] vdd gnd cell_6t
Xbit_r81_c132 bl[132] br[132] wl[81] vdd gnd cell_6t
Xbit_r82_c132 bl[132] br[132] wl[82] vdd gnd cell_6t
Xbit_r83_c132 bl[132] br[132] wl[83] vdd gnd cell_6t
Xbit_r84_c132 bl[132] br[132] wl[84] vdd gnd cell_6t
Xbit_r85_c132 bl[132] br[132] wl[85] vdd gnd cell_6t
Xbit_r86_c132 bl[132] br[132] wl[86] vdd gnd cell_6t
Xbit_r87_c132 bl[132] br[132] wl[87] vdd gnd cell_6t
Xbit_r88_c132 bl[132] br[132] wl[88] vdd gnd cell_6t
Xbit_r89_c132 bl[132] br[132] wl[89] vdd gnd cell_6t
Xbit_r90_c132 bl[132] br[132] wl[90] vdd gnd cell_6t
Xbit_r91_c132 bl[132] br[132] wl[91] vdd gnd cell_6t
Xbit_r92_c132 bl[132] br[132] wl[92] vdd gnd cell_6t
Xbit_r93_c132 bl[132] br[132] wl[93] vdd gnd cell_6t
Xbit_r94_c132 bl[132] br[132] wl[94] vdd gnd cell_6t
Xbit_r95_c132 bl[132] br[132] wl[95] vdd gnd cell_6t
Xbit_r96_c132 bl[132] br[132] wl[96] vdd gnd cell_6t
Xbit_r97_c132 bl[132] br[132] wl[97] vdd gnd cell_6t
Xbit_r98_c132 bl[132] br[132] wl[98] vdd gnd cell_6t
Xbit_r99_c132 bl[132] br[132] wl[99] vdd gnd cell_6t
Xbit_r100_c132 bl[132] br[132] wl[100] vdd gnd cell_6t
Xbit_r101_c132 bl[132] br[132] wl[101] vdd gnd cell_6t
Xbit_r102_c132 bl[132] br[132] wl[102] vdd gnd cell_6t
Xbit_r103_c132 bl[132] br[132] wl[103] vdd gnd cell_6t
Xbit_r104_c132 bl[132] br[132] wl[104] vdd gnd cell_6t
Xbit_r105_c132 bl[132] br[132] wl[105] vdd gnd cell_6t
Xbit_r106_c132 bl[132] br[132] wl[106] vdd gnd cell_6t
Xbit_r107_c132 bl[132] br[132] wl[107] vdd gnd cell_6t
Xbit_r108_c132 bl[132] br[132] wl[108] vdd gnd cell_6t
Xbit_r109_c132 bl[132] br[132] wl[109] vdd gnd cell_6t
Xbit_r110_c132 bl[132] br[132] wl[110] vdd gnd cell_6t
Xbit_r111_c132 bl[132] br[132] wl[111] vdd gnd cell_6t
Xbit_r112_c132 bl[132] br[132] wl[112] vdd gnd cell_6t
Xbit_r113_c132 bl[132] br[132] wl[113] vdd gnd cell_6t
Xbit_r114_c132 bl[132] br[132] wl[114] vdd gnd cell_6t
Xbit_r115_c132 bl[132] br[132] wl[115] vdd gnd cell_6t
Xbit_r116_c132 bl[132] br[132] wl[116] vdd gnd cell_6t
Xbit_r117_c132 bl[132] br[132] wl[117] vdd gnd cell_6t
Xbit_r118_c132 bl[132] br[132] wl[118] vdd gnd cell_6t
Xbit_r119_c132 bl[132] br[132] wl[119] vdd gnd cell_6t
Xbit_r120_c132 bl[132] br[132] wl[120] vdd gnd cell_6t
Xbit_r121_c132 bl[132] br[132] wl[121] vdd gnd cell_6t
Xbit_r122_c132 bl[132] br[132] wl[122] vdd gnd cell_6t
Xbit_r123_c132 bl[132] br[132] wl[123] vdd gnd cell_6t
Xbit_r124_c132 bl[132] br[132] wl[124] vdd gnd cell_6t
Xbit_r125_c132 bl[132] br[132] wl[125] vdd gnd cell_6t
Xbit_r126_c132 bl[132] br[132] wl[126] vdd gnd cell_6t
Xbit_r127_c132 bl[132] br[132] wl[127] vdd gnd cell_6t
Xbit_r128_c132 bl[132] br[132] wl[128] vdd gnd cell_6t
Xbit_r129_c132 bl[132] br[132] wl[129] vdd gnd cell_6t
Xbit_r130_c132 bl[132] br[132] wl[130] vdd gnd cell_6t
Xbit_r131_c132 bl[132] br[132] wl[131] vdd gnd cell_6t
Xbit_r132_c132 bl[132] br[132] wl[132] vdd gnd cell_6t
Xbit_r133_c132 bl[132] br[132] wl[133] vdd gnd cell_6t
Xbit_r134_c132 bl[132] br[132] wl[134] vdd gnd cell_6t
Xbit_r135_c132 bl[132] br[132] wl[135] vdd gnd cell_6t
Xbit_r136_c132 bl[132] br[132] wl[136] vdd gnd cell_6t
Xbit_r137_c132 bl[132] br[132] wl[137] vdd gnd cell_6t
Xbit_r138_c132 bl[132] br[132] wl[138] vdd gnd cell_6t
Xbit_r139_c132 bl[132] br[132] wl[139] vdd gnd cell_6t
Xbit_r140_c132 bl[132] br[132] wl[140] vdd gnd cell_6t
Xbit_r141_c132 bl[132] br[132] wl[141] vdd gnd cell_6t
Xbit_r142_c132 bl[132] br[132] wl[142] vdd gnd cell_6t
Xbit_r143_c132 bl[132] br[132] wl[143] vdd gnd cell_6t
Xbit_r144_c132 bl[132] br[132] wl[144] vdd gnd cell_6t
Xbit_r145_c132 bl[132] br[132] wl[145] vdd gnd cell_6t
Xbit_r146_c132 bl[132] br[132] wl[146] vdd gnd cell_6t
Xbit_r147_c132 bl[132] br[132] wl[147] vdd gnd cell_6t
Xbit_r148_c132 bl[132] br[132] wl[148] vdd gnd cell_6t
Xbit_r149_c132 bl[132] br[132] wl[149] vdd gnd cell_6t
Xbit_r150_c132 bl[132] br[132] wl[150] vdd gnd cell_6t
Xbit_r151_c132 bl[132] br[132] wl[151] vdd gnd cell_6t
Xbit_r152_c132 bl[132] br[132] wl[152] vdd gnd cell_6t
Xbit_r153_c132 bl[132] br[132] wl[153] vdd gnd cell_6t
Xbit_r154_c132 bl[132] br[132] wl[154] vdd gnd cell_6t
Xbit_r155_c132 bl[132] br[132] wl[155] vdd gnd cell_6t
Xbit_r156_c132 bl[132] br[132] wl[156] vdd gnd cell_6t
Xbit_r157_c132 bl[132] br[132] wl[157] vdd gnd cell_6t
Xbit_r158_c132 bl[132] br[132] wl[158] vdd gnd cell_6t
Xbit_r159_c132 bl[132] br[132] wl[159] vdd gnd cell_6t
Xbit_r160_c132 bl[132] br[132] wl[160] vdd gnd cell_6t
Xbit_r161_c132 bl[132] br[132] wl[161] vdd gnd cell_6t
Xbit_r162_c132 bl[132] br[132] wl[162] vdd gnd cell_6t
Xbit_r163_c132 bl[132] br[132] wl[163] vdd gnd cell_6t
Xbit_r164_c132 bl[132] br[132] wl[164] vdd gnd cell_6t
Xbit_r165_c132 bl[132] br[132] wl[165] vdd gnd cell_6t
Xbit_r166_c132 bl[132] br[132] wl[166] vdd gnd cell_6t
Xbit_r167_c132 bl[132] br[132] wl[167] vdd gnd cell_6t
Xbit_r168_c132 bl[132] br[132] wl[168] vdd gnd cell_6t
Xbit_r169_c132 bl[132] br[132] wl[169] vdd gnd cell_6t
Xbit_r170_c132 bl[132] br[132] wl[170] vdd gnd cell_6t
Xbit_r171_c132 bl[132] br[132] wl[171] vdd gnd cell_6t
Xbit_r172_c132 bl[132] br[132] wl[172] vdd gnd cell_6t
Xbit_r173_c132 bl[132] br[132] wl[173] vdd gnd cell_6t
Xbit_r174_c132 bl[132] br[132] wl[174] vdd gnd cell_6t
Xbit_r175_c132 bl[132] br[132] wl[175] vdd gnd cell_6t
Xbit_r176_c132 bl[132] br[132] wl[176] vdd gnd cell_6t
Xbit_r177_c132 bl[132] br[132] wl[177] vdd gnd cell_6t
Xbit_r178_c132 bl[132] br[132] wl[178] vdd gnd cell_6t
Xbit_r179_c132 bl[132] br[132] wl[179] vdd gnd cell_6t
Xbit_r180_c132 bl[132] br[132] wl[180] vdd gnd cell_6t
Xbit_r181_c132 bl[132] br[132] wl[181] vdd gnd cell_6t
Xbit_r182_c132 bl[132] br[132] wl[182] vdd gnd cell_6t
Xbit_r183_c132 bl[132] br[132] wl[183] vdd gnd cell_6t
Xbit_r184_c132 bl[132] br[132] wl[184] vdd gnd cell_6t
Xbit_r185_c132 bl[132] br[132] wl[185] vdd gnd cell_6t
Xbit_r186_c132 bl[132] br[132] wl[186] vdd gnd cell_6t
Xbit_r187_c132 bl[132] br[132] wl[187] vdd gnd cell_6t
Xbit_r188_c132 bl[132] br[132] wl[188] vdd gnd cell_6t
Xbit_r189_c132 bl[132] br[132] wl[189] vdd gnd cell_6t
Xbit_r190_c132 bl[132] br[132] wl[190] vdd gnd cell_6t
Xbit_r191_c132 bl[132] br[132] wl[191] vdd gnd cell_6t
Xbit_r192_c132 bl[132] br[132] wl[192] vdd gnd cell_6t
Xbit_r193_c132 bl[132] br[132] wl[193] vdd gnd cell_6t
Xbit_r194_c132 bl[132] br[132] wl[194] vdd gnd cell_6t
Xbit_r195_c132 bl[132] br[132] wl[195] vdd gnd cell_6t
Xbit_r196_c132 bl[132] br[132] wl[196] vdd gnd cell_6t
Xbit_r197_c132 bl[132] br[132] wl[197] vdd gnd cell_6t
Xbit_r198_c132 bl[132] br[132] wl[198] vdd gnd cell_6t
Xbit_r199_c132 bl[132] br[132] wl[199] vdd gnd cell_6t
Xbit_r200_c132 bl[132] br[132] wl[200] vdd gnd cell_6t
Xbit_r201_c132 bl[132] br[132] wl[201] vdd gnd cell_6t
Xbit_r202_c132 bl[132] br[132] wl[202] vdd gnd cell_6t
Xbit_r203_c132 bl[132] br[132] wl[203] vdd gnd cell_6t
Xbit_r204_c132 bl[132] br[132] wl[204] vdd gnd cell_6t
Xbit_r205_c132 bl[132] br[132] wl[205] vdd gnd cell_6t
Xbit_r206_c132 bl[132] br[132] wl[206] vdd gnd cell_6t
Xbit_r207_c132 bl[132] br[132] wl[207] vdd gnd cell_6t
Xbit_r208_c132 bl[132] br[132] wl[208] vdd gnd cell_6t
Xbit_r209_c132 bl[132] br[132] wl[209] vdd gnd cell_6t
Xbit_r210_c132 bl[132] br[132] wl[210] vdd gnd cell_6t
Xbit_r211_c132 bl[132] br[132] wl[211] vdd gnd cell_6t
Xbit_r212_c132 bl[132] br[132] wl[212] vdd gnd cell_6t
Xbit_r213_c132 bl[132] br[132] wl[213] vdd gnd cell_6t
Xbit_r214_c132 bl[132] br[132] wl[214] vdd gnd cell_6t
Xbit_r215_c132 bl[132] br[132] wl[215] vdd gnd cell_6t
Xbit_r216_c132 bl[132] br[132] wl[216] vdd gnd cell_6t
Xbit_r217_c132 bl[132] br[132] wl[217] vdd gnd cell_6t
Xbit_r218_c132 bl[132] br[132] wl[218] vdd gnd cell_6t
Xbit_r219_c132 bl[132] br[132] wl[219] vdd gnd cell_6t
Xbit_r220_c132 bl[132] br[132] wl[220] vdd gnd cell_6t
Xbit_r221_c132 bl[132] br[132] wl[221] vdd gnd cell_6t
Xbit_r222_c132 bl[132] br[132] wl[222] vdd gnd cell_6t
Xbit_r223_c132 bl[132] br[132] wl[223] vdd gnd cell_6t
Xbit_r224_c132 bl[132] br[132] wl[224] vdd gnd cell_6t
Xbit_r225_c132 bl[132] br[132] wl[225] vdd gnd cell_6t
Xbit_r226_c132 bl[132] br[132] wl[226] vdd gnd cell_6t
Xbit_r227_c132 bl[132] br[132] wl[227] vdd gnd cell_6t
Xbit_r228_c132 bl[132] br[132] wl[228] vdd gnd cell_6t
Xbit_r229_c132 bl[132] br[132] wl[229] vdd gnd cell_6t
Xbit_r230_c132 bl[132] br[132] wl[230] vdd gnd cell_6t
Xbit_r231_c132 bl[132] br[132] wl[231] vdd gnd cell_6t
Xbit_r232_c132 bl[132] br[132] wl[232] vdd gnd cell_6t
Xbit_r233_c132 bl[132] br[132] wl[233] vdd gnd cell_6t
Xbit_r234_c132 bl[132] br[132] wl[234] vdd gnd cell_6t
Xbit_r235_c132 bl[132] br[132] wl[235] vdd gnd cell_6t
Xbit_r236_c132 bl[132] br[132] wl[236] vdd gnd cell_6t
Xbit_r237_c132 bl[132] br[132] wl[237] vdd gnd cell_6t
Xbit_r238_c132 bl[132] br[132] wl[238] vdd gnd cell_6t
Xbit_r239_c132 bl[132] br[132] wl[239] vdd gnd cell_6t
Xbit_r240_c132 bl[132] br[132] wl[240] vdd gnd cell_6t
Xbit_r241_c132 bl[132] br[132] wl[241] vdd gnd cell_6t
Xbit_r242_c132 bl[132] br[132] wl[242] vdd gnd cell_6t
Xbit_r243_c132 bl[132] br[132] wl[243] vdd gnd cell_6t
Xbit_r244_c132 bl[132] br[132] wl[244] vdd gnd cell_6t
Xbit_r245_c132 bl[132] br[132] wl[245] vdd gnd cell_6t
Xbit_r246_c132 bl[132] br[132] wl[246] vdd gnd cell_6t
Xbit_r247_c132 bl[132] br[132] wl[247] vdd gnd cell_6t
Xbit_r248_c132 bl[132] br[132] wl[248] vdd gnd cell_6t
Xbit_r249_c132 bl[132] br[132] wl[249] vdd gnd cell_6t
Xbit_r250_c132 bl[132] br[132] wl[250] vdd gnd cell_6t
Xbit_r251_c132 bl[132] br[132] wl[251] vdd gnd cell_6t
Xbit_r252_c132 bl[132] br[132] wl[252] vdd gnd cell_6t
Xbit_r253_c132 bl[132] br[132] wl[253] vdd gnd cell_6t
Xbit_r254_c132 bl[132] br[132] wl[254] vdd gnd cell_6t
Xbit_r255_c132 bl[132] br[132] wl[255] vdd gnd cell_6t
Xbit_r0_c133 bl[133] br[133] wl[0] vdd gnd cell_6t
Xbit_r1_c133 bl[133] br[133] wl[1] vdd gnd cell_6t
Xbit_r2_c133 bl[133] br[133] wl[2] vdd gnd cell_6t
Xbit_r3_c133 bl[133] br[133] wl[3] vdd gnd cell_6t
Xbit_r4_c133 bl[133] br[133] wl[4] vdd gnd cell_6t
Xbit_r5_c133 bl[133] br[133] wl[5] vdd gnd cell_6t
Xbit_r6_c133 bl[133] br[133] wl[6] vdd gnd cell_6t
Xbit_r7_c133 bl[133] br[133] wl[7] vdd gnd cell_6t
Xbit_r8_c133 bl[133] br[133] wl[8] vdd gnd cell_6t
Xbit_r9_c133 bl[133] br[133] wl[9] vdd gnd cell_6t
Xbit_r10_c133 bl[133] br[133] wl[10] vdd gnd cell_6t
Xbit_r11_c133 bl[133] br[133] wl[11] vdd gnd cell_6t
Xbit_r12_c133 bl[133] br[133] wl[12] vdd gnd cell_6t
Xbit_r13_c133 bl[133] br[133] wl[13] vdd gnd cell_6t
Xbit_r14_c133 bl[133] br[133] wl[14] vdd gnd cell_6t
Xbit_r15_c133 bl[133] br[133] wl[15] vdd gnd cell_6t
Xbit_r16_c133 bl[133] br[133] wl[16] vdd gnd cell_6t
Xbit_r17_c133 bl[133] br[133] wl[17] vdd gnd cell_6t
Xbit_r18_c133 bl[133] br[133] wl[18] vdd gnd cell_6t
Xbit_r19_c133 bl[133] br[133] wl[19] vdd gnd cell_6t
Xbit_r20_c133 bl[133] br[133] wl[20] vdd gnd cell_6t
Xbit_r21_c133 bl[133] br[133] wl[21] vdd gnd cell_6t
Xbit_r22_c133 bl[133] br[133] wl[22] vdd gnd cell_6t
Xbit_r23_c133 bl[133] br[133] wl[23] vdd gnd cell_6t
Xbit_r24_c133 bl[133] br[133] wl[24] vdd gnd cell_6t
Xbit_r25_c133 bl[133] br[133] wl[25] vdd gnd cell_6t
Xbit_r26_c133 bl[133] br[133] wl[26] vdd gnd cell_6t
Xbit_r27_c133 bl[133] br[133] wl[27] vdd gnd cell_6t
Xbit_r28_c133 bl[133] br[133] wl[28] vdd gnd cell_6t
Xbit_r29_c133 bl[133] br[133] wl[29] vdd gnd cell_6t
Xbit_r30_c133 bl[133] br[133] wl[30] vdd gnd cell_6t
Xbit_r31_c133 bl[133] br[133] wl[31] vdd gnd cell_6t
Xbit_r32_c133 bl[133] br[133] wl[32] vdd gnd cell_6t
Xbit_r33_c133 bl[133] br[133] wl[33] vdd gnd cell_6t
Xbit_r34_c133 bl[133] br[133] wl[34] vdd gnd cell_6t
Xbit_r35_c133 bl[133] br[133] wl[35] vdd gnd cell_6t
Xbit_r36_c133 bl[133] br[133] wl[36] vdd gnd cell_6t
Xbit_r37_c133 bl[133] br[133] wl[37] vdd gnd cell_6t
Xbit_r38_c133 bl[133] br[133] wl[38] vdd gnd cell_6t
Xbit_r39_c133 bl[133] br[133] wl[39] vdd gnd cell_6t
Xbit_r40_c133 bl[133] br[133] wl[40] vdd gnd cell_6t
Xbit_r41_c133 bl[133] br[133] wl[41] vdd gnd cell_6t
Xbit_r42_c133 bl[133] br[133] wl[42] vdd gnd cell_6t
Xbit_r43_c133 bl[133] br[133] wl[43] vdd gnd cell_6t
Xbit_r44_c133 bl[133] br[133] wl[44] vdd gnd cell_6t
Xbit_r45_c133 bl[133] br[133] wl[45] vdd gnd cell_6t
Xbit_r46_c133 bl[133] br[133] wl[46] vdd gnd cell_6t
Xbit_r47_c133 bl[133] br[133] wl[47] vdd gnd cell_6t
Xbit_r48_c133 bl[133] br[133] wl[48] vdd gnd cell_6t
Xbit_r49_c133 bl[133] br[133] wl[49] vdd gnd cell_6t
Xbit_r50_c133 bl[133] br[133] wl[50] vdd gnd cell_6t
Xbit_r51_c133 bl[133] br[133] wl[51] vdd gnd cell_6t
Xbit_r52_c133 bl[133] br[133] wl[52] vdd gnd cell_6t
Xbit_r53_c133 bl[133] br[133] wl[53] vdd gnd cell_6t
Xbit_r54_c133 bl[133] br[133] wl[54] vdd gnd cell_6t
Xbit_r55_c133 bl[133] br[133] wl[55] vdd gnd cell_6t
Xbit_r56_c133 bl[133] br[133] wl[56] vdd gnd cell_6t
Xbit_r57_c133 bl[133] br[133] wl[57] vdd gnd cell_6t
Xbit_r58_c133 bl[133] br[133] wl[58] vdd gnd cell_6t
Xbit_r59_c133 bl[133] br[133] wl[59] vdd gnd cell_6t
Xbit_r60_c133 bl[133] br[133] wl[60] vdd gnd cell_6t
Xbit_r61_c133 bl[133] br[133] wl[61] vdd gnd cell_6t
Xbit_r62_c133 bl[133] br[133] wl[62] vdd gnd cell_6t
Xbit_r63_c133 bl[133] br[133] wl[63] vdd gnd cell_6t
Xbit_r64_c133 bl[133] br[133] wl[64] vdd gnd cell_6t
Xbit_r65_c133 bl[133] br[133] wl[65] vdd gnd cell_6t
Xbit_r66_c133 bl[133] br[133] wl[66] vdd gnd cell_6t
Xbit_r67_c133 bl[133] br[133] wl[67] vdd gnd cell_6t
Xbit_r68_c133 bl[133] br[133] wl[68] vdd gnd cell_6t
Xbit_r69_c133 bl[133] br[133] wl[69] vdd gnd cell_6t
Xbit_r70_c133 bl[133] br[133] wl[70] vdd gnd cell_6t
Xbit_r71_c133 bl[133] br[133] wl[71] vdd gnd cell_6t
Xbit_r72_c133 bl[133] br[133] wl[72] vdd gnd cell_6t
Xbit_r73_c133 bl[133] br[133] wl[73] vdd gnd cell_6t
Xbit_r74_c133 bl[133] br[133] wl[74] vdd gnd cell_6t
Xbit_r75_c133 bl[133] br[133] wl[75] vdd gnd cell_6t
Xbit_r76_c133 bl[133] br[133] wl[76] vdd gnd cell_6t
Xbit_r77_c133 bl[133] br[133] wl[77] vdd gnd cell_6t
Xbit_r78_c133 bl[133] br[133] wl[78] vdd gnd cell_6t
Xbit_r79_c133 bl[133] br[133] wl[79] vdd gnd cell_6t
Xbit_r80_c133 bl[133] br[133] wl[80] vdd gnd cell_6t
Xbit_r81_c133 bl[133] br[133] wl[81] vdd gnd cell_6t
Xbit_r82_c133 bl[133] br[133] wl[82] vdd gnd cell_6t
Xbit_r83_c133 bl[133] br[133] wl[83] vdd gnd cell_6t
Xbit_r84_c133 bl[133] br[133] wl[84] vdd gnd cell_6t
Xbit_r85_c133 bl[133] br[133] wl[85] vdd gnd cell_6t
Xbit_r86_c133 bl[133] br[133] wl[86] vdd gnd cell_6t
Xbit_r87_c133 bl[133] br[133] wl[87] vdd gnd cell_6t
Xbit_r88_c133 bl[133] br[133] wl[88] vdd gnd cell_6t
Xbit_r89_c133 bl[133] br[133] wl[89] vdd gnd cell_6t
Xbit_r90_c133 bl[133] br[133] wl[90] vdd gnd cell_6t
Xbit_r91_c133 bl[133] br[133] wl[91] vdd gnd cell_6t
Xbit_r92_c133 bl[133] br[133] wl[92] vdd gnd cell_6t
Xbit_r93_c133 bl[133] br[133] wl[93] vdd gnd cell_6t
Xbit_r94_c133 bl[133] br[133] wl[94] vdd gnd cell_6t
Xbit_r95_c133 bl[133] br[133] wl[95] vdd gnd cell_6t
Xbit_r96_c133 bl[133] br[133] wl[96] vdd gnd cell_6t
Xbit_r97_c133 bl[133] br[133] wl[97] vdd gnd cell_6t
Xbit_r98_c133 bl[133] br[133] wl[98] vdd gnd cell_6t
Xbit_r99_c133 bl[133] br[133] wl[99] vdd gnd cell_6t
Xbit_r100_c133 bl[133] br[133] wl[100] vdd gnd cell_6t
Xbit_r101_c133 bl[133] br[133] wl[101] vdd gnd cell_6t
Xbit_r102_c133 bl[133] br[133] wl[102] vdd gnd cell_6t
Xbit_r103_c133 bl[133] br[133] wl[103] vdd gnd cell_6t
Xbit_r104_c133 bl[133] br[133] wl[104] vdd gnd cell_6t
Xbit_r105_c133 bl[133] br[133] wl[105] vdd gnd cell_6t
Xbit_r106_c133 bl[133] br[133] wl[106] vdd gnd cell_6t
Xbit_r107_c133 bl[133] br[133] wl[107] vdd gnd cell_6t
Xbit_r108_c133 bl[133] br[133] wl[108] vdd gnd cell_6t
Xbit_r109_c133 bl[133] br[133] wl[109] vdd gnd cell_6t
Xbit_r110_c133 bl[133] br[133] wl[110] vdd gnd cell_6t
Xbit_r111_c133 bl[133] br[133] wl[111] vdd gnd cell_6t
Xbit_r112_c133 bl[133] br[133] wl[112] vdd gnd cell_6t
Xbit_r113_c133 bl[133] br[133] wl[113] vdd gnd cell_6t
Xbit_r114_c133 bl[133] br[133] wl[114] vdd gnd cell_6t
Xbit_r115_c133 bl[133] br[133] wl[115] vdd gnd cell_6t
Xbit_r116_c133 bl[133] br[133] wl[116] vdd gnd cell_6t
Xbit_r117_c133 bl[133] br[133] wl[117] vdd gnd cell_6t
Xbit_r118_c133 bl[133] br[133] wl[118] vdd gnd cell_6t
Xbit_r119_c133 bl[133] br[133] wl[119] vdd gnd cell_6t
Xbit_r120_c133 bl[133] br[133] wl[120] vdd gnd cell_6t
Xbit_r121_c133 bl[133] br[133] wl[121] vdd gnd cell_6t
Xbit_r122_c133 bl[133] br[133] wl[122] vdd gnd cell_6t
Xbit_r123_c133 bl[133] br[133] wl[123] vdd gnd cell_6t
Xbit_r124_c133 bl[133] br[133] wl[124] vdd gnd cell_6t
Xbit_r125_c133 bl[133] br[133] wl[125] vdd gnd cell_6t
Xbit_r126_c133 bl[133] br[133] wl[126] vdd gnd cell_6t
Xbit_r127_c133 bl[133] br[133] wl[127] vdd gnd cell_6t
Xbit_r128_c133 bl[133] br[133] wl[128] vdd gnd cell_6t
Xbit_r129_c133 bl[133] br[133] wl[129] vdd gnd cell_6t
Xbit_r130_c133 bl[133] br[133] wl[130] vdd gnd cell_6t
Xbit_r131_c133 bl[133] br[133] wl[131] vdd gnd cell_6t
Xbit_r132_c133 bl[133] br[133] wl[132] vdd gnd cell_6t
Xbit_r133_c133 bl[133] br[133] wl[133] vdd gnd cell_6t
Xbit_r134_c133 bl[133] br[133] wl[134] vdd gnd cell_6t
Xbit_r135_c133 bl[133] br[133] wl[135] vdd gnd cell_6t
Xbit_r136_c133 bl[133] br[133] wl[136] vdd gnd cell_6t
Xbit_r137_c133 bl[133] br[133] wl[137] vdd gnd cell_6t
Xbit_r138_c133 bl[133] br[133] wl[138] vdd gnd cell_6t
Xbit_r139_c133 bl[133] br[133] wl[139] vdd gnd cell_6t
Xbit_r140_c133 bl[133] br[133] wl[140] vdd gnd cell_6t
Xbit_r141_c133 bl[133] br[133] wl[141] vdd gnd cell_6t
Xbit_r142_c133 bl[133] br[133] wl[142] vdd gnd cell_6t
Xbit_r143_c133 bl[133] br[133] wl[143] vdd gnd cell_6t
Xbit_r144_c133 bl[133] br[133] wl[144] vdd gnd cell_6t
Xbit_r145_c133 bl[133] br[133] wl[145] vdd gnd cell_6t
Xbit_r146_c133 bl[133] br[133] wl[146] vdd gnd cell_6t
Xbit_r147_c133 bl[133] br[133] wl[147] vdd gnd cell_6t
Xbit_r148_c133 bl[133] br[133] wl[148] vdd gnd cell_6t
Xbit_r149_c133 bl[133] br[133] wl[149] vdd gnd cell_6t
Xbit_r150_c133 bl[133] br[133] wl[150] vdd gnd cell_6t
Xbit_r151_c133 bl[133] br[133] wl[151] vdd gnd cell_6t
Xbit_r152_c133 bl[133] br[133] wl[152] vdd gnd cell_6t
Xbit_r153_c133 bl[133] br[133] wl[153] vdd gnd cell_6t
Xbit_r154_c133 bl[133] br[133] wl[154] vdd gnd cell_6t
Xbit_r155_c133 bl[133] br[133] wl[155] vdd gnd cell_6t
Xbit_r156_c133 bl[133] br[133] wl[156] vdd gnd cell_6t
Xbit_r157_c133 bl[133] br[133] wl[157] vdd gnd cell_6t
Xbit_r158_c133 bl[133] br[133] wl[158] vdd gnd cell_6t
Xbit_r159_c133 bl[133] br[133] wl[159] vdd gnd cell_6t
Xbit_r160_c133 bl[133] br[133] wl[160] vdd gnd cell_6t
Xbit_r161_c133 bl[133] br[133] wl[161] vdd gnd cell_6t
Xbit_r162_c133 bl[133] br[133] wl[162] vdd gnd cell_6t
Xbit_r163_c133 bl[133] br[133] wl[163] vdd gnd cell_6t
Xbit_r164_c133 bl[133] br[133] wl[164] vdd gnd cell_6t
Xbit_r165_c133 bl[133] br[133] wl[165] vdd gnd cell_6t
Xbit_r166_c133 bl[133] br[133] wl[166] vdd gnd cell_6t
Xbit_r167_c133 bl[133] br[133] wl[167] vdd gnd cell_6t
Xbit_r168_c133 bl[133] br[133] wl[168] vdd gnd cell_6t
Xbit_r169_c133 bl[133] br[133] wl[169] vdd gnd cell_6t
Xbit_r170_c133 bl[133] br[133] wl[170] vdd gnd cell_6t
Xbit_r171_c133 bl[133] br[133] wl[171] vdd gnd cell_6t
Xbit_r172_c133 bl[133] br[133] wl[172] vdd gnd cell_6t
Xbit_r173_c133 bl[133] br[133] wl[173] vdd gnd cell_6t
Xbit_r174_c133 bl[133] br[133] wl[174] vdd gnd cell_6t
Xbit_r175_c133 bl[133] br[133] wl[175] vdd gnd cell_6t
Xbit_r176_c133 bl[133] br[133] wl[176] vdd gnd cell_6t
Xbit_r177_c133 bl[133] br[133] wl[177] vdd gnd cell_6t
Xbit_r178_c133 bl[133] br[133] wl[178] vdd gnd cell_6t
Xbit_r179_c133 bl[133] br[133] wl[179] vdd gnd cell_6t
Xbit_r180_c133 bl[133] br[133] wl[180] vdd gnd cell_6t
Xbit_r181_c133 bl[133] br[133] wl[181] vdd gnd cell_6t
Xbit_r182_c133 bl[133] br[133] wl[182] vdd gnd cell_6t
Xbit_r183_c133 bl[133] br[133] wl[183] vdd gnd cell_6t
Xbit_r184_c133 bl[133] br[133] wl[184] vdd gnd cell_6t
Xbit_r185_c133 bl[133] br[133] wl[185] vdd gnd cell_6t
Xbit_r186_c133 bl[133] br[133] wl[186] vdd gnd cell_6t
Xbit_r187_c133 bl[133] br[133] wl[187] vdd gnd cell_6t
Xbit_r188_c133 bl[133] br[133] wl[188] vdd gnd cell_6t
Xbit_r189_c133 bl[133] br[133] wl[189] vdd gnd cell_6t
Xbit_r190_c133 bl[133] br[133] wl[190] vdd gnd cell_6t
Xbit_r191_c133 bl[133] br[133] wl[191] vdd gnd cell_6t
Xbit_r192_c133 bl[133] br[133] wl[192] vdd gnd cell_6t
Xbit_r193_c133 bl[133] br[133] wl[193] vdd gnd cell_6t
Xbit_r194_c133 bl[133] br[133] wl[194] vdd gnd cell_6t
Xbit_r195_c133 bl[133] br[133] wl[195] vdd gnd cell_6t
Xbit_r196_c133 bl[133] br[133] wl[196] vdd gnd cell_6t
Xbit_r197_c133 bl[133] br[133] wl[197] vdd gnd cell_6t
Xbit_r198_c133 bl[133] br[133] wl[198] vdd gnd cell_6t
Xbit_r199_c133 bl[133] br[133] wl[199] vdd gnd cell_6t
Xbit_r200_c133 bl[133] br[133] wl[200] vdd gnd cell_6t
Xbit_r201_c133 bl[133] br[133] wl[201] vdd gnd cell_6t
Xbit_r202_c133 bl[133] br[133] wl[202] vdd gnd cell_6t
Xbit_r203_c133 bl[133] br[133] wl[203] vdd gnd cell_6t
Xbit_r204_c133 bl[133] br[133] wl[204] vdd gnd cell_6t
Xbit_r205_c133 bl[133] br[133] wl[205] vdd gnd cell_6t
Xbit_r206_c133 bl[133] br[133] wl[206] vdd gnd cell_6t
Xbit_r207_c133 bl[133] br[133] wl[207] vdd gnd cell_6t
Xbit_r208_c133 bl[133] br[133] wl[208] vdd gnd cell_6t
Xbit_r209_c133 bl[133] br[133] wl[209] vdd gnd cell_6t
Xbit_r210_c133 bl[133] br[133] wl[210] vdd gnd cell_6t
Xbit_r211_c133 bl[133] br[133] wl[211] vdd gnd cell_6t
Xbit_r212_c133 bl[133] br[133] wl[212] vdd gnd cell_6t
Xbit_r213_c133 bl[133] br[133] wl[213] vdd gnd cell_6t
Xbit_r214_c133 bl[133] br[133] wl[214] vdd gnd cell_6t
Xbit_r215_c133 bl[133] br[133] wl[215] vdd gnd cell_6t
Xbit_r216_c133 bl[133] br[133] wl[216] vdd gnd cell_6t
Xbit_r217_c133 bl[133] br[133] wl[217] vdd gnd cell_6t
Xbit_r218_c133 bl[133] br[133] wl[218] vdd gnd cell_6t
Xbit_r219_c133 bl[133] br[133] wl[219] vdd gnd cell_6t
Xbit_r220_c133 bl[133] br[133] wl[220] vdd gnd cell_6t
Xbit_r221_c133 bl[133] br[133] wl[221] vdd gnd cell_6t
Xbit_r222_c133 bl[133] br[133] wl[222] vdd gnd cell_6t
Xbit_r223_c133 bl[133] br[133] wl[223] vdd gnd cell_6t
Xbit_r224_c133 bl[133] br[133] wl[224] vdd gnd cell_6t
Xbit_r225_c133 bl[133] br[133] wl[225] vdd gnd cell_6t
Xbit_r226_c133 bl[133] br[133] wl[226] vdd gnd cell_6t
Xbit_r227_c133 bl[133] br[133] wl[227] vdd gnd cell_6t
Xbit_r228_c133 bl[133] br[133] wl[228] vdd gnd cell_6t
Xbit_r229_c133 bl[133] br[133] wl[229] vdd gnd cell_6t
Xbit_r230_c133 bl[133] br[133] wl[230] vdd gnd cell_6t
Xbit_r231_c133 bl[133] br[133] wl[231] vdd gnd cell_6t
Xbit_r232_c133 bl[133] br[133] wl[232] vdd gnd cell_6t
Xbit_r233_c133 bl[133] br[133] wl[233] vdd gnd cell_6t
Xbit_r234_c133 bl[133] br[133] wl[234] vdd gnd cell_6t
Xbit_r235_c133 bl[133] br[133] wl[235] vdd gnd cell_6t
Xbit_r236_c133 bl[133] br[133] wl[236] vdd gnd cell_6t
Xbit_r237_c133 bl[133] br[133] wl[237] vdd gnd cell_6t
Xbit_r238_c133 bl[133] br[133] wl[238] vdd gnd cell_6t
Xbit_r239_c133 bl[133] br[133] wl[239] vdd gnd cell_6t
Xbit_r240_c133 bl[133] br[133] wl[240] vdd gnd cell_6t
Xbit_r241_c133 bl[133] br[133] wl[241] vdd gnd cell_6t
Xbit_r242_c133 bl[133] br[133] wl[242] vdd gnd cell_6t
Xbit_r243_c133 bl[133] br[133] wl[243] vdd gnd cell_6t
Xbit_r244_c133 bl[133] br[133] wl[244] vdd gnd cell_6t
Xbit_r245_c133 bl[133] br[133] wl[245] vdd gnd cell_6t
Xbit_r246_c133 bl[133] br[133] wl[246] vdd gnd cell_6t
Xbit_r247_c133 bl[133] br[133] wl[247] vdd gnd cell_6t
Xbit_r248_c133 bl[133] br[133] wl[248] vdd gnd cell_6t
Xbit_r249_c133 bl[133] br[133] wl[249] vdd gnd cell_6t
Xbit_r250_c133 bl[133] br[133] wl[250] vdd gnd cell_6t
Xbit_r251_c133 bl[133] br[133] wl[251] vdd gnd cell_6t
Xbit_r252_c133 bl[133] br[133] wl[252] vdd gnd cell_6t
Xbit_r253_c133 bl[133] br[133] wl[253] vdd gnd cell_6t
Xbit_r254_c133 bl[133] br[133] wl[254] vdd gnd cell_6t
Xbit_r255_c133 bl[133] br[133] wl[255] vdd gnd cell_6t
Xbit_r0_c134 bl[134] br[134] wl[0] vdd gnd cell_6t
Xbit_r1_c134 bl[134] br[134] wl[1] vdd gnd cell_6t
Xbit_r2_c134 bl[134] br[134] wl[2] vdd gnd cell_6t
Xbit_r3_c134 bl[134] br[134] wl[3] vdd gnd cell_6t
Xbit_r4_c134 bl[134] br[134] wl[4] vdd gnd cell_6t
Xbit_r5_c134 bl[134] br[134] wl[5] vdd gnd cell_6t
Xbit_r6_c134 bl[134] br[134] wl[6] vdd gnd cell_6t
Xbit_r7_c134 bl[134] br[134] wl[7] vdd gnd cell_6t
Xbit_r8_c134 bl[134] br[134] wl[8] vdd gnd cell_6t
Xbit_r9_c134 bl[134] br[134] wl[9] vdd gnd cell_6t
Xbit_r10_c134 bl[134] br[134] wl[10] vdd gnd cell_6t
Xbit_r11_c134 bl[134] br[134] wl[11] vdd gnd cell_6t
Xbit_r12_c134 bl[134] br[134] wl[12] vdd gnd cell_6t
Xbit_r13_c134 bl[134] br[134] wl[13] vdd gnd cell_6t
Xbit_r14_c134 bl[134] br[134] wl[14] vdd gnd cell_6t
Xbit_r15_c134 bl[134] br[134] wl[15] vdd gnd cell_6t
Xbit_r16_c134 bl[134] br[134] wl[16] vdd gnd cell_6t
Xbit_r17_c134 bl[134] br[134] wl[17] vdd gnd cell_6t
Xbit_r18_c134 bl[134] br[134] wl[18] vdd gnd cell_6t
Xbit_r19_c134 bl[134] br[134] wl[19] vdd gnd cell_6t
Xbit_r20_c134 bl[134] br[134] wl[20] vdd gnd cell_6t
Xbit_r21_c134 bl[134] br[134] wl[21] vdd gnd cell_6t
Xbit_r22_c134 bl[134] br[134] wl[22] vdd gnd cell_6t
Xbit_r23_c134 bl[134] br[134] wl[23] vdd gnd cell_6t
Xbit_r24_c134 bl[134] br[134] wl[24] vdd gnd cell_6t
Xbit_r25_c134 bl[134] br[134] wl[25] vdd gnd cell_6t
Xbit_r26_c134 bl[134] br[134] wl[26] vdd gnd cell_6t
Xbit_r27_c134 bl[134] br[134] wl[27] vdd gnd cell_6t
Xbit_r28_c134 bl[134] br[134] wl[28] vdd gnd cell_6t
Xbit_r29_c134 bl[134] br[134] wl[29] vdd gnd cell_6t
Xbit_r30_c134 bl[134] br[134] wl[30] vdd gnd cell_6t
Xbit_r31_c134 bl[134] br[134] wl[31] vdd gnd cell_6t
Xbit_r32_c134 bl[134] br[134] wl[32] vdd gnd cell_6t
Xbit_r33_c134 bl[134] br[134] wl[33] vdd gnd cell_6t
Xbit_r34_c134 bl[134] br[134] wl[34] vdd gnd cell_6t
Xbit_r35_c134 bl[134] br[134] wl[35] vdd gnd cell_6t
Xbit_r36_c134 bl[134] br[134] wl[36] vdd gnd cell_6t
Xbit_r37_c134 bl[134] br[134] wl[37] vdd gnd cell_6t
Xbit_r38_c134 bl[134] br[134] wl[38] vdd gnd cell_6t
Xbit_r39_c134 bl[134] br[134] wl[39] vdd gnd cell_6t
Xbit_r40_c134 bl[134] br[134] wl[40] vdd gnd cell_6t
Xbit_r41_c134 bl[134] br[134] wl[41] vdd gnd cell_6t
Xbit_r42_c134 bl[134] br[134] wl[42] vdd gnd cell_6t
Xbit_r43_c134 bl[134] br[134] wl[43] vdd gnd cell_6t
Xbit_r44_c134 bl[134] br[134] wl[44] vdd gnd cell_6t
Xbit_r45_c134 bl[134] br[134] wl[45] vdd gnd cell_6t
Xbit_r46_c134 bl[134] br[134] wl[46] vdd gnd cell_6t
Xbit_r47_c134 bl[134] br[134] wl[47] vdd gnd cell_6t
Xbit_r48_c134 bl[134] br[134] wl[48] vdd gnd cell_6t
Xbit_r49_c134 bl[134] br[134] wl[49] vdd gnd cell_6t
Xbit_r50_c134 bl[134] br[134] wl[50] vdd gnd cell_6t
Xbit_r51_c134 bl[134] br[134] wl[51] vdd gnd cell_6t
Xbit_r52_c134 bl[134] br[134] wl[52] vdd gnd cell_6t
Xbit_r53_c134 bl[134] br[134] wl[53] vdd gnd cell_6t
Xbit_r54_c134 bl[134] br[134] wl[54] vdd gnd cell_6t
Xbit_r55_c134 bl[134] br[134] wl[55] vdd gnd cell_6t
Xbit_r56_c134 bl[134] br[134] wl[56] vdd gnd cell_6t
Xbit_r57_c134 bl[134] br[134] wl[57] vdd gnd cell_6t
Xbit_r58_c134 bl[134] br[134] wl[58] vdd gnd cell_6t
Xbit_r59_c134 bl[134] br[134] wl[59] vdd gnd cell_6t
Xbit_r60_c134 bl[134] br[134] wl[60] vdd gnd cell_6t
Xbit_r61_c134 bl[134] br[134] wl[61] vdd gnd cell_6t
Xbit_r62_c134 bl[134] br[134] wl[62] vdd gnd cell_6t
Xbit_r63_c134 bl[134] br[134] wl[63] vdd gnd cell_6t
Xbit_r64_c134 bl[134] br[134] wl[64] vdd gnd cell_6t
Xbit_r65_c134 bl[134] br[134] wl[65] vdd gnd cell_6t
Xbit_r66_c134 bl[134] br[134] wl[66] vdd gnd cell_6t
Xbit_r67_c134 bl[134] br[134] wl[67] vdd gnd cell_6t
Xbit_r68_c134 bl[134] br[134] wl[68] vdd gnd cell_6t
Xbit_r69_c134 bl[134] br[134] wl[69] vdd gnd cell_6t
Xbit_r70_c134 bl[134] br[134] wl[70] vdd gnd cell_6t
Xbit_r71_c134 bl[134] br[134] wl[71] vdd gnd cell_6t
Xbit_r72_c134 bl[134] br[134] wl[72] vdd gnd cell_6t
Xbit_r73_c134 bl[134] br[134] wl[73] vdd gnd cell_6t
Xbit_r74_c134 bl[134] br[134] wl[74] vdd gnd cell_6t
Xbit_r75_c134 bl[134] br[134] wl[75] vdd gnd cell_6t
Xbit_r76_c134 bl[134] br[134] wl[76] vdd gnd cell_6t
Xbit_r77_c134 bl[134] br[134] wl[77] vdd gnd cell_6t
Xbit_r78_c134 bl[134] br[134] wl[78] vdd gnd cell_6t
Xbit_r79_c134 bl[134] br[134] wl[79] vdd gnd cell_6t
Xbit_r80_c134 bl[134] br[134] wl[80] vdd gnd cell_6t
Xbit_r81_c134 bl[134] br[134] wl[81] vdd gnd cell_6t
Xbit_r82_c134 bl[134] br[134] wl[82] vdd gnd cell_6t
Xbit_r83_c134 bl[134] br[134] wl[83] vdd gnd cell_6t
Xbit_r84_c134 bl[134] br[134] wl[84] vdd gnd cell_6t
Xbit_r85_c134 bl[134] br[134] wl[85] vdd gnd cell_6t
Xbit_r86_c134 bl[134] br[134] wl[86] vdd gnd cell_6t
Xbit_r87_c134 bl[134] br[134] wl[87] vdd gnd cell_6t
Xbit_r88_c134 bl[134] br[134] wl[88] vdd gnd cell_6t
Xbit_r89_c134 bl[134] br[134] wl[89] vdd gnd cell_6t
Xbit_r90_c134 bl[134] br[134] wl[90] vdd gnd cell_6t
Xbit_r91_c134 bl[134] br[134] wl[91] vdd gnd cell_6t
Xbit_r92_c134 bl[134] br[134] wl[92] vdd gnd cell_6t
Xbit_r93_c134 bl[134] br[134] wl[93] vdd gnd cell_6t
Xbit_r94_c134 bl[134] br[134] wl[94] vdd gnd cell_6t
Xbit_r95_c134 bl[134] br[134] wl[95] vdd gnd cell_6t
Xbit_r96_c134 bl[134] br[134] wl[96] vdd gnd cell_6t
Xbit_r97_c134 bl[134] br[134] wl[97] vdd gnd cell_6t
Xbit_r98_c134 bl[134] br[134] wl[98] vdd gnd cell_6t
Xbit_r99_c134 bl[134] br[134] wl[99] vdd gnd cell_6t
Xbit_r100_c134 bl[134] br[134] wl[100] vdd gnd cell_6t
Xbit_r101_c134 bl[134] br[134] wl[101] vdd gnd cell_6t
Xbit_r102_c134 bl[134] br[134] wl[102] vdd gnd cell_6t
Xbit_r103_c134 bl[134] br[134] wl[103] vdd gnd cell_6t
Xbit_r104_c134 bl[134] br[134] wl[104] vdd gnd cell_6t
Xbit_r105_c134 bl[134] br[134] wl[105] vdd gnd cell_6t
Xbit_r106_c134 bl[134] br[134] wl[106] vdd gnd cell_6t
Xbit_r107_c134 bl[134] br[134] wl[107] vdd gnd cell_6t
Xbit_r108_c134 bl[134] br[134] wl[108] vdd gnd cell_6t
Xbit_r109_c134 bl[134] br[134] wl[109] vdd gnd cell_6t
Xbit_r110_c134 bl[134] br[134] wl[110] vdd gnd cell_6t
Xbit_r111_c134 bl[134] br[134] wl[111] vdd gnd cell_6t
Xbit_r112_c134 bl[134] br[134] wl[112] vdd gnd cell_6t
Xbit_r113_c134 bl[134] br[134] wl[113] vdd gnd cell_6t
Xbit_r114_c134 bl[134] br[134] wl[114] vdd gnd cell_6t
Xbit_r115_c134 bl[134] br[134] wl[115] vdd gnd cell_6t
Xbit_r116_c134 bl[134] br[134] wl[116] vdd gnd cell_6t
Xbit_r117_c134 bl[134] br[134] wl[117] vdd gnd cell_6t
Xbit_r118_c134 bl[134] br[134] wl[118] vdd gnd cell_6t
Xbit_r119_c134 bl[134] br[134] wl[119] vdd gnd cell_6t
Xbit_r120_c134 bl[134] br[134] wl[120] vdd gnd cell_6t
Xbit_r121_c134 bl[134] br[134] wl[121] vdd gnd cell_6t
Xbit_r122_c134 bl[134] br[134] wl[122] vdd gnd cell_6t
Xbit_r123_c134 bl[134] br[134] wl[123] vdd gnd cell_6t
Xbit_r124_c134 bl[134] br[134] wl[124] vdd gnd cell_6t
Xbit_r125_c134 bl[134] br[134] wl[125] vdd gnd cell_6t
Xbit_r126_c134 bl[134] br[134] wl[126] vdd gnd cell_6t
Xbit_r127_c134 bl[134] br[134] wl[127] vdd gnd cell_6t
Xbit_r128_c134 bl[134] br[134] wl[128] vdd gnd cell_6t
Xbit_r129_c134 bl[134] br[134] wl[129] vdd gnd cell_6t
Xbit_r130_c134 bl[134] br[134] wl[130] vdd gnd cell_6t
Xbit_r131_c134 bl[134] br[134] wl[131] vdd gnd cell_6t
Xbit_r132_c134 bl[134] br[134] wl[132] vdd gnd cell_6t
Xbit_r133_c134 bl[134] br[134] wl[133] vdd gnd cell_6t
Xbit_r134_c134 bl[134] br[134] wl[134] vdd gnd cell_6t
Xbit_r135_c134 bl[134] br[134] wl[135] vdd gnd cell_6t
Xbit_r136_c134 bl[134] br[134] wl[136] vdd gnd cell_6t
Xbit_r137_c134 bl[134] br[134] wl[137] vdd gnd cell_6t
Xbit_r138_c134 bl[134] br[134] wl[138] vdd gnd cell_6t
Xbit_r139_c134 bl[134] br[134] wl[139] vdd gnd cell_6t
Xbit_r140_c134 bl[134] br[134] wl[140] vdd gnd cell_6t
Xbit_r141_c134 bl[134] br[134] wl[141] vdd gnd cell_6t
Xbit_r142_c134 bl[134] br[134] wl[142] vdd gnd cell_6t
Xbit_r143_c134 bl[134] br[134] wl[143] vdd gnd cell_6t
Xbit_r144_c134 bl[134] br[134] wl[144] vdd gnd cell_6t
Xbit_r145_c134 bl[134] br[134] wl[145] vdd gnd cell_6t
Xbit_r146_c134 bl[134] br[134] wl[146] vdd gnd cell_6t
Xbit_r147_c134 bl[134] br[134] wl[147] vdd gnd cell_6t
Xbit_r148_c134 bl[134] br[134] wl[148] vdd gnd cell_6t
Xbit_r149_c134 bl[134] br[134] wl[149] vdd gnd cell_6t
Xbit_r150_c134 bl[134] br[134] wl[150] vdd gnd cell_6t
Xbit_r151_c134 bl[134] br[134] wl[151] vdd gnd cell_6t
Xbit_r152_c134 bl[134] br[134] wl[152] vdd gnd cell_6t
Xbit_r153_c134 bl[134] br[134] wl[153] vdd gnd cell_6t
Xbit_r154_c134 bl[134] br[134] wl[154] vdd gnd cell_6t
Xbit_r155_c134 bl[134] br[134] wl[155] vdd gnd cell_6t
Xbit_r156_c134 bl[134] br[134] wl[156] vdd gnd cell_6t
Xbit_r157_c134 bl[134] br[134] wl[157] vdd gnd cell_6t
Xbit_r158_c134 bl[134] br[134] wl[158] vdd gnd cell_6t
Xbit_r159_c134 bl[134] br[134] wl[159] vdd gnd cell_6t
Xbit_r160_c134 bl[134] br[134] wl[160] vdd gnd cell_6t
Xbit_r161_c134 bl[134] br[134] wl[161] vdd gnd cell_6t
Xbit_r162_c134 bl[134] br[134] wl[162] vdd gnd cell_6t
Xbit_r163_c134 bl[134] br[134] wl[163] vdd gnd cell_6t
Xbit_r164_c134 bl[134] br[134] wl[164] vdd gnd cell_6t
Xbit_r165_c134 bl[134] br[134] wl[165] vdd gnd cell_6t
Xbit_r166_c134 bl[134] br[134] wl[166] vdd gnd cell_6t
Xbit_r167_c134 bl[134] br[134] wl[167] vdd gnd cell_6t
Xbit_r168_c134 bl[134] br[134] wl[168] vdd gnd cell_6t
Xbit_r169_c134 bl[134] br[134] wl[169] vdd gnd cell_6t
Xbit_r170_c134 bl[134] br[134] wl[170] vdd gnd cell_6t
Xbit_r171_c134 bl[134] br[134] wl[171] vdd gnd cell_6t
Xbit_r172_c134 bl[134] br[134] wl[172] vdd gnd cell_6t
Xbit_r173_c134 bl[134] br[134] wl[173] vdd gnd cell_6t
Xbit_r174_c134 bl[134] br[134] wl[174] vdd gnd cell_6t
Xbit_r175_c134 bl[134] br[134] wl[175] vdd gnd cell_6t
Xbit_r176_c134 bl[134] br[134] wl[176] vdd gnd cell_6t
Xbit_r177_c134 bl[134] br[134] wl[177] vdd gnd cell_6t
Xbit_r178_c134 bl[134] br[134] wl[178] vdd gnd cell_6t
Xbit_r179_c134 bl[134] br[134] wl[179] vdd gnd cell_6t
Xbit_r180_c134 bl[134] br[134] wl[180] vdd gnd cell_6t
Xbit_r181_c134 bl[134] br[134] wl[181] vdd gnd cell_6t
Xbit_r182_c134 bl[134] br[134] wl[182] vdd gnd cell_6t
Xbit_r183_c134 bl[134] br[134] wl[183] vdd gnd cell_6t
Xbit_r184_c134 bl[134] br[134] wl[184] vdd gnd cell_6t
Xbit_r185_c134 bl[134] br[134] wl[185] vdd gnd cell_6t
Xbit_r186_c134 bl[134] br[134] wl[186] vdd gnd cell_6t
Xbit_r187_c134 bl[134] br[134] wl[187] vdd gnd cell_6t
Xbit_r188_c134 bl[134] br[134] wl[188] vdd gnd cell_6t
Xbit_r189_c134 bl[134] br[134] wl[189] vdd gnd cell_6t
Xbit_r190_c134 bl[134] br[134] wl[190] vdd gnd cell_6t
Xbit_r191_c134 bl[134] br[134] wl[191] vdd gnd cell_6t
Xbit_r192_c134 bl[134] br[134] wl[192] vdd gnd cell_6t
Xbit_r193_c134 bl[134] br[134] wl[193] vdd gnd cell_6t
Xbit_r194_c134 bl[134] br[134] wl[194] vdd gnd cell_6t
Xbit_r195_c134 bl[134] br[134] wl[195] vdd gnd cell_6t
Xbit_r196_c134 bl[134] br[134] wl[196] vdd gnd cell_6t
Xbit_r197_c134 bl[134] br[134] wl[197] vdd gnd cell_6t
Xbit_r198_c134 bl[134] br[134] wl[198] vdd gnd cell_6t
Xbit_r199_c134 bl[134] br[134] wl[199] vdd gnd cell_6t
Xbit_r200_c134 bl[134] br[134] wl[200] vdd gnd cell_6t
Xbit_r201_c134 bl[134] br[134] wl[201] vdd gnd cell_6t
Xbit_r202_c134 bl[134] br[134] wl[202] vdd gnd cell_6t
Xbit_r203_c134 bl[134] br[134] wl[203] vdd gnd cell_6t
Xbit_r204_c134 bl[134] br[134] wl[204] vdd gnd cell_6t
Xbit_r205_c134 bl[134] br[134] wl[205] vdd gnd cell_6t
Xbit_r206_c134 bl[134] br[134] wl[206] vdd gnd cell_6t
Xbit_r207_c134 bl[134] br[134] wl[207] vdd gnd cell_6t
Xbit_r208_c134 bl[134] br[134] wl[208] vdd gnd cell_6t
Xbit_r209_c134 bl[134] br[134] wl[209] vdd gnd cell_6t
Xbit_r210_c134 bl[134] br[134] wl[210] vdd gnd cell_6t
Xbit_r211_c134 bl[134] br[134] wl[211] vdd gnd cell_6t
Xbit_r212_c134 bl[134] br[134] wl[212] vdd gnd cell_6t
Xbit_r213_c134 bl[134] br[134] wl[213] vdd gnd cell_6t
Xbit_r214_c134 bl[134] br[134] wl[214] vdd gnd cell_6t
Xbit_r215_c134 bl[134] br[134] wl[215] vdd gnd cell_6t
Xbit_r216_c134 bl[134] br[134] wl[216] vdd gnd cell_6t
Xbit_r217_c134 bl[134] br[134] wl[217] vdd gnd cell_6t
Xbit_r218_c134 bl[134] br[134] wl[218] vdd gnd cell_6t
Xbit_r219_c134 bl[134] br[134] wl[219] vdd gnd cell_6t
Xbit_r220_c134 bl[134] br[134] wl[220] vdd gnd cell_6t
Xbit_r221_c134 bl[134] br[134] wl[221] vdd gnd cell_6t
Xbit_r222_c134 bl[134] br[134] wl[222] vdd gnd cell_6t
Xbit_r223_c134 bl[134] br[134] wl[223] vdd gnd cell_6t
Xbit_r224_c134 bl[134] br[134] wl[224] vdd gnd cell_6t
Xbit_r225_c134 bl[134] br[134] wl[225] vdd gnd cell_6t
Xbit_r226_c134 bl[134] br[134] wl[226] vdd gnd cell_6t
Xbit_r227_c134 bl[134] br[134] wl[227] vdd gnd cell_6t
Xbit_r228_c134 bl[134] br[134] wl[228] vdd gnd cell_6t
Xbit_r229_c134 bl[134] br[134] wl[229] vdd gnd cell_6t
Xbit_r230_c134 bl[134] br[134] wl[230] vdd gnd cell_6t
Xbit_r231_c134 bl[134] br[134] wl[231] vdd gnd cell_6t
Xbit_r232_c134 bl[134] br[134] wl[232] vdd gnd cell_6t
Xbit_r233_c134 bl[134] br[134] wl[233] vdd gnd cell_6t
Xbit_r234_c134 bl[134] br[134] wl[234] vdd gnd cell_6t
Xbit_r235_c134 bl[134] br[134] wl[235] vdd gnd cell_6t
Xbit_r236_c134 bl[134] br[134] wl[236] vdd gnd cell_6t
Xbit_r237_c134 bl[134] br[134] wl[237] vdd gnd cell_6t
Xbit_r238_c134 bl[134] br[134] wl[238] vdd gnd cell_6t
Xbit_r239_c134 bl[134] br[134] wl[239] vdd gnd cell_6t
Xbit_r240_c134 bl[134] br[134] wl[240] vdd gnd cell_6t
Xbit_r241_c134 bl[134] br[134] wl[241] vdd gnd cell_6t
Xbit_r242_c134 bl[134] br[134] wl[242] vdd gnd cell_6t
Xbit_r243_c134 bl[134] br[134] wl[243] vdd gnd cell_6t
Xbit_r244_c134 bl[134] br[134] wl[244] vdd gnd cell_6t
Xbit_r245_c134 bl[134] br[134] wl[245] vdd gnd cell_6t
Xbit_r246_c134 bl[134] br[134] wl[246] vdd gnd cell_6t
Xbit_r247_c134 bl[134] br[134] wl[247] vdd gnd cell_6t
Xbit_r248_c134 bl[134] br[134] wl[248] vdd gnd cell_6t
Xbit_r249_c134 bl[134] br[134] wl[249] vdd gnd cell_6t
Xbit_r250_c134 bl[134] br[134] wl[250] vdd gnd cell_6t
Xbit_r251_c134 bl[134] br[134] wl[251] vdd gnd cell_6t
Xbit_r252_c134 bl[134] br[134] wl[252] vdd gnd cell_6t
Xbit_r253_c134 bl[134] br[134] wl[253] vdd gnd cell_6t
Xbit_r254_c134 bl[134] br[134] wl[254] vdd gnd cell_6t
Xbit_r255_c134 bl[134] br[134] wl[255] vdd gnd cell_6t
Xbit_r0_c135 bl[135] br[135] wl[0] vdd gnd cell_6t
Xbit_r1_c135 bl[135] br[135] wl[1] vdd gnd cell_6t
Xbit_r2_c135 bl[135] br[135] wl[2] vdd gnd cell_6t
Xbit_r3_c135 bl[135] br[135] wl[3] vdd gnd cell_6t
Xbit_r4_c135 bl[135] br[135] wl[4] vdd gnd cell_6t
Xbit_r5_c135 bl[135] br[135] wl[5] vdd gnd cell_6t
Xbit_r6_c135 bl[135] br[135] wl[6] vdd gnd cell_6t
Xbit_r7_c135 bl[135] br[135] wl[7] vdd gnd cell_6t
Xbit_r8_c135 bl[135] br[135] wl[8] vdd gnd cell_6t
Xbit_r9_c135 bl[135] br[135] wl[9] vdd gnd cell_6t
Xbit_r10_c135 bl[135] br[135] wl[10] vdd gnd cell_6t
Xbit_r11_c135 bl[135] br[135] wl[11] vdd gnd cell_6t
Xbit_r12_c135 bl[135] br[135] wl[12] vdd gnd cell_6t
Xbit_r13_c135 bl[135] br[135] wl[13] vdd gnd cell_6t
Xbit_r14_c135 bl[135] br[135] wl[14] vdd gnd cell_6t
Xbit_r15_c135 bl[135] br[135] wl[15] vdd gnd cell_6t
Xbit_r16_c135 bl[135] br[135] wl[16] vdd gnd cell_6t
Xbit_r17_c135 bl[135] br[135] wl[17] vdd gnd cell_6t
Xbit_r18_c135 bl[135] br[135] wl[18] vdd gnd cell_6t
Xbit_r19_c135 bl[135] br[135] wl[19] vdd gnd cell_6t
Xbit_r20_c135 bl[135] br[135] wl[20] vdd gnd cell_6t
Xbit_r21_c135 bl[135] br[135] wl[21] vdd gnd cell_6t
Xbit_r22_c135 bl[135] br[135] wl[22] vdd gnd cell_6t
Xbit_r23_c135 bl[135] br[135] wl[23] vdd gnd cell_6t
Xbit_r24_c135 bl[135] br[135] wl[24] vdd gnd cell_6t
Xbit_r25_c135 bl[135] br[135] wl[25] vdd gnd cell_6t
Xbit_r26_c135 bl[135] br[135] wl[26] vdd gnd cell_6t
Xbit_r27_c135 bl[135] br[135] wl[27] vdd gnd cell_6t
Xbit_r28_c135 bl[135] br[135] wl[28] vdd gnd cell_6t
Xbit_r29_c135 bl[135] br[135] wl[29] vdd gnd cell_6t
Xbit_r30_c135 bl[135] br[135] wl[30] vdd gnd cell_6t
Xbit_r31_c135 bl[135] br[135] wl[31] vdd gnd cell_6t
Xbit_r32_c135 bl[135] br[135] wl[32] vdd gnd cell_6t
Xbit_r33_c135 bl[135] br[135] wl[33] vdd gnd cell_6t
Xbit_r34_c135 bl[135] br[135] wl[34] vdd gnd cell_6t
Xbit_r35_c135 bl[135] br[135] wl[35] vdd gnd cell_6t
Xbit_r36_c135 bl[135] br[135] wl[36] vdd gnd cell_6t
Xbit_r37_c135 bl[135] br[135] wl[37] vdd gnd cell_6t
Xbit_r38_c135 bl[135] br[135] wl[38] vdd gnd cell_6t
Xbit_r39_c135 bl[135] br[135] wl[39] vdd gnd cell_6t
Xbit_r40_c135 bl[135] br[135] wl[40] vdd gnd cell_6t
Xbit_r41_c135 bl[135] br[135] wl[41] vdd gnd cell_6t
Xbit_r42_c135 bl[135] br[135] wl[42] vdd gnd cell_6t
Xbit_r43_c135 bl[135] br[135] wl[43] vdd gnd cell_6t
Xbit_r44_c135 bl[135] br[135] wl[44] vdd gnd cell_6t
Xbit_r45_c135 bl[135] br[135] wl[45] vdd gnd cell_6t
Xbit_r46_c135 bl[135] br[135] wl[46] vdd gnd cell_6t
Xbit_r47_c135 bl[135] br[135] wl[47] vdd gnd cell_6t
Xbit_r48_c135 bl[135] br[135] wl[48] vdd gnd cell_6t
Xbit_r49_c135 bl[135] br[135] wl[49] vdd gnd cell_6t
Xbit_r50_c135 bl[135] br[135] wl[50] vdd gnd cell_6t
Xbit_r51_c135 bl[135] br[135] wl[51] vdd gnd cell_6t
Xbit_r52_c135 bl[135] br[135] wl[52] vdd gnd cell_6t
Xbit_r53_c135 bl[135] br[135] wl[53] vdd gnd cell_6t
Xbit_r54_c135 bl[135] br[135] wl[54] vdd gnd cell_6t
Xbit_r55_c135 bl[135] br[135] wl[55] vdd gnd cell_6t
Xbit_r56_c135 bl[135] br[135] wl[56] vdd gnd cell_6t
Xbit_r57_c135 bl[135] br[135] wl[57] vdd gnd cell_6t
Xbit_r58_c135 bl[135] br[135] wl[58] vdd gnd cell_6t
Xbit_r59_c135 bl[135] br[135] wl[59] vdd gnd cell_6t
Xbit_r60_c135 bl[135] br[135] wl[60] vdd gnd cell_6t
Xbit_r61_c135 bl[135] br[135] wl[61] vdd gnd cell_6t
Xbit_r62_c135 bl[135] br[135] wl[62] vdd gnd cell_6t
Xbit_r63_c135 bl[135] br[135] wl[63] vdd gnd cell_6t
Xbit_r64_c135 bl[135] br[135] wl[64] vdd gnd cell_6t
Xbit_r65_c135 bl[135] br[135] wl[65] vdd gnd cell_6t
Xbit_r66_c135 bl[135] br[135] wl[66] vdd gnd cell_6t
Xbit_r67_c135 bl[135] br[135] wl[67] vdd gnd cell_6t
Xbit_r68_c135 bl[135] br[135] wl[68] vdd gnd cell_6t
Xbit_r69_c135 bl[135] br[135] wl[69] vdd gnd cell_6t
Xbit_r70_c135 bl[135] br[135] wl[70] vdd gnd cell_6t
Xbit_r71_c135 bl[135] br[135] wl[71] vdd gnd cell_6t
Xbit_r72_c135 bl[135] br[135] wl[72] vdd gnd cell_6t
Xbit_r73_c135 bl[135] br[135] wl[73] vdd gnd cell_6t
Xbit_r74_c135 bl[135] br[135] wl[74] vdd gnd cell_6t
Xbit_r75_c135 bl[135] br[135] wl[75] vdd gnd cell_6t
Xbit_r76_c135 bl[135] br[135] wl[76] vdd gnd cell_6t
Xbit_r77_c135 bl[135] br[135] wl[77] vdd gnd cell_6t
Xbit_r78_c135 bl[135] br[135] wl[78] vdd gnd cell_6t
Xbit_r79_c135 bl[135] br[135] wl[79] vdd gnd cell_6t
Xbit_r80_c135 bl[135] br[135] wl[80] vdd gnd cell_6t
Xbit_r81_c135 bl[135] br[135] wl[81] vdd gnd cell_6t
Xbit_r82_c135 bl[135] br[135] wl[82] vdd gnd cell_6t
Xbit_r83_c135 bl[135] br[135] wl[83] vdd gnd cell_6t
Xbit_r84_c135 bl[135] br[135] wl[84] vdd gnd cell_6t
Xbit_r85_c135 bl[135] br[135] wl[85] vdd gnd cell_6t
Xbit_r86_c135 bl[135] br[135] wl[86] vdd gnd cell_6t
Xbit_r87_c135 bl[135] br[135] wl[87] vdd gnd cell_6t
Xbit_r88_c135 bl[135] br[135] wl[88] vdd gnd cell_6t
Xbit_r89_c135 bl[135] br[135] wl[89] vdd gnd cell_6t
Xbit_r90_c135 bl[135] br[135] wl[90] vdd gnd cell_6t
Xbit_r91_c135 bl[135] br[135] wl[91] vdd gnd cell_6t
Xbit_r92_c135 bl[135] br[135] wl[92] vdd gnd cell_6t
Xbit_r93_c135 bl[135] br[135] wl[93] vdd gnd cell_6t
Xbit_r94_c135 bl[135] br[135] wl[94] vdd gnd cell_6t
Xbit_r95_c135 bl[135] br[135] wl[95] vdd gnd cell_6t
Xbit_r96_c135 bl[135] br[135] wl[96] vdd gnd cell_6t
Xbit_r97_c135 bl[135] br[135] wl[97] vdd gnd cell_6t
Xbit_r98_c135 bl[135] br[135] wl[98] vdd gnd cell_6t
Xbit_r99_c135 bl[135] br[135] wl[99] vdd gnd cell_6t
Xbit_r100_c135 bl[135] br[135] wl[100] vdd gnd cell_6t
Xbit_r101_c135 bl[135] br[135] wl[101] vdd gnd cell_6t
Xbit_r102_c135 bl[135] br[135] wl[102] vdd gnd cell_6t
Xbit_r103_c135 bl[135] br[135] wl[103] vdd gnd cell_6t
Xbit_r104_c135 bl[135] br[135] wl[104] vdd gnd cell_6t
Xbit_r105_c135 bl[135] br[135] wl[105] vdd gnd cell_6t
Xbit_r106_c135 bl[135] br[135] wl[106] vdd gnd cell_6t
Xbit_r107_c135 bl[135] br[135] wl[107] vdd gnd cell_6t
Xbit_r108_c135 bl[135] br[135] wl[108] vdd gnd cell_6t
Xbit_r109_c135 bl[135] br[135] wl[109] vdd gnd cell_6t
Xbit_r110_c135 bl[135] br[135] wl[110] vdd gnd cell_6t
Xbit_r111_c135 bl[135] br[135] wl[111] vdd gnd cell_6t
Xbit_r112_c135 bl[135] br[135] wl[112] vdd gnd cell_6t
Xbit_r113_c135 bl[135] br[135] wl[113] vdd gnd cell_6t
Xbit_r114_c135 bl[135] br[135] wl[114] vdd gnd cell_6t
Xbit_r115_c135 bl[135] br[135] wl[115] vdd gnd cell_6t
Xbit_r116_c135 bl[135] br[135] wl[116] vdd gnd cell_6t
Xbit_r117_c135 bl[135] br[135] wl[117] vdd gnd cell_6t
Xbit_r118_c135 bl[135] br[135] wl[118] vdd gnd cell_6t
Xbit_r119_c135 bl[135] br[135] wl[119] vdd gnd cell_6t
Xbit_r120_c135 bl[135] br[135] wl[120] vdd gnd cell_6t
Xbit_r121_c135 bl[135] br[135] wl[121] vdd gnd cell_6t
Xbit_r122_c135 bl[135] br[135] wl[122] vdd gnd cell_6t
Xbit_r123_c135 bl[135] br[135] wl[123] vdd gnd cell_6t
Xbit_r124_c135 bl[135] br[135] wl[124] vdd gnd cell_6t
Xbit_r125_c135 bl[135] br[135] wl[125] vdd gnd cell_6t
Xbit_r126_c135 bl[135] br[135] wl[126] vdd gnd cell_6t
Xbit_r127_c135 bl[135] br[135] wl[127] vdd gnd cell_6t
Xbit_r128_c135 bl[135] br[135] wl[128] vdd gnd cell_6t
Xbit_r129_c135 bl[135] br[135] wl[129] vdd gnd cell_6t
Xbit_r130_c135 bl[135] br[135] wl[130] vdd gnd cell_6t
Xbit_r131_c135 bl[135] br[135] wl[131] vdd gnd cell_6t
Xbit_r132_c135 bl[135] br[135] wl[132] vdd gnd cell_6t
Xbit_r133_c135 bl[135] br[135] wl[133] vdd gnd cell_6t
Xbit_r134_c135 bl[135] br[135] wl[134] vdd gnd cell_6t
Xbit_r135_c135 bl[135] br[135] wl[135] vdd gnd cell_6t
Xbit_r136_c135 bl[135] br[135] wl[136] vdd gnd cell_6t
Xbit_r137_c135 bl[135] br[135] wl[137] vdd gnd cell_6t
Xbit_r138_c135 bl[135] br[135] wl[138] vdd gnd cell_6t
Xbit_r139_c135 bl[135] br[135] wl[139] vdd gnd cell_6t
Xbit_r140_c135 bl[135] br[135] wl[140] vdd gnd cell_6t
Xbit_r141_c135 bl[135] br[135] wl[141] vdd gnd cell_6t
Xbit_r142_c135 bl[135] br[135] wl[142] vdd gnd cell_6t
Xbit_r143_c135 bl[135] br[135] wl[143] vdd gnd cell_6t
Xbit_r144_c135 bl[135] br[135] wl[144] vdd gnd cell_6t
Xbit_r145_c135 bl[135] br[135] wl[145] vdd gnd cell_6t
Xbit_r146_c135 bl[135] br[135] wl[146] vdd gnd cell_6t
Xbit_r147_c135 bl[135] br[135] wl[147] vdd gnd cell_6t
Xbit_r148_c135 bl[135] br[135] wl[148] vdd gnd cell_6t
Xbit_r149_c135 bl[135] br[135] wl[149] vdd gnd cell_6t
Xbit_r150_c135 bl[135] br[135] wl[150] vdd gnd cell_6t
Xbit_r151_c135 bl[135] br[135] wl[151] vdd gnd cell_6t
Xbit_r152_c135 bl[135] br[135] wl[152] vdd gnd cell_6t
Xbit_r153_c135 bl[135] br[135] wl[153] vdd gnd cell_6t
Xbit_r154_c135 bl[135] br[135] wl[154] vdd gnd cell_6t
Xbit_r155_c135 bl[135] br[135] wl[155] vdd gnd cell_6t
Xbit_r156_c135 bl[135] br[135] wl[156] vdd gnd cell_6t
Xbit_r157_c135 bl[135] br[135] wl[157] vdd gnd cell_6t
Xbit_r158_c135 bl[135] br[135] wl[158] vdd gnd cell_6t
Xbit_r159_c135 bl[135] br[135] wl[159] vdd gnd cell_6t
Xbit_r160_c135 bl[135] br[135] wl[160] vdd gnd cell_6t
Xbit_r161_c135 bl[135] br[135] wl[161] vdd gnd cell_6t
Xbit_r162_c135 bl[135] br[135] wl[162] vdd gnd cell_6t
Xbit_r163_c135 bl[135] br[135] wl[163] vdd gnd cell_6t
Xbit_r164_c135 bl[135] br[135] wl[164] vdd gnd cell_6t
Xbit_r165_c135 bl[135] br[135] wl[165] vdd gnd cell_6t
Xbit_r166_c135 bl[135] br[135] wl[166] vdd gnd cell_6t
Xbit_r167_c135 bl[135] br[135] wl[167] vdd gnd cell_6t
Xbit_r168_c135 bl[135] br[135] wl[168] vdd gnd cell_6t
Xbit_r169_c135 bl[135] br[135] wl[169] vdd gnd cell_6t
Xbit_r170_c135 bl[135] br[135] wl[170] vdd gnd cell_6t
Xbit_r171_c135 bl[135] br[135] wl[171] vdd gnd cell_6t
Xbit_r172_c135 bl[135] br[135] wl[172] vdd gnd cell_6t
Xbit_r173_c135 bl[135] br[135] wl[173] vdd gnd cell_6t
Xbit_r174_c135 bl[135] br[135] wl[174] vdd gnd cell_6t
Xbit_r175_c135 bl[135] br[135] wl[175] vdd gnd cell_6t
Xbit_r176_c135 bl[135] br[135] wl[176] vdd gnd cell_6t
Xbit_r177_c135 bl[135] br[135] wl[177] vdd gnd cell_6t
Xbit_r178_c135 bl[135] br[135] wl[178] vdd gnd cell_6t
Xbit_r179_c135 bl[135] br[135] wl[179] vdd gnd cell_6t
Xbit_r180_c135 bl[135] br[135] wl[180] vdd gnd cell_6t
Xbit_r181_c135 bl[135] br[135] wl[181] vdd gnd cell_6t
Xbit_r182_c135 bl[135] br[135] wl[182] vdd gnd cell_6t
Xbit_r183_c135 bl[135] br[135] wl[183] vdd gnd cell_6t
Xbit_r184_c135 bl[135] br[135] wl[184] vdd gnd cell_6t
Xbit_r185_c135 bl[135] br[135] wl[185] vdd gnd cell_6t
Xbit_r186_c135 bl[135] br[135] wl[186] vdd gnd cell_6t
Xbit_r187_c135 bl[135] br[135] wl[187] vdd gnd cell_6t
Xbit_r188_c135 bl[135] br[135] wl[188] vdd gnd cell_6t
Xbit_r189_c135 bl[135] br[135] wl[189] vdd gnd cell_6t
Xbit_r190_c135 bl[135] br[135] wl[190] vdd gnd cell_6t
Xbit_r191_c135 bl[135] br[135] wl[191] vdd gnd cell_6t
Xbit_r192_c135 bl[135] br[135] wl[192] vdd gnd cell_6t
Xbit_r193_c135 bl[135] br[135] wl[193] vdd gnd cell_6t
Xbit_r194_c135 bl[135] br[135] wl[194] vdd gnd cell_6t
Xbit_r195_c135 bl[135] br[135] wl[195] vdd gnd cell_6t
Xbit_r196_c135 bl[135] br[135] wl[196] vdd gnd cell_6t
Xbit_r197_c135 bl[135] br[135] wl[197] vdd gnd cell_6t
Xbit_r198_c135 bl[135] br[135] wl[198] vdd gnd cell_6t
Xbit_r199_c135 bl[135] br[135] wl[199] vdd gnd cell_6t
Xbit_r200_c135 bl[135] br[135] wl[200] vdd gnd cell_6t
Xbit_r201_c135 bl[135] br[135] wl[201] vdd gnd cell_6t
Xbit_r202_c135 bl[135] br[135] wl[202] vdd gnd cell_6t
Xbit_r203_c135 bl[135] br[135] wl[203] vdd gnd cell_6t
Xbit_r204_c135 bl[135] br[135] wl[204] vdd gnd cell_6t
Xbit_r205_c135 bl[135] br[135] wl[205] vdd gnd cell_6t
Xbit_r206_c135 bl[135] br[135] wl[206] vdd gnd cell_6t
Xbit_r207_c135 bl[135] br[135] wl[207] vdd gnd cell_6t
Xbit_r208_c135 bl[135] br[135] wl[208] vdd gnd cell_6t
Xbit_r209_c135 bl[135] br[135] wl[209] vdd gnd cell_6t
Xbit_r210_c135 bl[135] br[135] wl[210] vdd gnd cell_6t
Xbit_r211_c135 bl[135] br[135] wl[211] vdd gnd cell_6t
Xbit_r212_c135 bl[135] br[135] wl[212] vdd gnd cell_6t
Xbit_r213_c135 bl[135] br[135] wl[213] vdd gnd cell_6t
Xbit_r214_c135 bl[135] br[135] wl[214] vdd gnd cell_6t
Xbit_r215_c135 bl[135] br[135] wl[215] vdd gnd cell_6t
Xbit_r216_c135 bl[135] br[135] wl[216] vdd gnd cell_6t
Xbit_r217_c135 bl[135] br[135] wl[217] vdd gnd cell_6t
Xbit_r218_c135 bl[135] br[135] wl[218] vdd gnd cell_6t
Xbit_r219_c135 bl[135] br[135] wl[219] vdd gnd cell_6t
Xbit_r220_c135 bl[135] br[135] wl[220] vdd gnd cell_6t
Xbit_r221_c135 bl[135] br[135] wl[221] vdd gnd cell_6t
Xbit_r222_c135 bl[135] br[135] wl[222] vdd gnd cell_6t
Xbit_r223_c135 bl[135] br[135] wl[223] vdd gnd cell_6t
Xbit_r224_c135 bl[135] br[135] wl[224] vdd gnd cell_6t
Xbit_r225_c135 bl[135] br[135] wl[225] vdd gnd cell_6t
Xbit_r226_c135 bl[135] br[135] wl[226] vdd gnd cell_6t
Xbit_r227_c135 bl[135] br[135] wl[227] vdd gnd cell_6t
Xbit_r228_c135 bl[135] br[135] wl[228] vdd gnd cell_6t
Xbit_r229_c135 bl[135] br[135] wl[229] vdd gnd cell_6t
Xbit_r230_c135 bl[135] br[135] wl[230] vdd gnd cell_6t
Xbit_r231_c135 bl[135] br[135] wl[231] vdd gnd cell_6t
Xbit_r232_c135 bl[135] br[135] wl[232] vdd gnd cell_6t
Xbit_r233_c135 bl[135] br[135] wl[233] vdd gnd cell_6t
Xbit_r234_c135 bl[135] br[135] wl[234] vdd gnd cell_6t
Xbit_r235_c135 bl[135] br[135] wl[235] vdd gnd cell_6t
Xbit_r236_c135 bl[135] br[135] wl[236] vdd gnd cell_6t
Xbit_r237_c135 bl[135] br[135] wl[237] vdd gnd cell_6t
Xbit_r238_c135 bl[135] br[135] wl[238] vdd gnd cell_6t
Xbit_r239_c135 bl[135] br[135] wl[239] vdd gnd cell_6t
Xbit_r240_c135 bl[135] br[135] wl[240] vdd gnd cell_6t
Xbit_r241_c135 bl[135] br[135] wl[241] vdd gnd cell_6t
Xbit_r242_c135 bl[135] br[135] wl[242] vdd gnd cell_6t
Xbit_r243_c135 bl[135] br[135] wl[243] vdd gnd cell_6t
Xbit_r244_c135 bl[135] br[135] wl[244] vdd gnd cell_6t
Xbit_r245_c135 bl[135] br[135] wl[245] vdd gnd cell_6t
Xbit_r246_c135 bl[135] br[135] wl[246] vdd gnd cell_6t
Xbit_r247_c135 bl[135] br[135] wl[247] vdd gnd cell_6t
Xbit_r248_c135 bl[135] br[135] wl[248] vdd gnd cell_6t
Xbit_r249_c135 bl[135] br[135] wl[249] vdd gnd cell_6t
Xbit_r250_c135 bl[135] br[135] wl[250] vdd gnd cell_6t
Xbit_r251_c135 bl[135] br[135] wl[251] vdd gnd cell_6t
Xbit_r252_c135 bl[135] br[135] wl[252] vdd gnd cell_6t
Xbit_r253_c135 bl[135] br[135] wl[253] vdd gnd cell_6t
Xbit_r254_c135 bl[135] br[135] wl[254] vdd gnd cell_6t
Xbit_r255_c135 bl[135] br[135] wl[255] vdd gnd cell_6t
Xbit_r0_c136 bl[136] br[136] wl[0] vdd gnd cell_6t
Xbit_r1_c136 bl[136] br[136] wl[1] vdd gnd cell_6t
Xbit_r2_c136 bl[136] br[136] wl[2] vdd gnd cell_6t
Xbit_r3_c136 bl[136] br[136] wl[3] vdd gnd cell_6t
Xbit_r4_c136 bl[136] br[136] wl[4] vdd gnd cell_6t
Xbit_r5_c136 bl[136] br[136] wl[5] vdd gnd cell_6t
Xbit_r6_c136 bl[136] br[136] wl[6] vdd gnd cell_6t
Xbit_r7_c136 bl[136] br[136] wl[7] vdd gnd cell_6t
Xbit_r8_c136 bl[136] br[136] wl[8] vdd gnd cell_6t
Xbit_r9_c136 bl[136] br[136] wl[9] vdd gnd cell_6t
Xbit_r10_c136 bl[136] br[136] wl[10] vdd gnd cell_6t
Xbit_r11_c136 bl[136] br[136] wl[11] vdd gnd cell_6t
Xbit_r12_c136 bl[136] br[136] wl[12] vdd gnd cell_6t
Xbit_r13_c136 bl[136] br[136] wl[13] vdd gnd cell_6t
Xbit_r14_c136 bl[136] br[136] wl[14] vdd gnd cell_6t
Xbit_r15_c136 bl[136] br[136] wl[15] vdd gnd cell_6t
Xbit_r16_c136 bl[136] br[136] wl[16] vdd gnd cell_6t
Xbit_r17_c136 bl[136] br[136] wl[17] vdd gnd cell_6t
Xbit_r18_c136 bl[136] br[136] wl[18] vdd gnd cell_6t
Xbit_r19_c136 bl[136] br[136] wl[19] vdd gnd cell_6t
Xbit_r20_c136 bl[136] br[136] wl[20] vdd gnd cell_6t
Xbit_r21_c136 bl[136] br[136] wl[21] vdd gnd cell_6t
Xbit_r22_c136 bl[136] br[136] wl[22] vdd gnd cell_6t
Xbit_r23_c136 bl[136] br[136] wl[23] vdd gnd cell_6t
Xbit_r24_c136 bl[136] br[136] wl[24] vdd gnd cell_6t
Xbit_r25_c136 bl[136] br[136] wl[25] vdd gnd cell_6t
Xbit_r26_c136 bl[136] br[136] wl[26] vdd gnd cell_6t
Xbit_r27_c136 bl[136] br[136] wl[27] vdd gnd cell_6t
Xbit_r28_c136 bl[136] br[136] wl[28] vdd gnd cell_6t
Xbit_r29_c136 bl[136] br[136] wl[29] vdd gnd cell_6t
Xbit_r30_c136 bl[136] br[136] wl[30] vdd gnd cell_6t
Xbit_r31_c136 bl[136] br[136] wl[31] vdd gnd cell_6t
Xbit_r32_c136 bl[136] br[136] wl[32] vdd gnd cell_6t
Xbit_r33_c136 bl[136] br[136] wl[33] vdd gnd cell_6t
Xbit_r34_c136 bl[136] br[136] wl[34] vdd gnd cell_6t
Xbit_r35_c136 bl[136] br[136] wl[35] vdd gnd cell_6t
Xbit_r36_c136 bl[136] br[136] wl[36] vdd gnd cell_6t
Xbit_r37_c136 bl[136] br[136] wl[37] vdd gnd cell_6t
Xbit_r38_c136 bl[136] br[136] wl[38] vdd gnd cell_6t
Xbit_r39_c136 bl[136] br[136] wl[39] vdd gnd cell_6t
Xbit_r40_c136 bl[136] br[136] wl[40] vdd gnd cell_6t
Xbit_r41_c136 bl[136] br[136] wl[41] vdd gnd cell_6t
Xbit_r42_c136 bl[136] br[136] wl[42] vdd gnd cell_6t
Xbit_r43_c136 bl[136] br[136] wl[43] vdd gnd cell_6t
Xbit_r44_c136 bl[136] br[136] wl[44] vdd gnd cell_6t
Xbit_r45_c136 bl[136] br[136] wl[45] vdd gnd cell_6t
Xbit_r46_c136 bl[136] br[136] wl[46] vdd gnd cell_6t
Xbit_r47_c136 bl[136] br[136] wl[47] vdd gnd cell_6t
Xbit_r48_c136 bl[136] br[136] wl[48] vdd gnd cell_6t
Xbit_r49_c136 bl[136] br[136] wl[49] vdd gnd cell_6t
Xbit_r50_c136 bl[136] br[136] wl[50] vdd gnd cell_6t
Xbit_r51_c136 bl[136] br[136] wl[51] vdd gnd cell_6t
Xbit_r52_c136 bl[136] br[136] wl[52] vdd gnd cell_6t
Xbit_r53_c136 bl[136] br[136] wl[53] vdd gnd cell_6t
Xbit_r54_c136 bl[136] br[136] wl[54] vdd gnd cell_6t
Xbit_r55_c136 bl[136] br[136] wl[55] vdd gnd cell_6t
Xbit_r56_c136 bl[136] br[136] wl[56] vdd gnd cell_6t
Xbit_r57_c136 bl[136] br[136] wl[57] vdd gnd cell_6t
Xbit_r58_c136 bl[136] br[136] wl[58] vdd gnd cell_6t
Xbit_r59_c136 bl[136] br[136] wl[59] vdd gnd cell_6t
Xbit_r60_c136 bl[136] br[136] wl[60] vdd gnd cell_6t
Xbit_r61_c136 bl[136] br[136] wl[61] vdd gnd cell_6t
Xbit_r62_c136 bl[136] br[136] wl[62] vdd gnd cell_6t
Xbit_r63_c136 bl[136] br[136] wl[63] vdd gnd cell_6t
Xbit_r64_c136 bl[136] br[136] wl[64] vdd gnd cell_6t
Xbit_r65_c136 bl[136] br[136] wl[65] vdd gnd cell_6t
Xbit_r66_c136 bl[136] br[136] wl[66] vdd gnd cell_6t
Xbit_r67_c136 bl[136] br[136] wl[67] vdd gnd cell_6t
Xbit_r68_c136 bl[136] br[136] wl[68] vdd gnd cell_6t
Xbit_r69_c136 bl[136] br[136] wl[69] vdd gnd cell_6t
Xbit_r70_c136 bl[136] br[136] wl[70] vdd gnd cell_6t
Xbit_r71_c136 bl[136] br[136] wl[71] vdd gnd cell_6t
Xbit_r72_c136 bl[136] br[136] wl[72] vdd gnd cell_6t
Xbit_r73_c136 bl[136] br[136] wl[73] vdd gnd cell_6t
Xbit_r74_c136 bl[136] br[136] wl[74] vdd gnd cell_6t
Xbit_r75_c136 bl[136] br[136] wl[75] vdd gnd cell_6t
Xbit_r76_c136 bl[136] br[136] wl[76] vdd gnd cell_6t
Xbit_r77_c136 bl[136] br[136] wl[77] vdd gnd cell_6t
Xbit_r78_c136 bl[136] br[136] wl[78] vdd gnd cell_6t
Xbit_r79_c136 bl[136] br[136] wl[79] vdd gnd cell_6t
Xbit_r80_c136 bl[136] br[136] wl[80] vdd gnd cell_6t
Xbit_r81_c136 bl[136] br[136] wl[81] vdd gnd cell_6t
Xbit_r82_c136 bl[136] br[136] wl[82] vdd gnd cell_6t
Xbit_r83_c136 bl[136] br[136] wl[83] vdd gnd cell_6t
Xbit_r84_c136 bl[136] br[136] wl[84] vdd gnd cell_6t
Xbit_r85_c136 bl[136] br[136] wl[85] vdd gnd cell_6t
Xbit_r86_c136 bl[136] br[136] wl[86] vdd gnd cell_6t
Xbit_r87_c136 bl[136] br[136] wl[87] vdd gnd cell_6t
Xbit_r88_c136 bl[136] br[136] wl[88] vdd gnd cell_6t
Xbit_r89_c136 bl[136] br[136] wl[89] vdd gnd cell_6t
Xbit_r90_c136 bl[136] br[136] wl[90] vdd gnd cell_6t
Xbit_r91_c136 bl[136] br[136] wl[91] vdd gnd cell_6t
Xbit_r92_c136 bl[136] br[136] wl[92] vdd gnd cell_6t
Xbit_r93_c136 bl[136] br[136] wl[93] vdd gnd cell_6t
Xbit_r94_c136 bl[136] br[136] wl[94] vdd gnd cell_6t
Xbit_r95_c136 bl[136] br[136] wl[95] vdd gnd cell_6t
Xbit_r96_c136 bl[136] br[136] wl[96] vdd gnd cell_6t
Xbit_r97_c136 bl[136] br[136] wl[97] vdd gnd cell_6t
Xbit_r98_c136 bl[136] br[136] wl[98] vdd gnd cell_6t
Xbit_r99_c136 bl[136] br[136] wl[99] vdd gnd cell_6t
Xbit_r100_c136 bl[136] br[136] wl[100] vdd gnd cell_6t
Xbit_r101_c136 bl[136] br[136] wl[101] vdd gnd cell_6t
Xbit_r102_c136 bl[136] br[136] wl[102] vdd gnd cell_6t
Xbit_r103_c136 bl[136] br[136] wl[103] vdd gnd cell_6t
Xbit_r104_c136 bl[136] br[136] wl[104] vdd gnd cell_6t
Xbit_r105_c136 bl[136] br[136] wl[105] vdd gnd cell_6t
Xbit_r106_c136 bl[136] br[136] wl[106] vdd gnd cell_6t
Xbit_r107_c136 bl[136] br[136] wl[107] vdd gnd cell_6t
Xbit_r108_c136 bl[136] br[136] wl[108] vdd gnd cell_6t
Xbit_r109_c136 bl[136] br[136] wl[109] vdd gnd cell_6t
Xbit_r110_c136 bl[136] br[136] wl[110] vdd gnd cell_6t
Xbit_r111_c136 bl[136] br[136] wl[111] vdd gnd cell_6t
Xbit_r112_c136 bl[136] br[136] wl[112] vdd gnd cell_6t
Xbit_r113_c136 bl[136] br[136] wl[113] vdd gnd cell_6t
Xbit_r114_c136 bl[136] br[136] wl[114] vdd gnd cell_6t
Xbit_r115_c136 bl[136] br[136] wl[115] vdd gnd cell_6t
Xbit_r116_c136 bl[136] br[136] wl[116] vdd gnd cell_6t
Xbit_r117_c136 bl[136] br[136] wl[117] vdd gnd cell_6t
Xbit_r118_c136 bl[136] br[136] wl[118] vdd gnd cell_6t
Xbit_r119_c136 bl[136] br[136] wl[119] vdd gnd cell_6t
Xbit_r120_c136 bl[136] br[136] wl[120] vdd gnd cell_6t
Xbit_r121_c136 bl[136] br[136] wl[121] vdd gnd cell_6t
Xbit_r122_c136 bl[136] br[136] wl[122] vdd gnd cell_6t
Xbit_r123_c136 bl[136] br[136] wl[123] vdd gnd cell_6t
Xbit_r124_c136 bl[136] br[136] wl[124] vdd gnd cell_6t
Xbit_r125_c136 bl[136] br[136] wl[125] vdd gnd cell_6t
Xbit_r126_c136 bl[136] br[136] wl[126] vdd gnd cell_6t
Xbit_r127_c136 bl[136] br[136] wl[127] vdd gnd cell_6t
Xbit_r128_c136 bl[136] br[136] wl[128] vdd gnd cell_6t
Xbit_r129_c136 bl[136] br[136] wl[129] vdd gnd cell_6t
Xbit_r130_c136 bl[136] br[136] wl[130] vdd gnd cell_6t
Xbit_r131_c136 bl[136] br[136] wl[131] vdd gnd cell_6t
Xbit_r132_c136 bl[136] br[136] wl[132] vdd gnd cell_6t
Xbit_r133_c136 bl[136] br[136] wl[133] vdd gnd cell_6t
Xbit_r134_c136 bl[136] br[136] wl[134] vdd gnd cell_6t
Xbit_r135_c136 bl[136] br[136] wl[135] vdd gnd cell_6t
Xbit_r136_c136 bl[136] br[136] wl[136] vdd gnd cell_6t
Xbit_r137_c136 bl[136] br[136] wl[137] vdd gnd cell_6t
Xbit_r138_c136 bl[136] br[136] wl[138] vdd gnd cell_6t
Xbit_r139_c136 bl[136] br[136] wl[139] vdd gnd cell_6t
Xbit_r140_c136 bl[136] br[136] wl[140] vdd gnd cell_6t
Xbit_r141_c136 bl[136] br[136] wl[141] vdd gnd cell_6t
Xbit_r142_c136 bl[136] br[136] wl[142] vdd gnd cell_6t
Xbit_r143_c136 bl[136] br[136] wl[143] vdd gnd cell_6t
Xbit_r144_c136 bl[136] br[136] wl[144] vdd gnd cell_6t
Xbit_r145_c136 bl[136] br[136] wl[145] vdd gnd cell_6t
Xbit_r146_c136 bl[136] br[136] wl[146] vdd gnd cell_6t
Xbit_r147_c136 bl[136] br[136] wl[147] vdd gnd cell_6t
Xbit_r148_c136 bl[136] br[136] wl[148] vdd gnd cell_6t
Xbit_r149_c136 bl[136] br[136] wl[149] vdd gnd cell_6t
Xbit_r150_c136 bl[136] br[136] wl[150] vdd gnd cell_6t
Xbit_r151_c136 bl[136] br[136] wl[151] vdd gnd cell_6t
Xbit_r152_c136 bl[136] br[136] wl[152] vdd gnd cell_6t
Xbit_r153_c136 bl[136] br[136] wl[153] vdd gnd cell_6t
Xbit_r154_c136 bl[136] br[136] wl[154] vdd gnd cell_6t
Xbit_r155_c136 bl[136] br[136] wl[155] vdd gnd cell_6t
Xbit_r156_c136 bl[136] br[136] wl[156] vdd gnd cell_6t
Xbit_r157_c136 bl[136] br[136] wl[157] vdd gnd cell_6t
Xbit_r158_c136 bl[136] br[136] wl[158] vdd gnd cell_6t
Xbit_r159_c136 bl[136] br[136] wl[159] vdd gnd cell_6t
Xbit_r160_c136 bl[136] br[136] wl[160] vdd gnd cell_6t
Xbit_r161_c136 bl[136] br[136] wl[161] vdd gnd cell_6t
Xbit_r162_c136 bl[136] br[136] wl[162] vdd gnd cell_6t
Xbit_r163_c136 bl[136] br[136] wl[163] vdd gnd cell_6t
Xbit_r164_c136 bl[136] br[136] wl[164] vdd gnd cell_6t
Xbit_r165_c136 bl[136] br[136] wl[165] vdd gnd cell_6t
Xbit_r166_c136 bl[136] br[136] wl[166] vdd gnd cell_6t
Xbit_r167_c136 bl[136] br[136] wl[167] vdd gnd cell_6t
Xbit_r168_c136 bl[136] br[136] wl[168] vdd gnd cell_6t
Xbit_r169_c136 bl[136] br[136] wl[169] vdd gnd cell_6t
Xbit_r170_c136 bl[136] br[136] wl[170] vdd gnd cell_6t
Xbit_r171_c136 bl[136] br[136] wl[171] vdd gnd cell_6t
Xbit_r172_c136 bl[136] br[136] wl[172] vdd gnd cell_6t
Xbit_r173_c136 bl[136] br[136] wl[173] vdd gnd cell_6t
Xbit_r174_c136 bl[136] br[136] wl[174] vdd gnd cell_6t
Xbit_r175_c136 bl[136] br[136] wl[175] vdd gnd cell_6t
Xbit_r176_c136 bl[136] br[136] wl[176] vdd gnd cell_6t
Xbit_r177_c136 bl[136] br[136] wl[177] vdd gnd cell_6t
Xbit_r178_c136 bl[136] br[136] wl[178] vdd gnd cell_6t
Xbit_r179_c136 bl[136] br[136] wl[179] vdd gnd cell_6t
Xbit_r180_c136 bl[136] br[136] wl[180] vdd gnd cell_6t
Xbit_r181_c136 bl[136] br[136] wl[181] vdd gnd cell_6t
Xbit_r182_c136 bl[136] br[136] wl[182] vdd gnd cell_6t
Xbit_r183_c136 bl[136] br[136] wl[183] vdd gnd cell_6t
Xbit_r184_c136 bl[136] br[136] wl[184] vdd gnd cell_6t
Xbit_r185_c136 bl[136] br[136] wl[185] vdd gnd cell_6t
Xbit_r186_c136 bl[136] br[136] wl[186] vdd gnd cell_6t
Xbit_r187_c136 bl[136] br[136] wl[187] vdd gnd cell_6t
Xbit_r188_c136 bl[136] br[136] wl[188] vdd gnd cell_6t
Xbit_r189_c136 bl[136] br[136] wl[189] vdd gnd cell_6t
Xbit_r190_c136 bl[136] br[136] wl[190] vdd gnd cell_6t
Xbit_r191_c136 bl[136] br[136] wl[191] vdd gnd cell_6t
Xbit_r192_c136 bl[136] br[136] wl[192] vdd gnd cell_6t
Xbit_r193_c136 bl[136] br[136] wl[193] vdd gnd cell_6t
Xbit_r194_c136 bl[136] br[136] wl[194] vdd gnd cell_6t
Xbit_r195_c136 bl[136] br[136] wl[195] vdd gnd cell_6t
Xbit_r196_c136 bl[136] br[136] wl[196] vdd gnd cell_6t
Xbit_r197_c136 bl[136] br[136] wl[197] vdd gnd cell_6t
Xbit_r198_c136 bl[136] br[136] wl[198] vdd gnd cell_6t
Xbit_r199_c136 bl[136] br[136] wl[199] vdd gnd cell_6t
Xbit_r200_c136 bl[136] br[136] wl[200] vdd gnd cell_6t
Xbit_r201_c136 bl[136] br[136] wl[201] vdd gnd cell_6t
Xbit_r202_c136 bl[136] br[136] wl[202] vdd gnd cell_6t
Xbit_r203_c136 bl[136] br[136] wl[203] vdd gnd cell_6t
Xbit_r204_c136 bl[136] br[136] wl[204] vdd gnd cell_6t
Xbit_r205_c136 bl[136] br[136] wl[205] vdd gnd cell_6t
Xbit_r206_c136 bl[136] br[136] wl[206] vdd gnd cell_6t
Xbit_r207_c136 bl[136] br[136] wl[207] vdd gnd cell_6t
Xbit_r208_c136 bl[136] br[136] wl[208] vdd gnd cell_6t
Xbit_r209_c136 bl[136] br[136] wl[209] vdd gnd cell_6t
Xbit_r210_c136 bl[136] br[136] wl[210] vdd gnd cell_6t
Xbit_r211_c136 bl[136] br[136] wl[211] vdd gnd cell_6t
Xbit_r212_c136 bl[136] br[136] wl[212] vdd gnd cell_6t
Xbit_r213_c136 bl[136] br[136] wl[213] vdd gnd cell_6t
Xbit_r214_c136 bl[136] br[136] wl[214] vdd gnd cell_6t
Xbit_r215_c136 bl[136] br[136] wl[215] vdd gnd cell_6t
Xbit_r216_c136 bl[136] br[136] wl[216] vdd gnd cell_6t
Xbit_r217_c136 bl[136] br[136] wl[217] vdd gnd cell_6t
Xbit_r218_c136 bl[136] br[136] wl[218] vdd gnd cell_6t
Xbit_r219_c136 bl[136] br[136] wl[219] vdd gnd cell_6t
Xbit_r220_c136 bl[136] br[136] wl[220] vdd gnd cell_6t
Xbit_r221_c136 bl[136] br[136] wl[221] vdd gnd cell_6t
Xbit_r222_c136 bl[136] br[136] wl[222] vdd gnd cell_6t
Xbit_r223_c136 bl[136] br[136] wl[223] vdd gnd cell_6t
Xbit_r224_c136 bl[136] br[136] wl[224] vdd gnd cell_6t
Xbit_r225_c136 bl[136] br[136] wl[225] vdd gnd cell_6t
Xbit_r226_c136 bl[136] br[136] wl[226] vdd gnd cell_6t
Xbit_r227_c136 bl[136] br[136] wl[227] vdd gnd cell_6t
Xbit_r228_c136 bl[136] br[136] wl[228] vdd gnd cell_6t
Xbit_r229_c136 bl[136] br[136] wl[229] vdd gnd cell_6t
Xbit_r230_c136 bl[136] br[136] wl[230] vdd gnd cell_6t
Xbit_r231_c136 bl[136] br[136] wl[231] vdd gnd cell_6t
Xbit_r232_c136 bl[136] br[136] wl[232] vdd gnd cell_6t
Xbit_r233_c136 bl[136] br[136] wl[233] vdd gnd cell_6t
Xbit_r234_c136 bl[136] br[136] wl[234] vdd gnd cell_6t
Xbit_r235_c136 bl[136] br[136] wl[235] vdd gnd cell_6t
Xbit_r236_c136 bl[136] br[136] wl[236] vdd gnd cell_6t
Xbit_r237_c136 bl[136] br[136] wl[237] vdd gnd cell_6t
Xbit_r238_c136 bl[136] br[136] wl[238] vdd gnd cell_6t
Xbit_r239_c136 bl[136] br[136] wl[239] vdd gnd cell_6t
Xbit_r240_c136 bl[136] br[136] wl[240] vdd gnd cell_6t
Xbit_r241_c136 bl[136] br[136] wl[241] vdd gnd cell_6t
Xbit_r242_c136 bl[136] br[136] wl[242] vdd gnd cell_6t
Xbit_r243_c136 bl[136] br[136] wl[243] vdd gnd cell_6t
Xbit_r244_c136 bl[136] br[136] wl[244] vdd gnd cell_6t
Xbit_r245_c136 bl[136] br[136] wl[245] vdd gnd cell_6t
Xbit_r246_c136 bl[136] br[136] wl[246] vdd gnd cell_6t
Xbit_r247_c136 bl[136] br[136] wl[247] vdd gnd cell_6t
Xbit_r248_c136 bl[136] br[136] wl[248] vdd gnd cell_6t
Xbit_r249_c136 bl[136] br[136] wl[249] vdd gnd cell_6t
Xbit_r250_c136 bl[136] br[136] wl[250] vdd gnd cell_6t
Xbit_r251_c136 bl[136] br[136] wl[251] vdd gnd cell_6t
Xbit_r252_c136 bl[136] br[136] wl[252] vdd gnd cell_6t
Xbit_r253_c136 bl[136] br[136] wl[253] vdd gnd cell_6t
Xbit_r254_c136 bl[136] br[136] wl[254] vdd gnd cell_6t
Xbit_r255_c136 bl[136] br[136] wl[255] vdd gnd cell_6t
Xbit_r0_c137 bl[137] br[137] wl[0] vdd gnd cell_6t
Xbit_r1_c137 bl[137] br[137] wl[1] vdd gnd cell_6t
Xbit_r2_c137 bl[137] br[137] wl[2] vdd gnd cell_6t
Xbit_r3_c137 bl[137] br[137] wl[3] vdd gnd cell_6t
Xbit_r4_c137 bl[137] br[137] wl[4] vdd gnd cell_6t
Xbit_r5_c137 bl[137] br[137] wl[5] vdd gnd cell_6t
Xbit_r6_c137 bl[137] br[137] wl[6] vdd gnd cell_6t
Xbit_r7_c137 bl[137] br[137] wl[7] vdd gnd cell_6t
Xbit_r8_c137 bl[137] br[137] wl[8] vdd gnd cell_6t
Xbit_r9_c137 bl[137] br[137] wl[9] vdd gnd cell_6t
Xbit_r10_c137 bl[137] br[137] wl[10] vdd gnd cell_6t
Xbit_r11_c137 bl[137] br[137] wl[11] vdd gnd cell_6t
Xbit_r12_c137 bl[137] br[137] wl[12] vdd gnd cell_6t
Xbit_r13_c137 bl[137] br[137] wl[13] vdd gnd cell_6t
Xbit_r14_c137 bl[137] br[137] wl[14] vdd gnd cell_6t
Xbit_r15_c137 bl[137] br[137] wl[15] vdd gnd cell_6t
Xbit_r16_c137 bl[137] br[137] wl[16] vdd gnd cell_6t
Xbit_r17_c137 bl[137] br[137] wl[17] vdd gnd cell_6t
Xbit_r18_c137 bl[137] br[137] wl[18] vdd gnd cell_6t
Xbit_r19_c137 bl[137] br[137] wl[19] vdd gnd cell_6t
Xbit_r20_c137 bl[137] br[137] wl[20] vdd gnd cell_6t
Xbit_r21_c137 bl[137] br[137] wl[21] vdd gnd cell_6t
Xbit_r22_c137 bl[137] br[137] wl[22] vdd gnd cell_6t
Xbit_r23_c137 bl[137] br[137] wl[23] vdd gnd cell_6t
Xbit_r24_c137 bl[137] br[137] wl[24] vdd gnd cell_6t
Xbit_r25_c137 bl[137] br[137] wl[25] vdd gnd cell_6t
Xbit_r26_c137 bl[137] br[137] wl[26] vdd gnd cell_6t
Xbit_r27_c137 bl[137] br[137] wl[27] vdd gnd cell_6t
Xbit_r28_c137 bl[137] br[137] wl[28] vdd gnd cell_6t
Xbit_r29_c137 bl[137] br[137] wl[29] vdd gnd cell_6t
Xbit_r30_c137 bl[137] br[137] wl[30] vdd gnd cell_6t
Xbit_r31_c137 bl[137] br[137] wl[31] vdd gnd cell_6t
Xbit_r32_c137 bl[137] br[137] wl[32] vdd gnd cell_6t
Xbit_r33_c137 bl[137] br[137] wl[33] vdd gnd cell_6t
Xbit_r34_c137 bl[137] br[137] wl[34] vdd gnd cell_6t
Xbit_r35_c137 bl[137] br[137] wl[35] vdd gnd cell_6t
Xbit_r36_c137 bl[137] br[137] wl[36] vdd gnd cell_6t
Xbit_r37_c137 bl[137] br[137] wl[37] vdd gnd cell_6t
Xbit_r38_c137 bl[137] br[137] wl[38] vdd gnd cell_6t
Xbit_r39_c137 bl[137] br[137] wl[39] vdd gnd cell_6t
Xbit_r40_c137 bl[137] br[137] wl[40] vdd gnd cell_6t
Xbit_r41_c137 bl[137] br[137] wl[41] vdd gnd cell_6t
Xbit_r42_c137 bl[137] br[137] wl[42] vdd gnd cell_6t
Xbit_r43_c137 bl[137] br[137] wl[43] vdd gnd cell_6t
Xbit_r44_c137 bl[137] br[137] wl[44] vdd gnd cell_6t
Xbit_r45_c137 bl[137] br[137] wl[45] vdd gnd cell_6t
Xbit_r46_c137 bl[137] br[137] wl[46] vdd gnd cell_6t
Xbit_r47_c137 bl[137] br[137] wl[47] vdd gnd cell_6t
Xbit_r48_c137 bl[137] br[137] wl[48] vdd gnd cell_6t
Xbit_r49_c137 bl[137] br[137] wl[49] vdd gnd cell_6t
Xbit_r50_c137 bl[137] br[137] wl[50] vdd gnd cell_6t
Xbit_r51_c137 bl[137] br[137] wl[51] vdd gnd cell_6t
Xbit_r52_c137 bl[137] br[137] wl[52] vdd gnd cell_6t
Xbit_r53_c137 bl[137] br[137] wl[53] vdd gnd cell_6t
Xbit_r54_c137 bl[137] br[137] wl[54] vdd gnd cell_6t
Xbit_r55_c137 bl[137] br[137] wl[55] vdd gnd cell_6t
Xbit_r56_c137 bl[137] br[137] wl[56] vdd gnd cell_6t
Xbit_r57_c137 bl[137] br[137] wl[57] vdd gnd cell_6t
Xbit_r58_c137 bl[137] br[137] wl[58] vdd gnd cell_6t
Xbit_r59_c137 bl[137] br[137] wl[59] vdd gnd cell_6t
Xbit_r60_c137 bl[137] br[137] wl[60] vdd gnd cell_6t
Xbit_r61_c137 bl[137] br[137] wl[61] vdd gnd cell_6t
Xbit_r62_c137 bl[137] br[137] wl[62] vdd gnd cell_6t
Xbit_r63_c137 bl[137] br[137] wl[63] vdd gnd cell_6t
Xbit_r64_c137 bl[137] br[137] wl[64] vdd gnd cell_6t
Xbit_r65_c137 bl[137] br[137] wl[65] vdd gnd cell_6t
Xbit_r66_c137 bl[137] br[137] wl[66] vdd gnd cell_6t
Xbit_r67_c137 bl[137] br[137] wl[67] vdd gnd cell_6t
Xbit_r68_c137 bl[137] br[137] wl[68] vdd gnd cell_6t
Xbit_r69_c137 bl[137] br[137] wl[69] vdd gnd cell_6t
Xbit_r70_c137 bl[137] br[137] wl[70] vdd gnd cell_6t
Xbit_r71_c137 bl[137] br[137] wl[71] vdd gnd cell_6t
Xbit_r72_c137 bl[137] br[137] wl[72] vdd gnd cell_6t
Xbit_r73_c137 bl[137] br[137] wl[73] vdd gnd cell_6t
Xbit_r74_c137 bl[137] br[137] wl[74] vdd gnd cell_6t
Xbit_r75_c137 bl[137] br[137] wl[75] vdd gnd cell_6t
Xbit_r76_c137 bl[137] br[137] wl[76] vdd gnd cell_6t
Xbit_r77_c137 bl[137] br[137] wl[77] vdd gnd cell_6t
Xbit_r78_c137 bl[137] br[137] wl[78] vdd gnd cell_6t
Xbit_r79_c137 bl[137] br[137] wl[79] vdd gnd cell_6t
Xbit_r80_c137 bl[137] br[137] wl[80] vdd gnd cell_6t
Xbit_r81_c137 bl[137] br[137] wl[81] vdd gnd cell_6t
Xbit_r82_c137 bl[137] br[137] wl[82] vdd gnd cell_6t
Xbit_r83_c137 bl[137] br[137] wl[83] vdd gnd cell_6t
Xbit_r84_c137 bl[137] br[137] wl[84] vdd gnd cell_6t
Xbit_r85_c137 bl[137] br[137] wl[85] vdd gnd cell_6t
Xbit_r86_c137 bl[137] br[137] wl[86] vdd gnd cell_6t
Xbit_r87_c137 bl[137] br[137] wl[87] vdd gnd cell_6t
Xbit_r88_c137 bl[137] br[137] wl[88] vdd gnd cell_6t
Xbit_r89_c137 bl[137] br[137] wl[89] vdd gnd cell_6t
Xbit_r90_c137 bl[137] br[137] wl[90] vdd gnd cell_6t
Xbit_r91_c137 bl[137] br[137] wl[91] vdd gnd cell_6t
Xbit_r92_c137 bl[137] br[137] wl[92] vdd gnd cell_6t
Xbit_r93_c137 bl[137] br[137] wl[93] vdd gnd cell_6t
Xbit_r94_c137 bl[137] br[137] wl[94] vdd gnd cell_6t
Xbit_r95_c137 bl[137] br[137] wl[95] vdd gnd cell_6t
Xbit_r96_c137 bl[137] br[137] wl[96] vdd gnd cell_6t
Xbit_r97_c137 bl[137] br[137] wl[97] vdd gnd cell_6t
Xbit_r98_c137 bl[137] br[137] wl[98] vdd gnd cell_6t
Xbit_r99_c137 bl[137] br[137] wl[99] vdd gnd cell_6t
Xbit_r100_c137 bl[137] br[137] wl[100] vdd gnd cell_6t
Xbit_r101_c137 bl[137] br[137] wl[101] vdd gnd cell_6t
Xbit_r102_c137 bl[137] br[137] wl[102] vdd gnd cell_6t
Xbit_r103_c137 bl[137] br[137] wl[103] vdd gnd cell_6t
Xbit_r104_c137 bl[137] br[137] wl[104] vdd gnd cell_6t
Xbit_r105_c137 bl[137] br[137] wl[105] vdd gnd cell_6t
Xbit_r106_c137 bl[137] br[137] wl[106] vdd gnd cell_6t
Xbit_r107_c137 bl[137] br[137] wl[107] vdd gnd cell_6t
Xbit_r108_c137 bl[137] br[137] wl[108] vdd gnd cell_6t
Xbit_r109_c137 bl[137] br[137] wl[109] vdd gnd cell_6t
Xbit_r110_c137 bl[137] br[137] wl[110] vdd gnd cell_6t
Xbit_r111_c137 bl[137] br[137] wl[111] vdd gnd cell_6t
Xbit_r112_c137 bl[137] br[137] wl[112] vdd gnd cell_6t
Xbit_r113_c137 bl[137] br[137] wl[113] vdd gnd cell_6t
Xbit_r114_c137 bl[137] br[137] wl[114] vdd gnd cell_6t
Xbit_r115_c137 bl[137] br[137] wl[115] vdd gnd cell_6t
Xbit_r116_c137 bl[137] br[137] wl[116] vdd gnd cell_6t
Xbit_r117_c137 bl[137] br[137] wl[117] vdd gnd cell_6t
Xbit_r118_c137 bl[137] br[137] wl[118] vdd gnd cell_6t
Xbit_r119_c137 bl[137] br[137] wl[119] vdd gnd cell_6t
Xbit_r120_c137 bl[137] br[137] wl[120] vdd gnd cell_6t
Xbit_r121_c137 bl[137] br[137] wl[121] vdd gnd cell_6t
Xbit_r122_c137 bl[137] br[137] wl[122] vdd gnd cell_6t
Xbit_r123_c137 bl[137] br[137] wl[123] vdd gnd cell_6t
Xbit_r124_c137 bl[137] br[137] wl[124] vdd gnd cell_6t
Xbit_r125_c137 bl[137] br[137] wl[125] vdd gnd cell_6t
Xbit_r126_c137 bl[137] br[137] wl[126] vdd gnd cell_6t
Xbit_r127_c137 bl[137] br[137] wl[127] vdd gnd cell_6t
Xbit_r128_c137 bl[137] br[137] wl[128] vdd gnd cell_6t
Xbit_r129_c137 bl[137] br[137] wl[129] vdd gnd cell_6t
Xbit_r130_c137 bl[137] br[137] wl[130] vdd gnd cell_6t
Xbit_r131_c137 bl[137] br[137] wl[131] vdd gnd cell_6t
Xbit_r132_c137 bl[137] br[137] wl[132] vdd gnd cell_6t
Xbit_r133_c137 bl[137] br[137] wl[133] vdd gnd cell_6t
Xbit_r134_c137 bl[137] br[137] wl[134] vdd gnd cell_6t
Xbit_r135_c137 bl[137] br[137] wl[135] vdd gnd cell_6t
Xbit_r136_c137 bl[137] br[137] wl[136] vdd gnd cell_6t
Xbit_r137_c137 bl[137] br[137] wl[137] vdd gnd cell_6t
Xbit_r138_c137 bl[137] br[137] wl[138] vdd gnd cell_6t
Xbit_r139_c137 bl[137] br[137] wl[139] vdd gnd cell_6t
Xbit_r140_c137 bl[137] br[137] wl[140] vdd gnd cell_6t
Xbit_r141_c137 bl[137] br[137] wl[141] vdd gnd cell_6t
Xbit_r142_c137 bl[137] br[137] wl[142] vdd gnd cell_6t
Xbit_r143_c137 bl[137] br[137] wl[143] vdd gnd cell_6t
Xbit_r144_c137 bl[137] br[137] wl[144] vdd gnd cell_6t
Xbit_r145_c137 bl[137] br[137] wl[145] vdd gnd cell_6t
Xbit_r146_c137 bl[137] br[137] wl[146] vdd gnd cell_6t
Xbit_r147_c137 bl[137] br[137] wl[147] vdd gnd cell_6t
Xbit_r148_c137 bl[137] br[137] wl[148] vdd gnd cell_6t
Xbit_r149_c137 bl[137] br[137] wl[149] vdd gnd cell_6t
Xbit_r150_c137 bl[137] br[137] wl[150] vdd gnd cell_6t
Xbit_r151_c137 bl[137] br[137] wl[151] vdd gnd cell_6t
Xbit_r152_c137 bl[137] br[137] wl[152] vdd gnd cell_6t
Xbit_r153_c137 bl[137] br[137] wl[153] vdd gnd cell_6t
Xbit_r154_c137 bl[137] br[137] wl[154] vdd gnd cell_6t
Xbit_r155_c137 bl[137] br[137] wl[155] vdd gnd cell_6t
Xbit_r156_c137 bl[137] br[137] wl[156] vdd gnd cell_6t
Xbit_r157_c137 bl[137] br[137] wl[157] vdd gnd cell_6t
Xbit_r158_c137 bl[137] br[137] wl[158] vdd gnd cell_6t
Xbit_r159_c137 bl[137] br[137] wl[159] vdd gnd cell_6t
Xbit_r160_c137 bl[137] br[137] wl[160] vdd gnd cell_6t
Xbit_r161_c137 bl[137] br[137] wl[161] vdd gnd cell_6t
Xbit_r162_c137 bl[137] br[137] wl[162] vdd gnd cell_6t
Xbit_r163_c137 bl[137] br[137] wl[163] vdd gnd cell_6t
Xbit_r164_c137 bl[137] br[137] wl[164] vdd gnd cell_6t
Xbit_r165_c137 bl[137] br[137] wl[165] vdd gnd cell_6t
Xbit_r166_c137 bl[137] br[137] wl[166] vdd gnd cell_6t
Xbit_r167_c137 bl[137] br[137] wl[167] vdd gnd cell_6t
Xbit_r168_c137 bl[137] br[137] wl[168] vdd gnd cell_6t
Xbit_r169_c137 bl[137] br[137] wl[169] vdd gnd cell_6t
Xbit_r170_c137 bl[137] br[137] wl[170] vdd gnd cell_6t
Xbit_r171_c137 bl[137] br[137] wl[171] vdd gnd cell_6t
Xbit_r172_c137 bl[137] br[137] wl[172] vdd gnd cell_6t
Xbit_r173_c137 bl[137] br[137] wl[173] vdd gnd cell_6t
Xbit_r174_c137 bl[137] br[137] wl[174] vdd gnd cell_6t
Xbit_r175_c137 bl[137] br[137] wl[175] vdd gnd cell_6t
Xbit_r176_c137 bl[137] br[137] wl[176] vdd gnd cell_6t
Xbit_r177_c137 bl[137] br[137] wl[177] vdd gnd cell_6t
Xbit_r178_c137 bl[137] br[137] wl[178] vdd gnd cell_6t
Xbit_r179_c137 bl[137] br[137] wl[179] vdd gnd cell_6t
Xbit_r180_c137 bl[137] br[137] wl[180] vdd gnd cell_6t
Xbit_r181_c137 bl[137] br[137] wl[181] vdd gnd cell_6t
Xbit_r182_c137 bl[137] br[137] wl[182] vdd gnd cell_6t
Xbit_r183_c137 bl[137] br[137] wl[183] vdd gnd cell_6t
Xbit_r184_c137 bl[137] br[137] wl[184] vdd gnd cell_6t
Xbit_r185_c137 bl[137] br[137] wl[185] vdd gnd cell_6t
Xbit_r186_c137 bl[137] br[137] wl[186] vdd gnd cell_6t
Xbit_r187_c137 bl[137] br[137] wl[187] vdd gnd cell_6t
Xbit_r188_c137 bl[137] br[137] wl[188] vdd gnd cell_6t
Xbit_r189_c137 bl[137] br[137] wl[189] vdd gnd cell_6t
Xbit_r190_c137 bl[137] br[137] wl[190] vdd gnd cell_6t
Xbit_r191_c137 bl[137] br[137] wl[191] vdd gnd cell_6t
Xbit_r192_c137 bl[137] br[137] wl[192] vdd gnd cell_6t
Xbit_r193_c137 bl[137] br[137] wl[193] vdd gnd cell_6t
Xbit_r194_c137 bl[137] br[137] wl[194] vdd gnd cell_6t
Xbit_r195_c137 bl[137] br[137] wl[195] vdd gnd cell_6t
Xbit_r196_c137 bl[137] br[137] wl[196] vdd gnd cell_6t
Xbit_r197_c137 bl[137] br[137] wl[197] vdd gnd cell_6t
Xbit_r198_c137 bl[137] br[137] wl[198] vdd gnd cell_6t
Xbit_r199_c137 bl[137] br[137] wl[199] vdd gnd cell_6t
Xbit_r200_c137 bl[137] br[137] wl[200] vdd gnd cell_6t
Xbit_r201_c137 bl[137] br[137] wl[201] vdd gnd cell_6t
Xbit_r202_c137 bl[137] br[137] wl[202] vdd gnd cell_6t
Xbit_r203_c137 bl[137] br[137] wl[203] vdd gnd cell_6t
Xbit_r204_c137 bl[137] br[137] wl[204] vdd gnd cell_6t
Xbit_r205_c137 bl[137] br[137] wl[205] vdd gnd cell_6t
Xbit_r206_c137 bl[137] br[137] wl[206] vdd gnd cell_6t
Xbit_r207_c137 bl[137] br[137] wl[207] vdd gnd cell_6t
Xbit_r208_c137 bl[137] br[137] wl[208] vdd gnd cell_6t
Xbit_r209_c137 bl[137] br[137] wl[209] vdd gnd cell_6t
Xbit_r210_c137 bl[137] br[137] wl[210] vdd gnd cell_6t
Xbit_r211_c137 bl[137] br[137] wl[211] vdd gnd cell_6t
Xbit_r212_c137 bl[137] br[137] wl[212] vdd gnd cell_6t
Xbit_r213_c137 bl[137] br[137] wl[213] vdd gnd cell_6t
Xbit_r214_c137 bl[137] br[137] wl[214] vdd gnd cell_6t
Xbit_r215_c137 bl[137] br[137] wl[215] vdd gnd cell_6t
Xbit_r216_c137 bl[137] br[137] wl[216] vdd gnd cell_6t
Xbit_r217_c137 bl[137] br[137] wl[217] vdd gnd cell_6t
Xbit_r218_c137 bl[137] br[137] wl[218] vdd gnd cell_6t
Xbit_r219_c137 bl[137] br[137] wl[219] vdd gnd cell_6t
Xbit_r220_c137 bl[137] br[137] wl[220] vdd gnd cell_6t
Xbit_r221_c137 bl[137] br[137] wl[221] vdd gnd cell_6t
Xbit_r222_c137 bl[137] br[137] wl[222] vdd gnd cell_6t
Xbit_r223_c137 bl[137] br[137] wl[223] vdd gnd cell_6t
Xbit_r224_c137 bl[137] br[137] wl[224] vdd gnd cell_6t
Xbit_r225_c137 bl[137] br[137] wl[225] vdd gnd cell_6t
Xbit_r226_c137 bl[137] br[137] wl[226] vdd gnd cell_6t
Xbit_r227_c137 bl[137] br[137] wl[227] vdd gnd cell_6t
Xbit_r228_c137 bl[137] br[137] wl[228] vdd gnd cell_6t
Xbit_r229_c137 bl[137] br[137] wl[229] vdd gnd cell_6t
Xbit_r230_c137 bl[137] br[137] wl[230] vdd gnd cell_6t
Xbit_r231_c137 bl[137] br[137] wl[231] vdd gnd cell_6t
Xbit_r232_c137 bl[137] br[137] wl[232] vdd gnd cell_6t
Xbit_r233_c137 bl[137] br[137] wl[233] vdd gnd cell_6t
Xbit_r234_c137 bl[137] br[137] wl[234] vdd gnd cell_6t
Xbit_r235_c137 bl[137] br[137] wl[235] vdd gnd cell_6t
Xbit_r236_c137 bl[137] br[137] wl[236] vdd gnd cell_6t
Xbit_r237_c137 bl[137] br[137] wl[237] vdd gnd cell_6t
Xbit_r238_c137 bl[137] br[137] wl[238] vdd gnd cell_6t
Xbit_r239_c137 bl[137] br[137] wl[239] vdd gnd cell_6t
Xbit_r240_c137 bl[137] br[137] wl[240] vdd gnd cell_6t
Xbit_r241_c137 bl[137] br[137] wl[241] vdd gnd cell_6t
Xbit_r242_c137 bl[137] br[137] wl[242] vdd gnd cell_6t
Xbit_r243_c137 bl[137] br[137] wl[243] vdd gnd cell_6t
Xbit_r244_c137 bl[137] br[137] wl[244] vdd gnd cell_6t
Xbit_r245_c137 bl[137] br[137] wl[245] vdd gnd cell_6t
Xbit_r246_c137 bl[137] br[137] wl[246] vdd gnd cell_6t
Xbit_r247_c137 bl[137] br[137] wl[247] vdd gnd cell_6t
Xbit_r248_c137 bl[137] br[137] wl[248] vdd gnd cell_6t
Xbit_r249_c137 bl[137] br[137] wl[249] vdd gnd cell_6t
Xbit_r250_c137 bl[137] br[137] wl[250] vdd gnd cell_6t
Xbit_r251_c137 bl[137] br[137] wl[251] vdd gnd cell_6t
Xbit_r252_c137 bl[137] br[137] wl[252] vdd gnd cell_6t
Xbit_r253_c137 bl[137] br[137] wl[253] vdd gnd cell_6t
Xbit_r254_c137 bl[137] br[137] wl[254] vdd gnd cell_6t
Xbit_r255_c137 bl[137] br[137] wl[255] vdd gnd cell_6t
Xbit_r0_c138 bl[138] br[138] wl[0] vdd gnd cell_6t
Xbit_r1_c138 bl[138] br[138] wl[1] vdd gnd cell_6t
Xbit_r2_c138 bl[138] br[138] wl[2] vdd gnd cell_6t
Xbit_r3_c138 bl[138] br[138] wl[3] vdd gnd cell_6t
Xbit_r4_c138 bl[138] br[138] wl[4] vdd gnd cell_6t
Xbit_r5_c138 bl[138] br[138] wl[5] vdd gnd cell_6t
Xbit_r6_c138 bl[138] br[138] wl[6] vdd gnd cell_6t
Xbit_r7_c138 bl[138] br[138] wl[7] vdd gnd cell_6t
Xbit_r8_c138 bl[138] br[138] wl[8] vdd gnd cell_6t
Xbit_r9_c138 bl[138] br[138] wl[9] vdd gnd cell_6t
Xbit_r10_c138 bl[138] br[138] wl[10] vdd gnd cell_6t
Xbit_r11_c138 bl[138] br[138] wl[11] vdd gnd cell_6t
Xbit_r12_c138 bl[138] br[138] wl[12] vdd gnd cell_6t
Xbit_r13_c138 bl[138] br[138] wl[13] vdd gnd cell_6t
Xbit_r14_c138 bl[138] br[138] wl[14] vdd gnd cell_6t
Xbit_r15_c138 bl[138] br[138] wl[15] vdd gnd cell_6t
Xbit_r16_c138 bl[138] br[138] wl[16] vdd gnd cell_6t
Xbit_r17_c138 bl[138] br[138] wl[17] vdd gnd cell_6t
Xbit_r18_c138 bl[138] br[138] wl[18] vdd gnd cell_6t
Xbit_r19_c138 bl[138] br[138] wl[19] vdd gnd cell_6t
Xbit_r20_c138 bl[138] br[138] wl[20] vdd gnd cell_6t
Xbit_r21_c138 bl[138] br[138] wl[21] vdd gnd cell_6t
Xbit_r22_c138 bl[138] br[138] wl[22] vdd gnd cell_6t
Xbit_r23_c138 bl[138] br[138] wl[23] vdd gnd cell_6t
Xbit_r24_c138 bl[138] br[138] wl[24] vdd gnd cell_6t
Xbit_r25_c138 bl[138] br[138] wl[25] vdd gnd cell_6t
Xbit_r26_c138 bl[138] br[138] wl[26] vdd gnd cell_6t
Xbit_r27_c138 bl[138] br[138] wl[27] vdd gnd cell_6t
Xbit_r28_c138 bl[138] br[138] wl[28] vdd gnd cell_6t
Xbit_r29_c138 bl[138] br[138] wl[29] vdd gnd cell_6t
Xbit_r30_c138 bl[138] br[138] wl[30] vdd gnd cell_6t
Xbit_r31_c138 bl[138] br[138] wl[31] vdd gnd cell_6t
Xbit_r32_c138 bl[138] br[138] wl[32] vdd gnd cell_6t
Xbit_r33_c138 bl[138] br[138] wl[33] vdd gnd cell_6t
Xbit_r34_c138 bl[138] br[138] wl[34] vdd gnd cell_6t
Xbit_r35_c138 bl[138] br[138] wl[35] vdd gnd cell_6t
Xbit_r36_c138 bl[138] br[138] wl[36] vdd gnd cell_6t
Xbit_r37_c138 bl[138] br[138] wl[37] vdd gnd cell_6t
Xbit_r38_c138 bl[138] br[138] wl[38] vdd gnd cell_6t
Xbit_r39_c138 bl[138] br[138] wl[39] vdd gnd cell_6t
Xbit_r40_c138 bl[138] br[138] wl[40] vdd gnd cell_6t
Xbit_r41_c138 bl[138] br[138] wl[41] vdd gnd cell_6t
Xbit_r42_c138 bl[138] br[138] wl[42] vdd gnd cell_6t
Xbit_r43_c138 bl[138] br[138] wl[43] vdd gnd cell_6t
Xbit_r44_c138 bl[138] br[138] wl[44] vdd gnd cell_6t
Xbit_r45_c138 bl[138] br[138] wl[45] vdd gnd cell_6t
Xbit_r46_c138 bl[138] br[138] wl[46] vdd gnd cell_6t
Xbit_r47_c138 bl[138] br[138] wl[47] vdd gnd cell_6t
Xbit_r48_c138 bl[138] br[138] wl[48] vdd gnd cell_6t
Xbit_r49_c138 bl[138] br[138] wl[49] vdd gnd cell_6t
Xbit_r50_c138 bl[138] br[138] wl[50] vdd gnd cell_6t
Xbit_r51_c138 bl[138] br[138] wl[51] vdd gnd cell_6t
Xbit_r52_c138 bl[138] br[138] wl[52] vdd gnd cell_6t
Xbit_r53_c138 bl[138] br[138] wl[53] vdd gnd cell_6t
Xbit_r54_c138 bl[138] br[138] wl[54] vdd gnd cell_6t
Xbit_r55_c138 bl[138] br[138] wl[55] vdd gnd cell_6t
Xbit_r56_c138 bl[138] br[138] wl[56] vdd gnd cell_6t
Xbit_r57_c138 bl[138] br[138] wl[57] vdd gnd cell_6t
Xbit_r58_c138 bl[138] br[138] wl[58] vdd gnd cell_6t
Xbit_r59_c138 bl[138] br[138] wl[59] vdd gnd cell_6t
Xbit_r60_c138 bl[138] br[138] wl[60] vdd gnd cell_6t
Xbit_r61_c138 bl[138] br[138] wl[61] vdd gnd cell_6t
Xbit_r62_c138 bl[138] br[138] wl[62] vdd gnd cell_6t
Xbit_r63_c138 bl[138] br[138] wl[63] vdd gnd cell_6t
Xbit_r64_c138 bl[138] br[138] wl[64] vdd gnd cell_6t
Xbit_r65_c138 bl[138] br[138] wl[65] vdd gnd cell_6t
Xbit_r66_c138 bl[138] br[138] wl[66] vdd gnd cell_6t
Xbit_r67_c138 bl[138] br[138] wl[67] vdd gnd cell_6t
Xbit_r68_c138 bl[138] br[138] wl[68] vdd gnd cell_6t
Xbit_r69_c138 bl[138] br[138] wl[69] vdd gnd cell_6t
Xbit_r70_c138 bl[138] br[138] wl[70] vdd gnd cell_6t
Xbit_r71_c138 bl[138] br[138] wl[71] vdd gnd cell_6t
Xbit_r72_c138 bl[138] br[138] wl[72] vdd gnd cell_6t
Xbit_r73_c138 bl[138] br[138] wl[73] vdd gnd cell_6t
Xbit_r74_c138 bl[138] br[138] wl[74] vdd gnd cell_6t
Xbit_r75_c138 bl[138] br[138] wl[75] vdd gnd cell_6t
Xbit_r76_c138 bl[138] br[138] wl[76] vdd gnd cell_6t
Xbit_r77_c138 bl[138] br[138] wl[77] vdd gnd cell_6t
Xbit_r78_c138 bl[138] br[138] wl[78] vdd gnd cell_6t
Xbit_r79_c138 bl[138] br[138] wl[79] vdd gnd cell_6t
Xbit_r80_c138 bl[138] br[138] wl[80] vdd gnd cell_6t
Xbit_r81_c138 bl[138] br[138] wl[81] vdd gnd cell_6t
Xbit_r82_c138 bl[138] br[138] wl[82] vdd gnd cell_6t
Xbit_r83_c138 bl[138] br[138] wl[83] vdd gnd cell_6t
Xbit_r84_c138 bl[138] br[138] wl[84] vdd gnd cell_6t
Xbit_r85_c138 bl[138] br[138] wl[85] vdd gnd cell_6t
Xbit_r86_c138 bl[138] br[138] wl[86] vdd gnd cell_6t
Xbit_r87_c138 bl[138] br[138] wl[87] vdd gnd cell_6t
Xbit_r88_c138 bl[138] br[138] wl[88] vdd gnd cell_6t
Xbit_r89_c138 bl[138] br[138] wl[89] vdd gnd cell_6t
Xbit_r90_c138 bl[138] br[138] wl[90] vdd gnd cell_6t
Xbit_r91_c138 bl[138] br[138] wl[91] vdd gnd cell_6t
Xbit_r92_c138 bl[138] br[138] wl[92] vdd gnd cell_6t
Xbit_r93_c138 bl[138] br[138] wl[93] vdd gnd cell_6t
Xbit_r94_c138 bl[138] br[138] wl[94] vdd gnd cell_6t
Xbit_r95_c138 bl[138] br[138] wl[95] vdd gnd cell_6t
Xbit_r96_c138 bl[138] br[138] wl[96] vdd gnd cell_6t
Xbit_r97_c138 bl[138] br[138] wl[97] vdd gnd cell_6t
Xbit_r98_c138 bl[138] br[138] wl[98] vdd gnd cell_6t
Xbit_r99_c138 bl[138] br[138] wl[99] vdd gnd cell_6t
Xbit_r100_c138 bl[138] br[138] wl[100] vdd gnd cell_6t
Xbit_r101_c138 bl[138] br[138] wl[101] vdd gnd cell_6t
Xbit_r102_c138 bl[138] br[138] wl[102] vdd gnd cell_6t
Xbit_r103_c138 bl[138] br[138] wl[103] vdd gnd cell_6t
Xbit_r104_c138 bl[138] br[138] wl[104] vdd gnd cell_6t
Xbit_r105_c138 bl[138] br[138] wl[105] vdd gnd cell_6t
Xbit_r106_c138 bl[138] br[138] wl[106] vdd gnd cell_6t
Xbit_r107_c138 bl[138] br[138] wl[107] vdd gnd cell_6t
Xbit_r108_c138 bl[138] br[138] wl[108] vdd gnd cell_6t
Xbit_r109_c138 bl[138] br[138] wl[109] vdd gnd cell_6t
Xbit_r110_c138 bl[138] br[138] wl[110] vdd gnd cell_6t
Xbit_r111_c138 bl[138] br[138] wl[111] vdd gnd cell_6t
Xbit_r112_c138 bl[138] br[138] wl[112] vdd gnd cell_6t
Xbit_r113_c138 bl[138] br[138] wl[113] vdd gnd cell_6t
Xbit_r114_c138 bl[138] br[138] wl[114] vdd gnd cell_6t
Xbit_r115_c138 bl[138] br[138] wl[115] vdd gnd cell_6t
Xbit_r116_c138 bl[138] br[138] wl[116] vdd gnd cell_6t
Xbit_r117_c138 bl[138] br[138] wl[117] vdd gnd cell_6t
Xbit_r118_c138 bl[138] br[138] wl[118] vdd gnd cell_6t
Xbit_r119_c138 bl[138] br[138] wl[119] vdd gnd cell_6t
Xbit_r120_c138 bl[138] br[138] wl[120] vdd gnd cell_6t
Xbit_r121_c138 bl[138] br[138] wl[121] vdd gnd cell_6t
Xbit_r122_c138 bl[138] br[138] wl[122] vdd gnd cell_6t
Xbit_r123_c138 bl[138] br[138] wl[123] vdd gnd cell_6t
Xbit_r124_c138 bl[138] br[138] wl[124] vdd gnd cell_6t
Xbit_r125_c138 bl[138] br[138] wl[125] vdd gnd cell_6t
Xbit_r126_c138 bl[138] br[138] wl[126] vdd gnd cell_6t
Xbit_r127_c138 bl[138] br[138] wl[127] vdd gnd cell_6t
Xbit_r128_c138 bl[138] br[138] wl[128] vdd gnd cell_6t
Xbit_r129_c138 bl[138] br[138] wl[129] vdd gnd cell_6t
Xbit_r130_c138 bl[138] br[138] wl[130] vdd gnd cell_6t
Xbit_r131_c138 bl[138] br[138] wl[131] vdd gnd cell_6t
Xbit_r132_c138 bl[138] br[138] wl[132] vdd gnd cell_6t
Xbit_r133_c138 bl[138] br[138] wl[133] vdd gnd cell_6t
Xbit_r134_c138 bl[138] br[138] wl[134] vdd gnd cell_6t
Xbit_r135_c138 bl[138] br[138] wl[135] vdd gnd cell_6t
Xbit_r136_c138 bl[138] br[138] wl[136] vdd gnd cell_6t
Xbit_r137_c138 bl[138] br[138] wl[137] vdd gnd cell_6t
Xbit_r138_c138 bl[138] br[138] wl[138] vdd gnd cell_6t
Xbit_r139_c138 bl[138] br[138] wl[139] vdd gnd cell_6t
Xbit_r140_c138 bl[138] br[138] wl[140] vdd gnd cell_6t
Xbit_r141_c138 bl[138] br[138] wl[141] vdd gnd cell_6t
Xbit_r142_c138 bl[138] br[138] wl[142] vdd gnd cell_6t
Xbit_r143_c138 bl[138] br[138] wl[143] vdd gnd cell_6t
Xbit_r144_c138 bl[138] br[138] wl[144] vdd gnd cell_6t
Xbit_r145_c138 bl[138] br[138] wl[145] vdd gnd cell_6t
Xbit_r146_c138 bl[138] br[138] wl[146] vdd gnd cell_6t
Xbit_r147_c138 bl[138] br[138] wl[147] vdd gnd cell_6t
Xbit_r148_c138 bl[138] br[138] wl[148] vdd gnd cell_6t
Xbit_r149_c138 bl[138] br[138] wl[149] vdd gnd cell_6t
Xbit_r150_c138 bl[138] br[138] wl[150] vdd gnd cell_6t
Xbit_r151_c138 bl[138] br[138] wl[151] vdd gnd cell_6t
Xbit_r152_c138 bl[138] br[138] wl[152] vdd gnd cell_6t
Xbit_r153_c138 bl[138] br[138] wl[153] vdd gnd cell_6t
Xbit_r154_c138 bl[138] br[138] wl[154] vdd gnd cell_6t
Xbit_r155_c138 bl[138] br[138] wl[155] vdd gnd cell_6t
Xbit_r156_c138 bl[138] br[138] wl[156] vdd gnd cell_6t
Xbit_r157_c138 bl[138] br[138] wl[157] vdd gnd cell_6t
Xbit_r158_c138 bl[138] br[138] wl[158] vdd gnd cell_6t
Xbit_r159_c138 bl[138] br[138] wl[159] vdd gnd cell_6t
Xbit_r160_c138 bl[138] br[138] wl[160] vdd gnd cell_6t
Xbit_r161_c138 bl[138] br[138] wl[161] vdd gnd cell_6t
Xbit_r162_c138 bl[138] br[138] wl[162] vdd gnd cell_6t
Xbit_r163_c138 bl[138] br[138] wl[163] vdd gnd cell_6t
Xbit_r164_c138 bl[138] br[138] wl[164] vdd gnd cell_6t
Xbit_r165_c138 bl[138] br[138] wl[165] vdd gnd cell_6t
Xbit_r166_c138 bl[138] br[138] wl[166] vdd gnd cell_6t
Xbit_r167_c138 bl[138] br[138] wl[167] vdd gnd cell_6t
Xbit_r168_c138 bl[138] br[138] wl[168] vdd gnd cell_6t
Xbit_r169_c138 bl[138] br[138] wl[169] vdd gnd cell_6t
Xbit_r170_c138 bl[138] br[138] wl[170] vdd gnd cell_6t
Xbit_r171_c138 bl[138] br[138] wl[171] vdd gnd cell_6t
Xbit_r172_c138 bl[138] br[138] wl[172] vdd gnd cell_6t
Xbit_r173_c138 bl[138] br[138] wl[173] vdd gnd cell_6t
Xbit_r174_c138 bl[138] br[138] wl[174] vdd gnd cell_6t
Xbit_r175_c138 bl[138] br[138] wl[175] vdd gnd cell_6t
Xbit_r176_c138 bl[138] br[138] wl[176] vdd gnd cell_6t
Xbit_r177_c138 bl[138] br[138] wl[177] vdd gnd cell_6t
Xbit_r178_c138 bl[138] br[138] wl[178] vdd gnd cell_6t
Xbit_r179_c138 bl[138] br[138] wl[179] vdd gnd cell_6t
Xbit_r180_c138 bl[138] br[138] wl[180] vdd gnd cell_6t
Xbit_r181_c138 bl[138] br[138] wl[181] vdd gnd cell_6t
Xbit_r182_c138 bl[138] br[138] wl[182] vdd gnd cell_6t
Xbit_r183_c138 bl[138] br[138] wl[183] vdd gnd cell_6t
Xbit_r184_c138 bl[138] br[138] wl[184] vdd gnd cell_6t
Xbit_r185_c138 bl[138] br[138] wl[185] vdd gnd cell_6t
Xbit_r186_c138 bl[138] br[138] wl[186] vdd gnd cell_6t
Xbit_r187_c138 bl[138] br[138] wl[187] vdd gnd cell_6t
Xbit_r188_c138 bl[138] br[138] wl[188] vdd gnd cell_6t
Xbit_r189_c138 bl[138] br[138] wl[189] vdd gnd cell_6t
Xbit_r190_c138 bl[138] br[138] wl[190] vdd gnd cell_6t
Xbit_r191_c138 bl[138] br[138] wl[191] vdd gnd cell_6t
Xbit_r192_c138 bl[138] br[138] wl[192] vdd gnd cell_6t
Xbit_r193_c138 bl[138] br[138] wl[193] vdd gnd cell_6t
Xbit_r194_c138 bl[138] br[138] wl[194] vdd gnd cell_6t
Xbit_r195_c138 bl[138] br[138] wl[195] vdd gnd cell_6t
Xbit_r196_c138 bl[138] br[138] wl[196] vdd gnd cell_6t
Xbit_r197_c138 bl[138] br[138] wl[197] vdd gnd cell_6t
Xbit_r198_c138 bl[138] br[138] wl[198] vdd gnd cell_6t
Xbit_r199_c138 bl[138] br[138] wl[199] vdd gnd cell_6t
Xbit_r200_c138 bl[138] br[138] wl[200] vdd gnd cell_6t
Xbit_r201_c138 bl[138] br[138] wl[201] vdd gnd cell_6t
Xbit_r202_c138 bl[138] br[138] wl[202] vdd gnd cell_6t
Xbit_r203_c138 bl[138] br[138] wl[203] vdd gnd cell_6t
Xbit_r204_c138 bl[138] br[138] wl[204] vdd gnd cell_6t
Xbit_r205_c138 bl[138] br[138] wl[205] vdd gnd cell_6t
Xbit_r206_c138 bl[138] br[138] wl[206] vdd gnd cell_6t
Xbit_r207_c138 bl[138] br[138] wl[207] vdd gnd cell_6t
Xbit_r208_c138 bl[138] br[138] wl[208] vdd gnd cell_6t
Xbit_r209_c138 bl[138] br[138] wl[209] vdd gnd cell_6t
Xbit_r210_c138 bl[138] br[138] wl[210] vdd gnd cell_6t
Xbit_r211_c138 bl[138] br[138] wl[211] vdd gnd cell_6t
Xbit_r212_c138 bl[138] br[138] wl[212] vdd gnd cell_6t
Xbit_r213_c138 bl[138] br[138] wl[213] vdd gnd cell_6t
Xbit_r214_c138 bl[138] br[138] wl[214] vdd gnd cell_6t
Xbit_r215_c138 bl[138] br[138] wl[215] vdd gnd cell_6t
Xbit_r216_c138 bl[138] br[138] wl[216] vdd gnd cell_6t
Xbit_r217_c138 bl[138] br[138] wl[217] vdd gnd cell_6t
Xbit_r218_c138 bl[138] br[138] wl[218] vdd gnd cell_6t
Xbit_r219_c138 bl[138] br[138] wl[219] vdd gnd cell_6t
Xbit_r220_c138 bl[138] br[138] wl[220] vdd gnd cell_6t
Xbit_r221_c138 bl[138] br[138] wl[221] vdd gnd cell_6t
Xbit_r222_c138 bl[138] br[138] wl[222] vdd gnd cell_6t
Xbit_r223_c138 bl[138] br[138] wl[223] vdd gnd cell_6t
Xbit_r224_c138 bl[138] br[138] wl[224] vdd gnd cell_6t
Xbit_r225_c138 bl[138] br[138] wl[225] vdd gnd cell_6t
Xbit_r226_c138 bl[138] br[138] wl[226] vdd gnd cell_6t
Xbit_r227_c138 bl[138] br[138] wl[227] vdd gnd cell_6t
Xbit_r228_c138 bl[138] br[138] wl[228] vdd gnd cell_6t
Xbit_r229_c138 bl[138] br[138] wl[229] vdd gnd cell_6t
Xbit_r230_c138 bl[138] br[138] wl[230] vdd gnd cell_6t
Xbit_r231_c138 bl[138] br[138] wl[231] vdd gnd cell_6t
Xbit_r232_c138 bl[138] br[138] wl[232] vdd gnd cell_6t
Xbit_r233_c138 bl[138] br[138] wl[233] vdd gnd cell_6t
Xbit_r234_c138 bl[138] br[138] wl[234] vdd gnd cell_6t
Xbit_r235_c138 bl[138] br[138] wl[235] vdd gnd cell_6t
Xbit_r236_c138 bl[138] br[138] wl[236] vdd gnd cell_6t
Xbit_r237_c138 bl[138] br[138] wl[237] vdd gnd cell_6t
Xbit_r238_c138 bl[138] br[138] wl[238] vdd gnd cell_6t
Xbit_r239_c138 bl[138] br[138] wl[239] vdd gnd cell_6t
Xbit_r240_c138 bl[138] br[138] wl[240] vdd gnd cell_6t
Xbit_r241_c138 bl[138] br[138] wl[241] vdd gnd cell_6t
Xbit_r242_c138 bl[138] br[138] wl[242] vdd gnd cell_6t
Xbit_r243_c138 bl[138] br[138] wl[243] vdd gnd cell_6t
Xbit_r244_c138 bl[138] br[138] wl[244] vdd gnd cell_6t
Xbit_r245_c138 bl[138] br[138] wl[245] vdd gnd cell_6t
Xbit_r246_c138 bl[138] br[138] wl[246] vdd gnd cell_6t
Xbit_r247_c138 bl[138] br[138] wl[247] vdd gnd cell_6t
Xbit_r248_c138 bl[138] br[138] wl[248] vdd gnd cell_6t
Xbit_r249_c138 bl[138] br[138] wl[249] vdd gnd cell_6t
Xbit_r250_c138 bl[138] br[138] wl[250] vdd gnd cell_6t
Xbit_r251_c138 bl[138] br[138] wl[251] vdd gnd cell_6t
Xbit_r252_c138 bl[138] br[138] wl[252] vdd gnd cell_6t
Xbit_r253_c138 bl[138] br[138] wl[253] vdd gnd cell_6t
Xbit_r254_c138 bl[138] br[138] wl[254] vdd gnd cell_6t
Xbit_r255_c138 bl[138] br[138] wl[255] vdd gnd cell_6t
Xbit_r0_c139 bl[139] br[139] wl[0] vdd gnd cell_6t
Xbit_r1_c139 bl[139] br[139] wl[1] vdd gnd cell_6t
Xbit_r2_c139 bl[139] br[139] wl[2] vdd gnd cell_6t
Xbit_r3_c139 bl[139] br[139] wl[3] vdd gnd cell_6t
Xbit_r4_c139 bl[139] br[139] wl[4] vdd gnd cell_6t
Xbit_r5_c139 bl[139] br[139] wl[5] vdd gnd cell_6t
Xbit_r6_c139 bl[139] br[139] wl[6] vdd gnd cell_6t
Xbit_r7_c139 bl[139] br[139] wl[7] vdd gnd cell_6t
Xbit_r8_c139 bl[139] br[139] wl[8] vdd gnd cell_6t
Xbit_r9_c139 bl[139] br[139] wl[9] vdd gnd cell_6t
Xbit_r10_c139 bl[139] br[139] wl[10] vdd gnd cell_6t
Xbit_r11_c139 bl[139] br[139] wl[11] vdd gnd cell_6t
Xbit_r12_c139 bl[139] br[139] wl[12] vdd gnd cell_6t
Xbit_r13_c139 bl[139] br[139] wl[13] vdd gnd cell_6t
Xbit_r14_c139 bl[139] br[139] wl[14] vdd gnd cell_6t
Xbit_r15_c139 bl[139] br[139] wl[15] vdd gnd cell_6t
Xbit_r16_c139 bl[139] br[139] wl[16] vdd gnd cell_6t
Xbit_r17_c139 bl[139] br[139] wl[17] vdd gnd cell_6t
Xbit_r18_c139 bl[139] br[139] wl[18] vdd gnd cell_6t
Xbit_r19_c139 bl[139] br[139] wl[19] vdd gnd cell_6t
Xbit_r20_c139 bl[139] br[139] wl[20] vdd gnd cell_6t
Xbit_r21_c139 bl[139] br[139] wl[21] vdd gnd cell_6t
Xbit_r22_c139 bl[139] br[139] wl[22] vdd gnd cell_6t
Xbit_r23_c139 bl[139] br[139] wl[23] vdd gnd cell_6t
Xbit_r24_c139 bl[139] br[139] wl[24] vdd gnd cell_6t
Xbit_r25_c139 bl[139] br[139] wl[25] vdd gnd cell_6t
Xbit_r26_c139 bl[139] br[139] wl[26] vdd gnd cell_6t
Xbit_r27_c139 bl[139] br[139] wl[27] vdd gnd cell_6t
Xbit_r28_c139 bl[139] br[139] wl[28] vdd gnd cell_6t
Xbit_r29_c139 bl[139] br[139] wl[29] vdd gnd cell_6t
Xbit_r30_c139 bl[139] br[139] wl[30] vdd gnd cell_6t
Xbit_r31_c139 bl[139] br[139] wl[31] vdd gnd cell_6t
Xbit_r32_c139 bl[139] br[139] wl[32] vdd gnd cell_6t
Xbit_r33_c139 bl[139] br[139] wl[33] vdd gnd cell_6t
Xbit_r34_c139 bl[139] br[139] wl[34] vdd gnd cell_6t
Xbit_r35_c139 bl[139] br[139] wl[35] vdd gnd cell_6t
Xbit_r36_c139 bl[139] br[139] wl[36] vdd gnd cell_6t
Xbit_r37_c139 bl[139] br[139] wl[37] vdd gnd cell_6t
Xbit_r38_c139 bl[139] br[139] wl[38] vdd gnd cell_6t
Xbit_r39_c139 bl[139] br[139] wl[39] vdd gnd cell_6t
Xbit_r40_c139 bl[139] br[139] wl[40] vdd gnd cell_6t
Xbit_r41_c139 bl[139] br[139] wl[41] vdd gnd cell_6t
Xbit_r42_c139 bl[139] br[139] wl[42] vdd gnd cell_6t
Xbit_r43_c139 bl[139] br[139] wl[43] vdd gnd cell_6t
Xbit_r44_c139 bl[139] br[139] wl[44] vdd gnd cell_6t
Xbit_r45_c139 bl[139] br[139] wl[45] vdd gnd cell_6t
Xbit_r46_c139 bl[139] br[139] wl[46] vdd gnd cell_6t
Xbit_r47_c139 bl[139] br[139] wl[47] vdd gnd cell_6t
Xbit_r48_c139 bl[139] br[139] wl[48] vdd gnd cell_6t
Xbit_r49_c139 bl[139] br[139] wl[49] vdd gnd cell_6t
Xbit_r50_c139 bl[139] br[139] wl[50] vdd gnd cell_6t
Xbit_r51_c139 bl[139] br[139] wl[51] vdd gnd cell_6t
Xbit_r52_c139 bl[139] br[139] wl[52] vdd gnd cell_6t
Xbit_r53_c139 bl[139] br[139] wl[53] vdd gnd cell_6t
Xbit_r54_c139 bl[139] br[139] wl[54] vdd gnd cell_6t
Xbit_r55_c139 bl[139] br[139] wl[55] vdd gnd cell_6t
Xbit_r56_c139 bl[139] br[139] wl[56] vdd gnd cell_6t
Xbit_r57_c139 bl[139] br[139] wl[57] vdd gnd cell_6t
Xbit_r58_c139 bl[139] br[139] wl[58] vdd gnd cell_6t
Xbit_r59_c139 bl[139] br[139] wl[59] vdd gnd cell_6t
Xbit_r60_c139 bl[139] br[139] wl[60] vdd gnd cell_6t
Xbit_r61_c139 bl[139] br[139] wl[61] vdd gnd cell_6t
Xbit_r62_c139 bl[139] br[139] wl[62] vdd gnd cell_6t
Xbit_r63_c139 bl[139] br[139] wl[63] vdd gnd cell_6t
Xbit_r64_c139 bl[139] br[139] wl[64] vdd gnd cell_6t
Xbit_r65_c139 bl[139] br[139] wl[65] vdd gnd cell_6t
Xbit_r66_c139 bl[139] br[139] wl[66] vdd gnd cell_6t
Xbit_r67_c139 bl[139] br[139] wl[67] vdd gnd cell_6t
Xbit_r68_c139 bl[139] br[139] wl[68] vdd gnd cell_6t
Xbit_r69_c139 bl[139] br[139] wl[69] vdd gnd cell_6t
Xbit_r70_c139 bl[139] br[139] wl[70] vdd gnd cell_6t
Xbit_r71_c139 bl[139] br[139] wl[71] vdd gnd cell_6t
Xbit_r72_c139 bl[139] br[139] wl[72] vdd gnd cell_6t
Xbit_r73_c139 bl[139] br[139] wl[73] vdd gnd cell_6t
Xbit_r74_c139 bl[139] br[139] wl[74] vdd gnd cell_6t
Xbit_r75_c139 bl[139] br[139] wl[75] vdd gnd cell_6t
Xbit_r76_c139 bl[139] br[139] wl[76] vdd gnd cell_6t
Xbit_r77_c139 bl[139] br[139] wl[77] vdd gnd cell_6t
Xbit_r78_c139 bl[139] br[139] wl[78] vdd gnd cell_6t
Xbit_r79_c139 bl[139] br[139] wl[79] vdd gnd cell_6t
Xbit_r80_c139 bl[139] br[139] wl[80] vdd gnd cell_6t
Xbit_r81_c139 bl[139] br[139] wl[81] vdd gnd cell_6t
Xbit_r82_c139 bl[139] br[139] wl[82] vdd gnd cell_6t
Xbit_r83_c139 bl[139] br[139] wl[83] vdd gnd cell_6t
Xbit_r84_c139 bl[139] br[139] wl[84] vdd gnd cell_6t
Xbit_r85_c139 bl[139] br[139] wl[85] vdd gnd cell_6t
Xbit_r86_c139 bl[139] br[139] wl[86] vdd gnd cell_6t
Xbit_r87_c139 bl[139] br[139] wl[87] vdd gnd cell_6t
Xbit_r88_c139 bl[139] br[139] wl[88] vdd gnd cell_6t
Xbit_r89_c139 bl[139] br[139] wl[89] vdd gnd cell_6t
Xbit_r90_c139 bl[139] br[139] wl[90] vdd gnd cell_6t
Xbit_r91_c139 bl[139] br[139] wl[91] vdd gnd cell_6t
Xbit_r92_c139 bl[139] br[139] wl[92] vdd gnd cell_6t
Xbit_r93_c139 bl[139] br[139] wl[93] vdd gnd cell_6t
Xbit_r94_c139 bl[139] br[139] wl[94] vdd gnd cell_6t
Xbit_r95_c139 bl[139] br[139] wl[95] vdd gnd cell_6t
Xbit_r96_c139 bl[139] br[139] wl[96] vdd gnd cell_6t
Xbit_r97_c139 bl[139] br[139] wl[97] vdd gnd cell_6t
Xbit_r98_c139 bl[139] br[139] wl[98] vdd gnd cell_6t
Xbit_r99_c139 bl[139] br[139] wl[99] vdd gnd cell_6t
Xbit_r100_c139 bl[139] br[139] wl[100] vdd gnd cell_6t
Xbit_r101_c139 bl[139] br[139] wl[101] vdd gnd cell_6t
Xbit_r102_c139 bl[139] br[139] wl[102] vdd gnd cell_6t
Xbit_r103_c139 bl[139] br[139] wl[103] vdd gnd cell_6t
Xbit_r104_c139 bl[139] br[139] wl[104] vdd gnd cell_6t
Xbit_r105_c139 bl[139] br[139] wl[105] vdd gnd cell_6t
Xbit_r106_c139 bl[139] br[139] wl[106] vdd gnd cell_6t
Xbit_r107_c139 bl[139] br[139] wl[107] vdd gnd cell_6t
Xbit_r108_c139 bl[139] br[139] wl[108] vdd gnd cell_6t
Xbit_r109_c139 bl[139] br[139] wl[109] vdd gnd cell_6t
Xbit_r110_c139 bl[139] br[139] wl[110] vdd gnd cell_6t
Xbit_r111_c139 bl[139] br[139] wl[111] vdd gnd cell_6t
Xbit_r112_c139 bl[139] br[139] wl[112] vdd gnd cell_6t
Xbit_r113_c139 bl[139] br[139] wl[113] vdd gnd cell_6t
Xbit_r114_c139 bl[139] br[139] wl[114] vdd gnd cell_6t
Xbit_r115_c139 bl[139] br[139] wl[115] vdd gnd cell_6t
Xbit_r116_c139 bl[139] br[139] wl[116] vdd gnd cell_6t
Xbit_r117_c139 bl[139] br[139] wl[117] vdd gnd cell_6t
Xbit_r118_c139 bl[139] br[139] wl[118] vdd gnd cell_6t
Xbit_r119_c139 bl[139] br[139] wl[119] vdd gnd cell_6t
Xbit_r120_c139 bl[139] br[139] wl[120] vdd gnd cell_6t
Xbit_r121_c139 bl[139] br[139] wl[121] vdd gnd cell_6t
Xbit_r122_c139 bl[139] br[139] wl[122] vdd gnd cell_6t
Xbit_r123_c139 bl[139] br[139] wl[123] vdd gnd cell_6t
Xbit_r124_c139 bl[139] br[139] wl[124] vdd gnd cell_6t
Xbit_r125_c139 bl[139] br[139] wl[125] vdd gnd cell_6t
Xbit_r126_c139 bl[139] br[139] wl[126] vdd gnd cell_6t
Xbit_r127_c139 bl[139] br[139] wl[127] vdd gnd cell_6t
Xbit_r128_c139 bl[139] br[139] wl[128] vdd gnd cell_6t
Xbit_r129_c139 bl[139] br[139] wl[129] vdd gnd cell_6t
Xbit_r130_c139 bl[139] br[139] wl[130] vdd gnd cell_6t
Xbit_r131_c139 bl[139] br[139] wl[131] vdd gnd cell_6t
Xbit_r132_c139 bl[139] br[139] wl[132] vdd gnd cell_6t
Xbit_r133_c139 bl[139] br[139] wl[133] vdd gnd cell_6t
Xbit_r134_c139 bl[139] br[139] wl[134] vdd gnd cell_6t
Xbit_r135_c139 bl[139] br[139] wl[135] vdd gnd cell_6t
Xbit_r136_c139 bl[139] br[139] wl[136] vdd gnd cell_6t
Xbit_r137_c139 bl[139] br[139] wl[137] vdd gnd cell_6t
Xbit_r138_c139 bl[139] br[139] wl[138] vdd gnd cell_6t
Xbit_r139_c139 bl[139] br[139] wl[139] vdd gnd cell_6t
Xbit_r140_c139 bl[139] br[139] wl[140] vdd gnd cell_6t
Xbit_r141_c139 bl[139] br[139] wl[141] vdd gnd cell_6t
Xbit_r142_c139 bl[139] br[139] wl[142] vdd gnd cell_6t
Xbit_r143_c139 bl[139] br[139] wl[143] vdd gnd cell_6t
Xbit_r144_c139 bl[139] br[139] wl[144] vdd gnd cell_6t
Xbit_r145_c139 bl[139] br[139] wl[145] vdd gnd cell_6t
Xbit_r146_c139 bl[139] br[139] wl[146] vdd gnd cell_6t
Xbit_r147_c139 bl[139] br[139] wl[147] vdd gnd cell_6t
Xbit_r148_c139 bl[139] br[139] wl[148] vdd gnd cell_6t
Xbit_r149_c139 bl[139] br[139] wl[149] vdd gnd cell_6t
Xbit_r150_c139 bl[139] br[139] wl[150] vdd gnd cell_6t
Xbit_r151_c139 bl[139] br[139] wl[151] vdd gnd cell_6t
Xbit_r152_c139 bl[139] br[139] wl[152] vdd gnd cell_6t
Xbit_r153_c139 bl[139] br[139] wl[153] vdd gnd cell_6t
Xbit_r154_c139 bl[139] br[139] wl[154] vdd gnd cell_6t
Xbit_r155_c139 bl[139] br[139] wl[155] vdd gnd cell_6t
Xbit_r156_c139 bl[139] br[139] wl[156] vdd gnd cell_6t
Xbit_r157_c139 bl[139] br[139] wl[157] vdd gnd cell_6t
Xbit_r158_c139 bl[139] br[139] wl[158] vdd gnd cell_6t
Xbit_r159_c139 bl[139] br[139] wl[159] vdd gnd cell_6t
Xbit_r160_c139 bl[139] br[139] wl[160] vdd gnd cell_6t
Xbit_r161_c139 bl[139] br[139] wl[161] vdd gnd cell_6t
Xbit_r162_c139 bl[139] br[139] wl[162] vdd gnd cell_6t
Xbit_r163_c139 bl[139] br[139] wl[163] vdd gnd cell_6t
Xbit_r164_c139 bl[139] br[139] wl[164] vdd gnd cell_6t
Xbit_r165_c139 bl[139] br[139] wl[165] vdd gnd cell_6t
Xbit_r166_c139 bl[139] br[139] wl[166] vdd gnd cell_6t
Xbit_r167_c139 bl[139] br[139] wl[167] vdd gnd cell_6t
Xbit_r168_c139 bl[139] br[139] wl[168] vdd gnd cell_6t
Xbit_r169_c139 bl[139] br[139] wl[169] vdd gnd cell_6t
Xbit_r170_c139 bl[139] br[139] wl[170] vdd gnd cell_6t
Xbit_r171_c139 bl[139] br[139] wl[171] vdd gnd cell_6t
Xbit_r172_c139 bl[139] br[139] wl[172] vdd gnd cell_6t
Xbit_r173_c139 bl[139] br[139] wl[173] vdd gnd cell_6t
Xbit_r174_c139 bl[139] br[139] wl[174] vdd gnd cell_6t
Xbit_r175_c139 bl[139] br[139] wl[175] vdd gnd cell_6t
Xbit_r176_c139 bl[139] br[139] wl[176] vdd gnd cell_6t
Xbit_r177_c139 bl[139] br[139] wl[177] vdd gnd cell_6t
Xbit_r178_c139 bl[139] br[139] wl[178] vdd gnd cell_6t
Xbit_r179_c139 bl[139] br[139] wl[179] vdd gnd cell_6t
Xbit_r180_c139 bl[139] br[139] wl[180] vdd gnd cell_6t
Xbit_r181_c139 bl[139] br[139] wl[181] vdd gnd cell_6t
Xbit_r182_c139 bl[139] br[139] wl[182] vdd gnd cell_6t
Xbit_r183_c139 bl[139] br[139] wl[183] vdd gnd cell_6t
Xbit_r184_c139 bl[139] br[139] wl[184] vdd gnd cell_6t
Xbit_r185_c139 bl[139] br[139] wl[185] vdd gnd cell_6t
Xbit_r186_c139 bl[139] br[139] wl[186] vdd gnd cell_6t
Xbit_r187_c139 bl[139] br[139] wl[187] vdd gnd cell_6t
Xbit_r188_c139 bl[139] br[139] wl[188] vdd gnd cell_6t
Xbit_r189_c139 bl[139] br[139] wl[189] vdd gnd cell_6t
Xbit_r190_c139 bl[139] br[139] wl[190] vdd gnd cell_6t
Xbit_r191_c139 bl[139] br[139] wl[191] vdd gnd cell_6t
Xbit_r192_c139 bl[139] br[139] wl[192] vdd gnd cell_6t
Xbit_r193_c139 bl[139] br[139] wl[193] vdd gnd cell_6t
Xbit_r194_c139 bl[139] br[139] wl[194] vdd gnd cell_6t
Xbit_r195_c139 bl[139] br[139] wl[195] vdd gnd cell_6t
Xbit_r196_c139 bl[139] br[139] wl[196] vdd gnd cell_6t
Xbit_r197_c139 bl[139] br[139] wl[197] vdd gnd cell_6t
Xbit_r198_c139 bl[139] br[139] wl[198] vdd gnd cell_6t
Xbit_r199_c139 bl[139] br[139] wl[199] vdd gnd cell_6t
Xbit_r200_c139 bl[139] br[139] wl[200] vdd gnd cell_6t
Xbit_r201_c139 bl[139] br[139] wl[201] vdd gnd cell_6t
Xbit_r202_c139 bl[139] br[139] wl[202] vdd gnd cell_6t
Xbit_r203_c139 bl[139] br[139] wl[203] vdd gnd cell_6t
Xbit_r204_c139 bl[139] br[139] wl[204] vdd gnd cell_6t
Xbit_r205_c139 bl[139] br[139] wl[205] vdd gnd cell_6t
Xbit_r206_c139 bl[139] br[139] wl[206] vdd gnd cell_6t
Xbit_r207_c139 bl[139] br[139] wl[207] vdd gnd cell_6t
Xbit_r208_c139 bl[139] br[139] wl[208] vdd gnd cell_6t
Xbit_r209_c139 bl[139] br[139] wl[209] vdd gnd cell_6t
Xbit_r210_c139 bl[139] br[139] wl[210] vdd gnd cell_6t
Xbit_r211_c139 bl[139] br[139] wl[211] vdd gnd cell_6t
Xbit_r212_c139 bl[139] br[139] wl[212] vdd gnd cell_6t
Xbit_r213_c139 bl[139] br[139] wl[213] vdd gnd cell_6t
Xbit_r214_c139 bl[139] br[139] wl[214] vdd gnd cell_6t
Xbit_r215_c139 bl[139] br[139] wl[215] vdd gnd cell_6t
Xbit_r216_c139 bl[139] br[139] wl[216] vdd gnd cell_6t
Xbit_r217_c139 bl[139] br[139] wl[217] vdd gnd cell_6t
Xbit_r218_c139 bl[139] br[139] wl[218] vdd gnd cell_6t
Xbit_r219_c139 bl[139] br[139] wl[219] vdd gnd cell_6t
Xbit_r220_c139 bl[139] br[139] wl[220] vdd gnd cell_6t
Xbit_r221_c139 bl[139] br[139] wl[221] vdd gnd cell_6t
Xbit_r222_c139 bl[139] br[139] wl[222] vdd gnd cell_6t
Xbit_r223_c139 bl[139] br[139] wl[223] vdd gnd cell_6t
Xbit_r224_c139 bl[139] br[139] wl[224] vdd gnd cell_6t
Xbit_r225_c139 bl[139] br[139] wl[225] vdd gnd cell_6t
Xbit_r226_c139 bl[139] br[139] wl[226] vdd gnd cell_6t
Xbit_r227_c139 bl[139] br[139] wl[227] vdd gnd cell_6t
Xbit_r228_c139 bl[139] br[139] wl[228] vdd gnd cell_6t
Xbit_r229_c139 bl[139] br[139] wl[229] vdd gnd cell_6t
Xbit_r230_c139 bl[139] br[139] wl[230] vdd gnd cell_6t
Xbit_r231_c139 bl[139] br[139] wl[231] vdd gnd cell_6t
Xbit_r232_c139 bl[139] br[139] wl[232] vdd gnd cell_6t
Xbit_r233_c139 bl[139] br[139] wl[233] vdd gnd cell_6t
Xbit_r234_c139 bl[139] br[139] wl[234] vdd gnd cell_6t
Xbit_r235_c139 bl[139] br[139] wl[235] vdd gnd cell_6t
Xbit_r236_c139 bl[139] br[139] wl[236] vdd gnd cell_6t
Xbit_r237_c139 bl[139] br[139] wl[237] vdd gnd cell_6t
Xbit_r238_c139 bl[139] br[139] wl[238] vdd gnd cell_6t
Xbit_r239_c139 bl[139] br[139] wl[239] vdd gnd cell_6t
Xbit_r240_c139 bl[139] br[139] wl[240] vdd gnd cell_6t
Xbit_r241_c139 bl[139] br[139] wl[241] vdd gnd cell_6t
Xbit_r242_c139 bl[139] br[139] wl[242] vdd gnd cell_6t
Xbit_r243_c139 bl[139] br[139] wl[243] vdd gnd cell_6t
Xbit_r244_c139 bl[139] br[139] wl[244] vdd gnd cell_6t
Xbit_r245_c139 bl[139] br[139] wl[245] vdd gnd cell_6t
Xbit_r246_c139 bl[139] br[139] wl[246] vdd gnd cell_6t
Xbit_r247_c139 bl[139] br[139] wl[247] vdd gnd cell_6t
Xbit_r248_c139 bl[139] br[139] wl[248] vdd gnd cell_6t
Xbit_r249_c139 bl[139] br[139] wl[249] vdd gnd cell_6t
Xbit_r250_c139 bl[139] br[139] wl[250] vdd gnd cell_6t
Xbit_r251_c139 bl[139] br[139] wl[251] vdd gnd cell_6t
Xbit_r252_c139 bl[139] br[139] wl[252] vdd gnd cell_6t
Xbit_r253_c139 bl[139] br[139] wl[253] vdd gnd cell_6t
Xbit_r254_c139 bl[139] br[139] wl[254] vdd gnd cell_6t
Xbit_r255_c139 bl[139] br[139] wl[255] vdd gnd cell_6t
Xbit_r0_c140 bl[140] br[140] wl[0] vdd gnd cell_6t
Xbit_r1_c140 bl[140] br[140] wl[1] vdd gnd cell_6t
Xbit_r2_c140 bl[140] br[140] wl[2] vdd gnd cell_6t
Xbit_r3_c140 bl[140] br[140] wl[3] vdd gnd cell_6t
Xbit_r4_c140 bl[140] br[140] wl[4] vdd gnd cell_6t
Xbit_r5_c140 bl[140] br[140] wl[5] vdd gnd cell_6t
Xbit_r6_c140 bl[140] br[140] wl[6] vdd gnd cell_6t
Xbit_r7_c140 bl[140] br[140] wl[7] vdd gnd cell_6t
Xbit_r8_c140 bl[140] br[140] wl[8] vdd gnd cell_6t
Xbit_r9_c140 bl[140] br[140] wl[9] vdd gnd cell_6t
Xbit_r10_c140 bl[140] br[140] wl[10] vdd gnd cell_6t
Xbit_r11_c140 bl[140] br[140] wl[11] vdd gnd cell_6t
Xbit_r12_c140 bl[140] br[140] wl[12] vdd gnd cell_6t
Xbit_r13_c140 bl[140] br[140] wl[13] vdd gnd cell_6t
Xbit_r14_c140 bl[140] br[140] wl[14] vdd gnd cell_6t
Xbit_r15_c140 bl[140] br[140] wl[15] vdd gnd cell_6t
Xbit_r16_c140 bl[140] br[140] wl[16] vdd gnd cell_6t
Xbit_r17_c140 bl[140] br[140] wl[17] vdd gnd cell_6t
Xbit_r18_c140 bl[140] br[140] wl[18] vdd gnd cell_6t
Xbit_r19_c140 bl[140] br[140] wl[19] vdd gnd cell_6t
Xbit_r20_c140 bl[140] br[140] wl[20] vdd gnd cell_6t
Xbit_r21_c140 bl[140] br[140] wl[21] vdd gnd cell_6t
Xbit_r22_c140 bl[140] br[140] wl[22] vdd gnd cell_6t
Xbit_r23_c140 bl[140] br[140] wl[23] vdd gnd cell_6t
Xbit_r24_c140 bl[140] br[140] wl[24] vdd gnd cell_6t
Xbit_r25_c140 bl[140] br[140] wl[25] vdd gnd cell_6t
Xbit_r26_c140 bl[140] br[140] wl[26] vdd gnd cell_6t
Xbit_r27_c140 bl[140] br[140] wl[27] vdd gnd cell_6t
Xbit_r28_c140 bl[140] br[140] wl[28] vdd gnd cell_6t
Xbit_r29_c140 bl[140] br[140] wl[29] vdd gnd cell_6t
Xbit_r30_c140 bl[140] br[140] wl[30] vdd gnd cell_6t
Xbit_r31_c140 bl[140] br[140] wl[31] vdd gnd cell_6t
Xbit_r32_c140 bl[140] br[140] wl[32] vdd gnd cell_6t
Xbit_r33_c140 bl[140] br[140] wl[33] vdd gnd cell_6t
Xbit_r34_c140 bl[140] br[140] wl[34] vdd gnd cell_6t
Xbit_r35_c140 bl[140] br[140] wl[35] vdd gnd cell_6t
Xbit_r36_c140 bl[140] br[140] wl[36] vdd gnd cell_6t
Xbit_r37_c140 bl[140] br[140] wl[37] vdd gnd cell_6t
Xbit_r38_c140 bl[140] br[140] wl[38] vdd gnd cell_6t
Xbit_r39_c140 bl[140] br[140] wl[39] vdd gnd cell_6t
Xbit_r40_c140 bl[140] br[140] wl[40] vdd gnd cell_6t
Xbit_r41_c140 bl[140] br[140] wl[41] vdd gnd cell_6t
Xbit_r42_c140 bl[140] br[140] wl[42] vdd gnd cell_6t
Xbit_r43_c140 bl[140] br[140] wl[43] vdd gnd cell_6t
Xbit_r44_c140 bl[140] br[140] wl[44] vdd gnd cell_6t
Xbit_r45_c140 bl[140] br[140] wl[45] vdd gnd cell_6t
Xbit_r46_c140 bl[140] br[140] wl[46] vdd gnd cell_6t
Xbit_r47_c140 bl[140] br[140] wl[47] vdd gnd cell_6t
Xbit_r48_c140 bl[140] br[140] wl[48] vdd gnd cell_6t
Xbit_r49_c140 bl[140] br[140] wl[49] vdd gnd cell_6t
Xbit_r50_c140 bl[140] br[140] wl[50] vdd gnd cell_6t
Xbit_r51_c140 bl[140] br[140] wl[51] vdd gnd cell_6t
Xbit_r52_c140 bl[140] br[140] wl[52] vdd gnd cell_6t
Xbit_r53_c140 bl[140] br[140] wl[53] vdd gnd cell_6t
Xbit_r54_c140 bl[140] br[140] wl[54] vdd gnd cell_6t
Xbit_r55_c140 bl[140] br[140] wl[55] vdd gnd cell_6t
Xbit_r56_c140 bl[140] br[140] wl[56] vdd gnd cell_6t
Xbit_r57_c140 bl[140] br[140] wl[57] vdd gnd cell_6t
Xbit_r58_c140 bl[140] br[140] wl[58] vdd gnd cell_6t
Xbit_r59_c140 bl[140] br[140] wl[59] vdd gnd cell_6t
Xbit_r60_c140 bl[140] br[140] wl[60] vdd gnd cell_6t
Xbit_r61_c140 bl[140] br[140] wl[61] vdd gnd cell_6t
Xbit_r62_c140 bl[140] br[140] wl[62] vdd gnd cell_6t
Xbit_r63_c140 bl[140] br[140] wl[63] vdd gnd cell_6t
Xbit_r64_c140 bl[140] br[140] wl[64] vdd gnd cell_6t
Xbit_r65_c140 bl[140] br[140] wl[65] vdd gnd cell_6t
Xbit_r66_c140 bl[140] br[140] wl[66] vdd gnd cell_6t
Xbit_r67_c140 bl[140] br[140] wl[67] vdd gnd cell_6t
Xbit_r68_c140 bl[140] br[140] wl[68] vdd gnd cell_6t
Xbit_r69_c140 bl[140] br[140] wl[69] vdd gnd cell_6t
Xbit_r70_c140 bl[140] br[140] wl[70] vdd gnd cell_6t
Xbit_r71_c140 bl[140] br[140] wl[71] vdd gnd cell_6t
Xbit_r72_c140 bl[140] br[140] wl[72] vdd gnd cell_6t
Xbit_r73_c140 bl[140] br[140] wl[73] vdd gnd cell_6t
Xbit_r74_c140 bl[140] br[140] wl[74] vdd gnd cell_6t
Xbit_r75_c140 bl[140] br[140] wl[75] vdd gnd cell_6t
Xbit_r76_c140 bl[140] br[140] wl[76] vdd gnd cell_6t
Xbit_r77_c140 bl[140] br[140] wl[77] vdd gnd cell_6t
Xbit_r78_c140 bl[140] br[140] wl[78] vdd gnd cell_6t
Xbit_r79_c140 bl[140] br[140] wl[79] vdd gnd cell_6t
Xbit_r80_c140 bl[140] br[140] wl[80] vdd gnd cell_6t
Xbit_r81_c140 bl[140] br[140] wl[81] vdd gnd cell_6t
Xbit_r82_c140 bl[140] br[140] wl[82] vdd gnd cell_6t
Xbit_r83_c140 bl[140] br[140] wl[83] vdd gnd cell_6t
Xbit_r84_c140 bl[140] br[140] wl[84] vdd gnd cell_6t
Xbit_r85_c140 bl[140] br[140] wl[85] vdd gnd cell_6t
Xbit_r86_c140 bl[140] br[140] wl[86] vdd gnd cell_6t
Xbit_r87_c140 bl[140] br[140] wl[87] vdd gnd cell_6t
Xbit_r88_c140 bl[140] br[140] wl[88] vdd gnd cell_6t
Xbit_r89_c140 bl[140] br[140] wl[89] vdd gnd cell_6t
Xbit_r90_c140 bl[140] br[140] wl[90] vdd gnd cell_6t
Xbit_r91_c140 bl[140] br[140] wl[91] vdd gnd cell_6t
Xbit_r92_c140 bl[140] br[140] wl[92] vdd gnd cell_6t
Xbit_r93_c140 bl[140] br[140] wl[93] vdd gnd cell_6t
Xbit_r94_c140 bl[140] br[140] wl[94] vdd gnd cell_6t
Xbit_r95_c140 bl[140] br[140] wl[95] vdd gnd cell_6t
Xbit_r96_c140 bl[140] br[140] wl[96] vdd gnd cell_6t
Xbit_r97_c140 bl[140] br[140] wl[97] vdd gnd cell_6t
Xbit_r98_c140 bl[140] br[140] wl[98] vdd gnd cell_6t
Xbit_r99_c140 bl[140] br[140] wl[99] vdd gnd cell_6t
Xbit_r100_c140 bl[140] br[140] wl[100] vdd gnd cell_6t
Xbit_r101_c140 bl[140] br[140] wl[101] vdd gnd cell_6t
Xbit_r102_c140 bl[140] br[140] wl[102] vdd gnd cell_6t
Xbit_r103_c140 bl[140] br[140] wl[103] vdd gnd cell_6t
Xbit_r104_c140 bl[140] br[140] wl[104] vdd gnd cell_6t
Xbit_r105_c140 bl[140] br[140] wl[105] vdd gnd cell_6t
Xbit_r106_c140 bl[140] br[140] wl[106] vdd gnd cell_6t
Xbit_r107_c140 bl[140] br[140] wl[107] vdd gnd cell_6t
Xbit_r108_c140 bl[140] br[140] wl[108] vdd gnd cell_6t
Xbit_r109_c140 bl[140] br[140] wl[109] vdd gnd cell_6t
Xbit_r110_c140 bl[140] br[140] wl[110] vdd gnd cell_6t
Xbit_r111_c140 bl[140] br[140] wl[111] vdd gnd cell_6t
Xbit_r112_c140 bl[140] br[140] wl[112] vdd gnd cell_6t
Xbit_r113_c140 bl[140] br[140] wl[113] vdd gnd cell_6t
Xbit_r114_c140 bl[140] br[140] wl[114] vdd gnd cell_6t
Xbit_r115_c140 bl[140] br[140] wl[115] vdd gnd cell_6t
Xbit_r116_c140 bl[140] br[140] wl[116] vdd gnd cell_6t
Xbit_r117_c140 bl[140] br[140] wl[117] vdd gnd cell_6t
Xbit_r118_c140 bl[140] br[140] wl[118] vdd gnd cell_6t
Xbit_r119_c140 bl[140] br[140] wl[119] vdd gnd cell_6t
Xbit_r120_c140 bl[140] br[140] wl[120] vdd gnd cell_6t
Xbit_r121_c140 bl[140] br[140] wl[121] vdd gnd cell_6t
Xbit_r122_c140 bl[140] br[140] wl[122] vdd gnd cell_6t
Xbit_r123_c140 bl[140] br[140] wl[123] vdd gnd cell_6t
Xbit_r124_c140 bl[140] br[140] wl[124] vdd gnd cell_6t
Xbit_r125_c140 bl[140] br[140] wl[125] vdd gnd cell_6t
Xbit_r126_c140 bl[140] br[140] wl[126] vdd gnd cell_6t
Xbit_r127_c140 bl[140] br[140] wl[127] vdd gnd cell_6t
Xbit_r128_c140 bl[140] br[140] wl[128] vdd gnd cell_6t
Xbit_r129_c140 bl[140] br[140] wl[129] vdd gnd cell_6t
Xbit_r130_c140 bl[140] br[140] wl[130] vdd gnd cell_6t
Xbit_r131_c140 bl[140] br[140] wl[131] vdd gnd cell_6t
Xbit_r132_c140 bl[140] br[140] wl[132] vdd gnd cell_6t
Xbit_r133_c140 bl[140] br[140] wl[133] vdd gnd cell_6t
Xbit_r134_c140 bl[140] br[140] wl[134] vdd gnd cell_6t
Xbit_r135_c140 bl[140] br[140] wl[135] vdd gnd cell_6t
Xbit_r136_c140 bl[140] br[140] wl[136] vdd gnd cell_6t
Xbit_r137_c140 bl[140] br[140] wl[137] vdd gnd cell_6t
Xbit_r138_c140 bl[140] br[140] wl[138] vdd gnd cell_6t
Xbit_r139_c140 bl[140] br[140] wl[139] vdd gnd cell_6t
Xbit_r140_c140 bl[140] br[140] wl[140] vdd gnd cell_6t
Xbit_r141_c140 bl[140] br[140] wl[141] vdd gnd cell_6t
Xbit_r142_c140 bl[140] br[140] wl[142] vdd gnd cell_6t
Xbit_r143_c140 bl[140] br[140] wl[143] vdd gnd cell_6t
Xbit_r144_c140 bl[140] br[140] wl[144] vdd gnd cell_6t
Xbit_r145_c140 bl[140] br[140] wl[145] vdd gnd cell_6t
Xbit_r146_c140 bl[140] br[140] wl[146] vdd gnd cell_6t
Xbit_r147_c140 bl[140] br[140] wl[147] vdd gnd cell_6t
Xbit_r148_c140 bl[140] br[140] wl[148] vdd gnd cell_6t
Xbit_r149_c140 bl[140] br[140] wl[149] vdd gnd cell_6t
Xbit_r150_c140 bl[140] br[140] wl[150] vdd gnd cell_6t
Xbit_r151_c140 bl[140] br[140] wl[151] vdd gnd cell_6t
Xbit_r152_c140 bl[140] br[140] wl[152] vdd gnd cell_6t
Xbit_r153_c140 bl[140] br[140] wl[153] vdd gnd cell_6t
Xbit_r154_c140 bl[140] br[140] wl[154] vdd gnd cell_6t
Xbit_r155_c140 bl[140] br[140] wl[155] vdd gnd cell_6t
Xbit_r156_c140 bl[140] br[140] wl[156] vdd gnd cell_6t
Xbit_r157_c140 bl[140] br[140] wl[157] vdd gnd cell_6t
Xbit_r158_c140 bl[140] br[140] wl[158] vdd gnd cell_6t
Xbit_r159_c140 bl[140] br[140] wl[159] vdd gnd cell_6t
Xbit_r160_c140 bl[140] br[140] wl[160] vdd gnd cell_6t
Xbit_r161_c140 bl[140] br[140] wl[161] vdd gnd cell_6t
Xbit_r162_c140 bl[140] br[140] wl[162] vdd gnd cell_6t
Xbit_r163_c140 bl[140] br[140] wl[163] vdd gnd cell_6t
Xbit_r164_c140 bl[140] br[140] wl[164] vdd gnd cell_6t
Xbit_r165_c140 bl[140] br[140] wl[165] vdd gnd cell_6t
Xbit_r166_c140 bl[140] br[140] wl[166] vdd gnd cell_6t
Xbit_r167_c140 bl[140] br[140] wl[167] vdd gnd cell_6t
Xbit_r168_c140 bl[140] br[140] wl[168] vdd gnd cell_6t
Xbit_r169_c140 bl[140] br[140] wl[169] vdd gnd cell_6t
Xbit_r170_c140 bl[140] br[140] wl[170] vdd gnd cell_6t
Xbit_r171_c140 bl[140] br[140] wl[171] vdd gnd cell_6t
Xbit_r172_c140 bl[140] br[140] wl[172] vdd gnd cell_6t
Xbit_r173_c140 bl[140] br[140] wl[173] vdd gnd cell_6t
Xbit_r174_c140 bl[140] br[140] wl[174] vdd gnd cell_6t
Xbit_r175_c140 bl[140] br[140] wl[175] vdd gnd cell_6t
Xbit_r176_c140 bl[140] br[140] wl[176] vdd gnd cell_6t
Xbit_r177_c140 bl[140] br[140] wl[177] vdd gnd cell_6t
Xbit_r178_c140 bl[140] br[140] wl[178] vdd gnd cell_6t
Xbit_r179_c140 bl[140] br[140] wl[179] vdd gnd cell_6t
Xbit_r180_c140 bl[140] br[140] wl[180] vdd gnd cell_6t
Xbit_r181_c140 bl[140] br[140] wl[181] vdd gnd cell_6t
Xbit_r182_c140 bl[140] br[140] wl[182] vdd gnd cell_6t
Xbit_r183_c140 bl[140] br[140] wl[183] vdd gnd cell_6t
Xbit_r184_c140 bl[140] br[140] wl[184] vdd gnd cell_6t
Xbit_r185_c140 bl[140] br[140] wl[185] vdd gnd cell_6t
Xbit_r186_c140 bl[140] br[140] wl[186] vdd gnd cell_6t
Xbit_r187_c140 bl[140] br[140] wl[187] vdd gnd cell_6t
Xbit_r188_c140 bl[140] br[140] wl[188] vdd gnd cell_6t
Xbit_r189_c140 bl[140] br[140] wl[189] vdd gnd cell_6t
Xbit_r190_c140 bl[140] br[140] wl[190] vdd gnd cell_6t
Xbit_r191_c140 bl[140] br[140] wl[191] vdd gnd cell_6t
Xbit_r192_c140 bl[140] br[140] wl[192] vdd gnd cell_6t
Xbit_r193_c140 bl[140] br[140] wl[193] vdd gnd cell_6t
Xbit_r194_c140 bl[140] br[140] wl[194] vdd gnd cell_6t
Xbit_r195_c140 bl[140] br[140] wl[195] vdd gnd cell_6t
Xbit_r196_c140 bl[140] br[140] wl[196] vdd gnd cell_6t
Xbit_r197_c140 bl[140] br[140] wl[197] vdd gnd cell_6t
Xbit_r198_c140 bl[140] br[140] wl[198] vdd gnd cell_6t
Xbit_r199_c140 bl[140] br[140] wl[199] vdd gnd cell_6t
Xbit_r200_c140 bl[140] br[140] wl[200] vdd gnd cell_6t
Xbit_r201_c140 bl[140] br[140] wl[201] vdd gnd cell_6t
Xbit_r202_c140 bl[140] br[140] wl[202] vdd gnd cell_6t
Xbit_r203_c140 bl[140] br[140] wl[203] vdd gnd cell_6t
Xbit_r204_c140 bl[140] br[140] wl[204] vdd gnd cell_6t
Xbit_r205_c140 bl[140] br[140] wl[205] vdd gnd cell_6t
Xbit_r206_c140 bl[140] br[140] wl[206] vdd gnd cell_6t
Xbit_r207_c140 bl[140] br[140] wl[207] vdd gnd cell_6t
Xbit_r208_c140 bl[140] br[140] wl[208] vdd gnd cell_6t
Xbit_r209_c140 bl[140] br[140] wl[209] vdd gnd cell_6t
Xbit_r210_c140 bl[140] br[140] wl[210] vdd gnd cell_6t
Xbit_r211_c140 bl[140] br[140] wl[211] vdd gnd cell_6t
Xbit_r212_c140 bl[140] br[140] wl[212] vdd gnd cell_6t
Xbit_r213_c140 bl[140] br[140] wl[213] vdd gnd cell_6t
Xbit_r214_c140 bl[140] br[140] wl[214] vdd gnd cell_6t
Xbit_r215_c140 bl[140] br[140] wl[215] vdd gnd cell_6t
Xbit_r216_c140 bl[140] br[140] wl[216] vdd gnd cell_6t
Xbit_r217_c140 bl[140] br[140] wl[217] vdd gnd cell_6t
Xbit_r218_c140 bl[140] br[140] wl[218] vdd gnd cell_6t
Xbit_r219_c140 bl[140] br[140] wl[219] vdd gnd cell_6t
Xbit_r220_c140 bl[140] br[140] wl[220] vdd gnd cell_6t
Xbit_r221_c140 bl[140] br[140] wl[221] vdd gnd cell_6t
Xbit_r222_c140 bl[140] br[140] wl[222] vdd gnd cell_6t
Xbit_r223_c140 bl[140] br[140] wl[223] vdd gnd cell_6t
Xbit_r224_c140 bl[140] br[140] wl[224] vdd gnd cell_6t
Xbit_r225_c140 bl[140] br[140] wl[225] vdd gnd cell_6t
Xbit_r226_c140 bl[140] br[140] wl[226] vdd gnd cell_6t
Xbit_r227_c140 bl[140] br[140] wl[227] vdd gnd cell_6t
Xbit_r228_c140 bl[140] br[140] wl[228] vdd gnd cell_6t
Xbit_r229_c140 bl[140] br[140] wl[229] vdd gnd cell_6t
Xbit_r230_c140 bl[140] br[140] wl[230] vdd gnd cell_6t
Xbit_r231_c140 bl[140] br[140] wl[231] vdd gnd cell_6t
Xbit_r232_c140 bl[140] br[140] wl[232] vdd gnd cell_6t
Xbit_r233_c140 bl[140] br[140] wl[233] vdd gnd cell_6t
Xbit_r234_c140 bl[140] br[140] wl[234] vdd gnd cell_6t
Xbit_r235_c140 bl[140] br[140] wl[235] vdd gnd cell_6t
Xbit_r236_c140 bl[140] br[140] wl[236] vdd gnd cell_6t
Xbit_r237_c140 bl[140] br[140] wl[237] vdd gnd cell_6t
Xbit_r238_c140 bl[140] br[140] wl[238] vdd gnd cell_6t
Xbit_r239_c140 bl[140] br[140] wl[239] vdd gnd cell_6t
Xbit_r240_c140 bl[140] br[140] wl[240] vdd gnd cell_6t
Xbit_r241_c140 bl[140] br[140] wl[241] vdd gnd cell_6t
Xbit_r242_c140 bl[140] br[140] wl[242] vdd gnd cell_6t
Xbit_r243_c140 bl[140] br[140] wl[243] vdd gnd cell_6t
Xbit_r244_c140 bl[140] br[140] wl[244] vdd gnd cell_6t
Xbit_r245_c140 bl[140] br[140] wl[245] vdd gnd cell_6t
Xbit_r246_c140 bl[140] br[140] wl[246] vdd gnd cell_6t
Xbit_r247_c140 bl[140] br[140] wl[247] vdd gnd cell_6t
Xbit_r248_c140 bl[140] br[140] wl[248] vdd gnd cell_6t
Xbit_r249_c140 bl[140] br[140] wl[249] vdd gnd cell_6t
Xbit_r250_c140 bl[140] br[140] wl[250] vdd gnd cell_6t
Xbit_r251_c140 bl[140] br[140] wl[251] vdd gnd cell_6t
Xbit_r252_c140 bl[140] br[140] wl[252] vdd gnd cell_6t
Xbit_r253_c140 bl[140] br[140] wl[253] vdd gnd cell_6t
Xbit_r254_c140 bl[140] br[140] wl[254] vdd gnd cell_6t
Xbit_r255_c140 bl[140] br[140] wl[255] vdd gnd cell_6t
Xbit_r0_c141 bl[141] br[141] wl[0] vdd gnd cell_6t
Xbit_r1_c141 bl[141] br[141] wl[1] vdd gnd cell_6t
Xbit_r2_c141 bl[141] br[141] wl[2] vdd gnd cell_6t
Xbit_r3_c141 bl[141] br[141] wl[3] vdd gnd cell_6t
Xbit_r4_c141 bl[141] br[141] wl[4] vdd gnd cell_6t
Xbit_r5_c141 bl[141] br[141] wl[5] vdd gnd cell_6t
Xbit_r6_c141 bl[141] br[141] wl[6] vdd gnd cell_6t
Xbit_r7_c141 bl[141] br[141] wl[7] vdd gnd cell_6t
Xbit_r8_c141 bl[141] br[141] wl[8] vdd gnd cell_6t
Xbit_r9_c141 bl[141] br[141] wl[9] vdd gnd cell_6t
Xbit_r10_c141 bl[141] br[141] wl[10] vdd gnd cell_6t
Xbit_r11_c141 bl[141] br[141] wl[11] vdd gnd cell_6t
Xbit_r12_c141 bl[141] br[141] wl[12] vdd gnd cell_6t
Xbit_r13_c141 bl[141] br[141] wl[13] vdd gnd cell_6t
Xbit_r14_c141 bl[141] br[141] wl[14] vdd gnd cell_6t
Xbit_r15_c141 bl[141] br[141] wl[15] vdd gnd cell_6t
Xbit_r16_c141 bl[141] br[141] wl[16] vdd gnd cell_6t
Xbit_r17_c141 bl[141] br[141] wl[17] vdd gnd cell_6t
Xbit_r18_c141 bl[141] br[141] wl[18] vdd gnd cell_6t
Xbit_r19_c141 bl[141] br[141] wl[19] vdd gnd cell_6t
Xbit_r20_c141 bl[141] br[141] wl[20] vdd gnd cell_6t
Xbit_r21_c141 bl[141] br[141] wl[21] vdd gnd cell_6t
Xbit_r22_c141 bl[141] br[141] wl[22] vdd gnd cell_6t
Xbit_r23_c141 bl[141] br[141] wl[23] vdd gnd cell_6t
Xbit_r24_c141 bl[141] br[141] wl[24] vdd gnd cell_6t
Xbit_r25_c141 bl[141] br[141] wl[25] vdd gnd cell_6t
Xbit_r26_c141 bl[141] br[141] wl[26] vdd gnd cell_6t
Xbit_r27_c141 bl[141] br[141] wl[27] vdd gnd cell_6t
Xbit_r28_c141 bl[141] br[141] wl[28] vdd gnd cell_6t
Xbit_r29_c141 bl[141] br[141] wl[29] vdd gnd cell_6t
Xbit_r30_c141 bl[141] br[141] wl[30] vdd gnd cell_6t
Xbit_r31_c141 bl[141] br[141] wl[31] vdd gnd cell_6t
Xbit_r32_c141 bl[141] br[141] wl[32] vdd gnd cell_6t
Xbit_r33_c141 bl[141] br[141] wl[33] vdd gnd cell_6t
Xbit_r34_c141 bl[141] br[141] wl[34] vdd gnd cell_6t
Xbit_r35_c141 bl[141] br[141] wl[35] vdd gnd cell_6t
Xbit_r36_c141 bl[141] br[141] wl[36] vdd gnd cell_6t
Xbit_r37_c141 bl[141] br[141] wl[37] vdd gnd cell_6t
Xbit_r38_c141 bl[141] br[141] wl[38] vdd gnd cell_6t
Xbit_r39_c141 bl[141] br[141] wl[39] vdd gnd cell_6t
Xbit_r40_c141 bl[141] br[141] wl[40] vdd gnd cell_6t
Xbit_r41_c141 bl[141] br[141] wl[41] vdd gnd cell_6t
Xbit_r42_c141 bl[141] br[141] wl[42] vdd gnd cell_6t
Xbit_r43_c141 bl[141] br[141] wl[43] vdd gnd cell_6t
Xbit_r44_c141 bl[141] br[141] wl[44] vdd gnd cell_6t
Xbit_r45_c141 bl[141] br[141] wl[45] vdd gnd cell_6t
Xbit_r46_c141 bl[141] br[141] wl[46] vdd gnd cell_6t
Xbit_r47_c141 bl[141] br[141] wl[47] vdd gnd cell_6t
Xbit_r48_c141 bl[141] br[141] wl[48] vdd gnd cell_6t
Xbit_r49_c141 bl[141] br[141] wl[49] vdd gnd cell_6t
Xbit_r50_c141 bl[141] br[141] wl[50] vdd gnd cell_6t
Xbit_r51_c141 bl[141] br[141] wl[51] vdd gnd cell_6t
Xbit_r52_c141 bl[141] br[141] wl[52] vdd gnd cell_6t
Xbit_r53_c141 bl[141] br[141] wl[53] vdd gnd cell_6t
Xbit_r54_c141 bl[141] br[141] wl[54] vdd gnd cell_6t
Xbit_r55_c141 bl[141] br[141] wl[55] vdd gnd cell_6t
Xbit_r56_c141 bl[141] br[141] wl[56] vdd gnd cell_6t
Xbit_r57_c141 bl[141] br[141] wl[57] vdd gnd cell_6t
Xbit_r58_c141 bl[141] br[141] wl[58] vdd gnd cell_6t
Xbit_r59_c141 bl[141] br[141] wl[59] vdd gnd cell_6t
Xbit_r60_c141 bl[141] br[141] wl[60] vdd gnd cell_6t
Xbit_r61_c141 bl[141] br[141] wl[61] vdd gnd cell_6t
Xbit_r62_c141 bl[141] br[141] wl[62] vdd gnd cell_6t
Xbit_r63_c141 bl[141] br[141] wl[63] vdd gnd cell_6t
Xbit_r64_c141 bl[141] br[141] wl[64] vdd gnd cell_6t
Xbit_r65_c141 bl[141] br[141] wl[65] vdd gnd cell_6t
Xbit_r66_c141 bl[141] br[141] wl[66] vdd gnd cell_6t
Xbit_r67_c141 bl[141] br[141] wl[67] vdd gnd cell_6t
Xbit_r68_c141 bl[141] br[141] wl[68] vdd gnd cell_6t
Xbit_r69_c141 bl[141] br[141] wl[69] vdd gnd cell_6t
Xbit_r70_c141 bl[141] br[141] wl[70] vdd gnd cell_6t
Xbit_r71_c141 bl[141] br[141] wl[71] vdd gnd cell_6t
Xbit_r72_c141 bl[141] br[141] wl[72] vdd gnd cell_6t
Xbit_r73_c141 bl[141] br[141] wl[73] vdd gnd cell_6t
Xbit_r74_c141 bl[141] br[141] wl[74] vdd gnd cell_6t
Xbit_r75_c141 bl[141] br[141] wl[75] vdd gnd cell_6t
Xbit_r76_c141 bl[141] br[141] wl[76] vdd gnd cell_6t
Xbit_r77_c141 bl[141] br[141] wl[77] vdd gnd cell_6t
Xbit_r78_c141 bl[141] br[141] wl[78] vdd gnd cell_6t
Xbit_r79_c141 bl[141] br[141] wl[79] vdd gnd cell_6t
Xbit_r80_c141 bl[141] br[141] wl[80] vdd gnd cell_6t
Xbit_r81_c141 bl[141] br[141] wl[81] vdd gnd cell_6t
Xbit_r82_c141 bl[141] br[141] wl[82] vdd gnd cell_6t
Xbit_r83_c141 bl[141] br[141] wl[83] vdd gnd cell_6t
Xbit_r84_c141 bl[141] br[141] wl[84] vdd gnd cell_6t
Xbit_r85_c141 bl[141] br[141] wl[85] vdd gnd cell_6t
Xbit_r86_c141 bl[141] br[141] wl[86] vdd gnd cell_6t
Xbit_r87_c141 bl[141] br[141] wl[87] vdd gnd cell_6t
Xbit_r88_c141 bl[141] br[141] wl[88] vdd gnd cell_6t
Xbit_r89_c141 bl[141] br[141] wl[89] vdd gnd cell_6t
Xbit_r90_c141 bl[141] br[141] wl[90] vdd gnd cell_6t
Xbit_r91_c141 bl[141] br[141] wl[91] vdd gnd cell_6t
Xbit_r92_c141 bl[141] br[141] wl[92] vdd gnd cell_6t
Xbit_r93_c141 bl[141] br[141] wl[93] vdd gnd cell_6t
Xbit_r94_c141 bl[141] br[141] wl[94] vdd gnd cell_6t
Xbit_r95_c141 bl[141] br[141] wl[95] vdd gnd cell_6t
Xbit_r96_c141 bl[141] br[141] wl[96] vdd gnd cell_6t
Xbit_r97_c141 bl[141] br[141] wl[97] vdd gnd cell_6t
Xbit_r98_c141 bl[141] br[141] wl[98] vdd gnd cell_6t
Xbit_r99_c141 bl[141] br[141] wl[99] vdd gnd cell_6t
Xbit_r100_c141 bl[141] br[141] wl[100] vdd gnd cell_6t
Xbit_r101_c141 bl[141] br[141] wl[101] vdd gnd cell_6t
Xbit_r102_c141 bl[141] br[141] wl[102] vdd gnd cell_6t
Xbit_r103_c141 bl[141] br[141] wl[103] vdd gnd cell_6t
Xbit_r104_c141 bl[141] br[141] wl[104] vdd gnd cell_6t
Xbit_r105_c141 bl[141] br[141] wl[105] vdd gnd cell_6t
Xbit_r106_c141 bl[141] br[141] wl[106] vdd gnd cell_6t
Xbit_r107_c141 bl[141] br[141] wl[107] vdd gnd cell_6t
Xbit_r108_c141 bl[141] br[141] wl[108] vdd gnd cell_6t
Xbit_r109_c141 bl[141] br[141] wl[109] vdd gnd cell_6t
Xbit_r110_c141 bl[141] br[141] wl[110] vdd gnd cell_6t
Xbit_r111_c141 bl[141] br[141] wl[111] vdd gnd cell_6t
Xbit_r112_c141 bl[141] br[141] wl[112] vdd gnd cell_6t
Xbit_r113_c141 bl[141] br[141] wl[113] vdd gnd cell_6t
Xbit_r114_c141 bl[141] br[141] wl[114] vdd gnd cell_6t
Xbit_r115_c141 bl[141] br[141] wl[115] vdd gnd cell_6t
Xbit_r116_c141 bl[141] br[141] wl[116] vdd gnd cell_6t
Xbit_r117_c141 bl[141] br[141] wl[117] vdd gnd cell_6t
Xbit_r118_c141 bl[141] br[141] wl[118] vdd gnd cell_6t
Xbit_r119_c141 bl[141] br[141] wl[119] vdd gnd cell_6t
Xbit_r120_c141 bl[141] br[141] wl[120] vdd gnd cell_6t
Xbit_r121_c141 bl[141] br[141] wl[121] vdd gnd cell_6t
Xbit_r122_c141 bl[141] br[141] wl[122] vdd gnd cell_6t
Xbit_r123_c141 bl[141] br[141] wl[123] vdd gnd cell_6t
Xbit_r124_c141 bl[141] br[141] wl[124] vdd gnd cell_6t
Xbit_r125_c141 bl[141] br[141] wl[125] vdd gnd cell_6t
Xbit_r126_c141 bl[141] br[141] wl[126] vdd gnd cell_6t
Xbit_r127_c141 bl[141] br[141] wl[127] vdd gnd cell_6t
Xbit_r128_c141 bl[141] br[141] wl[128] vdd gnd cell_6t
Xbit_r129_c141 bl[141] br[141] wl[129] vdd gnd cell_6t
Xbit_r130_c141 bl[141] br[141] wl[130] vdd gnd cell_6t
Xbit_r131_c141 bl[141] br[141] wl[131] vdd gnd cell_6t
Xbit_r132_c141 bl[141] br[141] wl[132] vdd gnd cell_6t
Xbit_r133_c141 bl[141] br[141] wl[133] vdd gnd cell_6t
Xbit_r134_c141 bl[141] br[141] wl[134] vdd gnd cell_6t
Xbit_r135_c141 bl[141] br[141] wl[135] vdd gnd cell_6t
Xbit_r136_c141 bl[141] br[141] wl[136] vdd gnd cell_6t
Xbit_r137_c141 bl[141] br[141] wl[137] vdd gnd cell_6t
Xbit_r138_c141 bl[141] br[141] wl[138] vdd gnd cell_6t
Xbit_r139_c141 bl[141] br[141] wl[139] vdd gnd cell_6t
Xbit_r140_c141 bl[141] br[141] wl[140] vdd gnd cell_6t
Xbit_r141_c141 bl[141] br[141] wl[141] vdd gnd cell_6t
Xbit_r142_c141 bl[141] br[141] wl[142] vdd gnd cell_6t
Xbit_r143_c141 bl[141] br[141] wl[143] vdd gnd cell_6t
Xbit_r144_c141 bl[141] br[141] wl[144] vdd gnd cell_6t
Xbit_r145_c141 bl[141] br[141] wl[145] vdd gnd cell_6t
Xbit_r146_c141 bl[141] br[141] wl[146] vdd gnd cell_6t
Xbit_r147_c141 bl[141] br[141] wl[147] vdd gnd cell_6t
Xbit_r148_c141 bl[141] br[141] wl[148] vdd gnd cell_6t
Xbit_r149_c141 bl[141] br[141] wl[149] vdd gnd cell_6t
Xbit_r150_c141 bl[141] br[141] wl[150] vdd gnd cell_6t
Xbit_r151_c141 bl[141] br[141] wl[151] vdd gnd cell_6t
Xbit_r152_c141 bl[141] br[141] wl[152] vdd gnd cell_6t
Xbit_r153_c141 bl[141] br[141] wl[153] vdd gnd cell_6t
Xbit_r154_c141 bl[141] br[141] wl[154] vdd gnd cell_6t
Xbit_r155_c141 bl[141] br[141] wl[155] vdd gnd cell_6t
Xbit_r156_c141 bl[141] br[141] wl[156] vdd gnd cell_6t
Xbit_r157_c141 bl[141] br[141] wl[157] vdd gnd cell_6t
Xbit_r158_c141 bl[141] br[141] wl[158] vdd gnd cell_6t
Xbit_r159_c141 bl[141] br[141] wl[159] vdd gnd cell_6t
Xbit_r160_c141 bl[141] br[141] wl[160] vdd gnd cell_6t
Xbit_r161_c141 bl[141] br[141] wl[161] vdd gnd cell_6t
Xbit_r162_c141 bl[141] br[141] wl[162] vdd gnd cell_6t
Xbit_r163_c141 bl[141] br[141] wl[163] vdd gnd cell_6t
Xbit_r164_c141 bl[141] br[141] wl[164] vdd gnd cell_6t
Xbit_r165_c141 bl[141] br[141] wl[165] vdd gnd cell_6t
Xbit_r166_c141 bl[141] br[141] wl[166] vdd gnd cell_6t
Xbit_r167_c141 bl[141] br[141] wl[167] vdd gnd cell_6t
Xbit_r168_c141 bl[141] br[141] wl[168] vdd gnd cell_6t
Xbit_r169_c141 bl[141] br[141] wl[169] vdd gnd cell_6t
Xbit_r170_c141 bl[141] br[141] wl[170] vdd gnd cell_6t
Xbit_r171_c141 bl[141] br[141] wl[171] vdd gnd cell_6t
Xbit_r172_c141 bl[141] br[141] wl[172] vdd gnd cell_6t
Xbit_r173_c141 bl[141] br[141] wl[173] vdd gnd cell_6t
Xbit_r174_c141 bl[141] br[141] wl[174] vdd gnd cell_6t
Xbit_r175_c141 bl[141] br[141] wl[175] vdd gnd cell_6t
Xbit_r176_c141 bl[141] br[141] wl[176] vdd gnd cell_6t
Xbit_r177_c141 bl[141] br[141] wl[177] vdd gnd cell_6t
Xbit_r178_c141 bl[141] br[141] wl[178] vdd gnd cell_6t
Xbit_r179_c141 bl[141] br[141] wl[179] vdd gnd cell_6t
Xbit_r180_c141 bl[141] br[141] wl[180] vdd gnd cell_6t
Xbit_r181_c141 bl[141] br[141] wl[181] vdd gnd cell_6t
Xbit_r182_c141 bl[141] br[141] wl[182] vdd gnd cell_6t
Xbit_r183_c141 bl[141] br[141] wl[183] vdd gnd cell_6t
Xbit_r184_c141 bl[141] br[141] wl[184] vdd gnd cell_6t
Xbit_r185_c141 bl[141] br[141] wl[185] vdd gnd cell_6t
Xbit_r186_c141 bl[141] br[141] wl[186] vdd gnd cell_6t
Xbit_r187_c141 bl[141] br[141] wl[187] vdd gnd cell_6t
Xbit_r188_c141 bl[141] br[141] wl[188] vdd gnd cell_6t
Xbit_r189_c141 bl[141] br[141] wl[189] vdd gnd cell_6t
Xbit_r190_c141 bl[141] br[141] wl[190] vdd gnd cell_6t
Xbit_r191_c141 bl[141] br[141] wl[191] vdd gnd cell_6t
Xbit_r192_c141 bl[141] br[141] wl[192] vdd gnd cell_6t
Xbit_r193_c141 bl[141] br[141] wl[193] vdd gnd cell_6t
Xbit_r194_c141 bl[141] br[141] wl[194] vdd gnd cell_6t
Xbit_r195_c141 bl[141] br[141] wl[195] vdd gnd cell_6t
Xbit_r196_c141 bl[141] br[141] wl[196] vdd gnd cell_6t
Xbit_r197_c141 bl[141] br[141] wl[197] vdd gnd cell_6t
Xbit_r198_c141 bl[141] br[141] wl[198] vdd gnd cell_6t
Xbit_r199_c141 bl[141] br[141] wl[199] vdd gnd cell_6t
Xbit_r200_c141 bl[141] br[141] wl[200] vdd gnd cell_6t
Xbit_r201_c141 bl[141] br[141] wl[201] vdd gnd cell_6t
Xbit_r202_c141 bl[141] br[141] wl[202] vdd gnd cell_6t
Xbit_r203_c141 bl[141] br[141] wl[203] vdd gnd cell_6t
Xbit_r204_c141 bl[141] br[141] wl[204] vdd gnd cell_6t
Xbit_r205_c141 bl[141] br[141] wl[205] vdd gnd cell_6t
Xbit_r206_c141 bl[141] br[141] wl[206] vdd gnd cell_6t
Xbit_r207_c141 bl[141] br[141] wl[207] vdd gnd cell_6t
Xbit_r208_c141 bl[141] br[141] wl[208] vdd gnd cell_6t
Xbit_r209_c141 bl[141] br[141] wl[209] vdd gnd cell_6t
Xbit_r210_c141 bl[141] br[141] wl[210] vdd gnd cell_6t
Xbit_r211_c141 bl[141] br[141] wl[211] vdd gnd cell_6t
Xbit_r212_c141 bl[141] br[141] wl[212] vdd gnd cell_6t
Xbit_r213_c141 bl[141] br[141] wl[213] vdd gnd cell_6t
Xbit_r214_c141 bl[141] br[141] wl[214] vdd gnd cell_6t
Xbit_r215_c141 bl[141] br[141] wl[215] vdd gnd cell_6t
Xbit_r216_c141 bl[141] br[141] wl[216] vdd gnd cell_6t
Xbit_r217_c141 bl[141] br[141] wl[217] vdd gnd cell_6t
Xbit_r218_c141 bl[141] br[141] wl[218] vdd gnd cell_6t
Xbit_r219_c141 bl[141] br[141] wl[219] vdd gnd cell_6t
Xbit_r220_c141 bl[141] br[141] wl[220] vdd gnd cell_6t
Xbit_r221_c141 bl[141] br[141] wl[221] vdd gnd cell_6t
Xbit_r222_c141 bl[141] br[141] wl[222] vdd gnd cell_6t
Xbit_r223_c141 bl[141] br[141] wl[223] vdd gnd cell_6t
Xbit_r224_c141 bl[141] br[141] wl[224] vdd gnd cell_6t
Xbit_r225_c141 bl[141] br[141] wl[225] vdd gnd cell_6t
Xbit_r226_c141 bl[141] br[141] wl[226] vdd gnd cell_6t
Xbit_r227_c141 bl[141] br[141] wl[227] vdd gnd cell_6t
Xbit_r228_c141 bl[141] br[141] wl[228] vdd gnd cell_6t
Xbit_r229_c141 bl[141] br[141] wl[229] vdd gnd cell_6t
Xbit_r230_c141 bl[141] br[141] wl[230] vdd gnd cell_6t
Xbit_r231_c141 bl[141] br[141] wl[231] vdd gnd cell_6t
Xbit_r232_c141 bl[141] br[141] wl[232] vdd gnd cell_6t
Xbit_r233_c141 bl[141] br[141] wl[233] vdd gnd cell_6t
Xbit_r234_c141 bl[141] br[141] wl[234] vdd gnd cell_6t
Xbit_r235_c141 bl[141] br[141] wl[235] vdd gnd cell_6t
Xbit_r236_c141 bl[141] br[141] wl[236] vdd gnd cell_6t
Xbit_r237_c141 bl[141] br[141] wl[237] vdd gnd cell_6t
Xbit_r238_c141 bl[141] br[141] wl[238] vdd gnd cell_6t
Xbit_r239_c141 bl[141] br[141] wl[239] vdd gnd cell_6t
Xbit_r240_c141 bl[141] br[141] wl[240] vdd gnd cell_6t
Xbit_r241_c141 bl[141] br[141] wl[241] vdd gnd cell_6t
Xbit_r242_c141 bl[141] br[141] wl[242] vdd gnd cell_6t
Xbit_r243_c141 bl[141] br[141] wl[243] vdd gnd cell_6t
Xbit_r244_c141 bl[141] br[141] wl[244] vdd gnd cell_6t
Xbit_r245_c141 bl[141] br[141] wl[245] vdd gnd cell_6t
Xbit_r246_c141 bl[141] br[141] wl[246] vdd gnd cell_6t
Xbit_r247_c141 bl[141] br[141] wl[247] vdd gnd cell_6t
Xbit_r248_c141 bl[141] br[141] wl[248] vdd gnd cell_6t
Xbit_r249_c141 bl[141] br[141] wl[249] vdd gnd cell_6t
Xbit_r250_c141 bl[141] br[141] wl[250] vdd gnd cell_6t
Xbit_r251_c141 bl[141] br[141] wl[251] vdd gnd cell_6t
Xbit_r252_c141 bl[141] br[141] wl[252] vdd gnd cell_6t
Xbit_r253_c141 bl[141] br[141] wl[253] vdd gnd cell_6t
Xbit_r254_c141 bl[141] br[141] wl[254] vdd gnd cell_6t
Xbit_r255_c141 bl[141] br[141] wl[255] vdd gnd cell_6t
Xbit_r0_c142 bl[142] br[142] wl[0] vdd gnd cell_6t
Xbit_r1_c142 bl[142] br[142] wl[1] vdd gnd cell_6t
Xbit_r2_c142 bl[142] br[142] wl[2] vdd gnd cell_6t
Xbit_r3_c142 bl[142] br[142] wl[3] vdd gnd cell_6t
Xbit_r4_c142 bl[142] br[142] wl[4] vdd gnd cell_6t
Xbit_r5_c142 bl[142] br[142] wl[5] vdd gnd cell_6t
Xbit_r6_c142 bl[142] br[142] wl[6] vdd gnd cell_6t
Xbit_r7_c142 bl[142] br[142] wl[7] vdd gnd cell_6t
Xbit_r8_c142 bl[142] br[142] wl[8] vdd gnd cell_6t
Xbit_r9_c142 bl[142] br[142] wl[9] vdd gnd cell_6t
Xbit_r10_c142 bl[142] br[142] wl[10] vdd gnd cell_6t
Xbit_r11_c142 bl[142] br[142] wl[11] vdd gnd cell_6t
Xbit_r12_c142 bl[142] br[142] wl[12] vdd gnd cell_6t
Xbit_r13_c142 bl[142] br[142] wl[13] vdd gnd cell_6t
Xbit_r14_c142 bl[142] br[142] wl[14] vdd gnd cell_6t
Xbit_r15_c142 bl[142] br[142] wl[15] vdd gnd cell_6t
Xbit_r16_c142 bl[142] br[142] wl[16] vdd gnd cell_6t
Xbit_r17_c142 bl[142] br[142] wl[17] vdd gnd cell_6t
Xbit_r18_c142 bl[142] br[142] wl[18] vdd gnd cell_6t
Xbit_r19_c142 bl[142] br[142] wl[19] vdd gnd cell_6t
Xbit_r20_c142 bl[142] br[142] wl[20] vdd gnd cell_6t
Xbit_r21_c142 bl[142] br[142] wl[21] vdd gnd cell_6t
Xbit_r22_c142 bl[142] br[142] wl[22] vdd gnd cell_6t
Xbit_r23_c142 bl[142] br[142] wl[23] vdd gnd cell_6t
Xbit_r24_c142 bl[142] br[142] wl[24] vdd gnd cell_6t
Xbit_r25_c142 bl[142] br[142] wl[25] vdd gnd cell_6t
Xbit_r26_c142 bl[142] br[142] wl[26] vdd gnd cell_6t
Xbit_r27_c142 bl[142] br[142] wl[27] vdd gnd cell_6t
Xbit_r28_c142 bl[142] br[142] wl[28] vdd gnd cell_6t
Xbit_r29_c142 bl[142] br[142] wl[29] vdd gnd cell_6t
Xbit_r30_c142 bl[142] br[142] wl[30] vdd gnd cell_6t
Xbit_r31_c142 bl[142] br[142] wl[31] vdd gnd cell_6t
Xbit_r32_c142 bl[142] br[142] wl[32] vdd gnd cell_6t
Xbit_r33_c142 bl[142] br[142] wl[33] vdd gnd cell_6t
Xbit_r34_c142 bl[142] br[142] wl[34] vdd gnd cell_6t
Xbit_r35_c142 bl[142] br[142] wl[35] vdd gnd cell_6t
Xbit_r36_c142 bl[142] br[142] wl[36] vdd gnd cell_6t
Xbit_r37_c142 bl[142] br[142] wl[37] vdd gnd cell_6t
Xbit_r38_c142 bl[142] br[142] wl[38] vdd gnd cell_6t
Xbit_r39_c142 bl[142] br[142] wl[39] vdd gnd cell_6t
Xbit_r40_c142 bl[142] br[142] wl[40] vdd gnd cell_6t
Xbit_r41_c142 bl[142] br[142] wl[41] vdd gnd cell_6t
Xbit_r42_c142 bl[142] br[142] wl[42] vdd gnd cell_6t
Xbit_r43_c142 bl[142] br[142] wl[43] vdd gnd cell_6t
Xbit_r44_c142 bl[142] br[142] wl[44] vdd gnd cell_6t
Xbit_r45_c142 bl[142] br[142] wl[45] vdd gnd cell_6t
Xbit_r46_c142 bl[142] br[142] wl[46] vdd gnd cell_6t
Xbit_r47_c142 bl[142] br[142] wl[47] vdd gnd cell_6t
Xbit_r48_c142 bl[142] br[142] wl[48] vdd gnd cell_6t
Xbit_r49_c142 bl[142] br[142] wl[49] vdd gnd cell_6t
Xbit_r50_c142 bl[142] br[142] wl[50] vdd gnd cell_6t
Xbit_r51_c142 bl[142] br[142] wl[51] vdd gnd cell_6t
Xbit_r52_c142 bl[142] br[142] wl[52] vdd gnd cell_6t
Xbit_r53_c142 bl[142] br[142] wl[53] vdd gnd cell_6t
Xbit_r54_c142 bl[142] br[142] wl[54] vdd gnd cell_6t
Xbit_r55_c142 bl[142] br[142] wl[55] vdd gnd cell_6t
Xbit_r56_c142 bl[142] br[142] wl[56] vdd gnd cell_6t
Xbit_r57_c142 bl[142] br[142] wl[57] vdd gnd cell_6t
Xbit_r58_c142 bl[142] br[142] wl[58] vdd gnd cell_6t
Xbit_r59_c142 bl[142] br[142] wl[59] vdd gnd cell_6t
Xbit_r60_c142 bl[142] br[142] wl[60] vdd gnd cell_6t
Xbit_r61_c142 bl[142] br[142] wl[61] vdd gnd cell_6t
Xbit_r62_c142 bl[142] br[142] wl[62] vdd gnd cell_6t
Xbit_r63_c142 bl[142] br[142] wl[63] vdd gnd cell_6t
Xbit_r64_c142 bl[142] br[142] wl[64] vdd gnd cell_6t
Xbit_r65_c142 bl[142] br[142] wl[65] vdd gnd cell_6t
Xbit_r66_c142 bl[142] br[142] wl[66] vdd gnd cell_6t
Xbit_r67_c142 bl[142] br[142] wl[67] vdd gnd cell_6t
Xbit_r68_c142 bl[142] br[142] wl[68] vdd gnd cell_6t
Xbit_r69_c142 bl[142] br[142] wl[69] vdd gnd cell_6t
Xbit_r70_c142 bl[142] br[142] wl[70] vdd gnd cell_6t
Xbit_r71_c142 bl[142] br[142] wl[71] vdd gnd cell_6t
Xbit_r72_c142 bl[142] br[142] wl[72] vdd gnd cell_6t
Xbit_r73_c142 bl[142] br[142] wl[73] vdd gnd cell_6t
Xbit_r74_c142 bl[142] br[142] wl[74] vdd gnd cell_6t
Xbit_r75_c142 bl[142] br[142] wl[75] vdd gnd cell_6t
Xbit_r76_c142 bl[142] br[142] wl[76] vdd gnd cell_6t
Xbit_r77_c142 bl[142] br[142] wl[77] vdd gnd cell_6t
Xbit_r78_c142 bl[142] br[142] wl[78] vdd gnd cell_6t
Xbit_r79_c142 bl[142] br[142] wl[79] vdd gnd cell_6t
Xbit_r80_c142 bl[142] br[142] wl[80] vdd gnd cell_6t
Xbit_r81_c142 bl[142] br[142] wl[81] vdd gnd cell_6t
Xbit_r82_c142 bl[142] br[142] wl[82] vdd gnd cell_6t
Xbit_r83_c142 bl[142] br[142] wl[83] vdd gnd cell_6t
Xbit_r84_c142 bl[142] br[142] wl[84] vdd gnd cell_6t
Xbit_r85_c142 bl[142] br[142] wl[85] vdd gnd cell_6t
Xbit_r86_c142 bl[142] br[142] wl[86] vdd gnd cell_6t
Xbit_r87_c142 bl[142] br[142] wl[87] vdd gnd cell_6t
Xbit_r88_c142 bl[142] br[142] wl[88] vdd gnd cell_6t
Xbit_r89_c142 bl[142] br[142] wl[89] vdd gnd cell_6t
Xbit_r90_c142 bl[142] br[142] wl[90] vdd gnd cell_6t
Xbit_r91_c142 bl[142] br[142] wl[91] vdd gnd cell_6t
Xbit_r92_c142 bl[142] br[142] wl[92] vdd gnd cell_6t
Xbit_r93_c142 bl[142] br[142] wl[93] vdd gnd cell_6t
Xbit_r94_c142 bl[142] br[142] wl[94] vdd gnd cell_6t
Xbit_r95_c142 bl[142] br[142] wl[95] vdd gnd cell_6t
Xbit_r96_c142 bl[142] br[142] wl[96] vdd gnd cell_6t
Xbit_r97_c142 bl[142] br[142] wl[97] vdd gnd cell_6t
Xbit_r98_c142 bl[142] br[142] wl[98] vdd gnd cell_6t
Xbit_r99_c142 bl[142] br[142] wl[99] vdd gnd cell_6t
Xbit_r100_c142 bl[142] br[142] wl[100] vdd gnd cell_6t
Xbit_r101_c142 bl[142] br[142] wl[101] vdd gnd cell_6t
Xbit_r102_c142 bl[142] br[142] wl[102] vdd gnd cell_6t
Xbit_r103_c142 bl[142] br[142] wl[103] vdd gnd cell_6t
Xbit_r104_c142 bl[142] br[142] wl[104] vdd gnd cell_6t
Xbit_r105_c142 bl[142] br[142] wl[105] vdd gnd cell_6t
Xbit_r106_c142 bl[142] br[142] wl[106] vdd gnd cell_6t
Xbit_r107_c142 bl[142] br[142] wl[107] vdd gnd cell_6t
Xbit_r108_c142 bl[142] br[142] wl[108] vdd gnd cell_6t
Xbit_r109_c142 bl[142] br[142] wl[109] vdd gnd cell_6t
Xbit_r110_c142 bl[142] br[142] wl[110] vdd gnd cell_6t
Xbit_r111_c142 bl[142] br[142] wl[111] vdd gnd cell_6t
Xbit_r112_c142 bl[142] br[142] wl[112] vdd gnd cell_6t
Xbit_r113_c142 bl[142] br[142] wl[113] vdd gnd cell_6t
Xbit_r114_c142 bl[142] br[142] wl[114] vdd gnd cell_6t
Xbit_r115_c142 bl[142] br[142] wl[115] vdd gnd cell_6t
Xbit_r116_c142 bl[142] br[142] wl[116] vdd gnd cell_6t
Xbit_r117_c142 bl[142] br[142] wl[117] vdd gnd cell_6t
Xbit_r118_c142 bl[142] br[142] wl[118] vdd gnd cell_6t
Xbit_r119_c142 bl[142] br[142] wl[119] vdd gnd cell_6t
Xbit_r120_c142 bl[142] br[142] wl[120] vdd gnd cell_6t
Xbit_r121_c142 bl[142] br[142] wl[121] vdd gnd cell_6t
Xbit_r122_c142 bl[142] br[142] wl[122] vdd gnd cell_6t
Xbit_r123_c142 bl[142] br[142] wl[123] vdd gnd cell_6t
Xbit_r124_c142 bl[142] br[142] wl[124] vdd gnd cell_6t
Xbit_r125_c142 bl[142] br[142] wl[125] vdd gnd cell_6t
Xbit_r126_c142 bl[142] br[142] wl[126] vdd gnd cell_6t
Xbit_r127_c142 bl[142] br[142] wl[127] vdd gnd cell_6t
Xbit_r128_c142 bl[142] br[142] wl[128] vdd gnd cell_6t
Xbit_r129_c142 bl[142] br[142] wl[129] vdd gnd cell_6t
Xbit_r130_c142 bl[142] br[142] wl[130] vdd gnd cell_6t
Xbit_r131_c142 bl[142] br[142] wl[131] vdd gnd cell_6t
Xbit_r132_c142 bl[142] br[142] wl[132] vdd gnd cell_6t
Xbit_r133_c142 bl[142] br[142] wl[133] vdd gnd cell_6t
Xbit_r134_c142 bl[142] br[142] wl[134] vdd gnd cell_6t
Xbit_r135_c142 bl[142] br[142] wl[135] vdd gnd cell_6t
Xbit_r136_c142 bl[142] br[142] wl[136] vdd gnd cell_6t
Xbit_r137_c142 bl[142] br[142] wl[137] vdd gnd cell_6t
Xbit_r138_c142 bl[142] br[142] wl[138] vdd gnd cell_6t
Xbit_r139_c142 bl[142] br[142] wl[139] vdd gnd cell_6t
Xbit_r140_c142 bl[142] br[142] wl[140] vdd gnd cell_6t
Xbit_r141_c142 bl[142] br[142] wl[141] vdd gnd cell_6t
Xbit_r142_c142 bl[142] br[142] wl[142] vdd gnd cell_6t
Xbit_r143_c142 bl[142] br[142] wl[143] vdd gnd cell_6t
Xbit_r144_c142 bl[142] br[142] wl[144] vdd gnd cell_6t
Xbit_r145_c142 bl[142] br[142] wl[145] vdd gnd cell_6t
Xbit_r146_c142 bl[142] br[142] wl[146] vdd gnd cell_6t
Xbit_r147_c142 bl[142] br[142] wl[147] vdd gnd cell_6t
Xbit_r148_c142 bl[142] br[142] wl[148] vdd gnd cell_6t
Xbit_r149_c142 bl[142] br[142] wl[149] vdd gnd cell_6t
Xbit_r150_c142 bl[142] br[142] wl[150] vdd gnd cell_6t
Xbit_r151_c142 bl[142] br[142] wl[151] vdd gnd cell_6t
Xbit_r152_c142 bl[142] br[142] wl[152] vdd gnd cell_6t
Xbit_r153_c142 bl[142] br[142] wl[153] vdd gnd cell_6t
Xbit_r154_c142 bl[142] br[142] wl[154] vdd gnd cell_6t
Xbit_r155_c142 bl[142] br[142] wl[155] vdd gnd cell_6t
Xbit_r156_c142 bl[142] br[142] wl[156] vdd gnd cell_6t
Xbit_r157_c142 bl[142] br[142] wl[157] vdd gnd cell_6t
Xbit_r158_c142 bl[142] br[142] wl[158] vdd gnd cell_6t
Xbit_r159_c142 bl[142] br[142] wl[159] vdd gnd cell_6t
Xbit_r160_c142 bl[142] br[142] wl[160] vdd gnd cell_6t
Xbit_r161_c142 bl[142] br[142] wl[161] vdd gnd cell_6t
Xbit_r162_c142 bl[142] br[142] wl[162] vdd gnd cell_6t
Xbit_r163_c142 bl[142] br[142] wl[163] vdd gnd cell_6t
Xbit_r164_c142 bl[142] br[142] wl[164] vdd gnd cell_6t
Xbit_r165_c142 bl[142] br[142] wl[165] vdd gnd cell_6t
Xbit_r166_c142 bl[142] br[142] wl[166] vdd gnd cell_6t
Xbit_r167_c142 bl[142] br[142] wl[167] vdd gnd cell_6t
Xbit_r168_c142 bl[142] br[142] wl[168] vdd gnd cell_6t
Xbit_r169_c142 bl[142] br[142] wl[169] vdd gnd cell_6t
Xbit_r170_c142 bl[142] br[142] wl[170] vdd gnd cell_6t
Xbit_r171_c142 bl[142] br[142] wl[171] vdd gnd cell_6t
Xbit_r172_c142 bl[142] br[142] wl[172] vdd gnd cell_6t
Xbit_r173_c142 bl[142] br[142] wl[173] vdd gnd cell_6t
Xbit_r174_c142 bl[142] br[142] wl[174] vdd gnd cell_6t
Xbit_r175_c142 bl[142] br[142] wl[175] vdd gnd cell_6t
Xbit_r176_c142 bl[142] br[142] wl[176] vdd gnd cell_6t
Xbit_r177_c142 bl[142] br[142] wl[177] vdd gnd cell_6t
Xbit_r178_c142 bl[142] br[142] wl[178] vdd gnd cell_6t
Xbit_r179_c142 bl[142] br[142] wl[179] vdd gnd cell_6t
Xbit_r180_c142 bl[142] br[142] wl[180] vdd gnd cell_6t
Xbit_r181_c142 bl[142] br[142] wl[181] vdd gnd cell_6t
Xbit_r182_c142 bl[142] br[142] wl[182] vdd gnd cell_6t
Xbit_r183_c142 bl[142] br[142] wl[183] vdd gnd cell_6t
Xbit_r184_c142 bl[142] br[142] wl[184] vdd gnd cell_6t
Xbit_r185_c142 bl[142] br[142] wl[185] vdd gnd cell_6t
Xbit_r186_c142 bl[142] br[142] wl[186] vdd gnd cell_6t
Xbit_r187_c142 bl[142] br[142] wl[187] vdd gnd cell_6t
Xbit_r188_c142 bl[142] br[142] wl[188] vdd gnd cell_6t
Xbit_r189_c142 bl[142] br[142] wl[189] vdd gnd cell_6t
Xbit_r190_c142 bl[142] br[142] wl[190] vdd gnd cell_6t
Xbit_r191_c142 bl[142] br[142] wl[191] vdd gnd cell_6t
Xbit_r192_c142 bl[142] br[142] wl[192] vdd gnd cell_6t
Xbit_r193_c142 bl[142] br[142] wl[193] vdd gnd cell_6t
Xbit_r194_c142 bl[142] br[142] wl[194] vdd gnd cell_6t
Xbit_r195_c142 bl[142] br[142] wl[195] vdd gnd cell_6t
Xbit_r196_c142 bl[142] br[142] wl[196] vdd gnd cell_6t
Xbit_r197_c142 bl[142] br[142] wl[197] vdd gnd cell_6t
Xbit_r198_c142 bl[142] br[142] wl[198] vdd gnd cell_6t
Xbit_r199_c142 bl[142] br[142] wl[199] vdd gnd cell_6t
Xbit_r200_c142 bl[142] br[142] wl[200] vdd gnd cell_6t
Xbit_r201_c142 bl[142] br[142] wl[201] vdd gnd cell_6t
Xbit_r202_c142 bl[142] br[142] wl[202] vdd gnd cell_6t
Xbit_r203_c142 bl[142] br[142] wl[203] vdd gnd cell_6t
Xbit_r204_c142 bl[142] br[142] wl[204] vdd gnd cell_6t
Xbit_r205_c142 bl[142] br[142] wl[205] vdd gnd cell_6t
Xbit_r206_c142 bl[142] br[142] wl[206] vdd gnd cell_6t
Xbit_r207_c142 bl[142] br[142] wl[207] vdd gnd cell_6t
Xbit_r208_c142 bl[142] br[142] wl[208] vdd gnd cell_6t
Xbit_r209_c142 bl[142] br[142] wl[209] vdd gnd cell_6t
Xbit_r210_c142 bl[142] br[142] wl[210] vdd gnd cell_6t
Xbit_r211_c142 bl[142] br[142] wl[211] vdd gnd cell_6t
Xbit_r212_c142 bl[142] br[142] wl[212] vdd gnd cell_6t
Xbit_r213_c142 bl[142] br[142] wl[213] vdd gnd cell_6t
Xbit_r214_c142 bl[142] br[142] wl[214] vdd gnd cell_6t
Xbit_r215_c142 bl[142] br[142] wl[215] vdd gnd cell_6t
Xbit_r216_c142 bl[142] br[142] wl[216] vdd gnd cell_6t
Xbit_r217_c142 bl[142] br[142] wl[217] vdd gnd cell_6t
Xbit_r218_c142 bl[142] br[142] wl[218] vdd gnd cell_6t
Xbit_r219_c142 bl[142] br[142] wl[219] vdd gnd cell_6t
Xbit_r220_c142 bl[142] br[142] wl[220] vdd gnd cell_6t
Xbit_r221_c142 bl[142] br[142] wl[221] vdd gnd cell_6t
Xbit_r222_c142 bl[142] br[142] wl[222] vdd gnd cell_6t
Xbit_r223_c142 bl[142] br[142] wl[223] vdd gnd cell_6t
Xbit_r224_c142 bl[142] br[142] wl[224] vdd gnd cell_6t
Xbit_r225_c142 bl[142] br[142] wl[225] vdd gnd cell_6t
Xbit_r226_c142 bl[142] br[142] wl[226] vdd gnd cell_6t
Xbit_r227_c142 bl[142] br[142] wl[227] vdd gnd cell_6t
Xbit_r228_c142 bl[142] br[142] wl[228] vdd gnd cell_6t
Xbit_r229_c142 bl[142] br[142] wl[229] vdd gnd cell_6t
Xbit_r230_c142 bl[142] br[142] wl[230] vdd gnd cell_6t
Xbit_r231_c142 bl[142] br[142] wl[231] vdd gnd cell_6t
Xbit_r232_c142 bl[142] br[142] wl[232] vdd gnd cell_6t
Xbit_r233_c142 bl[142] br[142] wl[233] vdd gnd cell_6t
Xbit_r234_c142 bl[142] br[142] wl[234] vdd gnd cell_6t
Xbit_r235_c142 bl[142] br[142] wl[235] vdd gnd cell_6t
Xbit_r236_c142 bl[142] br[142] wl[236] vdd gnd cell_6t
Xbit_r237_c142 bl[142] br[142] wl[237] vdd gnd cell_6t
Xbit_r238_c142 bl[142] br[142] wl[238] vdd gnd cell_6t
Xbit_r239_c142 bl[142] br[142] wl[239] vdd gnd cell_6t
Xbit_r240_c142 bl[142] br[142] wl[240] vdd gnd cell_6t
Xbit_r241_c142 bl[142] br[142] wl[241] vdd gnd cell_6t
Xbit_r242_c142 bl[142] br[142] wl[242] vdd gnd cell_6t
Xbit_r243_c142 bl[142] br[142] wl[243] vdd gnd cell_6t
Xbit_r244_c142 bl[142] br[142] wl[244] vdd gnd cell_6t
Xbit_r245_c142 bl[142] br[142] wl[245] vdd gnd cell_6t
Xbit_r246_c142 bl[142] br[142] wl[246] vdd gnd cell_6t
Xbit_r247_c142 bl[142] br[142] wl[247] vdd gnd cell_6t
Xbit_r248_c142 bl[142] br[142] wl[248] vdd gnd cell_6t
Xbit_r249_c142 bl[142] br[142] wl[249] vdd gnd cell_6t
Xbit_r250_c142 bl[142] br[142] wl[250] vdd gnd cell_6t
Xbit_r251_c142 bl[142] br[142] wl[251] vdd gnd cell_6t
Xbit_r252_c142 bl[142] br[142] wl[252] vdd gnd cell_6t
Xbit_r253_c142 bl[142] br[142] wl[253] vdd gnd cell_6t
Xbit_r254_c142 bl[142] br[142] wl[254] vdd gnd cell_6t
Xbit_r255_c142 bl[142] br[142] wl[255] vdd gnd cell_6t
Xbit_r0_c143 bl[143] br[143] wl[0] vdd gnd cell_6t
Xbit_r1_c143 bl[143] br[143] wl[1] vdd gnd cell_6t
Xbit_r2_c143 bl[143] br[143] wl[2] vdd gnd cell_6t
Xbit_r3_c143 bl[143] br[143] wl[3] vdd gnd cell_6t
Xbit_r4_c143 bl[143] br[143] wl[4] vdd gnd cell_6t
Xbit_r5_c143 bl[143] br[143] wl[5] vdd gnd cell_6t
Xbit_r6_c143 bl[143] br[143] wl[6] vdd gnd cell_6t
Xbit_r7_c143 bl[143] br[143] wl[7] vdd gnd cell_6t
Xbit_r8_c143 bl[143] br[143] wl[8] vdd gnd cell_6t
Xbit_r9_c143 bl[143] br[143] wl[9] vdd gnd cell_6t
Xbit_r10_c143 bl[143] br[143] wl[10] vdd gnd cell_6t
Xbit_r11_c143 bl[143] br[143] wl[11] vdd gnd cell_6t
Xbit_r12_c143 bl[143] br[143] wl[12] vdd gnd cell_6t
Xbit_r13_c143 bl[143] br[143] wl[13] vdd gnd cell_6t
Xbit_r14_c143 bl[143] br[143] wl[14] vdd gnd cell_6t
Xbit_r15_c143 bl[143] br[143] wl[15] vdd gnd cell_6t
Xbit_r16_c143 bl[143] br[143] wl[16] vdd gnd cell_6t
Xbit_r17_c143 bl[143] br[143] wl[17] vdd gnd cell_6t
Xbit_r18_c143 bl[143] br[143] wl[18] vdd gnd cell_6t
Xbit_r19_c143 bl[143] br[143] wl[19] vdd gnd cell_6t
Xbit_r20_c143 bl[143] br[143] wl[20] vdd gnd cell_6t
Xbit_r21_c143 bl[143] br[143] wl[21] vdd gnd cell_6t
Xbit_r22_c143 bl[143] br[143] wl[22] vdd gnd cell_6t
Xbit_r23_c143 bl[143] br[143] wl[23] vdd gnd cell_6t
Xbit_r24_c143 bl[143] br[143] wl[24] vdd gnd cell_6t
Xbit_r25_c143 bl[143] br[143] wl[25] vdd gnd cell_6t
Xbit_r26_c143 bl[143] br[143] wl[26] vdd gnd cell_6t
Xbit_r27_c143 bl[143] br[143] wl[27] vdd gnd cell_6t
Xbit_r28_c143 bl[143] br[143] wl[28] vdd gnd cell_6t
Xbit_r29_c143 bl[143] br[143] wl[29] vdd gnd cell_6t
Xbit_r30_c143 bl[143] br[143] wl[30] vdd gnd cell_6t
Xbit_r31_c143 bl[143] br[143] wl[31] vdd gnd cell_6t
Xbit_r32_c143 bl[143] br[143] wl[32] vdd gnd cell_6t
Xbit_r33_c143 bl[143] br[143] wl[33] vdd gnd cell_6t
Xbit_r34_c143 bl[143] br[143] wl[34] vdd gnd cell_6t
Xbit_r35_c143 bl[143] br[143] wl[35] vdd gnd cell_6t
Xbit_r36_c143 bl[143] br[143] wl[36] vdd gnd cell_6t
Xbit_r37_c143 bl[143] br[143] wl[37] vdd gnd cell_6t
Xbit_r38_c143 bl[143] br[143] wl[38] vdd gnd cell_6t
Xbit_r39_c143 bl[143] br[143] wl[39] vdd gnd cell_6t
Xbit_r40_c143 bl[143] br[143] wl[40] vdd gnd cell_6t
Xbit_r41_c143 bl[143] br[143] wl[41] vdd gnd cell_6t
Xbit_r42_c143 bl[143] br[143] wl[42] vdd gnd cell_6t
Xbit_r43_c143 bl[143] br[143] wl[43] vdd gnd cell_6t
Xbit_r44_c143 bl[143] br[143] wl[44] vdd gnd cell_6t
Xbit_r45_c143 bl[143] br[143] wl[45] vdd gnd cell_6t
Xbit_r46_c143 bl[143] br[143] wl[46] vdd gnd cell_6t
Xbit_r47_c143 bl[143] br[143] wl[47] vdd gnd cell_6t
Xbit_r48_c143 bl[143] br[143] wl[48] vdd gnd cell_6t
Xbit_r49_c143 bl[143] br[143] wl[49] vdd gnd cell_6t
Xbit_r50_c143 bl[143] br[143] wl[50] vdd gnd cell_6t
Xbit_r51_c143 bl[143] br[143] wl[51] vdd gnd cell_6t
Xbit_r52_c143 bl[143] br[143] wl[52] vdd gnd cell_6t
Xbit_r53_c143 bl[143] br[143] wl[53] vdd gnd cell_6t
Xbit_r54_c143 bl[143] br[143] wl[54] vdd gnd cell_6t
Xbit_r55_c143 bl[143] br[143] wl[55] vdd gnd cell_6t
Xbit_r56_c143 bl[143] br[143] wl[56] vdd gnd cell_6t
Xbit_r57_c143 bl[143] br[143] wl[57] vdd gnd cell_6t
Xbit_r58_c143 bl[143] br[143] wl[58] vdd gnd cell_6t
Xbit_r59_c143 bl[143] br[143] wl[59] vdd gnd cell_6t
Xbit_r60_c143 bl[143] br[143] wl[60] vdd gnd cell_6t
Xbit_r61_c143 bl[143] br[143] wl[61] vdd gnd cell_6t
Xbit_r62_c143 bl[143] br[143] wl[62] vdd gnd cell_6t
Xbit_r63_c143 bl[143] br[143] wl[63] vdd gnd cell_6t
Xbit_r64_c143 bl[143] br[143] wl[64] vdd gnd cell_6t
Xbit_r65_c143 bl[143] br[143] wl[65] vdd gnd cell_6t
Xbit_r66_c143 bl[143] br[143] wl[66] vdd gnd cell_6t
Xbit_r67_c143 bl[143] br[143] wl[67] vdd gnd cell_6t
Xbit_r68_c143 bl[143] br[143] wl[68] vdd gnd cell_6t
Xbit_r69_c143 bl[143] br[143] wl[69] vdd gnd cell_6t
Xbit_r70_c143 bl[143] br[143] wl[70] vdd gnd cell_6t
Xbit_r71_c143 bl[143] br[143] wl[71] vdd gnd cell_6t
Xbit_r72_c143 bl[143] br[143] wl[72] vdd gnd cell_6t
Xbit_r73_c143 bl[143] br[143] wl[73] vdd gnd cell_6t
Xbit_r74_c143 bl[143] br[143] wl[74] vdd gnd cell_6t
Xbit_r75_c143 bl[143] br[143] wl[75] vdd gnd cell_6t
Xbit_r76_c143 bl[143] br[143] wl[76] vdd gnd cell_6t
Xbit_r77_c143 bl[143] br[143] wl[77] vdd gnd cell_6t
Xbit_r78_c143 bl[143] br[143] wl[78] vdd gnd cell_6t
Xbit_r79_c143 bl[143] br[143] wl[79] vdd gnd cell_6t
Xbit_r80_c143 bl[143] br[143] wl[80] vdd gnd cell_6t
Xbit_r81_c143 bl[143] br[143] wl[81] vdd gnd cell_6t
Xbit_r82_c143 bl[143] br[143] wl[82] vdd gnd cell_6t
Xbit_r83_c143 bl[143] br[143] wl[83] vdd gnd cell_6t
Xbit_r84_c143 bl[143] br[143] wl[84] vdd gnd cell_6t
Xbit_r85_c143 bl[143] br[143] wl[85] vdd gnd cell_6t
Xbit_r86_c143 bl[143] br[143] wl[86] vdd gnd cell_6t
Xbit_r87_c143 bl[143] br[143] wl[87] vdd gnd cell_6t
Xbit_r88_c143 bl[143] br[143] wl[88] vdd gnd cell_6t
Xbit_r89_c143 bl[143] br[143] wl[89] vdd gnd cell_6t
Xbit_r90_c143 bl[143] br[143] wl[90] vdd gnd cell_6t
Xbit_r91_c143 bl[143] br[143] wl[91] vdd gnd cell_6t
Xbit_r92_c143 bl[143] br[143] wl[92] vdd gnd cell_6t
Xbit_r93_c143 bl[143] br[143] wl[93] vdd gnd cell_6t
Xbit_r94_c143 bl[143] br[143] wl[94] vdd gnd cell_6t
Xbit_r95_c143 bl[143] br[143] wl[95] vdd gnd cell_6t
Xbit_r96_c143 bl[143] br[143] wl[96] vdd gnd cell_6t
Xbit_r97_c143 bl[143] br[143] wl[97] vdd gnd cell_6t
Xbit_r98_c143 bl[143] br[143] wl[98] vdd gnd cell_6t
Xbit_r99_c143 bl[143] br[143] wl[99] vdd gnd cell_6t
Xbit_r100_c143 bl[143] br[143] wl[100] vdd gnd cell_6t
Xbit_r101_c143 bl[143] br[143] wl[101] vdd gnd cell_6t
Xbit_r102_c143 bl[143] br[143] wl[102] vdd gnd cell_6t
Xbit_r103_c143 bl[143] br[143] wl[103] vdd gnd cell_6t
Xbit_r104_c143 bl[143] br[143] wl[104] vdd gnd cell_6t
Xbit_r105_c143 bl[143] br[143] wl[105] vdd gnd cell_6t
Xbit_r106_c143 bl[143] br[143] wl[106] vdd gnd cell_6t
Xbit_r107_c143 bl[143] br[143] wl[107] vdd gnd cell_6t
Xbit_r108_c143 bl[143] br[143] wl[108] vdd gnd cell_6t
Xbit_r109_c143 bl[143] br[143] wl[109] vdd gnd cell_6t
Xbit_r110_c143 bl[143] br[143] wl[110] vdd gnd cell_6t
Xbit_r111_c143 bl[143] br[143] wl[111] vdd gnd cell_6t
Xbit_r112_c143 bl[143] br[143] wl[112] vdd gnd cell_6t
Xbit_r113_c143 bl[143] br[143] wl[113] vdd gnd cell_6t
Xbit_r114_c143 bl[143] br[143] wl[114] vdd gnd cell_6t
Xbit_r115_c143 bl[143] br[143] wl[115] vdd gnd cell_6t
Xbit_r116_c143 bl[143] br[143] wl[116] vdd gnd cell_6t
Xbit_r117_c143 bl[143] br[143] wl[117] vdd gnd cell_6t
Xbit_r118_c143 bl[143] br[143] wl[118] vdd gnd cell_6t
Xbit_r119_c143 bl[143] br[143] wl[119] vdd gnd cell_6t
Xbit_r120_c143 bl[143] br[143] wl[120] vdd gnd cell_6t
Xbit_r121_c143 bl[143] br[143] wl[121] vdd gnd cell_6t
Xbit_r122_c143 bl[143] br[143] wl[122] vdd gnd cell_6t
Xbit_r123_c143 bl[143] br[143] wl[123] vdd gnd cell_6t
Xbit_r124_c143 bl[143] br[143] wl[124] vdd gnd cell_6t
Xbit_r125_c143 bl[143] br[143] wl[125] vdd gnd cell_6t
Xbit_r126_c143 bl[143] br[143] wl[126] vdd gnd cell_6t
Xbit_r127_c143 bl[143] br[143] wl[127] vdd gnd cell_6t
Xbit_r128_c143 bl[143] br[143] wl[128] vdd gnd cell_6t
Xbit_r129_c143 bl[143] br[143] wl[129] vdd gnd cell_6t
Xbit_r130_c143 bl[143] br[143] wl[130] vdd gnd cell_6t
Xbit_r131_c143 bl[143] br[143] wl[131] vdd gnd cell_6t
Xbit_r132_c143 bl[143] br[143] wl[132] vdd gnd cell_6t
Xbit_r133_c143 bl[143] br[143] wl[133] vdd gnd cell_6t
Xbit_r134_c143 bl[143] br[143] wl[134] vdd gnd cell_6t
Xbit_r135_c143 bl[143] br[143] wl[135] vdd gnd cell_6t
Xbit_r136_c143 bl[143] br[143] wl[136] vdd gnd cell_6t
Xbit_r137_c143 bl[143] br[143] wl[137] vdd gnd cell_6t
Xbit_r138_c143 bl[143] br[143] wl[138] vdd gnd cell_6t
Xbit_r139_c143 bl[143] br[143] wl[139] vdd gnd cell_6t
Xbit_r140_c143 bl[143] br[143] wl[140] vdd gnd cell_6t
Xbit_r141_c143 bl[143] br[143] wl[141] vdd gnd cell_6t
Xbit_r142_c143 bl[143] br[143] wl[142] vdd gnd cell_6t
Xbit_r143_c143 bl[143] br[143] wl[143] vdd gnd cell_6t
Xbit_r144_c143 bl[143] br[143] wl[144] vdd gnd cell_6t
Xbit_r145_c143 bl[143] br[143] wl[145] vdd gnd cell_6t
Xbit_r146_c143 bl[143] br[143] wl[146] vdd gnd cell_6t
Xbit_r147_c143 bl[143] br[143] wl[147] vdd gnd cell_6t
Xbit_r148_c143 bl[143] br[143] wl[148] vdd gnd cell_6t
Xbit_r149_c143 bl[143] br[143] wl[149] vdd gnd cell_6t
Xbit_r150_c143 bl[143] br[143] wl[150] vdd gnd cell_6t
Xbit_r151_c143 bl[143] br[143] wl[151] vdd gnd cell_6t
Xbit_r152_c143 bl[143] br[143] wl[152] vdd gnd cell_6t
Xbit_r153_c143 bl[143] br[143] wl[153] vdd gnd cell_6t
Xbit_r154_c143 bl[143] br[143] wl[154] vdd gnd cell_6t
Xbit_r155_c143 bl[143] br[143] wl[155] vdd gnd cell_6t
Xbit_r156_c143 bl[143] br[143] wl[156] vdd gnd cell_6t
Xbit_r157_c143 bl[143] br[143] wl[157] vdd gnd cell_6t
Xbit_r158_c143 bl[143] br[143] wl[158] vdd gnd cell_6t
Xbit_r159_c143 bl[143] br[143] wl[159] vdd gnd cell_6t
Xbit_r160_c143 bl[143] br[143] wl[160] vdd gnd cell_6t
Xbit_r161_c143 bl[143] br[143] wl[161] vdd gnd cell_6t
Xbit_r162_c143 bl[143] br[143] wl[162] vdd gnd cell_6t
Xbit_r163_c143 bl[143] br[143] wl[163] vdd gnd cell_6t
Xbit_r164_c143 bl[143] br[143] wl[164] vdd gnd cell_6t
Xbit_r165_c143 bl[143] br[143] wl[165] vdd gnd cell_6t
Xbit_r166_c143 bl[143] br[143] wl[166] vdd gnd cell_6t
Xbit_r167_c143 bl[143] br[143] wl[167] vdd gnd cell_6t
Xbit_r168_c143 bl[143] br[143] wl[168] vdd gnd cell_6t
Xbit_r169_c143 bl[143] br[143] wl[169] vdd gnd cell_6t
Xbit_r170_c143 bl[143] br[143] wl[170] vdd gnd cell_6t
Xbit_r171_c143 bl[143] br[143] wl[171] vdd gnd cell_6t
Xbit_r172_c143 bl[143] br[143] wl[172] vdd gnd cell_6t
Xbit_r173_c143 bl[143] br[143] wl[173] vdd gnd cell_6t
Xbit_r174_c143 bl[143] br[143] wl[174] vdd gnd cell_6t
Xbit_r175_c143 bl[143] br[143] wl[175] vdd gnd cell_6t
Xbit_r176_c143 bl[143] br[143] wl[176] vdd gnd cell_6t
Xbit_r177_c143 bl[143] br[143] wl[177] vdd gnd cell_6t
Xbit_r178_c143 bl[143] br[143] wl[178] vdd gnd cell_6t
Xbit_r179_c143 bl[143] br[143] wl[179] vdd gnd cell_6t
Xbit_r180_c143 bl[143] br[143] wl[180] vdd gnd cell_6t
Xbit_r181_c143 bl[143] br[143] wl[181] vdd gnd cell_6t
Xbit_r182_c143 bl[143] br[143] wl[182] vdd gnd cell_6t
Xbit_r183_c143 bl[143] br[143] wl[183] vdd gnd cell_6t
Xbit_r184_c143 bl[143] br[143] wl[184] vdd gnd cell_6t
Xbit_r185_c143 bl[143] br[143] wl[185] vdd gnd cell_6t
Xbit_r186_c143 bl[143] br[143] wl[186] vdd gnd cell_6t
Xbit_r187_c143 bl[143] br[143] wl[187] vdd gnd cell_6t
Xbit_r188_c143 bl[143] br[143] wl[188] vdd gnd cell_6t
Xbit_r189_c143 bl[143] br[143] wl[189] vdd gnd cell_6t
Xbit_r190_c143 bl[143] br[143] wl[190] vdd gnd cell_6t
Xbit_r191_c143 bl[143] br[143] wl[191] vdd gnd cell_6t
Xbit_r192_c143 bl[143] br[143] wl[192] vdd gnd cell_6t
Xbit_r193_c143 bl[143] br[143] wl[193] vdd gnd cell_6t
Xbit_r194_c143 bl[143] br[143] wl[194] vdd gnd cell_6t
Xbit_r195_c143 bl[143] br[143] wl[195] vdd gnd cell_6t
Xbit_r196_c143 bl[143] br[143] wl[196] vdd gnd cell_6t
Xbit_r197_c143 bl[143] br[143] wl[197] vdd gnd cell_6t
Xbit_r198_c143 bl[143] br[143] wl[198] vdd gnd cell_6t
Xbit_r199_c143 bl[143] br[143] wl[199] vdd gnd cell_6t
Xbit_r200_c143 bl[143] br[143] wl[200] vdd gnd cell_6t
Xbit_r201_c143 bl[143] br[143] wl[201] vdd gnd cell_6t
Xbit_r202_c143 bl[143] br[143] wl[202] vdd gnd cell_6t
Xbit_r203_c143 bl[143] br[143] wl[203] vdd gnd cell_6t
Xbit_r204_c143 bl[143] br[143] wl[204] vdd gnd cell_6t
Xbit_r205_c143 bl[143] br[143] wl[205] vdd gnd cell_6t
Xbit_r206_c143 bl[143] br[143] wl[206] vdd gnd cell_6t
Xbit_r207_c143 bl[143] br[143] wl[207] vdd gnd cell_6t
Xbit_r208_c143 bl[143] br[143] wl[208] vdd gnd cell_6t
Xbit_r209_c143 bl[143] br[143] wl[209] vdd gnd cell_6t
Xbit_r210_c143 bl[143] br[143] wl[210] vdd gnd cell_6t
Xbit_r211_c143 bl[143] br[143] wl[211] vdd gnd cell_6t
Xbit_r212_c143 bl[143] br[143] wl[212] vdd gnd cell_6t
Xbit_r213_c143 bl[143] br[143] wl[213] vdd gnd cell_6t
Xbit_r214_c143 bl[143] br[143] wl[214] vdd gnd cell_6t
Xbit_r215_c143 bl[143] br[143] wl[215] vdd gnd cell_6t
Xbit_r216_c143 bl[143] br[143] wl[216] vdd gnd cell_6t
Xbit_r217_c143 bl[143] br[143] wl[217] vdd gnd cell_6t
Xbit_r218_c143 bl[143] br[143] wl[218] vdd gnd cell_6t
Xbit_r219_c143 bl[143] br[143] wl[219] vdd gnd cell_6t
Xbit_r220_c143 bl[143] br[143] wl[220] vdd gnd cell_6t
Xbit_r221_c143 bl[143] br[143] wl[221] vdd gnd cell_6t
Xbit_r222_c143 bl[143] br[143] wl[222] vdd gnd cell_6t
Xbit_r223_c143 bl[143] br[143] wl[223] vdd gnd cell_6t
Xbit_r224_c143 bl[143] br[143] wl[224] vdd gnd cell_6t
Xbit_r225_c143 bl[143] br[143] wl[225] vdd gnd cell_6t
Xbit_r226_c143 bl[143] br[143] wl[226] vdd gnd cell_6t
Xbit_r227_c143 bl[143] br[143] wl[227] vdd gnd cell_6t
Xbit_r228_c143 bl[143] br[143] wl[228] vdd gnd cell_6t
Xbit_r229_c143 bl[143] br[143] wl[229] vdd gnd cell_6t
Xbit_r230_c143 bl[143] br[143] wl[230] vdd gnd cell_6t
Xbit_r231_c143 bl[143] br[143] wl[231] vdd gnd cell_6t
Xbit_r232_c143 bl[143] br[143] wl[232] vdd gnd cell_6t
Xbit_r233_c143 bl[143] br[143] wl[233] vdd gnd cell_6t
Xbit_r234_c143 bl[143] br[143] wl[234] vdd gnd cell_6t
Xbit_r235_c143 bl[143] br[143] wl[235] vdd gnd cell_6t
Xbit_r236_c143 bl[143] br[143] wl[236] vdd gnd cell_6t
Xbit_r237_c143 bl[143] br[143] wl[237] vdd gnd cell_6t
Xbit_r238_c143 bl[143] br[143] wl[238] vdd gnd cell_6t
Xbit_r239_c143 bl[143] br[143] wl[239] vdd gnd cell_6t
Xbit_r240_c143 bl[143] br[143] wl[240] vdd gnd cell_6t
Xbit_r241_c143 bl[143] br[143] wl[241] vdd gnd cell_6t
Xbit_r242_c143 bl[143] br[143] wl[242] vdd gnd cell_6t
Xbit_r243_c143 bl[143] br[143] wl[243] vdd gnd cell_6t
Xbit_r244_c143 bl[143] br[143] wl[244] vdd gnd cell_6t
Xbit_r245_c143 bl[143] br[143] wl[245] vdd gnd cell_6t
Xbit_r246_c143 bl[143] br[143] wl[246] vdd gnd cell_6t
Xbit_r247_c143 bl[143] br[143] wl[247] vdd gnd cell_6t
Xbit_r248_c143 bl[143] br[143] wl[248] vdd gnd cell_6t
Xbit_r249_c143 bl[143] br[143] wl[249] vdd gnd cell_6t
Xbit_r250_c143 bl[143] br[143] wl[250] vdd gnd cell_6t
Xbit_r251_c143 bl[143] br[143] wl[251] vdd gnd cell_6t
Xbit_r252_c143 bl[143] br[143] wl[252] vdd gnd cell_6t
Xbit_r253_c143 bl[143] br[143] wl[253] vdd gnd cell_6t
Xbit_r254_c143 bl[143] br[143] wl[254] vdd gnd cell_6t
Xbit_r255_c143 bl[143] br[143] wl[255] vdd gnd cell_6t
Xbit_r0_c144 bl[144] br[144] wl[0] vdd gnd cell_6t
Xbit_r1_c144 bl[144] br[144] wl[1] vdd gnd cell_6t
Xbit_r2_c144 bl[144] br[144] wl[2] vdd gnd cell_6t
Xbit_r3_c144 bl[144] br[144] wl[3] vdd gnd cell_6t
Xbit_r4_c144 bl[144] br[144] wl[4] vdd gnd cell_6t
Xbit_r5_c144 bl[144] br[144] wl[5] vdd gnd cell_6t
Xbit_r6_c144 bl[144] br[144] wl[6] vdd gnd cell_6t
Xbit_r7_c144 bl[144] br[144] wl[7] vdd gnd cell_6t
Xbit_r8_c144 bl[144] br[144] wl[8] vdd gnd cell_6t
Xbit_r9_c144 bl[144] br[144] wl[9] vdd gnd cell_6t
Xbit_r10_c144 bl[144] br[144] wl[10] vdd gnd cell_6t
Xbit_r11_c144 bl[144] br[144] wl[11] vdd gnd cell_6t
Xbit_r12_c144 bl[144] br[144] wl[12] vdd gnd cell_6t
Xbit_r13_c144 bl[144] br[144] wl[13] vdd gnd cell_6t
Xbit_r14_c144 bl[144] br[144] wl[14] vdd gnd cell_6t
Xbit_r15_c144 bl[144] br[144] wl[15] vdd gnd cell_6t
Xbit_r16_c144 bl[144] br[144] wl[16] vdd gnd cell_6t
Xbit_r17_c144 bl[144] br[144] wl[17] vdd gnd cell_6t
Xbit_r18_c144 bl[144] br[144] wl[18] vdd gnd cell_6t
Xbit_r19_c144 bl[144] br[144] wl[19] vdd gnd cell_6t
Xbit_r20_c144 bl[144] br[144] wl[20] vdd gnd cell_6t
Xbit_r21_c144 bl[144] br[144] wl[21] vdd gnd cell_6t
Xbit_r22_c144 bl[144] br[144] wl[22] vdd gnd cell_6t
Xbit_r23_c144 bl[144] br[144] wl[23] vdd gnd cell_6t
Xbit_r24_c144 bl[144] br[144] wl[24] vdd gnd cell_6t
Xbit_r25_c144 bl[144] br[144] wl[25] vdd gnd cell_6t
Xbit_r26_c144 bl[144] br[144] wl[26] vdd gnd cell_6t
Xbit_r27_c144 bl[144] br[144] wl[27] vdd gnd cell_6t
Xbit_r28_c144 bl[144] br[144] wl[28] vdd gnd cell_6t
Xbit_r29_c144 bl[144] br[144] wl[29] vdd gnd cell_6t
Xbit_r30_c144 bl[144] br[144] wl[30] vdd gnd cell_6t
Xbit_r31_c144 bl[144] br[144] wl[31] vdd gnd cell_6t
Xbit_r32_c144 bl[144] br[144] wl[32] vdd gnd cell_6t
Xbit_r33_c144 bl[144] br[144] wl[33] vdd gnd cell_6t
Xbit_r34_c144 bl[144] br[144] wl[34] vdd gnd cell_6t
Xbit_r35_c144 bl[144] br[144] wl[35] vdd gnd cell_6t
Xbit_r36_c144 bl[144] br[144] wl[36] vdd gnd cell_6t
Xbit_r37_c144 bl[144] br[144] wl[37] vdd gnd cell_6t
Xbit_r38_c144 bl[144] br[144] wl[38] vdd gnd cell_6t
Xbit_r39_c144 bl[144] br[144] wl[39] vdd gnd cell_6t
Xbit_r40_c144 bl[144] br[144] wl[40] vdd gnd cell_6t
Xbit_r41_c144 bl[144] br[144] wl[41] vdd gnd cell_6t
Xbit_r42_c144 bl[144] br[144] wl[42] vdd gnd cell_6t
Xbit_r43_c144 bl[144] br[144] wl[43] vdd gnd cell_6t
Xbit_r44_c144 bl[144] br[144] wl[44] vdd gnd cell_6t
Xbit_r45_c144 bl[144] br[144] wl[45] vdd gnd cell_6t
Xbit_r46_c144 bl[144] br[144] wl[46] vdd gnd cell_6t
Xbit_r47_c144 bl[144] br[144] wl[47] vdd gnd cell_6t
Xbit_r48_c144 bl[144] br[144] wl[48] vdd gnd cell_6t
Xbit_r49_c144 bl[144] br[144] wl[49] vdd gnd cell_6t
Xbit_r50_c144 bl[144] br[144] wl[50] vdd gnd cell_6t
Xbit_r51_c144 bl[144] br[144] wl[51] vdd gnd cell_6t
Xbit_r52_c144 bl[144] br[144] wl[52] vdd gnd cell_6t
Xbit_r53_c144 bl[144] br[144] wl[53] vdd gnd cell_6t
Xbit_r54_c144 bl[144] br[144] wl[54] vdd gnd cell_6t
Xbit_r55_c144 bl[144] br[144] wl[55] vdd gnd cell_6t
Xbit_r56_c144 bl[144] br[144] wl[56] vdd gnd cell_6t
Xbit_r57_c144 bl[144] br[144] wl[57] vdd gnd cell_6t
Xbit_r58_c144 bl[144] br[144] wl[58] vdd gnd cell_6t
Xbit_r59_c144 bl[144] br[144] wl[59] vdd gnd cell_6t
Xbit_r60_c144 bl[144] br[144] wl[60] vdd gnd cell_6t
Xbit_r61_c144 bl[144] br[144] wl[61] vdd gnd cell_6t
Xbit_r62_c144 bl[144] br[144] wl[62] vdd gnd cell_6t
Xbit_r63_c144 bl[144] br[144] wl[63] vdd gnd cell_6t
Xbit_r64_c144 bl[144] br[144] wl[64] vdd gnd cell_6t
Xbit_r65_c144 bl[144] br[144] wl[65] vdd gnd cell_6t
Xbit_r66_c144 bl[144] br[144] wl[66] vdd gnd cell_6t
Xbit_r67_c144 bl[144] br[144] wl[67] vdd gnd cell_6t
Xbit_r68_c144 bl[144] br[144] wl[68] vdd gnd cell_6t
Xbit_r69_c144 bl[144] br[144] wl[69] vdd gnd cell_6t
Xbit_r70_c144 bl[144] br[144] wl[70] vdd gnd cell_6t
Xbit_r71_c144 bl[144] br[144] wl[71] vdd gnd cell_6t
Xbit_r72_c144 bl[144] br[144] wl[72] vdd gnd cell_6t
Xbit_r73_c144 bl[144] br[144] wl[73] vdd gnd cell_6t
Xbit_r74_c144 bl[144] br[144] wl[74] vdd gnd cell_6t
Xbit_r75_c144 bl[144] br[144] wl[75] vdd gnd cell_6t
Xbit_r76_c144 bl[144] br[144] wl[76] vdd gnd cell_6t
Xbit_r77_c144 bl[144] br[144] wl[77] vdd gnd cell_6t
Xbit_r78_c144 bl[144] br[144] wl[78] vdd gnd cell_6t
Xbit_r79_c144 bl[144] br[144] wl[79] vdd gnd cell_6t
Xbit_r80_c144 bl[144] br[144] wl[80] vdd gnd cell_6t
Xbit_r81_c144 bl[144] br[144] wl[81] vdd gnd cell_6t
Xbit_r82_c144 bl[144] br[144] wl[82] vdd gnd cell_6t
Xbit_r83_c144 bl[144] br[144] wl[83] vdd gnd cell_6t
Xbit_r84_c144 bl[144] br[144] wl[84] vdd gnd cell_6t
Xbit_r85_c144 bl[144] br[144] wl[85] vdd gnd cell_6t
Xbit_r86_c144 bl[144] br[144] wl[86] vdd gnd cell_6t
Xbit_r87_c144 bl[144] br[144] wl[87] vdd gnd cell_6t
Xbit_r88_c144 bl[144] br[144] wl[88] vdd gnd cell_6t
Xbit_r89_c144 bl[144] br[144] wl[89] vdd gnd cell_6t
Xbit_r90_c144 bl[144] br[144] wl[90] vdd gnd cell_6t
Xbit_r91_c144 bl[144] br[144] wl[91] vdd gnd cell_6t
Xbit_r92_c144 bl[144] br[144] wl[92] vdd gnd cell_6t
Xbit_r93_c144 bl[144] br[144] wl[93] vdd gnd cell_6t
Xbit_r94_c144 bl[144] br[144] wl[94] vdd gnd cell_6t
Xbit_r95_c144 bl[144] br[144] wl[95] vdd gnd cell_6t
Xbit_r96_c144 bl[144] br[144] wl[96] vdd gnd cell_6t
Xbit_r97_c144 bl[144] br[144] wl[97] vdd gnd cell_6t
Xbit_r98_c144 bl[144] br[144] wl[98] vdd gnd cell_6t
Xbit_r99_c144 bl[144] br[144] wl[99] vdd gnd cell_6t
Xbit_r100_c144 bl[144] br[144] wl[100] vdd gnd cell_6t
Xbit_r101_c144 bl[144] br[144] wl[101] vdd gnd cell_6t
Xbit_r102_c144 bl[144] br[144] wl[102] vdd gnd cell_6t
Xbit_r103_c144 bl[144] br[144] wl[103] vdd gnd cell_6t
Xbit_r104_c144 bl[144] br[144] wl[104] vdd gnd cell_6t
Xbit_r105_c144 bl[144] br[144] wl[105] vdd gnd cell_6t
Xbit_r106_c144 bl[144] br[144] wl[106] vdd gnd cell_6t
Xbit_r107_c144 bl[144] br[144] wl[107] vdd gnd cell_6t
Xbit_r108_c144 bl[144] br[144] wl[108] vdd gnd cell_6t
Xbit_r109_c144 bl[144] br[144] wl[109] vdd gnd cell_6t
Xbit_r110_c144 bl[144] br[144] wl[110] vdd gnd cell_6t
Xbit_r111_c144 bl[144] br[144] wl[111] vdd gnd cell_6t
Xbit_r112_c144 bl[144] br[144] wl[112] vdd gnd cell_6t
Xbit_r113_c144 bl[144] br[144] wl[113] vdd gnd cell_6t
Xbit_r114_c144 bl[144] br[144] wl[114] vdd gnd cell_6t
Xbit_r115_c144 bl[144] br[144] wl[115] vdd gnd cell_6t
Xbit_r116_c144 bl[144] br[144] wl[116] vdd gnd cell_6t
Xbit_r117_c144 bl[144] br[144] wl[117] vdd gnd cell_6t
Xbit_r118_c144 bl[144] br[144] wl[118] vdd gnd cell_6t
Xbit_r119_c144 bl[144] br[144] wl[119] vdd gnd cell_6t
Xbit_r120_c144 bl[144] br[144] wl[120] vdd gnd cell_6t
Xbit_r121_c144 bl[144] br[144] wl[121] vdd gnd cell_6t
Xbit_r122_c144 bl[144] br[144] wl[122] vdd gnd cell_6t
Xbit_r123_c144 bl[144] br[144] wl[123] vdd gnd cell_6t
Xbit_r124_c144 bl[144] br[144] wl[124] vdd gnd cell_6t
Xbit_r125_c144 bl[144] br[144] wl[125] vdd gnd cell_6t
Xbit_r126_c144 bl[144] br[144] wl[126] vdd gnd cell_6t
Xbit_r127_c144 bl[144] br[144] wl[127] vdd gnd cell_6t
Xbit_r128_c144 bl[144] br[144] wl[128] vdd gnd cell_6t
Xbit_r129_c144 bl[144] br[144] wl[129] vdd gnd cell_6t
Xbit_r130_c144 bl[144] br[144] wl[130] vdd gnd cell_6t
Xbit_r131_c144 bl[144] br[144] wl[131] vdd gnd cell_6t
Xbit_r132_c144 bl[144] br[144] wl[132] vdd gnd cell_6t
Xbit_r133_c144 bl[144] br[144] wl[133] vdd gnd cell_6t
Xbit_r134_c144 bl[144] br[144] wl[134] vdd gnd cell_6t
Xbit_r135_c144 bl[144] br[144] wl[135] vdd gnd cell_6t
Xbit_r136_c144 bl[144] br[144] wl[136] vdd gnd cell_6t
Xbit_r137_c144 bl[144] br[144] wl[137] vdd gnd cell_6t
Xbit_r138_c144 bl[144] br[144] wl[138] vdd gnd cell_6t
Xbit_r139_c144 bl[144] br[144] wl[139] vdd gnd cell_6t
Xbit_r140_c144 bl[144] br[144] wl[140] vdd gnd cell_6t
Xbit_r141_c144 bl[144] br[144] wl[141] vdd gnd cell_6t
Xbit_r142_c144 bl[144] br[144] wl[142] vdd gnd cell_6t
Xbit_r143_c144 bl[144] br[144] wl[143] vdd gnd cell_6t
Xbit_r144_c144 bl[144] br[144] wl[144] vdd gnd cell_6t
Xbit_r145_c144 bl[144] br[144] wl[145] vdd gnd cell_6t
Xbit_r146_c144 bl[144] br[144] wl[146] vdd gnd cell_6t
Xbit_r147_c144 bl[144] br[144] wl[147] vdd gnd cell_6t
Xbit_r148_c144 bl[144] br[144] wl[148] vdd gnd cell_6t
Xbit_r149_c144 bl[144] br[144] wl[149] vdd gnd cell_6t
Xbit_r150_c144 bl[144] br[144] wl[150] vdd gnd cell_6t
Xbit_r151_c144 bl[144] br[144] wl[151] vdd gnd cell_6t
Xbit_r152_c144 bl[144] br[144] wl[152] vdd gnd cell_6t
Xbit_r153_c144 bl[144] br[144] wl[153] vdd gnd cell_6t
Xbit_r154_c144 bl[144] br[144] wl[154] vdd gnd cell_6t
Xbit_r155_c144 bl[144] br[144] wl[155] vdd gnd cell_6t
Xbit_r156_c144 bl[144] br[144] wl[156] vdd gnd cell_6t
Xbit_r157_c144 bl[144] br[144] wl[157] vdd gnd cell_6t
Xbit_r158_c144 bl[144] br[144] wl[158] vdd gnd cell_6t
Xbit_r159_c144 bl[144] br[144] wl[159] vdd gnd cell_6t
Xbit_r160_c144 bl[144] br[144] wl[160] vdd gnd cell_6t
Xbit_r161_c144 bl[144] br[144] wl[161] vdd gnd cell_6t
Xbit_r162_c144 bl[144] br[144] wl[162] vdd gnd cell_6t
Xbit_r163_c144 bl[144] br[144] wl[163] vdd gnd cell_6t
Xbit_r164_c144 bl[144] br[144] wl[164] vdd gnd cell_6t
Xbit_r165_c144 bl[144] br[144] wl[165] vdd gnd cell_6t
Xbit_r166_c144 bl[144] br[144] wl[166] vdd gnd cell_6t
Xbit_r167_c144 bl[144] br[144] wl[167] vdd gnd cell_6t
Xbit_r168_c144 bl[144] br[144] wl[168] vdd gnd cell_6t
Xbit_r169_c144 bl[144] br[144] wl[169] vdd gnd cell_6t
Xbit_r170_c144 bl[144] br[144] wl[170] vdd gnd cell_6t
Xbit_r171_c144 bl[144] br[144] wl[171] vdd gnd cell_6t
Xbit_r172_c144 bl[144] br[144] wl[172] vdd gnd cell_6t
Xbit_r173_c144 bl[144] br[144] wl[173] vdd gnd cell_6t
Xbit_r174_c144 bl[144] br[144] wl[174] vdd gnd cell_6t
Xbit_r175_c144 bl[144] br[144] wl[175] vdd gnd cell_6t
Xbit_r176_c144 bl[144] br[144] wl[176] vdd gnd cell_6t
Xbit_r177_c144 bl[144] br[144] wl[177] vdd gnd cell_6t
Xbit_r178_c144 bl[144] br[144] wl[178] vdd gnd cell_6t
Xbit_r179_c144 bl[144] br[144] wl[179] vdd gnd cell_6t
Xbit_r180_c144 bl[144] br[144] wl[180] vdd gnd cell_6t
Xbit_r181_c144 bl[144] br[144] wl[181] vdd gnd cell_6t
Xbit_r182_c144 bl[144] br[144] wl[182] vdd gnd cell_6t
Xbit_r183_c144 bl[144] br[144] wl[183] vdd gnd cell_6t
Xbit_r184_c144 bl[144] br[144] wl[184] vdd gnd cell_6t
Xbit_r185_c144 bl[144] br[144] wl[185] vdd gnd cell_6t
Xbit_r186_c144 bl[144] br[144] wl[186] vdd gnd cell_6t
Xbit_r187_c144 bl[144] br[144] wl[187] vdd gnd cell_6t
Xbit_r188_c144 bl[144] br[144] wl[188] vdd gnd cell_6t
Xbit_r189_c144 bl[144] br[144] wl[189] vdd gnd cell_6t
Xbit_r190_c144 bl[144] br[144] wl[190] vdd gnd cell_6t
Xbit_r191_c144 bl[144] br[144] wl[191] vdd gnd cell_6t
Xbit_r192_c144 bl[144] br[144] wl[192] vdd gnd cell_6t
Xbit_r193_c144 bl[144] br[144] wl[193] vdd gnd cell_6t
Xbit_r194_c144 bl[144] br[144] wl[194] vdd gnd cell_6t
Xbit_r195_c144 bl[144] br[144] wl[195] vdd gnd cell_6t
Xbit_r196_c144 bl[144] br[144] wl[196] vdd gnd cell_6t
Xbit_r197_c144 bl[144] br[144] wl[197] vdd gnd cell_6t
Xbit_r198_c144 bl[144] br[144] wl[198] vdd gnd cell_6t
Xbit_r199_c144 bl[144] br[144] wl[199] vdd gnd cell_6t
Xbit_r200_c144 bl[144] br[144] wl[200] vdd gnd cell_6t
Xbit_r201_c144 bl[144] br[144] wl[201] vdd gnd cell_6t
Xbit_r202_c144 bl[144] br[144] wl[202] vdd gnd cell_6t
Xbit_r203_c144 bl[144] br[144] wl[203] vdd gnd cell_6t
Xbit_r204_c144 bl[144] br[144] wl[204] vdd gnd cell_6t
Xbit_r205_c144 bl[144] br[144] wl[205] vdd gnd cell_6t
Xbit_r206_c144 bl[144] br[144] wl[206] vdd gnd cell_6t
Xbit_r207_c144 bl[144] br[144] wl[207] vdd gnd cell_6t
Xbit_r208_c144 bl[144] br[144] wl[208] vdd gnd cell_6t
Xbit_r209_c144 bl[144] br[144] wl[209] vdd gnd cell_6t
Xbit_r210_c144 bl[144] br[144] wl[210] vdd gnd cell_6t
Xbit_r211_c144 bl[144] br[144] wl[211] vdd gnd cell_6t
Xbit_r212_c144 bl[144] br[144] wl[212] vdd gnd cell_6t
Xbit_r213_c144 bl[144] br[144] wl[213] vdd gnd cell_6t
Xbit_r214_c144 bl[144] br[144] wl[214] vdd gnd cell_6t
Xbit_r215_c144 bl[144] br[144] wl[215] vdd gnd cell_6t
Xbit_r216_c144 bl[144] br[144] wl[216] vdd gnd cell_6t
Xbit_r217_c144 bl[144] br[144] wl[217] vdd gnd cell_6t
Xbit_r218_c144 bl[144] br[144] wl[218] vdd gnd cell_6t
Xbit_r219_c144 bl[144] br[144] wl[219] vdd gnd cell_6t
Xbit_r220_c144 bl[144] br[144] wl[220] vdd gnd cell_6t
Xbit_r221_c144 bl[144] br[144] wl[221] vdd gnd cell_6t
Xbit_r222_c144 bl[144] br[144] wl[222] vdd gnd cell_6t
Xbit_r223_c144 bl[144] br[144] wl[223] vdd gnd cell_6t
Xbit_r224_c144 bl[144] br[144] wl[224] vdd gnd cell_6t
Xbit_r225_c144 bl[144] br[144] wl[225] vdd gnd cell_6t
Xbit_r226_c144 bl[144] br[144] wl[226] vdd gnd cell_6t
Xbit_r227_c144 bl[144] br[144] wl[227] vdd gnd cell_6t
Xbit_r228_c144 bl[144] br[144] wl[228] vdd gnd cell_6t
Xbit_r229_c144 bl[144] br[144] wl[229] vdd gnd cell_6t
Xbit_r230_c144 bl[144] br[144] wl[230] vdd gnd cell_6t
Xbit_r231_c144 bl[144] br[144] wl[231] vdd gnd cell_6t
Xbit_r232_c144 bl[144] br[144] wl[232] vdd gnd cell_6t
Xbit_r233_c144 bl[144] br[144] wl[233] vdd gnd cell_6t
Xbit_r234_c144 bl[144] br[144] wl[234] vdd gnd cell_6t
Xbit_r235_c144 bl[144] br[144] wl[235] vdd gnd cell_6t
Xbit_r236_c144 bl[144] br[144] wl[236] vdd gnd cell_6t
Xbit_r237_c144 bl[144] br[144] wl[237] vdd gnd cell_6t
Xbit_r238_c144 bl[144] br[144] wl[238] vdd gnd cell_6t
Xbit_r239_c144 bl[144] br[144] wl[239] vdd gnd cell_6t
Xbit_r240_c144 bl[144] br[144] wl[240] vdd gnd cell_6t
Xbit_r241_c144 bl[144] br[144] wl[241] vdd gnd cell_6t
Xbit_r242_c144 bl[144] br[144] wl[242] vdd gnd cell_6t
Xbit_r243_c144 bl[144] br[144] wl[243] vdd gnd cell_6t
Xbit_r244_c144 bl[144] br[144] wl[244] vdd gnd cell_6t
Xbit_r245_c144 bl[144] br[144] wl[245] vdd gnd cell_6t
Xbit_r246_c144 bl[144] br[144] wl[246] vdd gnd cell_6t
Xbit_r247_c144 bl[144] br[144] wl[247] vdd gnd cell_6t
Xbit_r248_c144 bl[144] br[144] wl[248] vdd gnd cell_6t
Xbit_r249_c144 bl[144] br[144] wl[249] vdd gnd cell_6t
Xbit_r250_c144 bl[144] br[144] wl[250] vdd gnd cell_6t
Xbit_r251_c144 bl[144] br[144] wl[251] vdd gnd cell_6t
Xbit_r252_c144 bl[144] br[144] wl[252] vdd gnd cell_6t
Xbit_r253_c144 bl[144] br[144] wl[253] vdd gnd cell_6t
Xbit_r254_c144 bl[144] br[144] wl[254] vdd gnd cell_6t
Xbit_r255_c144 bl[144] br[144] wl[255] vdd gnd cell_6t
Xbit_r0_c145 bl[145] br[145] wl[0] vdd gnd cell_6t
Xbit_r1_c145 bl[145] br[145] wl[1] vdd gnd cell_6t
Xbit_r2_c145 bl[145] br[145] wl[2] vdd gnd cell_6t
Xbit_r3_c145 bl[145] br[145] wl[3] vdd gnd cell_6t
Xbit_r4_c145 bl[145] br[145] wl[4] vdd gnd cell_6t
Xbit_r5_c145 bl[145] br[145] wl[5] vdd gnd cell_6t
Xbit_r6_c145 bl[145] br[145] wl[6] vdd gnd cell_6t
Xbit_r7_c145 bl[145] br[145] wl[7] vdd gnd cell_6t
Xbit_r8_c145 bl[145] br[145] wl[8] vdd gnd cell_6t
Xbit_r9_c145 bl[145] br[145] wl[9] vdd gnd cell_6t
Xbit_r10_c145 bl[145] br[145] wl[10] vdd gnd cell_6t
Xbit_r11_c145 bl[145] br[145] wl[11] vdd gnd cell_6t
Xbit_r12_c145 bl[145] br[145] wl[12] vdd gnd cell_6t
Xbit_r13_c145 bl[145] br[145] wl[13] vdd gnd cell_6t
Xbit_r14_c145 bl[145] br[145] wl[14] vdd gnd cell_6t
Xbit_r15_c145 bl[145] br[145] wl[15] vdd gnd cell_6t
Xbit_r16_c145 bl[145] br[145] wl[16] vdd gnd cell_6t
Xbit_r17_c145 bl[145] br[145] wl[17] vdd gnd cell_6t
Xbit_r18_c145 bl[145] br[145] wl[18] vdd gnd cell_6t
Xbit_r19_c145 bl[145] br[145] wl[19] vdd gnd cell_6t
Xbit_r20_c145 bl[145] br[145] wl[20] vdd gnd cell_6t
Xbit_r21_c145 bl[145] br[145] wl[21] vdd gnd cell_6t
Xbit_r22_c145 bl[145] br[145] wl[22] vdd gnd cell_6t
Xbit_r23_c145 bl[145] br[145] wl[23] vdd gnd cell_6t
Xbit_r24_c145 bl[145] br[145] wl[24] vdd gnd cell_6t
Xbit_r25_c145 bl[145] br[145] wl[25] vdd gnd cell_6t
Xbit_r26_c145 bl[145] br[145] wl[26] vdd gnd cell_6t
Xbit_r27_c145 bl[145] br[145] wl[27] vdd gnd cell_6t
Xbit_r28_c145 bl[145] br[145] wl[28] vdd gnd cell_6t
Xbit_r29_c145 bl[145] br[145] wl[29] vdd gnd cell_6t
Xbit_r30_c145 bl[145] br[145] wl[30] vdd gnd cell_6t
Xbit_r31_c145 bl[145] br[145] wl[31] vdd gnd cell_6t
Xbit_r32_c145 bl[145] br[145] wl[32] vdd gnd cell_6t
Xbit_r33_c145 bl[145] br[145] wl[33] vdd gnd cell_6t
Xbit_r34_c145 bl[145] br[145] wl[34] vdd gnd cell_6t
Xbit_r35_c145 bl[145] br[145] wl[35] vdd gnd cell_6t
Xbit_r36_c145 bl[145] br[145] wl[36] vdd gnd cell_6t
Xbit_r37_c145 bl[145] br[145] wl[37] vdd gnd cell_6t
Xbit_r38_c145 bl[145] br[145] wl[38] vdd gnd cell_6t
Xbit_r39_c145 bl[145] br[145] wl[39] vdd gnd cell_6t
Xbit_r40_c145 bl[145] br[145] wl[40] vdd gnd cell_6t
Xbit_r41_c145 bl[145] br[145] wl[41] vdd gnd cell_6t
Xbit_r42_c145 bl[145] br[145] wl[42] vdd gnd cell_6t
Xbit_r43_c145 bl[145] br[145] wl[43] vdd gnd cell_6t
Xbit_r44_c145 bl[145] br[145] wl[44] vdd gnd cell_6t
Xbit_r45_c145 bl[145] br[145] wl[45] vdd gnd cell_6t
Xbit_r46_c145 bl[145] br[145] wl[46] vdd gnd cell_6t
Xbit_r47_c145 bl[145] br[145] wl[47] vdd gnd cell_6t
Xbit_r48_c145 bl[145] br[145] wl[48] vdd gnd cell_6t
Xbit_r49_c145 bl[145] br[145] wl[49] vdd gnd cell_6t
Xbit_r50_c145 bl[145] br[145] wl[50] vdd gnd cell_6t
Xbit_r51_c145 bl[145] br[145] wl[51] vdd gnd cell_6t
Xbit_r52_c145 bl[145] br[145] wl[52] vdd gnd cell_6t
Xbit_r53_c145 bl[145] br[145] wl[53] vdd gnd cell_6t
Xbit_r54_c145 bl[145] br[145] wl[54] vdd gnd cell_6t
Xbit_r55_c145 bl[145] br[145] wl[55] vdd gnd cell_6t
Xbit_r56_c145 bl[145] br[145] wl[56] vdd gnd cell_6t
Xbit_r57_c145 bl[145] br[145] wl[57] vdd gnd cell_6t
Xbit_r58_c145 bl[145] br[145] wl[58] vdd gnd cell_6t
Xbit_r59_c145 bl[145] br[145] wl[59] vdd gnd cell_6t
Xbit_r60_c145 bl[145] br[145] wl[60] vdd gnd cell_6t
Xbit_r61_c145 bl[145] br[145] wl[61] vdd gnd cell_6t
Xbit_r62_c145 bl[145] br[145] wl[62] vdd gnd cell_6t
Xbit_r63_c145 bl[145] br[145] wl[63] vdd gnd cell_6t
Xbit_r64_c145 bl[145] br[145] wl[64] vdd gnd cell_6t
Xbit_r65_c145 bl[145] br[145] wl[65] vdd gnd cell_6t
Xbit_r66_c145 bl[145] br[145] wl[66] vdd gnd cell_6t
Xbit_r67_c145 bl[145] br[145] wl[67] vdd gnd cell_6t
Xbit_r68_c145 bl[145] br[145] wl[68] vdd gnd cell_6t
Xbit_r69_c145 bl[145] br[145] wl[69] vdd gnd cell_6t
Xbit_r70_c145 bl[145] br[145] wl[70] vdd gnd cell_6t
Xbit_r71_c145 bl[145] br[145] wl[71] vdd gnd cell_6t
Xbit_r72_c145 bl[145] br[145] wl[72] vdd gnd cell_6t
Xbit_r73_c145 bl[145] br[145] wl[73] vdd gnd cell_6t
Xbit_r74_c145 bl[145] br[145] wl[74] vdd gnd cell_6t
Xbit_r75_c145 bl[145] br[145] wl[75] vdd gnd cell_6t
Xbit_r76_c145 bl[145] br[145] wl[76] vdd gnd cell_6t
Xbit_r77_c145 bl[145] br[145] wl[77] vdd gnd cell_6t
Xbit_r78_c145 bl[145] br[145] wl[78] vdd gnd cell_6t
Xbit_r79_c145 bl[145] br[145] wl[79] vdd gnd cell_6t
Xbit_r80_c145 bl[145] br[145] wl[80] vdd gnd cell_6t
Xbit_r81_c145 bl[145] br[145] wl[81] vdd gnd cell_6t
Xbit_r82_c145 bl[145] br[145] wl[82] vdd gnd cell_6t
Xbit_r83_c145 bl[145] br[145] wl[83] vdd gnd cell_6t
Xbit_r84_c145 bl[145] br[145] wl[84] vdd gnd cell_6t
Xbit_r85_c145 bl[145] br[145] wl[85] vdd gnd cell_6t
Xbit_r86_c145 bl[145] br[145] wl[86] vdd gnd cell_6t
Xbit_r87_c145 bl[145] br[145] wl[87] vdd gnd cell_6t
Xbit_r88_c145 bl[145] br[145] wl[88] vdd gnd cell_6t
Xbit_r89_c145 bl[145] br[145] wl[89] vdd gnd cell_6t
Xbit_r90_c145 bl[145] br[145] wl[90] vdd gnd cell_6t
Xbit_r91_c145 bl[145] br[145] wl[91] vdd gnd cell_6t
Xbit_r92_c145 bl[145] br[145] wl[92] vdd gnd cell_6t
Xbit_r93_c145 bl[145] br[145] wl[93] vdd gnd cell_6t
Xbit_r94_c145 bl[145] br[145] wl[94] vdd gnd cell_6t
Xbit_r95_c145 bl[145] br[145] wl[95] vdd gnd cell_6t
Xbit_r96_c145 bl[145] br[145] wl[96] vdd gnd cell_6t
Xbit_r97_c145 bl[145] br[145] wl[97] vdd gnd cell_6t
Xbit_r98_c145 bl[145] br[145] wl[98] vdd gnd cell_6t
Xbit_r99_c145 bl[145] br[145] wl[99] vdd gnd cell_6t
Xbit_r100_c145 bl[145] br[145] wl[100] vdd gnd cell_6t
Xbit_r101_c145 bl[145] br[145] wl[101] vdd gnd cell_6t
Xbit_r102_c145 bl[145] br[145] wl[102] vdd gnd cell_6t
Xbit_r103_c145 bl[145] br[145] wl[103] vdd gnd cell_6t
Xbit_r104_c145 bl[145] br[145] wl[104] vdd gnd cell_6t
Xbit_r105_c145 bl[145] br[145] wl[105] vdd gnd cell_6t
Xbit_r106_c145 bl[145] br[145] wl[106] vdd gnd cell_6t
Xbit_r107_c145 bl[145] br[145] wl[107] vdd gnd cell_6t
Xbit_r108_c145 bl[145] br[145] wl[108] vdd gnd cell_6t
Xbit_r109_c145 bl[145] br[145] wl[109] vdd gnd cell_6t
Xbit_r110_c145 bl[145] br[145] wl[110] vdd gnd cell_6t
Xbit_r111_c145 bl[145] br[145] wl[111] vdd gnd cell_6t
Xbit_r112_c145 bl[145] br[145] wl[112] vdd gnd cell_6t
Xbit_r113_c145 bl[145] br[145] wl[113] vdd gnd cell_6t
Xbit_r114_c145 bl[145] br[145] wl[114] vdd gnd cell_6t
Xbit_r115_c145 bl[145] br[145] wl[115] vdd gnd cell_6t
Xbit_r116_c145 bl[145] br[145] wl[116] vdd gnd cell_6t
Xbit_r117_c145 bl[145] br[145] wl[117] vdd gnd cell_6t
Xbit_r118_c145 bl[145] br[145] wl[118] vdd gnd cell_6t
Xbit_r119_c145 bl[145] br[145] wl[119] vdd gnd cell_6t
Xbit_r120_c145 bl[145] br[145] wl[120] vdd gnd cell_6t
Xbit_r121_c145 bl[145] br[145] wl[121] vdd gnd cell_6t
Xbit_r122_c145 bl[145] br[145] wl[122] vdd gnd cell_6t
Xbit_r123_c145 bl[145] br[145] wl[123] vdd gnd cell_6t
Xbit_r124_c145 bl[145] br[145] wl[124] vdd gnd cell_6t
Xbit_r125_c145 bl[145] br[145] wl[125] vdd gnd cell_6t
Xbit_r126_c145 bl[145] br[145] wl[126] vdd gnd cell_6t
Xbit_r127_c145 bl[145] br[145] wl[127] vdd gnd cell_6t
Xbit_r128_c145 bl[145] br[145] wl[128] vdd gnd cell_6t
Xbit_r129_c145 bl[145] br[145] wl[129] vdd gnd cell_6t
Xbit_r130_c145 bl[145] br[145] wl[130] vdd gnd cell_6t
Xbit_r131_c145 bl[145] br[145] wl[131] vdd gnd cell_6t
Xbit_r132_c145 bl[145] br[145] wl[132] vdd gnd cell_6t
Xbit_r133_c145 bl[145] br[145] wl[133] vdd gnd cell_6t
Xbit_r134_c145 bl[145] br[145] wl[134] vdd gnd cell_6t
Xbit_r135_c145 bl[145] br[145] wl[135] vdd gnd cell_6t
Xbit_r136_c145 bl[145] br[145] wl[136] vdd gnd cell_6t
Xbit_r137_c145 bl[145] br[145] wl[137] vdd gnd cell_6t
Xbit_r138_c145 bl[145] br[145] wl[138] vdd gnd cell_6t
Xbit_r139_c145 bl[145] br[145] wl[139] vdd gnd cell_6t
Xbit_r140_c145 bl[145] br[145] wl[140] vdd gnd cell_6t
Xbit_r141_c145 bl[145] br[145] wl[141] vdd gnd cell_6t
Xbit_r142_c145 bl[145] br[145] wl[142] vdd gnd cell_6t
Xbit_r143_c145 bl[145] br[145] wl[143] vdd gnd cell_6t
Xbit_r144_c145 bl[145] br[145] wl[144] vdd gnd cell_6t
Xbit_r145_c145 bl[145] br[145] wl[145] vdd gnd cell_6t
Xbit_r146_c145 bl[145] br[145] wl[146] vdd gnd cell_6t
Xbit_r147_c145 bl[145] br[145] wl[147] vdd gnd cell_6t
Xbit_r148_c145 bl[145] br[145] wl[148] vdd gnd cell_6t
Xbit_r149_c145 bl[145] br[145] wl[149] vdd gnd cell_6t
Xbit_r150_c145 bl[145] br[145] wl[150] vdd gnd cell_6t
Xbit_r151_c145 bl[145] br[145] wl[151] vdd gnd cell_6t
Xbit_r152_c145 bl[145] br[145] wl[152] vdd gnd cell_6t
Xbit_r153_c145 bl[145] br[145] wl[153] vdd gnd cell_6t
Xbit_r154_c145 bl[145] br[145] wl[154] vdd gnd cell_6t
Xbit_r155_c145 bl[145] br[145] wl[155] vdd gnd cell_6t
Xbit_r156_c145 bl[145] br[145] wl[156] vdd gnd cell_6t
Xbit_r157_c145 bl[145] br[145] wl[157] vdd gnd cell_6t
Xbit_r158_c145 bl[145] br[145] wl[158] vdd gnd cell_6t
Xbit_r159_c145 bl[145] br[145] wl[159] vdd gnd cell_6t
Xbit_r160_c145 bl[145] br[145] wl[160] vdd gnd cell_6t
Xbit_r161_c145 bl[145] br[145] wl[161] vdd gnd cell_6t
Xbit_r162_c145 bl[145] br[145] wl[162] vdd gnd cell_6t
Xbit_r163_c145 bl[145] br[145] wl[163] vdd gnd cell_6t
Xbit_r164_c145 bl[145] br[145] wl[164] vdd gnd cell_6t
Xbit_r165_c145 bl[145] br[145] wl[165] vdd gnd cell_6t
Xbit_r166_c145 bl[145] br[145] wl[166] vdd gnd cell_6t
Xbit_r167_c145 bl[145] br[145] wl[167] vdd gnd cell_6t
Xbit_r168_c145 bl[145] br[145] wl[168] vdd gnd cell_6t
Xbit_r169_c145 bl[145] br[145] wl[169] vdd gnd cell_6t
Xbit_r170_c145 bl[145] br[145] wl[170] vdd gnd cell_6t
Xbit_r171_c145 bl[145] br[145] wl[171] vdd gnd cell_6t
Xbit_r172_c145 bl[145] br[145] wl[172] vdd gnd cell_6t
Xbit_r173_c145 bl[145] br[145] wl[173] vdd gnd cell_6t
Xbit_r174_c145 bl[145] br[145] wl[174] vdd gnd cell_6t
Xbit_r175_c145 bl[145] br[145] wl[175] vdd gnd cell_6t
Xbit_r176_c145 bl[145] br[145] wl[176] vdd gnd cell_6t
Xbit_r177_c145 bl[145] br[145] wl[177] vdd gnd cell_6t
Xbit_r178_c145 bl[145] br[145] wl[178] vdd gnd cell_6t
Xbit_r179_c145 bl[145] br[145] wl[179] vdd gnd cell_6t
Xbit_r180_c145 bl[145] br[145] wl[180] vdd gnd cell_6t
Xbit_r181_c145 bl[145] br[145] wl[181] vdd gnd cell_6t
Xbit_r182_c145 bl[145] br[145] wl[182] vdd gnd cell_6t
Xbit_r183_c145 bl[145] br[145] wl[183] vdd gnd cell_6t
Xbit_r184_c145 bl[145] br[145] wl[184] vdd gnd cell_6t
Xbit_r185_c145 bl[145] br[145] wl[185] vdd gnd cell_6t
Xbit_r186_c145 bl[145] br[145] wl[186] vdd gnd cell_6t
Xbit_r187_c145 bl[145] br[145] wl[187] vdd gnd cell_6t
Xbit_r188_c145 bl[145] br[145] wl[188] vdd gnd cell_6t
Xbit_r189_c145 bl[145] br[145] wl[189] vdd gnd cell_6t
Xbit_r190_c145 bl[145] br[145] wl[190] vdd gnd cell_6t
Xbit_r191_c145 bl[145] br[145] wl[191] vdd gnd cell_6t
Xbit_r192_c145 bl[145] br[145] wl[192] vdd gnd cell_6t
Xbit_r193_c145 bl[145] br[145] wl[193] vdd gnd cell_6t
Xbit_r194_c145 bl[145] br[145] wl[194] vdd gnd cell_6t
Xbit_r195_c145 bl[145] br[145] wl[195] vdd gnd cell_6t
Xbit_r196_c145 bl[145] br[145] wl[196] vdd gnd cell_6t
Xbit_r197_c145 bl[145] br[145] wl[197] vdd gnd cell_6t
Xbit_r198_c145 bl[145] br[145] wl[198] vdd gnd cell_6t
Xbit_r199_c145 bl[145] br[145] wl[199] vdd gnd cell_6t
Xbit_r200_c145 bl[145] br[145] wl[200] vdd gnd cell_6t
Xbit_r201_c145 bl[145] br[145] wl[201] vdd gnd cell_6t
Xbit_r202_c145 bl[145] br[145] wl[202] vdd gnd cell_6t
Xbit_r203_c145 bl[145] br[145] wl[203] vdd gnd cell_6t
Xbit_r204_c145 bl[145] br[145] wl[204] vdd gnd cell_6t
Xbit_r205_c145 bl[145] br[145] wl[205] vdd gnd cell_6t
Xbit_r206_c145 bl[145] br[145] wl[206] vdd gnd cell_6t
Xbit_r207_c145 bl[145] br[145] wl[207] vdd gnd cell_6t
Xbit_r208_c145 bl[145] br[145] wl[208] vdd gnd cell_6t
Xbit_r209_c145 bl[145] br[145] wl[209] vdd gnd cell_6t
Xbit_r210_c145 bl[145] br[145] wl[210] vdd gnd cell_6t
Xbit_r211_c145 bl[145] br[145] wl[211] vdd gnd cell_6t
Xbit_r212_c145 bl[145] br[145] wl[212] vdd gnd cell_6t
Xbit_r213_c145 bl[145] br[145] wl[213] vdd gnd cell_6t
Xbit_r214_c145 bl[145] br[145] wl[214] vdd gnd cell_6t
Xbit_r215_c145 bl[145] br[145] wl[215] vdd gnd cell_6t
Xbit_r216_c145 bl[145] br[145] wl[216] vdd gnd cell_6t
Xbit_r217_c145 bl[145] br[145] wl[217] vdd gnd cell_6t
Xbit_r218_c145 bl[145] br[145] wl[218] vdd gnd cell_6t
Xbit_r219_c145 bl[145] br[145] wl[219] vdd gnd cell_6t
Xbit_r220_c145 bl[145] br[145] wl[220] vdd gnd cell_6t
Xbit_r221_c145 bl[145] br[145] wl[221] vdd gnd cell_6t
Xbit_r222_c145 bl[145] br[145] wl[222] vdd gnd cell_6t
Xbit_r223_c145 bl[145] br[145] wl[223] vdd gnd cell_6t
Xbit_r224_c145 bl[145] br[145] wl[224] vdd gnd cell_6t
Xbit_r225_c145 bl[145] br[145] wl[225] vdd gnd cell_6t
Xbit_r226_c145 bl[145] br[145] wl[226] vdd gnd cell_6t
Xbit_r227_c145 bl[145] br[145] wl[227] vdd gnd cell_6t
Xbit_r228_c145 bl[145] br[145] wl[228] vdd gnd cell_6t
Xbit_r229_c145 bl[145] br[145] wl[229] vdd gnd cell_6t
Xbit_r230_c145 bl[145] br[145] wl[230] vdd gnd cell_6t
Xbit_r231_c145 bl[145] br[145] wl[231] vdd gnd cell_6t
Xbit_r232_c145 bl[145] br[145] wl[232] vdd gnd cell_6t
Xbit_r233_c145 bl[145] br[145] wl[233] vdd gnd cell_6t
Xbit_r234_c145 bl[145] br[145] wl[234] vdd gnd cell_6t
Xbit_r235_c145 bl[145] br[145] wl[235] vdd gnd cell_6t
Xbit_r236_c145 bl[145] br[145] wl[236] vdd gnd cell_6t
Xbit_r237_c145 bl[145] br[145] wl[237] vdd gnd cell_6t
Xbit_r238_c145 bl[145] br[145] wl[238] vdd gnd cell_6t
Xbit_r239_c145 bl[145] br[145] wl[239] vdd gnd cell_6t
Xbit_r240_c145 bl[145] br[145] wl[240] vdd gnd cell_6t
Xbit_r241_c145 bl[145] br[145] wl[241] vdd gnd cell_6t
Xbit_r242_c145 bl[145] br[145] wl[242] vdd gnd cell_6t
Xbit_r243_c145 bl[145] br[145] wl[243] vdd gnd cell_6t
Xbit_r244_c145 bl[145] br[145] wl[244] vdd gnd cell_6t
Xbit_r245_c145 bl[145] br[145] wl[245] vdd gnd cell_6t
Xbit_r246_c145 bl[145] br[145] wl[246] vdd gnd cell_6t
Xbit_r247_c145 bl[145] br[145] wl[247] vdd gnd cell_6t
Xbit_r248_c145 bl[145] br[145] wl[248] vdd gnd cell_6t
Xbit_r249_c145 bl[145] br[145] wl[249] vdd gnd cell_6t
Xbit_r250_c145 bl[145] br[145] wl[250] vdd gnd cell_6t
Xbit_r251_c145 bl[145] br[145] wl[251] vdd gnd cell_6t
Xbit_r252_c145 bl[145] br[145] wl[252] vdd gnd cell_6t
Xbit_r253_c145 bl[145] br[145] wl[253] vdd gnd cell_6t
Xbit_r254_c145 bl[145] br[145] wl[254] vdd gnd cell_6t
Xbit_r255_c145 bl[145] br[145] wl[255] vdd gnd cell_6t
Xbit_r0_c146 bl[146] br[146] wl[0] vdd gnd cell_6t
Xbit_r1_c146 bl[146] br[146] wl[1] vdd gnd cell_6t
Xbit_r2_c146 bl[146] br[146] wl[2] vdd gnd cell_6t
Xbit_r3_c146 bl[146] br[146] wl[3] vdd gnd cell_6t
Xbit_r4_c146 bl[146] br[146] wl[4] vdd gnd cell_6t
Xbit_r5_c146 bl[146] br[146] wl[5] vdd gnd cell_6t
Xbit_r6_c146 bl[146] br[146] wl[6] vdd gnd cell_6t
Xbit_r7_c146 bl[146] br[146] wl[7] vdd gnd cell_6t
Xbit_r8_c146 bl[146] br[146] wl[8] vdd gnd cell_6t
Xbit_r9_c146 bl[146] br[146] wl[9] vdd gnd cell_6t
Xbit_r10_c146 bl[146] br[146] wl[10] vdd gnd cell_6t
Xbit_r11_c146 bl[146] br[146] wl[11] vdd gnd cell_6t
Xbit_r12_c146 bl[146] br[146] wl[12] vdd gnd cell_6t
Xbit_r13_c146 bl[146] br[146] wl[13] vdd gnd cell_6t
Xbit_r14_c146 bl[146] br[146] wl[14] vdd gnd cell_6t
Xbit_r15_c146 bl[146] br[146] wl[15] vdd gnd cell_6t
Xbit_r16_c146 bl[146] br[146] wl[16] vdd gnd cell_6t
Xbit_r17_c146 bl[146] br[146] wl[17] vdd gnd cell_6t
Xbit_r18_c146 bl[146] br[146] wl[18] vdd gnd cell_6t
Xbit_r19_c146 bl[146] br[146] wl[19] vdd gnd cell_6t
Xbit_r20_c146 bl[146] br[146] wl[20] vdd gnd cell_6t
Xbit_r21_c146 bl[146] br[146] wl[21] vdd gnd cell_6t
Xbit_r22_c146 bl[146] br[146] wl[22] vdd gnd cell_6t
Xbit_r23_c146 bl[146] br[146] wl[23] vdd gnd cell_6t
Xbit_r24_c146 bl[146] br[146] wl[24] vdd gnd cell_6t
Xbit_r25_c146 bl[146] br[146] wl[25] vdd gnd cell_6t
Xbit_r26_c146 bl[146] br[146] wl[26] vdd gnd cell_6t
Xbit_r27_c146 bl[146] br[146] wl[27] vdd gnd cell_6t
Xbit_r28_c146 bl[146] br[146] wl[28] vdd gnd cell_6t
Xbit_r29_c146 bl[146] br[146] wl[29] vdd gnd cell_6t
Xbit_r30_c146 bl[146] br[146] wl[30] vdd gnd cell_6t
Xbit_r31_c146 bl[146] br[146] wl[31] vdd gnd cell_6t
Xbit_r32_c146 bl[146] br[146] wl[32] vdd gnd cell_6t
Xbit_r33_c146 bl[146] br[146] wl[33] vdd gnd cell_6t
Xbit_r34_c146 bl[146] br[146] wl[34] vdd gnd cell_6t
Xbit_r35_c146 bl[146] br[146] wl[35] vdd gnd cell_6t
Xbit_r36_c146 bl[146] br[146] wl[36] vdd gnd cell_6t
Xbit_r37_c146 bl[146] br[146] wl[37] vdd gnd cell_6t
Xbit_r38_c146 bl[146] br[146] wl[38] vdd gnd cell_6t
Xbit_r39_c146 bl[146] br[146] wl[39] vdd gnd cell_6t
Xbit_r40_c146 bl[146] br[146] wl[40] vdd gnd cell_6t
Xbit_r41_c146 bl[146] br[146] wl[41] vdd gnd cell_6t
Xbit_r42_c146 bl[146] br[146] wl[42] vdd gnd cell_6t
Xbit_r43_c146 bl[146] br[146] wl[43] vdd gnd cell_6t
Xbit_r44_c146 bl[146] br[146] wl[44] vdd gnd cell_6t
Xbit_r45_c146 bl[146] br[146] wl[45] vdd gnd cell_6t
Xbit_r46_c146 bl[146] br[146] wl[46] vdd gnd cell_6t
Xbit_r47_c146 bl[146] br[146] wl[47] vdd gnd cell_6t
Xbit_r48_c146 bl[146] br[146] wl[48] vdd gnd cell_6t
Xbit_r49_c146 bl[146] br[146] wl[49] vdd gnd cell_6t
Xbit_r50_c146 bl[146] br[146] wl[50] vdd gnd cell_6t
Xbit_r51_c146 bl[146] br[146] wl[51] vdd gnd cell_6t
Xbit_r52_c146 bl[146] br[146] wl[52] vdd gnd cell_6t
Xbit_r53_c146 bl[146] br[146] wl[53] vdd gnd cell_6t
Xbit_r54_c146 bl[146] br[146] wl[54] vdd gnd cell_6t
Xbit_r55_c146 bl[146] br[146] wl[55] vdd gnd cell_6t
Xbit_r56_c146 bl[146] br[146] wl[56] vdd gnd cell_6t
Xbit_r57_c146 bl[146] br[146] wl[57] vdd gnd cell_6t
Xbit_r58_c146 bl[146] br[146] wl[58] vdd gnd cell_6t
Xbit_r59_c146 bl[146] br[146] wl[59] vdd gnd cell_6t
Xbit_r60_c146 bl[146] br[146] wl[60] vdd gnd cell_6t
Xbit_r61_c146 bl[146] br[146] wl[61] vdd gnd cell_6t
Xbit_r62_c146 bl[146] br[146] wl[62] vdd gnd cell_6t
Xbit_r63_c146 bl[146] br[146] wl[63] vdd gnd cell_6t
Xbit_r64_c146 bl[146] br[146] wl[64] vdd gnd cell_6t
Xbit_r65_c146 bl[146] br[146] wl[65] vdd gnd cell_6t
Xbit_r66_c146 bl[146] br[146] wl[66] vdd gnd cell_6t
Xbit_r67_c146 bl[146] br[146] wl[67] vdd gnd cell_6t
Xbit_r68_c146 bl[146] br[146] wl[68] vdd gnd cell_6t
Xbit_r69_c146 bl[146] br[146] wl[69] vdd gnd cell_6t
Xbit_r70_c146 bl[146] br[146] wl[70] vdd gnd cell_6t
Xbit_r71_c146 bl[146] br[146] wl[71] vdd gnd cell_6t
Xbit_r72_c146 bl[146] br[146] wl[72] vdd gnd cell_6t
Xbit_r73_c146 bl[146] br[146] wl[73] vdd gnd cell_6t
Xbit_r74_c146 bl[146] br[146] wl[74] vdd gnd cell_6t
Xbit_r75_c146 bl[146] br[146] wl[75] vdd gnd cell_6t
Xbit_r76_c146 bl[146] br[146] wl[76] vdd gnd cell_6t
Xbit_r77_c146 bl[146] br[146] wl[77] vdd gnd cell_6t
Xbit_r78_c146 bl[146] br[146] wl[78] vdd gnd cell_6t
Xbit_r79_c146 bl[146] br[146] wl[79] vdd gnd cell_6t
Xbit_r80_c146 bl[146] br[146] wl[80] vdd gnd cell_6t
Xbit_r81_c146 bl[146] br[146] wl[81] vdd gnd cell_6t
Xbit_r82_c146 bl[146] br[146] wl[82] vdd gnd cell_6t
Xbit_r83_c146 bl[146] br[146] wl[83] vdd gnd cell_6t
Xbit_r84_c146 bl[146] br[146] wl[84] vdd gnd cell_6t
Xbit_r85_c146 bl[146] br[146] wl[85] vdd gnd cell_6t
Xbit_r86_c146 bl[146] br[146] wl[86] vdd gnd cell_6t
Xbit_r87_c146 bl[146] br[146] wl[87] vdd gnd cell_6t
Xbit_r88_c146 bl[146] br[146] wl[88] vdd gnd cell_6t
Xbit_r89_c146 bl[146] br[146] wl[89] vdd gnd cell_6t
Xbit_r90_c146 bl[146] br[146] wl[90] vdd gnd cell_6t
Xbit_r91_c146 bl[146] br[146] wl[91] vdd gnd cell_6t
Xbit_r92_c146 bl[146] br[146] wl[92] vdd gnd cell_6t
Xbit_r93_c146 bl[146] br[146] wl[93] vdd gnd cell_6t
Xbit_r94_c146 bl[146] br[146] wl[94] vdd gnd cell_6t
Xbit_r95_c146 bl[146] br[146] wl[95] vdd gnd cell_6t
Xbit_r96_c146 bl[146] br[146] wl[96] vdd gnd cell_6t
Xbit_r97_c146 bl[146] br[146] wl[97] vdd gnd cell_6t
Xbit_r98_c146 bl[146] br[146] wl[98] vdd gnd cell_6t
Xbit_r99_c146 bl[146] br[146] wl[99] vdd gnd cell_6t
Xbit_r100_c146 bl[146] br[146] wl[100] vdd gnd cell_6t
Xbit_r101_c146 bl[146] br[146] wl[101] vdd gnd cell_6t
Xbit_r102_c146 bl[146] br[146] wl[102] vdd gnd cell_6t
Xbit_r103_c146 bl[146] br[146] wl[103] vdd gnd cell_6t
Xbit_r104_c146 bl[146] br[146] wl[104] vdd gnd cell_6t
Xbit_r105_c146 bl[146] br[146] wl[105] vdd gnd cell_6t
Xbit_r106_c146 bl[146] br[146] wl[106] vdd gnd cell_6t
Xbit_r107_c146 bl[146] br[146] wl[107] vdd gnd cell_6t
Xbit_r108_c146 bl[146] br[146] wl[108] vdd gnd cell_6t
Xbit_r109_c146 bl[146] br[146] wl[109] vdd gnd cell_6t
Xbit_r110_c146 bl[146] br[146] wl[110] vdd gnd cell_6t
Xbit_r111_c146 bl[146] br[146] wl[111] vdd gnd cell_6t
Xbit_r112_c146 bl[146] br[146] wl[112] vdd gnd cell_6t
Xbit_r113_c146 bl[146] br[146] wl[113] vdd gnd cell_6t
Xbit_r114_c146 bl[146] br[146] wl[114] vdd gnd cell_6t
Xbit_r115_c146 bl[146] br[146] wl[115] vdd gnd cell_6t
Xbit_r116_c146 bl[146] br[146] wl[116] vdd gnd cell_6t
Xbit_r117_c146 bl[146] br[146] wl[117] vdd gnd cell_6t
Xbit_r118_c146 bl[146] br[146] wl[118] vdd gnd cell_6t
Xbit_r119_c146 bl[146] br[146] wl[119] vdd gnd cell_6t
Xbit_r120_c146 bl[146] br[146] wl[120] vdd gnd cell_6t
Xbit_r121_c146 bl[146] br[146] wl[121] vdd gnd cell_6t
Xbit_r122_c146 bl[146] br[146] wl[122] vdd gnd cell_6t
Xbit_r123_c146 bl[146] br[146] wl[123] vdd gnd cell_6t
Xbit_r124_c146 bl[146] br[146] wl[124] vdd gnd cell_6t
Xbit_r125_c146 bl[146] br[146] wl[125] vdd gnd cell_6t
Xbit_r126_c146 bl[146] br[146] wl[126] vdd gnd cell_6t
Xbit_r127_c146 bl[146] br[146] wl[127] vdd gnd cell_6t
Xbit_r128_c146 bl[146] br[146] wl[128] vdd gnd cell_6t
Xbit_r129_c146 bl[146] br[146] wl[129] vdd gnd cell_6t
Xbit_r130_c146 bl[146] br[146] wl[130] vdd gnd cell_6t
Xbit_r131_c146 bl[146] br[146] wl[131] vdd gnd cell_6t
Xbit_r132_c146 bl[146] br[146] wl[132] vdd gnd cell_6t
Xbit_r133_c146 bl[146] br[146] wl[133] vdd gnd cell_6t
Xbit_r134_c146 bl[146] br[146] wl[134] vdd gnd cell_6t
Xbit_r135_c146 bl[146] br[146] wl[135] vdd gnd cell_6t
Xbit_r136_c146 bl[146] br[146] wl[136] vdd gnd cell_6t
Xbit_r137_c146 bl[146] br[146] wl[137] vdd gnd cell_6t
Xbit_r138_c146 bl[146] br[146] wl[138] vdd gnd cell_6t
Xbit_r139_c146 bl[146] br[146] wl[139] vdd gnd cell_6t
Xbit_r140_c146 bl[146] br[146] wl[140] vdd gnd cell_6t
Xbit_r141_c146 bl[146] br[146] wl[141] vdd gnd cell_6t
Xbit_r142_c146 bl[146] br[146] wl[142] vdd gnd cell_6t
Xbit_r143_c146 bl[146] br[146] wl[143] vdd gnd cell_6t
Xbit_r144_c146 bl[146] br[146] wl[144] vdd gnd cell_6t
Xbit_r145_c146 bl[146] br[146] wl[145] vdd gnd cell_6t
Xbit_r146_c146 bl[146] br[146] wl[146] vdd gnd cell_6t
Xbit_r147_c146 bl[146] br[146] wl[147] vdd gnd cell_6t
Xbit_r148_c146 bl[146] br[146] wl[148] vdd gnd cell_6t
Xbit_r149_c146 bl[146] br[146] wl[149] vdd gnd cell_6t
Xbit_r150_c146 bl[146] br[146] wl[150] vdd gnd cell_6t
Xbit_r151_c146 bl[146] br[146] wl[151] vdd gnd cell_6t
Xbit_r152_c146 bl[146] br[146] wl[152] vdd gnd cell_6t
Xbit_r153_c146 bl[146] br[146] wl[153] vdd gnd cell_6t
Xbit_r154_c146 bl[146] br[146] wl[154] vdd gnd cell_6t
Xbit_r155_c146 bl[146] br[146] wl[155] vdd gnd cell_6t
Xbit_r156_c146 bl[146] br[146] wl[156] vdd gnd cell_6t
Xbit_r157_c146 bl[146] br[146] wl[157] vdd gnd cell_6t
Xbit_r158_c146 bl[146] br[146] wl[158] vdd gnd cell_6t
Xbit_r159_c146 bl[146] br[146] wl[159] vdd gnd cell_6t
Xbit_r160_c146 bl[146] br[146] wl[160] vdd gnd cell_6t
Xbit_r161_c146 bl[146] br[146] wl[161] vdd gnd cell_6t
Xbit_r162_c146 bl[146] br[146] wl[162] vdd gnd cell_6t
Xbit_r163_c146 bl[146] br[146] wl[163] vdd gnd cell_6t
Xbit_r164_c146 bl[146] br[146] wl[164] vdd gnd cell_6t
Xbit_r165_c146 bl[146] br[146] wl[165] vdd gnd cell_6t
Xbit_r166_c146 bl[146] br[146] wl[166] vdd gnd cell_6t
Xbit_r167_c146 bl[146] br[146] wl[167] vdd gnd cell_6t
Xbit_r168_c146 bl[146] br[146] wl[168] vdd gnd cell_6t
Xbit_r169_c146 bl[146] br[146] wl[169] vdd gnd cell_6t
Xbit_r170_c146 bl[146] br[146] wl[170] vdd gnd cell_6t
Xbit_r171_c146 bl[146] br[146] wl[171] vdd gnd cell_6t
Xbit_r172_c146 bl[146] br[146] wl[172] vdd gnd cell_6t
Xbit_r173_c146 bl[146] br[146] wl[173] vdd gnd cell_6t
Xbit_r174_c146 bl[146] br[146] wl[174] vdd gnd cell_6t
Xbit_r175_c146 bl[146] br[146] wl[175] vdd gnd cell_6t
Xbit_r176_c146 bl[146] br[146] wl[176] vdd gnd cell_6t
Xbit_r177_c146 bl[146] br[146] wl[177] vdd gnd cell_6t
Xbit_r178_c146 bl[146] br[146] wl[178] vdd gnd cell_6t
Xbit_r179_c146 bl[146] br[146] wl[179] vdd gnd cell_6t
Xbit_r180_c146 bl[146] br[146] wl[180] vdd gnd cell_6t
Xbit_r181_c146 bl[146] br[146] wl[181] vdd gnd cell_6t
Xbit_r182_c146 bl[146] br[146] wl[182] vdd gnd cell_6t
Xbit_r183_c146 bl[146] br[146] wl[183] vdd gnd cell_6t
Xbit_r184_c146 bl[146] br[146] wl[184] vdd gnd cell_6t
Xbit_r185_c146 bl[146] br[146] wl[185] vdd gnd cell_6t
Xbit_r186_c146 bl[146] br[146] wl[186] vdd gnd cell_6t
Xbit_r187_c146 bl[146] br[146] wl[187] vdd gnd cell_6t
Xbit_r188_c146 bl[146] br[146] wl[188] vdd gnd cell_6t
Xbit_r189_c146 bl[146] br[146] wl[189] vdd gnd cell_6t
Xbit_r190_c146 bl[146] br[146] wl[190] vdd gnd cell_6t
Xbit_r191_c146 bl[146] br[146] wl[191] vdd gnd cell_6t
Xbit_r192_c146 bl[146] br[146] wl[192] vdd gnd cell_6t
Xbit_r193_c146 bl[146] br[146] wl[193] vdd gnd cell_6t
Xbit_r194_c146 bl[146] br[146] wl[194] vdd gnd cell_6t
Xbit_r195_c146 bl[146] br[146] wl[195] vdd gnd cell_6t
Xbit_r196_c146 bl[146] br[146] wl[196] vdd gnd cell_6t
Xbit_r197_c146 bl[146] br[146] wl[197] vdd gnd cell_6t
Xbit_r198_c146 bl[146] br[146] wl[198] vdd gnd cell_6t
Xbit_r199_c146 bl[146] br[146] wl[199] vdd gnd cell_6t
Xbit_r200_c146 bl[146] br[146] wl[200] vdd gnd cell_6t
Xbit_r201_c146 bl[146] br[146] wl[201] vdd gnd cell_6t
Xbit_r202_c146 bl[146] br[146] wl[202] vdd gnd cell_6t
Xbit_r203_c146 bl[146] br[146] wl[203] vdd gnd cell_6t
Xbit_r204_c146 bl[146] br[146] wl[204] vdd gnd cell_6t
Xbit_r205_c146 bl[146] br[146] wl[205] vdd gnd cell_6t
Xbit_r206_c146 bl[146] br[146] wl[206] vdd gnd cell_6t
Xbit_r207_c146 bl[146] br[146] wl[207] vdd gnd cell_6t
Xbit_r208_c146 bl[146] br[146] wl[208] vdd gnd cell_6t
Xbit_r209_c146 bl[146] br[146] wl[209] vdd gnd cell_6t
Xbit_r210_c146 bl[146] br[146] wl[210] vdd gnd cell_6t
Xbit_r211_c146 bl[146] br[146] wl[211] vdd gnd cell_6t
Xbit_r212_c146 bl[146] br[146] wl[212] vdd gnd cell_6t
Xbit_r213_c146 bl[146] br[146] wl[213] vdd gnd cell_6t
Xbit_r214_c146 bl[146] br[146] wl[214] vdd gnd cell_6t
Xbit_r215_c146 bl[146] br[146] wl[215] vdd gnd cell_6t
Xbit_r216_c146 bl[146] br[146] wl[216] vdd gnd cell_6t
Xbit_r217_c146 bl[146] br[146] wl[217] vdd gnd cell_6t
Xbit_r218_c146 bl[146] br[146] wl[218] vdd gnd cell_6t
Xbit_r219_c146 bl[146] br[146] wl[219] vdd gnd cell_6t
Xbit_r220_c146 bl[146] br[146] wl[220] vdd gnd cell_6t
Xbit_r221_c146 bl[146] br[146] wl[221] vdd gnd cell_6t
Xbit_r222_c146 bl[146] br[146] wl[222] vdd gnd cell_6t
Xbit_r223_c146 bl[146] br[146] wl[223] vdd gnd cell_6t
Xbit_r224_c146 bl[146] br[146] wl[224] vdd gnd cell_6t
Xbit_r225_c146 bl[146] br[146] wl[225] vdd gnd cell_6t
Xbit_r226_c146 bl[146] br[146] wl[226] vdd gnd cell_6t
Xbit_r227_c146 bl[146] br[146] wl[227] vdd gnd cell_6t
Xbit_r228_c146 bl[146] br[146] wl[228] vdd gnd cell_6t
Xbit_r229_c146 bl[146] br[146] wl[229] vdd gnd cell_6t
Xbit_r230_c146 bl[146] br[146] wl[230] vdd gnd cell_6t
Xbit_r231_c146 bl[146] br[146] wl[231] vdd gnd cell_6t
Xbit_r232_c146 bl[146] br[146] wl[232] vdd gnd cell_6t
Xbit_r233_c146 bl[146] br[146] wl[233] vdd gnd cell_6t
Xbit_r234_c146 bl[146] br[146] wl[234] vdd gnd cell_6t
Xbit_r235_c146 bl[146] br[146] wl[235] vdd gnd cell_6t
Xbit_r236_c146 bl[146] br[146] wl[236] vdd gnd cell_6t
Xbit_r237_c146 bl[146] br[146] wl[237] vdd gnd cell_6t
Xbit_r238_c146 bl[146] br[146] wl[238] vdd gnd cell_6t
Xbit_r239_c146 bl[146] br[146] wl[239] vdd gnd cell_6t
Xbit_r240_c146 bl[146] br[146] wl[240] vdd gnd cell_6t
Xbit_r241_c146 bl[146] br[146] wl[241] vdd gnd cell_6t
Xbit_r242_c146 bl[146] br[146] wl[242] vdd gnd cell_6t
Xbit_r243_c146 bl[146] br[146] wl[243] vdd gnd cell_6t
Xbit_r244_c146 bl[146] br[146] wl[244] vdd gnd cell_6t
Xbit_r245_c146 bl[146] br[146] wl[245] vdd gnd cell_6t
Xbit_r246_c146 bl[146] br[146] wl[246] vdd gnd cell_6t
Xbit_r247_c146 bl[146] br[146] wl[247] vdd gnd cell_6t
Xbit_r248_c146 bl[146] br[146] wl[248] vdd gnd cell_6t
Xbit_r249_c146 bl[146] br[146] wl[249] vdd gnd cell_6t
Xbit_r250_c146 bl[146] br[146] wl[250] vdd gnd cell_6t
Xbit_r251_c146 bl[146] br[146] wl[251] vdd gnd cell_6t
Xbit_r252_c146 bl[146] br[146] wl[252] vdd gnd cell_6t
Xbit_r253_c146 bl[146] br[146] wl[253] vdd gnd cell_6t
Xbit_r254_c146 bl[146] br[146] wl[254] vdd gnd cell_6t
Xbit_r255_c146 bl[146] br[146] wl[255] vdd gnd cell_6t
Xbit_r0_c147 bl[147] br[147] wl[0] vdd gnd cell_6t
Xbit_r1_c147 bl[147] br[147] wl[1] vdd gnd cell_6t
Xbit_r2_c147 bl[147] br[147] wl[2] vdd gnd cell_6t
Xbit_r3_c147 bl[147] br[147] wl[3] vdd gnd cell_6t
Xbit_r4_c147 bl[147] br[147] wl[4] vdd gnd cell_6t
Xbit_r5_c147 bl[147] br[147] wl[5] vdd gnd cell_6t
Xbit_r6_c147 bl[147] br[147] wl[6] vdd gnd cell_6t
Xbit_r7_c147 bl[147] br[147] wl[7] vdd gnd cell_6t
Xbit_r8_c147 bl[147] br[147] wl[8] vdd gnd cell_6t
Xbit_r9_c147 bl[147] br[147] wl[9] vdd gnd cell_6t
Xbit_r10_c147 bl[147] br[147] wl[10] vdd gnd cell_6t
Xbit_r11_c147 bl[147] br[147] wl[11] vdd gnd cell_6t
Xbit_r12_c147 bl[147] br[147] wl[12] vdd gnd cell_6t
Xbit_r13_c147 bl[147] br[147] wl[13] vdd gnd cell_6t
Xbit_r14_c147 bl[147] br[147] wl[14] vdd gnd cell_6t
Xbit_r15_c147 bl[147] br[147] wl[15] vdd gnd cell_6t
Xbit_r16_c147 bl[147] br[147] wl[16] vdd gnd cell_6t
Xbit_r17_c147 bl[147] br[147] wl[17] vdd gnd cell_6t
Xbit_r18_c147 bl[147] br[147] wl[18] vdd gnd cell_6t
Xbit_r19_c147 bl[147] br[147] wl[19] vdd gnd cell_6t
Xbit_r20_c147 bl[147] br[147] wl[20] vdd gnd cell_6t
Xbit_r21_c147 bl[147] br[147] wl[21] vdd gnd cell_6t
Xbit_r22_c147 bl[147] br[147] wl[22] vdd gnd cell_6t
Xbit_r23_c147 bl[147] br[147] wl[23] vdd gnd cell_6t
Xbit_r24_c147 bl[147] br[147] wl[24] vdd gnd cell_6t
Xbit_r25_c147 bl[147] br[147] wl[25] vdd gnd cell_6t
Xbit_r26_c147 bl[147] br[147] wl[26] vdd gnd cell_6t
Xbit_r27_c147 bl[147] br[147] wl[27] vdd gnd cell_6t
Xbit_r28_c147 bl[147] br[147] wl[28] vdd gnd cell_6t
Xbit_r29_c147 bl[147] br[147] wl[29] vdd gnd cell_6t
Xbit_r30_c147 bl[147] br[147] wl[30] vdd gnd cell_6t
Xbit_r31_c147 bl[147] br[147] wl[31] vdd gnd cell_6t
Xbit_r32_c147 bl[147] br[147] wl[32] vdd gnd cell_6t
Xbit_r33_c147 bl[147] br[147] wl[33] vdd gnd cell_6t
Xbit_r34_c147 bl[147] br[147] wl[34] vdd gnd cell_6t
Xbit_r35_c147 bl[147] br[147] wl[35] vdd gnd cell_6t
Xbit_r36_c147 bl[147] br[147] wl[36] vdd gnd cell_6t
Xbit_r37_c147 bl[147] br[147] wl[37] vdd gnd cell_6t
Xbit_r38_c147 bl[147] br[147] wl[38] vdd gnd cell_6t
Xbit_r39_c147 bl[147] br[147] wl[39] vdd gnd cell_6t
Xbit_r40_c147 bl[147] br[147] wl[40] vdd gnd cell_6t
Xbit_r41_c147 bl[147] br[147] wl[41] vdd gnd cell_6t
Xbit_r42_c147 bl[147] br[147] wl[42] vdd gnd cell_6t
Xbit_r43_c147 bl[147] br[147] wl[43] vdd gnd cell_6t
Xbit_r44_c147 bl[147] br[147] wl[44] vdd gnd cell_6t
Xbit_r45_c147 bl[147] br[147] wl[45] vdd gnd cell_6t
Xbit_r46_c147 bl[147] br[147] wl[46] vdd gnd cell_6t
Xbit_r47_c147 bl[147] br[147] wl[47] vdd gnd cell_6t
Xbit_r48_c147 bl[147] br[147] wl[48] vdd gnd cell_6t
Xbit_r49_c147 bl[147] br[147] wl[49] vdd gnd cell_6t
Xbit_r50_c147 bl[147] br[147] wl[50] vdd gnd cell_6t
Xbit_r51_c147 bl[147] br[147] wl[51] vdd gnd cell_6t
Xbit_r52_c147 bl[147] br[147] wl[52] vdd gnd cell_6t
Xbit_r53_c147 bl[147] br[147] wl[53] vdd gnd cell_6t
Xbit_r54_c147 bl[147] br[147] wl[54] vdd gnd cell_6t
Xbit_r55_c147 bl[147] br[147] wl[55] vdd gnd cell_6t
Xbit_r56_c147 bl[147] br[147] wl[56] vdd gnd cell_6t
Xbit_r57_c147 bl[147] br[147] wl[57] vdd gnd cell_6t
Xbit_r58_c147 bl[147] br[147] wl[58] vdd gnd cell_6t
Xbit_r59_c147 bl[147] br[147] wl[59] vdd gnd cell_6t
Xbit_r60_c147 bl[147] br[147] wl[60] vdd gnd cell_6t
Xbit_r61_c147 bl[147] br[147] wl[61] vdd gnd cell_6t
Xbit_r62_c147 bl[147] br[147] wl[62] vdd gnd cell_6t
Xbit_r63_c147 bl[147] br[147] wl[63] vdd gnd cell_6t
Xbit_r64_c147 bl[147] br[147] wl[64] vdd gnd cell_6t
Xbit_r65_c147 bl[147] br[147] wl[65] vdd gnd cell_6t
Xbit_r66_c147 bl[147] br[147] wl[66] vdd gnd cell_6t
Xbit_r67_c147 bl[147] br[147] wl[67] vdd gnd cell_6t
Xbit_r68_c147 bl[147] br[147] wl[68] vdd gnd cell_6t
Xbit_r69_c147 bl[147] br[147] wl[69] vdd gnd cell_6t
Xbit_r70_c147 bl[147] br[147] wl[70] vdd gnd cell_6t
Xbit_r71_c147 bl[147] br[147] wl[71] vdd gnd cell_6t
Xbit_r72_c147 bl[147] br[147] wl[72] vdd gnd cell_6t
Xbit_r73_c147 bl[147] br[147] wl[73] vdd gnd cell_6t
Xbit_r74_c147 bl[147] br[147] wl[74] vdd gnd cell_6t
Xbit_r75_c147 bl[147] br[147] wl[75] vdd gnd cell_6t
Xbit_r76_c147 bl[147] br[147] wl[76] vdd gnd cell_6t
Xbit_r77_c147 bl[147] br[147] wl[77] vdd gnd cell_6t
Xbit_r78_c147 bl[147] br[147] wl[78] vdd gnd cell_6t
Xbit_r79_c147 bl[147] br[147] wl[79] vdd gnd cell_6t
Xbit_r80_c147 bl[147] br[147] wl[80] vdd gnd cell_6t
Xbit_r81_c147 bl[147] br[147] wl[81] vdd gnd cell_6t
Xbit_r82_c147 bl[147] br[147] wl[82] vdd gnd cell_6t
Xbit_r83_c147 bl[147] br[147] wl[83] vdd gnd cell_6t
Xbit_r84_c147 bl[147] br[147] wl[84] vdd gnd cell_6t
Xbit_r85_c147 bl[147] br[147] wl[85] vdd gnd cell_6t
Xbit_r86_c147 bl[147] br[147] wl[86] vdd gnd cell_6t
Xbit_r87_c147 bl[147] br[147] wl[87] vdd gnd cell_6t
Xbit_r88_c147 bl[147] br[147] wl[88] vdd gnd cell_6t
Xbit_r89_c147 bl[147] br[147] wl[89] vdd gnd cell_6t
Xbit_r90_c147 bl[147] br[147] wl[90] vdd gnd cell_6t
Xbit_r91_c147 bl[147] br[147] wl[91] vdd gnd cell_6t
Xbit_r92_c147 bl[147] br[147] wl[92] vdd gnd cell_6t
Xbit_r93_c147 bl[147] br[147] wl[93] vdd gnd cell_6t
Xbit_r94_c147 bl[147] br[147] wl[94] vdd gnd cell_6t
Xbit_r95_c147 bl[147] br[147] wl[95] vdd gnd cell_6t
Xbit_r96_c147 bl[147] br[147] wl[96] vdd gnd cell_6t
Xbit_r97_c147 bl[147] br[147] wl[97] vdd gnd cell_6t
Xbit_r98_c147 bl[147] br[147] wl[98] vdd gnd cell_6t
Xbit_r99_c147 bl[147] br[147] wl[99] vdd gnd cell_6t
Xbit_r100_c147 bl[147] br[147] wl[100] vdd gnd cell_6t
Xbit_r101_c147 bl[147] br[147] wl[101] vdd gnd cell_6t
Xbit_r102_c147 bl[147] br[147] wl[102] vdd gnd cell_6t
Xbit_r103_c147 bl[147] br[147] wl[103] vdd gnd cell_6t
Xbit_r104_c147 bl[147] br[147] wl[104] vdd gnd cell_6t
Xbit_r105_c147 bl[147] br[147] wl[105] vdd gnd cell_6t
Xbit_r106_c147 bl[147] br[147] wl[106] vdd gnd cell_6t
Xbit_r107_c147 bl[147] br[147] wl[107] vdd gnd cell_6t
Xbit_r108_c147 bl[147] br[147] wl[108] vdd gnd cell_6t
Xbit_r109_c147 bl[147] br[147] wl[109] vdd gnd cell_6t
Xbit_r110_c147 bl[147] br[147] wl[110] vdd gnd cell_6t
Xbit_r111_c147 bl[147] br[147] wl[111] vdd gnd cell_6t
Xbit_r112_c147 bl[147] br[147] wl[112] vdd gnd cell_6t
Xbit_r113_c147 bl[147] br[147] wl[113] vdd gnd cell_6t
Xbit_r114_c147 bl[147] br[147] wl[114] vdd gnd cell_6t
Xbit_r115_c147 bl[147] br[147] wl[115] vdd gnd cell_6t
Xbit_r116_c147 bl[147] br[147] wl[116] vdd gnd cell_6t
Xbit_r117_c147 bl[147] br[147] wl[117] vdd gnd cell_6t
Xbit_r118_c147 bl[147] br[147] wl[118] vdd gnd cell_6t
Xbit_r119_c147 bl[147] br[147] wl[119] vdd gnd cell_6t
Xbit_r120_c147 bl[147] br[147] wl[120] vdd gnd cell_6t
Xbit_r121_c147 bl[147] br[147] wl[121] vdd gnd cell_6t
Xbit_r122_c147 bl[147] br[147] wl[122] vdd gnd cell_6t
Xbit_r123_c147 bl[147] br[147] wl[123] vdd gnd cell_6t
Xbit_r124_c147 bl[147] br[147] wl[124] vdd gnd cell_6t
Xbit_r125_c147 bl[147] br[147] wl[125] vdd gnd cell_6t
Xbit_r126_c147 bl[147] br[147] wl[126] vdd gnd cell_6t
Xbit_r127_c147 bl[147] br[147] wl[127] vdd gnd cell_6t
Xbit_r128_c147 bl[147] br[147] wl[128] vdd gnd cell_6t
Xbit_r129_c147 bl[147] br[147] wl[129] vdd gnd cell_6t
Xbit_r130_c147 bl[147] br[147] wl[130] vdd gnd cell_6t
Xbit_r131_c147 bl[147] br[147] wl[131] vdd gnd cell_6t
Xbit_r132_c147 bl[147] br[147] wl[132] vdd gnd cell_6t
Xbit_r133_c147 bl[147] br[147] wl[133] vdd gnd cell_6t
Xbit_r134_c147 bl[147] br[147] wl[134] vdd gnd cell_6t
Xbit_r135_c147 bl[147] br[147] wl[135] vdd gnd cell_6t
Xbit_r136_c147 bl[147] br[147] wl[136] vdd gnd cell_6t
Xbit_r137_c147 bl[147] br[147] wl[137] vdd gnd cell_6t
Xbit_r138_c147 bl[147] br[147] wl[138] vdd gnd cell_6t
Xbit_r139_c147 bl[147] br[147] wl[139] vdd gnd cell_6t
Xbit_r140_c147 bl[147] br[147] wl[140] vdd gnd cell_6t
Xbit_r141_c147 bl[147] br[147] wl[141] vdd gnd cell_6t
Xbit_r142_c147 bl[147] br[147] wl[142] vdd gnd cell_6t
Xbit_r143_c147 bl[147] br[147] wl[143] vdd gnd cell_6t
Xbit_r144_c147 bl[147] br[147] wl[144] vdd gnd cell_6t
Xbit_r145_c147 bl[147] br[147] wl[145] vdd gnd cell_6t
Xbit_r146_c147 bl[147] br[147] wl[146] vdd gnd cell_6t
Xbit_r147_c147 bl[147] br[147] wl[147] vdd gnd cell_6t
Xbit_r148_c147 bl[147] br[147] wl[148] vdd gnd cell_6t
Xbit_r149_c147 bl[147] br[147] wl[149] vdd gnd cell_6t
Xbit_r150_c147 bl[147] br[147] wl[150] vdd gnd cell_6t
Xbit_r151_c147 bl[147] br[147] wl[151] vdd gnd cell_6t
Xbit_r152_c147 bl[147] br[147] wl[152] vdd gnd cell_6t
Xbit_r153_c147 bl[147] br[147] wl[153] vdd gnd cell_6t
Xbit_r154_c147 bl[147] br[147] wl[154] vdd gnd cell_6t
Xbit_r155_c147 bl[147] br[147] wl[155] vdd gnd cell_6t
Xbit_r156_c147 bl[147] br[147] wl[156] vdd gnd cell_6t
Xbit_r157_c147 bl[147] br[147] wl[157] vdd gnd cell_6t
Xbit_r158_c147 bl[147] br[147] wl[158] vdd gnd cell_6t
Xbit_r159_c147 bl[147] br[147] wl[159] vdd gnd cell_6t
Xbit_r160_c147 bl[147] br[147] wl[160] vdd gnd cell_6t
Xbit_r161_c147 bl[147] br[147] wl[161] vdd gnd cell_6t
Xbit_r162_c147 bl[147] br[147] wl[162] vdd gnd cell_6t
Xbit_r163_c147 bl[147] br[147] wl[163] vdd gnd cell_6t
Xbit_r164_c147 bl[147] br[147] wl[164] vdd gnd cell_6t
Xbit_r165_c147 bl[147] br[147] wl[165] vdd gnd cell_6t
Xbit_r166_c147 bl[147] br[147] wl[166] vdd gnd cell_6t
Xbit_r167_c147 bl[147] br[147] wl[167] vdd gnd cell_6t
Xbit_r168_c147 bl[147] br[147] wl[168] vdd gnd cell_6t
Xbit_r169_c147 bl[147] br[147] wl[169] vdd gnd cell_6t
Xbit_r170_c147 bl[147] br[147] wl[170] vdd gnd cell_6t
Xbit_r171_c147 bl[147] br[147] wl[171] vdd gnd cell_6t
Xbit_r172_c147 bl[147] br[147] wl[172] vdd gnd cell_6t
Xbit_r173_c147 bl[147] br[147] wl[173] vdd gnd cell_6t
Xbit_r174_c147 bl[147] br[147] wl[174] vdd gnd cell_6t
Xbit_r175_c147 bl[147] br[147] wl[175] vdd gnd cell_6t
Xbit_r176_c147 bl[147] br[147] wl[176] vdd gnd cell_6t
Xbit_r177_c147 bl[147] br[147] wl[177] vdd gnd cell_6t
Xbit_r178_c147 bl[147] br[147] wl[178] vdd gnd cell_6t
Xbit_r179_c147 bl[147] br[147] wl[179] vdd gnd cell_6t
Xbit_r180_c147 bl[147] br[147] wl[180] vdd gnd cell_6t
Xbit_r181_c147 bl[147] br[147] wl[181] vdd gnd cell_6t
Xbit_r182_c147 bl[147] br[147] wl[182] vdd gnd cell_6t
Xbit_r183_c147 bl[147] br[147] wl[183] vdd gnd cell_6t
Xbit_r184_c147 bl[147] br[147] wl[184] vdd gnd cell_6t
Xbit_r185_c147 bl[147] br[147] wl[185] vdd gnd cell_6t
Xbit_r186_c147 bl[147] br[147] wl[186] vdd gnd cell_6t
Xbit_r187_c147 bl[147] br[147] wl[187] vdd gnd cell_6t
Xbit_r188_c147 bl[147] br[147] wl[188] vdd gnd cell_6t
Xbit_r189_c147 bl[147] br[147] wl[189] vdd gnd cell_6t
Xbit_r190_c147 bl[147] br[147] wl[190] vdd gnd cell_6t
Xbit_r191_c147 bl[147] br[147] wl[191] vdd gnd cell_6t
Xbit_r192_c147 bl[147] br[147] wl[192] vdd gnd cell_6t
Xbit_r193_c147 bl[147] br[147] wl[193] vdd gnd cell_6t
Xbit_r194_c147 bl[147] br[147] wl[194] vdd gnd cell_6t
Xbit_r195_c147 bl[147] br[147] wl[195] vdd gnd cell_6t
Xbit_r196_c147 bl[147] br[147] wl[196] vdd gnd cell_6t
Xbit_r197_c147 bl[147] br[147] wl[197] vdd gnd cell_6t
Xbit_r198_c147 bl[147] br[147] wl[198] vdd gnd cell_6t
Xbit_r199_c147 bl[147] br[147] wl[199] vdd gnd cell_6t
Xbit_r200_c147 bl[147] br[147] wl[200] vdd gnd cell_6t
Xbit_r201_c147 bl[147] br[147] wl[201] vdd gnd cell_6t
Xbit_r202_c147 bl[147] br[147] wl[202] vdd gnd cell_6t
Xbit_r203_c147 bl[147] br[147] wl[203] vdd gnd cell_6t
Xbit_r204_c147 bl[147] br[147] wl[204] vdd gnd cell_6t
Xbit_r205_c147 bl[147] br[147] wl[205] vdd gnd cell_6t
Xbit_r206_c147 bl[147] br[147] wl[206] vdd gnd cell_6t
Xbit_r207_c147 bl[147] br[147] wl[207] vdd gnd cell_6t
Xbit_r208_c147 bl[147] br[147] wl[208] vdd gnd cell_6t
Xbit_r209_c147 bl[147] br[147] wl[209] vdd gnd cell_6t
Xbit_r210_c147 bl[147] br[147] wl[210] vdd gnd cell_6t
Xbit_r211_c147 bl[147] br[147] wl[211] vdd gnd cell_6t
Xbit_r212_c147 bl[147] br[147] wl[212] vdd gnd cell_6t
Xbit_r213_c147 bl[147] br[147] wl[213] vdd gnd cell_6t
Xbit_r214_c147 bl[147] br[147] wl[214] vdd gnd cell_6t
Xbit_r215_c147 bl[147] br[147] wl[215] vdd gnd cell_6t
Xbit_r216_c147 bl[147] br[147] wl[216] vdd gnd cell_6t
Xbit_r217_c147 bl[147] br[147] wl[217] vdd gnd cell_6t
Xbit_r218_c147 bl[147] br[147] wl[218] vdd gnd cell_6t
Xbit_r219_c147 bl[147] br[147] wl[219] vdd gnd cell_6t
Xbit_r220_c147 bl[147] br[147] wl[220] vdd gnd cell_6t
Xbit_r221_c147 bl[147] br[147] wl[221] vdd gnd cell_6t
Xbit_r222_c147 bl[147] br[147] wl[222] vdd gnd cell_6t
Xbit_r223_c147 bl[147] br[147] wl[223] vdd gnd cell_6t
Xbit_r224_c147 bl[147] br[147] wl[224] vdd gnd cell_6t
Xbit_r225_c147 bl[147] br[147] wl[225] vdd gnd cell_6t
Xbit_r226_c147 bl[147] br[147] wl[226] vdd gnd cell_6t
Xbit_r227_c147 bl[147] br[147] wl[227] vdd gnd cell_6t
Xbit_r228_c147 bl[147] br[147] wl[228] vdd gnd cell_6t
Xbit_r229_c147 bl[147] br[147] wl[229] vdd gnd cell_6t
Xbit_r230_c147 bl[147] br[147] wl[230] vdd gnd cell_6t
Xbit_r231_c147 bl[147] br[147] wl[231] vdd gnd cell_6t
Xbit_r232_c147 bl[147] br[147] wl[232] vdd gnd cell_6t
Xbit_r233_c147 bl[147] br[147] wl[233] vdd gnd cell_6t
Xbit_r234_c147 bl[147] br[147] wl[234] vdd gnd cell_6t
Xbit_r235_c147 bl[147] br[147] wl[235] vdd gnd cell_6t
Xbit_r236_c147 bl[147] br[147] wl[236] vdd gnd cell_6t
Xbit_r237_c147 bl[147] br[147] wl[237] vdd gnd cell_6t
Xbit_r238_c147 bl[147] br[147] wl[238] vdd gnd cell_6t
Xbit_r239_c147 bl[147] br[147] wl[239] vdd gnd cell_6t
Xbit_r240_c147 bl[147] br[147] wl[240] vdd gnd cell_6t
Xbit_r241_c147 bl[147] br[147] wl[241] vdd gnd cell_6t
Xbit_r242_c147 bl[147] br[147] wl[242] vdd gnd cell_6t
Xbit_r243_c147 bl[147] br[147] wl[243] vdd gnd cell_6t
Xbit_r244_c147 bl[147] br[147] wl[244] vdd gnd cell_6t
Xbit_r245_c147 bl[147] br[147] wl[245] vdd gnd cell_6t
Xbit_r246_c147 bl[147] br[147] wl[246] vdd gnd cell_6t
Xbit_r247_c147 bl[147] br[147] wl[247] vdd gnd cell_6t
Xbit_r248_c147 bl[147] br[147] wl[248] vdd gnd cell_6t
Xbit_r249_c147 bl[147] br[147] wl[249] vdd gnd cell_6t
Xbit_r250_c147 bl[147] br[147] wl[250] vdd gnd cell_6t
Xbit_r251_c147 bl[147] br[147] wl[251] vdd gnd cell_6t
Xbit_r252_c147 bl[147] br[147] wl[252] vdd gnd cell_6t
Xbit_r253_c147 bl[147] br[147] wl[253] vdd gnd cell_6t
Xbit_r254_c147 bl[147] br[147] wl[254] vdd gnd cell_6t
Xbit_r255_c147 bl[147] br[147] wl[255] vdd gnd cell_6t
Xbit_r0_c148 bl[148] br[148] wl[0] vdd gnd cell_6t
Xbit_r1_c148 bl[148] br[148] wl[1] vdd gnd cell_6t
Xbit_r2_c148 bl[148] br[148] wl[2] vdd gnd cell_6t
Xbit_r3_c148 bl[148] br[148] wl[3] vdd gnd cell_6t
Xbit_r4_c148 bl[148] br[148] wl[4] vdd gnd cell_6t
Xbit_r5_c148 bl[148] br[148] wl[5] vdd gnd cell_6t
Xbit_r6_c148 bl[148] br[148] wl[6] vdd gnd cell_6t
Xbit_r7_c148 bl[148] br[148] wl[7] vdd gnd cell_6t
Xbit_r8_c148 bl[148] br[148] wl[8] vdd gnd cell_6t
Xbit_r9_c148 bl[148] br[148] wl[9] vdd gnd cell_6t
Xbit_r10_c148 bl[148] br[148] wl[10] vdd gnd cell_6t
Xbit_r11_c148 bl[148] br[148] wl[11] vdd gnd cell_6t
Xbit_r12_c148 bl[148] br[148] wl[12] vdd gnd cell_6t
Xbit_r13_c148 bl[148] br[148] wl[13] vdd gnd cell_6t
Xbit_r14_c148 bl[148] br[148] wl[14] vdd gnd cell_6t
Xbit_r15_c148 bl[148] br[148] wl[15] vdd gnd cell_6t
Xbit_r16_c148 bl[148] br[148] wl[16] vdd gnd cell_6t
Xbit_r17_c148 bl[148] br[148] wl[17] vdd gnd cell_6t
Xbit_r18_c148 bl[148] br[148] wl[18] vdd gnd cell_6t
Xbit_r19_c148 bl[148] br[148] wl[19] vdd gnd cell_6t
Xbit_r20_c148 bl[148] br[148] wl[20] vdd gnd cell_6t
Xbit_r21_c148 bl[148] br[148] wl[21] vdd gnd cell_6t
Xbit_r22_c148 bl[148] br[148] wl[22] vdd gnd cell_6t
Xbit_r23_c148 bl[148] br[148] wl[23] vdd gnd cell_6t
Xbit_r24_c148 bl[148] br[148] wl[24] vdd gnd cell_6t
Xbit_r25_c148 bl[148] br[148] wl[25] vdd gnd cell_6t
Xbit_r26_c148 bl[148] br[148] wl[26] vdd gnd cell_6t
Xbit_r27_c148 bl[148] br[148] wl[27] vdd gnd cell_6t
Xbit_r28_c148 bl[148] br[148] wl[28] vdd gnd cell_6t
Xbit_r29_c148 bl[148] br[148] wl[29] vdd gnd cell_6t
Xbit_r30_c148 bl[148] br[148] wl[30] vdd gnd cell_6t
Xbit_r31_c148 bl[148] br[148] wl[31] vdd gnd cell_6t
Xbit_r32_c148 bl[148] br[148] wl[32] vdd gnd cell_6t
Xbit_r33_c148 bl[148] br[148] wl[33] vdd gnd cell_6t
Xbit_r34_c148 bl[148] br[148] wl[34] vdd gnd cell_6t
Xbit_r35_c148 bl[148] br[148] wl[35] vdd gnd cell_6t
Xbit_r36_c148 bl[148] br[148] wl[36] vdd gnd cell_6t
Xbit_r37_c148 bl[148] br[148] wl[37] vdd gnd cell_6t
Xbit_r38_c148 bl[148] br[148] wl[38] vdd gnd cell_6t
Xbit_r39_c148 bl[148] br[148] wl[39] vdd gnd cell_6t
Xbit_r40_c148 bl[148] br[148] wl[40] vdd gnd cell_6t
Xbit_r41_c148 bl[148] br[148] wl[41] vdd gnd cell_6t
Xbit_r42_c148 bl[148] br[148] wl[42] vdd gnd cell_6t
Xbit_r43_c148 bl[148] br[148] wl[43] vdd gnd cell_6t
Xbit_r44_c148 bl[148] br[148] wl[44] vdd gnd cell_6t
Xbit_r45_c148 bl[148] br[148] wl[45] vdd gnd cell_6t
Xbit_r46_c148 bl[148] br[148] wl[46] vdd gnd cell_6t
Xbit_r47_c148 bl[148] br[148] wl[47] vdd gnd cell_6t
Xbit_r48_c148 bl[148] br[148] wl[48] vdd gnd cell_6t
Xbit_r49_c148 bl[148] br[148] wl[49] vdd gnd cell_6t
Xbit_r50_c148 bl[148] br[148] wl[50] vdd gnd cell_6t
Xbit_r51_c148 bl[148] br[148] wl[51] vdd gnd cell_6t
Xbit_r52_c148 bl[148] br[148] wl[52] vdd gnd cell_6t
Xbit_r53_c148 bl[148] br[148] wl[53] vdd gnd cell_6t
Xbit_r54_c148 bl[148] br[148] wl[54] vdd gnd cell_6t
Xbit_r55_c148 bl[148] br[148] wl[55] vdd gnd cell_6t
Xbit_r56_c148 bl[148] br[148] wl[56] vdd gnd cell_6t
Xbit_r57_c148 bl[148] br[148] wl[57] vdd gnd cell_6t
Xbit_r58_c148 bl[148] br[148] wl[58] vdd gnd cell_6t
Xbit_r59_c148 bl[148] br[148] wl[59] vdd gnd cell_6t
Xbit_r60_c148 bl[148] br[148] wl[60] vdd gnd cell_6t
Xbit_r61_c148 bl[148] br[148] wl[61] vdd gnd cell_6t
Xbit_r62_c148 bl[148] br[148] wl[62] vdd gnd cell_6t
Xbit_r63_c148 bl[148] br[148] wl[63] vdd gnd cell_6t
Xbit_r64_c148 bl[148] br[148] wl[64] vdd gnd cell_6t
Xbit_r65_c148 bl[148] br[148] wl[65] vdd gnd cell_6t
Xbit_r66_c148 bl[148] br[148] wl[66] vdd gnd cell_6t
Xbit_r67_c148 bl[148] br[148] wl[67] vdd gnd cell_6t
Xbit_r68_c148 bl[148] br[148] wl[68] vdd gnd cell_6t
Xbit_r69_c148 bl[148] br[148] wl[69] vdd gnd cell_6t
Xbit_r70_c148 bl[148] br[148] wl[70] vdd gnd cell_6t
Xbit_r71_c148 bl[148] br[148] wl[71] vdd gnd cell_6t
Xbit_r72_c148 bl[148] br[148] wl[72] vdd gnd cell_6t
Xbit_r73_c148 bl[148] br[148] wl[73] vdd gnd cell_6t
Xbit_r74_c148 bl[148] br[148] wl[74] vdd gnd cell_6t
Xbit_r75_c148 bl[148] br[148] wl[75] vdd gnd cell_6t
Xbit_r76_c148 bl[148] br[148] wl[76] vdd gnd cell_6t
Xbit_r77_c148 bl[148] br[148] wl[77] vdd gnd cell_6t
Xbit_r78_c148 bl[148] br[148] wl[78] vdd gnd cell_6t
Xbit_r79_c148 bl[148] br[148] wl[79] vdd gnd cell_6t
Xbit_r80_c148 bl[148] br[148] wl[80] vdd gnd cell_6t
Xbit_r81_c148 bl[148] br[148] wl[81] vdd gnd cell_6t
Xbit_r82_c148 bl[148] br[148] wl[82] vdd gnd cell_6t
Xbit_r83_c148 bl[148] br[148] wl[83] vdd gnd cell_6t
Xbit_r84_c148 bl[148] br[148] wl[84] vdd gnd cell_6t
Xbit_r85_c148 bl[148] br[148] wl[85] vdd gnd cell_6t
Xbit_r86_c148 bl[148] br[148] wl[86] vdd gnd cell_6t
Xbit_r87_c148 bl[148] br[148] wl[87] vdd gnd cell_6t
Xbit_r88_c148 bl[148] br[148] wl[88] vdd gnd cell_6t
Xbit_r89_c148 bl[148] br[148] wl[89] vdd gnd cell_6t
Xbit_r90_c148 bl[148] br[148] wl[90] vdd gnd cell_6t
Xbit_r91_c148 bl[148] br[148] wl[91] vdd gnd cell_6t
Xbit_r92_c148 bl[148] br[148] wl[92] vdd gnd cell_6t
Xbit_r93_c148 bl[148] br[148] wl[93] vdd gnd cell_6t
Xbit_r94_c148 bl[148] br[148] wl[94] vdd gnd cell_6t
Xbit_r95_c148 bl[148] br[148] wl[95] vdd gnd cell_6t
Xbit_r96_c148 bl[148] br[148] wl[96] vdd gnd cell_6t
Xbit_r97_c148 bl[148] br[148] wl[97] vdd gnd cell_6t
Xbit_r98_c148 bl[148] br[148] wl[98] vdd gnd cell_6t
Xbit_r99_c148 bl[148] br[148] wl[99] vdd gnd cell_6t
Xbit_r100_c148 bl[148] br[148] wl[100] vdd gnd cell_6t
Xbit_r101_c148 bl[148] br[148] wl[101] vdd gnd cell_6t
Xbit_r102_c148 bl[148] br[148] wl[102] vdd gnd cell_6t
Xbit_r103_c148 bl[148] br[148] wl[103] vdd gnd cell_6t
Xbit_r104_c148 bl[148] br[148] wl[104] vdd gnd cell_6t
Xbit_r105_c148 bl[148] br[148] wl[105] vdd gnd cell_6t
Xbit_r106_c148 bl[148] br[148] wl[106] vdd gnd cell_6t
Xbit_r107_c148 bl[148] br[148] wl[107] vdd gnd cell_6t
Xbit_r108_c148 bl[148] br[148] wl[108] vdd gnd cell_6t
Xbit_r109_c148 bl[148] br[148] wl[109] vdd gnd cell_6t
Xbit_r110_c148 bl[148] br[148] wl[110] vdd gnd cell_6t
Xbit_r111_c148 bl[148] br[148] wl[111] vdd gnd cell_6t
Xbit_r112_c148 bl[148] br[148] wl[112] vdd gnd cell_6t
Xbit_r113_c148 bl[148] br[148] wl[113] vdd gnd cell_6t
Xbit_r114_c148 bl[148] br[148] wl[114] vdd gnd cell_6t
Xbit_r115_c148 bl[148] br[148] wl[115] vdd gnd cell_6t
Xbit_r116_c148 bl[148] br[148] wl[116] vdd gnd cell_6t
Xbit_r117_c148 bl[148] br[148] wl[117] vdd gnd cell_6t
Xbit_r118_c148 bl[148] br[148] wl[118] vdd gnd cell_6t
Xbit_r119_c148 bl[148] br[148] wl[119] vdd gnd cell_6t
Xbit_r120_c148 bl[148] br[148] wl[120] vdd gnd cell_6t
Xbit_r121_c148 bl[148] br[148] wl[121] vdd gnd cell_6t
Xbit_r122_c148 bl[148] br[148] wl[122] vdd gnd cell_6t
Xbit_r123_c148 bl[148] br[148] wl[123] vdd gnd cell_6t
Xbit_r124_c148 bl[148] br[148] wl[124] vdd gnd cell_6t
Xbit_r125_c148 bl[148] br[148] wl[125] vdd gnd cell_6t
Xbit_r126_c148 bl[148] br[148] wl[126] vdd gnd cell_6t
Xbit_r127_c148 bl[148] br[148] wl[127] vdd gnd cell_6t
Xbit_r128_c148 bl[148] br[148] wl[128] vdd gnd cell_6t
Xbit_r129_c148 bl[148] br[148] wl[129] vdd gnd cell_6t
Xbit_r130_c148 bl[148] br[148] wl[130] vdd gnd cell_6t
Xbit_r131_c148 bl[148] br[148] wl[131] vdd gnd cell_6t
Xbit_r132_c148 bl[148] br[148] wl[132] vdd gnd cell_6t
Xbit_r133_c148 bl[148] br[148] wl[133] vdd gnd cell_6t
Xbit_r134_c148 bl[148] br[148] wl[134] vdd gnd cell_6t
Xbit_r135_c148 bl[148] br[148] wl[135] vdd gnd cell_6t
Xbit_r136_c148 bl[148] br[148] wl[136] vdd gnd cell_6t
Xbit_r137_c148 bl[148] br[148] wl[137] vdd gnd cell_6t
Xbit_r138_c148 bl[148] br[148] wl[138] vdd gnd cell_6t
Xbit_r139_c148 bl[148] br[148] wl[139] vdd gnd cell_6t
Xbit_r140_c148 bl[148] br[148] wl[140] vdd gnd cell_6t
Xbit_r141_c148 bl[148] br[148] wl[141] vdd gnd cell_6t
Xbit_r142_c148 bl[148] br[148] wl[142] vdd gnd cell_6t
Xbit_r143_c148 bl[148] br[148] wl[143] vdd gnd cell_6t
Xbit_r144_c148 bl[148] br[148] wl[144] vdd gnd cell_6t
Xbit_r145_c148 bl[148] br[148] wl[145] vdd gnd cell_6t
Xbit_r146_c148 bl[148] br[148] wl[146] vdd gnd cell_6t
Xbit_r147_c148 bl[148] br[148] wl[147] vdd gnd cell_6t
Xbit_r148_c148 bl[148] br[148] wl[148] vdd gnd cell_6t
Xbit_r149_c148 bl[148] br[148] wl[149] vdd gnd cell_6t
Xbit_r150_c148 bl[148] br[148] wl[150] vdd gnd cell_6t
Xbit_r151_c148 bl[148] br[148] wl[151] vdd gnd cell_6t
Xbit_r152_c148 bl[148] br[148] wl[152] vdd gnd cell_6t
Xbit_r153_c148 bl[148] br[148] wl[153] vdd gnd cell_6t
Xbit_r154_c148 bl[148] br[148] wl[154] vdd gnd cell_6t
Xbit_r155_c148 bl[148] br[148] wl[155] vdd gnd cell_6t
Xbit_r156_c148 bl[148] br[148] wl[156] vdd gnd cell_6t
Xbit_r157_c148 bl[148] br[148] wl[157] vdd gnd cell_6t
Xbit_r158_c148 bl[148] br[148] wl[158] vdd gnd cell_6t
Xbit_r159_c148 bl[148] br[148] wl[159] vdd gnd cell_6t
Xbit_r160_c148 bl[148] br[148] wl[160] vdd gnd cell_6t
Xbit_r161_c148 bl[148] br[148] wl[161] vdd gnd cell_6t
Xbit_r162_c148 bl[148] br[148] wl[162] vdd gnd cell_6t
Xbit_r163_c148 bl[148] br[148] wl[163] vdd gnd cell_6t
Xbit_r164_c148 bl[148] br[148] wl[164] vdd gnd cell_6t
Xbit_r165_c148 bl[148] br[148] wl[165] vdd gnd cell_6t
Xbit_r166_c148 bl[148] br[148] wl[166] vdd gnd cell_6t
Xbit_r167_c148 bl[148] br[148] wl[167] vdd gnd cell_6t
Xbit_r168_c148 bl[148] br[148] wl[168] vdd gnd cell_6t
Xbit_r169_c148 bl[148] br[148] wl[169] vdd gnd cell_6t
Xbit_r170_c148 bl[148] br[148] wl[170] vdd gnd cell_6t
Xbit_r171_c148 bl[148] br[148] wl[171] vdd gnd cell_6t
Xbit_r172_c148 bl[148] br[148] wl[172] vdd gnd cell_6t
Xbit_r173_c148 bl[148] br[148] wl[173] vdd gnd cell_6t
Xbit_r174_c148 bl[148] br[148] wl[174] vdd gnd cell_6t
Xbit_r175_c148 bl[148] br[148] wl[175] vdd gnd cell_6t
Xbit_r176_c148 bl[148] br[148] wl[176] vdd gnd cell_6t
Xbit_r177_c148 bl[148] br[148] wl[177] vdd gnd cell_6t
Xbit_r178_c148 bl[148] br[148] wl[178] vdd gnd cell_6t
Xbit_r179_c148 bl[148] br[148] wl[179] vdd gnd cell_6t
Xbit_r180_c148 bl[148] br[148] wl[180] vdd gnd cell_6t
Xbit_r181_c148 bl[148] br[148] wl[181] vdd gnd cell_6t
Xbit_r182_c148 bl[148] br[148] wl[182] vdd gnd cell_6t
Xbit_r183_c148 bl[148] br[148] wl[183] vdd gnd cell_6t
Xbit_r184_c148 bl[148] br[148] wl[184] vdd gnd cell_6t
Xbit_r185_c148 bl[148] br[148] wl[185] vdd gnd cell_6t
Xbit_r186_c148 bl[148] br[148] wl[186] vdd gnd cell_6t
Xbit_r187_c148 bl[148] br[148] wl[187] vdd gnd cell_6t
Xbit_r188_c148 bl[148] br[148] wl[188] vdd gnd cell_6t
Xbit_r189_c148 bl[148] br[148] wl[189] vdd gnd cell_6t
Xbit_r190_c148 bl[148] br[148] wl[190] vdd gnd cell_6t
Xbit_r191_c148 bl[148] br[148] wl[191] vdd gnd cell_6t
Xbit_r192_c148 bl[148] br[148] wl[192] vdd gnd cell_6t
Xbit_r193_c148 bl[148] br[148] wl[193] vdd gnd cell_6t
Xbit_r194_c148 bl[148] br[148] wl[194] vdd gnd cell_6t
Xbit_r195_c148 bl[148] br[148] wl[195] vdd gnd cell_6t
Xbit_r196_c148 bl[148] br[148] wl[196] vdd gnd cell_6t
Xbit_r197_c148 bl[148] br[148] wl[197] vdd gnd cell_6t
Xbit_r198_c148 bl[148] br[148] wl[198] vdd gnd cell_6t
Xbit_r199_c148 bl[148] br[148] wl[199] vdd gnd cell_6t
Xbit_r200_c148 bl[148] br[148] wl[200] vdd gnd cell_6t
Xbit_r201_c148 bl[148] br[148] wl[201] vdd gnd cell_6t
Xbit_r202_c148 bl[148] br[148] wl[202] vdd gnd cell_6t
Xbit_r203_c148 bl[148] br[148] wl[203] vdd gnd cell_6t
Xbit_r204_c148 bl[148] br[148] wl[204] vdd gnd cell_6t
Xbit_r205_c148 bl[148] br[148] wl[205] vdd gnd cell_6t
Xbit_r206_c148 bl[148] br[148] wl[206] vdd gnd cell_6t
Xbit_r207_c148 bl[148] br[148] wl[207] vdd gnd cell_6t
Xbit_r208_c148 bl[148] br[148] wl[208] vdd gnd cell_6t
Xbit_r209_c148 bl[148] br[148] wl[209] vdd gnd cell_6t
Xbit_r210_c148 bl[148] br[148] wl[210] vdd gnd cell_6t
Xbit_r211_c148 bl[148] br[148] wl[211] vdd gnd cell_6t
Xbit_r212_c148 bl[148] br[148] wl[212] vdd gnd cell_6t
Xbit_r213_c148 bl[148] br[148] wl[213] vdd gnd cell_6t
Xbit_r214_c148 bl[148] br[148] wl[214] vdd gnd cell_6t
Xbit_r215_c148 bl[148] br[148] wl[215] vdd gnd cell_6t
Xbit_r216_c148 bl[148] br[148] wl[216] vdd gnd cell_6t
Xbit_r217_c148 bl[148] br[148] wl[217] vdd gnd cell_6t
Xbit_r218_c148 bl[148] br[148] wl[218] vdd gnd cell_6t
Xbit_r219_c148 bl[148] br[148] wl[219] vdd gnd cell_6t
Xbit_r220_c148 bl[148] br[148] wl[220] vdd gnd cell_6t
Xbit_r221_c148 bl[148] br[148] wl[221] vdd gnd cell_6t
Xbit_r222_c148 bl[148] br[148] wl[222] vdd gnd cell_6t
Xbit_r223_c148 bl[148] br[148] wl[223] vdd gnd cell_6t
Xbit_r224_c148 bl[148] br[148] wl[224] vdd gnd cell_6t
Xbit_r225_c148 bl[148] br[148] wl[225] vdd gnd cell_6t
Xbit_r226_c148 bl[148] br[148] wl[226] vdd gnd cell_6t
Xbit_r227_c148 bl[148] br[148] wl[227] vdd gnd cell_6t
Xbit_r228_c148 bl[148] br[148] wl[228] vdd gnd cell_6t
Xbit_r229_c148 bl[148] br[148] wl[229] vdd gnd cell_6t
Xbit_r230_c148 bl[148] br[148] wl[230] vdd gnd cell_6t
Xbit_r231_c148 bl[148] br[148] wl[231] vdd gnd cell_6t
Xbit_r232_c148 bl[148] br[148] wl[232] vdd gnd cell_6t
Xbit_r233_c148 bl[148] br[148] wl[233] vdd gnd cell_6t
Xbit_r234_c148 bl[148] br[148] wl[234] vdd gnd cell_6t
Xbit_r235_c148 bl[148] br[148] wl[235] vdd gnd cell_6t
Xbit_r236_c148 bl[148] br[148] wl[236] vdd gnd cell_6t
Xbit_r237_c148 bl[148] br[148] wl[237] vdd gnd cell_6t
Xbit_r238_c148 bl[148] br[148] wl[238] vdd gnd cell_6t
Xbit_r239_c148 bl[148] br[148] wl[239] vdd gnd cell_6t
Xbit_r240_c148 bl[148] br[148] wl[240] vdd gnd cell_6t
Xbit_r241_c148 bl[148] br[148] wl[241] vdd gnd cell_6t
Xbit_r242_c148 bl[148] br[148] wl[242] vdd gnd cell_6t
Xbit_r243_c148 bl[148] br[148] wl[243] vdd gnd cell_6t
Xbit_r244_c148 bl[148] br[148] wl[244] vdd gnd cell_6t
Xbit_r245_c148 bl[148] br[148] wl[245] vdd gnd cell_6t
Xbit_r246_c148 bl[148] br[148] wl[246] vdd gnd cell_6t
Xbit_r247_c148 bl[148] br[148] wl[247] vdd gnd cell_6t
Xbit_r248_c148 bl[148] br[148] wl[248] vdd gnd cell_6t
Xbit_r249_c148 bl[148] br[148] wl[249] vdd gnd cell_6t
Xbit_r250_c148 bl[148] br[148] wl[250] vdd gnd cell_6t
Xbit_r251_c148 bl[148] br[148] wl[251] vdd gnd cell_6t
Xbit_r252_c148 bl[148] br[148] wl[252] vdd gnd cell_6t
Xbit_r253_c148 bl[148] br[148] wl[253] vdd gnd cell_6t
Xbit_r254_c148 bl[148] br[148] wl[254] vdd gnd cell_6t
Xbit_r255_c148 bl[148] br[148] wl[255] vdd gnd cell_6t
Xbit_r0_c149 bl[149] br[149] wl[0] vdd gnd cell_6t
Xbit_r1_c149 bl[149] br[149] wl[1] vdd gnd cell_6t
Xbit_r2_c149 bl[149] br[149] wl[2] vdd gnd cell_6t
Xbit_r3_c149 bl[149] br[149] wl[3] vdd gnd cell_6t
Xbit_r4_c149 bl[149] br[149] wl[4] vdd gnd cell_6t
Xbit_r5_c149 bl[149] br[149] wl[5] vdd gnd cell_6t
Xbit_r6_c149 bl[149] br[149] wl[6] vdd gnd cell_6t
Xbit_r7_c149 bl[149] br[149] wl[7] vdd gnd cell_6t
Xbit_r8_c149 bl[149] br[149] wl[8] vdd gnd cell_6t
Xbit_r9_c149 bl[149] br[149] wl[9] vdd gnd cell_6t
Xbit_r10_c149 bl[149] br[149] wl[10] vdd gnd cell_6t
Xbit_r11_c149 bl[149] br[149] wl[11] vdd gnd cell_6t
Xbit_r12_c149 bl[149] br[149] wl[12] vdd gnd cell_6t
Xbit_r13_c149 bl[149] br[149] wl[13] vdd gnd cell_6t
Xbit_r14_c149 bl[149] br[149] wl[14] vdd gnd cell_6t
Xbit_r15_c149 bl[149] br[149] wl[15] vdd gnd cell_6t
Xbit_r16_c149 bl[149] br[149] wl[16] vdd gnd cell_6t
Xbit_r17_c149 bl[149] br[149] wl[17] vdd gnd cell_6t
Xbit_r18_c149 bl[149] br[149] wl[18] vdd gnd cell_6t
Xbit_r19_c149 bl[149] br[149] wl[19] vdd gnd cell_6t
Xbit_r20_c149 bl[149] br[149] wl[20] vdd gnd cell_6t
Xbit_r21_c149 bl[149] br[149] wl[21] vdd gnd cell_6t
Xbit_r22_c149 bl[149] br[149] wl[22] vdd gnd cell_6t
Xbit_r23_c149 bl[149] br[149] wl[23] vdd gnd cell_6t
Xbit_r24_c149 bl[149] br[149] wl[24] vdd gnd cell_6t
Xbit_r25_c149 bl[149] br[149] wl[25] vdd gnd cell_6t
Xbit_r26_c149 bl[149] br[149] wl[26] vdd gnd cell_6t
Xbit_r27_c149 bl[149] br[149] wl[27] vdd gnd cell_6t
Xbit_r28_c149 bl[149] br[149] wl[28] vdd gnd cell_6t
Xbit_r29_c149 bl[149] br[149] wl[29] vdd gnd cell_6t
Xbit_r30_c149 bl[149] br[149] wl[30] vdd gnd cell_6t
Xbit_r31_c149 bl[149] br[149] wl[31] vdd gnd cell_6t
Xbit_r32_c149 bl[149] br[149] wl[32] vdd gnd cell_6t
Xbit_r33_c149 bl[149] br[149] wl[33] vdd gnd cell_6t
Xbit_r34_c149 bl[149] br[149] wl[34] vdd gnd cell_6t
Xbit_r35_c149 bl[149] br[149] wl[35] vdd gnd cell_6t
Xbit_r36_c149 bl[149] br[149] wl[36] vdd gnd cell_6t
Xbit_r37_c149 bl[149] br[149] wl[37] vdd gnd cell_6t
Xbit_r38_c149 bl[149] br[149] wl[38] vdd gnd cell_6t
Xbit_r39_c149 bl[149] br[149] wl[39] vdd gnd cell_6t
Xbit_r40_c149 bl[149] br[149] wl[40] vdd gnd cell_6t
Xbit_r41_c149 bl[149] br[149] wl[41] vdd gnd cell_6t
Xbit_r42_c149 bl[149] br[149] wl[42] vdd gnd cell_6t
Xbit_r43_c149 bl[149] br[149] wl[43] vdd gnd cell_6t
Xbit_r44_c149 bl[149] br[149] wl[44] vdd gnd cell_6t
Xbit_r45_c149 bl[149] br[149] wl[45] vdd gnd cell_6t
Xbit_r46_c149 bl[149] br[149] wl[46] vdd gnd cell_6t
Xbit_r47_c149 bl[149] br[149] wl[47] vdd gnd cell_6t
Xbit_r48_c149 bl[149] br[149] wl[48] vdd gnd cell_6t
Xbit_r49_c149 bl[149] br[149] wl[49] vdd gnd cell_6t
Xbit_r50_c149 bl[149] br[149] wl[50] vdd gnd cell_6t
Xbit_r51_c149 bl[149] br[149] wl[51] vdd gnd cell_6t
Xbit_r52_c149 bl[149] br[149] wl[52] vdd gnd cell_6t
Xbit_r53_c149 bl[149] br[149] wl[53] vdd gnd cell_6t
Xbit_r54_c149 bl[149] br[149] wl[54] vdd gnd cell_6t
Xbit_r55_c149 bl[149] br[149] wl[55] vdd gnd cell_6t
Xbit_r56_c149 bl[149] br[149] wl[56] vdd gnd cell_6t
Xbit_r57_c149 bl[149] br[149] wl[57] vdd gnd cell_6t
Xbit_r58_c149 bl[149] br[149] wl[58] vdd gnd cell_6t
Xbit_r59_c149 bl[149] br[149] wl[59] vdd gnd cell_6t
Xbit_r60_c149 bl[149] br[149] wl[60] vdd gnd cell_6t
Xbit_r61_c149 bl[149] br[149] wl[61] vdd gnd cell_6t
Xbit_r62_c149 bl[149] br[149] wl[62] vdd gnd cell_6t
Xbit_r63_c149 bl[149] br[149] wl[63] vdd gnd cell_6t
Xbit_r64_c149 bl[149] br[149] wl[64] vdd gnd cell_6t
Xbit_r65_c149 bl[149] br[149] wl[65] vdd gnd cell_6t
Xbit_r66_c149 bl[149] br[149] wl[66] vdd gnd cell_6t
Xbit_r67_c149 bl[149] br[149] wl[67] vdd gnd cell_6t
Xbit_r68_c149 bl[149] br[149] wl[68] vdd gnd cell_6t
Xbit_r69_c149 bl[149] br[149] wl[69] vdd gnd cell_6t
Xbit_r70_c149 bl[149] br[149] wl[70] vdd gnd cell_6t
Xbit_r71_c149 bl[149] br[149] wl[71] vdd gnd cell_6t
Xbit_r72_c149 bl[149] br[149] wl[72] vdd gnd cell_6t
Xbit_r73_c149 bl[149] br[149] wl[73] vdd gnd cell_6t
Xbit_r74_c149 bl[149] br[149] wl[74] vdd gnd cell_6t
Xbit_r75_c149 bl[149] br[149] wl[75] vdd gnd cell_6t
Xbit_r76_c149 bl[149] br[149] wl[76] vdd gnd cell_6t
Xbit_r77_c149 bl[149] br[149] wl[77] vdd gnd cell_6t
Xbit_r78_c149 bl[149] br[149] wl[78] vdd gnd cell_6t
Xbit_r79_c149 bl[149] br[149] wl[79] vdd gnd cell_6t
Xbit_r80_c149 bl[149] br[149] wl[80] vdd gnd cell_6t
Xbit_r81_c149 bl[149] br[149] wl[81] vdd gnd cell_6t
Xbit_r82_c149 bl[149] br[149] wl[82] vdd gnd cell_6t
Xbit_r83_c149 bl[149] br[149] wl[83] vdd gnd cell_6t
Xbit_r84_c149 bl[149] br[149] wl[84] vdd gnd cell_6t
Xbit_r85_c149 bl[149] br[149] wl[85] vdd gnd cell_6t
Xbit_r86_c149 bl[149] br[149] wl[86] vdd gnd cell_6t
Xbit_r87_c149 bl[149] br[149] wl[87] vdd gnd cell_6t
Xbit_r88_c149 bl[149] br[149] wl[88] vdd gnd cell_6t
Xbit_r89_c149 bl[149] br[149] wl[89] vdd gnd cell_6t
Xbit_r90_c149 bl[149] br[149] wl[90] vdd gnd cell_6t
Xbit_r91_c149 bl[149] br[149] wl[91] vdd gnd cell_6t
Xbit_r92_c149 bl[149] br[149] wl[92] vdd gnd cell_6t
Xbit_r93_c149 bl[149] br[149] wl[93] vdd gnd cell_6t
Xbit_r94_c149 bl[149] br[149] wl[94] vdd gnd cell_6t
Xbit_r95_c149 bl[149] br[149] wl[95] vdd gnd cell_6t
Xbit_r96_c149 bl[149] br[149] wl[96] vdd gnd cell_6t
Xbit_r97_c149 bl[149] br[149] wl[97] vdd gnd cell_6t
Xbit_r98_c149 bl[149] br[149] wl[98] vdd gnd cell_6t
Xbit_r99_c149 bl[149] br[149] wl[99] vdd gnd cell_6t
Xbit_r100_c149 bl[149] br[149] wl[100] vdd gnd cell_6t
Xbit_r101_c149 bl[149] br[149] wl[101] vdd gnd cell_6t
Xbit_r102_c149 bl[149] br[149] wl[102] vdd gnd cell_6t
Xbit_r103_c149 bl[149] br[149] wl[103] vdd gnd cell_6t
Xbit_r104_c149 bl[149] br[149] wl[104] vdd gnd cell_6t
Xbit_r105_c149 bl[149] br[149] wl[105] vdd gnd cell_6t
Xbit_r106_c149 bl[149] br[149] wl[106] vdd gnd cell_6t
Xbit_r107_c149 bl[149] br[149] wl[107] vdd gnd cell_6t
Xbit_r108_c149 bl[149] br[149] wl[108] vdd gnd cell_6t
Xbit_r109_c149 bl[149] br[149] wl[109] vdd gnd cell_6t
Xbit_r110_c149 bl[149] br[149] wl[110] vdd gnd cell_6t
Xbit_r111_c149 bl[149] br[149] wl[111] vdd gnd cell_6t
Xbit_r112_c149 bl[149] br[149] wl[112] vdd gnd cell_6t
Xbit_r113_c149 bl[149] br[149] wl[113] vdd gnd cell_6t
Xbit_r114_c149 bl[149] br[149] wl[114] vdd gnd cell_6t
Xbit_r115_c149 bl[149] br[149] wl[115] vdd gnd cell_6t
Xbit_r116_c149 bl[149] br[149] wl[116] vdd gnd cell_6t
Xbit_r117_c149 bl[149] br[149] wl[117] vdd gnd cell_6t
Xbit_r118_c149 bl[149] br[149] wl[118] vdd gnd cell_6t
Xbit_r119_c149 bl[149] br[149] wl[119] vdd gnd cell_6t
Xbit_r120_c149 bl[149] br[149] wl[120] vdd gnd cell_6t
Xbit_r121_c149 bl[149] br[149] wl[121] vdd gnd cell_6t
Xbit_r122_c149 bl[149] br[149] wl[122] vdd gnd cell_6t
Xbit_r123_c149 bl[149] br[149] wl[123] vdd gnd cell_6t
Xbit_r124_c149 bl[149] br[149] wl[124] vdd gnd cell_6t
Xbit_r125_c149 bl[149] br[149] wl[125] vdd gnd cell_6t
Xbit_r126_c149 bl[149] br[149] wl[126] vdd gnd cell_6t
Xbit_r127_c149 bl[149] br[149] wl[127] vdd gnd cell_6t
Xbit_r128_c149 bl[149] br[149] wl[128] vdd gnd cell_6t
Xbit_r129_c149 bl[149] br[149] wl[129] vdd gnd cell_6t
Xbit_r130_c149 bl[149] br[149] wl[130] vdd gnd cell_6t
Xbit_r131_c149 bl[149] br[149] wl[131] vdd gnd cell_6t
Xbit_r132_c149 bl[149] br[149] wl[132] vdd gnd cell_6t
Xbit_r133_c149 bl[149] br[149] wl[133] vdd gnd cell_6t
Xbit_r134_c149 bl[149] br[149] wl[134] vdd gnd cell_6t
Xbit_r135_c149 bl[149] br[149] wl[135] vdd gnd cell_6t
Xbit_r136_c149 bl[149] br[149] wl[136] vdd gnd cell_6t
Xbit_r137_c149 bl[149] br[149] wl[137] vdd gnd cell_6t
Xbit_r138_c149 bl[149] br[149] wl[138] vdd gnd cell_6t
Xbit_r139_c149 bl[149] br[149] wl[139] vdd gnd cell_6t
Xbit_r140_c149 bl[149] br[149] wl[140] vdd gnd cell_6t
Xbit_r141_c149 bl[149] br[149] wl[141] vdd gnd cell_6t
Xbit_r142_c149 bl[149] br[149] wl[142] vdd gnd cell_6t
Xbit_r143_c149 bl[149] br[149] wl[143] vdd gnd cell_6t
Xbit_r144_c149 bl[149] br[149] wl[144] vdd gnd cell_6t
Xbit_r145_c149 bl[149] br[149] wl[145] vdd gnd cell_6t
Xbit_r146_c149 bl[149] br[149] wl[146] vdd gnd cell_6t
Xbit_r147_c149 bl[149] br[149] wl[147] vdd gnd cell_6t
Xbit_r148_c149 bl[149] br[149] wl[148] vdd gnd cell_6t
Xbit_r149_c149 bl[149] br[149] wl[149] vdd gnd cell_6t
Xbit_r150_c149 bl[149] br[149] wl[150] vdd gnd cell_6t
Xbit_r151_c149 bl[149] br[149] wl[151] vdd gnd cell_6t
Xbit_r152_c149 bl[149] br[149] wl[152] vdd gnd cell_6t
Xbit_r153_c149 bl[149] br[149] wl[153] vdd gnd cell_6t
Xbit_r154_c149 bl[149] br[149] wl[154] vdd gnd cell_6t
Xbit_r155_c149 bl[149] br[149] wl[155] vdd gnd cell_6t
Xbit_r156_c149 bl[149] br[149] wl[156] vdd gnd cell_6t
Xbit_r157_c149 bl[149] br[149] wl[157] vdd gnd cell_6t
Xbit_r158_c149 bl[149] br[149] wl[158] vdd gnd cell_6t
Xbit_r159_c149 bl[149] br[149] wl[159] vdd gnd cell_6t
Xbit_r160_c149 bl[149] br[149] wl[160] vdd gnd cell_6t
Xbit_r161_c149 bl[149] br[149] wl[161] vdd gnd cell_6t
Xbit_r162_c149 bl[149] br[149] wl[162] vdd gnd cell_6t
Xbit_r163_c149 bl[149] br[149] wl[163] vdd gnd cell_6t
Xbit_r164_c149 bl[149] br[149] wl[164] vdd gnd cell_6t
Xbit_r165_c149 bl[149] br[149] wl[165] vdd gnd cell_6t
Xbit_r166_c149 bl[149] br[149] wl[166] vdd gnd cell_6t
Xbit_r167_c149 bl[149] br[149] wl[167] vdd gnd cell_6t
Xbit_r168_c149 bl[149] br[149] wl[168] vdd gnd cell_6t
Xbit_r169_c149 bl[149] br[149] wl[169] vdd gnd cell_6t
Xbit_r170_c149 bl[149] br[149] wl[170] vdd gnd cell_6t
Xbit_r171_c149 bl[149] br[149] wl[171] vdd gnd cell_6t
Xbit_r172_c149 bl[149] br[149] wl[172] vdd gnd cell_6t
Xbit_r173_c149 bl[149] br[149] wl[173] vdd gnd cell_6t
Xbit_r174_c149 bl[149] br[149] wl[174] vdd gnd cell_6t
Xbit_r175_c149 bl[149] br[149] wl[175] vdd gnd cell_6t
Xbit_r176_c149 bl[149] br[149] wl[176] vdd gnd cell_6t
Xbit_r177_c149 bl[149] br[149] wl[177] vdd gnd cell_6t
Xbit_r178_c149 bl[149] br[149] wl[178] vdd gnd cell_6t
Xbit_r179_c149 bl[149] br[149] wl[179] vdd gnd cell_6t
Xbit_r180_c149 bl[149] br[149] wl[180] vdd gnd cell_6t
Xbit_r181_c149 bl[149] br[149] wl[181] vdd gnd cell_6t
Xbit_r182_c149 bl[149] br[149] wl[182] vdd gnd cell_6t
Xbit_r183_c149 bl[149] br[149] wl[183] vdd gnd cell_6t
Xbit_r184_c149 bl[149] br[149] wl[184] vdd gnd cell_6t
Xbit_r185_c149 bl[149] br[149] wl[185] vdd gnd cell_6t
Xbit_r186_c149 bl[149] br[149] wl[186] vdd gnd cell_6t
Xbit_r187_c149 bl[149] br[149] wl[187] vdd gnd cell_6t
Xbit_r188_c149 bl[149] br[149] wl[188] vdd gnd cell_6t
Xbit_r189_c149 bl[149] br[149] wl[189] vdd gnd cell_6t
Xbit_r190_c149 bl[149] br[149] wl[190] vdd gnd cell_6t
Xbit_r191_c149 bl[149] br[149] wl[191] vdd gnd cell_6t
Xbit_r192_c149 bl[149] br[149] wl[192] vdd gnd cell_6t
Xbit_r193_c149 bl[149] br[149] wl[193] vdd gnd cell_6t
Xbit_r194_c149 bl[149] br[149] wl[194] vdd gnd cell_6t
Xbit_r195_c149 bl[149] br[149] wl[195] vdd gnd cell_6t
Xbit_r196_c149 bl[149] br[149] wl[196] vdd gnd cell_6t
Xbit_r197_c149 bl[149] br[149] wl[197] vdd gnd cell_6t
Xbit_r198_c149 bl[149] br[149] wl[198] vdd gnd cell_6t
Xbit_r199_c149 bl[149] br[149] wl[199] vdd gnd cell_6t
Xbit_r200_c149 bl[149] br[149] wl[200] vdd gnd cell_6t
Xbit_r201_c149 bl[149] br[149] wl[201] vdd gnd cell_6t
Xbit_r202_c149 bl[149] br[149] wl[202] vdd gnd cell_6t
Xbit_r203_c149 bl[149] br[149] wl[203] vdd gnd cell_6t
Xbit_r204_c149 bl[149] br[149] wl[204] vdd gnd cell_6t
Xbit_r205_c149 bl[149] br[149] wl[205] vdd gnd cell_6t
Xbit_r206_c149 bl[149] br[149] wl[206] vdd gnd cell_6t
Xbit_r207_c149 bl[149] br[149] wl[207] vdd gnd cell_6t
Xbit_r208_c149 bl[149] br[149] wl[208] vdd gnd cell_6t
Xbit_r209_c149 bl[149] br[149] wl[209] vdd gnd cell_6t
Xbit_r210_c149 bl[149] br[149] wl[210] vdd gnd cell_6t
Xbit_r211_c149 bl[149] br[149] wl[211] vdd gnd cell_6t
Xbit_r212_c149 bl[149] br[149] wl[212] vdd gnd cell_6t
Xbit_r213_c149 bl[149] br[149] wl[213] vdd gnd cell_6t
Xbit_r214_c149 bl[149] br[149] wl[214] vdd gnd cell_6t
Xbit_r215_c149 bl[149] br[149] wl[215] vdd gnd cell_6t
Xbit_r216_c149 bl[149] br[149] wl[216] vdd gnd cell_6t
Xbit_r217_c149 bl[149] br[149] wl[217] vdd gnd cell_6t
Xbit_r218_c149 bl[149] br[149] wl[218] vdd gnd cell_6t
Xbit_r219_c149 bl[149] br[149] wl[219] vdd gnd cell_6t
Xbit_r220_c149 bl[149] br[149] wl[220] vdd gnd cell_6t
Xbit_r221_c149 bl[149] br[149] wl[221] vdd gnd cell_6t
Xbit_r222_c149 bl[149] br[149] wl[222] vdd gnd cell_6t
Xbit_r223_c149 bl[149] br[149] wl[223] vdd gnd cell_6t
Xbit_r224_c149 bl[149] br[149] wl[224] vdd gnd cell_6t
Xbit_r225_c149 bl[149] br[149] wl[225] vdd gnd cell_6t
Xbit_r226_c149 bl[149] br[149] wl[226] vdd gnd cell_6t
Xbit_r227_c149 bl[149] br[149] wl[227] vdd gnd cell_6t
Xbit_r228_c149 bl[149] br[149] wl[228] vdd gnd cell_6t
Xbit_r229_c149 bl[149] br[149] wl[229] vdd gnd cell_6t
Xbit_r230_c149 bl[149] br[149] wl[230] vdd gnd cell_6t
Xbit_r231_c149 bl[149] br[149] wl[231] vdd gnd cell_6t
Xbit_r232_c149 bl[149] br[149] wl[232] vdd gnd cell_6t
Xbit_r233_c149 bl[149] br[149] wl[233] vdd gnd cell_6t
Xbit_r234_c149 bl[149] br[149] wl[234] vdd gnd cell_6t
Xbit_r235_c149 bl[149] br[149] wl[235] vdd gnd cell_6t
Xbit_r236_c149 bl[149] br[149] wl[236] vdd gnd cell_6t
Xbit_r237_c149 bl[149] br[149] wl[237] vdd gnd cell_6t
Xbit_r238_c149 bl[149] br[149] wl[238] vdd gnd cell_6t
Xbit_r239_c149 bl[149] br[149] wl[239] vdd gnd cell_6t
Xbit_r240_c149 bl[149] br[149] wl[240] vdd gnd cell_6t
Xbit_r241_c149 bl[149] br[149] wl[241] vdd gnd cell_6t
Xbit_r242_c149 bl[149] br[149] wl[242] vdd gnd cell_6t
Xbit_r243_c149 bl[149] br[149] wl[243] vdd gnd cell_6t
Xbit_r244_c149 bl[149] br[149] wl[244] vdd gnd cell_6t
Xbit_r245_c149 bl[149] br[149] wl[245] vdd gnd cell_6t
Xbit_r246_c149 bl[149] br[149] wl[246] vdd gnd cell_6t
Xbit_r247_c149 bl[149] br[149] wl[247] vdd gnd cell_6t
Xbit_r248_c149 bl[149] br[149] wl[248] vdd gnd cell_6t
Xbit_r249_c149 bl[149] br[149] wl[249] vdd gnd cell_6t
Xbit_r250_c149 bl[149] br[149] wl[250] vdd gnd cell_6t
Xbit_r251_c149 bl[149] br[149] wl[251] vdd gnd cell_6t
Xbit_r252_c149 bl[149] br[149] wl[252] vdd gnd cell_6t
Xbit_r253_c149 bl[149] br[149] wl[253] vdd gnd cell_6t
Xbit_r254_c149 bl[149] br[149] wl[254] vdd gnd cell_6t
Xbit_r255_c149 bl[149] br[149] wl[255] vdd gnd cell_6t
Xbit_r0_c150 bl[150] br[150] wl[0] vdd gnd cell_6t
Xbit_r1_c150 bl[150] br[150] wl[1] vdd gnd cell_6t
Xbit_r2_c150 bl[150] br[150] wl[2] vdd gnd cell_6t
Xbit_r3_c150 bl[150] br[150] wl[3] vdd gnd cell_6t
Xbit_r4_c150 bl[150] br[150] wl[4] vdd gnd cell_6t
Xbit_r5_c150 bl[150] br[150] wl[5] vdd gnd cell_6t
Xbit_r6_c150 bl[150] br[150] wl[6] vdd gnd cell_6t
Xbit_r7_c150 bl[150] br[150] wl[7] vdd gnd cell_6t
Xbit_r8_c150 bl[150] br[150] wl[8] vdd gnd cell_6t
Xbit_r9_c150 bl[150] br[150] wl[9] vdd gnd cell_6t
Xbit_r10_c150 bl[150] br[150] wl[10] vdd gnd cell_6t
Xbit_r11_c150 bl[150] br[150] wl[11] vdd gnd cell_6t
Xbit_r12_c150 bl[150] br[150] wl[12] vdd gnd cell_6t
Xbit_r13_c150 bl[150] br[150] wl[13] vdd gnd cell_6t
Xbit_r14_c150 bl[150] br[150] wl[14] vdd gnd cell_6t
Xbit_r15_c150 bl[150] br[150] wl[15] vdd gnd cell_6t
Xbit_r16_c150 bl[150] br[150] wl[16] vdd gnd cell_6t
Xbit_r17_c150 bl[150] br[150] wl[17] vdd gnd cell_6t
Xbit_r18_c150 bl[150] br[150] wl[18] vdd gnd cell_6t
Xbit_r19_c150 bl[150] br[150] wl[19] vdd gnd cell_6t
Xbit_r20_c150 bl[150] br[150] wl[20] vdd gnd cell_6t
Xbit_r21_c150 bl[150] br[150] wl[21] vdd gnd cell_6t
Xbit_r22_c150 bl[150] br[150] wl[22] vdd gnd cell_6t
Xbit_r23_c150 bl[150] br[150] wl[23] vdd gnd cell_6t
Xbit_r24_c150 bl[150] br[150] wl[24] vdd gnd cell_6t
Xbit_r25_c150 bl[150] br[150] wl[25] vdd gnd cell_6t
Xbit_r26_c150 bl[150] br[150] wl[26] vdd gnd cell_6t
Xbit_r27_c150 bl[150] br[150] wl[27] vdd gnd cell_6t
Xbit_r28_c150 bl[150] br[150] wl[28] vdd gnd cell_6t
Xbit_r29_c150 bl[150] br[150] wl[29] vdd gnd cell_6t
Xbit_r30_c150 bl[150] br[150] wl[30] vdd gnd cell_6t
Xbit_r31_c150 bl[150] br[150] wl[31] vdd gnd cell_6t
Xbit_r32_c150 bl[150] br[150] wl[32] vdd gnd cell_6t
Xbit_r33_c150 bl[150] br[150] wl[33] vdd gnd cell_6t
Xbit_r34_c150 bl[150] br[150] wl[34] vdd gnd cell_6t
Xbit_r35_c150 bl[150] br[150] wl[35] vdd gnd cell_6t
Xbit_r36_c150 bl[150] br[150] wl[36] vdd gnd cell_6t
Xbit_r37_c150 bl[150] br[150] wl[37] vdd gnd cell_6t
Xbit_r38_c150 bl[150] br[150] wl[38] vdd gnd cell_6t
Xbit_r39_c150 bl[150] br[150] wl[39] vdd gnd cell_6t
Xbit_r40_c150 bl[150] br[150] wl[40] vdd gnd cell_6t
Xbit_r41_c150 bl[150] br[150] wl[41] vdd gnd cell_6t
Xbit_r42_c150 bl[150] br[150] wl[42] vdd gnd cell_6t
Xbit_r43_c150 bl[150] br[150] wl[43] vdd gnd cell_6t
Xbit_r44_c150 bl[150] br[150] wl[44] vdd gnd cell_6t
Xbit_r45_c150 bl[150] br[150] wl[45] vdd gnd cell_6t
Xbit_r46_c150 bl[150] br[150] wl[46] vdd gnd cell_6t
Xbit_r47_c150 bl[150] br[150] wl[47] vdd gnd cell_6t
Xbit_r48_c150 bl[150] br[150] wl[48] vdd gnd cell_6t
Xbit_r49_c150 bl[150] br[150] wl[49] vdd gnd cell_6t
Xbit_r50_c150 bl[150] br[150] wl[50] vdd gnd cell_6t
Xbit_r51_c150 bl[150] br[150] wl[51] vdd gnd cell_6t
Xbit_r52_c150 bl[150] br[150] wl[52] vdd gnd cell_6t
Xbit_r53_c150 bl[150] br[150] wl[53] vdd gnd cell_6t
Xbit_r54_c150 bl[150] br[150] wl[54] vdd gnd cell_6t
Xbit_r55_c150 bl[150] br[150] wl[55] vdd gnd cell_6t
Xbit_r56_c150 bl[150] br[150] wl[56] vdd gnd cell_6t
Xbit_r57_c150 bl[150] br[150] wl[57] vdd gnd cell_6t
Xbit_r58_c150 bl[150] br[150] wl[58] vdd gnd cell_6t
Xbit_r59_c150 bl[150] br[150] wl[59] vdd gnd cell_6t
Xbit_r60_c150 bl[150] br[150] wl[60] vdd gnd cell_6t
Xbit_r61_c150 bl[150] br[150] wl[61] vdd gnd cell_6t
Xbit_r62_c150 bl[150] br[150] wl[62] vdd gnd cell_6t
Xbit_r63_c150 bl[150] br[150] wl[63] vdd gnd cell_6t
Xbit_r64_c150 bl[150] br[150] wl[64] vdd gnd cell_6t
Xbit_r65_c150 bl[150] br[150] wl[65] vdd gnd cell_6t
Xbit_r66_c150 bl[150] br[150] wl[66] vdd gnd cell_6t
Xbit_r67_c150 bl[150] br[150] wl[67] vdd gnd cell_6t
Xbit_r68_c150 bl[150] br[150] wl[68] vdd gnd cell_6t
Xbit_r69_c150 bl[150] br[150] wl[69] vdd gnd cell_6t
Xbit_r70_c150 bl[150] br[150] wl[70] vdd gnd cell_6t
Xbit_r71_c150 bl[150] br[150] wl[71] vdd gnd cell_6t
Xbit_r72_c150 bl[150] br[150] wl[72] vdd gnd cell_6t
Xbit_r73_c150 bl[150] br[150] wl[73] vdd gnd cell_6t
Xbit_r74_c150 bl[150] br[150] wl[74] vdd gnd cell_6t
Xbit_r75_c150 bl[150] br[150] wl[75] vdd gnd cell_6t
Xbit_r76_c150 bl[150] br[150] wl[76] vdd gnd cell_6t
Xbit_r77_c150 bl[150] br[150] wl[77] vdd gnd cell_6t
Xbit_r78_c150 bl[150] br[150] wl[78] vdd gnd cell_6t
Xbit_r79_c150 bl[150] br[150] wl[79] vdd gnd cell_6t
Xbit_r80_c150 bl[150] br[150] wl[80] vdd gnd cell_6t
Xbit_r81_c150 bl[150] br[150] wl[81] vdd gnd cell_6t
Xbit_r82_c150 bl[150] br[150] wl[82] vdd gnd cell_6t
Xbit_r83_c150 bl[150] br[150] wl[83] vdd gnd cell_6t
Xbit_r84_c150 bl[150] br[150] wl[84] vdd gnd cell_6t
Xbit_r85_c150 bl[150] br[150] wl[85] vdd gnd cell_6t
Xbit_r86_c150 bl[150] br[150] wl[86] vdd gnd cell_6t
Xbit_r87_c150 bl[150] br[150] wl[87] vdd gnd cell_6t
Xbit_r88_c150 bl[150] br[150] wl[88] vdd gnd cell_6t
Xbit_r89_c150 bl[150] br[150] wl[89] vdd gnd cell_6t
Xbit_r90_c150 bl[150] br[150] wl[90] vdd gnd cell_6t
Xbit_r91_c150 bl[150] br[150] wl[91] vdd gnd cell_6t
Xbit_r92_c150 bl[150] br[150] wl[92] vdd gnd cell_6t
Xbit_r93_c150 bl[150] br[150] wl[93] vdd gnd cell_6t
Xbit_r94_c150 bl[150] br[150] wl[94] vdd gnd cell_6t
Xbit_r95_c150 bl[150] br[150] wl[95] vdd gnd cell_6t
Xbit_r96_c150 bl[150] br[150] wl[96] vdd gnd cell_6t
Xbit_r97_c150 bl[150] br[150] wl[97] vdd gnd cell_6t
Xbit_r98_c150 bl[150] br[150] wl[98] vdd gnd cell_6t
Xbit_r99_c150 bl[150] br[150] wl[99] vdd gnd cell_6t
Xbit_r100_c150 bl[150] br[150] wl[100] vdd gnd cell_6t
Xbit_r101_c150 bl[150] br[150] wl[101] vdd gnd cell_6t
Xbit_r102_c150 bl[150] br[150] wl[102] vdd gnd cell_6t
Xbit_r103_c150 bl[150] br[150] wl[103] vdd gnd cell_6t
Xbit_r104_c150 bl[150] br[150] wl[104] vdd gnd cell_6t
Xbit_r105_c150 bl[150] br[150] wl[105] vdd gnd cell_6t
Xbit_r106_c150 bl[150] br[150] wl[106] vdd gnd cell_6t
Xbit_r107_c150 bl[150] br[150] wl[107] vdd gnd cell_6t
Xbit_r108_c150 bl[150] br[150] wl[108] vdd gnd cell_6t
Xbit_r109_c150 bl[150] br[150] wl[109] vdd gnd cell_6t
Xbit_r110_c150 bl[150] br[150] wl[110] vdd gnd cell_6t
Xbit_r111_c150 bl[150] br[150] wl[111] vdd gnd cell_6t
Xbit_r112_c150 bl[150] br[150] wl[112] vdd gnd cell_6t
Xbit_r113_c150 bl[150] br[150] wl[113] vdd gnd cell_6t
Xbit_r114_c150 bl[150] br[150] wl[114] vdd gnd cell_6t
Xbit_r115_c150 bl[150] br[150] wl[115] vdd gnd cell_6t
Xbit_r116_c150 bl[150] br[150] wl[116] vdd gnd cell_6t
Xbit_r117_c150 bl[150] br[150] wl[117] vdd gnd cell_6t
Xbit_r118_c150 bl[150] br[150] wl[118] vdd gnd cell_6t
Xbit_r119_c150 bl[150] br[150] wl[119] vdd gnd cell_6t
Xbit_r120_c150 bl[150] br[150] wl[120] vdd gnd cell_6t
Xbit_r121_c150 bl[150] br[150] wl[121] vdd gnd cell_6t
Xbit_r122_c150 bl[150] br[150] wl[122] vdd gnd cell_6t
Xbit_r123_c150 bl[150] br[150] wl[123] vdd gnd cell_6t
Xbit_r124_c150 bl[150] br[150] wl[124] vdd gnd cell_6t
Xbit_r125_c150 bl[150] br[150] wl[125] vdd gnd cell_6t
Xbit_r126_c150 bl[150] br[150] wl[126] vdd gnd cell_6t
Xbit_r127_c150 bl[150] br[150] wl[127] vdd gnd cell_6t
Xbit_r128_c150 bl[150] br[150] wl[128] vdd gnd cell_6t
Xbit_r129_c150 bl[150] br[150] wl[129] vdd gnd cell_6t
Xbit_r130_c150 bl[150] br[150] wl[130] vdd gnd cell_6t
Xbit_r131_c150 bl[150] br[150] wl[131] vdd gnd cell_6t
Xbit_r132_c150 bl[150] br[150] wl[132] vdd gnd cell_6t
Xbit_r133_c150 bl[150] br[150] wl[133] vdd gnd cell_6t
Xbit_r134_c150 bl[150] br[150] wl[134] vdd gnd cell_6t
Xbit_r135_c150 bl[150] br[150] wl[135] vdd gnd cell_6t
Xbit_r136_c150 bl[150] br[150] wl[136] vdd gnd cell_6t
Xbit_r137_c150 bl[150] br[150] wl[137] vdd gnd cell_6t
Xbit_r138_c150 bl[150] br[150] wl[138] vdd gnd cell_6t
Xbit_r139_c150 bl[150] br[150] wl[139] vdd gnd cell_6t
Xbit_r140_c150 bl[150] br[150] wl[140] vdd gnd cell_6t
Xbit_r141_c150 bl[150] br[150] wl[141] vdd gnd cell_6t
Xbit_r142_c150 bl[150] br[150] wl[142] vdd gnd cell_6t
Xbit_r143_c150 bl[150] br[150] wl[143] vdd gnd cell_6t
Xbit_r144_c150 bl[150] br[150] wl[144] vdd gnd cell_6t
Xbit_r145_c150 bl[150] br[150] wl[145] vdd gnd cell_6t
Xbit_r146_c150 bl[150] br[150] wl[146] vdd gnd cell_6t
Xbit_r147_c150 bl[150] br[150] wl[147] vdd gnd cell_6t
Xbit_r148_c150 bl[150] br[150] wl[148] vdd gnd cell_6t
Xbit_r149_c150 bl[150] br[150] wl[149] vdd gnd cell_6t
Xbit_r150_c150 bl[150] br[150] wl[150] vdd gnd cell_6t
Xbit_r151_c150 bl[150] br[150] wl[151] vdd gnd cell_6t
Xbit_r152_c150 bl[150] br[150] wl[152] vdd gnd cell_6t
Xbit_r153_c150 bl[150] br[150] wl[153] vdd gnd cell_6t
Xbit_r154_c150 bl[150] br[150] wl[154] vdd gnd cell_6t
Xbit_r155_c150 bl[150] br[150] wl[155] vdd gnd cell_6t
Xbit_r156_c150 bl[150] br[150] wl[156] vdd gnd cell_6t
Xbit_r157_c150 bl[150] br[150] wl[157] vdd gnd cell_6t
Xbit_r158_c150 bl[150] br[150] wl[158] vdd gnd cell_6t
Xbit_r159_c150 bl[150] br[150] wl[159] vdd gnd cell_6t
Xbit_r160_c150 bl[150] br[150] wl[160] vdd gnd cell_6t
Xbit_r161_c150 bl[150] br[150] wl[161] vdd gnd cell_6t
Xbit_r162_c150 bl[150] br[150] wl[162] vdd gnd cell_6t
Xbit_r163_c150 bl[150] br[150] wl[163] vdd gnd cell_6t
Xbit_r164_c150 bl[150] br[150] wl[164] vdd gnd cell_6t
Xbit_r165_c150 bl[150] br[150] wl[165] vdd gnd cell_6t
Xbit_r166_c150 bl[150] br[150] wl[166] vdd gnd cell_6t
Xbit_r167_c150 bl[150] br[150] wl[167] vdd gnd cell_6t
Xbit_r168_c150 bl[150] br[150] wl[168] vdd gnd cell_6t
Xbit_r169_c150 bl[150] br[150] wl[169] vdd gnd cell_6t
Xbit_r170_c150 bl[150] br[150] wl[170] vdd gnd cell_6t
Xbit_r171_c150 bl[150] br[150] wl[171] vdd gnd cell_6t
Xbit_r172_c150 bl[150] br[150] wl[172] vdd gnd cell_6t
Xbit_r173_c150 bl[150] br[150] wl[173] vdd gnd cell_6t
Xbit_r174_c150 bl[150] br[150] wl[174] vdd gnd cell_6t
Xbit_r175_c150 bl[150] br[150] wl[175] vdd gnd cell_6t
Xbit_r176_c150 bl[150] br[150] wl[176] vdd gnd cell_6t
Xbit_r177_c150 bl[150] br[150] wl[177] vdd gnd cell_6t
Xbit_r178_c150 bl[150] br[150] wl[178] vdd gnd cell_6t
Xbit_r179_c150 bl[150] br[150] wl[179] vdd gnd cell_6t
Xbit_r180_c150 bl[150] br[150] wl[180] vdd gnd cell_6t
Xbit_r181_c150 bl[150] br[150] wl[181] vdd gnd cell_6t
Xbit_r182_c150 bl[150] br[150] wl[182] vdd gnd cell_6t
Xbit_r183_c150 bl[150] br[150] wl[183] vdd gnd cell_6t
Xbit_r184_c150 bl[150] br[150] wl[184] vdd gnd cell_6t
Xbit_r185_c150 bl[150] br[150] wl[185] vdd gnd cell_6t
Xbit_r186_c150 bl[150] br[150] wl[186] vdd gnd cell_6t
Xbit_r187_c150 bl[150] br[150] wl[187] vdd gnd cell_6t
Xbit_r188_c150 bl[150] br[150] wl[188] vdd gnd cell_6t
Xbit_r189_c150 bl[150] br[150] wl[189] vdd gnd cell_6t
Xbit_r190_c150 bl[150] br[150] wl[190] vdd gnd cell_6t
Xbit_r191_c150 bl[150] br[150] wl[191] vdd gnd cell_6t
Xbit_r192_c150 bl[150] br[150] wl[192] vdd gnd cell_6t
Xbit_r193_c150 bl[150] br[150] wl[193] vdd gnd cell_6t
Xbit_r194_c150 bl[150] br[150] wl[194] vdd gnd cell_6t
Xbit_r195_c150 bl[150] br[150] wl[195] vdd gnd cell_6t
Xbit_r196_c150 bl[150] br[150] wl[196] vdd gnd cell_6t
Xbit_r197_c150 bl[150] br[150] wl[197] vdd gnd cell_6t
Xbit_r198_c150 bl[150] br[150] wl[198] vdd gnd cell_6t
Xbit_r199_c150 bl[150] br[150] wl[199] vdd gnd cell_6t
Xbit_r200_c150 bl[150] br[150] wl[200] vdd gnd cell_6t
Xbit_r201_c150 bl[150] br[150] wl[201] vdd gnd cell_6t
Xbit_r202_c150 bl[150] br[150] wl[202] vdd gnd cell_6t
Xbit_r203_c150 bl[150] br[150] wl[203] vdd gnd cell_6t
Xbit_r204_c150 bl[150] br[150] wl[204] vdd gnd cell_6t
Xbit_r205_c150 bl[150] br[150] wl[205] vdd gnd cell_6t
Xbit_r206_c150 bl[150] br[150] wl[206] vdd gnd cell_6t
Xbit_r207_c150 bl[150] br[150] wl[207] vdd gnd cell_6t
Xbit_r208_c150 bl[150] br[150] wl[208] vdd gnd cell_6t
Xbit_r209_c150 bl[150] br[150] wl[209] vdd gnd cell_6t
Xbit_r210_c150 bl[150] br[150] wl[210] vdd gnd cell_6t
Xbit_r211_c150 bl[150] br[150] wl[211] vdd gnd cell_6t
Xbit_r212_c150 bl[150] br[150] wl[212] vdd gnd cell_6t
Xbit_r213_c150 bl[150] br[150] wl[213] vdd gnd cell_6t
Xbit_r214_c150 bl[150] br[150] wl[214] vdd gnd cell_6t
Xbit_r215_c150 bl[150] br[150] wl[215] vdd gnd cell_6t
Xbit_r216_c150 bl[150] br[150] wl[216] vdd gnd cell_6t
Xbit_r217_c150 bl[150] br[150] wl[217] vdd gnd cell_6t
Xbit_r218_c150 bl[150] br[150] wl[218] vdd gnd cell_6t
Xbit_r219_c150 bl[150] br[150] wl[219] vdd gnd cell_6t
Xbit_r220_c150 bl[150] br[150] wl[220] vdd gnd cell_6t
Xbit_r221_c150 bl[150] br[150] wl[221] vdd gnd cell_6t
Xbit_r222_c150 bl[150] br[150] wl[222] vdd gnd cell_6t
Xbit_r223_c150 bl[150] br[150] wl[223] vdd gnd cell_6t
Xbit_r224_c150 bl[150] br[150] wl[224] vdd gnd cell_6t
Xbit_r225_c150 bl[150] br[150] wl[225] vdd gnd cell_6t
Xbit_r226_c150 bl[150] br[150] wl[226] vdd gnd cell_6t
Xbit_r227_c150 bl[150] br[150] wl[227] vdd gnd cell_6t
Xbit_r228_c150 bl[150] br[150] wl[228] vdd gnd cell_6t
Xbit_r229_c150 bl[150] br[150] wl[229] vdd gnd cell_6t
Xbit_r230_c150 bl[150] br[150] wl[230] vdd gnd cell_6t
Xbit_r231_c150 bl[150] br[150] wl[231] vdd gnd cell_6t
Xbit_r232_c150 bl[150] br[150] wl[232] vdd gnd cell_6t
Xbit_r233_c150 bl[150] br[150] wl[233] vdd gnd cell_6t
Xbit_r234_c150 bl[150] br[150] wl[234] vdd gnd cell_6t
Xbit_r235_c150 bl[150] br[150] wl[235] vdd gnd cell_6t
Xbit_r236_c150 bl[150] br[150] wl[236] vdd gnd cell_6t
Xbit_r237_c150 bl[150] br[150] wl[237] vdd gnd cell_6t
Xbit_r238_c150 bl[150] br[150] wl[238] vdd gnd cell_6t
Xbit_r239_c150 bl[150] br[150] wl[239] vdd gnd cell_6t
Xbit_r240_c150 bl[150] br[150] wl[240] vdd gnd cell_6t
Xbit_r241_c150 bl[150] br[150] wl[241] vdd gnd cell_6t
Xbit_r242_c150 bl[150] br[150] wl[242] vdd gnd cell_6t
Xbit_r243_c150 bl[150] br[150] wl[243] vdd gnd cell_6t
Xbit_r244_c150 bl[150] br[150] wl[244] vdd gnd cell_6t
Xbit_r245_c150 bl[150] br[150] wl[245] vdd gnd cell_6t
Xbit_r246_c150 bl[150] br[150] wl[246] vdd gnd cell_6t
Xbit_r247_c150 bl[150] br[150] wl[247] vdd gnd cell_6t
Xbit_r248_c150 bl[150] br[150] wl[248] vdd gnd cell_6t
Xbit_r249_c150 bl[150] br[150] wl[249] vdd gnd cell_6t
Xbit_r250_c150 bl[150] br[150] wl[250] vdd gnd cell_6t
Xbit_r251_c150 bl[150] br[150] wl[251] vdd gnd cell_6t
Xbit_r252_c150 bl[150] br[150] wl[252] vdd gnd cell_6t
Xbit_r253_c150 bl[150] br[150] wl[253] vdd gnd cell_6t
Xbit_r254_c150 bl[150] br[150] wl[254] vdd gnd cell_6t
Xbit_r255_c150 bl[150] br[150] wl[255] vdd gnd cell_6t
Xbit_r0_c151 bl[151] br[151] wl[0] vdd gnd cell_6t
Xbit_r1_c151 bl[151] br[151] wl[1] vdd gnd cell_6t
Xbit_r2_c151 bl[151] br[151] wl[2] vdd gnd cell_6t
Xbit_r3_c151 bl[151] br[151] wl[3] vdd gnd cell_6t
Xbit_r4_c151 bl[151] br[151] wl[4] vdd gnd cell_6t
Xbit_r5_c151 bl[151] br[151] wl[5] vdd gnd cell_6t
Xbit_r6_c151 bl[151] br[151] wl[6] vdd gnd cell_6t
Xbit_r7_c151 bl[151] br[151] wl[7] vdd gnd cell_6t
Xbit_r8_c151 bl[151] br[151] wl[8] vdd gnd cell_6t
Xbit_r9_c151 bl[151] br[151] wl[9] vdd gnd cell_6t
Xbit_r10_c151 bl[151] br[151] wl[10] vdd gnd cell_6t
Xbit_r11_c151 bl[151] br[151] wl[11] vdd gnd cell_6t
Xbit_r12_c151 bl[151] br[151] wl[12] vdd gnd cell_6t
Xbit_r13_c151 bl[151] br[151] wl[13] vdd gnd cell_6t
Xbit_r14_c151 bl[151] br[151] wl[14] vdd gnd cell_6t
Xbit_r15_c151 bl[151] br[151] wl[15] vdd gnd cell_6t
Xbit_r16_c151 bl[151] br[151] wl[16] vdd gnd cell_6t
Xbit_r17_c151 bl[151] br[151] wl[17] vdd gnd cell_6t
Xbit_r18_c151 bl[151] br[151] wl[18] vdd gnd cell_6t
Xbit_r19_c151 bl[151] br[151] wl[19] vdd gnd cell_6t
Xbit_r20_c151 bl[151] br[151] wl[20] vdd gnd cell_6t
Xbit_r21_c151 bl[151] br[151] wl[21] vdd gnd cell_6t
Xbit_r22_c151 bl[151] br[151] wl[22] vdd gnd cell_6t
Xbit_r23_c151 bl[151] br[151] wl[23] vdd gnd cell_6t
Xbit_r24_c151 bl[151] br[151] wl[24] vdd gnd cell_6t
Xbit_r25_c151 bl[151] br[151] wl[25] vdd gnd cell_6t
Xbit_r26_c151 bl[151] br[151] wl[26] vdd gnd cell_6t
Xbit_r27_c151 bl[151] br[151] wl[27] vdd gnd cell_6t
Xbit_r28_c151 bl[151] br[151] wl[28] vdd gnd cell_6t
Xbit_r29_c151 bl[151] br[151] wl[29] vdd gnd cell_6t
Xbit_r30_c151 bl[151] br[151] wl[30] vdd gnd cell_6t
Xbit_r31_c151 bl[151] br[151] wl[31] vdd gnd cell_6t
Xbit_r32_c151 bl[151] br[151] wl[32] vdd gnd cell_6t
Xbit_r33_c151 bl[151] br[151] wl[33] vdd gnd cell_6t
Xbit_r34_c151 bl[151] br[151] wl[34] vdd gnd cell_6t
Xbit_r35_c151 bl[151] br[151] wl[35] vdd gnd cell_6t
Xbit_r36_c151 bl[151] br[151] wl[36] vdd gnd cell_6t
Xbit_r37_c151 bl[151] br[151] wl[37] vdd gnd cell_6t
Xbit_r38_c151 bl[151] br[151] wl[38] vdd gnd cell_6t
Xbit_r39_c151 bl[151] br[151] wl[39] vdd gnd cell_6t
Xbit_r40_c151 bl[151] br[151] wl[40] vdd gnd cell_6t
Xbit_r41_c151 bl[151] br[151] wl[41] vdd gnd cell_6t
Xbit_r42_c151 bl[151] br[151] wl[42] vdd gnd cell_6t
Xbit_r43_c151 bl[151] br[151] wl[43] vdd gnd cell_6t
Xbit_r44_c151 bl[151] br[151] wl[44] vdd gnd cell_6t
Xbit_r45_c151 bl[151] br[151] wl[45] vdd gnd cell_6t
Xbit_r46_c151 bl[151] br[151] wl[46] vdd gnd cell_6t
Xbit_r47_c151 bl[151] br[151] wl[47] vdd gnd cell_6t
Xbit_r48_c151 bl[151] br[151] wl[48] vdd gnd cell_6t
Xbit_r49_c151 bl[151] br[151] wl[49] vdd gnd cell_6t
Xbit_r50_c151 bl[151] br[151] wl[50] vdd gnd cell_6t
Xbit_r51_c151 bl[151] br[151] wl[51] vdd gnd cell_6t
Xbit_r52_c151 bl[151] br[151] wl[52] vdd gnd cell_6t
Xbit_r53_c151 bl[151] br[151] wl[53] vdd gnd cell_6t
Xbit_r54_c151 bl[151] br[151] wl[54] vdd gnd cell_6t
Xbit_r55_c151 bl[151] br[151] wl[55] vdd gnd cell_6t
Xbit_r56_c151 bl[151] br[151] wl[56] vdd gnd cell_6t
Xbit_r57_c151 bl[151] br[151] wl[57] vdd gnd cell_6t
Xbit_r58_c151 bl[151] br[151] wl[58] vdd gnd cell_6t
Xbit_r59_c151 bl[151] br[151] wl[59] vdd gnd cell_6t
Xbit_r60_c151 bl[151] br[151] wl[60] vdd gnd cell_6t
Xbit_r61_c151 bl[151] br[151] wl[61] vdd gnd cell_6t
Xbit_r62_c151 bl[151] br[151] wl[62] vdd gnd cell_6t
Xbit_r63_c151 bl[151] br[151] wl[63] vdd gnd cell_6t
Xbit_r64_c151 bl[151] br[151] wl[64] vdd gnd cell_6t
Xbit_r65_c151 bl[151] br[151] wl[65] vdd gnd cell_6t
Xbit_r66_c151 bl[151] br[151] wl[66] vdd gnd cell_6t
Xbit_r67_c151 bl[151] br[151] wl[67] vdd gnd cell_6t
Xbit_r68_c151 bl[151] br[151] wl[68] vdd gnd cell_6t
Xbit_r69_c151 bl[151] br[151] wl[69] vdd gnd cell_6t
Xbit_r70_c151 bl[151] br[151] wl[70] vdd gnd cell_6t
Xbit_r71_c151 bl[151] br[151] wl[71] vdd gnd cell_6t
Xbit_r72_c151 bl[151] br[151] wl[72] vdd gnd cell_6t
Xbit_r73_c151 bl[151] br[151] wl[73] vdd gnd cell_6t
Xbit_r74_c151 bl[151] br[151] wl[74] vdd gnd cell_6t
Xbit_r75_c151 bl[151] br[151] wl[75] vdd gnd cell_6t
Xbit_r76_c151 bl[151] br[151] wl[76] vdd gnd cell_6t
Xbit_r77_c151 bl[151] br[151] wl[77] vdd gnd cell_6t
Xbit_r78_c151 bl[151] br[151] wl[78] vdd gnd cell_6t
Xbit_r79_c151 bl[151] br[151] wl[79] vdd gnd cell_6t
Xbit_r80_c151 bl[151] br[151] wl[80] vdd gnd cell_6t
Xbit_r81_c151 bl[151] br[151] wl[81] vdd gnd cell_6t
Xbit_r82_c151 bl[151] br[151] wl[82] vdd gnd cell_6t
Xbit_r83_c151 bl[151] br[151] wl[83] vdd gnd cell_6t
Xbit_r84_c151 bl[151] br[151] wl[84] vdd gnd cell_6t
Xbit_r85_c151 bl[151] br[151] wl[85] vdd gnd cell_6t
Xbit_r86_c151 bl[151] br[151] wl[86] vdd gnd cell_6t
Xbit_r87_c151 bl[151] br[151] wl[87] vdd gnd cell_6t
Xbit_r88_c151 bl[151] br[151] wl[88] vdd gnd cell_6t
Xbit_r89_c151 bl[151] br[151] wl[89] vdd gnd cell_6t
Xbit_r90_c151 bl[151] br[151] wl[90] vdd gnd cell_6t
Xbit_r91_c151 bl[151] br[151] wl[91] vdd gnd cell_6t
Xbit_r92_c151 bl[151] br[151] wl[92] vdd gnd cell_6t
Xbit_r93_c151 bl[151] br[151] wl[93] vdd gnd cell_6t
Xbit_r94_c151 bl[151] br[151] wl[94] vdd gnd cell_6t
Xbit_r95_c151 bl[151] br[151] wl[95] vdd gnd cell_6t
Xbit_r96_c151 bl[151] br[151] wl[96] vdd gnd cell_6t
Xbit_r97_c151 bl[151] br[151] wl[97] vdd gnd cell_6t
Xbit_r98_c151 bl[151] br[151] wl[98] vdd gnd cell_6t
Xbit_r99_c151 bl[151] br[151] wl[99] vdd gnd cell_6t
Xbit_r100_c151 bl[151] br[151] wl[100] vdd gnd cell_6t
Xbit_r101_c151 bl[151] br[151] wl[101] vdd gnd cell_6t
Xbit_r102_c151 bl[151] br[151] wl[102] vdd gnd cell_6t
Xbit_r103_c151 bl[151] br[151] wl[103] vdd gnd cell_6t
Xbit_r104_c151 bl[151] br[151] wl[104] vdd gnd cell_6t
Xbit_r105_c151 bl[151] br[151] wl[105] vdd gnd cell_6t
Xbit_r106_c151 bl[151] br[151] wl[106] vdd gnd cell_6t
Xbit_r107_c151 bl[151] br[151] wl[107] vdd gnd cell_6t
Xbit_r108_c151 bl[151] br[151] wl[108] vdd gnd cell_6t
Xbit_r109_c151 bl[151] br[151] wl[109] vdd gnd cell_6t
Xbit_r110_c151 bl[151] br[151] wl[110] vdd gnd cell_6t
Xbit_r111_c151 bl[151] br[151] wl[111] vdd gnd cell_6t
Xbit_r112_c151 bl[151] br[151] wl[112] vdd gnd cell_6t
Xbit_r113_c151 bl[151] br[151] wl[113] vdd gnd cell_6t
Xbit_r114_c151 bl[151] br[151] wl[114] vdd gnd cell_6t
Xbit_r115_c151 bl[151] br[151] wl[115] vdd gnd cell_6t
Xbit_r116_c151 bl[151] br[151] wl[116] vdd gnd cell_6t
Xbit_r117_c151 bl[151] br[151] wl[117] vdd gnd cell_6t
Xbit_r118_c151 bl[151] br[151] wl[118] vdd gnd cell_6t
Xbit_r119_c151 bl[151] br[151] wl[119] vdd gnd cell_6t
Xbit_r120_c151 bl[151] br[151] wl[120] vdd gnd cell_6t
Xbit_r121_c151 bl[151] br[151] wl[121] vdd gnd cell_6t
Xbit_r122_c151 bl[151] br[151] wl[122] vdd gnd cell_6t
Xbit_r123_c151 bl[151] br[151] wl[123] vdd gnd cell_6t
Xbit_r124_c151 bl[151] br[151] wl[124] vdd gnd cell_6t
Xbit_r125_c151 bl[151] br[151] wl[125] vdd gnd cell_6t
Xbit_r126_c151 bl[151] br[151] wl[126] vdd gnd cell_6t
Xbit_r127_c151 bl[151] br[151] wl[127] vdd gnd cell_6t
Xbit_r128_c151 bl[151] br[151] wl[128] vdd gnd cell_6t
Xbit_r129_c151 bl[151] br[151] wl[129] vdd gnd cell_6t
Xbit_r130_c151 bl[151] br[151] wl[130] vdd gnd cell_6t
Xbit_r131_c151 bl[151] br[151] wl[131] vdd gnd cell_6t
Xbit_r132_c151 bl[151] br[151] wl[132] vdd gnd cell_6t
Xbit_r133_c151 bl[151] br[151] wl[133] vdd gnd cell_6t
Xbit_r134_c151 bl[151] br[151] wl[134] vdd gnd cell_6t
Xbit_r135_c151 bl[151] br[151] wl[135] vdd gnd cell_6t
Xbit_r136_c151 bl[151] br[151] wl[136] vdd gnd cell_6t
Xbit_r137_c151 bl[151] br[151] wl[137] vdd gnd cell_6t
Xbit_r138_c151 bl[151] br[151] wl[138] vdd gnd cell_6t
Xbit_r139_c151 bl[151] br[151] wl[139] vdd gnd cell_6t
Xbit_r140_c151 bl[151] br[151] wl[140] vdd gnd cell_6t
Xbit_r141_c151 bl[151] br[151] wl[141] vdd gnd cell_6t
Xbit_r142_c151 bl[151] br[151] wl[142] vdd gnd cell_6t
Xbit_r143_c151 bl[151] br[151] wl[143] vdd gnd cell_6t
Xbit_r144_c151 bl[151] br[151] wl[144] vdd gnd cell_6t
Xbit_r145_c151 bl[151] br[151] wl[145] vdd gnd cell_6t
Xbit_r146_c151 bl[151] br[151] wl[146] vdd gnd cell_6t
Xbit_r147_c151 bl[151] br[151] wl[147] vdd gnd cell_6t
Xbit_r148_c151 bl[151] br[151] wl[148] vdd gnd cell_6t
Xbit_r149_c151 bl[151] br[151] wl[149] vdd gnd cell_6t
Xbit_r150_c151 bl[151] br[151] wl[150] vdd gnd cell_6t
Xbit_r151_c151 bl[151] br[151] wl[151] vdd gnd cell_6t
Xbit_r152_c151 bl[151] br[151] wl[152] vdd gnd cell_6t
Xbit_r153_c151 bl[151] br[151] wl[153] vdd gnd cell_6t
Xbit_r154_c151 bl[151] br[151] wl[154] vdd gnd cell_6t
Xbit_r155_c151 bl[151] br[151] wl[155] vdd gnd cell_6t
Xbit_r156_c151 bl[151] br[151] wl[156] vdd gnd cell_6t
Xbit_r157_c151 bl[151] br[151] wl[157] vdd gnd cell_6t
Xbit_r158_c151 bl[151] br[151] wl[158] vdd gnd cell_6t
Xbit_r159_c151 bl[151] br[151] wl[159] vdd gnd cell_6t
Xbit_r160_c151 bl[151] br[151] wl[160] vdd gnd cell_6t
Xbit_r161_c151 bl[151] br[151] wl[161] vdd gnd cell_6t
Xbit_r162_c151 bl[151] br[151] wl[162] vdd gnd cell_6t
Xbit_r163_c151 bl[151] br[151] wl[163] vdd gnd cell_6t
Xbit_r164_c151 bl[151] br[151] wl[164] vdd gnd cell_6t
Xbit_r165_c151 bl[151] br[151] wl[165] vdd gnd cell_6t
Xbit_r166_c151 bl[151] br[151] wl[166] vdd gnd cell_6t
Xbit_r167_c151 bl[151] br[151] wl[167] vdd gnd cell_6t
Xbit_r168_c151 bl[151] br[151] wl[168] vdd gnd cell_6t
Xbit_r169_c151 bl[151] br[151] wl[169] vdd gnd cell_6t
Xbit_r170_c151 bl[151] br[151] wl[170] vdd gnd cell_6t
Xbit_r171_c151 bl[151] br[151] wl[171] vdd gnd cell_6t
Xbit_r172_c151 bl[151] br[151] wl[172] vdd gnd cell_6t
Xbit_r173_c151 bl[151] br[151] wl[173] vdd gnd cell_6t
Xbit_r174_c151 bl[151] br[151] wl[174] vdd gnd cell_6t
Xbit_r175_c151 bl[151] br[151] wl[175] vdd gnd cell_6t
Xbit_r176_c151 bl[151] br[151] wl[176] vdd gnd cell_6t
Xbit_r177_c151 bl[151] br[151] wl[177] vdd gnd cell_6t
Xbit_r178_c151 bl[151] br[151] wl[178] vdd gnd cell_6t
Xbit_r179_c151 bl[151] br[151] wl[179] vdd gnd cell_6t
Xbit_r180_c151 bl[151] br[151] wl[180] vdd gnd cell_6t
Xbit_r181_c151 bl[151] br[151] wl[181] vdd gnd cell_6t
Xbit_r182_c151 bl[151] br[151] wl[182] vdd gnd cell_6t
Xbit_r183_c151 bl[151] br[151] wl[183] vdd gnd cell_6t
Xbit_r184_c151 bl[151] br[151] wl[184] vdd gnd cell_6t
Xbit_r185_c151 bl[151] br[151] wl[185] vdd gnd cell_6t
Xbit_r186_c151 bl[151] br[151] wl[186] vdd gnd cell_6t
Xbit_r187_c151 bl[151] br[151] wl[187] vdd gnd cell_6t
Xbit_r188_c151 bl[151] br[151] wl[188] vdd gnd cell_6t
Xbit_r189_c151 bl[151] br[151] wl[189] vdd gnd cell_6t
Xbit_r190_c151 bl[151] br[151] wl[190] vdd gnd cell_6t
Xbit_r191_c151 bl[151] br[151] wl[191] vdd gnd cell_6t
Xbit_r192_c151 bl[151] br[151] wl[192] vdd gnd cell_6t
Xbit_r193_c151 bl[151] br[151] wl[193] vdd gnd cell_6t
Xbit_r194_c151 bl[151] br[151] wl[194] vdd gnd cell_6t
Xbit_r195_c151 bl[151] br[151] wl[195] vdd gnd cell_6t
Xbit_r196_c151 bl[151] br[151] wl[196] vdd gnd cell_6t
Xbit_r197_c151 bl[151] br[151] wl[197] vdd gnd cell_6t
Xbit_r198_c151 bl[151] br[151] wl[198] vdd gnd cell_6t
Xbit_r199_c151 bl[151] br[151] wl[199] vdd gnd cell_6t
Xbit_r200_c151 bl[151] br[151] wl[200] vdd gnd cell_6t
Xbit_r201_c151 bl[151] br[151] wl[201] vdd gnd cell_6t
Xbit_r202_c151 bl[151] br[151] wl[202] vdd gnd cell_6t
Xbit_r203_c151 bl[151] br[151] wl[203] vdd gnd cell_6t
Xbit_r204_c151 bl[151] br[151] wl[204] vdd gnd cell_6t
Xbit_r205_c151 bl[151] br[151] wl[205] vdd gnd cell_6t
Xbit_r206_c151 bl[151] br[151] wl[206] vdd gnd cell_6t
Xbit_r207_c151 bl[151] br[151] wl[207] vdd gnd cell_6t
Xbit_r208_c151 bl[151] br[151] wl[208] vdd gnd cell_6t
Xbit_r209_c151 bl[151] br[151] wl[209] vdd gnd cell_6t
Xbit_r210_c151 bl[151] br[151] wl[210] vdd gnd cell_6t
Xbit_r211_c151 bl[151] br[151] wl[211] vdd gnd cell_6t
Xbit_r212_c151 bl[151] br[151] wl[212] vdd gnd cell_6t
Xbit_r213_c151 bl[151] br[151] wl[213] vdd gnd cell_6t
Xbit_r214_c151 bl[151] br[151] wl[214] vdd gnd cell_6t
Xbit_r215_c151 bl[151] br[151] wl[215] vdd gnd cell_6t
Xbit_r216_c151 bl[151] br[151] wl[216] vdd gnd cell_6t
Xbit_r217_c151 bl[151] br[151] wl[217] vdd gnd cell_6t
Xbit_r218_c151 bl[151] br[151] wl[218] vdd gnd cell_6t
Xbit_r219_c151 bl[151] br[151] wl[219] vdd gnd cell_6t
Xbit_r220_c151 bl[151] br[151] wl[220] vdd gnd cell_6t
Xbit_r221_c151 bl[151] br[151] wl[221] vdd gnd cell_6t
Xbit_r222_c151 bl[151] br[151] wl[222] vdd gnd cell_6t
Xbit_r223_c151 bl[151] br[151] wl[223] vdd gnd cell_6t
Xbit_r224_c151 bl[151] br[151] wl[224] vdd gnd cell_6t
Xbit_r225_c151 bl[151] br[151] wl[225] vdd gnd cell_6t
Xbit_r226_c151 bl[151] br[151] wl[226] vdd gnd cell_6t
Xbit_r227_c151 bl[151] br[151] wl[227] vdd gnd cell_6t
Xbit_r228_c151 bl[151] br[151] wl[228] vdd gnd cell_6t
Xbit_r229_c151 bl[151] br[151] wl[229] vdd gnd cell_6t
Xbit_r230_c151 bl[151] br[151] wl[230] vdd gnd cell_6t
Xbit_r231_c151 bl[151] br[151] wl[231] vdd gnd cell_6t
Xbit_r232_c151 bl[151] br[151] wl[232] vdd gnd cell_6t
Xbit_r233_c151 bl[151] br[151] wl[233] vdd gnd cell_6t
Xbit_r234_c151 bl[151] br[151] wl[234] vdd gnd cell_6t
Xbit_r235_c151 bl[151] br[151] wl[235] vdd gnd cell_6t
Xbit_r236_c151 bl[151] br[151] wl[236] vdd gnd cell_6t
Xbit_r237_c151 bl[151] br[151] wl[237] vdd gnd cell_6t
Xbit_r238_c151 bl[151] br[151] wl[238] vdd gnd cell_6t
Xbit_r239_c151 bl[151] br[151] wl[239] vdd gnd cell_6t
Xbit_r240_c151 bl[151] br[151] wl[240] vdd gnd cell_6t
Xbit_r241_c151 bl[151] br[151] wl[241] vdd gnd cell_6t
Xbit_r242_c151 bl[151] br[151] wl[242] vdd gnd cell_6t
Xbit_r243_c151 bl[151] br[151] wl[243] vdd gnd cell_6t
Xbit_r244_c151 bl[151] br[151] wl[244] vdd gnd cell_6t
Xbit_r245_c151 bl[151] br[151] wl[245] vdd gnd cell_6t
Xbit_r246_c151 bl[151] br[151] wl[246] vdd gnd cell_6t
Xbit_r247_c151 bl[151] br[151] wl[247] vdd gnd cell_6t
Xbit_r248_c151 bl[151] br[151] wl[248] vdd gnd cell_6t
Xbit_r249_c151 bl[151] br[151] wl[249] vdd gnd cell_6t
Xbit_r250_c151 bl[151] br[151] wl[250] vdd gnd cell_6t
Xbit_r251_c151 bl[151] br[151] wl[251] vdd gnd cell_6t
Xbit_r252_c151 bl[151] br[151] wl[252] vdd gnd cell_6t
Xbit_r253_c151 bl[151] br[151] wl[253] vdd gnd cell_6t
Xbit_r254_c151 bl[151] br[151] wl[254] vdd gnd cell_6t
Xbit_r255_c151 bl[151] br[151] wl[255] vdd gnd cell_6t
Xbit_r0_c152 bl[152] br[152] wl[0] vdd gnd cell_6t
Xbit_r1_c152 bl[152] br[152] wl[1] vdd gnd cell_6t
Xbit_r2_c152 bl[152] br[152] wl[2] vdd gnd cell_6t
Xbit_r3_c152 bl[152] br[152] wl[3] vdd gnd cell_6t
Xbit_r4_c152 bl[152] br[152] wl[4] vdd gnd cell_6t
Xbit_r5_c152 bl[152] br[152] wl[5] vdd gnd cell_6t
Xbit_r6_c152 bl[152] br[152] wl[6] vdd gnd cell_6t
Xbit_r7_c152 bl[152] br[152] wl[7] vdd gnd cell_6t
Xbit_r8_c152 bl[152] br[152] wl[8] vdd gnd cell_6t
Xbit_r9_c152 bl[152] br[152] wl[9] vdd gnd cell_6t
Xbit_r10_c152 bl[152] br[152] wl[10] vdd gnd cell_6t
Xbit_r11_c152 bl[152] br[152] wl[11] vdd gnd cell_6t
Xbit_r12_c152 bl[152] br[152] wl[12] vdd gnd cell_6t
Xbit_r13_c152 bl[152] br[152] wl[13] vdd gnd cell_6t
Xbit_r14_c152 bl[152] br[152] wl[14] vdd gnd cell_6t
Xbit_r15_c152 bl[152] br[152] wl[15] vdd gnd cell_6t
Xbit_r16_c152 bl[152] br[152] wl[16] vdd gnd cell_6t
Xbit_r17_c152 bl[152] br[152] wl[17] vdd gnd cell_6t
Xbit_r18_c152 bl[152] br[152] wl[18] vdd gnd cell_6t
Xbit_r19_c152 bl[152] br[152] wl[19] vdd gnd cell_6t
Xbit_r20_c152 bl[152] br[152] wl[20] vdd gnd cell_6t
Xbit_r21_c152 bl[152] br[152] wl[21] vdd gnd cell_6t
Xbit_r22_c152 bl[152] br[152] wl[22] vdd gnd cell_6t
Xbit_r23_c152 bl[152] br[152] wl[23] vdd gnd cell_6t
Xbit_r24_c152 bl[152] br[152] wl[24] vdd gnd cell_6t
Xbit_r25_c152 bl[152] br[152] wl[25] vdd gnd cell_6t
Xbit_r26_c152 bl[152] br[152] wl[26] vdd gnd cell_6t
Xbit_r27_c152 bl[152] br[152] wl[27] vdd gnd cell_6t
Xbit_r28_c152 bl[152] br[152] wl[28] vdd gnd cell_6t
Xbit_r29_c152 bl[152] br[152] wl[29] vdd gnd cell_6t
Xbit_r30_c152 bl[152] br[152] wl[30] vdd gnd cell_6t
Xbit_r31_c152 bl[152] br[152] wl[31] vdd gnd cell_6t
Xbit_r32_c152 bl[152] br[152] wl[32] vdd gnd cell_6t
Xbit_r33_c152 bl[152] br[152] wl[33] vdd gnd cell_6t
Xbit_r34_c152 bl[152] br[152] wl[34] vdd gnd cell_6t
Xbit_r35_c152 bl[152] br[152] wl[35] vdd gnd cell_6t
Xbit_r36_c152 bl[152] br[152] wl[36] vdd gnd cell_6t
Xbit_r37_c152 bl[152] br[152] wl[37] vdd gnd cell_6t
Xbit_r38_c152 bl[152] br[152] wl[38] vdd gnd cell_6t
Xbit_r39_c152 bl[152] br[152] wl[39] vdd gnd cell_6t
Xbit_r40_c152 bl[152] br[152] wl[40] vdd gnd cell_6t
Xbit_r41_c152 bl[152] br[152] wl[41] vdd gnd cell_6t
Xbit_r42_c152 bl[152] br[152] wl[42] vdd gnd cell_6t
Xbit_r43_c152 bl[152] br[152] wl[43] vdd gnd cell_6t
Xbit_r44_c152 bl[152] br[152] wl[44] vdd gnd cell_6t
Xbit_r45_c152 bl[152] br[152] wl[45] vdd gnd cell_6t
Xbit_r46_c152 bl[152] br[152] wl[46] vdd gnd cell_6t
Xbit_r47_c152 bl[152] br[152] wl[47] vdd gnd cell_6t
Xbit_r48_c152 bl[152] br[152] wl[48] vdd gnd cell_6t
Xbit_r49_c152 bl[152] br[152] wl[49] vdd gnd cell_6t
Xbit_r50_c152 bl[152] br[152] wl[50] vdd gnd cell_6t
Xbit_r51_c152 bl[152] br[152] wl[51] vdd gnd cell_6t
Xbit_r52_c152 bl[152] br[152] wl[52] vdd gnd cell_6t
Xbit_r53_c152 bl[152] br[152] wl[53] vdd gnd cell_6t
Xbit_r54_c152 bl[152] br[152] wl[54] vdd gnd cell_6t
Xbit_r55_c152 bl[152] br[152] wl[55] vdd gnd cell_6t
Xbit_r56_c152 bl[152] br[152] wl[56] vdd gnd cell_6t
Xbit_r57_c152 bl[152] br[152] wl[57] vdd gnd cell_6t
Xbit_r58_c152 bl[152] br[152] wl[58] vdd gnd cell_6t
Xbit_r59_c152 bl[152] br[152] wl[59] vdd gnd cell_6t
Xbit_r60_c152 bl[152] br[152] wl[60] vdd gnd cell_6t
Xbit_r61_c152 bl[152] br[152] wl[61] vdd gnd cell_6t
Xbit_r62_c152 bl[152] br[152] wl[62] vdd gnd cell_6t
Xbit_r63_c152 bl[152] br[152] wl[63] vdd gnd cell_6t
Xbit_r64_c152 bl[152] br[152] wl[64] vdd gnd cell_6t
Xbit_r65_c152 bl[152] br[152] wl[65] vdd gnd cell_6t
Xbit_r66_c152 bl[152] br[152] wl[66] vdd gnd cell_6t
Xbit_r67_c152 bl[152] br[152] wl[67] vdd gnd cell_6t
Xbit_r68_c152 bl[152] br[152] wl[68] vdd gnd cell_6t
Xbit_r69_c152 bl[152] br[152] wl[69] vdd gnd cell_6t
Xbit_r70_c152 bl[152] br[152] wl[70] vdd gnd cell_6t
Xbit_r71_c152 bl[152] br[152] wl[71] vdd gnd cell_6t
Xbit_r72_c152 bl[152] br[152] wl[72] vdd gnd cell_6t
Xbit_r73_c152 bl[152] br[152] wl[73] vdd gnd cell_6t
Xbit_r74_c152 bl[152] br[152] wl[74] vdd gnd cell_6t
Xbit_r75_c152 bl[152] br[152] wl[75] vdd gnd cell_6t
Xbit_r76_c152 bl[152] br[152] wl[76] vdd gnd cell_6t
Xbit_r77_c152 bl[152] br[152] wl[77] vdd gnd cell_6t
Xbit_r78_c152 bl[152] br[152] wl[78] vdd gnd cell_6t
Xbit_r79_c152 bl[152] br[152] wl[79] vdd gnd cell_6t
Xbit_r80_c152 bl[152] br[152] wl[80] vdd gnd cell_6t
Xbit_r81_c152 bl[152] br[152] wl[81] vdd gnd cell_6t
Xbit_r82_c152 bl[152] br[152] wl[82] vdd gnd cell_6t
Xbit_r83_c152 bl[152] br[152] wl[83] vdd gnd cell_6t
Xbit_r84_c152 bl[152] br[152] wl[84] vdd gnd cell_6t
Xbit_r85_c152 bl[152] br[152] wl[85] vdd gnd cell_6t
Xbit_r86_c152 bl[152] br[152] wl[86] vdd gnd cell_6t
Xbit_r87_c152 bl[152] br[152] wl[87] vdd gnd cell_6t
Xbit_r88_c152 bl[152] br[152] wl[88] vdd gnd cell_6t
Xbit_r89_c152 bl[152] br[152] wl[89] vdd gnd cell_6t
Xbit_r90_c152 bl[152] br[152] wl[90] vdd gnd cell_6t
Xbit_r91_c152 bl[152] br[152] wl[91] vdd gnd cell_6t
Xbit_r92_c152 bl[152] br[152] wl[92] vdd gnd cell_6t
Xbit_r93_c152 bl[152] br[152] wl[93] vdd gnd cell_6t
Xbit_r94_c152 bl[152] br[152] wl[94] vdd gnd cell_6t
Xbit_r95_c152 bl[152] br[152] wl[95] vdd gnd cell_6t
Xbit_r96_c152 bl[152] br[152] wl[96] vdd gnd cell_6t
Xbit_r97_c152 bl[152] br[152] wl[97] vdd gnd cell_6t
Xbit_r98_c152 bl[152] br[152] wl[98] vdd gnd cell_6t
Xbit_r99_c152 bl[152] br[152] wl[99] vdd gnd cell_6t
Xbit_r100_c152 bl[152] br[152] wl[100] vdd gnd cell_6t
Xbit_r101_c152 bl[152] br[152] wl[101] vdd gnd cell_6t
Xbit_r102_c152 bl[152] br[152] wl[102] vdd gnd cell_6t
Xbit_r103_c152 bl[152] br[152] wl[103] vdd gnd cell_6t
Xbit_r104_c152 bl[152] br[152] wl[104] vdd gnd cell_6t
Xbit_r105_c152 bl[152] br[152] wl[105] vdd gnd cell_6t
Xbit_r106_c152 bl[152] br[152] wl[106] vdd gnd cell_6t
Xbit_r107_c152 bl[152] br[152] wl[107] vdd gnd cell_6t
Xbit_r108_c152 bl[152] br[152] wl[108] vdd gnd cell_6t
Xbit_r109_c152 bl[152] br[152] wl[109] vdd gnd cell_6t
Xbit_r110_c152 bl[152] br[152] wl[110] vdd gnd cell_6t
Xbit_r111_c152 bl[152] br[152] wl[111] vdd gnd cell_6t
Xbit_r112_c152 bl[152] br[152] wl[112] vdd gnd cell_6t
Xbit_r113_c152 bl[152] br[152] wl[113] vdd gnd cell_6t
Xbit_r114_c152 bl[152] br[152] wl[114] vdd gnd cell_6t
Xbit_r115_c152 bl[152] br[152] wl[115] vdd gnd cell_6t
Xbit_r116_c152 bl[152] br[152] wl[116] vdd gnd cell_6t
Xbit_r117_c152 bl[152] br[152] wl[117] vdd gnd cell_6t
Xbit_r118_c152 bl[152] br[152] wl[118] vdd gnd cell_6t
Xbit_r119_c152 bl[152] br[152] wl[119] vdd gnd cell_6t
Xbit_r120_c152 bl[152] br[152] wl[120] vdd gnd cell_6t
Xbit_r121_c152 bl[152] br[152] wl[121] vdd gnd cell_6t
Xbit_r122_c152 bl[152] br[152] wl[122] vdd gnd cell_6t
Xbit_r123_c152 bl[152] br[152] wl[123] vdd gnd cell_6t
Xbit_r124_c152 bl[152] br[152] wl[124] vdd gnd cell_6t
Xbit_r125_c152 bl[152] br[152] wl[125] vdd gnd cell_6t
Xbit_r126_c152 bl[152] br[152] wl[126] vdd gnd cell_6t
Xbit_r127_c152 bl[152] br[152] wl[127] vdd gnd cell_6t
Xbit_r128_c152 bl[152] br[152] wl[128] vdd gnd cell_6t
Xbit_r129_c152 bl[152] br[152] wl[129] vdd gnd cell_6t
Xbit_r130_c152 bl[152] br[152] wl[130] vdd gnd cell_6t
Xbit_r131_c152 bl[152] br[152] wl[131] vdd gnd cell_6t
Xbit_r132_c152 bl[152] br[152] wl[132] vdd gnd cell_6t
Xbit_r133_c152 bl[152] br[152] wl[133] vdd gnd cell_6t
Xbit_r134_c152 bl[152] br[152] wl[134] vdd gnd cell_6t
Xbit_r135_c152 bl[152] br[152] wl[135] vdd gnd cell_6t
Xbit_r136_c152 bl[152] br[152] wl[136] vdd gnd cell_6t
Xbit_r137_c152 bl[152] br[152] wl[137] vdd gnd cell_6t
Xbit_r138_c152 bl[152] br[152] wl[138] vdd gnd cell_6t
Xbit_r139_c152 bl[152] br[152] wl[139] vdd gnd cell_6t
Xbit_r140_c152 bl[152] br[152] wl[140] vdd gnd cell_6t
Xbit_r141_c152 bl[152] br[152] wl[141] vdd gnd cell_6t
Xbit_r142_c152 bl[152] br[152] wl[142] vdd gnd cell_6t
Xbit_r143_c152 bl[152] br[152] wl[143] vdd gnd cell_6t
Xbit_r144_c152 bl[152] br[152] wl[144] vdd gnd cell_6t
Xbit_r145_c152 bl[152] br[152] wl[145] vdd gnd cell_6t
Xbit_r146_c152 bl[152] br[152] wl[146] vdd gnd cell_6t
Xbit_r147_c152 bl[152] br[152] wl[147] vdd gnd cell_6t
Xbit_r148_c152 bl[152] br[152] wl[148] vdd gnd cell_6t
Xbit_r149_c152 bl[152] br[152] wl[149] vdd gnd cell_6t
Xbit_r150_c152 bl[152] br[152] wl[150] vdd gnd cell_6t
Xbit_r151_c152 bl[152] br[152] wl[151] vdd gnd cell_6t
Xbit_r152_c152 bl[152] br[152] wl[152] vdd gnd cell_6t
Xbit_r153_c152 bl[152] br[152] wl[153] vdd gnd cell_6t
Xbit_r154_c152 bl[152] br[152] wl[154] vdd gnd cell_6t
Xbit_r155_c152 bl[152] br[152] wl[155] vdd gnd cell_6t
Xbit_r156_c152 bl[152] br[152] wl[156] vdd gnd cell_6t
Xbit_r157_c152 bl[152] br[152] wl[157] vdd gnd cell_6t
Xbit_r158_c152 bl[152] br[152] wl[158] vdd gnd cell_6t
Xbit_r159_c152 bl[152] br[152] wl[159] vdd gnd cell_6t
Xbit_r160_c152 bl[152] br[152] wl[160] vdd gnd cell_6t
Xbit_r161_c152 bl[152] br[152] wl[161] vdd gnd cell_6t
Xbit_r162_c152 bl[152] br[152] wl[162] vdd gnd cell_6t
Xbit_r163_c152 bl[152] br[152] wl[163] vdd gnd cell_6t
Xbit_r164_c152 bl[152] br[152] wl[164] vdd gnd cell_6t
Xbit_r165_c152 bl[152] br[152] wl[165] vdd gnd cell_6t
Xbit_r166_c152 bl[152] br[152] wl[166] vdd gnd cell_6t
Xbit_r167_c152 bl[152] br[152] wl[167] vdd gnd cell_6t
Xbit_r168_c152 bl[152] br[152] wl[168] vdd gnd cell_6t
Xbit_r169_c152 bl[152] br[152] wl[169] vdd gnd cell_6t
Xbit_r170_c152 bl[152] br[152] wl[170] vdd gnd cell_6t
Xbit_r171_c152 bl[152] br[152] wl[171] vdd gnd cell_6t
Xbit_r172_c152 bl[152] br[152] wl[172] vdd gnd cell_6t
Xbit_r173_c152 bl[152] br[152] wl[173] vdd gnd cell_6t
Xbit_r174_c152 bl[152] br[152] wl[174] vdd gnd cell_6t
Xbit_r175_c152 bl[152] br[152] wl[175] vdd gnd cell_6t
Xbit_r176_c152 bl[152] br[152] wl[176] vdd gnd cell_6t
Xbit_r177_c152 bl[152] br[152] wl[177] vdd gnd cell_6t
Xbit_r178_c152 bl[152] br[152] wl[178] vdd gnd cell_6t
Xbit_r179_c152 bl[152] br[152] wl[179] vdd gnd cell_6t
Xbit_r180_c152 bl[152] br[152] wl[180] vdd gnd cell_6t
Xbit_r181_c152 bl[152] br[152] wl[181] vdd gnd cell_6t
Xbit_r182_c152 bl[152] br[152] wl[182] vdd gnd cell_6t
Xbit_r183_c152 bl[152] br[152] wl[183] vdd gnd cell_6t
Xbit_r184_c152 bl[152] br[152] wl[184] vdd gnd cell_6t
Xbit_r185_c152 bl[152] br[152] wl[185] vdd gnd cell_6t
Xbit_r186_c152 bl[152] br[152] wl[186] vdd gnd cell_6t
Xbit_r187_c152 bl[152] br[152] wl[187] vdd gnd cell_6t
Xbit_r188_c152 bl[152] br[152] wl[188] vdd gnd cell_6t
Xbit_r189_c152 bl[152] br[152] wl[189] vdd gnd cell_6t
Xbit_r190_c152 bl[152] br[152] wl[190] vdd gnd cell_6t
Xbit_r191_c152 bl[152] br[152] wl[191] vdd gnd cell_6t
Xbit_r192_c152 bl[152] br[152] wl[192] vdd gnd cell_6t
Xbit_r193_c152 bl[152] br[152] wl[193] vdd gnd cell_6t
Xbit_r194_c152 bl[152] br[152] wl[194] vdd gnd cell_6t
Xbit_r195_c152 bl[152] br[152] wl[195] vdd gnd cell_6t
Xbit_r196_c152 bl[152] br[152] wl[196] vdd gnd cell_6t
Xbit_r197_c152 bl[152] br[152] wl[197] vdd gnd cell_6t
Xbit_r198_c152 bl[152] br[152] wl[198] vdd gnd cell_6t
Xbit_r199_c152 bl[152] br[152] wl[199] vdd gnd cell_6t
Xbit_r200_c152 bl[152] br[152] wl[200] vdd gnd cell_6t
Xbit_r201_c152 bl[152] br[152] wl[201] vdd gnd cell_6t
Xbit_r202_c152 bl[152] br[152] wl[202] vdd gnd cell_6t
Xbit_r203_c152 bl[152] br[152] wl[203] vdd gnd cell_6t
Xbit_r204_c152 bl[152] br[152] wl[204] vdd gnd cell_6t
Xbit_r205_c152 bl[152] br[152] wl[205] vdd gnd cell_6t
Xbit_r206_c152 bl[152] br[152] wl[206] vdd gnd cell_6t
Xbit_r207_c152 bl[152] br[152] wl[207] vdd gnd cell_6t
Xbit_r208_c152 bl[152] br[152] wl[208] vdd gnd cell_6t
Xbit_r209_c152 bl[152] br[152] wl[209] vdd gnd cell_6t
Xbit_r210_c152 bl[152] br[152] wl[210] vdd gnd cell_6t
Xbit_r211_c152 bl[152] br[152] wl[211] vdd gnd cell_6t
Xbit_r212_c152 bl[152] br[152] wl[212] vdd gnd cell_6t
Xbit_r213_c152 bl[152] br[152] wl[213] vdd gnd cell_6t
Xbit_r214_c152 bl[152] br[152] wl[214] vdd gnd cell_6t
Xbit_r215_c152 bl[152] br[152] wl[215] vdd gnd cell_6t
Xbit_r216_c152 bl[152] br[152] wl[216] vdd gnd cell_6t
Xbit_r217_c152 bl[152] br[152] wl[217] vdd gnd cell_6t
Xbit_r218_c152 bl[152] br[152] wl[218] vdd gnd cell_6t
Xbit_r219_c152 bl[152] br[152] wl[219] vdd gnd cell_6t
Xbit_r220_c152 bl[152] br[152] wl[220] vdd gnd cell_6t
Xbit_r221_c152 bl[152] br[152] wl[221] vdd gnd cell_6t
Xbit_r222_c152 bl[152] br[152] wl[222] vdd gnd cell_6t
Xbit_r223_c152 bl[152] br[152] wl[223] vdd gnd cell_6t
Xbit_r224_c152 bl[152] br[152] wl[224] vdd gnd cell_6t
Xbit_r225_c152 bl[152] br[152] wl[225] vdd gnd cell_6t
Xbit_r226_c152 bl[152] br[152] wl[226] vdd gnd cell_6t
Xbit_r227_c152 bl[152] br[152] wl[227] vdd gnd cell_6t
Xbit_r228_c152 bl[152] br[152] wl[228] vdd gnd cell_6t
Xbit_r229_c152 bl[152] br[152] wl[229] vdd gnd cell_6t
Xbit_r230_c152 bl[152] br[152] wl[230] vdd gnd cell_6t
Xbit_r231_c152 bl[152] br[152] wl[231] vdd gnd cell_6t
Xbit_r232_c152 bl[152] br[152] wl[232] vdd gnd cell_6t
Xbit_r233_c152 bl[152] br[152] wl[233] vdd gnd cell_6t
Xbit_r234_c152 bl[152] br[152] wl[234] vdd gnd cell_6t
Xbit_r235_c152 bl[152] br[152] wl[235] vdd gnd cell_6t
Xbit_r236_c152 bl[152] br[152] wl[236] vdd gnd cell_6t
Xbit_r237_c152 bl[152] br[152] wl[237] vdd gnd cell_6t
Xbit_r238_c152 bl[152] br[152] wl[238] vdd gnd cell_6t
Xbit_r239_c152 bl[152] br[152] wl[239] vdd gnd cell_6t
Xbit_r240_c152 bl[152] br[152] wl[240] vdd gnd cell_6t
Xbit_r241_c152 bl[152] br[152] wl[241] vdd gnd cell_6t
Xbit_r242_c152 bl[152] br[152] wl[242] vdd gnd cell_6t
Xbit_r243_c152 bl[152] br[152] wl[243] vdd gnd cell_6t
Xbit_r244_c152 bl[152] br[152] wl[244] vdd gnd cell_6t
Xbit_r245_c152 bl[152] br[152] wl[245] vdd gnd cell_6t
Xbit_r246_c152 bl[152] br[152] wl[246] vdd gnd cell_6t
Xbit_r247_c152 bl[152] br[152] wl[247] vdd gnd cell_6t
Xbit_r248_c152 bl[152] br[152] wl[248] vdd gnd cell_6t
Xbit_r249_c152 bl[152] br[152] wl[249] vdd gnd cell_6t
Xbit_r250_c152 bl[152] br[152] wl[250] vdd gnd cell_6t
Xbit_r251_c152 bl[152] br[152] wl[251] vdd gnd cell_6t
Xbit_r252_c152 bl[152] br[152] wl[252] vdd gnd cell_6t
Xbit_r253_c152 bl[152] br[152] wl[253] vdd gnd cell_6t
Xbit_r254_c152 bl[152] br[152] wl[254] vdd gnd cell_6t
Xbit_r255_c152 bl[152] br[152] wl[255] vdd gnd cell_6t
Xbit_r0_c153 bl[153] br[153] wl[0] vdd gnd cell_6t
Xbit_r1_c153 bl[153] br[153] wl[1] vdd gnd cell_6t
Xbit_r2_c153 bl[153] br[153] wl[2] vdd gnd cell_6t
Xbit_r3_c153 bl[153] br[153] wl[3] vdd gnd cell_6t
Xbit_r4_c153 bl[153] br[153] wl[4] vdd gnd cell_6t
Xbit_r5_c153 bl[153] br[153] wl[5] vdd gnd cell_6t
Xbit_r6_c153 bl[153] br[153] wl[6] vdd gnd cell_6t
Xbit_r7_c153 bl[153] br[153] wl[7] vdd gnd cell_6t
Xbit_r8_c153 bl[153] br[153] wl[8] vdd gnd cell_6t
Xbit_r9_c153 bl[153] br[153] wl[9] vdd gnd cell_6t
Xbit_r10_c153 bl[153] br[153] wl[10] vdd gnd cell_6t
Xbit_r11_c153 bl[153] br[153] wl[11] vdd gnd cell_6t
Xbit_r12_c153 bl[153] br[153] wl[12] vdd gnd cell_6t
Xbit_r13_c153 bl[153] br[153] wl[13] vdd gnd cell_6t
Xbit_r14_c153 bl[153] br[153] wl[14] vdd gnd cell_6t
Xbit_r15_c153 bl[153] br[153] wl[15] vdd gnd cell_6t
Xbit_r16_c153 bl[153] br[153] wl[16] vdd gnd cell_6t
Xbit_r17_c153 bl[153] br[153] wl[17] vdd gnd cell_6t
Xbit_r18_c153 bl[153] br[153] wl[18] vdd gnd cell_6t
Xbit_r19_c153 bl[153] br[153] wl[19] vdd gnd cell_6t
Xbit_r20_c153 bl[153] br[153] wl[20] vdd gnd cell_6t
Xbit_r21_c153 bl[153] br[153] wl[21] vdd gnd cell_6t
Xbit_r22_c153 bl[153] br[153] wl[22] vdd gnd cell_6t
Xbit_r23_c153 bl[153] br[153] wl[23] vdd gnd cell_6t
Xbit_r24_c153 bl[153] br[153] wl[24] vdd gnd cell_6t
Xbit_r25_c153 bl[153] br[153] wl[25] vdd gnd cell_6t
Xbit_r26_c153 bl[153] br[153] wl[26] vdd gnd cell_6t
Xbit_r27_c153 bl[153] br[153] wl[27] vdd gnd cell_6t
Xbit_r28_c153 bl[153] br[153] wl[28] vdd gnd cell_6t
Xbit_r29_c153 bl[153] br[153] wl[29] vdd gnd cell_6t
Xbit_r30_c153 bl[153] br[153] wl[30] vdd gnd cell_6t
Xbit_r31_c153 bl[153] br[153] wl[31] vdd gnd cell_6t
Xbit_r32_c153 bl[153] br[153] wl[32] vdd gnd cell_6t
Xbit_r33_c153 bl[153] br[153] wl[33] vdd gnd cell_6t
Xbit_r34_c153 bl[153] br[153] wl[34] vdd gnd cell_6t
Xbit_r35_c153 bl[153] br[153] wl[35] vdd gnd cell_6t
Xbit_r36_c153 bl[153] br[153] wl[36] vdd gnd cell_6t
Xbit_r37_c153 bl[153] br[153] wl[37] vdd gnd cell_6t
Xbit_r38_c153 bl[153] br[153] wl[38] vdd gnd cell_6t
Xbit_r39_c153 bl[153] br[153] wl[39] vdd gnd cell_6t
Xbit_r40_c153 bl[153] br[153] wl[40] vdd gnd cell_6t
Xbit_r41_c153 bl[153] br[153] wl[41] vdd gnd cell_6t
Xbit_r42_c153 bl[153] br[153] wl[42] vdd gnd cell_6t
Xbit_r43_c153 bl[153] br[153] wl[43] vdd gnd cell_6t
Xbit_r44_c153 bl[153] br[153] wl[44] vdd gnd cell_6t
Xbit_r45_c153 bl[153] br[153] wl[45] vdd gnd cell_6t
Xbit_r46_c153 bl[153] br[153] wl[46] vdd gnd cell_6t
Xbit_r47_c153 bl[153] br[153] wl[47] vdd gnd cell_6t
Xbit_r48_c153 bl[153] br[153] wl[48] vdd gnd cell_6t
Xbit_r49_c153 bl[153] br[153] wl[49] vdd gnd cell_6t
Xbit_r50_c153 bl[153] br[153] wl[50] vdd gnd cell_6t
Xbit_r51_c153 bl[153] br[153] wl[51] vdd gnd cell_6t
Xbit_r52_c153 bl[153] br[153] wl[52] vdd gnd cell_6t
Xbit_r53_c153 bl[153] br[153] wl[53] vdd gnd cell_6t
Xbit_r54_c153 bl[153] br[153] wl[54] vdd gnd cell_6t
Xbit_r55_c153 bl[153] br[153] wl[55] vdd gnd cell_6t
Xbit_r56_c153 bl[153] br[153] wl[56] vdd gnd cell_6t
Xbit_r57_c153 bl[153] br[153] wl[57] vdd gnd cell_6t
Xbit_r58_c153 bl[153] br[153] wl[58] vdd gnd cell_6t
Xbit_r59_c153 bl[153] br[153] wl[59] vdd gnd cell_6t
Xbit_r60_c153 bl[153] br[153] wl[60] vdd gnd cell_6t
Xbit_r61_c153 bl[153] br[153] wl[61] vdd gnd cell_6t
Xbit_r62_c153 bl[153] br[153] wl[62] vdd gnd cell_6t
Xbit_r63_c153 bl[153] br[153] wl[63] vdd gnd cell_6t
Xbit_r64_c153 bl[153] br[153] wl[64] vdd gnd cell_6t
Xbit_r65_c153 bl[153] br[153] wl[65] vdd gnd cell_6t
Xbit_r66_c153 bl[153] br[153] wl[66] vdd gnd cell_6t
Xbit_r67_c153 bl[153] br[153] wl[67] vdd gnd cell_6t
Xbit_r68_c153 bl[153] br[153] wl[68] vdd gnd cell_6t
Xbit_r69_c153 bl[153] br[153] wl[69] vdd gnd cell_6t
Xbit_r70_c153 bl[153] br[153] wl[70] vdd gnd cell_6t
Xbit_r71_c153 bl[153] br[153] wl[71] vdd gnd cell_6t
Xbit_r72_c153 bl[153] br[153] wl[72] vdd gnd cell_6t
Xbit_r73_c153 bl[153] br[153] wl[73] vdd gnd cell_6t
Xbit_r74_c153 bl[153] br[153] wl[74] vdd gnd cell_6t
Xbit_r75_c153 bl[153] br[153] wl[75] vdd gnd cell_6t
Xbit_r76_c153 bl[153] br[153] wl[76] vdd gnd cell_6t
Xbit_r77_c153 bl[153] br[153] wl[77] vdd gnd cell_6t
Xbit_r78_c153 bl[153] br[153] wl[78] vdd gnd cell_6t
Xbit_r79_c153 bl[153] br[153] wl[79] vdd gnd cell_6t
Xbit_r80_c153 bl[153] br[153] wl[80] vdd gnd cell_6t
Xbit_r81_c153 bl[153] br[153] wl[81] vdd gnd cell_6t
Xbit_r82_c153 bl[153] br[153] wl[82] vdd gnd cell_6t
Xbit_r83_c153 bl[153] br[153] wl[83] vdd gnd cell_6t
Xbit_r84_c153 bl[153] br[153] wl[84] vdd gnd cell_6t
Xbit_r85_c153 bl[153] br[153] wl[85] vdd gnd cell_6t
Xbit_r86_c153 bl[153] br[153] wl[86] vdd gnd cell_6t
Xbit_r87_c153 bl[153] br[153] wl[87] vdd gnd cell_6t
Xbit_r88_c153 bl[153] br[153] wl[88] vdd gnd cell_6t
Xbit_r89_c153 bl[153] br[153] wl[89] vdd gnd cell_6t
Xbit_r90_c153 bl[153] br[153] wl[90] vdd gnd cell_6t
Xbit_r91_c153 bl[153] br[153] wl[91] vdd gnd cell_6t
Xbit_r92_c153 bl[153] br[153] wl[92] vdd gnd cell_6t
Xbit_r93_c153 bl[153] br[153] wl[93] vdd gnd cell_6t
Xbit_r94_c153 bl[153] br[153] wl[94] vdd gnd cell_6t
Xbit_r95_c153 bl[153] br[153] wl[95] vdd gnd cell_6t
Xbit_r96_c153 bl[153] br[153] wl[96] vdd gnd cell_6t
Xbit_r97_c153 bl[153] br[153] wl[97] vdd gnd cell_6t
Xbit_r98_c153 bl[153] br[153] wl[98] vdd gnd cell_6t
Xbit_r99_c153 bl[153] br[153] wl[99] vdd gnd cell_6t
Xbit_r100_c153 bl[153] br[153] wl[100] vdd gnd cell_6t
Xbit_r101_c153 bl[153] br[153] wl[101] vdd gnd cell_6t
Xbit_r102_c153 bl[153] br[153] wl[102] vdd gnd cell_6t
Xbit_r103_c153 bl[153] br[153] wl[103] vdd gnd cell_6t
Xbit_r104_c153 bl[153] br[153] wl[104] vdd gnd cell_6t
Xbit_r105_c153 bl[153] br[153] wl[105] vdd gnd cell_6t
Xbit_r106_c153 bl[153] br[153] wl[106] vdd gnd cell_6t
Xbit_r107_c153 bl[153] br[153] wl[107] vdd gnd cell_6t
Xbit_r108_c153 bl[153] br[153] wl[108] vdd gnd cell_6t
Xbit_r109_c153 bl[153] br[153] wl[109] vdd gnd cell_6t
Xbit_r110_c153 bl[153] br[153] wl[110] vdd gnd cell_6t
Xbit_r111_c153 bl[153] br[153] wl[111] vdd gnd cell_6t
Xbit_r112_c153 bl[153] br[153] wl[112] vdd gnd cell_6t
Xbit_r113_c153 bl[153] br[153] wl[113] vdd gnd cell_6t
Xbit_r114_c153 bl[153] br[153] wl[114] vdd gnd cell_6t
Xbit_r115_c153 bl[153] br[153] wl[115] vdd gnd cell_6t
Xbit_r116_c153 bl[153] br[153] wl[116] vdd gnd cell_6t
Xbit_r117_c153 bl[153] br[153] wl[117] vdd gnd cell_6t
Xbit_r118_c153 bl[153] br[153] wl[118] vdd gnd cell_6t
Xbit_r119_c153 bl[153] br[153] wl[119] vdd gnd cell_6t
Xbit_r120_c153 bl[153] br[153] wl[120] vdd gnd cell_6t
Xbit_r121_c153 bl[153] br[153] wl[121] vdd gnd cell_6t
Xbit_r122_c153 bl[153] br[153] wl[122] vdd gnd cell_6t
Xbit_r123_c153 bl[153] br[153] wl[123] vdd gnd cell_6t
Xbit_r124_c153 bl[153] br[153] wl[124] vdd gnd cell_6t
Xbit_r125_c153 bl[153] br[153] wl[125] vdd gnd cell_6t
Xbit_r126_c153 bl[153] br[153] wl[126] vdd gnd cell_6t
Xbit_r127_c153 bl[153] br[153] wl[127] vdd gnd cell_6t
Xbit_r128_c153 bl[153] br[153] wl[128] vdd gnd cell_6t
Xbit_r129_c153 bl[153] br[153] wl[129] vdd gnd cell_6t
Xbit_r130_c153 bl[153] br[153] wl[130] vdd gnd cell_6t
Xbit_r131_c153 bl[153] br[153] wl[131] vdd gnd cell_6t
Xbit_r132_c153 bl[153] br[153] wl[132] vdd gnd cell_6t
Xbit_r133_c153 bl[153] br[153] wl[133] vdd gnd cell_6t
Xbit_r134_c153 bl[153] br[153] wl[134] vdd gnd cell_6t
Xbit_r135_c153 bl[153] br[153] wl[135] vdd gnd cell_6t
Xbit_r136_c153 bl[153] br[153] wl[136] vdd gnd cell_6t
Xbit_r137_c153 bl[153] br[153] wl[137] vdd gnd cell_6t
Xbit_r138_c153 bl[153] br[153] wl[138] vdd gnd cell_6t
Xbit_r139_c153 bl[153] br[153] wl[139] vdd gnd cell_6t
Xbit_r140_c153 bl[153] br[153] wl[140] vdd gnd cell_6t
Xbit_r141_c153 bl[153] br[153] wl[141] vdd gnd cell_6t
Xbit_r142_c153 bl[153] br[153] wl[142] vdd gnd cell_6t
Xbit_r143_c153 bl[153] br[153] wl[143] vdd gnd cell_6t
Xbit_r144_c153 bl[153] br[153] wl[144] vdd gnd cell_6t
Xbit_r145_c153 bl[153] br[153] wl[145] vdd gnd cell_6t
Xbit_r146_c153 bl[153] br[153] wl[146] vdd gnd cell_6t
Xbit_r147_c153 bl[153] br[153] wl[147] vdd gnd cell_6t
Xbit_r148_c153 bl[153] br[153] wl[148] vdd gnd cell_6t
Xbit_r149_c153 bl[153] br[153] wl[149] vdd gnd cell_6t
Xbit_r150_c153 bl[153] br[153] wl[150] vdd gnd cell_6t
Xbit_r151_c153 bl[153] br[153] wl[151] vdd gnd cell_6t
Xbit_r152_c153 bl[153] br[153] wl[152] vdd gnd cell_6t
Xbit_r153_c153 bl[153] br[153] wl[153] vdd gnd cell_6t
Xbit_r154_c153 bl[153] br[153] wl[154] vdd gnd cell_6t
Xbit_r155_c153 bl[153] br[153] wl[155] vdd gnd cell_6t
Xbit_r156_c153 bl[153] br[153] wl[156] vdd gnd cell_6t
Xbit_r157_c153 bl[153] br[153] wl[157] vdd gnd cell_6t
Xbit_r158_c153 bl[153] br[153] wl[158] vdd gnd cell_6t
Xbit_r159_c153 bl[153] br[153] wl[159] vdd gnd cell_6t
Xbit_r160_c153 bl[153] br[153] wl[160] vdd gnd cell_6t
Xbit_r161_c153 bl[153] br[153] wl[161] vdd gnd cell_6t
Xbit_r162_c153 bl[153] br[153] wl[162] vdd gnd cell_6t
Xbit_r163_c153 bl[153] br[153] wl[163] vdd gnd cell_6t
Xbit_r164_c153 bl[153] br[153] wl[164] vdd gnd cell_6t
Xbit_r165_c153 bl[153] br[153] wl[165] vdd gnd cell_6t
Xbit_r166_c153 bl[153] br[153] wl[166] vdd gnd cell_6t
Xbit_r167_c153 bl[153] br[153] wl[167] vdd gnd cell_6t
Xbit_r168_c153 bl[153] br[153] wl[168] vdd gnd cell_6t
Xbit_r169_c153 bl[153] br[153] wl[169] vdd gnd cell_6t
Xbit_r170_c153 bl[153] br[153] wl[170] vdd gnd cell_6t
Xbit_r171_c153 bl[153] br[153] wl[171] vdd gnd cell_6t
Xbit_r172_c153 bl[153] br[153] wl[172] vdd gnd cell_6t
Xbit_r173_c153 bl[153] br[153] wl[173] vdd gnd cell_6t
Xbit_r174_c153 bl[153] br[153] wl[174] vdd gnd cell_6t
Xbit_r175_c153 bl[153] br[153] wl[175] vdd gnd cell_6t
Xbit_r176_c153 bl[153] br[153] wl[176] vdd gnd cell_6t
Xbit_r177_c153 bl[153] br[153] wl[177] vdd gnd cell_6t
Xbit_r178_c153 bl[153] br[153] wl[178] vdd gnd cell_6t
Xbit_r179_c153 bl[153] br[153] wl[179] vdd gnd cell_6t
Xbit_r180_c153 bl[153] br[153] wl[180] vdd gnd cell_6t
Xbit_r181_c153 bl[153] br[153] wl[181] vdd gnd cell_6t
Xbit_r182_c153 bl[153] br[153] wl[182] vdd gnd cell_6t
Xbit_r183_c153 bl[153] br[153] wl[183] vdd gnd cell_6t
Xbit_r184_c153 bl[153] br[153] wl[184] vdd gnd cell_6t
Xbit_r185_c153 bl[153] br[153] wl[185] vdd gnd cell_6t
Xbit_r186_c153 bl[153] br[153] wl[186] vdd gnd cell_6t
Xbit_r187_c153 bl[153] br[153] wl[187] vdd gnd cell_6t
Xbit_r188_c153 bl[153] br[153] wl[188] vdd gnd cell_6t
Xbit_r189_c153 bl[153] br[153] wl[189] vdd gnd cell_6t
Xbit_r190_c153 bl[153] br[153] wl[190] vdd gnd cell_6t
Xbit_r191_c153 bl[153] br[153] wl[191] vdd gnd cell_6t
Xbit_r192_c153 bl[153] br[153] wl[192] vdd gnd cell_6t
Xbit_r193_c153 bl[153] br[153] wl[193] vdd gnd cell_6t
Xbit_r194_c153 bl[153] br[153] wl[194] vdd gnd cell_6t
Xbit_r195_c153 bl[153] br[153] wl[195] vdd gnd cell_6t
Xbit_r196_c153 bl[153] br[153] wl[196] vdd gnd cell_6t
Xbit_r197_c153 bl[153] br[153] wl[197] vdd gnd cell_6t
Xbit_r198_c153 bl[153] br[153] wl[198] vdd gnd cell_6t
Xbit_r199_c153 bl[153] br[153] wl[199] vdd gnd cell_6t
Xbit_r200_c153 bl[153] br[153] wl[200] vdd gnd cell_6t
Xbit_r201_c153 bl[153] br[153] wl[201] vdd gnd cell_6t
Xbit_r202_c153 bl[153] br[153] wl[202] vdd gnd cell_6t
Xbit_r203_c153 bl[153] br[153] wl[203] vdd gnd cell_6t
Xbit_r204_c153 bl[153] br[153] wl[204] vdd gnd cell_6t
Xbit_r205_c153 bl[153] br[153] wl[205] vdd gnd cell_6t
Xbit_r206_c153 bl[153] br[153] wl[206] vdd gnd cell_6t
Xbit_r207_c153 bl[153] br[153] wl[207] vdd gnd cell_6t
Xbit_r208_c153 bl[153] br[153] wl[208] vdd gnd cell_6t
Xbit_r209_c153 bl[153] br[153] wl[209] vdd gnd cell_6t
Xbit_r210_c153 bl[153] br[153] wl[210] vdd gnd cell_6t
Xbit_r211_c153 bl[153] br[153] wl[211] vdd gnd cell_6t
Xbit_r212_c153 bl[153] br[153] wl[212] vdd gnd cell_6t
Xbit_r213_c153 bl[153] br[153] wl[213] vdd gnd cell_6t
Xbit_r214_c153 bl[153] br[153] wl[214] vdd gnd cell_6t
Xbit_r215_c153 bl[153] br[153] wl[215] vdd gnd cell_6t
Xbit_r216_c153 bl[153] br[153] wl[216] vdd gnd cell_6t
Xbit_r217_c153 bl[153] br[153] wl[217] vdd gnd cell_6t
Xbit_r218_c153 bl[153] br[153] wl[218] vdd gnd cell_6t
Xbit_r219_c153 bl[153] br[153] wl[219] vdd gnd cell_6t
Xbit_r220_c153 bl[153] br[153] wl[220] vdd gnd cell_6t
Xbit_r221_c153 bl[153] br[153] wl[221] vdd gnd cell_6t
Xbit_r222_c153 bl[153] br[153] wl[222] vdd gnd cell_6t
Xbit_r223_c153 bl[153] br[153] wl[223] vdd gnd cell_6t
Xbit_r224_c153 bl[153] br[153] wl[224] vdd gnd cell_6t
Xbit_r225_c153 bl[153] br[153] wl[225] vdd gnd cell_6t
Xbit_r226_c153 bl[153] br[153] wl[226] vdd gnd cell_6t
Xbit_r227_c153 bl[153] br[153] wl[227] vdd gnd cell_6t
Xbit_r228_c153 bl[153] br[153] wl[228] vdd gnd cell_6t
Xbit_r229_c153 bl[153] br[153] wl[229] vdd gnd cell_6t
Xbit_r230_c153 bl[153] br[153] wl[230] vdd gnd cell_6t
Xbit_r231_c153 bl[153] br[153] wl[231] vdd gnd cell_6t
Xbit_r232_c153 bl[153] br[153] wl[232] vdd gnd cell_6t
Xbit_r233_c153 bl[153] br[153] wl[233] vdd gnd cell_6t
Xbit_r234_c153 bl[153] br[153] wl[234] vdd gnd cell_6t
Xbit_r235_c153 bl[153] br[153] wl[235] vdd gnd cell_6t
Xbit_r236_c153 bl[153] br[153] wl[236] vdd gnd cell_6t
Xbit_r237_c153 bl[153] br[153] wl[237] vdd gnd cell_6t
Xbit_r238_c153 bl[153] br[153] wl[238] vdd gnd cell_6t
Xbit_r239_c153 bl[153] br[153] wl[239] vdd gnd cell_6t
Xbit_r240_c153 bl[153] br[153] wl[240] vdd gnd cell_6t
Xbit_r241_c153 bl[153] br[153] wl[241] vdd gnd cell_6t
Xbit_r242_c153 bl[153] br[153] wl[242] vdd gnd cell_6t
Xbit_r243_c153 bl[153] br[153] wl[243] vdd gnd cell_6t
Xbit_r244_c153 bl[153] br[153] wl[244] vdd gnd cell_6t
Xbit_r245_c153 bl[153] br[153] wl[245] vdd gnd cell_6t
Xbit_r246_c153 bl[153] br[153] wl[246] vdd gnd cell_6t
Xbit_r247_c153 bl[153] br[153] wl[247] vdd gnd cell_6t
Xbit_r248_c153 bl[153] br[153] wl[248] vdd gnd cell_6t
Xbit_r249_c153 bl[153] br[153] wl[249] vdd gnd cell_6t
Xbit_r250_c153 bl[153] br[153] wl[250] vdd gnd cell_6t
Xbit_r251_c153 bl[153] br[153] wl[251] vdd gnd cell_6t
Xbit_r252_c153 bl[153] br[153] wl[252] vdd gnd cell_6t
Xbit_r253_c153 bl[153] br[153] wl[253] vdd gnd cell_6t
Xbit_r254_c153 bl[153] br[153] wl[254] vdd gnd cell_6t
Xbit_r255_c153 bl[153] br[153] wl[255] vdd gnd cell_6t
Xbit_r0_c154 bl[154] br[154] wl[0] vdd gnd cell_6t
Xbit_r1_c154 bl[154] br[154] wl[1] vdd gnd cell_6t
Xbit_r2_c154 bl[154] br[154] wl[2] vdd gnd cell_6t
Xbit_r3_c154 bl[154] br[154] wl[3] vdd gnd cell_6t
Xbit_r4_c154 bl[154] br[154] wl[4] vdd gnd cell_6t
Xbit_r5_c154 bl[154] br[154] wl[5] vdd gnd cell_6t
Xbit_r6_c154 bl[154] br[154] wl[6] vdd gnd cell_6t
Xbit_r7_c154 bl[154] br[154] wl[7] vdd gnd cell_6t
Xbit_r8_c154 bl[154] br[154] wl[8] vdd gnd cell_6t
Xbit_r9_c154 bl[154] br[154] wl[9] vdd gnd cell_6t
Xbit_r10_c154 bl[154] br[154] wl[10] vdd gnd cell_6t
Xbit_r11_c154 bl[154] br[154] wl[11] vdd gnd cell_6t
Xbit_r12_c154 bl[154] br[154] wl[12] vdd gnd cell_6t
Xbit_r13_c154 bl[154] br[154] wl[13] vdd gnd cell_6t
Xbit_r14_c154 bl[154] br[154] wl[14] vdd gnd cell_6t
Xbit_r15_c154 bl[154] br[154] wl[15] vdd gnd cell_6t
Xbit_r16_c154 bl[154] br[154] wl[16] vdd gnd cell_6t
Xbit_r17_c154 bl[154] br[154] wl[17] vdd gnd cell_6t
Xbit_r18_c154 bl[154] br[154] wl[18] vdd gnd cell_6t
Xbit_r19_c154 bl[154] br[154] wl[19] vdd gnd cell_6t
Xbit_r20_c154 bl[154] br[154] wl[20] vdd gnd cell_6t
Xbit_r21_c154 bl[154] br[154] wl[21] vdd gnd cell_6t
Xbit_r22_c154 bl[154] br[154] wl[22] vdd gnd cell_6t
Xbit_r23_c154 bl[154] br[154] wl[23] vdd gnd cell_6t
Xbit_r24_c154 bl[154] br[154] wl[24] vdd gnd cell_6t
Xbit_r25_c154 bl[154] br[154] wl[25] vdd gnd cell_6t
Xbit_r26_c154 bl[154] br[154] wl[26] vdd gnd cell_6t
Xbit_r27_c154 bl[154] br[154] wl[27] vdd gnd cell_6t
Xbit_r28_c154 bl[154] br[154] wl[28] vdd gnd cell_6t
Xbit_r29_c154 bl[154] br[154] wl[29] vdd gnd cell_6t
Xbit_r30_c154 bl[154] br[154] wl[30] vdd gnd cell_6t
Xbit_r31_c154 bl[154] br[154] wl[31] vdd gnd cell_6t
Xbit_r32_c154 bl[154] br[154] wl[32] vdd gnd cell_6t
Xbit_r33_c154 bl[154] br[154] wl[33] vdd gnd cell_6t
Xbit_r34_c154 bl[154] br[154] wl[34] vdd gnd cell_6t
Xbit_r35_c154 bl[154] br[154] wl[35] vdd gnd cell_6t
Xbit_r36_c154 bl[154] br[154] wl[36] vdd gnd cell_6t
Xbit_r37_c154 bl[154] br[154] wl[37] vdd gnd cell_6t
Xbit_r38_c154 bl[154] br[154] wl[38] vdd gnd cell_6t
Xbit_r39_c154 bl[154] br[154] wl[39] vdd gnd cell_6t
Xbit_r40_c154 bl[154] br[154] wl[40] vdd gnd cell_6t
Xbit_r41_c154 bl[154] br[154] wl[41] vdd gnd cell_6t
Xbit_r42_c154 bl[154] br[154] wl[42] vdd gnd cell_6t
Xbit_r43_c154 bl[154] br[154] wl[43] vdd gnd cell_6t
Xbit_r44_c154 bl[154] br[154] wl[44] vdd gnd cell_6t
Xbit_r45_c154 bl[154] br[154] wl[45] vdd gnd cell_6t
Xbit_r46_c154 bl[154] br[154] wl[46] vdd gnd cell_6t
Xbit_r47_c154 bl[154] br[154] wl[47] vdd gnd cell_6t
Xbit_r48_c154 bl[154] br[154] wl[48] vdd gnd cell_6t
Xbit_r49_c154 bl[154] br[154] wl[49] vdd gnd cell_6t
Xbit_r50_c154 bl[154] br[154] wl[50] vdd gnd cell_6t
Xbit_r51_c154 bl[154] br[154] wl[51] vdd gnd cell_6t
Xbit_r52_c154 bl[154] br[154] wl[52] vdd gnd cell_6t
Xbit_r53_c154 bl[154] br[154] wl[53] vdd gnd cell_6t
Xbit_r54_c154 bl[154] br[154] wl[54] vdd gnd cell_6t
Xbit_r55_c154 bl[154] br[154] wl[55] vdd gnd cell_6t
Xbit_r56_c154 bl[154] br[154] wl[56] vdd gnd cell_6t
Xbit_r57_c154 bl[154] br[154] wl[57] vdd gnd cell_6t
Xbit_r58_c154 bl[154] br[154] wl[58] vdd gnd cell_6t
Xbit_r59_c154 bl[154] br[154] wl[59] vdd gnd cell_6t
Xbit_r60_c154 bl[154] br[154] wl[60] vdd gnd cell_6t
Xbit_r61_c154 bl[154] br[154] wl[61] vdd gnd cell_6t
Xbit_r62_c154 bl[154] br[154] wl[62] vdd gnd cell_6t
Xbit_r63_c154 bl[154] br[154] wl[63] vdd gnd cell_6t
Xbit_r64_c154 bl[154] br[154] wl[64] vdd gnd cell_6t
Xbit_r65_c154 bl[154] br[154] wl[65] vdd gnd cell_6t
Xbit_r66_c154 bl[154] br[154] wl[66] vdd gnd cell_6t
Xbit_r67_c154 bl[154] br[154] wl[67] vdd gnd cell_6t
Xbit_r68_c154 bl[154] br[154] wl[68] vdd gnd cell_6t
Xbit_r69_c154 bl[154] br[154] wl[69] vdd gnd cell_6t
Xbit_r70_c154 bl[154] br[154] wl[70] vdd gnd cell_6t
Xbit_r71_c154 bl[154] br[154] wl[71] vdd gnd cell_6t
Xbit_r72_c154 bl[154] br[154] wl[72] vdd gnd cell_6t
Xbit_r73_c154 bl[154] br[154] wl[73] vdd gnd cell_6t
Xbit_r74_c154 bl[154] br[154] wl[74] vdd gnd cell_6t
Xbit_r75_c154 bl[154] br[154] wl[75] vdd gnd cell_6t
Xbit_r76_c154 bl[154] br[154] wl[76] vdd gnd cell_6t
Xbit_r77_c154 bl[154] br[154] wl[77] vdd gnd cell_6t
Xbit_r78_c154 bl[154] br[154] wl[78] vdd gnd cell_6t
Xbit_r79_c154 bl[154] br[154] wl[79] vdd gnd cell_6t
Xbit_r80_c154 bl[154] br[154] wl[80] vdd gnd cell_6t
Xbit_r81_c154 bl[154] br[154] wl[81] vdd gnd cell_6t
Xbit_r82_c154 bl[154] br[154] wl[82] vdd gnd cell_6t
Xbit_r83_c154 bl[154] br[154] wl[83] vdd gnd cell_6t
Xbit_r84_c154 bl[154] br[154] wl[84] vdd gnd cell_6t
Xbit_r85_c154 bl[154] br[154] wl[85] vdd gnd cell_6t
Xbit_r86_c154 bl[154] br[154] wl[86] vdd gnd cell_6t
Xbit_r87_c154 bl[154] br[154] wl[87] vdd gnd cell_6t
Xbit_r88_c154 bl[154] br[154] wl[88] vdd gnd cell_6t
Xbit_r89_c154 bl[154] br[154] wl[89] vdd gnd cell_6t
Xbit_r90_c154 bl[154] br[154] wl[90] vdd gnd cell_6t
Xbit_r91_c154 bl[154] br[154] wl[91] vdd gnd cell_6t
Xbit_r92_c154 bl[154] br[154] wl[92] vdd gnd cell_6t
Xbit_r93_c154 bl[154] br[154] wl[93] vdd gnd cell_6t
Xbit_r94_c154 bl[154] br[154] wl[94] vdd gnd cell_6t
Xbit_r95_c154 bl[154] br[154] wl[95] vdd gnd cell_6t
Xbit_r96_c154 bl[154] br[154] wl[96] vdd gnd cell_6t
Xbit_r97_c154 bl[154] br[154] wl[97] vdd gnd cell_6t
Xbit_r98_c154 bl[154] br[154] wl[98] vdd gnd cell_6t
Xbit_r99_c154 bl[154] br[154] wl[99] vdd gnd cell_6t
Xbit_r100_c154 bl[154] br[154] wl[100] vdd gnd cell_6t
Xbit_r101_c154 bl[154] br[154] wl[101] vdd gnd cell_6t
Xbit_r102_c154 bl[154] br[154] wl[102] vdd gnd cell_6t
Xbit_r103_c154 bl[154] br[154] wl[103] vdd gnd cell_6t
Xbit_r104_c154 bl[154] br[154] wl[104] vdd gnd cell_6t
Xbit_r105_c154 bl[154] br[154] wl[105] vdd gnd cell_6t
Xbit_r106_c154 bl[154] br[154] wl[106] vdd gnd cell_6t
Xbit_r107_c154 bl[154] br[154] wl[107] vdd gnd cell_6t
Xbit_r108_c154 bl[154] br[154] wl[108] vdd gnd cell_6t
Xbit_r109_c154 bl[154] br[154] wl[109] vdd gnd cell_6t
Xbit_r110_c154 bl[154] br[154] wl[110] vdd gnd cell_6t
Xbit_r111_c154 bl[154] br[154] wl[111] vdd gnd cell_6t
Xbit_r112_c154 bl[154] br[154] wl[112] vdd gnd cell_6t
Xbit_r113_c154 bl[154] br[154] wl[113] vdd gnd cell_6t
Xbit_r114_c154 bl[154] br[154] wl[114] vdd gnd cell_6t
Xbit_r115_c154 bl[154] br[154] wl[115] vdd gnd cell_6t
Xbit_r116_c154 bl[154] br[154] wl[116] vdd gnd cell_6t
Xbit_r117_c154 bl[154] br[154] wl[117] vdd gnd cell_6t
Xbit_r118_c154 bl[154] br[154] wl[118] vdd gnd cell_6t
Xbit_r119_c154 bl[154] br[154] wl[119] vdd gnd cell_6t
Xbit_r120_c154 bl[154] br[154] wl[120] vdd gnd cell_6t
Xbit_r121_c154 bl[154] br[154] wl[121] vdd gnd cell_6t
Xbit_r122_c154 bl[154] br[154] wl[122] vdd gnd cell_6t
Xbit_r123_c154 bl[154] br[154] wl[123] vdd gnd cell_6t
Xbit_r124_c154 bl[154] br[154] wl[124] vdd gnd cell_6t
Xbit_r125_c154 bl[154] br[154] wl[125] vdd gnd cell_6t
Xbit_r126_c154 bl[154] br[154] wl[126] vdd gnd cell_6t
Xbit_r127_c154 bl[154] br[154] wl[127] vdd gnd cell_6t
Xbit_r128_c154 bl[154] br[154] wl[128] vdd gnd cell_6t
Xbit_r129_c154 bl[154] br[154] wl[129] vdd gnd cell_6t
Xbit_r130_c154 bl[154] br[154] wl[130] vdd gnd cell_6t
Xbit_r131_c154 bl[154] br[154] wl[131] vdd gnd cell_6t
Xbit_r132_c154 bl[154] br[154] wl[132] vdd gnd cell_6t
Xbit_r133_c154 bl[154] br[154] wl[133] vdd gnd cell_6t
Xbit_r134_c154 bl[154] br[154] wl[134] vdd gnd cell_6t
Xbit_r135_c154 bl[154] br[154] wl[135] vdd gnd cell_6t
Xbit_r136_c154 bl[154] br[154] wl[136] vdd gnd cell_6t
Xbit_r137_c154 bl[154] br[154] wl[137] vdd gnd cell_6t
Xbit_r138_c154 bl[154] br[154] wl[138] vdd gnd cell_6t
Xbit_r139_c154 bl[154] br[154] wl[139] vdd gnd cell_6t
Xbit_r140_c154 bl[154] br[154] wl[140] vdd gnd cell_6t
Xbit_r141_c154 bl[154] br[154] wl[141] vdd gnd cell_6t
Xbit_r142_c154 bl[154] br[154] wl[142] vdd gnd cell_6t
Xbit_r143_c154 bl[154] br[154] wl[143] vdd gnd cell_6t
Xbit_r144_c154 bl[154] br[154] wl[144] vdd gnd cell_6t
Xbit_r145_c154 bl[154] br[154] wl[145] vdd gnd cell_6t
Xbit_r146_c154 bl[154] br[154] wl[146] vdd gnd cell_6t
Xbit_r147_c154 bl[154] br[154] wl[147] vdd gnd cell_6t
Xbit_r148_c154 bl[154] br[154] wl[148] vdd gnd cell_6t
Xbit_r149_c154 bl[154] br[154] wl[149] vdd gnd cell_6t
Xbit_r150_c154 bl[154] br[154] wl[150] vdd gnd cell_6t
Xbit_r151_c154 bl[154] br[154] wl[151] vdd gnd cell_6t
Xbit_r152_c154 bl[154] br[154] wl[152] vdd gnd cell_6t
Xbit_r153_c154 bl[154] br[154] wl[153] vdd gnd cell_6t
Xbit_r154_c154 bl[154] br[154] wl[154] vdd gnd cell_6t
Xbit_r155_c154 bl[154] br[154] wl[155] vdd gnd cell_6t
Xbit_r156_c154 bl[154] br[154] wl[156] vdd gnd cell_6t
Xbit_r157_c154 bl[154] br[154] wl[157] vdd gnd cell_6t
Xbit_r158_c154 bl[154] br[154] wl[158] vdd gnd cell_6t
Xbit_r159_c154 bl[154] br[154] wl[159] vdd gnd cell_6t
Xbit_r160_c154 bl[154] br[154] wl[160] vdd gnd cell_6t
Xbit_r161_c154 bl[154] br[154] wl[161] vdd gnd cell_6t
Xbit_r162_c154 bl[154] br[154] wl[162] vdd gnd cell_6t
Xbit_r163_c154 bl[154] br[154] wl[163] vdd gnd cell_6t
Xbit_r164_c154 bl[154] br[154] wl[164] vdd gnd cell_6t
Xbit_r165_c154 bl[154] br[154] wl[165] vdd gnd cell_6t
Xbit_r166_c154 bl[154] br[154] wl[166] vdd gnd cell_6t
Xbit_r167_c154 bl[154] br[154] wl[167] vdd gnd cell_6t
Xbit_r168_c154 bl[154] br[154] wl[168] vdd gnd cell_6t
Xbit_r169_c154 bl[154] br[154] wl[169] vdd gnd cell_6t
Xbit_r170_c154 bl[154] br[154] wl[170] vdd gnd cell_6t
Xbit_r171_c154 bl[154] br[154] wl[171] vdd gnd cell_6t
Xbit_r172_c154 bl[154] br[154] wl[172] vdd gnd cell_6t
Xbit_r173_c154 bl[154] br[154] wl[173] vdd gnd cell_6t
Xbit_r174_c154 bl[154] br[154] wl[174] vdd gnd cell_6t
Xbit_r175_c154 bl[154] br[154] wl[175] vdd gnd cell_6t
Xbit_r176_c154 bl[154] br[154] wl[176] vdd gnd cell_6t
Xbit_r177_c154 bl[154] br[154] wl[177] vdd gnd cell_6t
Xbit_r178_c154 bl[154] br[154] wl[178] vdd gnd cell_6t
Xbit_r179_c154 bl[154] br[154] wl[179] vdd gnd cell_6t
Xbit_r180_c154 bl[154] br[154] wl[180] vdd gnd cell_6t
Xbit_r181_c154 bl[154] br[154] wl[181] vdd gnd cell_6t
Xbit_r182_c154 bl[154] br[154] wl[182] vdd gnd cell_6t
Xbit_r183_c154 bl[154] br[154] wl[183] vdd gnd cell_6t
Xbit_r184_c154 bl[154] br[154] wl[184] vdd gnd cell_6t
Xbit_r185_c154 bl[154] br[154] wl[185] vdd gnd cell_6t
Xbit_r186_c154 bl[154] br[154] wl[186] vdd gnd cell_6t
Xbit_r187_c154 bl[154] br[154] wl[187] vdd gnd cell_6t
Xbit_r188_c154 bl[154] br[154] wl[188] vdd gnd cell_6t
Xbit_r189_c154 bl[154] br[154] wl[189] vdd gnd cell_6t
Xbit_r190_c154 bl[154] br[154] wl[190] vdd gnd cell_6t
Xbit_r191_c154 bl[154] br[154] wl[191] vdd gnd cell_6t
Xbit_r192_c154 bl[154] br[154] wl[192] vdd gnd cell_6t
Xbit_r193_c154 bl[154] br[154] wl[193] vdd gnd cell_6t
Xbit_r194_c154 bl[154] br[154] wl[194] vdd gnd cell_6t
Xbit_r195_c154 bl[154] br[154] wl[195] vdd gnd cell_6t
Xbit_r196_c154 bl[154] br[154] wl[196] vdd gnd cell_6t
Xbit_r197_c154 bl[154] br[154] wl[197] vdd gnd cell_6t
Xbit_r198_c154 bl[154] br[154] wl[198] vdd gnd cell_6t
Xbit_r199_c154 bl[154] br[154] wl[199] vdd gnd cell_6t
Xbit_r200_c154 bl[154] br[154] wl[200] vdd gnd cell_6t
Xbit_r201_c154 bl[154] br[154] wl[201] vdd gnd cell_6t
Xbit_r202_c154 bl[154] br[154] wl[202] vdd gnd cell_6t
Xbit_r203_c154 bl[154] br[154] wl[203] vdd gnd cell_6t
Xbit_r204_c154 bl[154] br[154] wl[204] vdd gnd cell_6t
Xbit_r205_c154 bl[154] br[154] wl[205] vdd gnd cell_6t
Xbit_r206_c154 bl[154] br[154] wl[206] vdd gnd cell_6t
Xbit_r207_c154 bl[154] br[154] wl[207] vdd gnd cell_6t
Xbit_r208_c154 bl[154] br[154] wl[208] vdd gnd cell_6t
Xbit_r209_c154 bl[154] br[154] wl[209] vdd gnd cell_6t
Xbit_r210_c154 bl[154] br[154] wl[210] vdd gnd cell_6t
Xbit_r211_c154 bl[154] br[154] wl[211] vdd gnd cell_6t
Xbit_r212_c154 bl[154] br[154] wl[212] vdd gnd cell_6t
Xbit_r213_c154 bl[154] br[154] wl[213] vdd gnd cell_6t
Xbit_r214_c154 bl[154] br[154] wl[214] vdd gnd cell_6t
Xbit_r215_c154 bl[154] br[154] wl[215] vdd gnd cell_6t
Xbit_r216_c154 bl[154] br[154] wl[216] vdd gnd cell_6t
Xbit_r217_c154 bl[154] br[154] wl[217] vdd gnd cell_6t
Xbit_r218_c154 bl[154] br[154] wl[218] vdd gnd cell_6t
Xbit_r219_c154 bl[154] br[154] wl[219] vdd gnd cell_6t
Xbit_r220_c154 bl[154] br[154] wl[220] vdd gnd cell_6t
Xbit_r221_c154 bl[154] br[154] wl[221] vdd gnd cell_6t
Xbit_r222_c154 bl[154] br[154] wl[222] vdd gnd cell_6t
Xbit_r223_c154 bl[154] br[154] wl[223] vdd gnd cell_6t
Xbit_r224_c154 bl[154] br[154] wl[224] vdd gnd cell_6t
Xbit_r225_c154 bl[154] br[154] wl[225] vdd gnd cell_6t
Xbit_r226_c154 bl[154] br[154] wl[226] vdd gnd cell_6t
Xbit_r227_c154 bl[154] br[154] wl[227] vdd gnd cell_6t
Xbit_r228_c154 bl[154] br[154] wl[228] vdd gnd cell_6t
Xbit_r229_c154 bl[154] br[154] wl[229] vdd gnd cell_6t
Xbit_r230_c154 bl[154] br[154] wl[230] vdd gnd cell_6t
Xbit_r231_c154 bl[154] br[154] wl[231] vdd gnd cell_6t
Xbit_r232_c154 bl[154] br[154] wl[232] vdd gnd cell_6t
Xbit_r233_c154 bl[154] br[154] wl[233] vdd gnd cell_6t
Xbit_r234_c154 bl[154] br[154] wl[234] vdd gnd cell_6t
Xbit_r235_c154 bl[154] br[154] wl[235] vdd gnd cell_6t
Xbit_r236_c154 bl[154] br[154] wl[236] vdd gnd cell_6t
Xbit_r237_c154 bl[154] br[154] wl[237] vdd gnd cell_6t
Xbit_r238_c154 bl[154] br[154] wl[238] vdd gnd cell_6t
Xbit_r239_c154 bl[154] br[154] wl[239] vdd gnd cell_6t
Xbit_r240_c154 bl[154] br[154] wl[240] vdd gnd cell_6t
Xbit_r241_c154 bl[154] br[154] wl[241] vdd gnd cell_6t
Xbit_r242_c154 bl[154] br[154] wl[242] vdd gnd cell_6t
Xbit_r243_c154 bl[154] br[154] wl[243] vdd gnd cell_6t
Xbit_r244_c154 bl[154] br[154] wl[244] vdd gnd cell_6t
Xbit_r245_c154 bl[154] br[154] wl[245] vdd gnd cell_6t
Xbit_r246_c154 bl[154] br[154] wl[246] vdd gnd cell_6t
Xbit_r247_c154 bl[154] br[154] wl[247] vdd gnd cell_6t
Xbit_r248_c154 bl[154] br[154] wl[248] vdd gnd cell_6t
Xbit_r249_c154 bl[154] br[154] wl[249] vdd gnd cell_6t
Xbit_r250_c154 bl[154] br[154] wl[250] vdd gnd cell_6t
Xbit_r251_c154 bl[154] br[154] wl[251] vdd gnd cell_6t
Xbit_r252_c154 bl[154] br[154] wl[252] vdd gnd cell_6t
Xbit_r253_c154 bl[154] br[154] wl[253] vdd gnd cell_6t
Xbit_r254_c154 bl[154] br[154] wl[254] vdd gnd cell_6t
Xbit_r255_c154 bl[154] br[154] wl[255] vdd gnd cell_6t
Xbit_r0_c155 bl[155] br[155] wl[0] vdd gnd cell_6t
Xbit_r1_c155 bl[155] br[155] wl[1] vdd gnd cell_6t
Xbit_r2_c155 bl[155] br[155] wl[2] vdd gnd cell_6t
Xbit_r3_c155 bl[155] br[155] wl[3] vdd gnd cell_6t
Xbit_r4_c155 bl[155] br[155] wl[4] vdd gnd cell_6t
Xbit_r5_c155 bl[155] br[155] wl[5] vdd gnd cell_6t
Xbit_r6_c155 bl[155] br[155] wl[6] vdd gnd cell_6t
Xbit_r7_c155 bl[155] br[155] wl[7] vdd gnd cell_6t
Xbit_r8_c155 bl[155] br[155] wl[8] vdd gnd cell_6t
Xbit_r9_c155 bl[155] br[155] wl[9] vdd gnd cell_6t
Xbit_r10_c155 bl[155] br[155] wl[10] vdd gnd cell_6t
Xbit_r11_c155 bl[155] br[155] wl[11] vdd gnd cell_6t
Xbit_r12_c155 bl[155] br[155] wl[12] vdd gnd cell_6t
Xbit_r13_c155 bl[155] br[155] wl[13] vdd gnd cell_6t
Xbit_r14_c155 bl[155] br[155] wl[14] vdd gnd cell_6t
Xbit_r15_c155 bl[155] br[155] wl[15] vdd gnd cell_6t
Xbit_r16_c155 bl[155] br[155] wl[16] vdd gnd cell_6t
Xbit_r17_c155 bl[155] br[155] wl[17] vdd gnd cell_6t
Xbit_r18_c155 bl[155] br[155] wl[18] vdd gnd cell_6t
Xbit_r19_c155 bl[155] br[155] wl[19] vdd gnd cell_6t
Xbit_r20_c155 bl[155] br[155] wl[20] vdd gnd cell_6t
Xbit_r21_c155 bl[155] br[155] wl[21] vdd gnd cell_6t
Xbit_r22_c155 bl[155] br[155] wl[22] vdd gnd cell_6t
Xbit_r23_c155 bl[155] br[155] wl[23] vdd gnd cell_6t
Xbit_r24_c155 bl[155] br[155] wl[24] vdd gnd cell_6t
Xbit_r25_c155 bl[155] br[155] wl[25] vdd gnd cell_6t
Xbit_r26_c155 bl[155] br[155] wl[26] vdd gnd cell_6t
Xbit_r27_c155 bl[155] br[155] wl[27] vdd gnd cell_6t
Xbit_r28_c155 bl[155] br[155] wl[28] vdd gnd cell_6t
Xbit_r29_c155 bl[155] br[155] wl[29] vdd gnd cell_6t
Xbit_r30_c155 bl[155] br[155] wl[30] vdd gnd cell_6t
Xbit_r31_c155 bl[155] br[155] wl[31] vdd gnd cell_6t
Xbit_r32_c155 bl[155] br[155] wl[32] vdd gnd cell_6t
Xbit_r33_c155 bl[155] br[155] wl[33] vdd gnd cell_6t
Xbit_r34_c155 bl[155] br[155] wl[34] vdd gnd cell_6t
Xbit_r35_c155 bl[155] br[155] wl[35] vdd gnd cell_6t
Xbit_r36_c155 bl[155] br[155] wl[36] vdd gnd cell_6t
Xbit_r37_c155 bl[155] br[155] wl[37] vdd gnd cell_6t
Xbit_r38_c155 bl[155] br[155] wl[38] vdd gnd cell_6t
Xbit_r39_c155 bl[155] br[155] wl[39] vdd gnd cell_6t
Xbit_r40_c155 bl[155] br[155] wl[40] vdd gnd cell_6t
Xbit_r41_c155 bl[155] br[155] wl[41] vdd gnd cell_6t
Xbit_r42_c155 bl[155] br[155] wl[42] vdd gnd cell_6t
Xbit_r43_c155 bl[155] br[155] wl[43] vdd gnd cell_6t
Xbit_r44_c155 bl[155] br[155] wl[44] vdd gnd cell_6t
Xbit_r45_c155 bl[155] br[155] wl[45] vdd gnd cell_6t
Xbit_r46_c155 bl[155] br[155] wl[46] vdd gnd cell_6t
Xbit_r47_c155 bl[155] br[155] wl[47] vdd gnd cell_6t
Xbit_r48_c155 bl[155] br[155] wl[48] vdd gnd cell_6t
Xbit_r49_c155 bl[155] br[155] wl[49] vdd gnd cell_6t
Xbit_r50_c155 bl[155] br[155] wl[50] vdd gnd cell_6t
Xbit_r51_c155 bl[155] br[155] wl[51] vdd gnd cell_6t
Xbit_r52_c155 bl[155] br[155] wl[52] vdd gnd cell_6t
Xbit_r53_c155 bl[155] br[155] wl[53] vdd gnd cell_6t
Xbit_r54_c155 bl[155] br[155] wl[54] vdd gnd cell_6t
Xbit_r55_c155 bl[155] br[155] wl[55] vdd gnd cell_6t
Xbit_r56_c155 bl[155] br[155] wl[56] vdd gnd cell_6t
Xbit_r57_c155 bl[155] br[155] wl[57] vdd gnd cell_6t
Xbit_r58_c155 bl[155] br[155] wl[58] vdd gnd cell_6t
Xbit_r59_c155 bl[155] br[155] wl[59] vdd gnd cell_6t
Xbit_r60_c155 bl[155] br[155] wl[60] vdd gnd cell_6t
Xbit_r61_c155 bl[155] br[155] wl[61] vdd gnd cell_6t
Xbit_r62_c155 bl[155] br[155] wl[62] vdd gnd cell_6t
Xbit_r63_c155 bl[155] br[155] wl[63] vdd gnd cell_6t
Xbit_r64_c155 bl[155] br[155] wl[64] vdd gnd cell_6t
Xbit_r65_c155 bl[155] br[155] wl[65] vdd gnd cell_6t
Xbit_r66_c155 bl[155] br[155] wl[66] vdd gnd cell_6t
Xbit_r67_c155 bl[155] br[155] wl[67] vdd gnd cell_6t
Xbit_r68_c155 bl[155] br[155] wl[68] vdd gnd cell_6t
Xbit_r69_c155 bl[155] br[155] wl[69] vdd gnd cell_6t
Xbit_r70_c155 bl[155] br[155] wl[70] vdd gnd cell_6t
Xbit_r71_c155 bl[155] br[155] wl[71] vdd gnd cell_6t
Xbit_r72_c155 bl[155] br[155] wl[72] vdd gnd cell_6t
Xbit_r73_c155 bl[155] br[155] wl[73] vdd gnd cell_6t
Xbit_r74_c155 bl[155] br[155] wl[74] vdd gnd cell_6t
Xbit_r75_c155 bl[155] br[155] wl[75] vdd gnd cell_6t
Xbit_r76_c155 bl[155] br[155] wl[76] vdd gnd cell_6t
Xbit_r77_c155 bl[155] br[155] wl[77] vdd gnd cell_6t
Xbit_r78_c155 bl[155] br[155] wl[78] vdd gnd cell_6t
Xbit_r79_c155 bl[155] br[155] wl[79] vdd gnd cell_6t
Xbit_r80_c155 bl[155] br[155] wl[80] vdd gnd cell_6t
Xbit_r81_c155 bl[155] br[155] wl[81] vdd gnd cell_6t
Xbit_r82_c155 bl[155] br[155] wl[82] vdd gnd cell_6t
Xbit_r83_c155 bl[155] br[155] wl[83] vdd gnd cell_6t
Xbit_r84_c155 bl[155] br[155] wl[84] vdd gnd cell_6t
Xbit_r85_c155 bl[155] br[155] wl[85] vdd gnd cell_6t
Xbit_r86_c155 bl[155] br[155] wl[86] vdd gnd cell_6t
Xbit_r87_c155 bl[155] br[155] wl[87] vdd gnd cell_6t
Xbit_r88_c155 bl[155] br[155] wl[88] vdd gnd cell_6t
Xbit_r89_c155 bl[155] br[155] wl[89] vdd gnd cell_6t
Xbit_r90_c155 bl[155] br[155] wl[90] vdd gnd cell_6t
Xbit_r91_c155 bl[155] br[155] wl[91] vdd gnd cell_6t
Xbit_r92_c155 bl[155] br[155] wl[92] vdd gnd cell_6t
Xbit_r93_c155 bl[155] br[155] wl[93] vdd gnd cell_6t
Xbit_r94_c155 bl[155] br[155] wl[94] vdd gnd cell_6t
Xbit_r95_c155 bl[155] br[155] wl[95] vdd gnd cell_6t
Xbit_r96_c155 bl[155] br[155] wl[96] vdd gnd cell_6t
Xbit_r97_c155 bl[155] br[155] wl[97] vdd gnd cell_6t
Xbit_r98_c155 bl[155] br[155] wl[98] vdd gnd cell_6t
Xbit_r99_c155 bl[155] br[155] wl[99] vdd gnd cell_6t
Xbit_r100_c155 bl[155] br[155] wl[100] vdd gnd cell_6t
Xbit_r101_c155 bl[155] br[155] wl[101] vdd gnd cell_6t
Xbit_r102_c155 bl[155] br[155] wl[102] vdd gnd cell_6t
Xbit_r103_c155 bl[155] br[155] wl[103] vdd gnd cell_6t
Xbit_r104_c155 bl[155] br[155] wl[104] vdd gnd cell_6t
Xbit_r105_c155 bl[155] br[155] wl[105] vdd gnd cell_6t
Xbit_r106_c155 bl[155] br[155] wl[106] vdd gnd cell_6t
Xbit_r107_c155 bl[155] br[155] wl[107] vdd gnd cell_6t
Xbit_r108_c155 bl[155] br[155] wl[108] vdd gnd cell_6t
Xbit_r109_c155 bl[155] br[155] wl[109] vdd gnd cell_6t
Xbit_r110_c155 bl[155] br[155] wl[110] vdd gnd cell_6t
Xbit_r111_c155 bl[155] br[155] wl[111] vdd gnd cell_6t
Xbit_r112_c155 bl[155] br[155] wl[112] vdd gnd cell_6t
Xbit_r113_c155 bl[155] br[155] wl[113] vdd gnd cell_6t
Xbit_r114_c155 bl[155] br[155] wl[114] vdd gnd cell_6t
Xbit_r115_c155 bl[155] br[155] wl[115] vdd gnd cell_6t
Xbit_r116_c155 bl[155] br[155] wl[116] vdd gnd cell_6t
Xbit_r117_c155 bl[155] br[155] wl[117] vdd gnd cell_6t
Xbit_r118_c155 bl[155] br[155] wl[118] vdd gnd cell_6t
Xbit_r119_c155 bl[155] br[155] wl[119] vdd gnd cell_6t
Xbit_r120_c155 bl[155] br[155] wl[120] vdd gnd cell_6t
Xbit_r121_c155 bl[155] br[155] wl[121] vdd gnd cell_6t
Xbit_r122_c155 bl[155] br[155] wl[122] vdd gnd cell_6t
Xbit_r123_c155 bl[155] br[155] wl[123] vdd gnd cell_6t
Xbit_r124_c155 bl[155] br[155] wl[124] vdd gnd cell_6t
Xbit_r125_c155 bl[155] br[155] wl[125] vdd gnd cell_6t
Xbit_r126_c155 bl[155] br[155] wl[126] vdd gnd cell_6t
Xbit_r127_c155 bl[155] br[155] wl[127] vdd gnd cell_6t
Xbit_r128_c155 bl[155] br[155] wl[128] vdd gnd cell_6t
Xbit_r129_c155 bl[155] br[155] wl[129] vdd gnd cell_6t
Xbit_r130_c155 bl[155] br[155] wl[130] vdd gnd cell_6t
Xbit_r131_c155 bl[155] br[155] wl[131] vdd gnd cell_6t
Xbit_r132_c155 bl[155] br[155] wl[132] vdd gnd cell_6t
Xbit_r133_c155 bl[155] br[155] wl[133] vdd gnd cell_6t
Xbit_r134_c155 bl[155] br[155] wl[134] vdd gnd cell_6t
Xbit_r135_c155 bl[155] br[155] wl[135] vdd gnd cell_6t
Xbit_r136_c155 bl[155] br[155] wl[136] vdd gnd cell_6t
Xbit_r137_c155 bl[155] br[155] wl[137] vdd gnd cell_6t
Xbit_r138_c155 bl[155] br[155] wl[138] vdd gnd cell_6t
Xbit_r139_c155 bl[155] br[155] wl[139] vdd gnd cell_6t
Xbit_r140_c155 bl[155] br[155] wl[140] vdd gnd cell_6t
Xbit_r141_c155 bl[155] br[155] wl[141] vdd gnd cell_6t
Xbit_r142_c155 bl[155] br[155] wl[142] vdd gnd cell_6t
Xbit_r143_c155 bl[155] br[155] wl[143] vdd gnd cell_6t
Xbit_r144_c155 bl[155] br[155] wl[144] vdd gnd cell_6t
Xbit_r145_c155 bl[155] br[155] wl[145] vdd gnd cell_6t
Xbit_r146_c155 bl[155] br[155] wl[146] vdd gnd cell_6t
Xbit_r147_c155 bl[155] br[155] wl[147] vdd gnd cell_6t
Xbit_r148_c155 bl[155] br[155] wl[148] vdd gnd cell_6t
Xbit_r149_c155 bl[155] br[155] wl[149] vdd gnd cell_6t
Xbit_r150_c155 bl[155] br[155] wl[150] vdd gnd cell_6t
Xbit_r151_c155 bl[155] br[155] wl[151] vdd gnd cell_6t
Xbit_r152_c155 bl[155] br[155] wl[152] vdd gnd cell_6t
Xbit_r153_c155 bl[155] br[155] wl[153] vdd gnd cell_6t
Xbit_r154_c155 bl[155] br[155] wl[154] vdd gnd cell_6t
Xbit_r155_c155 bl[155] br[155] wl[155] vdd gnd cell_6t
Xbit_r156_c155 bl[155] br[155] wl[156] vdd gnd cell_6t
Xbit_r157_c155 bl[155] br[155] wl[157] vdd gnd cell_6t
Xbit_r158_c155 bl[155] br[155] wl[158] vdd gnd cell_6t
Xbit_r159_c155 bl[155] br[155] wl[159] vdd gnd cell_6t
Xbit_r160_c155 bl[155] br[155] wl[160] vdd gnd cell_6t
Xbit_r161_c155 bl[155] br[155] wl[161] vdd gnd cell_6t
Xbit_r162_c155 bl[155] br[155] wl[162] vdd gnd cell_6t
Xbit_r163_c155 bl[155] br[155] wl[163] vdd gnd cell_6t
Xbit_r164_c155 bl[155] br[155] wl[164] vdd gnd cell_6t
Xbit_r165_c155 bl[155] br[155] wl[165] vdd gnd cell_6t
Xbit_r166_c155 bl[155] br[155] wl[166] vdd gnd cell_6t
Xbit_r167_c155 bl[155] br[155] wl[167] vdd gnd cell_6t
Xbit_r168_c155 bl[155] br[155] wl[168] vdd gnd cell_6t
Xbit_r169_c155 bl[155] br[155] wl[169] vdd gnd cell_6t
Xbit_r170_c155 bl[155] br[155] wl[170] vdd gnd cell_6t
Xbit_r171_c155 bl[155] br[155] wl[171] vdd gnd cell_6t
Xbit_r172_c155 bl[155] br[155] wl[172] vdd gnd cell_6t
Xbit_r173_c155 bl[155] br[155] wl[173] vdd gnd cell_6t
Xbit_r174_c155 bl[155] br[155] wl[174] vdd gnd cell_6t
Xbit_r175_c155 bl[155] br[155] wl[175] vdd gnd cell_6t
Xbit_r176_c155 bl[155] br[155] wl[176] vdd gnd cell_6t
Xbit_r177_c155 bl[155] br[155] wl[177] vdd gnd cell_6t
Xbit_r178_c155 bl[155] br[155] wl[178] vdd gnd cell_6t
Xbit_r179_c155 bl[155] br[155] wl[179] vdd gnd cell_6t
Xbit_r180_c155 bl[155] br[155] wl[180] vdd gnd cell_6t
Xbit_r181_c155 bl[155] br[155] wl[181] vdd gnd cell_6t
Xbit_r182_c155 bl[155] br[155] wl[182] vdd gnd cell_6t
Xbit_r183_c155 bl[155] br[155] wl[183] vdd gnd cell_6t
Xbit_r184_c155 bl[155] br[155] wl[184] vdd gnd cell_6t
Xbit_r185_c155 bl[155] br[155] wl[185] vdd gnd cell_6t
Xbit_r186_c155 bl[155] br[155] wl[186] vdd gnd cell_6t
Xbit_r187_c155 bl[155] br[155] wl[187] vdd gnd cell_6t
Xbit_r188_c155 bl[155] br[155] wl[188] vdd gnd cell_6t
Xbit_r189_c155 bl[155] br[155] wl[189] vdd gnd cell_6t
Xbit_r190_c155 bl[155] br[155] wl[190] vdd gnd cell_6t
Xbit_r191_c155 bl[155] br[155] wl[191] vdd gnd cell_6t
Xbit_r192_c155 bl[155] br[155] wl[192] vdd gnd cell_6t
Xbit_r193_c155 bl[155] br[155] wl[193] vdd gnd cell_6t
Xbit_r194_c155 bl[155] br[155] wl[194] vdd gnd cell_6t
Xbit_r195_c155 bl[155] br[155] wl[195] vdd gnd cell_6t
Xbit_r196_c155 bl[155] br[155] wl[196] vdd gnd cell_6t
Xbit_r197_c155 bl[155] br[155] wl[197] vdd gnd cell_6t
Xbit_r198_c155 bl[155] br[155] wl[198] vdd gnd cell_6t
Xbit_r199_c155 bl[155] br[155] wl[199] vdd gnd cell_6t
Xbit_r200_c155 bl[155] br[155] wl[200] vdd gnd cell_6t
Xbit_r201_c155 bl[155] br[155] wl[201] vdd gnd cell_6t
Xbit_r202_c155 bl[155] br[155] wl[202] vdd gnd cell_6t
Xbit_r203_c155 bl[155] br[155] wl[203] vdd gnd cell_6t
Xbit_r204_c155 bl[155] br[155] wl[204] vdd gnd cell_6t
Xbit_r205_c155 bl[155] br[155] wl[205] vdd gnd cell_6t
Xbit_r206_c155 bl[155] br[155] wl[206] vdd gnd cell_6t
Xbit_r207_c155 bl[155] br[155] wl[207] vdd gnd cell_6t
Xbit_r208_c155 bl[155] br[155] wl[208] vdd gnd cell_6t
Xbit_r209_c155 bl[155] br[155] wl[209] vdd gnd cell_6t
Xbit_r210_c155 bl[155] br[155] wl[210] vdd gnd cell_6t
Xbit_r211_c155 bl[155] br[155] wl[211] vdd gnd cell_6t
Xbit_r212_c155 bl[155] br[155] wl[212] vdd gnd cell_6t
Xbit_r213_c155 bl[155] br[155] wl[213] vdd gnd cell_6t
Xbit_r214_c155 bl[155] br[155] wl[214] vdd gnd cell_6t
Xbit_r215_c155 bl[155] br[155] wl[215] vdd gnd cell_6t
Xbit_r216_c155 bl[155] br[155] wl[216] vdd gnd cell_6t
Xbit_r217_c155 bl[155] br[155] wl[217] vdd gnd cell_6t
Xbit_r218_c155 bl[155] br[155] wl[218] vdd gnd cell_6t
Xbit_r219_c155 bl[155] br[155] wl[219] vdd gnd cell_6t
Xbit_r220_c155 bl[155] br[155] wl[220] vdd gnd cell_6t
Xbit_r221_c155 bl[155] br[155] wl[221] vdd gnd cell_6t
Xbit_r222_c155 bl[155] br[155] wl[222] vdd gnd cell_6t
Xbit_r223_c155 bl[155] br[155] wl[223] vdd gnd cell_6t
Xbit_r224_c155 bl[155] br[155] wl[224] vdd gnd cell_6t
Xbit_r225_c155 bl[155] br[155] wl[225] vdd gnd cell_6t
Xbit_r226_c155 bl[155] br[155] wl[226] vdd gnd cell_6t
Xbit_r227_c155 bl[155] br[155] wl[227] vdd gnd cell_6t
Xbit_r228_c155 bl[155] br[155] wl[228] vdd gnd cell_6t
Xbit_r229_c155 bl[155] br[155] wl[229] vdd gnd cell_6t
Xbit_r230_c155 bl[155] br[155] wl[230] vdd gnd cell_6t
Xbit_r231_c155 bl[155] br[155] wl[231] vdd gnd cell_6t
Xbit_r232_c155 bl[155] br[155] wl[232] vdd gnd cell_6t
Xbit_r233_c155 bl[155] br[155] wl[233] vdd gnd cell_6t
Xbit_r234_c155 bl[155] br[155] wl[234] vdd gnd cell_6t
Xbit_r235_c155 bl[155] br[155] wl[235] vdd gnd cell_6t
Xbit_r236_c155 bl[155] br[155] wl[236] vdd gnd cell_6t
Xbit_r237_c155 bl[155] br[155] wl[237] vdd gnd cell_6t
Xbit_r238_c155 bl[155] br[155] wl[238] vdd gnd cell_6t
Xbit_r239_c155 bl[155] br[155] wl[239] vdd gnd cell_6t
Xbit_r240_c155 bl[155] br[155] wl[240] vdd gnd cell_6t
Xbit_r241_c155 bl[155] br[155] wl[241] vdd gnd cell_6t
Xbit_r242_c155 bl[155] br[155] wl[242] vdd gnd cell_6t
Xbit_r243_c155 bl[155] br[155] wl[243] vdd gnd cell_6t
Xbit_r244_c155 bl[155] br[155] wl[244] vdd gnd cell_6t
Xbit_r245_c155 bl[155] br[155] wl[245] vdd gnd cell_6t
Xbit_r246_c155 bl[155] br[155] wl[246] vdd gnd cell_6t
Xbit_r247_c155 bl[155] br[155] wl[247] vdd gnd cell_6t
Xbit_r248_c155 bl[155] br[155] wl[248] vdd gnd cell_6t
Xbit_r249_c155 bl[155] br[155] wl[249] vdd gnd cell_6t
Xbit_r250_c155 bl[155] br[155] wl[250] vdd gnd cell_6t
Xbit_r251_c155 bl[155] br[155] wl[251] vdd gnd cell_6t
Xbit_r252_c155 bl[155] br[155] wl[252] vdd gnd cell_6t
Xbit_r253_c155 bl[155] br[155] wl[253] vdd gnd cell_6t
Xbit_r254_c155 bl[155] br[155] wl[254] vdd gnd cell_6t
Xbit_r255_c155 bl[155] br[155] wl[255] vdd gnd cell_6t
Xbit_r0_c156 bl[156] br[156] wl[0] vdd gnd cell_6t
Xbit_r1_c156 bl[156] br[156] wl[1] vdd gnd cell_6t
Xbit_r2_c156 bl[156] br[156] wl[2] vdd gnd cell_6t
Xbit_r3_c156 bl[156] br[156] wl[3] vdd gnd cell_6t
Xbit_r4_c156 bl[156] br[156] wl[4] vdd gnd cell_6t
Xbit_r5_c156 bl[156] br[156] wl[5] vdd gnd cell_6t
Xbit_r6_c156 bl[156] br[156] wl[6] vdd gnd cell_6t
Xbit_r7_c156 bl[156] br[156] wl[7] vdd gnd cell_6t
Xbit_r8_c156 bl[156] br[156] wl[8] vdd gnd cell_6t
Xbit_r9_c156 bl[156] br[156] wl[9] vdd gnd cell_6t
Xbit_r10_c156 bl[156] br[156] wl[10] vdd gnd cell_6t
Xbit_r11_c156 bl[156] br[156] wl[11] vdd gnd cell_6t
Xbit_r12_c156 bl[156] br[156] wl[12] vdd gnd cell_6t
Xbit_r13_c156 bl[156] br[156] wl[13] vdd gnd cell_6t
Xbit_r14_c156 bl[156] br[156] wl[14] vdd gnd cell_6t
Xbit_r15_c156 bl[156] br[156] wl[15] vdd gnd cell_6t
Xbit_r16_c156 bl[156] br[156] wl[16] vdd gnd cell_6t
Xbit_r17_c156 bl[156] br[156] wl[17] vdd gnd cell_6t
Xbit_r18_c156 bl[156] br[156] wl[18] vdd gnd cell_6t
Xbit_r19_c156 bl[156] br[156] wl[19] vdd gnd cell_6t
Xbit_r20_c156 bl[156] br[156] wl[20] vdd gnd cell_6t
Xbit_r21_c156 bl[156] br[156] wl[21] vdd gnd cell_6t
Xbit_r22_c156 bl[156] br[156] wl[22] vdd gnd cell_6t
Xbit_r23_c156 bl[156] br[156] wl[23] vdd gnd cell_6t
Xbit_r24_c156 bl[156] br[156] wl[24] vdd gnd cell_6t
Xbit_r25_c156 bl[156] br[156] wl[25] vdd gnd cell_6t
Xbit_r26_c156 bl[156] br[156] wl[26] vdd gnd cell_6t
Xbit_r27_c156 bl[156] br[156] wl[27] vdd gnd cell_6t
Xbit_r28_c156 bl[156] br[156] wl[28] vdd gnd cell_6t
Xbit_r29_c156 bl[156] br[156] wl[29] vdd gnd cell_6t
Xbit_r30_c156 bl[156] br[156] wl[30] vdd gnd cell_6t
Xbit_r31_c156 bl[156] br[156] wl[31] vdd gnd cell_6t
Xbit_r32_c156 bl[156] br[156] wl[32] vdd gnd cell_6t
Xbit_r33_c156 bl[156] br[156] wl[33] vdd gnd cell_6t
Xbit_r34_c156 bl[156] br[156] wl[34] vdd gnd cell_6t
Xbit_r35_c156 bl[156] br[156] wl[35] vdd gnd cell_6t
Xbit_r36_c156 bl[156] br[156] wl[36] vdd gnd cell_6t
Xbit_r37_c156 bl[156] br[156] wl[37] vdd gnd cell_6t
Xbit_r38_c156 bl[156] br[156] wl[38] vdd gnd cell_6t
Xbit_r39_c156 bl[156] br[156] wl[39] vdd gnd cell_6t
Xbit_r40_c156 bl[156] br[156] wl[40] vdd gnd cell_6t
Xbit_r41_c156 bl[156] br[156] wl[41] vdd gnd cell_6t
Xbit_r42_c156 bl[156] br[156] wl[42] vdd gnd cell_6t
Xbit_r43_c156 bl[156] br[156] wl[43] vdd gnd cell_6t
Xbit_r44_c156 bl[156] br[156] wl[44] vdd gnd cell_6t
Xbit_r45_c156 bl[156] br[156] wl[45] vdd gnd cell_6t
Xbit_r46_c156 bl[156] br[156] wl[46] vdd gnd cell_6t
Xbit_r47_c156 bl[156] br[156] wl[47] vdd gnd cell_6t
Xbit_r48_c156 bl[156] br[156] wl[48] vdd gnd cell_6t
Xbit_r49_c156 bl[156] br[156] wl[49] vdd gnd cell_6t
Xbit_r50_c156 bl[156] br[156] wl[50] vdd gnd cell_6t
Xbit_r51_c156 bl[156] br[156] wl[51] vdd gnd cell_6t
Xbit_r52_c156 bl[156] br[156] wl[52] vdd gnd cell_6t
Xbit_r53_c156 bl[156] br[156] wl[53] vdd gnd cell_6t
Xbit_r54_c156 bl[156] br[156] wl[54] vdd gnd cell_6t
Xbit_r55_c156 bl[156] br[156] wl[55] vdd gnd cell_6t
Xbit_r56_c156 bl[156] br[156] wl[56] vdd gnd cell_6t
Xbit_r57_c156 bl[156] br[156] wl[57] vdd gnd cell_6t
Xbit_r58_c156 bl[156] br[156] wl[58] vdd gnd cell_6t
Xbit_r59_c156 bl[156] br[156] wl[59] vdd gnd cell_6t
Xbit_r60_c156 bl[156] br[156] wl[60] vdd gnd cell_6t
Xbit_r61_c156 bl[156] br[156] wl[61] vdd gnd cell_6t
Xbit_r62_c156 bl[156] br[156] wl[62] vdd gnd cell_6t
Xbit_r63_c156 bl[156] br[156] wl[63] vdd gnd cell_6t
Xbit_r64_c156 bl[156] br[156] wl[64] vdd gnd cell_6t
Xbit_r65_c156 bl[156] br[156] wl[65] vdd gnd cell_6t
Xbit_r66_c156 bl[156] br[156] wl[66] vdd gnd cell_6t
Xbit_r67_c156 bl[156] br[156] wl[67] vdd gnd cell_6t
Xbit_r68_c156 bl[156] br[156] wl[68] vdd gnd cell_6t
Xbit_r69_c156 bl[156] br[156] wl[69] vdd gnd cell_6t
Xbit_r70_c156 bl[156] br[156] wl[70] vdd gnd cell_6t
Xbit_r71_c156 bl[156] br[156] wl[71] vdd gnd cell_6t
Xbit_r72_c156 bl[156] br[156] wl[72] vdd gnd cell_6t
Xbit_r73_c156 bl[156] br[156] wl[73] vdd gnd cell_6t
Xbit_r74_c156 bl[156] br[156] wl[74] vdd gnd cell_6t
Xbit_r75_c156 bl[156] br[156] wl[75] vdd gnd cell_6t
Xbit_r76_c156 bl[156] br[156] wl[76] vdd gnd cell_6t
Xbit_r77_c156 bl[156] br[156] wl[77] vdd gnd cell_6t
Xbit_r78_c156 bl[156] br[156] wl[78] vdd gnd cell_6t
Xbit_r79_c156 bl[156] br[156] wl[79] vdd gnd cell_6t
Xbit_r80_c156 bl[156] br[156] wl[80] vdd gnd cell_6t
Xbit_r81_c156 bl[156] br[156] wl[81] vdd gnd cell_6t
Xbit_r82_c156 bl[156] br[156] wl[82] vdd gnd cell_6t
Xbit_r83_c156 bl[156] br[156] wl[83] vdd gnd cell_6t
Xbit_r84_c156 bl[156] br[156] wl[84] vdd gnd cell_6t
Xbit_r85_c156 bl[156] br[156] wl[85] vdd gnd cell_6t
Xbit_r86_c156 bl[156] br[156] wl[86] vdd gnd cell_6t
Xbit_r87_c156 bl[156] br[156] wl[87] vdd gnd cell_6t
Xbit_r88_c156 bl[156] br[156] wl[88] vdd gnd cell_6t
Xbit_r89_c156 bl[156] br[156] wl[89] vdd gnd cell_6t
Xbit_r90_c156 bl[156] br[156] wl[90] vdd gnd cell_6t
Xbit_r91_c156 bl[156] br[156] wl[91] vdd gnd cell_6t
Xbit_r92_c156 bl[156] br[156] wl[92] vdd gnd cell_6t
Xbit_r93_c156 bl[156] br[156] wl[93] vdd gnd cell_6t
Xbit_r94_c156 bl[156] br[156] wl[94] vdd gnd cell_6t
Xbit_r95_c156 bl[156] br[156] wl[95] vdd gnd cell_6t
Xbit_r96_c156 bl[156] br[156] wl[96] vdd gnd cell_6t
Xbit_r97_c156 bl[156] br[156] wl[97] vdd gnd cell_6t
Xbit_r98_c156 bl[156] br[156] wl[98] vdd gnd cell_6t
Xbit_r99_c156 bl[156] br[156] wl[99] vdd gnd cell_6t
Xbit_r100_c156 bl[156] br[156] wl[100] vdd gnd cell_6t
Xbit_r101_c156 bl[156] br[156] wl[101] vdd gnd cell_6t
Xbit_r102_c156 bl[156] br[156] wl[102] vdd gnd cell_6t
Xbit_r103_c156 bl[156] br[156] wl[103] vdd gnd cell_6t
Xbit_r104_c156 bl[156] br[156] wl[104] vdd gnd cell_6t
Xbit_r105_c156 bl[156] br[156] wl[105] vdd gnd cell_6t
Xbit_r106_c156 bl[156] br[156] wl[106] vdd gnd cell_6t
Xbit_r107_c156 bl[156] br[156] wl[107] vdd gnd cell_6t
Xbit_r108_c156 bl[156] br[156] wl[108] vdd gnd cell_6t
Xbit_r109_c156 bl[156] br[156] wl[109] vdd gnd cell_6t
Xbit_r110_c156 bl[156] br[156] wl[110] vdd gnd cell_6t
Xbit_r111_c156 bl[156] br[156] wl[111] vdd gnd cell_6t
Xbit_r112_c156 bl[156] br[156] wl[112] vdd gnd cell_6t
Xbit_r113_c156 bl[156] br[156] wl[113] vdd gnd cell_6t
Xbit_r114_c156 bl[156] br[156] wl[114] vdd gnd cell_6t
Xbit_r115_c156 bl[156] br[156] wl[115] vdd gnd cell_6t
Xbit_r116_c156 bl[156] br[156] wl[116] vdd gnd cell_6t
Xbit_r117_c156 bl[156] br[156] wl[117] vdd gnd cell_6t
Xbit_r118_c156 bl[156] br[156] wl[118] vdd gnd cell_6t
Xbit_r119_c156 bl[156] br[156] wl[119] vdd gnd cell_6t
Xbit_r120_c156 bl[156] br[156] wl[120] vdd gnd cell_6t
Xbit_r121_c156 bl[156] br[156] wl[121] vdd gnd cell_6t
Xbit_r122_c156 bl[156] br[156] wl[122] vdd gnd cell_6t
Xbit_r123_c156 bl[156] br[156] wl[123] vdd gnd cell_6t
Xbit_r124_c156 bl[156] br[156] wl[124] vdd gnd cell_6t
Xbit_r125_c156 bl[156] br[156] wl[125] vdd gnd cell_6t
Xbit_r126_c156 bl[156] br[156] wl[126] vdd gnd cell_6t
Xbit_r127_c156 bl[156] br[156] wl[127] vdd gnd cell_6t
Xbit_r128_c156 bl[156] br[156] wl[128] vdd gnd cell_6t
Xbit_r129_c156 bl[156] br[156] wl[129] vdd gnd cell_6t
Xbit_r130_c156 bl[156] br[156] wl[130] vdd gnd cell_6t
Xbit_r131_c156 bl[156] br[156] wl[131] vdd gnd cell_6t
Xbit_r132_c156 bl[156] br[156] wl[132] vdd gnd cell_6t
Xbit_r133_c156 bl[156] br[156] wl[133] vdd gnd cell_6t
Xbit_r134_c156 bl[156] br[156] wl[134] vdd gnd cell_6t
Xbit_r135_c156 bl[156] br[156] wl[135] vdd gnd cell_6t
Xbit_r136_c156 bl[156] br[156] wl[136] vdd gnd cell_6t
Xbit_r137_c156 bl[156] br[156] wl[137] vdd gnd cell_6t
Xbit_r138_c156 bl[156] br[156] wl[138] vdd gnd cell_6t
Xbit_r139_c156 bl[156] br[156] wl[139] vdd gnd cell_6t
Xbit_r140_c156 bl[156] br[156] wl[140] vdd gnd cell_6t
Xbit_r141_c156 bl[156] br[156] wl[141] vdd gnd cell_6t
Xbit_r142_c156 bl[156] br[156] wl[142] vdd gnd cell_6t
Xbit_r143_c156 bl[156] br[156] wl[143] vdd gnd cell_6t
Xbit_r144_c156 bl[156] br[156] wl[144] vdd gnd cell_6t
Xbit_r145_c156 bl[156] br[156] wl[145] vdd gnd cell_6t
Xbit_r146_c156 bl[156] br[156] wl[146] vdd gnd cell_6t
Xbit_r147_c156 bl[156] br[156] wl[147] vdd gnd cell_6t
Xbit_r148_c156 bl[156] br[156] wl[148] vdd gnd cell_6t
Xbit_r149_c156 bl[156] br[156] wl[149] vdd gnd cell_6t
Xbit_r150_c156 bl[156] br[156] wl[150] vdd gnd cell_6t
Xbit_r151_c156 bl[156] br[156] wl[151] vdd gnd cell_6t
Xbit_r152_c156 bl[156] br[156] wl[152] vdd gnd cell_6t
Xbit_r153_c156 bl[156] br[156] wl[153] vdd gnd cell_6t
Xbit_r154_c156 bl[156] br[156] wl[154] vdd gnd cell_6t
Xbit_r155_c156 bl[156] br[156] wl[155] vdd gnd cell_6t
Xbit_r156_c156 bl[156] br[156] wl[156] vdd gnd cell_6t
Xbit_r157_c156 bl[156] br[156] wl[157] vdd gnd cell_6t
Xbit_r158_c156 bl[156] br[156] wl[158] vdd gnd cell_6t
Xbit_r159_c156 bl[156] br[156] wl[159] vdd gnd cell_6t
Xbit_r160_c156 bl[156] br[156] wl[160] vdd gnd cell_6t
Xbit_r161_c156 bl[156] br[156] wl[161] vdd gnd cell_6t
Xbit_r162_c156 bl[156] br[156] wl[162] vdd gnd cell_6t
Xbit_r163_c156 bl[156] br[156] wl[163] vdd gnd cell_6t
Xbit_r164_c156 bl[156] br[156] wl[164] vdd gnd cell_6t
Xbit_r165_c156 bl[156] br[156] wl[165] vdd gnd cell_6t
Xbit_r166_c156 bl[156] br[156] wl[166] vdd gnd cell_6t
Xbit_r167_c156 bl[156] br[156] wl[167] vdd gnd cell_6t
Xbit_r168_c156 bl[156] br[156] wl[168] vdd gnd cell_6t
Xbit_r169_c156 bl[156] br[156] wl[169] vdd gnd cell_6t
Xbit_r170_c156 bl[156] br[156] wl[170] vdd gnd cell_6t
Xbit_r171_c156 bl[156] br[156] wl[171] vdd gnd cell_6t
Xbit_r172_c156 bl[156] br[156] wl[172] vdd gnd cell_6t
Xbit_r173_c156 bl[156] br[156] wl[173] vdd gnd cell_6t
Xbit_r174_c156 bl[156] br[156] wl[174] vdd gnd cell_6t
Xbit_r175_c156 bl[156] br[156] wl[175] vdd gnd cell_6t
Xbit_r176_c156 bl[156] br[156] wl[176] vdd gnd cell_6t
Xbit_r177_c156 bl[156] br[156] wl[177] vdd gnd cell_6t
Xbit_r178_c156 bl[156] br[156] wl[178] vdd gnd cell_6t
Xbit_r179_c156 bl[156] br[156] wl[179] vdd gnd cell_6t
Xbit_r180_c156 bl[156] br[156] wl[180] vdd gnd cell_6t
Xbit_r181_c156 bl[156] br[156] wl[181] vdd gnd cell_6t
Xbit_r182_c156 bl[156] br[156] wl[182] vdd gnd cell_6t
Xbit_r183_c156 bl[156] br[156] wl[183] vdd gnd cell_6t
Xbit_r184_c156 bl[156] br[156] wl[184] vdd gnd cell_6t
Xbit_r185_c156 bl[156] br[156] wl[185] vdd gnd cell_6t
Xbit_r186_c156 bl[156] br[156] wl[186] vdd gnd cell_6t
Xbit_r187_c156 bl[156] br[156] wl[187] vdd gnd cell_6t
Xbit_r188_c156 bl[156] br[156] wl[188] vdd gnd cell_6t
Xbit_r189_c156 bl[156] br[156] wl[189] vdd gnd cell_6t
Xbit_r190_c156 bl[156] br[156] wl[190] vdd gnd cell_6t
Xbit_r191_c156 bl[156] br[156] wl[191] vdd gnd cell_6t
Xbit_r192_c156 bl[156] br[156] wl[192] vdd gnd cell_6t
Xbit_r193_c156 bl[156] br[156] wl[193] vdd gnd cell_6t
Xbit_r194_c156 bl[156] br[156] wl[194] vdd gnd cell_6t
Xbit_r195_c156 bl[156] br[156] wl[195] vdd gnd cell_6t
Xbit_r196_c156 bl[156] br[156] wl[196] vdd gnd cell_6t
Xbit_r197_c156 bl[156] br[156] wl[197] vdd gnd cell_6t
Xbit_r198_c156 bl[156] br[156] wl[198] vdd gnd cell_6t
Xbit_r199_c156 bl[156] br[156] wl[199] vdd gnd cell_6t
Xbit_r200_c156 bl[156] br[156] wl[200] vdd gnd cell_6t
Xbit_r201_c156 bl[156] br[156] wl[201] vdd gnd cell_6t
Xbit_r202_c156 bl[156] br[156] wl[202] vdd gnd cell_6t
Xbit_r203_c156 bl[156] br[156] wl[203] vdd gnd cell_6t
Xbit_r204_c156 bl[156] br[156] wl[204] vdd gnd cell_6t
Xbit_r205_c156 bl[156] br[156] wl[205] vdd gnd cell_6t
Xbit_r206_c156 bl[156] br[156] wl[206] vdd gnd cell_6t
Xbit_r207_c156 bl[156] br[156] wl[207] vdd gnd cell_6t
Xbit_r208_c156 bl[156] br[156] wl[208] vdd gnd cell_6t
Xbit_r209_c156 bl[156] br[156] wl[209] vdd gnd cell_6t
Xbit_r210_c156 bl[156] br[156] wl[210] vdd gnd cell_6t
Xbit_r211_c156 bl[156] br[156] wl[211] vdd gnd cell_6t
Xbit_r212_c156 bl[156] br[156] wl[212] vdd gnd cell_6t
Xbit_r213_c156 bl[156] br[156] wl[213] vdd gnd cell_6t
Xbit_r214_c156 bl[156] br[156] wl[214] vdd gnd cell_6t
Xbit_r215_c156 bl[156] br[156] wl[215] vdd gnd cell_6t
Xbit_r216_c156 bl[156] br[156] wl[216] vdd gnd cell_6t
Xbit_r217_c156 bl[156] br[156] wl[217] vdd gnd cell_6t
Xbit_r218_c156 bl[156] br[156] wl[218] vdd gnd cell_6t
Xbit_r219_c156 bl[156] br[156] wl[219] vdd gnd cell_6t
Xbit_r220_c156 bl[156] br[156] wl[220] vdd gnd cell_6t
Xbit_r221_c156 bl[156] br[156] wl[221] vdd gnd cell_6t
Xbit_r222_c156 bl[156] br[156] wl[222] vdd gnd cell_6t
Xbit_r223_c156 bl[156] br[156] wl[223] vdd gnd cell_6t
Xbit_r224_c156 bl[156] br[156] wl[224] vdd gnd cell_6t
Xbit_r225_c156 bl[156] br[156] wl[225] vdd gnd cell_6t
Xbit_r226_c156 bl[156] br[156] wl[226] vdd gnd cell_6t
Xbit_r227_c156 bl[156] br[156] wl[227] vdd gnd cell_6t
Xbit_r228_c156 bl[156] br[156] wl[228] vdd gnd cell_6t
Xbit_r229_c156 bl[156] br[156] wl[229] vdd gnd cell_6t
Xbit_r230_c156 bl[156] br[156] wl[230] vdd gnd cell_6t
Xbit_r231_c156 bl[156] br[156] wl[231] vdd gnd cell_6t
Xbit_r232_c156 bl[156] br[156] wl[232] vdd gnd cell_6t
Xbit_r233_c156 bl[156] br[156] wl[233] vdd gnd cell_6t
Xbit_r234_c156 bl[156] br[156] wl[234] vdd gnd cell_6t
Xbit_r235_c156 bl[156] br[156] wl[235] vdd gnd cell_6t
Xbit_r236_c156 bl[156] br[156] wl[236] vdd gnd cell_6t
Xbit_r237_c156 bl[156] br[156] wl[237] vdd gnd cell_6t
Xbit_r238_c156 bl[156] br[156] wl[238] vdd gnd cell_6t
Xbit_r239_c156 bl[156] br[156] wl[239] vdd gnd cell_6t
Xbit_r240_c156 bl[156] br[156] wl[240] vdd gnd cell_6t
Xbit_r241_c156 bl[156] br[156] wl[241] vdd gnd cell_6t
Xbit_r242_c156 bl[156] br[156] wl[242] vdd gnd cell_6t
Xbit_r243_c156 bl[156] br[156] wl[243] vdd gnd cell_6t
Xbit_r244_c156 bl[156] br[156] wl[244] vdd gnd cell_6t
Xbit_r245_c156 bl[156] br[156] wl[245] vdd gnd cell_6t
Xbit_r246_c156 bl[156] br[156] wl[246] vdd gnd cell_6t
Xbit_r247_c156 bl[156] br[156] wl[247] vdd gnd cell_6t
Xbit_r248_c156 bl[156] br[156] wl[248] vdd gnd cell_6t
Xbit_r249_c156 bl[156] br[156] wl[249] vdd gnd cell_6t
Xbit_r250_c156 bl[156] br[156] wl[250] vdd gnd cell_6t
Xbit_r251_c156 bl[156] br[156] wl[251] vdd gnd cell_6t
Xbit_r252_c156 bl[156] br[156] wl[252] vdd gnd cell_6t
Xbit_r253_c156 bl[156] br[156] wl[253] vdd gnd cell_6t
Xbit_r254_c156 bl[156] br[156] wl[254] vdd gnd cell_6t
Xbit_r255_c156 bl[156] br[156] wl[255] vdd gnd cell_6t
Xbit_r0_c157 bl[157] br[157] wl[0] vdd gnd cell_6t
Xbit_r1_c157 bl[157] br[157] wl[1] vdd gnd cell_6t
Xbit_r2_c157 bl[157] br[157] wl[2] vdd gnd cell_6t
Xbit_r3_c157 bl[157] br[157] wl[3] vdd gnd cell_6t
Xbit_r4_c157 bl[157] br[157] wl[4] vdd gnd cell_6t
Xbit_r5_c157 bl[157] br[157] wl[5] vdd gnd cell_6t
Xbit_r6_c157 bl[157] br[157] wl[6] vdd gnd cell_6t
Xbit_r7_c157 bl[157] br[157] wl[7] vdd gnd cell_6t
Xbit_r8_c157 bl[157] br[157] wl[8] vdd gnd cell_6t
Xbit_r9_c157 bl[157] br[157] wl[9] vdd gnd cell_6t
Xbit_r10_c157 bl[157] br[157] wl[10] vdd gnd cell_6t
Xbit_r11_c157 bl[157] br[157] wl[11] vdd gnd cell_6t
Xbit_r12_c157 bl[157] br[157] wl[12] vdd gnd cell_6t
Xbit_r13_c157 bl[157] br[157] wl[13] vdd gnd cell_6t
Xbit_r14_c157 bl[157] br[157] wl[14] vdd gnd cell_6t
Xbit_r15_c157 bl[157] br[157] wl[15] vdd gnd cell_6t
Xbit_r16_c157 bl[157] br[157] wl[16] vdd gnd cell_6t
Xbit_r17_c157 bl[157] br[157] wl[17] vdd gnd cell_6t
Xbit_r18_c157 bl[157] br[157] wl[18] vdd gnd cell_6t
Xbit_r19_c157 bl[157] br[157] wl[19] vdd gnd cell_6t
Xbit_r20_c157 bl[157] br[157] wl[20] vdd gnd cell_6t
Xbit_r21_c157 bl[157] br[157] wl[21] vdd gnd cell_6t
Xbit_r22_c157 bl[157] br[157] wl[22] vdd gnd cell_6t
Xbit_r23_c157 bl[157] br[157] wl[23] vdd gnd cell_6t
Xbit_r24_c157 bl[157] br[157] wl[24] vdd gnd cell_6t
Xbit_r25_c157 bl[157] br[157] wl[25] vdd gnd cell_6t
Xbit_r26_c157 bl[157] br[157] wl[26] vdd gnd cell_6t
Xbit_r27_c157 bl[157] br[157] wl[27] vdd gnd cell_6t
Xbit_r28_c157 bl[157] br[157] wl[28] vdd gnd cell_6t
Xbit_r29_c157 bl[157] br[157] wl[29] vdd gnd cell_6t
Xbit_r30_c157 bl[157] br[157] wl[30] vdd gnd cell_6t
Xbit_r31_c157 bl[157] br[157] wl[31] vdd gnd cell_6t
Xbit_r32_c157 bl[157] br[157] wl[32] vdd gnd cell_6t
Xbit_r33_c157 bl[157] br[157] wl[33] vdd gnd cell_6t
Xbit_r34_c157 bl[157] br[157] wl[34] vdd gnd cell_6t
Xbit_r35_c157 bl[157] br[157] wl[35] vdd gnd cell_6t
Xbit_r36_c157 bl[157] br[157] wl[36] vdd gnd cell_6t
Xbit_r37_c157 bl[157] br[157] wl[37] vdd gnd cell_6t
Xbit_r38_c157 bl[157] br[157] wl[38] vdd gnd cell_6t
Xbit_r39_c157 bl[157] br[157] wl[39] vdd gnd cell_6t
Xbit_r40_c157 bl[157] br[157] wl[40] vdd gnd cell_6t
Xbit_r41_c157 bl[157] br[157] wl[41] vdd gnd cell_6t
Xbit_r42_c157 bl[157] br[157] wl[42] vdd gnd cell_6t
Xbit_r43_c157 bl[157] br[157] wl[43] vdd gnd cell_6t
Xbit_r44_c157 bl[157] br[157] wl[44] vdd gnd cell_6t
Xbit_r45_c157 bl[157] br[157] wl[45] vdd gnd cell_6t
Xbit_r46_c157 bl[157] br[157] wl[46] vdd gnd cell_6t
Xbit_r47_c157 bl[157] br[157] wl[47] vdd gnd cell_6t
Xbit_r48_c157 bl[157] br[157] wl[48] vdd gnd cell_6t
Xbit_r49_c157 bl[157] br[157] wl[49] vdd gnd cell_6t
Xbit_r50_c157 bl[157] br[157] wl[50] vdd gnd cell_6t
Xbit_r51_c157 bl[157] br[157] wl[51] vdd gnd cell_6t
Xbit_r52_c157 bl[157] br[157] wl[52] vdd gnd cell_6t
Xbit_r53_c157 bl[157] br[157] wl[53] vdd gnd cell_6t
Xbit_r54_c157 bl[157] br[157] wl[54] vdd gnd cell_6t
Xbit_r55_c157 bl[157] br[157] wl[55] vdd gnd cell_6t
Xbit_r56_c157 bl[157] br[157] wl[56] vdd gnd cell_6t
Xbit_r57_c157 bl[157] br[157] wl[57] vdd gnd cell_6t
Xbit_r58_c157 bl[157] br[157] wl[58] vdd gnd cell_6t
Xbit_r59_c157 bl[157] br[157] wl[59] vdd gnd cell_6t
Xbit_r60_c157 bl[157] br[157] wl[60] vdd gnd cell_6t
Xbit_r61_c157 bl[157] br[157] wl[61] vdd gnd cell_6t
Xbit_r62_c157 bl[157] br[157] wl[62] vdd gnd cell_6t
Xbit_r63_c157 bl[157] br[157] wl[63] vdd gnd cell_6t
Xbit_r64_c157 bl[157] br[157] wl[64] vdd gnd cell_6t
Xbit_r65_c157 bl[157] br[157] wl[65] vdd gnd cell_6t
Xbit_r66_c157 bl[157] br[157] wl[66] vdd gnd cell_6t
Xbit_r67_c157 bl[157] br[157] wl[67] vdd gnd cell_6t
Xbit_r68_c157 bl[157] br[157] wl[68] vdd gnd cell_6t
Xbit_r69_c157 bl[157] br[157] wl[69] vdd gnd cell_6t
Xbit_r70_c157 bl[157] br[157] wl[70] vdd gnd cell_6t
Xbit_r71_c157 bl[157] br[157] wl[71] vdd gnd cell_6t
Xbit_r72_c157 bl[157] br[157] wl[72] vdd gnd cell_6t
Xbit_r73_c157 bl[157] br[157] wl[73] vdd gnd cell_6t
Xbit_r74_c157 bl[157] br[157] wl[74] vdd gnd cell_6t
Xbit_r75_c157 bl[157] br[157] wl[75] vdd gnd cell_6t
Xbit_r76_c157 bl[157] br[157] wl[76] vdd gnd cell_6t
Xbit_r77_c157 bl[157] br[157] wl[77] vdd gnd cell_6t
Xbit_r78_c157 bl[157] br[157] wl[78] vdd gnd cell_6t
Xbit_r79_c157 bl[157] br[157] wl[79] vdd gnd cell_6t
Xbit_r80_c157 bl[157] br[157] wl[80] vdd gnd cell_6t
Xbit_r81_c157 bl[157] br[157] wl[81] vdd gnd cell_6t
Xbit_r82_c157 bl[157] br[157] wl[82] vdd gnd cell_6t
Xbit_r83_c157 bl[157] br[157] wl[83] vdd gnd cell_6t
Xbit_r84_c157 bl[157] br[157] wl[84] vdd gnd cell_6t
Xbit_r85_c157 bl[157] br[157] wl[85] vdd gnd cell_6t
Xbit_r86_c157 bl[157] br[157] wl[86] vdd gnd cell_6t
Xbit_r87_c157 bl[157] br[157] wl[87] vdd gnd cell_6t
Xbit_r88_c157 bl[157] br[157] wl[88] vdd gnd cell_6t
Xbit_r89_c157 bl[157] br[157] wl[89] vdd gnd cell_6t
Xbit_r90_c157 bl[157] br[157] wl[90] vdd gnd cell_6t
Xbit_r91_c157 bl[157] br[157] wl[91] vdd gnd cell_6t
Xbit_r92_c157 bl[157] br[157] wl[92] vdd gnd cell_6t
Xbit_r93_c157 bl[157] br[157] wl[93] vdd gnd cell_6t
Xbit_r94_c157 bl[157] br[157] wl[94] vdd gnd cell_6t
Xbit_r95_c157 bl[157] br[157] wl[95] vdd gnd cell_6t
Xbit_r96_c157 bl[157] br[157] wl[96] vdd gnd cell_6t
Xbit_r97_c157 bl[157] br[157] wl[97] vdd gnd cell_6t
Xbit_r98_c157 bl[157] br[157] wl[98] vdd gnd cell_6t
Xbit_r99_c157 bl[157] br[157] wl[99] vdd gnd cell_6t
Xbit_r100_c157 bl[157] br[157] wl[100] vdd gnd cell_6t
Xbit_r101_c157 bl[157] br[157] wl[101] vdd gnd cell_6t
Xbit_r102_c157 bl[157] br[157] wl[102] vdd gnd cell_6t
Xbit_r103_c157 bl[157] br[157] wl[103] vdd gnd cell_6t
Xbit_r104_c157 bl[157] br[157] wl[104] vdd gnd cell_6t
Xbit_r105_c157 bl[157] br[157] wl[105] vdd gnd cell_6t
Xbit_r106_c157 bl[157] br[157] wl[106] vdd gnd cell_6t
Xbit_r107_c157 bl[157] br[157] wl[107] vdd gnd cell_6t
Xbit_r108_c157 bl[157] br[157] wl[108] vdd gnd cell_6t
Xbit_r109_c157 bl[157] br[157] wl[109] vdd gnd cell_6t
Xbit_r110_c157 bl[157] br[157] wl[110] vdd gnd cell_6t
Xbit_r111_c157 bl[157] br[157] wl[111] vdd gnd cell_6t
Xbit_r112_c157 bl[157] br[157] wl[112] vdd gnd cell_6t
Xbit_r113_c157 bl[157] br[157] wl[113] vdd gnd cell_6t
Xbit_r114_c157 bl[157] br[157] wl[114] vdd gnd cell_6t
Xbit_r115_c157 bl[157] br[157] wl[115] vdd gnd cell_6t
Xbit_r116_c157 bl[157] br[157] wl[116] vdd gnd cell_6t
Xbit_r117_c157 bl[157] br[157] wl[117] vdd gnd cell_6t
Xbit_r118_c157 bl[157] br[157] wl[118] vdd gnd cell_6t
Xbit_r119_c157 bl[157] br[157] wl[119] vdd gnd cell_6t
Xbit_r120_c157 bl[157] br[157] wl[120] vdd gnd cell_6t
Xbit_r121_c157 bl[157] br[157] wl[121] vdd gnd cell_6t
Xbit_r122_c157 bl[157] br[157] wl[122] vdd gnd cell_6t
Xbit_r123_c157 bl[157] br[157] wl[123] vdd gnd cell_6t
Xbit_r124_c157 bl[157] br[157] wl[124] vdd gnd cell_6t
Xbit_r125_c157 bl[157] br[157] wl[125] vdd gnd cell_6t
Xbit_r126_c157 bl[157] br[157] wl[126] vdd gnd cell_6t
Xbit_r127_c157 bl[157] br[157] wl[127] vdd gnd cell_6t
Xbit_r128_c157 bl[157] br[157] wl[128] vdd gnd cell_6t
Xbit_r129_c157 bl[157] br[157] wl[129] vdd gnd cell_6t
Xbit_r130_c157 bl[157] br[157] wl[130] vdd gnd cell_6t
Xbit_r131_c157 bl[157] br[157] wl[131] vdd gnd cell_6t
Xbit_r132_c157 bl[157] br[157] wl[132] vdd gnd cell_6t
Xbit_r133_c157 bl[157] br[157] wl[133] vdd gnd cell_6t
Xbit_r134_c157 bl[157] br[157] wl[134] vdd gnd cell_6t
Xbit_r135_c157 bl[157] br[157] wl[135] vdd gnd cell_6t
Xbit_r136_c157 bl[157] br[157] wl[136] vdd gnd cell_6t
Xbit_r137_c157 bl[157] br[157] wl[137] vdd gnd cell_6t
Xbit_r138_c157 bl[157] br[157] wl[138] vdd gnd cell_6t
Xbit_r139_c157 bl[157] br[157] wl[139] vdd gnd cell_6t
Xbit_r140_c157 bl[157] br[157] wl[140] vdd gnd cell_6t
Xbit_r141_c157 bl[157] br[157] wl[141] vdd gnd cell_6t
Xbit_r142_c157 bl[157] br[157] wl[142] vdd gnd cell_6t
Xbit_r143_c157 bl[157] br[157] wl[143] vdd gnd cell_6t
Xbit_r144_c157 bl[157] br[157] wl[144] vdd gnd cell_6t
Xbit_r145_c157 bl[157] br[157] wl[145] vdd gnd cell_6t
Xbit_r146_c157 bl[157] br[157] wl[146] vdd gnd cell_6t
Xbit_r147_c157 bl[157] br[157] wl[147] vdd gnd cell_6t
Xbit_r148_c157 bl[157] br[157] wl[148] vdd gnd cell_6t
Xbit_r149_c157 bl[157] br[157] wl[149] vdd gnd cell_6t
Xbit_r150_c157 bl[157] br[157] wl[150] vdd gnd cell_6t
Xbit_r151_c157 bl[157] br[157] wl[151] vdd gnd cell_6t
Xbit_r152_c157 bl[157] br[157] wl[152] vdd gnd cell_6t
Xbit_r153_c157 bl[157] br[157] wl[153] vdd gnd cell_6t
Xbit_r154_c157 bl[157] br[157] wl[154] vdd gnd cell_6t
Xbit_r155_c157 bl[157] br[157] wl[155] vdd gnd cell_6t
Xbit_r156_c157 bl[157] br[157] wl[156] vdd gnd cell_6t
Xbit_r157_c157 bl[157] br[157] wl[157] vdd gnd cell_6t
Xbit_r158_c157 bl[157] br[157] wl[158] vdd gnd cell_6t
Xbit_r159_c157 bl[157] br[157] wl[159] vdd gnd cell_6t
Xbit_r160_c157 bl[157] br[157] wl[160] vdd gnd cell_6t
Xbit_r161_c157 bl[157] br[157] wl[161] vdd gnd cell_6t
Xbit_r162_c157 bl[157] br[157] wl[162] vdd gnd cell_6t
Xbit_r163_c157 bl[157] br[157] wl[163] vdd gnd cell_6t
Xbit_r164_c157 bl[157] br[157] wl[164] vdd gnd cell_6t
Xbit_r165_c157 bl[157] br[157] wl[165] vdd gnd cell_6t
Xbit_r166_c157 bl[157] br[157] wl[166] vdd gnd cell_6t
Xbit_r167_c157 bl[157] br[157] wl[167] vdd gnd cell_6t
Xbit_r168_c157 bl[157] br[157] wl[168] vdd gnd cell_6t
Xbit_r169_c157 bl[157] br[157] wl[169] vdd gnd cell_6t
Xbit_r170_c157 bl[157] br[157] wl[170] vdd gnd cell_6t
Xbit_r171_c157 bl[157] br[157] wl[171] vdd gnd cell_6t
Xbit_r172_c157 bl[157] br[157] wl[172] vdd gnd cell_6t
Xbit_r173_c157 bl[157] br[157] wl[173] vdd gnd cell_6t
Xbit_r174_c157 bl[157] br[157] wl[174] vdd gnd cell_6t
Xbit_r175_c157 bl[157] br[157] wl[175] vdd gnd cell_6t
Xbit_r176_c157 bl[157] br[157] wl[176] vdd gnd cell_6t
Xbit_r177_c157 bl[157] br[157] wl[177] vdd gnd cell_6t
Xbit_r178_c157 bl[157] br[157] wl[178] vdd gnd cell_6t
Xbit_r179_c157 bl[157] br[157] wl[179] vdd gnd cell_6t
Xbit_r180_c157 bl[157] br[157] wl[180] vdd gnd cell_6t
Xbit_r181_c157 bl[157] br[157] wl[181] vdd gnd cell_6t
Xbit_r182_c157 bl[157] br[157] wl[182] vdd gnd cell_6t
Xbit_r183_c157 bl[157] br[157] wl[183] vdd gnd cell_6t
Xbit_r184_c157 bl[157] br[157] wl[184] vdd gnd cell_6t
Xbit_r185_c157 bl[157] br[157] wl[185] vdd gnd cell_6t
Xbit_r186_c157 bl[157] br[157] wl[186] vdd gnd cell_6t
Xbit_r187_c157 bl[157] br[157] wl[187] vdd gnd cell_6t
Xbit_r188_c157 bl[157] br[157] wl[188] vdd gnd cell_6t
Xbit_r189_c157 bl[157] br[157] wl[189] vdd gnd cell_6t
Xbit_r190_c157 bl[157] br[157] wl[190] vdd gnd cell_6t
Xbit_r191_c157 bl[157] br[157] wl[191] vdd gnd cell_6t
Xbit_r192_c157 bl[157] br[157] wl[192] vdd gnd cell_6t
Xbit_r193_c157 bl[157] br[157] wl[193] vdd gnd cell_6t
Xbit_r194_c157 bl[157] br[157] wl[194] vdd gnd cell_6t
Xbit_r195_c157 bl[157] br[157] wl[195] vdd gnd cell_6t
Xbit_r196_c157 bl[157] br[157] wl[196] vdd gnd cell_6t
Xbit_r197_c157 bl[157] br[157] wl[197] vdd gnd cell_6t
Xbit_r198_c157 bl[157] br[157] wl[198] vdd gnd cell_6t
Xbit_r199_c157 bl[157] br[157] wl[199] vdd gnd cell_6t
Xbit_r200_c157 bl[157] br[157] wl[200] vdd gnd cell_6t
Xbit_r201_c157 bl[157] br[157] wl[201] vdd gnd cell_6t
Xbit_r202_c157 bl[157] br[157] wl[202] vdd gnd cell_6t
Xbit_r203_c157 bl[157] br[157] wl[203] vdd gnd cell_6t
Xbit_r204_c157 bl[157] br[157] wl[204] vdd gnd cell_6t
Xbit_r205_c157 bl[157] br[157] wl[205] vdd gnd cell_6t
Xbit_r206_c157 bl[157] br[157] wl[206] vdd gnd cell_6t
Xbit_r207_c157 bl[157] br[157] wl[207] vdd gnd cell_6t
Xbit_r208_c157 bl[157] br[157] wl[208] vdd gnd cell_6t
Xbit_r209_c157 bl[157] br[157] wl[209] vdd gnd cell_6t
Xbit_r210_c157 bl[157] br[157] wl[210] vdd gnd cell_6t
Xbit_r211_c157 bl[157] br[157] wl[211] vdd gnd cell_6t
Xbit_r212_c157 bl[157] br[157] wl[212] vdd gnd cell_6t
Xbit_r213_c157 bl[157] br[157] wl[213] vdd gnd cell_6t
Xbit_r214_c157 bl[157] br[157] wl[214] vdd gnd cell_6t
Xbit_r215_c157 bl[157] br[157] wl[215] vdd gnd cell_6t
Xbit_r216_c157 bl[157] br[157] wl[216] vdd gnd cell_6t
Xbit_r217_c157 bl[157] br[157] wl[217] vdd gnd cell_6t
Xbit_r218_c157 bl[157] br[157] wl[218] vdd gnd cell_6t
Xbit_r219_c157 bl[157] br[157] wl[219] vdd gnd cell_6t
Xbit_r220_c157 bl[157] br[157] wl[220] vdd gnd cell_6t
Xbit_r221_c157 bl[157] br[157] wl[221] vdd gnd cell_6t
Xbit_r222_c157 bl[157] br[157] wl[222] vdd gnd cell_6t
Xbit_r223_c157 bl[157] br[157] wl[223] vdd gnd cell_6t
Xbit_r224_c157 bl[157] br[157] wl[224] vdd gnd cell_6t
Xbit_r225_c157 bl[157] br[157] wl[225] vdd gnd cell_6t
Xbit_r226_c157 bl[157] br[157] wl[226] vdd gnd cell_6t
Xbit_r227_c157 bl[157] br[157] wl[227] vdd gnd cell_6t
Xbit_r228_c157 bl[157] br[157] wl[228] vdd gnd cell_6t
Xbit_r229_c157 bl[157] br[157] wl[229] vdd gnd cell_6t
Xbit_r230_c157 bl[157] br[157] wl[230] vdd gnd cell_6t
Xbit_r231_c157 bl[157] br[157] wl[231] vdd gnd cell_6t
Xbit_r232_c157 bl[157] br[157] wl[232] vdd gnd cell_6t
Xbit_r233_c157 bl[157] br[157] wl[233] vdd gnd cell_6t
Xbit_r234_c157 bl[157] br[157] wl[234] vdd gnd cell_6t
Xbit_r235_c157 bl[157] br[157] wl[235] vdd gnd cell_6t
Xbit_r236_c157 bl[157] br[157] wl[236] vdd gnd cell_6t
Xbit_r237_c157 bl[157] br[157] wl[237] vdd gnd cell_6t
Xbit_r238_c157 bl[157] br[157] wl[238] vdd gnd cell_6t
Xbit_r239_c157 bl[157] br[157] wl[239] vdd gnd cell_6t
Xbit_r240_c157 bl[157] br[157] wl[240] vdd gnd cell_6t
Xbit_r241_c157 bl[157] br[157] wl[241] vdd gnd cell_6t
Xbit_r242_c157 bl[157] br[157] wl[242] vdd gnd cell_6t
Xbit_r243_c157 bl[157] br[157] wl[243] vdd gnd cell_6t
Xbit_r244_c157 bl[157] br[157] wl[244] vdd gnd cell_6t
Xbit_r245_c157 bl[157] br[157] wl[245] vdd gnd cell_6t
Xbit_r246_c157 bl[157] br[157] wl[246] vdd gnd cell_6t
Xbit_r247_c157 bl[157] br[157] wl[247] vdd gnd cell_6t
Xbit_r248_c157 bl[157] br[157] wl[248] vdd gnd cell_6t
Xbit_r249_c157 bl[157] br[157] wl[249] vdd gnd cell_6t
Xbit_r250_c157 bl[157] br[157] wl[250] vdd gnd cell_6t
Xbit_r251_c157 bl[157] br[157] wl[251] vdd gnd cell_6t
Xbit_r252_c157 bl[157] br[157] wl[252] vdd gnd cell_6t
Xbit_r253_c157 bl[157] br[157] wl[253] vdd gnd cell_6t
Xbit_r254_c157 bl[157] br[157] wl[254] vdd gnd cell_6t
Xbit_r255_c157 bl[157] br[157] wl[255] vdd gnd cell_6t
Xbit_r0_c158 bl[158] br[158] wl[0] vdd gnd cell_6t
Xbit_r1_c158 bl[158] br[158] wl[1] vdd gnd cell_6t
Xbit_r2_c158 bl[158] br[158] wl[2] vdd gnd cell_6t
Xbit_r3_c158 bl[158] br[158] wl[3] vdd gnd cell_6t
Xbit_r4_c158 bl[158] br[158] wl[4] vdd gnd cell_6t
Xbit_r5_c158 bl[158] br[158] wl[5] vdd gnd cell_6t
Xbit_r6_c158 bl[158] br[158] wl[6] vdd gnd cell_6t
Xbit_r7_c158 bl[158] br[158] wl[7] vdd gnd cell_6t
Xbit_r8_c158 bl[158] br[158] wl[8] vdd gnd cell_6t
Xbit_r9_c158 bl[158] br[158] wl[9] vdd gnd cell_6t
Xbit_r10_c158 bl[158] br[158] wl[10] vdd gnd cell_6t
Xbit_r11_c158 bl[158] br[158] wl[11] vdd gnd cell_6t
Xbit_r12_c158 bl[158] br[158] wl[12] vdd gnd cell_6t
Xbit_r13_c158 bl[158] br[158] wl[13] vdd gnd cell_6t
Xbit_r14_c158 bl[158] br[158] wl[14] vdd gnd cell_6t
Xbit_r15_c158 bl[158] br[158] wl[15] vdd gnd cell_6t
Xbit_r16_c158 bl[158] br[158] wl[16] vdd gnd cell_6t
Xbit_r17_c158 bl[158] br[158] wl[17] vdd gnd cell_6t
Xbit_r18_c158 bl[158] br[158] wl[18] vdd gnd cell_6t
Xbit_r19_c158 bl[158] br[158] wl[19] vdd gnd cell_6t
Xbit_r20_c158 bl[158] br[158] wl[20] vdd gnd cell_6t
Xbit_r21_c158 bl[158] br[158] wl[21] vdd gnd cell_6t
Xbit_r22_c158 bl[158] br[158] wl[22] vdd gnd cell_6t
Xbit_r23_c158 bl[158] br[158] wl[23] vdd gnd cell_6t
Xbit_r24_c158 bl[158] br[158] wl[24] vdd gnd cell_6t
Xbit_r25_c158 bl[158] br[158] wl[25] vdd gnd cell_6t
Xbit_r26_c158 bl[158] br[158] wl[26] vdd gnd cell_6t
Xbit_r27_c158 bl[158] br[158] wl[27] vdd gnd cell_6t
Xbit_r28_c158 bl[158] br[158] wl[28] vdd gnd cell_6t
Xbit_r29_c158 bl[158] br[158] wl[29] vdd gnd cell_6t
Xbit_r30_c158 bl[158] br[158] wl[30] vdd gnd cell_6t
Xbit_r31_c158 bl[158] br[158] wl[31] vdd gnd cell_6t
Xbit_r32_c158 bl[158] br[158] wl[32] vdd gnd cell_6t
Xbit_r33_c158 bl[158] br[158] wl[33] vdd gnd cell_6t
Xbit_r34_c158 bl[158] br[158] wl[34] vdd gnd cell_6t
Xbit_r35_c158 bl[158] br[158] wl[35] vdd gnd cell_6t
Xbit_r36_c158 bl[158] br[158] wl[36] vdd gnd cell_6t
Xbit_r37_c158 bl[158] br[158] wl[37] vdd gnd cell_6t
Xbit_r38_c158 bl[158] br[158] wl[38] vdd gnd cell_6t
Xbit_r39_c158 bl[158] br[158] wl[39] vdd gnd cell_6t
Xbit_r40_c158 bl[158] br[158] wl[40] vdd gnd cell_6t
Xbit_r41_c158 bl[158] br[158] wl[41] vdd gnd cell_6t
Xbit_r42_c158 bl[158] br[158] wl[42] vdd gnd cell_6t
Xbit_r43_c158 bl[158] br[158] wl[43] vdd gnd cell_6t
Xbit_r44_c158 bl[158] br[158] wl[44] vdd gnd cell_6t
Xbit_r45_c158 bl[158] br[158] wl[45] vdd gnd cell_6t
Xbit_r46_c158 bl[158] br[158] wl[46] vdd gnd cell_6t
Xbit_r47_c158 bl[158] br[158] wl[47] vdd gnd cell_6t
Xbit_r48_c158 bl[158] br[158] wl[48] vdd gnd cell_6t
Xbit_r49_c158 bl[158] br[158] wl[49] vdd gnd cell_6t
Xbit_r50_c158 bl[158] br[158] wl[50] vdd gnd cell_6t
Xbit_r51_c158 bl[158] br[158] wl[51] vdd gnd cell_6t
Xbit_r52_c158 bl[158] br[158] wl[52] vdd gnd cell_6t
Xbit_r53_c158 bl[158] br[158] wl[53] vdd gnd cell_6t
Xbit_r54_c158 bl[158] br[158] wl[54] vdd gnd cell_6t
Xbit_r55_c158 bl[158] br[158] wl[55] vdd gnd cell_6t
Xbit_r56_c158 bl[158] br[158] wl[56] vdd gnd cell_6t
Xbit_r57_c158 bl[158] br[158] wl[57] vdd gnd cell_6t
Xbit_r58_c158 bl[158] br[158] wl[58] vdd gnd cell_6t
Xbit_r59_c158 bl[158] br[158] wl[59] vdd gnd cell_6t
Xbit_r60_c158 bl[158] br[158] wl[60] vdd gnd cell_6t
Xbit_r61_c158 bl[158] br[158] wl[61] vdd gnd cell_6t
Xbit_r62_c158 bl[158] br[158] wl[62] vdd gnd cell_6t
Xbit_r63_c158 bl[158] br[158] wl[63] vdd gnd cell_6t
Xbit_r64_c158 bl[158] br[158] wl[64] vdd gnd cell_6t
Xbit_r65_c158 bl[158] br[158] wl[65] vdd gnd cell_6t
Xbit_r66_c158 bl[158] br[158] wl[66] vdd gnd cell_6t
Xbit_r67_c158 bl[158] br[158] wl[67] vdd gnd cell_6t
Xbit_r68_c158 bl[158] br[158] wl[68] vdd gnd cell_6t
Xbit_r69_c158 bl[158] br[158] wl[69] vdd gnd cell_6t
Xbit_r70_c158 bl[158] br[158] wl[70] vdd gnd cell_6t
Xbit_r71_c158 bl[158] br[158] wl[71] vdd gnd cell_6t
Xbit_r72_c158 bl[158] br[158] wl[72] vdd gnd cell_6t
Xbit_r73_c158 bl[158] br[158] wl[73] vdd gnd cell_6t
Xbit_r74_c158 bl[158] br[158] wl[74] vdd gnd cell_6t
Xbit_r75_c158 bl[158] br[158] wl[75] vdd gnd cell_6t
Xbit_r76_c158 bl[158] br[158] wl[76] vdd gnd cell_6t
Xbit_r77_c158 bl[158] br[158] wl[77] vdd gnd cell_6t
Xbit_r78_c158 bl[158] br[158] wl[78] vdd gnd cell_6t
Xbit_r79_c158 bl[158] br[158] wl[79] vdd gnd cell_6t
Xbit_r80_c158 bl[158] br[158] wl[80] vdd gnd cell_6t
Xbit_r81_c158 bl[158] br[158] wl[81] vdd gnd cell_6t
Xbit_r82_c158 bl[158] br[158] wl[82] vdd gnd cell_6t
Xbit_r83_c158 bl[158] br[158] wl[83] vdd gnd cell_6t
Xbit_r84_c158 bl[158] br[158] wl[84] vdd gnd cell_6t
Xbit_r85_c158 bl[158] br[158] wl[85] vdd gnd cell_6t
Xbit_r86_c158 bl[158] br[158] wl[86] vdd gnd cell_6t
Xbit_r87_c158 bl[158] br[158] wl[87] vdd gnd cell_6t
Xbit_r88_c158 bl[158] br[158] wl[88] vdd gnd cell_6t
Xbit_r89_c158 bl[158] br[158] wl[89] vdd gnd cell_6t
Xbit_r90_c158 bl[158] br[158] wl[90] vdd gnd cell_6t
Xbit_r91_c158 bl[158] br[158] wl[91] vdd gnd cell_6t
Xbit_r92_c158 bl[158] br[158] wl[92] vdd gnd cell_6t
Xbit_r93_c158 bl[158] br[158] wl[93] vdd gnd cell_6t
Xbit_r94_c158 bl[158] br[158] wl[94] vdd gnd cell_6t
Xbit_r95_c158 bl[158] br[158] wl[95] vdd gnd cell_6t
Xbit_r96_c158 bl[158] br[158] wl[96] vdd gnd cell_6t
Xbit_r97_c158 bl[158] br[158] wl[97] vdd gnd cell_6t
Xbit_r98_c158 bl[158] br[158] wl[98] vdd gnd cell_6t
Xbit_r99_c158 bl[158] br[158] wl[99] vdd gnd cell_6t
Xbit_r100_c158 bl[158] br[158] wl[100] vdd gnd cell_6t
Xbit_r101_c158 bl[158] br[158] wl[101] vdd gnd cell_6t
Xbit_r102_c158 bl[158] br[158] wl[102] vdd gnd cell_6t
Xbit_r103_c158 bl[158] br[158] wl[103] vdd gnd cell_6t
Xbit_r104_c158 bl[158] br[158] wl[104] vdd gnd cell_6t
Xbit_r105_c158 bl[158] br[158] wl[105] vdd gnd cell_6t
Xbit_r106_c158 bl[158] br[158] wl[106] vdd gnd cell_6t
Xbit_r107_c158 bl[158] br[158] wl[107] vdd gnd cell_6t
Xbit_r108_c158 bl[158] br[158] wl[108] vdd gnd cell_6t
Xbit_r109_c158 bl[158] br[158] wl[109] vdd gnd cell_6t
Xbit_r110_c158 bl[158] br[158] wl[110] vdd gnd cell_6t
Xbit_r111_c158 bl[158] br[158] wl[111] vdd gnd cell_6t
Xbit_r112_c158 bl[158] br[158] wl[112] vdd gnd cell_6t
Xbit_r113_c158 bl[158] br[158] wl[113] vdd gnd cell_6t
Xbit_r114_c158 bl[158] br[158] wl[114] vdd gnd cell_6t
Xbit_r115_c158 bl[158] br[158] wl[115] vdd gnd cell_6t
Xbit_r116_c158 bl[158] br[158] wl[116] vdd gnd cell_6t
Xbit_r117_c158 bl[158] br[158] wl[117] vdd gnd cell_6t
Xbit_r118_c158 bl[158] br[158] wl[118] vdd gnd cell_6t
Xbit_r119_c158 bl[158] br[158] wl[119] vdd gnd cell_6t
Xbit_r120_c158 bl[158] br[158] wl[120] vdd gnd cell_6t
Xbit_r121_c158 bl[158] br[158] wl[121] vdd gnd cell_6t
Xbit_r122_c158 bl[158] br[158] wl[122] vdd gnd cell_6t
Xbit_r123_c158 bl[158] br[158] wl[123] vdd gnd cell_6t
Xbit_r124_c158 bl[158] br[158] wl[124] vdd gnd cell_6t
Xbit_r125_c158 bl[158] br[158] wl[125] vdd gnd cell_6t
Xbit_r126_c158 bl[158] br[158] wl[126] vdd gnd cell_6t
Xbit_r127_c158 bl[158] br[158] wl[127] vdd gnd cell_6t
Xbit_r128_c158 bl[158] br[158] wl[128] vdd gnd cell_6t
Xbit_r129_c158 bl[158] br[158] wl[129] vdd gnd cell_6t
Xbit_r130_c158 bl[158] br[158] wl[130] vdd gnd cell_6t
Xbit_r131_c158 bl[158] br[158] wl[131] vdd gnd cell_6t
Xbit_r132_c158 bl[158] br[158] wl[132] vdd gnd cell_6t
Xbit_r133_c158 bl[158] br[158] wl[133] vdd gnd cell_6t
Xbit_r134_c158 bl[158] br[158] wl[134] vdd gnd cell_6t
Xbit_r135_c158 bl[158] br[158] wl[135] vdd gnd cell_6t
Xbit_r136_c158 bl[158] br[158] wl[136] vdd gnd cell_6t
Xbit_r137_c158 bl[158] br[158] wl[137] vdd gnd cell_6t
Xbit_r138_c158 bl[158] br[158] wl[138] vdd gnd cell_6t
Xbit_r139_c158 bl[158] br[158] wl[139] vdd gnd cell_6t
Xbit_r140_c158 bl[158] br[158] wl[140] vdd gnd cell_6t
Xbit_r141_c158 bl[158] br[158] wl[141] vdd gnd cell_6t
Xbit_r142_c158 bl[158] br[158] wl[142] vdd gnd cell_6t
Xbit_r143_c158 bl[158] br[158] wl[143] vdd gnd cell_6t
Xbit_r144_c158 bl[158] br[158] wl[144] vdd gnd cell_6t
Xbit_r145_c158 bl[158] br[158] wl[145] vdd gnd cell_6t
Xbit_r146_c158 bl[158] br[158] wl[146] vdd gnd cell_6t
Xbit_r147_c158 bl[158] br[158] wl[147] vdd gnd cell_6t
Xbit_r148_c158 bl[158] br[158] wl[148] vdd gnd cell_6t
Xbit_r149_c158 bl[158] br[158] wl[149] vdd gnd cell_6t
Xbit_r150_c158 bl[158] br[158] wl[150] vdd gnd cell_6t
Xbit_r151_c158 bl[158] br[158] wl[151] vdd gnd cell_6t
Xbit_r152_c158 bl[158] br[158] wl[152] vdd gnd cell_6t
Xbit_r153_c158 bl[158] br[158] wl[153] vdd gnd cell_6t
Xbit_r154_c158 bl[158] br[158] wl[154] vdd gnd cell_6t
Xbit_r155_c158 bl[158] br[158] wl[155] vdd gnd cell_6t
Xbit_r156_c158 bl[158] br[158] wl[156] vdd gnd cell_6t
Xbit_r157_c158 bl[158] br[158] wl[157] vdd gnd cell_6t
Xbit_r158_c158 bl[158] br[158] wl[158] vdd gnd cell_6t
Xbit_r159_c158 bl[158] br[158] wl[159] vdd gnd cell_6t
Xbit_r160_c158 bl[158] br[158] wl[160] vdd gnd cell_6t
Xbit_r161_c158 bl[158] br[158] wl[161] vdd gnd cell_6t
Xbit_r162_c158 bl[158] br[158] wl[162] vdd gnd cell_6t
Xbit_r163_c158 bl[158] br[158] wl[163] vdd gnd cell_6t
Xbit_r164_c158 bl[158] br[158] wl[164] vdd gnd cell_6t
Xbit_r165_c158 bl[158] br[158] wl[165] vdd gnd cell_6t
Xbit_r166_c158 bl[158] br[158] wl[166] vdd gnd cell_6t
Xbit_r167_c158 bl[158] br[158] wl[167] vdd gnd cell_6t
Xbit_r168_c158 bl[158] br[158] wl[168] vdd gnd cell_6t
Xbit_r169_c158 bl[158] br[158] wl[169] vdd gnd cell_6t
Xbit_r170_c158 bl[158] br[158] wl[170] vdd gnd cell_6t
Xbit_r171_c158 bl[158] br[158] wl[171] vdd gnd cell_6t
Xbit_r172_c158 bl[158] br[158] wl[172] vdd gnd cell_6t
Xbit_r173_c158 bl[158] br[158] wl[173] vdd gnd cell_6t
Xbit_r174_c158 bl[158] br[158] wl[174] vdd gnd cell_6t
Xbit_r175_c158 bl[158] br[158] wl[175] vdd gnd cell_6t
Xbit_r176_c158 bl[158] br[158] wl[176] vdd gnd cell_6t
Xbit_r177_c158 bl[158] br[158] wl[177] vdd gnd cell_6t
Xbit_r178_c158 bl[158] br[158] wl[178] vdd gnd cell_6t
Xbit_r179_c158 bl[158] br[158] wl[179] vdd gnd cell_6t
Xbit_r180_c158 bl[158] br[158] wl[180] vdd gnd cell_6t
Xbit_r181_c158 bl[158] br[158] wl[181] vdd gnd cell_6t
Xbit_r182_c158 bl[158] br[158] wl[182] vdd gnd cell_6t
Xbit_r183_c158 bl[158] br[158] wl[183] vdd gnd cell_6t
Xbit_r184_c158 bl[158] br[158] wl[184] vdd gnd cell_6t
Xbit_r185_c158 bl[158] br[158] wl[185] vdd gnd cell_6t
Xbit_r186_c158 bl[158] br[158] wl[186] vdd gnd cell_6t
Xbit_r187_c158 bl[158] br[158] wl[187] vdd gnd cell_6t
Xbit_r188_c158 bl[158] br[158] wl[188] vdd gnd cell_6t
Xbit_r189_c158 bl[158] br[158] wl[189] vdd gnd cell_6t
Xbit_r190_c158 bl[158] br[158] wl[190] vdd gnd cell_6t
Xbit_r191_c158 bl[158] br[158] wl[191] vdd gnd cell_6t
Xbit_r192_c158 bl[158] br[158] wl[192] vdd gnd cell_6t
Xbit_r193_c158 bl[158] br[158] wl[193] vdd gnd cell_6t
Xbit_r194_c158 bl[158] br[158] wl[194] vdd gnd cell_6t
Xbit_r195_c158 bl[158] br[158] wl[195] vdd gnd cell_6t
Xbit_r196_c158 bl[158] br[158] wl[196] vdd gnd cell_6t
Xbit_r197_c158 bl[158] br[158] wl[197] vdd gnd cell_6t
Xbit_r198_c158 bl[158] br[158] wl[198] vdd gnd cell_6t
Xbit_r199_c158 bl[158] br[158] wl[199] vdd gnd cell_6t
Xbit_r200_c158 bl[158] br[158] wl[200] vdd gnd cell_6t
Xbit_r201_c158 bl[158] br[158] wl[201] vdd gnd cell_6t
Xbit_r202_c158 bl[158] br[158] wl[202] vdd gnd cell_6t
Xbit_r203_c158 bl[158] br[158] wl[203] vdd gnd cell_6t
Xbit_r204_c158 bl[158] br[158] wl[204] vdd gnd cell_6t
Xbit_r205_c158 bl[158] br[158] wl[205] vdd gnd cell_6t
Xbit_r206_c158 bl[158] br[158] wl[206] vdd gnd cell_6t
Xbit_r207_c158 bl[158] br[158] wl[207] vdd gnd cell_6t
Xbit_r208_c158 bl[158] br[158] wl[208] vdd gnd cell_6t
Xbit_r209_c158 bl[158] br[158] wl[209] vdd gnd cell_6t
Xbit_r210_c158 bl[158] br[158] wl[210] vdd gnd cell_6t
Xbit_r211_c158 bl[158] br[158] wl[211] vdd gnd cell_6t
Xbit_r212_c158 bl[158] br[158] wl[212] vdd gnd cell_6t
Xbit_r213_c158 bl[158] br[158] wl[213] vdd gnd cell_6t
Xbit_r214_c158 bl[158] br[158] wl[214] vdd gnd cell_6t
Xbit_r215_c158 bl[158] br[158] wl[215] vdd gnd cell_6t
Xbit_r216_c158 bl[158] br[158] wl[216] vdd gnd cell_6t
Xbit_r217_c158 bl[158] br[158] wl[217] vdd gnd cell_6t
Xbit_r218_c158 bl[158] br[158] wl[218] vdd gnd cell_6t
Xbit_r219_c158 bl[158] br[158] wl[219] vdd gnd cell_6t
Xbit_r220_c158 bl[158] br[158] wl[220] vdd gnd cell_6t
Xbit_r221_c158 bl[158] br[158] wl[221] vdd gnd cell_6t
Xbit_r222_c158 bl[158] br[158] wl[222] vdd gnd cell_6t
Xbit_r223_c158 bl[158] br[158] wl[223] vdd gnd cell_6t
Xbit_r224_c158 bl[158] br[158] wl[224] vdd gnd cell_6t
Xbit_r225_c158 bl[158] br[158] wl[225] vdd gnd cell_6t
Xbit_r226_c158 bl[158] br[158] wl[226] vdd gnd cell_6t
Xbit_r227_c158 bl[158] br[158] wl[227] vdd gnd cell_6t
Xbit_r228_c158 bl[158] br[158] wl[228] vdd gnd cell_6t
Xbit_r229_c158 bl[158] br[158] wl[229] vdd gnd cell_6t
Xbit_r230_c158 bl[158] br[158] wl[230] vdd gnd cell_6t
Xbit_r231_c158 bl[158] br[158] wl[231] vdd gnd cell_6t
Xbit_r232_c158 bl[158] br[158] wl[232] vdd gnd cell_6t
Xbit_r233_c158 bl[158] br[158] wl[233] vdd gnd cell_6t
Xbit_r234_c158 bl[158] br[158] wl[234] vdd gnd cell_6t
Xbit_r235_c158 bl[158] br[158] wl[235] vdd gnd cell_6t
Xbit_r236_c158 bl[158] br[158] wl[236] vdd gnd cell_6t
Xbit_r237_c158 bl[158] br[158] wl[237] vdd gnd cell_6t
Xbit_r238_c158 bl[158] br[158] wl[238] vdd gnd cell_6t
Xbit_r239_c158 bl[158] br[158] wl[239] vdd gnd cell_6t
Xbit_r240_c158 bl[158] br[158] wl[240] vdd gnd cell_6t
Xbit_r241_c158 bl[158] br[158] wl[241] vdd gnd cell_6t
Xbit_r242_c158 bl[158] br[158] wl[242] vdd gnd cell_6t
Xbit_r243_c158 bl[158] br[158] wl[243] vdd gnd cell_6t
Xbit_r244_c158 bl[158] br[158] wl[244] vdd gnd cell_6t
Xbit_r245_c158 bl[158] br[158] wl[245] vdd gnd cell_6t
Xbit_r246_c158 bl[158] br[158] wl[246] vdd gnd cell_6t
Xbit_r247_c158 bl[158] br[158] wl[247] vdd gnd cell_6t
Xbit_r248_c158 bl[158] br[158] wl[248] vdd gnd cell_6t
Xbit_r249_c158 bl[158] br[158] wl[249] vdd gnd cell_6t
Xbit_r250_c158 bl[158] br[158] wl[250] vdd gnd cell_6t
Xbit_r251_c158 bl[158] br[158] wl[251] vdd gnd cell_6t
Xbit_r252_c158 bl[158] br[158] wl[252] vdd gnd cell_6t
Xbit_r253_c158 bl[158] br[158] wl[253] vdd gnd cell_6t
Xbit_r254_c158 bl[158] br[158] wl[254] vdd gnd cell_6t
Xbit_r255_c158 bl[158] br[158] wl[255] vdd gnd cell_6t
Xbit_r0_c159 bl[159] br[159] wl[0] vdd gnd cell_6t
Xbit_r1_c159 bl[159] br[159] wl[1] vdd gnd cell_6t
Xbit_r2_c159 bl[159] br[159] wl[2] vdd gnd cell_6t
Xbit_r3_c159 bl[159] br[159] wl[3] vdd gnd cell_6t
Xbit_r4_c159 bl[159] br[159] wl[4] vdd gnd cell_6t
Xbit_r5_c159 bl[159] br[159] wl[5] vdd gnd cell_6t
Xbit_r6_c159 bl[159] br[159] wl[6] vdd gnd cell_6t
Xbit_r7_c159 bl[159] br[159] wl[7] vdd gnd cell_6t
Xbit_r8_c159 bl[159] br[159] wl[8] vdd gnd cell_6t
Xbit_r9_c159 bl[159] br[159] wl[9] vdd gnd cell_6t
Xbit_r10_c159 bl[159] br[159] wl[10] vdd gnd cell_6t
Xbit_r11_c159 bl[159] br[159] wl[11] vdd gnd cell_6t
Xbit_r12_c159 bl[159] br[159] wl[12] vdd gnd cell_6t
Xbit_r13_c159 bl[159] br[159] wl[13] vdd gnd cell_6t
Xbit_r14_c159 bl[159] br[159] wl[14] vdd gnd cell_6t
Xbit_r15_c159 bl[159] br[159] wl[15] vdd gnd cell_6t
Xbit_r16_c159 bl[159] br[159] wl[16] vdd gnd cell_6t
Xbit_r17_c159 bl[159] br[159] wl[17] vdd gnd cell_6t
Xbit_r18_c159 bl[159] br[159] wl[18] vdd gnd cell_6t
Xbit_r19_c159 bl[159] br[159] wl[19] vdd gnd cell_6t
Xbit_r20_c159 bl[159] br[159] wl[20] vdd gnd cell_6t
Xbit_r21_c159 bl[159] br[159] wl[21] vdd gnd cell_6t
Xbit_r22_c159 bl[159] br[159] wl[22] vdd gnd cell_6t
Xbit_r23_c159 bl[159] br[159] wl[23] vdd gnd cell_6t
Xbit_r24_c159 bl[159] br[159] wl[24] vdd gnd cell_6t
Xbit_r25_c159 bl[159] br[159] wl[25] vdd gnd cell_6t
Xbit_r26_c159 bl[159] br[159] wl[26] vdd gnd cell_6t
Xbit_r27_c159 bl[159] br[159] wl[27] vdd gnd cell_6t
Xbit_r28_c159 bl[159] br[159] wl[28] vdd gnd cell_6t
Xbit_r29_c159 bl[159] br[159] wl[29] vdd gnd cell_6t
Xbit_r30_c159 bl[159] br[159] wl[30] vdd gnd cell_6t
Xbit_r31_c159 bl[159] br[159] wl[31] vdd gnd cell_6t
Xbit_r32_c159 bl[159] br[159] wl[32] vdd gnd cell_6t
Xbit_r33_c159 bl[159] br[159] wl[33] vdd gnd cell_6t
Xbit_r34_c159 bl[159] br[159] wl[34] vdd gnd cell_6t
Xbit_r35_c159 bl[159] br[159] wl[35] vdd gnd cell_6t
Xbit_r36_c159 bl[159] br[159] wl[36] vdd gnd cell_6t
Xbit_r37_c159 bl[159] br[159] wl[37] vdd gnd cell_6t
Xbit_r38_c159 bl[159] br[159] wl[38] vdd gnd cell_6t
Xbit_r39_c159 bl[159] br[159] wl[39] vdd gnd cell_6t
Xbit_r40_c159 bl[159] br[159] wl[40] vdd gnd cell_6t
Xbit_r41_c159 bl[159] br[159] wl[41] vdd gnd cell_6t
Xbit_r42_c159 bl[159] br[159] wl[42] vdd gnd cell_6t
Xbit_r43_c159 bl[159] br[159] wl[43] vdd gnd cell_6t
Xbit_r44_c159 bl[159] br[159] wl[44] vdd gnd cell_6t
Xbit_r45_c159 bl[159] br[159] wl[45] vdd gnd cell_6t
Xbit_r46_c159 bl[159] br[159] wl[46] vdd gnd cell_6t
Xbit_r47_c159 bl[159] br[159] wl[47] vdd gnd cell_6t
Xbit_r48_c159 bl[159] br[159] wl[48] vdd gnd cell_6t
Xbit_r49_c159 bl[159] br[159] wl[49] vdd gnd cell_6t
Xbit_r50_c159 bl[159] br[159] wl[50] vdd gnd cell_6t
Xbit_r51_c159 bl[159] br[159] wl[51] vdd gnd cell_6t
Xbit_r52_c159 bl[159] br[159] wl[52] vdd gnd cell_6t
Xbit_r53_c159 bl[159] br[159] wl[53] vdd gnd cell_6t
Xbit_r54_c159 bl[159] br[159] wl[54] vdd gnd cell_6t
Xbit_r55_c159 bl[159] br[159] wl[55] vdd gnd cell_6t
Xbit_r56_c159 bl[159] br[159] wl[56] vdd gnd cell_6t
Xbit_r57_c159 bl[159] br[159] wl[57] vdd gnd cell_6t
Xbit_r58_c159 bl[159] br[159] wl[58] vdd gnd cell_6t
Xbit_r59_c159 bl[159] br[159] wl[59] vdd gnd cell_6t
Xbit_r60_c159 bl[159] br[159] wl[60] vdd gnd cell_6t
Xbit_r61_c159 bl[159] br[159] wl[61] vdd gnd cell_6t
Xbit_r62_c159 bl[159] br[159] wl[62] vdd gnd cell_6t
Xbit_r63_c159 bl[159] br[159] wl[63] vdd gnd cell_6t
Xbit_r64_c159 bl[159] br[159] wl[64] vdd gnd cell_6t
Xbit_r65_c159 bl[159] br[159] wl[65] vdd gnd cell_6t
Xbit_r66_c159 bl[159] br[159] wl[66] vdd gnd cell_6t
Xbit_r67_c159 bl[159] br[159] wl[67] vdd gnd cell_6t
Xbit_r68_c159 bl[159] br[159] wl[68] vdd gnd cell_6t
Xbit_r69_c159 bl[159] br[159] wl[69] vdd gnd cell_6t
Xbit_r70_c159 bl[159] br[159] wl[70] vdd gnd cell_6t
Xbit_r71_c159 bl[159] br[159] wl[71] vdd gnd cell_6t
Xbit_r72_c159 bl[159] br[159] wl[72] vdd gnd cell_6t
Xbit_r73_c159 bl[159] br[159] wl[73] vdd gnd cell_6t
Xbit_r74_c159 bl[159] br[159] wl[74] vdd gnd cell_6t
Xbit_r75_c159 bl[159] br[159] wl[75] vdd gnd cell_6t
Xbit_r76_c159 bl[159] br[159] wl[76] vdd gnd cell_6t
Xbit_r77_c159 bl[159] br[159] wl[77] vdd gnd cell_6t
Xbit_r78_c159 bl[159] br[159] wl[78] vdd gnd cell_6t
Xbit_r79_c159 bl[159] br[159] wl[79] vdd gnd cell_6t
Xbit_r80_c159 bl[159] br[159] wl[80] vdd gnd cell_6t
Xbit_r81_c159 bl[159] br[159] wl[81] vdd gnd cell_6t
Xbit_r82_c159 bl[159] br[159] wl[82] vdd gnd cell_6t
Xbit_r83_c159 bl[159] br[159] wl[83] vdd gnd cell_6t
Xbit_r84_c159 bl[159] br[159] wl[84] vdd gnd cell_6t
Xbit_r85_c159 bl[159] br[159] wl[85] vdd gnd cell_6t
Xbit_r86_c159 bl[159] br[159] wl[86] vdd gnd cell_6t
Xbit_r87_c159 bl[159] br[159] wl[87] vdd gnd cell_6t
Xbit_r88_c159 bl[159] br[159] wl[88] vdd gnd cell_6t
Xbit_r89_c159 bl[159] br[159] wl[89] vdd gnd cell_6t
Xbit_r90_c159 bl[159] br[159] wl[90] vdd gnd cell_6t
Xbit_r91_c159 bl[159] br[159] wl[91] vdd gnd cell_6t
Xbit_r92_c159 bl[159] br[159] wl[92] vdd gnd cell_6t
Xbit_r93_c159 bl[159] br[159] wl[93] vdd gnd cell_6t
Xbit_r94_c159 bl[159] br[159] wl[94] vdd gnd cell_6t
Xbit_r95_c159 bl[159] br[159] wl[95] vdd gnd cell_6t
Xbit_r96_c159 bl[159] br[159] wl[96] vdd gnd cell_6t
Xbit_r97_c159 bl[159] br[159] wl[97] vdd gnd cell_6t
Xbit_r98_c159 bl[159] br[159] wl[98] vdd gnd cell_6t
Xbit_r99_c159 bl[159] br[159] wl[99] vdd gnd cell_6t
Xbit_r100_c159 bl[159] br[159] wl[100] vdd gnd cell_6t
Xbit_r101_c159 bl[159] br[159] wl[101] vdd gnd cell_6t
Xbit_r102_c159 bl[159] br[159] wl[102] vdd gnd cell_6t
Xbit_r103_c159 bl[159] br[159] wl[103] vdd gnd cell_6t
Xbit_r104_c159 bl[159] br[159] wl[104] vdd gnd cell_6t
Xbit_r105_c159 bl[159] br[159] wl[105] vdd gnd cell_6t
Xbit_r106_c159 bl[159] br[159] wl[106] vdd gnd cell_6t
Xbit_r107_c159 bl[159] br[159] wl[107] vdd gnd cell_6t
Xbit_r108_c159 bl[159] br[159] wl[108] vdd gnd cell_6t
Xbit_r109_c159 bl[159] br[159] wl[109] vdd gnd cell_6t
Xbit_r110_c159 bl[159] br[159] wl[110] vdd gnd cell_6t
Xbit_r111_c159 bl[159] br[159] wl[111] vdd gnd cell_6t
Xbit_r112_c159 bl[159] br[159] wl[112] vdd gnd cell_6t
Xbit_r113_c159 bl[159] br[159] wl[113] vdd gnd cell_6t
Xbit_r114_c159 bl[159] br[159] wl[114] vdd gnd cell_6t
Xbit_r115_c159 bl[159] br[159] wl[115] vdd gnd cell_6t
Xbit_r116_c159 bl[159] br[159] wl[116] vdd gnd cell_6t
Xbit_r117_c159 bl[159] br[159] wl[117] vdd gnd cell_6t
Xbit_r118_c159 bl[159] br[159] wl[118] vdd gnd cell_6t
Xbit_r119_c159 bl[159] br[159] wl[119] vdd gnd cell_6t
Xbit_r120_c159 bl[159] br[159] wl[120] vdd gnd cell_6t
Xbit_r121_c159 bl[159] br[159] wl[121] vdd gnd cell_6t
Xbit_r122_c159 bl[159] br[159] wl[122] vdd gnd cell_6t
Xbit_r123_c159 bl[159] br[159] wl[123] vdd gnd cell_6t
Xbit_r124_c159 bl[159] br[159] wl[124] vdd gnd cell_6t
Xbit_r125_c159 bl[159] br[159] wl[125] vdd gnd cell_6t
Xbit_r126_c159 bl[159] br[159] wl[126] vdd gnd cell_6t
Xbit_r127_c159 bl[159] br[159] wl[127] vdd gnd cell_6t
Xbit_r128_c159 bl[159] br[159] wl[128] vdd gnd cell_6t
Xbit_r129_c159 bl[159] br[159] wl[129] vdd gnd cell_6t
Xbit_r130_c159 bl[159] br[159] wl[130] vdd gnd cell_6t
Xbit_r131_c159 bl[159] br[159] wl[131] vdd gnd cell_6t
Xbit_r132_c159 bl[159] br[159] wl[132] vdd gnd cell_6t
Xbit_r133_c159 bl[159] br[159] wl[133] vdd gnd cell_6t
Xbit_r134_c159 bl[159] br[159] wl[134] vdd gnd cell_6t
Xbit_r135_c159 bl[159] br[159] wl[135] vdd gnd cell_6t
Xbit_r136_c159 bl[159] br[159] wl[136] vdd gnd cell_6t
Xbit_r137_c159 bl[159] br[159] wl[137] vdd gnd cell_6t
Xbit_r138_c159 bl[159] br[159] wl[138] vdd gnd cell_6t
Xbit_r139_c159 bl[159] br[159] wl[139] vdd gnd cell_6t
Xbit_r140_c159 bl[159] br[159] wl[140] vdd gnd cell_6t
Xbit_r141_c159 bl[159] br[159] wl[141] vdd gnd cell_6t
Xbit_r142_c159 bl[159] br[159] wl[142] vdd gnd cell_6t
Xbit_r143_c159 bl[159] br[159] wl[143] vdd gnd cell_6t
Xbit_r144_c159 bl[159] br[159] wl[144] vdd gnd cell_6t
Xbit_r145_c159 bl[159] br[159] wl[145] vdd gnd cell_6t
Xbit_r146_c159 bl[159] br[159] wl[146] vdd gnd cell_6t
Xbit_r147_c159 bl[159] br[159] wl[147] vdd gnd cell_6t
Xbit_r148_c159 bl[159] br[159] wl[148] vdd gnd cell_6t
Xbit_r149_c159 bl[159] br[159] wl[149] vdd gnd cell_6t
Xbit_r150_c159 bl[159] br[159] wl[150] vdd gnd cell_6t
Xbit_r151_c159 bl[159] br[159] wl[151] vdd gnd cell_6t
Xbit_r152_c159 bl[159] br[159] wl[152] vdd gnd cell_6t
Xbit_r153_c159 bl[159] br[159] wl[153] vdd gnd cell_6t
Xbit_r154_c159 bl[159] br[159] wl[154] vdd gnd cell_6t
Xbit_r155_c159 bl[159] br[159] wl[155] vdd gnd cell_6t
Xbit_r156_c159 bl[159] br[159] wl[156] vdd gnd cell_6t
Xbit_r157_c159 bl[159] br[159] wl[157] vdd gnd cell_6t
Xbit_r158_c159 bl[159] br[159] wl[158] vdd gnd cell_6t
Xbit_r159_c159 bl[159] br[159] wl[159] vdd gnd cell_6t
Xbit_r160_c159 bl[159] br[159] wl[160] vdd gnd cell_6t
Xbit_r161_c159 bl[159] br[159] wl[161] vdd gnd cell_6t
Xbit_r162_c159 bl[159] br[159] wl[162] vdd gnd cell_6t
Xbit_r163_c159 bl[159] br[159] wl[163] vdd gnd cell_6t
Xbit_r164_c159 bl[159] br[159] wl[164] vdd gnd cell_6t
Xbit_r165_c159 bl[159] br[159] wl[165] vdd gnd cell_6t
Xbit_r166_c159 bl[159] br[159] wl[166] vdd gnd cell_6t
Xbit_r167_c159 bl[159] br[159] wl[167] vdd gnd cell_6t
Xbit_r168_c159 bl[159] br[159] wl[168] vdd gnd cell_6t
Xbit_r169_c159 bl[159] br[159] wl[169] vdd gnd cell_6t
Xbit_r170_c159 bl[159] br[159] wl[170] vdd gnd cell_6t
Xbit_r171_c159 bl[159] br[159] wl[171] vdd gnd cell_6t
Xbit_r172_c159 bl[159] br[159] wl[172] vdd gnd cell_6t
Xbit_r173_c159 bl[159] br[159] wl[173] vdd gnd cell_6t
Xbit_r174_c159 bl[159] br[159] wl[174] vdd gnd cell_6t
Xbit_r175_c159 bl[159] br[159] wl[175] vdd gnd cell_6t
Xbit_r176_c159 bl[159] br[159] wl[176] vdd gnd cell_6t
Xbit_r177_c159 bl[159] br[159] wl[177] vdd gnd cell_6t
Xbit_r178_c159 bl[159] br[159] wl[178] vdd gnd cell_6t
Xbit_r179_c159 bl[159] br[159] wl[179] vdd gnd cell_6t
Xbit_r180_c159 bl[159] br[159] wl[180] vdd gnd cell_6t
Xbit_r181_c159 bl[159] br[159] wl[181] vdd gnd cell_6t
Xbit_r182_c159 bl[159] br[159] wl[182] vdd gnd cell_6t
Xbit_r183_c159 bl[159] br[159] wl[183] vdd gnd cell_6t
Xbit_r184_c159 bl[159] br[159] wl[184] vdd gnd cell_6t
Xbit_r185_c159 bl[159] br[159] wl[185] vdd gnd cell_6t
Xbit_r186_c159 bl[159] br[159] wl[186] vdd gnd cell_6t
Xbit_r187_c159 bl[159] br[159] wl[187] vdd gnd cell_6t
Xbit_r188_c159 bl[159] br[159] wl[188] vdd gnd cell_6t
Xbit_r189_c159 bl[159] br[159] wl[189] vdd gnd cell_6t
Xbit_r190_c159 bl[159] br[159] wl[190] vdd gnd cell_6t
Xbit_r191_c159 bl[159] br[159] wl[191] vdd gnd cell_6t
Xbit_r192_c159 bl[159] br[159] wl[192] vdd gnd cell_6t
Xbit_r193_c159 bl[159] br[159] wl[193] vdd gnd cell_6t
Xbit_r194_c159 bl[159] br[159] wl[194] vdd gnd cell_6t
Xbit_r195_c159 bl[159] br[159] wl[195] vdd gnd cell_6t
Xbit_r196_c159 bl[159] br[159] wl[196] vdd gnd cell_6t
Xbit_r197_c159 bl[159] br[159] wl[197] vdd gnd cell_6t
Xbit_r198_c159 bl[159] br[159] wl[198] vdd gnd cell_6t
Xbit_r199_c159 bl[159] br[159] wl[199] vdd gnd cell_6t
Xbit_r200_c159 bl[159] br[159] wl[200] vdd gnd cell_6t
Xbit_r201_c159 bl[159] br[159] wl[201] vdd gnd cell_6t
Xbit_r202_c159 bl[159] br[159] wl[202] vdd gnd cell_6t
Xbit_r203_c159 bl[159] br[159] wl[203] vdd gnd cell_6t
Xbit_r204_c159 bl[159] br[159] wl[204] vdd gnd cell_6t
Xbit_r205_c159 bl[159] br[159] wl[205] vdd gnd cell_6t
Xbit_r206_c159 bl[159] br[159] wl[206] vdd gnd cell_6t
Xbit_r207_c159 bl[159] br[159] wl[207] vdd gnd cell_6t
Xbit_r208_c159 bl[159] br[159] wl[208] vdd gnd cell_6t
Xbit_r209_c159 bl[159] br[159] wl[209] vdd gnd cell_6t
Xbit_r210_c159 bl[159] br[159] wl[210] vdd gnd cell_6t
Xbit_r211_c159 bl[159] br[159] wl[211] vdd gnd cell_6t
Xbit_r212_c159 bl[159] br[159] wl[212] vdd gnd cell_6t
Xbit_r213_c159 bl[159] br[159] wl[213] vdd gnd cell_6t
Xbit_r214_c159 bl[159] br[159] wl[214] vdd gnd cell_6t
Xbit_r215_c159 bl[159] br[159] wl[215] vdd gnd cell_6t
Xbit_r216_c159 bl[159] br[159] wl[216] vdd gnd cell_6t
Xbit_r217_c159 bl[159] br[159] wl[217] vdd gnd cell_6t
Xbit_r218_c159 bl[159] br[159] wl[218] vdd gnd cell_6t
Xbit_r219_c159 bl[159] br[159] wl[219] vdd gnd cell_6t
Xbit_r220_c159 bl[159] br[159] wl[220] vdd gnd cell_6t
Xbit_r221_c159 bl[159] br[159] wl[221] vdd gnd cell_6t
Xbit_r222_c159 bl[159] br[159] wl[222] vdd gnd cell_6t
Xbit_r223_c159 bl[159] br[159] wl[223] vdd gnd cell_6t
Xbit_r224_c159 bl[159] br[159] wl[224] vdd gnd cell_6t
Xbit_r225_c159 bl[159] br[159] wl[225] vdd gnd cell_6t
Xbit_r226_c159 bl[159] br[159] wl[226] vdd gnd cell_6t
Xbit_r227_c159 bl[159] br[159] wl[227] vdd gnd cell_6t
Xbit_r228_c159 bl[159] br[159] wl[228] vdd gnd cell_6t
Xbit_r229_c159 bl[159] br[159] wl[229] vdd gnd cell_6t
Xbit_r230_c159 bl[159] br[159] wl[230] vdd gnd cell_6t
Xbit_r231_c159 bl[159] br[159] wl[231] vdd gnd cell_6t
Xbit_r232_c159 bl[159] br[159] wl[232] vdd gnd cell_6t
Xbit_r233_c159 bl[159] br[159] wl[233] vdd gnd cell_6t
Xbit_r234_c159 bl[159] br[159] wl[234] vdd gnd cell_6t
Xbit_r235_c159 bl[159] br[159] wl[235] vdd gnd cell_6t
Xbit_r236_c159 bl[159] br[159] wl[236] vdd gnd cell_6t
Xbit_r237_c159 bl[159] br[159] wl[237] vdd gnd cell_6t
Xbit_r238_c159 bl[159] br[159] wl[238] vdd gnd cell_6t
Xbit_r239_c159 bl[159] br[159] wl[239] vdd gnd cell_6t
Xbit_r240_c159 bl[159] br[159] wl[240] vdd gnd cell_6t
Xbit_r241_c159 bl[159] br[159] wl[241] vdd gnd cell_6t
Xbit_r242_c159 bl[159] br[159] wl[242] vdd gnd cell_6t
Xbit_r243_c159 bl[159] br[159] wl[243] vdd gnd cell_6t
Xbit_r244_c159 bl[159] br[159] wl[244] vdd gnd cell_6t
Xbit_r245_c159 bl[159] br[159] wl[245] vdd gnd cell_6t
Xbit_r246_c159 bl[159] br[159] wl[246] vdd gnd cell_6t
Xbit_r247_c159 bl[159] br[159] wl[247] vdd gnd cell_6t
Xbit_r248_c159 bl[159] br[159] wl[248] vdd gnd cell_6t
Xbit_r249_c159 bl[159] br[159] wl[249] vdd gnd cell_6t
Xbit_r250_c159 bl[159] br[159] wl[250] vdd gnd cell_6t
Xbit_r251_c159 bl[159] br[159] wl[251] vdd gnd cell_6t
Xbit_r252_c159 bl[159] br[159] wl[252] vdd gnd cell_6t
Xbit_r253_c159 bl[159] br[159] wl[253] vdd gnd cell_6t
Xbit_r254_c159 bl[159] br[159] wl[254] vdd gnd cell_6t
Xbit_r255_c159 bl[159] br[159] wl[255] vdd gnd cell_6t
Xbit_r0_c160 bl[160] br[160] wl[0] vdd gnd cell_6t
Xbit_r1_c160 bl[160] br[160] wl[1] vdd gnd cell_6t
Xbit_r2_c160 bl[160] br[160] wl[2] vdd gnd cell_6t
Xbit_r3_c160 bl[160] br[160] wl[3] vdd gnd cell_6t
Xbit_r4_c160 bl[160] br[160] wl[4] vdd gnd cell_6t
Xbit_r5_c160 bl[160] br[160] wl[5] vdd gnd cell_6t
Xbit_r6_c160 bl[160] br[160] wl[6] vdd gnd cell_6t
Xbit_r7_c160 bl[160] br[160] wl[7] vdd gnd cell_6t
Xbit_r8_c160 bl[160] br[160] wl[8] vdd gnd cell_6t
Xbit_r9_c160 bl[160] br[160] wl[9] vdd gnd cell_6t
Xbit_r10_c160 bl[160] br[160] wl[10] vdd gnd cell_6t
Xbit_r11_c160 bl[160] br[160] wl[11] vdd gnd cell_6t
Xbit_r12_c160 bl[160] br[160] wl[12] vdd gnd cell_6t
Xbit_r13_c160 bl[160] br[160] wl[13] vdd gnd cell_6t
Xbit_r14_c160 bl[160] br[160] wl[14] vdd gnd cell_6t
Xbit_r15_c160 bl[160] br[160] wl[15] vdd gnd cell_6t
Xbit_r16_c160 bl[160] br[160] wl[16] vdd gnd cell_6t
Xbit_r17_c160 bl[160] br[160] wl[17] vdd gnd cell_6t
Xbit_r18_c160 bl[160] br[160] wl[18] vdd gnd cell_6t
Xbit_r19_c160 bl[160] br[160] wl[19] vdd gnd cell_6t
Xbit_r20_c160 bl[160] br[160] wl[20] vdd gnd cell_6t
Xbit_r21_c160 bl[160] br[160] wl[21] vdd gnd cell_6t
Xbit_r22_c160 bl[160] br[160] wl[22] vdd gnd cell_6t
Xbit_r23_c160 bl[160] br[160] wl[23] vdd gnd cell_6t
Xbit_r24_c160 bl[160] br[160] wl[24] vdd gnd cell_6t
Xbit_r25_c160 bl[160] br[160] wl[25] vdd gnd cell_6t
Xbit_r26_c160 bl[160] br[160] wl[26] vdd gnd cell_6t
Xbit_r27_c160 bl[160] br[160] wl[27] vdd gnd cell_6t
Xbit_r28_c160 bl[160] br[160] wl[28] vdd gnd cell_6t
Xbit_r29_c160 bl[160] br[160] wl[29] vdd gnd cell_6t
Xbit_r30_c160 bl[160] br[160] wl[30] vdd gnd cell_6t
Xbit_r31_c160 bl[160] br[160] wl[31] vdd gnd cell_6t
Xbit_r32_c160 bl[160] br[160] wl[32] vdd gnd cell_6t
Xbit_r33_c160 bl[160] br[160] wl[33] vdd gnd cell_6t
Xbit_r34_c160 bl[160] br[160] wl[34] vdd gnd cell_6t
Xbit_r35_c160 bl[160] br[160] wl[35] vdd gnd cell_6t
Xbit_r36_c160 bl[160] br[160] wl[36] vdd gnd cell_6t
Xbit_r37_c160 bl[160] br[160] wl[37] vdd gnd cell_6t
Xbit_r38_c160 bl[160] br[160] wl[38] vdd gnd cell_6t
Xbit_r39_c160 bl[160] br[160] wl[39] vdd gnd cell_6t
Xbit_r40_c160 bl[160] br[160] wl[40] vdd gnd cell_6t
Xbit_r41_c160 bl[160] br[160] wl[41] vdd gnd cell_6t
Xbit_r42_c160 bl[160] br[160] wl[42] vdd gnd cell_6t
Xbit_r43_c160 bl[160] br[160] wl[43] vdd gnd cell_6t
Xbit_r44_c160 bl[160] br[160] wl[44] vdd gnd cell_6t
Xbit_r45_c160 bl[160] br[160] wl[45] vdd gnd cell_6t
Xbit_r46_c160 bl[160] br[160] wl[46] vdd gnd cell_6t
Xbit_r47_c160 bl[160] br[160] wl[47] vdd gnd cell_6t
Xbit_r48_c160 bl[160] br[160] wl[48] vdd gnd cell_6t
Xbit_r49_c160 bl[160] br[160] wl[49] vdd gnd cell_6t
Xbit_r50_c160 bl[160] br[160] wl[50] vdd gnd cell_6t
Xbit_r51_c160 bl[160] br[160] wl[51] vdd gnd cell_6t
Xbit_r52_c160 bl[160] br[160] wl[52] vdd gnd cell_6t
Xbit_r53_c160 bl[160] br[160] wl[53] vdd gnd cell_6t
Xbit_r54_c160 bl[160] br[160] wl[54] vdd gnd cell_6t
Xbit_r55_c160 bl[160] br[160] wl[55] vdd gnd cell_6t
Xbit_r56_c160 bl[160] br[160] wl[56] vdd gnd cell_6t
Xbit_r57_c160 bl[160] br[160] wl[57] vdd gnd cell_6t
Xbit_r58_c160 bl[160] br[160] wl[58] vdd gnd cell_6t
Xbit_r59_c160 bl[160] br[160] wl[59] vdd gnd cell_6t
Xbit_r60_c160 bl[160] br[160] wl[60] vdd gnd cell_6t
Xbit_r61_c160 bl[160] br[160] wl[61] vdd gnd cell_6t
Xbit_r62_c160 bl[160] br[160] wl[62] vdd gnd cell_6t
Xbit_r63_c160 bl[160] br[160] wl[63] vdd gnd cell_6t
Xbit_r64_c160 bl[160] br[160] wl[64] vdd gnd cell_6t
Xbit_r65_c160 bl[160] br[160] wl[65] vdd gnd cell_6t
Xbit_r66_c160 bl[160] br[160] wl[66] vdd gnd cell_6t
Xbit_r67_c160 bl[160] br[160] wl[67] vdd gnd cell_6t
Xbit_r68_c160 bl[160] br[160] wl[68] vdd gnd cell_6t
Xbit_r69_c160 bl[160] br[160] wl[69] vdd gnd cell_6t
Xbit_r70_c160 bl[160] br[160] wl[70] vdd gnd cell_6t
Xbit_r71_c160 bl[160] br[160] wl[71] vdd gnd cell_6t
Xbit_r72_c160 bl[160] br[160] wl[72] vdd gnd cell_6t
Xbit_r73_c160 bl[160] br[160] wl[73] vdd gnd cell_6t
Xbit_r74_c160 bl[160] br[160] wl[74] vdd gnd cell_6t
Xbit_r75_c160 bl[160] br[160] wl[75] vdd gnd cell_6t
Xbit_r76_c160 bl[160] br[160] wl[76] vdd gnd cell_6t
Xbit_r77_c160 bl[160] br[160] wl[77] vdd gnd cell_6t
Xbit_r78_c160 bl[160] br[160] wl[78] vdd gnd cell_6t
Xbit_r79_c160 bl[160] br[160] wl[79] vdd gnd cell_6t
Xbit_r80_c160 bl[160] br[160] wl[80] vdd gnd cell_6t
Xbit_r81_c160 bl[160] br[160] wl[81] vdd gnd cell_6t
Xbit_r82_c160 bl[160] br[160] wl[82] vdd gnd cell_6t
Xbit_r83_c160 bl[160] br[160] wl[83] vdd gnd cell_6t
Xbit_r84_c160 bl[160] br[160] wl[84] vdd gnd cell_6t
Xbit_r85_c160 bl[160] br[160] wl[85] vdd gnd cell_6t
Xbit_r86_c160 bl[160] br[160] wl[86] vdd gnd cell_6t
Xbit_r87_c160 bl[160] br[160] wl[87] vdd gnd cell_6t
Xbit_r88_c160 bl[160] br[160] wl[88] vdd gnd cell_6t
Xbit_r89_c160 bl[160] br[160] wl[89] vdd gnd cell_6t
Xbit_r90_c160 bl[160] br[160] wl[90] vdd gnd cell_6t
Xbit_r91_c160 bl[160] br[160] wl[91] vdd gnd cell_6t
Xbit_r92_c160 bl[160] br[160] wl[92] vdd gnd cell_6t
Xbit_r93_c160 bl[160] br[160] wl[93] vdd gnd cell_6t
Xbit_r94_c160 bl[160] br[160] wl[94] vdd gnd cell_6t
Xbit_r95_c160 bl[160] br[160] wl[95] vdd gnd cell_6t
Xbit_r96_c160 bl[160] br[160] wl[96] vdd gnd cell_6t
Xbit_r97_c160 bl[160] br[160] wl[97] vdd gnd cell_6t
Xbit_r98_c160 bl[160] br[160] wl[98] vdd gnd cell_6t
Xbit_r99_c160 bl[160] br[160] wl[99] vdd gnd cell_6t
Xbit_r100_c160 bl[160] br[160] wl[100] vdd gnd cell_6t
Xbit_r101_c160 bl[160] br[160] wl[101] vdd gnd cell_6t
Xbit_r102_c160 bl[160] br[160] wl[102] vdd gnd cell_6t
Xbit_r103_c160 bl[160] br[160] wl[103] vdd gnd cell_6t
Xbit_r104_c160 bl[160] br[160] wl[104] vdd gnd cell_6t
Xbit_r105_c160 bl[160] br[160] wl[105] vdd gnd cell_6t
Xbit_r106_c160 bl[160] br[160] wl[106] vdd gnd cell_6t
Xbit_r107_c160 bl[160] br[160] wl[107] vdd gnd cell_6t
Xbit_r108_c160 bl[160] br[160] wl[108] vdd gnd cell_6t
Xbit_r109_c160 bl[160] br[160] wl[109] vdd gnd cell_6t
Xbit_r110_c160 bl[160] br[160] wl[110] vdd gnd cell_6t
Xbit_r111_c160 bl[160] br[160] wl[111] vdd gnd cell_6t
Xbit_r112_c160 bl[160] br[160] wl[112] vdd gnd cell_6t
Xbit_r113_c160 bl[160] br[160] wl[113] vdd gnd cell_6t
Xbit_r114_c160 bl[160] br[160] wl[114] vdd gnd cell_6t
Xbit_r115_c160 bl[160] br[160] wl[115] vdd gnd cell_6t
Xbit_r116_c160 bl[160] br[160] wl[116] vdd gnd cell_6t
Xbit_r117_c160 bl[160] br[160] wl[117] vdd gnd cell_6t
Xbit_r118_c160 bl[160] br[160] wl[118] vdd gnd cell_6t
Xbit_r119_c160 bl[160] br[160] wl[119] vdd gnd cell_6t
Xbit_r120_c160 bl[160] br[160] wl[120] vdd gnd cell_6t
Xbit_r121_c160 bl[160] br[160] wl[121] vdd gnd cell_6t
Xbit_r122_c160 bl[160] br[160] wl[122] vdd gnd cell_6t
Xbit_r123_c160 bl[160] br[160] wl[123] vdd gnd cell_6t
Xbit_r124_c160 bl[160] br[160] wl[124] vdd gnd cell_6t
Xbit_r125_c160 bl[160] br[160] wl[125] vdd gnd cell_6t
Xbit_r126_c160 bl[160] br[160] wl[126] vdd gnd cell_6t
Xbit_r127_c160 bl[160] br[160] wl[127] vdd gnd cell_6t
Xbit_r128_c160 bl[160] br[160] wl[128] vdd gnd cell_6t
Xbit_r129_c160 bl[160] br[160] wl[129] vdd gnd cell_6t
Xbit_r130_c160 bl[160] br[160] wl[130] vdd gnd cell_6t
Xbit_r131_c160 bl[160] br[160] wl[131] vdd gnd cell_6t
Xbit_r132_c160 bl[160] br[160] wl[132] vdd gnd cell_6t
Xbit_r133_c160 bl[160] br[160] wl[133] vdd gnd cell_6t
Xbit_r134_c160 bl[160] br[160] wl[134] vdd gnd cell_6t
Xbit_r135_c160 bl[160] br[160] wl[135] vdd gnd cell_6t
Xbit_r136_c160 bl[160] br[160] wl[136] vdd gnd cell_6t
Xbit_r137_c160 bl[160] br[160] wl[137] vdd gnd cell_6t
Xbit_r138_c160 bl[160] br[160] wl[138] vdd gnd cell_6t
Xbit_r139_c160 bl[160] br[160] wl[139] vdd gnd cell_6t
Xbit_r140_c160 bl[160] br[160] wl[140] vdd gnd cell_6t
Xbit_r141_c160 bl[160] br[160] wl[141] vdd gnd cell_6t
Xbit_r142_c160 bl[160] br[160] wl[142] vdd gnd cell_6t
Xbit_r143_c160 bl[160] br[160] wl[143] vdd gnd cell_6t
Xbit_r144_c160 bl[160] br[160] wl[144] vdd gnd cell_6t
Xbit_r145_c160 bl[160] br[160] wl[145] vdd gnd cell_6t
Xbit_r146_c160 bl[160] br[160] wl[146] vdd gnd cell_6t
Xbit_r147_c160 bl[160] br[160] wl[147] vdd gnd cell_6t
Xbit_r148_c160 bl[160] br[160] wl[148] vdd gnd cell_6t
Xbit_r149_c160 bl[160] br[160] wl[149] vdd gnd cell_6t
Xbit_r150_c160 bl[160] br[160] wl[150] vdd gnd cell_6t
Xbit_r151_c160 bl[160] br[160] wl[151] vdd gnd cell_6t
Xbit_r152_c160 bl[160] br[160] wl[152] vdd gnd cell_6t
Xbit_r153_c160 bl[160] br[160] wl[153] vdd gnd cell_6t
Xbit_r154_c160 bl[160] br[160] wl[154] vdd gnd cell_6t
Xbit_r155_c160 bl[160] br[160] wl[155] vdd gnd cell_6t
Xbit_r156_c160 bl[160] br[160] wl[156] vdd gnd cell_6t
Xbit_r157_c160 bl[160] br[160] wl[157] vdd gnd cell_6t
Xbit_r158_c160 bl[160] br[160] wl[158] vdd gnd cell_6t
Xbit_r159_c160 bl[160] br[160] wl[159] vdd gnd cell_6t
Xbit_r160_c160 bl[160] br[160] wl[160] vdd gnd cell_6t
Xbit_r161_c160 bl[160] br[160] wl[161] vdd gnd cell_6t
Xbit_r162_c160 bl[160] br[160] wl[162] vdd gnd cell_6t
Xbit_r163_c160 bl[160] br[160] wl[163] vdd gnd cell_6t
Xbit_r164_c160 bl[160] br[160] wl[164] vdd gnd cell_6t
Xbit_r165_c160 bl[160] br[160] wl[165] vdd gnd cell_6t
Xbit_r166_c160 bl[160] br[160] wl[166] vdd gnd cell_6t
Xbit_r167_c160 bl[160] br[160] wl[167] vdd gnd cell_6t
Xbit_r168_c160 bl[160] br[160] wl[168] vdd gnd cell_6t
Xbit_r169_c160 bl[160] br[160] wl[169] vdd gnd cell_6t
Xbit_r170_c160 bl[160] br[160] wl[170] vdd gnd cell_6t
Xbit_r171_c160 bl[160] br[160] wl[171] vdd gnd cell_6t
Xbit_r172_c160 bl[160] br[160] wl[172] vdd gnd cell_6t
Xbit_r173_c160 bl[160] br[160] wl[173] vdd gnd cell_6t
Xbit_r174_c160 bl[160] br[160] wl[174] vdd gnd cell_6t
Xbit_r175_c160 bl[160] br[160] wl[175] vdd gnd cell_6t
Xbit_r176_c160 bl[160] br[160] wl[176] vdd gnd cell_6t
Xbit_r177_c160 bl[160] br[160] wl[177] vdd gnd cell_6t
Xbit_r178_c160 bl[160] br[160] wl[178] vdd gnd cell_6t
Xbit_r179_c160 bl[160] br[160] wl[179] vdd gnd cell_6t
Xbit_r180_c160 bl[160] br[160] wl[180] vdd gnd cell_6t
Xbit_r181_c160 bl[160] br[160] wl[181] vdd gnd cell_6t
Xbit_r182_c160 bl[160] br[160] wl[182] vdd gnd cell_6t
Xbit_r183_c160 bl[160] br[160] wl[183] vdd gnd cell_6t
Xbit_r184_c160 bl[160] br[160] wl[184] vdd gnd cell_6t
Xbit_r185_c160 bl[160] br[160] wl[185] vdd gnd cell_6t
Xbit_r186_c160 bl[160] br[160] wl[186] vdd gnd cell_6t
Xbit_r187_c160 bl[160] br[160] wl[187] vdd gnd cell_6t
Xbit_r188_c160 bl[160] br[160] wl[188] vdd gnd cell_6t
Xbit_r189_c160 bl[160] br[160] wl[189] vdd gnd cell_6t
Xbit_r190_c160 bl[160] br[160] wl[190] vdd gnd cell_6t
Xbit_r191_c160 bl[160] br[160] wl[191] vdd gnd cell_6t
Xbit_r192_c160 bl[160] br[160] wl[192] vdd gnd cell_6t
Xbit_r193_c160 bl[160] br[160] wl[193] vdd gnd cell_6t
Xbit_r194_c160 bl[160] br[160] wl[194] vdd gnd cell_6t
Xbit_r195_c160 bl[160] br[160] wl[195] vdd gnd cell_6t
Xbit_r196_c160 bl[160] br[160] wl[196] vdd gnd cell_6t
Xbit_r197_c160 bl[160] br[160] wl[197] vdd gnd cell_6t
Xbit_r198_c160 bl[160] br[160] wl[198] vdd gnd cell_6t
Xbit_r199_c160 bl[160] br[160] wl[199] vdd gnd cell_6t
Xbit_r200_c160 bl[160] br[160] wl[200] vdd gnd cell_6t
Xbit_r201_c160 bl[160] br[160] wl[201] vdd gnd cell_6t
Xbit_r202_c160 bl[160] br[160] wl[202] vdd gnd cell_6t
Xbit_r203_c160 bl[160] br[160] wl[203] vdd gnd cell_6t
Xbit_r204_c160 bl[160] br[160] wl[204] vdd gnd cell_6t
Xbit_r205_c160 bl[160] br[160] wl[205] vdd gnd cell_6t
Xbit_r206_c160 bl[160] br[160] wl[206] vdd gnd cell_6t
Xbit_r207_c160 bl[160] br[160] wl[207] vdd gnd cell_6t
Xbit_r208_c160 bl[160] br[160] wl[208] vdd gnd cell_6t
Xbit_r209_c160 bl[160] br[160] wl[209] vdd gnd cell_6t
Xbit_r210_c160 bl[160] br[160] wl[210] vdd gnd cell_6t
Xbit_r211_c160 bl[160] br[160] wl[211] vdd gnd cell_6t
Xbit_r212_c160 bl[160] br[160] wl[212] vdd gnd cell_6t
Xbit_r213_c160 bl[160] br[160] wl[213] vdd gnd cell_6t
Xbit_r214_c160 bl[160] br[160] wl[214] vdd gnd cell_6t
Xbit_r215_c160 bl[160] br[160] wl[215] vdd gnd cell_6t
Xbit_r216_c160 bl[160] br[160] wl[216] vdd gnd cell_6t
Xbit_r217_c160 bl[160] br[160] wl[217] vdd gnd cell_6t
Xbit_r218_c160 bl[160] br[160] wl[218] vdd gnd cell_6t
Xbit_r219_c160 bl[160] br[160] wl[219] vdd gnd cell_6t
Xbit_r220_c160 bl[160] br[160] wl[220] vdd gnd cell_6t
Xbit_r221_c160 bl[160] br[160] wl[221] vdd gnd cell_6t
Xbit_r222_c160 bl[160] br[160] wl[222] vdd gnd cell_6t
Xbit_r223_c160 bl[160] br[160] wl[223] vdd gnd cell_6t
Xbit_r224_c160 bl[160] br[160] wl[224] vdd gnd cell_6t
Xbit_r225_c160 bl[160] br[160] wl[225] vdd gnd cell_6t
Xbit_r226_c160 bl[160] br[160] wl[226] vdd gnd cell_6t
Xbit_r227_c160 bl[160] br[160] wl[227] vdd gnd cell_6t
Xbit_r228_c160 bl[160] br[160] wl[228] vdd gnd cell_6t
Xbit_r229_c160 bl[160] br[160] wl[229] vdd gnd cell_6t
Xbit_r230_c160 bl[160] br[160] wl[230] vdd gnd cell_6t
Xbit_r231_c160 bl[160] br[160] wl[231] vdd gnd cell_6t
Xbit_r232_c160 bl[160] br[160] wl[232] vdd gnd cell_6t
Xbit_r233_c160 bl[160] br[160] wl[233] vdd gnd cell_6t
Xbit_r234_c160 bl[160] br[160] wl[234] vdd gnd cell_6t
Xbit_r235_c160 bl[160] br[160] wl[235] vdd gnd cell_6t
Xbit_r236_c160 bl[160] br[160] wl[236] vdd gnd cell_6t
Xbit_r237_c160 bl[160] br[160] wl[237] vdd gnd cell_6t
Xbit_r238_c160 bl[160] br[160] wl[238] vdd gnd cell_6t
Xbit_r239_c160 bl[160] br[160] wl[239] vdd gnd cell_6t
Xbit_r240_c160 bl[160] br[160] wl[240] vdd gnd cell_6t
Xbit_r241_c160 bl[160] br[160] wl[241] vdd gnd cell_6t
Xbit_r242_c160 bl[160] br[160] wl[242] vdd gnd cell_6t
Xbit_r243_c160 bl[160] br[160] wl[243] vdd gnd cell_6t
Xbit_r244_c160 bl[160] br[160] wl[244] vdd gnd cell_6t
Xbit_r245_c160 bl[160] br[160] wl[245] vdd gnd cell_6t
Xbit_r246_c160 bl[160] br[160] wl[246] vdd gnd cell_6t
Xbit_r247_c160 bl[160] br[160] wl[247] vdd gnd cell_6t
Xbit_r248_c160 bl[160] br[160] wl[248] vdd gnd cell_6t
Xbit_r249_c160 bl[160] br[160] wl[249] vdd gnd cell_6t
Xbit_r250_c160 bl[160] br[160] wl[250] vdd gnd cell_6t
Xbit_r251_c160 bl[160] br[160] wl[251] vdd gnd cell_6t
Xbit_r252_c160 bl[160] br[160] wl[252] vdd gnd cell_6t
Xbit_r253_c160 bl[160] br[160] wl[253] vdd gnd cell_6t
Xbit_r254_c160 bl[160] br[160] wl[254] vdd gnd cell_6t
Xbit_r255_c160 bl[160] br[160] wl[255] vdd gnd cell_6t
Xbit_r0_c161 bl[161] br[161] wl[0] vdd gnd cell_6t
Xbit_r1_c161 bl[161] br[161] wl[1] vdd gnd cell_6t
Xbit_r2_c161 bl[161] br[161] wl[2] vdd gnd cell_6t
Xbit_r3_c161 bl[161] br[161] wl[3] vdd gnd cell_6t
Xbit_r4_c161 bl[161] br[161] wl[4] vdd gnd cell_6t
Xbit_r5_c161 bl[161] br[161] wl[5] vdd gnd cell_6t
Xbit_r6_c161 bl[161] br[161] wl[6] vdd gnd cell_6t
Xbit_r7_c161 bl[161] br[161] wl[7] vdd gnd cell_6t
Xbit_r8_c161 bl[161] br[161] wl[8] vdd gnd cell_6t
Xbit_r9_c161 bl[161] br[161] wl[9] vdd gnd cell_6t
Xbit_r10_c161 bl[161] br[161] wl[10] vdd gnd cell_6t
Xbit_r11_c161 bl[161] br[161] wl[11] vdd gnd cell_6t
Xbit_r12_c161 bl[161] br[161] wl[12] vdd gnd cell_6t
Xbit_r13_c161 bl[161] br[161] wl[13] vdd gnd cell_6t
Xbit_r14_c161 bl[161] br[161] wl[14] vdd gnd cell_6t
Xbit_r15_c161 bl[161] br[161] wl[15] vdd gnd cell_6t
Xbit_r16_c161 bl[161] br[161] wl[16] vdd gnd cell_6t
Xbit_r17_c161 bl[161] br[161] wl[17] vdd gnd cell_6t
Xbit_r18_c161 bl[161] br[161] wl[18] vdd gnd cell_6t
Xbit_r19_c161 bl[161] br[161] wl[19] vdd gnd cell_6t
Xbit_r20_c161 bl[161] br[161] wl[20] vdd gnd cell_6t
Xbit_r21_c161 bl[161] br[161] wl[21] vdd gnd cell_6t
Xbit_r22_c161 bl[161] br[161] wl[22] vdd gnd cell_6t
Xbit_r23_c161 bl[161] br[161] wl[23] vdd gnd cell_6t
Xbit_r24_c161 bl[161] br[161] wl[24] vdd gnd cell_6t
Xbit_r25_c161 bl[161] br[161] wl[25] vdd gnd cell_6t
Xbit_r26_c161 bl[161] br[161] wl[26] vdd gnd cell_6t
Xbit_r27_c161 bl[161] br[161] wl[27] vdd gnd cell_6t
Xbit_r28_c161 bl[161] br[161] wl[28] vdd gnd cell_6t
Xbit_r29_c161 bl[161] br[161] wl[29] vdd gnd cell_6t
Xbit_r30_c161 bl[161] br[161] wl[30] vdd gnd cell_6t
Xbit_r31_c161 bl[161] br[161] wl[31] vdd gnd cell_6t
Xbit_r32_c161 bl[161] br[161] wl[32] vdd gnd cell_6t
Xbit_r33_c161 bl[161] br[161] wl[33] vdd gnd cell_6t
Xbit_r34_c161 bl[161] br[161] wl[34] vdd gnd cell_6t
Xbit_r35_c161 bl[161] br[161] wl[35] vdd gnd cell_6t
Xbit_r36_c161 bl[161] br[161] wl[36] vdd gnd cell_6t
Xbit_r37_c161 bl[161] br[161] wl[37] vdd gnd cell_6t
Xbit_r38_c161 bl[161] br[161] wl[38] vdd gnd cell_6t
Xbit_r39_c161 bl[161] br[161] wl[39] vdd gnd cell_6t
Xbit_r40_c161 bl[161] br[161] wl[40] vdd gnd cell_6t
Xbit_r41_c161 bl[161] br[161] wl[41] vdd gnd cell_6t
Xbit_r42_c161 bl[161] br[161] wl[42] vdd gnd cell_6t
Xbit_r43_c161 bl[161] br[161] wl[43] vdd gnd cell_6t
Xbit_r44_c161 bl[161] br[161] wl[44] vdd gnd cell_6t
Xbit_r45_c161 bl[161] br[161] wl[45] vdd gnd cell_6t
Xbit_r46_c161 bl[161] br[161] wl[46] vdd gnd cell_6t
Xbit_r47_c161 bl[161] br[161] wl[47] vdd gnd cell_6t
Xbit_r48_c161 bl[161] br[161] wl[48] vdd gnd cell_6t
Xbit_r49_c161 bl[161] br[161] wl[49] vdd gnd cell_6t
Xbit_r50_c161 bl[161] br[161] wl[50] vdd gnd cell_6t
Xbit_r51_c161 bl[161] br[161] wl[51] vdd gnd cell_6t
Xbit_r52_c161 bl[161] br[161] wl[52] vdd gnd cell_6t
Xbit_r53_c161 bl[161] br[161] wl[53] vdd gnd cell_6t
Xbit_r54_c161 bl[161] br[161] wl[54] vdd gnd cell_6t
Xbit_r55_c161 bl[161] br[161] wl[55] vdd gnd cell_6t
Xbit_r56_c161 bl[161] br[161] wl[56] vdd gnd cell_6t
Xbit_r57_c161 bl[161] br[161] wl[57] vdd gnd cell_6t
Xbit_r58_c161 bl[161] br[161] wl[58] vdd gnd cell_6t
Xbit_r59_c161 bl[161] br[161] wl[59] vdd gnd cell_6t
Xbit_r60_c161 bl[161] br[161] wl[60] vdd gnd cell_6t
Xbit_r61_c161 bl[161] br[161] wl[61] vdd gnd cell_6t
Xbit_r62_c161 bl[161] br[161] wl[62] vdd gnd cell_6t
Xbit_r63_c161 bl[161] br[161] wl[63] vdd gnd cell_6t
Xbit_r64_c161 bl[161] br[161] wl[64] vdd gnd cell_6t
Xbit_r65_c161 bl[161] br[161] wl[65] vdd gnd cell_6t
Xbit_r66_c161 bl[161] br[161] wl[66] vdd gnd cell_6t
Xbit_r67_c161 bl[161] br[161] wl[67] vdd gnd cell_6t
Xbit_r68_c161 bl[161] br[161] wl[68] vdd gnd cell_6t
Xbit_r69_c161 bl[161] br[161] wl[69] vdd gnd cell_6t
Xbit_r70_c161 bl[161] br[161] wl[70] vdd gnd cell_6t
Xbit_r71_c161 bl[161] br[161] wl[71] vdd gnd cell_6t
Xbit_r72_c161 bl[161] br[161] wl[72] vdd gnd cell_6t
Xbit_r73_c161 bl[161] br[161] wl[73] vdd gnd cell_6t
Xbit_r74_c161 bl[161] br[161] wl[74] vdd gnd cell_6t
Xbit_r75_c161 bl[161] br[161] wl[75] vdd gnd cell_6t
Xbit_r76_c161 bl[161] br[161] wl[76] vdd gnd cell_6t
Xbit_r77_c161 bl[161] br[161] wl[77] vdd gnd cell_6t
Xbit_r78_c161 bl[161] br[161] wl[78] vdd gnd cell_6t
Xbit_r79_c161 bl[161] br[161] wl[79] vdd gnd cell_6t
Xbit_r80_c161 bl[161] br[161] wl[80] vdd gnd cell_6t
Xbit_r81_c161 bl[161] br[161] wl[81] vdd gnd cell_6t
Xbit_r82_c161 bl[161] br[161] wl[82] vdd gnd cell_6t
Xbit_r83_c161 bl[161] br[161] wl[83] vdd gnd cell_6t
Xbit_r84_c161 bl[161] br[161] wl[84] vdd gnd cell_6t
Xbit_r85_c161 bl[161] br[161] wl[85] vdd gnd cell_6t
Xbit_r86_c161 bl[161] br[161] wl[86] vdd gnd cell_6t
Xbit_r87_c161 bl[161] br[161] wl[87] vdd gnd cell_6t
Xbit_r88_c161 bl[161] br[161] wl[88] vdd gnd cell_6t
Xbit_r89_c161 bl[161] br[161] wl[89] vdd gnd cell_6t
Xbit_r90_c161 bl[161] br[161] wl[90] vdd gnd cell_6t
Xbit_r91_c161 bl[161] br[161] wl[91] vdd gnd cell_6t
Xbit_r92_c161 bl[161] br[161] wl[92] vdd gnd cell_6t
Xbit_r93_c161 bl[161] br[161] wl[93] vdd gnd cell_6t
Xbit_r94_c161 bl[161] br[161] wl[94] vdd gnd cell_6t
Xbit_r95_c161 bl[161] br[161] wl[95] vdd gnd cell_6t
Xbit_r96_c161 bl[161] br[161] wl[96] vdd gnd cell_6t
Xbit_r97_c161 bl[161] br[161] wl[97] vdd gnd cell_6t
Xbit_r98_c161 bl[161] br[161] wl[98] vdd gnd cell_6t
Xbit_r99_c161 bl[161] br[161] wl[99] vdd gnd cell_6t
Xbit_r100_c161 bl[161] br[161] wl[100] vdd gnd cell_6t
Xbit_r101_c161 bl[161] br[161] wl[101] vdd gnd cell_6t
Xbit_r102_c161 bl[161] br[161] wl[102] vdd gnd cell_6t
Xbit_r103_c161 bl[161] br[161] wl[103] vdd gnd cell_6t
Xbit_r104_c161 bl[161] br[161] wl[104] vdd gnd cell_6t
Xbit_r105_c161 bl[161] br[161] wl[105] vdd gnd cell_6t
Xbit_r106_c161 bl[161] br[161] wl[106] vdd gnd cell_6t
Xbit_r107_c161 bl[161] br[161] wl[107] vdd gnd cell_6t
Xbit_r108_c161 bl[161] br[161] wl[108] vdd gnd cell_6t
Xbit_r109_c161 bl[161] br[161] wl[109] vdd gnd cell_6t
Xbit_r110_c161 bl[161] br[161] wl[110] vdd gnd cell_6t
Xbit_r111_c161 bl[161] br[161] wl[111] vdd gnd cell_6t
Xbit_r112_c161 bl[161] br[161] wl[112] vdd gnd cell_6t
Xbit_r113_c161 bl[161] br[161] wl[113] vdd gnd cell_6t
Xbit_r114_c161 bl[161] br[161] wl[114] vdd gnd cell_6t
Xbit_r115_c161 bl[161] br[161] wl[115] vdd gnd cell_6t
Xbit_r116_c161 bl[161] br[161] wl[116] vdd gnd cell_6t
Xbit_r117_c161 bl[161] br[161] wl[117] vdd gnd cell_6t
Xbit_r118_c161 bl[161] br[161] wl[118] vdd gnd cell_6t
Xbit_r119_c161 bl[161] br[161] wl[119] vdd gnd cell_6t
Xbit_r120_c161 bl[161] br[161] wl[120] vdd gnd cell_6t
Xbit_r121_c161 bl[161] br[161] wl[121] vdd gnd cell_6t
Xbit_r122_c161 bl[161] br[161] wl[122] vdd gnd cell_6t
Xbit_r123_c161 bl[161] br[161] wl[123] vdd gnd cell_6t
Xbit_r124_c161 bl[161] br[161] wl[124] vdd gnd cell_6t
Xbit_r125_c161 bl[161] br[161] wl[125] vdd gnd cell_6t
Xbit_r126_c161 bl[161] br[161] wl[126] vdd gnd cell_6t
Xbit_r127_c161 bl[161] br[161] wl[127] vdd gnd cell_6t
Xbit_r128_c161 bl[161] br[161] wl[128] vdd gnd cell_6t
Xbit_r129_c161 bl[161] br[161] wl[129] vdd gnd cell_6t
Xbit_r130_c161 bl[161] br[161] wl[130] vdd gnd cell_6t
Xbit_r131_c161 bl[161] br[161] wl[131] vdd gnd cell_6t
Xbit_r132_c161 bl[161] br[161] wl[132] vdd gnd cell_6t
Xbit_r133_c161 bl[161] br[161] wl[133] vdd gnd cell_6t
Xbit_r134_c161 bl[161] br[161] wl[134] vdd gnd cell_6t
Xbit_r135_c161 bl[161] br[161] wl[135] vdd gnd cell_6t
Xbit_r136_c161 bl[161] br[161] wl[136] vdd gnd cell_6t
Xbit_r137_c161 bl[161] br[161] wl[137] vdd gnd cell_6t
Xbit_r138_c161 bl[161] br[161] wl[138] vdd gnd cell_6t
Xbit_r139_c161 bl[161] br[161] wl[139] vdd gnd cell_6t
Xbit_r140_c161 bl[161] br[161] wl[140] vdd gnd cell_6t
Xbit_r141_c161 bl[161] br[161] wl[141] vdd gnd cell_6t
Xbit_r142_c161 bl[161] br[161] wl[142] vdd gnd cell_6t
Xbit_r143_c161 bl[161] br[161] wl[143] vdd gnd cell_6t
Xbit_r144_c161 bl[161] br[161] wl[144] vdd gnd cell_6t
Xbit_r145_c161 bl[161] br[161] wl[145] vdd gnd cell_6t
Xbit_r146_c161 bl[161] br[161] wl[146] vdd gnd cell_6t
Xbit_r147_c161 bl[161] br[161] wl[147] vdd gnd cell_6t
Xbit_r148_c161 bl[161] br[161] wl[148] vdd gnd cell_6t
Xbit_r149_c161 bl[161] br[161] wl[149] vdd gnd cell_6t
Xbit_r150_c161 bl[161] br[161] wl[150] vdd gnd cell_6t
Xbit_r151_c161 bl[161] br[161] wl[151] vdd gnd cell_6t
Xbit_r152_c161 bl[161] br[161] wl[152] vdd gnd cell_6t
Xbit_r153_c161 bl[161] br[161] wl[153] vdd gnd cell_6t
Xbit_r154_c161 bl[161] br[161] wl[154] vdd gnd cell_6t
Xbit_r155_c161 bl[161] br[161] wl[155] vdd gnd cell_6t
Xbit_r156_c161 bl[161] br[161] wl[156] vdd gnd cell_6t
Xbit_r157_c161 bl[161] br[161] wl[157] vdd gnd cell_6t
Xbit_r158_c161 bl[161] br[161] wl[158] vdd gnd cell_6t
Xbit_r159_c161 bl[161] br[161] wl[159] vdd gnd cell_6t
Xbit_r160_c161 bl[161] br[161] wl[160] vdd gnd cell_6t
Xbit_r161_c161 bl[161] br[161] wl[161] vdd gnd cell_6t
Xbit_r162_c161 bl[161] br[161] wl[162] vdd gnd cell_6t
Xbit_r163_c161 bl[161] br[161] wl[163] vdd gnd cell_6t
Xbit_r164_c161 bl[161] br[161] wl[164] vdd gnd cell_6t
Xbit_r165_c161 bl[161] br[161] wl[165] vdd gnd cell_6t
Xbit_r166_c161 bl[161] br[161] wl[166] vdd gnd cell_6t
Xbit_r167_c161 bl[161] br[161] wl[167] vdd gnd cell_6t
Xbit_r168_c161 bl[161] br[161] wl[168] vdd gnd cell_6t
Xbit_r169_c161 bl[161] br[161] wl[169] vdd gnd cell_6t
Xbit_r170_c161 bl[161] br[161] wl[170] vdd gnd cell_6t
Xbit_r171_c161 bl[161] br[161] wl[171] vdd gnd cell_6t
Xbit_r172_c161 bl[161] br[161] wl[172] vdd gnd cell_6t
Xbit_r173_c161 bl[161] br[161] wl[173] vdd gnd cell_6t
Xbit_r174_c161 bl[161] br[161] wl[174] vdd gnd cell_6t
Xbit_r175_c161 bl[161] br[161] wl[175] vdd gnd cell_6t
Xbit_r176_c161 bl[161] br[161] wl[176] vdd gnd cell_6t
Xbit_r177_c161 bl[161] br[161] wl[177] vdd gnd cell_6t
Xbit_r178_c161 bl[161] br[161] wl[178] vdd gnd cell_6t
Xbit_r179_c161 bl[161] br[161] wl[179] vdd gnd cell_6t
Xbit_r180_c161 bl[161] br[161] wl[180] vdd gnd cell_6t
Xbit_r181_c161 bl[161] br[161] wl[181] vdd gnd cell_6t
Xbit_r182_c161 bl[161] br[161] wl[182] vdd gnd cell_6t
Xbit_r183_c161 bl[161] br[161] wl[183] vdd gnd cell_6t
Xbit_r184_c161 bl[161] br[161] wl[184] vdd gnd cell_6t
Xbit_r185_c161 bl[161] br[161] wl[185] vdd gnd cell_6t
Xbit_r186_c161 bl[161] br[161] wl[186] vdd gnd cell_6t
Xbit_r187_c161 bl[161] br[161] wl[187] vdd gnd cell_6t
Xbit_r188_c161 bl[161] br[161] wl[188] vdd gnd cell_6t
Xbit_r189_c161 bl[161] br[161] wl[189] vdd gnd cell_6t
Xbit_r190_c161 bl[161] br[161] wl[190] vdd gnd cell_6t
Xbit_r191_c161 bl[161] br[161] wl[191] vdd gnd cell_6t
Xbit_r192_c161 bl[161] br[161] wl[192] vdd gnd cell_6t
Xbit_r193_c161 bl[161] br[161] wl[193] vdd gnd cell_6t
Xbit_r194_c161 bl[161] br[161] wl[194] vdd gnd cell_6t
Xbit_r195_c161 bl[161] br[161] wl[195] vdd gnd cell_6t
Xbit_r196_c161 bl[161] br[161] wl[196] vdd gnd cell_6t
Xbit_r197_c161 bl[161] br[161] wl[197] vdd gnd cell_6t
Xbit_r198_c161 bl[161] br[161] wl[198] vdd gnd cell_6t
Xbit_r199_c161 bl[161] br[161] wl[199] vdd gnd cell_6t
Xbit_r200_c161 bl[161] br[161] wl[200] vdd gnd cell_6t
Xbit_r201_c161 bl[161] br[161] wl[201] vdd gnd cell_6t
Xbit_r202_c161 bl[161] br[161] wl[202] vdd gnd cell_6t
Xbit_r203_c161 bl[161] br[161] wl[203] vdd gnd cell_6t
Xbit_r204_c161 bl[161] br[161] wl[204] vdd gnd cell_6t
Xbit_r205_c161 bl[161] br[161] wl[205] vdd gnd cell_6t
Xbit_r206_c161 bl[161] br[161] wl[206] vdd gnd cell_6t
Xbit_r207_c161 bl[161] br[161] wl[207] vdd gnd cell_6t
Xbit_r208_c161 bl[161] br[161] wl[208] vdd gnd cell_6t
Xbit_r209_c161 bl[161] br[161] wl[209] vdd gnd cell_6t
Xbit_r210_c161 bl[161] br[161] wl[210] vdd gnd cell_6t
Xbit_r211_c161 bl[161] br[161] wl[211] vdd gnd cell_6t
Xbit_r212_c161 bl[161] br[161] wl[212] vdd gnd cell_6t
Xbit_r213_c161 bl[161] br[161] wl[213] vdd gnd cell_6t
Xbit_r214_c161 bl[161] br[161] wl[214] vdd gnd cell_6t
Xbit_r215_c161 bl[161] br[161] wl[215] vdd gnd cell_6t
Xbit_r216_c161 bl[161] br[161] wl[216] vdd gnd cell_6t
Xbit_r217_c161 bl[161] br[161] wl[217] vdd gnd cell_6t
Xbit_r218_c161 bl[161] br[161] wl[218] vdd gnd cell_6t
Xbit_r219_c161 bl[161] br[161] wl[219] vdd gnd cell_6t
Xbit_r220_c161 bl[161] br[161] wl[220] vdd gnd cell_6t
Xbit_r221_c161 bl[161] br[161] wl[221] vdd gnd cell_6t
Xbit_r222_c161 bl[161] br[161] wl[222] vdd gnd cell_6t
Xbit_r223_c161 bl[161] br[161] wl[223] vdd gnd cell_6t
Xbit_r224_c161 bl[161] br[161] wl[224] vdd gnd cell_6t
Xbit_r225_c161 bl[161] br[161] wl[225] vdd gnd cell_6t
Xbit_r226_c161 bl[161] br[161] wl[226] vdd gnd cell_6t
Xbit_r227_c161 bl[161] br[161] wl[227] vdd gnd cell_6t
Xbit_r228_c161 bl[161] br[161] wl[228] vdd gnd cell_6t
Xbit_r229_c161 bl[161] br[161] wl[229] vdd gnd cell_6t
Xbit_r230_c161 bl[161] br[161] wl[230] vdd gnd cell_6t
Xbit_r231_c161 bl[161] br[161] wl[231] vdd gnd cell_6t
Xbit_r232_c161 bl[161] br[161] wl[232] vdd gnd cell_6t
Xbit_r233_c161 bl[161] br[161] wl[233] vdd gnd cell_6t
Xbit_r234_c161 bl[161] br[161] wl[234] vdd gnd cell_6t
Xbit_r235_c161 bl[161] br[161] wl[235] vdd gnd cell_6t
Xbit_r236_c161 bl[161] br[161] wl[236] vdd gnd cell_6t
Xbit_r237_c161 bl[161] br[161] wl[237] vdd gnd cell_6t
Xbit_r238_c161 bl[161] br[161] wl[238] vdd gnd cell_6t
Xbit_r239_c161 bl[161] br[161] wl[239] vdd gnd cell_6t
Xbit_r240_c161 bl[161] br[161] wl[240] vdd gnd cell_6t
Xbit_r241_c161 bl[161] br[161] wl[241] vdd gnd cell_6t
Xbit_r242_c161 bl[161] br[161] wl[242] vdd gnd cell_6t
Xbit_r243_c161 bl[161] br[161] wl[243] vdd gnd cell_6t
Xbit_r244_c161 bl[161] br[161] wl[244] vdd gnd cell_6t
Xbit_r245_c161 bl[161] br[161] wl[245] vdd gnd cell_6t
Xbit_r246_c161 bl[161] br[161] wl[246] vdd gnd cell_6t
Xbit_r247_c161 bl[161] br[161] wl[247] vdd gnd cell_6t
Xbit_r248_c161 bl[161] br[161] wl[248] vdd gnd cell_6t
Xbit_r249_c161 bl[161] br[161] wl[249] vdd gnd cell_6t
Xbit_r250_c161 bl[161] br[161] wl[250] vdd gnd cell_6t
Xbit_r251_c161 bl[161] br[161] wl[251] vdd gnd cell_6t
Xbit_r252_c161 bl[161] br[161] wl[252] vdd gnd cell_6t
Xbit_r253_c161 bl[161] br[161] wl[253] vdd gnd cell_6t
Xbit_r254_c161 bl[161] br[161] wl[254] vdd gnd cell_6t
Xbit_r255_c161 bl[161] br[161] wl[255] vdd gnd cell_6t
Xbit_r0_c162 bl[162] br[162] wl[0] vdd gnd cell_6t
Xbit_r1_c162 bl[162] br[162] wl[1] vdd gnd cell_6t
Xbit_r2_c162 bl[162] br[162] wl[2] vdd gnd cell_6t
Xbit_r3_c162 bl[162] br[162] wl[3] vdd gnd cell_6t
Xbit_r4_c162 bl[162] br[162] wl[4] vdd gnd cell_6t
Xbit_r5_c162 bl[162] br[162] wl[5] vdd gnd cell_6t
Xbit_r6_c162 bl[162] br[162] wl[6] vdd gnd cell_6t
Xbit_r7_c162 bl[162] br[162] wl[7] vdd gnd cell_6t
Xbit_r8_c162 bl[162] br[162] wl[8] vdd gnd cell_6t
Xbit_r9_c162 bl[162] br[162] wl[9] vdd gnd cell_6t
Xbit_r10_c162 bl[162] br[162] wl[10] vdd gnd cell_6t
Xbit_r11_c162 bl[162] br[162] wl[11] vdd gnd cell_6t
Xbit_r12_c162 bl[162] br[162] wl[12] vdd gnd cell_6t
Xbit_r13_c162 bl[162] br[162] wl[13] vdd gnd cell_6t
Xbit_r14_c162 bl[162] br[162] wl[14] vdd gnd cell_6t
Xbit_r15_c162 bl[162] br[162] wl[15] vdd gnd cell_6t
Xbit_r16_c162 bl[162] br[162] wl[16] vdd gnd cell_6t
Xbit_r17_c162 bl[162] br[162] wl[17] vdd gnd cell_6t
Xbit_r18_c162 bl[162] br[162] wl[18] vdd gnd cell_6t
Xbit_r19_c162 bl[162] br[162] wl[19] vdd gnd cell_6t
Xbit_r20_c162 bl[162] br[162] wl[20] vdd gnd cell_6t
Xbit_r21_c162 bl[162] br[162] wl[21] vdd gnd cell_6t
Xbit_r22_c162 bl[162] br[162] wl[22] vdd gnd cell_6t
Xbit_r23_c162 bl[162] br[162] wl[23] vdd gnd cell_6t
Xbit_r24_c162 bl[162] br[162] wl[24] vdd gnd cell_6t
Xbit_r25_c162 bl[162] br[162] wl[25] vdd gnd cell_6t
Xbit_r26_c162 bl[162] br[162] wl[26] vdd gnd cell_6t
Xbit_r27_c162 bl[162] br[162] wl[27] vdd gnd cell_6t
Xbit_r28_c162 bl[162] br[162] wl[28] vdd gnd cell_6t
Xbit_r29_c162 bl[162] br[162] wl[29] vdd gnd cell_6t
Xbit_r30_c162 bl[162] br[162] wl[30] vdd gnd cell_6t
Xbit_r31_c162 bl[162] br[162] wl[31] vdd gnd cell_6t
Xbit_r32_c162 bl[162] br[162] wl[32] vdd gnd cell_6t
Xbit_r33_c162 bl[162] br[162] wl[33] vdd gnd cell_6t
Xbit_r34_c162 bl[162] br[162] wl[34] vdd gnd cell_6t
Xbit_r35_c162 bl[162] br[162] wl[35] vdd gnd cell_6t
Xbit_r36_c162 bl[162] br[162] wl[36] vdd gnd cell_6t
Xbit_r37_c162 bl[162] br[162] wl[37] vdd gnd cell_6t
Xbit_r38_c162 bl[162] br[162] wl[38] vdd gnd cell_6t
Xbit_r39_c162 bl[162] br[162] wl[39] vdd gnd cell_6t
Xbit_r40_c162 bl[162] br[162] wl[40] vdd gnd cell_6t
Xbit_r41_c162 bl[162] br[162] wl[41] vdd gnd cell_6t
Xbit_r42_c162 bl[162] br[162] wl[42] vdd gnd cell_6t
Xbit_r43_c162 bl[162] br[162] wl[43] vdd gnd cell_6t
Xbit_r44_c162 bl[162] br[162] wl[44] vdd gnd cell_6t
Xbit_r45_c162 bl[162] br[162] wl[45] vdd gnd cell_6t
Xbit_r46_c162 bl[162] br[162] wl[46] vdd gnd cell_6t
Xbit_r47_c162 bl[162] br[162] wl[47] vdd gnd cell_6t
Xbit_r48_c162 bl[162] br[162] wl[48] vdd gnd cell_6t
Xbit_r49_c162 bl[162] br[162] wl[49] vdd gnd cell_6t
Xbit_r50_c162 bl[162] br[162] wl[50] vdd gnd cell_6t
Xbit_r51_c162 bl[162] br[162] wl[51] vdd gnd cell_6t
Xbit_r52_c162 bl[162] br[162] wl[52] vdd gnd cell_6t
Xbit_r53_c162 bl[162] br[162] wl[53] vdd gnd cell_6t
Xbit_r54_c162 bl[162] br[162] wl[54] vdd gnd cell_6t
Xbit_r55_c162 bl[162] br[162] wl[55] vdd gnd cell_6t
Xbit_r56_c162 bl[162] br[162] wl[56] vdd gnd cell_6t
Xbit_r57_c162 bl[162] br[162] wl[57] vdd gnd cell_6t
Xbit_r58_c162 bl[162] br[162] wl[58] vdd gnd cell_6t
Xbit_r59_c162 bl[162] br[162] wl[59] vdd gnd cell_6t
Xbit_r60_c162 bl[162] br[162] wl[60] vdd gnd cell_6t
Xbit_r61_c162 bl[162] br[162] wl[61] vdd gnd cell_6t
Xbit_r62_c162 bl[162] br[162] wl[62] vdd gnd cell_6t
Xbit_r63_c162 bl[162] br[162] wl[63] vdd gnd cell_6t
Xbit_r64_c162 bl[162] br[162] wl[64] vdd gnd cell_6t
Xbit_r65_c162 bl[162] br[162] wl[65] vdd gnd cell_6t
Xbit_r66_c162 bl[162] br[162] wl[66] vdd gnd cell_6t
Xbit_r67_c162 bl[162] br[162] wl[67] vdd gnd cell_6t
Xbit_r68_c162 bl[162] br[162] wl[68] vdd gnd cell_6t
Xbit_r69_c162 bl[162] br[162] wl[69] vdd gnd cell_6t
Xbit_r70_c162 bl[162] br[162] wl[70] vdd gnd cell_6t
Xbit_r71_c162 bl[162] br[162] wl[71] vdd gnd cell_6t
Xbit_r72_c162 bl[162] br[162] wl[72] vdd gnd cell_6t
Xbit_r73_c162 bl[162] br[162] wl[73] vdd gnd cell_6t
Xbit_r74_c162 bl[162] br[162] wl[74] vdd gnd cell_6t
Xbit_r75_c162 bl[162] br[162] wl[75] vdd gnd cell_6t
Xbit_r76_c162 bl[162] br[162] wl[76] vdd gnd cell_6t
Xbit_r77_c162 bl[162] br[162] wl[77] vdd gnd cell_6t
Xbit_r78_c162 bl[162] br[162] wl[78] vdd gnd cell_6t
Xbit_r79_c162 bl[162] br[162] wl[79] vdd gnd cell_6t
Xbit_r80_c162 bl[162] br[162] wl[80] vdd gnd cell_6t
Xbit_r81_c162 bl[162] br[162] wl[81] vdd gnd cell_6t
Xbit_r82_c162 bl[162] br[162] wl[82] vdd gnd cell_6t
Xbit_r83_c162 bl[162] br[162] wl[83] vdd gnd cell_6t
Xbit_r84_c162 bl[162] br[162] wl[84] vdd gnd cell_6t
Xbit_r85_c162 bl[162] br[162] wl[85] vdd gnd cell_6t
Xbit_r86_c162 bl[162] br[162] wl[86] vdd gnd cell_6t
Xbit_r87_c162 bl[162] br[162] wl[87] vdd gnd cell_6t
Xbit_r88_c162 bl[162] br[162] wl[88] vdd gnd cell_6t
Xbit_r89_c162 bl[162] br[162] wl[89] vdd gnd cell_6t
Xbit_r90_c162 bl[162] br[162] wl[90] vdd gnd cell_6t
Xbit_r91_c162 bl[162] br[162] wl[91] vdd gnd cell_6t
Xbit_r92_c162 bl[162] br[162] wl[92] vdd gnd cell_6t
Xbit_r93_c162 bl[162] br[162] wl[93] vdd gnd cell_6t
Xbit_r94_c162 bl[162] br[162] wl[94] vdd gnd cell_6t
Xbit_r95_c162 bl[162] br[162] wl[95] vdd gnd cell_6t
Xbit_r96_c162 bl[162] br[162] wl[96] vdd gnd cell_6t
Xbit_r97_c162 bl[162] br[162] wl[97] vdd gnd cell_6t
Xbit_r98_c162 bl[162] br[162] wl[98] vdd gnd cell_6t
Xbit_r99_c162 bl[162] br[162] wl[99] vdd gnd cell_6t
Xbit_r100_c162 bl[162] br[162] wl[100] vdd gnd cell_6t
Xbit_r101_c162 bl[162] br[162] wl[101] vdd gnd cell_6t
Xbit_r102_c162 bl[162] br[162] wl[102] vdd gnd cell_6t
Xbit_r103_c162 bl[162] br[162] wl[103] vdd gnd cell_6t
Xbit_r104_c162 bl[162] br[162] wl[104] vdd gnd cell_6t
Xbit_r105_c162 bl[162] br[162] wl[105] vdd gnd cell_6t
Xbit_r106_c162 bl[162] br[162] wl[106] vdd gnd cell_6t
Xbit_r107_c162 bl[162] br[162] wl[107] vdd gnd cell_6t
Xbit_r108_c162 bl[162] br[162] wl[108] vdd gnd cell_6t
Xbit_r109_c162 bl[162] br[162] wl[109] vdd gnd cell_6t
Xbit_r110_c162 bl[162] br[162] wl[110] vdd gnd cell_6t
Xbit_r111_c162 bl[162] br[162] wl[111] vdd gnd cell_6t
Xbit_r112_c162 bl[162] br[162] wl[112] vdd gnd cell_6t
Xbit_r113_c162 bl[162] br[162] wl[113] vdd gnd cell_6t
Xbit_r114_c162 bl[162] br[162] wl[114] vdd gnd cell_6t
Xbit_r115_c162 bl[162] br[162] wl[115] vdd gnd cell_6t
Xbit_r116_c162 bl[162] br[162] wl[116] vdd gnd cell_6t
Xbit_r117_c162 bl[162] br[162] wl[117] vdd gnd cell_6t
Xbit_r118_c162 bl[162] br[162] wl[118] vdd gnd cell_6t
Xbit_r119_c162 bl[162] br[162] wl[119] vdd gnd cell_6t
Xbit_r120_c162 bl[162] br[162] wl[120] vdd gnd cell_6t
Xbit_r121_c162 bl[162] br[162] wl[121] vdd gnd cell_6t
Xbit_r122_c162 bl[162] br[162] wl[122] vdd gnd cell_6t
Xbit_r123_c162 bl[162] br[162] wl[123] vdd gnd cell_6t
Xbit_r124_c162 bl[162] br[162] wl[124] vdd gnd cell_6t
Xbit_r125_c162 bl[162] br[162] wl[125] vdd gnd cell_6t
Xbit_r126_c162 bl[162] br[162] wl[126] vdd gnd cell_6t
Xbit_r127_c162 bl[162] br[162] wl[127] vdd gnd cell_6t
Xbit_r128_c162 bl[162] br[162] wl[128] vdd gnd cell_6t
Xbit_r129_c162 bl[162] br[162] wl[129] vdd gnd cell_6t
Xbit_r130_c162 bl[162] br[162] wl[130] vdd gnd cell_6t
Xbit_r131_c162 bl[162] br[162] wl[131] vdd gnd cell_6t
Xbit_r132_c162 bl[162] br[162] wl[132] vdd gnd cell_6t
Xbit_r133_c162 bl[162] br[162] wl[133] vdd gnd cell_6t
Xbit_r134_c162 bl[162] br[162] wl[134] vdd gnd cell_6t
Xbit_r135_c162 bl[162] br[162] wl[135] vdd gnd cell_6t
Xbit_r136_c162 bl[162] br[162] wl[136] vdd gnd cell_6t
Xbit_r137_c162 bl[162] br[162] wl[137] vdd gnd cell_6t
Xbit_r138_c162 bl[162] br[162] wl[138] vdd gnd cell_6t
Xbit_r139_c162 bl[162] br[162] wl[139] vdd gnd cell_6t
Xbit_r140_c162 bl[162] br[162] wl[140] vdd gnd cell_6t
Xbit_r141_c162 bl[162] br[162] wl[141] vdd gnd cell_6t
Xbit_r142_c162 bl[162] br[162] wl[142] vdd gnd cell_6t
Xbit_r143_c162 bl[162] br[162] wl[143] vdd gnd cell_6t
Xbit_r144_c162 bl[162] br[162] wl[144] vdd gnd cell_6t
Xbit_r145_c162 bl[162] br[162] wl[145] vdd gnd cell_6t
Xbit_r146_c162 bl[162] br[162] wl[146] vdd gnd cell_6t
Xbit_r147_c162 bl[162] br[162] wl[147] vdd gnd cell_6t
Xbit_r148_c162 bl[162] br[162] wl[148] vdd gnd cell_6t
Xbit_r149_c162 bl[162] br[162] wl[149] vdd gnd cell_6t
Xbit_r150_c162 bl[162] br[162] wl[150] vdd gnd cell_6t
Xbit_r151_c162 bl[162] br[162] wl[151] vdd gnd cell_6t
Xbit_r152_c162 bl[162] br[162] wl[152] vdd gnd cell_6t
Xbit_r153_c162 bl[162] br[162] wl[153] vdd gnd cell_6t
Xbit_r154_c162 bl[162] br[162] wl[154] vdd gnd cell_6t
Xbit_r155_c162 bl[162] br[162] wl[155] vdd gnd cell_6t
Xbit_r156_c162 bl[162] br[162] wl[156] vdd gnd cell_6t
Xbit_r157_c162 bl[162] br[162] wl[157] vdd gnd cell_6t
Xbit_r158_c162 bl[162] br[162] wl[158] vdd gnd cell_6t
Xbit_r159_c162 bl[162] br[162] wl[159] vdd gnd cell_6t
Xbit_r160_c162 bl[162] br[162] wl[160] vdd gnd cell_6t
Xbit_r161_c162 bl[162] br[162] wl[161] vdd gnd cell_6t
Xbit_r162_c162 bl[162] br[162] wl[162] vdd gnd cell_6t
Xbit_r163_c162 bl[162] br[162] wl[163] vdd gnd cell_6t
Xbit_r164_c162 bl[162] br[162] wl[164] vdd gnd cell_6t
Xbit_r165_c162 bl[162] br[162] wl[165] vdd gnd cell_6t
Xbit_r166_c162 bl[162] br[162] wl[166] vdd gnd cell_6t
Xbit_r167_c162 bl[162] br[162] wl[167] vdd gnd cell_6t
Xbit_r168_c162 bl[162] br[162] wl[168] vdd gnd cell_6t
Xbit_r169_c162 bl[162] br[162] wl[169] vdd gnd cell_6t
Xbit_r170_c162 bl[162] br[162] wl[170] vdd gnd cell_6t
Xbit_r171_c162 bl[162] br[162] wl[171] vdd gnd cell_6t
Xbit_r172_c162 bl[162] br[162] wl[172] vdd gnd cell_6t
Xbit_r173_c162 bl[162] br[162] wl[173] vdd gnd cell_6t
Xbit_r174_c162 bl[162] br[162] wl[174] vdd gnd cell_6t
Xbit_r175_c162 bl[162] br[162] wl[175] vdd gnd cell_6t
Xbit_r176_c162 bl[162] br[162] wl[176] vdd gnd cell_6t
Xbit_r177_c162 bl[162] br[162] wl[177] vdd gnd cell_6t
Xbit_r178_c162 bl[162] br[162] wl[178] vdd gnd cell_6t
Xbit_r179_c162 bl[162] br[162] wl[179] vdd gnd cell_6t
Xbit_r180_c162 bl[162] br[162] wl[180] vdd gnd cell_6t
Xbit_r181_c162 bl[162] br[162] wl[181] vdd gnd cell_6t
Xbit_r182_c162 bl[162] br[162] wl[182] vdd gnd cell_6t
Xbit_r183_c162 bl[162] br[162] wl[183] vdd gnd cell_6t
Xbit_r184_c162 bl[162] br[162] wl[184] vdd gnd cell_6t
Xbit_r185_c162 bl[162] br[162] wl[185] vdd gnd cell_6t
Xbit_r186_c162 bl[162] br[162] wl[186] vdd gnd cell_6t
Xbit_r187_c162 bl[162] br[162] wl[187] vdd gnd cell_6t
Xbit_r188_c162 bl[162] br[162] wl[188] vdd gnd cell_6t
Xbit_r189_c162 bl[162] br[162] wl[189] vdd gnd cell_6t
Xbit_r190_c162 bl[162] br[162] wl[190] vdd gnd cell_6t
Xbit_r191_c162 bl[162] br[162] wl[191] vdd gnd cell_6t
Xbit_r192_c162 bl[162] br[162] wl[192] vdd gnd cell_6t
Xbit_r193_c162 bl[162] br[162] wl[193] vdd gnd cell_6t
Xbit_r194_c162 bl[162] br[162] wl[194] vdd gnd cell_6t
Xbit_r195_c162 bl[162] br[162] wl[195] vdd gnd cell_6t
Xbit_r196_c162 bl[162] br[162] wl[196] vdd gnd cell_6t
Xbit_r197_c162 bl[162] br[162] wl[197] vdd gnd cell_6t
Xbit_r198_c162 bl[162] br[162] wl[198] vdd gnd cell_6t
Xbit_r199_c162 bl[162] br[162] wl[199] vdd gnd cell_6t
Xbit_r200_c162 bl[162] br[162] wl[200] vdd gnd cell_6t
Xbit_r201_c162 bl[162] br[162] wl[201] vdd gnd cell_6t
Xbit_r202_c162 bl[162] br[162] wl[202] vdd gnd cell_6t
Xbit_r203_c162 bl[162] br[162] wl[203] vdd gnd cell_6t
Xbit_r204_c162 bl[162] br[162] wl[204] vdd gnd cell_6t
Xbit_r205_c162 bl[162] br[162] wl[205] vdd gnd cell_6t
Xbit_r206_c162 bl[162] br[162] wl[206] vdd gnd cell_6t
Xbit_r207_c162 bl[162] br[162] wl[207] vdd gnd cell_6t
Xbit_r208_c162 bl[162] br[162] wl[208] vdd gnd cell_6t
Xbit_r209_c162 bl[162] br[162] wl[209] vdd gnd cell_6t
Xbit_r210_c162 bl[162] br[162] wl[210] vdd gnd cell_6t
Xbit_r211_c162 bl[162] br[162] wl[211] vdd gnd cell_6t
Xbit_r212_c162 bl[162] br[162] wl[212] vdd gnd cell_6t
Xbit_r213_c162 bl[162] br[162] wl[213] vdd gnd cell_6t
Xbit_r214_c162 bl[162] br[162] wl[214] vdd gnd cell_6t
Xbit_r215_c162 bl[162] br[162] wl[215] vdd gnd cell_6t
Xbit_r216_c162 bl[162] br[162] wl[216] vdd gnd cell_6t
Xbit_r217_c162 bl[162] br[162] wl[217] vdd gnd cell_6t
Xbit_r218_c162 bl[162] br[162] wl[218] vdd gnd cell_6t
Xbit_r219_c162 bl[162] br[162] wl[219] vdd gnd cell_6t
Xbit_r220_c162 bl[162] br[162] wl[220] vdd gnd cell_6t
Xbit_r221_c162 bl[162] br[162] wl[221] vdd gnd cell_6t
Xbit_r222_c162 bl[162] br[162] wl[222] vdd gnd cell_6t
Xbit_r223_c162 bl[162] br[162] wl[223] vdd gnd cell_6t
Xbit_r224_c162 bl[162] br[162] wl[224] vdd gnd cell_6t
Xbit_r225_c162 bl[162] br[162] wl[225] vdd gnd cell_6t
Xbit_r226_c162 bl[162] br[162] wl[226] vdd gnd cell_6t
Xbit_r227_c162 bl[162] br[162] wl[227] vdd gnd cell_6t
Xbit_r228_c162 bl[162] br[162] wl[228] vdd gnd cell_6t
Xbit_r229_c162 bl[162] br[162] wl[229] vdd gnd cell_6t
Xbit_r230_c162 bl[162] br[162] wl[230] vdd gnd cell_6t
Xbit_r231_c162 bl[162] br[162] wl[231] vdd gnd cell_6t
Xbit_r232_c162 bl[162] br[162] wl[232] vdd gnd cell_6t
Xbit_r233_c162 bl[162] br[162] wl[233] vdd gnd cell_6t
Xbit_r234_c162 bl[162] br[162] wl[234] vdd gnd cell_6t
Xbit_r235_c162 bl[162] br[162] wl[235] vdd gnd cell_6t
Xbit_r236_c162 bl[162] br[162] wl[236] vdd gnd cell_6t
Xbit_r237_c162 bl[162] br[162] wl[237] vdd gnd cell_6t
Xbit_r238_c162 bl[162] br[162] wl[238] vdd gnd cell_6t
Xbit_r239_c162 bl[162] br[162] wl[239] vdd gnd cell_6t
Xbit_r240_c162 bl[162] br[162] wl[240] vdd gnd cell_6t
Xbit_r241_c162 bl[162] br[162] wl[241] vdd gnd cell_6t
Xbit_r242_c162 bl[162] br[162] wl[242] vdd gnd cell_6t
Xbit_r243_c162 bl[162] br[162] wl[243] vdd gnd cell_6t
Xbit_r244_c162 bl[162] br[162] wl[244] vdd gnd cell_6t
Xbit_r245_c162 bl[162] br[162] wl[245] vdd gnd cell_6t
Xbit_r246_c162 bl[162] br[162] wl[246] vdd gnd cell_6t
Xbit_r247_c162 bl[162] br[162] wl[247] vdd gnd cell_6t
Xbit_r248_c162 bl[162] br[162] wl[248] vdd gnd cell_6t
Xbit_r249_c162 bl[162] br[162] wl[249] vdd gnd cell_6t
Xbit_r250_c162 bl[162] br[162] wl[250] vdd gnd cell_6t
Xbit_r251_c162 bl[162] br[162] wl[251] vdd gnd cell_6t
Xbit_r252_c162 bl[162] br[162] wl[252] vdd gnd cell_6t
Xbit_r253_c162 bl[162] br[162] wl[253] vdd gnd cell_6t
Xbit_r254_c162 bl[162] br[162] wl[254] vdd gnd cell_6t
Xbit_r255_c162 bl[162] br[162] wl[255] vdd gnd cell_6t
Xbit_r0_c163 bl[163] br[163] wl[0] vdd gnd cell_6t
Xbit_r1_c163 bl[163] br[163] wl[1] vdd gnd cell_6t
Xbit_r2_c163 bl[163] br[163] wl[2] vdd gnd cell_6t
Xbit_r3_c163 bl[163] br[163] wl[3] vdd gnd cell_6t
Xbit_r4_c163 bl[163] br[163] wl[4] vdd gnd cell_6t
Xbit_r5_c163 bl[163] br[163] wl[5] vdd gnd cell_6t
Xbit_r6_c163 bl[163] br[163] wl[6] vdd gnd cell_6t
Xbit_r7_c163 bl[163] br[163] wl[7] vdd gnd cell_6t
Xbit_r8_c163 bl[163] br[163] wl[8] vdd gnd cell_6t
Xbit_r9_c163 bl[163] br[163] wl[9] vdd gnd cell_6t
Xbit_r10_c163 bl[163] br[163] wl[10] vdd gnd cell_6t
Xbit_r11_c163 bl[163] br[163] wl[11] vdd gnd cell_6t
Xbit_r12_c163 bl[163] br[163] wl[12] vdd gnd cell_6t
Xbit_r13_c163 bl[163] br[163] wl[13] vdd gnd cell_6t
Xbit_r14_c163 bl[163] br[163] wl[14] vdd gnd cell_6t
Xbit_r15_c163 bl[163] br[163] wl[15] vdd gnd cell_6t
Xbit_r16_c163 bl[163] br[163] wl[16] vdd gnd cell_6t
Xbit_r17_c163 bl[163] br[163] wl[17] vdd gnd cell_6t
Xbit_r18_c163 bl[163] br[163] wl[18] vdd gnd cell_6t
Xbit_r19_c163 bl[163] br[163] wl[19] vdd gnd cell_6t
Xbit_r20_c163 bl[163] br[163] wl[20] vdd gnd cell_6t
Xbit_r21_c163 bl[163] br[163] wl[21] vdd gnd cell_6t
Xbit_r22_c163 bl[163] br[163] wl[22] vdd gnd cell_6t
Xbit_r23_c163 bl[163] br[163] wl[23] vdd gnd cell_6t
Xbit_r24_c163 bl[163] br[163] wl[24] vdd gnd cell_6t
Xbit_r25_c163 bl[163] br[163] wl[25] vdd gnd cell_6t
Xbit_r26_c163 bl[163] br[163] wl[26] vdd gnd cell_6t
Xbit_r27_c163 bl[163] br[163] wl[27] vdd gnd cell_6t
Xbit_r28_c163 bl[163] br[163] wl[28] vdd gnd cell_6t
Xbit_r29_c163 bl[163] br[163] wl[29] vdd gnd cell_6t
Xbit_r30_c163 bl[163] br[163] wl[30] vdd gnd cell_6t
Xbit_r31_c163 bl[163] br[163] wl[31] vdd gnd cell_6t
Xbit_r32_c163 bl[163] br[163] wl[32] vdd gnd cell_6t
Xbit_r33_c163 bl[163] br[163] wl[33] vdd gnd cell_6t
Xbit_r34_c163 bl[163] br[163] wl[34] vdd gnd cell_6t
Xbit_r35_c163 bl[163] br[163] wl[35] vdd gnd cell_6t
Xbit_r36_c163 bl[163] br[163] wl[36] vdd gnd cell_6t
Xbit_r37_c163 bl[163] br[163] wl[37] vdd gnd cell_6t
Xbit_r38_c163 bl[163] br[163] wl[38] vdd gnd cell_6t
Xbit_r39_c163 bl[163] br[163] wl[39] vdd gnd cell_6t
Xbit_r40_c163 bl[163] br[163] wl[40] vdd gnd cell_6t
Xbit_r41_c163 bl[163] br[163] wl[41] vdd gnd cell_6t
Xbit_r42_c163 bl[163] br[163] wl[42] vdd gnd cell_6t
Xbit_r43_c163 bl[163] br[163] wl[43] vdd gnd cell_6t
Xbit_r44_c163 bl[163] br[163] wl[44] vdd gnd cell_6t
Xbit_r45_c163 bl[163] br[163] wl[45] vdd gnd cell_6t
Xbit_r46_c163 bl[163] br[163] wl[46] vdd gnd cell_6t
Xbit_r47_c163 bl[163] br[163] wl[47] vdd gnd cell_6t
Xbit_r48_c163 bl[163] br[163] wl[48] vdd gnd cell_6t
Xbit_r49_c163 bl[163] br[163] wl[49] vdd gnd cell_6t
Xbit_r50_c163 bl[163] br[163] wl[50] vdd gnd cell_6t
Xbit_r51_c163 bl[163] br[163] wl[51] vdd gnd cell_6t
Xbit_r52_c163 bl[163] br[163] wl[52] vdd gnd cell_6t
Xbit_r53_c163 bl[163] br[163] wl[53] vdd gnd cell_6t
Xbit_r54_c163 bl[163] br[163] wl[54] vdd gnd cell_6t
Xbit_r55_c163 bl[163] br[163] wl[55] vdd gnd cell_6t
Xbit_r56_c163 bl[163] br[163] wl[56] vdd gnd cell_6t
Xbit_r57_c163 bl[163] br[163] wl[57] vdd gnd cell_6t
Xbit_r58_c163 bl[163] br[163] wl[58] vdd gnd cell_6t
Xbit_r59_c163 bl[163] br[163] wl[59] vdd gnd cell_6t
Xbit_r60_c163 bl[163] br[163] wl[60] vdd gnd cell_6t
Xbit_r61_c163 bl[163] br[163] wl[61] vdd gnd cell_6t
Xbit_r62_c163 bl[163] br[163] wl[62] vdd gnd cell_6t
Xbit_r63_c163 bl[163] br[163] wl[63] vdd gnd cell_6t
Xbit_r64_c163 bl[163] br[163] wl[64] vdd gnd cell_6t
Xbit_r65_c163 bl[163] br[163] wl[65] vdd gnd cell_6t
Xbit_r66_c163 bl[163] br[163] wl[66] vdd gnd cell_6t
Xbit_r67_c163 bl[163] br[163] wl[67] vdd gnd cell_6t
Xbit_r68_c163 bl[163] br[163] wl[68] vdd gnd cell_6t
Xbit_r69_c163 bl[163] br[163] wl[69] vdd gnd cell_6t
Xbit_r70_c163 bl[163] br[163] wl[70] vdd gnd cell_6t
Xbit_r71_c163 bl[163] br[163] wl[71] vdd gnd cell_6t
Xbit_r72_c163 bl[163] br[163] wl[72] vdd gnd cell_6t
Xbit_r73_c163 bl[163] br[163] wl[73] vdd gnd cell_6t
Xbit_r74_c163 bl[163] br[163] wl[74] vdd gnd cell_6t
Xbit_r75_c163 bl[163] br[163] wl[75] vdd gnd cell_6t
Xbit_r76_c163 bl[163] br[163] wl[76] vdd gnd cell_6t
Xbit_r77_c163 bl[163] br[163] wl[77] vdd gnd cell_6t
Xbit_r78_c163 bl[163] br[163] wl[78] vdd gnd cell_6t
Xbit_r79_c163 bl[163] br[163] wl[79] vdd gnd cell_6t
Xbit_r80_c163 bl[163] br[163] wl[80] vdd gnd cell_6t
Xbit_r81_c163 bl[163] br[163] wl[81] vdd gnd cell_6t
Xbit_r82_c163 bl[163] br[163] wl[82] vdd gnd cell_6t
Xbit_r83_c163 bl[163] br[163] wl[83] vdd gnd cell_6t
Xbit_r84_c163 bl[163] br[163] wl[84] vdd gnd cell_6t
Xbit_r85_c163 bl[163] br[163] wl[85] vdd gnd cell_6t
Xbit_r86_c163 bl[163] br[163] wl[86] vdd gnd cell_6t
Xbit_r87_c163 bl[163] br[163] wl[87] vdd gnd cell_6t
Xbit_r88_c163 bl[163] br[163] wl[88] vdd gnd cell_6t
Xbit_r89_c163 bl[163] br[163] wl[89] vdd gnd cell_6t
Xbit_r90_c163 bl[163] br[163] wl[90] vdd gnd cell_6t
Xbit_r91_c163 bl[163] br[163] wl[91] vdd gnd cell_6t
Xbit_r92_c163 bl[163] br[163] wl[92] vdd gnd cell_6t
Xbit_r93_c163 bl[163] br[163] wl[93] vdd gnd cell_6t
Xbit_r94_c163 bl[163] br[163] wl[94] vdd gnd cell_6t
Xbit_r95_c163 bl[163] br[163] wl[95] vdd gnd cell_6t
Xbit_r96_c163 bl[163] br[163] wl[96] vdd gnd cell_6t
Xbit_r97_c163 bl[163] br[163] wl[97] vdd gnd cell_6t
Xbit_r98_c163 bl[163] br[163] wl[98] vdd gnd cell_6t
Xbit_r99_c163 bl[163] br[163] wl[99] vdd gnd cell_6t
Xbit_r100_c163 bl[163] br[163] wl[100] vdd gnd cell_6t
Xbit_r101_c163 bl[163] br[163] wl[101] vdd gnd cell_6t
Xbit_r102_c163 bl[163] br[163] wl[102] vdd gnd cell_6t
Xbit_r103_c163 bl[163] br[163] wl[103] vdd gnd cell_6t
Xbit_r104_c163 bl[163] br[163] wl[104] vdd gnd cell_6t
Xbit_r105_c163 bl[163] br[163] wl[105] vdd gnd cell_6t
Xbit_r106_c163 bl[163] br[163] wl[106] vdd gnd cell_6t
Xbit_r107_c163 bl[163] br[163] wl[107] vdd gnd cell_6t
Xbit_r108_c163 bl[163] br[163] wl[108] vdd gnd cell_6t
Xbit_r109_c163 bl[163] br[163] wl[109] vdd gnd cell_6t
Xbit_r110_c163 bl[163] br[163] wl[110] vdd gnd cell_6t
Xbit_r111_c163 bl[163] br[163] wl[111] vdd gnd cell_6t
Xbit_r112_c163 bl[163] br[163] wl[112] vdd gnd cell_6t
Xbit_r113_c163 bl[163] br[163] wl[113] vdd gnd cell_6t
Xbit_r114_c163 bl[163] br[163] wl[114] vdd gnd cell_6t
Xbit_r115_c163 bl[163] br[163] wl[115] vdd gnd cell_6t
Xbit_r116_c163 bl[163] br[163] wl[116] vdd gnd cell_6t
Xbit_r117_c163 bl[163] br[163] wl[117] vdd gnd cell_6t
Xbit_r118_c163 bl[163] br[163] wl[118] vdd gnd cell_6t
Xbit_r119_c163 bl[163] br[163] wl[119] vdd gnd cell_6t
Xbit_r120_c163 bl[163] br[163] wl[120] vdd gnd cell_6t
Xbit_r121_c163 bl[163] br[163] wl[121] vdd gnd cell_6t
Xbit_r122_c163 bl[163] br[163] wl[122] vdd gnd cell_6t
Xbit_r123_c163 bl[163] br[163] wl[123] vdd gnd cell_6t
Xbit_r124_c163 bl[163] br[163] wl[124] vdd gnd cell_6t
Xbit_r125_c163 bl[163] br[163] wl[125] vdd gnd cell_6t
Xbit_r126_c163 bl[163] br[163] wl[126] vdd gnd cell_6t
Xbit_r127_c163 bl[163] br[163] wl[127] vdd gnd cell_6t
Xbit_r128_c163 bl[163] br[163] wl[128] vdd gnd cell_6t
Xbit_r129_c163 bl[163] br[163] wl[129] vdd gnd cell_6t
Xbit_r130_c163 bl[163] br[163] wl[130] vdd gnd cell_6t
Xbit_r131_c163 bl[163] br[163] wl[131] vdd gnd cell_6t
Xbit_r132_c163 bl[163] br[163] wl[132] vdd gnd cell_6t
Xbit_r133_c163 bl[163] br[163] wl[133] vdd gnd cell_6t
Xbit_r134_c163 bl[163] br[163] wl[134] vdd gnd cell_6t
Xbit_r135_c163 bl[163] br[163] wl[135] vdd gnd cell_6t
Xbit_r136_c163 bl[163] br[163] wl[136] vdd gnd cell_6t
Xbit_r137_c163 bl[163] br[163] wl[137] vdd gnd cell_6t
Xbit_r138_c163 bl[163] br[163] wl[138] vdd gnd cell_6t
Xbit_r139_c163 bl[163] br[163] wl[139] vdd gnd cell_6t
Xbit_r140_c163 bl[163] br[163] wl[140] vdd gnd cell_6t
Xbit_r141_c163 bl[163] br[163] wl[141] vdd gnd cell_6t
Xbit_r142_c163 bl[163] br[163] wl[142] vdd gnd cell_6t
Xbit_r143_c163 bl[163] br[163] wl[143] vdd gnd cell_6t
Xbit_r144_c163 bl[163] br[163] wl[144] vdd gnd cell_6t
Xbit_r145_c163 bl[163] br[163] wl[145] vdd gnd cell_6t
Xbit_r146_c163 bl[163] br[163] wl[146] vdd gnd cell_6t
Xbit_r147_c163 bl[163] br[163] wl[147] vdd gnd cell_6t
Xbit_r148_c163 bl[163] br[163] wl[148] vdd gnd cell_6t
Xbit_r149_c163 bl[163] br[163] wl[149] vdd gnd cell_6t
Xbit_r150_c163 bl[163] br[163] wl[150] vdd gnd cell_6t
Xbit_r151_c163 bl[163] br[163] wl[151] vdd gnd cell_6t
Xbit_r152_c163 bl[163] br[163] wl[152] vdd gnd cell_6t
Xbit_r153_c163 bl[163] br[163] wl[153] vdd gnd cell_6t
Xbit_r154_c163 bl[163] br[163] wl[154] vdd gnd cell_6t
Xbit_r155_c163 bl[163] br[163] wl[155] vdd gnd cell_6t
Xbit_r156_c163 bl[163] br[163] wl[156] vdd gnd cell_6t
Xbit_r157_c163 bl[163] br[163] wl[157] vdd gnd cell_6t
Xbit_r158_c163 bl[163] br[163] wl[158] vdd gnd cell_6t
Xbit_r159_c163 bl[163] br[163] wl[159] vdd gnd cell_6t
Xbit_r160_c163 bl[163] br[163] wl[160] vdd gnd cell_6t
Xbit_r161_c163 bl[163] br[163] wl[161] vdd gnd cell_6t
Xbit_r162_c163 bl[163] br[163] wl[162] vdd gnd cell_6t
Xbit_r163_c163 bl[163] br[163] wl[163] vdd gnd cell_6t
Xbit_r164_c163 bl[163] br[163] wl[164] vdd gnd cell_6t
Xbit_r165_c163 bl[163] br[163] wl[165] vdd gnd cell_6t
Xbit_r166_c163 bl[163] br[163] wl[166] vdd gnd cell_6t
Xbit_r167_c163 bl[163] br[163] wl[167] vdd gnd cell_6t
Xbit_r168_c163 bl[163] br[163] wl[168] vdd gnd cell_6t
Xbit_r169_c163 bl[163] br[163] wl[169] vdd gnd cell_6t
Xbit_r170_c163 bl[163] br[163] wl[170] vdd gnd cell_6t
Xbit_r171_c163 bl[163] br[163] wl[171] vdd gnd cell_6t
Xbit_r172_c163 bl[163] br[163] wl[172] vdd gnd cell_6t
Xbit_r173_c163 bl[163] br[163] wl[173] vdd gnd cell_6t
Xbit_r174_c163 bl[163] br[163] wl[174] vdd gnd cell_6t
Xbit_r175_c163 bl[163] br[163] wl[175] vdd gnd cell_6t
Xbit_r176_c163 bl[163] br[163] wl[176] vdd gnd cell_6t
Xbit_r177_c163 bl[163] br[163] wl[177] vdd gnd cell_6t
Xbit_r178_c163 bl[163] br[163] wl[178] vdd gnd cell_6t
Xbit_r179_c163 bl[163] br[163] wl[179] vdd gnd cell_6t
Xbit_r180_c163 bl[163] br[163] wl[180] vdd gnd cell_6t
Xbit_r181_c163 bl[163] br[163] wl[181] vdd gnd cell_6t
Xbit_r182_c163 bl[163] br[163] wl[182] vdd gnd cell_6t
Xbit_r183_c163 bl[163] br[163] wl[183] vdd gnd cell_6t
Xbit_r184_c163 bl[163] br[163] wl[184] vdd gnd cell_6t
Xbit_r185_c163 bl[163] br[163] wl[185] vdd gnd cell_6t
Xbit_r186_c163 bl[163] br[163] wl[186] vdd gnd cell_6t
Xbit_r187_c163 bl[163] br[163] wl[187] vdd gnd cell_6t
Xbit_r188_c163 bl[163] br[163] wl[188] vdd gnd cell_6t
Xbit_r189_c163 bl[163] br[163] wl[189] vdd gnd cell_6t
Xbit_r190_c163 bl[163] br[163] wl[190] vdd gnd cell_6t
Xbit_r191_c163 bl[163] br[163] wl[191] vdd gnd cell_6t
Xbit_r192_c163 bl[163] br[163] wl[192] vdd gnd cell_6t
Xbit_r193_c163 bl[163] br[163] wl[193] vdd gnd cell_6t
Xbit_r194_c163 bl[163] br[163] wl[194] vdd gnd cell_6t
Xbit_r195_c163 bl[163] br[163] wl[195] vdd gnd cell_6t
Xbit_r196_c163 bl[163] br[163] wl[196] vdd gnd cell_6t
Xbit_r197_c163 bl[163] br[163] wl[197] vdd gnd cell_6t
Xbit_r198_c163 bl[163] br[163] wl[198] vdd gnd cell_6t
Xbit_r199_c163 bl[163] br[163] wl[199] vdd gnd cell_6t
Xbit_r200_c163 bl[163] br[163] wl[200] vdd gnd cell_6t
Xbit_r201_c163 bl[163] br[163] wl[201] vdd gnd cell_6t
Xbit_r202_c163 bl[163] br[163] wl[202] vdd gnd cell_6t
Xbit_r203_c163 bl[163] br[163] wl[203] vdd gnd cell_6t
Xbit_r204_c163 bl[163] br[163] wl[204] vdd gnd cell_6t
Xbit_r205_c163 bl[163] br[163] wl[205] vdd gnd cell_6t
Xbit_r206_c163 bl[163] br[163] wl[206] vdd gnd cell_6t
Xbit_r207_c163 bl[163] br[163] wl[207] vdd gnd cell_6t
Xbit_r208_c163 bl[163] br[163] wl[208] vdd gnd cell_6t
Xbit_r209_c163 bl[163] br[163] wl[209] vdd gnd cell_6t
Xbit_r210_c163 bl[163] br[163] wl[210] vdd gnd cell_6t
Xbit_r211_c163 bl[163] br[163] wl[211] vdd gnd cell_6t
Xbit_r212_c163 bl[163] br[163] wl[212] vdd gnd cell_6t
Xbit_r213_c163 bl[163] br[163] wl[213] vdd gnd cell_6t
Xbit_r214_c163 bl[163] br[163] wl[214] vdd gnd cell_6t
Xbit_r215_c163 bl[163] br[163] wl[215] vdd gnd cell_6t
Xbit_r216_c163 bl[163] br[163] wl[216] vdd gnd cell_6t
Xbit_r217_c163 bl[163] br[163] wl[217] vdd gnd cell_6t
Xbit_r218_c163 bl[163] br[163] wl[218] vdd gnd cell_6t
Xbit_r219_c163 bl[163] br[163] wl[219] vdd gnd cell_6t
Xbit_r220_c163 bl[163] br[163] wl[220] vdd gnd cell_6t
Xbit_r221_c163 bl[163] br[163] wl[221] vdd gnd cell_6t
Xbit_r222_c163 bl[163] br[163] wl[222] vdd gnd cell_6t
Xbit_r223_c163 bl[163] br[163] wl[223] vdd gnd cell_6t
Xbit_r224_c163 bl[163] br[163] wl[224] vdd gnd cell_6t
Xbit_r225_c163 bl[163] br[163] wl[225] vdd gnd cell_6t
Xbit_r226_c163 bl[163] br[163] wl[226] vdd gnd cell_6t
Xbit_r227_c163 bl[163] br[163] wl[227] vdd gnd cell_6t
Xbit_r228_c163 bl[163] br[163] wl[228] vdd gnd cell_6t
Xbit_r229_c163 bl[163] br[163] wl[229] vdd gnd cell_6t
Xbit_r230_c163 bl[163] br[163] wl[230] vdd gnd cell_6t
Xbit_r231_c163 bl[163] br[163] wl[231] vdd gnd cell_6t
Xbit_r232_c163 bl[163] br[163] wl[232] vdd gnd cell_6t
Xbit_r233_c163 bl[163] br[163] wl[233] vdd gnd cell_6t
Xbit_r234_c163 bl[163] br[163] wl[234] vdd gnd cell_6t
Xbit_r235_c163 bl[163] br[163] wl[235] vdd gnd cell_6t
Xbit_r236_c163 bl[163] br[163] wl[236] vdd gnd cell_6t
Xbit_r237_c163 bl[163] br[163] wl[237] vdd gnd cell_6t
Xbit_r238_c163 bl[163] br[163] wl[238] vdd gnd cell_6t
Xbit_r239_c163 bl[163] br[163] wl[239] vdd gnd cell_6t
Xbit_r240_c163 bl[163] br[163] wl[240] vdd gnd cell_6t
Xbit_r241_c163 bl[163] br[163] wl[241] vdd gnd cell_6t
Xbit_r242_c163 bl[163] br[163] wl[242] vdd gnd cell_6t
Xbit_r243_c163 bl[163] br[163] wl[243] vdd gnd cell_6t
Xbit_r244_c163 bl[163] br[163] wl[244] vdd gnd cell_6t
Xbit_r245_c163 bl[163] br[163] wl[245] vdd gnd cell_6t
Xbit_r246_c163 bl[163] br[163] wl[246] vdd gnd cell_6t
Xbit_r247_c163 bl[163] br[163] wl[247] vdd gnd cell_6t
Xbit_r248_c163 bl[163] br[163] wl[248] vdd gnd cell_6t
Xbit_r249_c163 bl[163] br[163] wl[249] vdd gnd cell_6t
Xbit_r250_c163 bl[163] br[163] wl[250] vdd gnd cell_6t
Xbit_r251_c163 bl[163] br[163] wl[251] vdd gnd cell_6t
Xbit_r252_c163 bl[163] br[163] wl[252] vdd gnd cell_6t
Xbit_r253_c163 bl[163] br[163] wl[253] vdd gnd cell_6t
Xbit_r254_c163 bl[163] br[163] wl[254] vdd gnd cell_6t
Xbit_r255_c163 bl[163] br[163] wl[255] vdd gnd cell_6t
Xbit_r0_c164 bl[164] br[164] wl[0] vdd gnd cell_6t
Xbit_r1_c164 bl[164] br[164] wl[1] vdd gnd cell_6t
Xbit_r2_c164 bl[164] br[164] wl[2] vdd gnd cell_6t
Xbit_r3_c164 bl[164] br[164] wl[3] vdd gnd cell_6t
Xbit_r4_c164 bl[164] br[164] wl[4] vdd gnd cell_6t
Xbit_r5_c164 bl[164] br[164] wl[5] vdd gnd cell_6t
Xbit_r6_c164 bl[164] br[164] wl[6] vdd gnd cell_6t
Xbit_r7_c164 bl[164] br[164] wl[7] vdd gnd cell_6t
Xbit_r8_c164 bl[164] br[164] wl[8] vdd gnd cell_6t
Xbit_r9_c164 bl[164] br[164] wl[9] vdd gnd cell_6t
Xbit_r10_c164 bl[164] br[164] wl[10] vdd gnd cell_6t
Xbit_r11_c164 bl[164] br[164] wl[11] vdd gnd cell_6t
Xbit_r12_c164 bl[164] br[164] wl[12] vdd gnd cell_6t
Xbit_r13_c164 bl[164] br[164] wl[13] vdd gnd cell_6t
Xbit_r14_c164 bl[164] br[164] wl[14] vdd gnd cell_6t
Xbit_r15_c164 bl[164] br[164] wl[15] vdd gnd cell_6t
Xbit_r16_c164 bl[164] br[164] wl[16] vdd gnd cell_6t
Xbit_r17_c164 bl[164] br[164] wl[17] vdd gnd cell_6t
Xbit_r18_c164 bl[164] br[164] wl[18] vdd gnd cell_6t
Xbit_r19_c164 bl[164] br[164] wl[19] vdd gnd cell_6t
Xbit_r20_c164 bl[164] br[164] wl[20] vdd gnd cell_6t
Xbit_r21_c164 bl[164] br[164] wl[21] vdd gnd cell_6t
Xbit_r22_c164 bl[164] br[164] wl[22] vdd gnd cell_6t
Xbit_r23_c164 bl[164] br[164] wl[23] vdd gnd cell_6t
Xbit_r24_c164 bl[164] br[164] wl[24] vdd gnd cell_6t
Xbit_r25_c164 bl[164] br[164] wl[25] vdd gnd cell_6t
Xbit_r26_c164 bl[164] br[164] wl[26] vdd gnd cell_6t
Xbit_r27_c164 bl[164] br[164] wl[27] vdd gnd cell_6t
Xbit_r28_c164 bl[164] br[164] wl[28] vdd gnd cell_6t
Xbit_r29_c164 bl[164] br[164] wl[29] vdd gnd cell_6t
Xbit_r30_c164 bl[164] br[164] wl[30] vdd gnd cell_6t
Xbit_r31_c164 bl[164] br[164] wl[31] vdd gnd cell_6t
Xbit_r32_c164 bl[164] br[164] wl[32] vdd gnd cell_6t
Xbit_r33_c164 bl[164] br[164] wl[33] vdd gnd cell_6t
Xbit_r34_c164 bl[164] br[164] wl[34] vdd gnd cell_6t
Xbit_r35_c164 bl[164] br[164] wl[35] vdd gnd cell_6t
Xbit_r36_c164 bl[164] br[164] wl[36] vdd gnd cell_6t
Xbit_r37_c164 bl[164] br[164] wl[37] vdd gnd cell_6t
Xbit_r38_c164 bl[164] br[164] wl[38] vdd gnd cell_6t
Xbit_r39_c164 bl[164] br[164] wl[39] vdd gnd cell_6t
Xbit_r40_c164 bl[164] br[164] wl[40] vdd gnd cell_6t
Xbit_r41_c164 bl[164] br[164] wl[41] vdd gnd cell_6t
Xbit_r42_c164 bl[164] br[164] wl[42] vdd gnd cell_6t
Xbit_r43_c164 bl[164] br[164] wl[43] vdd gnd cell_6t
Xbit_r44_c164 bl[164] br[164] wl[44] vdd gnd cell_6t
Xbit_r45_c164 bl[164] br[164] wl[45] vdd gnd cell_6t
Xbit_r46_c164 bl[164] br[164] wl[46] vdd gnd cell_6t
Xbit_r47_c164 bl[164] br[164] wl[47] vdd gnd cell_6t
Xbit_r48_c164 bl[164] br[164] wl[48] vdd gnd cell_6t
Xbit_r49_c164 bl[164] br[164] wl[49] vdd gnd cell_6t
Xbit_r50_c164 bl[164] br[164] wl[50] vdd gnd cell_6t
Xbit_r51_c164 bl[164] br[164] wl[51] vdd gnd cell_6t
Xbit_r52_c164 bl[164] br[164] wl[52] vdd gnd cell_6t
Xbit_r53_c164 bl[164] br[164] wl[53] vdd gnd cell_6t
Xbit_r54_c164 bl[164] br[164] wl[54] vdd gnd cell_6t
Xbit_r55_c164 bl[164] br[164] wl[55] vdd gnd cell_6t
Xbit_r56_c164 bl[164] br[164] wl[56] vdd gnd cell_6t
Xbit_r57_c164 bl[164] br[164] wl[57] vdd gnd cell_6t
Xbit_r58_c164 bl[164] br[164] wl[58] vdd gnd cell_6t
Xbit_r59_c164 bl[164] br[164] wl[59] vdd gnd cell_6t
Xbit_r60_c164 bl[164] br[164] wl[60] vdd gnd cell_6t
Xbit_r61_c164 bl[164] br[164] wl[61] vdd gnd cell_6t
Xbit_r62_c164 bl[164] br[164] wl[62] vdd gnd cell_6t
Xbit_r63_c164 bl[164] br[164] wl[63] vdd gnd cell_6t
Xbit_r64_c164 bl[164] br[164] wl[64] vdd gnd cell_6t
Xbit_r65_c164 bl[164] br[164] wl[65] vdd gnd cell_6t
Xbit_r66_c164 bl[164] br[164] wl[66] vdd gnd cell_6t
Xbit_r67_c164 bl[164] br[164] wl[67] vdd gnd cell_6t
Xbit_r68_c164 bl[164] br[164] wl[68] vdd gnd cell_6t
Xbit_r69_c164 bl[164] br[164] wl[69] vdd gnd cell_6t
Xbit_r70_c164 bl[164] br[164] wl[70] vdd gnd cell_6t
Xbit_r71_c164 bl[164] br[164] wl[71] vdd gnd cell_6t
Xbit_r72_c164 bl[164] br[164] wl[72] vdd gnd cell_6t
Xbit_r73_c164 bl[164] br[164] wl[73] vdd gnd cell_6t
Xbit_r74_c164 bl[164] br[164] wl[74] vdd gnd cell_6t
Xbit_r75_c164 bl[164] br[164] wl[75] vdd gnd cell_6t
Xbit_r76_c164 bl[164] br[164] wl[76] vdd gnd cell_6t
Xbit_r77_c164 bl[164] br[164] wl[77] vdd gnd cell_6t
Xbit_r78_c164 bl[164] br[164] wl[78] vdd gnd cell_6t
Xbit_r79_c164 bl[164] br[164] wl[79] vdd gnd cell_6t
Xbit_r80_c164 bl[164] br[164] wl[80] vdd gnd cell_6t
Xbit_r81_c164 bl[164] br[164] wl[81] vdd gnd cell_6t
Xbit_r82_c164 bl[164] br[164] wl[82] vdd gnd cell_6t
Xbit_r83_c164 bl[164] br[164] wl[83] vdd gnd cell_6t
Xbit_r84_c164 bl[164] br[164] wl[84] vdd gnd cell_6t
Xbit_r85_c164 bl[164] br[164] wl[85] vdd gnd cell_6t
Xbit_r86_c164 bl[164] br[164] wl[86] vdd gnd cell_6t
Xbit_r87_c164 bl[164] br[164] wl[87] vdd gnd cell_6t
Xbit_r88_c164 bl[164] br[164] wl[88] vdd gnd cell_6t
Xbit_r89_c164 bl[164] br[164] wl[89] vdd gnd cell_6t
Xbit_r90_c164 bl[164] br[164] wl[90] vdd gnd cell_6t
Xbit_r91_c164 bl[164] br[164] wl[91] vdd gnd cell_6t
Xbit_r92_c164 bl[164] br[164] wl[92] vdd gnd cell_6t
Xbit_r93_c164 bl[164] br[164] wl[93] vdd gnd cell_6t
Xbit_r94_c164 bl[164] br[164] wl[94] vdd gnd cell_6t
Xbit_r95_c164 bl[164] br[164] wl[95] vdd gnd cell_6t
Xbit_r96_c164 bl[164] br[164] wl[96] vdd gnd cell_6t
Xbit_r97_c164 bl[164] br[164] wl[97] vdd gnd cell_6t
Xbit_r98_c164 bl[164] br[164] wl[98] vdd gnd cell_6t
Xbit_r99_c164 bl[164] br[164] wl[99] vdd gnd cell_6t
Xbit_r100_c164 bl[164] br[164] wl[100] vdd gnd cell_6t
Xbit_r101_c164 bl[164] br[164] wl[101] vdd gnd cell_6t
Xbit_r102_c164 bl[164] br[164] wl[102] vdd gnd cell_6t
Xbit_r103_c164 bl[164] br[164] wl[103] vdd gnd cell_6t
Xbit_r104_c164 bl[164] br[164] wl[104] vdd gnd cell_6t
Xbit_r105_c164 bl[164] br[164] wl[105] vdd gnd cell_6t
Xbit_r106_c164 bl[164] br[164] wl[106] vdd gnd cell_6t
Xbit_r107_c164 bl[164] br[164] wl[107] vdd gnd cell_6t
Xbit_r108_c164 bl[164] br[164] wl[108] vdd gnd cell_6t
Xbit_r109_c164 bl[164] br[164] wl[109] vdd gnd cell_6t
Xbit_r110_c164 bl[164] br[164] wl[110] vdd gnd cell_6t
Xbit_r111_c164 bl[164] br[164] wl[111] vdd gnd cell_6t
Xbit_r112_c164 bl[164] br[164] wl[112] vdd gnd cell_6t
Xbit_r113_c164 bl[164] br[164] wl[113] vdd gnd cell_6t
Xbit_r114_c164 bl[164] br[164] wl[114] vdd gnd cell_6t
Xbit_r115_c164 bl[164] br[164] wl[115] vdd gnd cell_6t
Xbit_r116_c164 bl[164] br[164] wl[116] vdd gnd cell_6t
Xbit_r117_c164 bl[164] br[164] wl[117] vdd gnd cell_6t
Xbit_r118_c164 bl[164] br[164] wl[118] vdd gnd cell_6t
Xbit_r119_c164 bl[164] br[164] wl[119] vdd gnd cell_6t
Xbit_r120_c164 bl[164] br[164] wl[120] vdd gnd cell_6t
Xbit_r121_c164 bl[164] br[164] wl[121] vdd gnd cell_6t
Xbit_r122_c164 bl[164] br[164] wl[122] vdd gnd cell_6t
Xbit_r123_c164 bl[164] br[164] wl[123] vdd gnd cell_6t
Xbit_r124_c164 bl[164] br[164] wl[124] vdd gnd cell_6t
Xbit_r125_c164 bl[164] br[164] wl[125] vdd gnd cell_6t
Xbit_r126_c164 bl[164] br[164] wl[126] vdd gnd cell_6t
Xbit_r127_c164 bl[164] br[164] wl[127] vdd gnd cell_6t
Xbit_r128_c164 bl[164] br[164] wl[128] vdd gnd cell_6t
Xbit_r129_c164 bl[164] br[164] wl[129] vdd gnd cell_6t
Xbit_r130_c164 bl[164] br[164] wl[130] vdd gnd cell_6t
Xbit_r131_c164 bl[164] br[164] wl[131] vdd gnd cell_6t
Xbit_r132_c164 bl[164] br[164] wl[132] vdd gnd cell_6t
Xbit_r133_c164 bl[164] br[164] wl[133] vdd gnd cell_6t
Xbit_r134_c164 bl[164] br[164] wl[134] vdd gnd cell_6t
Xbit_r135_c164 bl[164] br[164] wl[135] vdd gnd cell_6t
Xbit_r136_c164 bl[164] br[164] wl[136] vdd gnd cell_6t
Xbit_r137_c164 bl[164] br[164] wl[137] vdd gnd cell_6t
Xbit_r138_c164 bl[164] br[164] wl[138] vdd gnd cell_6t
Xbit_r139_c164 bl[164] br[164] wl[139] vdd gnd cell_6t
Xbit_r140_c164 bl[164] br[164] wl[140] vdd gnd cell_6t
Xbit_r141_c164 bl[164] br[164] wl[141] vdd gnd cell_6t
Xbit_r142_c164 bl[164] br[164] wl[142] vdd gnd cell_6t
Xbit_r143_c164 bl[164] br[164] wl[143] vdd gnd cell_6t
Xbit_r144_c164 bl[164] br[164] wl[144] vdd gnd cell_6t
Xbit_r145_c164 bl[164] br[164] wl[145] vdd gnd cell_6t
Xbit_r146_c164 bl[164] br[164] wl[146] vdd gnd cell_6t
Xbit_r147_c164 bl[164] br[164] wl[147] vdd gnd cell_6t
Xbit_r148_c164 bl[164] br[164] wl[148] vdd gnd cell_6t
Xbit_r149_c164 bl[164] br[164] wl[149] vdd gnd cell_6t
Xbit_r150_c164 bl[164] br[164] wl[150] vdd gnd cell_6t
Xbit_r151_c164 bl[164] br[164] wl[151] vdd gnd cell_6t
Xbit_r152_c164 bl[164] br[164] wl[152] vdd gnd cell_6t
Xbit_r153_c164 bl[164] br[164] wl[153] vdd gnd cell_6t
Xbit_r154_c164 bl[164] br[164] wl[154] vdd gnd cell_6t
Xbit_r155_c164 bl[164] br[164] wl[155] vdd gnd cell_6t
Xbit_r156_c164 bl[164] br[164] wl[156] vdd gnd cell_6t
Xbit_r157_c164 bl[164] br[164] wl[157] vdd gnd cell_6t
Xbit_r158_c164 bl[164] br[164] wl[158] vdd gnd cell_6t
Xbit_r159_c164 bl[164] br[164] wl[159] vdd gnd cell_6t
Xbit_r160_c164 bl[164] br[164] wl[160] vdd gnd cell_6t
Xbit_r161_c164 bl[164] br[164] wl[161] vdd gnd cell_6t
Xbit_r162_c164 bl[164] br[164] wl[162] vdd gnd cell_6t
Xbit_r163_c164 bl[164] br[164] wl[163] vdd gnd cell_6t
Xbit_r164_c164 bl[164] br[164] wl[164] vdd gnd cell_6t
Xbit_r165_c164 bl[164] br[164] wl[165] vdd gnd cell_6t
Xbit_r166_c164 bl[164] br[164] wl[166] vdd gnd cell_6t
Xbit_r167_c164 bl[164] br[164] wl[167] vdd gnd cell_6t
Xbit_r168_c164 bl[164] br[164] wl[168] vdd gnd cell_6t
Xbit_r169_c164 bl[164] br[164] wl[169] vdd gnd cell_6t
Xbit_r170_c164 bl[164] br[164] wl[170] vdd gnd cell_6t
Xbit_r171_c164 bl[164] br[164] wl[171] vdd gnd cell_6t
Xbit_r172_c164 bl[164] br[164] wl[172] vdd gnd cell_6t
Xbit_r173_c164 bl[164] br[164] wl[173] vdd gnd cell_6t
Xbit_r174_c164 bl[164] br[164] wl[174] vdd gnd cell_6t
Xbit_r175_c164 bl[164] br[164] wl[175] vdd gnd cell_6t
Xbit_r176_c164 bl[164] br[164] wl[176] vdd gnd cell_6t
Xbit_r177_c164 bl[164] br[164] wl[177] vdd gnd cell_6t
Xbit_r178_c164 bl[164] br[164] wl[178] vdd gnd cell_6t
Xbit_r179_c164 bl[164] br[164] wl[179] vdd gnd cell_6t
Xbit_r180_c164 bl[164] br[164] wl[180] vdd gnd cell_6t
Xbit_r181_c164 bl[164] br[164] wl[181] vdd gnd cell_6t
Xbit_r182_c164 bl[164] br[164] wl[182] vdd gnd cell_6t
Xbit_r183_c164 bl[164] br[164] wl[183] vdd gnd cell_6t
Xbit_r184_c164 bl[164] br[164] wl[184] vdd gnd cell_6t
Xbit_r185_c164 bl[164] br[164] wl[185] vdd gnd cell_6t
Xbit_r186_c164 bl[164] br[164] wl[186] vdd gnd cell_6t
Xbit_r187_c164 bl[164] br[164] wl[187] vdd gnd cell_6t
Xbit_r188_c164 bl[164] br[164] wl[188] vdd gnd cell_6t
Xbit_r189_c164 bl[164] br[164] wl[189] vdd gnd cell_6t
Xbit_r190_c164 bl[164] br[164] wl[190] vdd gnd cell_6t
Xbit_r191_c164 bl[164] br[164] wl[191] vdd gnd cell_6t
Xbit_r192_c164 bl[164] br[164] wl[192] vdd gnd cell_6t
Xbit_r193_c164 bl[164] br[164] wl[193] vdd gnd cell_6t
Xbit_r194_c164 bl[164] br[164] wl[194] vdd gnd cell_6t
Xbit_r195_c164 bl[164] br[164] wl[195] vdd gnd cell_6t
Xbit_r196_c164 bl[164] br[164] wl[196] vdd gnd cell_6t
Xbit_r197_c164 bl[164] br[164] wl[197] vdd gnd cell_6t
Xbit_r198_c164 bl[164] br[164] wl[198] vdd gnd cell_6t
Xbit_r199_c164 bl[164] br[164] wl[199] vdd gnd cell_6t
Xbit_r200_c164 bl[164] br[164] wl[200] vdd gnd cell_6t
Xbit_r201_c164 bl[164] br[164] wl[201] vdd gnd cell_6t
Xbit_r202_c164 bl[164] br[164] wl[202] vdd gnd cell_6t
Xbit_r203_c164 bl[164] br[164] wl[203] vdd gnd cell_6t
Xbit_r204_c164 bl[164] br[164] wl[204] vdd gnd cell_6t
Xbit_r205_c164 bl[164] br[164] wl[205] vdd gnd cell_6t
Xbit_r206_c164 bl[164] br[164] wl[206] vdd gnd cell_6t
Xbit_r207_c164 bl[164] br[164] wl[207] vdd gnd cell_6t
Xbit_r208_c164 bl[164] br[164] wl[208] vdd gnd cell_6t
Xbit_r209_c164 bl[164] br[164] wl[209] vdd gnd cell_6t
Xbit_r210_c164 bl[164] br[164] wl[210] vdd gnd cell_6t
Xbit_r211_c164 bl[164] br[164] wl[211] vdd gnd cell_6t
Xbit_r212_c164 bl[164] br[164] wl[212] vdd gnd cell_6t
Xbit_r213_c164 bl[164] br[164] wl[213] vdd gnd cell_6t
Xbit_r214_c164 bl[164] br[164] wl[214] vdd gnd cell_6t
Xbit_r215_c164 bl[164] br[164] wl[215] vdd gnd cell_6t
Xbit_r216_c164 bl[164] br[164] wl[216] vdd gnd cell_6t
Xbit_r217_c164 bl[164] br[164] wl[217] vdd gnd cell_6t
Xbit_r218_c164 bl[164] br[164] wl[218] vdd gnd cell_6t
Xbit_r219_c164 bl[164] br[164] wl[219] vdd gnd cell_6t
Xbit_r220_c164 bl[164] br[164] wl[220] vdd gnd cell_6t
Xbit_r221_c164 bl[164] br[164] wl[221] vdd gnd cell_6t
Xbit_r222_c164 bl[164] br[164] wl[222] vdd gnd cell_6t
Xbit_r223_c164 bl[164] br[164] wl[223] vdd gnd cell_6t
Xbit_r224_c164 bl[164] br[164] wl[224] vdd gnd cell_6t
Xbit_r225_c164 bl[164] br[164] wl[225] vdd gnd cell_6t
Xbit_r226_c164 bl[164] br[164] wl[226] vdd gnd cell_6t
Xbit_r227_c164 bl[164] br[164] wl[227] vdd gnd cell_6t
Xbit_r228_c164 bl[164] br[164] wl[228] vdd gnd cell_6t
Xbit_r229_c164 bl[164] br[164] wl[229] vdd gnd cell_6t
Xbit_r230_c164 bl[164] br[164] wl[230] vdd gnd cell_6t
Xbit_r231_c164 bl[164] br[164] wl[231] vdd gnd cell_6t
Xbit_r232_c164 bl[164] br[164] wl[232] vdd gnd cell_6t
Xbit_r233_c164 bl[164] br[164] wl[233] vdd gnd cell_6t
Xbit_r234_c164 bl[164] br[164] wl[234] vdd gnd cell_6t
Xbit_r235_c164 bl[164] br[164] wl[235] vdd gnd cell_6t
Xbit_r236_c164 bl[164] br[164] wl[236] vdd gnd cell_6t
Xbit_r237_c164 bl[164] br[164] wl[237] vdd gnd cell_6t
Xbit_r238_c164 bl[164] br[164] wl[238] vdd gnd cell_6t
Xbit_r239_c164 bl[164] br[164] wl[239] vdd gnd cell_6t
Xbit_r240_c164 bl[164] br[164] wl[240] vdd gnd cell_6t
Xbit_r241_c164 bl[164] br[164] wl[241] vdd gnd cell_6t
Xbit_r242_c164 bl[164] br[164] wl[242] vdd gnd cell_6t
Xbit_r243_c164 bl[164] br[164] wl[243] vdd gnd cell_6t
Xbit_r244_c164 bl[164] br[164] wl[244] vdd gnd cell_6t
Xbit_r245_c164 bl[164] br[164] wl[245] vdd gnd cell_6t
Xbit_r246_c164 bl[164] br[164] wl[246] vdd gnd cell_6t
Xbit_r247_c164 bl[164] br[164] wl[247] vdd gnd cell_6t
Xbit_r248_c164 bl[164] br[164] wl[248] vdd gnd cell_6t
Xbit_r249_c164 bl[164] br[164] wl[249] vdd gnd cell_6t
Xbit_r250_c164 bl[164] br[164] wl[250] vdd gnd cell_6t
Xbit_r251_c164 bl[164] br[164] wl[251] vdd gnd cell_6t
Xbit_r252_c164 bl[164] br[164] wl[252] vdd gnd cell_6t
Xbit_r253_c164 bl[164] br[164] wl[253] vdd gnd cell_6t
Xbit_r254_c164 bl[164] br[164] wl[254] vdd gnd cell_6t
Xbit_r255_c164 bl[164] br[164] wl[255] vdd gnd cell_6t
Xbit_r0_c165 bl[165] br[165] wl[0] vdd gnd cell_6t
Xbit_r1_c165 bl[165] br[165] wl[1] vdd gnd cell_6t
Xbit_r2_c165 bl[165] br[165] wl[2] vdd gnd cell_6t
Xbit_r3_c165 bl[165] br[165] wl[3] vdd gnd cell_6t
Xbit_r4_c165 bl[165] br[165] wl[4] vdd gnd cell_6t
Xbit_r5_c165 bl[165] br[165] wl[5] vdd gnd cell_6t
Xbit_r6_c165 bl[165] br[165] wl[6] vdd gnd cell_6t
Xbit_r7_c165 bl[165] br[165] wl[7] vdd gnd cell_6t
Xbit_r8_c165 bl[165] br[165] wl[8] vdd gnd cell_6t
Xbit_r9_c165 bl[165] br[165] wl[9] vdd gnd cell_6t
Xbit_r10_c165 bl[165] br[165] wl[10] vdd gnd cell_6t
Xbit_r11_c165 bl[165] br[165] wl[11] vdd gnd cell_6t
Xbit_r12_c165 bl[165] br[165] wl[12] vdd gnd cell_6t
Xbit_r13_c165 bl[165] br[165] wl[13] vdd gnd cell_6t
Xbit_r14_c165 bl[165] br[165] wl[14] vdd gnd cell_6t
Xbit_r15_c165 bl[165] br[165] wl[15] vdd gnd cell_6t
Xbit_r16_c165 bl[165] br[165] wl[16] vdd gnd cell_6t
Xbit_r17_c165 bl[165] br[165] wl[17] vdd gnd cell_6t
Xbit_r18_c165 bl[165] br[165] wl[18] vdd gnd cell_6t
Xbit_r19_c165 bl[165] br[165] wl[19] vdd gnd cell_6t
Xbit_r20_c165 bl[165] br[165] wl[20] vdd gnd cell_6t
Xbit_r21_c165 bl[165] br[165] wl[21] vdd gnd cell_6t
Xbit_r22_c165 bl[165] br[165] wl[22] vdd gnd cell_6t
Xbit_r23_c165 bl[165] br[165] wl[23] vdd gnd cell_6t
Xbit_r24_c165 bl[165] br[165] wl[24] vdd gnd cell_6t
Xbit_r25_c165 bl[165] br[165] wl[25] vdd gnd cell_6t
Xbit_r26_c165 bl[165] br[165] wl[26] vdd gnd cell_6t
Xbit_r27_c165 bl[165] br[165] wl[27] vdd gnd cell_6t
Xbit_r28_c165 bl[165] br[165] wl[28] vdd gnd cell_6t
Xbit_r29_c165 bl[165] br[165] wl[29] vdd gnd cell_6t
Xbit_r30_c165 bl[165] br[165] wl[30] vdd gnd cell_6t
Xbit_r31_c165 bl[165] br[165] wl[31] vdd gnd cell_6t
Xbit_r32_c165 bl[165] br[165] wl[32] vdd gnd cell_6t
Xbit_r33_c165 bl[165] br[165] wl[33] vdd gnd cell_6t
Xbit_r34_c165 bl[165] br[165] wl[34] vdd gnd cell_6t
Xbit_r35_c165 bl[165] br[165] wl[35] vdd gnd cell_6t
Xbit_r36_c165 bl[165] br[165] wl[36] vdd gnd cell_6t
Xbit_r37_c165 bl[165] br[165] wl[37] vdd gnd cell_6t
Xbit_r38_c165 bl[165] br[165] wl[38] vdd gnd cell_6t
Xbit_r39_c165 bl[165] br[165] wl[39] vdd gnd cell_6t
Xbit_r40_c165 bl[165] br[165] wl[40] vdd gnd cell_6t
Xbit_r41_c165 bl[165] br[165] wl[41] vdd gnd cell_6t
Xbit_r42_c165 bl[165] br[165] wl[42] vdd gnd cell_6t
Xbit_r43_c165 bl[165] br[165] wl[43] vdd gnd cell_6t
Xbit_r44_c165 bl[165] br[165] wl[44] vdd gnd cell_6t
Xbit_r45_c165 bl[165] br[165] wl[45] vdd gnd cell_6t
Xbit_r46_c165 bl[165] br[165] wl[46] vdd gnd cell_6t
Xbit_r47_c165 bl[165] br[165] wl[47] vdd gnd cell_6t
Xbit_r48_c165 bl[165] br[165] wl[48] vdd gnd cell_6t
Xbit_r49_c165 bl[165] br[165] wl[49] vdd gnd cell_6t
Xbit_r50_c165 bl[165] br[165] wl[50] vdd gnd cell_6t
Xbit_r51_c165 bl[165] br[165] wl[51] vdd gnd cell_6t
Xbit_r52_c165 bl[165] br[165] wl[52] vdd gnd cell_6t
Xbit_r53_c165 bl[165] br[165] wl[53] vdd gnd cell_6t
Xbit_r54_c165 bl[165] br[165] wl[54] vdd gnd cell_6t
Xbit_r55_c165 bl[165] br[165] wl[55] vdd gnd cell_6t
Xbit_r56_c165 bl[165] br[165] wl[56] vdd gnd cell_6t
Xbit_r57_c165 bl[165] br[165] wl[57] vdd gnd cell_6t
Xbit_r58_c165 bl[165] br[165] wl[58] vdd gnd cell_6t
Xbit_r59_c165 bl[165] br[165] wl[59] vdd gnd cell_6t
Xbit_r60_c165 bl[165] br[165] wl[60] vdd gnd cell_6t
Xbit_r61_c165 bl[165] br[165] wl[61] vdd gnd cell_6t
Xbit_r62_c165 bl[165] br[165] wl[62] vdd gnd cell_6t
Xbit_r63_c165 bl[165] br[165] wl[63] vdd gnd cell_6t
Xbit_r64_c165 bl[165] br[165] wl[64] vdd gnd cell_6t
Xbit_r65_c165 bl[165] br[165] wl[65] vdd gnd cell_6t
Xbit_r66_c165 bl[165] br[165] wl[66] vdd gnd cell_6t
Xbit_r67_c165 bl[165] br[165] wl[67] vdd gnd cell_6t
Xbit_r68_c165 bl[165] br[165] wl[68] vdd gnd cell_6t
Xbit_r69_c165 bl[165] br[165] wl[69] vdd gnd cell_6t
Xbit_r70_c165 bl[165] br[165] wl[70] vdd gnd cell_6t
Xbit_r71_c165 bl[165] br[165] wl[71] vdd gnd cell_6t
Xbit_r72_c165 bl[165] br[165] wl[72] vdd gnd cell_6t
Xbit_r73_c165 bl[165] br[165] wl[73] vdd gnd cell_6t
Xbit_r74_c165 bl[165] br[165] wl[74] vdd gnd cell_6t
Xbit_r75_c165 bl[165] br[165] wl[75] vdd gnd cell_6t
Xbit_r76_c165 bl[165] br[165] wl[76] vdd gnd cell_6t
Xbit_r77_c165 bl[165] br[165] wl[77] vdd gnd cell_6t
Xbit_r78_c165 bl[165] br[165] wl[78] vdd gnd cell_6t
Xbit_r79_c165 bl[165] br[165] wl[79] vdd gnd cell_6t
Xbit_r80_c165 bl[165] br[165] wl[80] vdd gnd cell_6t
Xbit_r81_c165 bl[165] br[165] wl[81] vdd gnd cell_6t
Xbit_r82_c165 bl[165] br[165] wl[82] vdd gnd cell_6t
Xbit_r83_c165 bl[165] br[165] wl[83] vdd gnd cell_6t
Xbit_r84_c165 bl[165] br[165] wl[84] vdd gnd cell_6t
Xbit_r85_c165 bl[165] br[165] wl[85] vdd gnd cell_6t
Xbit_r86_c165 bl[165] br[165] wl[86] vdd gnd cell_6t
Xbit_r87_c165 bl[165] br[165] wl[87] vdd gnd cell_6t
Xbit_r88_c165 bl[165] br[165] wl[88] vdd gnd cell_6t
Xbit_r89_c165 bl[165] br[165] wl[89] vdd gnd cell_6t
Xbit_r90_c165 bl[165] br[165] wl[90] vdd gnd cell_6t
Xbit_r91_c165 bl[165] br[165] wl[91] vdd gnd cell_6t
Xbit_r92_c165 bl[165] br[165] wl[92] vdd gnd cell_6t
Xbit_r93_c165 bl[165] br[165] wl[93] vdd gnd cell_6t
Xbit_r94_c165 bl[165] br[165] wl[94] vdd gnd cell_6t
Xbit_r95_c165 bl[165] br[165] wl[95] vdd gnd cell_6t
Xbit_r96_c165 bl[165] br[165] wl[96] vdd gnd cell_6t
Xbit_r97_c165 bl[165] br[165] wl[97] vdd gnd cell_6t
Xbit_r98_c165 bl[165] br[165] wl[98] vdd gnd cell_6t
Xbit_r99_c165 bl[165] br[165] wl[99] vdd gnd cell_6t
Xbit_r100_c165 bl[165] br[165] wl[100] vdd gnd cell_6t
Xbit_r101_c165 bl[165] br[165] wl[101] vdd gnd cell_6t
Xbit_r102_c165 bl[165] br[165] wl[102] vdd gnd cell_6t
Xbit_r103_c165 bl[165] br[165] wl[103] vdd gnd cell_6t
Xbit_r104_c165 bl[165] br[165] wl[104] vdd gnd cell_6t
Xbit_r105_c165 bl[165] br[165] wl[105] vdd gnd cell_6t
Xbit_r106_c165 bl[165] br[165] wl[106] vdd gnd cell_6t
Xbit_r107_c165 bl[165] br[165] wl[107] vdd gnd cell_6t
Xbit_r108_c165 bl[165] br[165] wl[108] vdd gnd cell_6t
Xbit_r109_c165 bl[165] br[165] wl[109] vdd gnd cell_6t
Xbit_r110_c165 bl[165] br[165] wl[110] vdd gnd cell_6t
Xbit_r111_c165 bl[165] br[165] wl[111] vdd gnd cell_6t
Xbit_r112_c165 bl[165] br[165] wl[112] vdd gnd cell_6t
Xbit_r113_c165 bl[165] br[165] wl[113] vdd gnd cell_6t
Xbit_r114_c165 bl[165] br[165] wl[114] vdd gnd cell_6t
Xbit_r115_c165 bl[165] br[165] wl[115] vdd gnd cell_6t
Xbit_r116_c165 bl[165] br[165] wl[116] vdd gnd cell_6t
Xbit_r117_c165 bl[165] br[165] wl[117] vdd gnd cell_6t
Xbit_r118_c165 bl[165] br[165] wl[118] vdd gnd cell_6t
Xbit_r119_c165 bl[165] br[165] wl[119] vdd gnd cell_6t
Xbit_r120_c165 bl[165] br[165] wl[120] vdd gnd cell_6t
Xbit_r121_c165 bl[165] br[165] wl[121] vdd gnd cell_6t
Xbit_r122_c165 bl[165] br[165] wl[122] vdd gnd cell_6t
Xbit_r123_c165 bl[165] br[165] wl[123] vdd gnd cell_6t
Xbit_r124_c165 bl[165] br[165] wl[124] vdd gnd cell_6t
Xbit_r125_c165 bl[165] br[165] wl[125] vdd gnd cell_6t
Xbit_r126_c165 bl[165] br[165] wl[126] vdd gnd cell_6t
Xbit_r127_c165 bl[165] br[165] wl[127] vdd gnd cell_6t
Xbit_r128_c165 bl[165] br[165] wl[128] vdd gnd cell_6t
Xbit_r129_c165 bl[165] br[165] wl[129] vdd gnd cell_6t
Xbit_r130_c165 bl[165] br[165] wl[130] vdd gnd cell_6t
Xbit_r131_c165 bl[165] br[165] wl[131] vdd gnd cell_6t
Xbit_r132_c165 bl[165] br[165] wl[132] vdd gnd cell_6t
Xbit_r133_c165 bl[165] br[165] wl[133] vdd gnd cell_6t
Xbit_r134_c165 bl[165] br[165] wl[134] vdd gnd cell_6t
Xbit_r135_c165 bl[165] br[165] wl[135] vdd gnd cell_6t
Xbit_r136_c165 bl[165] br[165] wl[136] vdd gnd cell_6t
Xbit_r137_c165 bl[165] br[165] wl[137] vdd gnd cell_6t
Xbit_r138_c165 bl[165] br[165] wl[138] vdd gnd cell_6t
Xbit_r139_c165 bl[165] br[165] wl[139] vdd gnd cell_6t
Xbit_r140_c165 bl[165] br[165] wl[140] vdd gnd cell_6t
Xbit_r141_c165 bl[165] br[165] wl[141] vdd gnd cell_6t
Xbit_r142_c165 bl[165] br[165] wl[142] vdd gnd cell_6t
Xbit_r143_c165 bl[165] br[165] wl[143] vdd gnd cell_6t
Xbit_r144_c165 bl[165] br[165] wl[144] vdd gnd cell_6t
Xbit_r145_c165 bl[165] br[165] wl[145] vdd gnd cell_6t
Xbit_r146_c165 bl[165] br[165] wl[146] vdd gnd cell_6t
Xbit_r147_c165 bl[165] br[165] wl[147] vdd gnd cell_6t
Xbit_r148_c165 bl[165] br[165] wl[148] vdd gnd cell_6t
Xbit_r149_c165 bl[165] br[165] wl[149] vdd gnd cell_6t
Xbit_r150_c165 bl[165] br[165] wl[150] vdd gnd cell_6t
Xbit_r151_c165 bl[165] br[165] wl[151] vdd gnd cell_6t
Xbit_r152_c165 bl[165] br[165] wl[152] vdd gnd cell_6t
Xbit_r153_c165 bl[165] br[165] wl[153] vdd gnd cell_6t
Xbit_r154_c165 bl[165] br[165] wl[154] vdd gnd cell_6t
Xbit_r155_c165 bl[165] br[165] wl[155] vdd gnd cell_6t
Xbit_r156_c165 bl[165] br[165] wl[156] vdd gnd cell_6t
Xbit_r157_c165 bl[165] br[165] wl[157] vdd gnd cell_6t
Xbit_r158_c165 bl[165] br[165] wl[158] vdd gnd cell_6t
Xbit_r159_c165 bl[165] br[165] wl[159] vdd gnd cell_6t
Xbit_r160_c165 bl[165] br[165] wl[160] vdd gnd cell_6t
Xbit_r161_c165 bl[165] br[165] wl[161] vdd gnd cell_6t
Xbit_r162_c165 bl[165] br[165] wl[162] vdd gnd cell_6t
Xbit_r163_c165 bl[165] br[165] wl[163] vdd gnd cell_6t
Xbit_r164_c165 bl[165] br[165] wl[164] vdd gnd cell_6t
Xbit_r165_c165 bl[165] br[165] wl[165] vdd gnd cell_6t
Xbit_r166_c165 bl[165] br[165] wl[166] vdd gnd cell_6t
Xbit_r167_c165 bl[165] br[165] wl[167] vdd gnd cell_6t
Xbit_r168_c165 bl[165] br[165] wl[168] vdd gnd cell_6t
Xbit_r169_c165 bl[165] br[165] wl[169] vdd gnd cell_6t
Xbit_r170_c165 bl[165] br[165] wl[170] vdd gnd cell_6t
Xbit_r171_c165 bl[165] br[165] wl[171] vdd gnd cell_6t
Xbit_r172_c165 bl[165] br[165] wl[172] vdd gnd cell_6t
Xbit_r173_c165 bl[165] br[165] wl[173] vdd gnd cell_6t
Xbit_r174_c165 bl[165] br[165] wl[174] vdd gnd cell_6t
Xbit_r175_c165 bl[165] br[165] wl[175] vdd gnd cell_6t
Xbit_r176_c165 bl[165] br[165] wl[176] vdd gnd cell_6t
Xbit_r177_c165 bl[165] br[165] wl[177] vdd gnd cell_6t
Xbit_r178_c165 bl[165] br[165] wl[178] vdd gnd cell_6t
Xbit_r179_c165 bl[165] br[165] wl[179] vdd gnd cell_6t
Xbit_r180_c165 bl[165] br[165] wl[180] vdd gnd cell_6t
Xbit_r181_c165 bl[165] br[165] wl[181] vdd gnd cell_6t
Xbit_r182_c165 bl[165] br[165] wl[182] vdd gnd cell_6t
Xbit_r183_c165 bl[165] br[165] wl[183] vdd gnd cell_6t
Xbit_r184_c165 bl[165] br[165] wl[184] vdd gnd cell_6t
Xbit_r185_c165 bl[165] br[165] wl[185] vdd gnd cell_6t
Xbit_r186_c165 bl[165] br[165] wl[186] vdd gnd cell_6t
Xbit_r187_c165 bl[165] br[165] wl[187] vdd gnd cell_6t
Xbit_r188_c165 bl[165] br[165] wl[188] vdd gnd cell_6t
Xbit_r189_c165 bl[165] br[165] wl[189] vdd gnd cell_6t
Xbit_r190_c165 bl[165] br[165] wl[190] vdd gnd cell_6t
Xbit_r191_c165 bl[165] br[165] wl[191] vdd gnd cell_6t
Xbit_r192_c165 bl[165] br[165] wl[192] vdd gnd cell_6t
Xbit_r193_c165 bl[165] br[165] wl[193] vdd gnd cell_6t
Xbit_r194_c165 bl[165] br[165] wl[194] vdd gnd cell_6t
Xbit_r195_c165 bl[165] br[165] wl[195] vdd gnd cell_6t
Xbit_r196_c165 bl[165] br[165] wl[196] vdd gnd cell_6t
Xbit_r197_c165 bl[165] br[165] wl[197] vdd gnd cell_6t
Xbit_r198_c165 bl[165] br[165] wl[198] vdd gnd cell_6t
Xbit_r199_c165 bl[165] br[165] wl[199] vdd gnd cell_6t
Xbit_r200_c165 bl[165] br[165] wl[200] vdd gnd cell_6t
Xbit_r201_c165 bl[165] br[165] wl[201] vdd gnd cell_6t
Xbit_r202_c165 bl[165] br[165] wl[202] vdd gnd cell_6t
Xbit_r203_c165 bl[165] br[165] wl[203] vdd gnd cell_6t
Xbit_r204_c165 bl[165] br[165] wl[204] vdd gnd cell_6t
Xbit_r205_c165 bl[165] br[165] wl[205] vdd gnd cell_6t
Xbit_r206_c165 bl[165] br[165] wl[206] vdd gnd cell_6t
Xbit_r207_c165 bl[165] br[165] wl[207] vdd gnd cell_6t
Xbit_r208_c165 bl[165] br[165] wl[208] vdd gnd cell_6t
Xbit_r209_c165 bl[165] br[165] wl[209] vdd gnd cell_6t
Xbit_r210_c165 bl[165] br[165] wl[210] vdd gnd cell_6t
Xbit_r211_c165 bl[165] br[165] wl[211] vdd gnd cell_6t
Xbit_r212_c165 bl[165] br[165] wl[212] vdd gnd cell_6t
Xbit_r213_c165 bl[165] br[165] wl[213] vdd gnd cell_6t
Xbit_r214_c165 bl[165] br[165] wl[214] vdd gnd cell_6t
Xbit_r215_c165 bl[165] br[165] wl[215] vdd gnd cell_6t
Xbit_r216_c165 bl[165] br[165] wl[216] vdd gnd cell_6t
Xbit_r217_c165 bl[165] br[165] wl[217] vdd gnd cell_6t
Xbit_r218_c165 bl[165] br[165] wl[218] vdd gnd cell_6t
Xbit_r219_c165 bl[165] br[165] wl[219] vdd gnd cell_6t
Xbit_r220_c165 bl[165] br[165] wl[220] vdd gnd cell_6t
Xbit_r221_c165 bl[165] br[165] wl[221] vdd gnd cell_6t
Xbit_r222_c165 bl[165] br[165] wl[222] vdd gnd cell_6t
Xbit_r223_c165 bl[165] br[165] wl[223] vdd gnd cell_6t
Xbit_r224_c165 bl[165] br[165] wl[224] vdd gnd cell_6t
Xbit_r225_c165 bl[165] br[165] wl[225] vdd gnd cell_6t
Xbit_r226_c165 bl[165] br[165] wl[226] vdd gnd cell_6t
Xbit_r227_c165 bl[165] br[165] wl[227] vdd gnd cell_6t
Xbit_r228_c165 bl[165] br[165] wl[228] vdd gnd cell_6t
Xbit_r229_c165 bl[165] br[165] wl[229] vdd gnd cell_6t
Xbit_r230_c165 bl[165] br[165] wl[230] vdd gnd cell_6t
Xbit_r231_c165 bl[165] br[165] wl[231] vdd gnd cell_6t
Xbit_r232_c165 bl[165] br[165] wl[232] vdd gnd cell_6t
Xbit_r233_c165 bl[165] br[165] wl[233] vdd gnd cell_6t
Xbit_r234_c165 bl[165] br[165] wl[234] vdd gnd cell_6t
Xbit_r235_c165 bl[165] br[165] wl[235] vdd gnd cell_6t
Xbit_r236_c165 bl[165] br[165] wl[236] vdd gnd cell_6t
Xbit_r237_c165 bl[165] br[165] wl[237] vdd gnd cell_6t
Xbit_r238_c165 bl[165] br[165] wl[238] vdd gnd cell_6t
Xbit_r239_c165 bl[165] br[165] wl[239] vdd gnd cell_6t
Xbit_r240_c165 bl[165] br[165] wl[240] vdd gnd cell_6t
Xbit_r241_c165 bl[165] br[165] wl[241] vdd gnd cell_6t
Xbit_r242_c165 bl[165] br[165] wl[242] vdd gnd cell_6t
Xbit_r243_c165 bl[165] br[165] wl[243] vdd gnd cell_6t
Xbit_r244_c165 bl[165] br[165] wl[244] vdd gnd cell_6t
Xbit_r245_c165 bl[165] br[165] wl[245] vdd gnd cell_6t
Xbit_r246_c165 bl[165] br[165] wl[246] vdd gnd cell_6t
Xbit_r247_c165 bl[165] br[165] wl[247] vdd gnd cell_6t
Xbit_r248_c165 bl[165] br[165] wl[248] vdd gnd cell_6t
Xbit_r249_c165 bl[165] br[165] wl[249] vdd gnd cell_6t
Xbit_r250_c165 bl[165] br[165] wl[250] vdd gnd cell_6t
Xbit_r251_c165 bl[165] br[165] wl[251] vdd gnd cell_6t
Xbit_r252_c165 bl[165] br[165] wl[252] vdd gnd cell_6t
Xbit_r253_c165 bl[165] br[165] wl[253] vdd gnd cell_6t
Xbit_r254_c165 bl[165] br[165] wl[254] vdd gnd cell_6t
Xbit_r255_c165 bl[165] br[165] wl[255] vdd gnd cell_6t
Xbit_r0_c166 bl[166] br[166] wl[0] vdd gnd cell_6t
Xbit_r1_c166 bl[166] br[166] wl[1] vdd gnd cell_6t
Xbit_r2_c166 bl[166] br[166] wl[2] vdd gnd cell_6t
Xbit_r3_c166 bl[166] br[166] wl[3] vdd gnd cell_6t
Xbit_r4_c166 bl[166] br[166] wl[4] vdd gnd cell_6t
Xbit_r5_c166 bl[166] br[166] wl[5] vdd gnd cell_6t
Xbit_r6_c166 bl[166] br[166] wl[6] vdd gnd cell_6t
Xbit_r7_c166 bl[166] br[166] wl[7] vdd gnd cell_6t
Xbit_r8_c166 bl[166] br[166] wl[8] vdd gnd cell_6t
Xbit_r9_c166 bl[166] br[166] wl[9] vdd gnd cell_6t
Xbit_r10_c166 bl[166] br[166] wl[10] vdd gnd cell_6t
Xbit_r11_c166 bl[166] br[166] wl[11] vdd gnd cell_6t
Xbit_r12_c166 bl[166] br[166] wl[12] vdd gnd cell_6t
Xbit_r13_c166 bl[166] br[166] wl[13] vdd gnd cell_6t
Xbit_r14_c166 bl[166] br[166] wl[14] vdd gnd cell_6t
Xbit_r15_c166 bl[166] br[166] wl[15] vdd gnd cell_6t
Xbit_r16_c166 bl[166] br[166] wl[16] vdd gnd cell_6t
Xbit_r17_c166 bl[166] br[166] wl[17] vdd gnd cell_6t
Xbit_r18_c166 bl[166] br[166] wl[18] vdd gnd cell_6t
Xbit_r19_c166 bl[166] br[166] wl[19] vdd gnd cell_6t
Xbit_r20_c166 bl[166] br[166] wl[20] vdd gnd cell_6t
Xbit_r21_c166 bl[166] br[166] wl[21] vdd gnd cell_6t
Xbit_r22_c166 bl[166] br[166] wl[22] vdd gnd cell_6t
Xbit_r23_c166 bl[166] br[166] wl[23] vdd gnd cell_6t
Xbit_r24_c166 bl[166] br[166] wl[24] vdd gnd cell_6t
Xbit_r25_c166 bl[166] br[166] wl[25] vdd gnd cell_6t
Xbit_r26_c166 bl[166] br[166] wl[26] vdd gnd cell_6t
Xbit_r27_c166 bl[166] br[166] wl[27] vdd gnd cell_6t
Xbit_r28_c166 bl[166] br[166] wl[28] vdd gnd cell_6t
Xbit_r29_c166 bl[166] br[166] wl[29] vdd gnd cell_6t
Xbit_r30_c166 bl[166] br[166] wl[30] vdd gnd cell_6t
Xbit_r31_c166 bl[166] br[166] wl[31] vdd gnd cell_6t
Xbit_r32_c166 bl[166] br[166] wl[32] vdd gnd cell_6t
Xbit_r33_c166 bl[166] br[166] wl[33] vdd gnd cell_6t
Xbit_r34_c166 bl[166] br[166] wl[34] vdd gnd cell_6t
Xbit_r35_c166 bl[166] br[166] wl[35] vdd gnd cell_6t
Xbit_r36_c166 bl[166] br[166] wl[36] vdd gnd cell_6t
Xbit_r37_c166 bl[166] br[166] wl[37] vdd gnd cell_6t
Xbit_r38_c166 bl[166] br[166] wl[38] vdd gnd cell_6t
Xbit_r39_c166 bl[166] br[166] wl[39] vdd gnd cell_6t
Xbit_r40_c166 bl[166] br[166] wl[40] vdd gnd cell_6t
Xbit_r41_c166 bl[166] br[166] wl[41] vdd gnd cell_6t
Xbit_r42_c166 bl[166] br[166] wl[42] vdd gnd cell_6t
Xbit_r43_c166 bl[166] br[166] wl[43] vdd gnd cell_6t
Xbit_r44_c166 bl[166] br[166] wl[44] vdd gnd cell_6t
Xbit_r45_c166 bl[166] br[166] wl[45] vdd gnd cell_6t
Xbit_r46_c166 bl[166] br[166] wl[46] vdd gnd cell_6t
Xbit_r47_c166 bl[166] br[166] wl[47] vdd gnd cell_6t
Xbit_r48_c166 bl[166] br[166] wl[48] vdd gnd cell_6t
Xbit_r49_c166 bl[166] br[166] wl[49] vdd gnd cell_6t
Xbit_r50_c166 bl[166] br[166] wl[50] vdd gnd cell_6t
Xbit_r51_c166 bl[166] br[166] wl[51] vdd gnd cell_6t
Xbit_r52_c166 bl[166] br[166] wl[52] vdd gnd cell_6t
Xbit_r53_c166 bl[166] br[166] wl[53] vdd gnd cell_6t
Xbit_r54_c166 bl[166] br[166] wl[54] vdd gnd cell_6t
Xbit_r55_c166 bl[166] br[166] wl[55] vdd gnd cell_6t
Xbit_r56_c166 bl[166] br[166] wl[56] vdd gnd cell_6t
Xbit_r57_c166 bl[166] br[166] wl[57] vdd gnd cell_6t
Xbit_r58_c166 bl[166] br[166] wl[58] vdd gnd cell_6t
Xbit_r59_c166 bl[166] br[166] wl[59] vdd gnd cell_6t
Xbit_r60_c166 bl[166] br[166] wl[60] vdd gnd cell_6t
Xbit_r61_c166 bl[166] br[166] wl[61] vdd gnd cell_6t
Xbit_r62_c166 bl[166] br[166] wl[62] vdd gnd cell_6t
Xbit_r63_c166 bl[166] br[166] wl[63] vdd gnd cell_6t
Xbit_r64_c166 bl[166] br[166] wl[64] vdd gnd cell_6t
Xbit_r65_c166 bl[166] br[166] wl[65] vdd gnd cell_6t
Xbit_r66_c166 bl[166] br[166] wl[66] vdd gnd cell_6t
Xbit_r67_c166 bl[166] br[166] wl[67] vdd gnd cell_6t
Xbit_r68_c166 bl[166] br[166] wl[68] vdd gnd cell_6t
Xbit_r69_c166 bl[166] br[166] wl[69] vdd gnd cell_6t
Xbit_r70_c166 bl[166] br[166] wl[70] vdd gnd cell_6t
Xbit_r71_c166 bl[166] br[166] wl[71] vdd gnd cell_6t
Xbit_r72_c166 bl[166] br[166] wl[72] vdd gnd cell_6t
Xbit_r73_c166 bl[166] br[166] wl[73] vdd gnd cell_6t
Xbit_r74_c166 bl[166] br[166] wl[74] vdd gnd cell_6t
Xbit_r75_c166 bl[166] br[166] wl[75] vdd gnd cell_6t
Xbit_r76_c166 bl[166] br[166] wl[76] vdd gnd cell_6t
Xbit_r77_c166 bl[166] br[166] wl[77] vdd gnd cell_6t
Xbit_r78_c166 bl[166] br[166] wl[78] vdd gnd cell_6t
Xbit_r79_c166 bl[166] br[166] wl[79] vdd gnd cell_6t
Xbit_r80_c166 bl[166] br[166] wl[80] vdd gnd cell_6t
Xbit_r81_c166 bl[166] br[166] wl[81] vdd gnd cell_6t
Xbit_r82_c166 bl[166] br[166] wl[82] vdd gnd cell_6t
Xbit_r83_c166 bl[166] br[166] wl[83] vdd gnd cell_6t
Xbit_r84_c166 bl[166] br[166] wl[84] vdd gnd cell_6t
Xbit_r85_c166 bl[166] br[166] wl[85] vdd gnd cell_6t
Xbit_r86_c166 bl[166] br[166] wl[86] vdd gnd cell_6t
Xbit_r87_c166 bl[166] br[166] wl[87] vdd gnd cell_6t
Xbit_r88_c166 bl[166] br[166] wl[88] vdd gnd cell_6t
Xbit_r89_c166 bl[166] br[166] wl[89] vdd gnd cell_6t
Xbit_r90_c166 bl[166] br[166] wl[90] vdd gnd cell_6t
Xbit_r91_c166 bl[166] br[166] wl[91] vdd gnd cell_6t
Xbit_r92_c166 bl[166] br[166] wl[92] vdd gnd cell_6t
Xbit_r93_c166 bl[166] br[166] wl[93] vdd gnd cell_6t
Xbit_r94_c166 bl[166] br[166] wl[94] vdd gnd cell_6t
Xbit_r95_c166 bl[166] br[166] wl[95] vdd gnd cell_6t
Xbit_r96_c166 bl[166] br[166] wl[96] vdd gnd cell_6t
Xbit_r97_c166 bl[166] br[166] wl[97] vdd gnd cell_6t
Xbit_r98_c166 bl[166] br[166] wl[98] vdd gnd cell_6t
Xbit_r99_c166 bl[166] br[166] wl[99] vdd gnd cell_6t
Xbit_r100_c166 bl[166] br[166] wl[100] vdd gnd cell_6t
Xbit_r101_c166 bl[166] br[166] wl[101] vdd gnd cell_6t
Xbit_r102_c166 bl[166] br[166] wl[102] vdd gnd cell_6t
Xbit_r103_c166 bl[166] br[166] wl[103] vdd gnd cell_6t
Xbit_r104_c166 bl[166] br[166] wl[104] vdd gnd cell_6t
Xbit_r105_c166 bl[166] br[166] wl[105] vdd gnd cell_6t
Xbit_r106_c166 bl[166] br[166] wl[106] vdd gnd cell_6t
Xbit_r107_c166 bl[166] br[166] wl[107] vdd gnd cell_6t
Xbit_r108_c166 bl[166] br[166] wl[108] vdd gnd cell_6t
Xbit_r109_c166 bl[166] br[166] wl[109] vdd gnd cell_6t
Xbit_r110_c166 bl[166] br[166] wl[110] vdd gnd cell_6t
Xbit_r111_c166 bl[166] br[166] wl[111] vdd gnd cell_6t
Xbit_r112_c166 bl[166] br[166] wl[112] vdd gnd cell_6t
Xbit_r113_c166 bl[166] br[166] wl[113] vdd gnd cell_6t
Xbit_r114_c166 bl[166] br[166] wl[114] vdd gnd cell_6t
Xbit_r115_c166 bl[166] br[166] wl[115] vdd gnd cell_6t
Xbit_r116_c166 bl[166] br[166] wl[116] vdd gnd cell_6t
Xbit_r117_c166 bl[166] br[166] wl[117] vdd gnd cell_6t
Xbit_r118_c166 bl[166] br[166] wl[118] vdd gnd cell_6t
Xbit_r119_c166 bl[166] br[166] wl[119] vdd gnd cell_6t
Xbit_r120_c166 bl[166] br[166] wl[120] vdd gnd cell_6t
Xbit_r121_c166 bl[166] br[166] wl[121] vdd gnd cell_6t
Xbit_r122_c166 bl[166] br[166] wl[122] vdd gnd cell_6t
Xbit_r123_c166 bl[166] br[166] wl[123] vdd gnd cell_6t
Xbit_r124_c166 bl[166] br[166] wl[124] vdd gnd cell_6t
Xbit_r125_c166 bl[166] br[166] wl[125] vdd gnd cell_6t
Xbit_r126_c166 bl[166] br[166] wl[126] vdd gnd cell_6t
Xbit_r127_c166 bl[166] br[166] wl[127] vdd gnd cell_6t
Xbit_r128_c166 bl[166] br[166] wl[128] vdd gnd cell_6t
Xbit_r129_c166 bl[166] br[166] wl[129] vdd gnd cell_6t
Xbit_r130_c166 bl[166] br[166] wl[130] vdd gnd cell_6t
Xbit_r131_c166 bl[166] br[166] wl[131] vdd gnd cell_6t
Xbit_r132_c166 bl[166] br[166] wl[132] vdd gnd cell_6t
Xbit_r133_c166 bl[166] br[166] wl[133] vdd gnd cell_6t
Xbit_r134_c166 bl[166] br[166] wl[134] vdd gnd cell_6t
Xbit_r135_c166 bl[166] br[166] wl[135] vdd gnd cell_6t
Xbit_r136_c166 bl[166] br[166] wl[136] vdd gnd cell_6t
Xbit_r137_c166 bl[166] br[166] wl[137] vdd gnd cell_6t
Xbit_r138_c166 bl[166] br[166] wl[138] vdd gnd cell_6t
Xbit_r139_c166 bl[166] br[166] wl[139] vdd gnd cell_6t
Xbit_r140_c166 bl[166] br[166] wl[140] vdd gnd cell_6t
Xbit_r141_c166 bl[166] br[166] wl[141] vdd gnd cell_6t
Xbit_r142_c166 bl[166] br[166] wl[142] vdd gnd cell_6t
Xbit_r143_c166 bl[166] br[166] wl[143] vdd gnd cell_6t
Xbit_r144_c166 bl[166] br[166] wl[144] vdd gnd cell_6t
Xbit_r145_c166 bl[166] br[166] wl[145] vdd gnd cell_6t
Xbit_r146_c166 bl[166] br[166] wl[146] vdd gnd cell_6t
Xbit_r147_c166 bl[166] br[166] wl[147] vdd gnd cell_6t
Xbit_r148_c166 bl[166] br[166] wl[148] vdd gnd cell_6t
Xbit_r149_c166 bl[166] br[166] wl[149] vdd gnd cell_6t
Xbit_r150_c166 bl[166] br[166] wl[150] vdd gnd cell_6t
Xbit_r151_c166 bl[166] br[166] wl[151] vdd gnd cell_6t
Xbit_r152_c166 bl[166] br[166] wl[152] vdd gnd cell_6t
Xbit_r153_c166 bl[166] br[166] wl[153] vdd gnd cell_6t
Xbit_r154_c166 bl[166] br[166] wl[154] vdd gnd cell_6t
Xbit_r155_c166 bl[166] br[166] wl[155] vdd gnd cell_6t
Xbit_r156_c166 bl[166] br[166] wl[156] vdd gnd cell_6t
Xbit_r157_c166 bl[166] br[166] wl[157] vdd gnd cell_6t
Xbit_r158_c166 bl[166] br[166] wl[158] vdd gnd cell_6t
Xbit_r159_c166 bl[166] br[166] wl[159] vdd gnd cell_6t
Xbit_r160_c166 bl[166] br[166] wl[160] vdd gnd cell_6t
Xbit_r161_c166 bl[166] br[166] wl[161] vdd gnd cell_6t
Xbit_r162_c166 bl[166] br[166] wl[162] vdd gnd cell_6t
Xbit_r163_c166 bl[166] br[166] wl[163] vdd gnd cell_6t
Xbit_r164_c166 bl[166] br[166] wl[164] vdd gnd cell_6t
Xbit_r165_c166 bl[166] br[166] wl[165] vdd gnd cell_6t
Xbit_r166_c166 bl[166] br[166] wl[166] vdd gnd cell_6t
Xbit_r167_c166 bl[166] br[166] wl[167] vdd gnd cell_6t
Xbit_r168_c166 bl[166] br[166] wl[168] vdd gnd cell_6t
Xbit_r169_c166 bl[166] br[166] wl[169] vdd gnd cell_6t
Xbit_r170_c166 bl[166] br[166] wl[170] vdd gnd cell_6t
Xbit_r171_c166 bl[166] br[166] wl[171] vdd gnd cell_6t
Xbit_r172_c166 bl[166] br[166] wl[172] vdd gnd cell_6t
Xbit_r173_c166 bl[166] br[166] wl[173] vdd gnd cell_6t
Xbit_r174_c166 bl[166] br[166] wl[174] vdd gnd cell_6t
Xbit_r175_c166 bl[166] br[166] wl[175] vdd gnd cell_6t
Xbit_r176_c166 bl[166] br[166] wl[176] vdd gnd cell_6t
Xbit_r177_c166 bl[166] br[166] wl[177] vdd gnd cell_6t
Xbit_r178_c166 bl[166] br[166] wl[178] vdd gnd cell_6t
Xbit_r179_c166 bl[166] br[166] wl[179] vdd gnd cell_6t
Xbit_r180_c166 bl[166] br[166] wl[180] vdd gnd cell_6t
Xbit_r181_c166 bl[166] br[166] wl[181] vdd gnd cell_6t
Xbit_r182_c166 bl[166] br[166] wl[182] vdd gnd cell_6t
Xbit_r183_c166 bl[166] br[166] wl[183] vdd gnd cell_6t
Xbit_r184_c166 bl[166] br[166] wl[184] vdd gnd cell_6t
Xbit_r185_c166 bl[166] br[166] wl[185] vdd gnd cell_6t
Xbit_r186_c166 bl[166] br[166] wl[186] vdd gnd cell_6t
Xbit_r187_c166 bl[166] br[166] wl[187] vdd gnd cell_6t
Xbit_r188_c166 bl[166] br[166] wl[188] vdd gnd cell_6t
Xbit_r189_c166 bl[166] br[166] wl[189] vdd gnd cell_6t
Xbit_r190_c166 bl[166] br[166] wl[190] vdd gnd cell_6t
Xbit_r191_c166 bl[166] br[166] wl[191] vdd gnd cell_6t
Xbit_r192_c166 bl[166] br[166] wl[192] vdd gnd cell_6t
Xbit_r193_c166 bl[166] br[166] wl[193] vdd gnd cell_6t
Xbit_r194_c166 bl[166] br[166] wl[194] vdd gnd cell_6t
Xbit_r195_c166 bl[166] br[166] wl[195] vdd gnd cell_6t
Xbit_r196_c166 bl[166] br[166] wl[196] vdd gnd cell_6t
Xbit_r197_c166 bl[166] br[166] wl[197] vdd gnd cell_6t
Xbit_r198_c166 bl[166] br[166] wl[198] vdd gnd cell_6t
Xbit_r199_c166 bl[166] br[166] wl[199] vdd gnd cell_6t
Xbit_r200_c166 bl[166] br[166] wl[200] vdd gnd cell_6t
Xbit_r201_c166 bl[166] br[166] wl[201] vdd gnd cell_6t
Xbit_r202_c166 bl[166] br[166] wl[202] vdd gnd cell_6t
Xbit_r203_c166 bl[166] br[166] wl[203] vdd gnd cell_6t
Xbit_r204_c166 bl[166] br[166] wl[204] vdd gnd cell_6t
Xbit_r205_c166 bl[166] br[166] wl[205] vdd gnd cell_6t
Xbit_r206_c166 bl[166] br[166] wl[206] vdd gnd cell_6t
Xbit_r207_c166 bl[166] br[166] wl[207] vdd gnd cell_6t
Xbit_r208_c166 bl[166] br[166] wl[208] vdd gnd cell_6t
Xbit_r209_c166 bl[166] br[166] wl[209] vdd gnd cell_6t
Xbit_r210_c166 bl[166] br[166] wl[210] vdd gnd cell_6t
Xbit_r211_c166 bl[166] br[166] wl[211] vdd gnd cell_6t
Xbit_r212_c166 bl[166] br[166] wl[212] vdd gnd cell_6t
Xbit_r213_c166 bl[166] br[166] wl[213] vdd gnd cell_6t
Xbit_r214_c166 bl[166] br[166] wl[214] vdd gnd cell_6t
Xbit_r215_c166 bl[166] br[166] wl[215] vdd gnd cell_6t
Xbit_r216_c166 bl[166] br[166] wl[216] vdd gnd cell_6t
Xbit_r217_c166 bl[166] br[166] wl[217] vdd gnd cell_6t
Xbit_r218_c166 bl[166] br[166] wl[218] vdd gnd cell_6t
Xbit_r219_c166 bl[166] br[166] wl[219] vdd gnd cell_6t
Xbit_r220_c166 bl[166] br[166] wl[220] vdd gnd cell_6t
Xbit_r221_c166 bl[166] br[166] wl[221] vdd gnd cell_6t
Xbit_r222_c166 bl[166] br[166] wl[222] vdd gnd cell_6t
Xbit_r223_c166 bl[166] br[166] wl[223] vdd gnd cell_6t
Xbit_r224_c166 bl[166] br[166] wl[224] vdd gnd cell_6t
Xbit_r225_c166 bl[166] br[166] wl[225] vdd gnd cell_6t
Xbit_r226_c166 bl[166] br[166] wl[226] vdd gnd cell_6t
Xbit_r227_c166 bl[166] br[166] wl[227] vdd gnd cell_6t
Xbit_r228_c166 bl[166] br[166] wl[228] vdd gnd cell_6t
Xbit_r229_c166 bl[166] br[166] wl[229] vdd gnd cell_6t
Xbit_r230_c166 bl[166] br[166] wl[230] vdd gnd cell_6t
Xbit_r231_c166 bl[166] br[166] wl[231] vdd gnd cell_6t
Xbit_r232_c166 bl[166] br[166] wl[232] vdd gnd cell_6t
Xbit_r233_c166 bl[166] br[166] wl[233] vdd gnd cell_6t
Xbit_r234_c166 bl[166] br[166] wl[234] vdd gnd cell_6t
Xbit_r235_c166 bl[166] br[166] wl[235] vdd gnd cell_6t
Xbit_r236_c166 bl[166] br[166] wl[236] vdd gnd cell_6t
Xbit_r237_c166 bl[166] br[166] wl[237] vdd gnd cell_6t
Xbit_r238_c166 bl[166] br[166] wl[238] vdd gnd cell_6t
Xbit_r239_c166 bl[166] br[166] wl[239] vdd gnd cell_6t
Xbit_r240_c166 bl[166] br[166] wl[240] vdd gnd cell_6t
Xbit_r241_c166 bl[166] br[166] wl[241] vdd gnd cell_6t
Xbit_r242_c166 bl[166] br[166] wl[242] vdd gnd cell_6t
Xbit_r243_c166 bl[166] br[166] wl[243] vdd gnd cell_6t
Xbit_r244_c166 bl[166] br[166] wl[244] vdd gnd cell_6t
Xbit_r245_c166 bl[166] br[166] wl[245] vdd gnd cell_6t
Xbit_r246_c166 bl[166] br[166] wl[246] vdd gnd cell_6t
Xbit_r247_c166 bl[166] br[166] wl[247] vdd gnd cell_6t
Xbit_r248_c166 bl[166] br[166] wl[248] vdd gnd cell_6t
Xbit_r249_c166 bl[166] br[166] wl[249] vdd gnd cell_6t
Xbit_r250_c166 bl[166] br[166] wl[250] vdd gnd cell_6t
Xbit_r251_c166 bl[166] br[166] wl[251] vdd gnd cell_6t
Xbit_r252_c166 bl[166] br[166] wl[252] vdd gnd cell_6t
Xbit_r253_c166 bl[166] br[166] wl[253] vdd gnd cell_6t
Xbit_r254_c166 bl[166] br[166] wl[254] vdd gnd cell_6t
Xbit_r255_c166 bl[166] br[166] wl[255] vdd gnd cell_6t
Xbit_r0_c167 bl[167] br[167] wl[0] vdd gnd cell_6t
Xbit_r1_c167 bl[167] br[167] wl[1] vdd gnd cell_6t
Xbit_r2_c167 bl[167] br[167] wl[2] vdd gnd cell_6t
Xbit_r3_c167 bl[167] br[167] wl[3] vdd gnd cell_6t
Xbit_r4_c167 bl[167] br[167] wl[4] vdd gnd cell_6t
Xbit_r5_c167 bl[167] br[167] wl[5] vdd gnd cell_6t
Xbit_r6_c167 bl[167] br[167] wl[6] vdd gnd cell_6t
Xbit_r7_c167 bl[167] br[167] wl[7] vdd gnd cell_6t
Xbit_r8_c167 bl[167] br[167] wl[8] vdd gnd cell_6t
Xbit_r9_c167 bl[167] br[167] wl[9] vdd gnd cell_6t
Xbit_r10_c167 bl[167] br[167] wl[10] vdd gnd cell_6t
Xbit_r11_c167 bl[167] br[167] wl[11] vdd gnd cell_6t
Xbit_r12_c167 bl[167] br[167] wl[12] vdd gnd cell_6t
Xbit_r13_c167 bl[167] br[167] wl[13] vdd gnd cell_6t
Xbit_r14_c167 bl[167] br[167] wl[14] vdd gnd cell_6t
Xbit_r15_c167 bl[167] br[167] wl[15] vdd gnd cell_6t
Xbit_r16_c167 bl[167] br[167] wl[16] vdd gnd cell_6t
Xbit_r17_c167 bl[167] br[167] wl[17] vdd gnd cell_6t
Xbit_r18_c167 bl[167] br[167] wl[18] vdd gnd cell_6t
Xbit_r19_c167 bl[167] br[167] wl[19] vdd gnd cell_6t
Xbit_r20_c167 bl[167] br[167] wl[20] vdd gnd cell_6t
Xbit_r21_c167 bl[167] br[167] wl[21] vdd gnd cell_6t
Xbit_r22_c167 bl[167] br[167] wl[22] vdd gnd cell_6t
Xbit_r23_c167 bl[167] br[167] wl[23] vdd gnd cell_6t
Xbit_r24_c167 bl[167] br[167] wl[24] vdd gnd cell_6t
Xbit_r25_c167 bl[167] br[167] wl[25] vdd gnd cell_6t
Xbit_r26_c167 bl[167] br[167] wl[26] vdd gnd cell_6t
Xbit_r27_c167 bl[167] br[167] wl[27] vdd gnd cell_6t
Xbit_r28_c167 bl[167] br[167] wl[28] vdd gnd cell_6t
Xbit_r29_c167 bl[167] br[167] wl[29] vdd gnd cell_6t
Xbit_r30_c167 bl[167] br[167] wl[30] vdd gnd cell_6t
Xbit_r31_c167 bl[167] br[167] wl[31] vdd gnd cell_6t
Xbit_r32_c167 bl[167] br[167] wl[32] vdd gnd cell_6t
Xbit_r33_c167 bl[167] br[167] wl[33] vdd gnd cell_6t
Xbit_r34_c167 bl[167] br[167] wl[34] vdd gnd cell_6t
Xbit_r35_c167 bl[167] br[167] wl[35] vdd gnd cell_6t
Xbit_r36_c167 bl[167] br[167] wl[36] vdd gnd cell_6t
Xbit_r37_c167 bl[167] br[167] wl[37] vdd gnd cell_6t
Xbit_r38_c167 bl[167] br[167] wl[38] vdd gnd cell_6t
Xbit_r39_c167 bl[167] br[167] wl[39] vdd gnd cell_6t
Xbit_r40_c167 bl[167] br[167] wl[40] vdd gnd cell_6t
Xbit_r41_c167 bl[167] br[167] wl[41] vdd gnd cell_6t
Xbit_r42_c167 bl[167] br[167] wl[42] vdd gnd cell_6t
Xbit_r43_c167 bl[167] br[167] wl[43] vdd gnd cell_6t
Xbit_r44_c167 bl[167] br[167] wl[44] vdd gnd cell_6t
Xbit_r45_c167 bl[167] br[167] wl[45] vdd gnd cell_6t
Xbit_r46_c167 bl[167] br[167] wl[46] vdd gnd cell_6t
Xbit_r47_c167 bl[167] br[167] wl[47] vdd gnd cell_6t
Xbit_r48_c167 bl[167] br[167] wl[48] vdd gnd cell_6t
Xbit_r49_c167 bl[167] br[167] wl[49] vdd gnd cell_6t
Xbit_r50_c167 bl[167] br[167] wl[50] vdd gnd cell_6t
Xbit_r51_c167 bl[167] br[167] wl[51] vdd gnd cell_6t
Xbit_r52_c167 bl[167] br[167] wl[52] vdd gnd cell_6t
Xbit_r53_c167 bl[167] br[167] wl[53] vdd gnd cell_6t
Xbit_r54_c167 bl[167] br[167] wl[54] vdd gnd cell_6t
Xbit_r55_c167 bl[167] br[167] wl[55] vdd gnd cell_6t
Xbit_r56_c167 bl[167] br[167] wl[56] vdd gnd cell_6t
Xbit_r57_c167 bl[167] br[167] wl[57] vdd gnd cell_6t
Xbit_r58_c167 bl[167] br[167] wl[58] vdd gnd cell_6t
Xbit_r59_c167 bl[167] br[167] wl[59] vdd gnd cell_6t
Xbit_r60_c167 bl[167] br[167] wl[60] vdd gnd cell_6t
Xbit_r61_c167 bl[167] br[167] wl[61] vdd gnd cell_6t
Xbit_r62_c167 bl[167] br[167] wl[62] vdd gnd cell_6t
Xbit_r63_c167 bl[167] br[167] wl[63] vdd gnd cell_6t
Xbit_r64_c167 bl[167] br[167] wl[64] vdd gnd cell_6t
Xbit_r65_c167 bl[167] br[167] wl[65] vdd gnd cell_6t
Xbit_r66_c167 bl[167] br[167] wl[66] vdd gnd cell_6t
Xbit_r67_c167 bl[167] br[167] wl[67] vdd gnd cell_6t
Xbit_r68_c167 bl[167] br[167] wl[68] vdd gnd cell_6t
Xbit_r69_c167 bl[167] br[167] wl[69] vdd gnd cell_6t
Xbit_r70_c167 bl[167] br[167] wl[70] vdd gnd cell_6t
Xbit_r71_c167 bl[167] br[167] wl[71] vdd gnd cell_6t
Xbit_r72_c167 bl[167] br[167] wl[72] vdd gnd cell_6t
Xbit_r73_c167 bl[167] br[167] wl[73] vdd gnd cell_6t
Xbit_r74_c167 bl[167] br[167] wl[74] vdd gnd cell_6t
Xbit_r75_c167 bl[167] br[167] wl[75] vdd gnd cell_6t
Xbit_r76_c167 bl[167] br[167] wl[76] vdd gnd cell_6t
Xbit_r77_c167 bl[167] br[167] wl[77] vdd gnd cell_6t
Xbit_r78_c167 bl[167] br[167] wl[78] vdd gnd cell_6t
Xbit_r79_c167 bl[167] br[167] wl[79] vdd gnd cell_6t
Xbit_r80_c167 bl[167] br[167] wl[80] vdd gnd cell_6t
Xbit_r81_c167 bl[167] br[167] wl[81] vdd gnd cell_6t
Xbit_r82_c167 bl[167] br[167] wl[82] vdd gnd cell_6t
Xbit_r83_c167 bl[167] br[167] wl[83] vdd gnd cell_6t
Xbit_r84_c167 bl[167] br[167] wl[84] vdd gnd cell_6t
Xbit_r85_c167 bl[167] br[167] wl[85] vdd gnd cell_6t
Xbit_r86_c167 bl[167] br[167] wl[86] vdd gnd cell_6t
Xbit_r87_c167 bl[167] br[167] wl[87] vdd gnd cell_6t
Xbit_r88_c167 bl[167] br[167] wl[88] vdd gnd cell_6t
Xbit_r89_c167 bl[167] br[167] wl[89] vdd gnd cell_6t
Xbit_r90_c167 bl[167] br[167] wl[90] vdd gnd cell_6t
Xbit_r91_c167 bl[167] br[167] wl[91] vdd gnd cell_6t
Xbit_r92_c167 bl[167] br[167] wl[92] vdd gnd cell_6t
Xbit_r93_c167 bl[167] br[167] wl[93] vdd gnd cell_6t
Xbit_r94_c167 bl[167] br[167] wl[94] vdd gnd cell_6t
Xbit_r95_c167 bl[167] br[167] wl[95] vdd gnd cell_6t
Xbit_r96_c167 bl[167] br[167] wl[96] vdd gnd cell_6t
Xbit_r97_c167 bl[167] br[167] wl[97] vdd gnd cell_6t
Xbit_r98_c167 bl[167] br[167] wl[98] vdd gnd cell_6t
Xbit_r99_c167 bl[167] br[167] wl[99] vdd gnd cell_6t
Xbit_r100_c167 bl[167] br[167] wl[100] vdd gnd cell_6t
Xbit_r101_c167 bl[167] br[167] wl[101] vdd gnd cell_6t
Xbit_r102_c167 bl[167] br[167] wl[102] vdd gnd cell_6t
Xbit_r103_c167 bl[167] br[167] wl[103] vdd gnd cell_6t
Xbit_r104_c167 bl[167] br[167] wl[104] vdd gnd cell_6t
Xbit_r105_c167 bl[167] br[167] wl[105] vdd gnd cell_6t
Xbit_r106_c167 bl[167] br[167] wl[106] vdd gnd cell_6t
Xbit_r107_c167 bl[167] br[167] wl[107] vdd gnd cell_6t
Xbit_r108_c167 bl[167] br[167] wl[108] vdd gnd cell_6t
Xbit_r109_c167 bl[167] br[167] wl[109] vdd gnd cell_6t
Xbit_r110_c167 bl[167] br[167] wl[110] vdd gnd cell_6t
Xbit_r111_c167 bl[167] br[167] wl[111] vdd gnd cell_6t
Xbit_r112_c167 bl[167] br[167] wl[112] vdd gnd cell_6t
Xbit_r113_c167 bl[167] br[167] wl[113] vdd gnd cell_6t
Xbit_r114_c167 bl[167] br[167] wl[114] vdd gnd cell_6t
Xbit_r115_c167 bl[167] br[167] wl[115] vdd gnd cell_6t
Xbit_r116_c167 bl[167] br[167] wl[116] vdd gnd cell_6t
Xbit_r117_c167 bl[167] br[167] wl[117] vdd gnd cell_6t
Xbit_r118_c167 bl[167] br[167] wl[118] vdd gnd cell_6t
Xbit_r119_c167 bl[167] br[167] wl[119] vdd gnd cell_6t
Xbit_r120_c167 bl[167] br[167] wl[120] vdd gnd cell_6t
Xbit_r121_c167 bl[167] br[167] wl[121] vdd gnd cell_6t
Xbit_r122_c167 bl[167] br[167] wl[122] vdd gnd cell_6t
Xbit_r123_c167 bl[167] br[167] wl[123] vdd gnd cell_6t
Xbit_r124_c167 bl[167] br[167] wl[124] vdd gnd cell_6t
Xbit_r125_c167 bl[167] br[167] wl[125] vdd gnd cell_6t
Xbit_r126_c167 bl[167] br[167] wl[126] vdd gnd cell_6t
Xbit_r127_c167 bl[167] br[167] wl[127] vdd gnd cell_6t
Xbit_r128_c167 bl[167] br[167] wl[128] vdd gnd cell_6t
Xbit_r129_c167 bl[167] br[167] wl[129] vdd gnd cell_6t
Xbit_r130_c167 bl[167] br[167] wl[130] vdd gnd cell_6t
Xbit_r131_c167 bl[167] br[167] wl[131] vdd gnd cell_6t
Xbit_r132_c167 bl[167] br[167] wl[132] vdd gnd cell_6t
Xbit_r133_c167 bl[167] br[167] wl[133] vdd gnd cell_6t
Xbit_r134_c167 bl[167] br[167] wl[134] vdd gnd cell_6t
Xbit_r135_c167 bl[167] br[167] wl[135] vdd gnd cell_6t
Xbit_r136_c167 bl[167] br[167] wl[136] vdd gnd cell_6t
Xbit_r137_c167 bl[167] br[167] wl[137] vdd gnd cell_6t
Xbit_r138_c167 bl[167] br[167] wl[138] vdd gnd cell_6t
Xbit_r139_c167 bl[167] br[167] wl[139] vdd gnd cell_6t
Xbit_r140_c167 bl[167] br[167] wl[140] vdd gnd cell_6t
Xbit_r141_c167 bl[167] br[167] wl[141] vdd gnd cell_6t
Xbit_r142_c167 bl[167] br[167] wl[142] vdd gnd cell_6t
Xbit_r143_c167 bl[167] br[167] wl[143] vdd gnd cell_6t
Xbit_r144_c167 bl[167] br[167] wl[144] vdd gnd cell_6t
Xbit_r145_c167 bl[167] br[167] wl[145] vdd gnd cell_6t
Xbit_r146_c167 bl[167] br[167] wl[146] vdd gnd cell_6t
Xbit_r147_c167 bl[167] br[167] wl[147] vdd gnd cell_6t
Xbit_r148_c167 bl[167] br[167] wl[148] vdd gnd cell_6t
Xbit_r149_c167 bl[167] br[167] wl[149] vdd gnd cell_6t
Xbit_r150_c167 bl[167] br[167] wl[150] vdd gnd cell_6t
Xbit_r151_c167 bl[167] br[167] wl[151] vdd gnd cell_6t
Xbit_r152_c167 bl[167] br[167] wl[152] vdd gnd cell_6t
Xbit_r153_c167 bl[167] br[167] wl[153] vdd gnd cell_6t
Xbit_r154_c167 bl[167] br[167] wl[154] vdd gnd cell_6t
Xbit_r155_c167 bl[167] br[167] wl[155] vdd gnd cell_6t
Xbit_r156_c167 bl[167] br[167] wl[156] vdd gnd cell_6t
Xbit_r157_c167 bl[167] br[167] wl[157] vdd gnd cell_6t
Xbit_r158_c167 bl[167] br[167] wl[158] vdd gnd cell_6t
Xbit_r159_c167 bl[167] br[167] wl[159] vdd gnd cell_6t
Xbit_r160_c167 bl[167] br[167] wl[160] vdd gnd cell_6t
Xbit_r161_c167 bl[167] br[167] wl[161] vdd gnd cell_6t
Xbit_r162_c167 bl[167] br[167] wl[162] vdd gnd cell_6t
Xbit_r163_c167 bl[167] br[167] wl[163] vdd gnd cell_6t
Xbit_r164_c167 bl[167] br[167] wl[164] vdd gnd cell_6t
Xbit_r165_c167 bl[167] br[167] wl[165] vdd gnd cell_6t
Xbit_r166_c167 bl[167] br[167] wl[166] vdd gnd cell_6t
Xbit_r167_c167 bl[167] br[167] wl[167] vdd gnd cell_6t
Xbit_r168_c167 bl[167] br[167] wl[168] vdd gnd cell_6t
Xbit_r169_c167 bl[167] br[167] wl[169] vdd gnd cell_6t
Xbit_r170_c167 bl[167] br[167] wl[170] vdd gnd cell_6t
Xbit_r171_c167 bl[167] br[167] wl[171] vdd gnd cell_6t
Xbit_r172_c167 bl[167] br[167] wl[172] vdd gnd cell_6t
Xbit_r173_c167 bl[167] br[167] wl[173] vdd gnd cell_6t
Xbit_r174_c167 bl[167] br[167] wl[174] vdd gnd cell_6t
Xbit_r175_c167 bl[167] br[167] wl[175] vdd gnd cell_6t
Xbit_r176_c167 bl[167] br[167] wl[176] vdd gnd cell_6t
Xbit_r177_c167 bl[167] br[167] wl[177] vdd gnd cell_6t
Xbit_r178_c167 bl[167] br[167] wl[178] vdd gnd cell_6t
Xbit_r179_c167 bl[167] br[167] wl[179] vdd gnd cell_6t
Xbit_r180_c167 bl[167] br[167] wl[180] vdd gnd cell_6t
Xbit_r181_c167 bl[167] br[167] wl[181] vdd gnd cell_6t
Xbit_r182_c167 bl[167] br[167] wl[182] vdd gnd cell_6t
Xbit_r183_c167 bl[167] br[167] wl[183] vdd gnd cell_6t
Xbit_r184_c167 bl[167] br[167] wl[184] vdd gnd cell_6t
Xbit_r185_c167 bl[167] br[167] wl[185] vdd gnd cell_6t
Xbit_r186_c167 bl[167] br[167] wl[186] vdd gnd cell_6t
Xbit_r187_c167 bl[167] br[167] wl[187] vdd gnd cell_6t
Xbit_r188_c167 bl[167] br[167] wl[188] vdd gnd cell_6t
Xbit_r189_c167 bl[167] br[167] wl[189] vdd gnd cell_6t
Xbit_r190_c167 bl[167] br[167] wl[190] vdd gnd cell_6t
Xbit_r191_c167 bl[167] br[167] wl[191] vdd gnd cell_6t
Xbit_r192_c167 bl[167] br[167] wl[192] vdd gnd cell_6t
Xbit_r193_c167 bl[167] br[167] wl[193] vdd gnd cell_6t
Xbit_r194_c167 bl[167] br[167] wl[194] vdd gnd cell_6t
Xbit_r195_c167 bl[167] br[167] wl[195] vdd gnd cell_6t
Xbit_r196_c167 bl[167] br[167] wl[196] vdd gnd cell_6t
Xbit_r197_c167 bl[167] br[167] wl[197] vdd gnd cell_6t
Xbit_r198_c167 bl[167] br[167] wl[198] vdd gnd cell_6t
Xbit_r199_c167 bl[167] br[167] wl[199] vdd gnd cell_6t
Xbit_r200_c167 bl[167] br[167] wl[200] vdd gnd cell_6t
Xbit_r201_c167 bl[167] br[167] wl[201] vdd gnd cell_6t
Xbit_r202_c167 bl[167] br[167] wl[202] vdd gnd cell_6t
Xbit_r203_c167 bl[167] br[167] wl[203] vdd gnd cell_6t
Xbit_r204_c167 bl[167] br[167] wl[204] vdd gnd cell_6t
Xbit_r205_c167 bl[167] br[167] wl[205] vdd gnd cell_6t
Xbit_r206_c167 bl[167] br[167] wl[206] vdd gnd cell_6t
Xbit_r207_c167 bl[167] br[167] wl[207] vdd gnd cell_6t
Xbit_r208_c167 bl[167] br[167] wl[208] vdd gnd cell_6t
Xbit_r209_c167 bl[167] br[167] wl[209] vdd gnd cell_6t
Xbit_r210_c167 bl[167] br[167] wl[210] vdd gnd cell_6t
Xbit_r211_c167 bl[167] br[167] wl[211] vdd gnd cell_6t
Xbit_r212_c167 bl[167] br[167] wl[212] vdd gnd cell_6t
Xbit_r213_c167 bl[167] br[167] wl[213] vdd gnd cell_6t
Xbit_r214_c167 bl[167] br[167] wl[214] vdd gnd cell_6t
Xbit_r215_c167 bl[167] br[167] wl[215] vdd gnd cell_6t
Xbit_r216_c167 bl[167] br[167] wl[216] vdd gnd cell_6t
Xbit_r217_c167 bl[167] br[167] wl[217] vdd gnd cell_6t
Xbit_r218_c167 bl[167] br[167] wl[218] vdd gnd cell_6t
Xbit_r219_c167 bl[167] br[167] wl[219] vdd gnd cell_6t
Xbit_r220_c167 bl[167] br[167] wl[220] vdd gnd cell_6t
Xbit_r221_c167 bl[167] br[167] wl[221] vdd gnd cell_6t
Xbit_r222_c167 bl[167] br[167] wl[222] vdd gnd cell_6t
Xbit_r223_c167 bl[167] br[167] wl[223] vdd gnd cell_6t
Xbit_r224_c167 bl[167] br[167] wl[224] vdd gnd cell_6t
Xbit_r225_c167 bl[167] br[167] wl[225] vdd gnd cell_6t
Xbit_r226_c167 bl[167] br[167] wl[226] vdd gnd cell_6t
Xbit_r227_c167 bl[167] br[167] wl[227] vdd gnd cell_6t
Xbit_r228_c167 bl[167] br[167] wl[228] vdd gnd cell_6t
Xbit_r229_c167 bl[167] br[167] wl[229] vdd gnd cell_6t
Xbit_r230_c167 bl[167] br[167] wl[230] vdd gnd cell_6t
Xbit_r231_c167 bl[167] br[167] wl[231] vdd gnd cell_6t
Xbit_r232_c167 bl[167] br[167] wl[232] vdd gnd cell_6t
Xbit_r233_c167 bl[167] br[167] wl[233] vdd gnd cell_6t
Xbit_r234_c167 bl[167] br[167] wl[234] vdd gnd cell_6t
Xbit_r235_c167 bl[167] br[167] wl[235] vdd gnd cell_6t
Xbit_r236_c167 bl[167] br[167] wl[236] vdd gnd cell_6t
Xbit_r237_c167 bl[167] br[167] wl[237] vdd gnd cell_6t
Xbit_r238_c167 bl[167] br[167] wl[238] vdd gnd cell_6t
Xbit_r239_c167 bl[167] br[167] wl[239] vdd gnd cell_6t
Xbit_r240_c167 bl[167] br[167] wl[240] vdd gnd cell_6t
Xbit_r241_c167 bl[167] br[167] wl[241] vdd gnd cell_6t
Xbit_r242_c167 bl[167] br[167] wl[242] vdd gnd cell_6t
Xbit_r243_c167 bl[167] br[167] wl[243] vdd gnd cell_6t
Xbit_r244_c167 bl[167] br[167] wl[244] vdd gnd cell_6t
Xbit_r245_c167 bl[167] br[167] wl[245] vdd gnd cell_6t
Xbit_r246_c167 bl[167] br[167] wl[246] vdd gnd cell_6t
Xbit_r247_c167 bl[167] br[167] wl[247] vdd gnd cell_6t
Xbit_r248_c167 bl[167] br[167] wl[248] vdd gnd cell_6t
Xbit_r249_c167 bl[167] br[167] wl[249] vdd gnd cell_6t
Xbit_r250_c167 bl[167] br[167] wl[250] vdd gnd cell_6t
Xbit_r251_c167 bl[167] br[167] wl[251] vdd gnd cell_6t
Xbit_r252_c167 bl[167] br[167] wl[252] vdd gnd cell_6t
Xbit_r253_c167 bl[167] br[167] wl[253] vdd gnd cell_6t
Xbit_r254_c167 bl[167] br[167] wl[254] vdd gnd cell_6t
Xbit_r255_c167 bl[167] br[167] wl[255] vdd gnd cell_6t
Xbit_r0_c168 bl[168] br[168] wl[0] vdd gnd cell_6t
Xbit_r1_c168 bl[168] br[168] wl[1] vdd gnd cell_6t
Xbit_r2_c168 bl[168] br[168] wl[2] vdd gnd cell_6t
Xbit_r3_c168 bl[168] br[168] wl[3] vdd gnd cell_6t
Xbit_r4_c168 bl[168] br[168] wl[4] vdd gnd cell_6t
Xbit_r5_c168 bl[168] br[168] wl[5] vdd gnd cell_6t
Xbit_r6_c168 bl[168] br[168] wl[6] vdd gnd cell_6t
Xbit_r7_c168 bl[168] br[168] wl[7] vdd gnd cell_6t
Xbit_r8_c168 bl[168] br[168] wl[8] vdd gnd cell_6t
Xbit_r9_c168 bl[168] br[168] wl[9] vdd gnd cell_6t
Xbit_r10_c168 bl[168] br[168] wl[10] vdd gnd cell_6t
Xbit_r11_c168 bl[168] br[168] wl[11] vdd gnd cell_6t
Xbit_r12_c168 bl[168] br[168] wl[12] vdd gnd cell_6t
Xbit_r13_c168 bl[168] br[168] wl[13] vdd gnd cell_6t
Xbit_r14_c168 bl[168] br[168] wl[14] vdd gnd cell_6t
Xbit_r15_c168 bl[168] br[168] wl[15] vdd gnd cell_6t
Xbit_r16_c168 bl[168] br[168] wl[16] vdd gnd cell_6t
Xbit_r17_c168 bl[168] br[168] wl[17] vdd gnd cell_6t
Xbit_r18_c168 bl[168] br[168] wl[18] vdd gnd cell_6t
Xbit_r19_c168 bl[168] br[168] wl[19] vdd gnd cell_6t
Xbit_r20_c168 bl[168] br[168] wl[20] vdd gnd cell_6t
Xbit_r21_c168 bl[168] br[168] wl[21] vdd gnd cell_6t
Xbit_r22_c168 bl[168] br[168] wl[22] vdd gnd cell_6t
Xbit_r23_c168 bl[168] br[168] wl[23] vdd gnd cell_6t
Xbit_r24_c168 bl[168] br[168] wl[24] vdd gnd cell_6t
Xbit_r25_c168 bl[168] br[168] wl[25] vdd gnd cell_6t
Xbit_r26_c168 bl[168] br[168] wl[26] vdd gnd cell_6t
Xbit_r27_c168 bl[168] br[168] wl[27] vdd gnd cell_6t
Xbit_r28_c168 bl[168] br[168] wl[28] vdd gnd cell_6t
Xbit_r29_c168 bl[168] br[168] wl[29] vdd gnd cell_6t
Xbit_r30_c168 bl[168] br[168] wl[30] vdd gnd cell_6t
Xbit_r31_c168 bl[168] br[168] wl[31] vdd gnd cell_6t
Xbit_r32_c168 bl[168] br[168] wl[32] vdd gnd cell_6t
Xbit_r33_c168 bl[168] br[168] wl[33] vdd gnd cell_6t
Xbit_r34_c168 bl[168] br[168] wl[34] vdd gnd cell_6t
Xbit_r35_c168 bl[168] br[168] wl[35] vdd gnd cell_6t
Xbit_r36_c168 bl[168] br[168] wl[36] vdd gnd cell_6t
Xbit_r37_c168 bl[168] br[168] wl[37] vdd gnd cell_6t
Xbit_r38_c168 bl[168] br[168] wl[38] vdd gnd cell_6t
Xbit_r39_c168 bl[168] br[168] wl[39] vdd gnd cell_6t
Xbit_r40_c168 bl[168] br[168] wl[40] vdd gnd cell_6t
Xbit_r41_c168 bl[168] br[168] wl[41] vdd gnd cell_6t
Xbit_r42_c168 bl[168] br[168] wl[42] vdd gnd cell_6t
Xbit_r43_c168 bl[168] br[168] wl[43] vdd gnd cell_6t
Xbit_r44_c168 bl[168] br[168] wl[44] vdd gnd cell_6t
Xbit_r45_c168 bl[168] br[168] wl[45] vdd gnd cell_6t
Xbit_r46_c168 bl[168] br[168] wl[46] vdd gnd cell_6t
Xbit_r47_c168 bl[168] br[168] wl[47] vdd gnd cell_6t
Xbit_r48_c168 bl[168] br[168] wl[48] vdd gnd cell_6t
Xbit_r49_c168 bl[168] br[168] wl[49] vdd gnd cell_6t
Xbit_r50_c168 bl[168] br[168] wl[50] vdd gnd cell_6t
Xbit_r51_c168 bl[168] br[168] wl[51] vdd gnd cell_6t
Xbit_r52_c168 bl[168] br[168] wl[52] vdd gnd cell_6t
Xbit_r53_c168 bl[168] br[168] wl[53] vdd gnd cell_6t
Xbit_r54_c168 bl[168] br[168] wl[54] vdd gnd cell_6t
Xbit_r55_c168 bl[168] br[168] wl[55] vdd gnd cell_6t
Xbit_r56_c168 bl[168] br[168] wl[56] vdd gnd cell_6t
Xbit_r57_c168 bl[168] br[168] wl[57] vdd gnd cell_6t
Xbit_r58_c168 bl[168] br[168] wl[58] vdd gnd cell_6t
Xbit_r59_c168 bl[168] br[168] wl[59] vdd gnd cell_6t
Xbit_r60_c168 bl[168] br[168] wl[60] vdd gnd cell_6t
Xbit_r61_c168 bl[168] br[168] wl[61] vdd gnd cell_6t
Xbit_r62_c168 bl[168] br[168] wl[62] vdd gnd cell_6t
Xbit_r63_c168 bl[168] br[168] wl[63] vdd gnd cell_6t
Xbit_r64_c168 bl[168] br[168] wl[64] vdd gnd cell_6t
Xbit_r65_c168 bl[168] br[168] wl[65] vdd gnd cell_6t
Xbit_r66_c168 bl[168] br[168] wl[66] vdd gnd cell_6t
Xbit_r67_c168 bl[168] br[168] wl[67] vdd gnd cell_6t
Xbit_r68_c168 bl[168] br[168] wl[68] vdd gnd cell_6t
Xbit_r69_c168 bl[168] br[168] wl[69] vdd gnd cell_6t
Xbit_r70_c168 bl[168] br[168] wl[70] vdd gnd cell_6t
Xbit_r71_c168 bl[168] br[168] wl[71] vdd gnd cell_6t
Xbit_r72_c168 bl[168] br[168] wl[72] vdd gnd cell_6t
Xbit_r73_c168 bl[168] br[168] wl[73] vdd gnd cell_6t
Xbit_r74_c168 bl[168] br[168] wl[74] vdd gnd cell_6t
Xbit_r75_c168 bl[168] br[168] wl[75] vdd gnd cell_6t
Xbit_r76_c168 bl[168] br[168] wl[76] vdd gnd cell_6t
Xbit_r77_c168 bl[168] br[168] wl[77] vdd gnd cell_6t
Xbit_r78_c168 bl[168] br[168] wl[78] vdd gnd cell_6t
Xbit_r79_c168 bl[168] br[168] wl[79] vdd gnd cell_6t
Xbit_r80_c168 bl[168] br[168] wl[80] vdd gnd cell_6t
Xbit_r81_c168 bl[168] br[168] wl[81] vdd gnd cell_6t
Xbit_r82_c168 bl[168] br[168] wl[82] vdd gnd cell_6t
Xbit_r83_c168 bl[168] br[168] wl[83] vdd gnd cell_6t
Xbit_r84_c168 bl[168] br[168] wl[84] vdd gnd cell_6t
Xbit_r85_c168 bl[168] br[168] wl[85] vdd gnd cell_6t
Xbit_r86_c168 bl[168] br[168] wl[86] vdd gnd cell_6t
Xbit_r87_c168 bl[168] br[168] wl[87] vdd gnd cell_6t
Xbit_r88_c168 bl[168] br[168] wl[88] vdd gnd cell_6t
Xbit_r89_c168 bl[168] br[168] wl[89] vdd gnd cell_6t
Xbit_r90_c168 bl[168] br[168] wl[90] vdd gnd cell_6t
Xbit_r91_c168 bl[168] br[168] wl[91] vdd gnd cell_6t
Xbit_r92_c168 bl[168] br[168] wl[92] vdd gnd cell_6t
Xbit_r93_c168 bl[168] br[168] wl[93] vdd gnd cell_6t
Xbit_r94_c168 bl[168] br[168] wl[94] vdd gnd cell_6t
Xbit_r95_c168 bl[168] br[168] wl[95] vdd gnd cell_6t
Xbit_r96_c168 bl[168] br[168] wl[96] vdd gnd cell_6t
Xbit_r97_c168 bl[168] br[168] wl[97] vdd gnd cell_6t
Xbit_r98_c168 bl[168] br[168] wl[98] vdd gnd cell_6t
Xbit_r99_c168 bl[168] br[168] wl[99] vdd gnd cell_6t
Xbit_r100_c168 bl[168] br[168] wl[100] vdd gnd cell_6t
Xbit_r101_c168 bl[168] br[168] wl[101] vdd gnd cell_6t
Xbit_r102_c168 bl[168] br[168] wl[102] vdd gnd cell_6t
Xbit_r103_c168 bl[168] br[168] wl[103] vdd gnd cell_6t
Xbit_r104_c168 bl[168] br[168] wl[104] vdd gnd cell_6t
Xbit_r105_c168 bl[168] br[168] wl[105] vdd gnd cell_6t
Xbit_r106_c168 bl[168] br[168] wl[106] vdd gnd cell_6t
Xbit_r107_c168 bl[168] br[168] wl[107] vdd gnd cell_6t
Xbit_r108_c168 bl[168] br[168] wl[108] vdd gnd cell_6t
Xbit_r109_c168 bl[168] br[168] wl[109] vdd gnd cell_6t
Xbit_r110_c168 bl[168] br[168] wl[110] vdd gnd cell_6t
Xbit_r111_c168 bl[168] br[168] wl[111] vdd gnd cell_6t
Xbit_r112_c168 bl[168] br[168] wl[112] vdd gnd cell_6t
Xbit_r113_c168 bl[168] br[168] wl[113] vdd gnd cell_6t
Xbit_r114_c168 bl[168] br[168] wl[114] vdd gnd cell_6t
Xbit_r115_c168 bl[168] br[168] wl[115] vdd gnd cell_6t
Xbit_r116_c168 bl[168] br[168] wl[116] vdd gnd cell_6t
Xbit_r117_c168 bl[168] br[168] wl[117] vdd gnd cell_6t
Xbit_r118_c168 bl[168] br[168] wl[118] vdd gnd cell_6t
Xbit_r119_c168 bl[168] br[168] wl[119] vdd gnd cell_6t
Xbit_r120_c168 bl[168] br[168] wl[120] vdd gnd cell_6t
Xbit_r121_c168 bl[168] br[168] wl[121] vdd gnd cell_6t
Xbit_r122_c168 bl[168] br[168] wl[122] vdd gnd cell_6t
Xbit_r123_c168 bl[168] br[168] wl[123] vdd gnd cell_6t
Xbit_r124_c168 bl[168] br[168] wl[124] vdd gnd cell_6t
Xbit_r125_c168 bl[168] br[168] wl[125] vdd gnd cell_6t
Xbit_r126_c168 bl[168] br[168] wl[126] vdd gnd cell_6t
Xbit_r127_c168 bl[168] br[168] wl[127] vdd gnd cell_6t
Xbit_r128_c168 bl[168] br[168] wl[128] vdd gnd cell_6t
Xbit_r129_c168 bl[168] br[168] wl[129] vdd gnd cell_6t
Xbit_r130_c168 bl[168] br[168] wl[130] vdd gnd cell_6t
Xbit_r131_c168 bl[168] br[168] wl[131] vdd gnd cell_6t
Xbit_r132_c168 bl[168] br[168] wl[132] vdd gnd cell_6t
Xbit_r133_c168 bl[168] br[168] wl[133] vdd gnd cell_6t
Xbit_r134_c168 bl[168] br[168] wl[134] vdd gnd cell_6t
Xbit_r135_c168 bl[168] br[168] wl[135] vdd gnd cell_6t
Xbit_r136_c168 bl[168] br[168] wl[136] vdd gnd cell_6t
Xbit_r137_c168 bl[168] br[168] wl[137] vdd gnd cell_6t
Xbit_r138_c168 bl[168] br[168] wl[138] vdd gnd cell_6t
Xbit_r139_c168 bl[168] br[168] wl[139] vdd gnd cell_6t
Xbit_r140_c168 bl[168] br[168] wl[140] vdd gnd cell_6t
Xbit_r141_c168 bl[168] br[168] wl[141] vdd gnd cell_6t
Xbit_r142_c168 bl[168] br[168] wl[142] vdd gnd cell_6t
Xbit_r143_c168 bl[168] br[168] wl[143] vdd gnd cell_6t
Xbit_r144_c168 bl[168] br[168] wl[144] vdd gnd cell_6t
Xbit_r145_c168 bl[168] br[168] wl[145] vdd gnd cell_6t
Xbit_r146_c168 bl[168] br[168] wl[146] vdd gnd cell_6t
Xbit_r147_c168 bl[168] br[168] wl[147] vdd gnd cell_6t
Xbit_r148_c168 bl[168] br[168] wl[148] vdd gnd cell_6t
Xbit_r149_c168 bl[168] br[168] wl[149] vdd gnd cell_6t
Xbit_r150_c168 bl[168] br[168] wl[150] vdd gnd cell_6t
Xbit_r151_c168 bl[168] br[168] wl[151] vdd gnd cell_6t
Xbit_r152_c168 bl[168] br[168] wl[152] vdd gnd cell_6t
Xbit_r153_c168 bl[168] br[168] wl[153] vdd gnd cell_6t
Xbit_r154_c168 bl[168] br[168] wl[154] vdd gnd cell_6t
Xbit_r155_c168 bl[168] br[168] wl[155] vdd gnd cell_6t
Xbit_r156_c168 bl[168] br[168] wl[156] vdd gnd cell_6t
Xbit_r157_c168 bl[168] br[168] wl[157] vdd gnd cell_6t
Xbit_r158_c168 bl[168] br[168] wl[158] vdd gnd cell_6t
Xbit_r159_c168 bl[168] br[168] wl[159] vdd gnd cell_6t
Xbit_r160_c168 bl[168] br[168] wl[160] vdd gnd cell_6t
Xbit_r161_c168 bl[168] br[168] wl[161] vdd gnd cell_6t
Xbit_r162_c168 bl[168] br[168] wl[162] vdd gnd cell_6t
Xbit_r163_c168 bl[168] br[168] wl[163] vdd gnd cell_6t
Xbit_r164_c168 bl[168] br[168] wl[164] vdd gnd cell_6t
Xbit_r165_c168 bl[168] br[168] wl[165] vdd gnd cell_6t
Xbit_r166_c168 bl[168] br[168] wl[166] vdd gnd cell_6t
Xbit_r167_c168 bl[168] br[168] wl[167] vdd gnd cell_6t
Xbit_r168_c168 bl[168] br[168] wl[168] vdd gnd cell_6t
Xbit_r169_c168 bl[168] br[168] wl[169] vdd gnd cell_6t
Xbit_r170_c168 bl[168] br[168] wl[170] vdd gnd cell_6t
Xbit_r171_c168 bl[168] br[168] wl[171] vdd gnd cell_6t
Xbit_r172_c168 bl[168] br[168] wl[172] vdd gnd cell_6t
Xbit_r173_c168 bl[168] br[168] wl[173] vdd gnd cell_6t
Xbit_r174_c168 bl[168] br[168] wl[174] vdd gnd cell_6t
Xbit_r175_c168 bl[168] br[168] wl[175] vdd gnd cell_6t
Xbit_r176_c168 bl[168] br[168] wl[176] vdd gnd cell_6t
Xbit_r177_c168 bl[168] br[168] wl[177] vdd gnd cell_6t
Xbit_r178_c168 bl[168] br[168] wl[178] vdd gnd cell_6t
Xbit_r179_c168 bl[168] br[168] wl[179] vdd gnd cell_6t
Xbit_r180_c168 bl[168] br[168] wl[180] vdd gnd cell_6t
Xbit_r181_c168 bl[168] br[168] wl[181] vdd gnd cell_6t
Xbit_r182_c168 bl[168] br[168] wl[182] vdd gnd cell_6t
Xbit_r183_c168 bl[168] br[168] wl[183] vdd gnd cell_6t
Xbit_r184_c168 bl[168] br[168] wl[184] vdd gnd cell_6t
Xbit_r185_c168 bl[168] br[168] wl[185] vdd gnd cell_6t
Xbit_r186_c168 bl[168] br[168] wl[186] vdd gnd cell_6t
Xbit_r187_c168 bl[168] br[168] wl[187] vdd gnd cell_6t
Xbit_r188_c168 bl[168] br[168] wl[188] vdd gnd cell_6t
Xbit_r189_c168 bl[168] br[168] wl[189] vdd gnd cell_6t
Xbit_r190_c168 bl[168] br[168] wl[190] vdd gnd cell_6t
Xbit_r191_c168 bl[168] br[168] wl[191] vdd gnd cell_6t
Xbit_r192_c168 bl[168] br[168] wl[192] vdd gnd cell_6t
Xbit_r193_c168 bl[168] br[168] wl[193] vdd gnd cell_6t
Xbit_r194_c168 bl[168] br[168] wl[194] vdd gnd cell_6t
Xbit_r195_c168 bl[168] br[168] wl[195] vdd gnd cell_6t
Xbit_r196_c168 bl[168] br[168] wl[196] vdd gnd cell_6t
Xbit_r197_c168 bl[168] br[168] wl[197] vdd gnd cell_6t
Xbit_r198_c168 bl[168] br[168] wl[198] vdd gnd cell_6t
Xbit_r199_c168 bl[168] br[168] wl[199] vdd gnd cell_6t
Xbit_r200_c168 bl[168] br[168] wl[200] vdd gnd cell_6t
Xbit_r201_c168 bl[168] br[168] wl[201] vdd gnd cell_6t
Xbit_r202_c168 bl[168] br[168] wl[202] vdd gnd cell_6t
Xbit_r203_c168 bl[168] br[168] wl[203] vdd gnd cell_6t
Xbit_r204_c168 bl[168] br[168] wl[204] vdd gnd cell_6t
Xbit_r205_c168 bl[168] br[168] wl[205] vdd gnd cell_6t
Xbit_r206_c168 bl[168] br[168] wl[206] vdd gnd cell_6t
Xbit_r207_c168 bl[168] br[168] wl[207] vdd gnd cell_6t
Xbit_r208_c168 bl[168] br[168] wl[208] vdd gnd cell_6t
Xbit_r209_c168 bl[168] br[168] wl[209] vdd gnd cell_6t
Xbit_r210_c168 bl[168] br[168] wl[210] vdd gnd cell_6t
Xbit_r211_c168 bl[168] br[168] wl[211] vdd gnd cell_6t
Xbit_r212_c168 bl[168] br[168] wl[212] vdd gnd cell_6t
Xbit_r213_c168 bl[168] br[168] wl[213] vdd gnd cell_6t
Xbit_r214_c168 bl[168] br[168] wl[214] vdd gnd cell_6t
Xbit_r215_c168 bl[168] br[168] wl[215] vdd gnd cell_6t
Xbit_r216_c168 bl[168] br[168] wl[216] vdd gnd cell_6t
Xbit_r217_c168 bl[168] br[168] wl[217] vdd gnd cell_6t
Xbit_r218_c168 bl[168] br[168] wl[218] vdd gnd cell_6t
Xbit_r219_c168 bl[168] br[168] wl[219] vdd gnd cell_6t
Xbit_r220_c168 bl[168] br[168] wl[220] vdd gnd cell_6t
Xbit_r221_c168 bl[168] br[168] wl[221] vdd gnd cell_6t
Xbit_r222_c168 bl[168] br[168] wl[222] vdd gnd cell_6t
Xbit_r223_c168 bl[168] br[168] wl[223] vdd gnd cell_6t
Xbit_r224_c168 bl[168] br[168] wl[224] vdd gnd cell_6t
Xbit_r225_c168 bl[168] br[168] wl[225] vdd gnd cell_6t
Xbit_r226_c168 bl[168] br[168] wl[226] vdd gnd cell_6t
Xbit_r227_c168 bl[168] br[168] wl[227] vdd gnd cell_6t
Xbit_r228_c168 bl[168] br[168] wl[228] vdd gnd cell_6t
Xbit_r229_c168 bl[168] br[168] wl[229] vdd gnd cell_6t
Xbit_r230_c168 bl[168] br[168] wl[230] vdd gnd cell_6t
Xbit_r231_c168 bl[168] br[168] wl[231] vdd gnd cell_6t
Xbit_r232_c168 bl[168] br[168] wl[232] vdd gnd cell_6t
Xbit_r233_c168 bl[168] br[168] wl[233] vdd gnd cell_6t
Xbit_r234_c168 bl[168] br[168] wl[234] vdd gnd cell_6t
Xbit_r235_c168 bl[168] br[168] wl[235] vdd gnd cell_6t
Xbit_r236_c168 bl[168] br[168] wl[236] vdd gnd cell_6t
Xbit_r237_c168 bl[168] br[168] wl[237] vdd gnd cell_6t
Xbit_r238_c168 bl[168] br[168] wl[238] vdd gnd cell_6t
Xbit_r239_c168 bl[168] br[168] wl[239] vdd gnd cell_6t
Xbit_r240_c168 bl[168] br[168] wl[240] vdd gnd cell_6t
Xbit_r241_c168 bl[168] br[168] wl[241] vdd gnd cell_6t
Xbit_r242_c168 bl[168] br[168] wl[242] vdd gnd cell_6t
Xbit_r243_c168 bl[168] br[168] wl[243] vdd gnd cell_6t
Xbit_r244_c168 bl[168] br[168] wl[244] vdd gnd cell_6t
Xbit_r245_c168 bl[168] br[168] wl[245] vdd gnd cell_6t
Xbit_r246_c168 bl[168] br[168] wl[246] vdd gnd cell_6t
Xbit_r247_c168 bl[168] br[168] wl[247] vdd gnd cell_6t
Xbit_r248_c168 bl[168] br[168] wl[248] vdd gnd cell_6t
Xbit_r249_c168 bl[168] br[168] wl[249] vdd gnd cell_6t
Xbit_r250_c168 bl[168] br[168] wl[250] vdd gnd cell_6t
Xbit_r251_c168 bl[168] br[168] wl[251] vdd gnd cell_6t
Xbit_r252_c168 bl[168] br[168] wl[252] vdd gnd cell_6t
Xbit_r253_c168 bl[168] br[168] wl[253] vdd gnd cell_6t
Xbit_r254_c168 bl[168] br[168] wl[254] vdd gnd cell_6t
Xbit_r255_c168 bl[168] br[168] wl[255] vdd gnd cell_6t
Xbit_r0_c169 bl[169] br[169] wl[0] vdd gnd cell_6t
Xbit_r1_c169 bl[169] br[169] wl[1] vdd gnd cell_6t
Xbit_r2_c169 bl[169] br[169] wl[2] vdd gnd cell_6t
Xbit_r3_c169 bl[169] br[169] wl[3] vdd gnd cell_6t
Xbit_r4_c169 bl[169] br[169] wl[4] vdd gnd cell_6t
Xbit_r5_c169 bl[169] br[169] wl[5] vdd gnd cell_6t
Xbit_r6_c169 bl[169] br[169] wl[6] vdd gnd cell_6t
Xbit_r7_c169 bl[169] br[169] wl[7] vdd gnd cell_6t
Xbit_r8_c169 bl[169] br[169] wl[8] vdd gnd cell_6t
Xbit_r9_c169 bl[169] br[169] wl[9] vdd gnd cell_6t
Xbit_r10_c169 bl[169] br[169] wl[10] vdd gnd cell_6t
Xbit_r11_c169 bl[169] br[169] wl[11] vdd gnd cell_6t
Xbit_r12_c169 bl[169] br[169] wl[12] vdd gnd cell_6t
Xbit_r13_c169 bl[169] br[169] wl[13] vdd gnd cell_6t
Xbit_r14_c169 bl[169] br[169] wl[14] vdd gnd cell_6t
Xbit_r15_c169 bl[169] br[169] wl[15] vdd gnd cell_6t
Xbit_r16_c169 bl[169] br[169] wl[16] vdd gnd cell_6t
Xbit_r17_c169 bl[169] br[169] wl[17] vdd gnd cell_6t
Xbit_r18_c169 bl[169] br[169] wl[18] vdd gnd cell_6t
Xbit_r19_c169 bl[169] br[169] wl[19] vdd gnd cell_6t
Xbit_r20_c169 bl[169] br[169] wl[20] vdd gnd cell_6t
Xbit_r21_c169 bl[169] br[169] wl[21] vdd gnd cell_6t
Xbit_r22_c169 bl[169] br[169] wl[22] vdd gnd cell_6t
Xbit_r23_c169 bl[169] br[169] wl[23] vdd gnd cell_6t
Xbit_r24_c169 bl[169] br[169] wl[24] vdd gnd cell_6t
Xbit_r25_c169 bl[169] br[169] wl[25] vdd gnd cell_6t
Xbit_r26_c169 bl[169] br[169] wl[26] vdd gnd cell_6t
Xbit_r27_c169 bl[169] br[169] wl[27] vdd gnd cell_6t
Xbit_r28_c169 bl[169] br[169] wl[28] vdd gnd cell_6t
Xbit_r29_c169 bl[169] br[169] wl[29] vdd gnd cell_6t
Xbit_r30_c169 bl[169] br[169] wl[30] vdd gnd cell_6t
Xbit_r31_c169 bl[169] br[169] wl[31] vdd gnd cell_6t
Xbit_r32_c169 bl[169] br[169] wl[32] vdd gnd cell_6t
Xbit_r33_c169 bl[169] br[169] wl[33] vdd gnd cell_6t
Xbit_r34_c169 bl[169] br[169] wl[34] vdd gnd cell_6t
Xbit_r35_c169 bl[169] br[169] wl[35] vdd gnd cell_6t
Xbit_r36_c169 bl[169] br[169] wl[36] vdd gnd cell_6t
Xbit_r37_c169 bl[169] br[169] wl[37] vdd gnd cell_6t
Xbit_r38_c169 bl[169] br[169] wl[38] vdd gnd cell_6t
Xbit_r39_c169 bl[169] br[169] wl[39] vdd gnd cell_6t
Xbit_r40_c169 bl[169] br[169] wl[40] vdd gnd cell_6t
Xbit_r41_c169 bl[169] br[169] wl[41] vdd gnd cell_6t
Xbit_r42_c169 bl[169] br[169] wl[42] vdd gnd cell_6t
Xbit_r43_c169 bl[169] br[169] wl[43] vdd gnd cell_6t
Xbit_r44_c169 bl[169] br[169] wl[44] vdd gnd cell_6t
Xbit_r45_c169 bl[169] br[169] wl[45] vdd gnd cell_6t
Xbit_r46_c169 bl[169] br[169] wl[46] vdd gnd cell_6t
Xbit_r47_c169 bl[169] br[169] wl[47] vdd gnd cell_6t
Xbit_r48_c169 bl[169] br[169] wl[48] vdd gnd cell_6t
Xbit_r49_c169 bl[169] br[169] wl[49] vdd gnd cell_6t
Xbit_r50_c169 bl[169] br[169] wl[50] vdd gnd cell_6t
Xbit_r51_c169 bl[169] br[169] wl[51] vdd gnd cell_6t
Xbit_r52_c169 bl[169] br[169] wl[52] vdd gnd cell_6t
Xbit_r53_c169 bl[169] br[169] wl[53] vdd gnd cell_6t
Xbit_r54_c169 bl[169] br[169] wl[54] vdd gnd cell_6t
Xbit_r55_c169 bl[169] br[169] wl[55] vdd gnd cell_6t
Xbit_r56_c169 bl[169] br[169] wl[56] vdd gnd cell_6t
Xbit_r57_c169 bl[169] br[169] wl[57] vdd gnd cell_6t
Xbit_r58_c169 bl[169] br[169] wl[58] vdd gnd cell_6t
Xbit_r59_c169 bl[169] br[169] wl[59] vdd gnd cell_6t
Xbit_r60_c169 bl[169] br[169] wl[60] vdd gnd cell_6t
Xbit_r61_c169 bl[169] br[169] wl[61] vdd gnd cell_6t
Xbit_r62_c169 bl[169] br[169] wl[62] vdd gnd cell_6t
Xbit_r63_c169 bl[169] br[169] wl[63] vdd gnd cell_6t
Xbit_r64_c169 bl[169] br[169] wl[64] vdd gnd cell_6t
Xbit_r65_c169 bl[169] br[169] wl[65] vdd gnd cell_6t
Xbit_r66_c169 bl[169] br[169] wl[66] vdd gnd cell_6t
Xbit_r67_c169 bl[169] br[169] wl[67] vdd gnd cell_6t
Xbit_r68_c169 bl[169] br[169] wl[68] vdd gnd cell_6t
Xbit_r69_c169 bl[169] br[169] wl[69] vdd gnd cell_6t
Xbit_r70_c169 bl[169] br[169] wl[70] vdd gnd cell_6t
Xbit_r71_c169 bl[169] br[169] wl[71] vdd gnd cell_6t
Xbit_r72_c169 bl[169] br[169] wl[72] vdd gnd cell_6t
Xbit_r73_c169 bl[169] br[169] wl[73] vdd gnd cell_6t
Xbit_r74_c169 bl[169] br[169] wl[74] vdd gnd cell_6t
Xbit_r75_c169 bl[169] br[169] wl[75] vdd gnd cell_6t
Xbit_r76_c169 bl[169] br[169] wl[76] vdd gnd cell_6t
Xbit_r77_c169 bl[169] br[169] wl[77] vdd gnd cell_6t
Xbit_r78_c169 bl[169] br[169] wl[78] vdd gnd cell_6t
Xbit_r79_c169 bl[169] br[169] wl[79] vdd gnd cell_6t
Xbit_r80_c169 bl[169] br[169] wl[80] vdd gnd cell_6t
Xbit_r81_c169 bl[169] br[169] wl[81] vdd gnd cell_6t
Xbit_r82_c169 bl[169] br[169] wl[82] vdd gnd cell_6t
Xbit_r83_c169 bl[169] br[169] wl[83] vdd gnd cell_6t
Xbit_r84_c169 bl[169] br[169] wl[84] vdd gnd cell_6t
Xbit_r85_c169 bl[169] br[169] wl[85] vdd gnd cell_6t
Xbit_r86_c169 bl[169] br[169] wl[86] vdd gnd cell_6t
Xbit_r87_c169 bl[169] br[169] wl[87] vdd gnd cell_6t
Xbit_r88_c169 bl[169] br[169] wl[88] vdd gnd cell_6t
Xbit_r89_c169 bl[169] br[169] wl[89] vdd gnd cell_6t
Xbit_r90_c169 bl[169] br[169] wl[90] vdd gnd cell_6t
Xbit_r91_c169 bl[169] br[169] wl[91] vdd gnd cell_6t
Xbit_r92_c169 bl[169] br[169] wl[92] vdd gnd cell_6t
Xbit_r93_c169 bl[169] br[169] wl[93] vdd gnd cell_6t
Xbit_r94_c169 bl[169] br[169] wl[94] vdd gnd cell_6t
Xbit_r95_c169 bl[169] br[169] wl[95] vdd gnd cell_6t
Xbit_r96_c169 bl[169] br[169] wl[96] vdd gnd cell_6t
Xbit_r97_c169 bl[169] br[169] wl[97] vdd gnd cell_6t
Xbit_r98_c169 bl[169] br[169] wl[98] vdd gnd cell_6t
Xbit_r99_c169 bl[169] br[169] wl[99] vdd gnd cell_6t
Xbit_r100_c169 bl[169] br[169] wl[100] vdd gnd cell_6t
Xbit_r101_c169 bl[169] br[169] wl[101] vdd gnd cell_6t
Xbit_r102_c169 bl[169] br[169] wl[102] vdd gnd cell_6t
Xbit_r103_c169 bl[169] br[169] wl[103] vdd gnd cell_6t
Xbit_r104_c169 bl[169] br[169] wl[104] vdd gnd cell_6t
Xbit_r105_c169 bl[169] br[169] wl[105] vdd gnd cell_6t
Xbit_r106_c169 bl[169] br[169] wl[106] vdd gnd cell_6t
Xbit_r107_c169 bl[169] br[169] wl[107] vdd gnd cell_6t
Xbit_r108_c169 bl[169] br[169] wl[108] vdd gnd cell_6t
Xbit_r109_c169 bl[169] br[169] wl[109] vdd gnd cell_6t
Xbit_r110_c169 bl[169] br[169] wl[110] vdd gnd cell_6t
Xbit_r111_c169 bl[169] br[169] wl[111] vdd gnd cell_6t
Xbit_r112_c169 bl[169] br[169] wl[112] vdd gnd cell_6t
Xbit_r113_c169 bl[169] br[169] wl[113] vdd gnd cell_6t
Xbit_r114_c169 bl[169] br[169] wl[114] vdd gnd cell_6t
Xbit_r115_c169 bl[169] br[169] wl[115] vdd gnd cell_6t
Xbit_r116_c169 bl[169] br[169] wl[116] vdd gnd cell_6t
Xbit_r117_c169 bl[169] br[169] wl[117] vdd gnd cell_6t
Xbit_r118_c169 bl[169] br[169] wl[118] vdd gnd cell_6t
Xbit_r119_c169 bl[169] br[169] wl[119] vdd gnd cell_6t
Xbit_r120_c169 bl[169] br[169] wl[120] vdd gnd cell_6t
Xbit_r121_c169 bl[169] br[169] wl[121] vdd gnd cell_6t
Xbit_r122_c169 bl[169] br[169] wl[122] vdd gnd cell_6t
Xbit_r123_c169 bl[169] br[169] wl[123] vdd gnd cell_6t
Xbit_r124_c169 bl[169] br[169] wl[124] vdd gnd cell_6t
Xbit_r125_c169 bl[169] br[169] wl[125] vdd gnd cell_6t
Xbit_r126_c169 bl[169] br[169] wl[126] vdd gnd cell_6t
Xbit_r127_c169 bl[169] br[169] wl[127] vdd gnd cell_6t
Xbit_r128_c169 bl[169] br[169] wl[128] vdd gnd cell_6t
Xbit_r129_c169 bl[169] br[169] wl[129] vdd gnd cell_6t
Xbit_r130_c169 bl[169] br[169] wl[130] vdd gnd cell_6t
Xbit_r131_c169 bl[169] br[169] wl[131] vdd gnd cell_6t
Xbit_r132_c169 bl[169] br[169] wl[132] vdd gnd cell_6t
Xbit_r133_c169 bl[169] br[169] wl[133] vdd gnd cell_6t
Xbit_r134_c169 bl[169] br[169] wl[134] vdd gnd cell_6t
Xbit_r135_c169 bl[169] br[169] wl[135] vdd gnd cell_6t
Xbit_r136_c169 bl[169] br[169] wl[136] vdd gnd cell_6t
Xbit_r137_c169 bl[169] br[169] wl[137] vdd gnd cell_6t
Xbit_r138_c169 bl[169] br[169] wl[138] vdd gnd cell_6t
Xbit_r139_c169 bl[169] br[169] wl[139] vdd gnd cell_6t
Xbit_r140_c169 bl[169] br[169] wl[140] vdd gnd cell_6t
Xbit_r141_c169 bl[169] br[169] wl[141] vdd gnd cell_6t
Xbit_r142_c169 bl[169] br[169] wl[142] vdd gnd cell_6t
Xbit_r143_c169 bl[169] br[169] wl[143] vdd gnd cell_6t
Xbit_r144_c169 bl[169] br[169] wl[144] vdd gnd cell_6t
Xbit_r145_c169 bl[169] br[169] wl[145] vdd gnd cell_6t
Xbit_r146_c169 bl[169] br[169] wl[146] vdd gnd cell_6t
Xbit_r147_c169 bl[169] br[169] wl[147] vdd gnd cell_6t
Xbit_r148_c169 bl[169] br[169] wl[148] vdd gnd cell_6t
Xbit_r149_c169 bl[169] br[169] wl[149] vdd gnd cell_6t
Xbit_r150_c169 bl[169] br[169] wl[150] vdd gnd cell_6t
Xbit_r151_c169 bl[169] br[169] wl[151] vdd gnd cell_6t
Xbit_r152_c169 bl[169] br[169] wl[152] vdd gnd cell_6t
Xbit_r153_c169 bl[169] br[169] wl[153] vdd gnd cell_6t
Xbit_r154_c169 bl[169] br[169] wl[154] vdd gnd cell_6t
Xbit_r155_c169 bl[169] br[169] wl[155] vdd gnd cell_6t
Xbit_r156_c169 bl[169] br[169] wl[156] vdd gnd cell_6t
Xbit_r157_c169 bl[169] br[169] wl[157] vdd gnd cell_6t
Xbit_r158_c169 bl[169] br[169] wl[158] vdd gnd cell_6t
Xbit_r159_c169 bl[169] br[169] wl[159] vdd gnd cell_6t
Xbit_r160_c169 bl[169] br[169] wl[160] vdd gnd cell_6t
Xbit_r161_c169 bl[169] br[169] wl[161] vdd gnd cell_6t
Xbit_r162_c169 bl[169] br[169] wl[162] vdd gnd cell_6t
Xbit_r163_c169 bl[169] br[169] wl[163] vdd gnd cell_6t
Xbit_r164_c169 bl[169] br[169] wl[164] vdd gnd cell_6t
Xbit_r165_c169 bl[169] br[169] wl[165] vdd gnd cell_6t
Xbit_r166_c169 bl[169] br[169] wl[166] vdd gnd cell_6t
Xbit_r167_c169 bl[169] br[169] wl[167] vdd gnd cell_6t
Xbit_r168_c169 bl[169] br[169] wl[168] vdd gnd cell_6t
Xbit_r169_c169 bl[169] br[169] wl[169] vdd gnd cell_6t
Xbit_r170_c169 bl[169] br[169] wl[170] vdd gnd cell_6t
Xbit_r171_c169 bl[169] br[169] wl[171] vdd gnd cell_6t
Xbit_r172_c169 bl[169] br[169] wl[172] vdd gnd cell_6t
Xbit_r173_c169 bl[169] br[169] wl[173] vdd gnd cell_6t
Xbit_r174_c169 bl[169] br[169] wl[174] vdd gnd cell_6t
Xbit_r175_c169 bl[169] br[169] wl[175] vdd gnd cell_6t
Xbit_r176_c169 bl[169] br[169] wl[176] vdd gnd cell_6t
Xbit_r177_c169 bl[169] br[169] wl[177] vdd gnd cell_6t
Xbit_r178_c169 bl[169] br[169] wl[178] vdd gnd cell_6t
Xbit_r179_c169 bl[169] br[169] wl[179] vdd gnd cell_6t
Xbit_r180_c169 bl[169] br[169] wl[180] vdd gnd cell_6t
Xbit_r181_c169 bl[169] br[169] wl[181] vdd gnd cell_6t
Xbit_r182_c169 bl[169] br[169] wl[182] vdd gnd cell_6t
Xbit_r183_c169 bl[169] br[169] wl[183] vdd gnd cell_6t
Xbit_r184_c169 bl[169] br[169] wl[184] vdd gnd cell_6t
Xbit_r185_c169 bl[169] br[169] wl[185] vdd gnd cell_6t
Xbit_r186_c169 bl[169] br[169] wl[186] vdd gnd cell_6t
Xbit_r187_c169 bl[169] br[169] wl[187] vdd gnd cell_6t
Xbit_r188_c169 bl[169] br[169] wl[188] vdd gnd cell_6t
Xbit_r189_c169 bl[169] br[169] wl[189] vdd gnd cell_6t
Xbit_r190_c169 bl[169] br[169] wl[190] vdd gnd cell_6t
Xbit_r191_c169 bl[169] br[169] wl[191] vdd gnd cell_6t
Xbit_r192_c169 bl[169] br[169] wl[192] vdd gnd cell_6t
Xbit_r193_c169 bl[169] br[169] wl[193] vdd gnd cell_6t
Xbit_r194_c169 bl[169] br[169] wl[194] vdd gnd cell_6t
Xbit_r195_c169 bl[169] br[169] wl[195] vdd gnd cell_6t
Xbit_r196_c169 bl[169] br[169] wl[196] vdd gnd cell_6t
Xbit_r197_c169 bl[169] br[169] wl[197] vdd gnd cell_6t
Xbit_r198_c169 bl[169] br[169] wl[198] vdd gnd cell_6t
Xbit_r199_c169 bl[169] br[169] wl[199] vdd gnd cell_6t
Xbit_r200_c169 bl[169] br[169] wl[200] vdd gnd cell_6t
Xbit_r201_c169 bl[169] br[169] wl[201] vdd gnd cell_6t
Xbit_r202_c169 bl[169] br[169] wl[202] vdd gnd cell_6t
Xbit_r203_c169 bl[169] br[169] wl[203] vdd gnd cell_6t
Xbit_r204_c169 bl[169] br[169] wl[204] vdd gnd cell_6t
Xbit_r205_c169 bl[169] br[169] wl[205] vdd gnd cell_6t
Xbit_r206_c169 bl[169] br[169] wl[206] vdd gnd cell_6t
Xbit_r207_c169 bl[169] br[169] wl[207] vdd gnd cell_6t
Xbit_r208_c169 bl[169] br[169] wl[208] vdd gnd cell_6t
Xbit_r209_c169 bl[169] br[169] wl[209] vdd gnd cell_6t
Xbit_r210_c169 bl[169] br[169] wl[210] vdd gnd cell_6t
Xbit_r211_c169 bl[169] br[169] wl[211] vdd gnd cell_6t
Xbit_r212_c169 bl[169] br[169] wl[212] vdd gnd cell_6t
Xbit_r213_c169 bl[169] br[169] wl[213] vdd gnd cell_6t
Xbit_r214_c169 bl[169] br[169] wl[214] vdd gnd cell_6t
Xbit_r215_c169 bl[169] br[169] wl[215] vdd gnd cell_6t
Xbit_r216_c169 bl[169] br[169] wl[216] vdd gnd cell_6t
Xbit_r217_c169 bl[169] br[169] wl[217] vdd gnd cell_6t
Xbit_r218_c169 bl[169] br[169] wl[218] vdd gnd cell_6t
Xbit_r219_c169 bl[169] br[169] wl[219] vdd gnd cell_6t
Xbit_r220_c169 bl[169] br[169] wl[220] vdd gnd cell_6t
Xbit_r221_c169 bl[169] br[169] wl[221] vdd gnd cell_6t
Xbit_r222_c169 bl[169] br[169] wl[222] vdd gnd cell_6t
Xbit_r223_c169 bl[169] br[169] wl[223] vdd gnd cell_6t
Xbit_r224_c169 bl[169] br[169] wl[224] vdd gnd cell_6t
Xbit_r225_c169 bl[169] br[169] wl[225] vdd gnd cell_6t
Xbit_r226_c169 bl[169] br[169] wl[226] vdd gnd cell_6t
Xbit_r227_c169 bl[169] br[169] wl[227] vdd gnd cell_6t
Xbit_r228_c169 bl[169] br[169] wl[228] vdd gnd cell_6t
Xbit_r229_c169 bl[169] br[169] wl[229] vdd gnd cell_6t
Xbit_r230_c169 bl[169] br[169] wl[230] vdd gnd cell_6t
Xbit_r231_c169 bl[169] br[169] wl[231] vdd gnd cell_6t
Xbit_r232_c169 bl[169] br[169] wl[232] vdd gnd cell_6t
Xbit_r233_c169 bl[169] br[169] wl[233] vdd gnd cell_6t
Xbit_r234_c169 bl[169] br[169] wl[234] vdd gnd cell_6t
Xbit_r235_c169 bl[169] br[169] wl[235] vdd gnd cell_6t
Xbit_r236_c169 bl[169] br[169] wl[236] vdd gnd cell_6t
Xbit_r237_c169 bl[169] br[169] wl[237] vdd gnd cell_6t
Xbit_r238_c169 bl[169] br[169] wl[238] vdd gnd cell_6t
Xbit_r239_c169 bl[169] br[169] wl[239] vdd gnd cell_6t
Xbit_r240_c169 bl[169] br[169] wl[240] vdd gnd cell_6t
Xbit_r241_c169 bl[169] br[169] wl[241] vdd gnd cell_6t
Xbit_r242_c169 bl[169] br[169] wl[242] vdd gnd cell_6t
Xbit_r243_c169 bl[169] br[169] wl[243] vdd gnd cell_6t
Xbit_r244_c169 bl[169] br[169] wl[244] vdd gnd cell_6t
Xbit_r245_c169 bl[169] br[169] wl[245] vdd gnd cell_6t
Xbit_r246_c169 bl[169] br[169] wl[246] vdd gnd cell_6t
Xbit_r247_c169 bl[169] br[169] wl[247] vdd gnd cell_6t
Xbit_r248_c169 bl[169] br[169] wl[248] vdd gnd cell_6t
Xbit_r249_c169 bl[169] br[169] wl[249] vdd gnd cell_6t
Xbit_r250_c169 bl[169] br[169] wl[250] vdd gnd cell_6t
Xbit_r251_c169 bl[169] br[169] wl[251] vdd gnd cell_6t
Xbit_r252_c169 bl[169] br[169] wl[252] vdd gnd cell_6t
Xbit_r253_c169 bl[169] br[169] wl[253] vdd gnd cell_6t
Xbit_r254_c169 bl[169] br[169] wl[254] vdd gnd cell_6t
Xbit_r255_c169 bl[169] br[169] wl[255] vdd gnd cell_6t
Xbit_r0_c170 bl[170] br[170] wl[0] vdd gnd cell_6t
Xbit_r1_c170 bl[170] br[170] wl[1] vdd gnd cell_6t
Xbit_r2_c170 bl[170] br[170] wl[2] vdd gnd cell_6t
Xbit_r3_c170 bl[170] br[170] wl[3] vdd gnd cell_6t
Xbit_r4_c170 bl[170] br[170] wl[4] vdd gnd cell_6t
Xbit_r5_c170 bl[170] br[170] wl[5] vdd gnd cell_6t
Xbit_r6_c170 bl[170] br[170] wl[6] vdd gnd cell_6t
Xbit_r7_c170 bl[170] br[170] wl[7] vdd gnd cell_6t
Xbit_r8_c170 bl[170] br[170] wl[8] vdd gnd cell_6t
Xbit_r9_c170 bl[170] br[170] wl[9] vdd gnd cell_6t
Xbit_r10_c170 bl[170] br[170] wl[10] vdd gnd cell_6t
Xbit_r11_c170 bl[170] br[170] wl[11] vdd gnd cell_6t
Xbit_r12_c170 bl[170] br[170] wl[12] vdd gnd cell_6t
Xbit_r13_c170 bl[170] br[170] wl[13] vdd gnd cell_6t
Xbit_r14_c170 bl[170] br[170] wl[14] vdd gnd cell_6t
Xbit_r15_c170 bl[170] br[170] wl[15] vdd gnd cell_6t
Xbit_r16_c170 bl[170] br[170] wl[16] vdd gnd cell_6t
Xbit_r17_c170 bl[170] br[170] wl[17] vdd gnd cell_6t
Xbit_r18_c170 bl[170] br[170] wl[18] vdd gnd cell_6t
Xbit_r19_c170 bl[170] br[170] wl[19] vdd gnd cell_6t
Xbit_r20_c170 bl[170] br[170] wl[20] vdd gnd cell_6t
Xbit_r21_c170 bl[170] br[170] wl[21] vdd gnd cell_6t
Xbit_r22_c170 bl[170] br[170] wl[22] vdd gnd cell_6t
Xbit_r23_c170 bl[170] br[170] wl[23] vdd gnd cell_6t
Xbit_r24_c170 bl[170] br[170] wl[24] vdd gnd cell_6t
Xbit_r25_c170 bl[170] br[170] wl[25] vdd gnd cell_6t
Xbit_r26_c170 bl[170] br[170] wl[26] vdd gnd cell_6t
Xbit_r27_c170 bl[170] br[170] wl[27] vdd gnd cell_6t
Xbit_r28_c170 bl[170] br[170] wl[28] vdd gnd cell_6t
Xbit_r29_c170 bl[170] br[170] wl[29] vdd gnd cell_6t
Xbit_r30_c170 bl[170] br[170] wl[30] vdd gnd cell_6t
Xbit_r31_c170 bl[170] br[170] wl[31] vdd gnd cell_6t
Xbit_r32_c170 bl[170] br[170] wl[32] vdd gnd cell_6t
Xbit_r33_c170 bl[170] br[170] wl[33] vdd gnd cell_6t
Xbit_r34_c170 bl[170] br[170] wl[34] vdd gnd cell_6t
Xbit_r35_c170 bl[170] br[170] wl[35] vdd gnd cell_6t
Xbit_r36_c170 bl[170] br[170] wl[36] vdd gnd cell_6t
Xbit_r37_c170 bl[170] br[170] wl[37] vdd gnd cell_6t
Xbit_r38_c170 bl[170] br[170] wl[38] vdd gnd cell_6t
Xbit_r39_c170 bl[170] br[170] wl[39] vdd gnd cell_6t
Xbit_r40_c170 bl[170] br[170] wl[40] vdd gnd cell_6t
Xbit_r41_c170 bl[170] br[170] wl[41] vdd gnd cell_6t
Xbit_r42_c170 bl[170] br[170] wl[42] vdd gnd cell_6t
Xbit_r43_c170 bl[170] br[170] wl[43] vdd gnd cell_6t
Xbit_r44_c170 bl[170] br[170] wl[44] vdd gnd cell_6t
Xbit_r45_c170 bl[170] br[170] wl[45] vdd gnd cell_6t
Xbit_r46_c170 bl[170] br[170] wl[46] vdd gnd cell_6t
Xbit_r47_c170 bl[170] br[170] wl[47] vdd gnd cell_6t
Xbit_r48_c170 bl[170] br[170] wl[48] vdd gnd cell_6t
Xbit_r49_c170 bl[170] br[170] wl[49] vdd gnd cell_6t
Xbit_r50_c170 bl[170] br[170] wl[50] vdd gnd cell_6t
Xbit_r51_c170 bl[170] br[170] wl[51] vdd gnd cell_6t
Xbit_r52_c170 bl[170] br[170] wl[52] vdd gnd cell_6t
Xbit_r53_c170 bl[170] br[170] wl[53] vdd gnd cell_6t
Xbit_r54_c170 bl[170] br[170] wl[54] vdd gnd cell_6t
Xbit_r55_c170 bl[170] br[170] wl[55] vdd gnd cell_6t
Xbit_r56_c170 bl[170] br[170] wl[56] vdd gnd cell_6t
Xbit_r57_c170 bl[170] br[170] wl[57] vdd gnd cell_6t
Xbit_r58_c170 bl[170] br[170] wl[58] vdd gnd cell_6t
Xbit_r59_c170 bl[170] br[170] wl[59] vdd gnd cell_6t
Xbit_r60_c170 bl[170] br[170] wl[60] vdd gnd cell_6t
Xbit_r61_c170 bl[170] br[170] wl[61] vdd gnd cell_6t
Xbit_r62_c170 bl[170] br[170] wl[62] vdd gnd cell_6t
Xbit_r63_c170 bl[170] br[170] wl[63] vdd gnd cell_6t
Xbit_r64_c170 bl[170] br[170] wl[64] vdd gnd cell_6t
Xbit_r65_c170 bl[170] br[170] wl[65] vdd gnd cell_6t
Xbit_r66_c170 bl[170] br[170] wl[66] vdd gnd cell_6t
Xbit_r67_c170 bl[170] br[170] wl[67] vdd gnd cell_6t
Xbit_r68_c170 bl[170] br[170] wl[68] vdd gnd cell_6t
Xbit_r69_c170 bl[170] br[170] wl[69] vdd gnd cell_6t
Xbit_r70_c170 bl[170] br[170] wl[70] vdd gnd cell_6t
Xbit_r71_c170 bl[170] br[170] wl[71] vdd gnd cell_6t
Xbit_r72_c170 bl[170] br[170] wl[72] vdd gnd cell_6t
Xbit_r73_c170 bl[170] br[170] wl[73] vdd gnd cell_6t
Xbit_r74_c170 bl[170] br[170] wl[74] vdd gnd cell_6t
Xbit_r75_c170 bl[170] br[170] wl[75] vdd gnd cell_6t
Xbit_r76_c170 bl[170] br[170] wl[76] vdd gnd cell_6t
Xbit_r77_c170 bl[170] br[170] wl[77] vdd gnd cell_6t
Xbit_r78_c170 bl[170] br[170] wl[78] vdd gnd cell_6t
Xbit_r79_c170 bl[170] br[170] wl[79] vdd gnd cell_6t
Xbit_r80_c170 bl[170] br[170] wl[80] vdd gnd cell_6t
Xbit_r81_c170 bl[170] br[170] wl[81] vdd gnd cell_6t
Xbit_r82_c170 bl[170] br[170] wl[82] vdd gnd cell_6t
Xbit_r83_c170 bl[170] br[170] wl[83] vdd gnd cell_6t
Xbit_r84_c170 bl[170] br[170] wl[84] vdd gnd cell_6t
Xbit_r85_c170 bl[170] br[170] wl[85] vdd gnd cell_6t
Xbit_r86_c170 bl[170] br[170] wl[86] vdd gnd cell_6t
Xbit_r87_c170 bl[170] br[170] wl[87] vdd gnd cell_6t
Xbit_r88_c170 bl[170] br[170] wl[88] vdd gnd cell_6t
Xbit_r89_c170 bl[170] br[170] wl[89] vdd gnd cell_6t
Xbit_r90_c170 bl[170] br[170] wl[90] vdd gnd cell_6t
Xbit_r91_c170 bl[170] br[170] wl[91] vdd gnd cell_6t
Xbit_r92_c170 bl[170] br[170] wl[92] vdd gnd cell_6t
Xbit_r93_c170 bl[170] br[170] wl[93] vdd gnd cell_6t
Xbit_r94_c170 bl[170] br[170] wl[94] vdd gnd cell_6t
Xbit_r95_c170 bl[170] br[170] wl[95] vdd gnd cell_6t
Xbit_r96_c170 bl[170] br[170] wl[96] vdd gnd cell_6t
Xbit_r97_c170 bl[170] br[170] wl[97] vdd gnd cell_6t
Xbit_r98_c170 bl[170] br[170] wl[98] vdd gnd cell_6t
Xbit_r99_c170 bl[170] br[170] wl[99] vdd gnd cell_6t
Xbit_r100_c170 bl[170] br[170] wl[100] vdd gnd cell_6t
Xbit_r101_c170 bl[170] br[170] wl[101] vdd gnd cell_6t
Xbit_r102_c170 bl[170] br[170] wl[102] vdd gnd cell_6t
Xbit_r103_c170 bl[170] br[170] wl[103] vdd gnd cell_6t
Xbit_r104_c170 bl[170] br[170] wl[104] vdd gnd cell_6t
Xbit_r105_c170 bl[170] br[170] wl[105] vdd gnd cell_6t
Xbit_r106_c170 bl[170] br[170] wl[106] vdd gnd cell_6t
Xbit_r107_c170 bl[170] br[170] wl[107] vdd gnd cell_6t
Xbit_r108_c170 bl[170] br[170] wl[108] vdd gnd cell_6t
Xbit_r109_c170 bl[170] br[170] wl[109] vdd gnd cell_6t
Xbit_r110_c170 bl[170] br[170] wl[110] vdd gnd cell_6t
Xbit_r111_c170 bl[170] br[170] wl[111] vdd gnd cell_6t
Xbit_r112_c170 bl[170] br[170] wl[112] vdd gnd cell_6t
Xbit_r113_c170 bl[170] br[170] wl[113] vdd gnd cell_6t
Xbit_r114_c170 bl[170] br[170] wl[114] vdd gnd cell_6t
Xbit_r115_c170 bl[170] br[170] wl[115] vdd gnd cell_6t
Xbit_r116_c170 bl[170] br[170] wl[116] vdd gnd cell_6t
Xbit_r117_c170 bl[170] br[170] wl[117] vdd gnd cell_6t
Xbit_r118_c170 bl[170] br[170] wl[118] vdd gnd cell_6t
Xbit_r119_c170 bl[170] br[170] wl[119] vdd gnd cell_6t
Xbit_r120_c170 bl[170] br[170] wl[120] vdd gnd cell_6t
Xbit_r121_c170 bl[170] br[170] wl[121] vdd gnd cell_6t
Xbit_r122_c170 bl[170] br[170] wl[122] vdd gnd cell_6t
Xbit_r123_c170 bl[170] br[170] wl[123] vdd gnd cell_6t
Xbit_r124_c170 bl[170] br[170] wl[124] vdd gnd cell_6t
Xbit_r125_c170 bl[170] br[170] wl[125] vdd gnd cell_6t
Xbit_r126_c170 bl[170] br[170] wl[126] vdd gnd cell_6t
Xbit_r127_c170 bl[170] br[170] wl[127] vdd gnd cell_6t
Xbit_r128_c170 bl[170] br[170] wl[128] vdd gnd cell_6t
Xbit_r129_c170 bl[170] br[170] wl[129] vdd gnd cell_6t
Xbit_r130_c170 bl[170] br[170] wl[130] vdd gnd cell_6t
Xbit_r131_c170 bl[170] br[170] wl[131] vdd gnd cell_6t
Xbit_r132_c170 bl[170] br[170] wl[132] vdd gnd cell_6t
Xbit_r133_c170 bl[170] br[170] wl[133] vdd gnd cell_6t
Xbit_r134_c170 bl[170] br[170] wl[134] vdd gnd cell_6t
Xbit_r135_c170 bl[170] br[170] wl[135] vdd gnd cell_6t
Xbit_r136_c170 bl[170] br[170] wl[136] vdd gnd cell_6t
Xbit_r137_c170 bl[170] br[170] wl[137] vdd gnd cell_6t
Xbit_r138_c170 bl[170] br[170] wl[138] vdd gnd cell_6t
Xbit_r139_c170 bl[170] br[170] wl[139] vdd gnd cell_6t
Xbit_r140_c170 bl[170] br[170] wl[140] vdd gnd cell_6t
Xbit_r141_c170 bl[170] br[170] wl[141] vdd gnd cell_6t
Xbit_r142_c170 bl[170] br[170] wl[142] vdd gnd cell_6t
Xbit_r143_c170 bl[170] br[170] wl[143] vdd gnd cell_6t
Xbit_r144_c170 bl[170] br[170] wl[144] vdd gnd cell_6t
Xbit_r145_c170 bl[170] br[170] wl[145] vdd gnd cell_6t
Xbit_r146_c170 bl[170] br[170] wl[146] vdd gnd cell_6t
Xbit_r147_c170 bl[170] br[170] wl[147] vdd gnd cell_6t
Xbit_r148_c170 bl[170] br[170] wl[148] vdd gnd cell_6t
Xbit_r149_c170 bl[170] br[170] wl[149] vdd gnd cell_6t
Xbit_r150_c170 bl[170] br[170] wl[150] vdd gnd cell_6t
Xbit_r151_c170 bl[170] br[170] wl[151] vdd gnd cell_6t
Xbit_r152_c170 bl[170] br[170] wl[152] vdd gnd cell_6t
Xbit_r153_c170 bl[170] br[170] wl[153] vdd gnd cell_6t
Xbit_r154_c170 bl[170] br[170] wl[154] vdd gnd cell_6t
Xbit_r155_c170 bl[170] br[170] wl[155] vdd gnd cell_6t
Xbit_r156_c170 bl[170] br[170] wl[156] vdd gnd cell_6t
Xbit_r157_c170 bl[170] br[170] wl[157] vdd gnd cell_6t
Xbit_r158_c170 bl[170] br[170] wl[158] vdd gnd cell_6t
Xbit_r159_c170 bl[170] br[170] wl[159] vdd gnd cell_6t
Xbit_r160_c170 bl[170] br[170] wl[160] vdd gnd cell_6t
Xbit_r161_c170 bl[170] br[170] wl[161] vdd gnd cell_6t
Xbit_r162_c170 bl[170] br[170] wl[162] vdd gnd cell_6t
Xbit_r163_c170 bl[170] br[170] wl[163] vdd gnd cell_6t
Xbit_r164_c170 bl[170] br[170] wl[164] vdd gnd cell_6t
Xbit_r165_c170 bl[170] br[170] wl[165] vdd gnd cell_6t
Xbit_r166_c170 bl[170] br[170] wl[166] vdd gnd cell_6t
Xbit_r167_c170 bl[170] br[170] wl[167] vdd gnd cell_6t
Xbit_r168_c170 bl[170] br[170] wl[168] vdd gnd cell_6t
Xbit_r169_c170 bl[170] br[170] wl[169] vdd gnd cell_6t
Xbit_r170_c170 bl[170] br[170] wl[170] vdd gnd cell_6t
Xbit_r171_c170 bl[170] br[170] wl[171] vdd gnd cell_6t
Xbit_r172_c170 bl[170] br[170] wl[172] vdd gnd cell_6t
Xbit_r173_c170 bl[170] br[170] wl[173] vdd gnd cell_6t
Xbit_r174_c170 bl[170] br[170] wl[174] vdd gnd cell_6t
Xbit_r175_c170 bl[170] br[170] wl[175] vdd gnd cell_6t
Xbit_r176_c170 bl[170] br[170] wl[176] vdd gnd cell_6t
Xbit_r177_c170 bl[170] br[170] wl[177] vdd gnd cell_6t
Xbit_r178_c170 bl[170] br[170] wl[178] vdd gnd cell_6t
Xbit_r179_c170 bl[170] br[170] wl[179] vdd gnd cell_6t
Xbit_r180_c170 bl[170] br[170] wl[180] vdd gnd cell_6t
Xbit_r181_c170 bl[170] br[170] wl[181] vdd gnd cell_6t
Xbit_r182_c170 bl[170] br[170] wl[182] vdd gnd cell_6t
Xbit_r183_c170 bl[170] br[170] wl[183] vdd gnd cell_6t
Xbit_r184_c170 bl[170] br[170] wl[184] vdd gnd cell_6t
Xbit_r185_c170 bl[170] br[170] wl[185] vdd gnd cell_6t
Xbit_r186_c170 bl[170] br[170] wl[186] vdd gnd cell_6t
Xbit_r187_c170 bl[170] br[170] wl[187] vdd gnd cell_6t
Xbit_r188_c170 bl[170] br[170] wl[188] vdd gnd cell_6t
Xbit_r189_c170 bl[170] br[170] wl[189] vdd gnd cell_6t
Xbit_r190_c170 bl[170] br[170] wl[190] vdd gnd cell_6t
Xbit_r191_c170 bl[170] br[170] wl[191] vdd gnd cell_6t
Xbit_r192_c170 bl[170] br[170] wl[192] vdd gnd cell_6t
Xbit_r193_c170 bl[170] br[170] wl[193] vdd gnd cell_6t
Xbit_r194_c170 bl[170] br[170] wl[194] vdd gnd cell_6t
Xbit_r195_c170 bl[170] br[170] wl[195] vdd gnd cell_6t
Xbit_r196_c170 bl[170] br[170] wl[196] vdd gnd cell_6t
Xbit_r197_c170 bl[170] br[170] wl[197] vdd gnd cell_6t
Xbit_r198_c170 bl[170] br[170] wl[198] vdd gnd cell_6t
Xbit_r199_c170 bl[170] br[170] wl[199] vdd gnd cell_6t
Xbit_r200_c170 bl[170] br[170] wl[200] vdd gnd cell_6t
Xbit_r201_c170 bl[170] br[170] wl[201] vdd gnd cell_6t
Xbit_r202_c170 bl[170] br[170] wl[202] vdd gnd cell_6t
Xbit_r203_c170 bl[170] br[170] wl[203] vdd gnd cell_6t
Xbit_r204_c170 bl[170] br[170] wl[204] vdd gnd cell_6t
Xbit_r205_c170 bl[170] br[170] wl[205] vdd gnd cell_6t
Xbit_r206_c170 bl[170] br[170] wl[206] vdd gnd cell_6t
Xbit_r207_c170 bl[170] br[170] wl[207] vdd gnd cell_6t
Xbit_r208_c170 bl[170] br[170] wl[208] vdd gnd cell_6t
Xbit_r209_c170 bl[170] br[170] wl[209] vdd gnd cell_6t
Xbit_r210_c170 bl[170] br[170] wl[210] vdd gnd cell_6t
Xbit_r211_c170 bl[170] br[170] wl[211] vdd gnd cell_6t
Xbit_r212_c170 bl[170] br[170] wl[212] vdd gnd cell_6t
Xbit_r213_c170 bl[170] br[170] wl[213] vdd gnd cell_6t
Xbit_r214_c170 bl[170] br[170] wl[214] vdd gnd cell_6t
Xbit_r215_c170 bl[170] br[170] wl[215] vdd gnd cell_6t
Xbit_r216_c170 bl[170] br[170] wl[216] vdd gnd cell_6t
Xbit_r217_c170 bl[170] br[170] wl[217] vdd gnd cell_6t
Xbit_r218_c170 bl[170] br[170] wl[218] vdd gnd cell_6t
Xbit_r219_c170 bl[170] br[170] wl[219] vdd gnd cell_6t
Xbit_r220_c170 bl[170] br[170] wl[220] vdd gnd cell_6t
Xbit_r221_c170 bl[170] br[170] wl[221] vdd gnd cell_6t
Xbit_r222_c170 bl[170] br[170] wl[222] vdd gnd cell_6t
Xbit_r223_c170 bl[170] br[170] wl[223] vdd gnd cell_6t
Xbit_r224_c170 bl[170] br[170] wl[224] vdd gnd cell_6t
Xbit_r225_c170 bl[170] br[170] wl[225] vdd gnd cell_6t
Xbit_r226_c170 bl[170] br[170] wl[226] vdd gnd cell_6t
Xbit_r227_c170 bl[170] br[170] wl[227] vdd gnd cell_6t
Xbit_r228_c170 bl[170] br[170] wl[228] vdd gnd cell_6t
Xbit_r229_c170 bl[170] br[170] wl[229] vdd gnd cell_6t
Xbit_r230_c170 bl[170] br[170] wl[230] vdd gnd cell_6t
Xbit_r231_c170 bl[170] br[170] wl[231] vdd gnd cell_6t
Xbit_r232_c170 bl[170] br[170] wl[232] vdd gnd cell_6t
Xbit_r233_c170 bl[170] br[170] wl[233] vdd gnd cell_6t
Xbit_r234_c170 bl[170] br[170] wl[234] vdd gnd cell_6t
Xbit_r235_c170 bl[170] br[170] wl[235] vdd gnd cell_6t
Xbit_r236_c170 bl[170] br[170] wl[236] vdd gnd cell_6t
Xbit_r237_c170 bl[170] br[170] wl[237] vdd gnd cell_6t
Xbit_r238_c170 bl[170] br[170] wl[238] vdd gnd cell_6t
Xbit_r239_c170 bl[170] br[170] wl[239] vdd gnd cell_6t
Xbit_r240_c170 bl[170] br[170] wl[240] vdd gnd cell_6t
Xbit_r241_c170 bl[170] br[170] wl[241] vdd gnd cell_6t
Xbit_r242_c170 bl[170] br[170] wl[242] vdd gnd cell_6t
Xbit_r243_c170 bl[170] br[170] wl[243] vdd gnd cell_6t
Xbit_r244_c170 bl[170] br[170] wl[244] vdd gnd cell_6t
Xbit_r245_c170 bl[170] br[170] wl[245] vdd gnd cell_6t
Xbit_r246_c170 bl[170] br[170] wl[246] vdd gnd cell_6t
Xbit_r247_c170 bl[170] br[170] wl[247] vdd gnd cell_6t
Xbit_r248_c170 bl[170] br[170] wl[248] vdd gnd cell_6t
Xbit_r249_c170 bl[170] br[170] wl[249] vdd gnd cell_6t
Xbit_r250_c170 bl[170] br[170] wl[250] vdd gnd cell_6t
Xbit_r251_c170 bl[170] br[170] wl[251] vdd gnd cell_6t
Xbit_r252_c170 bl[170] br[170] wl[252] vdd gnd cell_6t
Xbit_r253_c170 bl[170] br[170] wl[253] vdd gnd cell_6t
Xbit_r254_c170 bl[170] br[170] wl[254] vdd gnd cell_6t
Xbit_r255_c170 bl[170] br[170] wl[255] vdd gnd cell_6t
Xbit_r0_c171 bl[171] br[171] wl[0] vdd gnd cell_6t
Xbit_r1_c171 bl[171] br[171] wl[1] vdd gnd cell_6t
Xbit_r2_c171 bl[171] br[171] wl[2] vdd gnd cell_6t
Xbit_r3_c171 bl[171] br[171] wl[3] vdd gnd cell_6t
Xbit_r4_c171 bl[171] br[171] wl[4] vdd gnd cell_6t
Xbit_r5_c171 bl[171] br[171] wl[5] vdd gnd cell_6t
Xbit_r6_c171 bl[171] br[171] wl[6] vdd gnd cell_6t
Xbit_r7_c171 bl[171] br[171] wl[7] vdd gnd cell_6t
Xbit_r8_c171 bl[171] br[171] wl[8] vdd gnd cell_6t
Xbit_r9_c171 bl[171] br[171] wl[9] vdd gnd cell_6t
Xbit_r10_c171 bl[171] br[171] wl[10] vdd gnd cell_6t
Xbit_r11_c171 bl[171] br[171] wl[11] vdd gnd cell_6t
Xbit_r12_c171 bl[171] br[171] wl[12] vdd gnd cell_6t
Xbit_r13_c171 bl[171] br[171] wl[13] vdd gnd cell_6t
Xbit_r14_c171 bl[171] br[171] wl[14] vdd gnd cell_6t
Xbit_r15_c171 bl[171] br[171] wl[15] vdd gnd cell_6t
Xbit_r16_c171 bl[171] br[171] wl[16] vdd gnd cell_6t
Xbit_r17_c171 bl[171] br[171] wl[17] vdd gnd cell_6t
Xbit_r18_c171 bl[171] br[171] wl[18] vdd gnd cell_6t
Xbit_r19_c171 bl[171] br[171] wl[19] vdd gnd cell_6t
Xbit_r20_c171 bl[171] br[171] wl[20] vdd gnd cell_6t
Xbit_r21_c171 bl[171] br[171] wl[21] vdd gnd cell_6t
Xbit_r22_c171 bl[171] br[171] wl[22] vdd gnd cell_6t
Xbit_r23_c171 bl[171] br[171] wl[23] vdd gnd cell_6t
Xbit_r24_c171 bl[171] br[171] wl[24] vdd gnd cell_6t
Xbit_r25_c171 bl[171] br[171] wl[25] vdd gnd cell_6t
Xbit_r26_c171 bl[171] br[171] wl[26] vdd gnd cell_6t
Xbit_r27_c171 bl[171] br[171] wl[27] vdd gnd cell_6t
Xbit_r28_c171 bl[171] br[171] wl[28] vdd gnd cell_6t
Xbit_r29_c171 bl[171] br[171] wl[29] vdd gnd cell_6t
Xbit_r30_c171 bl[171] br[171] wl[30] vdd gnd cell_6t
Xbit_r31_c171 bl[171] br[171] wl[31] vdd gnd cell_6t
Xbit_r32_c171 bl[171] br[171] wl[32] vdd gnd cell_6t
Xbit_r33_c171 bl[171] br[171] wl[33] vdd gnd cell_6t
Xbit_r34_c171 bl[171] br[171] wl[34] vdd gnd cell_6t
Xbit_r35_c171 bl[171] br[171] wl[35] vdd gnd cell_6t
Xbit_r36_c171 bl[171] br[171] wl[36] vdd gnd cell_6t
Xbit_r37_c171 bl[171] br[171] wl[37] vdd gnd cell_6t
Xbit_r38_c171 bl[171] br[171] wl[38] vdd gnd cell_6t
Xbit_r39_c171 bl[171] br[171] wl[39] vdd gnd cell_6t
Xbit_r40_c171 bl[171] br[171] wl[40] vdd gnd cell_6t
Xbit_r41_c171 bl[171] br[171] wl[41] vdd gnd cell_6t
Xbit_r42_c171 bl[171] br[171] wl[42] vdd gnd cell_6t
Xbit_r43_c171 bl[171] br[171] wl[43] vdd gnd cell_6t
Xbit_r44_c171 bl[171] br[171] wl[44] vdd gnd cell_6t
Xbit_r45_c171 bl[171] br[171] wl[45] vdd gnd cell_6t
Xbit_r46_c171 bl[171] br[171] wl[46] vdd gnd cell_6t
Xbit_r47_c171 bl[171] br[171] wl[47] vdd gnd cell_6t
Xbit_r48_c171 bl[171] br[171] wl[48] vdd gnd cell_6t
Xbit_r49_c171 bl[171] br[171] wl[49] vdd gnd cell_6t
Xbit_r50_c171 bl[171] br[171] wl[50] vdd gnd cell_6t
Xbit_r51_c171 bl[171] br[171] wl[51] vdd gnd cell_6t
Xbit_r52_c171 bl[171] br[171] wl[52] vdd gnd cell_6t
Xbit_r53_c171 bl[171] br[171] wl[53] vdd gnd cell_6t
Xbit_r54_c171 bl[171] br[171] wl[54] vdd gnd cell_6t
Xbit_r55_c171 bl[171] br[171] wl[55] vdd gnd cell_6t
Xbit_r56_c171 bl[171] br[171] wl[56] vdd gnd cell_6t
Xbit_r57_c171 bl[171] br[171] wl[57] vdd gnd cell_6t
Xbit_r58_c171 bl[171] br[171] wl[58] vdd gnd cell_6t
Xbit_r59_c171 bl[171] br[171] wl[59] vdd gnd cell_6t
Xbit_r60_c171 bl[171] br[171] wl[60] vdd gnd cell_6t
Xbit_r61_c171 bl[171] br[171] wl[61] vdd gnd cell_6t
Xbit_r62_c171 bl[171] br[171] wl[62] vdd gnd cell_6t
Xbit_r63_c171 bl[171] br[171] wl[63] vdd gnd cell_6t
Xbit_r64_c171 bl[171] br[171] wl[64] vdd gnd cell_6t
Xbit_r65_c171 bl[171] br[171] wl[65] vdd gnd cell_6t
Xbit_r66_c171 bl[171] br[171] wl[66] vdd gnd cell_6t
Xbit_r67_c171 bl[171] br[171] wl[67] vdd gnd cell_6t
Xbit_r68_c171 bl[171] br[171] wl[68] vdd gnd cell_6t
Xbit_r69_c171 bl[171] br[171] wl[69] vdd gnd cell_6t
Xbit_r70_c171 bl[171] br[171] wl[70] vdd gnd cell_6t
Xbit_r71_c171 bl[171] br[171] wl[71] vdd gnd cell_6t
Xbit_r72_c171 bl[171] br[171] wl[72] vdd gnd cell_6t
Xbit_r73_c171 bl[171] br[171] wl[73] vdd gnd cell_6t
Xbit_r74_c171 bl[171] br[171] wl[74] vdd gnd cell_6t
Xbit_r75_c171 bl[171] br[171] wl[75] vdd gnd cell_6t
Xbit_r76_c171 bl[171] br[171] wl[76] vdd gnd cell_6t
Xbit_r77_c171 bl[171] br[171] wl[77] vdd gnd cell_6t
Xbit_r78_c171 bl[171] br[171] wl[78] vdd gnd cell_6t
Xbit_r79_c171 bl[171] br[171] wl[79] vdd gnd cell_6t
Xbit_r80_c171 bl[171] br[171] wl[80] vdd gnd cell_6t
Xbit_r81_c171 bl[171] br[171] wl[81] vdd gnd cell_6t
Xbit_r82_c171 bl[171] br[171] wl[82] vdd gnd cell_6t
Xbit_r83_c171 bl[171] br[171] wl[83] vdd gnd cell_6t
Xbit_r84_c171 bl[171] br[171] wl[84] vdd gnd cell_6t
Xbit_r85_c171 bl[171] br[171] wl[85] vdd gnd cell_6t
Xbit_r86_c171 bl[171] br[171] wl[86] vdd gnd cell_6t
Xbit_r87_c171 bl[171] br[171] wl[87] vdd gnd cell_6t
Xbit_r88_c171 bl[171] br[171] wl[88] vdd gnd cell_6t
Xbit_r89_c171 bl[171] br[171] wl[89] vdd gnd cell_6t
Xbit_r90_c171 bl[171] br[171] wl[90] vdd gnd cell_6t
Xbit_r91_c171 bl[171] br[171] wl[91] vdd gnd cell_6t
Xbit_r92_c171 bl[171] br[171] wl[92] vdd gnd cell_6t
Xbit_r93_c171 bl[171] br[171] wl[93] vdd gnd cell_6t
Xbit_r94_c171 bl[171] br[171] wl[94] vdd gnd cell_6t
Xbit_r95_c171 bl[171] br[171] wl[95] vdd gnd cell_6t
Xbit_r96_c171 bl[171] br[171] wl[96] vdd gnd cell_6t
Xbit_r97_c171 bl[171] br[171] wl[97] vdd gnd cell_6t
Xbit_r98_c171 bl[171] br[171] wl[98] vdd gnd cell_6t
Xbit_r99_c171 bl[171] br[171] wl[99] vdd gnd cell_6t
Xbit_r100_c171 bl[171] br[171] wl[100] vdd gnd cell_6t
Xbit_r101_c171 bl[171] br[171] wl[101] vdd gnd cell_6t
Xbit_r102_c171 bl[171] br[171] wl[102] vdd gnd cell_6t
Xbit_r103_c171 bl[171] br[171] wl[103] vdd gnd cell_6t
Xbit_r104_c171 bl[171] br[171] wl[104] vdd gnd cell_6t
Xbit_r105_c171 bl[171] br[171] wl[105] vdd gnd cell_6t
Xbit_r106_c171 bl[171] br[171] wl[106] vdd gnd cell_6t
Xbit_r107_c171 bl[171] br[171] wl[107] vdd gnd cell_6t
Xbit_r108_c171 bl[171] br[171] wl[108] vdd gnd cell_6t
Xbit_r109_c171 bl[171] br[171] wl[109] vdd gnd cell_6t
Xbit_r110_c171 bl[171] br[171] wl[110] vdd gnd cell_6t
Xbit_r111_c171 bl[171] br[171] wl[111] vdd gnd cell_6t
Xbit_r112_c171 bl[171] br[171] wl[112] vdd gnd cell_6t
Xbit_r113_c171 bl[171] br[171] wl[113] vdd gnd cell_6t
Xbit_r114_c171 bl[171] br[171] wl[114] vdd gnd cell_6t
Xbit_r115_c171 bl[171] br[171] wl[115] vdd gnd cell_6t
Xbit_r116_c171 bl[171] br[171] wl[116] vdd gnd cell_6t
Xbit_r117_c171 bl[171] br[171] wl[117] vdd gnd cell_6t
Xbit_r118_c171 bl[171] br[171] wl[118] vdd gnd cell_6t
Xbit_r119_c171 bl[171] br[171] wl[119] vdd gnd cell_6t
Xbit_r120_c171 bl[171] br[171] wl[120] vdd gnd cell_6t
Xbit_r121_c171 bl[171] br[171] wl[121] vdd gnd cell_6t
Xbit_r122_c171 bl[171] br[171] wl[122] vdd gnd cell_6t
Xbit_r123_c171 bl[171] br[171] wl[123] vdd gnd cell_6t
Xbit_r124_c171 bl[171] br[171] wl[124] vdd gnd cell_6t
Xbit_r125_c171 bl[171] br[171] wl[125] vdd gnd cell_6t
Xbit_r126_c171 bl[171] br[171] wl[126] vdd gnd cell_6t
Xbit_r127_c171 bl[171] br[171] wl[127] vdd gnd cell_6t
Xbit_r128_c171 bl[171] br[171] wl[128] vdd gnd cell_6t
Xbit_r129_c171 bl[171] br[171] wl[129] vdd gnd cell_6t
Xbit_r130_c171 bl[171] br[171] wl[130] vdd gnd cell_6t
Xbit_r131_c171 bl[171] br[171] wl[131] vdd gnd cell_6t
Xbit_r132_c171 bl[171] br[171] wl[132] vdd gnd cell_6t
Xbit_r133_c171 bl[171] br[171] wl[133] vdd gnd cell_6t
Xbit_r134_c171 bl[171] br[171] wl[134] vdd gnd cell_6t
Xbit_r135_c171 bl[171] br[171] wl[135] vdd gnd cell_6t
Xbit_r136_c171 bl[171] br[171] wl[136] vdd gnd cell_6t
Xbit_r137_c171 bl[171] br[171] wl[137] vdd gnd cell_6t
Xbit_r138_c171 bl[171] br[171] wl[138] vdd gnd cell_6t
Xbit_r139_c171 bl[171] br[171] wl[139] vdd gnd cell_6t
Xbit_r140_c171 bl[171] br[171] wl[140] vdd gnd cell_6t
Xbit_r141_c171 bl[171] br[171] wl[141] vdd gnd cell_6t
Xbit_r142_c171 bl[171] br[171] wl[142] vdd gnd cell_6t
Xbit_r143_c171 bl[171] br[171] wl[143] vdd gnd cell_6t
Xbit_r144_c171 bl[171] br[171] wl[144] vdd gnd cell_6t
Xbit_r145_c171 bl[171] br[171] wl[145] vdd gnd cell_6t
Xbit_r146_c171 bl[171] br[171] wl[146] vdd gnd cell_6t
Xbit_r147_c171 bl[171] br[171] wl[147] vdd gnd cell_6t
Xbit_r148_c171 bl[171] br[171] wl[148] vdd gnd cell_6t
Xbit_r149_c171 bl[171] br[171] wl[149] vdd gnd cell_6t
Xbit_r150_c171 bl[171] br[171] wl[150] vdd gnd cell_6t
Xbit_r151_c171 bl[171] br[171] wl[151] vdd gnd cell_6t
Xbit_r152_c171 bl[171] br[171] wl[152] vdd gnd cell_6t
Xbit_r153_c171 bl[171] br[171] wl[153] vdd gnd cell_6t
Xbit_r154_c171 bl[171] br[171] wl[154] vdd gnd cell_6t
Xbit_r155_c171 bl[171] br[171] wl[155] vdd gnd cell_6t
Xbit_r156_c171 bl[171] br[171] wl[156] vdd gnd cell_6t
Xbit_r157_c171 bl[171] br[171] wl[157] vdd gnd cell_6t
Xbit_r158_c171 bl[171] br[171] wl[158] vdd gnd cell_6t
Xbit_r159_c171 bl[171] br[171] wl[159] vdd gnd cell_6t
Xbit_r160_c171 bl[171] br[171] wl[160] vdd gnd cell_6t
Xbit_r161_c171 bl[171] br[171] wl[161] vdd gnd cell_6t
Xbit_r162_c171 bl[171] br[171] wl[162] vdd gnd cell_6t
Xbit_r163_c171 bl[171] br[171] wl[163] vdd gnd cell_6t
Xbit_r164_c171 bl[171] br[171] wl[164] vdd gnd cell_6t
Xbit_r165_c171 bl[171] br[171] wl[165] vdd gnd cell_6t
Xbit_r166_c171 bl[171] br[171] wl[166] vdd gnd cell_6t
Xbit_r167_c171 bl[171] br[171] wl[167] vdd gnd cell_6t
Xbit_r168_c171 bl[171] br[171] wl[168] vdd gnd cell_6t
Xbit_r169_c171 bl[171] br[171] wl[169] vdd gnd cell_6t
Xbit_r170_c171 bl[171] br[171] wl[170] vdd gnd cell_6t
Xbit_r171_c171 bl[171] br[171] wl[171] vdd gnd cell_6t
Xbit_r172_c171 bl[171] br[171] wl[172] vdd gnd cell_6t
Xbit_r173_c171 bl[171] br[171] wl[173] vdd gnd cell_6t
Xbit_r174_c171 bl[171] br[171] wl[174] vdd gnd cell_6t
Xbit_r175_c171 bl[171] br[171] wl[175] vdd gnd cell_6t
Xbit_r176_c171 bl[171] br[171] wl[176] vdd gnd cell_6t
Xbit_r177_c171 bl[171] br[171] wl[177] vdd gnd cell_6t
Xbit_r178_c171 bl[171] br[171] wl[178] vdd gnd cell_6t
Xbit_r179_c171 bl[171] br[171] wl[179] vdd gnd cell_6t
Xbit_r180_c171 bl[171] br[171] wl[180] vdd gnd cell_6t
Xbit_r181_c171 bl[171] br[171] wl[181] vdd gnd cell_6t
Xbit_r182_c171 bl[171] br[171] wl[182] vdd gnd cell_6t
Xbit_r183_c171 bl[171] br[171] wl[183] vdd gnd cell_6t
Xbit_r184_c171 bl[171] br[171] wl[184] vdd gnd cell_6t
Xbit_r185_c171 bl[171] br[171] wl[185] vdd gnd cell_6t
Xbit_r186_c171 bl[171] br[171] wl[186] vdd gnd cell_6t
Xbit_r187_c171 bl[171] br[171] wl[187] vdd gnd cell_6t
Xbit_r188_c171 bl[171] br[171] wl[188] vdd gnd cell_6t
Xbit_r189_c171 bl[171] br[171] wl[189] vdd gnd cell_6t
Xbit_r190_c171 bl[171] br[171] wl[190] vdd gnd cell_6t
Xbit_r191_c171 bl[171] br[171] wl[191] vdd gnd cell_6t
Xbit_r192_c171 bl[171] br[171] wl[192] vdd gnd cell_6t
Xbit_r193_c171 bl[171] br[171] wl[193] vdd gnd cell_6t
Xbit_r194_c171 bl[171] br[171] wl[194] vdd gnd cell_6t
Xbit_r195_c171 bl[171] br[171] wl[195] vdd gnd cell_6t
Xbit_r196_c171 bl[171] br[171] wl[196] vdd gnd cell_6t
Xbit_r197_c171 bl[171] br[171] wl[197] vdd gnd cell_6t
Xbit_r198_c171 bl[171] br[171] wl[198] vdd gnd cell_6t
Xbit_r199_c171 bl[171] br[171] wl[199] vdd gnd cell_6t
Xbit_r200_c171 bl[171] br[171] wl[200] vdd gnd cell_6t
Xbit_r201_c171 bl[171] br[171] wl[201] vdd gnd cell_6t
Xbit_r202_c171 bl[171] br[171] wl[202] vdd gnd cell_6t
Xbit_r203_c171 bl[171] br[171] wl[203] vdd gnd cell_6t
Xbit_r204_c171 bl[171] br[171] wl[204] vdd gnd cell_6t
Xbit_r205_c171 bl[171] br[171] wl[205] vdd gnd cell_6t
Xbit_r206_c171 bl[171] br[171] wl[206] vdd gnd cell_6t
Xbit_r207_c171 bl[171] br[171] wl[207] vdd gnd cell_6t
Xbit_r208_c171 bl[171] br[171] wl[208] vdd gnd cell_6t
Xbit_r209_c171 bl[171] br[171] wl[209] vdd gnd cell_6t
Xbit_r210_c171 bl[171] br[171] wl[210] vdd gnd cell_6t
Xbit_r211_c171 bl[171] br[171] wl[211] vdd gnd cell_6t
Xbit_r212_c171 bl[171] br[171] wl[212] vdd gnd cell_6t
Xbit_r213_c171 bl[171] br[171] wl[213] vdd gnd cell_6t
Xbit_r214_c171 bl[171] br[171] wl[214] vdd gnd cell_6t
Xbit_r215_c171 bl[171] br[171] wl[215] vdd gnd cell_6t
Xbit_r216_c171 bl[171] br[171] wl[216] vdd gnd cell_6t
Xbit_r217_c171 bl[171] br[171] wl[217] vdd gnd cell_6t
Xbit_r218_c171 bl[171] br[171] wl[218] vdd gnd cell_6t
Xbit_r219_c171 bl[171] br[171] wl[219] vdd gnd cell_6t
Xbit_r220_c171 bl[171] br[171] wl[220] vdd gnd cell_6t
Xbit_r221_c171 bl[171] br[171] wl[221] vdd gnd cell_6t
Xbit_r222_c171 bl[171] br[171] wl[222] vdd gnd cell_6t
Xbit_r223_c171 bl[171] br[171] wl[223] vdd gnd cell_6t
Xbit_r224_c171 bl[171] br[171] wl[224] vdd gnd cell_6t
Xbit_r225_c171 bl[171] br[171] wl[225] vdd gnd cell_6t
Xbit_r226_c171 bl[171] br[171] wl[226] vdd gnd cell_6t
Xbit_r227_c171 bl[171] br[171] wl[227] vdd gnd cell_6t
Xbit_r228_c171 bl[171] br[171] wl[228] vdd gnd cell_6t
Xbit_r229_c171 bl[171] br[171] wl[229] vdd gnd cell_6t
Xbit_r230_c171 bl[171] br[171] wl[230] vdd gnd cell_6t
Xbit_r231_c171 bl[171] br[171] wl[231] vdd gnd cell_6t
Xbit_r232_c171 bl[171] br[171] wl[232] vdd gnd cell_6t
Xbit_r233_c171 bl[171] br[171] wl[233] vdd gnd cell_6t
Xbit_r234_c171 bl[171] br[171] wl[234] vdd gnd cell_6t
Xbit_r235_c171 bl[171] br[171] wl[235] vdd gnd cell_6t
Xbit_r236_c171 bl[171] br[171] wl[236] vdd gnd cell_6t
Xbit_r237_c171 bl[171] br[171] wl[237] vdd gnd cell_6t
Xbit_r238_c171 bl[171] br[171] wl[238] vdd gnd cell_6t
Xbit_r239_c171 bl[171] br[171] wl[239] vdd gnd cell_6t
Xbit_r240_c171 bl[171] br[171] wl[240] vdd gnd cell_6t
Xbit_r241_c171 bl[171] br[171] wl[241] vdd gnd cell_6t
Xbit_r242_c171 bl[171] br[171] wl[242] vdd gnd cell_6t
Xbit_r243_c171 bl[171] br[171] wl[243] vdd gnd cell_6t
Xbit_r244_c171 bl[171] br[171] wl[244] vdd gnd cell_6t
Xbit_r245_c171 bl[171] br[171] wl[245] vdd gnd cell_6t
Xbit_r246_c171 bl[171] br[171] wl[246] vdd gnd cell_6t
Xbit_r247_c171 bl[171] br[171] wl[247] vdd gnd cell_6t
Xbit_r248_c171 bl[171] br[171] wl[248] vdd gnd cell_6t
Xbit_r249_c171 bl[171] br[171] wl[249] vdd gnd cell_6t
Xbit_r250_c171 bl[171] br[171] wl[250] vdd gnd cell_6t
Xbit_r251_c171 bl[171] br[171] wl[251] vdd gnd cell_6t
Xbit_r252_c171 bl[171] br[171] wl[252] vdd gnd cell_6t
Xbit_r253_c171 bl[171] br[171] wl[253] vdd gnd cell_6t
Xbit_r254_c171 bl[171] br[171] wl[254] vdd gnd cell_6t
Xbit_r255_c171 bl[171] br[171] wl[255] vdd gnd cell_6t
Xbit_r0_c172 bl[172] br[172] wl[0] vdd gnd cell_6t
Xbit_r1_c172 bl[172] br[172] wl[1] vdd gnd cell_6t
Xbit_r2_c172 bl[172] br[172] wl[2] vdd gnd cell_6t
Xbit_r3_c172 bl[172] br[172] wl[3] vdd gnd cell_6t
Xbit_r4_c172 bl[172] br[172] wl[4] vdd gnd cell_6t
Xbit_r5_c172 bl[172] br[172] wl[5] vdd gnd cell_6t
Xbit_r6_c172 bl[172] br[172] wl[6] vdd gnd cell_6t
Xbit_r7_c172 bl[172] br[172] wl[7] vdd gnd cell_6t
Xbit_r8_c172 bl[172] br[172] wl[8] vdd gnd cell_6t
Xbit_r9_c172 bl[172] br[172] wl[9] vdd gnd cell_6t
Xbit_r10_c172 bl[172] br[172] wl[10] vdd gnd cell_6t
Xbit_r11_c172 bl[172] br[172] wl[11] vdd gnd cell_6t
Xbit_r12_c172 bl[172] br[172] wl[12] vdd gnd cell_6t
Xbit_r13_c172 bl[172] br[172] wl[13] vdd gnd cell_6t
Xbit_r14_c172 bl[172] br[172] wl[14] vdd gnd cell_6t
Xbit_r15_c172 bl[172] br[172] wl[15] vdd gnd cell_6t
Xbit_r16_c172 bl[172] br[172] wl[16] vdd gnd cell_6t
Xbit_r17_c172 bl[172] br[172] wl[17] vdd gnd cell_6t
Xbit_r18_c172 bl[172] br[172] wl[18] vdd gnd cell_6t
Xbit_r19_c172 bl[172] br[172] wl[19] vdd gnd cell_6t
Xbit_r20_c172 bl[172] br[172] wl[20] vdd gnd cell_6t
Xbit_r21_c172 bl[172] br[172] wl[21] vdd gnd cell_6t
Xbit_r22_c172 bl[172] br[172] wl[22] vdd gnd cell_6t
Xbit_r23_c172 bl[172] br[172] wl[23] vdd gnd cell_6t
Xbit_r24_c172 bl[172] br[172] wl[24] vdd gnd cell_6t
Xbit_r25_c172 bl[172] br[172] wl[25] vdd gnd cell_6t
Xbit_r26_c172 bl[172] br[172] wl[26] vdd gnd cell_6t
Xbit_r27_c172 bl[172] br[172] wl[27] vdd gnd cell_6t
Xbit_r28_c172 bl[172] br[172] wl[28] vdd gnd cell_6t
Xbit_r29_c172 bl[172] br[172] wl[29] vdd gnd cell_6t
Xbit_r30_c172 bl[172] br[172] wl[30] vdd gnd cell_6t
Xbit_r31_c172 bl[172] br[172] wl[31] vdd gnd cell_6t
Xbit_r32_c172 bl[172] br[172] wl[32] vdd gnd cell_6t
Xbit_r33_c172 bl[172] br[172] wl[33] vdd gnd cell_6t
Xbit_r34_c172 bl[172] br[172] wl[34] vdd gnd cell_6t
Xbit_r35_c172 bl[172] br[172] wl[35] vdd gnd cell_6t
Xbit_r36_c172 bl[172] br[172] wl[36] vdd gnd cell_6t
Xbit_r37_c172 bl[172] br[172] wl[37] vdd gnd cell_6t
Xbit_r38_c172 bl[172] br[172] wl[38] vdd gnd cell_6t
Xbit_r39_c172 bl[172] br[172] wl[39] vdd gnd cell_6t
Xbit_r40_c172 bl[172] br[172] wl[40] vdd gnd cell_6t
Xbit_r41_c172 bl[172] br[172] wl[41] vdd gnd cell_6t
Xbit_r42_c172 bl[172] br[172] wl[42] vdd gnd cell_6t
Xbit_r43_c172 bl[172] br[172] wl[43] vdd gnd cell_6t
Xbit_r44_c172 bl[172] br[172] wl[44] vdd gnd cell_6t
Xbit_r45_c172 bl[172] br[172] wl[45] vdd gnd cell_6t
Xbit_r46_c172 bl[172] br[172] wl[46] vdd gnd cell_6t
Xbit_r47_c172 bl[172] br[172] wl[47] vdd gnd cell_6t
Xbit_r48_c172 bl[172] br[172] wl[48] vdd gnd cell_6t
Xbit_r49_c172 bl[172] br[172] wl[49] vdd gnd cell_6t
Xbit_r50_c172 bl[172] br[172] wl[50] vdd gnd cell_6t
Xbit_r51_c172 bl[172] br[172] wl[51] vdd gnd cell_6t
Xbit_r52_c172 bl[172] br[172] wl[52] vdd gnd cell_6t
Xbit_r53_c172 bl[172] br[172] wl[53] vdd gnd cell_6t
Xbit_r54_c172 bl[172] br[172] wl[54] vdd gnd cell_6t
Xbit_r55_c172 bl[172] br[172] wl[55] vdd gnd cell_6t
Xbit_r56_c172 bl[172] br[172] wl[56] vdd gnd cell_6t
Xbit_r57_c172 bl[172] br[172] wl[57] vdd gnd cell_6t
Xbit_r58_c172 bl[172] br[172] wl[58] vdd gnd cell_6t
Xbit_r59_c172 bl[172] br[172] wl[59] vdd gnd cell_6t
Xbit_r60_c172 bl[172] br[172] wl[60] vdd gnd cell_6t
Xbit_r61_c172 bl[172] br[172] wl[61] vdd gnd cell_6t
Xbit_r62_c172 bl[172] br[172] wl[62] vdd gnd cell_6t
Xbit_r63_c172 bl[172] br[172] wl[63] vdd gnd cell_6t
Xbit_r64_c172 bl[172] br[172] wl[64] vdd gnd cell_6t
Xbit_r65_c172 bl[172] br[172] wl[65] vdd gnd cell_6t
Xbit_r66_c172 bl[172] br[172] wl[66] vdd gnd cell_6t
Xbit_r67_c172 bl[172] br[172] wl[67] vdd gnd cell_6t
Xbit_r68_c172 bl[172] br[172] wl[68] vdd gnd cell_6t
Xbit_r69_c172 bl[172] br[172] wl[69] vdd gnd cell_6t
Xbit_r70_c172 bl[172] br[172] wl[70] vdd gnd cell_6t
Xbit_r71_c172 bl[172] br[172] wl[71] vdd gnd cell_6t
Xbit_r72_c172 bl[172] br[172] wl[72] vdd gnd cell_6t
Xbit_r73_c172 bl[172] br[172] wl[73] vdd gnd cell_6t
Xbit_r74_c172 bl[172] br[172] wl[74] vdd gnd cell_6t
Xbit_r75_c172 bl[172] br[172] wl[75] vdd gnd cell_6t
Xbit_r76_c172 bl[172] br[172] wl[76] vdd gnd cell_6t
Xbit_r77_c172 bl[172] br[172] wl[77] vdd gnd cell_6t
Xbit_r78_c172 bl[172] br[172] wl[78] vdd gnd cell_6t
Xbit_r79_c172 bl[172] br[172] wl[79] vdd gnd cell_6t
Xbit_r80_c172 bl[172] br[172] wl[80] vdd gnd cell_6t
Xbit_r81_c172 bl[172] br[172] wl[81] vdd gnd cell_6t
Xbit_r82_c172 bl[172] br[172] wl[82] vdd gnd cell_6t
Xbit_r83_c172 bl[172] br[172] wl[83] vdd gnd cell_6t
Xbit_r84_c172 bl[172] br[172] wl[84] vdd gnd cell_6t
Xbit_r85_c172 bl[172] br[172] wl[85] vdd gnd cell_6t
Xbit_r86_c172 bl[172] br[172] wl[86] vdd gnd cell_6t
Xbit_r87_c172 bl[172] br[172] wl[87] vdd gnd cell_6t
Xbit_r88_c172 bl[172] br[172] wl[88] vdd gnd cell_6t
Xbit_r89_c172 bl[172] br[172] wl[89] vdd gnd cell_6t
Xbit_r90_c172 bl[172] br[172] wl[90] vdd gnd cell_6t
Xbit_r91_c172 bl[172] br[172] wl[91] vdd gnd cell_6t
Xbit_r92_c172 bl[172] br[172] wl[92] vdd gnd cell_6t
Xbit_r93_c172 bl[172] br[172] wl[93] vdd gnd cell_6t
Xbit_r94_c172 bl[172] br[172] wl[94] vdd gnd cell_6t
Xbit_r95_c172 bl[172] br[172] wl[95] vdd gnd cell_6t
Xbit_r96_c172 bl[172] br[172] wl[96] vdd gnd cell_6t
Xbit_r97_c172 bl[172] br[172] wl[97] vdd gnd cell_6t
Xbit_r98_c172 bl[172] br[172] wl[98] vdd gnd cell_6t
Xbit_r99_c172 bl[172] br[172] wl[99] vdd gnd cell_6t
Xbit_r100_c172 bl[172] br[172] wl[100] vdd gnd cell_6t
Xbit_r101_c172 bl[172] br[172] wl[101] vdd gnd cell_6t
Xbit_r102_c172 bl[172] br[172] wl[102] vdd gnd cell_6t
Xbit_r103_c172 bl[172] br[172] wl[103] vdd gnd cell_6t
Xbit_r104_c172 bl[172] br[172] wl[104] vdd gnd cell_6t
Xbit_r105_c172 bl[172] br[172] wl[105] vdd gnd cell_6t
Xbit_r106_c172 bl[172] br[172] wl[106] vdd gnd cell_6t
Xbit_r107_c172 bl[172] br[172] wl[107] vdd gnd cell_6t
Xbit_r108_c172 bl[172] br[172] wl[108] vdd gnd cell_6t
Xbit_r109_c172 bl[172] br[172] wl[109] vdd gnd cell_6t
Xbit_r110_c172 bl[172] br[172] wl[110] vdd gnd cell_6t
Xbit_r111_c172 bl[172] br[172] wl[111] vdd gnd cell_6t
Xbit_r112_c172 bl[172] br[172] wl[112] vdd gnd cell_6t
Xbit_r113_c172 bl[172] br[172] wl[113] vdd gnd cell_6t
Xbit_r114_c172 bl[172] br[172] wl[114] vdd gnd cell_6t
Xbit_r115_c172 bl[172] br[172] wl[115] vdd gnd cell_6t
Xbit_r116_c172 bl[172] br[172] wl[116] vdd gnd cell_6t
Xbit_r117_c172 bl[172] br[172] wl[117] vdd gnd cell_6t
Xbit_r118_c172 bl[172] br[172] wl[118] vdd gnd cell_6t
Xbit_r119_c172 bl[172] br[172] wl[119] vdd gnd cell_6t
Xbit_r120_c172 bl[172] br[172] wl[120] vdd gnd cell_6t
Xbit_r121_c172 bl[172] br[172] wl[121] vdd gnd cell_6t
Xbit_r122_c172 bl[172] br[172] wl[122] vdd gnd cell_6t
Xbit_r123_c172 bl[172] br[172] wl[123] vdd gnd cell_6t
Xbit_r124_c172 bl[172] br[172] wl[124] vdd gnd cell_6t
Xbit_r125_c172 bl[172] br[172] wl[125] vdd gnd cell_6t
Xbit_r126_c172 bl[172] br[172] wl[126] vdd gnd cell_6t
Xbit_r127_c172 bl[172] br[172] wl[127] vdd gnd cell_6t
Xbit_r128_c172 bl[172] br[172] wl[128] vdd gnd cell_6t
Xbit_r129_c172 bl[172] br[172] wl[129] vdd gnd cell_6t
Xbit_r130_c172 bl[172] br[172] wl[130] vdd gnd cell_6t
Xbit_r131_c172 bl[172] br[172] wl[131] vdd gnd cell_6t
Xbit_r132_c172 bl[172] br[172] wl[132] vdd gnd cell_6t
Xbit_r133_c172 bl[172] br[172] wl[133] vdd gnd cell_6t
Xbit_r134_c172 bl[172] br[172] wl[134] vdd gnd cell_6t
Xbit_r135_c172 bl[172] br[172] wl[135] vdd gnd cell_6t
Xbit_r136_c172 bl[172] br[172] wl[136] vdd gnd cell_6t
Xbit_r137_c172 bl[172] br[172] wl[137] vdd gnd cell_6t
Xbit_r138_c172 bl[172] br[172] wl[138] vdd gnd cell_6t
Xbit_r139_c172 bl[172] br[172] wl[139] vdd gnd cell_6t
Xbit_r140_c172 bl[172] br[172] wl[140] vdd gnd cell_6t
Xbit_r141_c172 bl[172] br[172] wl[141] vdd gnd cell_6t
Xbit_r142_c172 bl[172] br[172] wl[142] vdd gnd cell_6t
Xbit_r143_c172 bl[172] br[172] wl[143] vdd gnd cell_6t
Xbit_r144_c172 bl[172] br[172] wl[144] vdd gnd cell_6t
Xbit_r145_c172 bl[172] br[172] wl[145] vdd gnd cell_6t
Xbit_r146_c172 bl[172] br[172] wl[146] vdd gnd cell_6t
Xbit_r147_c172 bl[172] br[172] wl[147] vdd gnd cell_6t
Xbit_r148_c172 bl[172] br[172] wl[148] vdd gnd cell_6t
Xbit_r149_c172 bl[172] br[172] wl[149] vdd gnd cell_6t
Xbit_r150_c172 bl[172] br[172] wl[150] vdd gnd cell_6t
Xbit_r151_c172 bl[172] br[172] wl[151] vdd gnd cell_6t
Xbit_r152_c172 bl[172] br[172] wl[152] vdd gnd cell_6t
Xbit_r153_c172 bl[172] br[172] wl[153] vdd gnd cell_6t
Xbit_r154_c172 bl[172] br[172] wl[154] vdd gnd cell_6t
Xbit_r155_c172 bl[172] br[172] wl[155] vdd gnd cell_6t
Xbit_r156_c172 bl[172] br[172] wl[156] vdd gnd cell_6t
Xbit_r157_c172 bl[172] br[172] wl[157] vdd gnd cell_6t
Xbit_r158_c172 bl[172] br[172] wl[158] vdd gnd cell_6t
Xbit_r159_c172 bl[172] br[172] wl[159] vdd gnd cell_6t
Xbit_r160_c172 bl[172] br[172] wl[160] vdd gnd cell_6t
Xbit_r161_c172 bl[172] br[172] wl[161] vdd gnd cell_6t
Xbit_r162_c172 bl[172] br[172] wl[162] vdd gnd cell_6t
Xbit_r163_c172 bl[172] br[172] wl[163] vdd gnd cell_6t
Xbit_r164_c172 bl[172] br[172] wl[164] vdd gnd cell_6t
Xbit_r165_c172 bl[172] br[172] wl[165] vdd gnd cell_6t
Xbit_r166_c172 bl[172] br[172] wl[166] vdd gnd cell_6t
Xbit_r167_c172 bl[172] br[172] wl[167] vdd gnd cell_6t
Xbit_r168_c172 bl[172] br[172] wl[168] vdd gnd cell_6t
Xbit_r169_c172 bl[172] br[172] wl[169] vdd gnd cell_6t
Xbit_r170_c172 bl[172] br[172] wl[170] vdd gnd cell_6t
Xbit_r171_c172 bl[172] br[172] wl[171] vdd gnd cell_6t
Xbit_r172_c172 bl[172] br[172] wl[172] vdd gnd cell_6t
Xbit_r173_c172 bl[172] br[172] wl[173] vdd gnd cell_6t
Xbit_r174_c172 bl[172] br[172] wl[174] vdd gnd cell_6t
Xbit_r175_c172 bl[172] br[172] wl[175] vdd gnd cell_6t
Xbit_r176_c172 bl[172] br[172] wl[176] vdd gnd cell_6t
Xbit_r177_c172 bl[172] br[172] wl[177] vdd gnd cell_6t
Xbit_r178_c172 bl[172] br[172] wl[178] vdd gnd cell_6t
Xbit_r179_c172 bl[172] br[172] wl[179] vdd gnd cell_6t
Xbit_r180_c172 bl[172] br[172] wl[180] vdd gnd cell_6t
Xbit_r181_c172 bl[172] br[172] wl[181] vdd gnd cell_6t
Xbit_r182_c172 bl[172] br[172] wl[182] vdd gnd cell_6t
Xbit_r183_c172 bl[172] br[172] wl[183] vdd gnd cell_6t
Xbit_r184_c172 bl[172] br[172] wl[184] vdd gnd cell_6t
Xbit_r185_c172 bl[172] br[172] wl[185] vdd gnd cell_6t
Xbit_r186_c172 bl[172] br[172] wl[186] vdd gnd cell_6t
Xbit_r187_c172 bl[172] br[172] wl[187] vdd gnd cell_6t
Xbit_r188_c172 bl[172] br[172] wl[188] vdd gnd cell_6t
Xbit_r189_c172 bl[172] br[172] wl[189] vdd gnd cell_6t
Xbit_r190_c172 bl[172] br[172] wl[190] vdd gnd cell_6t
Xbit_r191_c172 bl[172] br[172] wl[191] vdd gnd cell_6t
Xbit_r192_c172 bl[172] br[172] wl[192] vdd gnd cell_6t
Xbit_r193_c172 bl[172] br[172] wl[193] vdd gnd cell_6t
Xbit_r194_c172 bl[172] br[172] wl[194] vdd gnd cell_6t
Xbit_r195_c172 bl[172] br[172] wl[195] vdd gnd cell_6t
Xbit_r196_c172 bl[172] br[172] wl[196] vdd gnd cell_6t
Xbit_r197_c172 bl[172] br[172] wl[197] vdd gnd cell_6t
Xbit_r198_c172 bl[172] br[172] wl[198] vdd gnd cell_6t
Xbit_r199_c172 bl[172] br[172] wl[199] vdd gnd cell_6t
Xbit_r200_c172 bl[172] br[172] wl[200] vdd gnd cell_6t
Xbit_r201_c172 bl[172] br[172] wl[201] vdd gnd cell_6t
Xbit_r202_c172 bl[172] br[172] wl[202] vdd gnd cell_6t
Xbit_r203_c172 bl[172] br[172] wl[203] vdd gnd cell_6t
Xbit_r204_c172 bl[172] br[172] wl[204] vdd gnd cell_6t
Xbit_r205_c172 bl[172] br[172] wl[205] vdd gnd cell_6t
Xbit_r206_c172 bl[172] br[172] wl[206] vdd gnd cell_6t
Xbit_r207_c172 bl[172] br[172] wl[207] vdd gnd cell_6t
Xbit_r208_c172 bl[172] br[172] wl[208] vdd gnd cell_6t
Xbit_r209_c172 bl[172] br[172] wl[209] vdd gnd cell_6t
Xbit_r210_c172 bl[172] br[172] wl[210] vdd gnd cell_6t
Xbit_r211_c172 bl[172] br[172] wl[211] vdd gnd cell_6t
Xbit_r212_c172 bl[172] br[172] wl[212] vdd gnd cell_6t
Xbit_r213_c172 bl[172] br[172] wl[213] vdd gnd cell_6t
Xbit_r214_c172 bl[172] br[172] wl[214] vdd gnd cell_6t
Xbit_r215_c172 bl[172] br[172] wl[215] vdd gnd cell_6t
Xbit_r216_c172 bl[172] br[172] wl[216] vdd gnd cell_6t
Xbit_r217_c172 bl[172] br[172] wl[217] vdd gnd cell_6t
Xbit_r218_c172 bl[172] br[172] wl[218] vdd gnd cell_6t
Xbit_r219_c172 bl[172] br[172] wl[219] vdd gnd cell_6t
Xbit_r220_c172 bl[172] br[172] wl[220] vdd gnd cell_6t
Xbit_r221_c172 bl[172] br[172] wl[221] vdd gnd cell_6t
Xbit_r222_c172 bl[172] br[172] wl[222] vdd gnd cell_6t
Xbit_r223_c172 bl[172] br[172] wl[223] vdd gnd cell_6t
Xbit_r224_c172 bl[172] br[172] wl[224] vdd gnd cell_6t
Xbit_r225_c172 bl[172] br[172] wl[225] vdd gnd cell_6t
Xbit_r226_c172 bl[172] br[172] wl[226] vdd gnd cell_6t
Xbit_r227_c172 bl[172] br[172] wl[227] vdd gnd cell_6t
Xbit_r228_c172 bl[172] br[172] wl[228] vdd gnd cell_6t
Xbit_r229_c172 bl[172] br[172] wl[229] vdd gnd cell_6t
Xbit_r230_c172 bl[172] br[172] wl[230] vdd gnd cell_6t
Xbit_r231_c172 bl[172] br[172] wl[231] vdd gnd cell_6t
Xbit_r232_c172 bl[172] br[172] wl[232] vdd gnd cell_6t
Xbit_r233_c172 bl[172] br[172] wl[233] vdd gnd cell_6t
Xbit_r234_c172 bl[172] br[172] wl[234] vdd gnd cell_6t
Xbit_r235_c172 bl[172] br[172] wl[235] vdd gnd cell_6t
Xbit_r236_c172 bl[172] br[172] wl[236] vdd gnd cell_6t
Xbit_r237_c172 bl[172] br[172] wl[237] vdd gnd cell_6t
Xbit_r238_c172 bl[172] br[172] wl[238] vdd gnd cell_6t
Xbit_r239_c172 bl[172] br[172] wl[239] vdd gnd cell_6t
Xbit_r240_c172 bl[172] br[172] wl[240] vdd gnd cell_6t
Xbit_r241_c172 bl[172] br[172] wl[241] vdd gnd cell_6t
Xbit_r242_c172 bl[172] br[172] wl[242] vdd gnd cell_6t
Xbit_r243_c172 bl[172] br[172] wl[243] vdd gnd cell_6t
Xbit_r244_c172 bl[172] br[172] wl[244] vdd gnd cell_6t
Xbit_r245_c172 bl[172] br[172] wl[245] vdd gnd cell_6t
Xbit_r246_c172 bl[172] br[172] wl[246] vdd gnd cell_6t
Xbit_r247_c172 bl[172] br[172] wl[247] vdd gnd cell_6t
Xbit_r248_c172 bl[172] br[172] wl[248] vdd gnd cell_6t
Xbit_r249_c172 bl[172] br[172] wl[249] vdd gnd cell_6t
Xbit_r250_c172 bl[172] br[172] wl[250] vdd gnd cell_6t
Xbit_r251_c172 bl[172] br[172] wl[251] vdd gnd cell_6t
Xbit_r252_c172 bl[172] br[172] wl[252] vdd gnd cell_6t
Xbit_r253_c172 bl[172] br[172] wl[253] vdd gnd cell_6t
Xbit_r254_c172 bl[172] br[172] wl[254] vdd gnd cell_6t
Xbit_r255_c172 bl[172] br[172] wl[255] vdd gnd cell_6t
Xbit_r0_c173 bl[173] br[173] wl[0] vdd gnd cell_6t
Xbit_r1_c173 bl[173] br[173] wl[1] vdd gnd cell_6t
Xbit_r2_c173 bl[173] br[173] wl[2] vdd gnd cell_6t
Xbit_r3_c173 bl[173] br[173] wl[3] vdd gnd cell_6t
Xbit_r4_c173 bl[173] br[173] wl[4] vdd gnd cell_6t
Xbit_r5_c173 bl[173] br[173] wl[5] vdd gnd cell_6t
Xbit_r6_c173 bl[173] br[173] wl[6] vdd gnd cell_6t
Xbit_r7_c173 bl[173] br[173] wl[7] vdd gnd cell_6t
Xbit_r8_c173 bl[173] br[173] wl[8] vdd gnd cell_6t
Xbit_r9_c173 bl[173] br[173] wl[9] vdd gnd cell_6t
Xbit_r10_c173 bl[173] br[173] wl[10] vdd gnd cell_6t
Xbit_r11_c173 bl[173] br[173] wl[11] vdd gnd cell_6t
Xbit_r12_c173 bl[173] br[173] wl[12] vdd gnd cell_6t
Xbit_r13_c173 bl[173] br[173] wl[13] vdd gnd cell_6t
Xbit_r14_c173 bl[173] br[173] wl[14] vdd gnd cell_6t
Xbit_r15_c173 bl[173] br[173] wl[15] vdd gnd cell_6t
Xbit_r16_c173 bl[173] br[173] wl[16] vdd gnd cell_6t
Xbit_r17_c173 bl[173] br[173] wl[17] vdd gnd cell_6t
Xbit_r18_c173 bl[173] br[173] wl[18] vdd gnd cell_6t
Xbit_r19_c173 bl[173] br[173] wl[19] vdd gnd cell_6t
Xbit_r20_c173 bl[173] br[173] wl[20] vdd gnd cell_6t
Xbit_r21_c173 bl[173] br[173] wl[21] vdd gnd cell_6t
Xbit_r22_c173 bl[173] br[173] wl[22] vdd gnd cell_6t
Xbit_r23_c173 bl[173] br[173] wl[23] vdd gnd cell_6t
Xbit_r24_c173 bl[173] br[173] wl[24] vdd gnd cell_6t
Xbit_r25_c173 bl[173] br[173] wl[25] vdd gnd cell_6t
Xbit_r26_c173 bl[173] br[173] wl[26] vdd gnd cell_6t
Xbit_r27_c173 bl[173] br[173] wl[27] vdd gnd cell_6t
Xbit_r28_c173 bl[173] br[173] wl[28] vdd gnd cell_6t
Xbit_r29_c173 bl[173] br[173] wl[29] vdd gnd cell_6t
Xbit_r30_c173 bl[173] br[173] wl[30] vdd gnd cell_6t
Xbit_r31_c173 bl[173] br[173] wl[31] vdd gnd cell_6t
Xbit_r32_c173 bl[173] br[173] wl[32] vdd gnd cell_6t
Xbit_r33_c173 bl[173] br[173] wl[33] vdd gnd cell_6t
Xbit_r34_c173 bl[173] br[173] wl[34] vdd gnd cell_6t
Xbit_r35_c173 bl[173] br[173] wl[35] vdd gnd cell_6t
Xbit_r36_c173 bl[173] br[173] wl[36] vdd gnd cell_6t
Xbit_r37_c173 bl[173] br[173] wl[37] vdd gnd cell_6t
Xbit_r38_c173 bl[173] br[173] wl[38] vdd gnd cell_6t
Xbit_r39_c173 bl[173] br[173] wl[39] vdd gnd cell_6t
Xbit_r40_c173 bl[173] br[173] wl[40] vdd gnd cell_6t
Xbit_r41_c173 bl[173] br[173] wl[41] vdd gnd cell_6t
Xbit_r42_c173 bl[173] br[173] wl[42] vdd gnd cell_6t
Xbit_r43_c173 bl[173] br[173] wl[43] vdd gnd cell_6t
Xbit_r44_c173 bl[173] br[173] wl[44] vdd gnd cell_6t
Xbit_r45_c173 bl[173] br[173] wl[45] vdd gnd cell_6t
Xbit_r46_c173 bl[173] br[173] wl[46] vdd gnd cell_6t
Xbit_r47_c173 bl[173] br[173] wl[47] vdd gnd cell_6t
Xbit_r48_c173 bl[173] br[173] wl[48] vdd gnd cell_6t
Xbit_r49_c173 bl[173] br[173] wl[49] vdd gnd cell_6t
Xbit_r50_c173 bl[173] br[173] wl[50] vdd gnd cell_6t
Xbit_r51_c173 bl[173] br[173] wl[51] vdd gnd cell_6t
Xbit_r52_c173 bl[173] br[173] wl[52] vdd gnd cell_6t
Xbit_r53_c173 bl[173] br[173] wl[53] vdd gnd cell_6t
Xbit_r54_c173 bl[173] br[173] wl[54] vdd gnd cell_6t
Xbit_r55_c173 bl[173] br[173] wl[55] vdd gnd cell_6t
Xbit_r56_c173 bl[173] br[173] wl[56] vdd gnd cell_6t
Xbit_r57_c173 bl[173] br[173] wl[57] vdd gnd cell_6t
Xbit_r58_c173 bl[173] br[173] wl[58] vdd gnd cell_6t
Xbit_r59_c173 bl[173] br[173] wl[59] vdd gnd cell_6t
Xbit_r60_c173 bl[173] br[173] wl[60] vdd gnd cell_6t
Xbit_r61_c173 bl[173] br[173] wl[61] vdd gnd cell_6t
Xbit_r62_c173 bl[173] br[173] wl[62] vdd gnd cell_6t
Xbit_r63_c173 bl[173] br[173] wl[63] vdd gnd cell_6t
Xbit_r64_c173 bl[173] br[173] wl[64] vdd gnd cell_6t
Xbit_r65_c173 bl[173] br[173] wl[65] vdd gnd cell_6t
Xbit_r66_c173 bl[173] br[173] wl[66] vdd gnd cell_6t
Xbit_r67_c173 bl[173] br[173] wl[67] vdd gnd cell_6t
Xbit_r68_c173 bl[173] br[173] wl[68] vdd gnd cell_6t
Xbit_r69_c173 bl[173] br[173] wl[69] vdd gnd cell_6t
Xbit_r70_c173 bl[173] br[173] wl[70] vdd gnd cell_6t
Xbit_r71_c173 bl[173] br[173] wl[71] vdd gnd cell_6t
Xbit_r72_c173 bl[173] br[173] wl[72] vdd gnd cell_6t
Xbit_r73_c173 bl[173] br[173] wl[73] vdd gnd cell_6t
Xbit_r74_c173 bl[173] br[173] wl[74] vdd gnd cell_6t
Xbit_r75_c173 bl[173] br[173] wl[75] vdd gnd cell_6t
Xbit_r76_c173 bl[173] br[173] wl[76] vdd gnd cell_6t
Xbit_r77_c173 bl[173] br[173] wl[77] vdd gnd cell_6t
Xbit_r78_c173 bl[173] br[173] wl[78] vdd gnd cell_6t
Xbit_r79_c173 bl[173] br[173] wl[79] vdd gnd cell_6t
Xbit_r80_c173 bl[173] br[173] wl[80] vdd gnd cell_6t
Xbit_r81_c173 bl[173] br[173] wl[81] vdd gnd cell_6t
Xbit_r82_c173 bl[173] br[173] wl[82] vdd gnd cell_6t
Xbit_r83_c173 bl[173] br[173] wl[83] vdd gnd cell_6t
Xbit_r84_c173 bl[173] br[173] wl[84] vdd gnd cell_6t
Xbit_r85_c173 bl[173] br[173] wl[85] vdd gnd cell_6t
Xbit_r86_c173 bl[173] br[173] wl[86] vdd gnd cell_6t
Xbit_r87_c173 bl[173] br[173] wl[87] vdd gnd cell_6t
Xbit_r88_c173 bl[173] br[173] wl[88] vdd gnd cell_6t
Xbit_r89_c173 bl[173] br[173] wl[89] vdd gnd cell_6t
Xbit_r90_c173 bl[173] br[173] wl[90] vdd gnd cell_6t
Xbit_r91_c173 bl[173] br[173] wl[91] vdd gnd cell_6t
Xbit_r92_c173 bl[173] br[173] wl[92] vdd gnd cell_6t
Xbit_r93_c173 bl[173] br[173] wl[93] vdd gnd cell_6t
Xbit_r94_c173 bl[173] br[173] wl[94] vdd gnd cell_6t
Xbit_r95_c173 bl[173] br[173] wl[95] vdd gnd cell_6t
Xbit_r96_c173 bl[173] br[173] wl[96] vdd gnd cell_6t
Xbit_r97_c173 bl[173] br[173] wl[97] vdd gnd cell_6t
Xbit_r98_c173 bl[173] br[173] wl[98] vdd gnd cell_6t
Xbit_r99_c173 bl[173] br[173] wl[99] vdd gnd cell_6t
Xbit_r100_c173 bl[173] br[173] wl[100] vdd gnd cell_6t
Xbit_r101_c173 bl[173] br[173] wl[101] vdd gnd cell_6t
Xbit_r102_c173 bl[173] br[173] wl[102] vdd gnd cell_6t
Xbit_r103_c173 bl[173] br[173] wl[103] vdd gnd cell_6t
Xbit_r104_c173 bl[173] br[173] wl[104] vdd gnd cell_6t
Xbit_r105_c173 bl[173] br[173] wl[105] vdd gnd cell_6t
Xbit_r106_c173 bl[173] br[173] wl[106] vdd gnd cell_6t
Xbit_r107_c173 bl[173] br[173] wl[107] vdd gnd cell_6t
Xbit_r108_c173 bl[173] br[173] wl[108] vdd gnd cell_6t
Xbit_r109_c173 bl[173] br[173] wl[109] vdd gnd cell_6t
Xbit_r110_c173 bl[173] br[173] wl[110] vdd gnd cell_6t
Xbit_r111_c173 bl[173] br[173] wl[111] vdd gnd cell_6t
Xbit_r112_c173 bl[173] br[173] wl[112] vdd gnd cell_6t
Xbit_r113_c173 bl[173] br[173] wl[113] vdd gnd cell_6t
Xbit_r114_c173 bl[173] br[173] wl[114] vdd gnd cell_6t
Xbit_r115_c173 bl[173] br[173] wl[115] vdd gnd cell_6t
Xbit_r116_c173 bl[173] br[173] wl[116] vdd gnd cell_6t
Xbit_r117_c173 bl[173] br[173] wl[117] vdd gnd cell_6t
Xbit_r118_c173 bl[173] br[173] wl[118] vdd gnd cell_6t
Xbit_r119_c173 bl[173] br[173] wl[119] vdd gnd cell_6t
Xbit_r120_c173 bl[173] br[173] wl[120] vdd gnd cell_6t
Xbit_r121_c173 bl[173] br[173] wl[121] vdd gnd cell_6t
Xbit_r122_c173 bl[173] br[173] wl[122] vdd gnd cell_6t
Xbit_r123_c173 bl[173] br[173] wl[123] vdd gnd cell_6t
Xbit_r124_c173 bl[173] br[173] wl[124] vdd gnd cell_6t
Xbit_r125_c173 bl[173] br[173] wl[125] vdd gnd cell_6t
Xbit_r126_c173 bl[173] br[173] wl[126] vdd gnd cell_6t
Xbit_r127_c173 bl[173] br[173] wl[127] vdd gnd cell_6t
Xbit_r128_c173 bl[173] br[173] wl[128] vdd gnd cell_6t
Xbit_r129_c173 bl[173] br[173] wl[129] vdd gnd cell_6t
Xbit_r130_c173 bl[173] br[173] wl[130] vdd gnd cell_6t
Xbit_r131_c173 bl[173] br[173] wl[131] vdd gnd cell_6t
Xbit_r132_c173 bl[173] br[173] wl[132] vdd gnd cell_6t
Xbit_r133_c173 bl[173] br[173] wl[133] vdd gnd cell_6t
Xbit_r134_c173 bl[173] br[173] wl[134] vdd gnd cell_6t
Xbit_r135_c173 bl[173] br[173] wl[135] vdd gnd cell_6t
Xbit_r136_c173 bl[173] br[173] wl[136] vdd gnd cell_6t
Xbit_r137_c173 bl[173] br[173] wl[137] vdd gnd cell_6t
Xbit_r138_c173 bl[173] br[173] wl[138] vdd gnd cell_6t
Xbit_r139_c173 bl[173] br[173] wl[139] vdd gnd cell_6t
Xbit_r140_c173 bl[173] br[173] wl[140] vdd gnd cell_6t
Xbit_r141_c173 bl[173] br[173] wl[141] vdd gnd cell_6t
Xbit_r142_c173 bl[173] br[173] wl[142] vdd gnd cell_6t
Xbit_r143_c173 bl[173] br[173] wl[143] vdd gnd cell_6t
Xbit_r144_c173 bl[173] br[173] wl[144] vdd gnd cell_6t
Xbit_r145_c173 bl[173] br[173] wl[145] vdd gnd cell_6t
Xbit_r146_c173 bl[173] br[173] wl[146] vdd gnd cell_6t
Xbit_r147_c173 bl[173] br[173] wl[147] vdd gnd cell_6t
Xbit_r148_c173 bl[173] br[173] wl[148] vdd gnd cell_6t
Xbit_r149_c173 bl[173] br[173] wl[149] vdd gnd cell_6t
Xbit_r150_c173 bl[173] br[173] wl[150] vdd gnd cell_6t
Xbit_r151_c173 bl[173] br[173] wl[151] vdd gnd cell_6t
Xbit_r152_c173 bl[173] br[173] wl[152] vdd gnd cell_6t
Xbit_r153_c173 bl[173] br[173] wl[153] vdd gnd cell_6t
Xbit_r154_c173 bl[173] br[173] wl[154] vdd gnd cell_6t
Xbit_r155_c173 bl[173] br[173] wl[155] vdd gnd cell_6t
Xbit_r156_c173 bl[173] br[173] wl[156] vdd gnd cell_6t
Xbit_r157_c173 bl[173] br[173] wl[157] vdd gnd cell_6t
Xbit_r158_c173 bl[173] br[173] wl[158] vdd gnd cell_6t
Xbit_r159_c173 bl[173] br[173] wl[159] vdd gnd cell_6t
Xbit_r160_c173 bl[173] br[173] wl[160] vdd gnd cell_6t
Xbit_r161_c173 bl[173] br[173] wl[161] vdd gnd cell_6t
Xbit_r162_c173 bl[173] br[173] wl[162] vdd gnd cell_6t
Xbit_r163_c173 bl[173] br[173] wl[163] vdd gnd cell_6t
Xbit_r164_c173 bl[173] br[173] wl[164] vdd gnd cell_6t
Xbit_r165_c173 bl[173] br[173] wl[165] vdd gnd cell_6t
Xbit_r166_c173 bl[173] br[173] wl[166] vdd gnd cell_6t
Xbit_r167_c173 bl[173] br[173] wl[167] vdd gnd cell_6t
Xbit_r168_c173 bl[173] br[173] wl[168] vdd gnd cell_6t
Xbit_r169_c173 bl[173] br[173] wl[169] vdd gnd cell_6t
Xbit_r170_c173 bl[173] br[173] wl[170] vdd gnd cell_6t
Xbit_r171_c173 bl[173] br[173] wl[171] vdd gnd cell_6t
Xbit_r172_c173 bl[173] br[173] wl[172] vdd gnd cell_6t
Xbit_r173_c173 bl[173] br[173] wl[173] vdd gnd cell_6t
Xbit_r174_c173 bl[173] br[173] wl[174] vdd gnd cell_6t
Xbit_r175_c173 bl[173] br[173] wl[175] vdd gnd cell_6t
Xbit_r176_c173 bl[173] br[173] wl[176] vdd gnd cell_6t
Xbit_r177_c173 bl[173] br[173] wl[177] vdd gnd cell_6t
Xbit_r178_c173 bl[173] br[173] wl[178] vdd gnd cell_6t
Xbit_r179_c173 bl[173] br[173] wl[179] vdd gnd cell_6t
Xbit_r180_c173 bl[173] br[173] wl[180] vdd gnd cell_6t
Xbit_r181_c173 bl[173] br[173] wl[181] vdd gnd cell_6t
Xbit_r182_c173 bl[173] br[173] wl[182] vdd gnd cell_6t
Xbit_r183_c173 bl[173] br[173] wl[183] vdd gnd cell_6t
Xbit_r184_c173 bl[173] br[173] wl[184] vdd gnd cell_6t
Xbit_r185_c173 bl[173] br[173] wl[185] vdd gnd cell_6t
Xbit_r186_c173 bl[173] br[173] wl[186] vdd gnd cell_6t
Xbit_r187_c173 bl[173] br[173] wl[187] vdd gnd cell_6t
Xbit_r188_c173 bl[173] br[173] wl[188] vdd gnd cell_6t
Xbit_r189_c173 bl[173] br[173] wl[189] vdd gnd cell_6t
Xbit_r190_c173 bl[173] br[173] wl[190] vdd gnd cell_6t
Xbit_r191_c173 bl[173] br[173] wl[191] vdd gnd cell_6t
Xbit_r192_c173 bl[173] br[173] wl[192] vdd gnd cell_6t
Xbit_r193_c173 bl[173] br[173] wl[193] vdd gnd cell_6t
Xbit_r194_c173 bl[173] br[173] wl[194] vdd gnd cell_6t
Xbit_r195_c173 bl[173] br[173] wl[195] vdd gnd cell_6t
Xbit_r196_c173 bl[173] br[173] wl[196] vdd gnd cell_6t
Xbit_r197_c173 bl[173] br[173] wl[197] vdd gnd cell_6t
Xbit_r198_c173 bl[173] br[173] wl[198] vdd gnd cell_6t
Xbit_r199_c173 bl[173] br[173] wl[199] vdd gnd cell_6t
Xbit_r200_c173 bl[173] br[173] wl[200] vdd gnd cell_6t
Xbit_r201_c173 bl[173] br[173] wl[201] vdd gnd cell_6t
Xbit_r202_c173 bl[173] br[173] wl[202] vdd gnd cell_6t
Xbit_r203_c173 bl[173] br[173] wl[203] vdd gnd cell_6t
Xbit_r204_c173 bl[173] br[173] wl[204] vdd gnd cell_6t
Xbit_r205_c173 bl[173] br[173] wl[205] vdd gnd cell_6t
Xbit_r206_c173 bl[173] br[173] wl[206] vdd gnd cell_6t
Xbit_r207_c173 bl[173] br[173] wl[207] vdd gnd cell_6t
Xbit_r208_c173 bl[173] br[173] wl[208] vdd gnd cell_6t
Xbit_r209_c173 bl[173] br[173] wl[209] vdd gnd cell_6t
Xbit_r210_c173 bl[173] br[173] wl[210] vdd gnd cell_6t
Xbit_r211_c173 bl[173] br[173] wl[211] vdd gnd cell_6t
Xbit_r212_c173 bl[173] br[173] wl[212] vdd gnd cell_6t
Xbit_r213_c173 bl[173] br[173] wl[213] vdd gnd cell_6t
Xbit_r214_c173 bl[173] br[173] wl[214] vdd gnd cell_6t
Xbit_r215_c173 bl[173] br[173] wl[215] vdd gnd cell_6t
Xbit_r216_c173 bl[173] br[173] wl[216] vdd gnd cell_6t
Xbit_r217_c173 bl[173] br[173] wl[217] vdd gnd cell_6t
Xbit_r218_c173 bl[173] br[173] wl[218] vdd gnd cell_6t
Xbit_r219_c173 bl[173] br[173] wl[219] vdd gnd cell_6t
Xbit_r220_c173 bl[173] br[173] wl[220] vdd gnd cell_6t
Xbit_r221_c173 bl[173] br[173] wl[221] vdd gnd cell_6t
Xbit_r222_c173 bl[173] br[173] wl[222] vdd gnd cell_6t
Xbit_r223_c173 bl[173] br[173] wl[223] vdd gnd cell_6t
Xbit_r224_c173 bl[173] br[173] wl[224] vdd gnd cell_6t
Xbit_r225_c173 bl[173] br[173] wl[225] vdd gnd cell_6t
Xbit_r226_c173 bl[173] br[173] wl[226] vdd gnd cell_6t
Xbit_r227_c173 bl[173] br[173] wl[227] vdd gnd cell_6t
Xbit_r228_c173 bl[173] br[173] wl[228] vdd gnd cell_6t
Xbit_r229_c173 bl[173] br[173] wl[229] vdd gnd cell_6t
Xbit_r230_c173 bl[173] br[173] wl[230] vdd gnd cell_6t
Xbit_r231_c173 bl[173] br[173] wl[231] vdd gnd cell_6t
Xbit_r232_c173 bl[173] br[173] wl[232] vdd gnd cell_6t
Xbit_r233_c173 bl[173] br[173] wl[233] vdd gnd cell_6t
Xbit_r234_c173 bl[173] br[173] wl[234] vdd gnd cell_6t
Xbit_r235_c173 bl[173] br[173] wl[235] vdd gnd cell_6t
Xbit_r236_c173 bl[173] br[173] wl[236] vdd gnd cell_6t
Xbit_r237_c173 bl[173] br[173] wl[237] vdd gnd cell_6t
Xbit_r238_c173 bl[173] br[173] wl[238] vdd gnd cell_6t
Xbit_r239_c173 bl[173] br[173] wl[239] vdd gnd cell_6t
Xbit_r240_c173 bl[173] br[173] wl[240] vdd gnd cell_6t
Xbit_r241_c173 bl[173] br[173] wl[241] vdd gnd cell_6t
Xbit_r242_c173 bl[173] br[173] wl[242] vdd gnd cell_6t
Xbit_r243_c173 bl[173] br[173] wl[243] vdd gnd cell_6t
Xbit_r244_c173 bl[173] br[173] wl[244] vdd gnd cell_6t
Xbit_r245_c173 bl[173] br[173] wl[245] vdd gnd cell_6t
Xbit_r246_c173 bl[173] br[173] wl[246] vdd gnd cell_6t
Xbit_r247_c173 bl[173] br[173] wl[247] vdd gnd cell_6t
Xbit_r248_c173 bl[173] br[173] wl[248] vdd gnd cell_6t
Xbit_r249_c173 bl[173] br[173] wl[249] vdd gnd cell_6t
Xbit_r250_c173 bl[173] br[173] wl[250] vdd gnd cell_6t
Xbit_r251_c173 bl[173] br[173] wl[251] vdd gnd cell_6t
Xbit_r252_c173 bl[173] br[173] wl[252] vdd gnd cell_6t
Xbit_r253_c173 bl[173] br[173] wl[253] vdd gnd cell_6t
Xbit_r254_c173 bl[173] br[173] wl[254] vdd gnd cell_6t
Xbit_r255_c173 bl[173] br[173] wl[255] vdd gnd cell_6t
Xbit_r0_c174 bl[174] br[174] wl[0] vdd gnd cell_6t
Xbit_r1_c174 bl[174] br[174] wl[1] vdd gnd cell_6t
Xbit_r2_c174 bl[174] br[174] wl[2] vdd gnd cell_6t
Xbit_r3_c174 bl[174] br[174] wl[3] vdd gnd cell_6t
Xbit_r4_c174 bl[174] br[174] wl[4] vdd gnd cell_6t
Xbit_r5_c174 bl[174] br[174] wl[5] vdd gnd cell_6t
Xbit_r6_c174 bl[174] br[174] wl[6] vdd gnd cell_6t
Xbit_r7_c174 bl[174] br[174] wl[7] vdd gnd cell_6t
Xbit_r8_c174 bl[174] br[174] wl[8] vdd gnd cell_6t
Xbit_r9_c174 bl[174] br[174] wl[9] vdd gnd cell_6t
Xbit_r10_c174 bl[174] br[174] wl[10] vdd gnd cell_6t
Xbit_r11_c174 bl[174] br[174] wl[11] vdd gnd cell_6t
Xbit_r12_c174 bl[174] br[174] wl[12] vdd gnd cell_6t
Xbit_r13_c174 bl[174] br[174] wl[13] vdd gnd cell_6t
Xbit_r14_c174 bl[174] br[174] wl[14] vdd gnd cell_6t
Xbit_r15_c174 bl[174] br[174] wl[15] vdd gnd cell_6t
Xbit_r16_c174 bl[174] br[174] wl[16] vdd gnd cell_6t
Xbit_r17_c174 bl[174] br[174] wl[17] vdd gnd cell_6t
Xbit_r18_c174 bl[174] br[174] wl[18] vdd gnd cell_6t
Xbit_r19_c174 bl[174] br[174] wl[19] vdd gnd cell_6t
Xbit_r20_c174 bl[174] br[174] wl[20] vdd gnd cell_6t
Xbit_r21_c174 bl[174] br[174] wl[21] vdd gnd cell_6t
Xbit_r22_c174 bl[174] br[174] wl[22] vdd gnd cell_6t
Xbit_r23_c174 bl[174] br[174] wl[23] vdd gnd cell_6t
Xbit_r24_c174 bl[174] br[174] wl[24] vdd gnd cell_6t
Xbit_r25_c174 bl[174] br[174] wl[25] vdd gnd cell_6t
Xbit_r26_c174 bl[174] br[174] wl[26] vdd gnd cell_6t
Xbit_r27_c174 bl[174] br[174] wl[27] vdd gnd cell_6t
Xbit_r28_c174 bl[174] br[174] wl[28] vdd gnd cell_6t
Xbit_r29_c174 bl[174] br[174] wl[29] vdd gnd cell_6t
Xbit_r30_c174 bl[174] br[174] wl[30] vdd gnd cell_6t
Xbit_r31_c174 bl[174] br[174] wl[31] vdd gnd cell_6t
Xbit_r32_c174 bl[174] br[174] wl[32] vdd gnd cell_6t
Xbit_r33_c174 bl[174] br[174] wl[33] vdd gnd cell_6t
Xbit_r34_c174 bl[174] br[174] wl[34] vdd gnd cell_6t
Xbit_r35_c174 bl[174] br[174] wl[35] vdd gnd cell_6t
Xbit_r36_c174 bl[174] br[174] wl[36] vdd gnd cell_6t
Xbit_r37_c174 bl[174] br[174] wl[37] vdd gnd cell_6t
Xbit_r38_c174 bl[174] br[174] wl[38] vdd gnd cell_6t
Xbit_r39_c174 bl[174] br[174] wl[39] vdd gnd cell_6t
Xbit_r40_c174 bl[174] br[174] wl[40] vdd gnd cell_6t
Xbit_r41_c174 bl[174] br[174] wl[41] vdd gnd cell_6t
Xbit_r42_c174 bl[174] br[174] wl[42] vdd gnd cell_6t
Xbit_r43_c174 bl[174] br[174] wl[43] vdd gnd cell_6t
Xbit_r44_c174 bl[174] br[174] wl[44] vdd gnd cell_6t
Xbit_r45_c174 bl[174] br[174] wl[45] vdd gnd cell_6t
Xbit_r46_c174 bl[174] br[174] wl[46] vdd gnd cell_6t
Xbit_r47_c174 bl[174] br[174] wl[47] vdd gnd cell_6t
Xbit_r48_c174 bl[174] br[174] wl[48] vdd gnd cell_6t
Xbit_r49_c174 bl[174] br[174] wl[49] vdd gnd cell_6t
Xbit_r50_c174 bl[174] br[174] wl[50] vdd gnd cell_6t
Xbit_r51_c174 bl[174] br[174] wl[51] vdd gnd cell_6t
Xbit_r52_c174 bl[174] br[174] wl[52] vdd gnd cell_6t
Xbit_r53_c174 bl[174] br[174] wl[53] vdd gnd cell_6t
Xbit_r54_c174 bl[174] br[174] wl[54] vdd gnd cell_6t
Xbit_r55_c174 bl[174] br[174] wl[55] vdd gnd cell_6t
Xbit_r56_c174 bl[174] br[174] wl[56] vdd gnd cell_6t
Xbit_r57_c174 bl[174] br[174] wl[57] vdd gnd cell_6t
Xbit_r58_c174 bl[174] br[174] wl[58] vdd gnd cell_6t
Xbit_r59_c174 bl[174] br[174] wl[59] vdd gnd cell_6t
Xbit_r60_c174 bl[174] br[174] wl[60] vdd gnd cell_6t
Xbit_r61_c174 bl[174] br[174] wl[61] vdd gnd cell_6t
Xbit_r62_c174 bl[174] br[174] wl[62] vdd gnd cell_6t
Xbit_r63_c174 bl[174] br[174] wl[63] vdd gnd cell_6t
Xbit_r64_c174 bl[174] br[174] wl[64] vdd gnd cell_6t
Xbit_r65_c174 bl[174] br[174] wl[65] vdd gnd cell_6t
Xbit_r66_c174 bl[174] br[174] wl[66] vdd gnd cell_6t
Xbit_r67_c174 bl[174] br[174] wl[67] vdd gnd cell_6t
Xbit_r68_c174 bl[174] br[174] wl[68] vdd gnd cell_6t
Xbit_r69_c174 bl[174] br[174] wl[69] vdd gnd cell_6t
Xbit_r70_c174 bl[174] br[174] wl[70] vdd gnd cell_6t
Xbit_r71_c174 bl[174] br[174] wl[71] vdd gnd cell_6t
Xbit_r72_c174 bl[174] br[174] wl[72] vdd gnd cell_6t
Xbit_r73_c174 bl[174] br[174] wl[73] vdd gnd cell_6t
Xbit_r74_c174 bl[174] br[174] wl[74] vdd gnd cell_6t
Xbit_r75_c174 bl[174] br[174] wl[75] vdd gnd cell_6t
Xbit_r76_c174 bl[174] br[174] wl[76] vdd gnd cell_6t
Xbit_r77_c174 bl[174] br[174] wl[77] vdd gnd cell_6t
Xbit_r78_c174 bl[174] br[174] wl[78] vdd gnd cell_6t
Xbit_r79_c174 bl[174] br[174] wl[79] vdd gnd cell_6t
Xbit_r80_c174 bl[174] br[174] wl[80] vdd gnd cell_6t
Xbit_r81_c174 bl[174] br[174] wl[81] vdd gnd cell_6t
Xbit_r82_c174 bl[174] br[174] wl[82] vdd gnd cell_6t
Xbit_r83_c174 bl[174] br[174] wl[83] vdd gnd cell_6t
Xbit_r84_c174 bl[174] br[174] wl[84] vdd gnd cell_6t
Xbit_r85_c174 bl[174] br[174] wl[85] vdd gnd cell_6t
Xbit_r86_c174 bl[174] br[174] wl[86] vdd gnd cell_6t
Xbit_r87_c174 bl[174] br[174] wl[87] vdd gnd cell_6t
Xbit_r88_c174 bl[174] br[174] wl[88] vdd gnd cell_6t
Xbit_r89_c174 bl[174] br[174] wl[89] vdd gnd cell_6t
Xbit_r90_c174 bl[174] br[174] wl[90] vdd gnd cell_6t
Xbit_r91_c174 bl[174] br[174] wl[91] vdd gnd cell_6t
Xbit_r92_c174 bl[174] br[174] wl[92] vdd gnd cell_6t
Xbit_r93_c174 bl[174] br[174] wl[93] vdd gnd cell_6t
Xbit_r94_c174 bl[174] br[174] wl[94] vdd gnd cell_6t
Xbit_r95_c174 bl[174] br[174] wl[95] vdd gnd cell_6t
Xbit_r96_c174 bl[174] br[174] wl[96] vdd gnd cell_6t
Xbit_r97_c174 bl[174] br[174] wl[97] vdd gnd cell_6t
Xbit_r98_c174 bl[174] br[174] wl[98] vdd gnd cell_6t
Xbit_r99_c174 bl[174] br[174] wl[99] vdd gnd cell_6t
Xbit_r100_c174 bl[174] br[174] wl[100] vdd gnd cell_6t
Xbit_r101_c174 bl[174] br[174] wl[101] vdd gnd cell_6t
Xbit_r102_c174 bl[174] br[174] wl[102] vdd gnd cell_6t
Xbit_r103_c174 bl[174] br[174] wl[103] vdd gnd cell_6t
Xbit_r104_c174 bl[174] br[174] wl[104] vdd gnd cell_6t
Xbit_r105_c174 bl[174] br[174] wl[105] vdd gnd cell_6t
Xbit_r106_c174 bl[174] br[174] wl[106] vdd gnd cell_6t
Xbit_r107_c174 bl[174] br[174] wl[107] vdd gnd cell_6t
Xbit_r108_c174 bl[174] br[174] wl[108] vdd gnd cell_6t
Xbit_r109_c174 bl[174] br[174] wl[109] vdd gnd cell_6t
Xbit_r110_c174 bl[174] br[174] wl[110] vdd gnd cell_6t
Xbit_r111_c174 bl[174] br[174] wl[111] vdd gnd cell_6t
Xbit_r112_c174 bl[174] br[174] wl[112] vdd gnd cell_6t
Xbit_r113_c174 bl[174] br[174] wl[113] vdd gnd cell_6t
Xbit_r114_c174 bl[174] br[174] wl[114] vdd gnd cell_6t
Xbit_r115_c174 bl[174] br[174] wl[115] vdd gnd cell_6t
Xbit_r116_c174 bl[174] br[174] wl[116] vdd gnd cell_6t
Xbit_r117_c174 bl[174] br[174] wl[117] vdd gnd cell_6t
Xbit_r118_c174 bl[174] br[174] wl[118] vdd gnd cell_6t
Xbit_r119_c174 bl[174] br[174] wl[119] vdd gnd cell_6t
Xbit_r120_c174 bl[174] br[174] wl[120] vdd gnd cell_6t
Xbit_r121_c174 bl[174] br[174] wl[121] vdd gnd cell_6t
Xbit_r122_c174 bl[174] br[174] wl[122] vdd gnd cell_6t
Xbit_r123_c174 bl[174] br[174] wl[123] vdd gnd cell_6t
Xbit_r124_c174 bl[174] br[174] wl[124] vdd gnd cell_6t
Xbit_r125_c174 bl[174] br[174] wl[125] vdd gnd cell_6t
Xbit_r126_c174 bl[174] br[174] wl[126] vdd gnd cell_6t
Xbit_r127_c174 bl[174] br[174] wl[127] vdd gnd cell_6t
Xbit_r128_c174 bl[174] br[174] wl[128] vdd gnd cell_6t
Xbit_r129_c174 bl[174] br[174] wl[129] vdd gnd cell_6t
Xbit_r130_c174 bl[174] br[174] wl[130] vdd gnd cell_6t
Xbit_r131_c174 bl[174] br[174] wl[131] vdd gnd cell_6t
Xbit_r132_c174 bl[174] br[174] wl[132] vdd gnd cell_6t
Xbit_r133_c174 bl[174] br[174] wl[133] vdd gnd cell_6t
Xbit_r134_c174 bl[174] br[174] wl[134] vdd gnd cell_6t
Xbit_r135_c174 bl[174] br[174] wl[135] vdd gnd cell_6t
Xbit_r136_c174 bl[174] br[174] wl[136] vdd gnd cell_6t
Xbit_r137_c174 bl[174] br[174] wl[137] vdd gnd cell_6t
Xbit_r138_c174 bl[174] br[174] wl[138] vdd gnd cell_6t
Xbit_r139_c174 bl[174] br[174] wl[139] vdd gnd cell_6t
Xbit_r140_c174 bl[174] br[174] wl[140] vdd gnd cell_6t
Xbit_r141_c174 bl[174] br[174] wl[141] vdd gnd cell_6t
Xbit_r142_c174 bl[174] br[174] wl[142] vdd gnd cell_6t
Xbit_r143_c174 bl[174] br[174] wl[143] vdd gnd cell_6t
Xbit_r144_c174 bl[174] br[174] wl[144] vdd gnd cell_6t
Xbit_r145_c174 bl[174] br[174] wl[145] vdd gnd cell_6t
Xbit_r146_c174 bl[174] br[174] wl[146] vdd gnd cell_6t
Xbit_r147_c174 bl[174] br[174] wl[147] vdd gnd cell_6t
Xbit_r148_c174 bl[174] br[174] wl[148] vdd gnd cell_6t
Xbit_r149_c174 bl[174] br[174] wl[149] vdd gnd cell_6t
Xbit_r150_c174 bl[174] br[174] wl[150] vdd gnd cell_6t
Xbit_r151_c174 bl[174] br[174] wl[151] vdd gnd cell_6t
Xbit_r152_c174 bl[174] br[174] wl[152] vdd gnd cell_6t
Xbit_r153_c174 bl[174] br[174] wl[153] vdd gnd cell_6t
Xbit_r154_c174 bl[174] br[174] wl[154] vdd gnd cell_6t
Xbit_r155_c174 bl[174] br[174] wl[155] vdd gnd cell_6t
Xbit_r156_c174 bl[174] br[174] wl[156] vdd gnd cell_6t
Xbit_r157_c174 bl[174] br[174] wl[157] vdd gnd cell_6t
Xbit_r158_c174 bl[174] br[174] wl[158] vdd gnd cell_6t
Xbit_r159_c174 bl[174] br[174] wl[159] vdd gnd cell_6t
Xbit_r160_c174 bl[174] br[174] wl[160] vdd gnd cell_6t
Xbit_r161_c174 bl[174] br[174] wl[161] vdd gnd cell_6t
Xbit_r162_c174 bl[174] br[174] wl[162] vdd gnd cell_6t
Xbit_r163_c174 bl[174] br[174] wl[163] vdd gnd cell_6t
Xbit_r164_c174 bl[174] br[174] wl[164] vdd gnd cell_6t
Xbit_r165_c174 bl[174] br[174] wl[165] vdd gnd cell_6t
Xbit_r166_c174 bl[174] br[174] wl[166] vdd gnd cell_6t
Xbit_r167_c174 bl[174] br[174] wl[167] vdd gnd cell_6t
Xbit_r168_c174 bl[174] br[174] wl[168] vdd gnd cell_6t
Xbit_r169_c174 bl[174] br[174] wl[169] vdd gnd cell_6t
Xbit_r170_c174 bl[174] br[174] wl[170] vdd gnd cell_6t
Xbit_r171_c174 bl[174] br[174] wl[171] vdd gnd cell_6t
Xbit_r172_c174 bl[174] br[174] wl[172] vdd gnd cell_6t
Xbit_r173_c174 bl[174] br[174] wl[173] vdd gnd cell_6t
Xbit_r174_c174 bl[174] br[174] wl[174] vdd gnd cell_6t
Xbit_r175_c174 bl[174] br[174] wl[175] vdd gnd cell_6t
Xbit_r176_c174 bl[174] br[174] wl[176] vdd gnd cell_6t
Xbit_r177_c174 bl[174] br[174] wl[177] vdd gnd cell_6t
Xbit_r178_c174 bl[174] br[174] wl[178] vdd gnd cell_6t
Xbit_r179_c174 bl[174] br[174] wl[179] vdd gnd cell_6t
Xbit_r180_c174 bl[174] br[174] wl[180] vdd gnd cell_6t
Xbit_r181_c174 bl[174] br[174] wl[181] vdd gnd cell_6t
Xbit_r182_c174 bl[174] br[174] wl[182] vdd gnd cell_6t
Xbit_r183_c174 bl[174] br[174] wl[183] vdd gnd cell_6t
Xbit_r184_c174 bl[174] br[174] wl[184] vdd gnd cell_6t
Xbit_r185_c174 bl[174] br[174] wl[185] vdd gnd cell_6t
Xbit_r186_c174 bl[174] br[174] wl[186] vdd gnd cell_6t
Xbit_r187_c174 bl[174] br[174] wl[187] vdd gnd cell_6t
Xbit_r188_c174 bl[174] br[174] wl[188] vdd gnd cell_6t
Xbit_r189_c174 bl[174] br[174] wl[189] vdd gnd cell_6t
Xbit_r190_c174 bl[174] br[174] wl[190] vdd gnd cell_6t
Xbit_r191_c174 bl[174] br[174] wl[191] vdd gnd cell_6t
Xbit_r192_c174 bl[174] br[174] wl[192] vdd gnd cell_6t
Xbit_r193_c174 bl[174] br[174] wl[193] vdd gnd cell_6t
Xbit_r194_c174 bl[174] br[174] wl[194] vdd gnd cell_6t
Xbit_r195_c174 bl[174] br[174] wl[195] vdd gnd cell_6t
Xbit_r196_c174 bl[174] br[174] wl[196] vdd gnd cell_6t
Xbit_r197_c174 bl[174] br[174] wl[197] vdd gnd cell_6t
Xbit_r198_c174 bl[174] br[174] wl[198] vdd gnd cell_6t
Xbit_r199_c174 bl[174] br[174] wl[199] vdd gnd cell_6t
Xbit_r200_c174 bl[174] br[174] wl[200] vdd gnd cell_6t
Xbit_r201_c174 bl[174] br[174] wl[201] vdd gnd cell_6t
Xbit_r202_c174 bl[174] br[174] wl[202] vdd gnd cell_6t
Xbit_r203_c174 bl[174] br[174] wl[203] vdd gnd cell_6t
Xbit_r204_c174 bl[174] br[174] wl[204] vdd gnd cell_6t
Xbit_r205_c174 bl[174] br[174] wl[205] vdd gnd cell_6t
Xbit_r206_c174 bl[174] br[174] wl[206] vdd gnd cell_6t
Xbit_r207_c174 bl[174] br[174] wl[207] vdd gnd cell_6t
Xbit_r208_c174 bl[174] br[174] wl[208] vdd gnd cell_6t
Xbit_r209_c174 bl[174] br[174] wl[209] vdd gnd cell_6t
Xbit_r210_c174 bl[174] br[174] wl[210] vdd gnd cell_6t
Xbit_r211_c174 bl[174] br[174] wl[211] vdd gnd cell_6t
Xbit_r212_c174 bl[174] br[174] wl[212] vdd gnd cell_6t
Xbit_r213_c174 bl[174] br[174] wl[213] vdd gnd cell_6t
Xbit_r214_c174 bl[174] br[174] wl[214] vdd gnd cell_6t
Xbit_r215_c174 bl[174] br[174] wl[215] vdd gnd cell_6t
Xbit_r216_c174 bl[174] br[174] wl[216] vdd gnd cell_6t
Xbit_r217_c174 bl[174] br[174] wl[217] vdd gnd cell_6t
Xbit_r218_c174 bl[174] br[174] wl[218] vdd gnd cell_6t
Xbit_r219_c174 bl[174] br[174] wl[219] vdd gnd cell_6t
Xbit_r220_c174 bl[174] br[174] wl[220] vdd gnd cell_6t
Xbit_r221_c174 bl[174] br[174] wl[221] vdd gnd cell_6t
Xbit_r222_c174 bl[174] br[174] wl[222] vdd gnd cell_6t
Xbit_r223_c174 bl[174] br[174] wl[223] vdd gnd cell_6t
Xbit_r224_c174 bl[174] br[174] wl[224] vdd gnd cell_6t
Xbit_r225_c174 bl[174] br[174] wl[225] vdd gnd cell_6t
Xbit_r226_c174 bl[174] br[174] wl[226] vdd gnd cell_6t
Xbit_r227_c174 bl[174] br[174] wl[227] vdd gnd cell_6t
Xbit_r228_c174 bl[174] br[174] wl[228] vdd gnd cell_6t
Xbit_r229_c174 bl[174] br[174] wl[229] vdd gnd cell_6t
Xbit_r230_c174 bl[174] br[174] wl[230] vdd gnd cell_6t
Xbit_r231_c174 bl[174] br[174] wl[231] vdd gnd cell_6t
Xbit_r232_c174 bl[174] br[174] wl[232] vdd gnd cell_6t
Xbit_r233_c174 bl[174] br[174] wl[233] vdd gnd cell_6t
Xbit_r234_c174 bl[174] br[174] wl[234] vdd gnd cell_6t
Xbit_r235_c174 bl[174] br[174] wl[235] vdd gnd cell_6t
Xbit_r236_c174 bl[174] br[174] wl[236] vdd gnd cell_6t
Xbit_r237_c174 bl[174] br[174] wl[237] vdd gnd cell_6t
Xbit_r238_c174 bl[174] br[174] wl[238] vdd gnd cell_6t
Xbit_r239_c174 bl[174] br[174] wl[239] vdd gnd cell_6t
Xbit_r240_c174 bl[174] br[174] wl[240] vdd gnd cell_6t
Xbit_r241_c174 bl[174] br[174] wl[241] vdd gnd cell_6t
Xbit_r242_c174 bl[174] br[174] wl[242] vdd gnd cell_6t
Xbit_r243_c174 bl[174] br[174] wl[243] vdd gnd cell_6t
Xbit_r244_c174 bl[174] br[174] wl[244] vdd gnd cell_6t
Xbit_r245_c174 bl[174] br[174] wl[245] vdd gnd cell_6t
Xbit_r246_c174 bl[174] br[174] wl[246] vdd gnd cell_6t
Xbit_r247_c174 bl[174] br[174] wl[247] vdd gnd cell_6t
Xbit_r248_c174 bl[174] br[174] wl[248] vdd gnd cell_6t
Xbit_r249_c174 bl[174] br[174] wl[249] vdd gnd cell_6t
Xbit_r250_c174 bl[174] br[174] wl[250] vdd gnd cell_6t
Xbit_r251_c174 bl[174] br[174] wl[251] vdd gnd cell_6t
Xbit_r252_c174 bl[174] br[174] wl[252] vdd gnd cell_6t
Xbit_r253_c174 bl[174] br[174] wl[253] vdd gnd cell_6t
Xbit_r254_c174 bl[174] br[174] wl[254] vdd gnd cell_6t
Xbit_r255_c174 bl[174] br[174] wl[255] vdd gnd cell_6t
Xbit_r0_c175 bl[175] br[175] wl[0] vdd gnd cell_6t
Xbit_r1_c175 bl[175] br[175] wl[1] vdd gnd cell_6t
Xbit_r2_c175 bl[175] br[175] wl[2] vdd gnd cell_6t
Xbit_r3_c175 bl[175] br[175] wl[3] vdd gnd cell_6t
Xbit_r4_c175 bl[175] br[175] wl[4] vdd gnd cell_6t
Xbit_r5_c175 bl[175] br[175] wl[5] vdd gnd cell_6t
Xbit_r6_c175 bl[175] br[175] wl[6] vdd gnd cell_6t
Xbit_r7_c175 bl[175] br[175] wl[7] vdd gnd cell_6t
Xbit_r8_c175 bl[175] br[175] wl[8] vdd gnd cell_6t
Xbit_r9_c175 bl[175] br[175] wl[9] vdd gnd cell_6t
Xbit_r10_c175 bl[175] br[175] wl[10] vdd gnd cell_6t
Xbit_r11_c175 bl[175] br[175] wl[11] vdd gnd cell_6t
Xbit_r12_c175 bl[175] br[175] wl[12] vdd gnd cell_6t
Xbit_r13_c175 bl[175] br[175] wl[13] vdd gnd cell_6t
Xbit_r14_c175 bl[175] br[175] wl[14] vdd gnd cell_6t
Xbit_r15_c175 bl[175] br[175] wl[15] vdd gnd cell_6t
Xbit_r16_c175 bl[175] br[175] wl[16] vdd gnd cell_6t
Xbit_r17_c175 bl[175] br[175] wl[17] vdd gnd cell_6t
Xbit_r18_c175 bl[175] br[175] wl[18] vdd gnd cell_6t
Xbit_r19_c175 bl[175] br[175] wl[19] vdd gnd cell_6t
Xbit_r20_c175 bl[175] br[175] wl[20] vdd gnd cell_6t
Xbit_r21_c175 bl[175] br[175] wl[21] vdd gnd cell_6t
Xbit_r22_c175 bl[175] br[175] wl[22] vdd gnd cell_6t
Xbit_r23_c175 bl[175] br[175] wl[23] vdd gnd cell_6t
Xbit_r24_c175 bl[175] br[175] wl[24] vdd gnd cell_6t
Xbit_r25_c175 bl[175] br[175] wl[25] vdd gnd cell_6t
Xbit_r26_c175 bl[175] br[175] wl[26] vdd gnd cell_6t
Xbit_r27_c175 bl[175] br[175] wl[27] vdd gnd cell_6t
Xbit_r28_c175 bl[175] br[175] wl[28] vdd gnd cell_6t
Xbit_r29_c175 bl[175] br[175] wl[29] vdd gnd cell_6t
Xbit_r30_c175 bl[175] br[175] wl[30] vdd gnd cell_6t
Xbit_r31_c175 bl[175] br[175] wl[31] vdd gnd cell_6t
Xbit_r32_c175 bl[175] br[175] wl[32] vdd gnd cell_6t
Xbit_r33_c175 bl[175] br[175] wl[33] vdd gnd cell_6t
Xbit_r34_c175 bl[175] br[175] wl[34] vdd gnd cell_6t
Xbit_r35_c175 bl[175] br[175] wl[35] vdd gnd cell_6t
Xbit_r36_c175 bl[175] br[175] wl[36] vdd gnd cell_6t
Xbit_r37_c175 bl[175] br[175] wl[37] vdd gnd cell_6t
Xbit_r38_c175 bl[175] br[175] wl[38] vdd gnd cell_6t
Xbit_r39_c175 bl[175] br[175] wl[39] vdd gnd cell_6t
Xbit_r40_c175 bl[175] br[175] wl[40] vdd gnd cell_6t
Xbit_r41_c175 bl[175] br[175] wl[41] vdd gnd cell_6t
Xbit_r42_c175 bl[175] br[175] wl[42] vdd gnd cell_6t
Xbit_r43_c175 bl[175] br[175] wl[43] vdd gnd cell_6t
Xbit_r44_c175 bl[175] br[175] wl[44] vdd gnd cell_6t
Xbit_r45_c175 bl[175] br[175] wl[45] vdd gnd cell_6t
Xbit_r46_c175 bl[175] br[175] wl[46] vdd gnd cell_6t
Xbit_r47_c175 bl[175] br[175] wl[47] vdd gnd cell_6t
Xbit_r48_c175 bl[175] br[175] wl[48] vdd gnd cell_6t
Xbit_r49_c175 bl[175] br[175] wl[49] vdd gnd cell_6t
Xbit_r50_c175 bl[175] br[175] wl[50] vdd gnd cell_6t
Xbit_r51_c175 bl[175] br[175] wl[51] vdd gnd cell_6t
Xbit_r52_c175 bl[175] br[175] wl[52] vdd gnd cell_6t
Xbit_r53_c175 bl[175] br[175] wl[53] vdd gnd cell_6t
Xbit_r54_c175 bl[175] br[175] wl[54] vdd gnd cell_6t
Xbit_r55_c175 bl[175] br[175] wl[55] vdd gnd cell_6t
Xbit_r56_c175 bl[175] br[175] wl[56] vdd gnd cell_6t
Xbit_r57_c175 bl[175] br[175] wl[57] vdd gnd cell_6t
Xbit_r58_c175 bl[175] br[175] wl[58] vdd gnd cell_6t
Xbit_r59_c175 bl[175] br[175] wl[59] vdd gnd cell_6t
Xbit_r60_c175 bl[175] br[175] wl[60] vdd gnd cell_6t
Xbit_r61_c175 bl[175] br[175] wl[61] vdd gnd cell_6t
Xbit_r62_c175 bl[175] br[175] wl[62] vdd gnd cell_6t
Xbit_r63_c175 bl[175] br[175] wl[63] vdd gnd cell_6t
Xbit_r64_c175 bl[175] br[175] wl[64] vdd gnd cell_6t
Xbit_r65_c175 bl[175] br[175] wl[65] vdd gnd cell_6t
Xbit_r66_c175 bl[175] br[175] wl[66] vdd gnd cell_6t
Xbit_r67_c175 bl[175] br[175] wl[67] vdd gnd cell_6t
Xbit_r68_c175 bl[175] br[175] wl[68] vdd gnd cell_6t
Xbit_r69_c175 bl[175] br[175] wl[69] vdd gnd cell_6t
Xbit_r70_c175 bl[175] br[175] wl[70] vdd gnd cell_6t
Xbit_r71_c175 bl[175] br[175] wl[71] vdd gnd cell_6t
Xbit_r72_c175 bl[175] br[175] wl[72] vdd gnd cell_6t
Xbit_r73_c175 bl[175] br[175] wl[73] vdd gnd cell_6t
Xbit_r74_c175 bl[175] br[175] wl[74] vdd gnd cell_6t
Xbit_r75_c175 bl[175] br[175] wl[75] vdd gnd cell_6t
Xbit_r76_c175 bl[175] br[175] wl[76] vdd gnd cell_6t
Xbit_r77_c175 bl[175] br[175] wl[77] vdd gnd cell_6t
Xbit_r78_c175 bl[175] br[175] wl[78] vdd gnd cell_6t
Xbit_r79_c175 bl[175] br[175] wl[79] vdd gnd cell_6t
Xbit_r80_c175 bl[175] br[175] wl[80] vdd gnd cell_6t
Xbit_r81_c175 bl[175] br[175] wl[81] vdd gnd cell_6t
Xbit_r82_c175 bl[175] br[175] wl[82] vdd gnd cell_6t
Xbit_r83_c175 bl[175] br[175] wl[83] vdd gnd cell_6t
Xbit_r84_c175 bl[175] br[175] wl[84] vdd gnd cell_6t
Xbit_r85_c175 bl[175] br[175] wl[85] vdd gnd cell_6t
Xbit_r86_c175 bl[175] br[175] wl[86] vdd gnd cell_6t
Xbit_r87_c175 bl[175] br[175] wl[87] vdd gnd cell_6t
Xbit_r88_c175 bl[175] br[175] wl[88] vdd gnd cell_6t
Xbit_r89_c175 bl[175] br[175] wl[89] vdd gnd cell_6t
Xbit_r90_c175 bl[175] br[175] wl[90] vdd gnd cell_6t
Xbit_r91_c175 bl[175] br[175] wl[91] vdd gnd cell_6t
Xbit_r92_c175 bl[175] br[175] wl[92] vdd gnd cell_6t
Xbit_r93_c175 bl[175] br[175] wl[93] vdd gnd cell_6t
Xbit_r94_c175 bl[175] br[175] wl[94] vdd gnd cell_6t
Xbit_r95_c175 bl[175] br[175] wl[95] vdd gnd cell_6t
Xbit_r96_c175 bl[175] br[175] wl[96] vdd gnd cell_6t
Xbit_r97_c175 bl[175] br[175] wl[97] vdd gnd cell_6t
Xbit_r98_c175 bl[175] br[175] wl[98] vdd gnd cell_6t
Xbit_r99_c175 bl[175] br[175] wl[99] vdd gnd cell_6t
Xbit_r100_c175 bl[175] br[175] wl[100] vdd gnd cell_6t
Xbit_r101_c175 bl[175] br[175] wl[101] vdd gnd cell_6t
Xbit_r102_c175 bl[175] br[175] wl[102] vdd gnd cell_6t
Xbit_r103_c175 bl[175] br[175] wl[103] vdd gnd cell_6t
Xbit_r104_c175 bl[175] br[175] wl[104] vdd gnd cell_6t
Xbit_r105_c175 bl[175] br[175] wl[105] vdd gnd cell_6t
Xbit_r106_c175 bl[175] br[175] wl[106] vdd gnd cell_6t
Xbit_r107_c175 bl[175] br[175] wl[107] vdd gnd cell_6t
Xbit_r108_c175 bl[175] br[175] wl[108] vdd gnd cell_6t
Xbit_r109_c175 bl[175] br[175] wl[109] vdd gnd cell_6t
Xbit_r110_c175 bl[175] br[175] wl[110] vdd gnd cell_6t
Xbit_r111_c175 bl[175] br[175] wl[111] vdd gnd cell_6t
Xbit_r112_c175 bl[175] br[175] wl[112] vdd gnd cell_6t
Xbit_r113_c175 bl[175] br[175] wl[113] vdd gnd cell_6t
Xbit_r114_c175 bl[175] br[175] wl[114] vdd gnd cell_6t
Xbit_r115_c175 bl[175] br[175] wl[115] vdd gnd cell_6t
Xbit_r116_c175 bl[175] br[175] wl[116] vdd gnd cell_6t
Xbit_r117_c175 bl[175] br[175] wl[117] vdd gnd cell_6t
Xbit_r118_c175 bl[175] br[175] wl[118] vdd gnd cell_6t
Xbit_r119_c175 bl[175] br[175] wl[119] vdd gnd cell_6t
Xbit_r120_c175 bl[175] br[175] wl[120] vdd gnd cell_6t
Xbit_r121_c175 bl[175] br[175] wl[121] vdd gnd cell_6t
Xbit_r122_c175 bl[175] br[175] wl[122] vdd gnd cell_6t
Xbit_r123_c175 bl[175] br[175] wl[123] vdd gnd cell_6t
Xbit_r124_c175 bl[175] br[175] wl[124] vdd gnd cell_6t
Xbit_r125_c175 bl[175] br[175] wl[125] vdd gnd cell_6t
Xbit_r126_c175 bl[175] br[175] wl[126] vdd gnd cell_6t
Xbit_r127_c175 bl[175] br[175] wl[127] vdd gnd cell_6t
Xbit_r128_c175 bl[175] br[175] wl[128] vdd gnd cell_6t
Xbit_r129_c175 bl[175] br[175] wl[129] vdd gnd cell_6t
Xbit_r130_c175 bl[175] br[175] wl[130] vdd gnd cell_6t
Xbit_r131_c175 bl[175] br[175] wl[131] vdd gnd cell_6t
Xbit_r132_c175 bl[175] br[175] wl[132] vdd gnd cell_6t
Xbit_r133_c175 bl[175] br[175] wl[133] vdd gnd cell_6t
Xbit_r134_c175 bl[175] br[175] wl[134] vdd gnd cell_6t
Xbit_r135_c175 bl[175] br[175] wl[135] vdd gnd cell_6t
Xbit_r136_c175 bl[175] br[175] wl[136] vdd gnd cell_6t
Xbit_r137_c175 bl[175] br[175] wl[137] vdd gnd cell_6t
Xbit_r138_c175 bl[175] br[175] wl[138] vdd gnd cell_6t
Xbit_r139_c175 bl[175] br[175] wl[139] vdd gnd cell_6t
Xbit_r140_c175 bl[175] br[175] wl[140] vdd gnd cell_6t
Xbit_r141_c175 bl[175] br[175] wl[141] vdd gnd cell_6t
Xbit_r142_c175 bl[175] br[175] wl[142] vdd gnd cell_6t
Xbit_r143_c175 bl[175] br[175] wl[143] vdd gnd cell_6t
Xbit_r144_c175 bl[175] br[175] wl[144] vdd gnd cell_6t
Xbit_r145_c175 bl[175] br[175] wl[145] vdd gnd cell_6t
Xbit_r146_c175 bl[175] br[175] wl[146] vdd gnd cell_6t
Xbit_r147_c175 bl[175] br[175] wl[147] vdd gnd cell_6t
Xbit_r148_c175 bl[175] br[175] wl[148] vdd gnd cell_6t
Xbit_r149_c175 bl[175] br[175] wl[149] vdd gnd cell_6t
Xbit_r150_c175 bl[175] br[175] wl[150] vdd gnd cell_6t
Xbit_r151_c175 bl[175] br[175] wl[151] vdd gnd cell_6t
Xbit_r152_c175 bl[175] br[175] wl[152] vdd gnd cell_6t
Xbit_r153_c175 bl[175] br[175] wl[153] vdd gnd cell_6t
Xbit_r154_c175 bl[175] br[175] wl[154] vdd gnd cell_6t
Xbit_r155_c175 bl[175] br[175] wl[155] vdd gnd cell_6t
Xbit_r156_c175 bl[175] br[175] wl[156] vdd gnd cell_6t
Xbit_r157_c175 bl[175] br[175] wl[157] vdd gnd cell_6t
Xbit_r158_c175 bl[175] br[175] wl[158] vdd gnd cell_6t
Xbit_r159_c175 bl[175] br[175] wl[159] vdd gnd cell_6t
Xbit_r160_c175 bl[175] br[175] wl[160] vdd gnd cell_6t
Xbit_r161_c175 bl[175] br[175] wl[161] vdd gnd cell_6t
Xbit_r162_c175 bl[175] br[175] wl[162] vdd gnd cell_6t
Xbit_r163_c175 bl[175] br[175] wl[163] vdd gnd cell_6t
Xbit_r164_c175 bl[175] br[175] wl[164] vdd gnd cell_6t
Xbit_r165_c175 bl[175] br[175] wl[165] vdd gnd cell_6t
Xbit_r166_c175 bl[175] br[175] wl[166] vdd gnd cell_6t
Xbit_r167_c175 bl[175] br[175] wl[167] vdd gnd cell_6t
Xbit_r168_c175 bl[175] br[175] wl[168] vdd gnd cell_6t
Xbit_r169_c175 bl[175] br[175] wl[169] vdd gnd cell_6t
Xbit_r170_c175 bl[175] br[175] wl[170] vdd gnd cell_6t
Xbit_r171_c175 bl[175] br[175] wl[171] vdd gnd cell_6t
Xbit_r172_c175 bl[175] br[175] wl[172] vdd gnd cell_6t
Xbit_r173_c175 bl[175] br[175] wl[173] vdd gnd cell_6t
Xbit_r174_c175 bl[175] br[175] wl[174] vdd gnd cell_6t
Xbit_r175_c175 bl[175] br[175] wl[175] vdd gnd cell_6t
Xbit_r176_c175 bl[175] br[175] wl[176] vdd gnd cell_6t
Xbit_r177_c175 bl[175] br[175] wl[177] vdd gnd cell_6t
Xbit_r178_c175 bl[175] br[175] wl[178] vdd gnd cell_6t
Xbit_r179_c175 bl[175] br[175] wl[179] vdd gnd cell_6t
Xbit_r180_c175 bl[175] br[175] wl[180] vdd gnd cell_6t
Xbit_r181_c175 bl[175] br[175] wl[181] vdd gnd cell_6t
Xbit_r182_c175 bl[175] br[175] wl[182] vdd gnd cell_6t
Xbit_r183_c175 bl[175] br[175] wl[183] vdd gnd cell_6t
Xbit_r184_c175 bl[175] br[175] wl[184] vdd gnd cell_6t
Xbit_r185_c175 bl[175] br[175] wl[185] vdd gnd cell_6t
Xbit_r186_c175 bl[175] br[175] wl[186] vdd gnd cell_6t
Xbit_r187_c175 bl[175] br[175] wl[187] vdd gnd cell_6t
Xbit_r188_c175 bl[175] br[175] wl[188] vdd gnd cell_6t
Xbit_r189_c175 bl[175] br[175] wl[189] vdd gnd cell_6t
Xbit_r190_c175 bl[175] br[175] wl[190] vdd gnd cell_6t
Xbit_r191_c175 bl[175] br[175] wl[191] vdd gnd cell_6t
Xbit_r192_c175 bl[175] br[175] wl[192] vdd gnd cell_6t
Xbit_r193_c175 bl[175] br[175] wl[193] vdd gnd cell_6t
Xbit_r194_c175 bl[175] br[175] wl[194] vdd gnd cell_6t
Xbit_r195_c175 bl[175] br[175] wl[195] vdd gnd cell_6t
Xbit_r196_c175 bl[175] br[175] wl[196] vdd gnd cell_6t
Xbit_r197_c175 bl[175] br[175] wl[197] vdd gnd cell_6t
Xbit_r198_c175 bl[175] br[175] wl[198] vdd gnd cell_6t
Xbit_r199_c175 bl[175] br[175] wl[199] vdd gnd cell_6t
Xbit_r200_c175 bl[175] br[175] wl[200] vdd gnd cell_6t
Xbit_r201_c175 bl[175] br[175] wl[201] vdd gnd cell_6t
Xbit_r202_c175 bl[175] br[175] wl[202] vdd gnd cell_6t
Xbit_r203_c175 bl[175] br[175] wl[203] vdd gnd cell_6t
Xbit_r204_c175 bl[175] br[175] wl[204] vdd gnd cell_6t
Xbit_r205_c175 bl[175] br[175] wl[205] vdd gnd cell_6t
Xbit_r206_c175 bl[175] br[175] wl[206] vdd gnd cell_6t
Xbit_r207_c175 bl[175] br[175] wl[207] vdd gnd cell_6t
Xbit_r208_c175 bl[175] br[175] wl[208] vdd gnd cell_6t
Xbit_r209_c175 bl[175] br[175] wl[209] vdd gnd cell_6t
Xbit_r210_c175 bl[175] br[175] wl[210] vdd gnd cell_6t
Xbit_r211_c175 bl[175] br[175] wl[211] vdd gnd cell_6t
Xbit_r212_c175 bl[175] br[175] wl[212] vdd gnd cell_6t
Xbit_r213_c175 bl[175] br[175] wl[213] vdd gnd cell_6t
Xbit_r214_c175 bl[175] br[175] wl[214] vdd gnd cell_6t
Xbit_r215_c175 bl[175] br[175] wl[215] vdd gnd cell_6t
Xbit_r216_c175 bl[175] br[175] wl[216] vdd gnd cell_6t
Xbit_r217_c175 bl[175] br[175] wl[217] vdd gnd cell_6t
Xbit_r218_c175 bl[175] br[175] wl[218] vdd gnd cell_6t
Xbit_r219_c175 bl[175] br[175] wl[219] vdd gnd cell_6t
Xbit_r220_c175 bl[175] br[175] wl[220] vdd gnd cell_6t
Xbit_r221_c175 bl[175] br[175] wl[221] vdd gnd cell_6t
Xbit_r222_c175 bl[175] br[175] wl[222] vdd gnd cell_6t
Xbit_r223_c175 bl[175] br[175] wl[223] vdd gnd cell_6t
Xbit_r224_c175 bl[175] br[175] wl[224] vdd gnd cell_6t
Xbit_r225_c175 bl[175] br[175] wl[225] vdd gnd cell_6t
Xbit_r226_c175 bl[175] br[175] wl[226] vdd gnd cell_6t
Xbit_r227_c175 bl[175] br[175] wl[227] vdd gnd cell_6t
Xbit_r228_c175 bl[175] br[175] wl[228] vdd gnd cell_6t
Xbit_r229_c175 bl[175] br[175] wl[229] vdd gnd cell_6t
Xbit_r230_c175 bl[175] br[175] wl[230] vdd gnd cell_6t
Xbit_r231_c175 bl[175] br[175] wl[231] vdd gnd cell_6t
Xbit_r232_c175 bl[175] br[175] wl[232] vdd gnd cell_6t
Xbit_r233_c175 bl[175] br[175] wl[233] vdd gnd cell_6t
Xbit_r234_c175 bl[175] br[175] wl[234] vdd gnd cell_6t
Xbit_r235_c175 bl[175] br[175] wl[235] vdd gnd cell_6t
Xbit_r236_c175 bl[175] br[175] wl[236] vdd gnd cell_6t
Xbit_r237_c175 bl[175] br[175] wl[237] vdd gnd cell_6t
Xbit_r238_c175 bl[175] br[175] wl[238] vdd gnd cell_6t
Xbit_r239_c175 bl[175] br[175] wl[239] vdd gnd cell_6t
Xbit_r240_c175 bl[175] br[175] wl[240] vdd gnd cell_6t
Xbit_r241_c175 bl[175] br[175] wl[241] vdd gnd cell_6t
Xbit_r242_c175 bl[175] br[175] wl[242] vdd gnd cell_6t
Xbit_r243_c175 bl[175] br[175] wl[243] vdd gnd cell_6t
Xbit_r244_c175 bl[175] br[175] wl[244] vdd gnd cell_6t
Xbit_r245_c175 bl[175] br[175] wl[245] vdd gnd cell_6t
Xbit_r246_c175 bl[175] br[175] wl[246] vdd gnd cell_6t
Xbit_r247_c175 bl[175] br[175] wl[247] vdd gnd cell_6t
Xbit_r248_c175 bl[175] br[175] wl[248] vdd gnd cell_6t
Xbit_r249_c175 bl[175] br[175] wl[249] vdd gnd cell_6t
Xbit_r250_c175 bl[175] br[175] wl[250] vdd gnd cell_6t
Xbit_r251_c175 bl[175] br[175] wl[251] vdd gnd cell_6t
Xbit_r252_c175 bl[175] br[175] wl[252] vdd gnd cell_6t
Xbit_r253_c175 bl[175] br[175] wl[253] vdd gnd cell_6t
Xbit_r254_c175 bl[175] br[175] wl[254] vdd gnd cell_6t
Xbit_r255_c175 bl[175] br[175] wl[255] vdd gnd cell_6t
Xbit_r0_c176 bl[176] br[176] wl[0] vdd gnd cell_6t
Xbit_r1_c176 bl[176] br[176] wl[1] vdd gnd cell_6t
Xbit_r2_c176 bl[176] br[176] wl[2] vdd gnd cell_6t
Xbit_r3_c176 bl[176] br[176] wl[3] vdd gnd cell_6t
Xbit_r4_c176 bl[176] br[176] wl[4] vdd gnd cell_6t
Xbit_r5_c176 bl[176] br[176] wl[5] vdd gnd cell_6t
Xbit_r6_c176 bl[176] br[176] wl[6] vdd gnd cell_6t
Xbit_r7_c176 bl[176] br[176] wl[7] vdd gnd cell_6t
Xbit_r8_c176 bl[176] br[176] wl[8] vdd gnd cell_6t
Xbit_r9_c176 bl[176] br[176] wl[9] vdd gnd cell_6t
Xbit_r10_c176 bl[176] br[176] wl[10] vdd gnd cell_6t
Xbit_r11_c176 bl[176] br[176] wl[11] vdd gnd cell_6t
Xbit_r12_c176 bl[176] br[176] wl[12] vdd gnd cell_6t
Xbit_r13_c176 bl[176] br[176] wl[13] vdd gnd cell_6t
Xbit_r14_c176 bl[176] br[176] wl[14] vdd gnd cell_6t
Xbit_r15_c176 bl[176] br[176] wl[15] vdd gnd cell_6t
Xbit_r16_c176 bl[176] br[176] wl[16] vdd gnd cell_6t
Xbit_r17_c176 bl[176] br[176] wl[17] vdd gnd cell_6t
Xbit_r18_c176 bl[176] br[176] wl[18] vdd gnd cell_6t
Xbit_r19_c176 bl[176] br[176] wl[19] vdd gnd cell_6t
Xbit_r20_c176 bl[176] br[176] wl[20] vdd gnd cell_6t
Xbit_r21_c176 bl[176] br[176] wl[21] vdd gnd cell_6t
Xbit_r22_c176 bl[176] br[176] wl[22] vdd gnd cell_6t
Xbit_r23_c176 bl[176] br[176] wl[23] vdd gnd cell_6t
Xbit_r24_c176 bl[176] br[176] wl[24] vdd gnd cell_6t
Xbit_r25_c176 bl[176] br[176] wl[25] vdd gnd cell_6t
Xbit_r26_c176 bl[176] br[176] wl[26] vdd gnd cell_6t
Xbit_r27_c176 bl[176] br[176] wl[27] vdd gnd cell_6t
Xbit_r28_c176 bl[176] br[176] wl[28] vdd gnd cell_6t
Xbit_r29_c176 bl[176] br[176] wl[29] vdd gnd cell_6t
Xbit_r30_c176 bl[176] br[176] wl[30] vdd gnd cell_6t
Xbit_r31_c176 bl[176] br[176] wl[31] vdd gnd cell_6t
Xbit_r32_c176 bl[176] br[176] wl[32] vdd gnd cell_6t
Xbit_r33_c176 bl[176] br[176] wl[33] vdd gnd cell_6t
Xbit_r34_c176 bl[176] br[176] wl[34] vdd gnd cell_6t
Xbit_r35_c176 bl[176] br[176] wl[35] vdd gnd cell_6t
Xbit_r36_c176 bl[176] br[176] wl[36] vdd gnd cell_6t
Xbit_r37_c176 bl[176] br[176] wl[37] vdd gnd cell_6t
Xbit_r38_c176 bl[176] br[176] wl[38] vdd gnd cell_6t
Xbit_r39_c176 bl[176] br[176] wl[39] vdd gnd cell_6t
Xbit_r40_c176 bl[176] br[176] wl[40] vdd gnd cell_6t
Xbit_r41_c176 bl[176] br[176] wl[41] vdd gnd cell_6t
Xbit_r42_c176 bl[176] br[176] wl[42] vdd gnd cell_6t
Xbit_r43_c176 bl[176] br[176] wl[43] vdd gnd cell_6t
Xbit_r44_c176 bl[176] br[176] wl[44] vdd gnd cell_6t
Xbit_r45_c176 bl[176] br[176] wl[45] vdd gnd cell_6t
Xbit_r46_c176 bl[176] br[176] wl[46] vdd gnd cell_6t
Xbit_r47_c176 bl[176] br[176] wl[47] vdd gnd cell_6t
Xbit_r48_c176 bl[176] br[176] wl[48] vdd gnd cell_6t
Xbit_r49_c176 bl[176] br[176] wl[49] vdd gnd cell_6t
Xbit_r50_c176 bl[176] br[176] wl[50] vdd gnd cell_6t
Xbit_r51_c176 bl[176] br[176] wl[51] vdd gnd cell_6t
Xbit_r52_c176 bl[176] br[176] wl[52] vdd gnd cell_6t
Xbit_r53_c176 bl[176] br[176] wl[53] vdd gnd cell_6t
Xbit_r54_c176 bl[176] br[176] wl[54] vdd gnd cell_6t
Xbit_r55_c176 bl[176] br[176] wl[55] vdd gnd cell_6t
Xbit_r56_c176 bl[176] br[176] wl[56] vdd gnd cell_6t
Xbit_r57_c176 bl[176] br[176] wl[57] vdd gnd cell_6t
Xbit_r58_c176 bl[176] br[176] wl[58] vdd gnd cell_6t
Xbit_r59_c176 bl[176] br[176] wl[59] vdd gnd cell_6t
Xbit_r60_c176 bl[176] br[176] wl[60] vdd gnd cell_6t
Xbit_r61_c176 bl[176] br[176] wl[61] vdd gnd cell_6t
Xbit_r62_c176 bl[176] br[176] wl[62] vdd gnd cell_6t
Xbit_r63_c176 bl[176] br[176] wl[63] vdd gnd cell_6t
Xbit_r64_c176 bl[176] br[176] wl[64] vdd gnd cell_6t
Xbit_r65_c176 bl[176] br[176] wl[65] vdd gnd cell_6t
Xbit_r66_c176 bl[176] br[176] wl[66] vdd gnd cell_6t
Xbit_r67_c176 bl[176] br[176] wl[67] vdd gnd cell_6t
Xbit_r68_c176 bl[176] br[176] wl[68] vdd gnd cell_6t
Xbit_r69_c176 bl[176] br[176] wl[69] vdd gnd cell_6t
Xbit_r70_c176 bl[176] br[176] wl[70] vdd gnd cell_6t
Xbit_r71_c176 bl[176] br[176] wl[71] vdd gnd cell_6t
Xbit_r72_c176 bl[176] br[176] wl[72] vdd gnd cell_6t
Xbit_r73_c176 bl[176] br[176] wl[73] vdd gnd cell_6t
Xbit_r74_c176 bl[176] br[176] wl[74] vdd gnd cell_6t
Xbit_r75_c176 bl[176] br[176] wl[75] vdd gnd cell_6t
Xbit_r76_c176 bl[176] br[176] wl[76] vdd gnd cell_6t
Xbit_r77_c176 bl[176] br[176] wl[77] vdd gnd cell_6t
Xbit_r78_c176 bl[176] br[176] wl[78] vdd gnd cell_6t
Xbit_r79_c176 bl[176] br[176] wl[79] vdd gnd cell_6t
Xbit_r80_c176 bl[176] br[176] wl[80] vdd gnd cell_6t
Xbit_r81_c176 bl[176] br[176] wl[81] vdd gnd cell_6t
Xbit_r82_c176 bl[176] br[176] wl[82] vdd gnd cell_6t
Xbit_r83_c176 bl[176] br[176] wl[83] vdd gnd cell_6t
Xbit_r84_c176 bl[176] br[176] wl[84] vdd gnd cell_6t
Xbit_r85_c176 bl[176] br[176] wl[85] vdd gnd cell_6t
Xbit_r86_c176 bl[176] br[176] wl[86] vdd gnd cell_6t
Xbit_r87_c176 bl[176] br[176] wl[87] vdd gnd cell_6t
Xbit_r88_c176 bl[176] br[176] wl[88] vdd gnd cell_6t
Xbit_r89_c176 bl[176] br[176] wl[89] vdd gnd cell_6t
Xbit_r90_c176 bl[176] br[176] wl[90] vdd gnd cell_6t
Xbit_r91_c176 bl[176] br[176] wl[91] vdd gnd cell_6t
Xbit_r92_c176 bl[176] br[176] wl[92] vdd gnd cell_6t
Xbit_r93_c176 bl[176] br[176] wl[93] vdd gnd cell_6t
Xbit_r94_c176 bl[176] br[176] wl[94] vdd gnd cell_6t
Xbit_r95_c176 bl[176] br[176] wl[95] vdd gnd cell_6t
Xbit_r96_c176 bl[176] br[176] wl[96] vdd gnd cell_6t
Xbit_r97_c176 bl[176] br[176] wl[97] vdd gnd cell_6t
Xbit_r98_c176 bl[176] br[176] wl[98] vdd gnd cell_6t
Xbit_r99_c176 bl[176] br[176] wl[99] vdd gnd cell_6t
Xbit_r100_c176 bl[176] br[176] wl[100] vdd gnd cell_6t
Xbit_r101_c176 bl[176] br[176] wl[101] vdd gnd cell_6t
Xbit_r102_c176 bl[176] br[176] wl[102] vdd gnd cell_6t
Xbit_r103_c176 bl[176] br[176] wl[103] vdd gnd cell_6t
Xbit_r104_c176 bl[176] br[176] wl[104] vdd gnd cell_6t
Xbit_r105_c176 bl[176] br[176] wl[105] vdd gnd cell_6t
Xbit_r106_c176 bl[176] br[176] wl[106] vdd gnd cell_6t
Xbit_r107_c176 bl[176] br[176] wl[107] vdd gnd cell_6t
Xbit_r108_c176 bl[176] br[176] wl[108] vdd gnd cell_6t
Xbit_r109_c176 bl[176] br[176] wl[109] vdd gnd cell_6t
Xbit_r110_c176 bl[176] br[176] wl[110] vdd gnd cell_6t
Xbit_r111_c176 bl[176] br[176] wl[111] vdd gnd cell_6t
Xbit_r112_c176 bl[176] br[176] wl[112] vdd gnd cell_6t
Xbit_r113_c176 bl[176] br[176] wl[113] vdd gnd cell_6t
Xbit_r114_c176 bl[176] br[176] wl[114] vdd gnd cell_6t
Xbit_r115_c176 bl[176] br[176] wl[115] vdd gnd cell_6t
Xbit_r116_c176 bl[176] br[176] wl[116] vdd gnd cell_6t
Xbit_r117_c176 bl[176] br[176] wl[117] vdd gnd cell_6t
Xbit_r118_c176 bl[176] br[176] wl[118] vdd gnd cell_6t
Xbit_r119_c176 bl[176] br[176] wl[119] vdd gnd cell_6t
Xbit_r120_c176 bl[176] br[176] wl[120] vdd gnd cell_6t
Xbit_r121_c176 bl[176] br[176] wl[121] vdd gnd cell_6t
Xbit_r122_c176 bl[176] br[176] wl[122] vdd gnd cell_6t
Xbit_r123_c176 bl[176] br[176] wl[123] vdd gnd cell_6t
Xbit_r124_c176 bl[176] br[176] wl[124] vdd gnd cell_6t
Xbit_r125_c176 bl[176] br[176] wl[125] vdd gnd cell_6t
Xbit_r126_c176 bl[176] br[176] wl[126] vdd gnd cell_6t
Xbit_r127_c176 bl[176] br[176] wl[127] vdd gnd cell_6t
Xbit_r128_c176 bl[176] br[176] wl[128] vdd gnd cell_6t
Xbit_r129_c176 bl[176] br[176] wl[129] vdd gnd cell_6t
Xbit_r130_c176 bl[176] br[176] wl[130] vdd gnd cell_6t
Xbit_r131_c176 bl[176] br[176] wl[131] vdd gnd cell_6t
Xbit_r132_c176 bl[176] br[176] wl[132] vdd gnd cell_6t
Xbit_r133_c176 bl[176] br[176] wl[133] vdd gnd cell_6t
Xbit_r134_c176 bl[176] br[176] wl[134] vdd gnd cell_6t
Xbit_r135_c176 bl[176] br[176] wl[135] vdd gnd cell_6t
Xbit_r136_c176 bl[176] br[176] wl[136] vdd gnd cell_6t
Xbit_r137_c176 bl[176] br[176] wl[137] vdd gnd cell_6t
Xbit_r138_c176 bl[176] br[176] wl[138] vdd gnd cell_6t
Xbit_r139_c176 bl[176] br[176] wl[139] vdd gnd cell_6t
Xbit_r140_c176 bl[176] br[176] wl[140] vdd gnd cell_6t
Xbit_r141_c176 bl[176] br[176] wl[141] vdd gnd cell_6t
Xbit_r142_c176 bl[176] br[176] wl[142] vdd gnd cell_6t
Xbit_r143_c176 bl[176] br[176] wl[143] vdd gnd cell_6t
Xbit_r144_c176 bl[176] br[176] wl[144] vdd gnd cell_6t
Xbit_r145_c176 bl[176] br[176] wl[145] vdd gnd cell_6t
Xbit_r146_c176 bl[176] br[176] wl[146] vdd gnd cell_6t
Xbit_r147_c176 bl[176] br[176] wl[147] vdd gnd cell_6t
Xbit_r148_c176 bl[176] br[176] wl[148] vdd gnd cell_6t
Xbit_r149_c176 bl[176] br[176] wl[149] vdd gnd cell_6t
Xbit_r150_c176 bl[176] br[176] wl[150] vdd gnd cell_6t
Xbit_r151_c176 bl[176] br[176] wl[151] vdd gnd cell_6t
Xbit_r152_c176 bl[176] br[176] wl[152] vdd gnd cell_6t
Xbit_r153_c176 bl[176] br[176] wl[153] vdd gnd cell_6t
Xbit_r154_c176 bl[176] br[176] wl[154] vdd gnd cell_6t
Xbit_r155_c176 bl[176] br[176] wl[155] vdd gnd cell_6t
Xbit_r156_c176 bl[176] br[176] wl[156] vdd gnd cell_6t
Xbit_r157_c176 bl[176] br[176] wl[157] vdd gnd cell_6t
Xbit_r158_c176 bl[176] br[176] wl[158] vdd gnd cell_6t
Xbit_r159_c176 bl[176] br[176] wl[159] vdd gnd cell_6t
Xbit_r160_c176 bl[176] br[176] wl[160] vdd gnd cell_6t
Xbit_r161_c176 bl[176] br[176] wl[161] vdd gnd cell_6t
Xbit_r162_c176 bl[176] br[176] wl[162] vdd gnd cell_6t
Xbit_r163_c176 bl[176] br[176] wl[163] vdd gnd cell_6t
Xbit_r164_c176 bl[176] br[176] wl[164] vdd gnd cell_6t
Xbit_r165_c176 bl[176] br[176] wl[165] vdd gnd cell_6t
Xbit_r166_c176 bl[176] br[176] wl[166] vdd gnd cell_6t
Xbit_r167_c176 bl[176] br[176] wl[167] vdd gnd cell_6t
Xbit_r168_c176 bl[176] br[176] wl[168] vdd gnd cell_6t
Xbit_r169_c176 bl[176] br[176] wl[169] vdd gnd cell_6t
Xbit_r170_c176 bl[176] br[176] wl[170] vdd gnd cell_6t
Xbit_r171_c176 bl[176] br[176] wl[171] vdd gnd cell_6t
Xbit_r172_c176 bl[176] br[176] wl[172] vdd gnd cell_6t
Xbit_r173_c176 bl[176] br[176] wl[173] vdd gnd cell_6t
Xbit_r174_c176 bl[176] br[176] wl[174] vdd gnd cell_6t
Xbit_r175_c176 bl[176] br[176] wl[175] vdd gnd cell_6t
Xbit_r176_c176 bl[176] br[176] wl[176] vdd gnd cell_6t
Xbit_r177_c176 bl[176] br[176] wl[177] vdd gnd cell_6t
Xbit_r178_c176 bl[176] br[176] wl[178] vdd gnd cell_6t
Xbit_r179_c176 bl[176] br[176] wl[179] vdd gnd cell_6t
Xbit_r180_c176 bl[176] br[176] wl[180] vdd gnd cell_6t
Xbit_r181_c176 bl[176] br[176] wl[181] vdd gnd cell_6t
Xbit_r182_c176 bl[176] br[176] wl[182] vdd gnd cell_6t
Xbit_r183_c176 bl[176] br[176] wl[183] vdd gnd cell_6t
Xbit_r184_c176 bl[176] br[176] wl[184] vdd gnd cell_6t
Xbit_r185_c176 bl[176] br[176] wl[185] vdd gnd cell_6t
Xbit_r186_c176 bl[176] br[176] wl[186] vdd gnd cell_6t
Xbit_r187_c176 bl[176] br[176] wl[187] vdd gnd cell_6t
Xbit_r188_c176 bl[176] br[176] wl[188] vdd gnd cell_6t
Xbit_r189_c176 bl[176] br[176] wl[189] vdd gnd cell_6t
Xbit_r190_c176 bl[176] br[176] wl[190] vdd gnd cell_6t
Xbit_r191_c176 bl[176] br[176] wl[191] vdd gnd cell_6t
Xbit_r192_c176 bl[176] br[176] wl[192] vdd gnd cell_6t
Xbit_r193_c176 bl[176] br[176] wl[193] vdd gnd cell_6t
Xbit_r194_c176 bl[176] br[176] wl[194] vdd gnd cell_6t
Xbit_r195_c176 bl[176] br[176] wl[195] vdd gnd cell_6t
Xbit_r196_c176 bl[176] br[176] wl[196] vdd gnd cell_6t
Xbit_r197_c176 bl[176] br[176] wl[197] vdd gnd cell_6t
Xbit_r198_c176 bl[176] br[176] wl[198] vdd gnd cell_6t
Xbit_r199_c176 bl[176] br[176] wl[199] vdd gnd cell_6t
Xbit_r200_c176 bl[176] br[176] wl[200] vdd gnd cell_6t
Xbit_r201_c176 bl[176] br[176] wl[201] vdd gnd cell_6t
Xbit_r202_c176 bl[176] br[176] wl[202] vdd gnd cell_6t
Xbit_r203_c176 bl[176] br[176] wl[203] vdd gnd cell_6t
Xbit_r204_c176 bl[176] br[176] wl[204] vdd gnd cell_6t
Xbit_r205_c176 bl[176] br[176] wl[205] vdd gnd cell_6t
Xbit_r206_c176 bl[176] br[176] wl[206] vdd gnd cell_6t
Xbit_r207_c176 bl[176] br[176] wl[207] vdd gnd cell_6t
Xbit_r208_c176 bl[176] br[176] wl[208] vdd gnd cell_6t
Xbit_r209_c176 bl[176] br[176] wl[209] vdd gnd cell_6t
Xbit_r210_c176 bl[176] br[176] wl[210] vdd gnd cell_6t
Xbit_r211_c176 bl[176] br[176] wl[211] vdd gnd cell_6t
Xbit_r212_c176 bl[176] br[176] wl[212] vdd gnd cell_6t
Xbit_r213_c176 bl[176] br[176] wl[213] vdd gnd cell_6t
Xbit_r214_c176 bl[176] br[176] wl[214] vdd gnd cell_6t
Xbit_r215_c176 bl[176] br[176] wl[215] vdd gnd cell_6t
Xbit_r216_c176 bl[176] br[176] wl[216] vdd gnd cell_6t
Xbit_r217_c176 bl[176] br[176] wl[217] vdd gnd cell_6t
Xbit_r218_c176 bl[176] br[176] wl[218] vdd gnd cell_6t
Xbit_r219_c176 bl[176] br[176] wl[219] vdd gnd cell_6t
Xbit_r220_c176 bl[176] br[176] wl[220] vdd gnd cell_6t
Xbit_r221_c176 bl[176] br[176] wl[221] vdd gnd cell_6t
Xbit_r222_c176 bl[176] br[176] wl[222] vdd gnd cell_6t
Xbit_r223_c176 bl[176] br[176] wl[223] vdd gnd cell_6t
Xbit_r224_c176 bl[176] br[176] wl[224] vdd gnd cell_6t
Xbit_r225_c176 bl[176] br[176] wl[225] vdd gnd cell_6t
Xbit_r226_c176 bl[176] br[176] wl[226] vdd gnd cell_6t
Xbit_r227_c176 bl[176] br[176] wl[227] vdd gnd cell_6t
Xbit_r228_c176 bl[176] br[176] wl[228] vdd gnd cell_6t
Xbit_r229_c176 bl[176] br[176] wl[229] vdd gnd cell_6t
Xbit_r230_c176 bl[176] br[176] wl[230] vdd gnd cell_6t
Xbit_r231_c176 bl[176] br[176] wl[231] vdd gnd cell_6t
Xbit_r232_c176 bl[176] br[176] wl[232] vdd gnd cell_6t
Xbit_r233_c176 bl[176] br[176] wl[233] vdd gnd cell_6t
Xbit_r234_c176 bl[176] br[176] wl[234] vdd gnd cell_6t
Xbit_r235_c176 bl[176] br[176] wl[235] vdd gnd cell_6t
Xbit_r236_c176 bl[176] br[176] wl[236] vdd gnd cell_6t
Xbit_r237_c176 bl[176] br[176] wl[237] vdd gnd cell_6t
Xbit_r238_c176 bl[176] br[176] wl[238] vdd gnd cell_6t
Xbit_r239_c176 bl[176] br[176] wl[239] vdd gnd cell_6t
Xbit_r240_c176 bl[176] br[176] wl[240] vdd gnd cell_6t
Xbit_r241_c176 bl[176] br[176] wl[241] vdd gnd cell_6t
Xbit_r242_c176 bl[176] br[176] wl[242] vdd gnd cell_6t
Xbit_r243_c176 bl[176] br[176] wl[243] vdd gnd cell_6t
Xbit_r244_c176 bl[176] br[176] wl[244] vdd gnd cell_6t
Xbit_r245_c176 bl[176] br[176] wl[245] vdd gnd cell_6t
Xbit_r246_c176 bl[176] br[176] wl[246] vdd gnd cell_6t
Xbit_r247_c176 bl[176] br[176] wl[247] vdd gnd cell_6t
Xbit_r248_c176 bl[176] br[176] wl[248] vdd gnd cell_6t
Xbit_r249_c176 bl[176] br[176] wl[249] vdd gnd cell_6t
Xbit_r250_c176 bl[176] br[176] wl[250] vdd gnd cell_6t
Xbit_r251_c176 bl[176] br[176] wl[251] vdd gnd cell_6t
Xbit_r252_c176 bl[176] br[176] wl[252] vdd gnd cell_6t
Xbit_r253_c176 bl[176] br[176] wl[253] vdd gnd cell_6t
Xbit_r254_c176 bl[176] br[176] wl[254] vdd gnd cell_6t
Xbit_r255_c176 bl[176] br[176] wl[255] vdd gnd cell_6t
Xbit_r0_c177 bl[177] br[177] wl[0] vdd gnd cell_6t
Xbit_r1_c177 bl[177] br[177] wl[1] vdd gnd cell_6t
Xbit_r2_c177 bl[177] br[177] wl[2] vdd gnd cell_6t
Xbit_r3_c177 bl[177] br[177] wl[3] vdd gnd cell_6t
Xbit_r4_c177 bl[177] br[177] wl[4] vdd gnd cell_6t
Xbit_r5_c177 bl[177] br[177] wl[5] vdd gnd cell_6t
Xbit_r6_c177 bl[177] br[177] wl[6] vdd gnd cell_6t
Xbit_r7_c177 bl[177] br[177] wl[7] vdd gnd cell_6t
Xbit_r8_c177 bl[177] br[177] wl[8] vdd gnd cell_6t
Xbit_r9_c177 bl[177] br[177] wl[9] vdd gnd cell_6t
Xbit_r10_c177 bl[177] br[177] wl[10] vdd gnd cell_6t
Xbit_r11_c177 bl[177] br[177] wl[11] vdd gnd cell_6t
Xbit_r12_c177 bl[177] br[177] wl[12] vdd gnd cell_6t
Xbit_r13_c177 bl[177] br[177] wl[13] vdd gnd cell_6t
Xbit_r14_c177 bl[177] br[177] wl[14] vdd gnd cell_6t
Xbit_r15_c177 bl[177] br[177] wl[15] vdd gnd cell_6t
Xbit_r16_c177 bl[177] br[177] wl[16] vdd gnd cell_6t
Xbit_r17_c177 bl[177] br[177] wl[17] vdd gnd cell_6t
Xbit_r18_c177 bl[177] br[177] wl[18] vdd gnd cell_6t
Xbit_r19_c177 bl[177] br[177] wl[19] vdd gnd cell_6t
Xbit_r20_c177 bl[177] br[177] wl[20] vdd gnd cell_6t
Xbit_r21_c177 bl[177] br[177] wl[21] vdd gnd cell_6t
Xbit_r22_c177 bl[177] br[177] wl[22] vdd gnd cell_6t
Xbit_r23_c177 bl[177] br[177] wl[23] vdd gnd cell_6t
Xbit_r24_c177 bl[177] br[177] wl[24] vdd gnd cell_6t
Xbit_r25_c177 bl[177] br[177] wl[25] vdd gnd cell_6t
Xbit_r26_c177 bl[177] br[177] wl[26] vdd gnd cell_6t
Xbit_r27_c177 bl[177] br[177] wl[27] vdd gnd cell_6t
Xbit_r28_c177 bl[177] br[177] wl[28] vdd gnd cell_6t
Xbit_r29_c177 bl[177] br[177] wl[29] vdd gnd cell_6t
Xbit_r30_c177 bl[177] br[177] wl[30] vdd gnd cell_6t
Xbit_r31_c177 bl[177] br[177] wl[31] vdd gnd cell_6t
Xbit_r32_c177 bl[177] br[177] wl[32] vdd gnd cell_6t
Xbit_r33_c177 bl[177] br[177] wl[33] vdd gnd cell_6t
Xbit_r34_c177 bl[177] br[177] wl[34] vdd gnd cell_6t
Xbit_r35_c177 bl[177] br[177] wl[35] vdd gnd cell_6t
Xbit_r36_c177 bl[177] br[177] wl[36] vdd gnd cell_6t
Xbit_r37_c177 bl[177] br[177] wl[37] vdd gnd cell_6t
Xbit_r38_c177 bl[177] br[177] wl[38] vdd gnd cell_6t
Xbit_r39_c177 bl[177] br[177] wl[39] vdd gnd cell_6t
Xbit_r40_c177 bl[177] br[177] wl[40] vdd gnd cell_6t
Xbit_r41_c177 bl[177] br[177] wl[41] vdd gnd cell_6t
Xbit_r42_c177 bl[177] br[177] wl[42] vdd gnd cell_6t
Xbit_r43_c177 bl[177] br[177] wl[43] vdd gnd cell_6t
Xbit_r44_c177 bl[177] br[177] wl[44] vdd gnd cell_6t
Xbit_r45_c177 bl[177] br[177] wl[45] vdd gnd cell_6t
Xbit_r46_c177 bl[177] br[177] wl[46] vdd gnd cell_6t
Xbit_r47_c177 bl[177] br[177] wl[47] vdd gnd cell_6t
Xbit_r48_c177 bl[177] br[177] wl[48] vdd gnd cell_6t
Xbit_r49_c177 bl[177] br[177] wl[49] vdd gnd cell_6t
Xbit_r50_c177 bl[177] br[177] wl[50] vdd gnd cell_6t
Xbit_r51_c177 bl[177] br[177] wl[51] vdd gnd cell_6t
Xbit_r52_c177 bl[177] br[177] wl[52] vdd gnd cell_6t
Xbit_r53_c177 bl[177] br[177] wl[53] vdd gnd cell_6t
Xbit_r54_c177 bl[177] br[177] wl[54] vdd gnd cell_6t
Xbit_r55_c177 bl[177] br[177] wl[55] vdd gnd cell_6t
Xbit_r56_c177 bl[177] br[177] wl[56] vdd gnd cell_6t
Xbit_r57_c177 bl[177] br[177] wl[57] vdd gnd cell_6t
Xbit_r58_c177 bl[177] br[177] wl[58] vdd gnd cell_6t
Xbit_r59_c177 bl[177] br[177] wl[59] vdd gnd cell_6t
Xbit_r60_c177 bl[177] br[177] wl[60] vdd gnd cell_6t
Xbit_r61_c177 bl[177] br[177] wl[61] vdd gnd cell_6t
Xbit_r62_c177 bl[177] br[177] wl[62] vdd gnd cell_6t
Xbit_r63_c177 bl[177] br[177] wl[63] vdd gnd cell_6t
Xbit_r64_c177 bl[177] br[177] wl[64] vdd gnd cell_6t
Xbit_r65_c177 bl[177] br[177] wl[65] vdd gnd cell_6t
Xbit_r66_c177 bl[177] br[177] wl[66] vdd gnd cell_6t
Xbit_r67_c177 bl[177] br[177] wl[67] vdd gnd cell_6t
Xbit_r68_c177 bl[177] br[177] wl[68] vdd gnd cell_6t
Xbit_r69_c177 bl[177] br[177] wl[69] vdd gnd cell_6t
Xbit_r70_c177 bl[177] br[177] wl[70] vdd gnd cell_6t
Xbit_r71_c177 bl[177] br[177] wl[71] vdd gnd cell_6t
Xbit_r72_c177 bl[177] br[177] wl[72] vdd gnd cell_6t
Xbit_r73_c177 bl[177] br[177] wl[73] vdd gnd cell_6t
Xbit_r74_c177 bl[177] br[177] wl[74] vdd gnd cell_6t
Xbit_r75_c177 bl[177] br[177] wl[75] vdd gnd cell_6t
Xbit_r76_c177 bl[177] br[177] wl[76] vdd gnd cell_6t
Xbit_r77_c177 bl[177] br[177] wl[77] vdd gnd cell_6t
Xbit_r78_c177 bl[177] br[177] wl[78] vdd gnd cell_6t
Xbit_r79_c177 bl[177] br[177] wl[79] vdd gnd cell_6t
Xbit_r80_c177 bl[177] br[177] wl[80] vdd gnd cell_6t
Xbit_r81_c177 bl[177] br[177] wl[81] vdd gnd cell_6t
Xbit_r82_c177 bl[177] br[177] wl[82] vdd gnd cell_6t
Xbit_r83_c177 bl[177] br[177] wl[83] vdd gnd cell_6t
Xbit_r84_c177 bl[177] br[177] wl[84] vdd gnd cell_6t
Xbit_r85_c177 bl[177] br[177] wl[85] vdd gnd cell_6t
Xbit_r86_c177 bl[177] br[177] wl[86] vdd gnd cell_6t
Xbit_r87_c177 bl[177] br[177] wl[87] vdd gnd cell_6t
Xbit_r88_c177 bl[177] br[177] wl[88] vdd gnd cell_6t
Xbit_r89_c177 bl[177] br[177] wl[89] vdd gnd cell_6t
Xbit_r90_c177 bl[177] br[177] wl[90] vdd gnd cell_6t
Xbit_r91_c177 bl[177] br[177] wl[91] vdd gnd cell_6t
Xbit_r92_c177 bl[177] br[177] wl[92] vdd gnd cell_6t
Xbit_r93_c177 bl[177] br[177] wl[93] vdd gnd cell_6t
Xbit_r94_c177 bl[177] br[177] wl[94] vdd gnd cell_6t
Xbit_r95_c177 bl[177] br[177] wl[95] vdd gnd cell_6t
Xbit_r96_c177 bl[177] br[177] wl[96] vdd gnd cell_6t
Xbit_r97_c177 bl[177] br[177] wl[97] vdd gnd cell_6t
Xbit_r98_c177 bl[177] br[177] wl[98] vdd gnd cell_6t
Xbit_r99_c177 bl[177] br[177] wl[99] vdd gnd cell_6t
Xbit_r100_c177 bl[177] br[177] wl[100] vdd gnd cell_6t
Xbit_r101_c177 bl[177] br[177] wl[101] vdd gnd cell_6t
Xbit_r102_c177 bl[177] br[177] wl[102] vdd gnd cell_6t
Xbit_r103_c177 bl[177] br[177] wl[103] vdd gnd cell_6t
Xbit_r104_c177 bl[177] br[177] wl[104] vdd gnd cell_6t
Xbit_r105_c177 bl[177] br[177] wl[105] vdd gnd cell_6t
Xbit_r106_c177 bl[177] br[177] wl[106] vdd gnd cell_6t
Xbit_r107_c177 bl[177] br[177] wl[107] vdd gnd cell_6t
Xbit_r108_c177 bl[177] br[177] wl[108] vdd gnd cell_6t
Xbit_r109_c177 bl[177] br[177] wl[109] vdd gnd cell_6t
Xbit_r110_c177 bl[177] br[177] wl[110] vdd gnd cell_6t
Xbit_r111_c177 bl[177] br[177] wl[111] vdd gnd cell_6t
Xbit_r112_c177 bl[177] br[177] wl[112] vdd gnd cell_6t
Xbit_r113_c177 bl[177] br[177] wl[113] vdd gnd cell_6t
Xbit_r114_c177 bl[177] br[177] wl[114] vdd gnd cell_6t
Xbit_r115_c177 bl[177] br[177] wl[115] vdd gnd cell_6t
Xbit_r116_c177 bl[177] br[177] wl[116] vdd gnd cell_6t
Xbit_r117_c177 bl[177] br[177] wl[117] vdd gnd cell_6t
Xbit_r118_c177 bl[177] br[177] wl[118] vdd gnd cell_6t
Xbit_r119_c177 bl[177] br[177] wl[119] vdd gnd cell_6t
Xbit_r120_c177 bl[177] br[177] wl[120] vdd gnd cell_6t
Xbit_r121_c177 bl[177] br[177] wl[121] vdd gnd cell_6t
Xbit_r122_c177 bl[177] br[177] wl[122] vdd gnd cell_6t
Xbit_r123_c177 bl[177] br[177] wl[123] vdd gnd cell_6t
Xbit_r124_c177 bl[177] br[177] wl[124] vdd gnd cell_6t
Xbit_r125_c177 bl[177] br[177] wl[125] vdd gnd cell_6t
Xbit_r126_c177 bl[177] br[177] wl[126] vdd gnd cell_6t
Xbit_r127_c177 bl[177] br[177] wl[127] vdd gnd cell_6t
Xbit_r128_c177 bl[177] br[177] wl[128] vdd gnd cell_6t
Xbit_r129_c177 bl[177] br[177] wl[129] vdd gnd cell_6t
Xbit_r130_c177 bl[177] br[177] wl[130] vdd gnd cell_6t
Xbit_r131_c177 bl[177] br[177] wl[131] vdd gnd cell_6t
Xbit_r132_c177 bl[177] br[177] wl[132] vdd gnd cell_6t
Xbit_r133_c177 bl[177] br[177] wl[133] vdd gnd cell_6t
Xbit_r134_c177 bl[177] br[177] wl[134] vdd gnd cell_6t
Xbit_r135_c177 bl[177] br[177] wl[135] vdd gnd cell_6t
Xbit_r136_c177 bl[177] br[177] wl[136] vdd gnd cell_6t
Xbit_r137_c177 bl[177] br[177] wl[137] vdd gnd cell_6t
Xbit_r138_c177 bl[177] br[177] wl[138] vdd gnd cell_6t
Xbit_r139_c177 bl[177] br[177] wl[139] vdd gnd cell_6t
Xbit_r140_c177 bl[177] br[177] wl[140] vdd gnd cell_6t
Xbit_r141_c177 bl[177] br[177] wl[141] vdd gnd cell_6t
Xbit_r142_c177 bl[177] br[177] wl[142] vdd gnd cell_6t
Xbit_r143_c177 bl[177] br[177] wl[143] vdd gnd cell_6t
Xbit_r144_c177 bl[177] br[177] wl[144] vdd gnd cell_6t
Xbit_r145_c177 bl[177] br[177] wl[145] vdd gnd cell_6t
Xbit_r146_c177 bl[177] br[177] wl[146] vdd gnd cell_6t
Xbit_r147_c177 bl[177] br[177] wl[147] vdd gnd cell_6t
Xbit_r148_c177 bl[177] br[177] wl[148] vdd gnd cell_6t
Xbit_r149_c177 bl[177] br[177] wl[149] vdd gnd cell_6t
Xbit_r150_c177 bl[177] br[177] wl[150] vdd gnd cell_6t
Xbit_r151_c177 bl[177] br[177] wl[151] vdd gnd cell_6t
Xbit_r152_c177 bl[177] br[177] wl[152] vdd gnd cell_6t
Xbit_r153_c177 bl[177] br[177] wl[153] vdd gnd cell_6t
Xbit_r154_c177 bl[177] br[177] wl[154] vdd gnd cell_6t
Xbit_r155_c177 bl[177] br[177] wl[155] vdd gnd cell_6t
Xbit_r156_c177 bl[177] br[177] wl[156] vdd gnd cell_6t
Xbit_r157_c177 bl[177] br[177] wl[157] vdd gnd cell_6t
Xbit_r158_c177 bl[177] br[177] wl[158] vdd gnd cell_6t
Xbit_r159_c177 bl[177] br[177] wl[159] vdd gnd cell_6t
Xbit_r160_c177 bl[177] br[177] wl[160] vdd gnd cell_6t
Xbit_r161_c177 bl[177] br[177] wl[161] vdd gnd cell_6t
Xbit_r162_c177 bl[177] br[177] wl[162] vdd gnd cell_6t
Xbit_r163_c177 bl[177] br[177] wl[163] vdd gnd cell_6t
Xbit_r164_c177 bl[177] br[177] wl[164] vdd gnd cell_6t
Xbit_r165_c177 bl[177] br[177] wl[165] vdd gnd cell_6t
Xbit_r166_c177 bl[177] br[177] wl[166] vdd gnd cell_6t
Xbit_r167_c177 bl[177] br[177] wl[167] vdd gnd cell_6t
Xbit_r168_c177 bl[177] br[177] wl[168] vdd gnd cell_6t
Xbit_r169_c177 bl[177] br[177] wl[169] vdd gnd cell_6t
Xbit_r170_c177 bl[177] br[177] wl[170] vdd gnd cell_6t
Xbit_r171_c177 bl[177] br[177] wl[171] vdd gnd cell_6t
Xbit_r172_c177 bl[177] br[177] wl[172] vdd gnd cell_6t
Xbit_r173_c177 bl[177] br[177] wl[173] vdd gnd cell_6t
Xbit_r174_c177 bl[177] br[177] wl[174] vdd gnd cell_6t
Xbit_r175_c177 bl[177] br[177] wl[175] vdd gnd cell_6t
Xbit_r176_c177 bl[177] br[177] wl[176] vdd gnd cell_6t
Xbit_r177_c177 bl[177] br[177] wl[177] vdd gnd cell_6t
Xbit_r178_c177 bl[177] br[177] wl[178] vdd gnd cell_6t
Xbit_r179_c177 bl[177] br[177] wl[179] vdd gnd cell_6t
Xbit_r180_c177 bl[177] br[177] wl[180] vdd gnd cell_6t
Xbit_r181_c177 bl[177] br[177] wl[181] vdd gnd cell_6t
Xbit_r182_c177 bl[177] br[177] wl[182] vdd gnd cell_6t
Xbit_r183_c177 bl[177] br[177] wl[183] vdd gnd cell_6t
Xbit_r184_c177 bl[177] br[177] wl[184] vdd gnd cell_6t
Xbit_r185_c177 bl[177] br[177] wl[185] vdd gnd cell_6t
Xbit_r186_c177 bl[177] br[177] wl[186] vdd gnd cell_6t
Xbit_r187_c177 bl[177] br[177] wl[187] vdd gnd cell_6t
Xbit_r188_c177 bl[177] br[177] wl[188] vdd gnd cell_6t
Xbit_r189_c177 bl[177] br[177] wl[189] vdd gnd cell_6t
Xbit_r190_c177 bl[177] br[177] wl[190] vdd gnd cell_6t
Xbit_r191_c177 bl[177] br[177] wl[191] vdd gnd cell_6t
Xbit_r192_c177 bl[177] br[177] wl[192] vdd gnd cell_6t
Xbit_r193_c177 bl[177] br[177] wl[193] vdd gnd cell_6t
Xbit_r194_c177 bl[177] br[177] wl[194] vdd gnd cell_6t
Xbit_r195_c177 bl[177] br[177] wl[195] vdd gnd cell_6t
Xbit_r196_c177 bl[177] br[177] wl[196] vdd gnd cell_6t
Xbit_r197_c177 bl[177] br[177] wl[197] vdd gnd cell_6t
Xbit_r198_c177 bl[177] br[177] wl[198] vdd gnd cell_6t
Xbit_r199_c177 bl[177] br[177] wl[199] vdd gnd cell_6t
Xbit_r200_c177 bl[177] br[177] wl[200] vdd gnd cell_6t
Xbit_r201_c177 bl[177] br[177] wl[201] vdd gnd cell_6t
Xbit_r202_c177 bl[177] br[177] wl[202] vdd gnd cell_6t
Xbit_r203_c177 bl[177] br[177] wl[203] vdd gnd cell_6t
Xbit_r204_c177 bl[177] br[177] wl[204] vdd gnd cell_6t
Xbit_r205_c177 bl[177] br[177] wl[205] vdd gnd cell_6t
Xbit_r206_c177 bl[177] br[177] wl[206] vdd gnd cell_6t
Xbit_r207_c177 bl[177] br[177] wl[207] vdd gnd cell_6t
Xbit_r208_c177 bl[177] br[177] wl[208] vdd gnd cell_6t
Xbit_r209_c177 bl[177] br[177] wl[209] vdd gnd cell_6t
Xbit_r210_c177 bl[177] br[177] wl[210] vdd gnd cell_6t
Xbit_r211_c177 bl[177] br[177] wl[211] vdd gnd cell_6t
Xbit_r212_c177 bl[177] br[177] wl[212] vdd gnd cell_6t
Xbit_r213_c177 bl[177] br[177] wl[213] vdd gnd cell_6t
Xbit_r214_c177 bl[177] br[177] wl[214] vdd gnd cell_6t
Xbit_r215_c177 bl[177] br[177] wl[215] vdd gnd cell_6t
Xbit_r216_c177 bl[177] br[177] wl[216] vdd gnd cell_6t
Xbit_r217_c177 bl[177] br[177] wl[217] vdd gnd cell_6t
Xbit_r218_c177 bl[177] br[177] wl[218] vdd gnd cell_6t
Xbit_r219_c177 bl[177] br[177] wl[219] vdd gnd cell_6t
Xbit_r220_c177 bl[177] br[177] wl[220] vdd gnd cell_6t
Xbit_r221_c177 bl[177] br[177] wl[221] vdd gnd cell_6t
Xbit_r222_c177 bl[177] br[177] wl[222] vdd gnd cell_6t
Xbit_r223_c177 bl[177] br[177] wl[223] vdd gnd cell_6t
Xbit_r224_c177 bl[177] br[177] wl[224] vdd gnd cell_6t
Xbit_r225_c177 bl[177] br[177] wl[225] vdd gnd cell_6t
Xbit_r226_c177 bl[177] br[177] wl[226] vdd gnd cell_6t
Xbit_r227_c177 bl[177] br[177] wl[227] vdd gnd cell_6t
Xbit_r228_c177 bl[177] br[177] wl[228] vdd gnd cell_6t
Xbit_r229_c177 bl[177] br[177] wl[229] vdd gnd cell_6t
Xbit_r230_c177 bl[177] br[177] wl[230] vdd gnd cell_6t
Xbit_r231_c177 bl[177] br[177] wl[231] vdd gnd cell_6t
Xbit_r232_c177 bl[177] br[177] wl[232] vdd gnd cell_6t
Xbit_r233_c177 bl[177] br[177] wl[233] vdd gnd cell_6t
Xbit_r234_c177 bl[177] br[177] wl[234] vdd gnd cell_6t
Xbit_r235_c177 bl[177] br[177] wl[235] vdd gnd cell_6t
Xbit_r236_c177 bl[177] br[177] wl[236] vdd gnd cell_6t
Xbit_r237_c177 bl[177] br[177] wl[237] vdd gnd cell_6t
Xbit_r238_c177 bl[177] br[177] wl[238] vdd gnd cell_6t
Xbit_r239_c177 bl[177] br[177] wl[239] vdd gnd cell_6t
Xbit_r240_c177 bl[177] br[177] wl[240] vdd gnd cell_6t
Xbit_r241_c177 bl[177] br[177] wl[241] vdd gnd cell_6t
Xbit_r242_c177 bl[177] br[177] wl[242] vdd gnd cell_6t
Xbit_r243_c177 bl[177] br[177] wl[243] vdd gnd cell_6t
Xbit_r244_c177 bl[177] br[177] wl[244] vdd gnd cell_6t
Xbit_r245_c177 bl[177] br[177] wl[245] vdd gnd cell_6t
Xbit_r246_c177 bl[177] br[177] wl[246] vdd gnd cell_6t
Xbit_r247_c177 bl[177] br[177] wl[247] vdd gnd cell_6t
Xbit_r248_c177 bl[177] br[177] wl[248] vdd gnd cell_6t
Xbit_r249_c177 bl[177] br[177] wl[249] vdd gnd cell_6t
Xbit_r250_c177 bl[177] br[177] wl[250] vdd gnd cell_6t
Xbit_r251_c177 bl[177] br[177] wl[251] vdd gnd cell_6t
Xbit_r252_c177 bl[177] br[177] wl[252] vdd gnd cell_6t
Xbit_r253_c177 bl[177] br[177] wl[253] vdd gnd cell_6t
Xbit_r254_c177 bl[177] br[177] wl[254] vdd gnd cell_6t
Xbit_r255_c177 bl[177] br[177] wl[255] vdd gnd cell_6t
Xbit_r0_c178 bl[178] br[178] wl[0] vdd gnd cell_6t
Xbit_r1_c178 bl[178] br[178] wl[1] vdd gnd cell_6t
Xbit_r2_c178 bl[178] br[178] wl[2] vdd gnd cell_6t
Xbit_r3_c178 bl[178] br[178] wl[3] vdd gnd cell_6t
Xbit_r4_c178 bl[178] br[178] wl[4] vdd gnd cell_6t
Xbit_r5_c178 bl[178] br[178] wl[5] vdd gnd cell_6t
Xbit_r6_c178 bl[178] br[178] wl[6] vdd gnd cell_6t
Xbit_r7_c178 bl[178] br[178] wl[7] vdd gnd cell_6t
Xbit_r8_c178 bl[178] br[178] wl[8] vdd gnd cell_6t
Xbit_r9_c178 bl[178] br[178] wl[9] vdd gnd cell_6t
Xbit_r10_c178 bl[178] br[178] wl[10] vdd gnd cell_6t
Xbit_r11_c178 bl[178] br[178] wl[11] vdd gnd cell_6t
Xbit_r12_c178 bl[178] br[178] wl[12] vdd gnd cell_6t
Xbit_r13_c178 bl[178] br[178] wl[13] vdd gnd cell_6t
Xbit_r14_c178 bl[178] br[178] wl[14] vdd gnd cell_6t
Xbit_r15_c178 bl[178] br[178] wl[15] vdd gnd cell_6t
Xbit_r16_c178 bl[178] br[178] wl[16] vdd gnd cell_6t
Xbit_r17_c178 bl[178] br[178] wl[17] vdd gnd cell_6t
Xbit_r18_c178 bl[178] br[178] wl[18] vdd gnd cell_6t
Xbit_r19_c178 bl[178] br[178] wl[19] vdd gnd cell_6t
Xbit_r20_c178 bl[178] br[178] wl[20] vdd gnd cell_6t
Xbit_r21_c178 bl[178] br[178] wl[21] vdd gnd cell_6t
Xbit_r22_c178 bl[178] br[178] wl[22] vdd gnd cell_6t
Xbit_r23_c178 bl[178] br[178] wl[23] vdd gnd cell_6t
Xbit_r24_c178 bl[178] br[178] wl[24] vdd gnd cell_6t
Xbit_r25_c178 bl[178] br[178] wl[25] vdd gnd cell_6t
Xbit_r26_c178 bl[178] br[178] wl[26] vdd gnd cell_6t
Xbit_r27_c178 bl[178] br[178] wl[27] vdd gnd cell_6t
Xbit_r28_c178 bl[178] br[178] wl[28] vdd gnd cell_6t
Xbit_r29_c178 bl[178] br[178] wl[29] vdd gnd cell_6t
Xbit_r30_c178 bl[178] br[178] wl[30] vdd gnd cell_6t
Xbit_r31_c178 bl[178] br[178] wl[31] vdd gnd cell_6t
Xbit_r32_c178 bl[178] br[178] wl[32] vdd gnd cell_6t
Xbit_r33_c178 bl[178] br[178] wl[33] vdd gnd cell_6t
Xbit_r34_c178 bl[178] br[178] wl[34] vdd gnd cell_6t
Xbit_r35_c178 bl[178] br[178] wl[35] vdd gnd cell_6t
Xbit_r36_c178 bl[178] br[178] wl[36] vdd gnd cell_6t
Xbit_r37_c178 bl[178] br[178] wl[37] vdd gnd cell_6t
Xbit_r38_c178 bl[178] br[178] wl[38] vdd gnd cell_6t
Xbit_r39_c178 bl[178] br[178] wl[39] vdd gnd cell_6t
Xbit_r40_c178 bl[178] br[178] wl[40] vdd gnd cell_6t
Xbit_r41_c178 bl[178] br[178] wl[41] vdd gnd cell_6t
Xbit_r42_c178 bl[178] br[178] wl[42] vdd gnd cell_6t
Xbit_r43_c178 bl[178] br[178] wl[43] vdd gnd cell_6t
Xbit_r44_c178 bl[178] br[178] wl[44] vdd gnd cell_6t
Xbit_r45_c178 bl[178] br[178] wl[45] vdd gnd cell_6t
Xbit_r46_c178 bl[178] br[178] wl[46] vdd gnd cell_6t
Xbit_r47_c178 bl[178] br[178] wl[47] vdd gnd cell_6t
Xbit_r48_c178 bl[178] br[178] wl[48] vdd gnd cell_6t
Xbit_r49_c178 bl[178] br[178] wl[49] vdd gnd cell_6t
Xbit_r50_c178 bl[178] br[178] wl[50] vdd gnd cell_6t
Xbit_r51_c178 bl[178] br[178] wl[51] vdd gnd cell_6t
Xbit_r52_c178 bl[178] br[178] wl[52] vdd gnd cell_6t
Xbit_r53_c178 bl[178] br[178] wl[53] vdd gnd cell_6t
Xbit_r54_c178 bl[178] br[178] wl[54] vdd gnd cell_6t
Xbit_r55_c178 bl[178] br[178] wl[55] vdd gnd cell_6t
Xbit_r56_c178 bl[178] br[178] wl[56] vdd gnd cell_6t
Xbit_r57_c178 bl[178] br[178] wl[57] vdd gnd cell_6t
Xbit_r58_c178 bl[178] br[178] wl[58] vdd gnd cell_6t
Xbit_r59_c178 bl[178] br[178] wl[59] vdd gnd cell_6t
Xbit_r60_c178 bl[178] br[178] wl[60] vdd gnd cell_6t
Xbit_r61_c178 bl[178] br[178] wl[61] vdd gnd cell_6t
Xbit_r62_c178 bl[178] br[178] wl[62] vdd gnd cell_6t
Xbit_r63_c178 bl[178] br[178] wl[63] vdd gnd cell_6t
Xbit_r64_c178 bl[178] br[178] wl[64] vdd gnd cell_6t
Xbit_r65_c178 bl[178] br[178] wl[65] vdd gnd cell_6t
Xbit_r66_c178 bl[178] br[178] wl[66] vdd gnd cell_6t
Xbit_r67_c178 bl[178] br[178] wl[67] vdd gnd cell_6t
Xbit_r68_c178 bl[178] br[178] wl[68] vdd gnd cell_6t
Xbit_r69_c178 bl[178] br[178] wl[69] vdd gnd cell_6t
Xbit_r70_c178 bl[178] br[178] wl[70] vdd gnd cell_6t
Xbit_r71_c178 bl[178] br[178] wl[71] vdd gnd cell_6t
Xbit_r72_c178 bl[178] br[178] wl[72] vdd gnd cell_6t
Xbit_r73_c178 bl[178] br[178] wl[73] vdd gnd cell_6t
Xbit_r74_c178 bl[178] br[178] wl[74] vdd gnd cell_6t
Xbit_r75_c178 bl[178] br[178] wl[75] vdd gnd cell_6t
Xbit_r76_c178 bl[178] br[178] wl[76] vdd gnd cell_6t
Xbit_r77_c178 bl[178] br[178] wl[77] vdd gnd cell_6t
Xbit_r78_c178 bl[178] br[178] wl[78] vdd gnd cell_6t
Xbit_r79_c178 bl[178] br[178] wl[79] vdd gnd cell_6t
Xbit_r80_c178 bl[178] br[178] wl[80] vdd gnd cell_6t
Xbit_r81_c178 bl[178] br[178] wl[81] vdd gnd cell_6t
Xbit_r82_c178 bl[178] br[178] wl[82] vdd gnd cell_6t
Xbit_r83_c178 bl[178] br[178] wl[83] vdd gnd cell_6t
Xbit_r84_c178 bl[178] br[178] wl[84] vdd gnd cell_6t
Xbit_r85_c178 bl[178] br[178] wl[85] vdd gnd cell_6t
Xbit_r86_c178 bl[178] br[178] wl[86] vdd gnd cell_6t
Xbit_r87_c178 bl[178] br[178] wl[87] vdd gnd cell_6t
Xbit_r88_c178 bl[178] br[178] wl[88] vdd gnd cell_6t
Xbit_r89_c178 bl[178] br[178] wl[89] vdd gnd cell_6t
Xbit_r90_c178 bl[178] br[178] wl[90] vdd gnd cell_6t
Xbit_r91_c178 bl[178] br[178] wl[91] vdd gnd cell_6t
Xbit_r92_c178 bl[178] br[178] wl[92] vdd gnd cell_6t
Xbit_r93_c178 bl[178] br[178] wl[93] vdd gnd cell_6t
Xbit_r94_c178 bl[178] br[178] wl[94] vdd gnd cell_6t
Xbit_r95_c178 bl[178] br[178] wl[95] vdd gnd cell_6t
Xbit_r96_c178 bl[178] br[178] wl[96] vdd gnd cell_6t
Xbit_r97_c178 bl[178] br[178] wl[97] vdd gnd cell_6t
Xbit_r98_c178 bl[178] br[178] wl[98] vdd gnd cell_6t
Xbit_r99_c178 bl[178] br[178] wl[99] vdd gnd cell_6t
Xbit_r100_c178 bl[178] br[178] wl[100] vdd gnd cell_6t
Xbit_r101_c178 bl[178] br[178] wl[101] vdd gnd cell_6t
Xbit_r102_c178 bl[178] br[178] wl[102] vdd gnd cell_6t
Xbit_r103_c178 bl[178] br[178] wl[103] vdd gnd cell_6t
Xbit_r104_c178 bl[178] br[178] wl[104] vdd gnd cell_6t
Xbit_r105_c178 bl[178] br[178] wl[105] vdd gnd cell_6t
Xbit_r106_c178 bl[178] br[178] wl[106] vdd gnd cell_6t
Xbit_r107_c178 bl[178] br[178] wl[107] vdd gnd cell_6t
Xbit_r108_c178 bl[178] br[178] wl[108] vdd gnd cell_6t
Xbit_r109_c178 bl[178] br[178] wl[109] vdd gnd cell_6t
Xbit_r110_c178 bl[178] br[178] wl[110] vdd gnd cell_6t
Xbit_r111_c178 bl[178] br[178] wl[111] vdd gnd cell_6t
Xbit_r112_c178 bl[178] br[178] wl[112] vdd gnd cell_6t
Xbit_r113_c178 bl[178] br[178] wl[113] vdd gnd cell_6t
Xbit_r114_c178 bl[178] br[178] wl[114] vdd gnd cell_6t
Xbit_r115_c178 bl[178] br[178] wl[115] vdd gnd cell_6t
Xbit_r116_c178 bl[178] br[178] wl[116] vdd gnd cell_6t
Xbit_r117_c178 bl[178] br[178] wl[117] vdd gnd cell_6t
Xbit_r118_c178 bl[178] br[178] wl[118] vdd gnd cell_6t
Xbit_r119_c178 bl[178] br[178] wl[119] vdd gnd cell_6t
Xbit_r120_c178 bl[178] br[178] wl[120] vdd gnd cell_6t
Xbit_r121_c178 bl[178] br[178] wl[121] vdd gnd cell_6t
Xbit_r122_c178 bl[178] br[178] wl[122] vdd gnd cell_6t
Xbit_r123_c178 bl[178] br[178] wl[123] vdd gnd cell_6t
Xbit_r124_c178 bl[178] br[178] wl[124] vdd gnd cell_6t
Xbit_r125_c178 bl[178] br[178] wl[125] vdd gnd cell_6t
Xbit_r126_c178 bl[178] br[178] wl[126] vdd gnd cell_6t
Xbit_r127_c178 bl[178] br[178] wl[127] vdd gnd cell_6t
Xbit_r128_c178 bl[178] br[178] wl[128] vdd gnd cell_6t
Xbit_r129_c178 bl[178] br[178] wl[129] vdd gnd cell_6t
Xbit_r130_c178 bl[178] br[178] wl[130] vdd gnd cell_6t
Xbit_r131_c178 bl[178] br[178] wl[131] vdd gnd cell_6t
Xbit_r132_c178 bl[178] br[178] wl[132] vdd gnd cell_6t
Xbit_r133_c178 bl[178] br[178] wl[133] vdd gnd cell_6t
Xbit_r134_c178 bl[178] br[178] wl[134] vdd gnd cell_6t
Xbit_r135_c178 bl[178] br[178] wl[135] vdd gnd cell_6t
Xbit_r136_c178 bl[178] br[178] wl[136] vdd gnd cell_6t
Xbit_r137_c178 bl[178] br[178] wl[137] vdd gnd cell_6t
Xbit_r138_c178 bl[178] br[178] wl[138] vdd gnd cell_6t
Xbit_r139_c178 bl[178] br[178] wl[139] vdd gnd cell_6t
Xbit_r140_c178 bl[178] br[178] wl[140] vdd gnd cell_6t
Xbit_r141_c178 bl[178] br[178] wl[141] vdd gnd cell_6t
Xbit_r142_c178 bl[178] br[178] wl[142] vdd gnd cell_6t
Xbit_r143_c178 bl[178] br[178] wl[143] vdd gnd cell_6t
Xbit_r144_c178 bl[178] br[178] wl[144] vdd gnd cell_6t
Xbit_r145_c178 bl[178] br[178] wl[145] vdd gnd cell_6t
Xbit_r146_c178 bl[178] br[178] wl[146] vdd gnd cell_6t
Xbit_r147_c178 bl[178] br[178] wl[147] vdd gnd cell_6t
Xbit_r148_c178 bl[178] br[178] wl[148] vdd gnd cell_6t
Xbit_r149_c178 bl[178] br[178] wl[149] vdd gnd cell_6t
Xbit_r150_c178 bl[178] br[178] wl[150] vdd gnd cell_6t
Xbit_r151_c178 bl[178] br[178] wl[151] vdd gnd cell_6t
Xbit_r152_c178 bl[178] br[178] wl[152] vdd gnd cell_6t
Xbit_r153_c178 bl[178] br[178] wl[153] vdd gnd cell_6t
Xbit_r154_c178 bl[178] br[178] wl[154] vdd gnd cell_6t
Xbit_r155_c178 bl[178] br[178] wl[155] vdd gnd cell_6t
Xbit_r156_c178 bl[178] br[178] wl[156] vdd gnd cell_6t
Xbit_r157_c178 bl[178] br[178] wl[157] vdd gnd cell_6t
Xbit_r158_c178 bl[178] br[178] wl[158] vdd gnd cell_6t
Xbit_r159_c178 bl[178] br[178] wl[159] vdd gnd cell_6t
Xbit_r160_c178 bl[178] br[178] wl[160] vdd gnd cell_6t
Xbit_r161_c178 bl[178] br[178] wl[161] vdd gnd cell_6t
Xbit_r162_c178 bl[178] br[178] wl[162] vdd gnd cell_6t
Xbit_r163_c178 bl[178] br[178] wl[163] vdd gnd cell_6t
Xbit_r164_c178 bl[178] br[178] wl[164] vdd gnd cell_6t
Xbit_r165_c178 bl[178] br[178] wl[165] vdd gnd cell_6t
Xbit_r166_c178 bl[178] br[178] wl[166] vdd gnd cell_6t
Xbit_r167_c178 bl[178] br[178] wl[167] vdd gnd cell_6t
Xbit_r168_c178 bl[178] br[178] wl[168] vdd gnd cell_6t
Xbit_r169_c178 bl[178] br[178] wl[169] vdd gnd cell_6t
Xbit_r170_c178 bl[178] br[178] wl[170] vdd gnd cell_6t
Xbit_r171_c178 bl[178] br[178] wl[171] vdd gnd cell_6t
Xbit_r172_c178 bl[178] br[178] wl[172] vdd gnd cell_6t
Xbit_r173_c178 bl[178] br[178] wl[173] vdd gnd cell_6t
Xbit_r174_c178 bl[178] br[178] wl[174] vdd gnd cell_6t
Xbit_r175_c178 bl[178] br[178] wl[175] vdd gnd cell_6t
Xbit_r176_c178 bl[178] br[178] wl[176] vdd gnd cell_6t
Xbit_r177_c178 bl[178] br[178] wl[177] vdd gnd cell_6t
Xbit_r178_c178 bl[178] br[178] wl[178] vdd gnd cell_6t
Xbit_r179_c178 bl[178] br[178] wl[179] vdd gnd cell_6t
Xbit_r180_c178 bl[178] br[178] wl[180] vdd gnd cell_6t
Xbit_r181_c178 bl[178] br[178] wl[181] vdd gnd cell_6t
Xbit_r182_c178 bl[178] br[178] wl[182] vdd gnd cell_6t
Xbit_r183_c178 bl[178] br[178] wl[183] vdd gnd cell_6t
Xbit_r184_c178 bl[178] br[178] wl[184] vdd gnd cell_6t
Xbit_r185_c178 bl[178] br[178] wl[185] vdd gnd cell_6t
Xbit_r186_c178 bl[178] br[178] wl[186] vdd gnd cell_6t
Xbit_r187_c178 bl[178] br[178] wl[187] vdd gnd cell_6t
Xbit_r188_c178 bl[178] br[178] wl[188] vdd gnd cell_6t
Xbit_r189_c178 bl[178] br[178] wl[189] vdd gnd cell_6t
Xbit_r190_c178 bl[178] br[178] wl[190] vdd gnd cell_6t
Xbit_r191_c178 bl[178] br[178] wl[191] vdd gnd cell_6t
Xbit_r192_c178 bl[178] br[178] wl[192] vdd gnd cell_6t
Xbit_r193_c178 bl[178] br[178] wl[193] vdd gnd cell_6t
Xbit_r194_c178 bl[178] br[178] wl[194] vdd gnd cell_6t
Xbit_r195_c178 bl[178] br[178] wl[195] vdd gnd cell_6t
Xbit_r196_c178 bl[178] br[178] wl[196] vdd gnd cell_6t
Xbit_r197_c178 bl[178] br[178] wl[197] vdd gnd cell_6t
Xbit_r198_c178 bl[178] br[178] wl[198] vdd gnd cell_6t
Xbit_r199_c178 bl[178] br[178] wl[199] vdd gnd cell_6t
Xbit_r200_c178 bl[178] br[178] wl[200] vdd gnd cell_6t
Xbit_r201_c178 bl[178] br[178] wl[201] vdd gnd cell_6t
Xbit_r202_c178 bl[178] br[178] wl[202] vdd gnd cell_6t
Xbit_r203_c178 bl[178] br[178] wl[203] vdd gnd cell_6t
Xbit_r204_c178 bl[178] br[178] wl[204] vdd gnd cell_6t
Xbit_r205_c178 bl[178] br[178] wl[205] vdd gnd cell_6t
Xbit_r206_c178 bl[178] br[178] wl[206] vdd gnd cell_6t
Xbit_r207_c178 bl[178] br[178] wl[207] vdd gnd cell_6t
Xbit_r208_c178 bl[178] br[178] wl[208] vdd gnd cell_6t
Xbit_r209_c178 bl[178] br[178] wl[209] vdd gnd cell_6t
Xbit_r210_c178 bl[178] br[178] wl[210] vdd gnd cell_6t
Xbit_r211_c178 bl[178] br[178] wl[211] vdd gnd cell_6t
Xbit_r212_c178 bl[178] br[178] wl[212] vdd gnd cell_6t
Xbit_r213_c178 bl[178] br[178] wl[213] vdd gnd cell_6t
Xbit_r214_c178 bl[178] br[178] wl[214] vdd gnd cell_6t
Xbit_r215_c178 bl[178] br[178] wl[215] vdd gnd cell_6t
Xbit_r216_c178 bl[178] br[178] wl[216] vdd gnd cell_6t
Xbit_r217_c178 bl[178] br[178] wl[217] vdd gnd cell_6t
Xbit_r218_c178 bl[178] br[178] wl[218] vdd gnd cell_6t
Xbit_r219_c178 bl[178] br[178] wl[219] vdd gnd cell_6t
Xbit_r220_c178 bl[178] br[178] wl[220] vdd gnd cell_6t
Xbit_r221_c178 bl[178] br[178] wl[221] vdd gnd cell_6t
Xbit_r222_c178 bl[178] br[178] wl[222] vdd gnd cell_6t
Xbit_r223_c178 bl[178] br[178] wl[223] vdd gnd cell_6t
Xbit_r224_c178 bl[178] br[178] wl[224] vdd gnd cell_6t
Xbit_r225_c178 bl[178] br[178] wl[225] vdd gnd cell_6t
Xbit_r226_c178 bl[178] br[178] wl[226] vdd gnd cell_6t
Xbit_r227_c178 bl[178] br[178] wl[227] vdd gnd cell_6t
Xbit_r228_c178 bl[178] br[178] wl[228] vdd gnd cell_6t
Xbit_r229_c178 bl[178] br[178] wl[229] vdd gnd cell_6t
Xbit_r230_c178 bl[178] br[178] wl[230] vdd gnd cell_6t
Xbit_r231_c178 bl[178] br[178] wl[231] vdd gnd cell_6t
Xbit_r232_c178 bl[178] br[178] wl[232] vdd gnd cell_6t
Xbit_r233_c178 bl[178] br[178] wl[233] vdd gnd cell_6t
Xbit_r234_c178 bl[178] br[178] wl[234] vdd gnd cell_6t
Xbit_r235_c178 bl[178] br[178] wl[235] vdd gnd cell_6t
Xbit_r236_c178 bl[178] br[178] wl[236] vdd gnd cell_6t
Xbit_r237_c178 bl[178] br[178] wl[237] vdd gnd cell_6t
Xbit_r238_c178 bl[178] br[178] wl[238] vdd gnd cell_6t
Xbit_r239_c178 bl[178] br[178] wl[239] vdd gnd cell_6t
Xbit_r240_c178 bl[178] br[178] wl[240] vdd gnd cell_6t
Xbit_r241_c178 bl[178] br[178] wl[241] vdd gnd cell_6t
Xbit_r242_c178 bl[178] br[178] wl[242] vdd gnd cell_6t
Xbit_r243_c178 bl[178] br[178] wl[243] vdd gnd cell_6t
Xbit_r244_c178 bl[178] br[178] wl[244] vdd gnd cell_6t
Xbit_r245_c178 bl[178] br[178] wl[245] vdd gnd cell_6t
Xbit_r246_c178 bl[178] br[178] wl[246] vdd gnd cell_6t
Xbit_r247_c178 bl[178] br[178] wl[247] vdd gnd cell_6t
Xbit_r248_c178 bl[178] br[178] wl[248] vdd gnd cell_6t
Xbit_r249_c178 bl[178] br[178] wl[249] vdd gnd cell_6t
Xbit_r250_c178 bl[178] br[178] wl[250] vdd gnd cell_6t
Xbit_r251_c178 bl[178] br[178] wl[251] vdd gnd cell_6t
Xbit_r252_c178 bl[178] br[178] wl[252] vdd gnd cell_6t
Xbit_r253_c178 bl[178] br[178] wl[253] vdd gnd cell_6t
Xbit_r254_c178 bl[178] br[178] wl[254] vdd gnd cell_6t
Xbit_r255_c178 bl[178] br[178] wl[255] vdd gnd cell_6t
Xbit_r0_c179 bl[179] br[179] wl[0] vdd gnd cell_6t
Xbit_r1_c179 bl[179] br[179] wl[1] vdd gnd cell_6t
Xbit_r2_c179 bl[179] br[179] wl[2] vdd gnd cell_6t
Xbit_r3_c179 bl[179] br[179] wl[3] vdd gnd cell_6t
Xbit_r4_c179 bl[179] br[179] wl[4] vdd gnd cell_6t
Xbit_r5_c179 bl[179] br[179] wl[5] vdd gnd cell_6t
Xbit_r6_c179 bl[179] br[179] wl[6] vdd gnd cell_6t
Xbit_r7_c179 bl[179] br[179] wl[7] vdd gnd cell_6t
Xbit_r8_c179 bl[179] br[179] wl[8] vdd gnd cell_6t
Xbit_r9_c179 bl[179] br[179] wl[9] vdd gnd cell_6t
Xbit_r10_c179 bl[179] br[179] wl[10] vdd gnd cell_6t
Xbit_r11_c179 bl[179] br[179] wl[11] vdd gnd cell_6t
Xbit_r12_c179 bl[179] br[179] wl[12] vdd gnd cell_6t
Xbit_r13_c179 bl[179] br[179] wl[13] vdd gnd cell_6t
Xbit_r14_c179 bl[179] br[179] wl[14] vdd gnd cell_6t
Xbit_r15_c179 bl[179] br[179] wl[15] vdd gnd cell_6t
Xbit_r16_c179 bl[179] br[179] wl[16] vdd gnd cell_6t
Xbit_r17_c179 bl[179] br[179] wl[17] vdd gnd cell_6t
Xbit_r18_c179 bl[179] br[179] wl[18] vdd gnd cell_6t
Xbit_r19_c179 bl[179] br[179] wl[19] vdd gnd cell_6t
Xbit_r20_c179 bl[179] br[179] wl[20] vdd gnd cell_6t
Xbit_r21_c179 bl[179] br[179] wl[21] vdd gnd cell_6t
Xbit_r22_c179 bl[179] br[179] wl[22] vdd gnd cell_6t
Xbit_r23_c179 bl[179] br[179] wl[23] vdd gnd cell_6t
Xbit_r24_c179 bl[179] br[179] wl[24] vdd gnd cell_6t
Xbit_r25_c179 bl[179] br[179] wl[25] vdd gnd cell_6t
Xbit_r26_c179 bl[179] br[179] wl[26] vdd gnd cell_6t
Xbit_r27_c179 bl[179] br[179] wl[27] vdd gnd cell_6t
Xbit_r28_c179 bl[179] br[179] wl[28] vdd gnd cell_6t
Xbit_r29_c179 bl[179] br[179] wl[29] vdd gnd cell_6t
Xbit_r30_c179 bl[179] br[179] wl[30] vdd gnd cell_6t
Xbit_r31_c179 bl[179] br[179] wl[31] vdd gnd cell_6t
Xbit_r32_c179 bl[179] br[179] wl[32] vdd gnd cell_6t
Xbit_r33_c179 bl[179] br[179] wl[33] vdd gnd cell_6t
Xbit_r34_c179 bl[179] br[179] wl[34] vdd gnd cell_6t
Xbit_r35_c179 bl[179] br[179] wl[35] vdd gnd cell_6t
Xbit_r36_c179 bl[179] br[179] wl[36] vdd gnd cell_6t
Xbit_r37_c179 bl[179] br[179] wl[37] vdd gnd cell_6t
Xbit_r38_c179 bl[179] br[179] wl[38] vdd gnd cell_6t
Xbit_r39_c179 bl[179] br[179] wl[39] vdd gnd cell_6t
Xbit_r40_c179 bl[179] br[179] wl[40] vdd gnd cell_6t
Xbit_r41_c179 bl[179] br[179] wl[41] vdd gnd cell_6t
Xbit_r42_c179 bl[179] br[179] wl[42] vdd gnd cell_6t
Xbit_r43_c179 bl[179] br[179] wl[43] vdd gnd cell_6t
Xbit_r44_c179 bl[179] br[179] wl[44] vdd gnd cell_6t
Xbit_r45_c179 bl[179] br[179] wl[45] vdd gnd cell_6t
Xbit_r46_c179 bl[179] br[179] wl[46] vdd gnd cell_6t
Xbit_r47_c179 bl[179] br[179] wl[47] vdd gnd cell_6t
Xbit_r48_c179 bl[179] br[179] wl[48] vdd gnd cell_6t
Xbit_r49_c179 bl[179] br[179] wl[49] vdd gnd cell_6t
Xbit_r50_c179 bl[179] br[179] wl[50] vdd gnd cell_6t
Xbit_r51_c179 bl[179] br[179] wl[51] vdd gnd cell_6t
Xbit_r52_c179 bl[179] br[179] wl[52] vdd gnd cell_6t
Xbit_r53_c179 bl[179] br[179] wl[53] vdd gnd cell_6t
Xbit_r54_c179 bl[179] br[179] wl[54] vdd gnd cell_6t
Xbit_r55_c179 bl[179] br[179] wl[55] vdd gnd cell_6t
Xbit_r56_c179 bl[179] br[179] wl[56] vdd gnd cell_6t
Xbit_r57_c179 bl[179] br[179] wl[57] vdd gnd cell_6t
Xbit_r58_c179 bl[179] br[179] wl[58] vdd gnd cell_6t
Xbit_r59_c179 bl[179] br[179] wl[59] vdd gnd cell_6t
Xbit_r60_c179 bl[179] br[179] wl[60] vdd gnd cell_6t
Xbit_r61_c179 bl[179] br[179] wl[61] vdd gnd cell_6t
Xbit_r62_c179 bl[179] br[179] wl[62] vdd gnd cell_6t
Xbit_r63_c179 bl[179] br[179] wl[63] vdd gnd cell_6t
Xbit_r64_c179 bl[179] br[179] wl[64] vdd gnd cell_6t
Xbit_r65_c179 bl[179] br[179] wl[65] vdd gnd cell_6t
Xbit_r66_c179 bl[179] br[179] wl[66] vdd gnd cell_6t
Xbit_r67_c179 bl[179] br[179] wl[67] vdd gnd cell_6t
Xbit_r68_c179 bl[179] br[179] wl[68] vdd gnd cell_6t
Xbit_r69_c179 bl[179] br[179] wl[69] vdd gnd cell_6t
Xbit_r70_c179 bl[179] br[179] wl[70] vdd gnd cell_6t
Xbit_r71_c179 bl[179] br[179] wl[71] vdd gnd cell_6t
Xbit_r72_c179 bl[179] br[179] wl[72] vdd gnd cell_6t
Xbit_r73_c179 bl[179] br[179] wl[73] vdd gnd cell_6t
Xbit_r74_c179 bl[179] br[179] wl[74] vdd gnd cell_6t
Xbit_r75_c179 bl[179] br[179] wl[75] vdd gnd cell_6t
Xbit_r76_c179 bl[179] br[179] wl[76] vdd gnd cell_6t
Xbit_r77_c179 bl[179] br[179] wl[77] vdd gnd cell_6t
Xbit_r78_c179 bl[179] br[179] wl[78] vdd gnd cell_6t
Xbit_r79_c179 bl[179] br[179] wl[79] vdd gnd cell_6t
Xbit_r80_c179 bl[179] br[179] wl[80] vdd gnd cell_6t
Xbit_r81_c179 bl[179] br[179] wl[81] vdd gnd cell_6t
Xbit_r82_c179 bl[179] br[179] wl[82] vdd gnd cell_6t
Xbit_r83_c179 bl[179] br[179] wl[83] vdd gnd cell_6t
Xbit_r84_c179 bl[179] br[179] wl[84] vdd gnd cell_6t
Xbit_r85_c179 bl[179] br[179] wl[85] vdd gnd cell_6t
Xbit_r86_c179 bl[179] br[179] wl[86] vdd gnd cell_6t
Xbit_r87_c179 bl[179] br[179] wl[87] vdd gnd cell_6t
Xbit_r88_c179 bl[179] br[179] wl[88] vdd gnd cell_6t
Xbit_r89_c179 bl[179] br[179] wl[89] vdd gnd cell_6t
Xbit_r90_c179 bl[179] br[179] wl[90] vdd gnd cell_6t
Xbit_r91_c179 bl[179] br[179] wl[91] vdd gnd cell_6t
Xbit_r92_c179 bl[179] br[179] wl[92] vdd gnd cell_6t
Xbit_r93_c179 bl[179] br[179] wl[93] vdd gnd cell_6t
Xbit_r94_c179 bl[179] br[179] wl[94] vdd gnd cell_6t
Xbit_r95_c179 bl[179] br[179] wl[95] vdd gnd cell_6t
Xbit_r96_c179 bl[179] br[179] wl[96] vdd gnd cell_6t
Xbit_r97_c179 bl[179] br[179] wl[97] vdd gnd cell_6t
Xbit_r98_c179 bl[179] br[179] wl[98] vdd gnd cell_6t
Xbit_r99_c179 bl[179] br[179] wl[99] vdd gnd cell_6t
Xbit_r100_c179 bl[179] br[179] wl[100] vdd gnd cell_6t
Xbit_r101_c179 bl[179] br[179] wl[101] vdd gnd cell_6t
Xbit_r102_c179 bl[179] br[179] wl[102] vdd gnd cell_6t
Xbit_r103_c179 bl[179] br[179] wl[103] vdd gnd cell_6t
Xbit_r104_c179 bl[179] br[179] wl[104] vdd gnd cell_6t
Xbit_r105_c179 bl[179] br[179] wl[105] vdd gnd cell_6t
Xbit_r106_c179 bl[179] br[179] wl[106] vdd gnd cell_6t
Xbit_r107_c179 bl[179] br[179] wl[107] vdd gnd cell_6t
Xbit_r108_c179 bl[179] br[179] wl[108] vdd gnd cell_6t
Xbit_r109_c179 bl[179] br[179] wl[109] vdd gnd cell_6t
Xbit_r110_c179 bl[179] br[179] wl[110] vdd gnd cell_6t
Xbit_r111_c179 bl[179] br[179] wl[111] vdd gnd cell_6t
Xbit_r112_c179 bl[179] br[179] wl[112] vdd gnd cell_6t
Xbit_r113_c179 bl[179] br[179] wl[113] vdd gnd cell_6t
Xbit_r114_c179 bl[179] br[179] wl[114] vdd gnd cell_6t
Xbit_r115_c179 bl[179] br[179] wl[115] vdd gnd cell_6t
Xbit_r116_c179 bl[179] br[179] wl[116] vdd gnd cell_6t
Xbit_r117_c179 bl[179] br[179] wl[117] vdd gnd cell_6t
Xbit_r118_c179 bl[179] br[179] wl[118] vdd gnd cell_6t
Xbit_r119_c179 bl[179] br[179] wl[119] vdd gnd cell_6t
Xbit_r120_c179 bl[179] br[179] wl[120] vdd gnd cell_6t
Xbit_r121_c179 bl[179] br[179] wl[121] vdd gnd cell_6t
Xbit_r122_c179 bl[179] br[179] wl[122] vdd gnd cell_6t
Xbit_r123_c179 bl[179] br[179] wl[123] vdd gnd cell_6t
Xbit_r124_c179 bl[179] br[179] wl[124] vdd gnd cell_6t
Xbit_r125_c179 bl[179] br[179] wl[125] vdd gnd cell_6t
Xbit_r126_c179 bl[179] br[179] wl[126] vdd gnd cell_6t
Xbit_r127_c179 bl[179] br[179] wl[127] vdd gnd cell_6t
Xbit_r128_c179 bl[179] br[179] wl[128] vdd gnd cell_6t
Xbit_r129_c179 bl[179] br[179] wl[129] vdd gnd cell_6t
Xbit_r130_c179 bl[179] br[179] wl[130] vdd gnd cell_6t
Xbit_r131_c179 bl[179] br[179] wl[131] vdd gnd cell_6t
Xbit_r132_c179 bl[179] br[179] wl[132] vdd gnd cell_6t
Xbit_r133_c179 bl[179] br[179] wl[133] vdd gnd cell_6t
Xbit_r134_c179 bl[179] br[179] wl[134] vdd gnd cell_6t
Xbit_r135_c179 bl[179] br[179] wl[135] vdd gnd cell_6t
Xbit_r136_c179 bl[179] br[179] wl[136] vdd gnd cell_6t
Xbit_r137_c179 bl[179] br[179] wl[137] vdd gnd cell_6t
Xbit_r138_c179 bl[179] br[179] wl[138] vdd gnd cell_6t
Xbit_r139_c179 bl[179] br[179] wl[139] vdd gnd cell_6t
Xbit_r140_c179 bl[179] br[179] wl[140] vdd gnd cell_6t
Xbit_r141_c179 bl[179] br[179] wl[141] vdd gnd cell_6t
Xbit_r142_c179 bl[179] br[179] wl[142] vdd gnd cell_6t
Xbit_r143_c179 bl[179] br[179] wl[143] vdd gnd cell_6t
Xbit_r144_c179 bl[179] br[179] wl[144] vdd gnd cell_6t
Xbit_r145_c179 bl[179] br[179] wl[145] vdd gnd cell_6t
Xbit_r146_c179 bl[179] br[179] wl[146] vdd gnd cell_6t
Xbit_r147_c179 bl[179] br[179] wl[147] vdd gnd cell_6t
Xbit_r148_c179 bl[179] br[179] wl[148] vdd gnd cell_6t
Xbit_r149_c179 bl[179] br[179] wl[149] vdd gnd cell_6t
Xbit_r150_c179 bl[179] br[179] wl[150] vdd gnd cell_6t
Xbit_r151_c179 bl[179] br[179] wl[151] vdd gnd cell_6t
Xbit_r152_c179 bl[179] br[179] wl[152] vdd gnd cell_6t
Xbit_r153_c179 bl[179] br[179] wl[153] vdd gnd cell_6t
Xbit_r154_c179 bl[179] br[179] wl[154] vdd gnd cell_6t
Xbit_r155_c179 bl[179] br[179] wl[155] vdd gnd cell_6t
Xbit_r156_c179 bl[179] br[179] wl[156] vdd gnd cell_6t
Xbit_r157_c179 bl[179] br[179] wl[157] vdd gnd cell_6t
Xbit_r158_c179 bl[179] br[179] wl[158] vdd gnd cell_6t
Xbit_r159_c179 bl[179] br[179] wl[159] vdd gnd cell_6t
Xbit_r160_c179 bl[179] br[179] wl[160] vdd gnd cell_6t
Xbit_r161_c179 bl[179] br[179] wl[161] vdd gnd cell_6t
Xbit_r162_c179 bl[179] br[179] wl[162] vdd gnd cell_6t
Xbit_r163_c179 bl[179] br[179] wl[163] vdd gnd cell_6t
Xbit_r164_c179 bl[179] br[179] wl[164] vdd gnd cell_6t
Xbit_r165_c179 bl[179] br[179] wl[165] vdd gnd cell_6t
Xbit_r166_c179 bl[179] br[179] wl[166] vdd gnd cell_6t
Xbit_r167_c179 bl[179] br[179] wl[167] vdd gnd cell_6t
Xbit_r168_c179 bl[179] br[179] wl[168] vdd gnd cell_6t
Xbit_r169_c179 bl[179] br[179] wl[169] vdd gnd cell_6t
Xbit_r170_c179 bl[179] br[179] wl[170] vdd gnd cell_6t
Xbit_r171_c179 bl[179] br[179] wl[171] vdd gnd cell_6t
Xbit_r172_c179 bl[179] br[179] wl[172] vdd gnd cell_6t
Xbit_r173_c179 bl[179] br[179] wl[173] vdd gnd cell_6t
Xbit_r174_c179 bl[179] br[179] wl[174] vdd gnd cell_6t
Xbit_r175_c179 bl[179] br[179] wl[175] vdd gnd cell_6t
Xbit_r176_c179 bl[179] br[179] wl[176] vdd gnd cell_6t
Xbit_r177_c179 bl[179] br[179] wl[177] vdd gnd cell_6t
Xbit_r178_c179 bl[179] br[179] wl[178] vdd gnd cell_6t
Xbit_r179_c179 bl[179] br[179] wl[179] vdd gnd cell_6t
Xbit_r180_c179 bl[179] br[179] wl[180] vdd gnd cell_6t
Xbit_r181_c179 bl[179] br[179] wl[181] vdd gnd cell_6t
Xbit_r182_c179 bl[179] br[179] wl[182] vdd gnd cell_6t
Xbit_r183_c179 bl[179] br[179] wl[183] vdd gnd cell_6t
Xbit_r184_c179 bl[179] br[179] wl[184] vdd gnd cell_6t
Xbit_r185_c179 bl[179] br[179] wl[185] vdd gnd cell_6t
Xbit_r186_c179 bl[179] br[179] wl[186] vdd gnd cell_6t
Xbit_r187_c179 bl[179] br[179] wl[187] vdd gnd cell_6t
Xbit_r188_c179 bl[179] br[179] wl[188] vdd gnd cell_6t
Xbit_r189_c179 bl[179] br[179] wl[189] vdd gnd cell_6t
Xbit_r190_c179 bl[179] br[179] wl[190] vdd gnd cell_6t
Xbit_r191_c179 bl[179] br[179] wl[191] vdd gnd cell_6t
Xbit_r192_c179 bl[179] br[179] wl[192] vdd gnd cell_6t
Xbit_r193_c179 bl[179] br[179] wl[193] vdd gnd cell_6t
Xbit_r194_c179 bl[179] br[179] wl[194] vdd gnd cell_6t
Xbit_r195_c179 bl[179] br[179] wl[195] vdd gnd cell_6t
Xbit_r196_c179 bl[179] br[179] wl[196] vdd gnd cell_6t
Xbit_r197_c179 bl[179] br[179] wl[197] vdd gnd cell_6t
Xbit_r198_c179 bl[179] br[179] wl[198] vdd gnd cell_6t
Xbit_r199_c179 bl[179] br[179] wl[199] vdd gnd cell_6t
Xbit_r200_c179 bl[179] br[179] wl[200] vdd gnd cell_6t
Xbit_r201_c179 bl[179] br[179] wl[201] vdd gnd cell_6t
Xbit_r202_c179 bl[179] br[179] wl[202] vdd gnd cell_6t
Xbit_r203_c179 bl[179] br[179] wl[203] vdd gnd cell_6t
Xbit_r204_c179 bl[179] br[179] wl[204] vdd gnd cell_6t
Xbit_r205_c179 bl[179] br[179] wl[205] vdd gnd cell_6t
Xbit_r206_c179 bl[179] br[179] wl[206] vdd gnd cell_6t
Xbit_r207_c179 bl[179] br[179] wl[207] vdd gnd cell_6t
Xbit_r208_c179 bl[179] br[179] wl[208] vdd gnd cell_6t
Xbit_r209_c179 bl[179] br[179] wl[209] vdd gnd cell_6t
Xbit_r210_c179 bl[179] br[179] wl[210] vdd gnd cell_6t
Xbit_r211_c179 bl[179] br[179] wl[211] vdd gnd cell_6t
Xbit_r212_c179 bl[179] br[179] wl[212] vdd gnd cell_6t
Xbit_r213_c179 bl[179] br[179] wl[213] vdd gnd cell_6t
Xbit_r214_c179 bl[179] br[179] wl[214] vdd gnd cell_6t
Xbit_r215_c179 bl[179] br[179] wl[215] vdd gnd cell_6t
Xbit_r216_c179 bl[179] br[179] wl[216] vdd gnd cell_6t
Xbit_r217_c179 bl[179] br[179] wl[217] vdd gnd cell_6t
Xbit_r218_c179 bl[179] br[179] wl[218] vdd gnd cell_6t
Xbit_r219_c179 bl[179] br[179] wl[219] vdd gnd cell_6t
Xbit_r220_c179 bl[179] br[179] wl[220] vdd gnd cell_6t
Xbit_r221_c179 bl[179] br[179] wl[221] vdd gnd cell_6t
Xbit_r222_c179 bl[179] br[179] wl[222] vdd gnd cell_6t
Xbit_r223_c179 bl[179] br[179] wl[223] vdd gnd cell_6t
Xbit_r224_c179 bl[179] br[179] wl[224] vdd gnd cell_6t
Xbit_r225_c179 bl[179] br[179] wl[225] vdd gnd cell_6t
Xbit_r226_c179 bl[179] br[179] wl[226] vdd gnd cell_6t
Xbit_r227_c179 bl[179] br[179] wl[227] vdd gnd cell_6t
Xbit_r228_c179 bl[179] br[179] wl[228] vdd gnd cell_6t
Xbit_r229_c179 bl[179] br[179] wl[229] vdd gnd cell_6t
Xbit_r230_c179 bl[179] br[179] wl[230] vdd gnd cell_6t
Xbit_r231_c179 bl[179] br[179] wl[231] vdd gnd cell_6t
Xbit_r232_c179 bl[179] br[179] wl[232] vdd gnd cell_6t
Xbit_r233_c179 bl[179] br[179] wl[233] vdd gnd cell_6t
Xbit_r234_c179 bl[179] br[179] wl[234] vdd gnd cell_6t
Xbit_r235_c179 bl[179] br[179] wl[235] vdd gnd cell_6t
Xbit_r236_c179 bl[179] br[179] wl[236] vdd gnd cell_6t
Xbit_r237_c179 bl[179] br[179] wl[237] vdd gnd cell_6t
Xbit_r238_c179 bl[179] br[179] wl[238] vdd gnd cell_6t
Xbit_r239_c179 bl[179] br[179] wl[239] vdd gnd cell_6t
Xbit_r240_c179 bl[179] br[179] wl[240] vdd gnd cell_6t
Xbit_r241_c179 bl[179] br[179] wl[241] vdd gnd cell_6t
Xbit_r242_c179 bl[179] br[179] wl[242] vdd gnd cell_6t
Xbit_r243_c179 bl[179] br[179] wl[243] vdd gnd cell_6t
Xbit_r244_c179 bl[179] br[179] wl[244] vdd gnd cell_6t
Xbit_r245_c179 bl[179] br[179] wl[245] vdd gnd cell_6t
Xbit_r246_c179 bl[179] br[179] wl[246] vdd gnd cell_6t
Xbit_r247_c179 bl[179] br[179] wl[247] vdd gnd cell_6t
Xbit_r248_c179 bl[179] br[179] wl[248] vdd gnd cell_6t
Xbit_r249_c179 bl[179] br[179] wl[249] vdd gnd cell_6t
Xbit_r250_c179 bl[179] br[179] wl[250] vdd gnd cell_6t
Xbit_r251_c179 bl[179] br[179] wl[251] vdd gnd cell_6t
Xbit_r252_c179 bl[179] br[179] wl[252] vdd gnd cell_6t
Xbit_r253_c179 bl[179] br[179] wl[253] vdd gnd cell_6t
Xbit_r254_c179 bl[179] br[179] wl[254] vdd gnd cell_6t
Xbit_r255_c179 bl[179] br[179] wl[255] vdd gnd cell_6t
Xbit_r0_c180 bl[180] br[180] wl[0] vdd gnd cell_6t
Xbit_r1_c180 bl[180] br[180] wl[1] vdd gnd cell_6t
Xbit_r2_c180 bl[180] br[180] wl[2] vdd gnd cell_6t
Xbit_r3_c180 bl[180] br[180] wl[3] vdd gnd cell_6t
Xbit_r4_c180 bl[180] br[180] wl[4] vdd gnd cell_6t
Xbit_r5_c180 bl[180] br[180] wl[5] vdd gnd cell_6t
Xbit_r6_c180 bl[180] br[180] wl[6] vdd gnd cell_6t
Xbit_r7_c180 bl[180] br[180] wl[7] vdd gnd cell_6t
Xbit_r8_c180 bl[180] br[180] wl[8] vdd gnd cell_6t
Xbit_r9_c180 bl[180] br[180] wl[9] vdd gnd cell_6t
Xbit_r10_c180 bl[180] br[180] wl[10] vdd gnd cell_6t
Xbit_r11_c180 bl[180] br[180] wl[11] vdd gnd cell_6t
Xbit_r12_c180 bl[180] br[180] wl[12] vdd gnd cell_6t
Xbit_r13_c180 bl[180] br[180] wl[13] vdd gnd cell_6t
Xbit_r14_c180 bl[180] br[180] wl[14] vdd gnd cell_6t
Xbit_r15_c180 bl[180] br[180] wl[15] vdd gnd cell_6t
Xbit_r16_c180 bl[180] br[180] wl[16] vdd gnd cell_6t
Xbit_r17_c180 bl[180] br[180] wl[17] vdd gnd cell_6t
Xbit_r18_c180 bl[180] br[180] wl[18] vdd gnd cell_6t
Xbit_r19_c180 bl[180] br[180] wl[19] vdd gnd cell_6t
Xbit_r20_c180 bl[180] br[180] wl[20] vdd gnd cell_6t
Xbit_r21_c180 bl[180] br[180] wl[21] vdd gnd cell_6t
Xbit_r22_c180 bl[180] br[180] wl[22] vdd gnd cell_6t
Xbit_r23_c180 bl[180] br[180] wl[23] vdd gnd cell_6t
Xbit_r24_c180 bl[180] br[180] wl[24] vdd gnd cell_6t
Xbit_r25_c180 bl[180] br[180] wl[25] vdd gnd cell_6t
Xbit_r26_c180 bl[180] br[180] wl[26] vdd gnd cell_6t
Xbit_r27_c180 bl[180] br[180] wl[27] vdd gnd cell_6t
Xbit_r28_c180 bl[180] br[180] wl[28] vdd gnd cell_6t
Xbit_r29_c180 bl[180] br[180] wl[29] vdd gnd cell_6t
Xbit_r30_c180 bl[180] br[180] wl[30] vdd gnd cell_6t
Xbit_r31_c180 bl[180] br[180] wl[31] vdd gnd cell_6t
Xbit_r32_c180 bl[180] br[180] wl[32] vdd gnd cell_6t
Xbit_r33_c180 bl[180] br[180] wl[33] vdd gnd cell_6t
Xbit_r34_c180 bl[180] br[180] wl[34] vdd gnd cell_6t
Xbit_r35_c180 bl[180] br[180] wl[35] vdd gnd cell_6t
Xbit_r36_c180 bl[180] br[180] wl[36] vdd gnd cell_6t
Xbit_r37_c180 bl[180] br[180] wl[37] vdd gnd cell_6t
Xbit_r38_c180 bl[180] br[180] wl[38] vdd gnd cell_6t
Xbit_r39_c180 bl[180] br[180] wl[39] vdd gnd cell_6t
Xbit_r40_c180 bl[180] br[180] wl[40] vdd gnd cell_6t
Xbit_r41_c180 bl[180] br[180] wl[41] vdd gnd cell_6t
Xbit_r42_c180 bl[180] br[180] wl[42] vdd gnd cell_6t
Xbit_r43_c180 bl[180] br[180] wl[43] vdd gnd cell_6t
Xbit_r44_c180 bl[180] br[180] wl[44] vdd gnd cell_6t
Xbit_r45_c180 bl[180] br[180] wl[45] vdd gnd cell_6t
Xbit_r46_c180 bl[180] br[180] wl[46] vdd gnd cell_6t
Xbit_r47_c180 bl[180] br[180] wl[47] vdd gnd cell_6t
Xbit_r48_c180 bl[180] br[180] wl[48] vdd gnd cell_6t
Xbit_r49_c180 bl[180] br[180] wl[49] vdd gnd cell_6t
Xbit_r50_c180 bl[180] br[180] wl[50] vdd gnd cell_6t
Xbit_r51_c180 bl[180] br[180] wl[51] vdd gnd cell_6t
Xbit_r52_c180 bl[180] br[180] wl[52] vdd gnd cell_6t
Xbit_r53_c180 bl[180] br[180] wl[53] vdd gnd cell_6t
Xbit_r54_c180 bl[180] br[180] wl[54] vdd gnd cell_6t
Xbit_r55_c180 bl[180] br[180] wl[55] vdd gnd cell_6t
Xbit_r56_c180 bl[180] br[180] wl[56] vdd gnd cell_6t
Xbit_r57_c180 bl[180] br[180] wl[57] vdd gnd cell_6t
Xbit_r58_c180 bl[180] br[180] wl[58] vdd gnd cell_6t
Xbit_r59_c180 bl[180] br[180] wl[59] vdd gnd cell_6t
Xbit_r60_c180 bl[180] br[180] wl[60] vdd gnd cell_6t
Xbit_r61_c180 bl[180] br[180] wl[61] vdd gnd cell_6t
Xbit_r62_c180 bl[180] br[180] wl[62] vdd gnd cell_6t
Xbit_r63_c180 bl[180] br[180] wl[63] vdd gnd cell_6t
Xbit_r64_c180 bl[180] br[180] wl[64] vdd gnd cell_6t
Xbit_r65_c180 bl[180] br[180] wl[65] vdd gnd cell_6t
Xbit_r66_c180 bl[180] br[180] wl[66] vdd gnd cell_6t
Xbit_r67_c180 bl[180] br[180] wl[67] vdd gnd cell_6t
Xbit_r68_c180 bl[180] br[180] wl[68] vdd gnd cell_6t
Xbit_r69_c180 bl[180] br[180] wl[69] vdd gnd cell_6t
Xbit_r70_c180 bl[180] br[180] wl[70] vdd gnd cell_6t
Xbit_r71_c180 bl[180] br[180] wl[71] vdd gnd cell_6t
Xbit_r72_c180 bl[180] br[180] wl[72] vdd gnd cell_6t
Xbit_r73_c180 bl[180] br[180] wl[73] vdd gnd cell_6t
Xbit_r74_c180 bl[180] br[180] wl[74] vdd gnd cell_6t
Xbit_r75_c180 bl[180] br[180] wl[75] vdd gnd cell_6t
Xbit_r76_c180 bl[180] br[180] wl[76] vdd gnd cell_6t
Xbit_r77_c180 bl[180] br[180] wl[77] vdd gnd cell_6t
Xbit_r78_c180 bl[180] br[180] wl[78] vdd gnd cell_6t
Xbit_r79_c180 bl[180] br[180] wl[79] vdd gnd cell_6t
Xbit_r80_c180 bl[180] br[180] wl[80] vdd gnd cell_6t
Xbit_r81_c180 bl[180] br[180] wl[81] vdd gnd cell_6t
Xbit_r82_c180 bl[180] br[180] wl[82] vdd gnd cell_6t
Xbit_r83_c180 bl[180] br[180] wl[83] vdd gnd cell_6t
Xbit_r84_c180 bl[180] br[180] wl[84] vdd gnd cell_6t
Xbit_r85_c180 bl[180] br[180] wl[85] vdd gnd cell_6t
Xbit_r86_c180 bl[180] br[180] wl[86] vdd gnd cell_6t
Xbit_r87_c180 bl[180] br[180] wl[87] vdd gnd cell_6t
Xbit_r88_c180 bl[180] br[180] wl[88] vdd gnd cell_6t
Xbit_r89_c180 bl[180] br[180] wl[89] vdd gnd cell_6t
Xbit_r90_c180 bl[180] br[180] wl[90] vdd gnd cell_6t
Xbit_r91_c180 bl[180] br[180] wl[91] vdd gnd cell_6t
Xbit_r92_c180 bl[180] br[180] wl[92] vdd gnd cell_6t
Xbit_r93_c180 bl[180] br[180] wl[93] vdd gnd cell_6t
Xbit_r94_c180 bl[180] br[180] wl[94] vdd gnd cell_6t
Xbit_r95_c180 bl[180] br[180] wl[95] vdd gnd cell_6t
Xbit_r96_c180 bl[180] br[180] wl[96] vdd gnd cell_6t
Xbit_r97_c180 bl[180] br[180] wl[97] vdd gnd cell_6t
Xbit_r98_c180 bl[180] br[180] wl[98] vdd gnd cell_6t
Xbit_r99_c180 bl[180] br[180] wl[99] vdd gnd cell_6t
Xbit_r100_c180 bl[180] br[180] wl[100] vdd gnd cell_6t
Xbit_r101_c180 bl[180] br[180] wl[101] vdd gnd cell_6t
Xbit_r102_c180 bl[180] br[180] wl[102] vdd gnd cell_6t
Xbit_r103_c180 bl[180] br[180] wl[103] vdd gnd cell_6t
Xbit_r104_c180 bl[180] br[180] wl[104] vdd gnd cell_6t
Xbit_r105_c180 bl[180] br[180] wl[105] vdd gnd cell_6t
Xbit_r106_c180 bl[180] br[180] wl[106] vdd gnd cell_6t
Xbit_r107_c180 bl[180] br[180] wl[107] vdd gnd cell_6t
Xbit_r108_c180 bl[180] br[180] wl[108] vdd gnd cell_6t
Xbit_r109_c180 bl[180] br[180] wl[109] vdd gnd cell_6t
Xbit_r110_c180 bl[180] br[180] wl[110] vdd gnd cell_6t
Xbit_r111_c180 bl[180] br[180] wl[111] vdd gnd cell_6t
Xbit_r112_c180 bl[180] br[180] wl[112] vdd gnd cell_6t
Xbit_r113_c180 bl[180] br[180] wl[113] vdd gnd cell_6t
Xbit_r114_c180 bl[180] br[180] wl[114] vdd gnd cell_6t
Xbit_r115_c180 bl[180] br[180] wl[115] vdd gnd cell_6t
Xbit_r116_c180 bl[180] br[180] wl[116] vdd gnd cell_6t
Xbit_r117_c180 bl[180] br[180] wl[117] vdd gnd cell_6t
Xbit_r118_c180 bl[180] br[180] wl[118] vdd gnd cell_6t
Xbit_r119_c180 bl[180] br[180] wl[119] vdd gnd cell_6t
Xbit_r120_c180 bl[180] br[180] wl[120] vdd gnd cell_6t
Xbit_r121_c180 bl[180] br[180] wl[121] vdd gnd cell_6t
Xbit_r122_c180 bl[180] br[180] wl[122] vdd gnd cell_6t
Xbit_r123_c180 bl[180] br[180] wl[123] vdd gnd cell_6t
Xbit_r124_c180 bl[180] br[180] wl[124] vdd gnd cell_6t
Xbit_r125_c180 bl[180] br[180] wl[125] vdd gnd cell_6t
Xbit_r126_c180 bl[180] br[180] wl[126] vdd gnd cell_6t
Xbit_r127_c180 bl[180] br[180] wl[127] vdd gnd cell_6t
Xbit_r128_c180 bl[180] br[180] wl[128] vdd gnd cell_6t
Xbit_r129_c180 bl[180] br[180] wl[129] vdd gnd cell_6t
Xbit_r130_c180 bl[180] br[180] wl[130] vdd gnd cell_6t
Xbit_r131_c180 bl[180] br[180] wl[131] vdd gnd cell_6t
Xbit_r132_c180 bl[180] br[180] wl[132] vdd gnd cell_6t
Xbit_r133_c180 bl[180] br[180] wl[133] vdd gnd cell_6t
Xbit_r134_c180 bl[180] br[180] wl[134] vdd gnd cell_6t
Xbit_r135_c180 bl[180] br[180] wl[135] vdd gnd cell_6t
Xbit_r136_c180 bl[180] br[180] wl[136] vdd gnd cell_6t
Xbit_r137_c180 bl[180] br[180] wl[137] vdd gnd cell_6t
Xbit_r138_c180 bl[180] br[180] wl[138] vdd gnd cell_6t
Xbit_r139_c180 bl[180] br[180] wl[139] vdd gnd cell_6t
Xbit_r140_c180 bl[180] br[180] wl[140] vdd gnd cell_6t
Xbit_r141_c180 bl[180] br[180] wl[141] vdd gnd cell_6t
Xbit_r142_c180 bl[180] br[180] wl[142] vdd gnd cell_6t
Xbit_r143_c180 bl[180] br[180] wl[143] vdd gnd cell_6t
Xbit_r144_c180 bl[180] br[180] wl[144] vdd gnd cell_6t
Xbit_r145_c180 bl[180] br[180] wl[145] vdd gnd cell_6t
Xbit_r146_c180 bl[180] br[180] wl[146] vdd gnd cell_6t
Xbit_r147_c180 bl[180] br[180] wl[147] vdd gnd cell_6t
Xbit_r148_c180 bl[180] br[180] wl[148] vdd gnd cell_6t
Xbit_r149_c180 bl[180] br[180] wl[149] vdd gnd cell_6t
Xbit_r150_c180 bl[180] br[180] wl[150] vdd gnd cell_6t
Xbit_r151_c180 bl[180] br[180] wl[151] vdd gnd cell_6t
Xbit_r152_c180 bl[180] br[180] wl[152] vdd gnd cell_6t
Xbit_r153_c180 bl[180] br[180] wl[153] vdd gnd cell_6t
Xbit_r154_c180 bl[180] br[180] wl[154] vdd gnd cell_6t
Xbit_r155_c180 bl[180] br[180] wl[155] vdd gnd cell_6t
Xbit_r156_c180 bl[180] br[180] wl[156] vdd gnd cell_6t
Xbit_r157_c180 bl[180] br[180] wl[157] vdd gnd cell_6t
Xbit_r158_c180 bl[180] br[180] wl[158] vdd gnd cell_6t
Xbit_r159_c180 bl[180] br[180] wl[159] vdd gnd cell_6t
Xbit_r160_c180 bl[180] br[180] wl[160] vdd gnd cell_6t
Xbit_r161_c180 bl[180] br[180] wl[161] vdd gnd cell_6t
Xbit_r162_c180 bl[180] br[180] wl[162] vdd gnd cell_6t
Xbit_r163_c180 bl[180] br[180] wl[163] vdd gnd cell_6t
Xbit_r164_c180 bl[180] br[180] wl[164] vdd gnd cell_6t
Xbit_r165_c180 bl[180] br[180] wl[165] vdd gnd cell_6t
Xbit_r166_c180 bl[180] br[180] wl[166] vdd gnd cell_6t
Xbit_r167_c180 bl[180] br[180] wl[167] vdd gnd cell_6t
Xbit_r168_c180 bl[180] br[180] wl[168] vdd gnd cell_6t
Xbit_r169_c180 bl[180] br[180] wl[169] vdd gnd cell_6t
Xbit_r170_c180 bl[180] br[180] wl[170] vdd gnd cell_6t
Xbit_r171_c180 bl[180] br[180] wl[171] vdd gnd cell_6t
Xbit_r172_c180 bl[180] br[180] wl[172] vdd gnd cell_6t
Xbit_r173_c180 bl[180] br[180] wl[173] vdd gnd cell_6t
Xbit_r174_c180 bl[180] br[180] wl[174] vdd gnd cell_6t
Xbit_r175_c180 bl[180] br[180] wl[175] vdd gnd cell_6t
Xbit_r176_c180 bl[180] br[180] wl[176] vdd gnd cell_6t
Xbit_r177_c180 bl[180] br[180] wl[177] vdd gnd cell_6t
Xbit_r178_c180 bl[180] br[180] wl[178] vdd gnd cell_6t
Xbit_r179_c180 bl[180] br[180] wl[179] vdd gnd cell_6t
Xbit_r180_c180 bl[180] br[180] wl[180] vdd gnd cell_6t
Xbit_r181_c180 bl[180] br[180] wl[181] vdd gnd cell_6t
Xbit_r182_c180 bl[180] br[180] wl[182] vdd gnd cell_6t
Xbit_r183_c180 bl[180] br[180] wl[183] vdd gnd cell_6t
Xbit_r184_c180 bl[180] br[180] wl[184] vdd gnd cell_6t
Xbit_r185_c180 bl[180] br[180] wl[185] vdd gnd cell_6t
Xbit_r186_c180 bl[180] br[180] wl[186] vdd gnd cell_6t
Xbit_r187_c180 bl[180] br[180] wl[187] vdd gnd cell_6t
Xbit_r188_c180 bl[180] br[180] wl[188] vdd gnd cell_6t
Xbit_r189_c180 bl[180] br[180] wl[189] vdd gnd cell_6t
Xbit_r190_c180 bl[180] br[180] wl[190] vdd gnd cell_6t
Xbit_r191_c180 bl[180] br[180] wl[191] vdd gnd cell_6t
Xbit_r192_c180 bl[180] br[180] wl[192] vdd gnd cell_6t
Xbit_r193_c180 bl[180] br[180] wl[193] vdd gnd cell_6t
Xbit_r194_c180 bl[180] br[180] wl[194] vdd gnd cell_6t
Xbit_r195_c180 bl[180] br[180] wl[195] vdd gnd cell_6t
Xbit_r196_c180 bl[180] br[180] wl[196] vdd gnd cell_6t
Xbit_r197_c180 bl[180] br[180] wl[197] vdd gnd cell_6t
Xbit_r198_c180 bl[180] br[180] wl[198] vdd gnd cell_6t
Xbit_r199_c180 bl[180] br[180] wl[199] vdd gnd cell_6t
Xbit_r200_c180 bl[180] br[180] wl[200] vdd gnd cell_6t
Xbit_r201_c180 bl[180] br[180] wl[201] vdd gnd cell_6t
Xbit_r202_c180 bl[180] br[180] wl[202] vdd gnd cell_6t
Xbit_r203_c180 bl[180] br[180] wl[203] vdd gnd cell_6t
Xbit_r204_c180 bl[180] br[180] wl[204] vdd gnd cell_6t
Xbit_r205_c180 bl[180] br[180] wl[205] vdd gnd cell_6t
Xbit_r206_c180 bl[180] br[180] wl[206] vdd gnd cell_6t
Xbit_r207_c180 bl[180] br[180] wl[207] vdd gnd cell_6t
Xbit_r208_c180 bl[180] br[180] wl[208] vdd gnd cell_6t
Xbit_r209_c180 bl[180] br[180] wl[209] vdd gnd cell_6t
Xbit_r210_c180 bl[180] br[180] wl[210] vdd gnd cell_6t
Xbit_r211_c180 bl[180] br[180] wl[211] vdd gnd cell_6t
Xbit_r212_c180 bl[180] br[180] wl[212] vdd gnd cell_6t
Xbit_r213_c180 bl[180] br[180] wl[213] vdd gnd cell_6t
Xbit_r214_c180 bl[180] br[180] wl[214] vdd gnd cell_6t
Xbit_r215_c180 bl[180] br[180] wl[215] vdd gnd cell_6t
Xbit_r216_c180 bl[180] br[180] wl[216] vdd gnd cell_6t
Xbit_r217_c180 bl[180] br[180] wl[217] vdd gnd cell_6t
Xbit_r218_c180 bl[180] br[180] wl[218] vdd gnd cell_6t
Xbit_r219_c180 bl[180] br[180] wl[219] vdd gnd cell_6t
Xbit_r220_c180 bl[180] br[180] wl[220] vdd gnd cell_6t
Xbit_r221_c180 bl[180] br[180] wl[221] vdd gnd cell_6t
Xbit_r222_c180 bl[180] br[180] wl[222] vdd gnd cell_6t
Xbit_r223_c180 bl[180] br[180] wl[223] vdd gnd cell_6t
Xbit_r224_c180 bl[180] br[180] wl[224] vdd gnd cell_6t
Xbit_r225_c180 bl[180] br[180] wl[225] vdd gnd cell_6t
Xbit_r226_c180 bl[180] br[180] wl[226] vdd gnd cell_6t
Xbit_r227_c180 bl[180] br[180] wl[227] vdd gnd cell_6t
Xbit_r228_c180 bl[180] br[180] wl[228] vdd gnd cell_6t
Xbit_r229_c180 bl[180] br[180] wl[229] vdd gnd cell_6t
Xbit_r230_c180 bl[180] br[180] wl[230] vdd gnd cell_6t
Xbit_r231_c180 bl[180] br[180] wl[231] vdd gnd cell_6t
Xbit_r232_c180 bl[180] br[180] wl[232] vdd gnd cell_6t
Xbit_r233_c180 bl[180] br[180] wl[233] vdd gnd cell_6t
Xbit_r234_c180 bl[180] br[180] wl[234] vdd gnd cell_6t
Xbit_r235_c180 bl[180] br[180] wl[235] vdd gnd cell_6t
Xbit_r236_c180 bl[180] br[180] wl[236] vdd gnd cell_6t
Xbit_r237_c180 bl[180] br[180] wl[237] vdd gnd cell_6t
Xbit_r238_c180 bl[180] br[180] wl[238] vdd gnd cell_6t
Xbit_r239_c180 bl[180] br[180] wl[239] vdd gnd cell_6t
Xbit_r240_c180 bl[180] br[180] wl[240] vdd gnd cell_6t
Xbit_r241_c180 bl[180] br[180] wl[241] vdd gnd cell_6t
Xbit_r242_c180 bl[180] br[180] wl[242] vdd gnd cell_6t
Xbit_r243_c180 bl[180] br[180] wl[243] vdd gnd cell_6t
Xbit_r244_c180 bl[180] br[180] wl[244] vdd gnd cell_6t
Xbit_r245_c180 bl[180] br[180] wl[245] vdd gnd cell_6t
Xbit_r246_c180 bl[180] br[180] wl[246] vdd gnd cell_6t
Xbit_r247_c180 bl[180] br[180] wl[247] vdd gnd cell_6t
Xbit_r248_c180 bl[180] br[180] wl[248] vdd gnd cell_6t
Xbit_r249_c180 bl[180] br[180] wl[249] vdd gnd cell_6t
Xbit_r250_c180 bl[180] br[180] wl[250] vdd gnd cell_6t
Xbit_r251_c180 bl[180] br[180] wl[251] vdd gnd cell_6t
Xbit_r252_c180 bl[180] br[180] wl[252] vdd gnd cell_6t
Xbit_r253_c180 bl[180] br[180] wl[253] vdd gnd cell_6t
Xbit_r254_c180 bl[180] br[180] wl[254] vdd gnd cell_6t
Xbit_r255_c180 bl[180] br[180] wl[255] vdd gnd cell_6t
Xbit_r0_c181 bl[181] br[181] wl[0] vdd gnd cell_6t
Xbit_r1_c181 bl[181] br[181] wl[1] vdd gnd cell_6t
Xbit_r2_c181 bl[181] br[181] wl[2] vdd gnd cell_6t
Xbit_r3_c181 bl[181] br[181] wl[3] vdd gnd cell_6t
Xbit_r4_c181 bl[181] br[181] wl[4] vdd gnd cell_6t
Xbit_r5_c181 bl[181] br[181] wl[5] vdd gnd cell_6t
Xbit_r6_c181 bl[181] br[181] wl[6] vdd gnd cell_6t
Xbit_r7_c181 bl[181] br[181] wl[7] vdd gnd cell_6t
Xbit_r8_c181 bl[181] br[181] wl[8] vdd gnd cell_6t
Xbit_r9_c181 bl[181] br[181] wl[9] vdd gnd cell_6t
Xbit_r10_c181 bl[181] br[181] wl[10] vdd gnd cell_6t
Xbit_r11_c181 bl[181] br[181] wl[11] vdd gnd cell_6t
Xbit_r12_c181 bl[181] br[181] wl[12] vdd gnd cell_6t
Xbit_r13_c181 bl[181] br[181] wl[13] vdd gnd cell_6t
Xbit_r14_c181 bl[181] br[181] wl[14] vdd gnd cell_6t
Xbit_r15_c181 bl[181] br[181] wl[15] vdd gnd cell_6t
Xbit_r16_c181 bl[181] br[181] wl[16] vdd gnd cell_6t
Xbit_r17_c181 bl[181] br[181] wl[17] vdd gnd cell_6t
Xbit_r18_c181 bl[181] br[181] wl[18] vdd gnd cell_6t
Xbit_r19_c181 bl[181] br[181] wl[19] vdd gnd cell_6t
Xbit_r20_c181 bl[181] br[181] wl[20] vdd gnd cell_6t
Xbit_r21_c181 bl[181] br[181] wl[21] vdd gnd cell_6t
Xbit_r22_c181 bl[181] br[181] wl[22] vdd gnd cell_6t
Xbit_r23_c181 bl[181] br[181] wl[23] vdd gnd cell_6t
Xbit_r24_c181 bl[181] br[181] wl[24] vdd gnd cell_6t
Xbit_r25_c181 bl[181] br[181] wl[25] vdd gnd cell_6t
Xbit_r26_c181 bl[181] br[181] wl[26] vdd gnd cell_6t
Xbit_r27_c181 bl[181] br[181] wl[27] vdd gnd cell_6t
Xbit_r28_c181 bl[181] br[181] wl[28] vdd gnd cell_6t
Xbit_r29_c181 bl[181] br[181] wl[29] vdd gnd cell_6t
Xbit_r30_c181 bl[181] br[181] wl[30] vdd gnd cell_6t
Xbit_r31_c181 bl[181] br[181] wl[31] vdd gnd cell_6t
Xbit_r32_c181 bl[181] br[181] wl[32] vdd gnd cell_6t
Xbit_r33_c181 bl[181] br[181] wl[33] vdd gnd cell_6t
Xbit_r34_c181 bl[181] br[181] wl[34] vdd gnd cell_6t
Xbit_r35_c181 bl[181] br[181] wl[35] vdd gnd cell_6t
Xbit_r36_c181 bl[181] br[181] wl[36] vdd gnd cell_6t
Xbit_r37_c181 bl[181] br[181] wl[37] vdd gnd cell_6t
Xbit_r38_c181 bl[181] br[181] wl[38] vdd gnd cell_6t
Xbit_r39_c181 bl[181] br[181] wl[39] vdd gnd cell_6t
Xbit_r40_c181 bl[181] br[181] wl[40] vdd gnd cell_6t
Xbit_r41_c181 bl[181] br[181] wl[41] vdd gnd cell_6t
Xbit_r42_c181 bl[181] br[181] wl[42] vdd gnd cell_6t
Xbit_r43_c181 bl[181] br[181] wl[43] vdd gnd cell_6t
Xbit_r44_c181 bl[181] br[181] wl[44] vdd gnd cell_6t
Xbit_r45_c181 bl[181] br[181] wl[45] vdd gnd cell_6t
Xbit_r46_c181 bl[181] br[181] wl[46] vdd gnd cell_6t
Xbit_r47_c181 bl[181] br[181] wl[47] vdd gnd cell_6t
Xbit_r48_c181 bl[181] br[181] wl[48] vdd gnd cell_6t
Xbit_r49_c181 bl[181] br[181] wl[49] vdd gnd cell_6t
Xbit_r50_c181 bl[181] br[181] wl[50] vdd gnd cell_6t
Xbit_r51_c181 bl[181] br[181] wl[51] vdd gnd cell_6t
Xbit_r52_c181 bl[181] br[181] wl[52] vdd gnd cell_6t
Xbit_r53_c181 bl[181] br[181] wl[53] vdd gnd cell_6t
Xbit_r54_c181 bl[181] br[181] wl[54] vdd gnd cell_6t
Xbit_r55_c181 bl[181] br[181] wl[55] vdd gnd cell_6t
Xbit_r56_c181 bl[181] br[181] wl[56] vdd gnd cell_6t
Xbit_r57_c181 bl[181] br[181] wl[57] vdd gnd cell_6t
Xbit_r58_c181 bl[181] br[181] wl[58] vdd gnd cell_6t
Xbit_r59_c181 bl[181] br[181] wl[59] vdd gnd cell_6t
Xbit_r60_c181 bl[181] br[181] wl[60] vdd gnd cell_6t
Xbit_r61_c181 bl[181] br[181] wl[61] vdd gnd cell_6t
Xbit_r62_c181 bl[181] br[181] wl[62] vdd gnd cell_6t
Xbit_r63_c181 bl[181] br[181] wl[63] vdd gnd cell_6t
Xbit_r64_c181 bl[181] br[181] wl[64] vdd gnd cell_6t
Xbit_r65_c181 bl[181] br[181] wl[65] vdd gnd cell_6t
Xbit_r66_c181 bl[181] br[181] wl[66] vdd gnd cell_6t
Xbit_r67_c181 bl[181] br[181] wl[67] vdd gnd cell_6t
Xbit_r68_c181 bl[181] br[181] wl[68] vdd gnd cell_6t
Xbit_r69_c181 bl[181] br[181] wl[69] vdd gnd cell_6t
Xbit_r70_c181 bl[181] br[181] wl[70] vdd gnd cell_6t
Xbit_r71_c181 bl[181] br[181] wl[71] vdd gnd cell_6t
Xbit_r72_c181 bl[181] br[181] wl[72] vdd gnd cell_6t
Xbit_r73_c181 bl[181] br[181] wl[73] vdd gnd cell_6t
Xbit_r74_c181 bl[181] br[181] wl[74] vdd gnd cell_6t
Xbit_r75_c181 bl[181] br[181] wl[75] vdd gnd cell_6t
Xbit_r76_c181 bl[181] br[181] wl[76] vdd gnd cell_6t
Xbit_r77_c181 bl[181] br[181] wl[77] vdd gnd cell_6t
Xbit_r78_c181 bl[181] br[181] wl[78] vdd gnd cell_6t
Xbit_r79_c181 bl[181] br[181] wl[79] vdd gnd cell_6t
Xbit_r80_c181 bl[181] br[181] wl[80] vdd gnd cell_6t
Xbit_r81_c181 bl[181] br[181] wl[81] vdd gnd cell_6t
Xbit_r82_c181 bl[181] br[181] wl[82] vdd gnd cell_6t
Xbit_r83_c181 bl[181] br[181] wl[83] vdd gnd cell_6t
Xbit_r84_c181 bl[181] br[181] wl[84] vdd gnd cell_6t
Xbit_r85_c181 bl[181] br[181] wl[85] vdd gnd cell_6t
Xbit_r86_c181 bl[181] br[181] wl[86] vdd gnd cell_6t
Xbit_r87_c181 bl[181] br[181] wl[87] vdd gnd cell_6t
Xbit_r88_c181 bl[181] br[181] wl[88] vdd gnd cell_6t
Xbit_r89_c181 bl[181] br[181] wl[89] vdd gnd cell_6t
Xbit_r90_c181 bl[181] br[181] wl[90] vdd gnd cell_6t
Xbit_r91_c181 bl[181] br[181] wl[91] vdd gnd cell_6t
Xbit_r92_c181 bl[181] br[181] wl[92] vdd gnd cell_6t
Xbit_r93_c181 bl[181] br[181] wl[93] vdd gnd cell_6t
Xbit_r94_c181 bl[181] br[181] wl[94] vdd gnd cell_6t
Xbit_r95_c181 bl[181] br[181] wl[95] vdd gnd cell_6t
Xbit_r96_c181 bl[181] br[181] wl[96] vdd gnd cell_6t
Xbit_r97_c181 bl[181] br[181] wl[97] vdd gnd cell_6t
Xbit_r98_c181 bl[181] br[181] wl[98] vdd gnd cell_6t
Xbit_r99_c181 bl[181] br[181] wl[99] vdd gnd cell_6t
Xbit_r100_c181 bl[181] br[181] wl[100] vdd gnd cell_6t
Xbit_r101_c181 bl[181] br[181] wl[101] vdd gnd cell_6t
Xbit_r102_c181 bl[181] br[181] wl[102] vdd gnd cell_6t
Xbit_r103_c181 bl[181] br[181] wl[103] vdd gnd cell_6t
Xbit_r104_c181 bl[181] br[181] wl[104] vdd gnd cell_6t
Xbit_r105_c181 bl[181] br[181] wl[105] vdd gnd cell_6t
Xbit_r106_c181 bl[181] br[181] wl[106] vdd gnd cell_6t
Xbit_r107_c181 bl[181] br[181] wl[107] vdd gnd cell_6t
Xbit_r108_c181 bl[181] br[181] wl[108] vdd gnd cell_6t
Xbit_r109_c181 bl[181] br[181] wl[109] vdd gnd cell_6t
Xbit_r110_c181 bl[181] br[181] wl[110] vdd gnd cell_6t
Xbit_r111_c181 bl[181] br[181] wl[111] vdd gnd cell_6t
Xbit_r112_c181 bl[181] br[181] wl[112] vdd gnd cell_6t
Xbit_r113_c181 bl[181] br[181] wl[113] vdd gnd cell_6t
Xbit_r114_c181 bl[181] br[181] wl[114] vdd gnd cell_6t
Xbit_r115_c181 bl[181] br[181] wl[115] vdd gnd cell_6t
Xbit_r116_c181 bl[181] br[181] wl[116] vdd gnd cell_6t
Xbit_r117_c181 bl[181] br[181] wl[117] vdd gnd cell_6t
Xbit_r118_c181 bl[181] br[181] wl[118] vdd gnd cell_6t
Xbit_r119_c181 bl[181] br[181] wl[119] vdd gnd cell_6t
Xbit_r120_c181 bl[181] br[181] wl[120] vdd gnd cell_6t
Xbit_r121_c181 bl[181] br[181] wl[121] vdd gnd cell_6t
Xbit_r122_c181 bl[181] br[181] wl[122] vdd gnd cell_6t
Xbit_r123_c181 bl[181] br[181] wl[123] vdd gnd cell_6t
Xbit_r124_c181 bl[181] br[181] wl[124] vdd gnd cell_6t
Xbit_r125_c181 bl[181] br[181] wl[125] vdd gnd cell_6t
Xbit_r126_c181 bl[181] br[181] wl[126] vdd gnd cell_6t
Xbit_r127_c181 bl[181] br[181] wl[127] vdd gnd cell_6t
Xbit_r128_c181 bl[181] br[181] wl[128] vdd gnd cell_6t
Xbit_r129_c181 bl[181] br[181] wl[129] vdd gnd cell_6t
Xbit_r130_c181 bl[181] br[181] wl[130] vdd gnd cell_6t
Xbit_r131_c181 bl[181] br[181] wl[131] vdd gnd cell_6t
Xbit_r132_c181 bl[181] br[181] wl[132] vdd gnd cell_6t
Xbit_r133_c181 bl[181] br[181] wl[133] vdd gnd cell_6t
Xbit_r134_c181 bl[181] br[181] wl[134] vdd gnd cell_6t
Xbit_r135_c181 bl[181] br[181] wl[135] vdd gnd cell_6t
Xbit_r136_c181 bl[181] br[181] wl[136] vdd gnd cell_6t
Xbit_r137_c181 bl[181] br[181] wl[137] vdd gnd cell_6t
Xbit_r138_c181 bl[181] br[181] wl[138] vdd gnd cell_6t
Xbit_r139_c181 bl[181] br[181] wl[139] vdd gnd cell_6t
Xbit_r140_c181 bl[181] br[181] wl[140] vdd gnd cell_6t
Xbit_r141_c181 bl[181] br[181] wl[141] vdd gnd cell_6t
Xbit_r142_c181 bl[181] br[181] wl[142] vdd gnd cell_6t
Xbit_r143_c181 bl[181] br[181] wl[143] vdd gnd cell_6t
Xbit_r144_c181 bl[181] br[181] wl[144] vdd gnd cell_6t
Xbit_r145_c181 bl[181] br[181] wl[145] vdd gnd cell_6t
Xbit_r146_c181 bl[181] br[181] wl[146] vdd gnd cell_6t
Xbit_r147_c181 bl[181] br[181] wl[147] vdd gnd cell_6t
Xbit_r148_c181 bl[181] br[181] wl[148] vdd gnd cell_6t
Xbit_r149_c181 bl[181] br[181] wl[149] vdd gnd cell_6t
Xbit_r150_c181 bl[181] br[181] wl[150] vdd gnd cell_6t
Xbit_r151_c181 bl[181] br[181] wl[151] vdd gnd cell_6t
Xbit_r152_c181 bl[181] br[181] wl[152] vdd gnd cell_6t
Xbit_r153_c181 bl[181] br[181] wl[153] vdd gnd cell_6t
Xbit_r154_c181 bl[181] br[181] wl[154] vdd gnd cell_6t
Xbit_r155_c181 bl[181] br[181] wl[155] vdd gnd cell_6t
Xbit_r156_c181 bl[181] br[181] wl[156] vdd gnd cell_6t
Xbit_r157_c181 bl[181] br[181] wl[157] vdd gnd cell_6t
Xbit_r158_c181 bl[181] br[181] wl[158] vdd gnd cell_6t
Xbit_r159_c181 bl[181] br[181] wl[159] vdd gnd cell_6t
Xbit_r160_c181 bl[181] br[181] wl[160] vdd gnd cell_6t
Xbit_r161_c181 bl[181] br[181] wl[161] vdd gnd cell_6t
Xbit_r162_c181 bl[181] br[181] wl[162] vdd gnd cell_6t
Xbit_r163_c181 bl[181] br[181] wl[163] vdd gnd cell_6t
Xbit_r164_c181 bl[181] br[181] wl[164] vdd gnd cell_6t
Xbit_r165_c181 bl[181] br[181] wl[165] vdd gnd cell_6t
Xbit_r166_c181 bl[181] br[181] wl[166] vdd gnd cell_6t
Xbit_r167_c181 bl[181] br[181] wl[167] vdd gnd cell_6t
Xbit_r168_c181 bl[181] br[181] wl[168] vdd gnd cell_6t
Xbit_r169_c181 bl[181] br[181] wl[169] vdd gnd cell_6t
Xbit_r170_c181 bl[181] br[181] wl[170] vdd gnd cell_6t
Xbit_r171_c181 bl[181] br[181] wl[171] vdd gnd cell_6t
Xbit_r172_c181 bl[181] br[181] wl[172] vdd gnd cell_6t
Xbit_r173_c181 bl[181] br[181] wl[173] vdd gnd cell_6t
Xbit_r174_c181 bl[181] br[181] wl[174] vdd gnd cell_6t
Xbit_r175_c181 bl[181] br[181] wl[175] vdd gnd cell_6t
Xbit_r176_c181 bl[181] br[181] wl[176] vdd gnd cell_6t
Xbit_r177_c181 bl[181] br[181] wl[177] vdd gnd cell_6t
Xbit_r178_c181 bl[181] br[181] wl[178] vdd gnd cell_6t
Xbit_r179_c181 bl[181] br[181] wl[179] vdd gnd cell_6t
Xbit_r180_c181 bl[181] br[181] wl[180] vdd gnd cell_6t
Xbit_r181_c181 bl[181] br[181] wl[181] vdd gnd cell_6t
Xbit_r182_c181 bl[181] br[181] wl[182] vdd gnd cell_6t
Xbit_r183_c181 bl[181] br[181] wl[183] vdd gnd cell_6t
Xbit_r184_c181 bl[181] br[181] wl[184] vdd gnd cell_6t
Xbit_r185_c181 bl[181] br[181] wl[185] vdd gnd cell_6t
Xbit_r186_c181 bl[181] br[181] wl[186] vdd gnd cell_6t
Xbit_r187_c181 bl[181] br[181] wl[187] vdd gnd cell_6t
Xbit_r188_c181 bl[181] br[181] wl[188] vdd gnd cell_6t
Xbit_r189_c181 bl[181] br[181] wl[189] vdd gnd cell_6t
Xbit_r190_c181 bl[181] br[181] wl[190] vdd gnd cell_6t
Xbit_r191_c181 bl[181] br[181] wl[191] vdd gnd cell_6t
Xbit_r192_c181 bl[181] br[181] wl[192] vdd gnd cell_6t
Xbit_r193_c181 bl[181] br[181] wl[193] vdd gnd cell_6t
Xbit_r194_c181 bl[181] br[181] wl[194] vdd gnd cell_6t
Xbit_r195_c181 bl[181] br[181] wl[195] vdd gnd cell_6t
Xbit_r196_c181 bl[181] br[181] wl[196] vdd gnd cell_6t
Xbit_r197_c181 bl[181] br[181] wl[197] vdd gnd cell_6t
Xbit_r198_c181 bl[181] br[181] wl[198] vdd gnd cell_6t
Xbit_r199_c181 bl[181] br[181] wl[199] vdd gnd cell_6t
Xbit_r200_c181 bl[181] br[181] wl[200] vdd gnd cell_6t
Xbit_r201_c181 bl[181] br[181] wl[201] vdd gnd cell_6t
Xbit_r202_c181 bl[181] br[181] wl[202] vdd gnd cell_6t
Xbit_r203_c181 bl[181] br[181] wl[203] vdd gnd cell_6t
Xbit_r204_c181 bl[181] br[181] wl[204] vdd gnd cell_6t
Xbit_r205_c181 bl[181] br[181] wl[205] vdd gnd cell_6t
Xbit_r206_c181 bl[181] br[181] wl[206] vdd gnd cell_6t
Xbit_r207_c181 bl[181] br[181] wl[207] vdd gnd cell_6t
Xbit_r208_c181 bl[181] br[181] wl[208] vdd gnd cell_6t
Xbit_r209_c181 bl[181] br[181] wl[209] vdd gnd cell_6t
Xbit_r210_c181 bl[181] br[181] wl[210] vdd gnd cell_6t
Xbit_r211_c181 bl[181] br[181] wl[211] vdd gnd cell_6t
Xbit_r212_c181 bl[181] br[181] wl[212] vdd gnd cell_6t
Xbit_r213_c181 bl[181] br[181] wl[213] vdd gnd cell_6t
Xbit_r214_c181 bl[181] br[181] wl[214] vdd gnd cell_6t
Xbit_r215_c181 bl[181] br[181] wl[215] vdd gnd cell_6t
Xbit_r216_c181 bl[181] br[181] wl[216] vdd gnd cell_6t
Xbit_r217_c181 bl[181] br[181] wl[217] vdd gnd cell_6t
Xbit_r218_c181 bl[181] br[181] wl[218] vdd gnd cell_6t
Xbit_r219_c181 bl[181] br[181] wl[219] vdd gnd cell_6t
Xbit_r220_c181 bl[181] br[181] wl[220] vdd gnd cell_6t
Xbit_r221_c181 bl[181] br[181] wl[221] vdd gnd cell_6t
Xbit_r222_c181 bl[181] br[181] wl[222] vdd gnd cell_6t
Xbit_r223_c181 bl[181] br[181] wl[223] vdd gnd cell_6t
Xbit_r224_c181 bl[181] br[181] wl[224] vdd gnd cell_6t
Xbit_r225_c181 bl[181] br[181] wl[225] vdd gnd cell_6t
Xbit_r226_c181 bl[181] br[181] wl[226] vdd gnd cell_6t
Xbit_r227_c181 bl[181] br[181] wl[227] vdd gnd cell_6t
Xbit_r228_c181 bl[181] br[181] wl[228] vdd gnd cell_6t
Xbit_r229_c181 bl[181] br[181] wl[229] vdd gnd cell_6t
Xbit_r230_c181 bl[181] br[181] wl[230] vdd gnd cell_6t
Xbit_r231_c181 bl[181] br[181] wl[231] vdd gnd cell_6t
Xbit_r232_c181 bl[181] br[181] wl[232] vdd gnd cell_6t
Xbit_r233_c181 bl[181] br[181] wl[233] vdd gnd cell_6t
Xbit_r234_c181 bl[181] br[181] wl[234] vdd gnd cell_6t
Xbit_r235_c181 bl[181] br[181] wl[235] vdd gnd cell_6t
Xbit_r236_c181 bl[181] br[181] wl[236] vdd gnd cell_6t
Xbit_r237_c181 bl[181] br[181] wl[237] vdd gnd cell_6t
Xbit_r238_c181 bl[181] br[181] wl[238] vdd gnd cell_6t
Xbit_r239_c181 bl[181] br[181] wl[239] vdd gnd cell_6t
Xbit_r240_c181 bl[181] br[181] wl[240] vdd gnd cell_6t
Xbit_r241_c181 bl[181] br[181] wl[241] vdd gnd cell_6t
Xbit_r242_c181 bl[181] br[181] wl[242] vdd gnd cell_6t
Xbit_r243_c181 bl[181] br[181] wl[243] vdd gnd cell_6t
Xbit_r244_c181 bl[181] br[181] wl[244] vdd gnd cell_6t
Xbit_r245_c181 bl[181] br[181] wl[245] vdd gnd cell_6t
Xbit_r246_c181 bl[181] br[181] wl[246] vdd gnd cell_6t
Xbit_r247_c181 bl[181] br[181] wl[247] vdd gnd cell_6t
Xbit_r248_c181 bl[181] br[181] wl[248] vdd gnd cell_6t
Xbit_r249_c181 bl[181] br[181] wl[249] vdd gnd cell_6t
Xbit_r250_c181 bl[181] br[181] wl[250] vdd gnd cell_6t
Xbit_r251_c181 bl[181] br[181] wl[251] vdd gnd cell_6t
Xbit_r252_c181 bl[181] br[181] wl[252] vdd gnd cell_6t
Xbit_r253_c181 bl[181] br[181] wl[253] vdd gnd cell_6t
Xbit_r254_c181 bl[181] br[181] wl[254] vdd gnd cell_6t
Xbit_r255_c181 bl[181] br[181] wl[255] vdd gnd cell_6t
Xbit_r0_c182 bl[182] br[182] wl[0] vdd gnd cell_6t
Xbit_r1_c182 bl[182] br[182] wl[1] vdd gnd cell_6t
Xbit_r2_c182 bl[182] br[182] wl[2] vdd gnd cell_6t
Xbit_r3_c182 bl[182] br[182] wl[3] vdd gnd cell_6t
Xbit_r4_c182 bl[182] br[182] wl[4] vdd gnd cell_6t
Xbit_r5_c182 bl[182] br[182] wl[5] vdd gnd cell_6t
Xbit_r6_c182 bl[182] br[182] wl[6] vdd gnd cell_6t
Xbit_r7_c182 bl[182] br[182] wl[7] vdd gnd cell_6t
Xbit_r8_c182 bl[182] br[182] wl[8] vdd gnd cell_6t
Xbit_r9_c182 bl[182] br[182] wl[9] vdd gnd cell_6t
Xbit_r10_c182 bl[182] br[182] wl[10] vdd gnd cell_6t
Xbit_r11_c182 bl[182] br[182] wl[11] vdd gnd cell_6t
Xbit_r12_c182 bl[182] br[182] wl[12] vdd gnd cell_6t
Xbit_r13_c182 bl[182] br[182] wl[13] vdd gnd cell_6t
Xbit_r14_c182 bl[182] br[182] wl[14] vdd gnd cell_6t
Xbit_r15_c182 bl[182] br[182] wl[15] vdd gnd cell_6t
Xbit_r16_c182 bl[182] br[182] wl[16] vdd gnd cell_6t
Xbit_r17_c182 bl[182] br[182] wl[17] vdd gnd cell_6t
Xbit_r18_c182 bl[182] br[182] wl[18] vdd gnd cell_6t
Xbit_r19_c182 bl[182] br[182] wl[19] vdd gnd cell_6t
Xbit_r20_c182 bl[182] br[182] wl[20] vdd gnd cell_6t
Xbit_r21_c182 bl[182] br[182] wl[21] vdd gnd cell_6t
Xbit_r22_c182 bl[182] br[182] wl[22] vdd gnd cell_6t
Xbit_r23_c182 bl[182] br[182] wl[23] vdd gnd cell_6t
Xbit_r24_c182 bl[182] br[182] wl[24] vdd gnd cell_6t
Xbit_r25_c182 bl[182] br[182] wl[25] vdd gnd cell_6t
Xbit_r26_c182 bl[182] br[182] wl[26] vdd gnd cell_6t
Xbit_r27_c182 bl[182] br[182] wl[27] vdd gnd cell_6t
Xbit_r28_c182 bl[182] br[182] wl[28] vdd gnd cell_6t
Xbit_r29_c182 bl[182] br[182] wl[29] vdd gnd cell_6t
Xbit_r30_c182 bl[182] br[182] wl[30] vdd gnd cell_6t
Xbit_r31_c182 bl[182] br[182] wl[31] vdd gnd cell_6t
Xbit_r32_c182 bl[182] br[182] wl[32] vdd gnd cell_6t
Xbit_r33_c182 bl[182] br[182] wl[33] vdd gnd cell_6t
Xbit_r34_c182 bl[182] br[182] wl[34] vdd gnd cell_6t
Xbit_r35_c182 bl[182] br[182] wl[35] vdd gnd cell_6t
Xbit_r36_c182 bl[182] br[182] wl[36] vdd gnd cell_6t
Xbit_r37_c182 bl[182] br[182] wl[37] vdd gnd cell_6t
Xbit_r38_c182 bl[182] br[182] wl[38] vdd gnd cell_6t
Xbit_r39_c182 bl[182] br[182] wl[39] vdd gnd cell_6t
Xbit_r40_c182 bl[182] br[182] wl[40] vdd gnd cell_6t
Xbit_r41_c182 bl[182] br[182] wl[41] vdd gnd cell_6t
Xbit_r42_c182 bl[182] br[182] wl[42] vdd gnd cell_6t
Xbit_r43_c182 bl[182] br[182] wl[43] vdd gnd cell_6t
Xbit_r44_c182 bl[182] br[182] wl[44] vdd gnd cell_6t
Xbit_r45_c182 bl[182] br[182] wl[45] vdd gnd cell_6t
Xbit_r46_c182 bl[182] br[182] wl[46] vdd gnd cell_6t
Xbit_r47_c182 bl[182] br[182] wl[47] vdd gnd cell_6t
Xbit_r48_c182 bl[182] br[182] wl[48] vdd gnd cell_6t
Xbit_r49_c182 bl[182] br[182] wl[49] vdd gnd cell_6t
Xbit_r50_c182 bl[182] br[182] wl[50] vdd gnd cell_6t
Xbit_r51_c182 bl[182] br[182] wl[51] vdd gnd cell_6t
Xbit_r52_c182 bl[182] br[182] wl[52] vdd gnd cell_6t
Xbit_r53_c182 bl[182] br[182] wl[53] vdd gnd cell_6t
Xbit_r54_c182 bl[182] br[182] wl[54] vdd gnd cell_6t
Xbit_r55_c182 bl[182] br[182] wl[55] vdd gnd cell_6t
Xbit_r56_c182 bl[182] br[182] wl[56] vdd gnd cell_6t
Xbit_r57_c182 bl[182] br[182] wl[57] vdd gnd cell_6t
Xbit_r58_c182 bl[182] br[182] wl[58] vdd gnd cell_6t
Xbit_r59_c182 bl[182] br[182] wl[59] vdd gnd cell_6t
Xbit_r60_c182 bl[182] br[182] wl[60] vdd gnd cell_6t
Xbit_r61_c182 bl[182] br[182] wl[61] vdd gnd cell_6t
Xbit_r62_c182 bl[182] br[182] wl[62] vdd gnd cell_6t
Xbit_r63_c182 bl[182] br[182] wl[63] vdd gnd cell_6t
Xbit_r64_c182 bl[182] br[182] wl[64] vdd gnd cell_6t
Xbit_r65_c182 bl[182] br[182] wl[65] vdd gnd cell_6t
Xbit_r66_c182 bl[182] br[182] wl[66] vdd gnd cell_6t
Xbit_r67_c182 bl[182] br[182] wl[67] vdd gnd cell_6t
Xbit_r68_c182 bl[182] br[182] wl[68] vdd gnd cell_6t
Xbit_r69_c182 bl[182] br[182] wl[69] vdd gnd cell_6t
Xbit_r70_c182 bl[182] br[182] wl[70] vdd gnd cell_6t
Xbit_r71_c182 bl[182] br[182] wl[71] vdd gnd cell_6t
Xbit_r72_c182 bl[182] br[182] wl[72] vdd gnd cell_6t
Xbit_r73_c182 bl[182] br[182] wl[73] vdd gnd cell_6t
Xbit_r74_c182 bl[182] br[182] wl[74] vdd gnd cell_6t
Xbit_r75_c182 bl[182] br[182] wl[75] vdd gnd cell_6t
Xbit_r76_c182 bl[182] br[182] wl[76] vdd gnd cell_6t
Xbit_r77_c182 bl[182] br[182] wl[77] vdd gnd cell_6t
Xbit_r78_c182 bl[182] br[182] wl[78] vdd gnd cell_6t
Xbit_r79_c182 bl[182] br[182] wl[79] vdd gnd cell_6t
Xbit_r80_c182 bl[182] br[182] wl[80] vdd gnd cell_6t
Xbit_r81_c182 bl[182] br[182] wl[81] vdd gnd cell_6t
Xbit_r82_c182 bl[182] br[182] wl[82] vdd gnd cell_6t
Xbit_r83_c182 bl[182] br[182] wl[83] vdd gnd cell_6t
Xbit_r84_c182 bl[182] br[182] wl[84] vdd gnd cell_6t
Xbit_r85_c182 bl[182] br[182] wl[85] vdd gnd cell_6t
Xbit_r86_c182 bl[182] br[182] wl[86] vdd gnd cell_6t
Xbit_r87_c182 bl[182] br[182] wl[87] vdd gnd cell_6t
Xbit_r88_c182 bl[182] br[182] wl[88] vdd gnd cell_6t
Xbit_r89_c182 bl[182] br[182] wl[89] vdd gnd cell_6t
Xbit_r90_c182 bl[182] br[182] wl[90] vdd gnd cell_6t
Xbit_r91_c182 bl[182] br[182] wl[91] vdd gnd cell_6t
Xbit_r92_c182 bl[182] br[182] wl[92] vdd gnd cell_6t
Xbit_r93_c182 bl[182] br[182] wl[93] vdd gnd cell_6t
Xbit_r94_c182 bl[182] br[182] wl[94] vdd gnd cell_6t
Xbit_r95_c182 bl[182] br[182] wl[95] vdd gnd cell_6t
Xbit_r96_c182 bl[182] br[182] wl[96] vdd gnd cell_6t
Xbit_r97_c182 bl[182] br[182] wl[97] vdd gnd cell_6t
Xbit_r98_c182 bl[182] br[182] wl[98] vdd gnd cell_6t
Xbit_r99_c182 bl[182] br[182] wl[99] vdd gnd cell_6t
Xbit_r100_c182 bl[182] br[182] wl[100] vdd gnd cell_6t
Xbit_r101_c182 bl[182] br[182] wl[101] vdd gnd cell_6t
Xbit_r102_c182 bl[182] br[182] wl[102] vdd gnd cell_6t
Xbit_r103_c182 bl[182] br[182] wl[103] vdd gnd cell_6t
Xbit_r104_c182 bl[182] br[182] wl[104] vdd gnd cell_6t
Xbit_r105_c182 bl[182] br[182] wl[105] vdd gnd cell_6t
Xbit_r106_c182 bl[182] br[182] wl[106] vdd gnd cell_6t
Xbit_r107_c182 bl[182] br[182] wl[107] vdd gnd cell_6t
Xbit_r108_c182 bl[182] br[182] wl[108] vdd gnd cell_6t
Xbit_r109_c182 bl[182] br[182] wl[109] vdd gnd cell_6t
Xbit_r110_c182 bl[182] br[182] wl[110] vdd gnd cell_6t
Xbit_r111_c182 bl[182] br[182] wl[111] vdd gnd cell_6t
Xbit_r112_c182 bl[182] br[182] wl[112] vdd gnd cell_6t
Xbit_r113_c182 bl[182] br[182] wl[113] vdd gnd cell_6t
Xbit_r114_c182 bl[182] br[182] wl[114] vdd gnd cell_6t
Xbit_r115_c182 bl[182] br[182] wl[115] vdd gnd cell_6t
Xbit_r116_c182 bl[182] br[182] wl[116] vdd gnd cell_6t
Xbit_r117_c182 bl[182] br[182] wl[117] vdd gnd cell_6t
Xbit_r118_c182 bl[182] br[182] wl[118] vdd gnd cell_6t
Xbit_r119_c182 bl[182] br[182] wl[119] vdd gnd cell_6t
Xbit_r120_c182 bl[182] br[182] wl[120] vdd gnd cell_6t
Xbit_r121_c182 bl[182] br[182] wl[121] vdd gnd cell_6t
Xbit_r122_c182 bl[182] br[182] wl[122] vdd gnd cell_6t
Xbit_r123_c182 bl[182] br[182] wl[123] vdd gnd cell_6t
Xbit_r124_c182 bl[182] br[182] wl[124] vdd gnd cell_6t
Xbit_r125_c182 bl[182] br[182] wl[125] vdd gnd cell_6t
Xbit_r126_c182 bl[182] br[182] wl[126] vdd gnd cell_6t
Xbit_r127_c182 bl[182] br[182] wl[127] vdd gnd cell_6t
Xbit_r128_c182 bl[182] br[182] wl[128] vdd gnd cell_6t
Xbit_r129_c182 bl[182] br[182] wl[129] vdd gnd cell_6t
Xbit_r130_c182 bl[182] br[182] wl[130] vdd gnd cell_6t
Xbit_r131_c182 bl[182] br[182] wl[131] vdd gnd cell_6t
Xbit_r132_c182 bl[182] br[182] wl[132] vdd gnd cell_6t
Xbit_r133_c182 bl[182] br[182] wl[133] vdd gnd cell_6t
Xbit_r134_c182 bl[182] br[182] wl[134] vdd gnd cell_6t
Xbit_r135_c182 bl[182] br[182] wl[135] vdd gnd cell_6t
Xbit_r136_c182 bl[182] br[182] wl[136] vdd gnd cell_6t
Xbit_r137_c182 bl[182] br[182] wl[137] vdd gnd cell_6t
Xbit_r138_c182 bl[182] br[182] wl[138] vdd gnd cell_6t
Xbit_r139_c182 bl[182] br[182] wl[139] vdd gnd cell_6t
Xbit_r140_c182 bl[182] br[182] wl[140] vdd gnd cell_6t
Xbit_r141_c182 bl[182] br[182] wl[141] vdd gnd cell_6t
Xbit_r142_c182 bl[182] br[182] wl[142] vdd gnd cell_6t
Xbit_r143_c182 bl[182] br[182] wl[143] vdd gnd cell_6t
Xbit_r144_c182 bl[182] br[182] wl[144] vdd gnd cell_6t
Xbit_r145_c182 bl[182] br[182] wl[145] vdd gnd cell_6t
Xbit_r146_c182 bl[182] br[182] wl[146] vdd gnd cell_6t
Xbit_r147_c182 bl[182] br[182] wl[147] vdd gnd cell_6t
Xbit_r148_c182 bl[182] br[182] wl[148] vdd gnd cell_6t
Xbit_r149_c182 bl[182] br[182] wl[149] vdd gnd cell_6t
Xbit_r150_c182 bl[182] br[182] wl[150] vdd gnd cell_6t
Xbit_r151_c182 bl[182] br[182] wl[151] vdd gnd cell_6t
Xbit_r152_c182 bl[182] br[182] wl[152] vdd gnd cell_6t
Xbit_r153_c182 bl[182] br[182] wl[153] vdd gnd cell_6t
Xbit_r154_c182 bl[182] br[182] wl[154] vdd gnd cell_6t
Xbit_r155_c182 bl[182] br[182] wl[155] vdd gnd cell_6t
Xbit_r156_c182 bl[182] br[182] wl[156] vdd gnd cell_6t
Xbit_r157_c182 bl[182] br[182] wl[157] vdd gnd cell_6t
Xbit_r158_c182 bl[182] br[182] wl[158] vdd gnd cell_6t
Xbit_r159_c182 bl[182] br[182] wl[159] vdd gnd cell_6t
Xbit_r160_c182 bl[182] br[182] wl[160] vdd gnd cell_6t
Xbit_r161_c182 bl[182] br[182] wl[161] vdd gnd cell_6t
Xbit_r162_c182 bl[182] br[182] wl[162] vdd gnd cell_6t
Xbit_r163_c182 bl[182] br[182] wl[163] vdd gnd cell_6t
Xbit_r164_c182 bl[182] br[182] wl[164] vdd gnd cell_6t
Xbit_r165_c182 bl[182] br[182] wl[165] vdd gnd cell_6t
Xbit_r166_c182 bl[182] br[182] wl[166] vdd gnd cell_6t
Xbit_r167_c182 bl[182] br[182] wl[167] vdd gnd cell_6t
Xbit_r168_c182 bl[182] br[182] wl[168] vdd gnd cell_6t
Xbit_r169_c182 bl[182] br[182] wl[169] vdd gnd cell_6t
Xbit_r170_c182 bl[182] br[182] wl[170] vdd gnd cell_6t
Xbit_r171_c182 bl[182] br[182] wl[171] vdd gnd cell_6t
Xbit_r172_c182 bl[182] br[182] wl[172] vdd gnd cell_6t
Xbit_r173_c182 bl[182] br[182] wl[173] vdd gnd cell_6t
Xbit_r174_c182 bl[182] br[182] wl[174] vdd gnd cell_6t
Xbit_r175_c182 bl[182] br[182] wl[175] vdd gnd cell_6t
Xbit_r176_c182 bl[182] br[182] wl[176] vdd gnd cell_6t
Xbit_r177_c182 bl[182] br[182] wl[177] vdd gnd cell_6t
Xbit_r178_c182 bl[182] br[182] wl[178] vdd gnd cell_6t
Xbit_r179_c182 bl[182] br[182] wl[179] vdd gnd cell_6t
Xbit_r180_c182 bl[182] br[182] wl[180] vdd gnd cell_6t
Xbit_r181_c182 bl[182] br[182] wl[181] vdd gnd cell_6t
Xbit_r182_c182 bl[182] br[182] wl[182] vdd gnd cell_6t
Xbit_r183_c182 bl[182] br[182] wl[183] vdd gnd cell_6t
Xbit_r184_c182 bl[182] br[182] wl[184] vdd gnd cell_6t
Xbit_r185_c182 bl[182] br[182] wl[185] vdd gnd cell_6t
Xbit_r186_c182 bl[182] br[182] wl[186] vdd gnd cell_6t
Xbit_r187_c182 bl[182] br[182] wl[187] vdd gnd cell_6t
Xbit_r188_c182 bl[182] br[182] wl[188] vdd gnd cell_6t
Xbit_r189_c182 bl[182] br[182] wl[189] vdd gnd cell_6t
Xbit_r190_c182 bl[182] br[182] wl[190] vdd gnd cell_6t
Xbit_r191_c182 bl[182] br[182] wl[191] vdd gnd cell_6t
Xbit_r192_c182 bl[182] br[182] wl[192] vdd gnd cell_6t
Xbit_r193_c182 bl[182] br[182] wl[193] vdd gnd cell_6t
Xbit_r194_c182 bl[182] br[182] wl[194] vdd gnd cell_6t
Xbit_r195_c182 bl[182] br[182] wl[195] vdd gnd cell_6t
Xbit_r196_c182 bl[182] br[182] wl[196] vdd gnd cell_6t
Xbit_r197_c182 bl[182] br[182] wl[197] vdd gnd cell_6t
Xbit_r198_c182 bl[182] br[182] wl[198] vdd gnd cell_6t
Xbit_r199_c182 bl[182] br[182] wl[199] vdd gnd cell_6t
Xbit_r200_c182 bl[182] br[182] wl[200] vdd gnd cell_6t
Xbit_r201_c182 bl[182] br[182] wl[201] vdd gnd cell_6t
Xbit_r202_c182 bl[182] br[182] wl[202] vdd gnd cell_6t
Xbit_r203_c182 bl[182] br[182] wl[203] vdd gnd cell_6t
Xbit_r204_c182 bl[182] br[182] wl[204] vdd gnd cell_6t
Xbit_r205_c182 bl[182] br[182] wl[205] vdd gnd cell_6t
Xbit_r206_c182 bl[182] br[182] wl[206] vdd gnd cell_6t
Xbit_r207_c182 bl[182] br[182] wl[207] vdd gnd cell_6t
Xbit_r208_c182 bl[182] br[182] wl[208] vdd gnd cell_6t
Xbit_r209_c182 bl[182] br[182] wl[209] vdd gnd cell_6t
Xbit_r210_c182 bl[182] br[182] wl[210] vdd gnd cell_6t
Xbit_r211_c182 bl[182] br[182] wl[211] vdd gnd cell_6t
Xbit_r212_c182 bl[182] br[182] wl[212] vdd gnd cell_6t
Xbit_r213_c182 bl[182] br[182] wl[213] vdd gnd cell_6t
Xbit_r214_c182 bl[182] br[182] wl[214] vdd gnd cell_6t
Xbit_r215_c182 bl[182] br[182] wl[215] vdd gnd cell_6t
Xbit_r216_c182 bl[182] br[182] wl[216] vdd gnd cell_6t
Xbit_r217_c182 bl[182] br[182] wl[217] vdd gnd cell_6t
Xbit_r218_c182 bl[182] br[182] wl[218] vdd gnd cell_6t
Xbit_r219_c182 bl[182] br[182] wl[219] vdd gnd cell_6t
Xbit_r220_c182 bl[182] br[182] wl[220] vdd gnd cell_6t
Xbit_r221_c182 bl[182] br[182] wl[221] vdd gnd cell_6t
Xbit_r222_c182 bl[182] br[182] wl[222] vdd gnd cell_6t
Xbit_r223_c182 bl[182] br[182] wl[223] vdd gnd cell_6t
Xbit_r224_c182 bl[182] br[182] wl[224] vdd gnd cell_6t
Xbit_r225_c182 bl[182] br[182] wl[225] vdd gnd cell_6t
Xbit_r226_c182 bl[182] br[182] wl[226] vdd gnd cell_6t
Xbit_r227_c182 bl[182] br[182] wl[227] vdd gnd cell_6t
Xbit_r228_c182 bl[182] br[182] wl[228] vdd gnd cell_6t
Xbit_r229_c182 bl[182] br[182] wl[229] vdd gnd cell_6t
Xbit_r230_c182 bl[182] br[182] wl[230] vdd gnd cell_6t
Xbit_r231_c182 bl[182] br[182] wl[231] vdd gnd cell_6t
Xbit_r232_c182 bl[182] br[182] wl[232] vdd gnd cell_6t
Xbit_r233_c182 bl[182] br[182] wl[233] vdd gnd cell_6t
Xbit_r234_c182 bl[182] br[182] wl[234] vdd gnd cell_6t
Xbit_r235_c182 bl[182] br[182] wl[235] vdd gnd cell_6t
Xbit_r236_c182 bl[182] br[182] wl[236] vdd gnd cell_6t
Xbit_r237_c182 bl[182] br[182] wl[237] vdd gnd cell_6t
Xbit_r238_c182 bl[182] br[182] wl[238] vdd gnd cell_6t
Xbit_r239_c182 bl[182] br[182] wl[239] vdd gnd cell_6t
Xbit_r240_c182 bl[182] br[182] wl[240] vdd gnd cell_6t
Xbit_r241_c182 bl[182] br[182] wl[241] vdd gnd cell_6t
Xbit_r242_c182 bl[182] br[182] wl[242] vdd gnd cell_6t
Xbit_r243_c182 bl[182] br[182] wl[243] vdd gnd cell_6t
Xbit_r244_c182 bl[182] br[182] wl[244] vdd gnd cell_6t
Xbit_r245_c182 bl[182] br[182] wl[245] vdd gnd cell_6t
Xbit_r246_c182 bl[182] br[182] wl[246] vdd gnd cell_6t
Xbit_r247_c182 bl[182] br[182] wl[247] vdd gnd cell_6t
Xbit_r248_c182 bl[182] br[182] wl[248] vdd gnd cell_6t
Xbit_r249_c182 bl[182] br[182] wl[249] vdd gnd cell_6t
Xbit_r250_c182 bl[182] br[182] wl[250] vdd gnd cell_6t
Xbit_r251_c182 bl[182] br[182] wl[251] vdd gnd cell_6t
Xbit_r252_c182 bl[182] br[182] wl[252] vdd gnd cell_6t
Xbit_r253_c182 bl[182] br[182] wl[253] vdd gnd cell_6t
Xbit_r254_c182 bl[182] br[182] wl[254] vdd gnd cell_6t
Xbit_r255_c182 bl[182] br[182] wl[255] vdd gnd cell_6t
Xbit_r0_c183 bl[183] br[183] wl[0] vdd gnd cell_6t
Xbit_r1_c183 bl[183] br[183] wl[1] vdd gnd cell_6t
Xbit_r2_c183 bl[183] br[183] wl[2] vdd gnd cell_6t
Xbit_r3_c183 bl[183] br[183] wl[3] vdd gnd cell_6t
Xbit_r4_c183 bl[183] br[183] wl[4] vdd gnd cell_6t
Xbit_r5_c183 bl[183] br[183] wl[5] vdd gnd cell_6t
Xbit_r6_c183 bl[183] br[183] wl[6] vdd gnd cell_6t
Xbit_r7_c183 bl[183] br[183] wl[7] vdd gnd cell_6t
Xbit_r8_c183 bl[183] br[183] wl[8] vdd gnd cell_6t
Xbit_r9_c183 bl[183] br[183] wl[9] vdd gnd cell_6t
Xbit_r10_c183 bl[183] br[183] wl[10] vdd gnd cell_6t
Xbit_r11_c183 bl[183] br[183] wl[11] vdd gnd cell_6t
Xbit_r12_c183 bl[183] br[183] wl[12] vdd gnd cell_6t
Xbit_r13_c183 bl[183] br[183] wl[13] vdd gnd cell_6t
Xbit_r14_c183 bl[183] br[183] wl[14] vdd gnd cell_6t
Xbit_r15_c183 bl[183] br[183] wl[15] vdd gnd cell_6t
Xbit_r16_c183 bl[183] br[183] wl[16] vdd gnd cell_6t
Xbit_r17_c183 bl[183] br[183] wl[17] vdd gnd cell_6t
Xbit_r18_c183 bl[183] br[183] wl[18] vdd gnd cell_6t
Xbit_r19_c183 bl[183] br[183] wl[19] vdd gnd cell_6t
Xbit_r20_c183 bl[183] br[183] wl[20] vdd gnd cell_6t
Xbit_r21_c183 bl[183] br[183] wl[21] vdd gnd cell_6t
Xbit_r22_c183 bl[183] br[183] wl[22] vdd gnd cell_6t
Xbit_r23_c183 bl[183] br[183] wl[23] vdd gnd cell_6t
Xbit_r24_c183 bl[183] br[183] wl[24] vdd gnd cell_6t
Xbit_r25_c183 bl[183] br[183] wl[25] vdd gnd cell_6t
Xbit_r26_c183 bl[183] br[183] wl[26] vdd gnd cell_6t
Xbit_r27_c183 bl[183] br[183] wl[27] vdd gnd cell_6t
Xbit_r28_c183 bl[183] br[183] wl[28] vdd gnd cell_6t
Xbit_r29_c183 bl[183] br[183] wl[29] vdd gnd cell_6t
Xbit_r30_c183 bl[183] br[183] wl[30] vdd gnd cell_6t
Xbit_r31_c183 bl[183] br[183] wl[31] vdd gnd cell_6t
Xbit_r32_c183 bl[183] br[183] wl[32] vdd gnd cell_6t
Xbit_r33_c183 bl[183] br[183] wl[33] vdd gnd cell_6t
Xbit_r34_c183 bl[183] br[183] wl[34] vdd gnd cell_6t
Xbit_r35_c183 bl[183] br[183] wl[35] vdd gnd cell_6t
Xbit_r36_c183 bl[183] br[183] wl[36] vdd gnd cell_6t
Xbit_r37_c183 bl[183] br[183] wl[37] vdd gnd cell_6t
Xbit_r38_c183 bl[183] br[183] wl[38] vdd gnd cell_6t
Xbit_r39_c183 bl[183] br[183] wl[39] vdd gnd cell_6t
Xbit_r40_c183 bl[183] br[183] wl[40] vdd gnd cell_6t
Xbit_r41_c183 bl[183] br[183] wl[41] vdd gnd cell_6t
Xbit_r42_c183 bl[183] br[183] wl[42] vdd gnd cell_6t
Xbit_r43_c183 bl[183] br[183] wl[43] vdd gnd cell_6t
Xbit_r44_c183 bl[183] br[183] wl[44] vdd gnd cell_6t
Xbit_r45_c183 bl[183] br[183] wl[45] vdd gnd cell_6t
Xbit_r46_c183 bl[183] br[183] wl[46] vdd gnd cell_6t
Xbit_r47_c183 bl[183] br[183] wl[47] vdd gnd cell_6t
Xbit_r48_c183 bl[183] br[183] wl[48] vdd gnd cell_6t
Xbit_r49_c183 bl[183] br[183] wl[49] vdd gnd cell_6t
Xbit_r50_c183 bl[183] br[183] wl[50] vdd gnd cell_6t
Xbit_r51_c183 bl[183] br[183] wl[51] vdd gnd cell_6t
Xbit_r52_c183 bl[183] br[183] wl[52] vdd gnd cell_6t
Xbit_r53_c183 bl[183] br[183] wl[53] vdd gnd cell_6t
Xbit_r54_c183 bl[183] br[183] wl[54] vdd gnd cell_6t
Xbit_r55_c183 bl[183] br[183] wl[55] vdd gnd cell_6t
Xbit_r56_c183 bl[183] br[183] wl[56] vdd gnd cell_6t
Xbit_r57_c183 bl[183] br[183] wl[57] vdd gnd cell_6t
Xbit_r58_c183 bl[183] br[183] wl[58] vdd gnd cell_6t
Xbit_r59_c183 bl[183] br[183] wl[59] vdd gnd cell_6t
Xbit_r60_c183 bl[183] br[183] wl[60] vdd gnd cell_6t
Xbit_r61_c183 bl[183] br[183] wl[61] vdd gnd cell_6t
Xbit_r62_c183 bl[183] br[183] wl[62] vdd gnd cell_6t
Xbit_r63_c183 bl[183] br[183] wl[63] vdd gnd cell_6t
Xbit_r64_c183 bl[183] br[183] wl[64] vdd gnd cell_6t
Xbit_r65_c183 bl[183] br[183] wl[65] vdd gnd cell_6t
Xbit_r66_c183 bl[183] br[183] wl[66] vdd gnd cell_6t
Xbit_r67_c183 bl[183] br[183] wl[67] vdd gnd cell_6t
Xbit_r68_c183 bl[183] br[183] wl[68] vdd gnd cell_6t
Xbit_r69_c183 bl[183] br[183] wl[69] vdd gnd cell_6t
Xbit_r70_c183 bl[183] br[183] wl[70] vdd gnd cell_6t
Xbit_r71_c183 bl[183] br[183] wl[71] vdd gnd cell_6t
Xbit_r72_c183 bl[183] br[183] wl[72] vdd gnd cell_6t
Xbit_r73_c183 bl[183] br[183] wl[73] vdd gnd cell_6t
Xbit_r74_c183 bl[183] br[183] wl[74] vdd gnd cell_6t
Xbit_r75_c183 bl[183] br[183] wl[75] vdd gnd cell_6t
Xbit_r76_c183 bl[183] br[183] wl[76] vdd gnd cell_6t
Xbit_r77_c183 bl[183] br[183] wl[77] vdd gnd cell_6t
Xbit_r78_c183 bl[183] br[183] wl[78] vdd gnd cell_6t
Xbit_r79_c183 bl[183] br[183] wl[79] vdd gnd cell_6t
Xbit_r80_c183 bl[183] br[183] wl[80] vdd gnd cell_6t
Xbit_r81_c183 bl[183] br[183] wl[81] vdd gnd cell_6t
Xbit_r82_c183 bl[183] br[183] wl[82] vdd gnd cell_6t
Xbit_r83_c183 bl[183] br[183] wl[83] vdd gnd cell_6t
Xbit_r84_c183 bl[183] br[183] wl[84] vdd gnd cell_6t
Xbit_r85_c183 bl[183] br[183] wl[85] vdd gnd cell_6t
Xbit_r86_c183 bl[183] br[183] wl[86] vdd gnd cell_6t
Xbit_r87_c183 bl[183] br[183] wl[87] vdd gnd cell_6t
Xbit_r88_c183 bl[183] br[183] wl[88] vdd gnd cell_6t
Xbit_r89_c183 bl[183] br[183] wl[89] vdd gnd cell_6t
Xbit_r90_c183 bl[183] br[183] wl[90] vdd gnd cell_6t
Xbit_r91_c183 bl[183] br[183] wl[91] vdd gnd cell_6t
Xbit_r92_c183 bl[183] br[183] wl[92] vdd gnd cell_6t
Xbit_r93_c183 bl[183] br[183] wl[93] vdd gnd cell_6t
Xbit_r94_c183 bl[183] br[183] wl[94] vdd gnd cell_6t
Xbit_r95_c183 bl[183] br[183] wl[95] vdd gnd cell_6t
Xbit_r96_c183 bl[183] br[183] wl[96] vdd gnd cell_6t
Xbit_r97_c183 bl[183] br[183] wl[97] vdd gnd cell_6t
Xbit_r98_c183 bl[183] br[183] wl[98] vdd gnd cell_6t
Xbit_r99_c183 bl[183] br[183] wl[99] vdd gnd cell_6t
Xbit_r100_c183 bl[183] br[183] wl[100] vdd gnd cell_6t
Xbit_r101_c183 bl[183] br[183] wl[101] vdd gnd cell_6t
Xbit_r102_c183 bl[183] br[183] wl[102] vdd gnd cell_6t
Xbit_r103_c183 bl[183] br[183] wl[103] vdd gnd cell_6t
Xbit_r104_c183 bl[183] br[183] wl[104] vdd gnd cell_6t
Xbit_r105_c183 bl[183] br[183] wl[105] vdd gnd cell_6t
Xbit_r106_c183 bl[183] br[183] wl[106] vdd gnd cell_6t
Xbit_r107_c183 bl[183] br[183] wl[107] vdd gnd cell_6t
Xbit_r108_c183 bl[183] br[183] wl[108] vdd gnd cell_6t
Xbit_r109_c183 bl[183] br[183] wl[109] vdd gnd cell_6t
Xbit_r110_c183 bl[183] br[183] wl[110] vdd gnd cell_6t
Xbit_r111_c183 bl[183] br[183] wl[111] vdd gnd cell_6t
Xbit_r112_c183 bl[183] br[183] wl[112] vdd gnd cell_6t
Xbit_r113_c183 bl[183] br[183] wl[113] vdd gnd cell_6t
Xbit_r114_c183 bl[183] br[183] wl[114] vdd gnd cell_6t
Xbit_r115_c183 bl[183] br[183] wl[115] vdd gnd cell_6t
Xbit_r116_c183 bl[183] br[183] wl[116] vdd gnd cell_6t
Xbit_r117_c183 bl[183] br[183] wl[117] vdd gnd cell_6t
Xbit_r118_c183 bl[183] br[183] wl[118] vdd gnd cell_6t
Xbit_r119_c183 bl[183] br[183] wl[119] vdd gnd cell_6t
Xbit_r120_c183 bl[183] br[183] wl[120] vdd gnd cell_6t
Xbit_r121_c183 bl[183] br[183] wl[121] vdd gnd cell_6t
Xbit_r122_c183 bl[183] br[183] wl[122] vdd gnd cell_6t
Xbit_r123_c183 bl[183] br[183] wl[123] vdd gnd cell_6t
Xbit_r124_c183 bl[183] br[183] wl[124] vdd gnd cell_6t
Xbit_r125_c183 bl[183] br[183] wl[125] vdd gnd cell_6t
Xbit_r126_c183 bl[183] br[183] wl[126] vdd gnd cell_6t
Xbit_r127_c183 bl[183] br[183] wl[127] vdd gnd cell_6t
Xbit_r128_c183 bl[183] br[183] wl[128] vdd gnd cell_6t
Xbit_r129_c183 bl[183] br[183] wl[129] vdd gnd cell_6t
Xbit_r130_c183 bl[183] br[183] wl[130] vdd gnd cell_6t
Xbit_r131_c183 bl[183] br[183] wl[131] vdd gnd cell_6t
Xbit_r132_c183 bl[183] br[183] wl[132] vdd gnd cell_6t
Xbit_r133_c183 bl[183] br[183] wl[133] vdd gnd cell_6t
Xbit_r134_c183 bl[183] br[183] wl[134] vdd gnd cell_6t
Xbit_r135_c183 bl[183] br[183] wl[135] vdd gnd cell_6t
Xbit_r136_c183 bl[183] br[183] wl[136] vdd gnd cell_6t
Xbit_r137_c183 bl[183] br[183] wl[137] vdd gnd cell_6t
Xbit_r138_c183 bl[183] br[183] wl[138] vdd gnd cell_6t
Xbit_r139_c183 bl[183] br[183] wl[139] vdd gnd cell_6t
Xbit_r140_c183 bl[183] br[183] wl[140] vdd gnd cell_6t
Xbit_r141_c183 bl[183] br[183] wl[141] vdd gnd cell_6t
Xbit_r142_c183 bl[183] br[183] wl[142] vdd gnd cell_6t
Xbit_r143_c183 bl[183] br[183] wl[143] vdd gnd cell_6t
Xbit_r144_c183 bl[183] br[183] wl[144] vdd gnd cell_6t
Xbit_r145_c183 bl[183] br[183] wl[145] vdd gnd cell_6t
Xbit_r146_c183 bl[183] br[183] wl[146] vdd gnd cell_6t
Xbit_r147_c183 bl[183] br[183] wl[147] vdd gnd cell_6t
Xbit_r148_c183 bl[183] br[183] wl[148] vdd gnd cell_6t
Xbit_r149_c183 bl[183] br[183] wl[149] vdd gnd cell_6t
Xbit_r150_c183 bl[183] br[183] wl[150] vdd gnd cell_6t
Xbit_r151_c183 bl[183] br[183] wl[151] vdd gnd cell_6t
Xbit_r152_c183 bl[183] br[183] wl[152] vdd gnd cell_6t
Xbit_r153_c183 bl[183] br[183] wl[153] vdd gnd cell_6t
Xbit_r154_c183 bl[183] br[183] wl[154] vdd gnd cell_6t
Xbit_r155_c183 bl[183] br[183] wl[155] vdd gnd cell_6t
Xbit_r156_c183 bl[183] br[183] wl[156] vdd gnd cell_6t
Xbit_r157_c183 bl[183] br[183] wl[157] vdd gnd cell_6t
Xbit_r158_c183 bl[183] br[183] wl[158] vdd gnd cell_6t
Xbit_r159_c183 bl[183] br[183] wl[159] vdd gnd cell_6t
Xbit_r160_c183 bl[183] br[183] wl[160] vdd gnd cell_6t
Xbit_r161_c183 bl[183] br[183] wl[161] vdd gnd cell_6t
Xbit_r162_c183 bl[183] br[183] wl[162] vdd gnd cell_6t
Xbit_r163_c183 bl[183] br[183] wl[163] vdd gnd cell_6t
Xbit_r164_c183 bl[183] br[183] wl[164] vdd gnd cell_6t
Xbit_r165_c183 bl[183] br[183] wl[165] vdd gnd cell_6t
Xbit_r166_c183 bl[183] br[183] wl[166] vdd gnd cell_6t
Xbit_r167_c183 bl[183] br[183] wl[167] vdd gnd cell_6t
Xbit_r168_c183 bl[183] br[183] wl[168] vdd gnd cell_6t
Xbit_r169_c183 bl[183] br[183] wl[169] vdd gnd cell_6t
Xbit_r170_c183 bl[183] br[183] wl[170] vdd gnd cell_6t
Xbit_r171_c183 bl[183] br[183] wl[171] vdd gnd cell_6t
Xbit_r172_c183 bl[183] br[183] wl[172] vdd gnd cell_6t
Xbit_r173_c183 bl[183] br[183] wl[173] vdd gnd cell_6t
Xbit_r174_c183 bl[183] br[183] wl[174] vdd gnd cell_6t
Xbit_r175_c183 bl[183] br[183] wl[175] vdd gnd cell_6t
Xbit_r176_c183 bl[183] br[183] wl[176] vdd gnd cell_6t
Xbit_r177_c183 bl[183] br[183] wl[177] vdd gnd cell_6t
Xbit_r178_c183 bl[183] br[183] wl[178] vdd gnd cell_6t
Xbit_r179_c183 bl[183] br[183] wl[179] vdd gnd cell_6t
Xbit_r180_c183 bl[183] br[183] wl[180] vdd gnd cell_6t
Xbit_r181_c183 bl[183] br[183] wl[181] vdd gnd cell_6t
Xbit_r182_c183 bl[183] br[183] wl[182] vdd gnd cell_6t
Xbit_r183_c183 bl[183] br[183] wl[183] vdd gnd cell_6t
Xbit_r184_c183 bl[183] br[183] wl[184] vdd gnd cell_6t
Xbit_r185_c183 bl[183] br[183] wl[185] vdd gnd cell_6t
Xbit_r186_c183 bl[183] br[183] wl[186] vdd gnd cell_6t
Xbit_r187_c183 bl[183] br[183] wl[187] vdd gnd cell_6t
Xbit_r188_c183 bl[183] br[183] wl[188] vdd gnd cell_6t
Xbit_r189_c183 bl[183] br[183] wl[189] vdd gnd cell_6t
Xbit_r190_c183 bl[183] br[183] wl[190] vdd gnd cell_6t
Xbit_r191_c183 bl[183] br[183] wl[191] vdd gnd cell_6t
Xbit_r192_c183 bl[183] br[183] wl[192] vdd gnd cell_6t
Xbit_r193_c183 bl[183] br[183] wl[193] vdd gnd cell_6t
Xbit_r194_c183 bl[183] br[183] wl[194] vdd gnd cell_6t
Xbit_r195_c183 bl[183] br[183] wl[195] vdd gnd cell_6t
Xbit_r196_c183 bl[183] br[183] wl[196] vdd gnd cell_6t
Xbit_r197_c183 bl[183] br[183] wl[197] vdd gnd cell_6t
Xbit_r198_c183 bl[183] br[183] wl[198] vdd gnd cell_6t
Xbit_r199_c183 bl[183] br[183] wl[199] vdd gnd cell_6t
Xbit_r200_c183 bl[183] br[183] wl[200] vdd gnd cell_6t
Xbit_r201_c183 bl[183] br[183] wl[201] vdd gnd cell_6t
Xbit_r202_c183 bl[183] br[183] wl[202] vdd gnd cell_6t
Xbit_r203_c183 bl[183] br[183] wl[203] vdd gnd cell_6t
Xbit_r204_c183 bl[183] br[183] wl[204] vdd gnd cell_6t
Xbit_r205_c183 bl[183] br[183] wl[205] vdd gnd cell_6t
Xbit_r206_c183 bl[183] br[183] wl[206] vdd gnd cell_6t
Xbit_r207_c183 bl[183] br[183] wl[207] vdd gnd cell_6t
Xbit_r208_c183 bl[183] br[183] wl[208] vdd gnd cell_6t
Xbit_r209_c183 bl[183] br[183] wl[209] vdd gnd cell_6t
Xbit_r210_c183 bl[183] br[183] wl[210] vdd gnd cell_6t
Xbit_r211_c183 bl[183] br[183] wl[211] vdd gnd cell_6t
Xbit_r212_c183 bl[183] br[183] wl[212] vdd gnd cell_6t
Xbit_r213_c183 bl[183] br[183] wl[213] vdd gnd cell_6t
Xbit_r214_c183 bl[183] br[183] wl[214] vdd gnd cell_6t
Xbit_r215_c183 bl[183] br[183] wl[215] vdd gnd cell_6t
Xbit_r216_c183 bl[183] br[183] wl[216] vdd gnd cell_6t
Xbit_r217_c183 bl[183] br[183] wl[217] vdd gnd cell_6t
Xbit_r218_c183 bl[183] br[183] wl[218] vdd gnd cell_6t
Xbit_r219_c183 bl[183] br[183] wl[219] vdd gnd cell_6t
Xbit_r220_c183 bl[183] br[183] wl[220] vdd gnd cell_6t
Xbit_r221_c183 bl[183] br[183] wl[221] vdd gnd cell_6t
Xbit_r222_c183 bl[183] br[183] wl[222] vdd gnd cell_6t
Xbit_r223_c183 bl[183] br[183] wl[223] vdd gnd cell_6t
Xbit_r224_c183 bl[183] br[183] wl[224] vdd gnd cell_6t
Xbit_r225_c183 bl[183] br[183] wl[225] vdd gnd cell_6t
Xbit_r226_c183 bl[183] br[183] wl[226] vdd gnd cell_6t
Xbit_r227_c183 bl[183] br[183] wl[227] vdd gnd cell_6t
Xbit_r228_c183 bl[183] br[183] wl[228] vdd gnd cell_6t
Xbit_r229_c183 bl[183] br[183] wl[229] vdd gnd cell_6t
Xbit_r230_c183 bl[183] br[183] wl[230] vdd gnd cell_6t
Xbit_r231_c183 bl[183] br[183] wl[231] vdd gnd cell_6t
Xbit_r232_c183 bl[183] br[183] wl[232] vdd gnd cell_6t
Xbit_r233_c183 bl[183] br[183] wl[233] vdd gnd cell_6t
Xbit_r234_c183 bl[183] br[183] wl[234] vdd gnd cell_6t
Xbit_r235_c183 bl[183] br[183] wl[235] vdd gnd cell_6t
Xbit_r236_c183 bl[183] br[183] wl[236] vdd gnd cell_6t
Xbit_r237_c183 bl[183] br[183] wl[237] vdd gnd cell_6t
Xbit_r238_c183 bl[183] br[183] wl[238] vdd gnd cell_6t
Xbit_r239_c183 bl[183] br[183] wl[239] vdd gnd cell_6t
Xbit_r240_c183 bl[183] br[183] wl[240] vdd gnd cell_6t
Xbit_r241_c183 bl[183] br[183] wl[241] vdd gnd cell_6t
Xbit_r242_c183 bl[183] br[183] wl[242] vdd gnd cell_6t
Xbit_r243_c183 bl[183] br[183] wl[243] vdd gnd cell_6t
Xbit_r244_c183 bl[183] br[183] wl[244] vdd gnd cell_6t
Xbit_r245_c183 bl[183] br[183] wl[245] vdd gnd cell_6t
Xbit_r246_c183 bl[183] br[183] wl[246] vdd gnd cell_6t
Xbit_r247_c183 bl[183] br[183] wl[247] vdd gnd cell_6t
Xbit_r248_c183 bl[183] br[183] wl[248] vdd gnd cell_6t
Xbit_r249_c183 bl[183] br[183] wl[249] vdd gnd cell_6t
Xbit_r250_c183 bl[183] br[183] wl[250] vdd gnd cell_6t
Xbit_r251_c183 bl[183] br[183] wl[251] vdd gnd cell_6t
Xbit_r252_c183 bl[183] br[183] wl[252] vdd gnd cell_6t
Xbit_r253_c183 bl[183] br[183] wl[253] vdd gnd cell_6t
Xbit_r254_c183 bl[183] br[183] wl[254] vdd gnd cell_6t
Xbit_r255_c183 bl[183] br[183] wl[255] vdd gnd cell_6t
Xbit_r0_c184 bl[184] br[184] wl[0] vdd gnd cell_6t
Xbit_r1_c184 bl[184] br[184] wl[1] vdd gnd cell_6t
Xbit_r2_c184 bl[184] br[184] wl[2] vdd gnd cell_6t
Xbit_r3_c184 bl[184] br[184] wl[3] vdd gnd cell_6t
Xbit_r4_c184 bl[184] br[184] wl[4] vdd gnd cell_6t
Xbit_r5_c184 bl[184] br[184] wl[5] vdd gnd cell_6t
Xbit_r6_c184 bl[184] br[184] wl[6] vdd gnd cell_6t
Xbit_r7_c184 bl[184] br[184] wl[7] vdd gnd cell_6t
Xbit_r8_c184 bl[184] br[184] wl[8] vdd gnd cell_6t
Xbit_r9_c184 bl[184] br[184] wl[9] vdd gnd cell_6t
Xbit_r10_c184 bl[184] br[184] wl[10] vdd gnd cell_6t
Xbit_r11_c184 bl[184] br[184] wl[11] vdd gnd cell_6t
Xbit_r12_c184 bl[184] br[184] wl[12] vdd gnd cell_6t
Xbit_r13_c184 bl[184] br[184] wl[13] vdd gnd cell_6t
Xbit_r14_c184 bl[184] br[184] wl[14] vdd gnd cell_6t
Xbit_r15_c184 bl[184] br[184] wl[15] vdd gnd cell_6t
Xbit_r16_c184 bl[184] br[184] wl[16] vdd gnd cell_6t
Xbit_r17_c184 bl[184] br[184] wl[17] vdd gnd cell_6t
Xbit_r18_c184 bl[184] br[184] wl[18] vdd gnd cell_6t
Xbit_r19_c184 bl[184] br[184] wl[19] vdd gnd cell_6t
Xbit_r20_c184 bl[184] br[184] wl[20] vdd gnd cell_6t
Xbit_r21_c184 bl[184] br[184] wl[21] vdd gnd cell_6t
Xbit_r22_c184 bl[184] br[184] wl[22] vdd gnd cell_6t
Xbit_r23_c184 bl[184] br[184] wl[23] vdd gnd cell_6t
Xbit_r24_c184 bl[184] br[184] wl[24] vdd gnd cell_6t
Xbit_r25_c184 bl[184] br[184] wl[25] vdd gnd cell_6t
Xbit_r26_c184 bl[184] br[184] wl[26] vdd gnd cell_6t
Xbit_r27_c184 bl[184] br[184] wl[27] vdd gnd cell_6t
Xbit_r28_c184 bl[184] br[184] wl[28] vdd gnd cell_6t
Xbit_r29_c184 bl[184] br[184] wl[29] vdd gnd cell_6t
Xbit_r30_c184 bl[184] br[184] wl[30] vdd gnd cell_6t
Xbit_r31_c184 bl[184] br[184] wl[31] vdd gnd cell_6t
Xbit_r32_c184 bl[184] br[184] wl[32] vdd gnd cell_6t
Xbit_r33_c184 bl[184] br[184] wl[33] vdd gnd cell_6t
Xbit_r34_c184 bl[184] br[184] wl[34] vdd gnd cell_6t
Xbit_r35_c184 bl[184] br[184] wl[35] vdd gnd cell_6t
Xbit_r36_c184 bl[184] br[184] wl[36] vdd gnd cell_6t
Xbit_r37_c184 bl[184] br[184] wl[37] vdd gnd cell_6t
Xbit_r38_c184 bl[184] br[184] wl[38] vdd gnd cell_6t
Xbit_r39_c184 bl[184] br[184] wl[39] vdd gnd cell_6t
Xbit_r40_c184 bl[184] br[184] wl[40] vdd gnd cell_6t
Xbit_r41_c184 bl[184] br[184] wl[41] vdd gnd cell_6t
Xbit_r42_c184 bl[184] br[184] wl[42] vdd gnd cell_6t
Xbit_r43_c184 bl[184] br[184] wl[43] vdd gnd cell_6t
Xbit_r44_c184 bl[184] br[184] wl[44] vdd gnd cell_6t
Xbit_r45_c184 bl[184] br[184] wl[45] vdd gnd cell_6t
Xbit_r46_c184 bl[184] br[184] wl[46] vdd gnd cell_6t
Xbit_r47_c184 bl[184] br[184] wl[47] vdd gnd cell_6t
Xbit_r48_c184 bl[184] br[184] wl[48] vdd gnd cell_6t
Xbit_r49_c184 bl[184] br[184] wl[49] vdd gnd cell_6t
Xbit_r50_c184 bl[184] br[184] wl[50] vdd gnd cell_6t
Xbit_r51_c184 bl[184] br[184] wl[51] vdd gnd cell_6t
Xbit_r52_c184 bl[184] br[184] wl[52] vdd gnd cell_6t
Xbit_r53_c184 bl[184] br[184] wl[53] vdd gnd cell_6t
Xbit_r54_c184 bl[184] br[184] wl[54] vdd gnd cell_6t
Xbit_r55_c184 bl[184] br[184] wl[55] vdd gnd cell_6t
Xbit_r56_c184 bl[184] br[184] wl[56] vdd gnd cell_6t
Xbit_r57_c184 bl[184] br[184] wl[57] vdd gnd cell_6t
Xbit_r58_c184 bl[184] br[184] wl[58] vdd gnd cell_6t
Xbit_r59_c184 bl[184] br[184] wl[59] vdd gnd cell_6t
Xbit_r60_c184 bl[184] br[184] wl[60] vdd gnd cell_6t
Xbit_r61_c184 bl[184] br[184] wl[61] vdd gnd cell_6t
Xbit_r62_c184 bl[184] br[184] wl[62] vdd gnd cell_6t
Xbit_r63_c184 bl[184] br[184] wl[63] vdd gnd cell_6t
Xbit_r64_c184 bl[184] br[184] wl[64] vdd gnd cell_6t
Xbit_r65_c184 bl[184] br[184] wl[65] vdd gnd cell_6t
Xbit_r66_c184 bl[184] br[184] wl[66] vdd gnd cell_6t
Xbit_r67_c184 bl[184] br[184] wl[67] vdd gnd cell_6t
Xbit_r68_c184 bl[184] br[184] wl[68] vdd gnd cell_6t
Xbit_r69_c184 bl[184] br[184] wl[69] vdd gnd cell_6t
Xbit_r70_c184 bl[184] br[184] wl[70] vdd gnd cell_6t
Xbit_r71_c184 bl[184] br[184] wl[71] vdd gnd cell_6t
Xbit_r72_c184 bl[184] br[184] wl[72] vdd gnd cell_6t
Xbit_r73_c184 bl[184] br[184] wl[73] vdd gnd cell_6t
Xbit_r74_c184 bl[184] br[184] wl[74] vdd gnd cell_6t
Xbit_r75_c184 bl[184] br[184] wl[75] vdd gnd cell_6t
Xbit_r76_c184 bl[184] br[184] wl[76] vdd gnd cell_6t
Xbit_r77_c184 bl[184] br[184] wl[77] vdd gnd cell_6t
Xbit_r78_c184 bl[184] br[184] wl[78] vdd gnd cell_6t
Xbit_r79_c184 bl[184] br[184] wl[79] vdd gnd cell_6t
Xbit_r80_c184 bl[184] br[184] wl[80] vdd gnd cell_6t
Xbit_r81_c184 bl[184] br[184] wl[81] vdd gnd cell_6t
Xbit_r82_c184 bl[184] br[184] wl[82] vdd gnd cell_6t
Xbit_r83_c184 bl[184] br[184] wl[83] vdd gnd cell_6t
Xbit_r84_c184 bl[184] br[184] wl[84] vdd gnd cell_6t
Xbit_r85_c184 bl[184] br[184] wl[85] vdd gnd cell_6t
Xbit_r86_c184 bl[184] br[184] wl[86] vdd gnd cell_6t
Xbit_r87_c184 bl[184] br[184] wl[87] vdd gnd cell_6t
Xbit_r88_c184 bl[184] br[184] wl[88] vdd gnd cell_6t
Xbit_r89_c184 bl[184] br[184] wl[89] vdd gnd cell_6t
Xbit_r90_c184 bl[184] br[184] wl[90] vdd gnd cell_6t
Xbit_r91_c184 bl[184] br[184] wl[91] vdd gnd cell_6t
Xbit_r92_c184 bl[184] br[184] wl[92] vdd gnd cell_6t
Xbit_r93_c184 bl[184] br[184] wl[93] vdd gnd cell_6t
Xbit_r94_c184 bl[184] br[184] wl[94] vdd gnd cell_6t
Xbit_r95_c184 bl[184] br[184] wl[95] vdd gnd cell_6t
Xbit_r96_c184 bl[184] br[184] wl[96] vdd gnd cell_6t
Xbit_r97_c184 bl[184] br[184] wl[97] vdd gnd cell_6t
Xbit_r98_c184 bl[184] br[184] wl[98] vdd gnd cell_6t
Xbit_r99_c184 bl[184] br[184] wl[99] vdd gnd cell_6t
Xbit_r100_c184 bl[184] br[184] wl[100] vdd gnd cell_6t
Xbit_r101_c184 bl[184] br[184] wl[101] vdd gnd cell_6t
Xbit_r102_c184 bl[184] br[184] wl[102] vdd gnd cell_6t
Xbit_r103_c184 bl[184] br[184] wl[103] vdd gnd cell_6t
Xbit_r104_c184 bl[184] br[184] wl[104] vdd gnd cell_6t
Xbit_r105_c184 bl[184] br[184] wl[105] vdd gnd cell_6t
Xbit_r106_c184 bl[184] br[184] wl[106] vdd gnd cell_6t
Xbit_r107_c184 bl[184] br[184] wl[107] vdd gnd cell_6t
Xbit_r108_c184 bl[184] br[184] wl[108] vdd gnd cell_6t
Xbit_r109_c184 bl[184] br[184] wl[109] vdd gnd cell_6t
Xbit_r110_c184 bl[184] br[184] wl[110] vdd gnd cell_6t
Xbit_r111_c184 bl[184] br[184] wl[111] vdd gnd cell_6t
Xbit_r112_c184 bl[184] br[184] wl[112] vdd gnd cell_6t
Xbit_r113_c184 bl[184] br[184] wl[113] vdd gnd cell_6t
Xbit_r114_c184 bl[184] br[184] wl[114] vdd gnd cell_6t
Xbit_r115_c184 bl[184] br[184] wl[115] vdd gnd cell_6t
Xbit_r116_c184 bl[184] br[184] wl[116] vdd gnd cell_6t
Xbit_r117_c184 bl[184] br[184] wl[117] vdd gnd cell_6t
Xbit_r118_c184 bl[184] br[184] wl[118] vdd gnd cell_6t
Xbit_r119_c184 bl[184] br[184] wl[119] vdd gnd cell_6t
Xbit_r120_c184 bl[184] br[184] wl[120] vdd gnd cell_6t
Xbit_r121_c184 bl[184] br[184] wl[121] vdd gnd cell_6t
Xbit_r122_c184 bl[184] br[184] wl[122] vdd gnd cell_6t
Xbit_r123_c184 bl[184] br[184] wl[123] vdd gnd cell_6t
Xbit_r124_c184 bl[184] br[184] wl[124] vdd gnd cell_6t
Xbit_r125_c184 bl[184] br[184] wl[125] vdd gnd cell_6t
Xbit_r126_c184 bl[184] br[184] wl[126] vdd gnd cell_6t
Xbit_r127_c184 bl[184] br[184] wl[127] vdd gnd cell_6t
Xbit_r128_c184 bl[184] br[184] wl[128] vdd gnd cell_6t
Xbit_r129_c184 bl[184] br[184] wl[129] vdd gnd cell_6t
Xbit_r130_c184 bl[184] br[184] wl[130] vdd gnd cell_6t
Xbit_r131_c184 bl[184] br[184] wl[131] vdd gnd cell_6t
Xbit_r132_c184 bl[184] br[184] wl[132] vdd gnd cell_6t
Xbit_r133_c184 bl[184] br[184] wl[133] vdd gnd cell_6t
Xbit_r134_c184 bl[184] br[184] wl[134] vdd gnd cell_6t
Xbit_r135_c184 bl[184] br[184] wl[135] vdd gnd cell_6t
Xbit_r136_c184 bl[184] br[184] wl[136] vdd gnd cell_6t
Xbit_r137_c184 bl[184] br[184] wl[137] vdd gnd cell_6t
Xbit_r138_c184 bl[184] br[184] wl[138] vdd gnd cell_6t
Xbit_r139_c184 bl[184] br[184] wl[139] vdd gnd cell_6t
Xbit_r140_c184 bl[184] br[184] wl[140] vdd gnd cell_6t
Xbit_r141_c184 bl[184] br[184] wl[141] vdd gnd cell_6t
Xbit_r142_c184 bl[184] br[184] wl[142] vdd gnd cell_6t
Xbit_r143_c184 bl[184] br[184] wl[143] vdd gnd cell_6t
Xbit_r144_c184 bl[184] br[184] wl[144] vdd gnd cell_6t
Xbit_r145_c184 bl[184] br[184] wl[145] vdd gnd cell_6t
Xbit_r146_c184 bl[184] br[184] wl[146] vdd gnd cell_6t
Xbit_r147_c184 bl[184] br[184] wl[147] vdd gnd cell_6t
Xbit_r148_c184 bl[184] br[184] wl[148] vdd gnd cell_6t
Xbit_r149_c184 bl[184] br[184] wl[149] vdd gnd cell_6t
Xbit_r150_c184 bl[184] br[184] wl[150] vdd gnd cell_6t
Xbit_r151_c184 bl[184] br[184] wl[151] vdd gnd cell_6t
Xbit_r152_c184 bl[184] br[184] wl[152] vdd gnd cell_6t
Xbit_r153_c184 bl[184] br[184] wl[153] vdd gnd cell_6t
Xbit_r154_c184 bl[184] br[184] wl[154] vdd gnd cell_6t
Xbit_r155_c184 bl[184] br[184] wl[155] vdd gnd cell_6t
Xbit_r156_c184 bl[184] br[184] wl[156] vdd gnd cell_6t
Xbit_r157_c184 bl[184] br[184] wl[157] vdd gnd cell_6t
Xbit_r158_c184 bl[184] br[184] wl[158] vdd gnd cell_6t
Xbit_r159_c184 bl[184] br[184] wl[159] vdd gnd cell_6t
Xbit_r160_c184 bl[184] br[184] wl[160] vdd gnd cell_6t
Xbit_r161_c184 bl[184] br[184] wl[161] vdd gnd cell_6t
Xbit_r162_c184 bl[184] br[184] wl[162] vdd gnd cell_6t
Xbit_r163_c184 bl[184] br[184] wl[163] vdd gnd cell_6t
Xbit_r164_c184 bl[184] br[184] wl[164] vdd gnd cell_6t
Xbit_r165_c184 bl[184] br[184] wl[165] vdd gnd cell_6t
Xbit_r166_c184 bl[184] br[184] wl[166] vdd gnd cell_6t
Xbit_r167_c184 bl[184] br[184] wl[167] vdd gnd cell_6t
Xbit_r168_c184 bl[184] br[184] wl[168] vdd gnd cell_6t
Xbit_r169_c184 bl[184] br[184] wl[169] vdd gnd cell_6t
Xbit_r170_c184 bl[184] br[184] wl[170] vdd gnd cell_6t
Xbit_r171_c184 bl[184] br[184] wl[171] vdd gnd cell_6t
Xbit_r172_c184 bl[184] br[184] wl[172] vdd gnd cell_6t
Xbit_r173_c184 bl[184] br[184] wl[173] vdd gnd cell_6t
Xbit_r174_c184 bl[184] br[184] wl[174] vdd gnd cell_6t
Xbit_r175_c184 bl[184] br[184] wl[175] vdd gnd cell_6t
Xbit_r176_c184 bl[184] br[184] wl[176] vdd gnd cell_6t
Xbit_r177_c184 bl[184] br[184] wl[177] vdd gnd cell_6t
Xbit_r178_c184 bl[184] br[184] wl[178] vdd gnd cell_6t
Xbit_r179_c184 bl[184] br[184] wl[179] vdd gnd cell_6t
Xbit_r180_c184 bl[184] br[184] wl[180] vdd gnd cell_6t
Xbit_r181_c184 bl[184] br[184] wl[181] vdd gnd cell_6t
Xbit_r182_c184 bl[184] br[184] wl[182] vdd gnd cell_6t
Xbit_r183_c184 bl[184] br[184] wl[183] vdd gnd cell_6t
Xbit_r184_c184 bl[184] br[184] wl[184] vdd gnd cell_6t
Xbit_r185_c184 bl[184] br[184] wl[185] vdd gnd cell_6t
Xbit_r186_c184 bl[184] br[184] wl[186] vdd gnd cell_6t
Xbit_r187_c184 bl[184] br[184] wl[187] vdd gnd cell_6t
Xbit_r188_c184 bl[184] br[184] wl[188] vdd gnd cell_6t
Xbit_r189_c184 bl[184] br[184] wl[189] vdd gnd cell_6t
Xbit_r190_c184 bl[184] br[184] wl[190] vdd gnd cell_6t
Xbit_r191_c184 bl[184] br[184] wl[191] vdd gnd cell_6t
Xbit_r192_c184 bl[184] br[184] wl[192] vdd gnd cell_6t
Xbit_r193_c184 bl[184] br[184] wl[193] vdd gnd cell_6t
Xbit_r194_c184 bl[184] br[184] wl[194] vdd gnd cell_6t
Xbit_r195_c184 bl[184] br[184] wl[195] vdd gnd cell_6t
Xbit_r196_c184 bl[184] br[184] wl[196] vdd gnd cell_6t
Xbit_r197_c184 bl[184] br[184] wl[197] vdd gnd cell_6t
Xbit_r198_c184 bl[184] br[184] wl[198] vdd gnd cell_6t
Xbit_r199_c184 bl[184] br[184] wl[199] vdd gnd cell_6t
Xbit_r200_c184 bl[184] br[184] wl[200] vdd gnd cell_6t
Xbit_r201_c184 bl[184] br[184] wl[201] vdd gnd cell_6t
Xbit_r202_c184 bl[184] br[184] wl[202] vdd gnd cell_6t
Xbit_r203_c184 bl[184] br[184] wl[203] vdd gnd cell_6t
Xbit_r204_c184 bl[184] br[184] wl[204] vdd gnd cell_6t
Xbit_r205_c184 bl[184] br[184] wl[205] vdd gnd cell_6t
Xbit_r206_c184 bl[184] br[184] wl[206] vdd gnd cell_6t
Xbit_r207_c184 bl[184] br[184] wl[207] vdd gnd cell_6t
Xbit_r208_c184 bl[184] br[184] wl[208] vdd gnd cell_6t
Xbit_r209_c184 bl[184] br[184] wl[209] vdd gnd cell_6t
Xbit_r210_c184 bl[184] br[184] wl[210] vdd gnd cell_6t
Xbit_r211_c184 bl[184] br[184] wl[211] vdd gnd cell_6t
Xbit_r212_c184 bl[184] br[184] wl[212] vdd gnd cell_6t
Xbit_r213_c184 bl[184] br[184] wl[213] vdd gnd cell_6t
Xbit_r214_c184 bl[184] br[184] wl[214] vdd gnd cell_6t
Xbit_r215_c184 bl[184] br[184] wl[215] vdd gnd cell_6t
Xbit_r216_c184 bl[184] br[184] wl[216] vdd gnd cell_6t
Xbit_r217_c184 bl[184] br[184] wl[217] vdd gnd cell_6t
Xbit_r218_c184 bl[184] br[184] wl[218] vdd gnd cell_6t
Xbit_r219_c184 bl[184] br[184] wl[219] vdd gnd cell_6t
Xbit_r220_c184 bl[184] br[184] wl[220] vdd gnd cell_6t
Xbit_r221_c184 bl[184] br[184] wl[221] vdd gnd cell_6t
Xbit_r222_c184 bl[184] br[184] wl[222] vdd gnd cell_6t
Xbit_r223_c184 bl[184] br[184] wl[223] vdd gnd cell_6t
Xbit_r224_c184 bl[184] br[184] wl[224] vdd gnd cell_6t
Xbit_r225_c184 bl[184] br[184] wl[225] vdd gnd cell_6t
Xbit_r226_c184 bl[184] br[184] wl[226] vdd gnd cell_6t
Xbit_r227_c184 bl[184] br[184] wl[227] vdd gnd cell_6t
Xbit_r228_c184 bl[184] br[184] wl[228] vdd gnd cell_6t
Xbit_r229_c184 bl[184] br[184] wl[229] vdd gnd cell_6t
Xbit_r230_c184 bl[184] br[184] wl[230] vdd gnd cell_6t
Xbit_r231_c184 bl[184] br[184] wl[231] vdd gnd cell_6t
Xbit_r232_c184 bl[184] br[184] wl[232] vdd gnd cell_6t
Xbit_r233_c184 bl[184] br[184] wl[233] vdd gnd cell_6t
Xbit_r234_c184 bl[184] br[184] wl[234] vdd gnd cell_6t
Xbit_r235_c184 bl[184] br[184] wl[235] vdd gnd cell_6t
Xbit_r236_c184 bl[184] br[184] wl[236] vdd gnd cell_6t
Xbit_r237_c184 bl[184] br[184] wl[237] vdd gnd cell_6t
Xbit_r238_c184 bl[184] br[184] wl[238] vdd gnd cell_6t
Xbit_r239_c184 bl[184] br[184] wl[239] vdd gnd cell_6t
Xbit_r240_c184 bl[184] br[184] wl[240] vdd gnd cell_6t
Xbit_r241_c184 bl[184] br[184] wl[241] vdd gnd cell_6t
Xbit_r242_c184 bl[184] br[184] wl[242] vdd gnd cell_6t
Xbit_r243_c184 bl[184] br[184] wl[243] vdd gnd cell_6t
Xbit_r244_c184 bl[184] br[184] wl[244] vdd gnd cell_6t
Xbit_r245_c184 bl[184] br[184] wl[245] vdd gnd cell_6t
Xbit_r246_c184 bl[184] br[184] wl[246] vdd gnd cell_6t
Xbit_r247_c184 bl[184] br[184] wl[247] vdd gnd cell_6t
Xbit_r248_c184 bl[184] br[184] wl[248] vdd gnd cell_6t
Xbit_r249_c184 bl[184] br[184] wl[249] vdd gnd cell_6t
Xbit_r250_c184 bl[184] br[184] wl[250] vdd gnd cell_6t
Xbit_r251_c184 bl[184] br[184] wl[251] vdd gnd cell_6t
Xbit_r252_c184 bl[184] br[184] wl[252] vdd gnd cell_6t
Xbit_r253_c184 bl[184] br[184] wl[253] vdd gnd cell_6t
Xbit_r254_c184 bl[184] br[184] wl[254] vdd gnd cell_6t
Xbit_r255_c184 bl[184] br[184] wl[255] vdd gnd cell_6t
Xbit_r0_c185 bl[185] br[185] wl[0] vdd gnd cell_6t
Xbit_r1_c185 bl[185] br[185] wl[1] vdd gnd cell_6t
Xbit_r2_c185 bl[185] br[185] wl[2] vdd gnd cell_6t
Xbit_r3_c185 bl[185] br[185] wl[3] vdd gnd cell_6t
Xbit_r4_c185 bl[185] br[185] wl[4] vdd gnd cell_6t
Xbit_r5_c185 bl[185] br[185] wl[5] vdd gnd cell_6t
Xbit_r6_c185 bl[185] br[185] wl[6] vdd gnd cell_6t
Xbit_r7_c185 bl[185] br[185] wl[7] vdd gnd cell_6t
Xbit_r8_c185 bl[185] br[185] wl[8] vdd gnd cell_6t
Xbit_r9_c185 bl[185] br[185] wl[9] vdd gnd cell_6t
Xbit_r10_c185 bl[185] br[185] wl[10] vdd gnd cell_6t
Xbit_r11_c185 bl[185] br[185] wl[11] vdd gnd cell_6t
Xbit_r12_c185 bl[185] br[185] wl[12] vdd gnd cell_6t
Xbit_r13_c185 bl[185] br[185] wl[13] vdd gnd cell_6t
Xbit_r14_c185 bl[185] br[185] wl[14] vdd gnd cell_6t
Xbit_r15_c185 bl[185] br[185] wl[15] vdd gnd cell_6t
Xbit_r16_c185 bl[185] br[185] wl[16] vdd gnd cell_6t
Xbit_r17_c185 bl[185] br[185] wl[17] vdd gnd cell_6t
Xbit_r18_c185 bl[185] br[185] wl[18] vdd gnd cell_6t
Xbit_r19_c185 bl[185] br[185] wl[19] vdd gnd cell_6t
Xbit_r20_c185 bl[185] br[185] wl[20] vdd gnd cell_6t
Xbit_r21_c185 bl[185] br[185] wl[21] vdd gnd cell_6t
Xbit_r22_c185 bl[185] br[185] wl[22] vdd gnd cell_6t
Xbit_r23_c185 bl[185] br[185] wl[23] vdd gnd cell_6t
Xbit_r24_c185 bl[185] br[185] wl[24] vdd gnd cell_6t
Xbit_r25_c185 bl[185] br[185] wl[25] vdd gnd cell_6t
Xbit_r26_c185 bl[185] br[185] wl[26] vdd gnd cell_6t
Xbit_r27_c185 bl[185] br[185] wl[27] vdd gnd cell_6t
Xbit_r28_c185 bl[185] br[185] wl[28] vdd gnd cell_6t
Xbit_r29_c185 bl[185] br[185] wl[29] vdd gnd cell_6t
Xbit_r30_c185 bl[185] br[185] wl[30] vdd gnd cell_6t
Xbit_r31_c185 bl[185] br[185] wl[31] vdd gnd cell_6t
Xbit_r32_c185 bl[185] br[185] wl[32] vdd gnd cell_6t
Xbit_r33_c185 bl[185] br[185] wl[33] vdd gnd cell_6t
Xbit_r34_c185 bl[185] br[185] wl[34] vdd gnd cell_6t
Xbit_r35_c185 bl[185] br[185] wl[35] vdd gnd cell_6t
Xbit_r36_c185 bl[185] br[185] wl[36] vdd gnd cell_6t
Xbit_r37_c185 bl[185] br[185] wl[37] vdd gnd cell_6t
Xbit_r38_c185 bl[185] br[185] wl[38] vdd gnd cell_6t
Xbit_r39_c185 bl[185] br[185] wl[39] vdd gnd cell_6t
Xbit_r40_c185 bl[185] br[185] wl[40] vdd gnd cell_6t
Xbit_r41_c185 bl[185] br[185] wl[41] vdd gnd cell_6t
Xbit_r42_c185 bl[185] br[185] wl[42] vdd gnd cell_6t
Xbit_r43_c185 bl[185] br[185] wl[43] vdd gnd cell_6t
Xbit_r44_c185 bl[185] br[185] wl[44] vdd gnd cell_6t
Xbit_r45_c185 bl[185] br[185] wl[45] vdd gnd cell_6t
Xbit_r46_c185 bl[185] br[185] wl[46] vdd gnd cell_6t
Xbit_r47_c185 bl[185] br[185] wl[47] vdd gnd cell_6t
Xbit_r48_c185 bl[185] br[185] wl[48] vdd gnd cell_6t
Xbit_r49_c185 bl[185] br[185] wl[49] vdd gnd cell_6t
Xbit_r50_c185 bl[185] br[185] wl[50] vdd gnd cell_6t
Xbit_r51_c185 bl[185] br[185] wl[51] vdd gnd cell_6t
Xbit_r52_c185 bl[185] br[185] wl[52] vdd gnd cell_6t
Xbit_r53_c185 bl[185] br[185] wl[53] vdd gnd cell_6t
Xbit_r54_c185 bl[185] br[185] wl[54] vdd gnd cell_6t
Xbit_r55_c185 bl[185] br[185] wl[55] vdd gnd cell_6t
Xbit_r56_c185 bl[185] br[185] wl[56] vdd gnd cell_6t
Xbit_r57_c185 bl[185] br[185] wl[57] vdd gnd cell_6t
Xbit_r58_c185 bl[185] br[185] wl[58] vdd gnd cell_6t
Xbit_r59_c185 bl[185] br[185] wl[59] vdd gnd cell_6t
Xbit_r60_c185 bl[185] br[185] wl[60] vdd gnd cell_6t
Xbit_r61_c185 bl[185] br[185] wl[61] vdd gnd cell_6t
Xbit_r62_c185 bl[185] br[185] wl[62] vdd gnd cell_6t
Xbit_r63_c185 bl[185] br[185] wl[63] vdd gnd cell_6t
Xbit_r64_c185 bl[185] br[185] wl[64] vdd gnd cell_6t
Xbit_r65_c185 bl[185] br[185] wl[65] vdd gnd cell_6t
Xbit_r66_c185 bl[185] br[185] wl[66] vdd gnd cell_6t
Xbit_r67_c185 bl[185] br[185] wl[67] vdd gnd cell_6t
Xbit_r68_c185 bl[185] br[185] wl[68] vdd gnd cell_6t
Xbit_r69_c185 bl[185] br[185] wl[69] vdd gnd cell_6t
Xbit_r70_c185 bl[185] br[185] wl[70] vdd gnd cell_6t
Xbit_r71_c185 bl[185] br[185] wl[71] vdd gnd cell_6t
Xbit_r72_c185 bl[185] br[185] wl[72] vdd gnd cell_6t
Xbit_r73_c185 bl[185] br[185] wl[73] vdd gnd cell_6t
Xbit_r74_c185 bl[185] br[185] wl[74] vdd gnd cell_6t
Xbit_r75_c185 bl[185] br[185] wl[75] vdd gnd cell_6t
Xbit_r76_c185 bl[185] br[185] wl[76] vdd gnd cell_6t
Xbit_r77_c185 bl[185] br[185] wl[77] vdd gnd cell_6t
Xbit_r78_c185 bl[185] br[185] wl[78] vdd gnd cell_6t
Xbit_r79_c185 bl[185] br[185] wl[79] vdd gnd cell_6t
Xbit_r80_c185 bl[185] br[185] wl[80] vdd gnd cell_6t
Xbit_r81_c185 bl[185] br[185] wl[81] vdd gnd cell_6t
Xbit_r82_c185 bl[185] br[185] wl[82] vdd gnd cell_6t
Xbit_r83_c185 bl[185] br[185] wl[83] vdd gnd cell_6t
Xbit_r84_c185 bl[185] br[185] wl[84] vdd gnd cell_6t
Xbit_r85_c185 bl[185] br[185] wl[85] vdd gnd cell_6t
Xbit_r86_c185 bl[185] br[185] wl[86] vdd gnd cell_6t
Xbit_r87_c185 bl[185] br[185] wl[87] vdd gnd cell_6t
Xbit_r88_c185 bl[185] br[185] wl[88] vdd gnd cell_6t
Xbit_r89_c185 bl[185] br[185] wl[89] vdd gnd cell_6t
Xbit_r90_c185 bl[185] br[185] wl[90] vdd gnd cell_6t
Xbit_r91_c185 bl[185] br[185] wl[91] vdd gnd cell_6t
Xbit_r92_c185 bl[185] br[185] wl[92] vdd gnd cell_6t
Xbit_r93_c185 bl[185] br[185] wl[93] vdd gnd cell_6t
Xbit_r94_c185 bl[185] br[185] wl[94] vdd gnd cell_6t
Xbit_r95_c185 bl[185] br[185] wl[95] vdd gnd cell_6t
Xbit_r96_c185 bl[185] br[185] wl[96] vdd gnd cell_6t
Xbit_r97_c185 bl[185] br[185] wl[97] vdd gnd cell_6t
Xbit_r98_c185 bl[185] br[185] wl[98] vdd gnd cell_6t
Xbit_r99_c185 bl[185] br[185] wl[99] vdd gnd cell_6t
Xbit_r100_c185 bl[185] br[185] wl[100] vdd gnd cell_6t
Xbit_r101_c185 bl[185] br[185] wl[101] vdd gnd cell_6t
Xbit_r102_c185 bl[185] br[185] wl[102] vdd gnd cell_6t
Xbit_r103_c185 bl[185] br[185] wl[103] vdd gnd cell_6t
Xbit_r104_c185 bl[185] br[185] wl[104] vdd gnd cell_6t
Xbit_r105_c185 bl[185] br[185] wl[105] vdd gnd cell_6t
Xbit_r106_c185 bl[185] br[185] wl[106] vdd gnd cell_6t
Xbit_r107_c185 bl[185] br[185] wl[107] vdd gnd cell_6t
Xbit_r108_c185 bl[185] br[185] wl[108] vdd gnd cell_6t
Xbit_r109_c185 bl[185] br[185] wl[109] vdd gnd cell_6t
Xbit_r110_c185 bl[185] br[185] wl[110] vdd gnd cell_6t
Xbit_r111_c185 bl[185] br[185] wl[111] vdd gnd cell_6t
Xbit_r112_c185 bl[185] br[185] wl[112] vdd gnd cell_6t
Xbit_r113_c185 bl[185] br[185] wl[113] vdd gnd cell_6t
Xbit_r114_c185 bl[185] br[185] wl[114] vdd gnd cell_6t
Xbit_r115_c185 bl[185] br[185] wl[115] vdd gnd cell_6t
Xbit_r116_c185 bl[185] br[185] wl[116] vdd gnd cell_6t
Xbit_r117_c185 bl[185] br[185] wl[117] vdd gnd cell_6t
Xbit_r118_c185 bl[185] br[185] wl[118] vdd gnd cell_6t
Xbit_r119_c185 bl[185] br[185] wl[119] vdd gnd cell_6t
Xbit_r120_c185 bl[185] br[185] wl[120] vdd gnd cell_6t
Xbit_r121_c185 bl[185] br[185] wl[121] vdd gnd cell_6t
Xbit_r122_c185 bl[185] br[185] wl[122] vdd gnd cell_6t
Xbit_r123_c185 bl[185] br[185] wl[123] vdd gnd cell_6t
Xbit_r124_c185 bl[185] br[185] wl[124] vdd gnd cell_6t
Xbit_r125_c185 bl[185] br[185] wl[125] vdd gnd cell_6t
Xbit_r126_c185 bl[185] br[185] wl[126] vdd gnd cell_6t
Xbit_r127_c185 bl[185] br[185] wl[127] vdd gnd cell_6t
Xbit_r128_c185 bl[185] br[185] wl[128] vdd gnd cell_6t
Xbit_r129_c185 bl[185] br[185] wl[129] vdd gnd cell_6t
Xbit_r130_c185 bl[185] br[185] wl[130] vdd gnd cell_6t
Xbit_r131_c185 bl[185] br[185] wl[131] vdd gnd cell_6t
Xbit_r132_c185 bl[185] br[185] wl[132] vdd gnd cell_6t
Xbit_r133_c185 bl[185] br[185] wl[133] vdd gnd cell_6t
Xbit_r134_c185 bl[185] br[185] wl[134] vdd gnd cell_6t
Xbit_r135_c185 bl[185] br[185] wl[135] vdd gnd cell_6t
Xbit_r136_c185 bl[185] br[185] wl[136] vdd gnd cell_6t
Xbit_r137_c185 bl[185] br[185] wl[137] vdd gnd cell_6t
Xbit_r138_c185 bl[185] br[185] wl[138] vdd gnd cell_6t
Xbit_r139_c185 bl[185] br[185] wl[139] vdd gnd cell_6t
Xbit_r140_c185 bl[185] br[185] wl[140] vdd gnd cell_6t
Xbit_r141_c185 bl[185] br[185] wl[141] vdd gnd cell_6t
Xbit_r142_c185 bl[185] br[185] wl[142] vdd gnd cell_6t
Xbit_r143_c185 bl[185] br[185] wl[143] vdd gnd cell_6t
Xbit_r144_c185 bl[185] br[185] wl[144] vdd gnd cell_6t
Xbit_r145_c185 bl[185] br[185] wl[145] vdd gnd cell_6t
Xbit_r146_c185 bl[185] br[185] wl[146] vdd gnd cell_6t
Xbit_r147_c185 bl[185] br[185] wl[147] vdd gnd cell_6t
Xbit_r148_c185 bl[185] br[185] wl[148] vdd gnd cell_6t
Xbit_r149_c185 bl[185] br[185] wl[149] vdd gnd cell_6t
Xbit_r150_c185 bl[185] br[185] wl[150] vdd gnd cell_6t
Xbit_r151_c185 bl[185] br[185] wl[151] vdd gnd cell_6t
Xbit_r152_c185 bl[185] br[185] wl[152] vdd gnd cell_6t
Xbit_r153_c185 bl[185] br[185] wl[153] vdd gnd cell_6t
Xbit_r154_c185 bl[185] br[185] wl[154] vdd gnd cell_6t
Xbit_r155_c185 bl[185] br[185] wl[155] vdd gnd cell_6t
Xbit_r156_c185 bl[185] br[185] wl[156] vdd gnd cell_6t
Xbit_r157_c185 bl[185] br[185] wl[157] vdd gnd cell_6t
Xbit_r158_c185 bl[185] br[185] wl[158] vdd gnd cell_6t
Xbit_r159_c185 bl[185] br[185] wl[159] vdd gnd cell_6t
Xbit_r160_c185 bl[185] br[185] wl[160] vdd gnd cell_6t
Xbit_r161_c185 bl[185] br[185] wl[161] vdd gnd cell_6t
Xbit_r162_c185 bl[185] br[185] wl[162] vdd gnd cell_6t
Xbit_r163_c185 bl[185] br[185] wl[163] vdd gnd cell_6t
Xbit_r164_c185 bl[185] br[185] wl[164] vdd gnd cell_6t
Xbit_r165_c185 bl[185] br[185] wl[165] vdd gnd cell_6t
Xbit_r166_c185 bl[185] br[185] wl[166] vdd gnd cell_6t
Xbit_r167_c185 bl[185] br[185] wl[167] vdd gnd cell_6t
Xbit_r168_c185 bl[185] br[185] wl[168] vdd gnd cell_6t
Xbit_r169_c185 bl[185] br[185] wl[169] vdd gnd cell_6t
Xbit_r170_c185 bl[185] br[185] wl[170] vdd gnd cell_6t
Xbit_r171_c185 bl[185] br[185] wl[171] vdd gnd cell_6t
Xbit_r172_c185 bl[185] br[185] wl[172] vdd gnd cell_6t
Xbit_r173_c185 bl[185] br[185] wl[173] vdd gnd cell_6t
Xbit_r174_c185 bl[185] br[185] wl[174] vdd gnd cell_6t
Xbit_r175_c185 bl[185] br[185] wl[175] vdd gnd cell_6t
Xbit_r176_c185 bl[185] br[185] wl[176] vdd gnd cell_6t
Xbit_r177_c185 bl[185] br[185] wl[177] vdd gnd cell_6t
Xbit_r178_c185 bl[185] br[185] wl[178] vdd gnd cell_6t
Xbit_r179_c185 bl[185] br[185] wl[179] vdd gnd cell_6t
Xbit_r180_c185 bl[185] br[185] wl[180] vdd gnd cell_6t
Xbit_r181_c185 bl[185] br[185] wl[181] vdd gnd cell_6t
Xbit_r182_c185 bl[185] br[185] wl[182] vdd gnd cell_6t
Xbit_r183_c185 bl[185] br[185] wl[183] vdd gnd cell_6t
Xbit_r184_c185 bl[185] br[185] wl[184] vdd gnd cell_6t
Xbit_r185_c185 bl[185] br[185] wl[185] vdd gnd cell_6t
Xbit_r186_c185 bl[185] br[185] wl[186] vdd gnd cell_6t
Xbit_r187_c185 bl[185] br[185] wl[187] vdd gnd cell_6t
Xbit_r188_c185 bl[185] br[185] wl[188] vdd gnd cell_6t
Xbit_r189_c185 bl[185] br[185] wl[189] vdd gnd cell_6t
Xbit_r190_c185 bl[185] br[185] wl[190] vdd gnd cell_6t
Xbit_r191_c185 bl[185] br[185] wl[191] vdd gnd cell_6t
Xbit_r192_c185 bl[185] br[185] wl[192] vdd gnd cell_6t
Xbit_r193_c185 bl[185] br[185] wl[193] vdd gnd cell_6t
Xbit_r194_c185 bl[185] br[185] wl[194] vdd gnd cell_6t
Xbit_r195_c185 bl[185] br[185] wl[195] vdd gnd cell_6t
Xbit_r196_c185 bl[185] br[185] wl[196] vdd gnd cell_6t
Xbit_r197_c185 bl[185] br[185] wl[197] vdd gnd cell_6t
Xbit_r198_c185 bl[185] br[185] wl[198] vdd gnd cell_6t
Xbit_r199_c185 bl[185] br[185] wl[199] vdd gnd cell_6t
Xbit_r200_c185 bl[185] br[185] wl[200] vdd gnd cell_6t
Xbit_r201_c185 bl[185] br[185] wl[201] vdd gnd cell_6t
Xbit_r202_c185 bl[185] br[185] wl[202] vdd gnd cell_6t
Xbit_r203_c185 bl[185] br[185] wl[203] vdd gnd cell_6t
Xbit_r204_c185 bl[185] br[185] wl[204] vdd gnd cell_6t
Xbit_r205_c185 bl[185] br[185] wl[205] vdd gnd cell_6t
Xbit_r206_c185 bl[185] br[185] wl[206] vdd gnd cell_6t
Xbit_r207_c185 bl[185] br[185] wl[207] vdd gnd cell_6t
Xbit_r208_c185 bl[185] br[185] wl[208] vdd gnd cell_6t
Xbit_r209_c185 bl[185] br[185] wl[209] vdd gnd cell_6t
Xbit_r210_c185 bl[185] br[185] wl[210] vdd gnd cell_6t
Xbit_r211_c185 bl[185] br[185] wl[211] vdd gnd cell_6t
Xbit_r212_c185 bl[185] br[185] wl[212] vdd gnd cell_6t
Xbit_r213_c185 bl[185] br[185] wl[213] vdd gnd cell_6t
Xbit_r214_c185 bl[185] br[185] wl[214] vdd gnd cell_6t
Xbit_r215_c185 bl[185] br[185] wl[215] vdd gnd cell_6t
Xbit_r216_c185 bl[185] br[185] wl[216] vdd gnd cell_6t
Xbit_r217_c185 bl[185] br[185] wl[217] vdd gnd cell_6t
Xbit_r218_c185 bl[185] br[185] wl[218] vdd gnd cell_6t
Xbit_r219_c185 bl[185] br[185] wl[219] vdd gnd cell_6t
Xbit_r220_c185 bl[185] br[185] wl[220] vdd gnd cell_6t
Xbit_r221_c185 bl[185] br[185] wl[221] vdd gnd cell_6t
Xbit_r222_c185 bl[185] br[185] wl[222] vdd gnd cell_6t
Xbit_r223_c185 bl[185] br[185] wl[223] vdd gnd cell_6t
Xbit_r224_c185 bl[185] br[185] wl[224] vdd gnd cell_6t
Xbit_r225_c185 bl[185] br[185] wl[225] vdd gnd cell_6t
Xbit_r226_c185 bl[185] br[185] wl[226] vdd gnd cell_6t
Xbit_r227_c185 bl[185] br[185] wl[227] vdd gnd cell_6t
Xbit_r228_c185 bl[185] br[185] wl[228] vdd gnd cell_6t
Xbit_r229_c185 bl[185] br[185] wl[229] vdd gnd cell_6t
Xbit_r230_c185 bl[185] br[185] wl[230] vdd gnd cell_6t
Xbit_r231_c185 bl[185] br[185] wl[231] vdd gnd cell_6t
Xbit_r232_c185 bl[185] br[185] wl[232] vdd gnd cell_6t
Xbit_r233_c185 bl[185] br[185] wl[233] vdd gnd cell_6t
Xbit_r234_c185 bl[185] br[185] wl[234] vdd gnd cell_6t
Xbit_r235_c185 bl[185] br[185] wl[235] vdd gnd cell_6t
Xbit_r236_c185 bl[185] br[185] wl[236] vdd gnd cell_6t
Xbit_r237_c185 bl[185] br[185] wl[237] vdd gnd cell_6t
Xbit_r238_c185 bl[185] br[185] wl[238] vdd gnd cell_6t
Xbit_r239_c185 bl[185] br[185] wl[239] vdd gnd cell_6t
Xbit_r240_c185 bl[185] br[185] wl[240] vdd gnd cell_6t
Xbit_r241_c185 bl[185] br[185] wl[241] vdd gnd cell_6t
Xbit_r242_c185 bl[185] br[185] wl[242] vdd gnd cell_6t
Xbit_r243_c185 bl[185] br[185] wl[243] vdd gnd cell_6t
Xbit_r244_c185 bl[185] br[185] wl[244] vdd gnd cell_6t
Xbit_r245_c185 bl[185] br[185] wl[245] vdd gnd cell_6t
Xbit_r246_c185 bl[185] br[185] wl[246] vdd gnd cell_6t
Xbit_r247_c185 bl[185] br[185] wl[247] vdd gnd cell_6t
Xbit_r248_c185 bl[185] br[185] wl[248] vdd gnd cell_6t
Xbit_r249_c185 bl[185] br[185] wl[249] vdd gnd cell_6t
Xbit_r250_c185 bl[185] br[185] wl[250] vdd gnd cell_6t
Xbit_r251_c185 bl[185] br[185] wl[251] vdd gnd cell_6t
Xbit_r252_c185 bl[185] br[185] wl[252] vdd gnd cell_6t
Xbit_r253_c185 bl[185] br[185] wl[253] vdd gnd cell_6t
Xbit_r254_c185 bl[185] br[185] wl[254] vdd gnd cell_6t
Xbit_r255_c185 bl[185] br[185] wl[255] vdd gnd cell_6t
Xbit_r0_c186 bl[186] br[186] wl[0] vdd gnd cell_6t
Xbit_r1_c186 bl[186] br[186] wl[1] vdd gnd cell_6t
Xbit_r2_c186 bl[186] br[186] wl[2] vdd gnd cell_6t
Xbit_r3_c186 bl[186] br[186] wl[3] vdd gnd cell_6t
Xbit_r4_c186 bl[186] br[186] wl[4] vdd gnd cell_6t
Xbit_r5_c186 bl[186] br[186] wl[5] vdd gnd cell_6t
Xbit_r6_c186 bl[186] br[186] wl[6] vdd gnd cell_6t
Xbit_r7_c186 bl[186] br[186] wl[7] vdd gnd cell_6t
Xbit_r8_c186 bl[186] br[186] wl[8] vdd gnd cell_6t
Xbit_r9_c186 bl[186] br[186] wl[9] vdd gnd cell_6t
Xbit_r10_c186 bl[186] br[186] wl[10] vdd gnd cell_6t
Xbit_r11_c186 bl[186] br[186] wl[11] vdd gnd cell_6t
Xbit_r12_c186 bl[186] br[186] wl[12] vdd gnd cell_6t
Xbit_r13_c186 bl[186] br[186] wl[13] vdd gnd cell_6t
Xbit_r14_c186 bl[186] br[186] wl[14] vdd gnd cell_6t
Xbit_r15_c186 bl[186] br[186] wl[15] vdd gnd cell_6t
Xbit_r16_c186 bl[186] br[186] wl[16] vdd gnd cell_6t
Xbit_r17_c186 bl[186] br[186] wl[17] vdd gnd cell_6t
Xbit_r18_c186 bl[186] br[186] wl[18] vdd gnd cell_6t
Xbit_r19_c186 bl[186] br[186] wl[19] vdd gnd cell_6t
Xbit_r20_c186 bl[186] br[186] wl[20] vdd gnd cell_6t
Xbit_r21_c186 bl[186] br[186] wl[21] vdd gnd cell_6t
Xbit_r22_c186 bl[186] br[186] wl[22] vdd gnd cell_6t
Xbit_r23_c186 bl[186] br[186] wl[23] vdd gnd cell_6t
Xbit_r24_c186 bl[186] br[186] wl[24] vdd gnd cell_6t
Xbit_r25_c186 bl[186] br[186] wl[25] vdd gnd cell_6t
Xbit_r26_c186 bl[186] br[186] wl[26] vdd gnd cell_6t
Xbit_r27_c186 bl[186] br[186] wl[27] vdd gnd cell_6t
Xbit_r28_c186 bl[186] br[186] wl[28] vdd gnd cell_6t
Xbit_r29_c186 bl[186] br[186] wl[29] vdd gnd cell_6t
Xbit_r30_c186 bl[186] br[186] wl[30] vdd gnd cell_6t
Xbit_r31_c186 bl[186] br[186] wl[31] vdd gnd cell_6t
Xbit_r32_c186 bl[186] br[186] wl[32] vdd gnd cell_6t
Xbit_r33_c186 bl[186] br[186] wl[33] vdd gnd cell_6t
Xbit_r34_c186 bl[186] br[186] wl[34] vdd gnd cell_6t
Xbit_r35_c186 bl[186] br[186] wl[35] vdd gnd cell_6t
Xbit_r36_c186 bl[186] br[186] wl[36] vdd gnd cell_6t
Xbit_r37_c186 bl[186] br[186] wl[37] vdd gnd cell_6t
Xbit_r38_c186 bl[186] br[186] wl[38] vdd gnd cell_6t
Xbit_r39_c186 bl[186] br[186] wl[39] vdd gnd cell_6t
Xbit_r40_c186 bl[186] br[186] wl[40] vdd gnd cell_6t
Xbit_r41_c186 bl[186] br[186] wl[41] vdd gnd cell_6t
Xbit_r42_c186 bl[186] br[186] wl[42] vdd gnd cell_6t
Xbit_r43_c186 bl[186] br[186] wl[43] vdd gnd cell_6t
Xbit_r44_c186 bl[186] br[186] wl[44] vdd gnd cell_6t
Xbit_r45_c186 bl[186] br[186] wl[45] vdd gnd cell_6t
Xbit_r46_c186 bl[186] br[186] wl[46] vdd gnd cell_6t
Xbit_r47_c186 bl[186] br[186] wl[47] vdd gnd cell_6t
Xbit_r48_c186 bl[186] br[186] wl[48] vdd gnd cell_6t
Xbit_r49_c186 bl[186] br[186] wl[49] vdd gnd cell_6t
Xbit_r50_c186 bl[186] br[186] wl[50] vdd gnd cell_6t
Xbit_r51_c186 bl[186] br[186] wl[51] vdd gnd cell_6t
Xbit_r52_c186 bl[186] br[186] wl[52] vdd gnd cell_6t
Xbit_r53_c186 bl[186] br[186] wl[53] vdd gnd cell_6t
Xbit_r54_c186 bl[186] br[186] wl[54] vdd gnd cell_6t
Xbit_r55_c186 bl[186] br[186] wl[55] vdd gnd cell_6t
Xbit_r56_c186 bl[186] br[186] wl[56] vdd gnd cell_6t
Xbit_r57_c186 bl[186] br[186] wl[57] vdd gnd cell_6t
Xbit_r58_c186 bl[186] br[186] wl[58] vdd gnd cell_6t
Xbit_r59_c186 bl[186] br[186] wl[59] vdd gnd cell_6t
Xbit_r60_c186 bl[186] br[186] wl[60] vdd gnd cell_6t
Xbit_r61_c186 bl[186] br[186] wl[61] vdd gnd cell_6t
Xbit_r62_c186 bl[186] br[186] wl[62] vdd gnd cell_6t
Xbit_r63_c186 bl[186] br[186] wl[63] vdd gnd cell_6t
Xbit_r64_c186 bl[186] br[186] wl[64] vdd gnd cell_6t
Xbit_r65_c186 bl[186] br[186] wl[65] vdd gnd cell_6t
Xbit_r66_c186 bl[186] br[186] wl[66] vdd gnd cell_6t
Xbit_r67_c186 bl[186] br[186] wl[67] vdd gnd cell_6t
Xbit_r68_c186 bl[186] br[186] wl[68] vdd gnd cell_6t
Xbit_r69_c186 bl[186] br[186] wl[69] vdd gnd cell_6t
Xbit_r70_c186 bl[186] br[186] wl[70] vdd gnd cell_6t
Xbit_r71_c186 bl[186] br[186] wl[71] vdd gnd cell_6t
Xbit_r72_c186 bl[186] br[186] wl[72] vdd gnd cell_6t
Xbit_r73_c186 bl[186] br[186] wl[73] vdd gnd cell_6t
Xbit_r74_c186 bl[186] br[186] wl[74] vdd gnd cell_6t
Xbit_r75_c186 bl[186] br[186] wl[75] vdd gnd cell_6t
Xbit_r76_c186 bl[186] br[186] wl[76] vdd gnd cell_6t
Xbit_r77_c186 bl[186] br[186] wl[77] vdd gnd cell_6t
Xbit_r78_c186 bl[186] br[186] wl[78] vdd gnd cell_6t
Xbit_r79_c186 bl[186] br[186] wl[79] vdd gnd cell_6t
Xbit_r80_c186 bl[186] br[186] wl[80] vdd gnd cell_6t
Xbit_r81_c186 bl[186] br[186] wl[81] vdd gnd cell_6t
Xbit_r82_c186 bl[186] br[186] wl[82] vdd gnd cell_6t
Xbit_r83_c186 bl[186] br[186] wl[83] vdd gnd cell_6t
Xbit_r84_c186 bl[186] br[186] wl[84] vdd gnd cell_6t
Xbit_r85_c186 bl[186] br[186] wl[85] vdd gnd cell_6t
Xbit_r86_c186 bl[186] br[186] wl[86] vdd gnd cell_6t
Xbit_r87_c186 bl[186] br[186] wl[87] vdd gnd cell_6t
Xbit_r88_c186 bl[186] br[186] wl[88] vdd gnd cell_6t
Xbit_r89_c186 bl[186] br[186] wl[89] vdd gnd cell_6t
Xbit_r90_c186 bl[186] br[186] wl[90] vdd gnd cell_6t
Xbit_r91_c186 bl[186] br[186] wl[91] vdd gnd cell_6t
Xbit_r92_c186 bl[186] br[186] wl[92] vdd gnd cell_6t
Xbit_r93_c186 bl[186] br[186] wl[93] vdd gnd cell_6t
Xbit_r94_c186 bl[186] br[186] wl[94] vdd gnd cell_6t
Xbit_r95_c186 bl[186] br[186] wl[95] vdd gnd cell_6t
Xbit_r96_c186 bl[186] br[186] wl[96] vdd gnd cell_6t
Xbit_r97_c186 bl[186] br[186] wl[97] vdd gnd cell_6t
Xbit_r98_c186 bl[186] br[186] wl[98] vdd gnd cell_6t
Xbit_r99_c186 bl[186] br[186] wl[99] vdd gnd cell_6t
Xbit_r100_c186 bl[186] br[186] wl[100] vdd gnd cell_6t
Xbit_r101_c186 bl[186] br[186] wl[101] vdd gnd cell_6t
Xbit_r102_c186 bl[186] br[186] wl[102] vdd gnd cell_6t
Xbit_r103_c186 bl[186] br[186] wl[103] vdd gnd cell_6t
Xbit_r104_c186 bl[186] br[186] wl[104] vdd gnd cell_6t
Xbit_r105_c186 bl[186] br[186] wl[105] vdd gnd cell_6t
Xbit_r106_c186 bl[186] br[186] wl[106] vdd gnd cell_6t
Xbit_r107_c186 bl[186] br[186] wl[107] vdd gnd cell_6t
Xbit_r108_c186 bl[186] br[186] wl[108] vdd gnd cell_6t
Xbit_r109_c186 bl[186] br[186] wl[109] vdd gnd cell_6t
Xbit_r110_c186 bl[186] br[186] wl[110] vdd gnd cell_6t
Xbit_r111_c186 bl[186] br[186] wl[111] vdd gnd cell_6t
Xbit_r112_c186 bl[186] br[186] wl[112] vdd gnd cell_6t
Xbit_r113_c186 bl[186] br[186] wl[113] vdd gnd cell_6t
Xbit_r114_c186 bl[186] br[186] wl[114] vdd gnd cell_6t
Xbit_r115_c186 bl[186] br[186] wl[115] vdd gnd cell_6t
Xbit_r116_c186 bl[186] br[186] wl[116] vdd gnd cell_6t
Xbit_r117_c186 bl[186] br[186] wl[117] vdd gnd cell_6t
Xbit_r118_c186 bl[186] br[186] wl[118] vdd gnd cell_6t
Xbit_r119_c186 bl[186] br[186] wl[119] vdd gnd cell_6t
Xbit_r120_c186 bl[186] br[186] wl[120] vdd gnd cell_6t
Xbit_r121_c186 bl[186] br[186] wl[121] vdd gnd cell_6t
Xbit_r122_c186 bl[186] br[186] wl[122] vdd gnd cell_6t
Xbit_r123_c186 bl[186] br[186] wl[123] vdd gnd cell_6t
Xbit_r124_c186 bl[186] br[186] wl[124] vdd gnd cell_6t
Xbit_r125_c186 bl[186] br[186] wl[125] vdd gnd cell_6t
Xbit_r126_c186 bl[186] br[186] wl[126] vdd gnd cell_6t
Xbit_r127_c186 bl[186] br[186] wl[127] vdd gnd cell_6t
Xbit_r128_c186 bl[186] br[186] wl[128] vdd gnd cell_6t
Xbit_r129_c186 bl[186] br[186] wl[129] vdd gnd cell_6t
Xbit_r130_c186 bl[186] br[186] wl[130] vdd gnd cell_6t
Xbit_r131_c186 bl[186] br[186] wl[131] vdd gnd cell_6t
Xbit_r132_c186 bl[186] br[186] wl[132] vdd gnd cell_6t
Xbit_r133_c186 bl[186] br[186] wl[133] vdd gnd cell_6t
Xbit_r134_c186 bl[186] br[186] wl[134] vdd gnd cell_6t
Xbit_r135_c186 bl[186] br[186] wl[135] vdd gnd cell_6t
Xbit_r136_c186 bl[186] br[186] wl[136] vdd gnd cell_6t
Xbit_r137_c186 bl[186] br[186] wl[137] vdd gnd cell_6t
Xbit_r138_c186 bl[186] br[186] wl[138] vdd gnd cell_6t
Xbit_r139_c186 bl[186] br[186] wl[139] vdd gnd cell_6t
Xbit_r140_c186 bl[186] br[186] wl[140] vdd gnd cell_6t
Xbit_r141_c186 bl[186] br[186] wl[141] vdd gnd cell_6t
Xbit_r142_c186 bl[186] br[186] wl[142] vdd gnd cell_6t
Xbit_r143_c186 bl[186] br[186] wl[143] vdd gnd cell_6t
Xbit_r144_c186 bl[186] br[186] wl[144] vdd gnd cell_6t
Xbit_r145_c186 bl[186] br[186] wl[145] vdd gnd cell_6t
Xbit_r146_c186 bl[186] br[186] wl[146] vdd gnd cell_6t
Xbit_r147_c186 bl[186] br[186] wl[147] vdd gnd cell_6t
Xbit_r148_c186 bl[186] br[186] wl[148] vdd gnd cell_6t
Xbit_r149_c186 bl[186] br[186] wl[149] vdd gnd cell_6t
Xbit_r150_c186 bl[186] br[186] wl[150] vdd gnd cell_6t
Xbit_r151_c186 bl[186] br[186] wl[151] vdd gnd cell_6t
Xbit_r152_c186 bl[186] br[186] wl[152] vdd gnd cell_6t
Xbit_r153_c186 bl[186] br[186] wl[153] vdd gnd cell_6t
Xbit_r154_c186 bl[186] br[186] wl[154] vdd gnd cell_6t
Xbit_r155_c186 bl[186] br[186] wl[155] vdd gnd cell_6t
Xbit_r156_c186 bl[186] br[186] wl[156] vdd gnd cell_6t
Xbit_r157_c186 bl[186] br[186] wl[157] vdd gnd cell_6t
Xbit_r158_c186 bl[186] br[186] wl[158] vdd gnd cell_6t
Xbit_r159_c186 bl[186] br[186] wl[159] vdd gnd cell_6t
Xbit_r160_c186 bl[186] br[186] wl[160] vdd gnd cell_6t
Xbit_r161_c186 bl[186] br[186] wl[161] vdd gnd cell_6t
Xbit_r162_c186 bl[186] br[186] wl[162] vdd gnd cell_6t
Xbit_r163_c186 bl[186] br[186] wl[163] vdd gnd cell_6t
Xbit_r164_c186 bl[186] br[186] wl[164] vdd gnd cell_6t
Xbit_r165_c186 bl[186] br[186] wl[165] vdd gnd cell_6t
Xbit_r166_c186 bl[186] br[186] wl[166] vdd gnd cell_6t
Xbit_r167_c186 bl[186] br[186] wl[167] vdd gnd cell_6t
Xbit_r168_c186 bl[186] br[186] wl[168] vdd gnd cell_6t
Xbit_r169_c186 bl[186] br[186] wl[169] vdd gnd cell_6t
Xbit_r170_c186 bl[186] br[186] wl[170] vdd gnd cell_6t
Xbit_r171_c186 bl[186] br[186] wl[171] vdd gnd cell_6t
Xbit_r172_c186 bl[186] br[186] wl[172] vdd gnd cell_6t
Xbit_r173_c186 bl[186] br[186] wl[173] vdd gnd cell_6t
Xbit_r174_c186 bl[186] br[186] wl[174] vdd gnd cell_6t
Xbit_r175_c186 bl[186] br[186] wl[175] vdd gnd cell_6t
Xbit_r176_c186 bl[186] br[186] wl[176] vdd gnd cell_6t
Xbit_r177_c186 bl[186] br[186] wl[177] vdd gnd cell_6t
Xbit_r178_c186 bl[186] br[186] wl[178] vdd gnd cell_6t
Xbit_r179_c186 bl[186] br[186] wl[179] vdd gnd cell_6t
Xbit_r180_c186 bl[186] br[186] wl[180] vdd gnd cell_6t
Xbit_r181_c186 bl[186] br[186] wl[181] vdd gnd cell_6t
Xbit_r182_c186 bl[186] br[186] wl[182] vdd gnd cell_6t
Xbit_r183_c186 bl[186] br[186] wl[183] vdd gnd cell_6t
Xbit_r184_c186 bl[186] br[186] wl[184] vdd gnd cell_6t
Xbit_r185_c186 bl[186] br[186] wl[185] vdd gnd cell_6t
Xbit_r186_c186 bl[186] br[186] wl[186] vdd gnd cell_6t
Xbit_r187_c186 bl[186] br[186] wl[187] vdd gnd cell_6t
Xbit_r188_c186 bl[186] br[186] wl[188] vdd gnd cell_6t
Xbit_r189_c186 bl[186] br[186] wl[189] vdd gnd cell_6t
Xbit_r190_c186 bl[186] br[186] wl[190] vdd gnd cell_6t
Xbit_r191_c186 bl[186] br[186] wl[191] vdd gnd cell_6t
Xbit_r192_c186 bl[186] br[186] wl[192] vdd gnd cell_6t
Xbit_r193_c186 bl[186] br[186] wl[193] vdd gnd cell_6t
Xbit_r194_c186 bl[186] br[186] wl[194] vdd gnd cell_6t
Xbit_r195_c186 bl[186] br[186] wl[195] vdd gnd cell_6t
Xbit_r196_c186 bl[186] br[186] wl[196] vdd gnd cell_6t
Xbit_r197_c186 bl[186] br[186] wl[197] vdd gnd cell_6t
Xbit_r198_c186 bl[186] br[186] wl[198] vdd gnd cell_6t
Xbit_r199_c186 bl[186] br[186] wl[199] vdd gnd cell_6t
Xbit_r200_c186 bl[186] br[186] wl[200] vdd gnd cell_6t
Xbit_r201_c186 bl[186] br[186] wl[201] vdd gnd cell_6t
Xbit_r202_c186 bl[186] br[186] wl[202] vdd gnd cell_6t
Xbit_r203_c186 bl[186] br[186] wl[203] vdd gnd cell_6t
Xbit_r204_c186 bl[186] br[186] wl[204] vdd gnd cell_6t
Xbit_r205_c186 bl[186] br[186] wl[205] vdd gnd cell_6t
Xbit_r206_c186 bl[186] br[186] wl[206] vdd gnd cell_6t
Xbit_r207_c186 bl[186] br[186] wl[207] vdd gnd cell_6t
Xbit_r208_c186 bl[186] br[186] wl[208] vdd gnd cell_6t
Xbit_r209_c186 bl[186] br[186] wl[209] vdd gnd cell_6t
Xbit_r210_c186 bl[186] br[186] wl[210] vdd gnd cell_6t
Xbit_r211_c186 bl[186] br[186] wl[211] vdd gnd cell_6t
Xbit_r212_c186 bl[186] br[186] wl[212] vdd gnd cell_6t
Xbit_r213_c186 bl[186] br[186] wl[213] vdd gnd cell_6t
Xbit_r214_c186 bl[186] br[186] wl[214] vdd gnd cell_6t
Xbit_r215_c186 bl[186] br[186] wl[215] vdd gnd cell_6t
Xbit_r216_c186 bl[186] br[186] wl[216] vdd gnd cell_6t
Xbit_r217_c186 bl[186] br[186] wl[217] vdd gnd cell_6t
Xbit_r218_c186 bl[186] br[186] wl[218] vdd gnd cell_6t
Xbit_r219_c186 bl[186] br[186] wl[219] vdd gnd cell_6t
Xbit_r220_c186 bl[186] br[186] wl[220] vdd gnd cell_6t
Xbit_r221_c186 bl[186] br[186] wl[221] vdd gnd cell_6t
Xbit_r222_c186 bl[186] br[186] wl[222] vdd gnd cell_6t
Xbit_r223_c186 bl[186] br[186] wl[223] vdd gnd cell_6t
Xbit_r224_c186 bl[186] br[186] wl[224] vdd gnd cell_6t
Xbit_r225_c186 bl[186] br[186] wl[225] vdd gnd cell_6t
Xbit_r226_c186 bl[186] br[186] wl[226] vdd gnd cell_6t
Xbit_r227_c186 bl[186] br[186] wl[227] vdd gnd cell_6t
Xbit_r228_c186 bl[186] br[186] wl[228] vdd gnd cell_6t
Xbit_r229_c186 bl[186] br[186] wl[229] vdd gnd cell_6t
Xbit_r230_c186 bl[186] br[186] wl[230] vdd gnd cell_6t
Xbit_r231_c186 bl[186] br[186] wl[231] vdd gnd cell_6t
Xbit_r232_c186 bl[186] br[186] wl[232] vdd gnd cell_6t
Xbit_r233_c186 bl[186] br[186] wl[233] vdd gnd cell_6t
Xbit_r234_c186 bl[186] br[186] wl[234] vdd gnd cell_6t
Xbit_r235_c186 bl[186] br[186] wl[235] vdd gnd cell_6t
Xbit_r236_c186 bl[186] br[186] wl[236] vdd gnd cell_6t
Xbit_r237_c186 bl[186] br[186] wl[237] vdd gnd cell_6t
Xbit_r238_c186 bl[186] br[186] wl[238] vdd gnd cell_6t
Xbit_r239_c186 bl[186] br[186] wl[239] vdd gnd cell_6t
Xbit_r240_c186 bl[186] br[186] wl[240] vdd gnd cell_6t
Xbit_r241_c186 bl[186] br[186] wl[241] vdd gnd cell_6t
Xbit_r242_c186 bl[186] br[186] wl[242] vdd gnd cell_6t
Xbit_r243_c186 bl[186] br[186] wl[243] vdd gnd cell_6t
Xbit_r244_c186 bl[186] br[186] wl[244] vdd gnd cell_6t
Xbit_r245_c186 bl[186] br[186] wl[245] vdd gnd cell_6t
Xbit_r246_c186 bl[186] br[186] wl[246] vdd gnd cell_6t
Xbit_r247_c186 bl[186] br[186] wl[247] vdd gnd cell_6t
Xbit_r248_c186 bl[186] br[186] wl[248] vdd gnd cell_6t
Xbit_r249_c186 bl[186] br[186] wl[249] vdd gnd cell_6t
Xbit_r250_c186 bl[186] br[186] wl[250] vdd gnd cell_6t
Xbit_r251_c186 bl[186] br[186] wl[251] vdd gnd cell_6t
Xbit_r252_c186 bl[186] br[186] wl[252] vdd gnd cell_6t
Xbit_r253_c186 bl[186] br[186] wl[253] vdd gnd cell_6t
Xbit_r254_c186 bl[186] br[186] wl[254] vdd gnd cell_6t
Xbit_r255_c186 bl[186] br[186] wl[255] vdd gnd cell_6t
Xbit_r0_c187 bl[187] br[187] wl[0] vdd gnd cell_6t
Xbit_r1_c187 bl[187] br[187] wl[1] vdd gnd cell_6t
Xbit_r2_c187 bl[187] br[187] wl[2] vdd gnd cell_6t
Xbit_r3_c187 bl[187] br[187] wl[3] vdd gnd cell_6t
Xbit_r4_c187 bl[187] br[187] wl[4] vdd gnd cell_6t
Xbit_r5_c187 bl[187] br[187] wl[5] vdd gnd cell_6t
Xbit_r6_c187 bl[187] br[187] wl[6] vdd gnd cell_6t
Xbit_r7_c187 bl[187] br[187] wl[7] vdd gnd cell_6t
Xbit_r8_c187 bl[187] br[187] wl[8] vdd gnd cell_6t
Xbit_r9_c187 bl[187] br[187] wl[9] vdd gnd cell_6t
Xbit_r10_c187 bl[187] br[187] wl[10] vdd gnd cell_6t
Xbit_r11_c187 bl[187] br[187] wl[11] vdd gnd cell_6t
Xbit_r12_c187 bl[187] br[187] wl[12] vdd gnd cell_6t
Xbit_r13_c187 bl[187] br[187] wl[13] vdd gnd cell_6t
Xbit_r14_c187 bl[187] br[187] wl[14] vdd gnd cell_6t
Xbit_r15_c187 bl[187] br[187] wl[15] vdd gnd cell_6t
Xbit_r16_c187 bl[187] br[187] wl[16] vdd gnd cell_6t
Xbit_r17_c187 bl[187] br[187] wl[17] vdd gnd cell_6t
Xbit_r18_c187 bl[187] br[187] wl[18] vdd gnd cell_6t
Xbit_r19_c187 bl[187] br[187] wl[19] vdd gnd cell_6t
Xbit_r20_c187 bl[187] br[187] wl[20] vdd gnd cell_6t
Xbit_r21_c187 bl[187] br[187] wl[21] vdd gnd cell_6t
Xbit_r22_c187 bl[187] br[187] wl[22] vdd gnd cell_6t
Xbit_r23_c187 bl[187] br[187] wl[23] vdd gnd cell_6t
Xbit_r24_c187 bl[187] br[187] wl[24] vdd gnd cell_6t
Xbit_r25_c187 bl[187] br[187] wl[25] vdd gnd cell_6t
Xbit_r26_c187 bl[187] br[187] wl[26] vdd gnd cell_6t
Xbit_r27_c187 bl[187] br[187] wl[27] vdd gnd cell_6t
Xbit_r28_c187 bl[187] br[187] wl[28] vdd gnd cell_6t
Xbit_r29_c187 bl[187] br[187] wl[29] vdd gnd cell_6t
Xbit_r30_c187 bl[187] br[187] wl[30] vdd gnd cell_6t
Xbit_r31_c187 bl[187] br[187] wl[31] vdd gnd cell_6t
Xbit_r32_c187 bl[187] br[187] wl[32] vdd gnd cell_6t
Xbit_r33_c187 bl[187] br[187] wl[33] vdd gnd cell_6t
Xbit_r34_c187 bl[187] br[187] wl[34] vdd gnd cell_6t
Xbit_r35_c187 bl[187] br[187] wl[35] vdd gnd cell_6t
Xbit_r36_c187 bl[187] br[187] wl[36] vdd gnd cell_6t
Xbit_r37_c187 bl[187] br[187] wl[37] vdd gnd cell_6t
Xbit_r38_c187 bl[187] br[187] wl[38] vdd gnd cell_6t
Xbit_r39_c187 bl[187] br[187] wl[39] vdd gnd cell_6t
Xbit_r40_c187 bl[187] br[187] wl[40] vdd gnd cell_6t
Xbit_r41_c187 bl[187] br[187] wl[41] vdd gnd cell_6t
Xbit_r42_c187 bl[187] br[187] wl[42] vdd gnd cell_6t
Xbit_r43_c187 bl[187] br[187] wl[43] vdd gnd cell_6t
Xbit_r44_c187 bl[187] br[187] wl[44] vdd gnd cell_6t
Xbit_r45_c187 bl[187] br[187] wl[45] vdd gnd cell_6t
Xbit_r46_c187 bl[187] br[187] wl[46] vdd gnd cell_6t
Xbit_r47_c187 bl[187] br[187] wl[47] vdd gnd cell_6t
Xbit_r48_c187 bl[187] br[187] wl[48] vdd gnd cell_6t
Xbit_r49_c187 bl[187] br[187] wl[49] vdd gnd cell_6t
Xbit_r50_c187 bl[187] br[187] wl[50] vdd gnd cell_6t
Xbit_r51_c187 bl[187] br[187] wl[51] vdd gnd cell_6t
Xbit_r52_c187 bl[187] br[187] wl[52] vdd gnd cell_6t
Xbit_r53_c187 bl[187] br[187] wl[53] vdd gnd cell_6t
Xbit_r54_c187 bl[187] br[187] wl[54] vdd gnd cell_6t
Xbit_r55_c187 bl[187] br[187] wl[55] vdd gnd cell_6t
Xbit_r56_c187 bl[187] br[187] wl[56] vdd gnd cell_6t
Xbit_r57_c187 bl[187] br[187] wl[57] vdd gnd cell_6t
Xbit_r58_c187 bl[187] br[187] wl[58] vdd gnd cell_6t
Xbit_r59_c187 bl[187] br[187] wl[59] vdd gnd cell_6t
Xbit_r60_c187 bl[187] br[187] wl[60] vdd gnd cell_6t
Xbit_r61_c187 bl[187] br[187] wl[61] vdd gnd cell_6t
Xbit_r62_c187 bl[187] br[187] wl[62] vdd gnd cell_6t
Xbit_r63_c187 bl[187] br[187] wl[63] vdd gnd cell_6t
Xbit_r64_c187 bl[187] br[187] wl[64] vdd gnd cell_6t
Xbit_r65_c187 bl[187] br[187] wl[65] vdd gnd cell_6t
Xbit_r66_c187 bl[187] br[187] wl[66] vdd gnd cell_6t
Xbit_r67_c187 bl[187] br[187] wl[67] vdd gnd cell_6t
Xbit_r68_c187 bl[187] br[187] wl[68] vdd gnd cell_6t
Xbit_r69_c187 bl[187] br[187] wl[69] vdd gnd cell_6t
Xbit_r70_c187 bl[187] br[187] wl[70] vdd gnd cell_6t
Xbit_r71_c187 bl[187] br[187] wl[71] vdd gnd cell_6t
Xbit_r72_c187 bl[187] br[187] wl[72] vdd gnd cell_6t
Xbit_r73_c187 bl[187] br[187] wl[73] vdd gnd cell_6t
Xbit_r74_c187 bl[187] br[187] wl[74] vdd gnd cell_6t
Xbit_r75_c187 bl[187] br[187] wl[75] vdd gnd cell_6t
Xbit_r76_c187 bl[187] br[187] wl[76] vdd gnd cell_6t
Xbit_r77_c187 bl[187] br[187] wl[77] vdd gnd cell_6t
Xbit_r78_c187 bl[187] br[187] wl[78] vdd gnd cell_6t
Xbit_r79_c187 bl[187] br[187] wl[79] vdd gnd cell_6t
Xbit_r80_c187 bl[187] br[187] wl[80] vdd gnd cell_6t
Xbit_r81_c187 bl[187] br[187] wl[81] vdd gnd cell_6t
Xbit_r82_c187 bl[187] br[187] wl[82] vdd gnd cell_6t
Xbit_r83_c187 bl[187] br[187] wl[83] vdd gnd cell_6t
Xbit_r84_c187 bl[187] br[187] wl[84] vdd gnd cell_6t
Xbit_r85_c187 bl[187] br[187] wl[85] vdd gnd cell_6t
Xbit_r86_c187 bl[187] br[187] wl[86] vdd gnd cell_6t
Xbit_r87_c187 bl[187] br[187] wl[87] vdd gnd cell_6t
Xbit_r88_c187 bl[187] br[187] wl[88] vdd gnd cell_6t
Xbit_r89_c187 bl[187] br[187] wl[89] vdd gnd cell_6t
Xbit_r90_c187 bl[187] br[187] wl[90] vdd gnd cell_6t
Xbit_r91_c187 bl[187] br[187] wl[91] vdd gnd cell_6t
Xbit_r92_c187 bl[187] br[187] wl[92] vdd gnd cell_6t
Xbit_r93_c187 bl[187] br[187] wl[93] vdd gnd cell_6t
Xbit_r94_c187 bl[187] br[187] wl[94] vdd gnd cell_6t
Xbit_r95_c187 bl[187] br[187] wl[95] vdd gnd cell_6t
Xbit_r96_c187 bl[187] br[187] wl[96] vdd gnd cell_6t
Xbit_r97_c187 bl[187] br[187] wl[97] vdd gnd cell_6t
Xbit_r98_c187 bl[187] br[187] wl[98] vdd gnd cell_6t
Xbit_r99_c187 bl[187] br[187] wl[99] vdd gnd cell_6t
Xbit_r100_c187 bl[187] br[187] wl[100] vdd gnd cell_6t
Xbit_r101_c187 bl[187] br[187] wl[101] vdd gnd cell_6t
Xbit_r102_c187 bl[187] br[187] wl[102] vdd gnd cell_6t
Xbit_r103_c187 bl[187] br[187] wl[103] vdd gnd cell_6t
Xbit_r104_c187 bl[187] br[187] wl[104] vdd gnd cell_6t
Xbit_r105_c187 bl[187] br[187] wl[105] vdd gnd cell_6t
Xbit_r106_c187 bl[187] br[187] wl[106] vdd gnd cell_6t
Xbit_r107_c187 bl[187] br[187] wl[107] vdd gnd cell_6t
Xbit_r108_c187 bl[187] br[187] wl[108] vdd gnd cell_6t
Xbit_r109_c187 bl[187] br[187] wl[109] vdd gnd cell_6t
Xbit_r110_c187 bl[187] br[187] wl[110] vdd gnd cell_6t
Xbit_r111_c187 bl[187] br[187] wl[111] vdd gnd cell_6t
Xbit_r112_c187 bl[187] br[187] wl[112] vdd gnd cell_6t
Xbit_r113_c187 bl[187] br[187] wl[113] vdd gnd cell_6t
Xbit_r114_c187 bl[187] br[187] wl[114] vdd gnd cell_6t
Xbit_r115_c187 bl[187] br[187] wl[115] vdd gnd cell_6t
Xbit_r116_c187 bl[187] br[187] wl[116] vdd gnd cell_6t
Xbit_r117_c187 bl[187] br[187] wl[117] vdd gnd cell_6t
Xbit_r118_c187 bl[187] br[187] wl[118] vdd gnd cell_6t
Xbit_r119_c187 bl[187] br[187] wl[119] vdd gnd cell_6t
Xbit_r120_c187 bl[187] br[187] wl[120] vdd gnd cell_6t
Xbit_r121_c187 bl[187] br[187] wl[121] vdd gnd cell_6t
Xbit_r122_c187 bl[187] br[187] wl[122] vdd gnd cell_6t
Xbit_r123_c187 bl[187] br[187] wl[123] vdd gnd cell_6t
Xbit_r124_c187 bl[187] br[187] wl[124] vdd gnd cell_6t
Xbit_r125_c187 bl[187] br[187] wl[125] vdd gnd cell_6t
Xbit_r126_c187 bl[187] br[187] wl[126] vdd gnd cell_6t
Xbit_r127_c187 bl[187] br[187] wl[127] vdd gnd cell_6t
Xbit_r128_c187 bl[187] br[187] wl[128] vdd gnd cell_6t
Xbit_r129_c187 bl[187] br[187] wl[129] vdd gnd cell_6t
Xbit_r130_c187 bl[187] br[187] wl[130] vdd gnd cell_6t
Xbit_r131_c187 bl[187] br[187] wl[131] vdd gnd cell_6t
Xbit_r132_c187 bl[187] br[187] wl[132] vdd gnd cell_6t
Xbit_r133_c187 bl[187] br[187] wl[133] vdd gnd cell_6t
Xbit_r134_c187 bl[187] br[187] wl[134] vdd gnd cell_6t
Xbit_r135_c187 bl[187] br[187] wl[135] vdd gnd cell_6t
Xbit_r136_c187 bl[187] br[187] wl[136] vdd gnd cell_6t
Xbit_r137_c187 bl[187] br[187] wl[137] vdd gnd cell_6t
Xbit_r138_c187 bl[187] br[187] wl[138] vdd gnd cell_6t
Xbit_r139_c187 bl[187] br[187] wl[139] vdd gnd cell_6t
Xbit_r140_c187 bl[187] br[187] wl[140] vdd gnd cell_6t
Xbit_r141_c187 bl[187] br[187] wl[141] vdd gnd cell_6t
Xbit_r142_c187 bl[187] br[187] wl[142] vdd gnd cell_6t
Xbit_r143_c187 bl[187] br[187] wl[143] vdd gnd cell_6t
Xbit_r144_c187 bl[187] br[187] wl[144] vdd gnd cell_6t
Xbit_r145_c187 bl[187] br[187] wl[145] vdd gnd cell_6t
Xbit_r146_c187 bl[187] br[187] wl[146] vdd gnd cell_6t
Xbit_r147_c187 bl[187] br[187] wl[147] vdd gnd cell_6t
Xbit_r148_c187 bl[187] br[187] wl[148] vdd gnd cell_6t
Xbit_r149_c187 bl[187] br[187] wl[149] vdd gnd cell_6t
Xbit_r150_c187 bl[187] br[187] wl[150] vdd gnd cell_6t
Xbit_r151_c187 bl[187] br[187] wl[151] vdd gnd cell_6t
Xbit_r152_c187 bl[187] br[187] wl[152] vdd gnd cell_6t
Xbit_r153_c187 bl[187] br[187] wl[153] vdd gnd cell_6t
Xbit_r154_c187 bl[187] br[187] wl[154] vdd gnd cell_6t
Xbit_r155_c187 bl[187] br[187] wl[155] vdd gnd cell_6t
Xbit_r156_c187 bl[187] br[187] wl[156] vdd gnd cell_6t
Xbit_r157_c187 bl[187] br[187] wl[157] vdd gnd cell_6t
Xbit_r158_c187 bl[187] br[187] wl[158] vdd gnd cell_6t
Xbit_r159_c187 bl[187] br[187] wl[159] vdd gnd cell_6t
Xbit_r160_c187 bl[187] br[187] wl[160] vdd gnd cell_6t
Xbit_r161_c187 bl[187] br[187] wl[161] vdd gnd cell_6t
Xbit_r162_c187 bl[187] br[187] wl[162] vdd gnd cell_6t
Xbit_r163_c187 bl[187] br[187] wl[163] vdd gnd cell_6t
Xbit_r164_c187 bl[187] br[187] wl[164] vdd gnd cell_6t
Xbit_r165_c187 bl[187] br[187] wl[165] vdd gnd cell_6t
Xbit_r166_c187 bl[187] br[187] wl[166] vdd gnd cell_6t
Xbit_r167_c187 bl[187] br[187] wl[167] vdd gnd cell_6t
Xbit_r168_c187 bl[187] br[187] wl[168] vdd gnd cell_6t
Xbit_r169_c187 bl[187] br[187] wl[169] vdd gnd cell_6t
Xbit_r170_c187 bl[187] br[187] wl[170] vdd gnd cell_6t
Xbit_r171_c187 bl[187] br[187] wl[171] vdd gnd cell_6t
Xbit_r172_c187 bl[187] br[187] wl[172] vdd gnd cell_6t
Xbit_r173_c187 bl[187] br[187] wl[173] vdd gnd cell_6t
Xbit_r174_c187 bl[187] br[187] wl[174] vdd gnd cell_6t
Xbit_r175_c187 bl[187] br[187] wl[175] vdd gnd cell_6t
Xbit_r176_c187 bl[187] br[187] wl[176] vdd gnd cell_6t
Xbit_r177_c187 bl[187] br[187] wl[177] vdd gnd cell_6t
Xbit_r178_c187 bl[187] br[187] wl[178] vdd gnd cell_6t
Xbit_r179_c187 bl[187] br[187] wl[179] vdd gnd cell_6t
Xbit_r180_c187 bl[187] br[187] wl[180] vdd gnd cell_6t
Xbit_r181_c187 bl[187] br[187] wl[181] vdd gnd cell_6t
Xbit_r182_c187 bl[187] br[187] wl[182] vdd gnd cell_6t
Xbit_r183_c187 bl[187] br[187] wl[183] vdd gnd cell_6t
Xbit_r184_c187 bl[187] br[187] wl[184] vdd gnd cell_6t
Xbit_r185_c187 bl[187] br[187] wl[185] vdd gnd cell_6t
Xbit_r186_c187 bl[187] br[187] wl[186] vdd gnd cell_6t
Xbit_r187_c187 bl[187] br[187] wl[187] vdd gnd cell_6t
Xbit_r188_c187 bl[187] br[187] wl[188] vdd gnd cell_6t
Xbit_r189_c187 bl[187] br[187] wl[189] vdd gnd cell_6t
Xbit_r190_c187 bl[187] br[187] wl[190] vdd gnd cell_6t
Xbit_r191_c187 bl[187] br[187] wl[191] vdd gnd cell_6t
Xbit_r192_c187 bl[187] br[187] wl[192] vdd gnd cell_6t
Xbit_r193_c187 bl[187] br[187] wl[193] vdd gnd cell_6t
Xbit_r194_c187 bl[187] br[187] wl[194] vdd gnd cell_6t
Xbit_r195_c187 bl[187] br[187] wl[195] vdd gnd cell_6t
Xbit_r196_c187 bl[187] br[187] wl[196] vdd gnd cell_6t
Xbit_r197_c187 bl[187] br[187] wl[197] vdd gnd cell_6t
Xbit_r198_c187 bl[187] br[187] wl[198] vdd gnd cell_6t
Xbit_r199_c187 bl[187] br[187] wl[199] vdd gnd cell_6t
Xbit_r200_c187 bl[187] br[187] wl[200] vdd gnd cell_6t
Xbit_r201_c187 bl[187] br[187] wl[201] vdd gnd cell_6t
Xbit_r202_c187 bl[187] br[187] wl[202] vdd gnd cell_6t
Xbit_r203_c187 bl[187] br[187] wl[203] vdd gnd cell_6t
Xbit_r204_c187 bl[187] br[187] wl[204] vdd gnd cell_6t
Xbit_r205_c187 bl[187] br[187] wl[205] vdd gnd cell_6t
Xbit_r206_c187 bl[187] br[187] wl[206] vdd gnd cell_6t
Xbit_r207_c187 bl[187] br[187] wl[207] vdd gnd cell_6t
Xbit_r208_c187 bl[187] br[187] wl[208] vdd gnd cell_6t
Xbit_r209_c187 bl[187] br[187] wl[209] vdd gnd cell_6t
Xbit_r210_c187 bl[187] br[187] wl[210] vdd gnd cell_6t
Xbit_r211_c187 bl[187] br[187] wl[211] vdd gnd cell_6t
Xbit_r212_c187 bl[187] br[187] wl[212] vdd gnd cell_6t
Xbit_r213_c187 bl[187] br[187] wl[213] vdd gnd cell_6t
Xbit_r214_c187 bl[187] br[187] wl[214] vdd gnd cell_6t
Xbit_r215_c187 bl[187] br[187] wl[215] vdd gnd cell_6t
Xbit_r216_c187 bl[187] br[187] wl[216] vdd gnd cell_6t
Xbit_r217_c187 bl[187] br[187] wl[217] vdd gnd cell_6t
Xbit_r218_c187 bl[187] br[187] wl[218] vdd gnd cell_6t
Xbit_r219_c187 bl[187] br[187] wl[219] vdd gnd cell_6t
Xbit_r220_c187 bl[187] br[187] wl[220] vdd gnd cell_6t
Xbit_r221_c187 bl[187] br[187] wl[221] vdd gnd cell_6t
Xbit_r222_c187 bl[187] br[187] wl[222] vdd gnd cell_6t
Xbit_r223_c187 bl[187] br[187] wl[223] vdd gnd cell_6t
Xbit_r224_c187 bl[187] br[187] wl[224] vdd gnd cell_6t
Xbit_r225_c187 bl[187] br[187] wl[225] vdd gnd cell_6t
Xbit_r226_c187 bl[187] br[187] wl[226] vdd gnd cell_6t
Xbit_r227_c187 bl[187] br[187] wl[227] vdd gnd cell_6t
Xbit_r228_c187 bl[187] br[187] wl[228] vdd gnd cell_6t
Xbit_r229_c187 bl[187] br[187] wl[229] vdd gnd cell_6t
Xbit_r230_c187 bl[187] br[187] wl[230] vdd gnd cell_6t
Xbit_r231_c187 bl[187] br[187] wl[231] vdd gnd cell_6t
Xbit_r232_c187 bl[187] br[187] wl[232] vdd gnd cell_6t
Xbit_r233_c187 bl[187] br[187] wl[233] vdd gnd cell_6t
Xbit_r234_c187 bl[187] br[187] wl[234] vdd gnd cell_6t
Xbit_r235_c187 bl[187] br[187] wl[235] vdd gnd cell_6t
Xbit_r236_c187 bl[187] br[187] wl[236] vdd gnd cell_6t
Xbit_r237_c187 bl[187] br[187] wl[237] vdd gnd cell_6t
Xbit_r238_c187 bl[187] br[187] wl[238] vdd gnd cell_6t
Xbit_r239_c187 bl[187] br[187] wl[239] vdd gnd cell_6t
Xbit_r240_c187 bl[187] br[187] wl[240] vdd gnd cell_6t
Xbit_r241_c187 bl[187] br[187] wl[241] vdd gnd cell_6t
Xbit_r242_c187 bl[187] br[187] wl[242] vdd gnd cell_6t
Xbit_r243_c187 bl[187] br[187] wl[243] vdd gnd cell_6t
Xbit_r244_c187 bl[187] br[187] wl[244] vdd gnd cell_6t
Xbit_r245_c187 bl[187] br[187] wl[245] vdd gnd cell_6t
Xbit_r246_c187 bl[187] br[187] wl[246] vdd gnd cell_6t
Xbit_r247_c187 bl[187] br[187] wl[247] vdd gnd cell_6t
Xbit_r248_c187 bl[187] br[187] wl[248] vdd gnd cell_6t
Xbit_r249_c187 bl[187] br[187] wl[249] vdd gnd cell_6t
Xbit_r250_c187 bl[187] br[187] wl[250] vdd gnd cell_6t
Xbit_r251_c187 bl[187] br[187] wl[251] vdd gnd cell_6t
Xbit_r252_c187 bl[187] br[187] wl[252] vdd gnd cell_6t
Xbit_r253_c187 bl[187] br[187] wl[253] vdd gnd cell_6t
Xbit_r254_c187 bl[187] br[187] wl[254] vdd gnd cell_6t
Xbit_r255_c187 bl[187] br[187] wl[255] vdd gnd cell_6t
Xbit_r0_c188 bl[188] br[188] wl[0] vdd gnd cell_6t
Xbit_r1_c188 bl[188] br[188] wl[1] vdd gnd cell_6t
Xbit_r2_c188 bl[188] br[188] wl[2] vdd gnd cell_6t
Xbit_r3_c188 bl[188] br[188] wl[3] vdd gnd cell_6t
Xbit_r4_c188 bl[188] br[188] wl[4] vdd gnd cell_6t
Xbit_r5_c188 bl[188] br[188] wl[5] vdd gnd cell_6t
Xbit_r6_c188 bl[188] br[188] wl[6] vdd gnd cell_6t
Xbit_r7_c188 bl[188] br[188] wl[7] vdd gnd cell_6t
Xbit_r8_c188 bl[188] br[188] wl[8] vdd gnd cell_6t
Xbit_r9_c188 bl[188] br[188] wl[9] vdd gnd cell_6t
Xbit_r10_c188 bl[188] br[188] wl[10] vdd gnd cell_6t
Xbit_r11_c188 bl[188] br[188] wl[11] vdd gnd cell_6t
Xbit_r12_c188 bl[188] br[188] wl[12] vdd gnd cell_6t
Xbit_r13_c188 bl[188] br[188] wl[13] vdd gnd cell_6t
Xbit_r14_c188 bl[188] br[188] wl[14] vdd gnd cell_6t
Xbit_r15_c188 bl[188] br[188] wl[15] vdd gnd cell_6t
Xbit_r16_c188 bl[188] br[188] wl[16] vdd gnd cell_6t
Xbit_r17_c188 bl[188] br[188] wl[17] vdd gnd cell_6t
Xbit_r18_c188 bl[188] br[188] wl[18] vdd gnd cell_6t
Xbit_r19_c188 bl[188] br[188] wl[19] vdd gnd cell_6t
Xbit_r20_c188 bl[188] br[188] wl[20] vdd gnd cell_6t
Xbit_r21_c188 bl[188] br[188] wl[21] vdd gnd cell_6t
Xbit_r22_c188 bl[188] br[188] wl[22] vdd gnd cell_6t
Xbit_r23_c188 bl[188] br[188] wl[23] vdd gnd cell_6t
Xbit_r24_c188 bl[188] br[188] wl[24] vdd gnd cell_6t
Xbit_r25_c188 bl[188] br[188] wl[25] vdd gnd cell_6t
Xbit_r26_c188 bl[188] br[188] wl[26] vdd gnd cell_6t
Xbit_r27_c188 bl[188] br[188] wl[27] vdd gnd cell_6t
Xbit_r28_c188 bl[188] br[188] wl[28] vdd gnd cell_6t
Xbit_r29_c188 bl[188] br[188] wl[29] vdd gnd cell_6t
Xbit_r30_c188 bl[188] br[188] wl[30] vdd gnd cell_6t
Xbit_r31_c188 bl[188] br[188] wl[31] vdd gnd cell_6t
Xbit_r32_c188 bl[188] br[188] wl[32] vdd gnd cell_6t
Xbit_r33_c188 bl[188] br[188] wl[33] vdd gnd cell_6t
Xbit_r34_c188 bl[188] br[188] wl[34] vdd gnd cell_6t
Xbit_r35_c188 bl[188] br[188] wl[35] vdd gnd cell_6t
Xbit_r36_c188 bl[188] br[188] wl[36] vdd gnd cell_6t
Xbit_r37_c188 bl[188] br[188] wl[37] vdd gnd cell_6t
Xbit_r38_c188 bl[188] br[188] wl[38] vdd gnd cell_6t
Xbit_r39_c188 bl[188] br[188] wl[39] vdd gnd cell_6t
Xbit_r40_c188 bl[188] br[188] wl[40] vdd gnd cell_6t
Xbit_r41_c188 bl[188] br[188] wl[41] vdd gnd cell_6t
Xbit_r42_c188 bl[188] br[188] wl[42] vdd gnd cell_6t
Xbit_r43_c188 bl[188] br[188] wl[43] vdd gnd cell_6t
Xbit_r44_c188 bl[188] br[188] wl[44] vdd gnd cell_6t
Xbit_r45_c188 bl[188] br[188] wl[45] vdd gnd cell_6t
Xbit_r46_c188 bl[188] br[188] wl[46] vdd gnd cell_6t
Xbit_r47_c188 bl[188] br[188] wl[47] vdd gnd cell_6t
Xbit_r48_c188 bl[188] br[188] wl[48] vdd gnd cell_6t
Xbit_r49_c188 bl[188] br[188] wl[49] vdd gnd cell_6t
Xbit_r50_c188 bl[188] br[188] wl[50] vdd gnd cell_6t
Xbit_r51_c188 bl[188] br[188] wl[51] vdd gnd cell_6t
Xbit_r52_c188 bl[188] br[188] wl[52] vdd gnd cell_6t
Xbit_r53_c188 bl[188] br[188] wl[53] vdd gnd cell_6t
Xbit_r54_c188 bl[188] br[188] wl[54] vdd gnd cell_6t
Xbit_r55_c188 bl[188] br[188] wl[55] vdd gnd cell_6t
Xbit_r56_c188 bl[188] br[188] wl[56] vdd gnd cell_6t
Xbit_r57_c188 bl[188] br[188] wl[57] vdd gnd cell_6t
Xbit_r58_c188 bl[188] br[188] wl[58] vdd gnd cell_6t
Xbit_r59_c188 bl[188] br[188] wl[59] vdd gnd cell_6t
Xbit_r60_c188 bl[188] br[188] wl[60] vdd gnd cell_6t
Xbit_r61_c188 bl[188] br[188] wl[61] vdd gnd cell_6t
Xbit_r62_c188 bl[188] br[188] wl[62] vdd gnd cell_6t
Xbit_r63_c188 bl[188] br[188] wl[63] vdd gnd cell_6t
Xbit_r64_c188 bl[188] br[188] wl[64] vdd gnd cell_6t
Xbit_r65_c188 bl[188] br[188] wl[65] vdd gnd cell_6t
Xbit_r66_c188 bl[188] br[188] wl[66] vdd gnd cell_6t
Xbit_r67_c188 bl[188] br[188] wl[67] vdd gnd cell_6t
Xbit_r68_c188 bl[188] br[188] wl[68] vdd gnd cell_6t
Xbit_r69_c188 bl[188] br[188] wl[69] vdd gnd cell_6t
Xbit_r70_c188 bl[188] br[188] wl[70] vdd gnd cell_6t
Xbit_r71_c188 bl[188] br[188] wl[71] vdd gnd cell_6t
Xbit_r72_c188 bl[188] br[188] wl[72] vdd gnd cell_6t
Xbit_r73_c188 bl[188] br[188] wl[73] vdd gnd cell_6t
Xbit_r74_c188 bl[188] br[188] wl[74] vdd gnd cell_6t
Xbit_r75_c188 bl[188] br[188] wl[75] vdd gnd cell_6t
Xbit_r76_c188 bl[188] br[188] wl[76] vdd gnd cell_6t
Xbit_r77_c188 bl[188] br[188] wl[77] vdd gnd cell_6t
Xbit_r78_c188 bl[188] br[188] wl[78] vdd gnd cell_6t
Xbit_r79_c188 bl[188] br[188] wl[79] vdd gnd cell_6t
Xbit_r80_c188 bl[188] br[188] wl[80] vdd gnd cell_6t
Xbit_r81_c188 bl[188] br[188] wl[81] vdd gnd cell_6t
Xbit_r82_c188 bl[188] br[188] wl[82] vdd gnd cell_6t
Xbit_r83_c188 bl[188] br[188] wl[83] vdd gnd cell_6t
Xbit_r84_c188 bl[188] br[188] wl[84] vdd gnd cell_6t
Xbit_r85_c188 bl[188] br[188] wl[85] vdd gnd cell_6t
Xbit_r86_c188 bl[188] br[188] wl[86] vdd gnd cell_6t
Xbit_r87_c188 bl[188] br[188] wl[87] vdd gnd cell_6t
Xbit_r88_c188 bl[188] br[188] wl[88] vdd gnd cell_6t
Xbit_r89_c188 bl[188] br[188] wl[89] vdd gnd cell_6t
Xbit_r90_c188 bl[188] br[188] wl[90] vdd gnd cell_6t
Xbit_r91_c188 bl[188] br[188] wl[91] vdd gnd cell_6t
Xbit_r92_c188 bl[188] br[188] wl[92] vdd gnd cell_6t
Xbit_r93_c188 bl[188] br[188] wl[93] vdd gnd cell_6t
Xbit_r94_c188 bl[188] br[188] wl[94] vdd gnd cell_6t
Xbit_r95_c188 bl[188] br[188] wl[95] vdd gnd cell_6t
Xbit_r96_c188 bl[188] br[188] wl[96] vdd gnd cell_6t
Xbit_r97_c188 bl[188] br[188] wl[97] vdd gnd cell_6t
Xbit_r98_c188 bl[188] br[188] wl[98] vdd gnd cell_6t
Xbit_r99_c188 bl[188] br[188] wl[99] vdd gnd cell_6t
Xbit_r100_c188 bl[188] br[188] wl[100] vdd gnd cell_6t
Xbit_r101_c188 bl[188] br[188] wl[101] vdd gnd cell_6t
Xbit_r102_c188 bl[188] br[188] wl[102] vdd gnd cell_6t
Xbit_r103_c188 bl[188] br[188] wl[103] vdd gnd cell_6t
Xbit_r104_c188 bl[188] br[188] wl[104] vdd gnd cell_6t
Xbit_r105_c188 bl[188] br[188] wl[105] vdd gnd cell_6t
Xbit_r106_c188 bl[188] br[188] wl[106] vdd gnd cell_6t
Xbit_r107_c188 bl[188] br[188] wl[107] vdd gnd cell_6t
Xbit_r108_c188 bl[188] br[188] wl[108] vdd gnd cell_6t
Xbit_r109_c188 bl[188] br[188] wl[109] vdd gnd cell_6t
Xbit_r110_c188 bl[188] br[188] wl[110] vdd gnd cell_6t
Xbit_r111_c188 bl[188] br[188] wl[111] vdd gnd cell_6t
Xbit_r112_c188 bl[188] br[188] wl[112] vdd gnd cell_6t
Xbit_r113_c188 bl[188] br[188] wl[113] vdd gnd cell_6t
Xbit_r114_c188 bl[188] br[188] wl[114] vdd gnd cell_6t
Xbit_r115_c188 bl[188] br[188] wl[115] vdd gnd cell_6t
Xbit_r116_c188 bl[188] br[188] wl[116] vdd gnd cell_6t
Xbit_r117_c188 bl[188] br[188] wl[117] vdd gnd cell_6t
Xbit_r118_c188 bl[188] br[188] wl[118] vdd gnd cell_6t
Xbit_r119_c188 bl[188] br[188] wl[119] vdd gnd cell_6t
Xbit_r120_c188 bl[188] br[188] wl[120] vdd gnd cell_6t
Xbit_r121_c188 bl[188] br[188] wl[121] vdd gnd cell_6t
Xbit_r122_c188 bl[188] br[188] wl[122] vdd gnd cell_6t
Xbit_r123_c188 bl[188] br[188] wl[123] vdd gnd cell_6t
Xbit_r124_c188 bl[188] br[188] wl[124] vdd gnd cell_6t
Xbit_r125_c188 bl[188] br[188] wl[125] vdd gnd cell_6t
Xbit_r126_c188 bl[188] br[188] wl[126] vdd gnd cell_6t
Xbit_r127_c188 bl[188] br[188] wl[127] vdd gnd cell_6t
Xbit_r128_c188 bl[188] br[188] wl[128] vdd gnd cell_6t
Xbit_r129_c188 bl[188] br[188] wl[129] vdd gnd cell_6t
Xbit_r130_c188 bl[188] br[188] wl[130] vdd gnd cell_6t
Xbit_r131_c188 bl[188] br[188] wl[131] vdd gnd cell_6t
Xbit_r132_c188 bl[188] br[188] wl[132] vdd gnd cell_6t
Xbit_r133_c188 bl[188] br[188] wl[133] vdd gnd cell_6t
Xbit_r134_c188 bl[188] br[188] wl[134] vdd gnd cell_6t
Xbit_r135_c188 bl[188] br[188] wl[135] vdd gnd cell_6t
Xbit_r136_c188 bl[188] br[188] wl[136] vdd gnd cell_6t
Xbit_r137_c188 bl[188] br[188] wl[137] vdd gnd cell_6t
Xbit_r138_c188 bl[188] br[188] wl[138] vdd gnd cell_6t
Xbit_r139_c188 bl[188] br[188] wl[139] vdd gnd cell_6t
Xbit_r140_c188 bl[188] br[188] wl[140] vdd gnd cell_6t
Xbit_r141_c188 bl[188] br[188] wl[141] vdd gnd cell_6t
Xbit_r142_c188 bl[188] br[188] wl[142] vdd gnd cell_6t
Xbit_r143_c188 bl[188] br[188] wl[143] vdd gnd cell_6t
Xbit_r144_c188 bl[188] br[188] wl[144] vdd gnd cell_6t
Xbit_r145_c188 bl[188] br[188] wl[145] vdd gnd cell_6t
Xbit_r146_c188 bl[188] br[188] wl[146] vdd gnd cell_6t
Xbit_r147_c188 bl[188] br[188] wl[147] vdd gnd cell_6t
Xbit_r148_c188 bl[188] br[188] wl[148] vdd gnd cell_6t
Xbit_r149_c188 bl[188] br[188] wl[149] vdd gnd cell_6t
Xbit_r150_c188 bl[188] br[188] wl[150] vdd gnd cell_6t
Xbit_r151_c188 bl[188] br[188] wl[151] vdd gnd cell_6t
Xbit_r152_c188 bl[188] br[188] wl[152] vdd gnd cell_6t
Xbit_r153_c188 bl[188] br[188] wl[153] vdd gnd cell_6t
Xbit_r154_c188 bl[188] br[188] wl[154] vdd gnd cell_6t
Xbit_r155_c188 bl[188] br[188] wl[155] vdd gnd cell_6t
Xbit_r156_c188 bl[188] br[188] wl[156] vdd gnd cell_6t
Xbit_r157_c188 bl[188] br[188] wl[157] vdd gnd cell_6t
Xbit_r158_c188 bl[188] br[188] wl[158] vdd gnd cell_6t
Xbit_r159_c188 bl[188] br[188] wl[159] vdd gnd cell_6t
Xbit_r160_c188 bl[188] br[188] wl[160] vdd gnd cell_6t
Xbit_r161_c188 bl[188] br[188] wl[161] vdd gnd cell_6t
Xbit_r162_c188 bl[188] br[188] wl[162] vdd gnd cell_6t
Xbit_r163_c188 bl[188] br[188] wl[163] vdd gnd cell_6t
Xbit_r164_c188 bl[188] br[188] wl[164] vdd gnd cell_6t
Xbit_r165_c188 bl[188] br[188] wl[165] vdd gnd cell_6t
Xbit_r166_c188 bl[188] br[188] wl[166] vdd gnd cell_6t
Xbit_r167_c188 bl[188] br[188] wl[167] vdd gnd cell_6t
Xbit_r168_c188 bl[188] br[188] wl[168] vdd gnd cell_6t
Xbit_r169_c188 bl[188] br[188] wl[169] vdd gnd cell_6t
Xbit_r170_c188 bl[188] br[188] wl[170] vdd gnd cell_6t
Xbit_r171_c188 bl[188] br[188] wl[171] vdd gnd cell_6t
Xbit_r172_c188 bl[188] br[188] wl[172] vdd gnd cell_6t
Xbit_r173_c188 bl[188] br[188] wl[173] vdd gnd cell_6t
Xbit_r174_c188 bl[188] br[188] wl[174] vdd gnd cell_6t
Xbit_r175_c188 bl[188] br[188] wl[175] vdd gnd cell_6t
Xbit_r176_c188 bl[188] br[188] wl[176] vdd gnd cell_6t
Xbit_r177_c188 bl[188] br[188] wl[177] vdd gnd cell_6t
Xbit_r178_c188 bl[188] br[188] wl[178] vdd gnd cell_6t
Xbit_r179_c188 bl[188] br[188] wl[179] vdd gnd cell_6t
Xbit_r180_c188 bl[188] br[188] wl[180] vdd gnd cell_6t
Xbit_r181_c188 bl[188] br[188] wl[181] vdd gnd cell_6t
Xbit_r182_c188 bl[188] br[188] wl[182] vdd gnd cell_6t
Xbit_r183_c188 bl[188] br[188] wl[183] vdd gnd cell_6t
Xbit_r184_c188 bl[188] br[188] wl[184] vdd gnd cell_6t
Xbit_r185_c188 bl[188] br[188] wl[185] vdd gnd cell_6t
Xbit_r186_c188 bl[188] br[188] wl[186] vdd gnd cell_6t
Xbit_r187_c188 bl[188] br[188] wl[187] vdd gnd cell_6t
Xbit_r188_c188 bl[188] br[188] wl[188] vdd gnd cell_6t
Xbit_r189_c188 bl[188] br[188] wl[189] vdd gnd cell_6t
Xbit_r190_c188 bl[188] br[188] wl[190] vdd gnd cell_6t
Xbit_r191_c188 bl[188] br[188] wl[191] vdd gnd cell_6t
Xbit_r192_c188 bl[188] br[188] wl[192] vdd gnd cell_6t
Xbit_r193_c188 bl[188] br[188] wl[193] vdd gnd cell_6t
Xbit_r194_c188 bl[188] br[188] wl[194] vdd gnd cell_6t
Xbit_r195_c188 bl[188] br[188] wl[195] vdd gnd cell_6t
Xbit_r196_c188 bl[188] br[188] wl[196] vdd gnd cell_6t
Xbit_r197_c188 bl[188] br[188] wl[197] vdd gnd cell_6t
Xbit_r198_c188 bl[188] br[188] wl[198] vdd gnd cell_6t
Xbit_r199_c188 bl[188] br[188] wl[199] vdd gnd cell_6t
Xbit_r200_c188 bl[188] br[188] wl[200] vdd gnd cell_6t
Xbit_r201_c188 bl[188] br[188] wl[201] vdd gnd cell_6t
Xbit_r202_c188 bl[188] br[188] wl[202] vdd gnd cell_6t
Xbit_r203_c188 bl[188] br[188] wl[203] vdd gnd cell_6t
Xbit_r204_c188 bl[188] br[188] wl[204] vdd gnd cell_6t
Xbit_r205_c188 bl[188] br[188] wl[205] vdd gnd cell_6t
Xbit_r206_c188 bl[188] br[188] wl[206] vdd gnd cell_6t
Xbit_r207_c188 bl[188] br[188] wl[207] vdd gnd cell_6t
Xbit_r208_c188 bl[188] br[188] wl[208] vdd gnd cell_6t
Xbit_r209_c188 bl[188] br[188] wl[209] vdd gnd cell_6t
Xbit_r210_c188 bl[188] br[188] wl[210] vdd gnd cell_6t
Xbit_r211_c188 bl[188] br[188] wl[211] vdd gnd cell_6t
Xbit_r212_c188 bl[188] br[188] wl[212] vdd gnd cell_6t
Xbit_r213_c188 bl[188] br[188] wl[213] vdd gnd cell_6t
Xbit_r214_c188 bl[188] br[188] wl[214] vdd gnd cell_6t
Xbit_r215_c188 bl[188] br[188] wl[215] vdd gnd cell_6t
Xbit_r216_c188 bl[188] br[188] wl[216] vdd gnd cell_6t
Xbit_r217_c188 bl[188] br[188] wl[217] vdd gnd cell_6t
Xbit_r218_c188 bl[188] br[188] wl[218] vdd gnd cell_6t
Xbit_r219_c188 bl[188] br[188] wl[219] vdd gnd cell_6t
Xbit_r220_c188 bl[188] br[188] wl[220] vdd gnd cell_6t
Xbit_r221_c188 bl[188] br[188] wl[221] vdd gnd cell_6t
Xbit_r222_c188 bl[188] br[188] wl[222] vdd gnd cell_6t
Xbit_r223_c188 bl[188] br[188] wl[223] vdd gnd cell_6t
Xbit_r224_c188 bl[188] br[188] wl[224] vdd gnd cell_6t
Xbit_r225_c188 bl[188] br[188] wl[225] vdd gnd cell_6t
Xbit_r226_c188 bl[188] br[188] wl[226] vdd gnd cell_6t
Xbit_r227_c188 bl[188] br[188] wl[227] vdd gnd cell_6t
Xbit_r228_c188 bl[188] br[188] wl[228] vdd gnd cell_6t
Xbit_r229_c188 bl[188] br[188] wl[229] vdd gnd cell_6t
Xbit_r230_c188 bl[188] br[188] wl[230] vdd gnd cell_6t
Xbit_r231_c188 bl[188] br[188] wl[231] vdd gnd cell_6t
Xbit_r232_c188 bl[188] br[188] wl[232] vdd gnd cell_6t
Xbit_r233_c188 bl[188] br[188] wl[233] vdd gnd cell_6t
Xbit_r234_c188 bl[188] br[188] wl[234] vdd gnd cell_6t
Xbit_r235_c188 bl[188] br[188] wl[235] vdd gnd cell_6t
Xbit_r236_c188 bl[188] br[188] wl[236] vdd gnd cell_6t
Xbit_r237_c188 bl[188] br[188] wl[237] vdd gnd cell_6t
Xbit_r238_c188 bl[188] br[188] wl[238] vdd gnd cell_6t
Xbit_r239_c188 bl[188] br[188] wl[239] vdd gnd cell_6t
Xbit_r240_c188 bl[188] br[188] wl[240] vdd gnd cell_6t
Xbit_r241_c188 bl[188] br[188] wl[241] vdd gnd cell_6t
Xbit_r242_c188 bl[188] br[188] wl[242] vdd gnd cell_6t
Xbit_r243_c188 bl[188] br[188] wl[243] vdd gnd cell_6t
Xbit_r244_c188 bl[188] br[188] wl[244] vdd gnd cell_6t
Xbit_r245_c188 bl[188] br[188] wl[245] vdd gnd cell_6t
Xbit_r246_c188 bl[188] br[188] wl[246] vdd gnd cell_6t
Xbit_r247_c188 bl[188] br[188] wl[247] vdd gnd cell_6t
Xbit_r248_c188 bl[188] br[188] wl[248] vdd gnd cell_6t
Xbit_r249_c188 bl[188] br[188] wl[249] vdd gnd cell_6t
Xbit_r250_c188 bl[188] br[188] wl[250] vdd gnd cell_6t
Xbit_r251_c188 bl[188] br[188] wl[251] vdd gnd cell_6t
Xbit_r252_c188 bl[188] br[188] wl[252] vdd gnd cell_6t
Xbit_r253_c188 bl[188] br[188] wl[253] vdd gnd cell_6t
Xbit_r254_c188 bl[188] br[188] wl[254] vdd gnd cell_6t
Xbit_r255_c188 bl[188] br[188] wl[255] vdd gnd cell_6t
Xbit_r0_c189 bl[189] br[189] wl[0] vdd gnd cell_6t
Xbit_r1_c189 bl[189] br[189] wl[1] vdd gnd cell_6t
Xbit_r2_c189 bl[189] br[189] wl[2] vdd gnd cell_6t
Xbit_r3_c189 bl[189] br[189] wl[3] vdd gnd cell_6t
Xbit_r4_c189 bl[189] br[189] wl[4] vdd gnd cell_6t
Xbit_r5_c189 bl[189] br[189] wl[5] vdd gnd cell_6t
Xbit_r6_c189 bl[189] br[189] wl[6] vdd gnd cell_6t
Xbit_r7_c189 bl[189] br[189] wl[7] vdd gnd cell_6t
Xbit_r8_c189 bl[189] br[189] wl[8] vdd gnd cell_6t
Xbit_r9_c189 bl[189] br[189] wl[9] vdd gnd cell_6t
Xbit_r10_c189 bl[189] br[189] wl[10] vdd gnd cell_6t
Xbit_r11_c189 bl[189] br[189] wl[11] vdd gnd cell_6t
Xbit_r12_c189 bl[189] br[189] wl[12] vdd gnd cell_6t
Xbit_r13_c189 bl[189] br[189] wl[13] vdd gnd cell_6t
Xbit_r14_c189 bl[189] br[189] wl[14] vdd gnd cell_6t
Xbit_r15_c189 bl[189] br[189] wl[15] vdd gnd cell_6t
Xbit_r16_c189 bl[189] br[189] wl[16] vdd gnd cell_6t
Xbit_r17_c189 bl[189] br[189] wl[17] vdd gnd cell_6t
Xbit_r18_c189 bl[189] br[189] wl[18] vdd gnd cell_6t
Xbit_r19_c189 bl[189] br[189] wl[19] vdd gnd cell_6t
Xbit_r20_c189 bl[189] br[189] wl[20] vdd gnd cell_6t
Xbit_r21_c189 bl[189] br[189] wl[21] vdd gnd cell_6t
Xbit_r22_c189 bl[189] br[189] wl[22] vdd gnd cell_6t
Xbit_r23_c189 bl[189] br[189] wl[23] vdd gnd cell_6t
Xbit_r24_c189 bl[189] br[189] wl[24] vdd gnd cell_6t
Xbit_r25_c189 bl[189] br[189] wl[25] vdd gnd cell_6t
Xbit_r26_c189 bl[189] br[189] wl[26] vdd gnd cell_6t
Xbit_r27_c189 bl[189] br[189] wl[27] vdd gnd cell_6t
Xbit_r28_c189 bl[189] br[189] wl[28] vdd gnd cell_6t
Xbit_r29_c189 bl[189] br[189] wl[29] vdd gnd cell_6t
Xbit_r30_c189 bl[189] br[189] wl[30] vdd gnd cell_6t
Xbit_r31_c189 bl[189] br[189] wl[31] vdd gnd cell_6t
Xbit_r32_c189 bl[189] br[189] wl[32] vdd gnd cell_6t
Xbit_r33_c189 bl[189] br[189] wl[33] vdd gnd cell_6t
Xbit_r34_c189 bl[189] br[189] wl[34] vdd gnd cell_6t
Xbit_r35_c189 bl[189] br[189] wl[35] vdd gnd cell_6t
Xbit_r36_c189 bl[189] br[189] wl[36] vdd gnd cell_6t
Xbit_r37_c189 bl[189] br[189] wl[37] vdd gnd cell_6t
Xbit_r38_c189 bl[189] br[189] wl[38] vdd gnd cell_6t
Xbit_r39_c189 bl[189] br[189] wl[39] vdd gnd cell_6t
Xbit_r40_c189 bl[189] br[189] wl[40] vdd gnd cell_6t
Xbit_r41_c189 bl[189] br[189] wl[41] vdd gnd cell_6t
Xbit_r42_c189 bl[189] br[189] wl[42] vdd gnd cell_6t
Xbit_r43_c189 bl[189] br[189] wl[43] vdd gnd cell_6t
Xbit_r44_c189 bl[189] br[189] wl[44] vdd gnd cell_6t
Xbit_r45_c189 bl[189] br[189] wl[45] vdd gnd cell_6t
Xbit_r46_c189 bl[189] br[189] wl[46] vdd gnd cell_6t
Xbit_r47_c189 bl[189] br[189] wl[47] vdd gnd cell_6t
Xbit_r48_c189 bl[189] br[189] wl[48] vdd gnd cell_6t
Xbit_r49_c189 bl[189] br[189] wl[49] vdd gnd cell_6t
Xbit_r50_c189 bl[189] br[189] wl[50] vdd gnd cell_6t
Xbit_r51_c189 bl[189] br[189] wl[51] vdd gnd cell_6t
Xbit_r52_c189 bl[189] br[189] wl[52] vdd gnd cell_6t
Xbit_r53_c189 bl[189] br[189] wl[53] vdd gnd cell_6t
Xbit_r54_c189 bl[189] br[189] wl[54] vdd gnd cell_6t
Xbit_r55_c189 bl[189] br[189] wl[55] vdd gnd cell_6t
Xbit_r56_c189 bl[189] br[189] wl[56] vdd gnd cell_6t
Xbit_r57_c189 bl[189] br[189] wl[57] vdd gnd cell_6t
Xbit_r58_c189 bl[189] br[189] wl[58] vdd gnd cell_6t
Xbit_r59_c189 bl[189] br[189] wl[59] vdd gnd cell_6t
Xbit_r60_c189 bl[189] br[189] wl[60] vdd gnd cell_6t
Xbit_r61_c189 bl[189] br[189] wl[61] vdd gnd cell_6t
Xbit_r62_c189 bl[189] br[189] wl[62] vdd gnd cell_6t
Xbit_r63_c189 bl[189] br[189] wl[63] vdd gnd cell_6t
Xbit_r64_c189 bl[189] br[189] wl[64] vdd gnd cell_6t
Xbit_r65_c189 bl[189] br[189] wl[65] vdd gnd cell_6t
Xbit_r66_c189 bl[189] br[189] wl[66] vdd gnd cell_6t
Xbit_r67_c189 bl[189] br[189] wl[67] vdd gnd cell_6t
Xbit_r68_c189 bl[189] br[189] wl[68] vdd gnd cell_6t
Xbit_r69_c189 bl[189] br[189] wl[69] vdd gnd cell_6t
Xbit_r70_c189 bl[189] br[189] wl[70] vdd gnd cell_6t
Xbit_r71_c189 bl[189] br[189] wl[71] vdd gnd cell_6t
Xbit_r72_c189 bl[189] br[189] wl[72] vdd gnd cell_6t
Xbit_r73_c189 bl[189] br[189] wl[73] vdd gnd cell_6t
Xbit_r74_c189 bl[189] br[189] wl[74] vdd gnd cell_6t
Xbit_r75_c189 bl[189] br[189] wl[75] vdd gnd cell_6t
Xbit_r76_c189 bl[189] br[189] wl[76] vdd gnd cell_6t
Xbit_r77_c189 bl[189] br[189] wl[77] vdd gnd cell_6t
Xbit_r78_c189 bl[189] br[189] wl[78] vdd gnd cell_6t
Xbit_r79_c189 bl[189] br[189] wl[79] vdd gnd cell_6t
Xbit_r80_c189 bl[189] br[189] wl[80] vdd gnd cell_6t
Xbit_r81_c189 bl[189] br[189] wl[81] vdd gnd cell_6t
Xbit_r82_c189 bl[189] br[189] wl[82] vdd gnd cell_6t
Xbit_r83_c189 bl[189] br[189] wl[83] vdd gnd cell_6t
Xbit_r84_c189 bl[189] br[189] wl[84] vdd gnd cell_6t
Xbit_r85_c189 bl[189] br[189] wl[85] vdd gnd cell_6t
Xbit_r86_c189 bl[189] br[189] wl[86] vdd gnd cell_6t
Xbit_r87_c189 bl[189] br[189] wl[87] vdd gnd cell_6t
Xbit_r88_c189 bl[189] br[189] wl[88] vdd gnd cell_6t
Xbit_r89_c189 bl[189] br[189] wl[89] vdd gnd cell_6t
Xbit_r90_c189 bl[189] br[189] wl[90] vdd gnd cell_6t
Xbit_r91_c189 bl[189] br[189] wl[91] vdd gnd cell_6t
Xbit_r92_c189 bl[189] br[189] wl[92] vdd gnd cell_6t
Xbit_r93_c189 bl[189] br[189] wl[93] vdd gnd cell_6t
Xbit_r94_c189 bl[189] br[189] wl[94] vdd gnd cell_6t
Xbit_r95_c189 bl[189] br[189] wl[95] vdd gnd cell_6t
Xbit_r96_c189 bl[189] br[189] wl[96] vdd gnd cell_6t
Xbit_r97_c189 bl[189] br[189] wl[97] vdd gnd cell_6t
Xbit_r98_c189 bl[189] br[189] wl[98] vdd gnd cell_6t
Xbit_r99_c189 bl[189] br[189] wl[99] vdd gnd cell_6t
Xbit_r100_c189 bl[189] br[189] wl[100] vdd gnd cell_6t
Xbit_r101_c189 bl[189] br[189] wl[101] vdd gnd cell_6t
Xbit_r102_c189 bl[189] br[189] wl[102] vdd gnd cell_6t
Xbit_r103_c189 bl[189] br[189] wl[103] vdd gnd cell_6t
Xbit_r104_c189 bl[189] br[189] wl[104] vdd gnd cell_6t
Xbit_r105_c189 bl[189] br[189] wl[105] vdd gnd cell_6t
Xbit_r106_c189 bl[189] br[189] wl[106] vdd gnd cell_6t
Xbit_r107_c189 bl[189] br[189] wl[107] vdd gnd cell_6t
Xbit_r108_c189 bl[189] br[189] wl[108] vdd gnd cell_6t
Xbit_r109_c189 bl[189] br[189] wl[109] vdd gnd cell_6t
Xbit_r110_c189 bl[189] br[189] wl[110] vdd gnd cell_6t
Xbit_r111_c189 bl[189] br[189] wl[111] vdd gnd cell_6t
Xbit_r112_c189 bl[189] br[189] wl[112] vdd gnd cell_6t
Xbit_r113_c189 bl[189] br[189] wl[113] vdd gnd cell_6t
Xbit_r114_c189 bl[189] br[189] wl[114] vdd gnd cell_6t
Xbit_r115_c189 bl[189] br[189] wl[115] vdd gnd cell_6t
Xbit_r116_c189 bl[189] br[189] wl[116] vdd gnd cell_6t
Xbit_r117_c189 bl[189] br[189] wl[117] vdd gnd cell_6t
Xbit_r118_c189 bl[189] br[189] wl[118] vdd gnd cell_6t
Xbit_r119_c189 bl[189] br[189] wl[119] vdd gnd cell_6t
Xbit_r120_c189 bl[189] br[189] wl[120] vdd gnd cell_6t
Xbit_r121_c189 bl[189] br[189] wl[121] vdd gnd cell_6t
Xbit_r122_c189 bl[189] br[189] wl[122] vdd gnd cell_6t
Xbit_r123_c189 bl[189] br[189] wl[123] vdd gnd cell_6t
Xbit_r124_c189 bl[189] br[189] wl[124] vdd gnd cell_6t
Xbit_r125_c189 bl[189] br[189] wl[125] vdd gnd cell_6t
Xbit_r126_c189 bl[189] br[189] wl[126] vdd gnd cell_6t
Xbit_r127_c189 bl[189] br[189] wl[127] vdd gnd cell_6t
Xbit_r128_c189 bl[189] br[189] wl[128] vdd gnd cell_6t
Xbit_r129_c189 bl[189] br[189] wl[129] vdd gnd cell_6t
Xbit_r130_c189 bl[189] br[189] wl[130] vdd gnd cell_6t
Xbit_r131_c189 bl[189] br[189] wl[131] vdd gnd cell_6t
Xbit_r132_c189 bl[189] br[189] wl[132] vdd gnd cell_6t
Xbit_r133_c189 bl[189] br[189] wl[133] vdd gnd cell_6t
Xbit_r134_c189 bl[189] br[189] wl[134] vdd gnd cell_6t
Xbit_r135_c189 bl[189] br[189] wl[135] vdd gnd cell_6t
Xbit_r136_c189 bl[189] br[189] wl[136] vdd gnd cell_6t
Xbit_r137_c189 bl[189] br[189] wl[137] vdd gnd cell_6t
Xbit_r138_c189 bl[189] br[189] wl[138] vdd gnd cell_6t
Xbit_r139_c189 bl[189] br[189] wl[139] vdd gnd cell_6t
Xbit_r140_c189 bl[189] br[189] wl[140] vdd gnd cell_6t
Xbit_r141_c189 bl[189] br[189] wl[141] vdd gnd cell_6t
Xbit_r142_c189 bl[189] br[189] wl[142] vdd gnd cell_6t
Xbit_r143_c189 bl[189] br[189] wl[143] vdd gnd cell_6t
Xbit_r144_c189 bl[189] br[189] wl[144] vdd gnd cell_6t
Xbit_r145_c189 bl[189] br[189] wl[145] vdd gnd cell_6t
Xbit_r146_c189 bl[189] br[189] wl[146] vdd gnd cell_6t
Xbit_r147_c189 bl[189] br[189] wl[147] vdd gnd cell_6t
Xbit_r148_c189 bl[189] br[189] wl[148] vdd gnd cell_6t
Xbit_r149_c189 bl[189] br[189] wl[149] vdd gnd cell_6t
Xbit_r150_c189 bl[189] br[189] wl[150] vdd gnd cell_6t
Xbit_r151_c189 bl[189] br[189] wl[151] vdd gnd cell_6t
Xbit_r152_c189 bl[189] br[189] wl[152] vdd gnd cell_6t
Xbit_r153_c189 bl[189] br[189] wl[153] vdd gnd cell_6t
Xbit_r154_c189 bl[189] br[189] wl[154] vdd gnd cell_6t
Xbit_r155_c189 bl[189] br[189] wl[155] vdd gnd cell_6t
Xbit_r156_c189 bl[189] br[189] wl[156] vdd gnd cell_6t
Xbit_r157_c189 bl[189] br[189] wl[157] vdd gnd cell_6t
Xbit_r158_c189 bl[189] br[189] wl[158] vdd gnd cell_6t
Xbit_r159_c189 bl[189] br[189] wl[159] vdd gnd cell_6t
Xbit_r160_c189 bl[189] br[189] wl[160] vdd gnd cell_6t
Xbit_r161_c189 bl[189] br[189] wl[161] vdd gnd cell_6t
Xbit_r162_c189 bl[189] br[189] wl[162] vdd gnd cell_6t
Xbit_r163_c189 bl[189] br[189] wl[163] vdd gnd cell_6t
Xbit_r164_c189 bl[189] br[189] wl[164] vdd gnd cell_6t
Xbit_r165_c189 bl[189] br[189] wl[165] vdd gnd cell_6t
Xbit_r166_c189 bl[189] br[189] wl[166] vdd gnd cell_6t
Xbit_r167_c189 bl[189] br[189] wl[167] vdd gnd cell_6t
Xbit_r168_c189 bl[189] br[189] wl[168] vdd gnd cell_6t
Xbit_r169_c189 bl[189] br[189] wl[169] vdd gnd cell_6t
Xbit_r170_c189 bl[189] br[189] wl[170] vdd gnd cell_6t
Xbit_r171_c189 bl[189] br[189] wl[171] vdd gnd cell_6t
Xbit_r172_c189 bl[189] br[189] wl[172] vdd gnd cell_6t
Xbit_r173_c189 bl[189] br[189] wl[173] vdd gnd cell_6t
Xbit_r174_c189 bl[189] br[189] wl[174] vdd gnd cell_6t
Xbit_r175_c189 bl[189] br[189] wl[175] vdd gnd cell_6t
Xbit_r176_c189 bl[189] br[189] wl[176] vdd gnd cell_6t
Xbit_r177_c189 bl[189] br[189] wl[177] vdd gnd cell_6t
Xbit_r178_c189 bl[189] br[189] wl[178] vdd gnd cell_6t
Xbit_r179_c189 bl[189] br[189] wl[179] vdd gnd cell_6t
Xbit_r180_c189 bl[189] br[189] wl[180] vdd gnd cell_6t
Xbit_r181_c189 bl[189] br[189] wl[181] vdd gnd cell_6t
Xbit_r182_c189 bl[189] br[189] wl[182] vdd gnd cell_6t
Xbit_r183_c189 bl[189] br[189] wl[183] vdd gnd cell_6t
Xbit_r184_c189 bl[189] br[189] wl[184] vdd gnd cell_6t
Xbit_r185_c189 bl[189] br[189] wl[185] vdd gnd cell_6t
Xbit_r186_c189 bl[189] br[189] wl[186] vdd gnd cell_6t
Xbit_r187_c189 bl[189] br[189] wl[187] vdd gnd cell_6t
Xbit_r188_c189 bl[189] br[189] wl[188] vdd gnd cell_6t
Xbit_r189_c189 bl[189] br[189] wl[189] vdd gnd cell_6t
Xbit_r190_c189 bl[189] br[189] wl[190] vdd gnd cell_6t
Xbit_r191_c189 bl[189] br[189] wl[191] vdd gnd cell_6t
Xbit_r192_c189 bl[189] br[189] wl[192] vdd gnd cell_6t
Xbit_r193_c189 bl[189] br[189] wl[193] vdd gnd cell_6t
Xbit_r194_c189 bl[189] br[189] wl[194] vdd gnd cell_6t
Xbit_r195_c189 bl[189] br[189] wl[195] vdd gnd cell_6t
Xbit_r196_c189 bl[189] br[189] wl[196] vdd gnd cell_6t
Xbit_r197_c189 bl[189] br[189] wl[197] vdd gnd cell_6t
Xbit_r198_c189 bl[189] br[189] wl[198] vdd gnd cell_6t
Xbit_r199_c189 bl[189] br[189] wl[199] vdd gnd cell_6t
Xbit_r200_c189 bl[189] br[189] wl[200] vdd gnd cell_6t
Xbit_r201_c189 bl[189] br[189] wl[201] vdd gnd cell_6t
Xbit_r202_c189 bl[189] br[189] wl[202] vdd gnd cell_6t
Xbit_r203_c189 bl[189] br[189] wl[203] vdd gnd cell_6t
Xbit_r204_c189 bl[189] br[189] wl[204] vdd gnd cell_6t
Xbit_r205_c189 bl[189] br[189] wl[205] vdd gnd cell_6t
Xbit_r206_c189 bl[189] br[189] wl[206] vdd gnd cell_6t
Xbit_r207_c189 bl[189] br[189] wl[207] vdd gnd cell_6t
Xbit_r208_c189 bl[189] br[189] wl[208] vdd gnd cell_6t
Xbit_r209_c189 bl[189] br[189] wl[209] vdd gnd cell_6t
Xbit_r210_c189 bl[189] br[189] wl[210] vdd gnd cell_6t
Xbit_r211_c189 bl[189] br[189] wl[211] vdd gnd cell_6t
Xbit_r212_c189 bl[189] br[189] wl[212] vdd gnd cell_6t
Xbit_r213_c189 bl[189] br[189] wl[213] vdd gnd cell_6t
Xbit_r214_c189 bl[189] br[189] wl[214] vdd gnd cell_6t
Xbit_r215_c189 bl[189] br[189] wl[215] vdd gnd cell_6t
Xbit_r216_c189 bl[189] br[189] wl[216] vdd gnd cell_6t
Xbit_r217_c189 bl[189] br[189] wl[217] vdd gnd cell_6t
Xbit_r218_c189 bl[189] br[189] wl[218] vdd gnd cell_6t
Xbit_r219_c189 bl[189] br[189] wl[219] vdd gnd cell_6t
Xbit_r220_c189 bl[189] br[189] wl[220] vdd gnd cell_6t
Xbit_r221_c189 bl[189] br[189] wl[221] vdd gnd cell_6t
Xbit_r222_c189 bl[189] br[189] wl[222] vdd gnd cell_6t
Xbit_r223_c189 bl[189] br[189] wl[223] vdd gnd cell_6t
Xbit_r224_c189 bl[189] br[189] wl[224] vdd gnd cell_6t
Xbit_r225_c189 bl[189] br[189] wl[225] vdd gnd cell_6t
Xbit_r226_c189 bl[189] br[189] wl[226] vdd gnd cell_6t
Xbit_r227_c189 bl[189] br[189] wl[227] vdd gnd cell_6t
Xbit_r228_c189 bl[189] br[189] wl[228] vdd gnd cell_6t
Xbit_r229_c189 bl[189] br[189] wl[229] vdd gnd cell_6t
Xbit_r230_c189 bl[189] br[189] wl[230] vdd gnd cell_6t
Xbit_r231_c189 bl[189] br[189] wl[231] vdd gnd cell_6t
Xbit_r232_c189 bl[189] br[189] wl[232] vdd gnd cell_6t
Xbit_r233_c189 bl[189] br[189] wl[233] vdd gnd cell_6t
Xbit_r234_c189 bl[189] br[189] wl[234] vdd gnd cell_6t
Xbit_r235_c189 bl[189] br[189] wl[235] vdd gnd cell_6t
Xbit_r236_c189 bl[189] br[189] wl[236] vdd gnd cell_6t
Xbit_r237_c189 bl[189] br[189] wl[237] vdd gnd cell_6t
Xbit_r238_c189 bl[189] br[189] wl[238] vdd gnd cell_6t
Xbit_r239_c189 bl[189] br[189] wl[239] vdd gnd cell_6t
Xbit_r240_c189 bl[189] br[189] wl[240] vdd gnd cell_6t
Xbit_r241_c189 bl[189] br[189] wl[241] vdd gnd cell_6t
Xbit_r242_c189 bl[189] br[189] wl[242] vdd gnd cell_6t
Xbit_r243_c189 bl[189] br[189] wl[243] vdd gnd cell_6t
Xbit_r244_c189 bl[189] br[189] wl[244] vdd gnd cell_6t
Xbit_r245_c189 bl[189] br[189] wl[245] vdd gnd cell_6t
Xbit_r246_c189 bl[189] br[189] wl[246] vdd gnd cell_6t
Xbit_r247_c189 bl[189] br[189] wl[247] vdd gnd cell_6t
Xbit_r248_c189 bl[189] br[189] wl[248] vdd gnd cell_6t
Xbit_r249_c189 bl[189] br[189] wl[249] vdd gnd cell_6t
Xbit_r250_c189 bl[189] br[189] wl[250] vdd gnd cell_6t
Xbit_r251_c189 bl[189] br[189] wl[251] vdd gnd cell_6t
Xbit_r252_c189 bl[189] br[189] wl[252] vdd gnd cell_6t
Xbit_r253_c189 bl[189] br[189] wl[253] vdd gnd cell_6t
Xbit_r254_c189 bl[189] br[189] wl[254] vdd gnd cell_6t
Xbit_r255_c189 bl[189] br[189] wl[255] vdd gnd cell_6t
Xbit_r0_c190 bl[190] br[190] wl[0] vdd gnd cell_6t
Xbit_r1_c190 bl[190] br[190] wl[1] vdd gnd cell_6t
Xbit_r2_c190 bl[190] br[190] wl[2] vdd gnd cell_6t
Xbit_r3_c190 bl[190] br[190] wl[3] vdd gnd cell_6t
Xbit_r4_c190 bl[190] br[190] wl[4] vdd gnd cell_6t
Xbit_r5_c190 bl[190] br[190] wl[5] vdd gnd cell_6t
Xbit_r6_c190 bl[190] br[190] wl[6] vdd gnd cell_6t
Xbit_r7_c190 bl[190] br[190] wl[7] vdd gnd cell_6t
Xbit_r8_c190 bl[190] br[190] wl[8] vdd gnd cell_6t
Xbit_r9_c190 bl[190] br[190] wl[9] vdd gnd cell_6t
Xbit_r10_c190 bl[190] br[190] wl[10] vdd gnd cell_6t
Xbit_r11_c190 bl[190] br[190] wl[11] vdd gnd cell_6t
Xbit_r12_c190 bl[190] br[190] wl[12] vdd gnd cell_6t
Xbit_r13_c190 bl[190] br[190] wl[13] vdd gnd cell_6t
Xbit_r14_c190 bl[190] br[190] wl[14] vdd gnd cell_6t
Xbit_r15_c190 bl[190] br[190] wl[15] vdd gnd cell_6t
Xbit_r16_c190 bl[190] br[190] wl[16] vdd gnd cell_6t
Xbit_r17_c190 bl[190] br[190] wl[17] vdd gnd cell_6t
Xbit_r18_c190 bl[190] br[190] wl[18] vdd gnd cell_6t
Xbit_r19_c190 bl[190] br[190] wl[19] vdd gnd cell_6t
Xbit_r20_c190 bl[190] br[190] wl[20] vdd gnd cell_6t
Xbit_r21_c190 bl[190] br[190] wl[21] vdd gnd cell_6t
Xbit_r22_c190 bl[190] br[190] wl[22] vdd gnd cell_6t
Xbit_r23_c190 bl[190] br[190] wl[23] vdd gnd cell_6t
Xbit_r24_c190 bl[190] br[190] wl[24] vdd gnd cell_6t
Xbit_r25_c190 bl[190] br[190] wl[25] vdd gnd cell_6t
Xbit_r26_c190 bl[190] br[190] wl[26] vdd gnd cell_6t
Xbit_r27_c190 bl[190] br[190] wl[27] vdd gnd cell_6t
Xbit_r28_c190 bl[190] br[190] wl[28] vdd gnd cell_6t
Xbit_r29_c190 bl[190] br[190] wl[29] vdd gnd cell_6t
Xbit_r30_c190 bl[190] br[190] wl[30] vdd gnd cell_6t
Xbit_r31_c190 bl[190] br[190] wl[31] vdd gnd cell_6t
Xbit_r32_c190 bl[190] br[190] wl[32] vdd gnd cell_6t
Xbit_r33_c190 bl[190] br[190] wl[33] vdd gnd cell_6t
Xbit_r34_c190 bl[190] br[190] wl[34] vdd gnd cell_6t
Xbit_r35_c190 bl[190] br[190] wl[35] vdd gnd cell_6t
Xbit_r36_c190 bl[190] br[190] wl[36] vdd gnd cell_6t
Xbit_r37_c190 bl[190] br[190] wl[37] vdd gnd cell_6t
Xbit_r38_c190 bl[190] br[190] wl[38] vdd gnd cell_6t
Xbit_r39_c190 bl[190] br[190] wl[39] vdd gnd cell_6t
Xbit_r40_c190 bl[190] br[190] wl[40] vdd gnd cell_6t
Xbit_r41_c190 bl[190] br[190] wl[41] vdd gnd cell_6t
Xbit_r42_c190 bl[190] br[190] wl[42] vdd gnd cell_6t
Xbit_r43_c190 bl[190] br[190] wl[43] vdd gnd cell_6t
Xbit_r44_c190 bl[190] br[190] wl[44] vdd gnd cell_6t
Xbit_r45_c190 bl[190] br[190] wl[45] vdd gnd cell_6t
Xbit_r46_c190 bl[190] br[190] wl[46] vdd gnd cell_6t
Xbit_r47_c190 bl[190] br[190] wl[47] vdd gnd cell_6t
Xbit_r48_c190 bl[190] br[190] wl[48] vdd gnd cell_6t
Xbit_r49_c190 bl[190] br[190] wl[49] vdd gnd cell_6t
Xbit_r50_c190 bl[190] br[190] wl[50] vdd gnd cell_6t
Xbit_r51_c190 bl[190] br[190] wl[51] vdd gnd cell_6t
Xbit_r52_c190 bl[190] br[190] wl[52] vdd gnd cell_6t
Xbit_r53_c190 bl[190] br[190] wl[53] vdd gnd cell_6t
Xbit_r54_c190 bl[190] br[190] wl[54] vdd gnd cell_6t
Xbit_r55_c190 bl[190] br[190] wl[55] vdd gnd cell_6t
Xbit_r56_c190 bl[190] br[190] wl[56] vdd gnd cell_6t
Xbit_r57_c190 bl[190] br[190] wl[57] vdd gnd cell_6t
Xbit_r58_c190 bl[190] br[190] wl[58] vdd gnd cell_6t
Xbit_r59_c190 bl[190] br[190] wl[59] vdd gnd cell_6t
Xbit_r60_c190 bl[190] br[190] wl[60] vdd gnd cell_6t
Xbit_r61_c190 bl[190] br[190] wl[61] vdd gnd cell_6t
Xbit_r62_c190 bl[190] br[190] wl[62] vdd gnd cell_6t
Xbit_r63_c190 bl[190] br[190] wl[63] vdd gnd cell_6t
Xbit_r64_c190 bl[190] br[190] wl[64] vdd gnd cell_6t
Xbit_r65_c190 bl[190] br[190] wl[65] vdd gnd cell_6t
Xbit_r66_c190 bl[190] br[190] wl[66] vdd gnd cell_6t
Xbit_r67_c190 bl[190] br[190] wl[67] vdd gnd cell_6t
Xbit_r68_c190 bl[190] br[190] wl[68] vdd gnd cell_6t
Xbit_r69_c190 bl[190] br[190] wl[69] vdd gnd cell_6t
Xbit_r70_c190 bl[190] br[190] wl[70] vdd gnd cell_6t
Xbit_r71_c190 bl[190] br[190] wl[71] vdd gnd cell_6t
Xbit_r72_c190 bl[190] br[190] wl[72] vdd gnd cell_6t
Xbit_r73_c190 bl[190] br[190] wl[73] vdd gnd cell_6t
Xbit_r74_c190 bl[190] br[190] wl[74] vdd gnd cell_6t
Xbit_r75_c190 bl[190] br[190] wl[75] vdd gnd cell_6t
Xbit_r76_c190 bl[190] br[190] wl[76] vdd gnd cell_6t
Xbit_r77_c190 bl[190] br[190] wl[77] vdd gnd cell_6t
Xbit_r78_c190 bl[190] br[190] wl[78] vdd gnd cell_6t
Xbit_r79_c190 bl[190] br[190] wl[79] vdd gnd cell_6t
Xbit_r80_c190 bl[190] br[190] wl[80] vdd gnd cell_6t
Xbit_r81_c190 bl[190] br[190] wl[81] vdd gnd cell_6t
Xbit_r82_c190 bl[190] br[190] wl[82] vdd gnd cell_6t
Xbit_r83_c190 bl[190] br[190] wl[83] vdd gnd cell_6t
Xbit_r84_c190 bl[190] br[190] wl[84] vdd gnd cell_6t
Xbit_r85_c190 bl[190] br[190] wl[85] vdd gnd cell_6t
Xbit_r86_c190 bl[190] br[190] wl[86] vdd gnd cell_6t
Xbit_r87_c190 bl[190] br[190] wl[87] vdd gnd cell_6t
Xbit_r88_c190 bl[190] br[190] wl[88] vdd gnd cell_6t
Xbit_r89_c190 bl[190] br[190] wl[89] vdd gnd cell_6t
Xbit_r90_c190 bl[190] br[190] wl[90] vdd gnd cell_6t
Xbit_r91_c190 bl[190] br[190] wl[91] vdd gnd cell_6t
Xbit_r92_c190 bl[190] br[190] wl[92] vdd gnd cell_6t
Xbit_r93_c190 bl[190] br[190] wl[93] vdd gnd cell_6t
Xbit_r94_c190 bl[190] br[190] wl[94] vdd gnd cell_6t
Xbit_r95_c190 bl[190] br[190] wl[95] vdd gnd cell_6t
Xbit_r96_c190 bl[190] br[190] wl[96] vdd gnd cell_6t
Xbit_r97_c190 bl[190] br[190] wl[97] vdd gnd cell_6t
Xbit_r98_c190 bl[190] br[190] wl[98] vdd gnd cell_6t
Xbit_r99_c190 bl[190] br[190] wl[99] vdd gnd cell_6t
Xbit_r100_c190 bl[190] br[190] wl[100] vdd gnd cell_6t
Xbit_r101_c190 bl[190] br[190] wl[101] vdd gnd cell_6t
Xbit_r102_c190 bl[190] br[190] wl[102] vdd gnd cell_6t
Xbit_r103_c190 bl[190] br[190] wl[103] vdd gnd cell_6t
Xbit_r104_c190 bl[190] br[190] wl[104] vdd gnd cell_6t
Xbit_r105_c190 bl[190] br[190] wl[105] vdd gnd cell_6t
Xbit_r106_c190 bl[190] br[190] wl[106] vdd gnd cell_6t
Xbit_r107_c190 bl[190] br[190] wl[107] vdd gnd cell_6t
Xbit_r108_c190 bl[190] br[190] wl[108] vdd gnd cell_6t
Xbit_r109_c190 bl[190] br[190] wl[109] vdd gnd cell_6t
Xbit_r110_c190 bl[190] br[190] wl[110] vdd gnd cell_6t
Xbit_r111_c190 bl[190] br[190] wl[111] vdd gnd cell_6t
Xbit_r112_c190 bl[190] br[190] wl[112] vdd gnd cell_6t
Xbit_r113_c190 bl[190] br[190] wl[113] vdd gnd cell_6t
Xbit_r114_c190 bl[190] br[190] wl[114] vdd gnd cell_6t
Xbit_r115_c190 bl[190] br[190] wl[115] vdd gnd cell_6t
Xbit_r116_c190 bl[190] br[190] wl[116] vdd gnd cell_6t
Xbit_r117_c190 bl[190] br[190] wl[117] vdd gnd cell_6t
Xbit_r118_c190 bl[190] br[190] wl[118] vdd gnd cell_6t
Xbit_r119_c190 bl[190] br[190] wl[119] vdd gnd cell_6t
Xbit_r120_c190 bl[190] br[190] wl[120] vdd gnd cell_6t
Xbit_r121_c190 bl[190] br[190] wl[121] vdd gnd cell_6t
Xbit_r122_c190 bl[190] br[190] wl[122] vdd gnd cell_6t
Xbit_r123_c190 bl[190] br[190] wl[123] vdd gnd cell_6t
Xbit_r124_c190 bl[190] br[190] wl[124] vdd gnd cell_6t
Xbit_r125_c190 bl[190] br[190] wl[125] vdd gnd cell_6t
Xbit_r126_c190 bl[190] br[190] wl[126] vdd gnd cell_6t
Xbit_r127_c190 bl[190] br[190] wl[127] vdd gnd cell_6t
Xbit_r128_c190 bl[190] br[190] wl[128] vdd gnd cell_6t
Xbit_r129_c190 bl[190] br[190] wl[129] vdd gnd cell_6t
Xbit_r130_c190 bl[190] br[190] wl[130] vdd gnd cell_6t
Xbit_r131_c190 bl[190] br[190] wl[131] vdd gnd cell_6t
Xbit_r132_c190 bl[190] br[190] wl[132] vdd gnd cell_6t
Xbit_r133_c190 bl[190] br[190] wl[133] vdd gnd cell_6t
Xbit_r134_c190 bl[190] br[190] wl[134] vdd gnd cell_6t
Xbit_r135_c190 bl[190] br[190] wl[135] vdd gnd cell_6t
Xbit_r136_c190 bl[190] br[190] wl[136] vdd gnd cell_6t
Xbit_r137_c190 bl[190] br[190] wl[137] vdd gnd cell_6t
Xbit_r138_c190 bl[190] br[190] wl[138] vdd gnd cell_6t
Xbit_r139_c190 bl[190] br[190] wl[139] vdd gnd cell_6t
Xbit_r140_c190 bl[190] br[190] wl[140] vdd gnd cell_6t
Xbit_r141_c190 bl[190] br[190] wl[141] vdd gnd cell_6t
Xbit_r142_c190 bl[190] br[190] wl[142] vdd gnd cell_6t
Xbit_r143_c190 bl[190] br[190] wl[143] vdd gnd cell_6t
Xbit_r144_c190 bl[190] br[190] wl[144] vdd gnd cell_6t
Xbit_r145_c190 bl[190] br[190] wl[145] vdd gnd cell_6t
Xbit_r146_c190 bl[190] br[190] wl[146] vdd gnd cell_6t
Xbit_r147_c190 bl[190] br[190] wl[147] vdd gnd cell_6t
Xbit_r148_c190 bl[190] br[190] wl[148] vdd gnd cell_6t
Xbit_r149_c190 bl[190] br[190] wl[149] vdd gnd cell_6t
Xbit_r150_c190 bl[190] br[190] wl[150] vdd gnd cell_6t
Xbit_r151_c190 bl[190] br[190] wl[151] vdd gnd cell_6t
Xbit_r152_c190 bl[190] br[190] wl[152] vdd gnd cell_6t
Xbit_r153_c190 bl[190] br[190] wl[153] vdd gnd cell_6t
Xbit_r154_c190 bl[190] br[190] wl[154] vdd gnd cell_6t
Xbit_r155_c190 bl[190] br[190] wl[155] vdd gnd cell_6t
Xbit_r156_c190 bl[190] br[190] wl[156] vdd gnd cell_6t
Xbit_r157_c190 bl[190] br[190] wl[157] vdd gnd cell_6t
Xbit_r158_c190 bl[190] br[190] wl[158] vdd gnd cell_6t
Xbit_r159_c190 bl[190] br[190] wl[159] vdd gnd cell_6t
Xbit_r160_c190 bl[190] br[190] wl[160] vdd gnd cell_6t
Xbit_r161_c190 bl[190] br[190] wl[161] vdd gnd cell_6t
Xbit_r162_c190 bl[190] br[190] wl[162] vdd gnd cell_6t
Xbit_r163_c190 bl[190] br[190] wl[163] vdd gnd cell_6t
Xbit_r164_c190 bl[190] br[190] wl[164] vdd gnd cell_6t
Xbit_r165_c190 bl[190] br[190] wl[165] vdd gnd cell_6t
Xbit_r166_c190 bl[190] br[190] wl[166] vdd gnd cell_6t
Xbit_r167_c190 bl[190] br[190] wl[167] vdd gnd cell_6t
Xbit_r168_c190 bl[190] br[190] wl[168] vdd gnd cell_6t
Xbit_r169_c190 bl[190] br[190] wl[169] vdd gnd cell_6t
Xbit_r170_c190 bl[190] br[190] wl[170] vdd gnd cell_6t
Xbit_r171_c190 bl[190] br[190] wl[171] vdd gnd cell_6t
Xbit_r172_c190 bl[190] br[190] wl[172] vdd gnd cell_6t
Xbit_r173_c190 bl[190] br[190] wl[173] vdd gnd cell_6t
Xbit_r174_c190 bl[190] br[190] wl[174] vdd gnd cell_6t
Xbit_r175_c190 bl[190] br[190] wl[175] vdd gnd cell_6t
Xbit_r176_c190 bl[190] br[190] wl[176] vdd gnd cell_6t
Xbit_r177_c190 bl[190] br[190] wl[177] vdd gnd cell_6t
Xbit_r178_c190 bl[190] br[190] wl[178] vdd gnd cell_6t
Xbit_r179_c190 bl[190] br[190] wl[179] vdd gnd cell_6t
Xbit_r180_c190 bl[190] br[190] wl[180] vdd gnd cell_6t
Xbit_r181_c190 bl[190] br[190] wl[181] vdd gnd cell_6t
Xbit_r182_c190 bl[190] br[190] wl[182] vdd gnd cell_6t
Xbit_r183_c190 bl[190] br[190] wl[183] vdd gnd cell_6t
Xbit_r184_c190 bl[190] br[190] wl[184] vdd gnd cell_6t
Xbit_r185_c190 bl[190] br[190] wl[185] vdd gnd cell_6t
Xbit_r186_c190 bl[190] br[190] wl[186] vdd gnd cell_6t
Xbit_r187_c190 bl[190] br[190] wl[187] vdd gnd cell_6t
Xbit_r188_c190 bl[190] br[190] wl[188] vdd gnd cell_6t
Xbit_r189_c190 bl[190] br[190] wl[189] vdd gnd cell_6t
Xbit_r190_c190 bl[190] br[190] wl[190] vdd gnd cell_6t
Xbit_r191_c190 bl[190] br[190] wl[191] vdd gnd cell_6t
Xbit_r192_c190 bl[190] br[190] wl[192] vdd gnd cell_6t
Xbit_r193_c190 bl[190] br[190] wl[193] vdd gnd cell_6t
Xbit_r194_c190 bl[190] br[190] wl[194] vdd gnd cell_6t
Xbit_r195_c190 bl[190] br[190] wl[195] vdd gnd cell_6t
Xbit_r196_c190 bl[190] br[190] wl[196] vdd gnd cell_6t
Xbit_r197_c190 bl[190] br[190] wl[197] vdd gnd cell_6t
Xbit_r198_c190 bl[190] br[190] wl[198] vdd gnd cell_6t
Xbit_r199_c190 bl[190] br[190] wl[199] vdd gnd cell_6t
Xbit_r200_c190 bl[190] br[190] wl[200] vdd gnd cell_6t
Xbit_r201_c190 bl[190] br[190] wl[201] vdd gnd cell_6t
Xbit_r202_c190 bl[190] br[190] wl[202] vdd gnd cell_6t
Xbit_r203_c190 bl[190] br[190] wl[203] vdd gnd cell_6t
Xbit_r204_c190 bl[190] br[190] wl[204] vdd gnd cell_6t
Xbit_r205_c190 bl[190] br[190] wl[205] vdd gnd cell_6t
Xbit_r206_c190 bl[190] br[190] wl[206] vdd gnd cell_6t
Xbit_r207_c190 bl[190] br[190] wl[207] vdd gnd cell_6t
Xbit_r208_c190 bl[190] br[190] wl[208] vdd gnd cell_6t
Xbit_r209_c190 bl[190] br[190] wl[209] vdd gnd cell_6t
Xbit_r210_c190 bl[190] br[190] wl[210] vdd gnd cell_6t
Xbit_r211_c190 bl[190] br[190] wl[211] vdd gnd cell_6t
Xbit_r212_c190 bl[190] br[190] wl[212] vdd gnd cell_6t
Xbit_r213_c190 bl[190] br[190] wl[213] vdd gnd cell_6t
Xbit_r214_c190 bl[190] br[190] wl[214] vdd gnd cell_6t
Xbit_r215_c190 bl[190] br[190] wl[215] vdd gnd cell_6t
Xbit_r216_c190 bl[190] br[190] wl[216] vdd gnd cell_6t
Xbit_r217_c190 bl[190] br[190] wl[217] vdd gnd cell_6t
Xbit_r218_c190 bl[190] br[190] wl[218] vdd gnd cell_6t
Xbit_r219_c190 bl[190] br[190] wl[219] vdd gnd cell_6t
Xbit_r220_c190 bl[190] br[190] wl[220] vdd gnd cell_6t
Xbit_r221_c190 bl[190] br[190] wl[221] vdd gnd cell_6t
Xbit_r222_c190 bl[190] br[190] wl[222] vdd gnd cell_6t
Xbit_r223_c190 bl[190] br[190] wl[223] vdd gnd cell_6t
Xbit_r224_c190 bl[190] br[190] wl[224] vdd gnd cell_6t
Xbit_r225_c190 bl[190] br[190] wl[225] vdd gnd cell_6t
Xbit_r226_c190 bl[190] br[190] wl[226] vdd gnd cell_6t
Xbit_r227_c190 bl[190] br[190] wl[227] vdd gnd cell_6t
Xbit_r228_c190 bl[190] br[190] wl[228] vdd gnd cell_6t
Xbit_r229_c190 bl[190] br[190] wl[229] vdd gnd cell_6t
Xbit_r230_c190 bl[190] br[190] wl[230] vdd gnd cell_6t
Xbit_r231_c190 bl[190] br[190] wl[231] vdd gnd cell_6t
Xbit_r232_c190 bl[190] br[190] wl[232] vdd gnd cell_6t
Xbit_r233_c190 bl[190] br[190] wl[233] vdd gnd cell_6t
Xbit_r234_c190 bl[190] br[190] wl[234] vdd gnd cell_6t
Xbit_r235_c190 bl[190] br[190] wl[235] vdd gnd cell_6t
Xbit_r236_c190 bl[190] br[190] wl[236] vdd gnd cell_6t
Xbit_r237_c190 bl[190] br[190] wl[237] vdd gnd cell_6t
Xbit_r238_c190 bl[190] br[190] wl[238] vdd gnd cell_6t
Xbit_r239_c190 bl[190] br[190] wl[239] vdd gnd cell_6t
Xbit_r240_c190 bl[190] br[190] wl[240] vdd gnd cell_6t
Xbit_r241_c190 bl[190] br[190] wl[241] vdd gnd cell_6t
Xbit_r242_c190 bl[190] br[190] wl[242] vdd gnd cell_6t
Xbit_r243_c190 bl[190] br[190] wl[243] vdd gnd cell_6t
Xbit_r244_c190 bl[190] br[190] wl[244] vdd gnd cell_6t
Xbit_r245_c190 bl[190] br[190] wl[245] vdd gnd cell_6t
Xbit_r246_c190 bl[190] br[190] wl[246] vdd gnd cell_6t
Xbit_r247_c190 bl[190] br[190] wl[247] vdd gnd cell_6t
Xbit_r248_c190 bl[190] br[190] wl[248] vdd gnd cell_6t
Xbit_r249_c190 bl[190] br[190] wl[249] vdd gnd cell_6t
Xbit_r250_c190 bl[190] br[190] wl[250] vdd gnd cell_6t
Xbit_r251_c190 bl[190] br[190] wl[251] vdd gnd cell_6t
Xbit_r252_c190 bl[190] br[190] wl[252] vdd gnd cell_6t
Xbit_r253_c190 bl[190] br[190] wl[253] vdd gnd cell_6t
Xbit_r254_c190 bl[190] br[190] wl[254] vdd gnd cell_6t
Xbit_r255_c190 bl[190] br[190] wl[255] vdd gnd cell_6t
Xbit_r0_c191 bl[191] br[191] wl[0] vdd gnd cell_6t
Xbit_r1_c191 bl[191] br[191] wl[1] vdd gnd cell_6t
Xbit_r2_c191 bl[191] br[191] wl[2] vdd gnd cell_6t
Xbit_r3_c191 bl[191] br[191] wl[3] vdd gnd cell_6t
Xbit_r4_c191 bl[191] br[191] wl[4] vdd gnd cell_6t
Xbit_r5_c191 bl[191] br[191] wl[5] vdd gnd cell_6t
Xbit_r6_c191 bl[191] br[191] wl[6] vdd gnd cell_6t
Xbit_r7_c191 bl[191] br[191] wl[7] vdd gnd cell_6t
Xbit_r8_c191 bl[191] br[191] wl[8] vdd gnd cell_6t
Xbit_r9_c191 bl[191] br[191] wl[9] vdd gnd cell_6t
Xbit_r10_c191 bl[191] br[191] wl[10] vdd gnd cell_6t
Xbit_r11_c191 bl[191] br[191] wl[11] vdd gnd cell_6t
Xbit_r12_c191 bl[191] br[191] wl[12] vdd gnd cell_6t
Xbit_r13_c191 bl[191] br[191] wl[13] vdd gnd cell_6t
Xbit_r14_c191 bl[191] br[191] wl[14] vdd gnd cell_6t
Xbit_r15_c191 bl[191] br[191] wl[15] vdd gnd cell_6t
Xbit_r16_c191 bl[191] br[191] wl[16] vdd gnd cell_6t
Xbit_r17_c191 bl[191] br[191] wl[17] vdd gnd cell_6t
Xbit_r18_c191 bl[191] br[191] wl[18] vdd gnd cell_6t
Xbit_r19_c191 bl[191] br[191] wl[19] vdd gnd cell_6t
Xbit_r20_c191 bl[191] br[191] wl[20] vdd gnd cell_6t
Xbit_r21_c191 bl[191] br[191] wl[21] vdd gnd cell_6t
Xbit_r22_c191 bl[191] br[191] wl[22] vdd gnd cell_6t
Xbit_r23_c191 bl[191] br[191] wl[23] vdd gnd cell_6t
Xbit_r24_c191 bl[191] br[191] wl[24] vdd gnd cell_6t
Xbit_r25_c191 bl[191] br[191] wl[25] vdd gnd cell_6t
Xbit_r26_c191 bl[191] br[191] wl[26] vdd gnd cell_6t
Xbit_r27_c191 bl[191] br[191] wl[27] vdd gnd cell_6t
Xbit_r28_c191 bl[191] br[191] wl[28] vdd gnd cell_6t
Xbit_r29_c191 bl[191] br[191] wl[29] vdd gnd cell_6t
Xbit_r30_c191 bl[191] br[191] wl[30] vdd gnd cell_6t
Xbit_r31_c191 bl[191] br[191] wl[31] vdd gnd cell_6t
Xbit_r32_c191 bl[191] br[191] wl[32] vdd gnd cell_6t
Xbit_r33_c191 bl[191] br[191] wl[33] vdd gnd cell_6t
Xbit_r34_c191 bl[191] br[191] wl[34] vdd gnd cell_6t
Xbit_r35_c191 bl[191] br[191] wl[35] vdd gnd cell_6t
Xbit_r36_c191 bl[191] br[191] wl[36] vdd gnd cell_6t
Xbit_r37_c191 bl[191] br[191] wl[37] vdd gnd cell_6t
Xbit_r38_c191 bl[191] br[191] wl[38] vdd gnd cell_6t
Xbit_r39_c191 bl[191] br[191] wl[39] vdd gnd cell_6t
Xbit_r40_c191 bl[191] br[191] wl[40] vdd gnd cell_6t
Xbit_r41_c191 bl[191] br[191] wl[41] vdd gnd cell_6t
Xbit_r42_c191 bl[191] br[191] wl[42] vdd gnd cell_6t
Xbit_r43_c191 bl[191] br[191] wl[43] vdd gnd cell_6t
Xbit_r44_c191 bl[191] br[191] wl[44] vdd gnd cell_6t
Xbit_r45_c191 bl[191] br[191] wl[45] vdd gnd cell_6t
Xbit_r46_c191 bl[191] br[191] wl[46] vdd gnd cell_6t
Xbit_r47_c191 bl[191] br[191] wl[47] vdd gnd cell_6t
Xbit_r48_c191 bl[191] br[191] wl[48] vdd gnd cell_6t
Xbit_r49_c191 bl[191] br[191] wl[49] vdd gnd cell_6t
Xbit_r50_c191 bl[191] br[191] wl[50] vdd gnd cell_6t
Xbit_r51_c191 bl[191] br[191] wl[51] vdd gnd cell_6t
Xbit_r52_c191 bl[191] br[191] wl[52] vdd gnd cell_6t
Xbit_r53_c191 bl[191] br[191] wl[53] vdd gnd cell_6t
Xbit_r54_c191 bl[191] br[191] wl[54] vdd gnd cell_6t
Xbit_r55_c191 bl[191] br[191] wl[55] vdd gnd cell_6t
Xbit_r56_c191 bl[191] br[191] wl[56] vdd gnd cell_6t
Xbit_r57_c191 bl[191] br[191] wl[57] vdd gnd cell_6t
Xbit_r58_c191 bl[191] br[191] wl[58] vdd gnd cell_6t
Xbit_r59_c191 bl[191] br[191] wl[59] vdd gnd cell_6t
Xbit_r60_c191 bl[191] br[191] wl[60] vdd gnd cell_6t
Xbit_r61_c191 bl[191] br[191] wl[61] vdd gnd cell_6t
Xbit_r62_c191 bl[191] br[191] wl[62] vdd gnd cell_6t
Xbit_r63_c191 bl[191] br[191] wl[63] vdd gnd cell_6t
Xbit_r64_c191 bl[191] br[191] wl[64] vdd gnd cell_6t
Xbit_r65_c191 bl[191] br[191] wl[65] vdd gnd cell_6t
Xbit_r66_c191 bl[191] br[191] wl[66] vdd gnd cell_6t
Xbit_r67_c191 bl[191] br[191] wl[67] vdd gnd cell_6t
Xbit_r68_c191 bl[191] br[191] wl[68] vdd gnd cell_6t
Xbit_r69_c191 bl[191] br[191] wl[69] vdd gnd cell_6t
Xbit_r70_c191 bl[191] br[191] wl[70] vdd gnd cell_6t
Xbit_r71_c191 bl[191] br[191] wl[71] vdd gnd cell_6t
Xbit_r72_c191 bl[191] br[191] wl[72] vdd gnd cell_6t
Xbit_r73_c191 bl[191] br[191] wl[73] vdd gnd cell_6t
Xbit_r74_c191 bl[191] br[191] wl[74] vdd gnd cell_6t
Xbit_r75_c191 bl[191] br[191] wl[75] vdd gnd cell_6t
Xbit_r76_c191 bl[191] br[191] wl[76] vdd gnd cell_6t
Xbit_r77_c191 bl[191] br[191] wl[77] vdd gnd cell_6t
Xbit_r78_c191 bl[191] br[191] wl[78] vdd gnd cell_6t
Xbit_r79_c191 bl[191] br[191] wl[79] vdd gnd cell_6t
Xbit_r80_c191 bl[191] br[191] wl[80] vdd gnd cell_6t
Xbit_r81_c191 bl[191] br[191] wl[81] vdd gnd cell_6t
Xbit_r82_c191 bl[191] br[191] wl[82] vdd gnd cell_6t
Xbit_r83_c191 bl[191] br[191] wl[83] vdd gnd cell_6t
Xbit_r84_c191 bl[191] br[191] wl[84] vdd gnd cell_6t
Xbit_r85_c191 bl[191] br[191] wl[85] vdd gnd cell_6t
Xbit_r86_c191 bl[191] br[191] wl[86] vdd gnd cell_6t
Xbit_r87_c191 bl[191] br[191] wl[87] vdd gnd cell_6t
Xbit_r88_c191 bl[191] br[191] wl[88] vdd gnd cell_6t
Xbit_r89_c191 bl[191] br[191] wl[89] vdd gnd cell_6t
Xbit_r90_c191 bl[191] br[191] wl[90] vdd gnd cell_6t
Xbit_r91_c191 bl[191] br[191] wl[91] vdd gnd cell_6t
Xbit_r92_c191 bl[191] br[191] wl[92] vdd gnd cell_6t
Xbit_r93_c191 bl[191] br[191] wl[93] vdd gnd cell_6t
Xbit_r94_c191 bl[191] br[191] wl[94] vdd gnd cell_6t
Xbit_r95_c191 bl[191] br[191] wl[95] vdd gnd cell_6t
Xbit_r96_c191 bl[191] br[191] wl[96] vdd gnd cell_6t
Xbit_r97_c191 bl[191] br[191] wl[97] vdd gnd cell_6t
Xbit_r98_c191 bl[191] br[191] wl[98] vdd gnd cell_6t
Xbit_r99_c191 bl[191] br[191] wl[99] vdd gnd cell_6t
Xbit_r100_c191 bl[191] br[191] wl[100] vdd gnd cell_6t
Xbit_r101_c191 bl[191] br[191] wl[101] vdd gnd cell_6t
Xbit_r102_c191 bl[191] br[191] wl[102] vdd gnd cell_6t
Xbit_r103_c191 bl[191] br[191] wl[103] vdd gnd cell_6t
Xbit_r104_c191 bl[191] br[191] wl[104] vdd gnd cell_6t
Xbit_r105_c191 bl[191] br[191] wl[105] vdd gnd cell_6t
Xbit_r106_c191 bl[191] br[191] wl[106] vdd gnd cell_6t
Xbit_r107_c191 bl[191] br[191] wl[107] vdd gnd cell_6t
Xbit_r108_c191 bl[191] br[191] wl[108] vdd gnd cell_6t
Xbit_r109_c191 bl[191] br[191] wl[109] vdd gnd cell_6t
Xbit_r110_c191 bl[191] br[191] wl[110] vdd gnd cell_6t
Xbit_r111_c191 bl[191] br[191] wl[111] vdd gnd cell_6t
Xbit_r112_c191 bl[191] br[191] wl[112] vdd gnd cell_6t
Xbit_r113_c191 bl[191] br[191] wl[113] vdd gnd cell_6t
Xbit_r114_c191 bl[191] br[191] wl[114] vdd gnd cell_6t
Xbit_r115_c191 bl[191] br[191] wl[115] vdd gnd cell_6t
Xbit_r116_c191 bl[191] br[191] wl[116] vdd gnd cell_6t
Xbit_r117_c191 bl[191] br[191] wl[117] vdd gnd cell_6t
Xbit_r118_c191 bl[191] br[191] wl[118] vdd gnd cell_6t
Xbit_r119_c191 bl[191] br[191] wl[119] vdd gnd cell_6t
Xbit_r120_c191 bl[191] br[191] wl[120] vdd gnd cell_6t
Xbit_r121_c191 bl[191] br[191] wl[121] vdd gnd cell_6t
Xbit_r122_c191 bl[191] br[191] wl[122] vdd gnd cell_6t
Xbit_r123_c191 bl[191] br[191] wl[123] vdd gnd cell_6t
Xbit_r124_c191 bl[191] br[191] wl[124] vdd gnd cell_6t
Xbit_r125_c191 bl[191] br[191] wl[125] vdd gnd cell_6t
Xbit_r126_c191 bl[191] br[191] wl[126] vdd gnd cell_6t
Xbit_r127_c191 bl[191] br[191] wl[127] vdd gnd cell_6t
Xbit_r128_c191 bl[191] br[191] wl[128] vdd gnd cell_6t
Xbit_r129_c191 bl[191] br[191] wl[129] vdd gnd cell_6t
Xbit_r130_c191 bl[191] br[191] wl[130] vdd gnd cell_6t
Xbit_r131_c191 bl[191] br[191] wl[131] vdd gnd cell_6t
Xbit_r132_c191 bl[191] br[191] wl[132] vdd gnd cell_6t
Xbit_r133_c191 bl[191] br[191] wl[133] vdd gnd cell_6t
Xbit_r134_c191 bl[191] br[191] wl[134] vdd gnd cell_6t
Xbit_r135_c191 bl[191] br[191] wl[135] vdd gnd cell_6t
Xbit_r136_c191 bl[191] br[191] wl[136] vdd gnd cell_6t
Xbit_r137_c191 bl[191] br[191] wl[137] vdd gnd cell_6t
Xbit_r138_c191 bl[191] br[191] wl[138] vdd gnd cell_6t
Xbit_r139_c191 bl[191] br[191] wl[139] vdd gnd cell_6t
Xbit_r140_c191 bl[191] br[191] wl[140] vdd gnd cell_6t
Xbit_r141_c191 bl[191] br[191] wl[141] vdd gnd cell_6t
Xbit_r142_c191 bl[191] br[191] wl[142] vdd gnd cell_6t
Xbit_r143_c191 bl[191] br[191] wl[143] vdd gnd cell_6t
Xbit_r144_c191 bl[191] br[191] wl[144] vdd gnd cell_6t
Xbit_r145_c191 bl[191] br[191] wl[145] vdd gnd cell_6t
Xbit_r146_c191 bl[191] br[191] wl[146] vdd gnd cell_6t
Xbit_r147_c191 bl[191] br[191] wl[147] vdd gnd cell_6t
Xbit_r148_c191 bl[191] br[191] wl[148] vdd gnd cell_6t
Xbit_r149_c191 bl[191] br[191] wl[149] vdd gnd cell_6t
Xbit_r150_c191 bl[191] br[191] wl[150] vdd gnd cell_6t
Xbit_r151_c191 bl[191] br[191] wl[151] vdd gnd cell_6t
Xbit_r152_c191 bl[191] br[191] wl[152] vdd gnd cell_6t
Xbit_r153_c191 bl[191] br[191] wl[153] vdd gnd cell_6t
Xbit_r154_c191 bl[191] br[191] wl[154] vdd gnd cell_6t
Xbit_r155_c191 bl[191] br[191] wl[155] vdd gnd cell_6t
Xbit_r156_c191 bl[191] br[191] wl[156] vdd gnd cell_6t
Xbit_r157_c191 bl[191] br[191] wl[157] vdd gnd cell_6t
Xbit_r158_c191 bl[191] br[191] wl[158] vdd gnd cell_6t
Xbit_r159_c191 bl[191] br[191] wl[159] vdd gnd cell_6t
Xbit_r160_c191 bl[191] br[191] wl[160] vdd gnd cell_6t
Xbit_r161_c191 bl[191] br[191] wl[161] vdd gnd cell_6t
Xbit_r162_c191 bl[191] br[191] wl[162] vdd gnd cell_6t
Xbit_r163_c191 bl[191] br[191] wl[163] vdd gnd cell_6t
Xbit_r164_c191 bl[191] br[191] wl[164] vdd gnd cell_6t
Xbit_r165_c191 bl[191] br[191] wl[165] vdd gnd cell_6t
Xbit_r166_c191 bl[191] br[191] wl[166] vdd gnd cell_6t
Xbit_r167_c191 bl[191] br[191] wl[167] vdd gnd cell_6t
Xbit_r168_c191 bl[191] br[191] wl[168] vdd gnd cell_6t
Xbit_r169_c191 bl[191] br[191] wl[169] vdd gnd cell_6t
Xbit_r170_c191 bl[191] br[191] wl[170] vdd gnd cell_6t
Xbit_r171_c191 bl[191] br[191] wl[171] vdd gnd cell_6t
Xbit_r172_c191 bl[191] br[191] wl[172] vdd gnd cell_6t
Xbit_r173_c191 bl[191] br[191] wl[173] vdd gnd cell_6t
Xbit_r174_c191 bl[191] br[191] wl[174] vdd gnd cell_6t
Xbit_r175_c191 bl[191] br[191] wl[175] vdd gnd cell_6t
Xbit_r176_c191 bl[191] br[191] wl[176] vdd gnd cell_6t
Xbit_r177_c191 bl[191] br[191] wl[177] vdd gnd cell_6t
Xbit_r178_c191 bl[191] br[191] wl[178] vdd gnd cell_6t
Xbit_r179_c191 bl[191] br[191] wl[179] vdd gnd cell_6t
Xbit_r180_c191 bl[191] br[191] wl[180] vdd gnd cell_6t
Xbit_r181_c191 bl[191] br[191] wl[181] vdd gnd cell_6t
Xbit_r182_c191 bl[191] br[191] wl[182] vdd gnd cell_6t
Xbit_r183_c191 bl[191] br[191] wl[183] vdd gnd cell_6t
Xbit_r184_c191 bl[191] br[191] wl[184] vdd gnd cell_6t
Xbit_r185_c191 bl[191] br[191] wl[185] vdd gnd cell_6t
Xbit_r186_c191 bl[191] br[191] wl[186] vdd gnd cell_6t
Xbit_r187_c191 bl[191] br[191] wl[187] vdd gnd cell_6t
Xbit_r188_c191 bl[191] br[191] wl[188] vdd gnd cell_6t
Xbit_r189_c191 bl[191] br[191] wl[189] vdd gnd cell_6t
Xbit_r190_c191 bl[191] br[191] wl[190] vdd gnd cell_6t
Xbit_r191_c191 bl[191] br[191] wl[191] vdd gnd cell_6t
Xbit_r192_c191 bl[191] br[191] wl[192] vdd gnd cell_6t
Xbit_r193_c191 bl[191] br[191] wl[193] vdd gnd cell_6t
Xbit_r194_c191 bl[191] br[191] wl[194] vdd gnd cell_6t
Xbit_r195_c191 bl[191] br[191] wl[195] vdd gnd cell_6t
Xbit_r196_c191 bl[191] br[191] wl[196] vdd gnd cell_6t
Xbit_r197_c191 bl[191] br[191] wl[197] vdd gnd cell_6t
Xbit_r198_c191 bl[191] br[191] wl[198] vdd gnd cell_6t
Xbit_r199_c191 bl[191] br[191] wl[199] vdd gnd cell_6t
Xbit_r200_c191 bl[191] br[191] wl[200] vdd gnd cell_6t
Xbit_r201_c191 bl[191] br[191] wl[201] vdd gnd cell_6t
Xbit_r202_c191 bl[191] br[191] wl[202] vdd gnd cell_6t
Xbit_r203_c191 bl[191] br[191] wl[203] vdd gnd cell_6t
Xbit_r204_c191 bl[191] br[191] wl[204] vdd gnd cell_6t
Xbit_r205_c191 bl[191] br[191] wl[205] vdd gnd cell_6t
Xbit_r206_c191 bl[191] br[191] wl[206] vdd gnd cell_6t
Xbit_r207_c191 bl[191] br[191] wl[207] vdd gnd cell_6t
Xbit_r208_c191 bl[191] br[191] wl[208] vdd gnd cell_6t
Xbit_r209_c191 bl[191] br[191] wl[209] vdd gnd cell_6t
Xbit_r210_c191 bl[191] br[191] wl[210] vdd gnd cell_6t
Xbit_r211_c191 bl[191] br[191] wl[211] vdd gnd cell_6t
Xbit_r212_c191 bl[191] br[191] wl[212] vdd gnd cell_6t
Xbit_r213_c191 bl[191] br[191] wl[213] vdd gnd cell_6t
Xbit_r214_c191 bl[191] br[191] wl[214] vdd gnd cell_6t
Xbit_r215_c191 bl[191] br[191] wl[215] vdd gnd cell_6t
Xbit_r216_c191 bl[191] br[191] wl[216] vdd gnd cell_6t
Xbit_r217_c191 bl[191] br[191] wl[217] vdd gnd cell_6t
Xbit_r218_c191 bl[191] br[191] wl[218] vdd gnd cell_6t
Xbit_r219_c191 bl[191] br[191] wl[219] vdd gnd cell_6t
Xbit_r220_c191 bl[191] br[191] wl[220] vdd gnd cell_6t
Xbit_r221_c191 bl[191] br[191] wl[221] vdd gnd cell_6t
Xbit_r222_c191 bl[191] br[191] wl[222] vdd gnd cell_6t
Xbit_r223_c191 bl[191] br[191] wl[223] vdd gnd cell_6t
Xbit_r224_c191 bl[191] br[191] wl[224] vdd gnd cell_6t
Xbit_r225_c191 bl[191] br[191] wl[225] vdd gnd cell_6t
Xbit_r226_c191 bl[191] br[191] wl[226] vdd gnd cell_6t
Xbit_r227_c191 bl[191] br[191] wl[227] vdd gnd cell_6t
Xbit_r228_c191 bl[191] br[191] wl[228] vdd gnd cell_6t
Xbit_r229_c191 bl[191] br[191] wl[229] vdd gnd cell_6t
Xbit_r230_c191 bl[191] br[191] wl[230] vdd gnd cell_6t
Xbit_r231_c191 bl[191] br[191] wl[231] vdd gnd cell_6t
Xbit_r232_c191 bl[191] br[191] wl[232] vdd gnd cell_6t
Xbit_r233_c191 bl[191] br[191] wl[233] vdd gnd cell_6t
Xbit_r234_c191 bl[191] br[191] wl[234] vdd gnd cell_6t
Xbit_r235_c191 bl[191] br[191] wl[235] vdd gnd cell_6t
Xbit_r236_c191 bl[191] br[191] wl[236] vdd gnd cell_6t
Xbit_r237_c191 bl[191] br[191] wl[237] vdd gnd cell_6t
Xbit_r238_c191 bl[191] br[191] wl[238] vdd gnd cell_6t
Xbit_r239_c191 bl[191] br[191] wl[239] vdd gnd cell_6t
Xbit_r240_c191 bl[191] br[191] wl[240] vdd gnd cell_6t
Xbit_r241_c191 bl[191] br[191] wl[241] vdd gnd cell_6t
Xbit_r242_c191 bl[191] br[191] wl[242] vdd gnd cell_6t
Xbit_r243_c191 bl[191] br[191] wl[243] vdd gnd cell_6t
Xbit_r244_c191 bl[191] br[191] wl[244] vdd gnd cell_6t
Xbit_r245_c191 bl[191] br[191] wl[245] vdd gnd cell_6t
Xbit_r246_c191 bl[191] br[191] wl[246] vdd gnd cell_6t
Xbit_r247_c191 bl[191] br[191] wl[247] vdd gnd cell_6t
Xbit_r248_c191 bl[191] br[191] wl[248] vdd gnd cell_6t
Xbit_r249_c191 bl[191] br[191] wl[249] vdd gnd cell_6t
Xbit_r250_c191 bl[191] br[191] wl[250] vdd gnd cell_6t
Xbit_r251_c191 bl[191] br[191] wl[251] vdd gnd cell_6t
Xbit_r252_c191 bl[191] br[191] wl[252] vdd gnd cell_6t
Xbit_r253_c191 bl[191] br[191] wl[253] vdd gnd cell_6t
Xbit_r254_c191 bl[191] br[191] wl[254] vdd gnd cell_6t
Xbit_r255_c191 bl[191] br[191] wl[255] vdd gnd cell_6t
Xbit_r0_c192 bl[192] br[192] wl[0] vdd gnd cell_6t
Xbit_r1_c192 bl[192] br[192] wl[1] vdd gnd cell_6t
Xbit_r2_c192 bl[192] br[192] wl[2] vdd gnd cell_6t
Xbit_r3_c192 bl[192] br[192] wl[3] vdd gnd cell_6t
Xbit_r4_c192 bl[192] br[192] wl[4] vdd gnd cell_6t
Xbit_r5_c192 bl[192] br[192] wl[5] vdd gnd cell_6t
Xbit_r6_c192 bl[192] br[192] wl[6] vdd gnd cell_6t
Xbit_r7_c192 bl[192] br[192] wl[7] vdd gnd cell_6t
Xbit_r8_c192 bl[192] br[192] wl[8] vdd gnd cell_6t
Xbit_r9_c192 bl[192] br[192] wl[9] vdd gnd cell_6t
Xbit_r10_c192 bl[192] br[192] wl[10] vdd gnd cell_6t
Xbit_r11_c192 bl[192] br[192] wl[11] vdd gnd cell_6t
Xbit_r12_c192 bl[192] br[192] wl[12] vdd gnd cell_6t
Xbit_r13_c192 bl[192] br[192] wl[13] vdd gnd cell_6t
Xbit_r14_c192 bl[192] br[192] wl[14] vdd gnd cell_6t
Xbit_r15_c192 bl[192] br[192] wl[15] vdd gnd cell_6t
Xbit_r16_c192 bl[192] br[192] wl[16] vdd gnd cell_6t
Xbit_r17_c192 bl[192] br[192] wl[17] vdd gnd cell_6t
Xbit_r18_c192 bl[192] br[192] wl[18] vdd gnd cell_6t
Xbit_r19_c192 bl[192] br[192] wl[19] vdd gnd cell_6t
Xbit_r20_c192 bl[192] br[192] wl[20] vdd gnd cell_6t
Xbit_r21_c192 bl[192] br[192] wl[21] vdd gnd cell_6t
Xbit_r22_c192 bl[192] br[192] wl[22] vdd gnd cell_6t
Xbit_r23_c192 bl[192] br[192] wl[23] vdd gnd cell_6t
Xbit_r24_c192 bl[192] br[192] wl[24] vdd gnd cell_6t
Xbit_r25_c192 bl[192] br[192] wl[25] vdd gnd cell_6t
Xbit_r26_c192 bl[192] br[192] wl[26] vdd gnd cell_6t
Xbit_r27_c192 bl[192] br[192] wl[27] vdd gnd cell_6t
Xbit_r28_c192 bl[192] br[192] wl[28] vdd gnd cell_6t
Xbit_r29_c192 bl[192] br[192] wl[29] vdd gnd cell_6t
Xbit_r30_c192 bl[192] br[192] wl[30] vdd gnd cell_6t
Xbit_r31_c192 bl[192] br[192] wl[31] vdd gnd cell_6t
Xbit_r32_c192 bl[192] br[192] wl[32] vdd gnd cell_6t
Xbit_r33_c192 bl[192] br[192] wl[33] vdd gnd cell_6t
Xbit_r34_c192 bl[192] br[192] wl[34] vdd gnd cell_6t
Xbit_r35_c192 bl[192] br[192] wl[35] vdd gnd cell_6t
Xbit_r36_c192 bl[192] br[192] wl[36] vdd gnd cell_6t
Xbit_r37_c192 bl[192] br[192] wl[37] vdd gnd cell_6t
Xbit_r38_c192 bl[192] br[192] wl[38] vdd gnd cell_6t
Xbit_r39_c192 bl[192] br[192] wl[39] vdd gnd cell_6t
Xbit_r40_c192 bl[192] br[192] wl[40] vdd gnd cell_6t
Xbit_r41_c192 bl[192] br[192] wl[41] vdd gnd cell_6t
Xbit_r42_c192 bl[192] br[192] wl[42] vdd gnd cell_6t
Xbit_r43_c192 bl[192] br[192] wl[43] vdd gnd cell_6t
Xbit_r44_c192 bl[192] br[192] wl[44] vdd gnd cell_6t
Xbit_r45_c192 bl[192] br[192] wl[45] vdd gnd cell_6t
Xbit_r46_c192 bl[192] br[192] wl[46] vdd gnd cell_6t
Xbit_r47_c192 bl[192] br[192] wl[47] vdd gnd cell_6t
Xbit_r48_c192 bl[192] br[192] wl[48] vdd gnd cell_6t
Xbit_r49_c192 bl[192] br[192] wl[49] vdd gnd cell_6t
Xbit_r50_c192 bl[192] br[192] wl[50] vdd gnd cell_6t
Xbit_r51_c192 bl[192] br[192] wl[51] vdd gnd cell_6t
Xbit_r52_c192 bl[192] br[192] wl[52] vdd gnd cell_6t
Xbit_r53_c192 bl[192] br[192] wl[53] vdd gnd cell_6t
Xbit_r54_c192 bl[192] br[192] wl[54] vdd gnd cell_6t
Xbit_r55_c192 bl[192] br[192] wl[55] vdd gnd cell_6t
Xbit_r56_c192 bl[192] br[192] wl[56] vdd gnd cell_6t
Xbit_r57_c192 bl[192] br[192] wl[57] vdd gnd cell_6t
Xbit_r58_c192 bl[192] br[192] wl[58] vdd gnd cell_6t
Xbit_r59_c192 bl[192] br[192] wl[59] vdd gnd cell_6t
Xbit_r60_c192 bl[192] br[192] wl[60] vdd gnd cell_6t
Xbit_r61_c192 bl[192] br[192] wl[61] vdd gnd cell_6t
Xbit_r62_c192 bl[192] br[192] wl[62] vdd gnd cell_6t
Xbit_r63_c192 bl[192] br[192] wl[63] vdd gnd cell_6t
Xbit_r64_c192 bl[192] br[192] wl[64] vdd gnd cell_6t
Xbit_r65_c192 bl[192] br[192] wl[65] vdd gnd cell_6t
Xbit_r66_c192 bl[192] br[192] wl[66] vdd gnd cell_6t
Xbit_r67_c192 bl[192] br[192] wl[67] vdd gnd cell_6t
Xbit_r68_c192 bl[192] br[192] wl[68] vdd gnd cell_6t
Xbit_r69_c192 bl[192] br[192] wl[69] vdd gnd cell_6t
Xbit_r70_c192 bl[192] br[192] wl[70] vdd gnd cell_6t
Xbit_r71_c192 bl[192] br[192] wl[71] vdd gnd cell_6t
Xbit_r72_c192 bl[192] br[192] wl[72] vdd gnd cell_6t
Xbit_r73_c192 bl[192] br[192] wl[73] vdd gnd cell_6t
Xbit_r74_c192 bl[192] br[192] wl[74] vdd gnd cell_6t
Xbit_r75_c192 bl[192] br[192] wl[75] vdd gnd cell_6t
Xbit_r76_c192 bl[192] br[192] wl[76] vdd gnd cell_6t
Xbit_r77_c192 bl[192] br[192] wl[77] vdd gnd cell_6t
Xbit_r78_c192 bl[192] br[192] wl[78] vdd gnd cell_6t
Xbit_r79_c192 bl[192] br[192] wl[79] vdd gnd cell_6t
Xbit_r80_c192 bl[192] br[192] wl[80] vdd gnd cell_6t
Xbit_r81_c192 bl[192] br[192] wl[81] vdd gnd cell_6t
Xbit_r82_c192 bl[192] br[192] wl[82] vdd gnd cell_6t
Xbit_r83_c192 bl[192] br[192] wl[83] vdd gnd cell_6t
Xbit_r84_c192 bl[192] br[192] wl[84] vdd gnd cell_6t
Xbit_r85_c192 bl[192] br[192] wl[85] vdd gnd cell_6t
Xbit_r86_c192 bl[192] br[192] wl[86] vdd gnd cell_6t
Xbit_r87_c192 bl[192] br[192] wl[87] vdd gnd cell_6t
Xbit_r88_c192 bl[192] br[192] wl[88] vdd gnd cell_6t
Xbit_r89_c192 bl[192] br[192] wl[89] vdd gnd cell_6t
Xbit_r90_c192 bl[192] br[192] wl[90] vdd gnd cell_6t
Xbit_r91_c192 bl[192] br[192] wl[91] vdd gnd cell_6t
Xbit_r92_c192 bl[192] br[192] wl[92] vdd gnd cell_6t
Xbit_r93_c192 bl[192] br[192] wl[93] vdd gnd cell_6t
Xbit_r94_c192 bl[192] br[192] wl[94] vdd gnd cell_6t
Xbit_r95_c192 bl[192] br[192] wl[95] vdd gnd cell_6t
Xbit_r96_c192 bl[192] br[192] wl[96] vdd gnd cell_6t
Xbit_r97_c192 bl[192] br[192] wl[97] vdd gnd cell_6t
Xbit_r98_c192 bl[192] br[192] wl[98] vdd gnd cell_6t
Xbit_r99_c192 bl[192] br[192] wl[99] vdd gnd cell_6t
Xbit_r100_c192 bl[192] br[192] wl[100] vdd gnd cell_6t
Xbit_r101_c192 bl[192] br[192] wl[101] vdd gnd cell_6t
Xbit_r102_c192 bl[192] br[192] wl[102] vdd gnd cell_6t
Xbit_r103_c192 bl[192] br[192] wl[103] vdd gnd cell_6t
Xbit_r104_c192 bl[192] br[192] wl[104] vdd gnd cell_6t
Xbit_r105_c192 bl[192] br[192] wl[105] vdd gnd cell_6t
Xbit_r106_c192 bl[192] br[192] wl[106] vdd gnd cell_6t
Xbit_r107_c192 bl[192] br[192] wl[107] vdd gnd cell_6t
Xbit_r108_c192 bl[192] br[192] wl[108] vdd gnd cell_6t
Xbit_r109_c192 bl[192] br[192] wl[109] vdd gnd cell_6t
Xbit_r110_c192 bl[192] br[192] wl[110] vdd gnd cell_6t
Xbit_r111_c192 bl[192] br[192] wl[111] vdd gnd cell_6t
Xbit_r112_c192 bl[192] br[192] wl[112] vdd gnd cell_6t
Xbit_r113_c192 bl[192] br[192] wl[113] vdd gnd cell_6t
Xbit_r114_c192 bl[192] br[192] wl[114] vdd gnd cell_6t
Xbit_r115_c192 bl[192] br[192] wl[115] vdd gnd cell_6t
Xbit_r116_c192 bl[192] br[192] wl[116] vdd gnd cell_6t
Xbit_r117_c192 bl[192] br[192] wl[117] vdd gnd cell_6t
Xbit_r118_c192 bl[192] br[192] wl[118] vdd gnd cell_6t
Xbit_r119_c192 bl[192] br[192] wl[119] vdd gnd cell_6t
Xbit_r120_c192 bl[192] br[192] wl[120] vdd gnd cell_6t
Xbit_r121_c192 bl[192] br[192] wl[121] vdd gnd cell_6t
Xbit_r122_c192 bl[192] br[192] wl[122] vdd gnd cell_6t
Xbit_r123_c192 bl[192] br[192] wl[123] vdd gnd cell_6t
Xbit_r124_c192 bl[192] br[192] wl[124] vdd gnd cell_6t
Xbit_r125_c192 bl[192] br[192] wl[125] vdd gnd cell_6t
Xbit_r126_c192 bl[192] br[192] wl[126] vdd gnd cell_6t
Xbit_r127_c192 bl[192] br[192] wl[127] vdd gnd cell_6t
Xbit_r128_c192 bl[192] br[192] wl[128] vdd gnd cell_6t
Xbit_r129_c192 bl[192] br[192] wl[129] vdd gnd cell_6t
Xbit_r130_c192 bl[192] br[192] wl[130] vdd gnd cell_6t
Xbit_r131_c192 bl[192] br[192] wl[131] vdd gnd cell_6t
Xbit_r132_c192 bl[192] br[192] wl[132] vdd gnd cell_6t
Xbit_r133_c192 bl[192] br[192] wl[133] vdd gnd cell_6t
Xbit_r134_c192 bl[192] br[192] wl[134] vdd gnd cell_6t
Xbit_r135_c192 bl[192] br[192] wl[135] vdd gnd cell_6t
Xbit_r136_c192 bl[192] br[192] wl[136] vdd gnd cell_6t
Xbit_r137_c192 bl[192] br[192] wl[137] vdd gnd cell_6t
Xbit_r138_c192 bl[192] br[192] wl[138] vdd gnd cell_6t
Xbit_r139_c192 bl[192] br[192] wl[139] vdd gnd cell_6t
Xbit_r140_c192 bl[192] br[192] wl[140] vdd gnd cell_6t
Xbit_r141_c192 bl[192] br[192] wl[141] vdd gnd cell_6t
Xbit_r142_c192 bl[192] br[192] wl[142] vdd gnd cell_6t
Xbit_r143_c192 bl[192] br[192] wl[143] vdd gnd cell_6t
Xbit_r144_c192 bl[192] br[192] wl[144] vdd gnd cell_6t
Xbit_r145_c192 bl[192] br[192] wl[145] vdd gnd cell_6t
Xbit_r146_c192 bl[192] br[192] wl[146] vdd gnd cell_6t
Xbit_r147_c192 bl[192] br[192] wl[147] vdd gnd cell_6t
Xbit_r148_c192 bl[192] br[192] wl[148] vdd gnd cell_6t
Xbit_r149_c192 bl[192] br[192] wl[149] vdd gnd cell_6t
Xbit_r150_c192 bl[192] br[192] wl[150] vdd gnd cell_6t
Xbit_r151_c192 bl[192] br[192] wl[151] vdd gnd cell_6t
Xbit_r152_c192 bl[192] br[192] wl[152] vdd gnd cell_6t
Xbit_r153_c192 bl[192] br[192] wl[153] vdd gnd cell_6t
Xbit_r154_c192 bl[192] br[192] wl[154] vdd gnd cell_6t
Xbit_r155_c192 bl[192] br[192] wl[155] vdd gnd cell_6t
Xbit_r156_c192 bl[192] br[192] wl[156] vdd gnd cell_6t
Xbit_r157_c192 bl[192] br[192] wl[157] vdd gnd cell_6t
Xbit_r158_c192 bl[192] br[192] wl[158] vdd gnd cell_6t
Xbit_r159_c192 bl[192] br[192] wl[159] vdd gnd cell_6t
Xbit_r160_c192 bl[192] br[192] wl[160] vdd gnd cell_6t
Xbit_r161_c192 bl[192] br[192] wl[161] vdd gnd cell_6t
Xbit_r162_c192 bl[192] br[192] wl[162] vdd gnd cell_6t
Xbit_r163_c192 bl[192] br[192] wl[163] vdd gnd cell_6t
Xbit_r164_c192 bl[192] br[192] wl[164] vdd gnd cell_6t
Xbit_r165_c192 bl[192] br[192] wl[165] vdd gnd cell_6t
Xbit_r166_c192 bl[192] br[192] wl[166] vdd gnd cell_6t
Xbit_r167_c192 bl[192] br[192] wl[167] vdd gnd cell_6t
Xbit_r168_c192 bl[192] br[192] wl[168] vdd gnd cell_6t
Xbit_r169_c192 bl[192] br[192] wl[169] vdd gnd cell_6t
Xbit_r170_c192 bl[192] br[192] wl[170] vdd gnd cell_6t
Xbit_r171_c192 bl[192] br[192] wl[171] vdd gnd cell_6t
Xbit_r172_c192 bl[192] br[192] wl[172] vdd gnd cell_6t
Xbit_r173_c192 bl[192] br[192] wl[173] vdd gnd cell_6t
Xbit_r174_c192 bl[192] br[192] wl[174] vdd gnd cell_6t
Xbit_r175_c192 bl[192] br[192] wl[175] vdd gnd cell_6t
Xbit_r176_c192 bl[192] br[192] wl[176] vdd gnd cell_6t
Xbit_r177_c192 bl[192] br[192] wl[177] vdd gnd cell_6t
Xbit_r178_c192 bl[192] br[192] wl[178] vdd gnd cell_6t
Xbit_r179_c192 bl[192] br[192] wl[179] vdd gnd cell_6t
Xbit_r180_c192 bl[192] br[192] wl[180] vdd gnd cell_6t
Xbit_r181_c192 bl[192] br[192] wl[181] vdd gnd cell_6t
Xbit_r182_c192 bl[192] br[192] wl[182] vdd gnd cell_6t
Xbit_r183_c192 bl[192] br[192] wl[183] vdd gnd cell_6t
Xbit_r184_c192 bl[192] br[192] wl[184] vdd gnd cell_6t
Xbit_r185_c192 bl[192] br[192] wl[185] vdd gnd cell_6t
Xbit_r186_c192 bl[192] br[192] wl[186] vdd gnd cell_6t
Xbit_r187_c192 bl[192] br[192] wl[187] vdd gnd cell_6t
Xbit_r188_c192 bl[192] br[192] wl[188] vdd gnd cell_6t
Xbit_r189_c192 bl[192] br[192] wl[189] vdd gnd cell_6t
Xbit_r190_c192 bl[192] br[192] wl[190] vdd gnd cell_6t
Xbit_r191_c192 bl[192] br[192] wl[191] vdd gnd cell_6t
Xbit_r192_c192 bl[192] br[192] wl[192] vdd gnd cell_6t
Xbit_r193_c192 bl[192] br[192] wl[193] vdd gnd cell_6t
Xbit_r194_c192 bl[192] br[192] wl[194] vdd gnd cell_6t
Xbit_r195_c192 bl[192] br[192] wl[195] vdd gnd cell_6t
Xbit_r196_c192 bl[192] br[192] wl[196] vdd gnd cell_6t
Xbit_r197_c192 bl[192] br[192] wl[197] vdd gnd cell_6t
Xbit_r198_c192 bl[192] br[192] wl[198] vdd gnd cell_6t
Xbit_r199_c192 bl[192] br[192] wl[199] vdd gnd cell_6t
Xbit_r200_c192 bl[192] br[192] wl[200] vdd gnd cell_6t
Xbit_r201_c192 bl[192] br[192] wl[201] vdd gnd cell_6t
Xbit_r202_c192 bl[192] br[192] wl[202] vdd gnd cell_6t
Xbit_r203_c192 bl[192] br[192] wl[203] vdd gnd cell_6t
Xbit_r204_c192 bl[192] br[192] wl[204] vdd gnd cell_6t
Xbit_r205_c192 bl[192] br[192] wl[205] vdd gnd cell_6t
Xbit_r206_c192 bl[192] br[192] wl[206] vdd gnd cell_6t
Xbit_r207_c192 bl[192] br[192] wl[207] vdd gnd cell_6t
Xbit_r208_c192 bl[192] br[192] wl[208] vdd gnd cell_6t
Xbit_r209_c192 bl[192] br[192] wl[209] vdd gnd cell_6t
Xbit_r210_c192 bl[192] br[192] wl[210] vdd gnd cell_6t
Xbit_r211_c192 bl[192] br[192] wl[211] vdd gnd cell_6t
Xbit_r212_c192 bl[192] br[192] wl[212] vdd gnd cell_6t
Xbit_r213_c192 bl[192] br[192] wl[213] vdd gnd cell_6t
Xbit_r214_c192 bl[192] br[192] wl[214] vdd gnd cell_6t
Xbit_r215_c192 bl[192] br[192] wl[215] vdd gnd cell_6t
Xbit_r216_c192 bl[192] br[192] wl[216] vdd gnd cell_6t
Xbit_r217_c192 bl[192] br[192] wl[217] vdd gnd cell_6t
Xbit_r218_c192 bl[192] br[192] wl[218] vdd gnd cell_6t
Xbit_r219_c192 bl[192] br[192] wl[219] vdd gnd cell_6t
Xbit_r220_c192 bl[192] br[192] wl[220] vdd gnd cell_6t
Xbit_r221_c192 bl[192] br[192] wl[221] vdd gnd cell_6t
Xbit_r222_c192 bl[192] br[192] wl[222] vdd gnd cell_6t
Xbit_r223_c192 bl[192] br[192] wl[223] vdd gnd cell_6t
Xbit_r224_c192 bl[192] br[192] wl[224] vdd gnd cell_6t
Xbit_r225_c192 bl[192] br[192] wl[225] vdd gnd cell_6t
Xbit_r226_c192 bl[192] br[192] wl[226] vdd gnd cell_6t
Xbit_r227_c192 bl[192] br[192] wl[227] vdd gnd cell_6t
Xbit_r228_c192 bl[192] br[192] wl[228] vdd gnd cell_6t
Xbit_r229_c192 bl[192] br[192] wl[229] vdd gnd cell_6t
Xbit_r230_c192 bl[192] br[192] wl[230] vdd gnd cell_6t
Xbit_r231_c192 bl[192] br[192] wl[231] vdd gnd cell_6t
Xbit_r232_c192 bl[192] br[192] wl[232] vdd gnd cell_6t
Xbit_r233_c192 bl[192] br[192] wl[233] vdd gnd cell_6t
Xbit_r234_c192 bl[192] br[192] wl[234] vdd gnd cell_6t
Xbit_r235_c192 bl[192] br[192] wl[235] vdd gnd cell_6t
Xbit_r236_c192 bl[192] br[192] wl[236] vdd gnd cell_6t
Xbit_r237_c192 bl[192] br[192] wl[237] vdd gnd cell_6t
Xbit_r238_c192 bl[192] br[192] wl[238] vdd gnd cell_6t
Xbit_r239_c192 bl[192] br[192] wl[239] vdd gnd cell_6t
Xbit_r240_c192 bl[192] br[192] wl[240] vdd gnd cell_6t
Xbit_r241_c192 bl[192] br[192] wl[241] vdd gnd cell_6t
Xbit_r242_c192 bl[192] br[192] wl[242] vdd gnd cell_6t
Xbit_r243_c192 bl[192] br[192] wl[243] vdd gnd cell_6t
Xbit_r244_c192 bl[192] br[192] wl[244] vdd gnd cell_6t
Xbit_r245_c192 bl[192] br[192] wl[245] vdd gnd cell_6t
Xbit_r246_c192 bl[192] br[192] wl[246] vdd gnd cell_6t
Xbit_r247_c192 bl[192] br[192] wl[247] vdd gnd cell_6t
Xbit_r248_c192 bl[192] br[192] wl[248] vdd gnd cell_6t
Xbit_r249_c192 bl[192] br[192] wl[249] vdd gnd cell_6t
Xbit_r250_c192 bl[192] br[192] wl[250] vdd gnd cell_6t
Xbit_r251_c192 bl[192] br[192] wl[251] vdd gnd cell_6t
Xbit_r252_c192 bl[192] br[192] wl[252] vdd gnd cell_6t
Xbit_r253_c192 bl[192] br[192] wl[253] vdd gnd cell_6t
Xbit_r254_c192 bl[192] br[192] wl[254] vdd gnd cell_6t
Xbit_r255_c192 bl[192] br[192] wl[255] vdd gnd cell_6t
Xbit_r0_c193 bl[193] br[193] wl[0] vdd gnd cell_6t
Xbit_r1_c193 bl[193] br[193] wl[1] vdd gnd cell_6t
Xbit_r2_c193 bl[193] br[193] wl[2] vdd gnd cell_6t
Xbit_r3_c193 bl[193] br[193] wl[3] vdd gnd cell_6t
Xbit_r4_c193 bl[193] br[193] wl[4] vdd gnd cell_6t
Xbit_r5_c193 bl[193] br[193] wl[5] vdd gnd cell_6t
Xbit_r6_c193 bl[193] br[193] wl[6] vdd gnd cell_6t
Xbit_r7_c193 bl[193] br[193] wl[7] vdd gnd cell_6t
Xbit_r8_c193 bl[193] br[193] wl[8] vdd gnd cell_6t
Xbit_r9_c193 bl[193] br[193] wl[9] vdd gnd cell_6t
Xbit_r10_c193 bl[193] br[193] wl[10] vdd gnd cell_6t
Xbit_r11_c193 bl[193] br[193] wl[11] vdd gnd cell_6t
Xbit_r12_c193 bl[193] br[193] wl[12] vdd gnd cell_6t
Xbit_r13_c193 bl[193] br[193] wl[13] vdd gnd cell_6t
Xbit_r14_c193 bl[193] br[193] wl[14] vdd gnd cell_6t
Xbit_r15_c193 bl[193] br[193] wl[15] vdd gnd cell_6t
Xbit_r16_c193 bl[193] br[193] wl[16] vdd gnd cell_6t
Xbit_r17_c193 bl[193] br[193] wl[17] vdd gnd cell_6t
Xbit_r18_c193 bl[193] br[193] wl[18] vdd gnd cell_6t
Xbit_r19_c193 bl[193] br[193] wl[19] vdd gnd cell_6t
Xbit_r20_c193 bl[193] br[193] wl[20] vdd gnd cell_6t
Xbit_r21_c193 bl[193] br[193] wl[21] vdd gnd cell_6t
Xbit_r22_c193 bl[193] br[193] wl[22] vdd gnd cell_6t
Xbit_r23_c193 bl[193] br[193] wl[23] vdd gnd cell_6t
Xbit_r24_c193 bl[193] br[193] wl[24] vdd gnd cell_6t
Xbit_r25_c193 bl[193] br[193] wl[25] vdd gnd cell_6t
Xbit_r26_c193 bl[193] br[193] wl[26] vdd gnd cell_6t
Xbit_r27_c193 bl[193] br[193] wl[27] vdd gnd cell_6t
Xbit_r28_c193 bl[193] br[193] wl[28] vdd gnd cell_6t
Xbit_r29_c193 bl[193] br[193] wl[29] vdd gnd cell_6t
Xbit_r30_c193 bl[193] br[193] wl[30] vdd gnd cell_6t
Xbit_r31_c193 bl[193] br[193] wl[31] vdd gnd cell_6t
Xbit_r32_c193 bl[193] br[193] wl[32] vdd gnd cell_6t
Xbit_r33_c193 bl[193] br[193] wl[33] vdd gnd cell_6t
Xbit_r34_c193 bl[193] br[193] wl[34] vdd gnd cell_6t
Xbit_r35_c193 bl[193] br[193] wl[35] vdd gnd cell_6t
Xbit_r36_c193 bl[193] br[193] wl[36] vdd gnd cell_6t
Xbit_r37_c193 bl[193] br[193] wl[37] vdd gnd cell_6t
Xbit_r38_c193 bl[193] br[193] wl[38] vdd gnd cell_6t
Xbit_r39_c193 bl[193] br[193] wl[39] vdd gnd cell_6t
Xbit_r40_c193 bl[193] br[193] wl[40] vdd gnd cell_6t
Xbit_r41_c193 bl[193] br[193] wl[41] vdd gnd cell_6t
Xbit_r42_c193 bl[193] br[193] wl[42] vdd gnd cell_6t
Xbit_r43_c193 bl[193] br[193] wl[43] vdd gnd cell_6t
Xbit_r44_c193 bl[193] br[193] wl[44] vdd gnd cell_6t
Xbit_r45_c193 bl[193] br[193] wl[45] vdd gnd cell_6t
Xbit_r46_c193 bl[193] br[193] wl[46] vdd gnd cell_6t
Xbit_r47_c193 bl[193] br[193] wl[47] vdd gnd cell_6t
Xbit_r48_c193 bl[193] br[193] wl[48] vdd gnd cell_6t
Xbit_r49_c193 bl[193] br[193] wl[49] vdd gnd cell_6t
Xbit_r50_c193 bl[193] br[193] wl[50] vdd gnd cell_6t
Xbit_r51_c193 bl[193] br[193] wl[51] vdd gnd cell_6t
Xbit_r52_c193 bl[193] br[193] wl[52] vdd gnd cell_6t
Xbit_r53_c193 bl[193] br[193] wl[53] vdd gnd cell_6t
Xbit_r54_c193 bl[193] br[193] wl[54] vdd gnd cell_6t
Xbit_r55_c193 bl[193] br[193] wl[55] vdd gnd cell_6t
Xbit_r56_c193 bl[193] br[193] wl[56] vdd gnd cell_6t
Xbit_r57_c193 bl[193] br[193] wl[57] vdd gnd cell_6t
Xbit_r58_c193 bl[193] br[193] wl[58] vdd gnd cell_6t
Xbit_r59_c193 bl[193] br[193] wl[59] vdd gnd cell_6t
Xbit_r60_c193 bl[193] br[193] wl[60] vdd gnd cell_6t
Xbit_r61_c193 bl[193] br[193] wl[61] vdd gnd cell_6t
Xbit_r62_c193 bl[193] br[193] wl[62] vdd gnd cell_6t
Xbit_r63_c193 bl[193] br[193] wl[63] vdd gnd cell_6t
Xbit_r64_c193 bl[193] br[193] wl[64] vdd gnd cell_6t
Xbit_r65_c193 bl[193] br[193] wl[65] vdd gnd cell_6t
Xbit_r66_c193 bl[193] br[193] wl[66] vdd gnd cell_6t
Xbit_r67_c193 bl[193] br[193] wl[67] vdd gnd cell_6t
Xbit_r68_c193 bl[193] br[193] wl[68] vdd gnd cell_6t
Xbit_r69_c193 bl[193] br[193] wl[69] vdd gnd cell_6t
Xbit_r70_c193 bl[193] br[193] wl[70] vdd gnd cell_6t
Xbit_r71_c193 bl[193] br[193] wl[71] vdd gnd cell_6t
Xbit_r72_c193 bl[193] br[193] wl[72] vdd gnd cell_6t
Xbit_r73_c193 bl[193] br[193] wl[73] vdd gnd cell_6t
Xbit_r74_c193 bl[193] br[193] wl[74] vdd gnd cell_6t
Xbit_r75_c193 bl[193] br[193] wl[75] vdd gnd cell_6t
Xbit_r76_c193 bl[193] br[193] wl[76] vdd gnd cell_6t
Xbit_r77_c193 bl[193] br[193] wl[77] vdd gnd cell_6t
Xbit_r78_c193 bl[193] br[193] wl[78] vdd gnd cell_6t
Xbit_r79_c193 bl[193] br[193] wl[79] vdd gnd cell_6t
Xbit_r80_c193 bl[193] br[193] wl[80] vdd gnd cell_6t
Xbit_r81_c193 bl[193] br[193] wl[81] vdd gnd cell_6t
Xbit_r82_c193 bl[193] br[193] wl[82] vdd gnd cell_6t
Xbit_r83_c193 bl[193] br[193] wl[83] vdd gnd cell_6t
Xbit_r84_c193 bl[193] br[193] wl[84] vdd gnd cell_6t
Xbit_r85_c193 bl[193] br[193] wl[85] vdd gnd cell_6t
Xbit_r86_c193 bl[193] br[193] wl[86] vdd gnd cell_6t
Xbit_r87_c193 bl[193] br[193] wl[87] vdd gnd cell_6t
Xbit_r88_c193 bl[193] br[193] wl[88] vdd gnd cell_6t
Xbit_r89_c193 bl[193] br[193] wl[89] vdd gnd cell_6t
Xbit_r90_c193 bl[193] br[193] wl[90] vdd gnd cell_6t
Xbit_r91_c193 bl[193] br[193] wl[91] vdd gnd cell_6t
Xbit_r92_c193 bl[193] br[193] wl[92] vdd gnd cell_6t
Xbit_r93_c193 bl[193] br[193] wl[93] vdd gnd cell_6t
Xbit_r94_c193 bl[193] br[193] wl[94] vdd gnd cell_6t
Xbit_r95_c193 bl[193] br[193] wl[95] vdd gnd cell_6t
Xbit_r96_c193 bl[193] br[193] wl[96] vdd gnd cell_6t
Xbit_r97_c193 bl[193] br[193] wl[97] vdd gnd cell_6t
Xbit_r98_c193 bl[193] br[193] wl[98] vdd gnd cell_6t
Xbit_r99_c193 bl[193] br[193] wl[99] vdd gnd cell_6t
Xbit_r100_c193 bl[193] br[193] wl[100] vdd gnd cell_6t
Xbit_r101_c193 bl[193] br[193] wl[101] vdd gnd cell_6t
Xbit_r102_c193 bl[193] br[193] wl[102] vdd gnd cell_6t
Xbit_r103_c193 bl[193] br[193] wl[103] vdd gnd cell_6t
Xbit_r104_c193 bl[193] br[193] wl[104] vdd gnd cell_6t
Xbit_r105_c193 bl[193] br[193] wl[105] vdd gnd cell_6t
Xbit_r106_c193 bl[193] br[193] wl[106] vdd gnd cell_6t
Xbit_r107_c193 bl[193] br[193] wl[107] vdd gnd cell_6t
Xbit_r108_c193 bl[193] br[193] wl[108] vdd gnd cell_6t
Xbit_r109_c193 bl[193] br[193] wl[109] vdd gnd cell_6t
Xbit_r110_c193 bl[193] br[193] wl[110] vdd gnd cell_6t
Xbit_r111_c193 bl[193] br[193] wl[111] vdd gnd cell_6t
Xbit_r112_c193 bl[193] br[193] wl[112] vdd gnd cell_6t
Xbit_r113_c193 bl[193] br[193] wl[113] vdd gnd cell_6t
Xbit_r114_c193 bl[193] br[193] wl[114] vdd gnd cell_6t
Xbit_r115_c193 bl[193] br[193] wl[115] vdd gnd cell_6t
Xbit_r116_c193 bl[193] br[193] wl[116] vdd gnd cell_6t
Xbit_r117_c193 bl[193] br[193] wl[117] vdd gnd cell_6t
Xbit_r118_c193 bl[193] br[193] wl[118] vdd gnd cell_6t
Xbit_r119_c193 bl[193] br[193] wl[119] vdd gnd cell_6t
Xbit_r120_c193 bl[193] br[193] wl[120] vdd gnd cell_6t
Xbit_r121_c193 bl[193] br[193] wl[121] vdd gnd cell_6t
Xbit_r122_c193 bl[193] br[193] wl[122] vdd gnd cell_6t
Xbit_r123_c193 bl[193] br[193] wl[123] vdd gnd cell_6t
Xbit_r124_c193 bl[193] br[193] wl[124] vdd gnd cell_6t
Xbit_r125_c193 bl[193] br[193] wl[125] vdd gnd cell_6t
Xbit_r126_c193 bl[193] br[193] wl[126] vdd gnd cell_6t
Xbit_r127_c193 bl[193] br[193] wl[127] vdd gnd cell_6t
Xbit_r128_c193 bl[193] br[193] wl[128] vdd gnd cell_6t
Xbit_r129_c193 bl[193] br[193] wl[129] vdd gnd cell_6t
Xbit_r130_c193 bl[193] br[193] wl[130] vdd gnd cell_6t
Xbit_r131_c193 bl[193] br[193] wl[131] vdd gnd cell_6t
Xbit_r132_c193 bl[193] br[193] wl[132] vdd gnd cell_6t
Xbit_r133_c193 bl[193] br[193] wl[133] vdd gnd cell_6t
Xbit_r134_c193 bl[193] br[193] wl[134] vdd gnd cell_6t
Xbit_r135_c193 bl[193] br[193] wl[135] vdd gnd cell_6t
Xbit_r136_c193 bl[193] br[193] wl[136] vdd gnd cell_6t
Xbit_r137_c193 bl[193] br[193] wl[137] vdd gnd cell_6t
Xbit_r138_c193 bl[193] br[193] wl[138] vdd gnd cell_6t
Xbit_r139_c193 bl[193] br[193] wl[139] vdd gnd cell_6t
Xbit_r140_c193 bl[193] br[193] wl[140] vdd gnd cell_6t
Xbit_r141_c193 bl[193] br[193] wl[141] vdd gnd cell_6t
Xbit_r142_c193 bl[193] br[193] wl[142] vdd gnd cell_6t
Xbit_r143_c193 bl[193] br[193] wl[143] vdd gnd cell_6t
Xbit_r144_c193 bl[193] br[193] wl[144] vdd gnd cell_6t
Xbit_r145_c193 bl[193] br[193] wl[145] vdd gnd cell_6t
Xbit_r146_c193 bl[193] br[193] wl[146] vdd gnd cell_6t
Xbit_r147_c193 bl[193] br[193] wl[147] vdd gnd cell_6t
Xbit_r148_c193 bl[193] br[193] wl[148] vdd gnd cell_6t
Xbit_r149_c193 bl[193] br[193] wl[149] vdd gnd cell_6t
Xbit_r150_c193 bl[193] br[193] wl[150] vdd gnd cell_6t
Xbit_r151_c193 bl[193] br[193] wl[151] vdd gnd cell_6t
Xbit_r152_c193 bl[193] br[193] wl[152] vdd gnd cell_6t
Xbit_r153_c193 bl[193] br[193] wl[153] vdd gnd cell_6t
Xbit_r154_c193 bl[193] br[193] wl[154] vdd gnd cell_6t
Xbit_r155_c193 bl[193] br[193] wl[155] vdd gnd cell_6t
Xbit_r156_c193 bl[193] br[193] wl[156] vdd gnd cell_6t
Xbit_r157_c193 bl[193] br[193] wl[157] vdd gnd cell_6t
Xbit_r158_c193 bl[193] br[193] wl[158] vdd gnd cell_6t
Xbit_r159_c193 bl[193] br[193] wl[159] vdd gnd cell_6t
Xbit_r160_c193 bl[193] br[193] wl[160] vdd gnd cell_6t
Xbit_r161_c193 bl[193] br[193] wl[161] vdd gnd cell_6t
Xbit_r162_c193 bl[193] br[193] wl[162] vdd gnd cell_6t
Xbit_r163_c193 bl[193] br[193] wl[163] vdd gnd cell_6t
Xbit_r164_c193 bl[193] br[193] wl[164] vdd gnd cell_6t
Xbit_r165_c193 bl[193] br[193] wl[165] vdd gnd cell_6t
Xbit_r166_c193 bl[193] br[193] wl[166] vdd gnd cell_6t
Xbit_r167_c193 bl[193] br[193] wl[167] vdd gnd cell_6t
Xbit_r168_c193 bl[193] br[193] wl[168] vdd gnd cell_6t
Xbit_r169_c193 bl[193] br[193] wl[169] vdd gnd cell_6t
Xbit_r170_c193 bl[193] br[193] wl[170] vdd gnd cell_6t
Xbit_r171_c193 bl[193] br[193] wl[171] vdd gnd cell_6t
Xbit_r172_c193 bl[193] br[193] wl[172] vdd gnd cell_6t
Xbit_r173_c193 bl[193] br[193] wl[173] vdd gnd cell_6t
Xbit_r174_c193 bl[193] br[193] wl[174] vdd gnd cell_6t
Xbit_r175_c193 bl[193] br[193] wl[175] vdd gnd cell_6t
Xbit_r176_c193 bl[193] br[193] wl[176] vdd gnd cell_6t
Xbit_r177_c193 bl[193] br[193] wl[177] vdd gnd cell_6t
Xbit_r178_c193 bl[193] br[193] wl[178] vdd gnd cell_6t
Xbit_r179_c193 bl[193] br[193] wl[179] vdd gnd cell_6t
Xbit_r180_c193 bl[193] br[193] wl[180] vdd gnd cell_6t
Xbit_r181_c193 bl[193] br[193] wl[181] vdd gnd cell_6t
Xbit_r182_c193 bl[193] br[193] wl[182] vdd gnd cell_6t
Xbit_r183_c193 bl[193] br[193] wl[183] vdd gnd cell_6t
Xbit_r184_c193 bl[193] br[193] wl[184] vdd gnd cell_6t
Xbit_r185_c193 bl[193] br[193] wl[185] vdd gnd cell_6t
Xbit_r186_c193 bl[193] br[193] wl[186] vdd gnd cell_6t
Xbit_r187_c193 bl[193] br[193] wl[187] vdd gnd cell_6t
Xbit_r188_c193 bl[193] br[193] wl[188] vdd gnd cell_6t
Xbit_r189_c193 bl[193] br[193] wl[189] vdd gnd cell_6t
Xbit_r190_c193 bl[193] br[193] wl[190] vdd gnd cell_6t
Xbit_r191_c193 bl[193] br[193] wl[191] vdd gnd cell_6t
Xbit_r192_c193 bl[193] br[193] wl[192] vdd gnd cell_6t
Xbit_r193_c193 bl[193] br[193] wl[193] vdd gnd cell_6t
Xbit_r194_c193 bl[193] br[193] wl[194] vdd gnd cell_6t
Xbit_r195_c193 bl[193] br[193] wl[195] vdd gnd cell_6t
Xbit_r196_c193 bl[193] br[193] wl[196] vdd gnd cell_6t
Xbit_r197_c193 bl[193] br[193] wl[197] vdd gnd cell_6t
Xbit_r198_c193 bl[193] br[193] wl[198] vdd gnd cell_6t
Xbit_r199_c193 bl[193] br[193] wl[199] vdd gnd cell_6t
Xbit_r200_c193 bl[193] br[193] wl[200] vdd gnd cell_6t
Xbit_r201_c193 bl[193] br[193] wl[201] vdd gnd cell_6t
Xbit_r202_c193 bl[193] br[193] wl[202] vdd gnd cell_6t
Xbit_r203_c193 bl[193] br[193] wl[203] vdd gnd cell_6t
Xbit_r204_c193 bl[193] br[193] wl[204] vdd gnd cell_6t
Xbit_r205_c193 bl[193] br[193] wl[205] vdd gnd cell_6t
Xbit_r206_c193 bl[193] br[193] wl[206] vdd gnd cell_6t
Xbit_r207_c193 bl[193] br[193] wl[207] vdd gnd cell_6t
Xbit_r208_c193 bl[193] br[193] wl[208] vdd gnd cell_6t
Xbit_r209_c193 bl[193] br[193] wl[209] vdd gnd cell_6t
Xbit_r210_c193 bl[193] br[193] wl[210] vdd gnd cell_6t
Xbit_r211_c193 bl[193] br[193] wl[211] vdd gnd cell_6t
Xbit_r212_c193 bl[193] br[193] wl[212] vdd gnd cell_6t
Xbit_r213_c193 bl[193] br[193] wl[213] vdd gnd cell_6t
Xbit_r214_c193 bl[193] br[193] wl[214] vdd gnd cell_6t
Xbit_r215_c193 bl[193] br[193] wl[215] vdd gnd cell_6t
Xbit_r216_c193 bl[193] br[193] wl[216] vdd gnd cell_6t
Xbit_r217_c193 bl[193] br[193] wl[217] vdd gnd cell_6t
Xbit_r218_c193 bl[193] br[193] wl[218] vdd gnd cell_6t
Xbit_r219_c193 bl[193] br[193] wl[219] vdd gnd cell_6t
Xbit_r220_c193 bl[193] br[193] wl[220] vdd gnd cell_6t
Xbit_r221_c193 bl[193] br[193] wl[221] vdd gnd cell_6t
Xbit_r222_c193 bl[193] br[193] wl[222] vdd gnd cell_6t
Xbit_r223_c193 bl[193] br[193] wl[223] vdd gnd cell_6t
Xbit_r224_c193 bl[193] br[193] wl[224] vdd gnd cell_6t
Xbit_r225_c193 bl[193] br[193] wl[225] vdd gnd cell_6t
Xbit_r226_c193 bl[193] br[193] wl[226] vdd gnd cell_6t
Xbit_r227_c193 bl[193] br[193] wl[227] vdd gnd cell_6t
Xbit_r228_c193 bl[193] br[193] wl[228] vdd gnd cell_6t
Xbit_r229_c193 bl[193] br[193] wl[229] vdd gnd cell_6t
Xbit_r230_c193 bl[193] br[193] wl[230] vdd gnd cell_6t
Xbit_r231_c193 bl[193] br[193] wl[231] vdd gnd cell_6t
Xbit_r232_c193 bl[193] br[193] wl[232] vdd gnd cell_6t
Xbit_r233_c193 bl[193] br[193] wl[233] vdd gnd cell_6t
Xbit_r234_c193 bl[193] br[193] wl[234] vdd gnd cell_6t
Xbit_r235_c193 bl[193] br[193] wl[235] vdd gnd cell_6t
Xbit_r236_c193 bl[193] br[193] wl[236] vdd gnd cell_6t
Xbit_r237_c193 bl[193] br[193] wl[237] vdd gnd cell_6t
Xbit_r238_c193 bl[193] br[193] wl[238] vdd gnd cell_6t
Xbit_r239_c193 bl[193] br[193] wl[239] vdd gnd cell_6t
Xbit_r240_c193 bl[193] br[193] wl[240] vdd gnd cell_6t
Xbit_r241_c193 bl[193] br[193] wl[241] vdd gnd cell_6t
Xbit_r242_c193 bl[193] br[193] wl[242] vdd gnd cell_6t
Xbit_r243_c193 bl[193] br[193] wl[243] vdd gnd cell_6t
Xbit_r244_c193 bl[193] br[193] wl[244] vdd gnd cell_6t
Xbit_r245_c193 bl[193] br[193] wl[245] vdd gnd cell_6t
Xbit_r246_c193 bl[193] br[193] wl[246] vdd gnd cell_6t
Xbit_r247_c193 bl[193] br[193] wl[247] vdd gnd cell_6t
Xbit_r248_c193 bl[193] br[193] wl[248] vdd gnd cell_6t
Xbit_r249_c193 bl[193] br[193] wl[249] vdd gnd cell_6t
Xbit_r250_c193 bl[193] br[193] wl[250] vdd gnd cell_6t
Xbit_r251_c193 bl[193] br[193] wl[251] vdd gnd cell_6t
Xbit_r252_c193 bl[193] br[193] wl[252] vdd gnd cell_6t
Xbit_r253_c193 bl[193] br[193] wl[253] vdd gnd cell_6t
Xbit_r254_c193 bl[193] br[193] wl[254] vdd gnd cell_6t
Xbit_r255_c193 bl[193] br[193] wl[255] vdd gnd cell_6t
Xbit_r0_c194 bl[194] br[194] wl[0] vdd gnd cell_6t
Xbit_r1_c194 bl[194] br[194] wl[1] vdd gnd cell_6t
Xbit_r2_c194 bl[194] br[194] wl[2] vdd gnd cell_6t
Xbit_r3_c194 bl[194] br[194] wl[3] vdd gnd cell_6t
Xbit_r4_c194 bl[194] br[194] wl[4] vdd gnd cell_6t
Xbit_r5_c194 bl[194] br[194] wl[5] vdd gnd cell_6t
Xbit_r6_c194 bl[194] br[194] wl[6] vdd gnd cell_6t
Xbit_r7_c194 bl[194] br[194] wl[7] vdd gnd cell_6t
Xbit_r8_c194 bl[194] br[194] wl[8] vdd gnd cell_6t
Xbit_r9_c194 bl[194] br[194] wl[9] vdd gnd cell_6t
Xbit_r10_c194 bl[194] br[194] wl[10] vdd gnd cell_6t
Xbit_r11_c194 bl[194] br[194] wl[11] vdd gnd cell_6t
Xbit_r12_c194 bl[194] br[194] wl[12] vdd gnd cell_6t
Xbit_r13_c194 bl[194] br[194] wl[13] vdd gnd cell_6t
Xbit_r14_c194 bl[194] br[194] wl[14] vdd gnd cell_6t
Xbit_r15_c194 bl[194] br[194] wl[15] vdd gnd cell_6t
Xbit_r16_c194 bl[194] br[194] wl[16] vdd gnd cell_6t
Xbit_r17_c194 bl[194] br[194] wl[17] vdd gnd cell_6t
Xbit_r18_c194 bl[194] br[194] wl[18] vdd gnd cell_6t
Xbit_r19_c194 bl[194] br[194] wl[19] vdd gnd cell_6t
Xbit_r20_c194 bl[194] br[194] wl[20] vdd gnd cell_6t
Xbit_r21_c194 bl[194] br[194] wl[21] vdd gnd cell_6t
Xbit_r22_c194 bl[194] br[194] wl[22] vdd gnd cell_6t
Xbit_r23_c194 bl[194] br[194] wl[23] vdd gnd cell_6t
Xbit_r24_c194 bl[194] br[194] wl[24] vdd gnd cell_6t
Xbit_r25_c194 bl[194] br[194] wl[25] vdd gnd cell_6t
Xbit_r26_c194 bl[194] br[194] wl[26] vdd gnd cell_6t
Xbit_r27_c194 bl[194] br[194] wl[27] vdd gnd cell_6t
Xbit_r28_c194 bl[194] br[194] wl[28] vdd gnd cell_6t
Xbit_r29_c194 bl[194] br[194] wl[29] vdd gnd cell_6t
Xbit_r30_c194 bl[194] br[194] wl[30] vdd gnd cell_6t
Xbit_r31_c194 bl[194] br[194] wl[31] vdd gnd cell_6t
Xbit_r32_c194 bl[194] br[194] wl[32] vdd gnd cell_6t
Xbit_r33_c194 bl[194] br[194] wl[33] vdd gnd cell_6t
Xbit_r34_c194 bl[194] br[194] wl[34] vdd gnd cell_6t
Xbit_r35_c194 bl[194] br[194] wl[35] vdd gnd cell_6t
Xbit_r36_c194 bl[194] br[194] wl[36] vdd gnd cell_6t
Xbit_r37_c194 bl[194] br[194] wl[37] vdd gnd cell_6t
Xbit_r38_c194 bl[194] br[194] wl[38] vdd gnd cell_6t
Xbit_r39_c194 bl[194] br[194] wl[39] vdd gnd cell_6t
Xbit_r40_c194 bl[194] br[194] wl[40] vdd gnd cell_6t
Xbit_r41_c194 bl[194] br[194] wl[41] vdd gnd cell_6t
Xbit_r42_c194 bl[194] br[194] wl[42] vdd gnd cell_6t
Xbit_r43_c194 bl[194] br[194] wl[43] vdd gnd cell_6t
Xbit_r44_c194 bl[194] br[194] wl[44] vdd gnd cell_6t
Xbit_r45_c194 bl[194] br[194] wl[45] vdd gnd cell_6t
Xbit_r46_c194 bl[194] br[194] wl[46] vdd gnd cell_6t
Xbit_r47_c194 bl[194] br[194] wl[47] vdd gnd cell_6t
Xbit_r48_c194 bl[194] br[194] wl[48] vdd gnd cell_6t
Xbit_r49_c194 bl[194] br[194] wl[49] vdd gnd cell_6t
Xbit_r50_c194 bl[194] br[194] wl[50] vdd gnd cell_6t
Xbit_r51_c194 bl[194] br[194] wl[51] vdd gnd cell_6t
Xbit_r52_c194 bl[194] br[194] wl[52] vdd gnd cell_6t
Xbit_r53_c194 bl[194] br[194] wl[53] vdd gnd cell_6t
Xbit_r54_c194 bl[194] br[194] wl[54] vdd gnd cell_6t
Xbit_r55_c194 bl[194] br[194] wl[55] vdd gnd cell_6t
Xbit_r56_c194 bl[194] br[194] wl[56] vdd gnd cell_6t
Xbit_r57_c194 bl[194] br[194] wl[57] vdd gnd cell_6t
Xbit_r58_c194 bl[194] br[194] wl[58] vdd gnd cell_6t
Xbit_r59_c194 bl[194] br[194] wl[59] vdd gnd cell_6t
Xbit_r60_c194 bl[194] br[194] wl[60] vdd gnd cell_6t
Xbit_r61_c194 bl[194] br[194] wl[61] vdd gnd cell_6t
Xbit_r62_c194 bl[194] br[194] wl[62] vdd gnd cell_6t
Xbit_r63_c194 bl[194] br[194] wl[63] vdd gnd cell_6t
Xbit_r64_c194 bl[194] br[194] wl[64] vdd gnd cell_6t
Xbit_r65_c194 bl[194] br[194] wl[65] vdd gnd cell_6t
Xbit_r66_c194 bl[194] br[194] wl[66] vdd gnd cell_6t
Xbit_r67_c194 bl[194] br[194] wl[67] vdd gnd cell_6t
Xbit_r68_c194 bl[194] br[194] wl[68] vdd gnd cell_6t
Xbit_r69_c194 bl[194] br[194] wl[69] vdd gnd cell_6t
Xbit_r70_c194 bl[194] br[194] wl[70] vdd gnd cell_6t
Xbit_r71_c194 bl[194] br[194] wl[71] vdd gnd cell_6t
Xbit_r72_c194 bl[194] br[194] wl[72] vdd gnd cell_6t
Xbit_r73_c194 bl[194] br[194] wl[73] vdd gnd cell_6t
Xbit_r74_c194 bl[194] br[194] wl[74] vdd gnd cell_6t
Xbit_r75_c194 bl[194] br[194] wl[75] vdd gnd cell_6t
Xbit_r76_c194 bl[194] br[194] wl[76] vdd gnd cell_6t
Xbit_r77_c194 bl[194] br[194] wl[77] vdd gnd cell_6t
Xbit_r78_c194 bl[194] br[194] wl[78] vdd gnd cell_6t
Xbit_r79_c194 bl[194] br[194] wl[79] vdd gnd cell_6t
Xbit_r80_c194 bl[194] br[194] wl[80] vdd gnd cell_6t
Xbit_r81_c194 bl[194] br[194] wl[81] vdd gnd cell_6t
Xbit_r82_c194 bl[194] br[194] wl[82] vdd gnd cell_6t
Xbit_r83_c194 bl[194] br[194] wl[83] vdd gnd cell_6t
Xbit_r84_c194 bl[194] br[194] wl[84] vdd gnd cell_6t
Xbit_r85_c194 bl[194] br[194] wl[85] vdd gnd cell_6t
Xbit_r86_c194 bl[194] br[194] wl[86] vdd gnd cell_6t
Xbit_r87_c194 bl[194] br[194] wl[87] vdd gnd cell_6t
Xbit_r88_c194 bl[194] br[194] wl[88] vdd gnd cell_6t
Xbit_r89_c194 bl[194] br[194] wl[89] vdd gnd cell_6t
Xbit_r90_c194 bl[194] br[194] wl[90] vdd gnd cell_6t
Xbit_r91_c194 bl[194] br[194] wl[91] vdd gnd cell_6t
Xbit_r92_c194 bl[194] br[194] wl[92] vdd gnd cell_6t
Xbit_r93_c194 bl[194] br[194] wl[93] vdd gnd cell_6t
Xbit_r94_c194 bl[194] br[194] wl[94] vdd gnd cell_6t
Xbit_r95_c194 bl[194] br[194] wl[95] vdd gnd cell_6t
Xbit_r96_c194 bl[194] br[194] wl[96] vdd gnd cell_6t
Xbit_r97_c194 bl[194] br[194] wl[97] vdd gnd cell_6t
Xbit_r98_c194 bl[194] br[194] wl[98] vdd gnd cell_6t
Xbit_r99_c194 bl[194] br[194] wl[99] vdd gnd cell_6t
Xbit_r100_c194 bl[194] br[194] wl[100] vdd gnd cell_6t
Xbit_r101_c194 bl[194] br[194] wl[101] vdd gnd cell_6t
Xbit_r102_c194 bl[194] br[194] wl[102] vdd gnd cell_6t
Xbit_r103_c194 bl[194] br[194] wl[103] vdd gnd cell_6t
Xbit_r104_c194 bl[194] br[194] wl[104] vdd gnd cell_6t
Xbit_r105_c194 bl[194] br[194] wl[105] vdd gnd cell_6t
Xbit_r106_c194 bl[194] br[194] wl[106] vdd gnd cell_6t
Xbit_r107_c194 bl[194] br[194] wl[107] vdd gnd cell_6t
Xbit_r108_c194 bl[194] br[194] wl[108] vdd gnd cell_6t
Xbit_r109_c194 bl[194] br[194] wl[109] vdd gnd cell_6t
Xbit_r110_c194 bl[194] br[194] wl[110] vdd gnd cell_6t
Xbit_r111_c194 bl[194] br[194] wl[111] vdd gnd cell_6t
Xbit_r112_c194 bl[194] br[194] wl[112] vdd gnd cell_6t
Xbit_r113_c194 bl[194] br[194] wl[113] vdd gnd cell_6t
Xbit_r114_c194 bl[194] br[194] wl[114] vdd gnd cell_6t
Xbit_r115_c194 bl[194] br[194] wl[115] vdd gnd cell_6t
Xbit_r116_c194 bl[194] br[194] wl[116] vdd gnd cell_6t
Xbit_r117_c194 bl[194] br[194] wl[117] vdd gnd cell_6t
Xbit_r118_c194 bl[194] br[194] wl[118] vdd gnd cell_6t
Xbit_r119_c194 bl[194] br[194] wl[119] vdd gnd cell_6t
Xbit_r120_c194 bl[194] br[194] wl[120] vdd gnd cell_6t
Xbit_r121_c194 bl[194] br[194] wl[121] vdd gnd cell_6t
Xbit_r122_c194 bl[194] br[194] wl[122] vdd gnd cell_6t
Xbit_r123_c194 bl[194] br[194] wl[123] vdd gnd cell_6t
Xbit_r124_c194 bl[194] br[194] wl[124] vdd gnd cell_6t
Xbit_r125_c194 bl[194] br[194] wl[125] vdd gnd cell_6t
Xbit_r126_c194 bl[194] br[194] wl[126] vdd gnd cell_6t
Xbit_r127_c194 bl[194] br[194] wl[127] vdd gnd cell_6t
Xbit_r128_c194 bl[194] br[194] wl[128] vdd gnd cell_6t
Xbit_r129_c194 bl[194] br[194] wl[129] vdd gnd cell_6t
Xbit_r130_c194 bl[194] br[194] wl[130] vdd gnd cell_6t
Xbit_r131_c194 bl[194] br[194] wl[131] vdd gnd cell_6t
Xbit_r132_c194 bl[194] br[194] wl[132] vdd gnd cell_6t
Xbit_r133_c194 bl[194] br[194] wl[133] vdd gnd cell_6t
Xbit_r134_c194 bl[194] br[194] wl[134] vdd gnd cell_6t
Xbit_r135_c194 bl[194] br[194] wl[135] vdd gnd cell_6t
Xbit_r136_c194 bl[194] br[194] wl[136] vdd gnd cell_6t
Xbit_r137_c194 bl[194] br[194] wl[137] vdd gnd cell_6t
Xbit_r138_c194 bl[194] br[194] wl[138] vdd gnd cell_6t
Xbit_r139_c194 bl[194] br[194] wl[139] vdd gnd cell_6t
Xbit_r140_c194 bl[194] br[194] wl[140] vdd gnd cell_6t
Xbit_r141_c194 bl[194] br[194] wl[141] vdd gnd cell_6t
Xbit_r142_c194 bl[194] br[194] wl[142] vdd gnd cell_6t
Xbit_r143_c194 bl[194] br[194] wl[143] vdd gnd cell_6t
Xbit_r144_c194 bl[194] br[194] wl[144] vdd gnd cell_6t
Xbit_r145_c194 bl[194] br[194] wl[145] vdd gnd cell_6t
Xbit_r146_c194 bl[194] br[194] wl[146] vdd gnd cell_6t
Xbit_r147_c194 bl[194] br[194] wl[147] vdd gnd cell_6t
Xbit_r148_c194 bl[194] br[194] wl[148] vdd gnd cell_6t
Xbit_r149_c194 bl[194] br[194] wl[149] vdd gnd cell_6t
Xbit_r150_c194 bl[194] br[194] wl[150] vdd gnd cell_6t
Xbit_r151_c194 bl[194] br[194] wl[151] vdd gnd cell_6t
Xbit_r152_c194 bl[194] br[194] wl[152] vdd gnd cell_6t
Xbit_r153_c194 bl[194] br[194] wl[153] vdd gnd cell_6t
Xbit_r154_c194 bl[194] br[194] wl[154] vdd gnd cell_6t
Xbit_r155_c194 bl[194] br[194] wl[155] vdd gnd cell_6t
Xbit_r156_c194 bl[194] br[194] wl[156] vdd gnd cell_6t
Xbit_r157_c194 bl[194] br[194] wl[157] vdd gnd cell_6t
Xbit_r158_c194 bl[194] br[194] wl[158] vdd gnd cell_6t
Xbit_r159_c194 bl[194] br[194] wl[159] vdd gnd cell_6t
Xbit_r160_c194 bl[194] br[194] wl[160] vdd gnd cell_6t
Xbit_r161_c194 bl[194] br[194] wl[161] vdd gnd cell_6t
Xbit_r162_c194 bl[194] br[194] wl[162] vdd gnd cell_6t
Xbit_r163_c194 bl[194] br[194] wl[163] vdd gnd cell_6t
Xbit_r164_c194 bl[194] br[194] wl[164] vdd gnd cell_6t
Xbit_r165_c194 bl[194] br[194] wl[165] vdd gnd cell_6t
Xbit_r166_c194 bl[194] br[194] wl[166] vdd gnd cell_6t
Xbit_r167_c194 bl[194] br[194] wl[167] vdd gnd cell_6t
Xbit_r168_c194 bl[194] br[194] wl[168] vdd gnd cell_6t
Xbit_r169_c194 bl[194] br[194] wl[169] vdd gnd cell_6t
Xbit_r170_c194 bl[194] br[194] wl[170] vdd gnd cell_6t
Xbit_r171_c194 bl[194] br[194] wl[171] vdd gnd cell_6t
Xbit_r172_c194 bl[194] br[194] wl[172] vdd gnd cell_6t
Xbit_r173_c194 bl[194] br[194] wl[173] vdd gnd cell_6t
Xbit_r174_c194 bl[194] br[194] wl[174] vdd gnd cell_6t
Xbit_r175_c194 bl[194] br[194] wl[175] vdd gnd cell_6t
Xbit_r176_c194 bl[194] br[194] wl[176] vdd gnd cell_6t
Xbit_r177_c194 bl[194] br[194] wl[177] vdd gnd cell_6t
Xbit_r178_c194 bl[194] br[194] wl[178] vdd gnd cell_6t
Xbit_r179_c194 bl[194] br[194] wl[179] vdd gnd cell_6t
Xbit_r180_c194 bl[194] br[194] wl[180] vdd gnd cell_6t
Xbit_r181_c194 bl[194] br[194] wl[181] vdd gnd cell_6t
Xbit_r182_c194 bl[194] br[194] wl[182] vdd gnd cell_6t
Xbit_r183_c194 bl[194] br[194] wl[183] vdd gnd cell_6t
Xbit_r184_c194 bl[194] br[194] wl[184] vdd gnd cell_6t
Xbit_r185_c194 bl[194] br[194] wl[185] vdd gnd cell_6t
Xbit_r186_c194 bl[194] br[194] wl[186] vdd gnd cell_6t
Xbit_r187_c194 bl[194] br[194] wl[187] vdd gnd cell_6t
Xbit_r188_c194 bl[194] br[194] wl[188] vdd gnd cell_6t
Xbit_r189_c194 bl[194] br[194] wl[189] vdd gnd cell_6t
Xbit_r190_c194 bl[194] br[194] wl[190] vdd gnd cell_6t
Xbit_r191_c194 bl[194] br[194] wl[191] vdd gnd cell_6t
Xbit_r192_c194 bl[194] br[194] wl[192] vdd gnd cell_6t
Xbit_r193_c194 bl[194] br[194] wl[193] vdd gnd cell_6t
Xbit_r194_c194 bl[194] br[194] wl[194] vdd gnd cell_6t
Xbit_r195_c194 bl[194] br[194] wl[195] vdd gnd cell_6t
Xbit_r196_c194 bl[194] br[194] wl[196] vdd gnd cell_6t
Xbit_r197_c194 bl[194] br[194] wl[197] vdd gnd cell_6t
Xbit_r198_c194 bl[194] br[194] wl[198] vdd gnd cell_6t
Xbit_r199_c194 bl[194] br[194] wl[199] vdd gnd cell_6t
Xbit_r200_c194 bl[194] br[194] wl[200] vdd gnd cell_6t
Xbit_r201_c194 bl[194] br[194] wl[201] vdd gnd cell_6t
Xbit_r202_c194 bl[194] br[194] wl[202] vdd gnd cell_6t
Xbit_r203_c194 bl[194] br[194] wl[203] vdd gnd cell_6t
Xbit_r204_c194 bl[194] br[194] wl[204] vdd gnd cell_6t
Xbit_r205_c194 bl[194] br[194] wl[205] vdd gnd cell_6t
Xbit_r206_c194 bl[194] br[194] wl[206] vdd gnd cell_6t
Xbit_r207_c194 bl[194] br[194] wl[207] vdd gnd cell_6t
Xbit_r208_c194 bl[194] br[194] wl[208] vdd gnd cell_6t
Xbit_r209_c194 bl[194] br[194] wl[209] vdd gnd cell_6t
Xbit_r210_c194 bl[194] br[194] wl[210] vdd gnd cell_6t
Xbit_r211_c194 bl[194] br[194] wl[211] vdd gnd cell_6t
Xbit_r212_c194 bl[194] br[194] wl[212] vdd gnd cell_6t
Xbit_r213_c194 bl[194] br[194] wl[213] vdd gnd cell_6t
Xbit_r214_c194 bl[194] br[194] wl[214] vdd gnd cell_6t
Xbit_r215_c194 bl[194] br[194] wl[215] vdd gnd cell_6t
Xbit_r216_c194 bl[194] br[194] wl[216] vdd gnd cell_6t
Xbit_r217_c194 bl[194] br[194] wl[217] vdd gnd cell_6t
Xbit_r218_c194 bl[194] br[194] wl[218] vdd gnd cell_6t
Xbit_r219_c194 bl[194] br[194] wl[219] vdd gnd cell_6t
Xbit_r220_c194 bl[194] br[194] wl[220] vdd gnd cell_6t
Xbit_r221_c194 bl[194] br[194] wl[221] vdd gnd cell_6t
Xbit_r222_c194 bl[194] br[194] wl[222] vdd gnd cell_6t
Xbit_r223_c194 bl[194] br[194] wl[223] vdd gnd cell_6t
Xbit_r224_c194 bl[194] br[194] wl[224] vdd gnd cell_6t
Xbit_r225_c194 bl[194] br[194] wl[225] vdd gnd cell_6t
Xbit_r226_c194 bl[194] br[194] wl[226] vdd gnd cell_6t
Xbit_r227_c194 bl[194] br[194] wl[227] vdd gnd cell_6t
Xbit_r228_c194 bl[194] br[194] wl[228] vdd gnd cell_6t
Xbit_r229_c194 bl[194] br[194] wl[229] vdd gnd cell_6t
Xbit_r230_c194 bl[194] br[194] wl[230] vdd gnd cell_6t
Xbit_r231_c194 bl[194] br[194] wl[231] vdd gnd cell_6t
Xbit_r232_c194 bl[194] br[194] wl[232] vdd gnd cell_6t
Xbit_r233_c194 bl[194] br[194] wl[233] vdd gnd cell_6t
Xbit_r234_c194 bl[194] br[194] wl[234] vdd gnd cell_6t
Xbit_r235_c194 bl[194] br[194] wl[235] vdd gnd cell_6t
Xbit_r236_c194 bl[194] br[194] wl[236] vdd gnd cell_6t
Xbit_r237_c194 bl[194] br[194] wl[237] vdd gnd cell_6t
Xbit_r238_c194 bl[194] br[194] wl[238] vdd gnd cell_6t
Xbit_r239_c194 bl[194] br[194] wl[239] vdd gnd cell_6t
Xbit_r240_c194 bl[194] br[194] wl[240] vdd gnd cell_6t
Xbit_r241_c194 bl[194] br[194] wl[241] vdd gnd cell_6t
Xbit_r242_c194 bl[194] br[194] wl[242] vdd gnd cell_6t
Xbit_r243_c194 bl[194] br[194] wl[243] vdd gnd cell_6t
Xbit_r244_c194 bl[194] br[194] wl[244] vdd gnd cell_6t
Xbit_r245_c194 bl[194] br[194] wl[245] vdd gnd cell_6t
Xbit_r246_c194 bl[194] br[194] wl[246] vdd gnd cell_6t
Xbit_r247_c194 bl[194] br[194] wl[247] vdd gnd cell_6t
Xbit_r248_c194 bl[194] br[194] wl[248] vdd gnd cell_6t
Xbit_r249_c194 bl[194] br[194] wl[249] vdd gnd cell_6t
Xbit_r250_c194 bl[194] br[194] wl[250] vdd gnd cell_6t
Xbit_r251_c194 bl[194] br[194] wl[251] vdd gnd cell_6t
Xbit_r252_c194 bl[194] br[194] wl[252] vdd gnd cell_6t
Xbit_r253_c194 bl[194] br[194] wl[253] vdd gnd cell_6t
Xbit_r254_c194 bl[194] br[194] wl[254] vdd gnd cell_6t
Xbit_r255_c194 bl[194] br[194] wl[255] vdd gnd cell_6t
Xbit_r0_c195 bl[195] br[195] wl[0] vdd gnd cell_6t
Xbit_r1_c195 bl[195] br[195] wl[1] vdd gnd cell_6t
Xbit_r2_c195 bl[195] br[195] wl[2] vdd gnd cell_6t
Xbit_r3_c195 bl[195] br[195] wl[3] vdd gnd cell_6t
Xbit_r4_c195 bl[195] br[195] wl[4] vdd gnd cell_6t
Xbit_r5_c195 bl[195] br[195] wl[5] vdd gnd cell_6t
Xbit_r6_c195 bl[195] br[195] wl[6] vdd gnd cell_6t
Xbit_r7_c195 bl[195] br[195] wl[7] vdd gnd cell_6t
Xbit_r8_c195 bl[195] br[195] wl[8] vdd gnd cell_6t
Xbit_r9_c195 bl[195] br[195] wl[9] vdd gnd cell_6t
Xbit_r10_c195 bl[195] br[195] wl[10] vdd gnd cell_6t
Xbit_r11_c195 bl[195] br[195] wl[11] vdd gnd cell_6t
Xbit_r12_c195 bl[195] br[195] wl[12] vdd gnd cell_6t
Xbit_r13_c195 bl[195] br[195] wl[13] vdd gnd cell_6t
Xbit_r14_c195 bl[195] br[195] wl[14] vdd gnd cell_6t
Xbit_r15_c195 bl[195] br[195] wl[15] vdd gnd cell_6t
Xbit_r16_c195 bl[195] br[195] wl[16] vdd gnd cell_6t
Xbit_r17_c195 bl[195] br[195] wl[17] vdd gnd cell_6t
Xbit_r18_c195 bl[195] br[195] wl[18] vdd gnd cell_6t
Xbit_r19_c195 bl[195] br[195] wl[19] vdd gnd cell_6t
Xbit_r20_c195 bl[195] br[195] wl[20] vdd gnd cell_6t
Xbit_r21_c195 bl[195] br[195] wl[21] vdd gnd cell_6t
Xbit_r22_c195 bl[195] br[195] wl[22] vdd gnd cell_6t
Xbit_r23_c195 bl[195] br[195] wl[23] vdd gnd cell_6t
Xbit_r24_c195 bl[195] br[195] wl[24] vdd gnd cell_6t
Xbit_r25_c195 bl[195] br[195] wl[25] vdd gnd cell_6t
Xbit_r26_c195 bl[195] br[195] wl[26] vdd gnd cell_6t
Xbit_r27_c195 bl[195] br[195] wl[27] vdd gnd cell_6t
Xbit_r28_c195 bl[195] br[195] wl[28] vdd gnd cell_6t
Xbit_r29_c195 bl[195] br[195] wl[29] vdd gnd cell_6t
Xbit_r30_c195 bl[195] br[195] wl[30] vdd gnd cell_6t
Xbit_r31_c195 bl[195] br[195] wl[31] vdd gnd cell_6t
Xbit_r32_c195 bl[195] br[195] wl[32] vdd gnd cell_6t
Xbit_r33_c195 bl[195] br[195] wl[33] vdd gnd cell_6t
Xbit_r34_c195 bl[195] br[195] wl[34] vdd gnd cell_6t
Xbit_r35_c195 bl[195] br[195] wl[35] vdd gnd cell_6t
Xbit_r36_c195 bl[195] br[195] wl[36] vdd gnd cell_6t
Xbit_r37_c195 bl[195] br[195] wl[37] vdd gnd cell_6t
Xbit_r38_c195 bl[195] br[195] wl[38] vdd gnd cell_6t
Xbit_r39_c195 bl[195] br[195] wl[39] vdd gnd cell_6t
Xbit_r40_c195 bl[195] br[195] wl[40] vdd gnd cell_6t
Xbit_r41_c195 bl[195] br[195] wl[41] vdd gnd cell_6t
Xbit_r42_c195 bl[195] br[195] wl[42] vdd gnd cell_6t
Xbit_r43_c195 bl[195] br[195] wl[43] vdd gnd cell_6t
Xbit_r44_c195 bl[195] br[195] wl[44] vdd gnd cell_6t
Xbit_r45_c195 bl[195] br[195] wl[45] vdd gnd cell_6t
Xbit_r46_c195 bl[195] br[195] wl[46] vdd gnd cell_6t
Xbit_r47_c195 bl[195] br[195] wl[47] vdd gnd cell_6t
Xbit_r48_c195 bl[195] br[195] wl[48] vdd gnd cell_6t
Xbit_r49_c195 bl[195] br[195] wl[49] vdd gnd cell_6t
Xbit_r50_c195 bl[195] br[195] wl[50] vdd gnd cell_6t
Xbit_r51_c195 bl[195] br[195] wl[51] vdd gnd cell_6t
Xbit_r52_c195 bl[195] br[195] wl[52] vdd gnd cell_6t
Xbit_r53_c195 bl[195] br[195] wl[53] vdd gnd cell_6t
Xbit_r54_c195 bl[195] br[195] wl[54] vdd gnd cell_6t
Xbit_r55_c195 bl[195] br[195] wl[55] vdd gnd cell_6t
Xbit_r56_c195 bl[195] br[195] wl[56] vdd gnd cell_6t
Xbit_r57_c195 bl[195] br[195] wl[57] vdd gnd cell_6t
Xbit_r58_c195 bl[195] br[195] wl[58] vdd gnd cell_6t
Xbit_r59_c195 bl[195] br[195] wl[59] vdd gnd cell_6t
Xbit_r60_c195 bl[195] br[195] wl[60] vdd gnd cell_6t
Xbit_r61_c195 bl[195] br[195] wl[61] vdd gnd cell_6t
Xbit_r62_c195 bl[195] br[195] wl[62] vdd gnd cell_6t
Xbit_r63_c195 bl[195] br[195] wl[63] vdd gnd cell_6t
Xbit_r64_c195 bl[195] br[195] wl[64] vdd gnd cell_6t
Xbit_r65_c195 bl[195] br[195] wl[65] vdd gnd cell_6t
Xbit_r66_c195 bl[195] br[195] wl[66] vdd gnd cell_6t
Xbit_r67_c195 bl[195] br[195] wl[67] vdd gnd cell_6t
Xbit_r68_c195 bl[195] br[195] wl[68] vdd gnd cell_6t
Xbit_r69_c195 bl[195] br[195] wl[69] vdd gnd cell_6t
Xbit_r70_c195 bl[195] br[195] wl[70] vdd gnd cell_6t
Xbit_r71_c195 bl[195] br[195] wl[71] vdd gnd cell_6t
Xbit_r72_c195 bl[195] br[195] wl[72] vdd gnd cell_6t
Xbit_r73_c195 bl[195] br[195] wl[73] vdd gnd cell_6t
Xbit_r74_c195 bl[195] br[195] wl[74] vdd gnd cell_6t
Xbit_r75_c195 bl[195] br[195] wl[75] vdd gnd cell_6t
Xbit_r76_c195 bl[195] br[195] wl[76] vdd gnd cell_6t
Xbit_r77_c195 bl[195] br[195] wl[77] vdd gnd cell_6t
Xbit_r78_c195 bl[195] br[195] wl[78] vdd gnd cell_6t
Xbit_r79_c195 bl[195] br[195] wl[79] vdd gnd cell_6t
Xbit_r80_c195 bl[195] br[195] wl[80] vdd gnd cell_6t
Xbit_r81_c195 bl[195] br[195] wl[81] vdd gnd cell_6t
Xbit_r82_c195 bl[195] br[195] wl[82] vdd gnd cell_6t
Xbit_r83_c195 bl[195] br[195] wl[83] vdd gnd cell_6t
Xbit_r84_c195 bl[195] br[195] wl[84] vdd gnd cell_6t
Xbit_r85_c195 bl[195] br[195] wl[85] vdd gnd cell_6t
Xbit_r86_c195 bl[195] br[195] wl[86] vdd gnd cell_6t
Xbit_r87_c195 bl[195] br[195] wl[87] vdd gnd cell_6t
Xbit_r88_c195 bl[195] br[195] wl[88] vdd gnd cell_6t
Xbit_r89_c195 bl[195] br[195] wl[89] vdd gnd cell_6t
Xbit_r90_c195 bl[195] br[195] wl[90] vdd gnd cell_6t
Xbit_r91_c195 bl[195] br[195] wl[91] vdd gnd cell_6t
Xbit_r92_c195 bl[195] br[195] wl[92] vdd gnd cell_6t
Xbit_r93_c195 bl[195] br[195] wl[93] vdd gnd cell_6t
Xbit_r94_c195 bl[195] br[195] wl[94] vdd gnd cell_6t
Xbit_r95_c195 bl[195] br[195] wl[95] vdd gnd cell_6t
Xbit_r96_c195 bl[195] br[195] wl[96] vdd gnd cell_6t
Xbit_r97_c195 bl[195] br[195] wl[97] vdd gnd cell_6t
Xbit_r98_c195 bl[195] br[195] wl[98] vdd gnd cell_6t
Xbit_r99_c195 bl[195] br[195] wl[99] vdd gnd cell_6t
Xbit_r100_c195 bl[195] br[195] wl[100] vdd gnd cell_6t
Xbit_r101_c195 bl[195] br[195] wl[101] vdd gnd cell_6t
Xbit_r102_c195 bl[195] br[195] wl[102] vdd gnd cell_6t
Xbit_r103_c195 bl[195] br[195] wl[103] vdd gnd cell_6t
Xbit_r104_c195 bl[195] br[195] wl[104] vdd gnd cell_6t
Xbit_r105_c195 bl[195] br[195] wl[105] vdd gnd cell_6t
Xbit_r106_c195 bl[195] br[195] wl[106] vdd gnd cell_6t
Xbit_r107_c195 bl[195] br[195] wl[107] vdd gnd cell_6t
Xbit_r108_c195 bl[195] br[195] wl[108] vdd gnd cell_6t
Xbit_r109_c195 bl[195] br[195] wl[109] vdd gnd cell_6t
Xbit_r110_c195 bl[195] br[195] wl[110] vdd gnd cell_6t
Xbit_r111_c195 bl[195] br[195] wl[111] vdd gnd cell_6t
Xbit_r112_c195 bl[195] br[195] wl[112] vdd gnd cell_6t
Xbit_r113_c195 bl[195] br[195] wl[113] vdd gnd cell_6t
Xbit_r114_c195 bl[195] br[195] wl[114] vdd gnd cell_6t
Xbit_r115_c195 bl[195] br[195] wl[115] vdd gnd cell_6t
Xbit_r116_c195 bl[195] br[195] wl[116] vdd gnd cell_6t
Xbit_r117_c195 bl[195] br[195] wl[117] vdd gnd cell_6t
Xbit_r118_c195 bl[195] br[195] wl[118] vdd gnd cell_6t
Xbit_r119_c195 bl[195] br[195] wl[119] vdd gnd cell_6t
Xbit_r120_c195 bl[195] br[195] wl[120] vdd gnd cell_6t
Xbit_r121_c195 bl[195] br[195] wl[121] vdd gnd cell_6t
Xbit_r122_c195 bl[195] br[195] wl[122] vdd gnd cell_6t
Xbit_r123_c195 bl[195] br[195] wl[123] vdd gnd cell_6t
Xbit_r124_c195 bl[195] br[195] wl[124] vdd gnd cell_6t
Xbit_r125_c195 bl[195] br[195] wl[125] vdd gnd cell_6t
Xbit_r126_c195 bl[195] br[195] wl[126] vdd gnd cell_6t
Xbit_r127_c195 bl[195] br[195] wl[127] vdd gnd cell_6t
Xbit_r128_c195 bl[195] br[195] wl[128] vdd gnd cell_6t
Xbit_r129_c195 bl[195] br[195] wl[129] vdd gnd cell_6t
Xbit_r130_c195 bl[195] br[195] wl[130] vdd gnd cell_6t
Xbit_r131_c195 bl[195] br[195] wl[131] vdd gnd cell_6t
Xbit_r132_c195 bl[195] br[195] wl[132] vdd gnd cell_6t
Xbit_r133_c195 bl[195] br[195] wl[133] vdd gnd cell_6t
Xbit_r134_c195 bl[195] br[195] wl[134] vdd gnd cell_6t
Xbit_r135_c195 bl[195] br[195] wl[135] vdd gnd cell_6t
Xbit_r136_c195 bl[195] br[195] wl[136] vdd gnd cell_6t
Xbit_r137_c195 bl[195] br[195] wl[137] vdd gnd cell_6t
Xbit_r138_c195 bl[195] br[195] wl[138] vdd gnd cell_6t
Xbit_r139_c195 bl[195] br[195] wl[139] vdd gnd cell_6t
Xbit_r140_c195 bl[195] br[195] wl[140] vdd gnd cell_6t
Xbit_r141_c195 bl[195] br[195] wl[141] vdd gnd cell_6t
Xbit_r142_c195 bl[195] br[195] wl[142] vdd gnd cell_6t
Xbit_r143_c195 bl[195] br[195] wl[143] vdd gnd cell_6t
Xbit_r144_c195 bl[195] br[195] wl[144] vdd gnd cell_6t
Xbit_r145_c195 bl[195] br[195] wl[145] vdd gnd cell_6t
Xbit_r146_c195 bl[195] br[195] wl[146] vdd gnd cell_6t
Xbit_r147_c195 bl[195] br[195] wl[147] vdd gnd cell_6t
Xbit_r148_c195 bl[195] br[195] wl[148] vdd gnd cell_6t
Xbit_r149_c195 bl[195] br[195] wl[149] vdd gnd cell_6t
Xbit_r150_c195 bl[195] br[195] wl[150] vdd gnd cell_6t
Xbit_r151_c195 bl[195] br[195] wl[151] vdd gnd cell_6t
Xbit_r152_c195 bl[195] br[195] wl[152] vdd gnd cell_6t
Xbit_r153_c195 bl[195] br[195] wl[153] vdd gnd cell_6t
Xbit_r154_c195 bl[195] br[195] wl[154] vdd gnd cell_6t
Xbit_r155_c195 bl[195] br[195] wl[155] vdd gnd cell_6t
Xbit_r156_c195 bl[195] br[195] wl[156] vdd gnd cell_6t
Xbit_r157_c195 bl[195] br[195] wl[157] vdd gnd cell_6t
Xbit_r158_c195 bl[195] br[195] wl[158] vdd gnd cell_6t
Xbit_r159_c195 bl[195] br[195] wl[159] vdd gnd cell_6t
Xbit_r160_c195 bl[195] br[195] wl[160] vdd gnd cell_6t
Xbit_r161_c195 bl[195] br[195] wl[161] vdd gnd cell_6t
Xbit_r162_c195 bl[195] br[195] wl[162] vdd gnd cell_6t
Xbit_r163_c195 bl[195] br[195] wl[163] vdd gnd cell_6t
Xbit_r164_c195 bl[195] br[195] wl[164] vdd gnd cell_6t
Xbit_r165_c195 bl[195] br[195] wl[165] vdd gnd cell_6t
Xbit_r166_c195 bl[195] br[195] wl[166] vdd gnd cell_6t
Xbit_r167_c195 bl[195] br[195] wl[167] vdd gnd cell_6t
Xbit_r168_c195 bl[195] br[195] wl[168] vdd gnd cell_6t
Xbit_r169_c195 bl[195] br[195] wl[169] vdd gnd cell_6t
Xbit_r170_c195 bl[195] br[195] wl[170] vdd gnd cell_6t
Xbit_r171_c195 bl[195] br[195] wl[171] vdd gnd cell_6t
Xbit_r172_c195 bl[195] br[195] wl[172] vdd gnd cell_6t
Xbit_r173_c195 bl[195] br[195] wl[173] vdd gnd cell_6t
Xbit_r174_c195 bl[195] br[195] wl[174] vdd gnd cell_6t
Xbit_r175_c195 bl[195] br[195] wl[175] vdd gnd cell_6t
Xbit_r176_c195 bl[195] br[195] wl[176] vdd gnd cell_6t
Xbit_r177_c195 bl[195] br[195] wl[177] vdd gnd cell_6t
Xbit_r178_c195 bl[195] br[195] wl[178] vdd gnd cell_6t
Xbit_r179_c195 bl[195] br[195] wl[179] vdd gnd cell_6t
Xbit_r180_c195 bl[195] br[195] wl[180] vdd gnd cell_6t
Xbit_r181_c195 bl[195] br[195] wl[181] vdd gnd cell_6t
Xbit_r182_c195 bl[195] br[195] wl[182] vdd gnd cell_6t
Xbit_r183_c195 bl[195] br[195] wl[183] vdd gnd cell_6t
Xbit_r184_c195 bl[195] br[195] wl[184] vdd gnd cell_6t
Xbit_r185_c195 bl[195] br[195] wl[185] vdd gnd cell_6t
Xbit_r186_c195 bl[195] br[195] wl[186] vdd gnd cell_6t
Xbit_r187_c195 bl[195] br[195] wl[187] vdd gnd cell_6t
Xbit_r188_c195 bl[195] br[195] wl[188] vdd gnd cell_6t
Xbit_r189_c195 bl[195] br[195] wl[189] vdd gnd cell_6t
Xbit_r190_c195 bl[195] br[195] wl[190] vdd gnd cell_6t
Xbit_r191_c195 bl[195] br[195] wl[191] vdd gnd cell_6t
Xbit_r192_c195 bl[195] br[195] wl[192] vdd gnd cell_6t
Xbit_r193_c195 bl[195] br[195] wl[193] vdd gnd cell_6t
Xbit_r194_c195 bl[195] br[195] wl[194] vdd gnd cell_6t
Xbit_r195_c195 bl[195] br[195] wl[195] vdd gnd cell_6t
Xbit_r196_c195 bl[195] br[195] wl[196] vdd gnd cell_6t
Xbit_r197_c195 bl[195] br[195] wl[197] vdd gnd cell_6t
Xbit_r198_c195 bl[195] br[195] wl[198] vdd gnd cell_6t
Xbit_r199_c195 bl[195] br[195] wl[199] vdd gnd cell_6t
Xbit_r200_c195 bl[195] br[195] wl[200] vdd gnd cell_6t
Xbit_r201_c195 bl[195] br[195] wl[201] vdd gnd cell_6t
Xbit_r202_c195 bl[195] br[195] wl[202] vdd gnd cell_6t
Xbit_r203_c195 bl[195] br[195] wl[203] vdd gnd cell_6t
Xbit_r204_c195 bl[195] br[195] wl[204] vdd gnd cell_6t
Xbit_r205_c195 bl[195] br[195] wl[205] vdd gnd cell_6t
Xbit_r206_c195 bl[195] br[195] wl[206] vdd gnd cell_6t
Xbit_r207_c195 bl[195] br[195] wl[207] vdd gnd cell_6t
Xbit_r208_c195 bl[195] br[195] wl[208] vdd gnd cell_6t
Xbit_r209_c195 bl[195] br[195] wl[209] vdd gnd cell_6t
Xbit_r210_c195 bl[195] br[195] wl[210] vdd gnd cell_6t
Xbit_r211_c195 bl[195] br[195] wl[211] vdd gnd cell_6t
Xbit_r212_c195 bl[195] br[195] wl[212] vdd gnd cell_6t
Xbit_r213_c195 bl[195] br[195] wl[213] vdd gnd cell_6t
Xbit_r214_c195 bl[195] br[195] wl[214] vdd gnd cell_6t
Xbit_r215_c195 bl[195] br[195] wl[215] vdd gnd cell_6t
Xbit_r216_c195 bl[195] br[195] wl[216] vdd gnd cell_6t
Xbit_r217_c195 bl[195] br[195] wl[217] vdd gnd cell_6t
Xbit_r218_c195 bl[195] br[195] wl[218] vdd gnd cell_6t
Xbit_r219_c195 bl[195] br[195] wl[219] vdd gnd cell_6t
Xbit_r220_c195 bl[195] br[195] wl[220] vdd gnd cell_6t
Xbit_r221_c195 bl[195] br[195] wl[221] vdd gnd cell_6t
Xbit_r222_c195 bl[195] br[195] wl[222] vdd gnd cell_6t
Xbit_r223_c195 bl[195] br[195] wl[223] vdd gnd cell_6t
Xbit_r224_c195 bl[195] br[195] wl[224] vdd gnd cell_6t
Xbit_r225_c195 bl[195] br[195] wl[225] vdd gnd cell_6t
Xbit_r226_c195 bl[195] br[195] wl[226] vdd gnd cell_6t
Xbit_r227_c195 bl[195] br[195] wl[227] vdd gnd cell_6t
Xbit_r228_c195 bl[195] br[195] wl[228] vdd gnd cell_6t
Xbit_r229_c195 bl[195] br[195] wl[229] vdd gnd cell_6t
Xbit_r230_c195 bl[195] br[195] wl[230] vdd gnd cell_6t
Xbit_r231_c195 bl[195] br[195] wl[231] vdd gnd cell_6t
Xbit_r232_c195 bl[195] br[195] wl[232] vdd gnd cell_6t
Xbit_r233_c195 bl[195] br[195] wl[233] vdd gnd cell_6t
Xbit_r234_c195 bl[195] br[195] wl[234] vdd gnd cell_6t
Xbit_r235_c195 bl[195] br[195] wl[235] vdd gnd cell_6t
Xbit_r236_c195 bl[195] br[195] wl[236] vdd gnd cell_6t
Xbit_r237_c195 bl[195] br[195] wl[237] vdd gnd cell_6t
Xbit_r238_c195 bl[195] br[195] wl[238] vdd gnd cell_6t
Xbit_r239_c195 bl[195] br[195] wl[239] vdd gnd cell_6t
Xbit_r240_c195 bl[195] br[195] wl[240] vdd gnd cell_6t
Xbit_r241_c195 bl[195] br[195] wl[241] vdd gnd cell_6t
Xbit_r242_c195 bl[195] br[195] wl[242] vdd gnd cell_6t
Xbit_r243_c195 bl[195] br[195] wl[243] vdd gnd cell_6t
Xbit_r244_c195 bl[195] br[195] wl[244] vdd gnd cell_6t
Xbit_r245_c195 bl[195] br[195] wl[245] vdd gnd cell_6t
Xbit_r246_c195 bl[195] br[195] wl[246] vdd gnd cell_6t
Xbit_r247_c195 bl[195] br[195] wl[247] vdd gnd cell_6t
Xbit_r248_c195 bl[195] br[195] wl[248] vdd gnd cell_6t
Xbit_r249_c195 bl[195] br[195] wl[249] vdd gnd cell_6t
Xbit_r250_c195 bl[195] br[195] wl[250] vdd gnd cell_6t
Xbit_r251_c195 bl[195] br[195] wl[251] vdd gnd cell_6t
Xbit_r252_c195 bl[195] br[195] wl[252] vdd gnd cell_6t
Xbit_r253_c195 bl[195] br[195] wl[253] vdd gnd cell_6t
Xbit_r254_c195 bl[195] br[195] wl[254] vdd gnd cell_6t
Xbit_r255_c195 bl[195] br[195] wl[255] vdd gnd cell_6t
Xbit_r0_c196 bl[196] br[196] wl[0] vdd gnd cell_6t
Xbit_r1_c196 bl[196] br[196] wl[1] vdd gnd cell_6t
Xbit_r2_c196 bl[196] br[196] wl[2] vdd gnd cell_6t
Xbit_r3_c196 bl[196] br[196] wl[3] vdd gnd cell_6t
Xbit_r4_c196 bl[196] br[196] wl[4] vdd gnd cell_6t
Xbit_r5_c196 bl[196] br[196] wl[5] vdd gnd cell_6t
Xbit_r6_c196 bl[196] br[196] wl[6] vdd gnd cell_6t
Xbit_r7_c196 bl[196] br[196] wl[7] vdd gnd cell_6t
Xbit_r8_c196 bl[196] br[196] wl[8] vdd gnd cell_6t
Xbit_r9_c196 bl[196] br[196] wl[9] vdd gnd cell_6t
Xbit_r10_c196 bl[196] br[196] wl[10] vdd gnd cell_6t
Xbit_r11_c196 bl[196] br[196] wl[11] vdd gnd cell_6t
Xbit_r12_c196 bl[196] br[196] wl[12] vdd gnd cell_6t
Xbit_r13_c196 bl[196] br[196] wl[13] vdd gnd cell_6t
Xbit_r14_c196 bl[196] br[196] wl[14] vdd gnd cell_6t
Xbit_r15_c196 bl[196] br[196] wl[15] vdd gnd cell_6t
Xbit_r16_c196 bl[196] br[196] wl[16] vdd gnd cell_6t
Xbit_r17_c196 bl[196] br[196] wl[17] vdd gnd cell_6t
Xbit_r18_c196 bl[196] br[196] wl[18] vdd gnd cell_6t
Xbit_r19_c196 bl[196] br[196] wl[19] vdd gnd cell_6t
Xbit_r20_c196 bl[196] br[196] wl[20] vdd gnd cell_6t
Xbit_r21_c196 bl[196] br[196] wl[21] vdd gnd cell_6t
Xbit_r22_c196 bl[196] br[196] wl[22] vdd gnd cell_6t
Xbit_r23_c196 bl[196] br[196] wl[23] vdd gnd cell_6t
Xbit_r24_c196 bl[196] br[196] wl[24] vdd gnd cell_6t
Xbit_r25_c196 bl[196] br[196] wl[25] vdd gnd cell_6t
Xbit_r26_c196 bl[196] br[196] wl[26] vdd gnd cell_6t
Xbit_r27_c196 bl[196] br[196] wl[27] vdd gnd cell_6t
Xbit_r28_c196 bl[196] br[196] wl[28] vdd gnd cell_6t
Xbit_r29_c196 bl[196] br[196] wl[29] vdd gnd cell_6t
Xbit_r30_c196 bl[196] br[196] wl[30] vdd gnd cell_6t
Xbit_r31_c196 bl[196] br[196] wl[31] vdd gnd cell_6t
Xbit_r32_c196 bl[196] br[196] wl[32] vdd gnd cell_6t
Xbit_r33_c196 bl[196] br[196] wl[33] vdd gnd cell_6t
Xbit_r34_c196 bl[196] br[196] wl[34] vdd gnd cell_6t
Xbit_r35_c196 bl[196] br[196] wl[35] vdd gnd cell_6t
Xbit_r36_c196 bl[196] br[196] wl[36] vdd gnd cell_6t
Xbit_r37_c196 bl[196] br[196] wl[37] vdd gnd cell_6t
Xbit_r38_c196 bl[196] br[196] wl[38] vdd gnd cell_6t
Xbit_r39_c196 bl[196] br[196] wl[39] vdd gnd cell_6t
Xbit_r40_c196 bl[196] br[196] wl[40] vdd gnd cell_6t
Xbit_r41_c196 bl[196] br[196] wl[41] vdd gnd cell_6t
Xbit_r42_c196 bl[196] br[196] wl[42] vdd gnd cell_6t
Xbit_r43_c196 bl[196] br[196] wl[43] vdd gnd cell_6t
Xbit_r44_c196 bl[196] br[196] wl[44] vdd gnd cell_6t
Xbit_r45_c196 bl[196] br[196] wl[45] vdd gnd cell_6t
Xbit_r46_c196 bl[196] br[196] wl[46] vdd gnd cell_6t
Xbit_r47_c196 bl[196] br[196] wl[47] vdd gnd cell_6t
Xbit_r48_c196 bl[196] br[196] wl[48] vdd gnd cell_6t
Xbit_r49_c196 bl[196] br[196] wl[49] vdd gnd cell_6t
Xbit_r50_c196 bl[196] br[196] wl[50] vdd gnd cell_6t
Xbit_r51_c196 bl[196] br[196] wl[51] vdd gnd cell_6t
Xbit_r52_c196 bl[196] br[196] wl[52] vdd gnd cell_6t
Xbit_r53_c196 bl[196] br[196] wl[53] vdd gnd cell_6t
Xbit_r54_c196 bl[196] br[196] wl[54] vdd gnd cell_6t
Xbit_r55_c196 bl[196] br[196] wl[55] vdd gnd cell_6t
Xbit_r56_c196 bl[196] br[196] wl[56] vdd gnd cell_6t
Xbit_r57_c196 bl[196] br[196] wl[57] vdd gnd cell_6t
Xbit_r58_c196 bl[196] br[196] wl[58] vdd gnd cell_6t
Xbit_r59_c196 bl[196] br[196] wl[59] vdd gnd cell_6t
Xbit_r60_c196 bl[196] br[196] wl[60] vdd gnd cell_6t
Xbit_r61_c196 bl[196] br[196] wl[61] vdd gnd cell_6t
Xbit_r62_c196 bl[196] br[196] wl[62] vdd gnd cell_6t
Xbit_r63_c196 bl[196] br[196] wl[63] vdd gnd cell_6t
Xbit_r64_c196 bl[196] br[196] wl[64] vdd gnd cell_6t
Xbit_r65_c196 bl[196] br[196] wl[65] vdd gnd cell_6t
Xbit_r66_c196 bl[196] br[196] wl[66] vdd gnd cell_6t
Xbit_r67_c196 bl[196] br[196] wl[67] vdd gnd cell_6t
Xbit_r68_c196 bl[196] br[196] wl[68] vdd gnd cell_6t
Xbit_r69_c196 bl[196] br[196] wl[69] vdd gnd cell_6t
Xbit_r70_c196 bl[196] br[196] wl[70] vdd gnd cell_6t
Xbit_r71_c196 bl[196] br[196] wl[71] vdd gnd cell_6t
Xbit_r72_c196 bl[196] br[196] wl[72] vdd gnd cell_6t
Xbit_r73_c196 bl[196] br[196] wl[73] vdd gnd cell_6t
Xbit_r74_c196 bl[196] br[196] wl[74] vdd gnd cell_6t
Xbit_r75_c196 bl[196] br[196] wl[75] vdd gnd cell_6t
Xbit_r76_c196 bl[196] br[196] wl[76] vdd gnd cell_6t
Xbit_r77_c196 bl[196] br[196] wl[77] vdd gnd cell_6t
Xbit_r78_c196 bl[196] br[196] wl[78] vdd gnd cell_6t
Xbit_r79_c196 bl[196] br[196] wl[79] vdd gnd cell_6t
Xbit_r80_c196 bl[196] br[196] wl[80] vdd gnd cell_6t
Xbit_r81_c196 bl[196] br[196] wl[81] vdd gnd cell_6t
Xbit_r82_c196 bl[196] br[196] wl[82] vdd gnd cell_6t
Xbit_r83_c196 bl[196] br[196] wl[83] vdd gnd cell_6t
Xbit_r84_c196 bl[196] br[196] wl[84] vdd gnd cell_6t
Xbit_r85_c196 bl[196] br[196] wl[85] vdd gnd cell_6t
Xbit_r86_c196 bl[196] br[196] wl[86] vdd gnd cell_6t
Xbit_r87_c196 bl[196] br[196] wl[87] vdd gnd cell_6t
Xbit_r88_c196 bl[196] br[196] wl[88] vdd gnd cell_6t
Xbit_r89_c196 bl[196] br[196] wl[89] vdd gnd cell_6t
Xbit_r90_c196 bl[196] br[196] wl[90] vdd gnd cell_6t
Xbit_r91_c196 bl[196] br[196] wl[91] vdd gnd cell_6t
Xbit_r92_c196 bl[196] br[196] wl[92] vdd gnd cell_6t
Xbit_r93_c196 bl[196] br[196] wl[93] vdd gnd cell_6t
Xbit_r94_c196 bl[196] br[196] wl[94] vdd gnd cell_6t
Xbit_r95_c196 bl[196] br[196] wl[95] vdd gnd cell_6t
Xbit_r96_c196 bl[196] br[196] wl[96] vdd gnd cell_6t
Xbit_r97_c196 bl[196] br[196] wl[97] vdd gnd cell_6t
Xbit_r98_c196 bl[196] br[196] wl[98] vdd gnd cell_6t
Xbit_r99_c196 bl[196] br[196] wl[99] vdd gnd cell_6t
Xbit_r100_c196 bl[196] br[196] wl[100] vdd gnd cell_6t
Xbit_r101_c196 bl[196] br[196] wl[101] vdd gnd cell_6t
Xbit_r102_c196 bl[196] br[196] wl[102] vdd gnd cell_6t
Xbit_r103_c196 bl[196] br[196] wl[103] vdd gnd cell_6t
Xbit_r104_c196 bl[196] br[196] wl[104] vdd gnd cell_6t
Xbit_r105_c196 bl[196] br[196] wl[105] vdd gnd cell_6t
Xbit_r106_c196 bl[196] br[196] wl[106] vdd gnd cell_6t
Xbit_r107_c196 bl[196] br[196] wl[107] vdd gnd cell_6t
Xbit_r108_c196 bl[196] br[196] wl[108] vdd gnd cell_6t
Xbit_r109_c196 bl[196] br[196] wl[109] vdd gnd cell_6t
Xbit_r110_c196 bl[196] br[196] wl[110] vdd gnd cell_6t
Xbit_r111_c196 bl[196] br[196] wl[111] vdd gnd cell_6t
Xbit_r112_c196 bl[196] br[196] wl[112] vdd gnd cell_6t
Xbit_r113_c196 bl[196] br[196] wl[113] vdd gnd cell_6t
Xbit_r114_c196 bl[196] br[196] wl[114] vdd gnd cell_6t
Xbit_r115_c196 bl[196] br[196] wl[115] vdd gnd cell_6t
Xbit_r116_c196 bl[196] br[196] wl[116] vdd gnd cell_6t
Xbit_r117_c196 bl[196] br[196] wl[117] vdd gnd cell_6t
Xbit_r118_c196 bl[196] br[196] wl[118] vdd gnd cell_6t
Xbit_r119_c196 bl[196] br[196] wl[119] vdd gnd cell_6t
Xbit_r120_c196 bl[196] br[196] wl[120] vdd gnd cell_6t
Xbit_r121_c196 bl[196] br[196] wl[121] vdd gnd cell_6t
Xbit_r122_c196 bl[196] br[196] wl[122] vdd gnd cell_6t
Xbit_r123_c196 bl[196] br[196] wl[123] vdd gnd cell_6t
Xbit_r124_c196 bl[196] br[196] wl[124] vdd gnd cell_6t
Xbit_r125_c196 bl[196] br[196] wl[125] vdd gnd cell_6t
Xbit_r126_c196 bl[196] br[196] wl[126] vdd gnd cell_6t
Xbit_r127_c196 bl[196] br[196] wl[127] vdd gnd cell_6t
Xbit_r128_c196 bl[196] br[196] wl[128] vdd gnd cell_6t
Xbit_r129_c196 bl[196] br[196] wl[129] vdd gnd cell_6t
Xbit_r130_c196 bl[196] br[196] wl[130] vdd gnd cell_6t
Xbit_r131_c196 bl[196] br[196] wl[131] vdd gnd cell_6t
Xbit_r132_c196 bl[196] br[196] wl[132] vdd gnd cell_6t
Xbit_r133_c196 bl[196] br[196] wl[133] vdd gnd cell_6t
Xbit_r134_c196 bl[196] br[196] wl[134] vdd gnd cell_6t
Xbit_r135_c196 bl[196] br[196] wl[135] vdd gnd cell_6t
Xbit_r136_c196 bl[196] br[196] wl[136] vdd gnd cell_6t
Xbit_r137_c196 bl[196] br[196] wl[137] vdd gnd cell_6t
Xbit_r138_c196 bl[196] br[196] wl[138] vdd gnd cell_6t
Xbit_r139_c196 bl[196] br[196] wl[139] vdd gnd cell_6t
Xbit_r140_c196 bl[196] br[196] wl[140] vdd gnd cell_6t
Xbit_r141_c196 bl[196] br[196] wl[141] vdd gnd cell_6t
Xbit_r142_c196 bl[196] br[196] wl[142] vdd gnd cell_6t
Xbit_r143_c196 bl[196] br[196] wl[143] vdd gnd cell_6t
Xbit_r144_c196 bl[196] br[196] wl[144] vdd gnd cell_6t
Xbit_r145_c196 bl[196] br[196] wl[145] vdd gnd cell_6t
Xbit_r146_c196 bl[196] br[196] wl[146] vdd gnd cell_6t
Xbit_r147_c196 bl[196] br[196] wl[147] vdd gnd cell_6t
Xbit_r148_c196 bl[196] br[196] wl[148] vdd gnd cell_6t
Xbit_r149_c196 bl[196] br[196] wl[149] vdd gnd cell_6t
Xbit_r150_c196 bl[196] br[196] wl[150] vdd gnd cell_6t
Xbit_r151_c196 bl[196] br[196] wl[151] vdd gnd cell_6t
Xbit_r152_c196 bl[196] br[196] wl[152] vdd gnd cell_6t
Xbit_r153_c196 bl[196] br[196] wl[153] vdd gnd cell_6t
Xbit_r154_c196 bl[196] br[196] wl[154] vdd gnd cell_6t
Xbit_r155_c196 bl[196] br[196] wl[155] vdd gnd cell_6t
Xbit_r156_c196 bl[196] br[196] wl[156] vdd gnd cell_6t
Xbit_r157_c196 bl[196] br[196] wl[157] vdd gnd cell_6t
Xbit_r158_c196 bl[196] br[196] wl[158] vdd gnd cell_6t
Xbit_r159_c196 bl[196] br[196] wl[159] vdd gnd cell_6t
Xbit_r160_c196 bl[196] br[196] wl[160] vdd gnd cell_6t
Xbit_r161_c196 bl[196] br[196] wl[161] vdd gnd cell_6t
Xbit_r162_c196 bl[196] br[196] wl[162] vdd gnd cell_6t
Xbit_r163_c196 bl[196] br[196] wl[163] vdd gnd cell_6t
Xbit_r164_c196 bl[196] br[196] wl[164] vdd gnd cell_6t
Xbit_r165_c196 bl[196] br[196] wl[165] vdd gnd cell_6t
Xbit_r166_c196 bl[196] br[196] wl[166] vdd gnd cell_6t
Xbit_r167_c196 bl[196] br[196] wl[167] vdd gnd cell_6t
Xbit_r168_c196 bl[196] br[196] wl[168] vdd gnd cell_6t
Xbit_r169_c196 bl[196] br[196] wl[169] vdd gnd cell_6t
Xbit_r170_c196 bl[196] br[196] wl[170] vdd gnd cell_6t
Xbit_r171_c196 bl[196] br[196] wl[171] vdd gnd cell_6t
Xbit_r172_c196 bl[196] br[196] wl[172] vdd gnd cell_6t
Xbit_r173_c196 bl[196] br[196] wl[173] vdd gnd cell_6t
Xbit_r174_c196 bl[196] br[196] wl[174] vdd gnd cell_6t
Xbit_r175_c196 bl[196] br[196] wl[175] vdd gnd cell_6t
Xbit_r176_c196 bl[196] br[196] wl[176] vdd gnd cell_6t
Xbit_r177_c196 bl[196] br[196] wl[177] vdd gnd cell_6t
Xbit_r178_c196 bl[196] br[196] wl[178] vdd gnd cell_6t
Xbit_r179_c196 bl[196] br[196] wl[179] vdd gnd cell_6t
Xbit_r180_c196 bl[196] br[196] wl[180] vdd gnd cell_6t
Xbit_r181_c196 bl[196] br[196] wl[181] vdd gnd cell_6t
Xbit_r182_c196 bl[196] br[196] wl[182] vdd gnd cell_6t
Xbit_r183_c196 bl[196] br[196] wl[183] vdd gnd cell_6t
Xbit_r184_c196 bl[196] br[196] wl[184] vdd gnd cell_6t
Xbit_r185_c196 bl[196] br[196] wl[185] vdd gnd cell_6t
Xbit_r186_c196 bl[196] br[196] wl[186] vdd gnd cell_6t
Xbit_r187_c196 bl[196] br[196] wl[187] vdd gnd cell_6t
Xbit_r188_c196 bl[196] br[196] wl[188] vdd gnd cell_6t
Xbit_r189_c196 bl[196] br[196] wl[189] vdd gnd cell_6t
Xbit_r190_c196 bl[196] br[196] wl[190] vdd gnd cell_6t
Xbit_r191_c196 bl[196] br[196] wl[191] vdd gnd cell_6t
Xbit_r192_c196 bl[196] br[196] wl[192] vdd gnd cell_6t
Xbit_r193_c196 bl[196] br[196] wl[193] vdd gnd cell_6t
Xbit_r194_c196 bl[196] br[196] wl[194] vdd gnd cell_6t
Xbit_r195_c196 bl[196] br[196] wl[195] vdd gnd cell_6t
Xbit_r196_c196 bl[196] br[196] wl[196] vdd gnd cell_6t
Xbit_r197_c196 bl[196] br[196] wl[197] vdd gnd cell_6t
Xbit_r198_c196 bl[196] br[196] wl[198] vdd gnd cell_6t
Xbit_r199_c196 bl[196] br[196] wl[199] vdd gnd cell_6t
Xbit_r200_c196 bl[196] br[196] wl[200] vdd gnd cell_6t
Xbit_r201_c196 bl[196] br[196] wl[201] vdd gnd cell_6t
Xbit_r202_c196 bl[196] br[196] wl[202] vdd gnd cell_6t
Xbit_r203_c196 bl[196] br[196] wl[203] vdd gnd cell_6t
Xbit_r204_c196 bl[196] br[196] wl[204] vdd gnd cell_6t
Xbit_r205_c196 bl[196] br[196] wl[205] vdd gnd cell_6t
Xbit_r206_c196 bl[196] br[196] wl[206] vdd gnd cell_6t
Xbit_r207_c196 bl[196] br[196] wl[207] vdd gnd cell_6t
Xbit_r208_c196 bl[196] br[196] wl[208] vdd gnd cell_6t
Xbit_r209_c196 bl[196] br[196] wl[209] vdd gnd cell_6t
Xbit_r210_c196 bl[196] br[196] wl[210] vdd gnd cell_6t
Xbit_r211_c196 bl[196] br[196] wl[211] vdd gnd cell_6t
Xbit_r212_c196 bl[196] br[196] wl[212] vdd gnd cell_6t
Xbit_r213_c196 bl[196] br[196] wl[213] vdd gnd cell_6t
Xbit_r214_c196 bl[196] br[196] wl[214] vdd gnd cell_6t
Xbit_r215_c196 bl[196] br[196] wl[215] vdd gnd cell_6t
Xbit_r216_c196 bl[196] br[196] wl[216] vdd gnd cell_6t
Xbit_r217_c196 bl[196] br[196] wl[217] vdd gnd cell_6t
Xbit_r218_c196 bl[196] br[196] wl[218] vdd gnd cell_6t
Xbit_r219_c196 bl[196] br[196] wl[219] vdd gnd cell_6t
Xbit_r220_c196 bl[196] br[196] wl[220] vdd gnd cell_6t
Xbit_r221_c196 bl[196] br[196] wl[221] vdd gnd cell_6t
Xbit_r222_c196 bl[196] br[196] wl[222] vdd gnd cell_6t
Xbit_r223_c196 bl[196] br[196] wl[223] vdd gnd cell_6t
Xbit_r224_c196 bl[196] br[196] wl[224] vdd gnd cell_6t
Xbit_r225_c196 bl[196] br[196] wl[225] vdd gnd cell_6t
Xbit_r226_c196 bl[196] br[196] wl[226] vdd gnd cell_6t
Xbit_r227_c196 bl[196] br[196] wl[227] vdd gnd cell_6t
Xbit_r228_c196 bl[196] br[196] wl[228] vdd gnd cell_6t
Xbit_r229_c196 bl[196] br[196] wl[229] vdd gnd cell_6t
Xbit_r230_c196 bl[196] br[196] wl[230] vdd gnd cell_6t
Xbit_r231_c196 bl[196] br[196] wl[231] vdd gnd cell_6t
Xbit_r232_c196 bl[196] br[196] wl[232] vdd gnd cell_6t
Xbit_r233_c196 bl[196] br[196] wl[233] vdd gnd cell_6t
Xbit_r234_c196 bl[196] br[196] wl[234] vdd gnd cell_6t
Xbit_r235_c196 bl[196] br[196] wl[235] vdd gnd cell_6t
Xbit_r236_c196 bl[196] br[196] wl[236] vdd gnd cell_6t
Xbit_r237_c196 bl[196] br[196] wl[237] vdd gnd cell_6t
Xbit_r238_c196 bl[196] br[196] wl[238] vdd gnd cell_6t
Xbit_r239_c196 bl[196] br[196] wl[239] vdd gnd cell_6t
Xbit_r240_c196 bl[196] br[196] wl[240] vdd gnd cell_6t
Xbit_r241_c196 bl[196] br[196] wl[241] vdd gnd cell_6t
Xbit_r242_c196 bl[196] br[196] wl[242] vdd gnd cell_6t
Xbit_r243_c196 bl[196] br[196] wl[243] vdd gnd cell_6t
Xbit_r244_c196 bl[196] br[196] wl[244] vdd gnd cell_6t
Xbit_r245_c196 bl[196] br[196] wl[245] vdd gnd cell_6t
Xbit_r246_c196 bl[196] br[196] wl[246] vdd gnd cell_6t
Xbit_r247_c196 bl[196] br[196] wl[247] vdd gnd cell_6t
Xbit_r248_c196 bl[196] br[196] wl[248] vdd gnd cell_6t
Xbit_r249_c196 bl[196] br[196] wl[249] vdd gnd cell_6t
Xbit_r250_c196 bl[196] br[196] wl[250] vdd gnd cell_6t
Xbit_r251_c196 bl[196] br[196] wl[251] vdd gnd cell_6t
Xbit_r252_c196 bl[196] br[196] wl[252] vdd gnd cell_6t
Xbit_r253_c196 bl[196] br[196] wl[253] vdd gnd cell_6t
Xbit_r254_c196 bl[196] br[196] wl[254] vdd gnd cell_6t
Xbit_r255_c196 bl[196] br[196] wl[255] vdd gnd cell_6t
Xbit_r0_c197 bl[197] br[197] wl[0] vdd gnd cell_6t
Xbit_r1_c197 bl[197] br[197] wl[1] vdd gnd cell_6t
Xbit_r2_c197 bl[197] br[197] wl[2] vdd gnd cell_6t
Xbit_r3_c197 bl[197] br[197] wl[3] vdd gnd cell_6t
Xbit_r4_c197 bl[197] br[197] wl[4] vdd gnd cell_6t
Xbit_r5_c197 bl[197] br[197] wl[5] vdd gnd cell_6t
Xbit_r6_c197 bl[197] br[197] wl[6] vdd gnd cell_6t
Xbit_r7_c197 bl[197] br[197] wl[7] vdd gnd cell_6t
Xbit_r8_c197 bl[197] br[197] wl[8] vdd gnd cell_6t
Xbit_r9_c197 bl[197] br[197] wl[9] vdd gnd cell_6t
Xbit_r10_c197 bl[197] br[197] wl[10] vdd gnd cell_6t
Xbit_r11_c197 bl[197] br[197] wl[11] vdd gnd cell_6t
Xbit_r12_c197 bl[197] br[197] wl[12] vdd gnd cell_6t
Xbit_r13_c197 bl[197] br[197] wl[13] vdd gnd cell_6t
Xbit_r14_c197 bl[197] br[197] wl[14] vdd gnd cell_6t
Xbit_r15_c197 bl[197] br[197] wl[15] vdd gnd cell_6t
Xbit_r16_c197 bl[197] br[197] wl[16] vdd gnd cell_6t
Xbit_r17_c197 bl[197] br[197] wl[17] vdd gnd cell_6t
Xbit_r18_c197 bl[197] br[197] wl[18] vdd gnd cell_6t
Xbit_r19_c197 bl[197] br[197] wl[19] vdd gnd cell_6t
Xbit_r20_c197 bl[197] br[197] wl[20] vdd gnd cell_6t
Xbit_r21_c197 bl[197] br[197] wl[21] vdd gnd cell_6t
Xbit_r22_c197 bl[197] br[197] wl[22] vdd gnd cell_6t
Xbit_r23_c197 bl[197] br[197] wl[23] vdd gnd cell_6t
Xbit_r24_c197 bl[197] br[197] wl[24] vdd gnd cell_6t
Xbit_r25_c197 bl[197] br[197] wl[25] vdd gnd cell_6t
Xbit_r26_c197 bl[197] br[197] wl[26] vdd gnd cell_6t
Xbit_r27_c197 bl[197] br[197] wl[27] vdd gnd cell_6t
Xbit_r28_c197 bl[197] br[197] wl[28] vdd gnd cell_6t
Xbit_r29_c197 bl[197] br[197] wl[29] vdd gnd cell_6t
Xbit_r30_c197 bl[197] br[197] wl[30] vdd gnd cell_6t
Xbit_r31_c197 bl[197] br[197] wl[31] vdd gnd cell_6t
Xbit_r32_c197 bl[197] br[197] wl[32] vdd gnd cell_6t
Xbit_r33_c197 bl[197] br[197] wl[33] vdd gnd cell_6t
Xbit_r34_c197 bl[197] br[197] wl[34] vdd gnd cell_6t
Xbit_r35_c197 bl[197] br[197] wl[35] vdd gnd cell_6t
Xbit_r36_c197 bl[197] br[197] wl[36] vdd gnd cell_6t
Xbit_r37_c197 bl[197] br[197] wl[37] vdd gnd cell_6t
Xbit_r38_c197 bl[197] br[197] wl[38] vdd gnd cell_6t
Xbit_r39_c197 bl[197] br[197] wl[39] vdd gnd cell_6t
Xbit_r40_c197 bl[197] br[197] wl[40] vdd gnd cell_6t
Xbit_r41_c197 bl[197] br[197] wl[41] vdd gnd cell_6t
Xbit_r42_c197 bl[197] br[197] wl[42] vdd gnd cell_6t
Xbit_r43_c197 bl[197] br[197] wl[43] vdd gnd cell_6t
Xbit_r44_c197 bl[197] br[197] wl[44] vdd gnd cell_6t
Xbit_r45_c197 bl[197] br[197] wl[45] vdd gnd cell_6t
Xbit_r46_c197 bl[197] br[197] wl[46] vdd gnd cell_6t
Xbit_r47_c197 bl[197] br[197] wl[47] vdd gnd cell_6t
Xbit_r48_c197 bl[197] br[197] wl[48] vdd gnd cell_6t
Xbit_r49_c197 bl[197] br[197] wl[49] vdd gnd cell_6t
Xbit_r50_c197 bl[197] br[197] wl[50] vdd gnd cell_6t
Xbit_r51_c197 bl[197] br[197] wl[51] vdd gnd cell_6t
Xbit_r52_c197 bl[197] br[197] wl[52] vdd gnd cell_6t
Xbit_r53_c197 bl[197] br[197] wl[53] vdd gnd cell_6t
Xbit_r54_c197 bl[197] br[197] wl[54] vdd gnd cell_6t
Xbit_r55_c197 bl[197] br[197] wl[55] vdd gnd cell_6t
Xbit_r56_c197 bl[197] br[197] wl[56] vdd gnd cell_6t
Xbit_r57_c197 bl[197] br[197] wl[57] vdd gnd cell_6t
Xbit_r58_c197 bl[197] br[197] wl[58] vdd gnd cell_6t
Xbit_r59_c197 bl[197] br[197] wl[59] vdd gnd cell_6t
Xbit_r60_c197 bl[197] br[197] wl[60] vdd gnd cell_6t
Xbit_r61_c197 bl[197] br[197] wl[61] vdd gnd cell_6t
Xbit_r62_c197 bl[197] br[197] wl[62] vdd gnd cell_6t
Xbit_r63_c197 bl[197] br[197] wl[63] vdd gnd cell_6t
Xbit_r64_c197 bl[197] br[197] wl[64] vdd gnd cell_6t
Xbit_r65_c197 bl[197] br[197] wl[65] vdd gnd cell_6t
Xbit_r66_c197 bl[197] br[197] wl[66] vdd gnd cell_6t
Xbit_r67_c197 bl[197] br[197] wl[67] vdd gnd cell_6t
Xbit_r68_c197 bl[197] br[197] wl[68] vdd gnd cell_6t
Xbit_r69_c197 bl[197] br[197] wl[69] vdd gnd cell_6t
Xbit_r70_c197 bl[197] br[197] wl[70] vdd gnd cell_6t
Xbit_r71_c197 bl[197] br[197] wl[71] vdd gnd cell_6t
Xbit_r72_c197 bl[197] br[197] wl[72] vdd gnd cell_6t
Xbit_r73_c197 bl[197] br[197] wl[73] vdd gnd cell_6t
Xbit_r74_c197 bl[197] br[197] wl[74] vdd gnd cell_6t
Xbit_r75_c197 bl[197] br[197] wl[75] vdd gnd cell_6t
Xbit_r76_c197 bl[197] br[197] wl[76] vdd gnd cell_6t
Xbit_r77_c197 bl[197] br[197] wl[77] vdd gnd cell_6t
Xbit_r78_c197 bl[197] br[197] wl[78] vdd gnd cell_6t
Xbit_r79_c197 bl[197] br[197] wl[79] vdd gnd cell_6t
Xbit_r80_c197 bl[197] br[197] wl[80] vdd gnd cell_6t
Xbit_r81_c197 bl[197] br[197] wl[81] vdd gnd cell_6t
Xbit_r82_c197 bl[197] br[197] wl[82] vdd gnd cell_6t
Xbit_r83_c197 bl[197] br[197] wl[83] vdd gnd cell_6t
Xbit_r84_c197 bl[197] br[197] wl[84] vdd gnd cell_6t
Xbit_r85_c197 bl[197] br[197] wl[85] vdd gnd cell_6t
Xbit_r86_c197 bl[197] br[197] wl[86] vdd gnd cell_6t
Xbit_r87_c197 bl[197] br[197] wl[87] vdd gnd cell_6t
Xbit_r88_c197 bl[197] br[197] wl[88] vdd gnd cell_6t
Xbit_r89_c197 bl[197] br[197] wl[89] vdd gnd cell_6t
Xbit_r90_c197 bl[197] br[197] wl[90] vdd gnd cell_6t
Xbit_r91_c197 bl[197] br[197] wl[91] vdd gnd cell_6t
Xbit_r92_c197 bl[197] br[197] wl[92] vdd gnd cell_6t
Xbit_r93_c197 bl[197] br[197] wl[93] vdd gnd cell_6t
Xbit_r94_c197 bl[197] br[197] wl[94] vdd gnd cell_6t
Xbit_r95_c197 bl[197] br[197] wl[95] vdd gnd cell_6t
Xbit_r96_c197 bl[197] br[197] wl[96] vdd gnd cell_6t
Xbit_r97_c197 bl[197] br[197] wl[97] vdd gnd cell_6t
Xbit_r98_c197 bl[197] br[197] wl[98] vdd gnd cell_6t
Xbit_r99_c197 bl[197] br[197] wl[99] vdd gnd cell_6t
Xbit_r100_c197 bl[197] br[197] wl[100] vdd gnd cell_6t
Xbit_r101_c197 bl[197] br[197] wl[101] vdd gnd cell_6t
Xbit_r102_c197 bl[197] br[197] wl[102] vdd gnd cell_6t
Xbit_r103_c197 bl[197] br[197] wl[103] vdd gnd cell_6t
Xbit_r104_c197 bl[197] br[197] wl[104] vdd gnd cell_6t
Xbit_r105_c197 bl[197] br[197] wl[105] vdd gnd cell_6t
Xbit_r106_c197 bl[197] br[197] wl[106] vdd gnd cell_6t
Xbit_r107_c197 bl[197] br[197] wl[107] vdd gnd cell_6t
Xbit_r108_c197 bl[197] br[197] wl[108] vdd gnd cell_6t
Xbit_r109_c197 bl[197] br[197] wl[109] vdd gnd cell_6t
Xbit_r110_c197 bl[197] br[197] wl[110] vdd gnd cell_6t
Xbit_r111_c197 bl[197] br[197] wl[111] vdd gnd cell_6t
Xbit_r112_c197 bl[197] br[197] wl[112] vdd gnd cell_6t
Xbit_r113_c197 bl[197] br[197] wl[113] vdd gnd cell_6t
Xbit_r114_c197 bl[197] br[197] wl[114] vdd gnd cell_6t
Xbit_r115_c197 bl[197] br[197] wl[115] vdd gnd cell_6t
Xbit_r116_c197 bl[197] br[197] wl[116] vdd gnd cell_6t
Xbit_r117_c197 bl[197] br[197] wl[117] vdd gnd cell_6t
Xbit_r118_c197 bl[197] br[197] wl[118] vdd gnd cell_6t
Xbit_r119_c197 bl[197] br[197] wl[119] vdd gnd cell_6t
Xbit_r120_c197 bl[197] br[197] wl[120] vdd gnd cell_6t
Xbit_r121_c197 bl[197] br[197] wl[121] vdd gnd cell_6t
Xbit_r122_c197 bl[197] br[197] wl[122] vdd gnd cell_6t
Xbit_r123_c197 bl[197] br[197] wl[123] vdd gnd cell_6t
Xbit_r124_c197 bl[197] br[197] wl[124] vdd gnd cell_6t
Xbit_r125_c197 bl[197] br[197] wl[125] vdd gnd cell_6t
Xbit_r126_c197 bl[197] br[197] wl[126] vdd gnd cell_6t
Xbit_r127_c197 bl[197] br[197] wl[127] vdd gnd cell_6t
Xbit_r128_c197 bl[197] br[197] wl[128] vdd gnd cell_6t
Xbit_r129_c197 bl[197] br[197] wl[129] vdd gnd cell_6t
Xbit_r130_c197 bl[197] br[197] wl[130] vdd gnd cell_6t
Xbit_r131_c197 bl[197] br[197] wl[131] vdd gnd cell_6t
Xbit_r132_c197 bl[197] br[197] wl[132] vdd gnd cell_6t
Xbit_r133_c197 bl[197] br[197] wl[133] vdd gnd cell_6t
Xbit_r134_c197 bl[197] br[197] wl[134] vdd gnd cell_6t
Xbit_r135_c197 bl[197] br[197] wl[135] vdd gnd cell_6t
Xbit_r136_c197 bl[197] br[197] wl[136] vdd gnd cell_6t
Xbit_r137_c197 bl[197] br[197] wl[137] vdd gnd cell_6t
Xbit_r138_c197 bl[197] br[197] wl[138] vdd gnd cell_6t
Xbit_r139_c197 bl[197] br[197] wl[139] vdd gnd cell_6t
Xbit_r140_c197 bl[197] br[197] wl[140] vdd gnd cell_6t
Xbit_r141_c197 bl[197] br[197] wl[141] vdd gnd cell_6t
Xbit_r142_c197 bl[197] br[197] wl[142] vdd gnd cell_6t
Xbit_r143_c197 bl[197] br[197] wl[143] vdd gnd cell_6t
Xbit_r144_c197 bl[197] br[197] wl[144] vdd gnd cell_6t
Xbit_r145_c197 bl[197] br[197] wl[145] vdd gnd cell_6t
Xbit_r146_c197 bl[197] br[197] wl[146] vdd gnd cell_6t
Xbit_r147_c197 bl[197] br[197] wl[147] vdd gnd cell_6t
Xbit_r148_c197 bl[197] br[197] wl[148] vdd gnd cell_6t
Xbit_r149_c197 bl[197] br[197] wl[149] vdd gnd cell_6t
Xbit_r150_c197 bl[197] br[197] wl[150] vdd gnd cell_6t
Xbit_r151_c197 bl[197] br[197] wl[151] vdd gnd cell_6t
Xbit_r152_c197 bl[197] br[197] wl[152] vdd gnd cell_6t
Xbit_r153_c197 bl[197] br[197] wl[153] vdd gnd cell_6t
Xbit_r154_c197 bl[197] br[197] wl[154] vdd gnd cell_6t
Xbit_r155_c197 bl[197] br[197] wl[155] vdd gnd cell_6t
Xbit_r156_c197 bl[197] br[197] wl[156] vdd gnd cell_6t
Xbit_r157_c197 bl[197] br[197] wl[157] vdd gnd cell_6t
Xbit_r158_c197 bl[197] br[197] wl[158] vdd gnd cell_6t
Xbit_r159_c197 bl[197] br[197] wl[159] vdd gnd cell_6t
Xbit_r160_c197 bl[197] br[197] wl[160] vdd gnd cell_6t
Xbit_r161_c197 bl[197] br[197] wl[161] vdd gnd cell_6t
Xbit_r162_c197 bl[197] br[197] wl[162] vdd gnd cell_6t
Xbit_r163_c197 bl[197] br[197] wl[163] vdd gnd cell_6t
Xbit_r164_c197 bl[197] br[197] wl[164] vdd gnd cell_6t
Xbit_r165_c197 bl[197] br[197] wl[165] vdd gnd cell_6t
Xbit_r166_c197 bl[197] br[197] wl[166] vdd gnd cell_6t
Xbit_r167_c197 bl[197] br[197] wl[167] vdd gnd cell_6t
Xbit_r168_c197 bl[197] br[197] wl[168] vdd gnd cell_6t
Xbit_r169_c197 bl[197] br[197] wl[169] vdd gnd cell_6t
Xbit_r170_c197 bl[197] br[197] wl[170] vdd gnd cell_6t
Xbit_r171_c197 bl[197] br[197] wl[171] vdd gnd cell_6t
Xbit_r172_c197 bl[197] br[197] wl[172] vdd gnd cell_6t
Xbit_r173_c197 bl[197] br[197] wl[173] vdd gnd cell_6t
Xbit_r174_c197 bl[197] br[197] wl[174] vdd gnd cell_6t
Xbit_r175_c197 bl[197] br[197] wl[175] vdd gnd cell_6t
Xbit_r176_c197 bl[197] br[197] wl[176] vdd gnd cell_6t
Xbit_r177_c197 bl[197] br[197] wl[177] vdd gnd cell_6t
Xbit_r178_c197 bl[197] br[197] wl[178] vdd gnd cell_6t
Xbit_r179_c197 bl[197] br[197] wl[179] vdd gnd cell_6t
Xbit_r180_c197 bl[197] br[197] wl[180] vdd gnd cell_6t
Xbit_r181_c197 bl[197] br[197] wl[181] vdd gnd cell_6t
Xbit_r182_c197 bl[197] br[197] wl[182] vdd gnd cell_6t
Xbit_r183_c197 bl[197] br[197] wl[183] vdd gnd cell_6t
Xbit_r184_c197 bl[197] br[197] wl[184] vdd gnd cell_6t
Xbit_r185_c197 bl[197] br[197] wl[185] vdd gnd cell_6t
Xbit_r186_c197 bl[197] br[197] wl[186] vdd gnd cell_6t
Xbit_r187_c197 bl[197] br[197] wl[187] vdd gnd cell_6t
Xbit_r188_c197 bl[197] br[197] wl[188] vdd gnd cell_6t
Xbit_r189_c197 bl[197] br[197] wl[189] vdd gnd cell_6t
Xbit_r190_c197 bl[197] br[197] wl[190] vdd gnd cell_6t
Xbit_r191_c197 bl[197] br[197] wl[191] vdd gnd cell_6t
Xbit_r192_c197 bl[197] br[197] wl[192] vdd gnd cell_6t
Xbit_r193_c197 bl[197] br[197] wl[193] vdd gnd cell_6t
Xbit_r194_c197 bl[197] br[197] wl[194] vdd gnd cell_6t
Xbit_r195_c197 bl[197] br[197] wl[195] vdd gnd cell_6t
Xbit_r196_c197 bl[197] br[197] wl[196] vdd gnd cell_6t
Xbit_r197_c197 bl[197] br[197] wl[197] vdd gnd cell_6t
Xbit_r198_c197 bl[197] br[197] wl[198] vdd gnd cell_6t
Xbit_r199_c197 bl[197] br[197] wl[199] vdd gnd cell_6t
Xbit_r200_c197 bl[197] br[197] wl[200] vdd gnd cell_6t
Xbit_r201_c197 bl[197] br[197] wl[201] vdd gnd cell_6t
Xbit_r202_c197 bl[197] br[197] wl[202] vdd gnd cell_6t
Xbit_r203_c197 bl[197] br[197] wl[203] vdd gnd cell_6t
Xbit_r204_c197 bl[197] br[197] wl[204] vdd gnd cell_6t
Xbit_r205_c197 bl[197] br[197] wl[205] vdd gnd cell_6t
Xbit_r206_c197 bl[197] br[197] wl[206] vdd gnd cell_6t
Xbit_r207_c197 bl[197] br[197] wl[207] vdd gnd cell_6t
Xbit_r208_c197 bl[197] br[197] wl[208] vdd gnd cell_6t
Xbit_r209_c197 bl[197] br[197] wl[209] vdd gnd cell_6t
Xbit_r210_c197 bl[197] br[197] wl[210] vdd gnd cell_6t
Xbit_r211_c197 bl[197] br[197] wl[211] vdd gnd cell_6t
Xbit_r212_c197 bl[197] br[197] wl[212] vdd gnd cell_6t
Xbit_r213_c197 bl[197] br[197] wl[213] vdd gnd cell_6t
Xbit_r214_c197 bl[197] br[197] wl[214] vdd gnd cell_6t
Xbit_r215_c197 bl[197] br[197] wl[215] vdd gnd cell_6t
Xbit_r216_c197 bl[197] br[197] wl[216] vdd gnd cell_6t
Xbit_r217_c197 bl[197] br[197] wl[217] vdd gnd cell_6t
Xbit_r218_c197 bl[197] br[197] wl[218] vdd gnd cell_6t
Xbit_r219_c197 bl[197] br[197] wl[219] vdd gnd cell_6t
Xbit_r220_c197 bl[197] br[197] wl[220] vdd gnd cell_6t
Xbit_r221_c197 bl[197] br[197] wl[221] vdd gnd cell_6t
Xbit_r222_c197 bl[197] br[197] wl[222] vdd gnd cell_6t
Xbit_r223_c197 bl[197] br[197] wl[223] vdd gnd cell_6t
Xbit_r224_c197 bl[197] br[197] wl[224] vdd gnd cell_6t
Xbit_r225_c197 bl[197] br[197] wl[225] vdd gnd cell_6t
Xbit_r226_c197 bl[197] br[197] wl[226] vdd gnd cell_6t
Xbit_r227_c197 bl[197] br[197] wl[227] vdd gnd cell_6t
Xbit_r228_c197 bl[197] br[197] wl[228] vdd gnd cell_6t
Xbit_r229_c197 bl[197] br[197] wl[229] vdd gnd cell_6t
Xbit_r230_c197 bl[197] br[197] wl[230] vdd gnd cell_6t
Xbit_r231_c197 bl[197] br[197] wl[231] vdd gnd cell_6t
Xbit_r232_c197 bl[197] br[197] wl[232] vdd gnd cell_6t
Xbit_r233_c197 bl[197] br[197] wl[233] vdd gnd cell_6t
Xbit_r234_c197 bl[197] br[197] wl[234] vdd gnd cell_6t
Xbit_r235_c197 bl[197] br[197] wl[235] vdd gnd cell_6t
Xbit_r236_c197 bl[197] br[197] wl[236] vdd gnd cell_6t
Xbit_r237_c197 bl[197] br[197] wl[237] vdd gnd cell_6t
Xbit_r238_c197 bl[197] br[197] wl[238] vdd gnd cell_6t
Xbit_r239_c197 bl[197] br[197] wl[239] vdd gnd cell_6t
Xbit_r240_c197 bl[197] br[197] wl[240] vdd gnd cell_6t
Xbit_r241_c197 bl[197] br[197] wl[241] vdd gnd cell_6t
Xbit_r242_c197 bl[197] br[197] wl[242] vdd gnd cell_6t
Xbit_r243_c197 bl[197] br[197] wl[243] vdd gnd cell_6t
Xbit_r244_c197 bl[197] br[197] wl[244] vdd gnd cell_6t
Xbit_r245_c197 bl[197] br[197] wl[245] vdd gnd cell_6t
Xbit_r246_c197 bl[197] br[197] wl[246] vdd gnd cell_6t
Xbit_r247_c197 bl[197] br[197] wl[247] vdd gnd cell_6t
Xbit_r248_c197 bl[197] br[197] wl[248] vdd gnd cell_6t
Xbit_r249_c197 bl[197] br[197] wl[249] vdd gnd cell_6t
Xbit_r250_c197 bl[197] br[197] wl[250] vdd gnd cell_6t
Xbit_r251_c197 bl[197] br[197] wl[251] vdd gnd cell_6t
Xbit_r252_c197 bl[197] br[197] wl[252] vdd gnd cell_6t
Xbit_r253_c197 bl[197] br[197] wl[253] vdd gnd cell_6t
Xbit_r254_c197 bl[197] br[197] wl[254] vdd gnd cell_6t
Xbit_r255_c197 bl[197] br[197] wl[255] vdd gnd cell_6t
Xbit_r0_c198 bl[198] br[198] wl[0] vdd gnd cell_6t
Xbit_r1_c198 bl[198] br[198] wl[1] vdd gnd cell_6t
Xbit_r2_c198 bl[198] br[198] wl[2] vdd gnd cell_6t
Xbit_r3_c198 bl[198] br[198] wl[3] vdd gnd cell_6t
Xbit_r4_c198 bl[198] br[198] wl[4] vdd gnd cell_6t
Xbit_r5_c198 bl[198] br[198] wl[5] vdd gnd cell_6t
Xbit_r6_c198 bl[198] br[198] wl[6] vdd gnd cell_6t
Xbit_r7_c198 bl[198] br[198] wl[7] vdd gnd cell_6t
Xbit_r8_c198 bl[198] br[198] wl[8] vdd gnd cell_6t
Xbit_r9_c198 bl[198] br[198] wl[9] vdd gnd cell_6t
Xbit_r10_c198 bl[198] br[198] wl[10] vdd gnd cell_6t
Xbit_r11_c198 bl[198] br[198] wl[11] vdd gnd cell_6t
Xbit_r12_c198 bl[198] br[198] wl[12] vdd gnd cell_6t
Xbit_r13_c198 bl[198] br[198] wl[13] vdd gnd cell_6t
Xbit_r14_c198 bl[198] br[198] wl[14] vdd gnd cell_6t
Xbit_r15_c198 bl[198] br[198] wl[15] vdd gnd cell_6t
Xbit_r16_c198 bl[198] br[198] wl[16] vdd gnd cell_6t
Xbit_r17_c198 bl[198] br[198] wl[17] vdd gnd cell_6t
Xbit_r18_c198 bl[198] br[198] wl[18] vdd gnd cell_6t
Xbit_r19_c198 bl[198] br[198] wl[19] vdd gnd cell_6t
Xbit_r20_c198 bl[198] br[198] wl[20] vdd gnd cell_6t
Xbit_r21_c198 bl[198] br[198] wl[21] vdd gnd cell_6t
Xbit_r22_c198 bl[198] br[198] wl[22] vdd gnd cell_6t
Xbit_r23_c198 bl[198] br[198] wl[23] vdd gnd cell_6t
Xbit_r24_c198 bl[198] br[198] wl[24] vdd gnd cell_6t
Xbit_r25_c198 bl[198] br[198] wl[25] vdd gnd cell_6t
Xbit_r26_c198 bl[198] br[198] wl[26] vdd gnd cell_6t
Xbit_r27_c198 bl[198] br[198] wl[27] vdd gnd cell_6t
Xbit_r28_c198 bl[198] br[198] wl[28] vdd gnd cell_6t
Xbit_r29_c198 bl[198] br[198] wl[29] vdd gnd cell_6t
Xbit_r30_c198 bl[198] br[198] wl[30] vdd gnd cell_6t
Xbit_r31_c198 bl[198] br[198] wl[31] vdd gnd cell_6t
Xbit_r32_c198 bl[198] br[198] wl[32] vdd gnd cell_6t
Xbit_r33_c198 bl[198] br[198] wl[33] vdd gnd cell_6t
Xbit_r34_c198 bl[198] br[198] wl[34] vdd gnd cell_6t
Xbit_r35_c198 bl[198] br[198] wl[35] vdd gnd cell_6t
Xbit_r36_c198 bl[198] br[198] wl[36] vdd gnd cell_6t
Xbit_r37_c198 bl[198] br[198] wl[37] vdd gnd cell_6t
Xbit_r38_c198 bl[198] br[198] wl[38] vdd gnd cell_6t
Xbit_r39_c198 bl[198] br[198] wl[39] vdd gnd cell_6t
Xbit_r40_c198 bl[198] br[198] wl[40] vdd gnd cell_6t
Xbit_r41_c198 bl[198] br[198] wl[41] vdd gnd cell_6t
Xbit_r42_c198 bl[198] br[198] wl[42] vdd gnd cell_6t
Xbit_r43_c198 bl[198] br[198] wl[43] vdd gnd cell_6t
Xbit_r44_c198 bl[198] br[198] wl[44] vdd gnd cell_6t
Xbit_r45_c198 bl[198] br[198] wl[45] vdd gnd cell_6t
Xbit_r46_c198 bl[198] br[198] wl[46] vdd gnd cell_6t
Xbit_r47_c198 bl[198] br[198] wl[47] vdd gnd cell_6t
Xbit_r48_c198 bl[198] br[198] wl[48] vdd gnd cell_6t
Xbit_r49_c198 bl[198] br[198] wl[49] vdd gnd cell_6t
Xbit_r50_c198 bl[198] br[198] wl[50] vdd gnd cell_6t
Xbit_r51_c198 bl[198] br[198] wl[51] vdd gnd cell_6t
Xbit_r52_c198 bl[198] br[198] wl[52] vdd gnd cell_6t
Xbit_r53_c198 bl[198] br[198] wl[53] vdd gnd cell_6t
Xbit_r54_c198 bl[198] br[198] wl[54] vdd gnd cell_6t
Xbit_r55_c198 bl[198] br[198] wl[55] vdd gnd cell_6t
Xbit_r56_c198 bl[198] br[198] wl[56] vdd gnd cell_6t
Xbit_r57_c198 bl[198] br[198] wl[57] vdd gnd cell_6t
Xbit_r58_c198 bl[198] br[198] wl[58] vdd gnd cell_6t
Xbit_r59_c198 bl[198] br[198] wl[59] vdd gnd cell_6t
Xbit_r60_c198 bl[198] br[198] wl[60] vdd gnd cell_6t
Xbit_r61_c198 bl[198] br[198] wl[61] vdd gnd cell_6t
Xbit_r62_c198 bl[198] br[198] wl[62] vdd gnd cell_6t
Xbit_r63_c198 bl[198] br[198] wl[63] vdd gnd cell_6t
Xbit_r64_c198 bl[198] br[198] wl[64] vdd gnd cell_6t
Xbit_r65_c198 bl[198] br[198] wl[65] vdd gnd cell_6t
Xbit_r66_c198 bl[198] br[198] wl[66] vdd gnd cell_6t
Xbit_r67_c198 bl[198] br[198] wl[67] vdd gnd cell_6t
Xbit_r68_c198 bl[198] br[198] wl[68] vdd gnd cell_6t
Xbit_r69_c198 bl[198] br[198] wl[69] vdd gnd cell_6t
Xbit_r70_c198 bl[198] br[198] wl[70] vdd gnd cell_6t
Xbit_r71_c198 bl[198] br[198] wl[71] vdd gnd cell_6t
Xbit_r72_c198 bl[198] br[198] wl[72] vdd gnd cell_6t
Xbit_r73_c198 bl[198] br[198] wl[73] vdd gnd cell_6t
Xbit_r74_c198 bl[198] br[198] wl[74] vdd gnd cell_6t
Xbit_r75_c198 bl[198] br[198] wl[75] vdd gnd cell_6t
Xbit_r76_c198 bl[198] br[198] wl[76] vdd gnd cell_6t
Xbit_r77_c198 bl[198] br[198] wl[77] vdd gnd cell_6t
Xbit_r78_c198 bl[198] br[198] wl[78] vdd gnd cell_6t
Xbit_r79_c198 bl[198] br[198] wl[79] vdd gnd cell_6t
Xbit_r80_c198 bl[198] br[198] wl[80] vdd gnd cell_6t
Xbit_r81_c198 bl[198] br[198] wl[81] vdd gnd cell_6t
Xbit_r82_c198 bl[198] br[198] wl[82] vdd gnd cell_6t
Xbit_r83_c198 bl[198] br[198] wl[83] vdd gnd cell_6t
Xbit_r84_c198 bl[198] br[198] wl[84] vdd gnd cell_6t
Xbit_r85_c198 bl[198] br[198] wl[85] vdd gnd cell_6t
Xbit_r86_c198 bl[198] br[198] wl[86] vdd gnd cell_6t
Xbit_r87_c198 bl[198] br[198] wl[87] vdd gnd cell_6t
Xbit_r88_c198 bl[198] br[198] wl[88] vdd gnd cell_6t
Xbit_r89_c198 bl[198] br[198] wl[89] vdd gnd cell_6t
Xbit_r90_c198 bl[198] br[198] wl[90] vdd gnd cell_6t
Xbit_r91_c198 bl[198] br[198] wl[91] vdd gnd cell_6t
Xbit_r92_c198 bl[198] br[198] wl[92] vdd gnd cell_6t
Xbit_r93_c198 bl[198] br[198] wl[93] vdd gnd cell_6t
Xbit_r94_c198 bl[198] br[198] wl[94] vdd gnd cell_6t
Xbit_r95_c198 bl[198] br[198] wl[95] vdd gnd cell_6t
Xbit_r96_c198 bl[198] br[198] wl[96] vdd gnd cell_6t
Xbit_r97_c198 bl[198] br[198] wl[97] vdd gnd cell_6t
Xbit_r98_c198 bl[198] br[198] wl[98] vdd gnd cell_6t
Xbit_r99_c198 bl[198] br[198] wl[99] vdd gnd cell_6t
Xbit_r100_c198 bl[198] br[198] wl[100] vdd gnd cell_6t
Xbit_r101_c198 bl[198] br[198] wl[101] vdd gnd cell_6t
Xbit_r102_c198 bl[198] br[198] wl[102] vdd gnd cell_6t
Xbit_r103_c198 bl[198] br[198] wl[103] vdd gnd cell_6t
Xbit_r104_c198 bl[198] br[198] wl[104] vdd gnd cell_6t
Xbit_r105_c198 bl[198] br[198] wl[105] vdd gnd cell_6t
Xbit_r106_c198 bl[198] br[198] wl[106] vdd gnd cell_6t
Xbit_r107_c198 bl[198] br[198] wl[107] vdd gnd cell_6t
Xbit_r108_c198 bl[198] br[198] wl[108] vdd gnd cell_6t
Xbit_r109_c198 bl[198] br[198] wl[109] vdd gnd cell_6t
Xbit_r110_c198 bl[198] br[198] wl[110] vdd gnd cell_6t
Xbit_r111_c198 bl[198] br[198] wl[111] vdd gnd cell_6t
Xbit_r112_c198 bl[198] br[198] wl[112] vdd gnd cell_6t
Xbit_r113_c198 bl[198] br[198] wl[113] vdd gnd cell_6t
Xbit_r114_c198 bl[198] br[198] wl[114] vdd gnd cell_6t
Xbit_r115_c198 bl[198] br[198] wl[115] vdd gnd cell_6t
Xbit_r116_c198 bl[198] br[198] wl[116] vdd gnd cell_6t
Xbit_r117_c198 bl[198] br[198] wl[117] vdd gnd cell_6t
Xbit_r118_c198 bl[198] br[198] wl[118] vdd gnd cell_6t
Xbit_r119_c198 bl[198] br[198] wl[119] vdd gnd cell_6t
Xbit_r120_c198 bl[198] br[198] wl[120] vdd gnd cell_6t
Xbit_r121_c198 bl[198] br[198] wl[121] vdd gnd cell_6t
Xbit_r122_c198 bl[198] br[198] wl[122] vdd gnd cell_6t
Xbit_r123_c198 bl[198] br[198] wl[123] vdd gnd cell_6t
Xbit_r124_c198 bl[198] br[198] wl[124] vdd gnd cell_6t
Xbit_r125_c198 bl[198] br[198] wl[125] vdd gnd cell_6t
Xbit_r126_c198 bl[198] br[198] wl[126] vdd gnd cell_6t
Xbit_r127_c198 bl[198] br[198] wl[127] vdd gnd cell_6t
Xbit_r128_c198 bl[198] br[198] wl[128] vdd gnd cell_6t
Xbit_r129_c198 bl[198] br[198] wl[129] vdd gnd cell_6t
Xbit_r130_c198 bl[198] br[198] wl[130] vdd gnd cell_6t
Xbit_r131_c198 bl[198] br[198] wl[131] vdd gnd cell_6t
Xbit_r132_c198 bl[198] br[198] wl[132] vdd gnd cell_6t
Xbit_r133_c198 bl[198] br[198] wl[133] vdd gnd cell_6t
Xbit_r134_c198 bl[198] br[198] wl[134] vdd gnd cell_6t
Xbit_r135_c198 bl[198] br[198] wl[135] vdd gnd cell_6t
Xbit_r136_c198 bl[198] br[198] wl[136] vdd gnd cell_6t
Xbit_r137_c198 bl[198] br[198] wl[137] vdd gnd cell_6t
Xbit_r138_c198 bl[198] br[198] wl[138] vdd gnd cell_6t
Xbit_r139_c198 bl[198] br[198] wl[139] vdd gnd cell_6t
Xbit_r140_c198 bl[198] br[198] wl[140] vdd gnd cell_6t
Xbit_r141_c198 bl[198] br[198] wl[141] vdd gnd cell_6t
Xbit_r142_c198 bl[198] br[198] wl[142] vdd gnd cell_6t
Xbit_r143_c198 bl[198] br[198] wl[143] vdd gnd cell_6t
Xbit_r144_c198 bl[198] br[198] wl[144] vdd gnd cell_6t
Xbit_r145_c198 bl[198] br[198] wl[145] vdd gnd cell_6t
Xbit_r146_c198 bl[198] br[198] wl[146] vdd gnd cell_6t
Xbit_r147_c198 bl[198] br[198] wl[147] vdd gnd cell_6t
Xbit_r148_c198 bl[198] br[198] wl[148] vdd gnd cell_6t
Xbit_r149_c198 bl[198] br[198] wl[149] vdd gnd cell_6t
Xbit_r150_c198 bl[198] br[198] wl[150] vdd gnd cell_6t
Xbit_r151_c198 bl[198] br[198] wl[151] vdd gnd cell_6t
Xbit_r152_c198 bl[198] br[198] wl[152] vdd gnd cell_6t
Xbit_r153_c198 bl[198] br[198] wl[153] vdd gnd cell_6t
Xbit_r154_c198 bl[198] br[198] wl[154] vdd gnd cell_6t
Xbit_r155_c198 bl[198] br[198] wl[155] vdd gnd cell_6t
Xbit_r156_c198 bl[198] br[198] wl[156] vdd gnd cell_6t
Xbit_r157_c198 bl[198] br[198] wl[157] vdd gnd cell_6t
Xbit_r158_c198 bl[198] br[198] wl[158] vdd gnd cell_6t
Xbit_r159_c198 bl[198] br[198] wl[159] vdd gnd cell_6t
Xbit_r160_c198 bl[198] br[198] wl[160] vdd gnd cell_6t
Xbit_r161_c198 bl[198] br[198] wl[161] vdd gnd cell_6t
Xbit_r162_c198 bl[198] br[198] wl[162] vdd gnd cell_6t
Xbit_r163_c198 bl[198] br[198] wl[163] vdd gnd cell_6t
Xbit_r164_c198 bl[198] br[198] wl[164] vdd gnd cell_6t
Xbit_r165_c198 bl[198] br[198] wl[165] vdd gnd cell_6t
Xbit_r166_c198 bl[198] br[198] wl[166] vdd gnd cell_6t
Xbit_r167_c198 bl[198] br[198] wl[167] vdd gnd cell_6t
Xbit_r168_c198 bl[198] br[198] wl[168] vdd gnd cell_6t
Xbit_r169_c198 bl[198] br[198] wl[169] vdd gnd cell_6t
Xbit_r170_c198 bl[198] br[198] wl[170] vdd gnd cell_6t
Xbit_r171_c198 bl[198] br[198] wl[171] vdd gnd cell_6t
Xbit_r172_c198 bl[198] br[198] wl[172] vdd gnd cell_6t
Xbit_r173_c198 bl[198] br[198] wl[173] vdd gnd cell_6t
Xbit_r174_c198 bl[198] br[198] wl[174] vdd gnd cell_6t
Xbit_r175_c198 bl[198] br[198] wl[175] vdd gnd cell_6t
Xbit_r176_c198 bl[198] br[198] wl[176] vdd gnd cell_6t
Xbit_r177_c198 bl[198] br[198] wl[177] vdd gnd cell_6t
Xbit_r178_c198 bl[198] br[198] wl[178] vdd gnd cell_6t
Xbit_r179_c198 bl[198] br[198] wl[179] vdd gnd cell_6t
Xbit_r180_c198 bl[198] br[198] wl[180] vdd gnd cell_6t
Xbit_r181_c198 bl[198] br[198] wl[181] vdd gnd cell_6t
Xbit_r182_c198 bl[198] br[198] wl[182] vdd gnd cell_6t
Xbit_r183_c198 bl[198] br[198] wl[183] vdd gnd cell_6t
Xbit_r184_c198 bl[198] br[198] wl[184] vdd gnd cell_6t
Xbit_r185_c198 bl[198] br[198] wl[185] vdd gnd cell_6t
Xbit_r186_c198 bl[198] br[198] wl[186] vdd gnd cell_6t
Xbit_r187_c198 bl[198] br[198] wl[187] vdd gnd cell_6t
Xbit_r188_c198 bl[198] br[198] wl[188] vdd gnd cell_6t
Xbit_r189_c198 bl[198] br[198] wl[189] vdd gnd cell_6t
Xbit_r190_c198 bl[198] br[198] wl[190] vdd gnd cell_6t
Xbit_r191_c198 bl[198] br[198] wl[191] vdd gnd cell_6t
Xbit_r192_c198 bl[198] br[198] wl[192] vdd gnd cell_6t
Xbit_r193_c198 bl[198] br[198] wl[193] vdd gnd cell_6t
Xbit_r194_c198 bl[198] br[198] wl[194] vdd gnd cell_6t
Xbit_r195_c198 bl[198] br[198] wl[195] vdd gnd cell_6t
Xbit_r196_c198 bl[198] br[198] wl[196] vdd gnd cell_6t
Xbit_r197_c198 bl[198] br[198] wl[197] vdd gnd cell_6t
Xbit_r198_c198 bl[198] br[198] wl[198] vdd gnd cell_6t
Xbit_r199_c198 bl[198] br[198] wl[199] vdd gnd cell_6t
Xbit_r200_c198 bl[198] br[198] wl[200] vdd gnd cell_6t
Xbit_r201_c198 bl[198] br[198] wl[201] vdd gnd cell_6t
Xbit_r202_c198 bl[198] br[198] wl[202] vdd gnd cell_6t
Xbit_r203_c198 bl[198] br[198] wl[203] vdd gnd cell_6t
Xbit_r204_c198 bl[198] br[198] wl[204] vdd gnd cell_6t
Xbit_r205_c198 bl[198] br[198] wl[205] vdd gnd cell_6t
Xbit_r206_c198 bl[198] br[198] wl[206] vdd gnd cell_6t
Xbit_r207_c198 bl[198] br[198] wl[207] vdd gnd cell_6t
Xbit_r208_c198 bl[198] br[198] wl[208] vdd gnd cell_6t
Xbit_r209_c198 bl[198] br[198] wl[209] vdd gnd cell_6t
Xbit_r210_c198 bl[198] br[198] wl[210] vdd gnd cell_6t
Xbit_r211_c198 bl[198] br[198] wl[211] vdd gnd cell_6t
Xbit_r212_c198 bl[198] br[198] wl[212] vdd gnd cell_6t
Xbit_r213_c198 bl[198] br[198] wl[213] vdd gnd cell_6t
Xbit_r214_c198 bl[198] br[198] wl[214] vdd gnd cell_6t
Xbit_r215_c198 bl[198] br[198] wl[215] vdd gnd cell_6t
Xbit_r216_c198 bl[198] br[198] wl[216] vdd gnd cell_6t
Xbit_r217_c198 bl[198] br[198] wl[217] vdd gnd cell_6t
Xbit_r218_c198 bl[198] br[198] wl[218] vdd gnd cell_6t
Xbit_r219_c198 bl[198] br[198] wl[219] vdd gnd cell_6t
Xbit_r220_c198 bl[198] br[198] wl[220] vdd gnd cell_6t
Xbit_r221_c198 bl[198] br[198] wl[221] vdd gnd cell_6t
Xbit_r222_c198 bl[198] br[198] wl[222] vdd gnd cell_6t
Xbit_r223_c198 bl[198] br[198] wl[223] vdd gnd cell_6t
Xbit_r224_c198 bl[198] br[198] wl[224] vdd gnd cell_6t
Xbit_r225_c198 bl[198] br[198] wl[225] vdd gnd cell_6t
Xbit_r226_c198 bl[198] br[198] wl[226] vdd gnd cell_6t
Xbit_r227_c198 bl[198] br[198] wl[227] vdd gnd cell_6t
Xbit_r228_c198 bl[198] br[198] wl[228] vdd gnd cell_6t
Xbit_r229_c198 bl[198] br[198] wl[229] vdd gnd cell_6t
Xbit_r230_c198 bl[198] br[198] wl[230] vdd gnd cell_6t
Xbit_r231_c198 bl[198] br[198] wl[231] vdd gnd cell_6t
Xbit_r232_c198 bl[198] br[198] wl[232] vdd gnd cell_6t
Xbit_r233_c198 bl[198] br[198] wl[233] vdd gnd cell_6t
Xbit_r234_c198 bl[198] br[198] wl[234] vdd gnd cell_6t
Xbit_r235_c198 bl[198] br[198] wl[235] vdd gnd cell_6t
Xbit_r236_c198 bl[198] br[198] wl[236] vdd gnd cell_6t
Xbit_r237_c198 bl[198] br[198] wl[237] vdd gnd cell_6t
Xbit_r238_c198 bl[198] br[198] wl[238] vdd gnd cell_6t
Xbit_r239_c198 bl[198] br[198] wl[239] vdd gnd cell_6t
Xbit_r240_c198 bl[198] br[198] wl[240] vdd gnd cell_6t
Xbit_r241_c198 bl[198] br[198] wl[241] vdd gnd cell_6t
Xbit_r242_c198 bl[198] br[198] wl[242] vdd gnd cell_6t
Xbit_r243_c198 bl[198] br[198] wl[243] vdd gnd cell_6t
Xbit_r244_c198 bl[198] br[198] wl[244] vdd gnd cell_6t
Xbit_r245_c198 bl[198] br[198] wl[245] vdd gnd cell_6t
Xbit_r246_c198 bl[198] br[198] wl[246] vdd gnd cell_6t
Xbit_r247_c198 bl[198] br[198] wl[247] vdd gnd cell_6t
Xbit_r248_c198 bl[198] br[198] wl[248] vdd gnd cell_6t
Xbit_r249_c198 bl[198] br[198] wl[249] vdd gnd cell_6t
Xbit_r250_c198 bl[198] br[198] wl[250] vdd gnd cell_6t
Xbit_r251_c198 bl[198] br[198] wl[251] vdd gnd cell_6t
Xbit_r252_c198 bl[198] br[198] wl[252] vdd gnd cell_6t
Xbit_r253_c198 bl[198] br[198] wl[253] vdd gnd cell_6t
Xbit_r254_c198 bl[198] br[198] wl[254] vdd gnd cell_6t
Xbit_r255_c198 bl[198] br[198] wl[255] vdd gnd cell_6t
Xbit_r0_c199 bl[199] br[199] wl[0] vdd gnd cell_6t
Xbit_r1_c199 bl[199] br[199] wl[1] vdd gnd cell_6t
Xbit_r2_c199 bl[199] br[199] wl[2] vdd gnd cell_6t
Xbit_r3_c199 bl[199] br[199] wl[3] vdd gnd cell_6t
Xbit_r4_c199 bl[199] br[199] wl[4] vdd gnd cell_6t
Xbit_r5_c199 bl[199] br[199] wl[5] vdd gnd cell_6t
Xbit_r6_c199 bl[199] br[199] wl[6] vdd gnd cell_6t
Xbit_r7_c199 bl[199] br[199] wl[7] vdd gnd cell_6t
Xbit_r8_c199 bl[199] br[199] wl[8] vdd gnd cell_6t
Xbit_r9_c199 bl[199] br[199] wl[9] vdd gnd cell_6t
Xbit_r10_c199 bl[199] br[199] wl[10] vdd gnd cell_6t
Xbit_r11_c199 bl[199] br[199] wl[11] vdd gnd cell_6t
Xbit_r12_c199 bl[199] br[199] wl[12] vdd gnd cell_6t
Xbit_r13_c199 bl[199] br[199] wl[13] vdd gnd cell_6t
Xbit_r14_c199 bl[199] br[199] wl[14] vdd gnd cell_6t
Xbit_r15_c199 bl[199] br[199] wl[15] vdd gnd cell_6t
Xbit_r16_c199 bl[199] br[199] wl[16] vdd gnd cell_6t
Xbit_r17_c199 bl[199] br[199] wl[17] vdd gnd cell_6t
Xbit_r18_c199 bl[199] br[199] wl[18] vdd gnd cell_6t
Xbit_r19_c199 bl[199] br[199] wl[19] vdd gnd cell_6t
Xbit_r20_c199 bl[199] br[199] wl[20] vdd gnd cell_6t
Xbit_r21_c199 bl[199] br[199] wl[21] vdd gnd cell_6t
Xbit_r22_c199 bl[199] br[199] wl[22] vdd gnd cell_6t
Xbit_r23_c199 bl[199] br[199] wl[23] vdd gnd cell_6t
Xbit_r24_c199 bl[199] br[199] wl[24] vdd gnd cell_6t
Xbit_r25_c199 bl[199] br[199] wl[25] vdd gnd cell_6t
Xbit_r26_c199 bl[199] br[199] wl[26] vdd gnd cell_6t
Xbit_r27_c199 bl[199] br[199] wl[27] vdd gnd cell_6t
Xbit_r28_c199 bl[199] br[199] wl[28] vdd gnd cell_6t
Xbit_r29_c199 bl[199] br[199] wl[29] vdd gnd cell_6t
Xbit_r30_c199 bl[199] br[199] wl[30] vdd gnd cell_6t
Xbit_r31_c199 bl[199] br[199] wl[31] vdd gnd cell_6t
Xbit_r32_c199 bl[199] br[199] wl[32] vdd gnd cell_6t
Xbit_r33_c199 bl[199] br[199] wl[33] vdd gnd cell_6t
Xbit_r34_c199 bl[199] br[199] wl[34] vdd gnd cell_6t
Xbit_r35_c199 bl[199] br[199] wl[35] vdd gnd cell_6t
Xbit_r36_c199 bl[199] br[199] wl[36] vdd gnd cell_6t
Xbit_r37_c199 bl[199] br[199] wl[37] vdd gnd cell_6t
Xbit_r38_c199 bl[199] br[199] wl[38] vdd gnd cell_6t
Xbit_r39_c199 bl[199] br[199] wl[39] vdd gnd cell_6t
Xbit_r40_c199 bl[199] br[199] wl[40] vdd gnd cell_6t
Xbit_r41_c199 bl[199] br[199] wl[41] vdd gnd cell_6t
Xbit_r42_c199 bl[199] br[199] wl[42] vdd gnd cell_6t
Xbit_r43_c199 bl[199] br[199] wl[43] vdd gnd cell_6t
Xbit_r44_c199 bl[199] br[199] wl[44] vdd gnd cell_6t
Xbit_r45_c199 bl[199] br[199] wl[45] vdd gnd cell_6t
Xbit_r46_c199 bl[199] br[199] wl[46] vdd gnd cell_6t
Xbit_r47_c199 bl[199] br[199] wl[47] vdd gnd cell_6t
Xbit_r48_c199 bl[199] br[199] wl[48] vdd gnd cell_6t
Xbit_r49_c199 bl[199] br[199] wl[49] vdd gnd cell_6t
Xbit_r50_c199 bl[199] br[199] wl[50] vdd gnd cell_6t
Xbit_r51_c199 bl[199] br[199] wl[51] vdd gnd cell_6t
Xbit_r52_c199 bl[199] br[199] wl[52] vdd gnd cell_6t
Xbit_r53_c199 bl[199] br[199] wl[53] vdd gnd cell_6t
Xbit_r54_c199 bl[199] br[199] wl[54] vdd gnd cell_6t
Xbit_r55_c199 bl[199] br[199] wl[55] vdd gnd cell_6t
Xbit_r56_c199 bl[199] br[199] wl[56] vdd gnd cell_6t
Xbit_r57_c199 bl[199] br[199] wl[57] vdd gnd cell_6t
Xbit_r58_c199 bl[199] br[199] wl[58] vdd gnd cell_6t
Xbit_r59_c199 bl[199] br[199] wl[59] vdd gnd cell_6t
Xbit_r60_c199 bl[199] br[199] wl[60] vdd gnd cell_6t
Xbit_r61_c199 bl[199] br[199] wl[61] vdd gnd cell_6t
Xbit_r62_c199 bl[199] br[199] wl[62] vdd gnd cell_6t
Xbit_r63_c199 bl[199] br[199] wl[63] vdd gnd cell_6t
Xbit_r64_c199 bl[199] br[199] wl[64] vdd gnd cell_6t
Xbit_r65_c199 bl[199] br[199] wl[65] vdd gnd cell_6t
Xbit_r66_c199 bl[199] br[199] wl[66] vdd gnd cell_6t
Xbit_r67_c199 bl[199] br[199] wl[67] vdd gnd cell_6t
Xbit_r68_c199 bl[199] br[199] wl[68] vdd gnd cell_6t
Xbit_r69_c199 bl[199] br[199] wl[69] vdd gnd cell_6t
Xbit_r70_c199 bl[199] br[199] wl[70] vdd gnd cell_6t
Xbit_r71_c199 bl[199] br[199] wl[71] vdd gnd cell_6t
Xbit_r72_c199 bl[199] br[199] wl[72] vdd gnd cell_6t
Xbit_r73_c199 bl[199] br[199] wl[73] vdd gnd cell_6t
Xbit_r74_c199 bl[199] br[199] wl[74] vdd gnd cell_6t
Xbit_r75_c199 bl[199] br[199] wl[75] vdd gnd cell_6t
Xbit_r76_c199 bl[199] br[199] wl[76] vdd gnd cell_6t
Xbit_r77_c199 bl[199] br[199] wl[77] vdd gnd cell_6t
Xbit_r78_c199 bl[199] br[199] wl[78] vdd gnd cell_6t
Xbit_r79_c199 bl[199] br[199] wl[79] vdd gnd cell_6t
Xbit_r80_c199 bl[199] br[199] wl[80] vdd gnd cell_6t
Xbit_r81_c199 bl[199] br[199] wl[81] vdd gnd cell_6t
Xbit_r82_c199 bl[199] br[199] wl[82] vdd gnd cell_6t
Xbit_r83_c199 bl[199] br[199] wl[83] vdd gnd cell_6t
Xbit_r84_c199 bl[199] br[199] wl[84] vdd gnd cell_6t
Xbit_r85_c199 bl[199] br[199] wl[85] vdd gnd cell_6t
Xbit_r86_c199 bl[199] br[199] wl[86] vdd gnd cell_6t
Xbit_r87_c199 bl[199] br[199] wl[87] vdd gnd cell_6t
Xbit_r88_c199 bl[199] br[199] wl[88] vdd gnd cell_6t
Xbit_r89_c199 bl[199] br[199] wl[89] vdd gnd cell_6t
Xbit_r90_c199 bl[199] br[199] wl[90] vdd gnd cell_6t
Xbit_r91_c199 bl[199] br[199] wl[91] vdd gnd cell_6t
Xbit_r92_c199 bl[199] br[199] wl[92] vdd gnd cell_6t
Xbit_r93_c199 bl[199] br[199] wl[93] vdd gnd cell_6t
Xbit_r94_c199 bl[199] br[199] wl[94] vdd gnd cell_6t
Xbit_r95_c199 bl[199] br[199] wl[95] vdd gnd cell_6t
Xbit_r96_c199 bl[199] br[199] wl[96] vdd gnd cell_6t
Xbit_r97_c199 bl[199] br[199] wl[97] vdd gnd cell_6t
Xbit_r98_c199 bl[199] br[199] wl[98] vdd gnd cell_6t
Xbit_r99_c199 bl[199] br[199] wl[99] vdd gnd cell_6t
Xbit_r100_c199 bl[199] br[199] wl[100] vdd gnd cell_6t
Xbit_r101_c199 bl[199] br[199] wl[101] vdd gnd cell_6t
Xbit_r102_c199 bl[199] br[199] wl[102] vdd gnd cell_6t
Xbit_r103_c199 bl[199] br[199] wl[103] vdd gnd cell_6t
Xbit_r104_c199 bl[199] br[199] wl[104] vdd gnd cell_6t
Xbit_r105_c199 bl[199] br[199] wl[105] vdd gnd cell_6t
Xbit_r106_c199 bl[199] br[199] wl[106] vdd gnd cell_6t
Xbit_r107_c199 bl[199] br[199] wl[107] vdd gnd cell_6t
Xbit_r108_c199 bl[199] br[199] wl[108] vdd gnd cell_6t
Xbit_r109_c199 bl[199] br[199] wl[109] vdd gnd cell_6t
Xbit_r110_c199 bl[199] br[199] wl[110] vdd gnd cell_6t
Xbit_r111_c199 bl[199] br[199] wl[111] vdd gnd cell_6t
Xbit_r112_c199 bl[199] br[199] wl[112] vdd gnd cell_6t
Xbit_r113_c199 bl[199] br[199] wl[113] vdd gnd cell_6t
Xbit_r114_c199 bl[199] br[199] wl[114] vdd gnd cell_6t
Xbit_r115_c199 bl[199] br[199] wl[115] vdd gnd cell_6t
Xbit_r116_c199 bl[199] br[199] wl[116] vdd gnd cell_6t
Xbit_r117_c199 bl[199] br[199] wl[117] vdd gnd cell_6t
Xbit_r118_c199 bl[199] br[199] wl[118] vdd gnd cell_6t
Xbit_r119_c199 bl[199] br[199] wl[119] vdd gnd cell_6t
Xbit_r120_c199 bl[199] br[199] wl[120] vdd gnd cell_6t
Xbit_r121_c199 bl[199] br[199] wl[121] vdd gnd cell_6t
Xbit_r122_c199 bl[199] br[199] wl[122] vdd gnd cell_6t
Xbit_r123_c199 bl[199] br[199] wl[123] vdd gnd cell_6t
Xbit_r124_c199 bl[199] br[199] wl[124] vdd gnd cell_6t
Xbit_r125_c199 bl[199] br[199] wl[125] vdd gnd cell_6t
Xbit_r126_c199 bl[199] br[199] wl[126] vdd gnd cell_6t
Xbit_r127_c199 bl[199] br[199] wl[127] vdd gnd cell_6t
Xbit_r128_c199 bl[199] br[199] wl[128] vdd gnd cell_6t
Xbit_r129_c199 bl[199] br[199] wl[129] vdd gnd cell_6t
Xbit_r130_c199 bl[199] br[199] wl[130] vdd gnd cell_6t
Xbit_r131_c199 bl[199] br[199] wl[131] vdd gnd cell_6t
Xbit_r132_c199 bl[199] br[199] wl[132] vdd gnd cell_6t
Xbit_r133_c199 bl[199] br[199] wl[133] vdd gnd cell_6t
Xbit_r134_c199 bl[199] br[199] wl[134] vdd gnd cell_6t
Xbit_r135_c199 bl[199] br[199] wl[135] vdd gnd cell_6t
Xbit_r136_c199 bl[199] br[199] wl[136] vdd gnd cell_6t
Xbit_r137_c199 bl[199] br[199] wl[137] vdd gnd cell_6t
Xbit_r138_c199 bl[199] br[199] wl[138] vdd gnd cell_6t
Xbit_r139_c199 bl[199] br[199] wl[139] vdd gnd cell_6t
Xbit_r140_c199 bl[199] br[199] wl[140] vdd gnd cell_6t
Xbit_r141_c199 bl[199] br[199] wl[141] vdd gnd cell_6t
Xbit_r142_c199 bl[199] br[199] wl[142] vdd gnd cell_6t
Xbit_r143_c199 bl[199] br[199] wl[143] vdd gnd cell_6t
Xbit_r144_c199 bl[199] br[199] wl[144] vdd gnd cell_6t
Xbit_r145_c199 bl[199] br[199] wl[145] vdd gnd cell_6t
Xbit_r146_c199 bl[199] br[199] wl[146] vdd gnd cell_6t
Xbit_r147_c199 bl[199] br[199] wl[147] vdd gnd cell_6t
Xbit_r148_c199 bl[199] br[199] wl[148] vdd gnd cell_6t
Xbit_r149_c199 bl[199] br[199] wl[149] vdd gnd cell_6t
Xbit_r150_c199 bl[199] br[199] wl[150] vdd gnd cell_6t
Xbit_r151_c199 bl[199] br[199] wl[151] vdd gnd cell_6t
Xbit_r152_c199 bl[199] br[199] wl[152] vdd gnd cell_6t
Xbit_r153_c199 bl[199] br[199] wl[153] vdd gnd cell_6t
Xbit_r154_c199 bl[199] br[199] wl[154] vdd gnd cell_6t
Xbit_r155_c199 bl[199] br[199] wl[155] vdd gnd cell_6t
Xbit_r156_c199 bl[199] br[199] wl[156] vdd gnd cell_6t
Xbit_r157_c199 bl[199] br[199] wl[157] vdd gnd cell_6t
Xbit_r158_c199 bl[199] br[199] wl[158] vdd gnd cell_6t
Xbit_r159_c199 bl[199] br[199] wl[159] vdd gnd cell_6t
Xbit_r160_c199 bl[199] br[199] wl[160] vdd gnd cell_6t
Xbit_r161_c199 bl[199] br[199] wl[161] vdd gnd cell_6t
Xbit_r162_c199 bl[199] br[199] wl[162] vdd gnd cell_6t
Xbit_r163_c199 bl[199] br[199] wl[163] vdd gnd cell_6t
Xbit_r164_c199 bl[199] br[199] wl[164] vdd gnd cell_6t
Xbit_r165_c199 bl[199] br[199] wl[165] vdd gnd cell_6t
Xbit_r166_c199 bl[199] br[199] wl[166] vdd gnd cell_6t
Xbit_r167_c199 bl[199] br[199] wl[167] vdd gnd cell_6t
Xbit_r168_c199 bl[199] br[199] wl[168] vdd gnd cell_6t
Xbit_r169_c199 bl[199] br[199] wl[169] vdd gnd cell_6t
Xbit_r170_c199 bl[199] br[199] wl[170] vdd gnd cell_6t
Xbit_r171_c199 bl[199] br[199] wl[171] vdd gnd cell_6t
Xbit_r172_c199 bl[199] br[199] wl[172] vdd gnd cell_6t
Xbit_r173_c199 bl[199] br[199] wl[173] vdd gnd cell_6t
Xbit_r174_c199 bl[199] br[199] wl[174] vdd gnd cell_6t
Xbit_r175_c199 bl[199] br[199] wl[175] vdd gnd cell_6t
Xbit_r176_c199 bl[199] br[199] wl[176] vdd gnd cell_6t
Xbit_r177_c199 bl[199] br[199] wl[177] vdd gnd cell_6t
Xbit_r178_c199 bl[199] br[199] wl[178] vdd gnd cell_6t
Xbit_r179_c199 bl[199] br[199] wl[179] vdd gnd cell_6t
Xbit_r180_c199 bl[199] br[199] wl[180] vdd gnd cell_6t
Xbit_r181_c199 bl[199] br[199] wl[181] vdd gnd cell_6t
Xbit_r182_c199 bl[199] br[199] wl[182] vdd gnd cell_6t
Xbit_r183_c199 bl[199] br[199] wl[183] vdd gnd cell_6t
Xbit_r184_c199 bl[199] br[199] wl[184] vdd gnd cell_6t
Xbit_r185_c199 bl[199] br[199] wl[185] vdd gnd cell_6t
Xbit_r186_c199 bl[199] br[199] wl[186] vdd gnd cell_6t
Xbit_r187_c199 bl[199] br[199] wl[187] vdd gnd cell_6t
Xbit_r188_c199 bl[199] br[199] wl[188] vdd gnd cell_6t
Xbit_r189_c199 bl[199] br[199] wl[189] vdd gnd cell_6t
Xbit_r190_c199 bl[199] br[199] wl[190] vdd gnd cell_6t
Xbit_r191_c199 bl[199] br[199] wl[191] vdd gnd cell_6t
Xbit_r192_c199 bl[199] br[199] wl[192] vdd gnd cell_6t
Xbit_r193_c199 bl[199] br[199] wl[193] vdd gnd cell_6t
Xbit_r194_c199 bl[199] br[199] wl[194] vdd gnd cell_6t
Xbit_r195_c199 bl[199] br[199] wl[195] vdd gnd cell_6t
Xbit_r196_c199 bl[199] br[199] wl[196] vdd gnd cell_6t
Xbit_r197_c199 bl[199] br[199] wl[197] vdd gnd cell_6t
Xbit_r198_c199 bl[199] br[199] wl[198] vdd gnd cell_6t
Xbit_r199_c199 bl[199] br[199] wl[199] vdd gnd cell_6t
Xbit_r200_c199 bl[199] br[199] wl[200] vdd gnd cell_6t
Xbit_r201_c199 bl[199] br[199] wl[201] vdd gnd cell_6t
Xbit_r202_c199 bl[199] br[199] wl[202] vdd gnd cell_6t
Xbit_r203_c199 bl[199] br[199] wl[203] vdd gnd cell_6t
Xbit_r204_c199 bl[199] br[199] wl[204] vdd gnd cell_6t
Xbit_r205_c199 bl[199] br[199] wl[205] vdd gnd cell_6t
Xbit_r206_c199 bl[199] br[199] wl[206] vdd gnd cell_6t
Xbit_r207_c199 bl[199] br[199] wl[207] vdd gnd cell_6t
Xbit_r208_c199 bl[199] br[199] wl[208] vdd gnd cell_6t
Xbit_r209_c199 bl[199] br[199] wl[209] vdd gnd cell_6t
Xbit_r210_c199 bl[199] br[199] wl[210] vdd gnd cell_6t
Xbit_r211_c199 bl[199] br[199] wl[211] vdd gnd cell_6t
Xbit_r212_c199 bl[199] br[199] wl[212] vdd gnd cell_6t
Xbit_r213_c199 bl[199] br[199] wl[213] vdd gnd cell_6t
Xbit_r214_c199 bl[199] br[199] wl[214] vdd gnd cell_6t
Xbit_r215_c199 bl[199] br[199] wl[215] vdd gnd cell_6t
Xbit_r216_c199 bl[199] br[199] wl[216] vdd gnd cell_6t
Xbit_r217_c199 bl[199] br[199] wl[217] vdd gnd cell_6t
Xbit_r218_c199 bl[199] br[199] wl[218] vdd gnd cell_6t
Xbit_r219_c199 bl[199] br[199] wl[219] vdd gnd cell_6t
Xbit_r220_c199 bl[199] br[199] wl[220] vdd gnd cell_6t
Xbit_r221_c199 bl[199] br[199] wl[221] vdd gnd cell_6t
Xbit_r222_c199 bl[199] br[199] wl[222] vdd gnd cell_6t
Xbit_r223_c199 bl[199] br[199] wl[223] vdd gnd cell_6t
Xbit_r224_c199 bl[199] br[199] wl[224] vdd gnd cell_6t
Xbit_r225_c199 bl[199] br[199] wl[225] vdd gnd cell_6t
Xbit_r226_c199 bl[199] br[199] wl[226] vdd gnd cell_6t
Xbit_r227_c199 bl[199] br[199] wl[227] vdd gnd cell_6t
Xbit_r228_c199 bl[199] br[199] wl[228] vdd gnd cell_6t
Xbit_r229_c199 bl[199] br[199] wl[229] vdd gnd cell_6t
Xbit_r230_c199 bl[199] br[199] wl[230] vdd gnd cell_6t
Xbit_r231_c199 bl[199] br[199] wl[231] vdd gnd cell_6t
Xbit_r232_c199 bl[199] br[199] wl[232] vdd gnd cell_6t
Xbit_r233_c199 bl[199] br[199] wl[233] vdd gnd cell_6t
Xbit_r234_c199 bl[199] br[199] wl[234] vdd gnd cell_6t
Xbit_r235_c199 bl[199] br[199] wl[235] vdd gnd cell_6t
Xbit_r236_c199 bl[199] br[199] wl[236] vdd gnd cell_6t
Xbit_r237_c199 bl[199] br[199] wl[237] vdd gnd cell_6t
Xbit_r238_c199 bl[199] br[199] wl[238] vdd gnd cell_6t
Xbit_r239_c199 bl[199] br[199] wl[239] vdd gnd cell_6t
Xbit_r240_c199 bl[199] br[199] wl[240] vdd gnd cell_6t
Xbit_r241_c199 bl[199] br[199] wl[241] vdd gnd cell_6t
Xbit_r242_c199 bl[199] br[199] wl[242] vdd gnd cell_6t
Xbit_r243_c199 bl[199] br[199] wl[243] vdd gnd cell_6t
Xbit_r244_c199 bl[199] br[199] wl[244] vdd gnd cell_6t
Xbit_r245_c199 bl[199] br[199] wl[245] vdd gnd cell_6t
Xbit_r246_c199 bl[199] br[199] wl[246] vdd gnd cell_6t
Xbit_r247_c199 bl[199] br[199] wl[247] vdd gnd cell_6t
Xbit_r248_c199 bl[199] br[199] wl[248] vdd gnd cell_6t
Xbit_r249_c199 bl[199] br[199] wl[249] vdd gnd cell_6t
Xbit_r250_c199 bl[199] br[199] wl[250] vdd gnd cell_6t
Xbit_r251_c199 bl[199] br[199] wl[251] vdd gnd cell_6t
Xbit_r252_c199 bl[199] br[199] wl[252] vdd gnd cell_6t
Xbit_r253_c199 bl[199] br[199] wl[253] vdd gnd cell_6t
Xbit_r254_c199 bl[199] br[199] wl[254] vdd gnd cell_6t
Xbit_r255_c199 bl[199] br[199] wl[255] vdd gnd cell_6t
Xbit_r0_c200 bl[200] br[200] wl[0] vdd gnd cell_6t
Xbit_r1_c200 bl[200] br[200] wl[1] vdd gnd cell_6t
Xbit_r2_c200 bl[200] br[200] wl[2] vdd gnd cell_6t
Xbit_r3_c200 bl[200] br[200] wl[3] vdd gnd cell_6t
Xbit_r4_c200 bl[200] br[200] wl[4] vdd gnd cell_6t
Xbit_r5_c200 bl[200] br[200] wl[5] vdd gnd cell_6t
Xbit_r6_c200 bl[200] br[200] wl[6] vdd gnd cell_6t
Xbit_r7_c200 bl[200] br[200] wl[7] vdd gnd cell_6t
Xbit_r8_c200 bl[200] br[200] wl[8] vdd gnd cell_6t
Xbit_r9_c200 bl[200] br[200] wl[9] vdd gnd cell_6t
Xbit_r10_c200 bl[200] br[200] wl[10] vdd gnd cell_6t
Xbit_r11_c200 bl[200] br[200] wl[11] vdd gnd cell_6t
Xbit_r12_c200 bl[200] br[200] wl[12] vdd gnd cell_6t
Xbit_r13_c200 bl[200] br[200] wl[13] vdd gnd cell_6t
Xbit_r14_c200 bl[200] br[200] wl[14] vdd gnd cell_6t
Xbit_r15_c200 bl[200] br[200] wl[15] vdd gnd cell_6t
Xbit_r16_c200 bl[200] br[200] wl[16] vdd gnd cell_6t
Xbit_r17_c200 bl[200] br[200] wl[17] vdd gnd cell_6t
Xbit_r18_c200 bl[200] br[200] wl[18] vdd gnd cell_6t
Xbit_r19_c200 bl[200] br[200] wl[19] vdd gnd cell_6t
Xbit_r20_c200 bl[200] br[200] wl[20] vdd gnd cell_6t
Xbit_r21_c200 bl[200] br[200] wl[21] vdd gnd cell_6t
Xbit_r22_c200 bl[200] br[200] wl[22] vdd gnd cell_6t
Xbit_r23_c200 bl[200] br[200] wl[23] vdd gnd cell_6t
Xbit_r24_c200 bl[200] br[200] wl[24] vdd gnd cell_6t
Xbit_r25_c200 bl[200] br[200] wl[25] vdd gnd cell_6t
Xbit_r26_c200 bl[200] br[200] wl[26] vdd gnd cell_6t
Xbit_r27_c200 bl[200] br[200] wl[27] vdd gnd cell_6t
Xbit_r28_c200 bl[200] br[200] wl[28] vdd gnd cell_6t
Xbit_r29_c200 bl[200] br[200] wl[29] vdd gnd cell_6t
Xbit_r30_c200 bl[200] br[200] wl[30] vdd gnd cell_6t
Xbit_r31_c200 bl[200] br[200] wl[31] vdd gnd cell_6t
Xbit_r32_c200 bl[200] br[200] wl[32] vdd gnd cell_6t
Xbit_r33_c200 bl[200] br[200] wl[33] vdd gnd cell_6t
Xbit_r34_c200 bl[200] br[200] wl[34] vdd gnd cell_6t
Xbit_r35_c200 bl[200] br[200] wl[35] vdd gnd cell_6t
Xbit_r36_c200 bl[200] br[200] wl[36] vdd gnd cell_6t
Xbit_r37_c200 bl[200] br[200] wl[37] vdd gnd cell_6t
Xbit_r38_c200 bl[200] br[200] wl[38] vdd gnd cell_6t
Xbit_r39_c200 bl[200] br[200] wl[39] vdd gnd cell_6t
Xbit_r40_c200 bl[200] br[200] wl[40] vdd gnd cell_6t
Xbit_r41_c200 bl[200] br[200] wl[41] vdd gnd cell_6t
Xbit_r42_c200 bl[200] br[200] wl[42] vdd gnd cell_6t
Xbit_r43_c200 bl[200] br[200] wl[43] vdd gnd cell_6t
Xbit_r44_c200 bl[200] br[200] wl[44] vdd gnd cell_6t
Xbit_r45_c200 bl[200] br[200] wl[45] vdd gnd cell_6t
Xbit_r46_c200 bl[200] br[200] wl[46] vdd gnd cell_6t
Xbit_r47_c200 bl[200] br[200] wl[47] vdd gnd cell_6t
Xbit_r48_c200 bl[200] br[200] wl[48] vdd gnd cell_6t
Xbit_r49_c200 bl[200] br[200] wl[49] vdd gnd cell_6t
Xbit_r50_c200 bl[200] br[200] wl[50] vdd gnd cell_6t
Xbit_r51_c200 bl[200] br[200] wl[51] vdd gnd cell_6t
Xbit_r52_c200 bl[200] br[200] wl[52] vdd gnd cell_6t
Xbit_r53_c200 bl[200] br[200] wl[53] vdd gnd cell_6t
Xbit_r54_c200 bl[200] br[200] wl[54] vdd gnd cell_6t
Xbit_r55_c200 bl[200] br[200] wl[55] vdd gnd cell_6t
Xbit_r56_c200 bl[200] br[200] wl[56] vdd gnd cell_6t
Xbit_r57_c200 bl[200] br[200] wl[57] vdd gnd cell_6t
Xbit_r58_c200 bl[200] br[200] wl[58] vdd gnd cell_6t
Xbit_r59_c200 bl[200] br[200] wl[59] vdd gnd cell_6t
Xbit_r60_c200 bl[200] br[200] wl[60] vdd gnd cell_6t
Xbit_r61_c200 bl[200] br[200] wl[61] vdd gnd cell_6t
Xbit_r62_c200 bl[200] br[200] wl[62] vdd gnd cell_6t
Xbit_r63_c200 bl[200] br[200] wl[63] vdd gnd cell_6t
Xbit_r64_c200 bl[200] br[200] wl[64] vdd gnd cell_6t
Xbit_r65_c200 bl[200] br[200] wl[65] vdd gnd cell_6t
Xbit_r66_c200 bl[200] br[200] wl[66] vdd gnd cell_6t
Xbit_r67_c200 bl[200] br[200] wl[67] vdd gnd cell_6t
Xbit_r68_c200 bl[200] br[200] wl[68] vdd gnd cell_6t
Xbit_r69_c200 bl[200] br[200] wl[69] vdd gnd cell_6t
Xbit_r70_c200 bl[200] br[200] wl[70] vdd gnd cell_6t
Xbit_r71_c200 bl[200] br[200] wl[71] vdd gnd cell_6t
Xbit_r72_c200 bl[200] br[200] wl[72] vdd gnd cell_6t
Xbit_r73_c200 bl[200] br[200] wl[73] vdd gnd cell_6t
Xbit_r74_c200 bl[200] br[200] wl[74] vdd gnd cell_6t
Xbit_r75_c200 bl[200] br[200] wl[75] vdd gnd cell_6t
Xbit_r76_c200 bl[200] br[200] wl[76] vdd gnd cell_6t
Xbit_r77_c200 bl[200] br[200] wl[77] vdd gnd cell_6t
Xbit_r78_c200 bl[200] br[200] wl[78] vdd gnd cell_6t
Xbit_r79_c200 bl[200] br[200] wl[79] vdd gnd cell_6t
Xbit_r80_c200 bl[200] br[200] wl[80] vdd gnd cell_6t
Xbit_r81_c200 bl[200] br[200] wl[81] vdd gnd cell_6t
Xbit_r82_c200 bl[200] br[200] wl[82] vdd gnd cell_6t
Xbit_r83_c200 bl[200] br[200] wl[83] vdd gnd cell_6t
Xbit_r84_c200 bl[200] br[200] wl[84] vdd gnd cell_6t
Xbit_r85_c200 bl[200] br[200] wl[85] vdd gnd cell_6t
Xbit_r86_c200 bl[200] br[200] wl[86] vdd gnd cell_6t
Xbit_r87_c200 bl[200] br[200] wl[87] vdd gnd cell_6t
Xbit_r88_c200 bl[200] br[200] wl[88] vdd gnd cell_6t
Xbit_r89_c200 bl[200] br[200] wl[89] vdd gnd cell_6t
Xbit_r90_c200 bl[200] br[200] wl[90] vdd gnd cell_6t
Xbit_r91_c200 bl[200] br[200] wl[91] vdd gnd cell_6t
Xbit_r92_c200 bl[200] br[200] wl[92] vdd gnd cell_6t
Xbit_r93_c200 bl[200] br[200] wl[93] vdd gnd cell_6t
Xbit_r94_c200 bl[200] br[200] wl[94] vdd gnd cell_6t
Xbit_r95_c200 bl[200] br[200] wl[95] vdd gnd cell_6t
Xbit_r96_c200 bl[200] br[200] wl[96] vdd gnd cell_6t
Xbit_r97_c200 bl[200] br[200] wl[97] vdd gnd cell_6t
Xbit_r98_c200 bl[200] br[200] wl[98] vdd gnd cell_6t
Xbit_r99_c200 bl[200] br[200] wl[99] vdd gnd cell_6t
Xbit_r100_c200 bl[200] br[200] wl[100] vdd gnd cell_6t
Xbit_r101_c200 bl[200] br[200] wl[101] vdd gnd cell_6t
Xbit_r102_c200 bl[200] br[200] wl[102] vdd gnd cell_6t
Xbit_r103_c200 bl[200] br[200] wl[103] vdd gnd cell_6t
Xbit_r104_c200 bl[200] br[200] wl[104] vdd gnd cell_6t
Xbit_r105_c200 bl[200] br[200] wl[105] vdd gnd cell_6t
Xbit_r106_c200 bl[200] br[200] wl[106] vdd gnd cell_6t
Xbit_r107_c200 bl[200] br[200] wl[107] vdd gnd cell_6t
Xbit_r108_c200 bl[200] br[200] wl[108] vdd gnd cell_6t
Xbit_r109_c200 bl[200] br[200] wl[109] vdd gnd cell_6t
Xbit_r110_c200 bl[200] br[200] wl[110] vdd gnd cell_6t
Xbit_r111_c200 bl[200] br[200] wl[111] vdd gnd cell_6t
Xbit_r112_c200 bl[200] br[200] wl[112] vdd gnd cell_6t
Xbit_r113_c200 bl[200] br[200] wl[113] vdd gnd cell_6t
Xbit_r114_c200 bl[200] br[200] wl[114] vdd gnd cell_6t
Xbit_r115_c200 bl[200] br[200] wl[115] vdd gnd cell_6t
Xbit_r116_c200 bl[200] br[200] wl[116] vdd gnd cell_6t
Xbit_r117_c200 bl[200] br[200] wl[117] vdd gnd cell_6t
Xbit_r118_c200 bl[200] br[200] wl[118] vdd gnd cell_6t
Xbit_r119_c200 bl[200] br[200] wl[119] vdd gnd cell_6t
Xbit_r120_c200 bl[200] br[200] wl[120] vdd gnd cell_6t
Xbit_r121_c200 bl[200] br[200] wl[121] vdd gnd cell_6t
Xbit_r122_c200 bl[200] br[200] wl[122] vdd gnd cell_6t
Xbit_r123_c200 bl[200] br[200] wl[123] vdd gnd cell_6t
Xbit_r124_c200 bl[200] br[200] wl[124] vdd gnd cell_6t
Xbit_r125_c200 bl[200] br[200] wl[125] vdd gnd cell_6t
Xbit_r126_c200 bl[200] br[200] wl[126] vdd gnd cell_6t
Xbit_r127_c200 bl[200] br[200] wl[127] vdd gnd cell_6t
Xbit_r128_c200 bl[200] br[200] wl[128] vdd gnd cell_6t
Xbit_r129_c200 bl[200] br[200] wl[129] vdd gnd cell_6t
Xbit_r130_c200 bl[200] br[200] wl[130] vdd gnd cell_6t
Xbit_r131_c200 bl[200] br[200] wl[131] vdd gnd cell_6t
Xbit_r132_c200 bl[200] br[200] wl[132] vdd gnd cell_6t
Xbit_r133_c200 bl[200] br[200] wl[133] vdd gnd cell_6t
Xbit_r134_c200 bl[200] br[200] wl[134] vdd gnd cell_6t
Xbit_r135_c200 bl[200] br[200] wl[135] vdd gnd cell_6t
Xbit_r136_c200 bl[200] br[200] wl[136] vdd gnd cell_6t
Xbit_r137_c200 bl[200] br[200] wl[137] vdd gnd cell_6t
Xbit_r138_c200 bl[200] br[200] wl[138] vdd gnd cell_6t
Xbit_r139_c200 bl[200] br[200] wl[139] vdd gnd cell_6t
Xbit_r140_c200 bl[200] br[200] wl[140] vdd gnd cell_6t
Xbit_r141_c200 bl[200] br[200] wl[141] vdd gnd cell_6t
Xbit_r142_c200 bl[200] br[200] wl[142] vdd gnd cell_6t
Xbit_r143_c200 bl[200] br[200] wl[143] vdd gnd cell_6t
Xbit_r144_c200 bl[200] br[200] wl[144] vdd gnd cell_6t
Xbit_r145_c200 bl[200] br[200] wl[145] vdd gnd cell_6t
Xbit_r146_c200 bl[200] br[200] wl[146] vdd gnd cell_6t
Xbit_r147_c200 bl[200] br[200] wl[147] vdd gnd cell_6t
Xbit_r148_c200 bl[200] br[200] wl[148] vdd gnd cell_6t
Xbit_r149_c200 bl[200] br[200] wl[149] vdd gnd cell_6t
Xbit_r150_c200 bl[200] br[200] wl[150] vdd gnd cell_6t
Xbit_r151_c200 bl[200] br[200] wl[151] vdd gnd cell_6t
Xbit_r152_c200 bl[200] br[200] wl[152] vdd gnd cell_6t
Xbit_r153_c200 bl[200] br[200] wl[153] vdd gnd cell_6t
Xbit_r154_c200 bl[200] br[200] wl[154] vdd gnd cell_6t
Xbit_r155_c200 bl[200] br[200] wl[155] vdd gnd cell_6t
Xbit_r156_c200 bl[200] br[200] wl[156] vdd gnd cell_6t
Xbit_r157_c200 bl[200] br[200] wl[157] vdd gnd cell_6t
Xbit_r158_c200 bl[200] br[200] wl[158] vdd gnd cell_6t
Xbit_r159_c200 bl[200] br[200] wl[159] vdd gnd cell_6t
Xbit_r160_c200 bl[200] br[200] wl[160] vdd gnd cell_6t
Xbit_r161_c200 bl[200] br[200] wl[161] vdd gnd cell_6t
Xbit_r162_c200 bl[200] br[200] wl[162] vdd gnd cell_6t
Xbit_r163_c200 bl[200] br[200] wl[163] vdd gnd cell_6t
Xbit_r164_c200 bl[200] br[200] wl[164] vdd gnd cell_6t
Xbit_r165_c200 bl[200] br[200] wl[165] vdd gnd cell_6t
Xbit_r166_c200 bl[200] br[200] wl[166] vdd gnd cell_6t
Xbit_r167_c200 bl[200] br[200] wl[167] vdd gnd cell_6t
Xbit_r168_c200 bl[200] br[200] wl[168] vdd gnd cell_6t
Xbit_r169_c200 bl[200] br[200] wl[169] vdd gnd cell_6t
Xbit_r170_c200 bl[200] br[200] wl[170] vdd gnd cell_6t
Xbit_r171_c200 bl[200] br[200] wl[171] vdd gnd cell_6t
Xbit_r172_c200 bl[200] br[200] wl[172] vdd gnd cell_6t
Xbit_r173_c200 bl[200] br[200] wl[173] vdd gnd cell_6t
Xbit_r174_c200 bl[200] br[200] wl[174] vdd gnd cell_6t
Xbit_r175_c200 bl[200] br[200] wl[175] vdd gnd cell_6t
Xbit_r176_c200 bl[200] br[200] wl[176] vdd gnd cell_6t
Xbit_r177_c200 bl[200] br[200] wl[177] vdd gnd cell_6t
Xbit_r178_c200 bl[200] br[200] wl[178] vdd gnd cell_6t
Xbit_r179_c200 bl[200] br[200] wl[179] vdd gnd cell_6t
Xbit_r180_c200 bl[200] br[200] wl[180] vdd gnd cell_6t
Xbit_r181_c200 bl[200] br[200] wl[181] vdd gnd cell_6t
Xbit_r182_c200 bl[200] br[200] wl[182] vdd gnd cell_6t
Xbit_r183_c200 bl[200] br[200] wl[183] vdd gnd cell_6t
Xbit_r184_c200 bl[200] br[200] wl[184] vdd gnd cell_6t
Xbit_r185_c200 bl[200] br[200] wl[185] vdd gnd cell_6t
Xbit_r186_c200 bl[200] br[200] wl[186] vdd gnd cell_6t
Xbit_r187_c200 bl[200] br[200] wl[187] vdd gnd cell_6t
Xbit_r188_c200 bl[200] br[200] wl[188] vdd gnd cell_6t
Xbit_r189_c200 bl[200] br[200] wl[189] vdd gnd cell_6t
Xbit_r190_c200 bl[200] br[200] wl[190] vdd gnd cell_6t
Xbit_r191_c200 bl[200] br[200] wl[191] vdd gnd cell_6t
Xbit_r192_c200 bl[200] br[200] wl[192] vdd gnd cell_6t
Xbit_r193_c200 bl[200] br[200] wl[193] vdd gnd cell_6t
Xbit_r194_c200 bl[200] br[200] wl[194] vdd gnd cell_6t
Xbit_r195_c200 bl[200] br[200] wl[195] vdd gnd cell_6t
Xbit_r196_c200 bl[200] br[200] wl[196] vdd gnd cell_6t
Xbit_r197_c200 bl[200] br[200] wl[197] vdd gnd cell_6t
Xbit_r198_c200 bl[200] br[200] wl[198] vdd gnd cell_6t
Xbit_r199_c200 bl[200] br[200] wl[199] vdd gnd cell_6t
Xbit_r200_c200 bl[200] br[200] wl[200] vdd gnd cell_6t
Xbit_r201_c200 bl[200] br[200] wl[201] vdd gnd cell_6t
Xbit_r202_c200 bl[200] br[200] wl[202] vdd gnd cell_6t
Xbit_r203_c200 bl[200] br[200] wl[203] vdd gnd cell_6t
Xbit_r204_c200 bl[200] br[200] wl[204] vdd gnd cell_6t
Xbit_r205_c200 bl[200] br[200] wl[205] vdd gnd cell_6t
Xbit_r206_c200 bl[200] br[200] wl[206] vdd gnd cell_6t
Xbit_r207_c200 bl[200] br[200] wl[207] vdd gnd cell_6t
Xbit_r208_c200 bl[200] br[200] wl[208] vdd gnd cell_6t
Xbit_r209_c200 bl[200] br[200] wl[209] vdd gnd cell_6t
Xbit_r210_c200 bl[200] br[200] wl[210] vdd gnd cell_6t
Xbit_r211_c200 bl[200] br[200] wl[211] vdd gnd cell_6t
Xbit_r212_c200 bl[200] br[200] wl[212] vdd gnd cell_6t
Xbit_r213_c200 bl[200] br[200] wl[213] vdd gnd cell_6t
Xbit_r214_c200 bl[200] br[200] wl[214] vdd gnd cell_6t
Xbit_r215_c200 bl[200] br[200] wl[215] vdd gnd cell_6t
Xbit_r216_c200 bl[200] br[200] wl[216] vdd gnd cell_6t
Xbit_r217_c200 bl[200] br[200] wl[217] vdd gnd cell_6t
Xbit_r218_c200 bl[200] br[200] wl[218] vdd gnd cell_6t
Xbit_r219_c200 bl[200] br[200] wl[219] vdd gnd cell_6t
Xbit_r220_c200 bl[200] br[200] wl[220] vdd gnd cell_6t
Xbit_r221_c200 bl[200] br[200] wl[221] vdd gnd cell_6t
Xbit_r222_c200 bl[200] br[200] wl[222] vdd gnd cell_6t
Xbit_r223_c200 bl[200] br[200] wl[223] vdd gnd cell_6t
Xbit_r224_c200 bl[200] br[200] wl[224] vdd gnd cell_6t
Xbit_r225_c200 bl[200] br[200] wl[225] vdd gnd cell_6t
Xbit_r226_c200 bl[200] br[200] wl[226] vdd gnd cell_6t
Xbit_r227_c200 bl[200] br[200] wl[227] vdd gnd cell_6t
Xbit_r228_c200 bl[200] br[200] wl[228] vdd gnd cell_6t
Xbit_r229_c200 bl[200] br[200] wl[229] vdd gnd cell_6t
Xbit_r230_c200 bl[200] br[200] wl[230] vdd gnd cell_6t
Xbit_r231_c200 bl[200] br[200] wl[231] vdd gnd cell_6t
Xbit_r232_c200 bl[200] br[200] wl[232] vdd gnd cell_6t
Xbit_r233_c200 bl[200] br[200] wl[233] vdd gnd cell_6t
Xbit_r234_c200 bl[200] br[200] wl[234] vdd gnd cell_6t
Xbit_r235_c200 bl[200] br[200] wl[235] vdd gnd cell_6t
Xbit_r236_c200 bl[200] br[200] wl[236] vdd gnd cell_6t
Xbit_r237_c200 bl[200] br[200] wl[237] vdd gnd cell_6t
Xbit_r238_c200 bl[200] br[200] wl[238] vdd gnd cell_6t
Xbit_r239_c200 bl[200] br[200] wl[239] vdd gnd cell_6t
Xbit_r240_c200 bl[200] br[200] wl[240] vdd gnd cell_6t
Xbit_r241_c200 bl[200] br[200] wl[241] vdd gnd cell_6t
Xbit_r242_c200 bl[200] br[200] wl[242] vdd gnd cell_6t
Xbit_r243_c200 bl[200] br[200] wl[243] vdd gnd cell_6t
Xbit_r244_c200 bl[200] br[200] wl[244] vdd gnd cell_6t
Xbit_r245_c200 bl[200] br[200] wl[245] vdd gnd cell_6t
Xbit_r246_c200 bl[200] br[200] wl[246] vdd gnd cell_6t
Xbit_r247_c200 bl[200] br[200] wl[247] vdd gnd cell_6t
Xbit_r248_c200 bl[200] br[200] wl[248] vdd gnd cell_6t
Xbit_r249_c200 bl[200] br[200] wl[249] vdd gnd cell_6t
Xbit_r250_c200 bl[200] br[200] wl[250] vdd gnd cell_6t
Xbit_r251_c200 bl[200] br[200] wl[251] vdd gnd cell_6t
Xbit_r252_c200 bl[200] br[200] wl[252] vdd gnd cell_6t
Xbit_r253_c200 bl[200] br[200] wl[253] vdd gnd cell_6t
Xbit_r254_c200 bl[200] br[200] wl[254] vdd gnd cell_6t
Xbit_r255_c200 bl[200] br[200] wl[255] vdd gnd cell_6t
Xbit_r0_c201 bl[201] br[201] wl[0] vdd gnd cell_6t
Xbit_r1_c201 bl[201] br[201] wl[1] vdd gnd cell_6t
Xbit_r2_c201 bl[201] br[201] wl[2] vdd gnd cell_6t
Xbit_r3_c201 bl[201] br[201] wl[3] vdd gnd cell_6t
Xbit_r4_c201 bl[201] br[201] wl[4] vdd gnd cell_6t
Xbit_r5_c201 bl[201] br[201] wl[5] vdd gnd cell_6t
Xbit_r6_c201 bl[201] br[201] wl[6] vdd gnd cell_6t
Xbit_r7_c201 bl[201] br[201] wl[7] vdd gnd cell_6t
Xbit_r8_c201 bl[201] br[201] wl[8] vdd gnd cell_6t
Xbit_r9_c201 bl[201] br[201] wl[9] vdd gnd cell_6t
Xbit_r10_c201 bl[201] br[201] wl[10] vdd gnd cell_6t
Xbit_r11_c201 bl[201] br[201] wl[11] vdd gnd cell_6t
Xbit_r12_c201 bl[201] br[201] wl[12] vdd gnd cell_6t
Xbit_r13_c201 bl[201] br[201] wl[13] vdd gnd cell_6t
Xbit_r14_c201 bl[201] br[201] wl[14] vdd gnd cell_6t
Xbit_r15_c201 bl[201] br[201] wl[15] vdd gnd cell_6t
Xbit_r16_c201 bl[201] br[201] wl[16] vdd gnd cell_6t
Xbit_r17_c201 bl[201] br[201] wl[17] vdd gnd cell_6t
Xbit_r18_c201 bl[201] br[201] wl[18] vdd gnd cell_6t
Xbit_r19_c201 bl[201] br[201] wl[19] vdd gnd cell_6t
Xbit_r20_c201 bl[201] br[201] wl[20] vdd gnd cell_6t
Xbit_r21_c201 bl[201] br[201] wl[21] vdd gnd cell_6t
Xbit_r22_c201 bl[201] br[201] wl[22] vdd gnd cell_6t
Xbit_r23_c201 bl[201] br[201] wl[23] vdd gnd cell_6t
Xbit_r24_c201 bl[201] br[201] wl[24] vdd gnd cell_6t
Xbit_r25_c201 bl[201] br[201] wl[25] vdd gnd cell_6t
Xbit_r26_c201 bl[201] br[201] wl[26] vdd gnd cell_6t
Xbit_r27_c201 bl[201] br[201] wl[27] vdd gnd cell_6t
Xbit_r28_c201 bl[201] br[201] wl[28] vdd gnd cell_6t
Xbit_r29_c201 bl[201] br[201] wl[29] vdd gnd cell_6t
Xbit_r30_c201 bl[201] br[201] wl[30] vdd gnd cell_6t
Xbit_r31_c201 bl[201] br[201] wl[31] vdd gnd cell_6t
Xbit_r32_c201 bl[201] br[201] wl[32] vdd gnd cell_6t
Xbit_r33_c201 bl[201] br[201] wl[33] vdd gnd cell_6t
Xbit_r34_c201 bl[201] br[201] wl[34] vdd gnd cell_6t
Xbit_r35_c201 bl[201] br[201] wl[35] vdd gnd cell_6t
Xbit_r36_c201 bl[201] br[201] wl[36] vdd gnd cell_6t
Xbit_r37_c201 bl[201] br[201] wl[37] vdd gnd cell_6t
Xbit_r38_c201 bl[201] br[201] wl[38] vdd gnd cell_6t
Xbit_r39_c201 bl[201] br[201] wl[39] vdd gnd cell_6t
Xbit_r40_c201 bl[201] br[201] wl[40] vdd gnd cell_6t
Xbit_r41_c201 bl[201] br[201] wl[41] vdd gnd cell_6t
Xbit_r42_c201 bl[201] br[201] wl[42] vdd gnd cell_6t
Xbit_r43_c201 bl[201] br[201] wl[43] vdd gnd cell_6t
Xbit_r44_c201 bl[201] br[201] wl[44] vdd gnd cell_6t
Xbit_r45_c201 bl[201] br[201] wl[45] vdd gnd cell_6t
Xbit_r46_c201 bl[201] br[201] wl[46] vdd gnd cell_6t
Xbit_r47_c201 bl[201] br[201] wl[47] vdd gnd cell_6t
Xbit_r48_c201 bl[201] br[201] wl[48] vdd gnd cell_6t
Xbit_r49_c201 bl[201] br[201] wl[49] vdd gnd cell_6t
Xbit_r50_c201 bl[201] br[201] wl[50] vdd gnd cell_6t
Xbit_r51_c201 bl[201] br[201] wl[51] vdd gnd cell_6t
Xbit_r52_c201 bl[201] br[201] wl[52] vdd gnd cell_6t
Xbit_r53_c201 bl[201] br[201] wl[53] vdd gnd cell_6t
Xbit_r54_c201 bl[201] br[201] wl[54] vdd gnd cell_6t
Xbit_r55_c201 bl[201] br[201] wl[55] vdd gnd cell_6t
Xbit_r56_c201 bl[201] br[201] wl[56] vdd gnd cell_6t
Xbit_r57_c201 bl[201] br[201] wl[57] vdd gnd cell_6t
Xbit_r58_c201 bl[201] br[201] wl[58] vdd gnd cell_6t
Xbit_r59_c201 bl[201] br[201] wl[59] vdd gnd cell_6t
Xbit_r60_c201 bl[201] br[201] wl[60] vdd gnd cell_6t
Xbit_r61_c201 bl[201] br[201] wl[61] vdd gnd cell_6t
Xbit_r62_c201 bl[201] br[201] wl[62] vdd gnd cell_6t
Xbit_r63_c201 bl[201] br[201] wl[63] vdd gnd cell_6t
Xbit_r64_c201 bl[201] br[201] wl[64] vdd gnd cell_6t
Xbit_r65_c201 bl[201] br[201] wl[65] vdd gnd cell_6t
Xbit_r66_c201 bl[201] br[201] wl[66] vdd gnd cell_6t
Xbit_r67_c201 bl[201] br[201] wl[67] vdd gnd cell_6t
Xbit_r68_c201 bl[201] br[201] wl[68] vdd gnd cell_6t
Xbit_r69_c201 bl[201] br[201] wl[69] vdd gnd cell_6t
Xbit_r70_c201 bl[201] br[201] wl[70] vdd gnd cell_6t
Xbit_r71_c201 bl[201] br[201] wl[71] vdd gnd cell_6t
Xbit_r72_c201 bl[201] br[201] wl[72] vdd gnd cell_6t
Xbit_r73_c201 bl[201] br[201] wl[73] vdd gnd cell_6t
Xbit_r74_c201 bl[201] br[201] wl[74] vdd gnd cell_6t
Xbit_r75_c201 bl[201] br[201] wl[75] vdd gnd cell_6t
Xbit_r76_c201 bl[201] br[201] wl[76] vdd gnd cell_6t
Xbit_r77_c201 bl[201] br[201] wl[77] vdd gnd cell_6t
Xbit_r78_c201 bl[201] br[201] wl[78] vdd gnd cell_6t
Xbit_r79_c201 bl[201] br[201] wl[79] vdd gnd cell_6t
Xbit_r80_c201 bl[201] br[201] wl[80] vdd gnd cell_6t
Xbit_r81_c201 bl[201] br[201] wl[81] vdd gnd cell_6t
Xbit_r82_c201 bl[201] br[201] wl[82] vdd gnd cell_6t
Xbit_r83_c201 bl[201] br[201] wl[83] vdd gnd cell_6t
Xbit_r84_c201 bl[201] br[201] wl[84] vdd gnd cell_6t
Xbit_r85_c201 bl[201] br[201] wl[85] vdd gnd cell_6t
Xbit_r86_c201 bl[201] br[201] wl[86] vdd gnd cell_6t
Xbit_r87_c201 bl[201] br[201] wl[87] vdd gnd cell_6t
Xbit_r88_c201 bl[201] br[201] wl[88] vdd gnd cell_6t
Xbit_r89_c201 bl[201] br[201] wl[89] vdd gnd cell_6t
Xbit_r90_c201 bl[201] br[201] wl[90] vdd gnd cell_6t
Xbit_r91_c201 bl[201] br[201] wl[91] vdd gnd cell_6t
Xbit_r92_c201 bl[201] br[201] wl[92] vdd gnd cell_6t
Xbit_r93_c201 bl[201] br[201] wl[93] vdd gnd cell_6t
Xbit_r94_c201 bl[201] br[201] wl[94] vdd gnd cell_6t
Xbit_r95_c201 bl[201] br[201] wl[95] vdd gnd cell_6t
Xbit_r96_c201 bl[201] br[201] wl[96] vdd gnd cell_6t
Xbit_r97_c201 bl[201] br[201] wl[97] vdd gnd cell_6t
Xbit_r98_c201 bl[201] br[201] wl[98] vdd gnd cell_6t
Xbit_r99_c201 bl[201] br[201] wl[99] vdd gnd cell_6t
Xbit_r100_c201 bl[201] br[201] wl[100] vdd gnd cell_6t
Xbit_r101_c201 bl[201] br[201] wl[101] vdd gnd cell_6t
Xbit_r102_c201 bl[201] br[201] wl[102] vdd gnd cell_6t
Xbit_r103_c201 bl[201] br[201] wl[103] vdd gnd cell_6t
Xbit_r104_c201 bl[201] br[201] wl[104] vdd gnd cell_6t
Xbit_r105_c201 bl[201] br[201] wl[105] vdd gnd cell_6t
Xbit_r106_c201 bl[201] br[201] wl[106] vdd gnd cell_6t
Xbit_r107_c201 bl[201] br[201] wl[107] vdd gnd cell_6t
Xbit_r108_c201 bl[201] br[201] wl[108] vdd gnd cell_6t
Xbit_r109_c201 bl[201] br[201] wl[109] vdd gnd cell_6t
Xbit_r110_c201 bl[201] br[201] wl[110] vdd gnd cell_6t
Xbit_r111_c201 bl[201] br[201] wl[111] vdd gnd cell_6t
Xbit_r112_c201 bl[201] br[201] wl[112] vdd gnd cell_6t
Xbit_r113_c201 bl[201] br[201] wl[113] vdd gnd cell_6t
Xbit_r114_c201 bl[201] br[201] wl[114] vdd gnd cell_6t
Xbit_r115_c201 bl[201] br[201] wl[115] vdd gnd cell_6t
Xbit_r116_c201 bl[201] br[201] wl[116] vdd gnd cell_6t
Xbit_r117_c201 bl[201] br[201] wl[117] vdd gnd cell_6t
Xbit_r118_c201 bl[201] br[201] wl[118] vdd gnd cell_6t
Xbit_r119_c201 bl[201] br[201] wl[119] vdd gnd cell_6t
Xbit_r120_c201 bl[201] br[201] wl[120] vdd gnd cell_6t
Xbit_r121_c201 bl[201] br[201] wl[121] vdd gnd cell_6t
Xbit_r122_c201 bl[201] br[201] wl[122] vdd gnd cell_6t
Xbit_r123_c201 bl[201] br[201] wl[123] vdd gnd cell_6t
Xbit_r124_c201 bl[201] br[201] wl[124] vdd gnd cell_6t
Xbit_r125_c201 bl[201] br[201] wl[125] vdd gnd cell_6t
Xbit_r126_c201 bl[201] br[201] wl[126] vdd gnd cell_6t
Xbit_r127_c201 bl[201] br[201] wl[127] vdd gnd cell_6t
Xbit_r128_c201 bl[201] br[201] wl[128] vdd gnd cell_6t
Xbit_r129_c201 bl[201] br[201] wl[129] vdd gnd cell_6t
Xbit_r130_c201 bl[201] br[201] wl[130] vdd gnd cell_6t
Xbit_r131_c201 bl[201] br[201] wl[131] vdd gnd cell_6t
Xbit_r132_c201 bl[201] br[201] wl[132] vdd gnd cell_6t
Xbit_r133_c201 bl[201] br[201] wl[133] vdd gnd cell_6t
Xbit_r134_c201 bl[201] br[201] wl[134] vdd gnd cell_6t
Xbit_r135_c201 bl[201] br[201] wl[135] vdd gnd cell_6t
Xbit_r136_c201 bl[201] br[201] wl[136] vdd gnd cell_6t
Xbit_r137_c201 bl[201] br[201] wl[137] vdd gnd cell_6t
Xbit_r138_c201 bl[201] br[201] wl[138] vdd gnd cell_6t
Xbit_r139_c201 bl[201] br[201] wl[139] vdd gnd cell_6t
Xbit_r140_c201 bl[201] br[201] wl[140] vdd gnd cell_6t
Xbit_r141_c201 bl[201] br[201] wl[141] vdd gnd cell_6t
Xbit_r142_c201 bl[201] br[201] wl[142] vdd gnd cell_6t
Xbit_r143_c201 bl[201] br[201] wl[143] vdd gnd cell_6t
Xbit_r144_c201 bl[201] br[201] wl[144] vdd gnd cell_6t
Xbit_r145_c201 bl[201] br[201] wl[145] vdd gnd cell_6t
Xbit_r146_c201 bl[201] br[201] wl[146] vdd gnd cell_6t
Xbit_r147_c201 bl[201] br[201] wl[147] vdd gnd cell_6t
Xbit_r148_c201 bl[201] br[201] wl[148] vdd gnd cell_6t
Xbit_r149_c201 bl[201] br[201] wl[149] vdd gnd cell_6t
Xbit_r150_c201 bl[201] br[201] wl[150] vdd gnd cell_6t
Xbit_r151_c201 bl[201] br[201] wl[151] vdd gnd cell_6t
Xbit_r152_c201 bl[201] br[201] wl[152] vdd gnd cell_6t
Xbit_r153_c201 bl[201] br[201] wl[153] vdd gnd cell_6t
Xbit_r154_c201 bl[201] br[201] wl[154] vdd gnd cell_6t
Xbit_r155_c201 bl[201] br[201] wl[155] vdd gnd cell_6t
Xbit_r156_c201 bl[201] br[201] wl[156] vdd gnd cell_6t
Xbit_r157_c201 bl[201] br[201] wl[157] vdd gnd cell_6t
Xbit_r158_c201 bl[201] br[201] wl[158] vdd gnd cell_6t
Xbit_r159_c201 bl[201] br[201] wl[159] vdd gnd cell_6t
Xbit_r160_c201 bl[201] br[201] wl[160] vdd gnd cell_6t
Xbit_r161_c201 bl[201] br[201] wl[161] vdd gnd cell_6t
Xbit_r162_c201 bl[201] br[201] wl[162] vdd gnd cell_6t
Xbit_r163_c201 bl[201] br[201] wl[163] vdd gnd cell_6t
Xbit_r164_c201 bl[201] br[201] wl[164] vdd gnd cell_6t
Xbit_r165_c201 bl[201] br[201] wl[165] vdd gnd cell_6t
Xbit_r166_c201 bl[201] br[201] wl[166] vdd gnd cell_6t
Xbit_r167_c201 bl[201] br[201] wl[167] vdd gnd cell_6t
Xbit_r168_c201 bl[201] br[201] wl[168] vdd gnd cell_6t
Xbit_r169_c201 bl[201] br[201] wl[169] vdd gnd cell_6t
Xbit_r170_c201 bl[201] br[201] wl[170] vdd gnd cell_6t
Xbit_r171_c201 bl[201] br[201] wl[171] vdd gnd cell_6t
Xbit_r172_c201 bl[201] br[201] wl[172] vdd gnd cell_6t
Xbit_r173_c201 bl[201] br[201] wl[173] vdd gnd cell_6t
Xbit_r174_c201 bl[201] br[201] wl[174] vdd gnd cell_6t
Xbit_r175_c201 bl[201] br[201] wl[175] vdd gnd cell_6t
Xbit_r176_c201 bl[201] br[201] wl[176] vdd gnd cell_6t
Xbit_r177_c201 bl[201] br[201] wl[177] vdd gnd cell_6t
Xbit_r178_c201 bl[201] br[201] wl[178] vdd gnd cell_6t
Xbit_r179_c201 bl[201] br[201] wl[179] vdd gnd cell_6t
Xbit_r180_c201 bl[201] br[201] wl[180] vdd gnd cell_6t
Xbit_r181_c201 bl[201] br[201] wl[181] vdd gnd cell_6t
Xbit_r182_c201 bl[201] br[201] wl[182] vdd gnd cell_6t
Xbit_r183_c201 bl[201] br[201] wl[183] vdd gnd cell_6t
Xbit_r184_c201 bl[201] br[201] wl[184] vdd gnd cell_6t
Xbit_r185_c201 bl[201] br[201] wl[185] vdd gnd cell_6t
Xbit_r186_c201 bl[201] br[201] wl[186] vdd gnd cell_6t
Xbit_r187_c201 bl[201] br[201] wl[187] vdd gnd cell_6t
Xbit_r188_c201 bl[201] br[201] wl[188] vdd gnd cell_6t
Xbit_r189_c201 bl[201] br[201] wl[189] vdd gnd cell_6t
Xbit_r190_c201 bl[201] br[201] wl[190] vdd gnd cell_6t
Xbit_r191_c201 bl[201] br[201] wl[191] vdd gnd cell_6t
Xbit_r192_c201 bl[201] br[201] wl[192] vdd gnd cell_6t
Xbit_r193_c201 bl[201] br[201] wl[193] vdd gnd cell_6t
Xbit_r194_c201 bl[201] br[201] wl[194] vdd gnd cell_6t
Xbit_r195_c201 bl[201] br[201] wl[195] vdd gnd cell_6t
Xbit_r196_c201 bl[201] br[201] wl[196] vdd gnd cell_6t
Xbit_r197_c201 bl[201] br[201] wl[197] vdd gnd cell_6t
Xbit_r198_c201 bl[201] br[201] wl[198] vdd gnd cell_6t
Xbit_r199_c201 bl[201] br[201] wl[199] vdd gnd cell_6t
Xbit_r200_c201 bl[201] br[201] wl[200] vdd gnd cell_6t
Xbit_r201_c201 bl[201] br[201] wl[201] vdd gnd cell_6t
Xbit_r202_c201 bl[201] br[201] wl[202] vdd gnd cell_6t
Xbit_r203_c201 bl[201] br[201] wl[203] vdd gnd cell_6t
Xbit_r204_c201 bl[201] br[201] wl[204] vdd gnd cell_6t
Xbit_r205_c201 bl[201] br[201] wl[205] vdd gnd cell_6t
Xbit_r206_c201 bl[201] br[201] wl[206] vdd gnd cell_6t
Xbit_r207_c201 bl[201] br[201] wl[207] vdd gnd cell_6t
Xbit_r208_c201 bl[201] br[201] wl[208] vdd gnd cell_6t
Xbit_r209_c201 bl[201] br[201] wl[209] vdd gnd cell_6t
Xbit_r210_c201 bl[201] br[201] wl[210] vdd gnd cell_6t
Xbit_r211_c201 bl[201] br[201] wl[211] vdd gnd cell_6t
Xbit_r212_c201 bl[201] br[201] wl[212] vdd gnd cell_6t
Xbit_r213_c201 bl[201] br[201] wl[213] vdd gnd cell_6t
Xbit_r214_c201 bl[201] br[201] wl[214] vdd gnd cell_6t
Xbit_r215_c201 bl[201] br[201] wl[215] vdd gnd cell_6t
Xbit_r216_c201 bl[201] br[201] wl[216] vdd gnd cell_6t
Xbit_r217_c201 bl[201] br[201] wl[217] vdd gnd cell_6t
Xbit_r218_c201 bl[201] br[201] wl[218] vdd gnd cell_6t
Xbit_r219_c201 bl[201] br[201] wl[219] vdd gnd cell_6t
Xbit_r220_c201 bl[201] br[201] wl[220] vdd gnd cell_6t
Xbit_r221_c201 bl[201] br[201] wl[221] vdd gnd cell_6t
Xbit_r222_c201 bl[201] br[201] wl[222] vdd gnd cell_6t
Xbit_r223_c201 bl[201] br[201] wl[223] vdd gnd cell_6t
Xbit_r224_c201 bl[201] br[201] wl[224] vdd gnd cell_6t
Xbit_r225_c201 bl[201] br[201] wl[225] vdd gnd cell_6t
Xbit_r226_c201 bl[201] br[201] wl[226] vdd gnd cell_6t
Xbit_r227_c201 bl[201] br[201] wl[227] vdd gnd cell_6t
Xbit_r228_c201 bl[201] br[201] wl[228] vdd gnd cell_6t
Xbit_r229_c201 bl[201] br[201] wl[229] vdd gnd cell_6t
Xbit_r230_c201 bl[201] br[201] wl[230] vdd gnd cell_6t
Xbit_r231_c201 bl[201] br[201] wl[231] vdd gnd cell_6t
Xbit_r232_c201 bl[201] br[201] wl[232] vdd gnd cell_6t
Xbit_r233_c201 bl[201] br[201] wl[233] vdd gnd cell_6t
Xbit_r234_c201 bl[201] br[201] wl[234] vdd gnd cell_6t
Xbit_r235_c201 bl[201] br[201] wl[235] vdd gnd cell_6t
Xbit_r236_c201 bl[201] br[201] wl[236] vdd gnd cell_6t
Xbit_r237_c201 bl[201] br[201] wl[237] vdd gnd cell_6t
Xbit_r238_c201 bl[201] br[201] wl[238] vdd gnd cell_6t
Xbit_r239_c201 bl[201] br[201] wl[239] vdd gnd cell_6t
Xbit_r240_c201 bl[201] br[201] wl[240] vdd gnd cell_6t
Xbit_r241_c201 bl[201] br[201] wl[241] vdd gnd cell_6t
Xbit_r242_c201 bl[201] br[201] wl[242] vdd gnd cell_6t
Xbit_r243_c201 bl[201] br[201] wl[243] vdd gnd cell_6t
Xbit_r244_c201 bl[201] br[201] wl[244] vdd gnd cell_6t
Xbit_r245_c201 bl[201] br[201] wl[245] vdd gnd cell_6t
Xbit_r246_c201 bl[201] br[201] wl[246] vdd gnd cell_6t
Xbit_r247_c201 bl[201] br[201] wl[247] vdd gnd cell_6t
Xbit_r248_c201 bl[201] br[201] wl[248] vdd gnd cell_6t
Xbit_r249_c201 bl[201] br[201] wl[249] vdd gnd cell_6t
Xbit_r250_c201 bl[201] br[201] wl[250] vdd gnd cell_6t
Xbit_r251_c201 bl[201] br[201] wl[251] vdd gnd cell_6t
Xbit_r252_c201 bl[201] br[201] wl[252] vdd gnd cell_6t
Xbit_r253_c201 bl[201] br[201] wl[253] vdd gnd cell_6t
Xbit_r254_c201 bl[201] br[201] wl[254] vdd gnd cell_6t
Xbit_r255_c201 bl[201] br[201] wl[255] vdd gnd cell_6t
Xbit_r0_c202 bl[202] br[202] wl[0] vdd gnd cell_6t
Xbit_r1_c202 bl[202] br[202] wl[1] vdd gnd cell_6t
Xbit_r2_c202 bl[202] br[202] wl[2] vdd gnd cell_6t
Xbit_r3_c202 bl[202] br[202] wl[3] vdd gnd cell_6t
Xbit_r4_c202 bl[202] br[202] wl[4] vdd gnd cell_6t
Xbit_r5_c202 bl[202] br[202] wl[5] vdd gnd cell_6t
Xbit_r6_c202 bl[202] br[202] wl[6] vdd gnd cell_6t
Xbit_r7_c202 bl[202] br[202] wl[7] vdd gnd cell_6t
Xbit_r8_c202 bl[202] br[202] wl[8] vdd gnd cell_6t
Xbit_r9_c202 bl[202] br[202] wl[9] vdd gnd cell_6t
Xbit_r10_c202 bl[202] br[202] wl[10] vdd gnd cell_6t
Xbit_r11_c202 bl[202] br[202] wl[11] vdd gnd cell_6t
Xbit_r12_c202 bl[202] br[202] wl[12] vdd gnd cell_6t
Xbit_r13_c202 bl[202] br[202] wl[13] vdd gnd cell_6t
Xbit_r14_c202 bl[202] br[202] wl[14] vdd gnd cell_6t
Xbit_r15_c202 bl[202] br[202] wl[15] vdd gnd cell_6t
Xbit_r16_c202 bl[202] br[202] wl[16] vdd gnd cell_6t
Xbit_r17_c202 bl[202] br[202] wl[17] vdd gnd cell_6t
Xbit_r18_c202 bl[202] br[202] wl[18] vdd gnd cell_6t
Xbit_r19_c202 bl[202] br[202] wl[19] vdd gnd cell_6t
Xbit_r20_c202 bl[202] br[202] wl[20] vdd gnd cell_6t
Xbit_r21_c202 bl[202] br[202] wl[21] vdd gnd cell_6t
Xbit_r22_c202 bl[202] br[202] wl[22] vdd gnd cell_6t
Xbit_r23_c202 bl[202] br[202] wl[23] vdd gnd cell_6t
Xbit_r24_c202 bl[202] br[202] wl[24] vdd gnd cell_6t
Xbit_r25_c202 bl[202] br[202] wl[25] vdd gnd cell_6t
Xbit_r26_c202 bl[202] br[202] wl[26] vdd gnd cell_6t
Xbit_r27_c202 bl[202] br[202] wl[27] vdd gnd cell_6t
Xbit_r28_c202 bl[202] br[202] wl[28] vdd gnd cell_6t
Xbit_r29_c202 bl[202] br[202] wl[29] vdd gnd cell_6t
Xbit_r30_c202 bl[202] br[202] wl[30] vdd gnd cell_6t
Xbit_r31_c202 bl[202] br[202] wl[31] vdd gnd cell_6t
Xbit_r32_c202 bl[202] br[202] wl[32] vdd gnd cell_6t
Xbit_r33_c202 bl[202] br[202] wl[33] vdd gnd cell_6t
Xbit_r34_c202 bl[202] br[202] wl[34] vdd gnd cell_6t
Xbit_r35_c202 bl[202] br[202] wl[35] vdd gnd cell_6t
Xbit_r36_c202 bl[202] br[202] wl[36] vdd gnd cell_6t
Xbit_r37_c202 bl[202] br[202] wl[37] vdd gnd cell_6t
Xbit_r38_c202 bl[202] br[202] wl[38] vdd gnd cell_6t
Xbit_r39_c202 bl[202] br[202] wl[39] vdd gnd cell_6t
Xbit_r40_c202 bl[202] br[202] wl[40] vdd gnd cell_6t
Xbit_r41_c202 bl[202] br[202] wl[41] vdd gnd cell_6t
Xbit_r42_c202 bl[202] br[202] wl[42] vdd gnd cell_6t
Xbit_r43_c202 bl[202] br[202] wl[43] vdd gnd cell_6t
Xbit_r44_c202 bl[202] br[202] wl[44] vdd gnd cell_6t
Xbit_r45_c202 bl[202] br[202] wl[45] vdd gnd cell_6t
Xbit_r46_c202 bl[202] br[202] wl[46] vdd gnd cell_6t
Xbit_r47_c202 bl[202] br[202] wl[47] vdd gnd cell_6t
Xbit_r48_c202 bl[202] br[202] wl[48] vdd gnd cell_6t
Xbit_r49_c202 bl[202] br[202] wl[49] vdd gnd cell_6t
Xbit_r50_c202 bl[202] br[202] wl[50] vdd gnd cell_6t
Xbit_r51_c202 bl[202] br[202] wl[51] vdd gnd cell_6t
Xbit_r52_c202 bl[202] br[202] wl[52] vdd gnd cell_6t
Xbit_r53_c202 bl[202] br[202] wl[53] vdd gnd cell_6t
Xbit_r54_c202 bl[202] br[202] wl[54] vdd gnd cell_6t
Xbit_r55_c202 bl[202] br[202] wl[55] vdd gnd cell_6t
Xbit_r56_c202 bl[202] br[202] wl[56] vdd gnd cell_6t
Xbit_r57_c202 bl[202] br[202] wl[57] vdd gnd cell_6t
Xbit_r58_c202 bl[202] br[202] wl[58] vdd gnd cell_6t
Xbit_r59_c202 bl[202] br[202] wl[59] vdd gnd cell_6t
Xbit_r60_c202 bl[202] br[202] wl[60] vdd gnd cell_6t
Xbit_r61_c202 bl[202] br[202] wl[61] vdd gnd cell_6t
Xbit_r62_c202 bl[202] br[202] wl[62] vdd gnd cell_6t
Xbit_r63_c202 bl[202] br[202] wl[63] vdd gnd cell_6t
Xbit_r64_c202 bl[202] br[202] wl[64] vdd gnd cell_6t
Xbit_r65_c202 bl[202] br[202] wl[65] vdd gnd cell_6t
Xbit_r66_c202 bl[202] br[202] wl[66] vdd gnd cell_6t
Xbit_r67_c202 bl[202] br[202] wl[67] vdd gnd cell_6t
Xbit_r68_c202 bl[202] br[202] wl[68] vdd gnd cell_6t
Xbit_r69_c202 bl[202] br[202] wl[69] vdd gnd cell_6t
Xbit_r70_c202 bl[202] br[202] wl[70] vdd gnd cell_6t
Xbit_r71_c202 bl[202] br[202] wl[71] vdd gnd cell_6t
Xbit_r72_c202 bl[202] br[202] wl[72] vdd gnd cell_6t
Xbit_r73_c202 bl[202] br[202] wl[73] vdd gnd cell_6t
Xbit_r74_c202 bl[202] br[202] wl[74] vdd gnd cell_6t
Xbit_r75_c202 bl[202] br[202] wl[75] vdd gnd cell_6t
Xbit_r76_c202 bl[202] br[202] wl[76] vdd gnd cell_6t
Xbit_r77_c202 bl[202] br[202] wl[77] vdd gnd cell_6t
Xbit_r78_c202 bl[202] br[202] wl[78] vdd gnd cell_6t
Xbit_r79_c202 bl[202] br[202] wl[79] vdd gnd cell_6t
Xbit_r80_c202 bl[202] br[202] wl[80] vdd gnd cell_6t
Xbit_r81_c202 bl[202] br[202] wl[81] vdd gnd cell_6t
Xbit_r82_c202 bl[202] br[202] wl[82] vdd gnd cell_6t
Xbit_r83_c202 bl[202] br[202] wl[83] vdd gnd cell_6t
Xbit_r84_c202 bl[202] br[202] wl[84] vdd gnd cell_6t
Xbit_r85_c202 bl[202] br[202] wl[85] vdd gnd cell_6t
Xbit_r86_c202 bl[202] br[202] wl[86] vdd gnd cell_6t
Xbit_r87_c202 bl[202] br[202] wl[87] vdd gnd cell_6t
Xbit_r88_c202 bl[202] br[202] wl[88] vdd gnd cell_6t
Xbit_r89_c202 bl[202] br[202] wl[89] vdd gnd cell_6t
Xbit_r90_c202 bl[202] br[202] wl[90] vdd gnd cell_6t
Xbit_r91_c202 bl[202] br[202] wl[91] vdd gnd cell_6t
Xbit_r92_c202 bl[202] br[202] wl[92] vdd gnd cell_6t
Xbit_r93_c202 bl[202] br[202] wl[93] vdd gnd cell_6t
Xbit_r94_c202 bl[202] br[202] wl[94] vdd gnd cell_6t
Xbit_r95_c202 bl[202] br[202] wl[95] vdd gnd cell_6t
Xbit_r96_c202 bl[202] br[202] wl[96] vdd gnd cell_6t
Xbit_r97_c202 bl[202] br[202] wl[97] vdd gnd cell_6t
Xbit_r98_c202 bl[202] br[202] wl[98] vdd gnd cell_6t
Xbit_r99_c202 bl[202] br[202] wl[99] vdd gnd cell_6t
Xbit_r100_c202 bl[202] br[202] wl[100] vdd gnd cell_6t
Xbit_r101_c202 bl[202] br[202] wl[101] vdd gnd cell_6t
Xbit_r102_c202 bl[202] br[202] wl[102] vdd gnd cell_6t
Xbit_r103_c202 bl[202] br[202] wl[103] vdd gnd cell_6t
Xbit_r104_c202 bl[202] br[202] wl[104] vdd gnd cell_6t
Xbit_r105_c202 bl[202] br[202] wl[105] vdd gnd cell_6t
Xbit_r106_c202 bl[202] br[202] wl[106] vdd gnd cell_6t
Xbit_r107_c202 bl[202] br[202] wl[107] vdd gnd cell_6t
Xbit_r108_c202 bl[202] br[202] wl[108] vdd gnd cell_6t
Xbit_r109_c202 bl[202] br[202] wl[109] vdd gnd cell_6t
Xbit_r110_c202 bl[202] br[202] wl[110] vdd gnd cell_6t
Xbit_r111_c202 bl[202] br[202] wl[111] vdd gnd cell_6t
Xbit_r112_c202 bl[202] br[202] wl[112] vdd gnd cell_6t
Xbit_r113_c202 bl[202] br[202] wl[113] vdd gnd cell_6t
Xbit_r114_c202 bl[202] br[202] wl[114] vdd gnd cell_6t
Xbit_r115_c202 bl[202] br[202] wl[115] vdd gnd cell_6t
Xbit_r116_c202 bl[202] br[202] wl[116] vdd gnd cell_6t
Xbit_r117_c202 bl[202] br[202] wl[117] vdd gnd cell_6t
Xbit_r118_c202 bl[202] br[202] wl[118] vdd gnd cell_6t
Xbit_r119_c202 bl[202] br[202] wl[119] vdd gnd cell_6t
Xbit_r120_c202 bl[202] br[202] wl[120] vdd gnd cell_6t
Xbit_r121_c202 bl[202] br[202] wl[121] vdd gnd cell_6t
Xbit_r122_c202 bl[202] br[202] wl[122] vdd gnd cell_6t
Xbit_r123_c202 bl[202] br[202] wl[123] vdd gnd cell_6t
Xbit_r124_c202 bl[202] br[202] wl[124] vdd gnd cell_6t
Xbit_r125_c202 bl[202] br[202] wl[125] vdd gnd cell_6t
Xbit_r126_c202 bl[202] br[202] wl[126] vdd gnd cell_6t
Xbit_r127_c202 bl[202] br[202] wl[127] vdd gnd cell_6t
Xbit_r128_c202 bl[202] br[202] wl[128] vdd gnd cell_6t
Xbit_r129_c202 bl[202] br[202] wl[129] vdd gnd cell_6t
Xbit_r130_c202 bl[202] br[202] wl[130] vdd gnd cell_6t
Xbit_r131_c202 bl[202] br[202] wl[131] vdd gnd cell_6t
Xbit_r132_c202 bl[202] br[202] wl[132] vdd gnd cell_6t
Xbit_r133_c202 bl[202] br[202] wl[133] vdd gnd cell_6t
Xbit_r134_c202 bl[202] br[202] wl[134] vdd gnd cell_6t
Xbit_r135_c202 bl[202] br[202] wl[135] vdd gnd cell_6t
Xbit_r136_c202 bl[202] br[202] wl[136] vdd gnd cell_6t
Xbit_r137_c202 bl[202] br[202] wl[137] vdd gnd cell_6t
Xbit_r138_c202 bl[202] br[202] wl[138] vdd gnd cell_6t
Xbit_r139_c202 bl[202] br[202] wl[139] vdd gnd cell_6t
Xbit_r140_c202 bl[202] br[202] wl[140] vdd gnd cell_6t
Xbit_r141_c202 bl[202] br[202] wl[141] vdd gnd cell_6t
Xbit_r142_c202 bl[202] br[202] wl[142] vdd gnd cell_6t
Xbit_r143_c202 bl[202] br[202] wl[143] vdd gnd cell_6t
Xbit_r144_c202 bl[202] br[202] wl[144] vdd gnd cell_6t
Xbit_r145_c202 bl[202] br[202] wl[145] vdd gnd cell_6t
Xbit_r146_c202 bl[202] br[202] wl[146] vdd gnd cell_6t
Xbit_r147_c202 bl[202] br[202] wl[147] vdd gnd cell_6t
Xbit_r148_c202 bl[202] br[202] wl[148] vdd gnd cell_6t
Xbit_r149_c202 bl[202] br[202] wl[149] vdd gnd cell_6t
Xbit_r150_c202 bl[202] br[202] wl[150] vdd gnd cell_6t
Xbit_r151_c202 bl[202] br[202] wl[151] vdd gnd cell_6t
Xbit_r152_c202 bl[202] br[202] wl[152] vdd gnd cell_6t
Xbit_r153_c202 bl[202] br[202] wl[153] vdd gnd cell_6t
Xbit_r154_c202 bl[202] br[202] wl[154] vdd gnd cell_6t
Xbit_r155_c202 bl[202] br[202] wl[155] vdd gnd cell_6t
Xbit_r156_c202 bl[202] br[202] wl[156] vdd gnd cell_6t
Xbit_r157_c202 bl[202] br[202] wl[157] vdd gnd cell_6t
Xbit_r158_c202 bl[202] br[202] wl[158] vdd gnd cell_6t
Xbit_r159_c202 bl[202] br[202] wl[159] vdd gnd cell_6t
Xbit_r160_c202 bl[202] br[202] wl[160] vdd gnd cell_6t
Xbit_r161_c202 bl[202] br[202] wl[161] vdd gnd cell_6t
Xbit_r162_c202 bl[202] br[202] wl[162] vdd gnd cell_6t
Xbit_r163_c202 bl[202] br[202] wl[163] vdd gnd cell_6t
Xbit_r164_c202 bl[202] br[202] wl[164] vdd gnd cell_6t
Xbit_r165_c202 bl[202] br[202] wl[165] vdd gnd cell_6t
Xbit_r166_c202 bl[202] br[202] wl[166] vdd gnd cell_6t
Xbit_r167_c202 bl[202] br[202] wl[167] vdd gnd cell_6t
Xbit_r168_c202 bl[202] br[202] wl[168] vdd gnd cell_6t
Xbit_r169_c202 bl[202] br[202] wl[169] vdd gnd cell_6t
Xbit_r170_c202 bl[202] br[202] wl[170] vdd gnd cell_6t
Xbit_r171_c202 bl[202] br[202] wl[171] vdd gnd cell_6t
Xbit_r172_c202 bl[202] br[202] wl[172] vdd gnd cell_6t
Xbit_r173_c202 bl[202] br[202] wl[173] vdd gnd cell_6t
Xbit_r174_c202 bl[202] br[202] wl[174] vdd gnd cell_6t
Xbit_r175_c202 bl[202] br[202] wl[175] vdd gnd cell_6t
Xbit_r176_c202 bl[202] br[202] wl[176] vdd gnd cell_6t
Xbit_r177_c202 bl[202] br[202] wl[177] vdd gnd cell_6t
Xbit_r178_c202 bl[202] br[202] wl[178] vdd gnd cell_6t
Xbit_r179_c202 bl[202] br[202] wl[179] vdd gnd cell_6t
Xbit_r180_c202 bl[202] br[202] wl[180] vdd gnd cell_6t
Xbit_r181_c202 bl[202] br[202] wl[181] vdd gnd cell_6t
Xbit_r182_c202 bl[202] br[202] wl[182] vdd gnd cell_6t
Xbit_r183_c202 bl[202] br[202] wl[183] vdd gnd cell_6t
Xbit_r184_c202 bl[202] br[202] wl[184] vdd gnd cell_6t
Xbit_r185_c202 bl[202] br[202] wl[185] vdd gnd cell_6t
Xbit_r186_c202 bl[202] br[202] wl[186] vdd gnd cell_6t
Xbit_r187_c202 bl[202] br[202] wl[187] vdd gnd cell_6t
Xbit_r188_c202 bl[202] br[202] wl[188] vdd gnd cell_6t
Xbit_r189_c202 bl[202] br[202] wl[189] vdd gnd cell_6t
Xbit_r190_c202 bl[202] br[202] wl[190] vdd gnd cell_6t
Xbit_r191_c202 bl[202] br[202] wl[191] vdd gnd cell_6t
Xbit_r192_c202 bl[202] br[202] wl[192] vdd gnd cell_6t
Xbit_r193_c202 bl[202] br[202] wl[193] vdd gnd cell_6t
Xbit_r194_c202 bl[202] br[202] wl[194] vdd gnd cell_6t
Xbit_r195_c202 bl[202] br[202] wl[195] vdd gnd cell_6t
Xbit_r196_c202 bl[202] br[202] wl[196] vdd gnd cell_6t
Xbit_r197_c202 bl[202] br[202] wl[197] vdd gnd cell_6t
Xbit_r198_c202 bl[202] br[202] wl[198] vdd gnd cell_6t
Xbit_r199_c202 bl[202] br[202] wl[199] vdd gnd cell_6t
Xbit_r200_c202 bl[202] br[202] wl[200] vdd gnd cell_6t
Xbit_r201_c202 bl[202] br[202] wl[201] vdd gnd cell_6t
Xbit_r202_c202 bl[202] br[202] wl[202] vdd gnd cell_6t
Xbit_r203_c202 bl[202] br[202] wl[203] vdd gnd cell_6t
Xbit_r204_c202 bl[202] br[202] wl[204] vdd gnd cell_6t
Xbit_r205_c202 bl[202] br[202] wl[205] vdd gnd cell_6t
Xbit_r206_c202 bl[202] br[202] wl[206] vdd gnd cell_6t
Xbit_r207_c202 bl[202] br[202] wl[207] vdd gnd cell_6t
Xbit_r208_c202 bl[202] br[202] wl[208] vdd gnd cell_6t
Xbit_r209_c202 bl[202] br[202] wl[209] vdd gnd cell_6t
Xbit_r210_c202 bl[202] br[202] wl[210] vdd gnd cell_6t
Xbit_r211_c202 bl[202] br[202] wl[211] vdd gnd cell_6t
Xbit_r212_c202 bl[202] br[202] wl[212] vdd gnd cell_6t
Xbit_r213_c202 bl[202] br[202] wl[213] vdd gnd cell_6t
Xbit_r214_c202 bl[202] br[202] wl[214] vdd gnd cell_6t
Xbit_r215_c202 bl[202] br[202] wl[215] vdd gnd cell_6t
Xbit_r216_c202 bl[202] br[202] wl[216] vdd gnd cell_6t
Xbit_r217_c202 bl[202] br[202] wl[217] vdd gnd cell_6t
Xbit_r218_c202 bl[202] br[202] wl[218] vdd gnd cell_6t
Xbit_r219_c202 bl[202] br[202] wl[219] vdd gnd cell_6t
Xbit_r220_c202 bl[202] br[202] wl[220] vdd gnd cell_6t
Xbit_r221_c202 bl[202] br[202] wl[221] vdd gnd cell_6t
Xbit_r222_c202 bl[202] br[202] wl[222] vdd gnd cell_6t
Xbit_r223_c202 bl[202] br[202] wl[223] vdd gnd cell_6t
Xbit_r224_c202 bl[202] br[202] wl[224] vdd gnd cell_6t
Xbit_r225_c202 bl[202] br[202] wl[225] vdd gnd cell_6t
Xbit_r226_c202 bl[202] br[202] wl[226] vdd gnd cell_6t
Xbit_r227_c202 bl[202] br[202] wl[227] vdd gnd cell_6t
Xbit_r228_c202 bl[202] br[202] wl[228] vdd gnd cell_6t
Xbit_r229_c202 bl[202] br[202] wl[229] vdd gnd cell_6t
Xbit_r230_c202 bl[202] br[202] wl[230] vdd gnd cell_6t
Xbit_r231_c202 bl[202] br[202] wl[231] vdd gnd cell_6t
Xbit_r232_c202 bl[202] br[202] wl[232] vdd gnd cell_6t
Xbit_r233_c202 bl[202] br[202] wl[233] vdd gnd cell_6t
Xbit_r234_c202 bl[202] br[202] wl[234] vdd gnd cell_6t
Xbit_r235_c202 bl[202] br[202] wl[235] vdd gnd cell_6t
Xbit_r236_c202 bl[202] br[202] wl[236] vdd gnd cell_6t
Xbit_r237_c202 bl[202] br[202] wl[237] vdd gnd cell_6t
Xbit_r238_c202 bl[202] br[202] wl[238] vdd gnd cell_6t
Xbit_r239_c202 bl[202] br[202] wl[239] vdd gnd cell_6t
Xbit_r240_c202 bl[202] br[202] wl[240] vdd gnd cell_6t
Xbit_r241_c202 bl[202] br[202] wl[241] vdd gnd cell_6t
Xbit_r242_c202 bl[202] br[202] wl[242] vdd gnd cell_6t
Xbit_r243_c202 bl[202] br[202] wl[243] vdd gnd cell_6t
Xbit_r244_c202 bl[202] br[202] wl[244] vdd gnd cell_6t
Xbit_r245_c202 bl[202] br[202] wl[245] vdd gnd cell_6t
Xbit_r246_c202 bl[202] br[202] wl[246] vdd gnd cell_6t
Xbit_r247_c202 bl[202] br[202] wl[247] vdd gnd cell_6t
Xbit_r248_c202 bl[202] br[202] wl[248] vdd gnd cell_6t
Xbit_r249_c202 bl[202] br[202] wl[249] vdd gnd cell_6t
Xbit_r250_c202 bl[202] br[202] wl[250] vdd gnd cell_6t
Xbit_r251_c202 bl[202] br[202] wl[251] vdd gnd cell_6t
Xbit_r252_c202 bl[202] br[202] wl[252] vdd gnd cell_6t
Xbit_r253_c202 bl[202] br[202] wl[253] vdd gnd cell_6t
Xbit_r254_c202 bl[202] br[202] wl[254] vdd gnd cell_6t
Xbit_r255_c202 bl[202] br[202] wl[255] vdd gnd cell_6t
Xbit_r0_c203 bl[203] br[203] wl[0] vdd gnd cell_6t
Xbit_r1_c203 bl[203] br[203] wl[1] vdd gnd cell_6t
Xbit_r2_c203 bl[203] br[203] wl[2] vdd gnd cell_6t
Xbit_r3_c203 bl[203] br[203] wl[3] vdd gnd cell_6t
Xbit_r4_c203 bl[203] br[203] wl[4] vdd gnd cell_6t
Xbit_r5_c203 bl[203] br[203] wl[5] vdd gnd cell_6t
Xbit_r6_c203 bl[203] br[203] wl[6] vdd gnd cell_6t
Xbit_r7_c203 bl[203] br[203] wl[7] vdd gnd cell_6t
Xbit_r8_c203 bl[203] br[203] wl[8] vdd gnd cell_6t
Xbit_r9_c203 bl[203] br[203] wl[9] vdd gnd cell_6t
Xbit_r10_c203 bl[203] br[203] wl[10] vdd gnd cell_6t
Xbit_r11_c203 bl[203] br[203] wl[11] vdd gnd cell_6t
Xbit_r12_c203 bl[203] br[203] wl[12] vdd gnd cell_6t
Xbit_r13_c203 bl[203] br[203] wl[13] vdd gnd cell_6t
Xbit_r14_c203 bl[203] br[203] wl[14] vdd gnd cell_6t
Xbit_r15_c203 bl[203] br[203] wl[15] vdd gnd cell_6t
Xbit_r16_c203 bl[203] br[203] wl[16] vdd gnd cell_6t
Xbit_r17_c203 bl[203] br[203] wl[17] vdd gnd cell_6t
Xbit_r18_c203 bl[203] br[203] wl[18] vdd gnd cell_6t
Xbit_r19_c203 bl[203] br[203] wl[19] vdd gnd cell_6t
Xbit_r20_c203 bl[203] br[203] wl[20] vdd gnd cell_6t
Xbit_r21_c203 bl[203] br[203] wl[21] vdd gnd cell_6t
Xbit_r22_c203 bl[203] br[203] wl[22] vdd gnd cell_6t
Xbit_r23_c203 bl[203] br[203] wl[23] vdd gnd cell_6t
Xbit_r24_c203 bl[203] br[203] wl[24] vdd gnd cell_6t
Xbit_r25_c203 bl[203] br[203] wl[25] vdd gnd cell_6t
Xbit_r26_c203 bl[203] br[203] wl[26] vdd gnd cell_6t
Xbit_r27_c203 bl[203] br[203] wl[27] vdd gnd cell_6t
Xbit_r28_c203 bl[203] br[203] wl[28] vdd gnd cell_6t
Xbit_r29_c203 bl[203] br[203] wl[29] vdd gnd cell_6t
Xbit_r30_c203 bl[203] br[203] wl[30] vdd gnd cell_6t
Xbit_r31_c203 bl[203] br[203] wl[31] vdd gnd cell_6t
Xbit_r32_c203 bl[203] br[203] wl[32] vdd gnd cell_6t
Xbit_r33_c203 bl[203] br[203] wl[33] vdd gnd cell_6t
Xbit_r34_c203 bl[203] br[203] wl[34] vdd gnd cell_6t
Xbit_r35_c203 bl[203] br[203] wl[35] vdd gnd cell_6t
Xbit_r36_c203 bl[203] br[203] wl[36] vdd gnd cell_6t
Xbit_r37_c203 bl[203] br[203] wl[37] vdd gnd cell_6t
Xbit_r38_c203 bl[203] br[203] wl[38] vdd gnd cell_6t
Xbit_r39_c203 bl[203] br[203] wl[39] vdd gnd cell_6t
Xbit_r40_c203 bl[203] br[203] wl[40] vdd gnd cell_6t
Xbit_r41_c203 bl[203] br[203] wl[41] vdd gnd cell_6t
Xbit_r42_c203 bl[203] br[203] wl[42] vdd gnd cell_6t
Xbit_r43_c203 bl[203] br[203] wl[43] vdd gnd cell_6t
Xbit_r44_c203 bl[203] br[203] wl[44] vdd gnd cell_6t
Xbit_r45_c203 bl[203] br[203] wl[45] vdd gnd cell_6t
Xbit_r46_c203 bl[203] br[203] wl[46] vdd gnd cell_6t
Xbit_r47_c203 bl[203] br[203] wl[47] vdd gnd cell_6t
Xbit_r48_c203 bl[203] br[203] wl[48] vdd gnd cell_6t
Xbit_r49_c203 bl[203] br[203] wl[49] vdd gnd cell_6t
Xbit_r50_c203 bl[203] br[203] wl[50] vdd gnd cell_6t
Xbit_r51_c203 bl[203] br[203] wl[51] vdd gnd cell_6t
Xbit_r52_c203 bl[203] br[203] wl[52] vdd gnd cell_6t
Xbit_r53_c203 bl[203] br[203] wl[53] vdd gnd cell_6t
Xbit_r54_c203 bl[203] br[203] wl[54] vdd gnd cell_6t
Xbit_r55_c203 bl[203] br[203] wl[55] vdd gnd cell_6t
Xbit_r56_c203 bl[203] br[203] wl[56] vdd gnd cell_6t
Xbit_r57_c203 bl[203] br[203] wl[57] vdd gnd cell_6t
Xbit_r58_c203 bl[203] br[203] wl[58] vdd gnd cell_6t
Xbit_r59_c203 bl[203] br[203] wl[59] vdd gnd cell_6t
Xbit_r60_c203 bl[203] br[203] wl[60] vdd gnd cell_6t
Xbit_r61_c203 bl[203] br[203] wl[61] vdd gnd cell_6t
Xbit_r62_c203 bl[203] br[203] wl[62] vdd gnd cell_6t
Xbit_r63_c203 bl[203] br[203] wl[63] vdd gnd cell_6t
Xbit_r64_c203 bl[203] br[203] wl[64] vdd gnd cell_6t
Xbit_r65_c203 bl[203] br[203] wl[65] vdd gnd cell_6t
Xbit_r66_c203 bl[203] br[203] wl[66] vdd gnd cell_6t
Xbit_r67_c203 bl[203] br[203] wl[67] vdd gnd cell_6t
Xbit_r68_c203 bl[203] br[203] wl[68] vdd gnd cell_6t
Xbit_r69_c203 bl[203] br[203] wl[69] vdd gnd cell_6t
Xbit_r70_c203 bl[203] br[203] wl[70] vdd gnd cell_6t
Xbit_r71_c203 bl[203] br[203] wl[71] vdd gnd cell_6t
Xbit_r72_c203 bl[203] br[203] wl[72] vdd gnd cell_6t
Xbit_r73_c203 bl[203] br[203] wl[73] vdd gnd cell_6t
Xbit_r74_c203 bl[203] br[203] wl[74] vdd gnd cell_6t
Xbit_r75_c203 bl[203] br[203] wl[75] vdd gnd cell_6t
Xbit_r76_c203 bl[203] br[203] wl[76] vdd gnd cell_6t
Xbit_r77_c203 bl[203] br[203] wl[77] vdd gnd cell_6t
Xbit_r78_c203 bl[203] br[203] wl[78] vdd gnd cell_6t
Xbit_r79_c203 bl[203] br[203] wl[79] vdd gnd cell_6t
Xbit_r80_c203 bl[203] br[203] wl[80] vdd gnd cell_6t
Xbit_r81_c203 bl[203] br[203] wl[81] vdd gnd cell_6t
Xbit_r82_c203 bl[203] br[203] wl[82] vdd gnd cell_6t
Xbit_r83_c203 bl[203] br[203] wl[83] vdd gnd cell_6t
Xbit_r84_c203 bl[203] br[203] wl[84] vdd gnd cell_6t
Xbit_r85_c203 bl[203] br[203] wl[85] vdd gnd cell_6t
Xbit_r86_c203 bl[203] br[203] wl[86] vdd gnd cell_6t
Xbit_r87_c203 bl[203] br[203] wl[87] vdd gnd cell_6t
Xbit_r88_c203 bl[203] br[203] wl[88] vdd gnd cell_6t
Xbit_r89_c203 bl[203] br[203] wl[89] vdd gnd cell_6t
Xbit_r90_c203 bl[203] br[203] wl[90] vdd gnd cell_6t
Xbit_r91_c203 bl[203] br[203] wl[91] vdd gnd cell_6t
Xbit_r92_c203 bl[203] br[203] wl[92] vdd gnd cell_6t
Xbit_r93_c203 bl[203] br[203] wl[93] vdd gnd cell_6t
Xbit_r94_c203 bl[203] br[203] wl[94] vdd gnd cell_6t
Xbit_r95_c203 bl[203] br[203] wl[95] vdd gnd cell_6t
Xbit_r96_c203 bl[203] br[203] wl[96] vdd gnd cell_6t
Xbit_r97_c203 bl[203] br[203] wl[97] vdd gnd cell_6t
Xbit_r98_c203 bl[203] br[203] wl[98] vdd gnd cell_6t
Xbit_r99_c203 bl[203] br[203] wl[99] vdd gnd cell_6t
Xbit_r100_c203 bl[203] br[203] wl[100] vdd gnd cell_6t
Xbit_r101_c203 bl[203] br[203] wl[101] vdd gnd cell_6t
Xbit_r102_c203 bl[203] br[203] wl[102] vdd gnd cell_6t
Xbit_r103_c203 bl[203] br[203] wl[103] vdd gnd cell_6t
Xbit_r104_c203 bl[203] br[203] wl[104] vdd gnd cell_6t
Xbit_r105_c203 bl[203] br[203] wl[105] vdd gnd cell_6t
Xbit_r106_c203 bl[203] br[203] wl[106] vdd gnd cell_6t
Xbit_r107_c203 bl[203] br[203] wl[107] vdd gnd cell_6t
Xbit_r108_c203 bl[203] br[203] wl[108] vdd gnd cell_6t
Xbit_r109_c203 bl[203] br[203] wl[109] vdd gnd cell_6t
Xbit_r110_c203 bl[203] br[203] wl[110] vdd gnd cell_6t
Xbit_r111_c203 bl[203] br[203] wl[111] vdd gnd cell_6t
Xbit_r112_c203 bl[203] br[203] wl[112] vdd gnd cell_6t
Xbit_r113_c203 bl[203] br[203] wl[113] vdd gnd cell_6t
Xbit_r114_c203 bl[203] br[203] wl[114] vdd gnd cell_6t
Xbit_r115_c203 bl[203] br[203] wl[115] vdd gnd cell_6t
Xbit_r116_c203 bl[203] br[203] wl[116] vdd gnd cell_6t
Xbit_r117_c203 bl[203] br[203] wl[117] vdd gnd cell_6t
Xbit_r118_c203 bl[203] br[203] wl[118] vdd gnd cell_6t
Xbit_r119_c203 bl[203] br[203] wl[119] vdd gnd cell_6t
Xbit_r120_c203 bl[203] br[203] wl[120] vdd gnd cell_6t
Xbit_r121_c203 bl[203] br[203] wl[121] vdd gnd cell_6t
Xbit_r122_c203 bl[203] br[203] wl[122] vdd gnd cell_6t
Xbit_r123_c203 bl[203] br[203] wl[123] vdd gnd cell_6t
Xbit_r124_c203 bl[203] br[203] wl[124] vdd gnd cell_6t
Xbit_r125_c203 bl[203] br[203] wl[125] vdd gnd cell_6t
Xbit_r126_c203 bl[203] br[203] wl[126] vdd gnd cell_6t
Xbit_r127_c203 bl[203] br[203] wl[127] vdd gnd cell_6t
Xbit_r128_c203 bl[203] br[203] wl[128] vdd gnd cell_6t
Xbit_r129_c203 bl[203] br[203] wl[129] vdd gnd cell_6t
Xbit_r130_c203 bl[203] br[203] wl[130] vdd gnd cell_6t
Xbit_r131_c203 bl[203] br[203] wl[131] vdd gnd cell_6t
Xbit_r132_c203 bl[203] br[203] wl[132] vdd gnd cell_6t
Xbit_r133_c203 bl[203] br[203] wl[133] vdd gnd cell_6t
Xbit_r134_c203 bl[203] br[203] wl[134] vdd gnd cell_6t
Xbit_r135_c203 bl[203] br[203] wl[135] vdd gnd cell_6t
Xbit_r136_c203 bl[203] br[203] wl[136] vdd gnd cell_6t
Xbit_r137_c203 bl[203] br[203] wl[137] vdd gnd cell_6t
Xbit_r138_c203 bl[203] br[203] wl[138] vdd gnd cell_6t
Xbit_r139_c203 bl[203] br[203] wl[139] vdd gnd cell_6t
Xbit_r140_c203 bl[203] br[203] wl[140] vdd gnd cell_6t
Xbit_r141_c203 bl[203] br[203] wl[141] vdd gnd cell_6t
Xbit_r142_c203 bl[203] br[203] wl[142] vdd gnd cell_6t
Xbit_r143_c203 bl[203] br[203] wl[143] vdd gnd cell_6t
Xbit_r144_c203 bl[203] br[203] wl[144] vdd gnd cell_6t
Xbit_r145_c203 bl[203] br[203] wl[145] vdd gnd cell_6t
Xbit_r146_c203 bl[203] br[203] wl[146] vdd gnd cell_6t
Xbit_r147_c203 bl[203] br[203] wl[147] vdd gnd cell_6t
Xbit_r148_c203 bl[203] br[203] wl[148] vdd gnd cell_6t
Xbit_r149_c203 bl[203] br[203] wl[149] vdd gnd cell_6t
Xbit_r150_c203 bl[203] br[203] wl[150] vdd gnd cell_6t
Xbit_r151_c203 bl[203] br[203] wl[151] vdd gnd cell_6t
Xbit_r152_c203 bl[203] br[203] wl[152] vdd gnd cell_6t
Xbit_r153_c203 bl[203] br[203] wl[153] vdd gnd cell_6t
Xbit_r154_c203 bl[203] br[203] wl[154] vdd gnd cell_6t
Xbit_r155_c203 bl[203] br[203] wl[155] vdd gnd cell_6t
Xbit_r156_c203 bl[203] br[203] wl[156] vdd gnd cell_6t
Xbit_r157_c203 bl[203] br[203] wl[157] vdd gnd cell_6t
Xbit_r158_c203 bl[203] br[203] wl[158] vdd gnd cell_6t
Xbit_r159_c203 bl[203] br[203] wl[159] vdd gnd cell_6t
Xbit_r160_c203 bl[203] br[203] wl[160] vdd gnd cell_6t
Xbit_r161_c203 bl[203] br[203] wl[161] vdd gnd cell_6t
Xbit_r162_c203 bl[203] br[203] wl[162] vdd gnd cell_6t
Xbit_r163_c203 bl[203] br[203] wl[163] vdd gnd cell_6t
Xbit_r164_c203 bl[203] br[203] wl[164] vdd gnd cell_6t
Xbit_r165_c203 bl[203] br[203] wl[165] vdd gnd cell_6t
Xbit_r166_c203 bl[203] br[203] wl[166] vdd gnd cell_6t
Xbit_r167_c203 bl[203] br[203] wl[167] vdd gnd cell_6t
Xbit_r168_c203 bl[203] br[203] wl[168] vdd gnd cell_6t
Xbit_r169_c203 bl[203] br[203] wl[169] vdd gnd cell_6t
Xbit_r170_c203 bl[203] br[203] wl[170] vdd gnd cell_6t
Xbit_r171_c203 bl[203] br[203] wl[171] vdd gnd cell_6t
Xbit_r172_c203 bl[203] br[203] wl[172] vdd gnd cell_6t
Xbit_r173_c203 bl[203] br[203] wl[173] vdd gnd cell_6t
Xbit_r174_c203 bl[203] br[203] wl[174] vdd gnd cell_6t
Xbit_r175_c203 bl[203] br[203] wl[175] vdd gnd cell_6t
Xbit_r176_c203 bl[203] br[203] wl[176] vdd gnd cell_6t
Xbit_r177_c203 bl[203] br[203] wl[177] vdd gnd cell_6t
Xbit_r178_c203 bl[203] br[203] wl[178] vdd gnd cell_6t
Xbit_r179_c203 bl[203] br[203] wl[179] vdd gnd cell_6t
Xbit_r180_c203 bl[203] br[203] wl[180] vdd gnd cell_6t
Xbit_r181_c203 bl[203] br[203] wl[181] vdd gnd cell_6t
Xbit_r182_c203 bl[203] br[203] wl[182] vdd gnd cell_6t
Xbit_r183_c203 bl[203] br[203] wl[183] vdd gnd cell_6t
Xbit_r184_c203 bl[203] br[203] wl[184] vdd gnd cell_6t
Xbit_r185_c203 bl[203] br[203] wl[185] vdd gnd cell_6t
Xbit_r186_c203 bl[203] br[203] wl[186] vdd gnd cell_6t
Xbit_r187_c203 bl[203] br[203] wl[187] vdd gnd cell_6t
Xbit_r188_c203 bl[203] br[203] wl[188] vdd gnd cell_6t
Xbit_r189_c203 bl[203] br[203] wl[189] vdd gnd cell_6t
Xbit_r190_c203 bl[203] br[203] wl[190] vdd gnd cell_6t
Xbit_r191_c203 bl[203] br[203] wl[191] vdd gnd cell_6t
Xbit_r192_c203 bl[203] br[203] wl[192] vdd gnd cell_6t
Xbit_r193_c203 bl[203] br[203] wl[193] vdd gnd cell_6t
Xbit_r194_c203 bl[203] br[203] wl[194] vdd gnd cell_6t
Xbit_r195_c203 bl[203] br[203] wl[195] vdd gnd cell_6t
Xbit_r196_c203 bl[203] br[203] wl[196] vdd gnd cell_6t
Xbit_r197_c203 bl[203] br[203] wl[197] vdd gnd cell_6t
Xbit_r198_c203 bl[203] br[203] wl[198] vdd gnd cell_6t
Xbit_r199_c203 bl[203] br[203] wl[199] vdd gnd cell_6t
Xbit_r200_c203 bl[203] br[203] wl[200] vdd gnd cell_6t
Xbit_r201_c203 bl[203] br[203] wl[201] vdd gnd cell_6t
Xbit_r202_c203 bl[203] br[203] wl[202] vdd gnd cell_6t
Xbit_r203_c203 bl[203] br[203] wl[203] vdd gnd cell_6t
Xbit_r204_c203 bl[203] br[203] wl[204] vdd gnd cell_6t
Xbit_r205_c203 bl[203] br[203] wl[205] vdd gnd cell_6t
Xbit_r206_c203 bl[203] br[203] wl[206] vdd gnd cell_6t
Xbit_r207_c203 bl[203] br[203] wl[207] vdd gnd cell_6t
Xbit_r208_c203 bl[203] br[203] wl[208] vdd gnd cell_6t
Xbit_r209_c203 bl[203] br[203] wl[209] vdd gnd cell_6t
Xbit_r210_c203 bl[203] br[203] wl[210] vdd gnd cell_6t
Xbit_r211_c203 bl[203] br[203] wl[211] vdd gnd cell_6t
Xbit_r212_c203 bl[203] br[203] wl[212] vdd gnd cell_6t
Xbit_r213_c203 bl[203] br[203] wl[213] vdd gnd cell_6t
Xbit_r214_c203 bl[203] br[203] wl[214] vdd gnd cell_6t
Xbit_r215_c203 bl[203] br[203] wl[215] vdd gnd cell_6t
Xbit_r216_c203 bl[203] br[203] wl[216] vdd gnd cell_6t
Xbit_r217_c203 bl[203] br[203] wl[217] vdd gnd cell_6t
Xbit_r218_c203 bl[203] br[203] wl[218] vdd gnd cell_6t
Xbit_r219_c203 bl[203] br[203] wl[219] vdd gnd cell_6t
Xbit_r220_c203 bl[203] br[203] wl[220] vdd gnd cell_6t
Xbit_r221_c203 bl[203] br[203] wl[221] vdd gnd cell_6t
Xbit_r222_c203 bl[203] br[203] wl[222] vdd gnd cell_6t
Xbit_r223_c203 bl[203] br[203] wl[223] vdd gnd cell_6t
Xbit_r224_c203 bl[203] br[203] wl[224] vdd gnd cell_6t
Xbit_r225_c203 bl[203] br[203] wl[225] vdd gnd cell_6t
Xbit_r226_c203 bl[203] br[203] wl[226] vdd gnd cell_6t
Xbit_r227_c203 bl[203] br[203] wl[227] vdd gnd cell_6t
Xbit_r228_c203 bl[203] br[203] wl[228] vdd gnd cell_6t
Xbit_r229_c203 bl[203] br[203] wl[229] vdd gnd cell_6t
Xbit_r230_c203 bl[203] br[203] wl[230] vdd gnd cell_6t
Xbit_r231_c203 bl[203] br[203] wl[231] vdd gnd cell_6t
Xbit_r232_c203 bl[203] br[203] wl[232] vdd gnd cell_6t
Xbit_r233_c203 bl[203] br[203] wl[233] vdd gnd cell_6t
Xbit_r234_c203 bl[203] br[203] wl[234] vdd gnd cell_6t
Xbit_r235_c203 bl[203] br[203] wl[235] vdd gnd cell_6t
Xbit_r236_c203 bl[203] br[203] wl[236] vdd gnd cell_6t
Xbit_r237_c203 bl[203] br[203] wl[237] vdd gnd cell_6t
Xbit_r238_c203 bl[203] br[203] wl[238] vdd gnd cell_6t
Xbit_r239_c203 bl[203] br[203] wl[239] vdd gnd cell_6t
Xbit_r240_c203 bl[203] br[203] wl[240] vdd gnd cell_6t
Xbit_r241_c203 bl[203] br[203] wl[241] vdd gnd cell_6t
Xbit_r242_c203 bl[203] br[203] wl[242] vdd gnd cell_6t
Xbit_r243_c203 bl[203] br[203] wl[243] vdd gnd cell_6t
Xbit_r244_c203 bl[203] br[203] wl[244] vdd gnd cell_6t
Xbit_r245_c203 bl[203] br[203] wl[245] vdd gnd cell_6t
Xbit_r246_c203 bl[203] br[203] wl[246] vdd gnd cell_6t
Xbit_r247_c203 bl[203] br[203] wl[247] vdd gnd cell_6t
Xbit_r248_c203 bl[203] br[203] wl[248] vdd gnd cell_6t
Xbit_r249_c203 bl[203] br[203] wl[249] vdd gnd cell_6t
Xbit_r250_c203 bl[203] br[203] wl[250] vdd gnd cell_6t
Xbit_r251_c203 bl[203] br[203] wl[251] vdd gnd cell_6t
Xbit_r252_c203 bl[203] br[203] wl[252] vdd gnd cell_6t
Xbit_r253_c203 bl[203] br[203] wl[253] vdd gnd cell_6t
Xbit_r254_c203 bl[203] br[203] wl[254] vdd gnd cell_6t
Xbit_r255_c203 bl[203] br[203] wl[255] vdd gnd cell_6t
Xbit_r0_c204 bl[204] br[204] wl[0] vdd gnd cell_6t
Xbit_r1_c204 bl[204] br[204] wl[1] vdd gnd cell_6t
Xbit_r2_c204 bl[204] br[204] wl[2] vdd gnd cell_6t
Xbit_r3_c204 bl[204] br[204] wl[3] vdd gnd cell_6t
Xbit_r4_c204 bl[204] br[204] wl[4] vdd gnd cell_6t
Xbit_r5_c204 bl[204] br[204] wl[5] vdd gnd cell_6t
Xbit_r6_c204 bl[204] br[204] wl[6] vdd gnd cell_6t
Xbit_r7_c204 bl[204] br[204] wl[7] vdd gnd cell_6t
Xbit_r8_c204 bl[204] br[204] wl[8] vdd gnd cell_6t
Xbit_r9_c204 bl[204] br[204] wl[9] vdd gnd cell_6t
Xbit_r10_c204 bl[204] br[204] wl[10] vdd gnd cell_6t
Xbit_r11_c204 bl[204] br[204] wl[11] vdd gnd cell_6t
Xbit_r12_c204 bl[204] br[204] wl[12] vdd gnd cell_6t
Xbit_r13_c204 bl[204] br[204] wl[13] vdd gnd cell_6t
Xbit_r14_c204 bl[204] br[204] wl[14] vdd gnd cell_6t
Xbit_r15_c204 bl[204] br[204] wl[15] vdd gnd cell_6t
Xbit_r16_c204 bl[204] br[204] wl[16] vdd gnd cell_6t
Xbit_r17_c204 bl[204] br[204] wl[17] vdd gnd cell_6t
Xbit_r18_c204 bl[204] br[204] wl[18] vdd gnd cell_6t
Xbit_r19_c204 bl[204] br[204] wl[19] vdd gnd cell_6t
Xbit_r20_c204 bl[204] br[204] wl[20] vdd gnd cell_6t
Xbit_r21_c204 bl[204] br[204] wl[21] vdd gnd cell_6t
Xbit_r22_c204 bl[204] br[204] wl[22] vdd gnd cell_6t
Xbit_r23_c204 bl[204] br[204] wl[23] vdd gnd cell_6t
Xbit_r24_c204 bl[204] br[204] wl[24] vdd gnd cell_6t
Xbit_r25_c204 bl[204] br[204] wl[25] vdd gnd cell_6t
Xbit_r26_c204 bl[204] br[204] wl[26] vdd gnd cell_6t
Xbit_r27_c204 bl[204] br[204] wl[27] vdd gnd cell_6t
Xbit_r28_c204 bl[204] br[204] wl[28] vdd gnd cell_6t
Xbit_r29_c204 bl[204] br[204] wl[29] vdd gnd cell_6t
Xbit_r30_c204 bl[204] br[204] wl[30] vdd gnd cell_6t
Xbit_r31_c204 bl[204] br[204] wl[31] vdd gnd cell_6t
Xbit_r32_c204 bl[204] br[204] wl[32] vdd gnd cell_6t
Xbit_r33_c204 bl[204] br[204] wl[33] vdd gnd cell_6t
Xbit_r34_c204 bl[204] br[204] wl[34] vdd gnd cell_6t
Xbit_r35_c204 bl[204] br[204] wl[35] vdd gnd cell_6t
Xbit_r36_c204 bl[204] br[204] wl[36] vdd gnd cell_6t
Xbit_r37_c204 bl[204] br[204] wl[37] vdd gnd cell_6t
Xbit_r38_c204 bl[204] br[204] wl[38] vdd gnd cell_6t
Xbit_r39_c204 bl[204] br[204] wl[39] vdd gnd cell_6t
Xbit_r40_c204 bl[204] br[204] wl[40] vdd gnd cell_6t
Xbit_r41_c204 bl[204] br[204] wl[41] vdd gnd cell_6t
Xbit_r42_c204 bl[204] br[204] wl[42] vdd gnd cell_6t
Xbit_r43_c204 bl[204] br[204] wl[43] vdd gnd cell_6t
Xbit_r44_c204 bl[204] br[204] wl[44] vdd gnd cell_6t
Xbit_r45_c204 bl[204] br[204] wl[45] vdd gnd cell_6t
Xbit_r46_c204 bl[204] br[204] wl[46] vdd gnd cell_6t
Xbit_r47_c204 bl[204] br[204] wl[47] vdd gnd cell_6t
Xbit_r48_c204 bl[204] br[204] wl[48] vdd gnd cell_6t
Xbit_r49_c204 bl[204] br[204] wl[49] vdd gnd cell_6t
Xbit_r50_c204 bl[204] br[204] wl[50] vdd gnd cell_6t
Xbit_r51_c204 bl[204] br[204] wl[51] vdd gnd cell_6t
Xbit_r52_c204 bl[204] br[204] wl[52] vdd gnd cell_6t
Xbit_r53_c204 bl[204] br[204] wl[53] vdd gnd cell_6t
Xbit_r54_c204 bl[204] br[204] wl[54] vdd gnd cell_6t
Xbit_r55_c204 bl[204] br[204] wl[55] vdd gnd cell_6t
Xbit_r56_c204 bl[204] br[204] wl[56] vdd gnd cell_6t
Xbit_r57_c204 bl[204] br[204] wl[57] vdd gnd cell_6t
Xbit_r58_c204 bl[204] br[204] wl[58] vdd gnd cell_6t
Xbit_r59_c204 bl[204] br[204] wl[59] vdd gnd cell_6t
Xbit_r60_c204 bl[204] br[204] wl[60] vdd gnd cell_6t
Xbit_r61_c204 bl[204] br[204] wl[61] vdd gnd cell_6t
Xbit_r62_c204 bl[204] br[204] wl[62] vdd gnd cell_6t
Xbit_r63_c204 bl[204] br[204] wl[63] vdd gnd cell_6t
Xbit_r64_c204 bl[204] br[204] wl[64] vdd gnd cell_6t
Xbit_r65_c204 bl[204] br[204] wl[65] vdd gnd cell_6t
Xbit_r66_c204 bl[204] br[204] wl[66] vdd gnd cell_6t
Xbit_r67_c204 bl[204] br[204] wl[67] vdd gnd cell_6t
Xbit_r68_c204 bl[204] br[204] wl[68] vdd gnd cell_6t
Xbit_r69_c204 bl[204] br[204] wl[69] vdd gnd cell_6t
Xbit_r70_c204 bl[204] br[204] wl[70] vdd gnd cell_6t
Xbit_r71_c204 bl[204] br[204] wl[71] vdd gnd cell_6t
Xbit_r72_c204 bl[204] br[204] wl[72] vdd gnd cell_6t
Xbit_r73_c204 bl[204] br[204] wl[73] vdd gnd cell_6t
Xbit_r74_c204 bl[204] br[204] wl[74] vdd gnd cell_6t
Xbit_r75_c204 bl[204] br[204] wl[75] vdd gnd cell_6t
Xbit_r76_c204 bl[204] br[204] wl[76] vdd gnd cell_6t
Xbit_r77_c204 bl[204] br[204] wl[77] vdd gnd cell_6t
Xbit_r78_c204 bl[204] br[204] wl[78] vdd gnd cell_6t
Xbit_r79_c204 bl[204] br[204] wl[79] vdd gnd cell_6t
Xbit_r80_c204 bl[204] br[204] wl[80] vdd gnd cell_6t
Xbit_r81_c204 bl[204] br[204] wl[81] vdd gnd cell_6t
Xbit_r82_c204 bl[204] br[204] wl[82] vdd gnd cell_6t
Xbit_r83_c204 bl[204] br[204] wl[83] vdd gnd cell_6t
Xbit_r84_c204 bl[204] br[204] wl[84] vdd gnd cell_6t
Xbit_r85_c204 bl[204] br[204] wl[85] vdd gnd cell_6t
Xbit_r86_c204 bl[204] br[204] wl[86] vdd gnd cell_6t
Xbit_r87_c204 bl[204] br[204] wl[87] vdd gnd cell_6t
Xbit_r88_c204 bl[204] br[204] wl[88] vdd gnd cell_6t
Xbit_r89_c204 bl[204] br[204] wl[89] vdd gnd cell_6t
Xbit_r90_c204 bl[204] br[204] wl[90] vdd gnd cell_6t
Xbit_r91_c204 bl[204] br[204] wl[91] vdd gnd cell_6t
Xbit_r92_c204 bl[204] br[204] wl[92] vdd gnd cell_6t
Xbit_r93_c204 bl[204] br[204] wl[93] vdd gnd cell_6t
Xbit_r94_c204 bl[204] br[204] wl[94] vdd gnd cell_6t
Xbit_r95_c204 bl[204] br[204] wl[95] vdd gnd cell_6t
Xbit_r96_c204 bl[204] br[204] wl[96] vdd gnd cell_6t
Xbit_r97_c204 bl[204] br[204] wl[97] vdd gnd cell_6t
Xbit_r98_c204 bl[204] br[204] wl[98] vdd gnd cell_6t
Xbit_r99_c204 bl[204] br[204] wl[99] vdd gnd cell_6t
Xbit_r100_c204 bl[204] br[204] wl[100] vdd gnd cell_6t
Xbit_r101_c204 bl[204] br[204] wl[101] vdd gnd cell_6t
Xbit_r102_c204 bl[204] br[204] wl[102] vdd gnd cell_6t
Xbit_r103_c204 bl[204] br[204] wl[103] vdd gnd cell_6t
Xbit_r104_c204 bl[204] br[204] wl[104] vdd gnd cell_6t
Xbit_r105_c204 bl[204] br[204] wl[105] vdd gnd cell_6t
Xbit_r106_c204 bl[204] br[204] wl[106] vdd gnd cell_6t
Xbit_r107_c204 bl[204] br[204] wl[107] vdd gnd cell_6t
Xbit_r108_c204 bl[204] br[204] wl[108] vdd gnd cell_6t
Xbit_r109_c204 bl[204] br[204] wl[109] vdd gnd cell_6t
Xbit_r110_c204 bl[204] br[204] wl[110] vdd gnd cell_6t
Xbit_r111_c204 bl[204] br[204] wl[111] vdd gnd cell_6t
Xbit_r112_c204 bl[204] br[204] wl[112] vdd gnd cell_6t
Xbit_r113_c204 bl[204] br[204] wl[113] vdd gnd cell_6t
Xbit_r114_c204 bl[204] br[204] wl[114] vdd gnd cell_6t
Xbit_r115_c204 bl[204] br[204] wl[115] vdd gnd cell_6t
Xbit_r116_c204 bl[204] br[204] wl[116] vdd gnd cell_6t
Xbit_r117_c204 bl[204] br[204] wl[117] vdd gnd cell_6t
Xbit_r118_c204 bl[204] br[204] wl[118] vdd gnd cell_6t
Xbit_r119_c204 bl[204] br[204] wl[119] vdd gnd cell_6t
Xbit_r120_c204 bl[204] br[204] wl[120] vdd gnd cell_6t
Xbit_r121_c204 bl[204] br[204] wl[121] vdd gnd cell_6t
Xbit_r122_c204 bl[204] br[204] wl[122] vdd gnd cell_6t
Xbit_r123_c204 bl[204] br[204] wl[123] vdd gnd cell_6t
Xbit_r124_c204 bl[204] br[204] wl[124] vdd gnd cell_6t
Xbit_r125_c204 bl[204] br[204] wl[125] vdd gnd cell_6t
Xbit_r126_c204 bl[204] br[204] wl[126] vdd gnd cell_6t
Xbit_r127_c204 bl[204] br[204] wl[127] vdd gnd cell_6t
Xbit_r128_c204 bl[204] br[204] wl[128] vdd gnd cell_6t
Xbit_r129_c204 bl[204] br[204] wl[129] vdd gnd cell_6t
Xbit_r130_c204 bl[204] br[204] wl[130] vdd gnd cell_6t
Xbit_r131_c204 bl[204] br[204] wl[131] vdd gnd cell_6t
Xbit_r132_c204 bl[204] br[204] wl[132] vdd gnd cell_6t
Xbit_r133_c204 bl[204] br[204] wl[133] vdd gnd cell_6t
Xbit_r134_c204 bl[204] br[204] wl[134] vdd gnd cell_6t
Xbit_r135_c204 bl[204] br[204] wl[135] vdd gnd cell_6t
Xbit_r136_c204 bl[204] br[204] wl[136] vdd gnd cell_6t
Xbit_r137_c204 bl[204] br[204] wl[137] vdd gnd cell_6t
Xbit_r138_c204 bl[204] br[204] wl[138] vdd gnd cell_6t
Xbit_r139_c204 bl[204] br[204] wl[139] vdd gnd cell_6t
Xbit_r140_c204 bl[204] br[204] wl[140] vdd gnd cell_6t
Xbit_r141_c204 bl[204] br[204] wl[141] vdd gnd cell_6t
Xbit_r142_c204 bl[204] br[204] wl[142] vdd gnd cell_6t
Xbit_r143_c204 bl[204] br[204] wl[143] vdd gnd cell_6t
Xbit_r144_c204 bl[204] br[204] wl[144] vdd gnd cell_6t
Xbit_r145_c204 bl[204] br[204] wl[145] vdd gnd cell_6t
Xbit_r146_c204 bl[204] br[204] wl[146] vdd gnd cell_6t
Xbit_r147_c204 bl[204] br[204] wl[147] vdd gnd cell_6t
Xbit_r148_c204 bl[204] br[204] wl[148] vdd gnd cell_6t
Xbit_r149_c204 bl[204] br[204] wl[149] vdd gnd cell_6t
Xbit_r150_c204 bl[204] br[204] wl[150] vdd gnd cell_6t
Xbit_r151_c204 bl[204] br[204] wl[151] vdd gnd cell_6t
Xbit_r152_c204 bl[204] br[204] wl[152] vdd gnd cell_6t
Xbit_r153_c204 bl[204] br[204] wl[153] vdd gnd cell_6t
Xbit_r154_c204 bl[204] br[204] wl[154] vdd gnd cell_6t
Xbit_r155_c204 bl[204] br[204] wl[155] vdd gnd cell_6t
Xbit_r156_c204 bl[204] br[204] wl[156] vdd gnd cell_6t
Xbit_r157_c204 bl[204] br[204] wl[157] vdd gnd cell_6t
Xbit_r158_c204 bl[204] br[204] wl[158] vdd gnd cell_6t
Xbit_r159_c204 bl[204] br[204] wl[159] vdd gnd cell_6t
Xbit_r160_c204 bl[204] br[204] wl[160] vdd gnd cell_6t
Xbit_r161_c204 bl[204] br[204] wl[161] vdd gnd cell_6t
Xbit_r162_c204 bl[204] br[204] wl[162] vdd gnd cell_6t
Xbit_r163_c204 bl[204] br[204] wl[163] vdd gnd cell_6t
Xbit_r164_c204 bl[204] br[204] wl[164] vdd gnd cell_6t
Xbit_r165_c204 bl[204] br[204] wl[165] vdd gnd cell_6t
Xbit_r166_c204 bl[204] br[204] wl[166] vdd gnd cell_6t
Xbit_r167_c204 bl[204] br[204] wl[167] vdd gnd cell_6t
Xbit_r168_c204 bl[204] br[204] wl[168] vdd gnd cell_6t
Xbit_r169_c204 bl[204] br[204] wl[169] vdd gnd cell_6t
Xbit_r170_c204 bl[204] br[204] wl[170] vdd gnd cell_6t
Xbit_r171_c204 bl[204] br[204] wl[171] vdd gnd cell_6t
Xbit_r172_c204 bl[204] br[204] wl[172] vdd gnd cell_6t
Xbit_r173_c204 bl[204] br[204] wl[173] vdd gnd cell_6t
Xbit_r174_c204 bl[204] br[204] wl[174] vdd gnd cell_6t
Xbit_r175_c204 bl[204] br[204] wl[175] vdd gnd cell_6t
Xbit_r176_c204 bl[204] br[204] wl[176] vdd gnd cell_6t
Xbit_r177_c204 bl[204] br[204] wl[177] vdd gnd cell_6t
Xbit_r178_c204 bl[204] br[204] wl[178] vdd gnd cell_6t
Xbit_r179_c204 bl[204] br[204] wl[179] vdd gnd cell_6t
Xbit_r180_c204 bl[204] br[204] wl[180] vdd gnd cell_6t
Xbit_r181_c204 bl[204] br[204] wl[181] vdd gnd cell_6t
Xbit_r182_c204 bl[204] br[204] wl[182] vdd gnd cell_6t
Xbit_r183_c204 bl[204] br[204] wl[183] vdd gnd cell_6t
Xbit_r184_c204 bl[204] br[204] wl[184] vdd gnd cell_6t
Xbit_r185_c204 bl[204] br[204] wl[185] vdd gnd cell_6t
Xbit_r186_c204 bl[204] br[204] wl[186] vdd gnd cell_6t
Xbit_r187_c204 bl[204] br[204] wl[187] vdd gnd cell_6t
Xbit_r188_c204 bl[204] br[204] wl[188] vdd gnd cell_6t
Xbit_r189_c204 bl[204] br[204] wl[189] vdd gnd cell_6t
Xbit_r190_c204 bl[204] br[204] wl[190] vdd gnd cell_6t
Xbit_r191_c204 bl[204] br[204] wl[191] vdd gnd cell_6t
Xbit_r192_c204 bl[204] br[204] wl[192] vdd gnd cell_6t
Xbit_r193_c204 bl[204] br[204] wl[193] vdd gnd cell_6t
Xbit_r194_c204 bl[204] br[204] wl[194] vdd gnd cell_6t
Xbit_r195_c204 bl[204] br[204] wl[195] vdd gnd cell_6t
Xbit_r196_c204 bl[204] br[204] wl[196] vdd gnd cell_6t
Xbit_r197_c204 bl[204] br[204] wl[197] vdd gnd cell_6t
Xbit_r198_c204 bl[204] br[204] wl[198] vdd gnd cell_6t
Xbit_r199_c204 bl[204] br[204] wl[199] vdd gnd cell_6t
Xbit_r200_c204 bl[204] br[204] wl[200] vdd gnd cell_6t
Xbit_r201_c204 bl[204] br[204] wl[201] vdd gnd cell_6t
Xbit_r202_c204 bl[204] br[204] wl[202] vdd gnd cell_6t
Xbit_r203_c204 bl[204] br[204] wl[203] vdd gnd cell_6t
Xbit_r204_c204 bl[204] br[204] wl[204] vdd gnd cell_6t
Xbit_r205_c204 bl[204] br[204] wl[205] vdd gnd cell_6t
Xbit_r206_c204 bl[204] br[204] wl[206] vdd gnd cell_6t
Xbit_r207_c204 bl[204] br[204] wl[207] vdd gnd cell_6t
Xbit_r208_c204 bl[204] br[204] wl[208] vdd gnd cell_6t
Xbit_r209_c204 bl[204] br[204] wl[209] vdd gnd cell_6t
Xbit_r210_c204 bl[204] br[204] wl[210] vdd gnd cell_6t
Xbit_r211_c204 bl[204] br[204] wl[211] vdd gnd cell_6t
Xbit_r212_c204 bl[204] br[204] wl[212] vdd gnd cell_6t
Xbit_r213_c204 bl[204] br[204] wl[213] vdd gnd cell_6t
Xbit_r214_c204 bl[204] br[204] wl[214] vdd gnd cell_6t
Xbit_r215_c204 bl[204] br[204] wl[215] vdd gnd cell_6t
Xbit_r216_c204 bl[204] br[204] wl[216] vdd gnd cell_6t
Xbit_r217_c204 bl[204] br[204] wl[217] vdd gnd cell_6t
Xbit_r218_c204 bl[204] br[204] wl[218] vdd gnd cell_6t
Xbit_r219_c204 bl[204] br[204] wl[219] vdd gnd cell_6t
Xbit_r220_c204 bl[204] br[204] wl[220] vdd gnd cell_6t
Xbit_r221_c204 bl[204] br[204] wl[221] vdd gnd cell_6t
Xbit_r222_c204 bl[204] br[204] wl[222] vdd gnd cell_6t
Xbit_r223_c204 bl[204] br[204] wl[223] vdd gnd cell_6t
Xbit_r224_c204 bl[204] br[204] wl[224] vdd gnd cell_6t
Xbit_r225_c204 bl[204] br[204] wl[225] vdd gnd cell_6t
Xbit_r226_c204 bl[204] br[204] wl[226] vdd gnd cell_6t
Xbit_r227_c204 bl[204] br[204] wl[227] vdd gnd cell_6t
Xbit_r228_c204 bl[204] br[204] wl[228] vdd gnd cell_6t
Xbit_r229_c204 bl[204] br[204] wl[229] vdd gnd cell_6t
Xbit_r230_c204 bl[204] br[204] wl[230] vdd gnd cell_6t
Xbit_r231_c204 bl[204] br[204] wl[231] vdd gnd cell_6t
Xbit_r232_c204 bl[204] br[204] wl[232] vdd gnd cell_6t
Xbit_r233_c204 bl[204] br[204] wl[233] vdd gnd cell_6t
Xbit_r234_c204 bl[204] br[204] wl[234] vdd gnd cell_6t
Xbit_r235_c204 bl[204] br[204] wl[235] vdd gnd cell_6t
Xbit_r236_c204 bl[204] br[204] wl[236] vdd gnd cell_6t
Xbit_r237_c204 bl[204] br[204] wl[237] vdd gnd cell_6t
Xbit_r238_c204 bl[204] br[204] wl[238] vdd gnd cell_6t
Xbit_r239_c204 bl[204] br[204] wl[239] vdd gnd cell_6t
Xbit_r240_c204 bl[204] br[204] wl[240] vdd gnd cell_6t
Xbit_r241_c204 bl[204] br[204] wl[241] vdd gnd cell_6t
Xbit_r242_c204 bl[204] br[204] wl[242] vdd gnd cell_6t
Xbit_r243_c204 bl[204] br[204] wl[243] vdd gnd cell_6t
Xbit_r244_c204 bl[204] br[204] wl[244] vdd gnd cell_6t
Xbit_r245_c204 bl[204] br[204] wl[245] vdd gnd cell_6t
Xbit_r246_c204 bl[204] br[204] wl[246] vdd gnd cell_6t
Xbit_r247_c204 bl[204] br[204] wl[247] vdd gnd cell_6t
Xbit_r248_c204 bl[204] br[204] wl[248] vdd gnd cell_6t
Xbit_r249_c204 bl[204] br[204] wl[249] vdd gnd cell_6t
Xbit_r250_c204 bl[204] br[204] wl[250] vdd gnd cell_6t
Xbit_r251_c204 bl[204] br[204] wl[251] vdd gnd cell_6t
Xbit_r252_c204 bl[204] br[204] wl[252] vdd gnd cell_6t
Xbit_r253_c204 bl[204] br[204] wl[253] vdd gnd cell_6t
Xbit_r254_c204 bl[204] br[204] wl[254] vdd gnd cell_6t
Xbit_r255_c204 bl[204] br[204] wl[255] vdd gnd cell_6t
Xbit_r0_c205 bl[205] br[205] wl[0] vdd gnd cell_6t
Xbit_r1_c205 bl[205] br[205] wl[1] vdd gnd cell_6t
Xbit_r2_c205 bl[205] br[205] wl[2] vdd gnd cell_6t
Xbit_r3_c205 bl[205] br[205] wl[3] vdd gnd cell_6t
Xbit_r4_c205 bl[205] br[205] wl[4] vdd gnd cell_6t
Xbit_r5_c205 bl[205] br[205] wl[5] vdd gnd cell_6t
Xbit_r6_c205 bl[205] br[205] wl[6] vdd gnd cell_6t
Xbit_r7_c205 bl[205] br[205] wl[7] vdd gnd cell_6t
Xbit_r8_c205 bl[205] br[205] wl[8] vdd gnd cell_6t
Xbit_r9_c205 bl[205] br[205] wl[9] vdd gnd cell_6t
Xbit_r10_c205 bl[205] br[205] wl[10] vdd gnd cell_6t
Xbit_r11_c205 bl[205] br[205] wl[11] vdd gnd cell_6t
Xbit_r12_c205 bl[205] br[205] wl[12] vdd gnd cell_6t
Xbit_r13_c205 bl[205] br[205] wl[13] vdd gnd cell_6t
Xbit_r14_c205 bl[205] br[205] wl[14] vdd gnd cell_6t
Xbit_r15_c205 bl[205] br[205] wl[15] vdd gnd cell_6t
Xbit_r16_c205 bl[205] br[205] wl[16] vdd gnd cell_6t
Xbit_r17_c205 bl[205] br[205] wl[17] vdd gnd cell_6t
Xbit_r18_c205 bl[205] br[205] wl[18] vdd gnd cell_6t
Xbit_r19_c205 bl[205] br[205] wl[19] vdd gnd cell_6t
Xbit_r20_c205 bl[205] br[205] wl[20] vdd gnd cell_6t
Xbit_r21_c205 bl[205] br[205] wl[21] vdd gnd cell_6t
Xbit_r22_c205 bl[205] br[205] wl[22] vdd gnd cell_6t
Xbit_r23_c205 bl[205] br[205] wl[23] vdd gnd cell_6t
Xbit_r24_c205 bl[205] br[205] wl[24] vdd gnd cell_6t
Xbit_r25_c205 bl[205] br[205] wl[25] vdd gnd cell_6t
Xbit_r26_c205 bl[205] br[205] wl[26] vdd gnd cell_6t
Xbit_r27_c205 bl[205] br[205] wl[27] vdd gnd cell_6t
Xbit_r28_c205 bl[205] br[205] wl[28] vdd gnd cell_6t
Xbit_r29_c205 bl[205] br[205] wl[29] vdd gnd cell_6t
Xbit_r30_c205 bl[205] br[205] wl[30] vdd gnd cell_6t
Xbit_r31_c205 bl[205] br[205] wl[31] vdd gnd cell_6t
Xbit_r32_c205 bl[205] br[205] wl[32] vdd gnd cell_6t
Xbit_r33_c205 bl[205] br[205] wl[33] vdd gnd cell_6t
Xbit_r34_c205 bl[205] br[205] wl[34] vdd gnd cell_6t
Xbit_r35_c205 bl[205] br[205] wl[35] vdd gnd cell_6t
Xbit_r36_c205 bl[205] br[205] wl[36] vdd gnd cell_6t
Xbit_r37_c205 bl[205] br[205] wl[37] vdd gnd cell_6t
Xbit_r38_c205 bl[205] br[205] wl[38] vdd gnd cell_6t
Xbit_r39_c205 bl[205] br[205] wl[39] vdd gnd cell_6t
Xbit_r40_c205 bl[205] br[205] wl[40] vdd gnd cell_6t
Xbit_r41_c205 bl[205] br[205] wl[41] vdd gnd cell_6t
Xbit_r42_c205 bl[205] br[205] wl[42] vdd gnd cell_6t
Xbit_r43_c205 bl[205] br[205] wl[43] vdd gnd cell_6t
Xbit_r44_c205 bl[205] br[205] wl[44] vdd gnd cell_6t
Xbit_r45_c205 bl[205] br[205] wl[45] vdd gnd cell_6t
Xbit_r46_c205 bl[205] br[205] wl[46] vdd gnd cell_6t
Xbit_r47_c205 bl[205] br[205] wl[47] vdd gnd cell_6t
Xbit_r48_c205 bl[205] br[205] wl[48] vdd gnd cell_6t
Xbit_r49_c205 bl[205] br[205] wl[49] vdd gnd cell_6t
Xbit_r50_c205 bl[205] br[205] wl[50] vdd gnd cell_6t
Xbit_r51_c205 bl[205] br[205] wl[51] vdd gnd cell_6t
Xbit_r52_c205 bl[205] br[205] wl[52] vdd gnd cell_6t
Xbit_r53_c205 bl[205] br[205] wl[53] vdd gnd cell_6t
Xbit_r54_c205 bl[205] br[205] wl[54] vdd gnd cell_6t
Xbit_r55_c205 bl[205] br[205] wl[55] vdd gnd cell_6t
Xbit_r56_c205 bl[205] br[205] wl[56] vdd gnd cell_6t
Xbit_r57_c205 bl[205] br[205] wl[57] vdd gnd cell_6t
Xbit_r58_c205 bl[205] br[205] wl[58] vdd gnd cell_6t
Xbit_r59_c205 bl[205] br[205] wl[59] vdd gnd cell_6t
Xbit_r60_c205 bl[205] br[205] wl[60] vdd gnd cell_6t
Xbit_r61_c205 bl[205] br[205] wl[61] vdd gnd cell_6t
Xbit_r62_c205 bl[205] br[205] wl[62] vdd gnd cell_6t
Xbit_r63_c205 bl[205] br[205] wl[63] vdd gnd cell_6t
Xbit_r64_c205 bl[205] br[205] wl[64] vdd gnd cell_6t
Xbit_r65_c205 bl[205] br[205] wl[65] vdd gnd cell_6t
Xbit_r66_c205 bl[205] br[205] wl[66] vdd gnd cell_6t
Xbit_r67_c205 bl[205] br[205] wl[67] vdd gnd cell_6t
Xbit_r68_c205 bl[205] br[205] wl[68] vdd gnd cell_6t
Xbit_r69_c205 bl[205] br[205] wl[69] vdd gnd cell_6t
Xbit_r70_c205 bl[205] br[205] wl[70] vdd gnd cell_6t
Xbit_r71_c205 bl[205] br[205] wl[71] vdd gnd cell_6t
Xbit_r72_c205 bl[205] br[205] wl[72] vdd gnd cell_6t
Xbit_r73_c205 bl[205] br[205] wl[73] vdd gnd cell_6t
Xbit_r74_c205 bl[205] br[205] wl[74] vdd gnd cell_6t
Xbit_r75_c205 bl[205] br[205] wl[75] vdd gnd cell_6t
Xbit_r76_c205 bl[205] br[205] wl[76] vdd gnd cell_6t
Xbit_r77_c205 bl[205] br[205] wl[77] vdd gnd cell_6t
Xbit_r78_c205 bl[205] br[205] wl[78] vdd gnd cell_6t
Xbit_r79_c205 bl[205] br[205] wl[79] vdd gnd cell_6t
Xbit_r80_c205 bl[205] br[205] wl[80] vdd gnd cell_6t
Xbit_r81_c205 bl[205] br[205] wl[81] vdd gnd cell_6t
Xbit_r82_c205 bl[205] br[205] wl[82] vdd gnd cell_6t
Xbit_r83_c205 bl[205] br[205] wl[83] vdd gnd cell_6t
Xbit_r84_c205 bl[205] br[205] wl[84] vdd gnd cell_6t
Xbit_r85_c205 bl[205] br[205] wl[85] vdd gnd cell_6t
Xbit_r86_c205 bl[205] br[205] wl[86] vdd gnd cell_6t
Xbit_r87_c205 bl[205] br[205] wl[87] vdd gnd cell_6t
Xbit_r88_c205 bl[205] br[205] wl[88] vdd gnd cell_6t
Xbit_r89_c205 bl[205] br[205] wl[89] vdd gnd cell_6t
Xbit_r90_c205 bl[205] br[205] wl[90] vdd gnd cell_6t
Xbit_r91_c205 bl[205] br[205] wl[91] vdd gnd cell_6t
Xbit_r92_c205 bl[205] br[205] wl[92] vdd gnd cell_6t
Xbit_r93_c205 bl[205] br[205] wl[93] vdd gnd cell_6t
Xbit_r94_c205 bl[205] br[205] wl[94] vdd gnd cell_6t
Xbit_r95_c205 bl[205] br[205] wl[95] vdd gnd cell_6t
Xbit_r96_c205 bl[205] br[205] wl[96] vdd gnd cell_6t
Xbit_r97_c205 bl[205] br[205] wl[97] vdd gnd cell_6t
Xbit_r98_c205 bl[205] br[205] wl[98] vdd gnd cell_6t
Xbit_r99_c205 bl[205] br[205] wl[99] vdd gnd cell_6t
Xbit_r100_c205 bl[205] br[205] wl[100] vdd gnd cell_6t
Xbit_r101_c205 bl[205] br[205] wl[101] vdd gnd cell_6t
Xbit_r102_c205 bl[205] br[205] wl[102] vdd gnd cell_6t
Xbit_r103_c205 bl[205] br[205] wl[103] vdd gnd cell_6t
Xbit_r104_c205 bl[205] br[205] wl[104] vdd gnd cell_6t
Xbit_r105_c205 bl[205] br[205] wl[105] vdd gnd cell_6t
Xbit_r106_c205 bl[205] br[205] wl[106] vdd gnd cell_6t
Xbit_r107_c205 bl[205] br[205] wl[107] vdd gnd cell_6t
Xbit_r108_c205 bl[205] br[205] wl[108] vdd gnd cell_6t
Xbit_r109_c205 bl[205] br[205] wl[109] vdd gnd cell_6t
Xbit_r110_c205 bl[205] br[205] wl[110] vdd gnd cell_6t
Xbit_r111_c205 bl[205] br[205] wl[111] vdd gnd cell_6t
Xbit_r112_c205 bl[205] br[205] wl[112] vdd gnd cell_6t
Xbit_r113_c205 bl[205] br[205] wl[113] vdd gnd cell_6t
Xbit_r114_c205 bl[205] br[205] wl[114] vdd gnd cell_6t
Xbit_r115_c205 bl[205] br[205] wl[115] vdd gnd cell_6t
Xbit_r116_c205 bl[205] br[205] wl[116] vdd gnd cell_6t
Xbit_r117_c205 bl[205] br[205] wl[117] vdd gnd cell_6t
Xbit_r118_c205 bl[205] br[205] wl[118] vdd gnd cell_6t
Xbit_r119_c205 bl[205] br[205] wl[119] vdd gnd cell_6t
Xbit_r120_c205 bl[205] br[205] wl[120] vdd gnd cell_6t
Xbit_r121_c205 bl[205] br[205] wl[121] vdd gnd cell_6t
Xbit_r122_c205 bl[205] br[205] wl[122] vdd gnd cell_6t
Xbit_r123_c205 bl[205] br[205] wl[123] vdd gnd cell_6t
Xbit_r124_c205 bl[205] br[205] wl[124] vdd gnd cell_6t
Xbit_r125_c205 bl[205] br[205] wl[125] vdd gnd cell_6t
Xbit_r126_c205 bl[205] br[205] wl[126] vdd gnd cell_6t
Xbit_r127_c205 bl[205] br[205] wl[127] vdd gnd cell_6t
Xbit_r128_c205 bl[205] br[205] wl[128] vdd gnd cell_6t
Xbit_r129_c205 bl[205] br[205] wl[129] vdd gnd cell_6t
Xbit_r130_c205 bl[205] br[205] wl[130] vdd gnd cell_6t
Xbit_r131_c205 bl[205] br[205] wl[131] vdd gnd cell_6t
Xbit_r132_c205 bl[205] br[205] wl[132] vdd gnd cell_6t
Xbit_r133_c205 bl[205] br[205] wl[133] vdd gnd cell_6t
Xbit_r134_c205 bl[205] br[205] wl[134] vdd gnd cell_6t
Xbit_r135_c205 bl[205] br[205] wl[135] vdd gnd cell_6t
Xbit_r136_c205 bl[205] br[205] wl[136] vdd gnd cell_6t
Xbit_r137_c205 bl[205] br[205] wl[137] vdd gnd cell_6t
Xbit_r138_c205 bl[205] br[205] wl[138] vdd gnd cell_6t
Xbit_r139_c205 bl[205] br[205] wl[139] vdd gnd cell_6t
Xbit_r140_c205 bl[205] br[205] wl[140] vdd gnd cell_6t
Xbit_r141_c205 bl[205] br[205] wl[141] vdd gnd cell_6t
Xbit_r142_c205 bl[205] br[205] wl[142] vdd gnd cell_6t
Xbit_r143_c205 bl[205] br[205] wl[143] vdd gnd cell_6t
Xbit_r144_c205 bl[205] br[205] wl[144] vdd gnd cell_6t
Xbit_r145_c205 bl[205] br[205] wl[145] vdd gnd cell_6t
Xbit_r146_c205 bl[205] br[205] wl[146] vdd gnd cell_6t
Xbit_r147_c205 bl[205] br[205] wl[147] vdd gnd cell_6t
Xbit_r148_c205 bl[205] br[205] wl[148] vdd gnd cell_6t
Xbit_r149_c205 bl[205] br[205] wl[149] vdd gnd cell_6t
Xbit_r150_c205 bl[205] br[205] wl[150] vdd gnd cell_6t
Xbit_r151_c205 bl[205] br[205] wl[151] vdd gnd cell_6t
Xbit_r152_c205 bl[205] br[205] wl[152] vdd gnd cell_6t
Xbit_r153_c205 bl[205] br[205] wl[153] vdd gnd cell_6t
Xbit_r154_c205 bl[205] br[205] wl[154] vdd gnd cell_6t
Xbit_r155_c205 bl[205] br[205] wl[155] vdd gnd cell_6t
Xbit_r156_c205 bl[205] br[205] wl[156] vdd gnd cell_6t
Xbit_r157_c205 bl[205] br[205] wl[157] vdd gnd cell_6t
Xbit_r158_c205 bl[205] br[205] wl[158] vdd gnd cell_6t
Xbit_r159_c205 bl[205] br[205] wl[159] vdd gnd cell_6t
Xbit_r160_c205 bl[205] br[205] wl[160] vdd gnd cell_6t
Xbit_r161_c205 bl[205] br[205] wl[161] vdd gnd cell_6t
Xbit_r162_c205 bl[205] br[205] wl[162] vdd gnd cell_6t
Xbit_r163_c205 bl[205] br[205] wl[163] vdd gnd cell_6t
Xbit_r164_c205 bl[205] br[205] wl[164] vdd gnd cell_6t
Xbit_r165_c205 bl[205] br[205] wl[165] vdd gnd cell_6t
Xbit_r166_c205 bl[205] br[205] wl[166] vdd gnd cell_6t
Xbit_r167_c205 bl[205] br[205] wl[167] vdd gnd cell_6t
Xbit_r168_c205 bl[205] br[205] wl[168] vdd gnd cell_6t
Xbit_r169_c205 bl[205] br[205] wl[169] vdd gnd cell_6t
Xbit_r170_c205 bl[205] br[205] wl[170] vdd gnd cell_6t
Xbit_r171_c205 bl[205] br[205] wl[171] vdd gnd cell_6t
Xbit_r172_c205 bl[205] br[205] wl[172] vdd gnd cell_6t
Xbit_r173_c205 bl[205] br[205] wl[173] vdd gnd cell_6t
Xbit_r174_c205 bl[205] br[205] wl[174] vdd gnd cell_6t
Xbit_r175_c205 bl[205] br[205] wl[175] vdd gnd cell_6t
Xbit_r176_c205 bl[205] br[205] wl[176] vdd gnd cell_6t
Xbit_r177_c205 bl[205] br[205] wl[177] vdd gnd cell_6t
Xbit_r178_c205 bl[205] br[205] wl[178] vdd gnd cell_6t
Xbit_r179_c205 bl[205] br[205] wl[179] vdd gnd cell_6t
Xbit_r180_c205 bl[205] br[205] wl[180] vdd gnd cell_6t
Xbit_r181_c205 bl[205] br[205] wl[181] vdd gnd cell_6t
Xbit_r182_c205 bl[205] br[205] wl[182] vdd gnd cell_6t
Xbit_r183_c205 bl[205] br[205] wl[183] vdd gnd cell_6t
Xbit_r184_c205 bl[205] br[205] wl[184] vdd gnd cell_6t
Xbit_r185_c205 bl[205] br[205] wl[185] vdd gnd cell_6t
Xbit_r186_c205 bl[205] br[205] wl[186] vdd gnd cell_6t
Xbit_r187_c205 bl[205] br[205] wl[187] vdd gnd cell_6t
Xbit_r188_c205 bl[205] br[205] wl[188] vdd gnd cell_6t
Xbit_r189_c205 bl[205] br[205] wl[189] vdd gnd cell_6t
Xbit_r190_c205 bl[205] br[205] wl[190] vdd gnd cell_6t
Xbit_r191_c205 bl[205] br[205] wl[191] vdd gnd cell_6t
Xbit_r192_c205 bl[205] br[205] wl[192] vdd gnd cell_6t
Xbit_r193_c205 bl[205] br[205] wl[193] vdd gnd cell_6t
Xbit_r194_c205 bl[205] br[205] wl[194] vdd gnd cell_6t
Xbit_r195_c205 bl[205] br[205] wl[195] vdd gnd cell_6t
Xbit_r196_c205 bl[205] br[205] wl[196] vdd gnd cell_6t
Xbit_r197_c205 bl[205] br[205] wl[197] vdd gnd cell_6t
Xbit_r198_c205 bl[205] br[205] wl[198] vdd gnd cell_6t
Xbit_r199_c205 bl[205] br[205] wl[199] vdd gnd cell_6t
Xbit_r200_c205 bl[205] br[205] wl[200] vdd gnd cell_6t
Xbit_r201_c205 bl[205] br[205] wl[201] vdd gnd cell_6t
Xbit_r202_c205 bl[205] br[205] wl[202] vdd gnd cell_6t
Xbit_r203_c205 bl[205] br[205] wl[203] vdd gnd cell_6t
Xbit_r204_c205 bl[205] br[205] wl[204] vdd gnd cell_6t
Xbit_r205_c205 bl[205] br[205] wl[205] vdd gnd cell_6t
Xbit_r206_c205 bl[205] br[205] wl[206] vdd gnd cell_6t
Xbit_r207_c205 bl[205] br[205] wl[207] vdd gnd cell_6t
Xbit_r208_c205 bl[205] br[205] wl[208] vdd gnd cell_6t
Xbit_r209_c205 bl[205] br[205] wl[209] vdd gnd cell_6t
Xbit_r210_c205 bl[205] br[205] wl[210] vdd gnd cell_6t
Xbit_r211_c205 bl[205] br[205] wl[211] vdd gnd cell_6t
Xbit_r212_c205 bl[205] br[205] wl[212] vdd gnd cell_6t
Xbit_r213_c205 bl[205] br[205] wl[213] vdd gnd cell_6t
Xbit_r214_c205 bl[205] br[205] wl[214] vdd gnd cell_6t
Xbit_r215_c205 bl[205] br[205] wl[215] vdd gnd cell_6t
Xbit_r216_c205 bl[205] br[205] wl[216] vdd gnd cell_6t
Xbit_r217_c205 bl[205] br[205] wl[217] vdd gnd cell_6t
Xbit_r218_c205 bl[205] br[205] wl[218] vdd gnd cell_6t
Xbit_r219_c205 bl[205] br[205] wl[219] vdd gnd cell_6t
Xbit_r220_c205 bl[205] br[205] wl[220] vdd gnd cell_6t
Xbit_r221_c205 bl[205] br[205] wl[221] vdd gnd cell_6t
Xbit_r222_c205 bl[205] br[205] wl[222] vdd gnd cell_6t
Xbit_r223_c205 bl[205] br[205] wl[223] vdd gnd cell_6t
Xbit_r224_c205 bl[205] br[205] wl[224] vdd gnd cell_6t
Xbit_r225_c205 bl[205] br[205] wl[225] vdd gnd cell_6t
Xbit_r226_c205 bl[205] br[205] wl[226] vdd gnd cell_6t
Xbit_r227_c205 bl[205] br[205] wl[227] vdd gnd cell_6t
Xbit_r228_c205 bl[205] br[205] wl[228] vdd gnd cell_6t
Xbit_r229_c205 bl[205] br[205] wl[229] vdd gnd cell_6t
Xbit_r230_c205 bl[205] br[205] wl[230] vdd gnd cell_6t
Xbit_r231_c205 bl[205] br[205] wl[231] vdd gnd cell_6t
Xbit_r232_c205 bl[205] br[205] wl[232] vdd gnd cell_6t
Xbit_r233_c205 bl[205] br[205] wl[233] vdd gnd cell_6t
Xbit_r234_c205 bl[205] br[205] wl[234] vdd gnd cell_6t
Xbit_r235_c205 bl[205] br[205] wl[235] vdd gnd cell_6t
Xbit_r236_c205 bl[205] br[205] wl[236] vdd gnd cell_6t
Xbit_r237_c205 bl[205] br[205] wl[237] vdd gnd cell_6t
Xbit_r238_c205 bl[205] br[205] wl[238] vdd gnd cell_6t
Xbit_r239_c205 bl[205] br[205] wl[239] vdd gnd cell_6t
Xbit_r240_c205 bl[205] br[205] wl[240] vdd gnd cell_6t
Xbit_r241_c205 bl[205] br[205] wl[241] vdd gnd cell_6t
Xbit_r242_c205 bl[205] br[205] wl[242] vdd gnd cell_6t
Xbit_r243_c205 bl[205] br[205] wl[243] vdd gnd cell_6t
Xbit_r244_c205 bl[205] br[205] wl[244] vdd gnd cell_6t
Xbit_r245_c205 bl[205] br[205] wl[245] vdd gnd cell_6t
Xbit_r246_c205 bl[205] br[205] wl[246] vdd gnd cell_6t
Xbit_r247_c205 bl[205] br[205] wl[247] vdd gnd cell_6t
Xbit_r248_c205 bl[205] br[205] wl[248] vdd gnd cell_6t
Xbit_r249_c205 bl[205] br[205] wl[249] vdd gnd cell_6t
Xbit_r250_c205 bl[205] br[205] wl[250] vdd gnd cell_6t
Xbit_r251_c205 bl[205] br[205] wl[251] vdd gnd cell_6t
Xbit_r252_c205 bl[205] br[205] wl[252] vdd gnd cell_6t
Xbit_r253_c205 bl[205] br[205] wl[253] vdd gnd cell_6t
Xbit_r254_c205 bl[205] br[205] wl[254] vdd gnd cell_6t
Xbit_r255_c205 bl[205] br[205] wl[255] vdd gnd cell_6t
Xbit_r0_c206 bl[206] br[206] wl[0] vdd gnd cell_6t
Xbit_r1_c206 bl[206] br[206] wl[1] vdd gnd cell_6t
Xbit_r2_c206 bl[206] br[206] wl[2] vdd gnd cell_6t
Xbit_r3_c206 bl[206] br[206] wl[3] vdd gnd cell_6t
Xbit_r4_c206 bl[206] br[206] wl[4] vdd gnd cell_6t
Xbit_r5_c206 bl[206] br[206] wl[5] vdd gnd cell_6t
Xbit_r6_c206 bl[206] br[206] wl[6] vdd gnd cell_6t
Xbit_r7_c206 bl[206] br[206] wl[7] vdd gnd cell_6t
Xbit_r8_c206 bl[206] br[206] wl[8] vdd gnd cell_6t
Xbit_r9_c206 bl[206] br[206] wl[9] vdd gnd cell_6t
Xbit_r10_c206 bl[206] br[206] wl[10] vdd gnd cell_6t
Xbit_r11_c206 bl[206] br[206] wl[11] vdd gnd cell_6t
Xbit_r12_c206 bl[206] br[206] wl[12] vdd gnd cell_6t
Xbit_r13_c206 bl[206] br[206] wl[13] vdd gnd cell_6t
Xbit_r14_c206 bl[206] br[206] wl[14] vdd gnd cell_6t
Xbit_r15_c206 bl[206] br[206] wl[15] vdd gnd cell_6t
Xbit_r16_c206 bl[206] br[206] wl[16] vdd gnd cell_6t
Xbit_r17_c206 bl[206] br[206] wl[17] vdd gnd cell_6t
Xbit_r18_c206 bl[206] br[206] wl[18] vdd gnd cell_6t
Xbit_r19_c206 bl[206] br[206] wl[19] vdd gnd cell_6t
Xbit_r20_c206 bl[206] br[206] wl[20] vdd gnd cell_6t
Xbit_r21_c206 bl[206] br[206] wl[21] vdd gnd cell_6t
Xbit_r22_c206 bl[206] br[206] wl[22] vdd gnd cell_6t
Xbit_r23_c206 bl[206] br[206] wl[23] vdd gnd cell_6t
Xbit_r24_c206 bl[206] br[206] wl[24] vdd gnd cell_6t
Xbit_r25_c206 bl[206] br[206] wl[25] vdd gnd cell_6t
Xbit_r26_c206 bl[206] br[206] wl[26] vdd gnd cell_6t
Xbit_r27_c206 bl[206] br[206] wl[27] vdd gnd cell_6t
Xbit_r28_c206 bl[206] br[206] wl[28] vdd gnd cell_6t
Xbit_r29_c206 bl[206] br[206] wl[29] vdd gnd cell_6t
Xbit_r30_c206 bl[206] br[206] wl[30] vdd gnd cell_6t
Xbit_r31_c206 bl[206] br[206] wl[31] vdd gnd cell_6t
Xbit_r32_c206 bl[206] br[206] wl[32] vdd gnd cell_6t
Xbit_r33_c206 bl[206] br[206] wl[33] vdd gnd cell_6t
Xbit_r34_c206 bl[206] br[206] wl[34] vdd gnd cell_6t
Xbit_r35_c206 bl[206] br[206] wl[35] vdd gnd cell_6t
Xbit_r36_c206 bl[206] br[206] wl[36] vdd gnd cell_6t
Xbit_r37_c206 bl[206] br[206] wl[37] vdd gnd cell_6t
Xbit_r38_c206 bl[206] br[206] wl[38] vdd gnd cell_6t
Xbit_r39_c206 bl[206] br[206] wl[39] vdd gnd cell_6t
Xbit_r40_c206 bl[206] br[206] wl[40] vdd gnd cell_6t
Xbit_r41_c206 bl[206] br[206] wl[41] vdd gnd cell_6t
Xbit_r42_c206 bl[206] br[206] wl[42] vdd gnd cell_6t
Xbit_r43_c206 bl[206] br[206] wl[43] vdd gnd cell_6t
Xbit_r44_c206 bl[206] br[206] wl[44] vdd gnd cell_6t
Xbit_r45_c206 bl[206] br[206] wl[45] vdd gnd cell_6t
Xbit_r46_c206 bl[206] br[206] wl[46] vdd gnd cell_6t
Xbit_r47_c206 bl[206] br[206] wl[47] vdd gnd cell_6t
Xbit_r48_c206 bl[206] br[206] wl[48] vdd gnd cell_6t
Xbit_r49_c206 bl[206] br[206] wl[49] vdd gnd cell_6t
Xbit_r50_c206 bl[206] br[206] wl[50] vdd gnd cell_6t
Xbit_r51_c206 bl[206] br[206] wl[51] vdd gnd cell_6t
Xbit_r52_c206 bl[206] br[206] wl[52] vdd gnd cell_6t
Xbit_r53_c206 bl[206] br[206] wl[53] vdd gnd cell_6t
Xbit_r54_c206 bl[206] br[206] wl[54] vdd gnd cell_6t
Xbit_r55_c206 bl[206] br[206] wl[55] vdd gnd cell_6t
Xbit_r56_c206 bl[206] br[206] wl[56] vdd gnd cell_6t
Xbit_r57_c206 bl[206] br[206] wl[57] vdd gnd cell_6t
Xbit_r58_c206 bl[206] br[206] wl[58] vdd gnd cell_6t
Xbit_r59_c206 bl[206] br[206] wl[59] vdd gnd cell_6t
Xbit_r60_c206 bl[206] br[206] wl[60] vdd gnd cell_6t
Xbit_r61_c206 bl[206] br[206] wl[61] vdd gnd cell_6t
Xbit_r62_c206 bl[206] br[206] wl[62] vdd gnd cell_6t
Xbit_r63_c206 bl[206] br[206] wl[63] vdd gnd cell_6t
Xbit_r64_c206 bl[206] br[206] wl[64] vdd gnd cell_6t
Xbit_r65_c206 bl[206] br[206] wl[65] vdd gnd cell_6t
Xbit_r66_c206 bl[206] br[206] wl[66] vdd gnd cell_6t
Xbit_r67_c206 bl[206] br[206] wl[67] vdd gnd cell_6t
Xbit_r68_c206 bl[206] br[206] wl[68] vdd gnd cell_6t
Xbit_r69_c206 bl[206] br[206] wl[69] vdd gnd cell_6t
Xbit_r70_c206 bl[206] br[206] wl[70] vdd gnd cell_6t
Xbit_r71_c206 bl[206] br[206] wl[71] vdd gnd cell_6t
Xbit_r72_c206 bl[206] br[206] wl[72] vdd gnd cell_6t
Xbit_r73_c206 bl[206] br[206] wl[73] vdd gnd cell_6t
Xbit_r74_c206 bl[206] br[206] wl[74] vdd gnd cell_6t
Xbit_r75_c206 bl[206] br[206] wl[75] vdd gnd cell_6t
Xbit_r76_c206 bl[206] br[206] wl[76] vdd gnd cell_6t
Xbit_r77_c206 bl[206] br[206] wl[77] vdd gnd cell_6t
Xbit_r78_c206 bl[206] br[206] wl[78] vdd gnd cell_6t
Xbit_r79_c206 bl[206] br[206] wl[79] vdd gnd cell_6t
Xbit_r80_c206 bl[206] br[206] wl[80] vdd gnd cell_6t
Xbit_r81_c206 bl[206] br[206] wl[81] vdd gnd cell_6t
Xbit_r82_c206 bl[206] br[206] wl[82] vdd gnd cell_6t
Xbit_r83_c206 bl[206] br[206] wl[83] vdd gnd cell_6t
Xbit_r84_c206 bl[206] br[206] wl[84] vdd gnd cell_6t
Xbit_r85_c206 bl[206] br[206] wl[85] vdd gnd cell_6t
Xbit_r86_c206 bl[206] br[206] wl[86] vdd gnd cell_6t
Xbit_r87_c206 bl[206] br[206] wl[87] vdd gnd cell_6t
Xbit_r88_c206 bl[206] br[206] wl[88] vdd gnd cell_6t
Xbit_r89_c206 bl[206] br[206] wl[89] vdd gnd cell_6t
Xbit_r90_c206 bl[206] br[206] wl[90] vdd gnd cell_6t
Xbit_r91_c206 bl[206] br[206] wl[91] vdd gnd cell_6t
Xbit_r92_c206 bl[206] br[206] wl[92] vdd gnd cell_6t
Xbit_r93_c206 bl[206] br[206] wl[93] vdd gnd cell_6t
Xbit_r94_c206 bl[206] br[206] wl[94] vdd gnd cell_6t
Xbit_r95_c206 bl[206] br[206] wl[95] vdd gnd cell_6t
Xbit_r96_c206 bl[206] br[206] wl[96] vdd gnd cell_6t
Xbit_r97_c206 bl[206] br[206] wl[97] vdd gnd cell_6t
Xbit_r98_c206 bl[206] br[206] wl[98] vdd gnd cell_6t
Xbit_r99_c206 bl[206] br[206] wl[99] vdd gnd cell_6t
Xbit_r100_c206 bl[206] br[206] wl[100] vdd gnd cell_6t
Xbit_r101_c206 bl[206] br[206] wl[101] vdd gnd cell_6t
Xbit_r102_c206 bl[206] br[206] wl[102] vdd gnd cell_6t
Xbit_r103_c206 bl[206] br[206] wl[103] vdd gnd cell_6t
Xbit_r104_c206 bl[206] br[206] wl[104] vdd gnd cell_6t
Xbit_r105_c206 bl[206] br[206] wl[105] vdd gnd cell_6t
Xbit_r106_c206 bl[206] br[206] wl[106] vdd gnd cell_6t
Xbit_r107_c206 bl[206] br[206] wl[107] vdd gnd cell_6t
Xbit_r108_c206 bl[206] br[206] wl[108] vdd gnd cell_6t
Xbit_r109_c206 bl[206] br[206] wl[109] vdd gnd cell_6t
Xbit_r110_c206 bl[206] br[206] wl[110] vdd gnd cell_6t
Xbit_r111_c206 bl[206] br[206] wl[111] vdd gnd cell_6t
Xbit_r112_c206 bl[206] br[206] wl[112] vdd gnd cell_6t
Xbit_r113_c206 bl[206] br[206] wl[113] vdd gnd cell_6t
Xbit_r114_c206 bl[206] br[206] wl[114] vdd gnd cell_6t
Xbit_r115_c206 bl[206] br[206] wl[115] vdd gnd cell_6t
Xbit_r116_c206 bl[206] br[206] wl[116] vdd gnd cell_6t
Xbit_r117_c206 bl[206] br[206] wl[117] vdd gnd cell_6t
Xbit_r118_c206 bl[206] br[206] wl[118] vdd gnd cell_6t
Xbit_r119_c206 bl[206] br[206] wl[119] vdd gnd cell_6t
Xbit_r120_c206 bl[206] br[206] wl[120] vdd gnd cell_6t
Xbit_r121_c206 bl[206] br[206] wl[121] vdd gnd cell_6t
Xbit_r122_c206 bl[206] br[206] wl[122] vdd gnd cell_6t
Xbit_r123_c206 bl[206] br[206] wl[123] vdd gnd cell_6t
Xbit_r124_c206 bl[206] br[206] wl[124] vdd gnd cell_6t
Xbit_r125_c206 bl[206] br[206] wl[125] vdd gnd cell_6t
Xbit_r126_c206 bl[206] br[206] wl[126] vdd gnd cell_6t
Xbit_r127_c206 bl[206] br[206] wl[127] vdd gnd cell_6t
Xbit_r128_c206 bl[206] br[206] wl[128] vdd gnd cell_6t
Xbit_r129_c206 bl[206] br[206] wl[129] vdd gnd cell_6t
Xbit_r130_c206 bl[206] br[206] wl[130] vdd gnd cell_6t
Xbit_r131_c206 bl[206] br[206] wl[131] vdd gnd cell_6t
Xbit_r132_c206 bl[206] br[206] wl[132] vdd gnd cell_6t
Xbit_r133_c206 bl[206] br[206] wl[133] vdd gnd cell_6t
Xbit_r134_c206 bl[206] br[206] wl[134] vdd gnd cell_6t
Xbit_r135_c206 bl[206] br[206] wl[135] vdd gnd cell_6t
Xbit_r136_c206 bl[206] br[206] wl[136] vdd gnd cell_6t
Xbit_r137_c206 bl[206] br[206] wl[137] vdd gnd cell_6t
Xbit_r138_c206 bl[206] br[206] wl[138] vdd gnd cell_6t
Xbit_r139_c206 bl[206] br[206] wl[139] vdd gnd cell_6t
Xbit_r140_c206 bl[206] br[206] wl[140] vdd gnd cell_6t
Xbit_r141_c206 bl[206] br[206] wl[141] vdd gnd cell_6t
Xbit_r142_c206 bl[206] br[206] wl[142] vdd gnd cell_6t
Xbit_r143_c206 bl[206] br[206] wl[143] vdd gnd cell_6t
Xbit_r144_c206 bl[206] br[206] wl[144] vdd gnd cell_6t
Xbit_r145_c206 bl[206] br[206] wl[145] vdd gnd cell_6t
Xbit_r146_c206 bl[206] br[206] wl[146] vdd gnd cell_6t
Xbit_r147_c206 bl[206] br[206] wl[147] vdd gnd cell_6t
Xbit_r148_c206 bl[206] br[206] wl[148] vdd gnd cell_6t
Xbit_r149_c206 bl[206] br[206] wl[149] vdd gnd cell_6t
Xbit_r150_c206 bl[206] br[206] wl[150] vdd gnd cell_6t
Xbit_r151_c206 bl[206] br[206] wl[151] vdd gnd cell_6t
Xbit_r152_c206 bl[206] br[206] wl[152] vdd gnd cell_6t
Xbit_r153_c206 bl[206] br[206] wl[153] vdd gnd cell_6t
Xbit_r154_c206 bl[206] br[206] wl[154] vdd gnd cell_6t
Xbit_r155_c206 bl[206] br[206] wl[155] vdd gnd cell_6t
Xbit_r156_c206 bl[206] br[206] wl[156] vdd gnd cell_6t
Xbit_r157_c206 bl[206] br[206] wl[157] vdd gnd cell_6t
Xbit_r158_c206 bl[206] br[206] wl[158] vdd gnd cell_6t
Xbit_r159_c206 bl[206] br[206] wl[159] vdd gnd cell_6t
Xbit_r160_c206 bl[206] br[206] wl[160] vdd gnd cell_6t
Xbit_r161_c206 bl[206] br[206] wl[161] vdd gnd cell_6t
Xbit_r162_c206 bl[206] br[206] wl[162] vdd gnd cell_6t
Xbit_r163_c206 bl[206] br[206] wl[163] vdd gnd cell_6t
Xbit_r164_c206 bl[206] br[206] wl[164] vdd gnd cell_6t
Xbit_r165_c206 bl[206] br[206] wl[165] vdd gnd cell_6t
Xbit_r166_c206 bl[206] br[206] wl[166] vdd gnd cell_6t
Xbit_r167_c206 bl[206] br[206] wl[167] vdd gnd cell_6t
Xbit_r168_c206 bl[206] br[206] wl[168] vdd gnd cell_6t
Xbit_r169_c206 bl[206] br[206] wl[169] vdd gnd cell_6t
Xbit_r170_c206 bl[206] br[206] wl[170] vdd gnd cell_6t
Xbit_r171_c206 bl[206] br[206] wl[171] vdd gnd cell_6t
Xbit_r172_c206 bl[206] br[206] wl[172] vdd gnd cell_6t
Xbit_r173_c206 bl[206] br[206] wl[173] vdd gnd cell_6t
Xbit_r174_c206 bl[206] br[206] wl[174] vdd gnd cell_6t
Xbit_r175_c206 bl[206] br[206] wl[175] vdd gnd cell_6t
Xbit_r176_c206 bl[206] br[206] wl[176] vdd gnd cell_6t
Xbit_r177_c206 bl[206] br[206] wl[177] vdd gnd cell_6t
Xbit_r178_c206 bl[206] br[206] wl[178] vdd gnd cell_6t
Xbit_r179_c206 bl[206] br[206] wl[179] vdd gnd cell_6t
Xbit_r180_c206 bl[206] br[206] wl[180] vdd gnd cell_6t
Xbit_r181_c206 bl[206] br[206] wl[181] vdd gnd cell_6t
Xbit_r182_c206 bl[206] br[206] wl[182] vdd gnd cell_6t
Xbit_r183_c206 bl[206] br[206] wl[183] vdd gnd cell_6t
Xbit_r184_c206 bl[206] br[206] wl[184] vdd gnd cell_6t
Xbit_r185_c206 bl[206] br[206] wl[185] vdd gnd cell_6t
Xbit_r186_c206 bl[206] br[206] wl[186] vdd gnd cell_6t
Xbit_r187_c206 bl[206] br[206] wl[187] vdd gnd cell_6t
Xbit_r188_c206 bl[206] br[206] wl[188] vdd gnd cell_6t
Xbit_r189_c206 bl[206] br[206] wl[189] vdd gnd cell_6t
Xbit_r190_c206 bl[206] br[206] wl[190] vdd gnd cell_6t
Xbit_r191_c206 bl[206] br[206] wl[191] vdd gnd cell_6t
Xbit_r192_c206 bl[206] br[206] wl[192] vdd gnd cell_6t
Xbit_r193_c206 bl[206] br[206] wl[193] vdd gnd cell_6t
Xbit_r194_c206 bl[206] br[206] wl[194] vdd gnd cell_6t
Xbit_r195_c206 bl[206] br[206] wl[195] vdd gnd cell_6t
Xbit_r196_c206 bl[206] br[206] wl[196] vdd gnd cell_6t
Xbit_r197_c206 bl[206] br[206] wl[197] vdd gnd cell_6t
Xbit_r198_c206 bl[206] br[206] wl[198] vdd gnd cell_6t
Xbit_r199_c206 bl[206] br[206] wl[199] vdd gnd cell_6t
Xbit_r200_c206 bl[206] br[206] wl[200] vdd gnd cell_6t
Xbit_r201_c206 bl[206] br[206] wl[201] vdd gnd cell_6t
Xbit_r202_c206 bl[206] br[206] wl[202] vdd gnd cell_6t
Xbit_r203_c206 bl[206] br[206] wl[203] vdd gnd cell_6t
Xbit_r204_c206 bl[206] br[206] wl[204] vdd gnd cell_6t
Xbit_r205_c206 bl[206] br[206] wl[205] vdd gnd cell_6t
Xbit_r206_c206 bl[206] br[206] wl[206] vdd gnd cell_6t
Xbit_r207_c206 bl[206] br[206] wl[207] vdd gnd cell_6t
Xbit_r208_c206 bl[206] br[206] wl[208] vdd gnd cell_6t
Xbit_r209_c206 bl[206] br[206] wl[209] vdd gnd cell_6t
Xbit_r210_c206 bl[206] br[206] wl[210] vdd gnd cell_6t
Xbit_r211_c206 bl[206] br[206] wl[211] vdd gnd cell_6t
Xbit_r212_c206 bl[206] br[206] wl[212] vdd gnd cell_6t
Xbit_r213_c206 bl[206] br[206] wl[213] vdd gnd cell_6t
Xbit_r214_c206 bl[206] br[206] wl[214] vdd gnd cell_6t
Xbit_r215_c206 bl[206] br[206] wl[215] vdd gnd cell_6t
Xbit_r216_c206 bl[206] br[206] wl[216] vdd gnd cell_6t
Xbit_r217_c206 bl[206] br[206] wl[217] vdd gnd cell_6t
Xbit_r218_c206 bl[206] br[206] wl[218] vdd gnd cell_6t
Xbit_r219_c206 bl[206] br[206] wl[219] vdd gnd cell_6t
Xbit_r220_c206 bl[206] br[206] wl[220] vdd gnd cell_6t
Xbit_r221_c206 bl[206] br[206] wl[221] vdd gnd cell_6t
Xbit_r222_c206 bl[206] br[206] wl[222] vdd gnd cell_6t
Xbit_r223_c206 bl[206] br[206] wl[223] vdd gnd cell_6t
Xbit_r224_c206 bl[206] br[206] wl[224] vdd gnd cell_6t
Xbit_r225_c206 bl[206] br[206] wl[225] vdd gnd cell_6t
Xbit_r226_c206 bl[206] br[206] wl[226] vdd gnd cell_6t
Xbit_r227_c206 bl[206] br[206] wl[227] vdd gnd cell_6t
Xbit_r228_c206 bl[206] br[206] wl[228] vdd gnd cell_6t
Xbit_r229_c206 bl[206] br[206] wl[229] vdd gnd cell_6t
Xbit_r230_c206 bl[206] br[206] wl[230] vdd gnd cell_6t
Xbit_r231_c206 bl[206] br[206] wl[231] vdd gnd cell_6t
Xbit_r232_c206 bl[206] br[206] wl[232] vdd gnd cell_6t
Xbit_r233_c206 bl[206] br[206] wl[233] vdd gnd cell_6t
Xbit_r234_c206 bl[206] br[206] wl[234] vdd gnd cell_6t
Xbit_r235_c206 bl[206] br[206] wl[235] vdd gnd cell_6t
Xbit_r236_c206 bl[206] br[206] wl[236] vdd gnd cell_6t
Xbit_r237_c206 bl[206] br[206] wl[237] vdd gnd cell_6t
Xbit_r238_c206 bl[206] br[206] wl[238] vdd gnd cell_6t
Xbit_r239_c206 bl[206] br[206] wl[239] vdd gnd cell_6t
Xbit_r240_c206 bl[206] br[206] wl[240] vdd gnd cell_6t
Xbit_r241_c206 bl[206] br[206] wl[241] vdd gnd cell_6t
Xbit_r242_c206 bl[206] br[206] wl[242] vdd gnd cell_6t
Xbit_r243_c206 bl[206] br[206] wl[243] vdd gnd cell_6t
Xbit_r244_c206 bl[206] br[206] wl[244] vdd gnd cell_6t
Xbit_r245_c206 bl[206] br[206] wl[245] vdd gnd cell_6t
Xbit_r246_c206 bl[206] br[206] wl[246] vdd gnd cell_6t
Xbit_r247_c206 bl[206] br[206] wl[247] vdd gnd cell_6t
Xbit_r248_c206 bl[206] br[206] wl[248] vdd gnd cell_6t
Xbit_r249_c206 bl[206] br[206] wl[249] vdd gnd cell_6t
Xbit_r250_c206 bl[206] br[206] wl[250] vdd gnd cell_6t
Xbit_r251_c206 bl[206] br[206] wl[251] vdd gnd cell_6t
Xbit_r252_c206 bl[206] br[206] wl[252] vdd gnd cell_6t
Xbit_r253_c206 bl[206] br[206] wl[253] vdd gnd cell_6t
Xbit_r254_c206 bl[206] br[206] wl[254] vdd gnd cell_6t
Xbit_r255_c206 bl[206] br[206] wl[255] vdd gnd cell_6t
Xbit_r0_c207 bl[207] br[207] wl[0] vdd gnd cell_6t
Xbit_r1_c207 bl[207] br[207] wl[1] vdd gnd cell_6t
Xbit_r2_c207 bl[207] br[207] wl[2] vdd gnd cell_6t
Xbit_r3_c207 bl[207] br[207] wl[3] vdd gnd cell_6t
Xbit_r4_c207 bl[207] br[207] wl[4] vdd gnd cell_6t
Xbit_r5_c207 bl[207] br[207] wl[5] vdd gnd cell_6t
Xbit_r6_c207 bl[207] br[207] wl[6] vdd gnd cell_6t
Xbit_r7_c207 bl[207] br[207] wl[7] vdd gnd cell_6t
Xbit_r8_c207 bl[207] br[207] wl[8] vdd gnd cell_6t
Xbit_r9_c207 bl[207] br[207] wl[9] vdd gnd cell_6t
Xbit_r10_c207 bl[207] br[207] wl[10] vdd gnd cell_6t
Xbit_r11_c207 bl[207] br[207] wl[11] vdd gnd cell_6t
Xbit_r12_c207 bl[207] br[207] wl[12] vdd gnd cell_6t
Xbit_r13_c207 bl[207] br[207] wl[13] vdd gnd cell_6t
Xbit_r14_c207 bl[207] br[207] wl[14] vdd gnd cell_6t
Xbit_r15_c207 bl[207] br[207] wl[15] vdd gnd cell_6t
Xbit_r16_c207 bl[207] br[207] wl[16] vdd gnd cell_6t
Xbit_r17_c207 bl[207] br[207] wl[17] vdd gnd cell_6t
Xbit_r18_c207 bl[207] br[207] wl[18] vdd gnd cell_6t
Xbit_r19_c207 bl[207] br[207] wl[19] vdd gnd cell_6t
Xbit_r20_c207 bl[207] br[207] wl[20] vdd gnd cell_6t
Xbit_r21_c207 bl[207] br[207] wl[21] vdd gnd cell_6t
Xbit_r22_c207 bl[207] br[207] wl[22] vdd gnd cell_6t
Xbit_r23_c207 bl[207] br[207] wl[23] vdd gnd cell_6t
Xbit_r24_c207 bl[207] br[207] wl[24] vdd gnd cell_6t
Xbit_r25_c207 bl[207] br[207] wl[25] vdd gnd cell_6t
Xbit_r26_c207 bl[207] br[207] wl[26] vdd gnd cell_6t
Xbit_r27_c207 bl[207] br[207] wl[27] vdd gnd cell_6t
Xbit_r28_c207 bl[207] br[207] wl[28] vdd gnd cell_6t
Xbit_r29_c207 bl[207] br[207] wl[29] vdd gnd cell_6t
Xbit_r30_c207 bl[207] br[207] wl[30] vdd gnd cell_6t
Xbit_r31_c207 bl[207] br[207] wl[31] vdd gnd cell_6t
Xbit_r32_c207 bl[207] br[207] wl[32] vdd gnd cell_6t
Xbit_r33_c207 bl[207] br[207] wl[33] vdd gnd cell_6t
Xbit_r34_c207 bl[207] br[207] wl[34] vdd gnd cell_6t
Xbit_r35_c207 bl[207] br[207] wl[35] vdd gnd cell_6t
Xbit_r36_c207 bl[207] br[207] wl[36] vdd gnd cell_6t
Xbit_r37_c207 bl[207] br[207] wl[37] vdd gnd cell_6t
Xbit_r38_c207 bl[207] br[207] wl[38] vdd gnd cell_6t
Xbit_r39_c207 bl[207] br[207] wl[39] vdd gnd cell_6t
Xbit_r40_c207 bl[207] br[207] wl[40] vdd gnd cell_6t
Xbit_r41_c207 bl[207] br[207] wl[41] vdd gnd cell_6t
Xbit_r42_c207 bl[207] br[207] wl[42] vdd gnd cell_6t
Xbit_r43_c207 bl[207] br[207] wl[43] vdd gnd cell_6t
Xbit_r44_c207 bl[207] br[207] wl[44] vdd gnd cell_6t
Xbit_r45_c207 bl[207] br[207] wl[45] vdd gnd cell_6t
Xbit_r46_c207 bl[207] br[207] wl[46] vdd gnd cell_6t
Xbit_r47_c207 bl[207] br[207] wl[47] vdd gnd cell_6t
Xbit_r48_c207 bl[207] br[207] wl[48] vdd gnd cell_6t
Xbit_r49_c207 bl[207] br[207] wl[49] vdd gnd cell_6t
Xbit_r50_c207 bl[207] br[207] wl[50] vdd gnd cell_6t
Xbit_r51_c207 bl[207] br[207] wl[51] vdd gnd cell_6t
Xbit_r52_c207 bl[207] br[207] wl[52] vdd gnd cell_6t
Xbit_r53_c207 bl[207] br[207] wl[53] vdd gnd cell_6t
Xbit_r54_c207 bl[207] br[207] wl[54] vdd gnd cell_6t
Xbit_r55_c207 bl[207] br[207] wl[55] vdd gnd cell_6t
Xbit_r56_c207 bl[207] br[207] wl[56] vdd gnd cell_6t
Xbit_r57_c207 bl[207] br[207] wl[57] vdd gnd cell_6t
Xbit_r58_c207 bl[207] br[207] wl[58] vdd gnd cell_6t
Xbit_r59_c207 bl[207] br[207] wl[59] vdd gnd cell_6t
Xbit_r60_c207 bl[207] br[207] wl[60] vdd gnd cell_6t
Xbit_r61_c207 bl[207] br[207] wl[61] vdd gnd cell_6t
Xbit_r62_c207 bl[207] br[207] wl[62] vdd gnd cell_6t
Xbit_r63_c207 bl[207] br[207] wl[63] vdd gnd cell_6t
Xbit_r64_c207 bl[207] br[207] wl[64] vdd gnd cell_6t
Xbit_r65_c207 bl[207] br[207] wl[65] vdd gnd cell_6t
Xbit_r66_c207 bl[207] br[207] wl[66] vdd gnd cell_6t
Xbit_r67_c207 bl[207] br[207] wl[67] vdd gnd cell_6t
Xbit_r68_c207 bl[207] br[207] wl[68] vdd gnd cell_6t
Xbit_r69_c207 bl[207] br[207] wl[69] vdd gnd cell_6t
Xbit_r70_c207 bl[207] br[207] wl[70] vdd gnd cell_6t
Xbit_r71_c207 bl[207] br[207] wl[71] vdd gnd cell_6t
Xbit_r72_c207 bl[207] br[207] wl[72] vdd gnd cell_6t
Xbit_r73_c207 bl[207] br[207] wl[73] vdd gnd cell_6t
Xbit_r74_c207 bl[207] br[207] wl[74] vdd gnd cell_6t
Xbit_r75_c207 bl[207] br[207] wl[75] vdd gnd cell_6t
Xbit_r76_c207 bl[207] br[207] wl[76] vdd gnd cell_6t
Xbit_r77_c207 bl[207] br[207] wl[77] vdd gnd cell_6t
Xbit_r78_c207 bl[207] br[207] wl[78] vdd gnd cell_6t
Xbit_r79_c207 bl[207] br[207] wl[79] vdd gnd cell_6t
Xbit_r80_c207 bl[207] br[207] wl[80] vdd gnd cell_6t
Xbit_r81_c207 bl[207] br[207] wl[81] vdd gnd cell_6t
Xbit_r82_c207 bl[207] br[207] wl[82] vdd gnd cell_6t
Xbit_r83_c207 bl[207] br[207] wl[83] vdd gnd cell_6t
Xbit_r84_c207 bl[207] br[207] wl[84] vdd gnd cell_6t
Xbit_r85_c207 bl[207] br[207] wl[85] vdd gnd cell_6t
Xbit_r86_c207 bl[207] br[207] wl[86] vdd gnd cell_6t
Xbit_r87_c207 bl[207] br[207] wl[87] vdd gnd cell_6t
Xbit_r88_c207 bl[207] br[207] wl[88] vdd gnd cell_6t
Xbit_r89_c207 bl[207] br[207] wl[89] vdd gnd cell_6t
Xbit_r90_c207 bl[207] br[207] wl[90] vdd gnd cell_6t
Xbit_r91_c207 bl[207] br[207] wl[91] vdd gnd cell_6t
Xbit_r92_c207 bl[207] br[207] wl[92] vdd gnd cell_6t
Xbit_r93_c207 bl[207] br[207] wl[93] vdd gnd cell_6t
Xbit_r94_c207 bl[207] br[207] wl[94] vdd gnd cell_6t
Xbit_r95_c207 bl[207] br[207] wl[95] vdd gnd cell_6t
Xbit_r96_c207 bl[207] br[207] wl[96] vdd gnd cell_6t
Xbit_r97_c207 bl[207] br[207] wl[97] vdd gnd cell_6t
Xbit_r98_c207 bl[207] br[207] wl[98] vdd gnd cell_6t
Xbit_r99_c207 bl[207] br[207] wl[99] vdd gnd cell_6t
Xbit_r100_c207 bl[207] br[207] wl[100] vdd gnd cell_6t
Xbit_r101_c207 bl[207] br[207] wl[101] vdd gnd cell_6t
Xbit_r102_c207 bl[207] br[207] wl[102] vdd gnd cell_6t
Xbit_r103_c207 bl[207] br[207] wl[103] vdd gnd cell_6t
Xbit_r104_c207 bl[207] br[207] wl[104] vdd gnd cell_6t
Xbit_r105_c207 bl[207] br[207] wl[105] vdd gnd cell_6t
Xbit_r106_c207 bl[207] br[207] wl[106] vdd gnd cell_6t
Xbit_r107_c207 bl[207] br[207] wl[107] vdd gnd cell_6t
Xbit_r108_c207 bl[207] br[207] wl[108] vdd gnd cell_6t
Xbit_r109_c207 bl[207] br[207] wl[109] vdd gnd cell_6t
Xbit_r110_c207 bl[207] br[207] wl[110] vdd gnd cell_6t
Xbit_r111_c207 bl[207] br[207] wl[111] vdd gnd cell_6t
Xbit_r112_c207 bl[207] br[207] wl[112] vdd gnd cell_6t
Xbit_r113_c207 bl[207] br[207] wl[113] vdd gnd cell_6t
Xbit_r114_c207 bl[207] br[207] wl[114] vdd gnd cell_6t
Xbit_r115_c207 bl[207] br[207] wl[115] vdd gnd cell_6t
Xbit_r116_c207 bl[207] br[207] wl[116] vdd gnd cell_6t
Xbit_r117_c207 bl[207] br[207] wl[117] vdd gnd cell_6t
Xbit_r118_c207 bl[207] br[207] wl[118] vdd gnd cell_6t
Xbit_r119_c207 bl[207] br[207] wl[119] vdd gnd cell_6t
Xbit_r120_c207 bl[207] br[207] wl[120] vdd gnd cell_6t
Xbit_r121_c207 bl[207] br[207] wl[121] vdd gnd cell_6t
Xbit_r122_c207 bl[207] br[207] wl[122] vdd gnd cell_6t
Xbit_r123_c207 bl[207] br[207] wl[123] vdd gnd cell_6t
Xbit_r124_c207 bl[207] br[207] wl[124] vdd gnd cell_6t
Xbit_r125_c207 bl[207] br[207] wl[125] vdd gnd cell_6t
Xbit_r126_c207 bl[207] br[207] wl[126] vdd gnd cell_6t
Xbit_r127_c207 bl[207] br[207] wl[127] vdd gnd cell_6t
Xbit_r128_c207 bl[207] br[207] wl[128] vdd gnd cell_6t
Xbit_r129_c207 bl[207] br[207] wl[129] vdd gnd cell_6t
Xbit_r130_c207 bl[207] br[207] wl[130] vdd gnd cell_6t
Xbit_r131_c207 bl[207] br[207] wl[131] vdd gnd cell_6t
Xbit_r132_c207 bl[207] br[207] wl[132] vdd gnd cell_6t
Xbit_r133_c207 bl[207] br[207] wl[133] vdd gnd cell_6t
Xbit_r134_c207 bl[207] br[207] wl[134] vdd gnd cell_6t
Xbit_r135_c207 bl[207] br[207] wl[135] vdd gnd cell_6t
Xbit_r136_c207 bl[207] br[207] wl[136] vdd gnd cell_6t
Xbit_r137_c207 bl[207] br[207] wl[137] vdd gnd cell_6t
Xbit_r138_c207 bl[207] br[207] wl[138] vdd gnd cell_6t
Xbit_r139_c207 bl[207] br[207] wl[139] vdd gnd cell_6t
Xbit_r140_c207 bl[207] br[207] wl[140] vdd gnd cell_6t
Xbit_r141_c207 bl[207] br[207] wl[141] vdd gnd cell_6t
Xbit_r142_c207 bl[207] br[207] wl[142] vdd gnd cell_6t
Xbit_r143_c207 bl[207] br[207] wl[143] vdd gnd cell_6t
Xbit_r144_c207 bl[207] br[207] wl[144] vdd gnd cell_6t
Xbit_r145_c207 bl[207] br[207] wl[145] vdd gnd cell_6t
Xbit_r146_c207 bl[207] br[207] wl[146] vdd gnd cell_6t
Xbit_r147_c207 bl[207] br[207] wl[147] vdd gnd cell_6t
Xbit_r148_c207 bl[207] br[207] wl[148] vdd gnd cell_6t
Xbit_r149_c207 bl[207] br[207] wl[149] vdd gnd cell_6t
Xbit_r150_c207 bl[207] br[207] wl[150] vdd gnd cell_6t
Xbit_r151_c207 bl[207] br[207] wl[151] vdd gnd cell_6t
Xbit_r152_c207 bl[207] br[207] wl[152] vdd gnd cell_6t
Xbit_r153_c207 bl[207] br[207] wl[153] vdd gnd cell_6t
Xbit_r154_c207 bl[207] br[207] wl[154] vdd gnd cell_6t
Xbit_r155_c207 bl[207] br[207] wl[155] vdd gnd cell_6t
Xbit_r156_c207 bl[207] br[207] wl[156] vdd gnd cell_6t
Xbit_r157_c207 bl[207] br[207] wl[157] vdd gnd cell_6t
Xbit_r158_c207 bl[207] br[207] wl[158] vdd gnd cell_6t
Xbit_r159_c207 bl[207] br[207] wl[159] vdd gnd cell_6t
Xbit_r160_c207 bl[207] br[207] wl[160] vdd gnd cell_6t
Xbit_r161_c207 bl[207] br[207] wl[161] vdd gnd cell_6t
Xbit_r162_c207 bl[207] br[207] wl[162] vdd gnd cell_6t
Xbit_r163_c207 bl[207] br[207] wl[163] vdd gnd cell_6t
Xbit_r164_c207 bl[207] br[207] wl[164] vdd gnd cell_6t
Xbit_r165_c207 bl[207] br[207] wl[165] vdd gnd cell_6t
Xbit_r166_c207 bl[207] br[207] wl[166] vdd gnd cell_6t
Xbit_r167_c207 bl[207] br[207] wl[167] vdd gnd cell_6t
Xbit_r168_c207 bl[207] br[207] wl[168] vdd gnd cell_6t
Xbit_r169_c207 bl[207] br[207] wl[169] vdd gnd cell_6t
Xbit_r170_c207 bl[207] br[207] wl[170] vdd gnd cell_6t
Xbit_r171_c207 bl[207] br[207] wl[171] vdd gnd cell_6t
Xbit_r172_c207 bl[207] br[207] wl[172] vdd gnd cell_6t
Xbit_r173_c207 bl[207] br[207] wl[173] vdd gnd cell_6t
Xbit_r174_c207 bl[207] br[207] wl[174] vdd gnd cell_6t
Xbit_r175_c207 bl[207] br[207] wl[175] vdd gnd cell_6t
Xbit_r176_c207 bl[207] br[207] wl[176] vdd gnd cell_6t
Xbit_r177_c207 bl[207] br[207] wl[177] vdd gnd cell_6t
Xbit_r178_c207 bl[207] br[207] wl[178] vdd gnd cell_6t
Xbit_r179_c207 bl[207] br[207] wl[179] vdd gnd cell_6t
Xbit_r180_c207 bl[207] br[207] wl[180] vdd gnd cell_6t
Xbit_r181_c207 bl[207] br[207] wl[181] vdd gnd cell_6t
Xbit_r182_c207 bl[207] br[207] wl[182] vdd gnd cell_6t
Xbit_r183_c207 bl[207] br[207] wl[183] vdd gnd cell_6t
Xbit_r184_c207 bl[207] br[207] wl[184] vdd gnd cell_6t
Xbit_r185_c207 bl[207] br[207] wl[185] vdd gnd cell_6t
Xbit_r186_c207 bl[207] br[207] wl[186] vdd gnd cell_6t
Xbit_r187_c207 bl[207] br[207] wl[187] vdd gnd cell_6t
Xbit_r188_c207 bl[207] br[207] wl[188] vdd gnd cell_6t
Xbit_r189_c207 bl[207] br[207] wl[189] vdd gnd cell_6t
Xbit_r190_c207 bl[207] br[207] wl[190] vdd gnd cell_6t
Xbit_r191_c207 bl[207] br[207] wl[191] vdd gnd cell_6t
Xbit_r192_c207 bl[207] br[207] wl[192] vdd gnd cell_6t
Xbit_r193_c207 bl[207] br[207] wl[193] vdd gnd cell_6t
Xbit_r194_c207 bl[207] br[207] wl[194] vdd gnd cell_6t
Xbit_r195_c207 bl[207] br[207] wl[195] vdd gnd cell_6t
Xbit_r196_c207 bl[207] br[207] wl[196] vdd gnd cell_6t
Xbit_r197_c207 bl[207] br[207] wl[197] vdd gnd cell_6t
Xbit_r198_c207 bl[207] br[207] wl[198] vdd gnd cell_6t
Xbit_r199_c207 bl[207] br[207] wl[199] vdd gnd cell_6t
Xbit_r200_c207 bl[207] br[207] wl[200] vdd gnd cell_6t
Xbit_r201_c207 bl[207] br[207] wl[201] vdd gnd cell_6t
Xbit_r202_c207 bl[207] br[207] wl[202] vdd gnd cell_6t
Xbit_r203_c207 bl[207] br[207] wl[203] vdd gnd cell_6t
Xbit_r204_c207 bl[207] br[207] wl[204] vdd gnd cell_6t
Xbit_r205_c207 bl[207] br[207] wl[205] vdd gnd cell_6t
Xbit_r206_c207 bl[207] br[207] wl[206] vdd gnd cell_6t
Xbit_r207_c207 bl[207] br[207] wl[207] vdd gnd cell_6t
Xbit_r208_c207 bl[207] br[207] wl[208] vdd gnd cell_6t
Xbit_r209_c207 bl[207] br[207] wl[209] vdd gnd cell_6t
Xbit_r210_c207 bl[207] br[207] wl[210] vdd gnd cell_6t
Xbit_r211_c207 bl[207] br[207] wl[211] vdd gnd cell_6t
Xbit_r212_c207 bl[207] br[207] wl[212] vdd gnd cell_6t
Xbit_r213_c207 bl[207] br[207] wl[213] vdd gnd cell_6t
Xbit_r214_c207 bl[207] br[207] wl[214] vdd gnd cell_6t
Xbit_r215_c207 bl[207] br[207] wl[215] vdd gnd cell_6t
Xbit_r216_c207 bl[207] br[207] wl[216] vdd gnd cell_6t
Xbit_r217_c207 bl[207] br[207] wl[217] vdd gnd cell_6t
Xbit_r218_c207 bl[207] br[207] wl[218] vdd gnd cell_6t
Xbit_r219_c207 bl[207] br[207] wl[219] vdd gnd cell_6t
Xbit_r220_c207 bl[207] br[207] wl[220] vdd gnd cell_6t
Xbit_r221_c207 bl[207] br[207] wl[221] vdd gnd cell_6t
Xbit_r222_c207 bl[207] br[207] wl[222] vdd gnd cell_6t
Xbit_r223_c207 bl[207] br[207] wl[223] vdd gnd cell_6t
Xbit_r224_c207 bl[207] br[207] wl[224] vdd gnd cell_6t
Xbit_r225_c207 bl[207] br[207] wl[225] vdd gnd cell_6t
Xbit_r226_c207 bl[207] br[207] wl[226] vdd gnd cell_6t
Xbit_r227_c207 bl[207] br[207] wl[227] vdd gnd cell_6t
Xbit_r228_c207 bl[207] br[207] wl[228] vdd gnd cell_6t
Xbit_r229_c207 bl[207] br[207] wl[229] vdd gnd cell_6t
Xbit_r230_c207 bl[207] br[207] wl[230] vdd gnd cell_6t
Xbit_r231_c207 bl[207] br[207] wl[231] vdd gnd cell_6t
Xbit_r232_c207 bl[207] br[207] wl[232] vdd gnd cell_6t
Xbit_r233_c207 bl[207] br[207] wl[233] vdd gnd cell_6t
Xbit_r234_c207 bl[207] br[207] wl[234] vdd gnd cell_6t
Xbit_r235_c207 bl[207] br[207] wl[235] vdd gnd cell_6t
Xbit_r236_c207 bl[207] br[207] wl[236] vdd gnd cell_6t
Xbit_r237_c207 bl[207] br[207] wl[237] vdd gnd cell_6t
Xbit_r238_c207 bl[207] br[207] wl[238] vdd gnd cell_6t
Xbit_r239_c207 bl[207] br[207] wl[239] vdd gnd cell_6t
Xbit_r240_c207 bl[207] br[207] wl[240] vdd gnd cell_6t
Xbit_r241_c207 bl[207] br[207] wl[241] vdd gnd cell_6t
Xbit_r242_c207 bl[207] br[207] wl[242] vdd gnd cell_6t
Xbit_r243_c207 bl[207] br[207] wl[243] vdd gnd cell_6t
Xbit_r244_c207 bl[207] br[207] wl[244] vdd gnd cell_6t
Xbit_r245_c207 bl[207] br[207] wl[245] vdd gnd cell_6t
Xbit_r246_c207 bl[207] br[207] wl[246] vdd gnd cell_6t
Xbit_r247_c207 bl[207] br[207] wl[247] vdd gnd cell_6t
Xbit_r248_c207 bl[207] br[207] wl[248] vdd gnd cell_6t
Xbit_r249_c207 bl[207] br[207] wl[249] vdd gnd cell_6t
Xbit_r250_c207 bl[207] br[207] wl[250] vdd gnd cell_6t
Xbit_r251_c207 bl[207] br[207] wl[251] vdd gnd cell_6t
Xbit_r252_c207 bl[207] br[207] wl[252] vdd gnd cell_6t
Xbit_r253_c207 bl[207] br[207] wl[253] vdd gnd cell_6t
Xbit_r254_c207 bl[207] br[207] wl[254] vdd gnd cell_6t
Xbit_r255_c207 bl[207] br[207] wl[255] vdd gnd cell_6t
Xbit_r0_c208 bl[208] br[208] wl[0] vdd gnd cell_6t
Xbit_r1_c208 bl[208] br[208] wl[1] vdd gnd cell_6t
Xbit_r2_c208 bl[208] br[208] wl[2] vdd gnd cell_6t
Xbit_r3_c208 bl[208] br[208] wl[3] vdd gnd cell_6t
Xbit_r4_c208 bl[208] br[208] wl[4] vdd gnd cell_6t
Xbit_r5_c208 bl[208] br[208] wl[5] vdd gnd cell_6t
Xbit_r6_c208 bl[208] br[208] wl[6] vdd gnd cell_6t
Xbit_r7_c208 bl[208] br[208] wl[7] vdd gnd cell_6t
Xbit_r8_c208 bl[208] br[208] wl[8] vdd gnd cell_6t
Xbit_r9_c208 bl[208] br[208] wl[9] vdd gnd cell_6t
Xbit_r10_c208 bl[208] br[208] wl[10] vdd gnd cell_6t
Xbit_r11_c208 bl[208] br[208] wl[11] vdd gnd cell_6t
Xbit_r12_c208 bl[208] br[208] wl[12] vdd gnd cell_6t
Xbit_r13_c208 bl[208] br[208] wl[13] vdd gnd cell_6t
Xbit_r14_c208 bl[208] br[208] wl[14] vdd gnd cell_6t
Xbit_r15_c208 bl[208] br[208] wl[15] vdd gnd cell_6t
Xbit_r16_c208 bl[208] br[208] wl[16] vdd gnd cell_6t
Xbit_r17_c208 bl[208] br[208] wl[17] vdd gnd cell_6t
Xbit_r18_c208 bl[208] br[208] wl[18] vdd gnd cell_6t
Xbit_r19_c208 bl[208] br[208] wl[19] vdd gnd cell_6t
Xbit_r20_c208 bl[208] br[208] wl[20] vdd gnd cell_6t
Xbit_r21_c208 bl[208] br[208] wl[21] vdd gnd cell_6t
Xbit_r22_c208 bl[208] br[208] wl[22] vdd gnd cell_6t
Xbit_r23_c208 bl[208] br[208] wl[23] vdd gnd cell_6t
Xbit_r24_c208 bl[208] br[208] wl[24] vdd gnd cell_6t
Xbit_r25_c208 bl[208] br[208] wl[25] vdd gnd cell_6t
Xbit_r26_c208 bl[208] br[208] wl[26] vdd gnd cell_6t
Xbit_r27_c208 bl[208] br[208] wl[27] vdd gnd cell_6t
Xbit_r28_c208 bl[208] br[208] wl[28] vdd gnd cell_6t
Xbit_r29_c208 bl[208] br[208] wl[29] vdd gnd cell_6t
Xbit_r30_c208 bl[208] br[208] wl[30] vdd gnd cell_6t
Xbit_r31_c208 bl[208] br[208] wl[31] vdd gnd cell_6t
Xbit_r32_c208 bl[208] br[208] wl[32] vdd gnd cell_6t
Xbit_r33_c208 bl[208] br[208] wl[33] vdd gnd cell_6t
Xbit_r34_c208 bl[208] br[208] wl[34] vdd gnd cell_6t
Xbit_r35_c208 bl[208] br[208] wl[35] vdd gnd cell_6t
Xbit_r36_c208 bl[208] br[208] wl[36] vdd gnd cell_6t
Xbit_r37_c208 bl[208] br[208] wl[37] vdd gnd cell_6t
Xbit_r38_c208 bl[208] br[208] wl[38] vdd gnd cell_6t
Xbit_r39_c208 bl[208] br[208] wl[39] vdd gnd cell_6t
Xbit_r40_c208 bl[208] br[208] wl[40] vdd gnd cell_6t
Xbit_r41_c208 bl[208] br[208] wl[41] vdd gnd cell_6t
Xbit_r42_c208 bl[208] br[208] wl[42] vdd gnd cell_6t
Xbit_r43_c208 bl[208] br[208] wl[43] vdd gnd cell_6t
Xbit_r44_c208 bl[208] br[208] wl[44] vdd gnd cell_6t
Xbit_r45_c208 bl[208] br[208] wl[45] vdd gnd cell_6t
Xbit_r46_c208 bl[208] br[208] wl[46] vdd gnd cell_6t
Xbit_r47_c208 bl[208] br[208] wl[47] vdd gnd cell_6t
Xbit_r48_c208 bl[208] br[208] wl[48] vdd gnd cell_6t
Xbit_r49_c208 bl[208] br[208] wl[49] vdd gnd cell_6t
Xbit_r50_c208 bl[208] br[208] wl[50] vdd gnd cell_6t
Xbit_r51_c208 bl[208] br[208] wl[51] vdd gnd cell_6t
Xbit_r52_c208 bl[208] br[208] wl[52] vdd gnd cell_6t
Xbit_r53_c208 bl[208] br[208] wl[53] vdd gnd cell_6t
Xbit_r54_c208 bl[208] br[208] wl[54] vdd gnd cell_6t
Xbit_r55_c208 bl[208] br[208] wl[55] vdd gnd cell_6t
Xbit_r56_c208 bl[208] br[208] wl[56] vdd gnd cell_6t
Xbit_r57_c208 bl[208] br[208] wl[57] vdd gnd cell_6t
Xbit_r58_c208 bl[208] br[208] wl[58] vdd gnd cell_6t
Xbit_r59_c208 bl[208] br[208] wl[59] vdd gnd cell_6t
Xbit_r60_c208 bl[208] br[208] wl[60] vdd gnd cell_6t
Xbit_r61_c208 bl[208] br[208] wl[61] vdd gnd cell_6t
Xbit_r62_c208 bl[208] br[208] wl[62] vdd gnd cell_6t
Xbit_r63_c208 bl[208] br[208] wl[63] vdd gnd cell_6t
Xbit_r64_c208 bl[208] br[208] wl[64] vdd gnd cell_6t
Xbit_r65_c208 bl[208] br[208] wl[65] vdd gnd cell_6t
Xbit_r66_c208 bl[208] br[208] wl[66] vdd gnd cell_6t
Xbit_r67_c208 bl[208] br[208] wl[67] vdd gnd cell_6t
Xbit_r68_c208 bl[208] br[208] wl[68] vdd gnd cell_6t
Xbit_r69_c208 bl[208] br[208] wl[69] vdd gnd cell_6t
Xbit_r70_c208 bl[208] br[208] wl[70] vdd gnd cell_6t
Xbit_r71_c208 bl[208] br[208] wl[71] vdd gnd cell_6t
Xbit_r72_c208 bl[208] br[208] wl[72] vdd gnd cell_6t
Xbit_r73_c208 bl[208] br[208] wl[73] vdd gnd cell_6t
Xbit_r74_c208 bl[208] br[208] wl[74] vdd gnd cell_6t
Xbit_r75_c208 bl[208] br[208] wl[75] vdd gnd cell_6t
Xbit_r76_c208 bl[208] br[208] wl[76] vdd gnd cell_6t
Xbit_r77_c208 bl[208] br[208] wl[77] vdd gnd cell_6t
Xbit_r78_c208 bl[208] br[208] wl[78] vdd gnd cell_6t
Xbit_r79_c208 bl[208] br[208] wl[79] vdd gnd cell_6t
Xbit_r80_c208 bl[208] br[208] wl[80] vdd gnd cell_6t
Xbit_r81_c208 bl[208] br[208] wl[81] vdd gnd cell_6t
Xbit_r82_c208 bl[208] br[208] wl[82] vdd gnd cell_6t
Xbit_r83_c208 bl[208] br[208] wl[83] vdd gnd cell_6t
Xbit_r84_c208 bl[208] br[208] wl[84] vdd gnd cell_6t
Xbit_r85_c208 bl[208] br[208] wl[85] vdd gnd cell_6t
Xbit_r86_c208 bl[208] br[208] wl[86] vdd gnd cell_6t
Xbit_r87_c208 bl[208] br[208] wl[87] vdd gnd cell_6t
Xbit_r88_c208 bl[208] br[208] wl[88] vdd gnd cell_6t
Xbit_r89_c208 bl[208] br[208] wl[89] vdd gnd cell_6t
Xbit_r90_c208 bl[208] br[208] wl[90] vdd gnd cell_6t
Xbit_r91_c208 bl[208] br[208] wl[91] vdd gnd cell_6t
Xbit_r92_c208 bl[208] br[208] wl[92] vdd gnd cell_6t
Xbit_r93_c208 bl[208] br[208] wl[93] vdd gnd cell_6t
Xbit_r94_c208 bl[208] br[208] wl[94] vdd gnd cell_6t
Xbit_r95_c208 bl[208] br[208] wl[95] vdd gnd cell_6t
Xbit_r96_c208 bl[208] br[208] wl[96] vdd gnd cell_6t
Xbit_r97_c208 bl[208] br[208] wl[97] vdd gnd cell_6t
Xbit_r98_c208 bl[208] br[208] wl[98] vdd gnd cell_6t
Xbit_r99_c208 bl[208] br[208] wl[99] vdd gnd cell_6t
Xbit_r100_c208 bl[208] br[208] wl[100] vdd gnd cell_6t
Xbit_r101_c208 bl[208] br[208] wl[101] vdd gnd cell_6t
Xbit_r102_c208 bl[208] br[208] wl[102] vdd gnd cell_6t
Xbit_r103_c208 bl[208] br[208] wl[103] vdd gnd cell_6t
Xbit_r104_c208 bl[208] br[208] wl[104] vdd gnd cell_6t
Xbit_r105_c208 bl[208] br[208] wl[105] vdd gnd cell_6t
Xbit_r106_c208 bl[208] br[208] wl[106] vdd gnd cell_6t
Xbit_r107_c208 bl[208] br[208] wl[107] vdd gnd cell_6t
Xbit_r108_c208 bl[208] br[208] wl[108] vdd gnd cell_6t
Xbit_r109_c208 bl[208] br[208] wl[109] vdd gnd cell_6t
Xbit_r110_c208 bl[208] br[208] wl[110] vdd gnd cell_6t
Xbit_r111_c208 bl[208] br[208] wl[111] vdd gnd cell_6t
Xbit_r112_c208 bl[208] br[208] wl[112] vdd gnd cell_6t
Xbit_r113_c208 bl[208] br[208] wl[113] vdd gnd cell_6t
Xbit_r114_c208 bl[208] br[208] wl[114] vdd gnd cell_6t
Xbit_r115_c208 bl[208] br[208] wl[115] vdd gnd cell_6t
Xbit_r116_c208 bl[208] br[208] wl[116] vdd gnd cell_6t
Xbit_r117_c208 bl[208] br[208] wl[117] vdd gnd cell_6t
Xbit_r118_c208 bl[208] br[208] wl[118] vdd gnd cell_6t
Xbit_r119_c208 bl[208] br[208] wl[119] vdd gnd cell_6t
Xbit_r120_c208 bl[208] br[208] wl[120] vdd gnd cell_6t
Xbit_r121_c208 bl[208] br[208] wl[121] vdd gnd cell_6t
Xbit_r122_c208 bl[208] br[208] wl[122] vdd gnd cell_6t
Xbit_r123_c208 bl[208] br[208] wl[123] vdd gnd cell_6t
Xbit_r124_c208 bl[208] br[208] wl[124] vdd gnd cell_6t
Xbit_r125_c208 bl[208] br[208] wl[125] vdd gnd cell_6t
Xbit_r126_c208 bl[208] br[208] wl[126] vdd gnd cell_6t
Xbit_r127_c208 bl[208] br[208] wl[127] vdd gnd cell_6t
Xbit_r128_c208 bl[208] br[208] wl[128] vdd gnd cell_6t
Xbit_r129_c208 bl[208] br[208] wl[129] vdd gnd cell_6t
Xbit_r130_c208 bl[208] br[208] wl[130] vdd gnd cell_6t
Xbit_r131_c208 bl[208] br[208] wl[131] vdd gnd cell_6t
Xbit_r132_c208 bl[208] br[208] wl[132] vdd gnd cell_6t
Xbit_r133_c208 bl[208] br[208] wl[133] vdd gnd cell_6t
Xbit_r134_c208 bl[208] br[208] wl[134] vdd gnd cell_6t
Xbit_r135_c208 bl[208] br[208] wl[135] vdd gnd cell_6t
Xbit_r136_c208 bl[208] br[208] wl[136] vdd gnd cell_6t
Xbit_r137_c208 bl[208] br[208] wl[137] vdd gnd cell_6t
Xbit_r138_c208 bl[208] br[208] wl[138] vdd gnd cell_6t
Xbit_r139_c208 bl[208] br[208] wl[139] vdd gnd cell_6t
Xbit_r140_c208 bl[208] br[208] wl[140] vdd gnd cell_6t
Xbit_r141_c208 bl[208] br[208] wl[141] vdd gnd cell_6t
Xbit_r142_c208 bl[208] br[208] wl[142] vdd gnd cell_6t
Xbit_r143_c208 bl[208] br[208] wl[143] vdd gnd cell_6t
Xbit_r144_c208 bl[208] br[208] wl[144] vdd gnd cell_6t
Xbit_r145_c208 bl[208] br[208] wl[145] vdd gnd cell_6t
Xbit_r146_c208 bl[208] br[208] wl[146] vdd gnd cell_6t
Xbit_r147_c208 bl[208] br[208] wl[147] vdd gnd cell_6t
Xbit_r148_c208 bl[208] br[208] wl[148] vdd gnd cell_6t
Xbit_r149_c208 bl[208] br[208] wl[149] vdd gnd cell_6t
Xbit_r150_c208 bl[208] br[208] wl[150] vdd gnd cell_6t
Xbit_r151_c208 bl[208] br[208] wl[151] vdd gnd cell_6t
Xbit_r152_c208 bl[208] br[208] wl[152] vdd gnd cell_6t
Xbit_r153_c208 bl[208] br[208] wl[153] vdd gnd cell_6t
Xbit_r154_c208 bl[208] br[208] wl[154] vdd gnd cell_6t
Xbit_r155_c208 bl[208] br[208] wl[155] vdd gnd cell_6t
Xbit_r156_c208 bl[208] br[208] wl[156] vdd gnd cell_6t
Xbit_r157_c208 bl[208] br[208] wl[157] vdd gnd cell_6t
Xbit_r158_c208 bl[208] br[208] wl[158] vdd gnd cell_6t
Xbit_r159_c208 bl[208] br[208] wl[159] vdd gnd cell_6t
Xbit_r160_c208 bl[208] br[208] wl[160] vdd gnd cell_6t
Xbit_r161_c208 bl[208] br[208] wl[161] vdd gnd cell_6t
Xbit_r162_c208 bl[208] br[208] wl[162] vdd gnd cell_6t
Xbit_r163_c208 bl[208] br[208] wl[163] vdd gnd cell_6t
Xbit_r164_c208 bl[208] br[208] wl[164] vdd gnd cell_6t
Xbit_r165_c208 bl[208] br[208] wl[165] vdd gnd cell_6t
Xbit_r166_c208 bl[208] br[208] wl[166] vdd gnd cell_6t
Xbit_r167_c208 bl[208] br[208] wl[167] vdd gnd cell_6t
Xbit_r168_c208 bl[208] br[208] wl[168] vdd gnd cell_6t
Xbit_r169_c208 bl[208] br[208] wl[169] vdd gnd cell_6t
Xbit_r170_c208 bl[208] br[208] wl[170] vdd gnd cell_6t
Xbit_r171_c208 bl[208] br[208] wl[171] vdd gnd cell_6t
Xbit_r172_c208 bl[208] br[208] wl[172] vdd gnd cell_6t
Xbit_r173_c208 bl[208] br[208] wl[173] vdd gnd cell_6t
Xbit_r174_c208 bl[208] br[208] wl[174] vdd gnd cell_6t
Xbit_r175_c208 bl[208] br[208] wl[175] vdd gnd cell_6t
Xbit_r176_c208 bl[208] br[208] wl[176] vdd gnd cell_6t
Xbit_r177_c208 bl[208] br[208] wl[177] vdd gnd cell_6t
Xbit_r178_c208 bl[208] br[208] wl[178] vdd gnd cell_6t
Xbit_r179_c208 bl[208] br[208] wl[179] vdd gnd cell_6t
Xbit_r180_c208 bl[208] br[208] wl[180] vdd gnd cell_6t
Xbit_r181_c208 bl[208] br[208] wl[181] vdd gnd cell_6t
Xbit_r182_c208 bl[208] br[208] wl[182] vdd gnd cell_6t
Xbit_r183_c208 bl[208] br[208] wl[183] vdd gnd cell_6t
Xbit_r184_c208 bl[208] br[208] wl[184] vdd gnd cell_6t
Xbit_r185_c208 bl[208] br[208] wl[185] vdd gnd cell_6t
Xbit_r186_c208 bl[208] br[208] wl[186] vdd gnd cell_6t
Xbit_r187_c208 bl[208] br[208] wl[187] vdd gnd cell_6t
Xbit_r188_c208 bl[208] br[208] wl[188] vdd gnd cell_6t
Xbit_r189_c208 bl[208] br[208] wl[189] vdd gnd cell_6t
Xbit_r190_c208 bl[208] br[208] wl[190] vdd gnd cell_6t
Xbit_r191_c208 bl[208] br[208] wl[191] vdd gnd cell_6t
Xbit_r192_c208 bl[208] br[208] wl[192] vdd gnd cell_6t
Xbit_r193_c208 bl[208] br[208] wl[193] vdd gnd cell_6t
Xbit_r194_c208 bl[208] br[208] wl[194] vdd gnd cell_6t
Xbit_r195_c208 bl[208] br[208] wl[195] vdd gnd cell_6t
Xbit_r196_c208 bl[208] br[208] wl[196] vdd gnd cell_6t
Xbit_r197_c208 bl[208] br[208] wl[197] vdd gnd cell_6t
Xbit_r198_c208 bl[208] br[208] wl[198] vdd gnd cell_6t
Xbit_r199_c208 bl[208] br[208] wl[199] vdd gnd cell_6t
Xbit_r200_c208 bl[208] br[208] wl[200] vdd gnd cell_6t
Xbit_r201_c208 bl[208] br[208] wl[201] vdd gnd cell_6t
Xbit_r202_c208 bl[208] br[208] wl[202] vdd gnd cell_6t
Xbit_r203_c208 bl[208] br[208] wl[203] vdd gnd cell_6t
Xbit_r204_c208 bl[208] br[208] wl[204] vdd gnd cell_6t
Xbit_r205_c208 bl[208] br[208] wl[205] vdd gnd cell_6t
Xbit_r206_c208 bl[208] br[208] wl[206] vdd gnd cell_6t
Xbit_r207_c208 bl[208] br[208] wl[207] vdd gnd cell_6t
Xbit_r208_c208 bl[208] br[208] wl[208] vdd gnd cell_6t
Xbit_r209_c208 bl[208] br[208] wl[209] vdd gnd cell_6t
Xbit_r210_c208 bl[208] br[208] wl[210] vdd gnd cell_6t
Xbit_r211_c208 bl[208] br[208] wl[211] vdd gnd cell_6t
Xbit_r212_c208 bl[208] br[208] wl[212] vdd gnd cell_6t
Xbit_r213_c208 bl[208] br[208] wl[213] vdd gnd cell_6t
Xbit_r214_c208 bl[208] br[208] wl[214] vdd gnd cell_6t
Xbit_r215_c208 bl[208] br[208] wl[215] vdd gnd cell_6t
Xbit_r216_c208 bl[208] br[208] wl[216] vdd gnd cell_6t
Xbit_r217_c208 bl[208] br[208] wl[217] vdd gnd cell_6t
Xbit_r218_c208 bl[208] br[208] wl[218] vdd gnd cell_6t
Xbit_r219_c208 bl[208] br[208] wl[219] vdd gnd cell_6t
Xbit_r220_c208 bl[208] br[208] wl[220] vdd gnd cell_6t
Xbit_r221_c208 bl[208] br[208] wl[221] vdd gnd cell_6t
Xbit_r222_c208 bl[208] br[208] wl[222] vdd gnd cell_6t
Xbit_r223_c208 bl[208] br[208] wl[223] vdd gnd cell_6t
Xbit_r224_c208 bl[208] br[208] wl[224] vdd gnd cell_6t
Xbit_r225_c208 bl[208] br[208] wl[225] vdd gnd cell_6t
Xbit_r226_c208 bl[208] br[208] wl[226] vdd gnd cell_6t
Xbit_r227_c208 bl[208] br[208] wl[227] vdd gnd cell_6t
Xbit_r228_c208 bl[208] br[208] wl[228] vdd gnd cell_6t
Xbit_r229_c208 bl[208] br[208] wl[229] vdd gnd cell_6t
Xbit_r230_c208 bl[208] br[208] wl[230] vdd gnd cell_6t
Xbit_r231_c208 bl[208] br[208] wl[231] vdd gnd cell_6t
Xbit_r232_c208 bl[208] br[208] wl[232] vdd gnd cell_6t
Xbit_r233_c208 bl[208] br[208] wl[233] vdd gnd cell_6t
Xbit_r234_c208 bl[208] br[208] wl[234] vdd gnd cell_6t
Xbit_r235_c208 bl[208] br[208] wl[235] vdd gnd cell_6t
Xbit_r236_c208 bl[208] br[208] wl[236] vdd gnd cell_6t
Xbit_r237_c208 bl[208] br[208] wl[237] vdd gnd cell_6t
Xbit_r238_c208 bl[208] br[208] wl[238] vdd gnd cell_6t
Xbit_r239_c208 bl[208] br[208] wl[239] vdd gnd cell_6t
Xbit_r240_c208 bl[208] br[208] wl[240] vdd gnd cell_6t
Xbit_r241_c208 bl[208] br[208] wl[241] vdd gnd cell_6t
Xbit_r242_c208 bl[208] br[208] wl[242] vdd gnd cell_6t
Xbit_r243_c208 bl[208] br[208] wl[243] vdd gnd cell_6t
Xbit_r244_c208 bl[208] br[208] wl[244] vdd gnd cell_6t
Xbit_r245_c208 bl[208] br[208] wl[245] vdd gnd cell_6t
Xbit_r246_c208 bl[208] br[208] wl[246] vdd gnd cell_6t
Xbit_r247_c208 bl[208] br[208] wl[247] vdd gnd cell_6t
Xbit_r248_c208 bl[208] br[208] wl[248] vdd gnd cell_6t
Xbit_r249_c208 bl[208] br[208] wl[249] vdd gnd cell_6t
Xbit_r250_c208 bl[208] br[208] wl[250] vdd gnd cell_6t
Xbit_r251_c208 bl[208] br[208] wl[251] vdd gnd cell_6t
Xbit_r252_c208 bl[208] br[208] wl[252] vdd gnd cell_6t
Xbit_r253_c208 bl[208] br[208] wl[253] vdd gnd cell_6t
Xbit_r254_c208 bl[208] br[208] wl[254] vdd gnd cell_6t
Xbit_r255_c208 bl[208] br[208] wl[255] vdd gnd cell_6t
Xbit_r0_c209 bl[209] br[209] wl[0] vdd gnd cell_6t
Xbit_r1_c209 bl[209] br[209] wl[1] vdd gnd cell_6t
Xbit_r2_c209 bl[209] br[209] wl[2] vdd gnd cell_6t
Xbit_r3_c209 bl[209] br[209] wl[3] vdd gnd cell_6t
Xbit_r4_c209 bl[209] br[209] wl[4] vdd gnd cell_6t
Xbit_r5_c209 bl[209] br[209] wl[5] vdd gnd cell_6t
Xbit_r6_c209 bl[209] br[209] wl[6] vdd gnd cell_6t
Xbit_r7_c209 bl[209] br[209] wl[7] vdd gnd cell_6t
Xbit_r8_c209 bl[209] br[209] wl[8] vdd gnd cell_6t
Xbit_r9_c209 bl[209] br[209] wl[9] vdd gnd cell_6t
Xbit_r10_c209 bl[209] br[209] wl[10] vdd gnd cell_6t
Xbit_r11_c209 bl[209] br[209] wl[11] vdd gnd cell_6t
Xbit_r12_c209 bl[209] br[209] wl[12] vdd gnd cell_6t
Xbit_r13_c209 bl[209] br[209] wl[13] vdd gnd cell_6t
Xbit_r14_c209 bl[209] br[209] wl[14] vdd gnd cell_6t
Xbit_r15_c209 bl[209] br[209] wl[15] vdd gnd cell_6t
Xbit_r16_c209 bl[209] br[209] wl[16] vdd gnd cell_6t
Xbit_r17_c209 bl[209] br[209] wl[17] vdd gnd cell_6t
Xbit_r18_c209 bl[209] br[209] wl[18] vdd gnd cell_6t
Xbit_r19_c209 bl[209] br[209] wl[19] vdd gnd cell_6t
Xbit_r20_c209 bl[209] br[209] wl[20] vdd gnd cell_6t
Xbit_r21_c209 bl[209] br[209] wl[21] vdd gnd cell_6t
Xbit_r22_c209 bl[209] br[209] wl[22] vdd gnd cell_6t
Xbit_r23_c209 bl[209] br[209] wl[23] vdd gnd cell_6t
Xbit_r24_c209 bl[209] br[209] wl[24] vdd gnd cell_6t
Xbit_r25_c209 bl[209] br[209] wl[25] vdd gnd cell_6t
Xbit_r26_c209 bl[209] br[209] wl[26] vdd gnd cell_6t
Xbit_r27_c209 bl[209] br[209] wl[27] vdd gnd cell_6t
Xbit_r28_c209 bl[209] br[209] wl[28] vdd gnd cell_6t
Xbit_r29_c209 bl[209] br[209] wl[29] vdd gnd cell_6t
Xbit_r30_c209 bl[209] br[209] wl[30] vdd gnd cell_6t
Xbit_r31_c209 bl[209] br[209] wl[31] vdd gnd cell_6t
Xbit_r32_c209 bl[209] br[209] wl[32] vdd gnd cell_6t
Xbit_r33_c209 bl[209] br[209] wl[33] vdd gnd cell_6t
Xbit_r34_c209 bl[209] br[209] wl[34] vdd gnd cell_6t
Xbit_r35_c209 bl[209] br[209] wl[35] vdd gnd cell_6t
Xbit_r36_c209 bl[209] br[209] wl[36] vdd gnd cell_6t
Xbit_r37_c209 bl[209] br[209] wl[37] vdd gnd cell_6t
Xbit_r38_c209 bl[209] br[209] wl[38] vdd gnd cell_6t
Xbit_r39_c209 bl[209] br[209] wl[39] vdd gnd cell_6t
Xbit_r40_c209 bl[209] br[209] wl[40] vdd gnd cell_6t
Xbit_r41_c209 bl[209] br[209] wl[41] vdd gnd cell_6t
Xbit_r42_c209 bl[209] br[209] wl[42] vdd gnd cell_6t
Xbit_r43_c209 bl[209] br[209] wl[43] vdd gnd cell_6t
Xbit_r44_c209 bl[209] br[209] wl[44] vdd gnd cell_6t
Xbit_r45_c209 bl[209] br[209] wl[45] vdd gnd cell_6t
Xbit_r46_c209 bl[209] br[209] wl[46] vdd gnd cell_6t
Xbit_r47_c209 bl[209] br[209] wl[47] vdd gnd cell_6t
Xbit_r48_c209 bl[209] br[209] wl[48] vdd gnd cell_6t
Xbit_r49_c209 bl[209] br[209] wl[49] vdd gnd cell_6t
Xbit_r50_c209 bl[209] br[209] wl[50] vdd gnd cell_6t
Xbit_r51_c209 bl[209] br[209] wl[51] vdd gnd cell_6t
Xbit_r52_c209 bl[209] br[209] wl[52] vdd gnd cell_6t
Xbit_r53_c209 bl[209] br[209] wl[53] vdd gnd cell_6t
Xbit_r54_c209 bl[209] br[209] wl[54] vdd gnd cell_6t
Xbit_r55_c209 bl[209] br[209] wl[55] vdd gnd cell_6t
Xbit_r56_c209 bl[209] br[209] wl[56] vdd gnd cell_6t
Xbit_r57_c209 bl[209] br[209] wl[57] vdd gnd cell_6t
Xbit_r58_c209 bl[209] br[209] wl[58] vdd gnd cell_6t
Xbit_r59_c209 bl[209] br[209] wl[59] vdd gnd cell_6t
Xbit_r60_c209 bl[209] br[209] wl[60] vdd gnd cell_6t
Xbit_r61_c209 bl[209] br[209] wl[61] vdd gnd cell_6t
Xbit_r62_c209 bl[209] br[209] wl[62] vdd gnd cell_6t
Xbit_r63_c209 bl[209] br[209] wl[63] vdd gnd cell_6t
Xbit_r64_c209 bl[209] br[209] wl[64] vdd gnd cell_6t
Xbit_r65_c209 bl[209] br[209] wl[65] vdd gnd cell_6t
Xbit_r66_c209 bl[209] br[209] wl[66] vdd gnd cell_6t
Xbit_r67_c209 bl[209] br[209] wl[67] vdd gnd cell_6t
Xbit_r68_c209 bl[209] br[209] wl[68] vdd gnd cell_6t
Xbit_r69_c209 bl[209] br[209] wl[69] vdd gnd cell_6t
Xbit_r70_c209 bl[209] br[209] wl[70] vdd gnd cell_6t
Xbit_r71_c209 bl[209] br[209] wl[71] vdd gnd cell_6t
Xbit_r72_c209 bl[209] br[209] wl[72] vdd gnd cell_6t
Xbit_r73_c209 bl[209] br[209] wl[73] vdd gnd cell_6t
Xbit_r74_c209 bl[209] br[209] wl[74] vdd gnd cell_6t
Xbit_r75_c209 bl[209] br[209] wl[75] vdd gnd cell_6t
Xbit_r76_c209 bl[209] br[209] wl[76] vdd gnd cell_6t
Xbit_r77_c209 bl[209] br[209] wl[77] vdd gnd cell_6t
Xbit_r78_c209 bl[209] br[209] wl[78] vdd gnd cell_6t
Xbit_r79_c209 bl[209] br[209] wl[79] vdd gnd cell_6t
Xbit_r80_c209 bl[209] br[209] wl[80] vdd gnd cell_6t
Xbit_r81_c209 bl[209] br[209] wl[81] vdd gnd cell_6t
Xbit_r82_c209 bl[209] br[209] wl[82] vdd gnd cell_6t
Xbit_r83_c209 bl[209] br[209] wl[83] vdd gnd cell_6t
Xbit_r84_c209 bl[209] br[209] wl[84] vdd gnd cell_6t
Xbit_r85_c209 bl[209] br[209] wl[85] vdd gnd cell_6t
Xbit_r86_c209 bl[209] br[209] wl[86] vdd gnd cell_6t
Xbit_r87_c209 bl[209] br[209] wl[87] vdd gnd cell_6t
Xbit_r88_c209 bl[209] br[209] wl[88] vdd gnd cell_6t
Xbit_r89_c209 bl[209] br[209] wl[89] vdd gnd cell_6t
Xbit_r90_c209 bl[209] br[209] wl[90] vdd gnd cell_6t
Xbit_r91_c209 bl[209] br[209] wl[91] vdd gnd cell_6t
Xbit_r92_c209 bl[209] br[209] wl[92] vdd gnd cell_6t
Xbit_r93_c209 bl[209] br[209] wl[93] vdd gnd cell_6t
Xbit_r94_c209 bl[209] br[209] wl[94] vdd gnd cell_6t
Xbit_r95_c209 bl[209] br[209] wl[95] vdd gnd cell_6t
Xbit_r96_c209 bl[209] br[209] wl[96] vdd gnd cell_6t
Xbit_r97_c209 bl[209] br[209] wl[97] vdd gnd cell_6t
Xbit_r98_c209 bl[209] br[209] wl[98] vdd gnd cell_6t
Xbit_r99_c209 bl[209] br[209] wl[99] vdd gnd cell_6t
Xbit_r100_c209 bl[209] br[209] wl[100] vdd gnd cell_6t
Xbit_r101_c209 bl[209] br[209] wl[101] vdd gnd cell_6t
Xbit_r102_c209 bl[209] br[209] wl[102] vdd gnd cell_6t
Xbit_r103_c209 bl[209] br[209] wl[103] vdd gnd cell_6t
Xbit_r104_c209 bl[209] br[209] wl[104] vdd gnd cell_6t
Xbit_r105_c209 bl[209] br[209] wl[105] vdd gnd cell_6t
Xbit_r106_c209 bl[209] br[209] wl[106] vdd gnd cell_6t
Xbit_r107_c209 bl[209] br[209] wl[107] vdd gnd cell_6t
Xbit_r108_c209 bl[209] br[209] wl[108] vdd gnd cell_6t
Xbit_r109_c209 bl[209] br[209] wl[109] vdd gnd cell_6t
Xbit_r110_c209 bl[209] br[209] wl[110] vdd gnd cell_6t
Xbit_r111_c209 bl[209] br[209] wl[111] vdd gnd cell_6t
Xbit_r112_c209 bl[209] br[209] wl[112] vdd gnd cell_6t
Xbit_r113_c209 bl[209] br[209] wl[113] vdd gnd cell_6t
Xbit_r114_c209 bl[209] br[209] wl[114] vdd gnd cell_6t
Xbit_r115_c209 bl[209] br[209] wl[115] vdd gnd cell_6t
Xbit_r116_c209 bl[209] br[209] wl[116] vdd gnd cell_6t
Xbit_r117_c209 bl[209] br[209] wl[117] vdd gnd cell_6t
Xbit_r118_c209 bl[209] br[209] wl[118] vdd gnd cell_6t
Xbit_r119_c209 bl[209] br[209] wl[119] vdd gnd cell_6t
Xbit_r120_c209 bl[209] br[209] wl[120] vdd gnd cell_6t
Xbit_r121_c209 bl[209] br[209] wl[121] vdd gnd cell_6t
Xbit_r122_c209 bl[209] br[209] wl[122] vdd gnd cell_6t
Xbit_r123_c209 bl[209] br[209] wl[123] vdd gnd cell_6t
Xbit_r124_c209 bl[209] br[209] wl[124] vdd gnd cell_6t
Xbit_r125_c209 bl[209] br[209] wl[125] vdd gnd cell_6t
Xbit_r126_c209 bl[209] br[209] wl[126] vdd gnd cell_6t
Xbit_r127_c209 bl[209] br[209] wl[127] vdd gnd cell_6t
Xbit_r128_c209 bl[209] br[209] wl[128] vdd gnd cell_6t
Xbit_r129_c209 bl[209] br[209] wl[129] vdd gnd cell_6t
Xbit_r130_c209 bl[209] br[209] wl[130] vdd gnd cell_6t
Xbit_r131_c209 bl[209] br[209] wl[131] vdd gnd cell_6t
Xbit_r132_c209 bl[209] br[209] wl[132] vdd gnd cell_6t
Xbit_r133_c209 bl[209] br[209] wl[133] vdd gnd cell_6t
Xbit_r134_c209 bl[209] br[209] wl[134] vdd gnd cell_6t
Xbit_r135_c209 bl[209] br[209] wl[135] vdd gnd cell_6t
Xbit_r136_c209 bl[209] br[209] wl[136] vdd gnd cell_6t
Xbit_r137_c209 bl[209] br[209] wl[137] vdd gnd cell_6t
Xbit_r138_c209 bl[209] br[209] wl[138] vdd gnd cell_6t
Xbit_r139_c209 bl[209] br[209] wl[139] vdd gnd cell_6t
Xbit_r140_c209 bl[209] br[209] wl[140] vdd gnd cell_6t
Xbit_r141_c209 bl[209] br[209] wl[141] vdd gnd cell_6t
Xbit_r142_c209 bl[209] br[209] wl[142] vdd gnd cell_6t
Xbit_r143_c209 bl[209] br[209] wl[143] vdd gnd cell_6t
Xbit_r144_c209 bl[209] br[209] wl[144] vdd gnd cell_6t
Xbit_r145_c209 bl[209] br[209] wl[145] vdd gnd cell_6t
Xbit_r146_c209 bl[209] br[209] wl[146] vdd gnd cell_6t
Xbit_r147_c209 bl[209] br[209] wl[147] vdd gnd cell_6t
Xbit_r148_c209 bl[209] br[209] wl[148] vdd gnd cell_6t
Xbit_r149_c209 bl[209] br[209] wl[149] vdd gnd cell_6t
Xbit_r150_c209 bl[209] br[209] wl[150] vdd gnd cell_6t
Xbit_r151_c209 bl[209] br[209] wl[151] vdd gnd cell_6t
Xbit_r152_c209 bl[209] br[209] wl[152] vdd gnd cell_6t
Xbit_r153_c209 bl[209] br[209] wl[153] vdd gnd cell_6t
Xbit_r154_c209 bl[209] br[209] wl[154] vdd gnd cell_6t
Xbit_r155_c209 bl[209] br[209] wl[155] vdd gnd cell_6t
Xbit_r156_c209 bl[209] br[209] wl[156] vdd gnd cell_6t
Xbit_r157_c209 bl[209] br[209] wl[157] vdd gnd cell_6t
Xbit_r158_c209 bl[209] br[209] wl[158] vdd gnd cell_6t
Xbit_r159_c209 bl[209] br[209] wl[159] vdd gnd cell_6t
Xbit_r160_c209 bl[209] br[209] wl[160] vdd gnd cell_6t
Xbit_r161_c209 bl[209] br[209] wl[161] vdd gnd cell_6t
Xbit_r162_c209 bl[209] br[209] wl[162] vdd gnd cell_6t
Xbit_r163_c209 bl[209] br[209] wl[163] vdd gnd cell_6t
Xbit_r164_c209 bl[209] br[209] wl[164] vdd gnd cell_6t
Xbit_r165_c209 bl[209] br[209] wl[165] vdd gnd cell_6t
Xbit_r166_c209 bl[209] br[209] wl[166] vdd gnd cell_6t
Xbit_r167_c209 bl[209] br[209] wl[167] vdd gnd cell_6t
Xbit_r168_c209 bl[209] br[209] wl[168] vdd gnd cell_6t
Xbit_r169_c209 bl[209] br[209] wl[169] vdd gnd cell_6t
Xbit_r170_c209 bl[209] br[209] wl[170] vdd gnd cell_6t
Xbit_r171_c209 bl[209] br[209] wl[171] vdd gnd cell_6t
Xbit_r172_c209 bl[209] br[209] wl[172] vdd gnd cell_6t
Xbit_r173_c209 bl[209] br[209] wl[173] vdd gnd cell_6t
Xbit_r174_c209 bl[209] br[209] wl[174] vdd gnd cell_6t
Xbit_r175_c209 bl[209] br[209] wl[175] vdd gnd cell_6t
Xbit_r176_c209 bl[209] br[209] wl[176] vdd gnd cell_6t
Xbit_r177_c209 bl[209] br[209] wl[177] vdd gnd cell_6t
Xbit_r178_c209 bl[209] br[209] wl[178] vdd gnd cell_6t
Xbit_r179_c209 bl[209] br[209] wl[179] vdd gnd cell_6t
Xbit_r180_c209 bl[209] br[209] wl[180] vdd gnd cell_6t
Xbit_r181_c209 bl[209] br[209] wl[181] vdd gnd cell_6t
Xbit_r182_c209 bl[209] br[209] wl[182] vdd gnd cell_6t
Xbit_r183_c209 bl[209] br[209] wl[183] vdd gnd cell_6t
Xbit_r184_c209 bl[209] br[209] wl[184] vdd gnd cell_6t
Xbit_r185_c209 bl[209] br[209] wl[185] vdd gnd cell_6t
Xbit_r186_c209 bl[209] br[209] wl[186] vdd gnd cell_6t
Xbit_r187_c209 bl[209] br[209] wl[187] vdd gnd cell_6t
Xbit_r188_c209 bl[209] br[209] wl[188] vdd gnd cell_6t
Xbit_r189_c209 bl[209] br[209] wl[189] vdd gnd cell_6t
Xbit_r190_c209 bl[209] br[209] wl[190] vdd gnd cell_6t
Xbit_r191_c209 bl[209] br[209] wl[191] vdd gnd cell_6t
Xbit_r192_c209 bl[209] br[209] wl[192] vdd gnd cell_6t
Xbit_r193_c209 bl[209] br[209] wl[193] vdd gnd cell_6t
Xbit_r194_c209 bl[209] br[209] wl[194] vdd gnd cell_6t
Xbit_r195_c209 bl[209] br[209] wl[195] vdd gnd cell_6t
Xbit_r196_c209 bl[209] br[209] wl[196] vdd gnd cell_6t
Xbit_r197_c209 bl[209] br[209] wl[197] vdd gnd cell_6t
Xbit_r198_c209 bl[209] br[209] wl[198] vdd gnd cell_6t
Xbit_r199_c209 bl[209] br[209] wl[199] vdd gnd cell_6t
Xbit_r200_c209 bl[209] br[209] wl[200] vdd gnd cell_6t
Xbit_r201_c209 bl[209] br[209] wl[201] vdd gnd cell_6t
Xbit_r202_c209 bl[209] br[209] wl[202] vdd gnd cell_6t
Xbit_r203_c209 bl[209] br[209] wl[203] vdd gnd cell_6t
Xbit_r204_c209 bl[209] br[209] wl[204] vdd gnd cell_6t
Xbit_r205_c209 bl[209] br[209] wl[205] vdd gnd cell_6t
Xbit_r206_c209 bl[209] br[209] wl[206] vdd gnd cell_6t
Xbit_r207_c209 bl[209] br[209] wl[207] vdd gnd cell_6t
Xbit_r208_c209 bl[209] br[209] wl[208] vdd gnd cell_6t
Xbit_r209_c209 bl[209] br[209] wl[209] vdd gnd cell_6t
Xbit_r210_c209 bl[209] br[209] wl[210] vdd gnd cell_6t
Xbit_r211_c209 bl[209] br[209] wl[211] vdd gnd cell_6t
Xbit_r212_c209 bl[209] br[209] wl[212] vdd gnd cell_6t
Xbit_r213_c209 bl[209] br[209] wl[213] vdd gnd cell_6t
Xbit_r214_c209 bl[209] br[209] wl[214] vdd gnd cell_6t
Xbit_r215_c209 bl[209] br[209] wl[215] vdd gnd cell_6t
Xbit_r216_c209 bl[209] br[209] wl[216] vdd gnd cell_6t
Xbit_r217_c209 bl[209] br[209] wl[217] vdd gnd cell_6t
Xbit_r218_c209 bl[209] br[209] wl[218] vdd gnd cell_6t
Xbit_r219_c209 bl[209] br[209] wl[219] vdd gnd cell_6t
Xbit_r220_c209 bl[209] br[209] wl[220] vdd gnd cell_6t
Xbit_r221_c209 bl[209] br[209] wl[221] vdd gnd cell_6t
Xbit_r222_c209 bl[209] br[209] wl[222] vdd gnd cell_6t
Xbit_r223_c209 bl[209] br[209] wl[223] vdd gnd cell_6t
Xbit_r224_c209 bl[209] br[209] wl[224] vdd gnd cell_6t
Xbit_r225_c209 bl[209] br[209] wl[225] vdd gnd cell_6t
Xbit_r226_c209 bl[209] br[209] wl[226] vdd gnd cell_6t
Xbit_r227_c209 bl[209] br[209] wl[227] vdd gnd cell_6t
Xbit_r228_c209 bl[209] br[209] wl[228] vdd gnd cell_6t
Xbit_r229_c209 bl[209] br[209] wl[229] vdd gnd cell_6t
Xbit_r230_c209 bl[209] br[209] wl[230] vdd gnd cell_6t
Xbit_r231_c209 bl[209] br[209] wl[231] vdd gnd cell_6t
Xbit_r232_c209 bl[209] br[209] wl[232] vdd gnd cell_6t
Xbit_r233_c209 bl[209] br[209] wl[233] vdd gnd cell_6t
Xbit_r234_c209 bl[209] br[209] wl[234] vdd gnd cell_6t
Xbit_r235_c209 bl[209] br[209] wl[235] vdd gnd cell_6t
Xbit_r236_c209 bl[209] br[209] wl[236] vdd gnd cell_6t
Xbit_r237_c209 bl[209] br[209] wl[237] vdd gnd cell_6t
Xbit_r238_c209 bl[209] br[209] wl[238] vdd gnd cell_6t
Xbit_r239_c209 bl[209] br[209] wl[239] vdd gnd cell_6t
Xbit_r240_c209 bl[209] br[209] wl[240] vdd gnd cell_6t
Xbit_r241_c209 bl[209] br[209] wl[241] vdd gnd cell_6t
Xbit_r242_c209 bl[209] br[209] wl[242] vdd gnd cell_6t
Xbit_r243_c209 bl[209] br[209] wl[243] vdd gnd cell_6t
Xbit_r244_c209 bl[209] br[209] wl[244] vdd gnd cell_6t
Xbit_r245_c209 bl[209] br[209] wl[245] vdd gnd cell_6t
Xbit_r246_c209 bl[209] br[209] wl[246] vdd gnd cell_6t
Xbit_r247_c209 bl[209] br[209] wl[247] vdd gnd cell_6t
Xbit_r248_c209 bl[209] br[209] wl[248] vdd gnd cell_6t
Xbit_r249_c209 bl[209] br[209] wl[249] vdd gnd cell_6t
Xbit_r250_c209 bl[209] br[209] wl[250] vdd gnd cell_6t
Xbit_r251_c209 bl[209] br[209] wl[251] vdd gnd cell_6t
Xbit_r252_c209 bl[209] br[209] wl[252] vdd gnd cell_6t
Xbit_r253_c209 bl[209] br[209] wl[253] vdd gnd cell_6t
Xbit_r254_c209 bl[209] br[209] wl[254] vdd gnd cell_6t
Xbit_r255_c209 bl[209] br[209] wl[255] vdd gnd cell_6t
Xbit_r0_c210 bl[210] br[210] wl[0] vdd gnd cell_6t
Xbit_r1_c210 bl[210] br[210] wl[1] vdd gnd cell_6t
Xbit_r2_c210 bl[210] br[210] wl[2] vdd gnd cell_6t
Xbit_r3_c210 bl[210] br[210] wl[3] vdd gnd cell_6t
Xbit_r4_c210 bl[210] br[210] wl[4] vdd gnd cell_6t
Xbit_r5_c210 bl[210] br[210] wl[5] vdd gnd cell_6t
Xbit_r6_c210 bl[210] br[210] wl[6] vdd gnd cell_6t
Xbit_r7_c210 bl[210] br[210] wl[7] vdd gnd cell_6t
Xbit_r8_c210 bl[210] br[210] wl[8] vdd gnd cell_6t
Xbit_r9_c210 bl[210] br[210] wl[9] vdd gnd cell_6t
Xbit_r10_c210 bl[210] br[210] wl[10] vdd gnd cell_6t
Xbit_r11_c210 bl[210] br[210] wl[11] vdd gnd cell_6t
Xbit_r12_c210 bl[210] br[210] wl[12] vdd gnd cell_6t
Xbit_r13_c210 bl[210] br[210] wl[13] vdd gnd cell_6t
Xbit_r14_c210 bl[210] br[210] wl[14] vdd gnd cell_6t
Xbit_r15_c210 bl[210] br[210] wl[15] vdd gnd cell_6t
Xbit_r16_c210 bl[210] br[210] wl[16] vdd gnd cell_6t
Xbit_r17_c210 bl[210] br[210] wl[17] vdd gnd cell_6t
Xbit_r18_c210 bl[210] br[210] wl[18] vdd gnd cell_6t
Xbit_r19_c210 bl[210] br[210] wl[19] vdd gnd cell_6t
Xbit_r20_c210 bl[210] br[210] wl[20] vdd gnd cell_6t
Xbit_r21_c210 bl[210] br[210] wl[21] vdd gnd cell_6t
Xbit_r22_c210 bl[210] br[210] wl[22] vdd gnd cell_6t
Xbit_r23_c210 bl[210] br[210] wl[23] vdd gnd cell_6t
Xbit_r24_c210 bl[210] br[210] wl[24] vdd gnd cell_6t
Xbit_r25_c210 bl[210] br[210] wl[25] vdd gnd cell_6t
Xbit_r26_c210 bl[210] br[210] wl[26] vdd gnd cell_6t
Xbit_r27_c210 bl[210] br[210] wl[27] vdd gnd cell_6t
Xbit_r28_c210 bl[210] br[210] wl[28] vdd gnd cell_6t
Xbit_r29_c210 bl[210] br[210] wl[29] vdd gnd cell_6t
Xbit_r30_c210 bl[210] br[210] wl[30] vdd gnd cell_6t
Xbit_r31_c210 bl[210] br[210] wl[31] vdd gnd cell_6t
Xbit_r32_c210 bl[210] br[210] wl[32] vdd gnd cell_6t
Xbit_r33_c210 bl[210] br[210] wl[33] vdd gnd cell_6t
Xbit_r34_c210 bl[210] br[210] wl[34] vdd gnd cell_6t
Xbit_r35_c210 bl[210] br[210] wl[35] vdd gnd cell_6t
Xbit_r36_c210 bl[210] br[210] wl[36] vdd gnd cell_6t
Xbit_r37_c210 bl[210] br[210] wl[37] vdd gnd cell_6t
Xbit_r38_c210 bl[210] br[210] wl[38] vdd gnd cell_6t
Xbit_r39_c210 bl[210] br[210] wl[39] vdd gnd cell_6t
Xbit_r40_c210 bl[210] br[210] wl[40] vdd gnd cell_6t
Xbit_r41_c210 bl[210] br[210] wl[41] vdd gnd cell_6t
Xbit_r42_c210 bl[210] br[210] wl[42] vdd gnd cell_6t
Xbit_r43_c210 bl[210] br[210] wl[43] vdd gnd cell_6t
Xbit_r44_c210 bl[210] br[210] wl[44] vdd gnd cell_6t
Xbit_r45_c210 bl[210] br[210] wl[45] vdd gnd cell_6t
Xbit_r46_c210 bl[210] br[210] wl[46] vdd gnd cell_6t
Xbit_r47_c210 bl[210] br[210] wl[47] vdd gnd cell_6t
Xbit_r48_c210 bl[210] br[210] wl[48] vdd gnd cell_6t
Xbit_r49_c210 bl[210] br[210] wl[49] vdd gnd cell_6t
Xbit_r50_c210 bl[210] br[210] wl[50] vdd gnd cell_6t
Xbit_r51_c210 bl[210] br[210] wl[51] vdd gnd cell_6t
Xbit_r52_c210 bl[210] br[210] wl[52] vdd gnd cell_6t
Xbit_r53_c210 bl[210] br[210] wl[53] vdd gnd cell_6t
Xbit_r54_c210 bl[210] br[210] wl[54] vdd gnd cell_6t
Xbit_r55_c210 bl[210] br[210] wl[55] vdd gnd cell_6t
Xbit_r56_c210 bl[210] br[210] wl[56] vdd gnd cell_6t
Xbit_r57_c210 bl[210] br[210] wl[57] vdd gnd cell_6t
Xbit_r58_c210 bl[210] br[210] wl[58] vdd gnd cell_6t
Xbit_r59_c210 bl[210] br[210] wl[59] vdd gnd cell_6t
Xbit_r60_c210 bl[210] br[210] wl[60] vdd gnd cell_6t
Xbit_r61_c210 bl[210] br[210] wl[61] vdd gnd cell_6t
Xbit_r62_c210 bl[210] br[210] wl[62] vdd gnd cell_6t
Xbit_r63_c210 bl[210] br[210] wl[63] vdd gnd cell_6t
Xbit_r64_c210 bl[210] br[210] wl[64] vdd gnd cell_6t
Xbit_r65_c210 bl[210] br[210] wl[65] vdd gnd cell_6t
Xbit_r66_c210 bl[210] br[210] wl[66] vdd gnd cell_6t
Xbit_r67_c210 bl[210] br[210] wl[67] vdd gnd cell_6t
Xbit_r68_c210 bl[210] br[210] wl[68] vdd gnd cell_6t
Xbit_r69_c210 bl[210] br[210] wl[69] vdd gnd cell_6t
Xbit_r70_c210 bl[210] br[210] wl[70] vdd gnd cell_6t
Xbit_r71_c210 bl[210] br[210] wl[71] vdd gnd cell_6t
Xbit_r72_c210 bl[210] br[210] wl[72] vdd gnd cell_6t
Xbit_r73_c210 bl[210] br[210] wl[73] vdd gnd cell_6t
Xbit_r74_c210 bl[210] br[210] wl[74] vdd gnd cell_6t
Xbit_r75_c210 bl[210] br[210] wl[75] vdd gnd cell_6t
Xbit_r76_c210 bl[210] br[210] wl[76] vdd gnd cell_6t
Xbit_r77_c210 bl[210] br[210] wl[77] vdd gnd cell_6t
Xbit_r78_c210 bl[210] br[210] wl[78] vdd gnd cell_6t
Xbit_r79_c210 bl[210] br[210] wl[79] vdd gnd cell_6t
Xbit_r80_c210 bl[210] br[210] wl[80] vdd gnd cell_6t
Xbit_r81_c210 bl[210] br[210] wl[81] vdd gnd cell_6t
Xbit_r82_c210 bl[210] br[210] wl[82] vdd gnd cell_6t
Xbit_r83_c210 bl[210] br[210] wl[83] vdd gnd cell_6t
Xbit_r84_c210 bl[210] br[210] wl[84] vdd gnd cell_6t
Xbit_r85_c210 bl[210] br[210] wl[85] vdd gnd cell_6t
Xbit_r86_c210 bl[210] br[210] wl[86] vdd gnd cell_6t
Xbit_r87_c210 bl[210] br[210] wl[87] vdd gnd cell_6t
Xbit_r88_c210 bl[210] br[210] wl[88] vdd gnd cell_6t
Xbit_r89_c210 bl[210] br[210] wl[89] vdd gnd cell_6t
Xbit_r90_c210 bl[210] br[210] wl[90] vdd gnd cell_6t
Xbit_r91_c210 bl[210] br[210] wl[91] vdd gnd cell_6t
Xbit_r92_c210 bl[210] br[210] wl[92] vdd gnd cell_6t
Xbit_r93_c210 bl[210] br[210] wl[93] vdd gnd cell_6t
Xbit_r94_c210 bl[210] br[210] wl[94] vdd gnd cell_6t
Xbit_r95_c210 bl[210] br[210] wl[95] vdd gnd cell_6t
Xbit_r96_c210 bl[210] br[210] wl[96] vdd gnd cell_6t
Xbit_r97_c210 bl[210] br[210] wl[97] vdd gnd cell_6t
Xbit_r98_c210 bl[210] br[210] wl[98] vdd gnd cell_6t
Xbit_r99_c210 bl[210] br[210] wl[99] vdd gnd cell_6t
Xbit_r100_c210 bl[210] br[210] wl[100] vdd gnd cell_6t
Xbit_r101_c210 bl[210] br[210] wl[101] vdd gnd cell_6t
Xbit_r102_c210 bl[210] br[210] wl[102] vdd gnd cell_6t
Xbit_r103_c210 bl[210] br[210] wl[103] vdd gnd cell_6t
Xbit_r104_c210 bl[210] br[210] wl[104] vdd gnd cell_6t
Xbit_r105_c210 bl[210] br[210] wl[105] vdd gnd cell_6t
Xbit_r106_c210 bl[210] br[210] wl[106] vdd gnd cell_6t
Xbit_r107_c210 bl[210] br[210] wl[107] vdd gnd cell_6t
Xbit_r108_c210 bl[210] br[210] wl[108] vdd gnd cell_6t
Xbit_r109_c210 bl[210] br[210] wl[109] vdd gnd cell_6t
Xbit_r110_c210 bl[210] br[210] wl[110] vdd gnd cell_6t
Xbit_r111_c210 bl[210] br[210] wl[111] vdd gnd cell_6t
Xbit_r112_c210 bl[210] br[210] wl[112] vdd gnd cell_6t
Xbit_r113_c210 bl[210] br[210] wl[113] vdd gnd cell_6t
Xbit_r114_c210 bl[210] br[210] wl[114] vdd gnd cell_6t
Xbit_r115_c210 bl[210] br[210] wl[115] vdd gnd cell_6t
Xbit_r116_c210 bl[210] br[210] wl[116] vdd gnd cell_6t
Xbit_r117_c210 bl[210] br[210] wl[117] vdd gnd cell_6t
Xbit_r118_c210 bl[210] br[210] wl[118] vdd gnd cell_6t
Xbit_r119_c210 bl[210] br[210] wl[119] vdd gnd cell_6t
Xbit_r120_c210 bl[210] br[210] wl[120] vdd gnd cell_6t
Xbit_r121_c210 bl[210] br[210] wl[121] vdd gnd cell_6t
Xbit_r122_c210 bl[210] br[210] wl[122] vdd gnd cell_6t
Xbit_r123_c210 bl[210] br[210] wl[123] vdd gnd cell_6t
Xbit_r124_c210 bl[210] br[210] wl[124] vdd gnd cell_6t
Xbit_r125_c210 bl[210] br[210] wl[125] vdd gnd cell_6t
Xbit_r126_c210 bl[210] br[210] wl[126] vdd gnd cell_6t
Xbit_r127_c210 bl[210] br[210] wl[127] vdd gnd cell_6t
Xbit_r128_c210 bl[210] br[210] wl[128] vdd gnd cell_6t
Xbit_r129_c210 bl[210] br[210] wl[129] vdd gnd cell_6t
Xbit_r130_c210 bl[210] br[210] wl[130] vdd gnd cell_6t
Xbit_r131_c210 bl[210] br[210] wl[131] vdd gnd cell_6t
Xbit_r132_c210 bl[210] br[210] wl[132] vdd gnd cell_6t
Xbit_r133_c210 bl[210] br[210] wl[133] vdd gnd cell_6t
Xbit_r134_c210 bl[210] br[210] wl[134] vdd gnd cell_6t
Xbit_r135_c210 bl[210] br[210] wl[135] vdd gnd cell_6t
Xbit_r136_c210 bl[210] br[210] wl[136] vdd gnd cell_6t
Xbit_r137_c210 bl[210] br[210] wl[137] vdd gnd cell_6t
Xbit_r138_c210 bl[210] br[210] wl[138] vdd gnd cell_6t
Xbit_r139_c210 bl[210] br[210] wl[139] vdd gnd cell_6t
Xbit_r140_c210 bl[210] br[210] wl[140] vdd gnd cell_6t
Xbit_r141_c210 bl[210] br[210] wl[141] vdd gnd cell_6t
Xbit_r142_c210 bl[210] br[210] wl[142] vdd gnd cell_6t
Xbit_r143_c210 bl[210] br[210] wl[143] vdd gnd cell_6t
Xbit_r144_c210 bl[210] br[210] wl[144] vdd gnd cell_6t
Xbit_r145_c210 bl[210] br[210] wl[145] vdd gnd cell_6t
Xbit_r146_c210 bl[210] br[210] wl[146] vdd gnd cell_6t
Xbit_r147_c210 bl[210] br[210] wl[147] vdd gnd cell_6t
Xbit_r148_c210 bl[210] br[210] wl[148] vdd gnd cell_6t
Xbit_r149_c210 bl[210] br[210] wl[149] vdd gnd cell_6t
Xbit_r150_c210 bl[210] br[210] wl[150] vdd gnd cell_6t
Xbit_r151_c210 bl[210] br[210] wl[151] vdd gnd cell_6t
Xbit_r152_c210 bl[210] br[210] wl[152] vdd gnd cell_6t
Xbit_r153_c210 bl[210] br[210] wl[153] vdd gnd cell_6t
Xbit_r154_c210 bl[210] br[210] wl[154] vdd gnd cell_6t
Xbit_r155_c210 bl[210] br[210] wl[155] vdd gnd cell_6t
Xbit_r156_c210 bl[210] br[210] wl[156] vdd gnd cell_6t
Xbit_r157_c210 bl[210] br[210] wl[157] vdd gnd cell_6t
Xbit_r158_c210 bl[210] br[210] wl[158] vdd gnd cell_6t
Xbit_r159_c210 bl[210] br[210] wl[159] vdd gnd cell_6t
Xbit_r160_c210 bl[210] br[210] wl[160] vdd gnd cell_6t
Xbit_r161_c210 bl[210] br[210] wl[161] vdd gnd cell_6t
Xbit_r162_c210 bl[210] br[210] wl[162] vdd gnd cell_6t
Xbit_r163_c210 bl[210] br[210] wl[163] vdd gnd cell_6t
Xbit_r164_c210 bl[210] br[210] wl[164] vdd gnd cell_6t
Xbit_r165_c210 bl[210] br[210] wl[165] vdd gnd cell_6t
Xbit_r166_c210 bl[210] br[210] wl[166] vdd gnd cell_6t
Xbit_r167_c210 bl[210] br[210] wl[167] vdd gnd cell_6t
Xbit_r168_c210 bl[210] br[210] wl[168] vdd gnd cell_6t
Xbit_r169_c210 bl[210] br[210] wl[169] vdd gnd cell_6t
Xbit_r170_c210 bl[210] br[210] wl[170] vdd gnd cell_6t
Xbit_r171_c210 bl[210] br[210] wl[171] vdd gnd cell_6t
Xbit_r172_c210 bl[210] br[210] wl[172] vdd gnd cell_6t
Xbit_r173_c210 bl[210] br[210] wl[173] vdd gnd cell_6t
Xbit_r174_c210 bl[210] br[210] wl[174] vdd gnd cell_6t
Xbit_r175_c210 bl[210] br[210] wl[175] vdd gnd cell_6t
Xbit_r176_c210 bl[210] br[210] wl[176] vdd gnd cell_6t
Xbit_r177_c210 bl[210] br[210] wl[177] vdd gnd cell_6t
Xbit_r178_c210 bl[210] br[210] wl[178] vdd gnd cell_6t
Xbit_r179_c210 bl[210] br[210] wl[179] vdd gnd cell_6t
Xbit_r180_c210 bl[210] br[210] wl[180] vdd gnd cell_6t
Xbit_r181_c210 bl[210] br[210] wl[181] vdd gnd cell_6t
Xbit_r182_c210 bl[210] br[210] wl[182] vdd gnd cell_6t
Xbit_r183_c210 bl[210] br[210] wl[183] vdd gnd cell_6t
Xbit_r184_c210 bl[210] br[210] wl[184] vdd gnd cell_6t
Xbit_r185_c210 bl[210] br[210] wl[185] vdd gnd cell_6t
Xbit_r186_c210 bl[210] br[210] wl[186] vdd gnd cell_6t
Xbit_r187_c210 bl[210] br[210] wl[187] vdd gnd cell_6t
Xbit_r188_c210 bl[210] br[210] wl[188] vdd gnd cell_6t
Xbit_r189_c210 bl[210] br[210] wl[189] vdd gnd cell_6t
Xbit_r190_c210 bl[210] br[210] wl[190] vdd gnd cell_6t
Xbit_r191_c210 bl[210] br[210] wl[191] vdd gnd cell_6t
Xbit_r192_c210 bl[210] br[210] wl[192] vdd gnd cell_6t
Xbit_r193_c210 bl[210] br[210] wl[193] vdd gnd cell_6t
Xbit_r194_c210 bl[210] br[210] wl[194] vdd gnd cell_6t
Xbit_r195_c210 bl[210] br[210] wl[195] vdd gnd cell_6t
Xbit_r196_c210 bl[210] br[210] wl[196] vdd gnd cell_6t
Xbit_r197_c210 bl[210] br[210] wl[197] vdd gnd cell_6t
Xbit_r198_c210 bl[210] br[210] wl[198] vdd gnd cell_6t
Xbit_r199_c210 bl[210] br[210] wl[199] vdd gnd cell_6t
Xbit_r200_c210 bl[210] br[210] wl[200] vdd gnd cell_6t
Xbit_r201_c210 bl[210] br[210] wl[201] vdd gnd cell_6t
Xbit_r202_c210 bl[210] br[210] wl[202] vdd gnd cell_6t
Xbit_r203_c210 bl[210] br[210] wl[203] vdd gnd cell_6t
Xbit_r204_c210 bl[210] br[210] wl[204] vdd gnd cell_6t
Xbit_r205_c210 bl[210] br[210] wl[205] vdd gnd cell_6t
Xbit_r206_c210 bl[210] br[210] wl[206] vdd gnd cell_6t
Xbit_r207_c210 bl[210] br[210] wl[207] vdd gnd cell_6t
Xbit_r208_c210 bl[210] br[210] wl[208] vdd gnd cell_6t
Xbit_r209_c210 bl[210] br[210] wl[209] vdd gnd cell_6t
Xbit_r210_c210 bl[210] br[210] wl[210] vdd gnd cell_6t
Xbit_r211_c210 bl[210] br[210] wl[211] vdd gnd cell_6t
Xbit_r212_c210 bl[210] br[210] wl[212] vdd gnd cell_6t
Xbit_r213_c210 bl[210] br[210] wl[213] vdd gnd cell_6t
Xbit_r214_c210 bl[210] br[210] wl[214] vdd gnd cell_6t
Xbit_r215_c210 bl[210] br[210] wl[215] vdd gnd cell_6t
Xbit_r216_c210 bl[210] br[210] wl[216] vdd gnd cell_6t
Xbit_r217_c210 bl[210] br[210] wl[217] vdd gnd cell_6t
Xbit_r218_c210 bl[210] br[210] wl[218] vdd gnd cell_6t
Xbit_r219_c210 bl[210] br[210] wl[219] vdd gnd cell_6t
Xbit_r220_c210 bl[210] br[210] wl[220] vdd gnd cell_6t
Xbit_r221_c210 bl[210] br[210] wl[221] vdd gnd cell_6t
Xbit_r222_c210 bl[210] br[210] wl[222] vdd gnd cell_6t
Xbit_r223_c210 bl[210] br[210] wl[223] vdd gnd cell_6t
Xbit_r224_c210 bl[210] br[210] wl[224] vdd gnd cell_6t
Xbit_r225_c210 bl[210] br[210] wl[225] vdd gnd cell_6t
Xbit_r226_c210 bl[210] br[210] wl[226] vdd gnd cell_6t
Xbit_r227_c210 bl[210] br[210] wl[227] vdd gnd cell_6t
Xbit_r228_c210 bl[210] br[210] wl[228] vdd gnd cell_6t
Xbit_r229_c210 bl[210] br[210] wl[229] vdd gnd cell_6t
Xbit_r230_c210 bl[210] br[210] wl[230] vdd gnd cell_6t
Xbit_r231_c210 bl[210] br[210] wl[231] vdd gnd cell_6t
Xbit_r232_c210 bl[210] br[210] wl[232] vdd gnd cell_6t
Xbit_r233_c210 bl[210] br[210] wl[233] vdd gnd cell_6t
Xbit_r234_c210 bl[210] br[210] wl[234] vdd gnd cell_6t
Xbit_r235_c210 bl[210] br[210] wl[235] vdd gnd cell_6t
Xbit_r236_c210 bl[210] br[210] wl[236] vdd gnd cell_6t
Xbit_r237_c210 bl[210] br[210] wl[237] vdd gnd cell_6t
Xbit_r238_c210 bl[210] br[210] wl[238] vdd gnd cell_6t
Xbit_r239_c210 bl[210] br[210] wl[239] vdd gnd cell_6t
Xbit_r240_c210 bl[210] br[210] wl[240] vdd gnd cell_6t
Xbit_r241_c210 bl[210] br[210] wl[241] vdd gnd cell_6t
Xbit_r242_c210 bl[210] br[210] wl[242] vdd gnd cell_6t
Xbit_r243_c210 bl[210] br[210] wl[243] vdd gnd cell_6t
Xbit_r244_c210 bl[210] br[210] wl[244] vdd gnd cell_6t
Xbit_r245_c210 bl[210] br[210] wl[245] vdd gnd cell_6t
Xbit_r246_c210 bl[210] br[210] wl[246] vdd gnd cell_6t
Xbit_r247_c210 bl[210] br[210] wl[247] vdd gnd cell_6t
Xbit_r248_c210 bl[210] br[210] wl[248] vdd gnd cell_6t
Xbit_r249_c210 bl[210] br[210] wl[249] vdd gnd cell_6t
Xbit_r250_c210 bl[210] br[210] wl[250] vdd gnd cell_6t
Xbit_r251_c210 bl[210] br[210] wl[251] vdd gnd cell_6t
Xbit_r252_c210 bl[210] br[210] wl[252] vdd gnd cell_6t
Xbit_r253_c210 bl[210] br[210] wl[253] vdd gnd cell_6t
Xbit_r254_c210 bl[210] br[210] wl[254] vdd gnd cell_6t
Xbit_r255_c210 bl[210] br[210] wl[255] vdd gnd cell_6t
Xbit_r0_c211 bl[211] br[211] wl[0] vdd gnd cell_6t
Xbit_r1_c211 bl[211] br[211] wl[1] vdd gnd cell_6t
Xbit_r2_c211 bl[211] br[211] wl[2] vdd gnd cell_6t
Xbit_r3_c211 bl[211] br[211] wl[3] vdd gnd cell_6t
Xbit_r4_c211 bl[211] br[211] wl[4] vdd gnd cell_6t
Xbit_r5_c211 bl[211] br[211] wl[5] vdd gnd cell_6t
Xbit_r6_c211 bl[211] br[211] wl[6] vdd gnd cell_6t
Xbit_r7_c211 bl[211] br[211] wl[7] vdd gnd cell_6t
Xbit_r8_c211 bl[211] br[211] wl[8] vdd gnd cell_6t
Xbit_r9_c211 bl[211] br[211] wl[9] vdd gnd cell_6t
Xbit_r10_c211 bl[211] br[211] wl[10] vdd gnd cell_6t
Xbit_r11_c211 bl[211] br[211] wl[11] vdd gnd cell_6t
Xbit_r12_c211 bl[211] br[211] wl[12] vdd gnd cell_6t
Xbit_r13_c211 bl[211] br[211] wl[13] vdd gnd cell_6t
Xbit_r14_c211 bl[211] br[211] wl[14] vdd gnd cell_6t
Xbit_r15_c211 bl[211] br[211] wl[15] vdd gnd cell_6t
Xbit_r16_c211 bl[211] br[211] wl[16] vdd gnd cell_6t
Xbit_r17_c211 bl[211] br[211] wl[17] vdd gnd cell_6t
Xbit_r18_c211 bl[211] br[211] wl[18] vdd gnd cell_6t
Xbit_r19_c211 bl[211] br[211] wl[19] vdd gnd cell_6t
Xbit_r20_c211 bl[211] br[211] wl[20] vdd gnd cell_6t
Xbit_r21_c211 bl[211] br[211] wl[21] vdd gnd cell_6t
Xbit_r22_c211 bl[211] br[211] wl[22] vdd gnd cell_6t
Xbit_r23_c211 bl[211] br[211] wl[23] vdd gnd cell_6t
Xbit_r24_c211 bl[211] br[211] wl[24] vdd gnd cell_6t
Xbit_r25_c211 bl[211] br[211] wl[25] vdd gnd cell_6t
Xbit_r26_c211 bl[211] br[211] wl[26] vdd gnd cell_6t
Xbit_r27_c211 bl[211] br[211] wl[27] vdd gnd cell_6t
Xbit_r28_c211 bl[211] br[211] wl[28] vdd gnd cell_6t
Xbit_r29_c211 bl[211] br[211] wl[29] vdd gnd cell_6t
Xbit_r30_c211 bl[211] br[211] wl[30] vdd gnd cell_6t
Xbit_r31_c211 bl[211] br[211] wl[31] vdd gnd cell_6t
Xbit_r32_c211 bl[211] br[211] wl[32] vdd gnd cell_6t
Xbit_r33_c211 bl[211] br[211] wl[33] vdd gnd cell_6t
Xbit_r34_c211 bl[211] br[211] wl[34] vdd gnd cell_6t
Xbit_r35_c211 bl[211] br[211] wl[35] vdd gnd cell_6t
Xbit_r36_c211 bl[211] br[211] wl[36] vdd gnd cell_6t
Xbit_r37_c211 bl[211] br[211] wl[37] vdd gnd cell_6t
Xbit_r38_c211 bl[211] br[211] wl[38] vdd gnd cell_6t
Xbit_r39_c211 bl[211] br[211] wl[39] vdd gnd cell_6t
Xbit_r40_c211 bl[211] br[211] wl[40] vdd gnd cell_6t
Xbit_r41_c211 bl[211] br[211] wl[41] vdd gnd cell_6t
Xbit_r42_c211 bl[211] br[211] wl[42] vdd gnd cell_6t
Xbit_r43_c211 bl[211] br[211] wl[43] vdd gnd cell_6t
Xbit_r44_c211 bl[211] br[211] wl[44] vdd gnd cell_6t
Xbit_r45_c211 bl[211] br[211] wl[45] vdd gnd cell_6t
Xbit_r46_c211 bl[211] br[211] wl[46] vdd gnd cell_6t
Xbit_r47_c211 bl[211] br[211] wl[47] vdd gnd cell_6t
Xbit_r48_c211 bl[211] br[211] wl[48] vdd gnd cell_6t
Xbit_r49_c211 bl[211] br[211] wl[49] vdd gnd cell_6t
Xbit_r50_c211 bl[211] br[211] wl[50] vdd gnd cell_6t
Xbit_r51_c211 bl[211] br[211] wl[51] vdd gnd cell_6t
Xbit_r52_c211 bl[211] br[211] wl[52] vdd gnd cell_6t
Xbit_r53_c211 bl[211] br[211] wl[53] vdd gnd cell_6t
Xbit_r54_c211 bl[211] br[211] wl[54] vdd gnd cell_6t
Xbit_r55_c211 bl[211] br[211] wl[55] vdd gnd cell_6t
Xbit_r56_c211 bl[211] br[211] wl[56] vdd gnd cell_6t
Xbit_r57_c211 bl[211] br[211] wl[57] vdd gnd cell_6t
Xbit_r58_c211 bl[211] br[211] wl[58] vdd gnd cell_6t
Xbit_r59_c211 bl[211] br[211] wl[59] vdd gnd cell_6t
Xbit_r60_c211 bl[211] br[211] wl[60] vdd gnd cell_6t
Xbit_r61_c211 bl[211] br[211] wl[61] vdd gnd cell_6t
Xbit_r62_c211 bl[211] br[211] wl[62] vdd gnd cell_6t
Xbit_r63_c211 bl[211] br[211] wl[63] vdd gnd cell_6t
Xbit_r64_c211 bl[211] br[211] wl[64] vdd gnd cell_6t
Xbit_r65_c211 bl[211] br[211] wl[65] vdd gnd cell_6t
Xbit_r66_c211 bl[211] br[211] wl[66] vdd gnd cell_6t
Xbit_r67_c211 bl[211] br[211] wl[67] vdd gnd cell_6t
Xbit_r68_c211 bl[211] br[211] wl[68] vdd gnd cell_6t
Xbit_r69_c211 bl[211] br[211] wl[69] vdd gnd cell_6t
Xbit_r70_c211 bl[211] br[211] wl[70] vdd gnd cell_6t
Xbit_r71_c211 bl[211] br[211] wl[71] vdd gnd cell_6t
Xbit_r72_c211 bl[211] br[211] wl[72] vdd gnd cell_6t
Xbit_r73_c211 bl[211] br[211] wl[73] vdd gnd cell_6t
Xbit_r74_c211 bl[211] br[211] wl[74] vdd gnd cell_6t
Xbit_r75_c211 bl[211] br[211] wl[75] vdd gnd cell_6t
Xbit_r76_c211 bl[211] br[211] wl[76] vdd gnd cell_6t
Xbit_r77_c211 bl[211] br[211] wl[77] vdd gnd cell_6t
Xbit_r78_c211 bl[211] br[211] wl[78] vdd gnd cell_6t
Xbit_r79_c211 bl[211] br[211] wl[79] vdd gnd cell_6t
Xbit_r80_c211 bl[211] br[211] wl[80] vdd gnd cell_6t
Xbit_r81_c211 bl[211] br[211] wl[81] vdd gnd cell_6t
Xbit_r82_c211 bl[211] br[211] wl[82] vdd gnd cell_6t
Xbit_r83_c211 bl[211] br[211] wl[83] vdd gnd cell_6t
Xbit_r84_c211 bl[211] br[211] wl[84] vdd gnd cell_6t
Xbit_r85_c211 bl[211] br[211] wl[85] vdd gnd cell_6t
Xbit_r86_c211 bl[211] br[211] wl[86] vdd gnd cell_6t
Xbit_r87_c211 bl[211] br[211] wl[87] vdd gnd cell_6t
Xbit_r88_c211 bl[211] br[211] wl[88] vdd gnd cell_6t
Xbit_r89_c211 bl[211] br[211] wl[89] vdd gnd cell_6t
Xbit_r90_c211 bl[211] br[211] wl[90] vdd gnd cell_6t
Xbit_r91_c211 bl[211] br[211] wl[91] vdd gnd cell_6t
Xbit_r92_c211 bl[211] br[211] wl[92] vdd gnd cell_6t
Xbit_r93_c211 bl[211] br[211] wl[93] vdd gnd cell_6t
Xbit_r94_c211 bl[211] br[211] wl[94] vdd gnd cell_6t
Xbit_r95_c211 bl[211] br[211] wl[95] vdd gnd cell_6t
Xbit_r96_c211 bl[211] br[211] wl[96] vdd gnd cell_6t
Xbit_r97_c211 bl[211] br[211] wl[97] vdd gnd cell_6t
Xbit_r98_c211 bl[211] br[211] wl[98] vdd gnd cell_6t
Xbit_r99_c211 bl[211] br[211] wl[99] vdd gnd cell_6t
Xbit_r100_c211 bl[211] br[211] wl[100] vdd gnd cell_6t
Xbit_r101_c211 bl[211] br[211] wl[101] vdd gnd cell_6t
Xbit_r102_c211 bl[211] br[211] wl[102] vdd gnd cell_6t
Xbit_r103_c211 bl[211] br[211] wl[103] vdd gnd cell_6t
Xbit_r104_c211 bl[211] br[211] wl[104] vdd gnd cell_6t
Xbit_r105_c211 bl[211] br[211] wl[105] vdd gnd cell_6t
Xbit_r106_c211 bl[211] br[211] wl[106] vdd gnd cell_6t
Xbit_r107_c211 bl[211] br[211] wl[107] vdd gnd cell_6t
Xbit_r108_c211 bl[211] br[211] wl[108] vdd gnd cell_6t
Xbit_r109_c211 bl[211] br[211] wl[109] vdd gnd cell_6t
Xbit_r110_c211 bl[211] br[211] wl[110] vdd gnd cell_6t
Xbit_r111_c211 bl[211] br[211] wl[111] vdd gnd cell_6t
Xbit_r112_c211 bl[211] br[211] wl[112] vdd gnd cell_6t
Xbit_r113_c211 bl[211] br[211] wl[113] vdd gnd cell_6t
Xbit_r114_c211 bl[211] br[211] wl[114] vdd gnd cell_6t
Xbit_r115_c211 bl[211] br[211] wl[115] vdd gnd cell_6t
Xbit_r116_c211 bl[211] br[211] wl[116] vdd gnd cell_6t
Xbit_r117_c211 bl[211] br[211] wl[117] vdd gnd cell_6t
Xbit_r118_c211 bl[211] br[211] wl[118] vdd gnd cell_6t
Xbit_r119_c211 bl[211] br[211] wl[119] vdd gnd cell_6t
Xbit_r120_c211 bl[211] br[211] wl[120] vdd gnd cell_6t
Xbit_r121_c211 bl[211] br[211] wl[121] vdd gnd cell_6t
Xbit_r122_c211 bl[211] br[211] wl[122] vdd gnd cell_6t
Xbit_r123_c211 bl[211] br[211] wl[123] vdd gnd cell_6t
Xbit_r124_c211 bl[211] br[211] wl[124] vdd gnd cell_6t
Xbit_r125_c211 bl[211] br[211] wl[125] vdd gnd cell_6t
Xbit_r126_c211 bl[211] br[211] wl[126] vdd gnd cell_6t
Xbit_r127_c211 bl[211] br[211] wl[127] vdd gnd cell_6t
Xbit_r128_c211 bl[211] br[211] wl[128] vdd gnd cell_6t
Xbit_r129_c211 bl[211] br[211] wl[129] vdd gnd cell_6t
Xbit_r130_c211 bl[211] br[211] wl[130] vdd gnd cell_6t
Xbit_r131_c211 bl[211] br[211] wl[131] vdd gnd cell_6t
Xbit_r132_c211 bl[211] br[211] wl[132] vdd gnd cell_6t
Xbit_r133_c211 bl[211] br[211] wl[133] vdd gnd cell_6t
Xbit_r134_c211 bl[211] br[211] wl[134] vdd gnd cell_6t
Xbit_r135_c211 bl[211] br[211] wl[135] vdd gnd cell_6t
Xbit_r136_c211 bl[211] br[211] wl[136] vdd gnd cell_6t
Xbit_r137_c211 bl[211] br[211] wl[137] vdd gnd cell_6t
Xbit_r138_c211 bl[211] br[211] wl[138] vdd gnd cell_6t
Xbit_r139_c211 bl[211] br[211] wl[139] vdd gnd cell_6t
Xbit_r140_c211 bl[211] br[211] wl[140] vdd gnd cell_6t
Xbit_r141_c211 bl[211] br[211] wl[141] vdd gnd cell_6t
Xbit_r142_c211 bl[211] br[211] wl[142] vdd gnd cell_6t
Xbit_r143_c211 bl[211] br[211] wl[143] vdd gnd cell_6t
Xbit_r144_c211 bl[211] br[211] wl[144] vdd gnd cell_6t
Xbit_r145_c211 bl[211] br[211] wl[145] vdd gnd cell_6t
Xbit_r146_c211 bl[211] br[211] wl[146] vdd gnd cell_6t
Xbit_r147_c211 bl[211] br[211] wl[147] vdd gnd cell_6t
Xbit_r148_c211 bl[211] br[211] wl[148] vdd gnd cell_6t
Xbit_r149_c211 bl[211] br[211] wl[149] vdd gnd cell_6t
Xbit_r150_c211 bl[211] br[211] wl[150] vdd gnd cell_6t
Xbit_r151_c211 bl[211] br[211] wl[151] vdd gnd cell_6t
Xbit_r152_c211 bl[211] br[211] wl[152] vdd gnd cell_6t
Xbit_r153_c211 bl[211] br[211] wl[153] vdd gnd cell_6t
Xbit_r154_c211 bl[211] br[211] wl[154] vdd gnd cell_6t
Xbit_r155_c211 bl[211] br[211] wl[155] vdd gnd cell_6t
Xbit_r156_c211 bl[211] br[211] wl[156] vdd gnd cell_6t
Xbit_r157_c211 bl[211] br[211] wl[157] vdd gnd cell_6t
Xbit_r158_c211 bl[211] br[211] wl[158] vdd gnd cell_6t
Xbit_r159_c211 bl[211] br[211] wl[159] vdd gnd cell_6t
Xbit_r160_c211 bl[211] br[211] wl[160] vdd gnd cell_6t
Xbit_r161_c211 bl[211] br[211] wl[161] vdd gnd cell_6t
Xbit_r162_c211 bl[211] br[211] wl[162] vdd gnd cell_6t
Xbit_r163_c211 bl[211] br[211] wl[163] vdd gnd cell_6t
Xbit_r164_c211 bl[211] br[211] wl[164] vdd gnd cell_6t
Xbit_r165_c211 bl[211] br[211] wl[165] vdd gnd cell_6t
Xbit_r166_c211 bl[211] br[211] wl[166] vdd gnd cell_6t
Xbit_r167_c211 bl[211] br[211] wl[167] vdd gnd cell_6t
Xbit_r168_c211 bl[211] br[211] wl[168] vdd gnd cell_6t
Xbit_r169_c211 bl[211] br[211] wl[169] vdd gnd cell_6t
Xbit_r170_c211 bl[211] br[211] wl[170] vdd gnd cell_6t
Xbit_r171_c211 bl[211] br[211] wl[171] vdd gnd cell_6t
Xbit_r172_c211 bl[211] br[211] wl[172] vdd gnd cell_6t
Xbit_r173_c211 bl[211] br[211] wl[173] vdd gnd cell_6t
Xbit_r174_c211 bl[211] br[211] wl[174] vdd gnd cell_6t
Xbit_r175_c211 bl[211] br[211] wl[175] vdd gnd cell_6t
Xbit_r176_c211 bl[211] br[211] wl[176] vdd gnd cell_6t
Xbit_r177_c211 bl[211] br[211] wl[177] vdd gnd cell_6t
Xbit_r178_c211 bl[211] br[211] wl[178] vdd gnd cell_6t
Xbit_r179_c211 bl[211] br[211] wl[179] vdd gnd cell_6t
Xbit_r180_c211 bl[211] br[211] wl[180] vdd gnd cell_6t
Xbit_r181_c211 bl[211] br[211] wl[181] vdd gnd cell_6t
Xbit_r182_c211 bl[211] br[211] wl[182] vdd gnd cell_6t
Xbit_r183_c211 bl[211] br[211] wl[183] vdd gnd cell_6t
Xbit_r184_c211 bl[211] br[211] wl[184] vdd gnd cell_6t
Xbit_r185_c211 bl[211] br[211] wl[185] vdd gnd cell_6t
Xbit_r186_c211 bl[211] br[211] wl[186] vdd gnd cell_6t
Xbit_r187_c211 bl[211] br[211] wl[187] vdd gnd cell_6t
Xbit_r188_c211 bl[211] br[211] wl[188] vdd gnd cell_6t
Xbit_r189_c211 bl[211] br[211] wl[189] vdd gnd cell_6t
Xbit_r190_c211 bl[211] br[211] wl[190] vdd gnd cell_6t
Xbit_r191_c211 bl[211] br[211] wl[191] vdd gnd cell_6t
Xbit_r192_c211 bl[211] br[211] wl[192] vdd gnd cell_6t
Xbit_r193_c211 bl[211] br[211] wl[193] vdd gnd cell_6t
Xbit_r194_c211 bl[211] br[211] wl[194] vdd gnd cell_6t
Xbit_r195_c211 bl[211] br[211] wl[195] vdd gnd cell_6t
Xbit_r196_c211 bl[211] br[211] wl[196] vdd gnd cell_6t
Xbit_r197_c211 bl[211] br[211] wl[197] vdd gnd cell_6t
Xbit_r198_c211 bl[211] br[211] wl[198] vdd gnd cell_6t
Xbit_r199_c211 bl[211] br[211] wl[199] vdd gnd cell_6t
Xbit_r200_c211 bl[211] br[211] wl[200] vdd gnd cell_6t
Xbit_r201_c211 bl[211] br[211] wl[201] vdd gnd cell_6t
Xbit_r202_c211 bl[211] br[211] wl[202] vdd gnd cell_6t
Xbit_r203_c211 bl[211] br[211] wl[203] vdd gnd cell_6t
Xbit_r204_c211 bl[211] br[211] wl[204] vdd gnd cell_6t
Xbit_r205_c211 bl[211] br[211] wl[205] vdd gnd cell_6t
Xbit_r206_c211 bl[211] br[211] wl[206] vdd gnd cell_6t
Xbit_r207_c211 bl[211] br[211] wl[207] vdd gnd cell_6t
Xbit_r208_c211 bl[211] br[211] wl[208] vdd gnd cell_6t
Xbit_r209_c211 bl[211] br[211] wl[209] vdd gnd cell_6t
Xbit_r210_c211 bl[211] br[211] wl[210] vdd gnd cell_6t
Xbit_r211_c211 bl[211] br[211] wl[211] vdd gnd cell_6t
Xbit_r212_c211 bl[211] br[211] wl[212] vdd gnd cell_6t
Xbit_r213_c211 bl[211] br[211] wl[213] vdd gnd cell_6t
Xbit_r214_c211 bl[211] br[211] wl[214] vdd gnd cell_6t
Xbit_r215_c211 bl[211] br[211] wl[215] vdd gnd cell_6t
Xbit_r216_c211 bl[211] br[211] wl[216] vdd gnd cell_6t
Xbit_r217_c211 bl[211] br[211] wl[217] vdd gnd cell_6t
Xbit_r218_c211 bl[211] br[211] wl[218] vdd gnd cell_6t
Xbit_r219_c211 bl[211] br[211] wl[219] vdd gnd cell_6t
Xbit_r220_c211 bl[211] br[211] wl[220] vdd gnd cell_6t
Xbit_r221_c211 bl[211] br[211] wl[221] vdd gnd cell_6t
Xbit_r222_c211 bl[211] br[211] wl[222] vdd gnd cell_6t
Xbit_r223_c211 bl[211] br[211] wl[223] vdd gnd cell_6t
Xbit_r224_c211 bl[211] br[211] wl[224] vdd gnd cell_6t
Xbit_r225_c211 bl[211] br[211] wl[225] vdd gnd cell_6t
Xbit_r226_c211 bl[211] br[211] wl[226] vdd gnd cell_6t
Xbit_r227_c211 bl[211] br[211] wl[227] vdd gnd cell_6t
Xbit_r228_c211 bl[211] br[211] wl[228] vdd gnd cell_6t
Xbit_r229_c211 bl[211] br[211] wl[229] vdd gnd cell_6t
Xbit_r230_c211 bl[211] br[211] wl[230] vdd gnd cell_6t
Xbit_r231_c211 bl[211] br[211] wl[231] vdd gnd cell_6t
Xbit_r232_c211 bl[211] br[211] wl[232] vdd gnd cell_6t
Xbit_r233_c211 bl[211] br[211] wl[233] vdd gnd cell_6t
Xbit_r234_c211 bl[211] br[211] wl[234] vdd gnd cell_6t
Xbit_r235_c211 bl[211] br[211] wl[235] vdd gnd cell_6t
Xbit_r236_c211 bl[211] br[211] wl[236] vdd gnd cell_6t
Xbit_r237_c211 bl[211] br[211] wl[237] vdd gnd cell_6t
Xbit_r238_c211 bl[211] br[211] wl[238] vdd gnd cell_6t
Xbit_r239_c211 bl[211] br[211] wl[239] vdd gnd cell_6t
Xbit_r240_c211 bl[211] br[211] wl[240] vdd gnd cell_6t
Xbit_r241_c211 bl[211] br[211] wl[241] vdd gnd cell_6t
Xbit_r242_c211 bl[211] br[211] wl[242] vdd gnd cell_6t
Xbit_r243_c211 bl[211] br[211] wl[243] vdd gnd cell_6t
Xbit_r244_c211 bl[211] br[211] wl[244] vdd gnd cell_6t
Xbit_r245_c211 bl[211] br[211] wl[245] vdd gnd cell_6t
Xbit_r246_c211 bl[211] br[211] wl[246] vdd gnd cell_6t
Xbit_r247_c211 bl[211] br[211] wl[247] vdd gnd cell_6t
Xbit_r248_c211 bl[211] br[211] wl[248] vdd gnd cell_6t
Xbit_r249_c211 bl[211] br[211] wl[249] vdd gnd cell_6t
Xbit_r250_c211 bl[211] br[211] wl[250] vdd gnd cell_6t
Xbit_r251_c211 bl[211] br[211] wl[251] vdd gnd cell_6t
Xbit_r252_c211 bl[211] br[211] wl[252] vdd gnd cell_6t
Xbit_r253_c211 bl[211] br[211] wl[253] vdd gnd cell_6t
Xbit_r254_c211 bl[211] br[211] wl[254] vdd gnd cell_6t
Xbit_r255_c211 bl[211] br[211] wl[255] vdd gnd cell_6t
Xbit_r0_c212 bl[212] br[212] wl[0] vdd gnd cell_6t
Xbit_r1_c212 bl[212] br[212] wl[1] vdd gnd cell_6t
Xbit_r2_c212 bl[212] br[212] wl[2] vdd gnd cell_6t
Xbit_r3_c212 bl[212] br[212] wl[3] vdd gnd cell_6t
Xbit_r4_c212 bl[212] br[212] wl[4] vdd gnd cell_6t
Xbit_r5_c212 bl[212] br[212] wl[5] vdd gnd cell_6t
Xbit_r6_c212 bl[212] br[212] wl[6] vdd gnd cell_6t
Xbit_r7_c212 bl[212] br[212] wl[7] vdd gnd cell_6t
Xbit_r8_c212 bl[212] br[212] wl[8] vdd gnd cell_6t
Xbit_r9_c212 bl[212] br[212] wl[9] vdd gnd cell_6t
Xbit_r10_c212 bl[212] br[212] wl[10] vdd gnd cell_6t
Xbit_r11_c212 bl[212] br[212] wl[11] vdd gnd cell_6t
Xbit_r12_c212 bl[212] br[212] wl[12] vdd gnd cell_6t
Xbit_r13_c212 bl[212] br[212] wl[13] vdd gnd cell_6t
Xbit_r14_c212 bl[212] br[212] wl[14] vdd gnd cell_6t
Xbit_r15_c212 bl[212] br[212] wl[15] vdd gnd cell_6t
Xbit_r16_c212 bl[212] br[212] wl[16] vdd gnd cell_6t
Xbit_r17_c212 bl[212] br[212] wl[17] vdd gnd cell_6t
Xbit_r18_c212 bl[212] br[212] wl[18] vdd gnd cell_6t
Xbit_r19_c212 bl[212] br[212] wl[19] vdd gnd cell_6t
Xbit_r20_c212 bl[212] br[212] wl[20] vdd gnd cell_6t
Xbit_r21_c212 bl[212] br[212] wl[21] vdd gnd cell_6t
Xbit_r22_c212 bl[212] br[212] wl[22] vdd gnd cell_6t
Xbit_r23_c212 bl[212] br[212] wl[23] vdd gnd cell_6t
Xbit_r24_c212 bl[212] br[212] wl[24] vdd gnd cell_6t
Xbit_r25_c212 bl[212] br[212] wl[25] vdd gnd cell_6t
Xbit_r26_c212 bl[212] br[212] wl[26] vdd gnd cell_6t
Xbit_r27_c212 bl[212] br[212] wl[27] vdd gnd cell_6t
Xbit_r28_c212 bl[212] br[212] wl[28] vdd gnd cell_6t
Xbit_r29_c212 bl[212] br[212] wl[29] vdd gnd cell_6t
Xbit_r30_c212 bl[212] br[212] wl[30] vdd gnd cell_6t
Xbit_r31_c212 bl[212] br[212] wl[31] vdd gnd cell_6t
Xbit_r32_c212 bl[212] br[212] wl[32] vdd gnd cell_6t
Xbit_r33_c212 bl[212] br[212] wl[33] vdd gnd cell_6t
Xbit_r34_c212 bl[212] br[212] wl[34] vdd gnd cell_6t
Xbit_r35_c212 bl[212] br[212] wl[35] vdd gnd cell_6t
Xbit_r36_c212 bl[212] br[212] wl[36] vdd gnd cell_6t
Xbit_r37_c212 bl[212] br[212] wl[37] vdd gnd cell_6t
Xbit_r38_c212 bl[212] br[212] wl[38] vdd gnd cell_6t
Xbit_r39_c212 bl[212] br[212] wl[39] vdd gnd cell_6t
Xbit_r40_c212 bl[212] br[212] wl[40] vdd gnd cell_6t
Xbit_r41_c212 bl[212] br[212] wl[41] vdd gnd cell_6t
Xbit_r42_c212 bl[212] br[212] wl[42] vdd gnd cell_6t
Xbit_r43_c212 bl[212] br[212] wl[43] vdd gnd cell_6t
Xbit_r44_c212 bl[212] br[212] wl[44] vdd gnd cell_6t
Xbit_r45_c212 bl[212] br[212] wl[45] vdd gnd cell_6t
Xbit_r46_c212 bl[212] br[212] wl[46] vdd gnd cell_6t
Xbit_r47_c212 bl[212] br[212] wl[47] vdd gnd cell_6t
Xbit_r48_c212 bl[212] br[212] wl[48] vdd gnd cell_6t
Xbit_r49_c212 bl[212] br[212] wl[49] vdd gnd cell_6t
Xbit_r50_c212 bl[212] br[212] wl[50] vdd gnd cell_6t
Xbit_r51_c212 bl[212] br[212] wl[51] vdd gnd cell_6t
Xbit_r52_c212 bl[212] br[212] wl[52] vdd gnd cell_6t
Xbit_r53_c212 bl[212] br[212] wl[53] vdd gnd cell_6t
Xbit_r54_c212 bl[212] br[212] wl[54] vdd gnd cell_6t
Xbit_r55_c212 bl[212] br[212] wl[55] vdd gnd cell_6t
Xbit_r56_c212 bl[212] br[212] wl[56] vdd gnd cell_6t
Xbit_r57_c212 bl[212] br[212] wl[57] vdd gnd cell_6t
Xbit_r58_c212 bl[212] br[212] wl[58] vdd gnd cell_6t
Xbit_r59_c212 bl[212] br[212] wl[59] vdd gnd cell_6t
Xbit_r60_c212 bl[212] br[212] wl[60] vdd gnd cell_6t
Xbit_r61_c212 bl[212] br[212] wl[61] vdd gnd cell_6t
Xbit_r62_c212 bl[212] br[212] wl[62] vdd gnd cell_6t
Xbit_r63_c212 bl[212] br[212] wl[63] vdd gnd cell_6t
Xbit_r64_c212 bl[212] br[212] wl[64] vdd gnd cell_6t
Xbit_r65_c212 bl[212] br[212] wl[65] vdd gnd cell_6t
Xbit_r66_c212 bl[212] br[212] wl[66] vdd gnd cell_6t
Xbit_r67_c212 bl[212] br[212] wl[67] vdd gnd cell_6t
Xbit_r68_c212 bl[212] br[212] wl[68] vdd gnd cell_6t
Xbit_r69_c212 bl[212] br[212] wl[69] vdd gnd cell_6t
Xbit_r70_c212 bl[212] br[212] wl[70] vdd gnd cell_6t
Xbit_r71_c212 bl[212] br[212] wl[71] vdd gnd cell_6t
Xbit_r72_c212 bl[212] br[212] wl[72] vdd gnd cell_6t
Xbit_r73_c212 bl[212] br[212] wl[73] vdd gnd cell_6t
Xbit_r74_c212 bl[212] br[212] wl[74] vdd gnd cell_6t
Xbit_r75_c212 bl[212] br[212] wl[75] vdd gnd cell_6t
Xbit_r76_c212 bl[212] br[212] wl[76] vdd gnd cell_6t
Xbit_r77_c212 bl[212] br[212] wl[77] vdd gnd cell_6t
Xbit_r78_c212 bl[212] br[212] wl[78] vdd gnd cell_6t
Xbit_r79_c212 bl[212] br[212] wl[79] vdd gnd cell_6t
Xbit_r80_c212 bl[212] br[212] wl[80] vdd gnd cell_6t
Xbit_r81_c212 bl[212] br[212] wl[81] vdd gnd cell_6t
Xbit_r82_c212 bl[212] br[212] wl[82] vdd gnd cell_6t
Xbit_r83_c212 bl[212] br[212] wl[83] vdd gnd cell_6t
Xbit_r84_c212 bl[212] br[212] wl[84] vdd gnd cell_6t
Xbit_r85_c212 bl[212] br[212] wl[85] vdd gnd cell_6t
Xbit_r86_c212 bl[212] br[212] wl[86] vdd gnd cell_6t
Xbit_r87_c212 bl[212] br[212] wl[87] vdd gnd cell_6t
Xbit_r88_c212 bl[212] br[212] wl[88] vdd gnd cell_6t
Xbit_r89_c212 bl[212] br[212] wl[89] vdd gnd cell_6t
Xbit_r90_c212 bl[212] br[212] wl[90] vdd gnd cell_6t
Xbit_r91_c212 bl[212] br[212] wl[91] vdd gnd cell_6t
Xbit_r92_c212 bl[212] br[212] wl[92] vdd gnd cell_6t
Xbit_r93_c212 bl[212] br[212] wl[93] vdd gnd cell_6t
Xbit_r94_c212 bl[212] br[212] wl[94] vdd gnd cell_6t
Xbit_r95_c212 bl[212] br[212] wl[95] vdd gnd cell_6t
Xbit_r96_c212 bl[212] br[212] wl[96] vdd gnd cell_6t
Xbit_r97_c212 bl[212] br[212] wl[97] vdd gnd cell_6t
Xbit_r98_c212 bl[212] br[212] wl[98] vdd gnd cell_6t
Xbit_r99_c212 bl[212] br[212] wl[99] vdd gnd cell_6t
Xbit_r100_c212 bl[212] br[212] wl[100] vdd gnd cell_6t
Xbit_r101_c212 bl[212] br[212] wl[101] vdd gnd cell_6t
Xbit_r102_c212 bl[212] br[212] wl[102] vdd gnd cell_6t
Xbit_r103_c212 bl[212] br[212] wl[103] vdd gnd cell_6t
Xbit_r104_c212 bl[212] br[212] wl[104] vdd gnd cell_6t
Xbit_r105_c212 bl[212] br[212] wl[105] vdd gnd cell_6t
Xbit_r106_c212 bl[212] br[212] wl[106] vdd gnd cell_6t
Xbit_r107_c212 bl[212] br[212] wl[107] vdd gnd cell_6t
Xbit_r108_c212 bl[212] br[212] wl[108] vdd gnd cell_6t
Xbit_r109_c212 bl[212] br[212] wl[109] vdd gnd cell_6t
Xbit_r110_c212 bl[212] br[212] wl[110] vdd gnd cell_6t
Xbit_r111_c212 bl[212] br[212] wl[111] vdd gnd cell_6t
Xbit_r112_c212 bl[212] br[212] wl[112] vdd gnd cell_6t
Xbit_r113_c212 bl[212] br[212] wl[113] vdd gnd cell_6t
Xbit_r114_c212 bl[212] br[212] wl[114] vdd gnd cell_6t
Xbit_r115_c212 bl[212] br[212] wl[115] vdd gnd cell_6t
Xbit_r116_c212 bl[212] br[212] wl[116] vdd gnd cell_6t
Xbit_r117_c212 bl[212] br[212] wl[117] vdd gnd cell_6t
Xbit_r118_c212 bl[212] br[212] wl[118] vdd gnd cell_6t
Xbit_r119_c212 bl[212] br[212] wl[119] vdd gnd cell_6t
Xbit_r120_c212 bl[212] br[212] wl[120] vdd gnd cell_6t
Xbit_r121_c212 bl[212] br[212] wl[121] vdd gnd cell_6t
Xbit_r122_c212 bl[212] br[212] wl[122] vdd gnd cell_6t
Xbit_r123_c212 bl[212] br[212] wl[123] vdd gnd cell_6t
Xbit_r124_c212 bl[212] br[212] wl[124] vdd gnd cell_6t
Xbit_r125_c212 bl[212] br[212] wl[125] vdd gnd cell_6t
Xbit_r126_c212 bl[212] br[212] wl[126] vdd gnd cell_6t
Xbit_r127_c212 bl[212] br[212] wl[127] vdd gnd cell_6t
Xbit_r128_c212 bl[212] br[212] wl[128] vdd gnd cell_6t
Xbit_r129_c212 bl[212] br[212] wl[129] vdd gnd cell_6t
Xbit_r130_c212 bl[212] br[212] wl[130] vdd gnd cell_6t
Xbit_r131_c212 bl[212] br[212] wl[131] vdd gnd cell_6t
Xbit_r132_c212 bl[212] br[212] wl[132] vdd gnd cell_6t
Xbit_r133_c212 bl[212] br[212] wl[133] vdd gnd cell_6t
Xbit_r134_c212 bl[212] br[212] wl[134] vdd gnd cell_6t
Xbit_r135_c212 bl[212] br[212] wl[135] vdd gnd cell_6t
Xbit_r136_c212 bl[212] br[212] wl[136] vdd gnd cell_6t
Xbit_r137_c212 bl[212] br[212] wl[137] vdd gnd cell_6t
Xbit_r138_c212 bl[212] br[212] wl[138] vdd gnd cell_6t
Xbit_r139_c212 bl[212] br[212] wl[139] vdd gnd cell_6t
Xbit_r140_c212 bl[212] br[212] wl[140] vdd gnd cell_6t
Xbit_r141_c212 bl[212] br[212] wl[141] vdd gnd cell_6t
Xbit_r142_c212 bl[212] br[212] wl[142] vdd gnd cell_6t
Xbit_r143_c212 bl[212] br[212] wl[143] vdd gnd cell_6t
Xbit_r144_c212 bl[212] br[212] wl[144] vdd gnd cell_6t
Xbit_r145_c212 bl[212] br[212] wl[145] vdd gnd cell_6t
Xbit_r146_c212 bl[212] br[212] wl[146] vdd gnd cell_6t
Xbit_r147_c212 bl[212] br[212] wl[147] vdd gnd cell_6t
Xbit_r148_c212 bl[212] br[212] wl[148] vdd gnd cell_6t
Xbit_r149_c212 bl[212] br[212] wl[149] vdd gnd cell_6t
Xbit_r150_c212 bl[212] br[212] wl[150] vdd gnd cell_6t
Xbit_r151_c212 bl[212] br[212] wl[151] vdd gnd cell_6t
Xbit_r152_c212 bl[212] br[212] wl[152] vdd gnd cell_6t
Xbit_r153_c212 bl[212] br[212] wl[153] vdd gnd cell_6t
Xbit_r154_c212 bl[212] br[212] wl[154] vdd gnd cell_6t
Xbit_r155_c212 bl[212] br[212] wl[155] vdd gnd cell_6t
Xbit_r156_c212 bl[212] br[212] wl[156] vdd gnd cell_6t
Xbit_r157_c212 bl[212] br[212] wl[157] vdd gnd cell_6t
Xbit_r158_c212 bl[212] br[212] wl[158] vdd gnd cell_6t
Xbit_r159_c212 bl[212] br[212] wl[159] vdd gnd cell_6t
Xbit_r160_c212 bl[212] br[212] wl[160] vdd gnd cell_6t
Xbit_r161_c212 bl[212] br[212] wl[161] vdd gnd cell_6t
Xbit_r162_c212 bl[212] br[212] wl[162] vdd gnd cell_6t
Xbit_r163_c212 bl[212] br[212] wl[163] vdd gnd cell_6t
Xbit_r164_c212 bl[212] br[212] wl[164] vdd gnd cell_6t
Xbit_r165_c212 bl[212] br[212] wl[165] vdd gnd cell_6t
Xbit_r166_c212 bl[212] br[212] wl[166] vdd gnd cell_6t
Xbit_r167_c212 bl[212] br[212] wl[167] vdd gnd cell_6t
Xbit_r168_c212 bl[212] br[212] wl[168] vdd gnd cell_6t
Xbit_r169_c212 bl[212] br[212] wl[169] vdd gnd cell_6t
Xbit_r170_c212 bl[212] br[212] wl[170] vdd gnd cell_6t
Xbit_r171_c212 bl[212] br[212] wl[171] vdd gnd cell_6t
Xbit_r172_c212 bl[212] br[212] wl[172] vdd gnd cell_6t
Xbit_r173_c212 bl[212] br[212] wl[173] vdd gnd cell_6t
Xbit_r174_c212 bl[212] br[212] wl[174] vdd gnd cell_6t
Xbit_r175_c212 bl[212] br[212] wl[175] vdd gnd cell_6t
Xbit_r176_c212 bl[212] br[212] wl[176] vdd gnd cell_6t
Xbit_r177_c212 bl[212] br[212] wl[177] vdd gnd cell_6t
Xbit_r178_c212 bl[212] br[212] wl[178] vdd gnd cell_6t
Xbit_r179_c212 bl[212] br[212] wl[179] vdd gnd cell_6t
Xbit_r180_c212 bl[212] br[212] wl[180] vdd gnd cell_6t
Xbit_r181_c212 bl[212] br[212] wl[181] vdd gnd cell_6t
Xbit_r182_c212 bl[212] br[212] wl[182] vdd gnd cell_6t
Xbit_r183_c212 bl[212] br[212] wl[183] vdd gnd cell_6t
Xbit_r184_c212 bl[212] br[212] wl[184] vdd gnd cell_6t
Xbit_r185_c212 bl[212] br[212] wl[185] vdd gnd cell_6t
Xbit_r186_c212 bl[212] br[212] wl[186] vdd gnd cell_6t
Xbit_r187_c212 bl[212] br[212] wl[187] vdd gnd cell_6t
Xbit_r188_c212 bl[212] br[212] wl[188] vdd gnd cell_6t
Xbit_r189_c212 bl[212] br[212] wl[189] vdd gnd cell_6t
Xbit_r190_c212 bl[212] br[212] wl[190] vdd gnd cell_6t
Xbit_r191_c212 bl[212] br[212] wl[191] vdd gnd cell_6t
Xbit_r192_c212 bl[212] br[212] wl[192] vdd gnd cell_6t
Xbit_r193_c212 bl[212] br[212] wl[193] vdd gnd cell_6t
Xbit_r194_c212 bl[212] br[212] wl[194] vdd gnd cell_6t
Xbit_r195_c212 bl[212] br[212] wl[195] vdd gnd cell_6t
Xbit_r196_c212 bl[212] br[212] wl[196] vdd gnd cell_6t
Xbit_r197_c212 bl[212] br[212] wl[197] vdd gnd cell_6t
Xbit_r198_c212 bl[212] br[212] wl[198] vdd gnd cell_6t
Xbit_r199_c212 bl[212] br[212] wl[199] vdd gnd cell_6t
Xbit_r200_c212 bl[212] br[212] wl[200] vdd gnd cell_6t
Xbit_r201_c212 bl[212] br[212] wl[201] vdd gnd cell_6t
Xbit_r202_c212 bl[212] br[212] wl[202] vdd gnd cell_6t
Xbit_r203_c212 bl[212] br[212] wl[203] vdd gnd cell_6t
Xbit_r204_c212 bl[212] br[212] wl[204] vdd gnd cell_6t
Xbit_r205_c212 bl[212] br[212] wl[205] vdd gnd cell_6t
Xbit_r206_c212 bl[212] br[212] wl[206] vdd gnd cell_6t
Xbit_r207_c212 bl[212] br[212] wl[207] vdd gnd cell_6t
Xbit_r208_c212 bl[212] br[212] wl[208] vdd gnd cell_6t
Xbit_r209_c212 bl[212] br[212] wl[209] vdd gnd cell_6t
Xbit_r210_c212 bl[212] br[212] wl[210] vdd gnd cell_6t
Xbit_r211_c212 bl[212] br[212] wl[211] vdd gnd cell_6t
Xbit_r212_c212 bl[212] br[212] wl[212] vdd gnd cell_6t
Xbit_r213_c212 bl[212] br[212] wl[213] vdd gnd cell_6t
Xbit_r214_c212 bl[212] br[212] wl[214] vdd gnd cell_6t
Xbit_r215_c212 bl[212] br[212] wl[215] vdd gnd cell_6t
Xbit_r216_c212 bl[212] br[212] wl[216] vdd gnd cell_6t
Xbit_r217_c212 bl[212] br[212] wl[217] vdd gnd cell_6t
Xbit_r218_c212 bl[212] br[212] wl[218] vdd gnd cell_6t
Xbit_r219_c212 bl[212] br[212] wl[219] vdd gnd cell_6t
Xbit_r220_c212 bl[212] br[212] wl[220] vdd gnd cell_6t
Xbit_r221_c212 bl[212] br[212] wl[221] vdd gnd cell_6t
Xbit_r222_c212 bl[212] br[212] wl[222] vdd gnd cell_6t
Xbit_r223_c212 bl[212] br[212] wl[223] vdd gnd cell_6t
Xbit_r224_c212 bl[212] br[212] wl[224] vdd gnd cell_6t
Xbit_r225_c212 bl[212] br[212] wl[225] vdd gnd cell_6t
Xbit_r226_c212 bl[212] br[212] wl[226] vdd gnd cell_6t
Xbit_r227_c212 bl[212] br[212] wl[227] vdd gnd cell_6t
Xbit_r228_c212 bl[212] br[212] wl[228] vdd gnd cell_6t
Xbit_r229_c212 bl[212] br[212] wl[229] vdd gnd cell_6t
Xbit_r230_c212 bl[212] br[212] wl[230] vdd gnd cell_6t
Xbit_r231_c212 bl[212] br[212] wl[231] vdd gnd cell_6t
Xbit_r232_c212 bl[212] br[212] wl[232] vdd gnd cell_6t
Xbit_r233_c212 bl[212] br[212] wl[233] vdd gnd cell_6t
Xbit_r234_c212 bl[212] br[212] wl[234] vdd gnd cell_6t
Xbit_r235_c212 bl[212] br[212] wl[235] vdd gnd cell_6t
Xbit_r236_c212 bl[212] br[212] wl[236] vdd gnd cell_6t
Xbit_r237_c212 bl[212] br[212] wl[237] vdd gnd cell_6t
Xbit_r238_c212 bl[212] br[212] wl[238] vdd gnd cell_6t
Xbit_r239_c212 bl[212] br[212] wl[239] vdd gnd cell_6t
Xbit_r240_c212 bl[212] br[212] wl[240] vdd gnd cell_6t
Xbit_r241_c212 bl[212] br[212] wl[241] vdd gnd cell_6t
Xbit_r242_c212 bl[212] br[212] wl[242] vdd gnd cell_6t
Xbit_r243_c212 bl[212] br[212] wl[243] vdd gnd cell_6t
Xbit_r244_c212 bl[212] br[212] wl[244] vdd gnd cell_6t
Xbit_r245_c212 bl[212] br[212] wl[245] vdd gnd cell_6t
Xbit_r246_c212 bl[212] br[212] wl[246] vdd gnd cell_6t
Xbit_r247_c212 bl[212] br[212] wl[247] vdd gnd cell_6t
Xbit_r248_c212 bl[212] br[212] wl[248] vdd gnd cell_6t
Xbit_r249_c212 bl[212] br[212] wl[249] vdd gnd cell_6t
Xbit_r250_c212 bl[212] br[212] wl[250] vdd gnd cell_6t
Xbit_r251_c212 bl[212] br[212] wl[251] vdd gnd cell_6t
Xbit_r252_c212 bl[212] br[212] wl[252] vdd gnd cell_6t
Xbit_r253_c212 bl[212] br[212] wl[253] vdd gnd cell_6t
Xbit_r254_c212 bl[212] br[212] wl[254] vdd gnd cell_6t
Xbit_r255_c212 bl[212] br[212] wl[255] vdd gnd cell_6t
Xbit_r0_c213 bl[213] br[213] wl[0] vdd gnd cell_6t
Xbit_r1_c213 bl[213] br[213] wl[1] vdd gnd cell_6t
Xbit_r2_c213 bl[213] br[213] wl[2] vdd gnd cell_6t
Xbit_r3_c213 bl[213] br[213] wl[3] vdd gnd cell_6t
Xbit_r4_c213 bl[213] br[213] wl[4] vdd gnd cell_6t
Xbit_r5_c213 bl[213] br[213] wl[5] vdd gnd cell_6t
Xbit_r6_c213 bl[213] br[213] wl[6] vdd gnd cell_6t
Xbit_r7_c213 bl[213] br[213] wl[7] vdd gnd cell_6t
Xbit_r8_c213 bl[213] br[213] wl[8] vdd gnd cell_6t
Xbit_r9_c213 bl[213] br[213] wl[9] vdd gnd cell_6t
Xbit_r10_c213 bl[213] br[213] wl[10] vdd gnd cell_6t
Xbit_r11_c213 bl[213] br[213] wl[11] vdd gnd cell_6t
Xbit_r12_c213 bl[213] br[213] wl[12] vdd gnd cell_6t
Xbit_r13_c213 bl[213] br[213] wl[13] vdd gnd cell_6t
Xbit_r14_c213 bl[213] br[213] wl[14] vdd gnd cell_6t
Xbit_r15_c213 bl[213] br[213] wl[15] vdd gnd cell_6t
Xbit_r16_c213 bl[213] br[213] wl[16] vdd gnd cell_6t
Xbit_r17_c213 bl[213] br[213] wl[17] vdd gnd cell_6t
Xbit_r18_c213 bl[213] br[213] wl[18] vdd gnd cell_6t
Xbit_r19_c213 bl[213] br[213] wl[19] vdd gnd cell_6t
Xbit_r20_c213 bl[213] br[213] wl[20] vdd gnd cell_6t
Xbit_r21_c213 bl[213] br[213] wl[21] vdd gnd cell_6t
Xbit_r22_c213 bl[213] br[213] wl[22] vdd gnd cell_6t
Xbit_r23_c213 bl[213] br[213] wl[23] vdd gnd cell_6t
Xbit_r24_c213 bl[213] br[213] wl[24] vdd gnd cell_6t
Xbit_r25_c213 bl[213] br[213] wl[25] vdd gnd cell_6t
Xbit_r26_c213 bl[213] br[213] wl[26] vdd gnd cell_6t
Xbit_r27_c213 bl[213] br[213] wl[27] vdd gnd cell_6t
Xbit_r28_c213 bl[213] br[213] wl[28] vdd gnd cell_6t
Xbit_r29_c213 bl[213] br[213] wl[29] vdd gnd cell_6t
Xbit_r30_c213 bl[213] br[213] wl[30] vdd gnd cell_6t
Xbit_r31_c213 bl[213] br[213] wl[31] vdd gnd cell_6t
Xbit_r32_c213 bl[213] br[213] wl[32] vdd gnd cell_6t
Xbit_r33_c213 bl[213] br[213] wl[33] vdd gnd cell_6t
Xbit_r34_c213 bl[213] br[213] wl[34] vdd gnd cell_6t
Xbit_r35_c213 bl[213] br[213] wl[35] vdd gnd cell_6t
Xbit_r36_c213 bl[213] br[213] wl[36] vdd gnd cell_6t
Xbit_r37_c213 bl[213] br[213] wl[37] vdd gnd cell_6t
Xbit_r38_c213 bl[213] br[213] wl[38] vdd gnd cell_6t
Xbit_r39_c213 bl[213] br[213] wl[39] vdd gnd cell_6t
Xbit_r40_c213 bl[213] br[213] wl[40] vdd gnd cell_6t
Xbit_r41_c213 bl[213] br[213] wl[41] vdd gnd cell_6t
Xbit_r42_c213 bl[213] br[213] wl[42] vdd gnd cell_6t
Xbit_r43_c213 bl[213] br[213] wl[43] vdd gnd cell_6t
Xbit_r44_c213 bl[213] br[213] wl[44] vdd gnd cell_6t
Xbit_r45_c213 bl[213] br[213] wl[45] vdd gnd cell_6t
Xbit_r46_c213 bl[213] br[213] wl[46] vdd gnd cell_6t
Xbit_r47_c213 bl[213] br[213] wl[47] vdd gnd cell_6t
Xbit_r48_c213 bl[213] br[213] wl[48] vdd gnd cell_6t
Xbit_r49_c213 bl[213] br[213] wl[49] vdd gnd cell_6t
Xbit_r50_c213 bl[213] br[213] wl[50] vdd gnd cell_6t
Xbit_r51_c213 bl[213] br[213] wl[51] vdd gnd cell_6t
Xbit_r52_c213 bl[213] br[213] wl[52] vdd gnd cell_6t
Xbit_r53_c213 bl[213] br[213] wl[53] vdd gnd cell_6t
Xbit_r54_c213 bl[213] br[213] wl[54] vdd gnd cell_6t
Xbit_r55_c213 bl[213] br[213] wl[55] vdd gnd cell_6t
Xbit_r56_c213 bl[213] br[213] wl[56] vdd gnd cell_6t
Xbit_r57_c213 bl[213] br[213] wl[57] vdd gnd cell_6t
Xbit_r58_c213 bl[213] br[213] wl[58] vdd gnd cell_6t
Xbit_r59_c213 bl[213] br[213] wl[59] vdd gnd cell_6t
Xbit_r60_c213 bl[213] br[213] wl[60] vdd gnd cell_6t
Xbit_r61_c213 bl[213] br[213] wl[61] vdd gnd cell_6t
Xbit_r62_c213 bl[213] br[213] wl[62] vdd gnd cell_6t
Xbit_r63_c213 bl[213] br[213] wl[63] vdd gnd cell_6t
Xbit_r64_c213 bl[213] br[213] wl[64] vdd gnd cell_6t
Xbit_r65_c213 bl[213] br[213] wl[65] vdd gnd cell_6t
Xbit_r66_c213 bl[213] br[213] wl[66] vdd gnd cell_6t
Xbit_r67_c213 bl[213] br[213] wl[67] vdd gnd cell_6t
Xbit_r68_c213 bl[213] br[213] wl[68] vdd gnd cell_6t
Xbit_r69_c213 bl[213] br[213] wl[69] vdd gnd cell_6t
Xbit_r70_c213 bl[213] br[213] wl[70] vdd gnd cell_6t
Xbit_r71_c213 bl[213] br[213] wl[71] vdd gnd cell_6t
Xbit_r72_c213 bl[213] br[213] wl[72] vdd gnd cell_6t
Xbit_r73_c213 bl[213] br[213] wl[73] vdd gnd cell_6t
Xbit_r74_c213 bl[213] br[213] wl[74] vdd gnd cell_6t
Xbit_r75_c213 bl[213] br[213] wl[75] vdd gnd cell_6t
Xbit_r76_c213 bl[213] br[213] wl[76] vdd gnd cell_6t
Xbit_r77_c213 bl[213] br[213] wl[77] vdd gnd cell_6t
Xbit_r78_c213 bl[213] br[213] wl[78] vdd gnd cell_6t
Xbit_r79_c213 bl[213] br[213] wl[79] vdd gnd cell_6t
Xbit_r80_c213 bl[213] br[213] wl[80] vdd gnd cell_6t
Xbit_r81_c213 bl[213] br[213] wl[81] vdd gnd cell_6t
Xbit_r82_c213 bl[213] br[213] wl[82] vdd gnd cell_6t
Xbit_r83_c213 bl[213] br[213] wl[83] vdd gnd cell_6t
Xbit_r84_c213 bl[213] br[213] wl[84] vdd gnd cell_6t
Xbit_r85_c213 bl[213] br[213] wl[85] vdd gnd cell_6t
Xbit_r86_c213 bl[213] br[213] wl[86] vdd gnd cell_6t
Xbit_r87_c213 bl[213] br[213] wl[87] vdd gnd cell_6t
Xbit_r88_c213 bl[213] br[213] wl[88] vdd gnd cell_6t
Xbit_r89_c213 bl[213] br[213] wl[89] vdd gnd cell_6t
Xbit_r90_c213 bl[213] br[213] wl[90] vdd gnd cell_6t
Xbit_r91_c213 bl[213] br[213] wl[91] vdd gnd cell_6t
Xbit_r92_c213 bl[213] br[213] wl[92] vdd gnd cell_6t
Xbit_r93_c213 bl[213] br[213] wl[93] vdd gnd cell_6t
Xbit_r94_c213 bl[213] br[213] wl[94] vdd gnd cell_6t
Xbit_r95_c213 bl[213] br[213] wl[95] vdd gnd cell_6t
Xbit_r96_c213 bl[213] br[213] wl[96] vdd gnd cell_6t
Xbit_r97_c213 bl[213] br[213] wl[97] vdd gnd cell_6t
Xbit_r98_c213 bl[213] br[213] wl[98] vdd gnd cell_6t
Xbit_r99_c213 bl[213] br[213] wl[99] vdd gnd cell_6t
Xbit_r100_c213 bl[213] br[213] wl[100] vdd gnd cell_6t
Xbit_r101_c213 bl[213] br[213] wl[101] vdd gnd cell_6t
Xbit_r102_c213 bl[213] br[213] wl[102] vdd gnd cell_6t
Xbit_r103_c213 bl[213] br[213] wl[103] vdd gnd cell_6t
Xbit_r104_c213 bl[213] br[213] wl[104] vdd gnd cell_6t
Xbit_r105_c213 bl[213] br[213] wl[105] vdd gnd cell_6t
Xbit_r106_c213 bl[213] br[213] wl[106] vdd gnd cell_6t
Xbit_r107_c213 bl[213] br[213] wl[107] vdd gnd cell_6t
Xbit_r108_c213 bl[213] br[213] wl[108] vdd gnd cell_6t
Xbit_r109_c213 bl[213] br[213] wl[109] vdd gnd cell_6t
Xbit_r110_c213 bl[213] br[213] wl[110] vdd gnd cell_6t
Xbit_r111_c213 bl[213] br[213] wl[111] vdd gnd cell_6t
Xbit_r112_c213 bl[213] br[213] wl[112] vdd gnd cell_6t
Xbit_r113_c213 bl[213] br[213] wl[113] vdd gnd cell_6t
Xbit_r114_c213 bl[213] br[213] wl[114] vdd gnd cell_6t
Xbit_r115_c213 bl[213] br[213] wl[115] vdd gnd cell_6t
Xbit_r116_c213 bl[213] br[213] wl[116] vdd gnd cell_6t
Xbit_r117_c213 bl[213] br[213] wl[117] vdd gnd cell_6t
Xbit_r118_c213 bl[213] br[213] wl[118] vdd gnd cell_6t
Xbit_r119_c213 bl[213] br[213] wl[119] vdd gnd cell_6t
Xbit_r120_c213 bl[213] br[213] wl[120] vdd gnd cell_6t
Xbit_r121_c213 bl[213] br[213] wl[121] vdd gnd cell_6t
Xbit_r122_c213 bl[213] br[213] wl[122] vdd gnd cell_6t
Xbit_r123_c213 bl[213] br[213] wl[123] vdd gnd cell_6t
Xbit_r124_c213 bl[213] br[213] wl[124] vdd gnd cell_6t
Xbit_r125_c213 bl[213] br[213] wl[125] vdd gnd cell_6t
Xbit_r126_c213 bl[213] br[213] wl[126] vdd gnd cell_6t
Xbit_r127_c213 bl[213] br[213] wl[127] vdd gnd cell_6t
Xbit_r128_c213 bl[213] br[213] wl[128] vdd gnd cell_6t
Xbit_r129_c213 bl[213] br[213] wl[129] vdd gnd cell_6t
Xbit_r130_c213 bl[213] br[213] wl[130] vdd gnd cell_6t
Xbit_r131_c213 bl[213] br[213] wl[131] vdd gnd cell_6t
Xbit_r132_c213 bl[213] br[213] wl[132] vdd gnd cell_6t
Xbit_r133_c213 bl[213] br[213] wl[133] vdd gnd cell_6t
Xbit_r134_c213 bl[213] br[213] wl[134] vdd gnd cell_6t
Xbit_r135_c213 bl[213] br[213] wl[135] vdd gnd cell_6t
Xbit_r136_c213 bl[213] br[213] wl[136] vdd gnd cell_6t
Xbit_r137_c213 bl[213] br[213] wl[137] vdd gnd cell_6t
Xbit_r138_c213 bl[213] br[213] wl[138] vdd gnd cell_6t
Xbit_r139_c213 bl[213] br[213] wl[139] vdd gnd cell_6t
Xbit_r140_c213 bl[213] br[213] wl[140] vdd gnd cell_6t
Xbit_r141_c213 bl[213] br[213] wl[141] vdd gnd cell_6t
Xbit_r142_c213 bl[213] br[213] wl[142] vdd gnd cell_6t
Xbit_r143_c213 bl[213] br[213] wl[143] vdd gnd cell_6t
Xbit_r144_c213 bl[213] br[213] wl[144] vdd gnd cell_6t
Xbit_r145_c213 bl[213] br[213] wl[145] vdd gnd cell_6t
Xbit_r146_c213 bl[213] br[213] wl[146] vdd gnd cell_6t
Xbit_r147_c213 bl[213] br[213] wl[147] vdd gnd cell_6t
Xbit_r148_c213 bl[213] br[213] wl[148] vdd gnd cell_6t
Xbit_r149_c213 bl[213] br[213] wl[149] vdd gnd cell_6t
Xbit_r150_c213 bl[213] br[213] wl[150] vdd gnd cell_6t
Xbit_r151_c213 bl[213] br[213] wl[151] vdd gnd cell_6t
Xbit_r152_c213 bl[213] br[213] wl[152] vdd gnd cell_6t
Xbit_r153_c213 bl[213] br[213] wl[153] vdd gnd cell_6t
Xbit_r154_c213 bl[213] br[213] wl[154] vdd gnd cell_6t
Xbit_r155_c213 bl[213] br[213] wl[155] vdd gnd cell_6t
Xbit_r156_c213 bl[213] br[213] wl[156] vdd gnd cell_6t
Xbit_r157_c213 bl[213] br[213] wl[157] vdd gnd cell_6t
Xbit_r158_c213 bl[213] br[213] wl[158] vdd gnd cell_6t
Xbit_r159_c213 bl[213] br[213] wl[159] vdd gnd cell_6t
Xbit_r160_c213 bl[213] br[213] wl[160] vdd gnd cell_6t
Xbit_r161_c213 bl[213] br[213] wl[161] vdd gnd cell_6t
Xbit_r162_c213 bl[213] br[213] wl[162] vdd gnd cell_6t
Xbit_r163_c213 bl[213] br[213] wl[163] vdd gnd cell_6t
Xbit_r164_c213 bl[213] br[213] wl[164] vdd gnd cell_6t
Xbit_r165_c213 bl[213] br[213] wl[165] vdd gnd cell_6t
Xbit_r166_c213 bl[213] br[213] wl[166] vdd gnd cell_6t
Xbit_r167_c213 bl[213] br[213] wl[167] vdd gnd cell_6t
Xbit_r168_c213 bl[213] br[213] wl[168] vdd gnd cell_6t
Xbit_r169_c213 bl[213] br[213] wl[169] vdd gnd cell_6t
Xbit_r170_c213 bl[213] br[213] wl[170] vdd gnd cell_6t
Xbit_r171_c213 bl[213] br[213] wl[171] vdd gnd cell_6t
Xbit_r172_c213 bl[213] br[213] wl[172] vdd gnd cell_6t
Xbit_r173_c213 bl[213] br[213] wl[173] vdd gnd cell_6t
Xbit_r174_c213 bl[213] br[213] wl[174] vdd gnd cell_6t
Xbit_r175_c213 bl[213] br[213] wl[175] vdd gnd cell_6t
Xbit_r176_c213 bl[213] br[213] wl[176] vdd gnd cell_6t
Xbit_r177_c213 bl[213] br[213] wl[177] vdd gnd cell_6t
Xbit_r178_c213 bl[213] br[213] wl[178] vdd gnd cell_6t
Xbit_r179_c213 bl[213] br[213] wl[179] vdd gnd cell_6t
Xbit_r180_c213 bl[213] br[213] wl[180] vdd gnd cell_6t
Xbit_r181_c213 bl[213] br[213] wl[181] vdd gnd cell_6t
Xbit_r182_c213 bl[213] br[213] wl[182] vdd gnd cell_6t
Xbit_r183_c213 bl[213] br[213] wl[183] vdd gnd cell_6t
Xbit_r184_c213 bl[213] br[213] wl[184] vdd gnd cell_6t
Xbit_r185_c213 bl[213] br[213] wl[185] vdd gnd cell_6t
Xbit_r186_c213 bl[213] br[213] wl[186] vdd gnd cell_6t
Xbit_r187_c213 bl[213] br[213] wl[187] vdd gnd cell_6t
Xbit_r188_c213 bl[213] br[213] wl[188] vdd gnd cell_6t
Xbit_r189_c213 bl[213] br[213] wl[189] vdd gnd cell_6t
Xbit_r190_c213 bl[213] br[213] wl[190] vdd gnd cell_6t
Xbit_r191_c213 bl[213] br[213] wl[191] vdd gnd cell_6t
Xbit_r192_c213 bl[213] br[213] wl[192] vdd gnd cell_6t
Xbit_r193_c213 bl[213] br[213] wl[193] vdd gnd cell_6t
Xbit_r194_c213 bl[213] br[213] wl[194] vdd gnd cell_6t
Xbit_r195_c213 bl[213] br[213] wl[195] vdd gnd cell_6t
Xbit_r196_c213 bl[213] br[213] wl[196] vdd gnd cell_6t
Xbit_r197_c213 bl[213] br[213] wl[197] vdd gnd cell_6t
Xbit_r198_c213 bl[213] br[213] wl[198] vdd gnd cell_6t
Xbit_r199_c213 bl[213] br[213] wl[199] vdd gnd cell_6t
Xbit_r200_c213 bl[213] br[213] wl[200] vdd gnd cell_6t
Xbit_r201_c213 bl[213] br[213] wl[201] vdd gnd cell_6t
Xbit_r202_c213 bl[213] br[213] wl[202] vdd gnd cell_6t
Xbit_r203_c213 bl[213] br[213] wl[203] vdd gnd cell_6t
Xbit_r204_c213 bl[213] br[213] wl[204] vdd gnd cell_6t
Xbit_r205_c213 bl[213] br[213] wl[205] vdd gnd cell_6t
Xbit_r206_c213 bl[213] br[213] wl[206] vdd gnd cell_6t
Xbit_r207_c213 bl[213] br[213] wl[207] vdd gnd cell_6t
Xbit_r208_c213 bl[213] br[213] wl[208] vdd gnd cell_6t
Xbit_r209_c213 bl[213] br[213] wl[209] vdd gnd cell_6t
Xbit_r210_c213 bl[213] br[213] wl[210] vdd gnd cell_6t
Xbit_r211_c213 bl[213] br[213] wl[211] vdd gnd cell_6t
Xbit_r212_c213 bl[213] br[213] wl[212] vdd gnd cell_6t
Xbit_r213_c213 bl[213] br[213] wl[213] vdd gnd cell_6t
Xbit_r214_c213 bl[213] br[213] wl[214] vdd gnd cell_6t
Xbit_r215_c213 bl[213] br[213] wl[215] vdd gnd cell_6t
Xbit_r216_c213 bl[213] br[213] wl[216] vdd gnd cell_6t
Xbit_r217_c213 bl[213] br[213] wl[217] vdd gnd cell_6t
Xbit_r218_c213 bl[213] br[213] wl[218] vdd gnd cell_6t
Xbit_r219_c213 bl[213] br[213] wl[219] vdd gnd cell_6t
Xbit_r220_c213 bl[213] br[213] wl[220] vdd gnd cell_6t
Xbit_r221_c213 bl[213] br[213] wl[221] vdd gnd cell_6t
Xbit_r222_c213 bl[213] br[213] wl[222] vdd gnd cell_6t
Xbit_r223_c213 bl[213] br[213] wl[223] vdd gnd cell_6t
Xbit_r224_c213 bl[213] br[213] wl[224] vdd gnd cell_6t
Xbit_r225_c213 bl[213] br[213] wl[225] vdd gnd cell_6t
Xbit_r226_c213 bl[213] br[213] wl[226] vdd gnd cell_6t
Xbit_r227_c213 bl[213] br[213] wl[227] vdd gnd cell_6t
Xbit_r228_c213 bl[213] br[213] wl[228] vdd gnd cell_6t
Xbit_r229_c213 bl[213] br[213] wl[229] vdd gnd cell_6t
Xbit_r230_c213 bl[213] br[213] wl[230] vdd gnd cell_6t
Xbit_r231_c213 bl[213] br[213] wl[231] vdd gnd cell_6t
Xbit_r232_c213 bl[213] br[213] wl[232] vdd gnd cell_6t
Xbit_r233_c213 bl[213] br[213] wl[233] vdd gnd cell_6t
Xbit_r234_c213 bl[213] br[213] wl[234] vdd gnd cell_6t
Xbit_r235_c213 bl[213] br[213] wl[235] vdd gnd cell_6t
Xbit_r236_c213 bl[213] br[213] wl[236] vdd gnd cell_6t
Xbit_r237_c213 bl[213] br[213] wl[237] vdd gnd cell_6t
Xbit_r238_c213 bl[213] br[213] wl[238] vdd gnd cell_6t
Xbit_r239_c213 bl[213] br[213] wl[239] vdd gnd cell_6t
Xbit_r240_c213 bl[213] br[213] wl[240] vdd gnd cell_6t
Xbit_r241_c213 bl[213] br[213] wl[241] vdd gnd cell_6t
Xbit_r242_c213 bl[213] br[213] wl[242] vdd gnd cell_6t
Xbit_r243_c213 bl[213] br[213] wl[243] vdd gnd cell_6t
Xbit_r244_c213 bl[213] br[213] wl[244] vdd gnd cell_6t
Xbit_r245_c213 bl[213] br[213] wl[245] vdd gnd cell_6t
Xbit_r246_c213 bl[213] br[213] wl[246] vdd gnd cell_6t
Xbit_r247_c213 bl[213] br[213] wl[247] vdd gnd cell_6t
Xbit_r248_c213 bl[213] br[213] wl[248] vdd gnd cell_6t
Xbit_r249_c213 bl[213] br[213] wl[249] vdd gnd cell_6t
Xbit_r250_c213 bl[213] br[213] wl[250] vdd gnd cell_6t
Xbit_r251_c213 bl[213] br[213] wl[251] vdd gnd cell_6t
Xbit_r252_c213 bl[213] br[213] wl[252] vdd gnd cell_6t
Xbit_r253_c213 bl[213] br[213] wl[253] vdd gnd cell_6t
Xbit_r254_c213 bl[213] br[213] wl[254] vdd gnd cell_6t
Xbit_r255_c213 bl[213] br[213] wl[255] vdd gnd cell_6t
Xbit_r0_c214 bl[214] br[214] wl[0] vdd gnd cell_6t
Xbit_r1_c214 bl[214] br[214] wl[1] vdd gnd cell_6t
Xbit_r2_c214 bl[214] br[214] wl[2] vdd gnd cell_6t
Xbit_r3_c214 bl[214] br[214] wl[3] vdd gnd cell_6t
Xbit_r4_c214 bl[214] br[214] wl[4] vdd gnd cell_6t
Xbit_r5_c214 bl[214] br[214] wl[5] vdd gnd cell_6t
Xbit_r6_c214 bl[214] br[214] wl[6] vdd gnd cell_6t
Xbit_r7_c214 bl[214] br[214] wl[7] vdd gnd cell_6t
Xbit_r8_c214 bl[214] br[214] wl[8] vdd gnd cell_6t
Xbit_r9_c214 bl[214] br[214] wl[9] vdd gnd cell_6t
Xbit_r10_c214 bl[214] br[214] wl[10] vdd gnd cell_6t
Xbit_r11_c214 bl[214] br[214] wl[11] vdd gnd cell_6t
Xbit_r12_c214 bl[214] br[214] wl[12] vdd gnd cell_6t
Xbit_r13_c214 bl[214] br[214] wl[13] vdd gnd cell_6t
Xbit_r14_c214 bl[214] br[214] wl[14] vdd gnd cell_6t
Xbit_r15_c214 bl[214] br[214] wl[15] vdd gnd cell_6t
Xbit_r16_c214 bl[214] br[214] wl[16] vdd gnd cell_6t
Xbit_r17_c214 bl[214] br[214] wl[17] vdd gnd cell_6t
Xbit_r18_c214 bl[214] br[214] wl[18] vdd gnd cell_6t
Xbit_r19_c214 bl[214] br[214] wl[19] vdd gnd cell_6t
Xbit_r20_c214 bl[214] br[214] wl[20] vdd gnd cell_6t
Xbit_r21_c214 bl[214] br[214] wl[21] vdd gnd cell_6t
Xbit_r22_c214 bl[214] br[214] wl[22] vdd gnd cell_6t
Xbit_r23_c214 bl[214] br[214] wl[23] vdd gnd cell_6t
Xbit_r24_c214 bl[214] br[214] wl[24] vdd gnd cell_6t
Xbit_r25_c214 bl[214] br[214] wl[25] vdd gnd cell_6t
Xbit_r26_c214 bl[214] br[214] wl[26] vdd gnd cell_6t
Xbit_r27_c214 bl[214] br[214] wl[27] vdd gnd cell_6t
Xbit_r28_c214 bl[214] br[214] wl[28] vdd gnd cell_6t
Xbit_r29_c214 bl[214] br[214] wl[29] vdd gnd cell_6t
Xbit_r30_c214 bl[214] br[214] wl[30] vdd gnd cell_6t
Xbit_r31_c214 bl[214] br[214] wl[31] vdd gnd cell_6t
Xbit_r32_c214 bl[214] br[214] wl[32] vdd gnd cell_6t
Xbit_r33_c214 bl[214] br[214] wl[33] vdd gnd cell_6t
Xbit_r34_c214 bl[214] br[214] wl[34] vdd gnd cell_6t
Xbit_r35_c214 bl[214] br[214] wl[35] vdd gnd cell_6t
Xbit_r36_c214 bl[214] br[214] wl[36] vdd gnd cell_6t
Xbit_r37_c214 bl[214] br[214] wl[37] vdd gnd cell_6t
Xbit_r38_c214 bl[214] br[214] wl[38] vdd gnd cell_6t
Xbit_r39_c214 bl[214] br[214] wl[39] vdd gnd cell_6t
Xbit_r40_c214 bl[214] br[214] wl[40] vdd gnd cell_6t
Xbit_r41_c214 bl[214] br[214] wl[41] vdd gnd cell_6t
Xbit_r42_c214 bl[214] br[214] wl[42] vdd gnd cell_6t
Xbit_r43_c214 bl[214] br[214] wl[43] vdd gnd cell_6t
Xbit_r44_c214 bl[214] br[214] wl[44] vdd gnd cell_6t
Xbit_r45_c214 bl[214] br[214] wl[45] vdd gnd cell_6t
Xbit_r46_c214 bl[214] br[214] wl[46] vdd gnd cell_6t
Xbit_r47_c214 bl[214] br[214] wl[47] vdd gnd cell_6t
Xbit_r48_c214 bl[214] br[214] wl[48] vdd gnd cell_6t
Xbit_r49_c214 bl[214] br[214] wl[49] vdd gnd cell_6t
Xbit_r50_c214 bl[214] br[214] wl[50] vdd gnd cell_6t
Xbit_r51_c214 bl[214] br[214] wl[51] vdd gnd cell_6t
Xbit_r52_c214 bl[214] br[214] wl[52] vdd gnd cell_6t
Xbit_r53_c214 bl[214] br[214] wl[53] vdd gnd cell_6t
Xbit_r54_c214 bl[214] br[214] wl[54] vdd gnd cell_6t
Xbit_r55_c214 bl[214] br[214] wl[55] vdd gnd cell_6t
Xbit_r56_c214 bl[214] br[214] wl[56] vdd gnd cell_6t
Xbit_r57_c214 bl[214] br[214] wl[57] vdd gnd cell_6t
Xbit_r58_c214 bl[214] br[214] wl[58] vdd gnd cell_6t
Xbit_r59_c214 bl[214] br[214] wl[59] vdd gnd cell_6t
Xbit_r60_c214 bl[214] br[214] wl[60] vdd gnd cell_6t
Xbit_r61_c214 bl[214] br[214] wl[61] vdd gnd cell_6t
Xbit_r62_c214 bl[214] br[214] wl[62] vdd gnd cell_6t
Xbit_r63_c214 bl[214] br[214] wl[63] vdd gnd cell_6t
Xbit_r64_c214 bl[214] br[214] wl[64] vdd gnd cell_6t
Xbit_r65_c214 bl[214] br[214] wl[65] vdd gnd cell_6t
Xbit_r66_c214 bl[214] br[214] wl[66] vdd gnd cell_6t
Xbit_r67_c214 bl[214] br[214] wl[67] vdd gnd cell_6t
Xbit_r68_c214 bl[214] br[214] wl[68] vdd gnd cell_6t
Xbit_r69_c214 bl[214] br[214] wl[69] vdd gnd cell_6t
Xbit_r70_c214 bl[214] br[214] wl[70] vdd gnd cell_6t
Xbit_r71_c214 bl[214] br[214] wl[71] vdd gnd cell_6t
Xbit_r72_c214 bl[214] br[214] wl[72] vdd gnd cell_6t
Xbit_r73_c214 bl[214] br[214] wl[73] vdd gnd cell_6t
Xbit_r74_c214 bl[214] br[214] wl[74] vdd gnd cell_6t
Xbit_r75_c214 bl[214] br[214] wl[75] vdd gnd cell_6t
Xbit_r76_c214 bl[214] br[214] wl[76] vdd gnd cell_6t
Xbit_r77_c214 bl[214] br[214] wl[77] vdd gnd cell_6t
Xbit_r78_c214 bl[214] br[214] wl[78] vdd gnd cell_6t
Xbit_r79_c214 bl[214] br[214] wl[79] vdd gnd cell_6t
Xbit_r80_c214 bl[214] br[214] wl[80] vdd gnd cell_6t
Xbit_r81_c214 bl[214] br[214] wl[81] vdd gnd cell_6t
Xbit_r82_c214 bl[214] br[214] wl[82] vdd gnd cell_6t
Xbit_r83_c214 bl[214] br[214] wl[83] vdd gnd cell_6t
Xbit_r84_c214 bl[214] br[214] wl[84] vdd gnd cell_6t
Xbit_r85_c214 bl[214] br[214] wl[85] vdd gnd cell_6t
Xbit_r86_c214 bl[214] br[214] wl[86] vdd gnd cell_6t
Xbit_r87_c214 bl[214] br[214] wl[87] vdd gnd cell_6t
Xbit_r88_c214 bl[214] br[214] wl[88] vdd gnd cell_6t
Xbit_r89_c214 bl[214] br[214] wl[89] vdd gnd cell_6t
Xbit_r90_c214 bl[214] br[214] wl[90] vdd gnd cell_6t
Xbit_r91_c214 bl[214] br[214] wl[91] vdd gnd cell_6t
Xbit_r92_c214 bl[214] br[214] wl[92] vdd gnd cell_6t
Xbit_r93_c214 bl[214] br[214] wl[93] vdd gnd cell_6t
Xbit_r94_c214 bl[214] br[214] wl[94] vdd gnd cell_6t
Xbit_r95_c214 bl[214] br[214] wl[95] vdd gnd cell_6t
Xbit_r96_c214 bl[214] br[214] wl[96] vdd gnd cell_6t
Xbit_r97_c214 bl[214] br[214] wl[97] vdd gnd cell_6t
Xbit_r98_c214 bl[214] br[214] wl[98] vdd gnd cell_6t
Xbit_r99_c214 bl[214] br[214] wl[99] vdd gnd cell_6t
Xbit_r100_c214 bl[214] br[214] wl[100] vdd gnd cell_6t
Xbit_r101_c214 bl[214] br[214] wl[101] vdd gnd cell_6t
Xbit_r102_c214 bl[214] br[214] wl[102] vdd gnd cell_6t
Xbit_r103_c214 bl[214] br[214] wl[103] vdd gnd cell_6t
Xbit_r104_c214 bl[214] br[214] wl[104] vdd gnd cell_6t
Xbit_r105_c214 bl[214] br[214] wl[105] vdd gnd cell_6t
Xbit_r106_c214 bl[214] br[214] wl[106] vdd gnd cell_6t
Xbit_r107_c214 bl[214] br[214] wl[107] vdd gnd cell_6t
Xbit_r108_c214 bl[214] br[214] wl[108] vdd gnd cell_6t
Xbit_r109_c214 bl[214] br[214] wl[109] vdd gnd cell_6t
Xbit_r110_c214 bl[214] br[214] wl[110] vdd gnd cell_6t
Xbit_r111_c214 bl[214] br[214] wl[111] vdd gnd cell_6t
Xbit_r112_c214 bl[214] br[214] wl[112] vdd gnd cell_6t
Xbit_r113_c214 bl[214] br[214] wl[113] vdd gnd cell_6t
Xbit_r114_c214 bl[214] br[214] wl[114] vdd gnd cell_6t
Xbit_r115_c214 bl[214] br[214] wl[115] vdd gnd cell_6t
Xbit_r116_c214 bl[214] br[214] wl[116] vdd gnd cell_6t
Xbit_r117_c214 bl[214] br[214] wl[117] vdd gnd cell_6t
Xbit_r118_c214 bl[214] br[214] wl[118] vdd gnd cell_6t
Xbit_r119_c214 bl[214] br[214] wl[119] vdd gnd cell_6t
Xbit_r120_c214 bl[214] br[214] wl[120] vdd gnd cell_6t
Xbit_r121_c214 bl[214] br[214] wl[121] vdd gnd cell_6t
Xbit_r122_c214 bl[214] br[214] wl[122] vdd gnd cell_6t
Xbit_r123_c214 bl[214] br[214] wl[123] vdd gnd cell_6t
Xbit_r124_c214 bl[214] br[214] wl[124] vdd gnd cell_6t
Xbit_r125_c214 bl[214] br[214] wl[125] vdd gnd cell_6t
Xbit_r126_c214 bl[214] br[214] wl[126] vdd gnd cell_6t
Xbit_r127_c214 bl[214] br[214] wl[127] vdd gnd cell_6t
Xbit_r128_c214 bl[214] br[214] wl[128] vdd gnd cell_6t
Xbit_r129_c214 bl[214] br[214] wl[129] vdd gnd cell_6t
Xbit_r130_c214 bl[214] br[214] wl[130] vdd gnd cell_6t
Xbit_r131_c214 bl[214] br[214] wl[131] vdd gnd cell_6t
Xbit_r132_c214 bl[214] br[214] wl[132] vdd gnd cell_6t
Xbit_r133_c214 bl[214] br[214] wl[133] vdd gnd cell_6t
Xbit_r134_c214 bl[214] br[214] wl[134] vdd gnd cell_6t
Xbit_r135_c214 bl[214] br[214] wl[135] vdd gnd cell_6t
Xbit_r136_c214 bl[214] br[214] wl[136] vdd gnd cell_6t
Xbit_r137_c214 bl[214] br[214] wl[137] vdd gnd cell_6t
Xbit_r138_c214 bl[214] br[214] wl[138] vdd gnd cell_6t
Xbit_r139_c214 bl[214] br[214] wl[139] vdd gnd cell_6t
Xbit_r140_c214 bl[214] br[214] wl[140] vdd gnd cell_6t
Xbit_r141_c214 bl[214] br[214] wl[141] vdd gnd cell_6t
Xbit_r142_c214 bl[214] br[214] wl[142] vdd gnd cell_6t
Xbit_r143_c214 bl[214] br[214] wl[143] vdd gnd cell_6t
Xbit_r144_c214 bl[214] br[214] wl[144] vdd gnd cell_6t
Xbit_r145_c214 bl[214] br[214] wl[145] vdd gnd cell_6t
Xbit_r146_c214 bl[214] br[214] wl[146] vdd gnd cell_6t
Xbit_r147_c214 bl[214] br[214] wl[147] vdd gnd cell_6t
Xbit_r148_c214 bl[214] br[214] wl[148] vdd gnd cell_6t
Xbit_r149_c214 bl[214] br[214] wl[149] vdd gnd cell_6t
Xbit_r150_c214 bl[214] br[214] wl[150] vdd gnd cell_6t
Xbit_r151_c214 bl[214] br[214] wl[151] vdd gnd cell_6t
Xbit_r152_c214 bl[214] br[214] wl[152] vdd gnd cell_6t
Xbit_r153_c214 bl[214] br[214] wl[153] vdd gnd cell_6t
Xbit_r154_c214 bl[214] br[214] wl[154] vdd gnd cell_6t
Xbit_r155_c214 bl[214] br[214] wl[155] vdd gnd cell_6t
Xbit_r156_c214 bl[214] br[214] wl[156] vdd gnd cell_6t
Xbit_r157_c214 bl[214] br[214] wl[157] vdd gnd cell_6t
Xbit_r158_c214 bl[214] br[214] wl[158] vdd gnd cell_6t
Xbit_r159_c214 bl[214] br[214] wl[159] vdd gnd cell_6t
Xbit_r160_c214 bl[214] br[214] wl[160] vdd gnd cell_6t
Xbit_r161_c214 bl[214] br[214] wl[161] vdd gnd cell_6t
Xbit_r162_c214 bl[214] br[214] wl[162] vdd gnd cell_6t
Xbit_r163_c214 bl[214] br[214] wl[163] vdd gnd cell_6t
Xbit_r164_c214 bl[214] br[214] wl[164] vdd gnd cell_6t
Xbit_r165_c214 bl[214] br[214] wl[165] vdd gnd cell_6t
Xbit_r166_c214 bl[214] br[214] wl[166] vdd gnd cell_6t
Xbit_r167_c214 bl[214] br[214] wl[167] vdd gnd cell_6t
Xbit_r168_c214 bl[214] br[214] wl[168] vdd gnd cell_6t
Xbit_r169_c214 bl[214] br[214] wl[169] vdd gnd cell_6t
Xbit_r170_c214 bl[214] br[214] wl[170] vdd gnd cell_6t
Xbit_r171_c214 bl[214] br[214] wl[171] vdd gnd cell_6t
Xbit_r172_c214 bl[214] br[214] wl[172] vdd gnd cell_6t
Xbit_r173_c214 bl[214] br[214] wl[173] vdd gnd cell_6t
Xbit_r174_c214 bl[214] br[214] wl[174] vdd gnd cell_6t
Xbit_r175_c214 bl[214] br[214] wl[175] vdd gnd cell_6t
Xbit_r176_c214 bl[214] br[214] wl[176] vdd gnd cell_6t
Xbit_r177_c214 bl[214] br[214] wl[177] vdd gnd cell_6t
Xbit_r178_c214 bl[214] br[214] wl[178] vdd gnd cell_6t
Xbit_r179_c214 bl[214] br[214] wl[179] vdd gnd cell_6t
Xbit_r180_c214 bl[214] br[214] wl[180] vdd gnd cell_6t
Xbit_r181_c214 bl[214] br[214] wl[181] vdd gnd cell_6t
Xbit_r182_c214 bl[214] br[214] wl[182] vdd gnd cell_6t
Xbit_r183_c214 bl[214] br[214] wl[183] vdd gnd cell_6t
Xbit_r184_c214 bl[214] br[214] wl[184] vdd gnd cell_6t
Xbit_r185_c214 bl[214] br[214] wl[185] vdd gnd cell_6t
Xbit_r186_c214 bl[214] br[214] wl[186] vdd gnd cell_6t
Xbit_r187_c214 bl[214] br[214] wl[187] vdd gnd cell_6t
Xbit_r188_c214 bl[214] br[214] wl[188] vdd gnd cell_6t
Xbit_r189_c214 bl[214] br[214] wl[189] vdd gnd cell_6t
Xbit_r190_c214 bl[214] br[214] wl[190] vdd gnd cell_6t
Xbit_r191_c214 bl[214] br[214] wl[191] vdd gnd cell_6t
Xbit_r192_c214 bl[214] br[214] wl[192] vdd gnd cell_6t
Xbit_r193_c214 bl[214] br[214] wl[193] vdd gnd cell_6t
Xbit_r194_c214 bl[214] br[214] wl[194] vdd gnd cell_6t
Xbit_r195_c214 bl[214] br[214] wl[195] vdd gnd cell_6t
Xbit_r196_c214 bl[214] br[214] wl[196] vdd gnd cell_6t
Xbit_r197_c214 bl[214] br[214] wl[197] vdd gnd cell_6t
Xbit_r198_c214 bl[214] br[214] wl[198] vdd gnd cell_6t
Xbit_r199_c214 bl[214] br[214] wl[199] vdd gnd cell_6t
Xbit_r200_c214 bl[214] br[214] wl[200] vdd gnd cell_6t
Xbit_r201_c214 bl[214] br[214] wl[201] vdd gnd cell_6t
Xbit_r202_c214 bl[214] br[214] wl[202] vdd gnd cell_6t
Xbit_r203_c214 bl[214] br[214] wl[203] vdd gnd cell_6t
Xbit_r204_c214 bl[214] br[214] wl[204] vdd gnd cell_6t
Xbit_r205_c214 bl[214] br[214] wl[205] vdd gnd cell_6t
Xbit_r206_c214 bl[214] br[214] wl[206] vdd gnd cell_6t
Xbit_r207_c214 bl[214] br[214] wl[207] vdd gnd cell_6t
Xbit_r208_c214 bl[214] br[214] wl[208] vdd gnd cell_6t
Xbit_r209_c214 bl[214] br[214] wl[209] vdd gnd cell_6t
Xbit_r210_c214 bl[214] br[214] wl[210] vdd gnd cell_6t
Xbit_r211_c214 bl[214] br[214] wl[211] vdd gnd cell_6t
Xbit_r212_c214 bl[214] br[214] wl[212] vdd gnd cell_6t
Xbit_r213_c214 bl[214] br[214] wl[213] vdd gnd cell_6t
Xbit_r214_c214 bl[214] br[214] wl[214] vdd gnd cell_6t
Xbit_r215_c214 bl[214] br[214] wl[215] vdd gnd cell_6t
Xbit_r216_c214 bl[214] br[214] wl[216] vdd gnd cell_6t
Xbit_r217_c214 bl[214] br[214] wl[217] vdd gnd cell_6t
Xbit_r218_c214 bl[214] br[214] wl[218] vdd gnd cell_6t
Xbit_r219_c214 bl[214] br[214] wl[219] vdd gnd cell_6t
Xbit_r220_c214 bl[214] br[214] wl[220] vdd gnd cell_6t
Xbit_r221_c214 bl[214] br[214] wl[221] vdd gnd cell_6t
Xbit_r222_c214 bl[214] br[214] wl[222] vdd gnd cell_6t
Xbit_r223_c214 bl[214] br[214] wl[223] vdd gnd cell_6t
Xbit_r224_c214 bl[214] br[214] wl[224] vdd gnd cell_6t
Xbit_r225_c214 bl[214] br[214] wl[225] vdd gnd cell_6t
Xbit_r226_c214 bl[214] br[214] wl[226] vdd gnd cell_6t
Xbit_r227_c214 bl[214] br[214] wl[227] vdd gnd cell_6t
Xbit_r228_c214 bl[214] br[214] wl[228] vdd gnd cell_6t
Xbit_r229_c214 bl[214] br[214] wl[229] vdd gnd cell_6t
Xbit_r230_c214 bl[214] br[214] wl[230] vdd gnd cell_6t
Xbit_r231_c214 bl[214] br[214] wl[231] vdd gnd cell_6t
Xbit_r232_c214 bl[214] br[214] wl[232] vdd gnd cell_6t
Xbit_r233_c214 bl[214] br[214] wl[233] vdd gnd cell_6t
Xbit_r234_c214 bl[214] br[214] wl[234] vdd gnd cell_6t
Xbit_r235_c214 bl[214] br[214] wl[235] vdd gnd cell_6t
Xbit_r236_c214 bl[214] br[214] wl[236] vdd gnd cell_6t
Xbit_r237_c214 bl[214] br[214] wl[237] vdd gnd cell_6t
Xbit_r238_c214 bl[214] br[214] wl[238] vdd gnd cell_6t
Xbit_r239_c214 bl[214] br[214] wl[239] vdd gnd cell_6t
Xbit_r240_c214 bl[214] br[214] wl[240] vdd gnd cell_6t
Xbit_r241_c214 bl[214] br[214] wl[241] vdd gnd cell_6t
Xbit_r242_c214 bl[214] br[214] wl[242] vdd gnd cell_6t
Xbit_r243_c214 bl[214] br[214] wl[243] vdd gnd cell_6t
Xbit_r244_c214 bl[214] br[214] wl[244] vdd gnd cell_6t
Xbit_r245_c214 bl[214] br[214] wl[245] vdd gnd cell_6t
Xbit_r246_c214 bl[214] br[214] wl[246] vdd gnd cell_6t
Xbit_r247_c214 bl[214] br[214] wl[247] vdd gnd cell_6t
Xbit_r248_c214 bl[214] br[214] wl[248] vdd gnd cell_6t
Xbit_r249_c214 bl[214] br[214] wl[249] vdd gnd cell_6t
Xbit_r250_c214 bl[214] br[214] wl[250] vdd gnd cell_6t
Xbit_r251_c214 bl[214] br[214] wl[251] vdd gnd cell_6t
Xbit_r252_c214 bl[214] br[214] wl[252] vdd gnd cell_6t
Xbit_r253_c214 bl[214] br[214] wl[253] vdd gnd cell_6t
Xbit_r254_c214 bl[214] br[214] wl[254] vdd gnd cell_6t
Xbit_r255_c214 bl[214] br[214] wl[255] vdd gnd cell_6t
Xbit_r0_c215 bl[215] br[215] wl[0] vdd gnd cell_6t
Xbit_r1_c215 bl[215] br[215] wl[1] vdd gnd cell_6t
Xbit_r2_c215 bl[215] br[215] wl[2] vdd gnd cell_6t
Xbit_r3_c215 bl[215] br[215] wl[3] vdd gnd cell_6t
Xbit_r4_c215 bl[215] br[215] wl[4] vdd gnd cell_6t
Xbit_r5_c215 bl[215] br[215] wl[5] vdd gnd cell_6t
Xbit_r6_c215 bl[215] br[215] wl[6] vdd gnd cell_6t
Xbit_r7_c215 bl[215] br[215] wl[7] vdd gnd cell_6t
Xbit_r8_c215 bl[215] br[215] wl[8] vdd gnd cell_6t
Xbit_r9_c215 bl[215] br[215] wl[9] vdd gnd cell_6t
Xbit_r10_c215 bl[215] br[215] wl[10] vdd gnd cell_6t
Xbit_r11_c215 bl[215] br[215] wl[11] vdd gnd cell_6t
Xbit_r12_c215 bl[215] br[215] wl[12] vdd gnd cell_6t
Xbit_r13_c215 bl[215] br[215] wl[13] vdd gnd cell_6t
Xbit_r14_c215 bl[215] br[215] wl[14] vdd gnd cell_6t
Xbit_r15_c215 bl[215] br[215] wl[15] vdd gnd cell_6t
Xbit_r16_c215 bl[215] br[215] wl[16] vdd gnd cell_6t
Xbit_r17_c215 bl[215] br[215] wl[17] vdd gnd cell_6t
Xbit_r18_c215 bl[215] br[215] wl[18] vdd gnd cell_6t
Xbit_r19_c215 bl[215] br[215] wl[19] vdd gnd cell_6t
Xbit_r20_c215 bl[215] br[215] wl[20] vdd gnd cell_6t
Xbit_r21_c215 bl[215] br[215] wl[21] vdd gnd cell_6t
Xbit_r22_c215 bl[215] br[215] wl[22] vdd gnd cell_6t
Xbit_r23_c215 bl[215] br[215] wl[23] vdd gnd cell_6t
Xbit_r24_c215 bl[215] br[215] wl[24] vdd gnd cell_6t
Xbit_r25_c215 bl[215] br[215] wl[25] vdd gnd cell_6t
Xbit_r26_c215 bl[215] br[215] wl[26] vdd gnd cell_6t
Xbit_r27_c215 bl[215] br[215] wl[27] vdd gnd cell_6t
Xbit_r28_c215 bl[215] br[215] wl[28] vdd gnd cell_6t
Xbit_r29_c215 bl[215] br[215] wl[29] vdd gnd cell_6t
Xbit_r30_c215 bl[215] br[215] wl[30] vdd gnd cell_6t
Xbit_r31_c215 bl[215] br[215] wl[31] vdd gnd cell_6t
Xbit_r32_c215 bl[215] br[215] wl[32] vdd gnd cell_6t
Xbit_r33_c215 bl[215] br[215] wl[33] vdd gnd cell_6t
Xbit_r34_c215 bl[215] br[215] wl[34] vdd gnd cell_6t
Xbit_r35_c215 bl[215] br[215] wl[35] vdd gnd cell_6t
Xbit_r36_c215 bl[215] br[215] wl[36] vdd gnd cell_6t
Xbit_r37_c215 bl[215] br[215] wl[37] vdd gnd cell_6t
Xbit_r38_c215 bl[215] br[215] wl[38] vdd gnd cell_6t
Xbit_r39_c215 bl[215] br[215] wl[39] vdd gnd cell_6t
Xbit_r40_c215 bl[215] br[215] wl[40] vdd gnd cell_6t
Xbit_r41_c215 bl[215] br[215] wl[41] vdd gnd cell_6t
Xbit_r42_c215 bl[215] br[215] wl[42] vdd gnd cell_6t
Xbit_r43_c215 bl[215] br[215] wl[43] vdd gnd cell_6t
Xbit_r44_c215 bl[215] br[215] wl[44] vdd gnd cell_6t
Xbit_r45_c215 bl[215] br[215] wl[45] vdd gnd cell_6t
Xbit_r46_c215 bl[215] br[215] wl[46] vdd gnd cell_6t
Xbit_r47_c215 bl[215] br[215] wl[47] vdd gnd cell_6t
Xbit_r48_c215 bl[215] br[215] wl[48] vdd gnd cell_6t
Xbit_r49_c215 bl[215] br[215] wl[49] vdd gnd cell_6t
Xbit_r50_c215 bl[215] br[215] wl[50] vdd gnd cell_6t
Xbit_r51_c215 bl[215] br[215] wl[51] vdd gnd cell_6t
Xbit_r52_c215 bl[215] br[215] wl[52] vdd gnd cell_6t
Xbit_r53_c215 bl[215] br[215] wl[53] vdd gnd cell_6t
Xbit_r54_c215 bl[215] br[215] wl[54] vdd gnd cell_6t
Xbit_r55_c215 bl[215] br[215] wl[55] vdd gnd cell_6t
Xbit_r56_c215 bl[215] br[215] wl[56] vdd gnd cell_6t
Xbit_r57_c215 bl[215] br[215] wl[57] vdd gnd cell_6t
Xbit_r58_c215 bl[215] br[215] wl[58] vdd gnd cell_6t
Xbit_r59_c215 bl[215] br[215] wl[59] vdd gnd cell_6t
Xbit_r60_c215 bl[215] br[215] wl[60] vdd gnd cell_6t
Xbit_r61_c215 bl[215] br[215] wl[61] vdd gnd cell_6t
Xbit_r62_c215 bl[215] br[215] wl[62] vdd gnd cell_6t
Xbit_r63_c215 bl[215] br[215] wl[63] vdd gnd cell_6t
Xbit_r64_c215 bl[215] br[215] wl[64] vdd gnd cell_6t
Xbit_r65_c215 bl[215] br[215] wl[65] vdd gnd cell_6t
Xbit_r66_c215 bl[215] br[215] wl[66] vdd gnd cell_6t
Xbit_r67_c215 bl[215] br[215] wl[67] vdd gnd cell_6t
Xbit_r68_c215 bl[215] br[215] wl[68] vdd gnd cell_6t
Xbit_r69_c215 bl[215] br[215] wl[69] vdd gnd cell_6t
Xbit_r70_c215 bl[215] br[215] wl[70] vdd gnd cell_6t
Xbit_r71_c215 bl[215] br[215] wl[71] vdd gnd cell_6t
Xbit_r72_c215 bl[215] br[215] wl[72] vdd gnd cell_6t
Xbit_r73_c215 bl[215] br[215] wl[73] vdd gnd cell_6t
Xbit_r74_c215 bl[215] br[215] wl[74] vdd gnd cell_6t
Xbit_r75_c215 bl[215] br[215] wl[75] vdd gnd cell_6t
Xbit_r76_c215 bl[215] br[215] wl[76] vdd gnd cell_6t
Xbit_r77_c215 bl[215] br[215] wl[77] vdd gnd cell_6t
Xbit_r78_c215 bl[215] br[215] wl[78] vdd gnd cell_6t
Xbit_r79_c215 bl[215] br[215] wl[79] vdd gnd cell_6t
Xbit_r80_c215 bl[215] br[215] wl[80] vdd gnd cell_6t
Xbit_r81_c215 bl[215] br[215] wl[81] vdd gnd cell_6t
Xbit_r82_c215 bl[215] br[215] wl[82] vdd gnd cell_6t
Xbit_r83_c215 bl[215] br[215] wl[83] vdd gnd cell_6t
Xbit_r84_c215 bl[215] br[215] wl[84] vdd gnd cell_6t
Xbit_r85_c215 bl[215] br[215] wl[85] vdd gnd cell_6t
Xbit_r86_c215 bl[215] br[215] wl[86] vdd gnd cell_6t
Xbit_r87_c215 bl[215] br[215] wl[87] vdd gnd cell_6t
Xbit_r88_c215 bl[215] br[215] wl[88] vdd gnd cell_6t
Xbit_r89_c215 bl[215] br[215] wl[89] vdd gnd cell_6t
Xbit_r90_c215 bl[215] br[215] wl[90] vdd gnd cell_6t
Xbit_r91_c215 bl[215] br[215] wl[91] vdd gnd cell_6t
Xbit_r92_c215 bl[215] br[215] wl[92] vdd gnd cell_6t
Xbit_r93_c215 bl[215] br[215] wl[93] vdd gnd cell_6t
Xbit_r94_c215 bl[215] br[215] wl[94] vdd gnd cell_6t
Xbit_r95_c215 bl[215] br[215] wl[95] vdd gnd cell_6t
Xbit_r96_c215 bl[215] br[215] wl[96] vdd gnd cell_6t
Xbit_r97_c215 bl[215] br[215] wl[97] vdd gnd cell_6t
Xbit_r98_c215 bl[215] br[215] wl[98] vdd gnd cell_6t
Xbit_r99_c215 bl[215] br[215] wl[99] vdd gnd cell_6t
Xbit_r100_c215 bl[215] br[215] wl[100] vdd gnd cell_6t
Xbit_r101_c215 bl[215] br[215] wl[101] vdd gnd cell_6t
Xbit_r102_c215 bl[215] br[215] wl[102] vdd gnd cell_6t
Xbit_r103_c215 bl[215] br[215] wl[103] vdd gnd cell_6t
Xbit_r104_c215 bl[215] br[215] wl[104] vdd gnd cell_6t
Xbit_r105_c215 bl[215] br[215] wl[105] vdd gnd cell_6t
Xbit_r106_c215 bl[215] br[215] wl[106] vdd gnd cell_6t
Xbit_r107_c215 bl[215] br[215] wl[107] vdd gnd cell_6t
Xbit_r108_c215 bl[215] br[215] wl[108] vdd gnd cell_6t
Xbit_r109_c215 bl[215] br[215] wl[109] vdd gnd cell_6t
Xbit_r110_c215 bl[215] br[215] wl[110] vdd gnd cell_6t
Xbit_r111_c215 bl[215] br[215] wl[111] vdd gnd cell_6t
Xbit_r112_c215 bl[215] br[215] wl[112] vdd gnd cell_6t
Xbit_r113_c215 bl[215] br[215] wl[113] vdd gnd cell_6t
Xbit_r114_c215 bl[215] br[215] wl[114] vdd gnd cell_6t
Xbit_r115_c215 bl[215] br[215] wl[115] vdd gnd cell_6t
Xbit_r116_c215 bl[215] br[215] wl[116] vdd gnd cell_6t
Xbit_r117_c215 bl[215] br[215] wl[117] vdd gnd cell_6t
Xbit_r118_c215 bl[215] br[215] wl[118] vdd gnd cell_6t
Xbit_r119_c215 bl[215] br[215] wl[119] vdd gnd cell_6t
Xbit_r120_c215 bl[215] br[215] wl[120] vdd gnd cell_6t
Xbit_r121_c215 bl[215] br[215] wl[121] vdd gnd cell_6t
Xbit_r122_c215 bl[215] br[215] wl[122] vdd gnd cell_6t
Xbit_r123_c215 bl[215] br[215] wl[123] vdd gnd cell_6t
Xbit_r124_c215 bl[215] br[215] wl[124] vdd gnd cell_6t
Xbit_r125_c215 bl[215] br[215] wl[125] vdd gnd cell_6t
Xbit_r126_c215 bl[215] br[215] wl[126] vdd gnd cell_6t
Xbit_r127_c215 bl[215] br[215] wl[127] vdd gnd cell_6t
Xbit_r128_c215 bl[215] br[215] wl[128] vdd gnd cell_6t
Xbit_r129_c215 bl[215] br[215] wl[129] vdd gnd cell_6t
Xbit_r130_c215 bl[215] br[215] wl[130] vdd gnd cell_6t
Xbit_r131_c215 bl[215] br[215] wl[131] vdd gnd cell_6t
Xbit_r132_c215 bl[215] br[215] wl[132] vdd gnd cell_6t
Xbit_r133_c215 bl[215] br[215] wl[133] vdd gnd cell_6t
Xbit_r134_c215 bl[215] br[215] wl[134] vdd gnd cell_6t
Xbit_r135_c215 bl[215] br[215] wl[135] vdd gnd cell_6t
Xbit_r136_c215 bl[215] br[215] wl[136] vdd gnd cell_6t
Xbit_r137_c215 bl[215] br[215] wl[137] vdd gnd cell_6t
Xbit_r138_c215 bl[215] br[215] wl[138] vdd gnd cell_6t
Xbit_r139_c215 bl[215] br[215] wl[139] vdd gnd cell_6t
Xbit_r140_c215 bl[215] br[215] wl[140] vdd gnd cell_6t
Xbit_r141_c215 bl[215] br[215] wl[141] vdd gnd cell_6t
Xbit_r142_c215 bl[215] br[215] wl[142] vdd gnd cell_6t
Xbit_r143_c215 bl[215] br[215] wl[143] vdd gnd cell_6t
Xbit_r144_c215 bl[215] br[215] wl[144] vdd gnd cell_6t
Xbit_r145_c215 bl[215] br[215] wl[145] vdd gnd cell_6t
Xbit_r146_c215 bl[215] br[215] wl[146] vdd gnd cell_6t
Xbit_r147_c215 bl[215] br[215] wl[147] vdd gnd cell_6t
Xbit_r148_c215 bl[215] br[215] wl[148] vdd gnd cell_6t
Xbit_r149_c215 bl[215] br[215] wl[149] vdd gnd cell_6t
Xbit_r150_c215 bl[215] br[215] wl[150] vdd gnd cell_6t
Xbit_r151_c215 bl[215] br[215] wl[151] vdd gnd cell_6t
Xbit_r152_c215 bl[215] br[215] wl[152] vdd gnd cell_6t
Xbit_r153_c215 bl[215] br[215] wl[153] vdd gnd cell_6t
Xbit_r154_c215 bl[215] br[215] wl[154] vdd gnd cell_6t
Xbit_r155_c215 bl[215] br[215] wl[155] vdd gnd cell_6t
Xbit_r156_c215 bl[215] br[215] wl[156] vdd gnd cell_6t
Xbit_r157_c215 bl[215] br[215] wl[157] vdd gnd cell_6t
Xbit_r158_c215 bl[215] br[215] wl[158] vdd gnd cell_6t
Xbit_r159_c215 bl[215] br[215] wl[159] vdd gnd cell_6t
Xbit_r160_c215 bl[215] br[215] wl[160] vdd gnd cell_6t
Xbit_r161_c215 bl[215] br[215] wl[161] vdd gnd cell_6t
Xbit_r162_c215 bl[215] br[215] wl[162] vdd gnd cell_6t
Xbit_r163_c215 bl[215] br[215] wl[163] vdd gnd cell_6t
Xbit_r164_c215 bl[215] br[215] wl[164] vdd gnd cell_6t
Xbit_r165_c215 bl[215] br[215] wl[165] vdd gnd cell_6t
Xbit_r166_c215 bl[215] br[215] wl[166] vdd gnd cell_6t
Xbit_r167_c215 bl[215] br[215] wl[167] vdd gnd cell_6t
Xbit_r168_c215 bl[215] br[215] wl[168] vdd gnd cell_6t
Xbit_r169_c215 bl[215] br[215] wl[169] vdd gnd cell_6t
Xbit_r170_c215 bl[215] br[215] wl[170] vdd gnd cell_6t
Xbit_r171_c215 bl[215] br[215] wl[171] vdd gnd cell_6t
Xbit_r172_c215 bl[215] br[215] wl[172] vdd gnd cell_6t
Xbit_r173_c215 bl[215] br[215] wl[173] vdd gnd cell_6t
Xbit_r174_c215 bl[215] br[215] wl[174] vdd gnd cell_6t
Xbit_r175_c215 bl[215] br[215] wl[175] vdd gnd cell_6t
Xbit_r176_c215 bl[215] br[215] wl[176] vdd gnd cell_6t
Xbit_r177_c215 bl[215] br[215] wl[177] vdd gnd cell_6t
Xbit_r178_c215 bl[215] br[215] wl[178] vdd gnd cell_6t
Xbit_r179_c215 bl[215] br[215] wl[179] vdd gnd cell_6t
Xbit_r180_c215 bl[215] br[215] wl[180] vdd gnd cell_6t
Xbit_r181_c215 bl[215] br[215] wl[181] vdd gnd cell_6t
Xbit_r182_c215 bl[215] br[215] wl[182] vdd gnd cell_6t
Xbit_r183_c215 bl[215] br[215] wl[183] vdd gnd cell_6t
Xbit_r184_c215 bl[215] br[215] wl[184] vdd gnd cell_6t
Xbit_r185_c215 bl[215] br[215] wl[185] vdd gnd cell_6t
Xbit_r186_c215 bl[215] br[215] wl[186] vdd gnd cell_6t
Xbit_r187_c215 bl[215] br[215] wl[187] vdd gnd cell_6t
Xbit_r188_c215 bl[215] br[215] wl[188] vdd gnd cell_6t
Xbit_r189_c215 bl[215] br[215] wl[189] vdd gnd cell_6t
Xbit_r190_c215 bl[215] br[215] wl[190] vdd gnd cell_6t
Xbit_r191_c215 bl[215] br[215] wl[191] vdd gnd cell_6t
Xbit_r192_c215 bl[215] br[215] wl[192] vdd gnd cell_6t
Xbit_r193_c215 bl[215] br[215] wl[193] vdd gnd cell_6t
Xbit_r194_c215 bl[215] br[215] wl[194] vdd gnd cell_6t
Xbit_r195_c215 bl[215] br[215] wl[195] vdd gnd cell_6t
Xbit_r196_c215 bl[215] br[215] wl[196] vdd gnd cell_6t
Xbit_r197_c215 bl[215] br[215] wl[197] vdd gnd cell_6t
Xbit_r198_c215 bl[215] br[215] wl[198] vdd gnd cell_6t
Xbit_r199_c215 bl[215] br[215] wl[199] vdd gnd cell_6t
Xbit_r200_c215 bl[215] br[215] wl[200] vdd gnd cell_6t
Xbit_r201_c215 bl[215] br[215] wl[201] vdd gnd cell_6t
Xbit_r202_c215 bl[215] br[215] wl[202] vdd gnd cell_6t
Xbit_r203_c215 bl[215] br[215] wl[203] vdd gnd cell_6t
Xbit_r204_c215 bl[215] br[215] wl[204] vdd gnd cell_6t
Xbit_r205_c215 bl[215] br[215] wl[205] vdd gnd cell_6t
Xbit_r206_c215 bl[215] br[215] wl[206] vdd gnd cell_6t
Xbit_r207_c215 bl[215] br[215] wl[207] vdd gnd cell_6t
Xbit_r208_c215 bl[215] br[215] wl[208] vdd gnd cell_6t
Xbit_r209_c215 bl[215] br[215] wl[209] vdd gnd cell_6t
Xbit_r210_c215 bl[215] br[215] wl[210] vdd gnd cell_6t
Xbit_r211_c215 bl[215] br[215] wl[211] vdd gnd cell_6t
Xbit_r212_c215 bl[215] br[215] wl[212] vdd gnd cell_6t
Xbit_r213_c215 bl[215] br[215] wl[213] vdd gnd cell_6t
Xbit_r214_c215 bl[215] br[215] wl[214] vdd gnd cell_6t
Xbit_r215_c215 bl[215] br[215] wl[215] vdd gnd cell_6t
Xbit_r216_c215 bl[215] br[215] wl[216] vdd gnd cell_6t
Xbit_r217_c215 bl[215] br[215] wl[217] vdd gnd cell_6t
Xbit_r218_c215 bl[215] br[215] wl[218] vdd gnd cell_6t
Xbit_r219_c215 bl[215] br[215] wl[219] vdd gnd cell_6t
Xbit_r220_c215 bl[215] br[215] wl[220] vdd gnd cell_6t
Xbit_r221_c215 bl[215] br[215] wl[221] vdd gnd cell_6t
Xbit_r222_c215 bl[215] br[215] wl[222] vdd gnd cell_6t
Xbit_r223_c215 bl[215] br[215] wl[223] vdd gnd cell_6t
Xbit_r224_c215 bl[215] br[215] wl[224] vdd gnd cell_6t
Xbit_r225_c215 bl[215] br[215] wl[225] vdd gnd cell_6t
Xbit_r226_c215 bl[215] br[215] wl[226] vdd gnd cell_6t
Xbit_r227_c215 bl[215] br[215] wl[227] vdd gnd cell_6t
Xbit_r228_c215 bl[215] br[215] wl[228] vdd gnd cell_6t
Xbit_r229_c215 bl[215] br[215] wl[229] vdd gnd cell_6t
Xbit_r230_c215 bl[215] br[215] wl[230] vdd gnd cell_6t
Xbit_r231_c215 bl[215] br[215] wl[231] vdd gnd cell_6t
Xbit_r232_c215 bl[215] br[215] wl[232] vdd gnd cell_6t
Xbit_r233_c215 bl[215] br[215] wl[233] vdd gnd cell_6t
Xbit_r234_c215 bl[215] br[215] wl[234] vdd gnd cell_6t
Xbit_r235_c215 bl[215] br[215] wl[235] vdd gnd cell_6t
Xbit_r236_c215 bl[215] br[215] wl[236] vdd gnd cell_6t
Xbit_r237_c215 bl[215] br[215] wl[237] vdd gnd cell_6t
Xbit_r238_c215 bl[215] br[215] wl[238] vdd gnd cell_6t
Xbit_r239_c215 bl[215] br[215] wl[239] vdd gnd cell_6t
Xbit_r240_c215 bl[215] br[215] wl[240] vdd gnd cell_6t
Xbit_r241_c215 bl[215] br[215] wl[241] vdd gnd cell_6t
Xbit_r242_c215 bl[215] br[215] wl[242] vdd gnd cell_6t
Xbit_r243_c215 bl[215] br[215] wl[243] vdd gnd cell_6t
Xbit_r244_c215 bl[215] br[215] wl[244] vdd gnd cell_6t
Xbit_r245_c215 bl[215] br[215] wl[245] vdd gnd cell_6t
Xbit_r246_c215 bl[215] br[215] wl[246] vdd gnd cell_6t
Xbit_r247_c215 bl[215] br[215] wl[247] vdd gnd cell_6t
Xbit_r248_c215 bl[215] br[215] wl[248] vdd gnd cell_6t
Xbit_r249_c215 bl[215] br[215] wl[249] vdd gnd cell_6t
Xbit_r250_c215 bl[215] br[215] wl[250] vdd gnd cell_6t
Xbit_r251_c215 bl[215] br[215] wl[251] vdd gnd cell_6t
Xbit_r252_c215 bl[215] br[215] wl[252] vdd gnd cell_6t
Xbit_r253_c215 bl[215] br[215] wl[253] vdd gnd cell_6t
Xbit_r254_c215 bl[215] br[215] wl[254] vdd gnd cell_6t
Xbit_r255_c215 bl[215] br[215] wl[255] vdd gnd cell_6t
Xbit_r0_c216 bl[216] br[216] wl[0] vdd gnd cell_6t
Xbit_r1_c216 bl[216] br[216] wl[1] vdd gnd cell_6t
Xbit_r2_c216 bl[216] br[216] wl[2] vdd gnd cell_6t
Xbit_r3_c216 bl[216] br[216] wl[3] vdd gnd cell_6t
Xbit_r4_c216 bl[216] br[216] wl[4] vdd gnd cell_6t
Xbit_r5_c216 bl[216] br[216] wl[5] vdd gnd cell_6t
Xbit_r6_c216 bl[216] br[216] wl[6] vdd gnd cell_6t
Xbit_r7_c216 bl[216] br[216] wl[7] vdd gnd cell_6t
Xbit_r8_c216 bl[216] br[216] wl[8] vdd gnd cell_6t
Xbit_r9_c216 bl[216] br[216] wl[9] vdd gnd cell_6t
Xbit_r10_c216 bl[216] br[216] wl[10] vdd gnd cell_6t
Xbit_r11_c216 bl[216] br[216] wl[11] vdd gnd cell_6t
Xbit_r12_c216 bl[216] br[216] wl[12] vdd gnd cell_6t
Xbit_r13_c216 bl[216] br[216] wl[13] vdd gnd cell_6t
Xbit_r14_c216 bl[216] br[216] wl[14] vdd gnd cell_6t
Xbit_r15_c216 bl[216] br[216] wl[15] vdd gnd cell_6t
Xbit_r16_c216 bl[216] br[216] wl[16] vdd gnd cell_6t
Xbit_r17_c216 bl[216] br[216] wl[17] vdd gnd cell_6t
Xbit_r18_c216 bl[216] br[216] wl[18] vdd gnd cell_6t
Xbit_r19_c216 bl[216] br[216] wl[19] vdd gnd cell_6t
Xbit_r20_c216 bl[216] br[216] wl[20] vdd gnd cell_6t
Xbit_r21_c216 bl[216] br[216] wl[21] vdd gnd cell_6t
Xbit_r22_c216 bl[216] br[216] wl[22] vdd gnd cell_6t
Xbit_r23_c216 bl[216] br[216] wl[23] vdd gnd cell_6t
Xbit_r24_c216 bl[216] br[216] wl[24] vdd gnd cell_6t
Xbit_r25_c216 bl[216] br[216] wl[25] vdd gnd cell_6t
Xbit_r26_c216 bl[216] br[216] wl[26] vdd gnd cell_6t
Xbit_r27_c216 bl[216] br[216] wl[27] vdd gnd cell_6t
Xbit_r28_c216 bl[216] br[216] wl[28] vdd gnd cell_6t
Xbit_r29_c216 bl[216] br[216] wl[29] vdd gnd cell_6t
Xbit_r30_c216 bl[216] br[216] wl[30] vdd gnd cell_6t
Xbit_r31_c216 bl[216] br[216] wl[31] vdd gnd cell_6t
Xbit_r32_c216 bl[216] br[216] wl[32] vdd gnd cell_6t
Xbit_r33_c216 bl[216] br[216] wl[33] vdd gnd cell_6t
Xbit_r34_c216 bl[216] br[216] wl[34] vdd gnd cell_6t
Xbit_r35_c216 bl[216] br[216] wl[35] vdd gnd cell_6t
Xbit_r36_c216 bl[216] br[216] wl[36] vdd gnd cell_6t
Xbit_r37_c216 bl[216] br[216] wl[37] vdd gnd cell_6t
Xbit_r38_c216 bl[216] br[216] wl[38] vdd gnd cell_6t
Xbit_r39_c216 bl[216] br[216] wl[39] vdd gnd cell_6t
Xbit_r40_c216 bl[216] br[216] wl[40] vdd gnd cell_6t
Xbit_r41_c216 bl[216] br[216] wl[41] vdd gnd cell_6t
Xbit_r42_c216 bl[216] br[216] wl[42] vdd gnd cell_6t
Xbit_r43_c216 bl[216] br[216] wl[43] vdd gnd cell_6t
Xbit_r44_c216 bl[216] br[216] wl[44] vdd gnd cell_6t
Xbit_r45_c216 bl[216] br[216] wl[45] vdd gnd cell_6t
Xbit_r46_c216 bl[216] br[216] wl[46] vdd gnd cell_6t
Xbit_r47_c216 bl[216] br[216] wl[47] vdd gnd cell_6t
Xbit_r48_c216 bl[216] br[216] wl[48] vdd gnd cell_6t
Xbit_r49_c216 bl[216] br[216] wl[49] vdd gnd cell_6t
Xbit_r50_c216 bl[216] br[216] wl[50] vdd gnd cell_6t
Xbit_r51_c216 bl[216] br[216] wl[51] vdd gnd cell_6t
Xbit_r52_c216 bl[216] br[216] wl[52] vdd gnd cell_6t
Xbit_r53_c216 bl[216] br[216] wl[53] vdd gnd cell_6t
Xbit_r54_c216 bl[216] br[216] wl[54] vdd gnd cell_6t
Xbit_r55_c216 bl[216] br[216] wl[55] vdd gnd cell_6t
Xbit_r56_c216 bl[216] br[216] wl[56] vdd gnd cell_6t
Xbit_r57_c216 bl[216] br[216] wl[57] vdd gnd cell_6t
Xbit_r58_c216 bl[216] br[216] wl[58] vdd gnd cell_6t
Xbit_r59_c216 bl[216] br[216] wl[59] vdd gnd cell_6t
Xbit_r60_c216 bl[216] br[216] wl[60] vdd gnd cell_6t
Xbit_r61_c216 bl[216] br[216] wl[61] vdd gnd cell_6t
Xbit_r62_c216 bl[216] br[216] wl[62] vdd gnd cell_6t
Xbit_r63_c216 bl[216] br[216] wl[63] vdd gnd cell_6t
Xbit_r64_c216 bl[216] br[216] wl[64] vdd gnd cell_6t
Xbit_r65_c216 bl[216] br[216] wl[65] vdd gnd cell_6t
Xbit_r66_c216 bl[216] br[216] wl[66] vdd gnd cell_6t
Xbit_r67_c216 bl[216] br[216] wl[67] vdd gnd cell_6t
Xbit_r68_c216 bl[216] br[216] wl[68] vdd gnd cell_6t
Xbit_r69_c216 bl[216] br[216] wl[69] vdd gnd cell_6t
Xbit_r70_c216 bl[216] br[216] wl[70] vdd gnd cell_6t
Xbit_r71_c216 bl[216] br[216] wl[71] vdd gnd cell_6t
Xbit_r72_c216 bl[216] br[216] wl[72] vdd gnd cell_6t
Xbit_r73_c216 bl[216] br[216] wl[73] vdd gnd cell_6t
Xbit_r74_c216 bl[216] br[216] wl[74] vdd gnd cell_6t
Xbit_r75_c216 bl[216] br[216] wl[75] vdd gnd cell_6t
Xbit_r76_c216 bl[216] br[216] wl[76] vdd gnd cell_6t
Xbit_r77_c216 bl[216] br[216] wl[77] vdd gnd cell_6t
Xbit_r78_c216 bl[216] br[216] wl[78] vdd gnd cell_6t
Xbit_r79_c216 bl[216] br[216] wl[79] vdd gnd cell_6t
Xbit_r80_c216 bl[216] br[216] wl[80] vdd gnd cell_6t
Xbit_r81_c216 bl[216] br[216] wl[81] vdd gnd cell_6t
Xbit_r82_c216 bl[216] br[216] wl[82] vdd gnd cell_6t
Xbit_r83_c216 bl[216] br[216] wl[83] vdd gnd cell_6t
Xbit_r84_c216 bl[216] br[216] wl[84] vdd gnd cell_6t
Xbit_r85_c216 bl[216] br[216] wl[85] vdd gnd cell_6t
Xbit_r86_c216 bl[216] br[216] wl[86] vdd gnd cell_6t
Xbit_r87_c216 bl[216] br[216] wl[87] vdd gnd cell_6t
Xbit_r88_c216 bl[216] br[216] wl[88] vdd gnd cell_6t
Xbit_r89_c216 bl[216] br[216] wl[89] vdd gnd cell_6t
Xbit_r90_c216 bl[216] br[216] wl[90] vdd gnd cell_6t
Xbit_r91_c216 bl[216] br[216] wl[91] vdd gnd cell_6t
Xbit_r92_c216 bl[216] br[216] wl[92] vdd gnd cell_6t
Xbit_r93_c216 bl[216] br[216] wl[93] vdd gnd cell_6t
Xbit_r94_c216 bl[216] br[216] wl[94] vdd gnd cell_6t
Xbit_r95_c216 bl[216] br[216] wl[95] vdd gnd cell_6t
Xbit_r96_c216 bl[216] br[216] wl[96] vdd gnd cell_6t
Xbit_r97_c216 bl[216] br[216] wl[97] vdd gnd cell_6t
Xbit_r98_c216 bl[216] br[216] wl[98] vdd gnd cell_6t
Xbit_r99_c216 bl[216] br[216] wl[99] vdd gnd cell_6t
Xbit_r100_c216 bl[216] br[216] wl[100] vdd gnd cell_6t
Xbit_r101_c216 bl[216] br[216] wl[101] vdd gnd cell_6t
Xbit_r102_c216 bl[216] br[216] wl[102] vdd gnd cell_6t
Xbit_r103_c216 bl[216] br[216] wl[103] vdd gnd cell_6t
Xbit_r104_c216 bl[216] br[216] wl[104] vdd gnd cell_6t
Xbit_r105_c216 bl[216] br[216] wl[105] vdd gnd cell_6t
Xbit_r106_c216 bl[216] br[216] wl[106] vdd gnd cell_6t
Xbit_r107_c216 bl[216] br[216] wl[107] vdd gnd cell_6t
Xbit_r108_c216 bl[216] br[216] wl[108] vdd gnd cell_6t
Xbit_r109_c216 bl[216] br[216] wl[109] vdd gnd cell_6t
Xbit_r110_c216 bl[216] br[216] wl[110] vdd gnd cell_6t
Xbit_r111_c216 bl[216] br[216] wl[111] vdd gnd cell_6t
Xbit_r112_c216 bl[216] br[216] wl[112] vdd gnd cell_6t
Xbit_r113_c216 bl[216] br[216] wl[113] vdd gnd cell_6t
Xbit_r114_c216 bl[216] br[216] wl[114] vdd gnd cell_6t
Xbit_r115_c216 bl[216] br[216] wl[115] vdd gnd cell_6t
Xbit_r116_c216 bl[216] br[216] wl[116] vdd gnd cell_6t
Xbit_r117_c216 bl[216] br[216] wl[117] vdd gnd cell_6t
Xbit_r118_c216 bl[216] br[216] wl[118] vdd gnd cell_6t
Xbit_r119_c216 bl[216] br[216] wl[119] vdd gnd cell_6t
Xbit_r120_c216 bl[216] br[216] wl[120] vdd gnd cell_6t
Xbit_r121_c216 bl[216] br[216] wl[121] vdd gnd cell_6t
Xbit_r122_c216 bl[216] br[216] wl[122] vdd gnd cell_6t
Xbit_r123_c216 bl[216] br[216] wl[123] vdd gnd cell_6t
Xbit_r124_c216 bl[216] br[216] wl[124] vdd gnd cell_6t
Xbit_r125_c216 bl[216] br[216] wl[125] vdd gnd cell_6t
Xbit_r126_c216 bl[216] br[216] wl[126] vdd gnd cell_6t
Xbit_r127_c216 bl[216] br[216] wl[127] vdd gnd cell_6t
Xbit_r128_c216 bl[216] br[216] wl[128] vdd gnd cell_6t
Xbit_r129_c216 bl[216] br[216] wl[129] vdd gnd cell_6t
Xbit_r130_c216 bl[216] br[216] wl[130] vdd gnd cell_6t
Xbit_r131_c216 bl[216] br[216] wl[131] vdd gnd cell_6t
Xbit_r132_c216 bl[216] br[216] wl[132] vdd gnd cell_6t
Xbit_r133_c216 bl[216] br[216] wl[133] vdd gnd cell_6t
Xbit_r134_c216 bl[216] br[216] wl[134] vdd gnd cell_6t
Xbit_r135_c216 bl[216] br[216] wl[135] vdd gnd cell_6t
Xbit_r136_c216 bl[216] br[216] wl[136] vdd gnd cell_6t
Xbit_r137_c216 bl[216] br[216] wl[137] vdd gnd cell_6t
Xbit_r138_c216 bl[216] br[216] wl[138] vdd gnd cell_6t
Xbit_r139_c216 bl[216] br[216] wl[139] vdd gnd cell_6t
Xbit_r140_c216 bl[216] br[216] wl[140] vdd gnd cell_6t
Xbit_r141_c216 bl[216] br[216] wl[141] vdd gnd cell_6t
Xbit_r142_c216 bl[216] br[216] wl[142] vdd gnd cell_6t
Xbit_r143_c216 bl[216] br[216] wl[143] vdd gnd cell_6t
Xbit_r144_c216 bl[216] br[216] wl[144] vdd gnd cell_6t
Xbit_r145_c216 bl[216] br[216] wl[145] vdd gnd cell_6t
Xbit_r146_c216 bl[216] br[216] wl[146] vdd gnd cell_6t
Xbit_r147_c216 bl[216] br[216] wl[147] vdd gnd cell_6t
Xbit_r148_c216 bl[216] br[216] wl[148] vdd gnd cell_6t
Xbit_r149_c216 bl[216] br[216] wl[149] vdd gnd cell_6t
Xbit_r150_c216 bl[216] br[216] wl[150] vdd gnd cell_6t
Xbit_r151_c216 bl[216] br[216] wl[151] vdd gnd cell_6t
Xbit_r152_c216 bl[216] br[216] wl[152] vdd gnd cell_6t
Xbit_r153_c216 bl[216] br[216] wl[153] vdd gnd cell_6t
Xbit_r154_c216 bl[216] br[216] wl[154] vdd gnd cell_6t
Xbit_r155_c216 bl[216] br[216] wl[155] vdd gnd cell_6t
Xbit_r156_c216 bl[216] br[216] wl[156] vdd gnd cell_6t
Xbit_r157_c216 bl[216] br[216] wl[157] vdd gnd cell_6t
Xbit_r158_c216 bl[216] br[216] wl[158] vdd gnd cell_6t
Xbit_r159_c216 bl[216] br[216] wl[159] vdd gnd cell_6t
Xbit_r160_c216 bl[216] br[216] wl[160] vdd gnd cell_6t
Xbit_r161_c216 bl[216] br[216] wl[161] vdd gnd cell_6t
Xbit_r162_c216 bl[216] br[216] wl[162] vdd gnd cell_6t
Xbit_r163_c216 bl[216] br[216] wl[163] vdd gnd cell_6t
Xbit_r164_c216 bl[216] br[216] wl[164] vdd gnd cell_6t
Xbit_r165_c216 bl[216] br[216] wl[165] vdd gnd cell_6t
Xbit_r166_c216 bl[216] br[216] wl[166] vdd gnd cell_6t
Xbit_r167_c216 bl[216] br[216] wl[167] vdd gnd cell_6t
Xbit_r168_c216 bl[216] br[216] wl[168] vdd gnd cell_6t
Xbit_r169_c216 bl[216] br[216] wl[169] vdd gnd cell_6t
Xbit_r170_c216 bl[216] br[216] wl[170] vdd gnd cell_6t
Xbit_r171_c216 bl[216] br[216] wl[171] vdd gnd cell_6t
Xbit_r172_c216 bl[216] br[216] wl[172] vdd gnd cell_6t
Xbit_r173_c216 bl[216] br[216] wl[173] vdd gnd cell_6t
Xbit_r174_c216 bl[216] br[216] wl[174] vdd gnd cell_6t
Xbit_r175_c216 bl[216] br[216] wl[175] vdd gnd cell_6t
Xbit_r176_c216 bl[216] br[216] wl[176] vdd gnd cell_6t
Xbit_r177_c216 bl[216] br[216] wl[177] vdd gnd cell_6t
Xbit_r178_c216 bl[216] br[216] wl[178] vdd gnd cell_6t
Xbit_r179_c216 bl[216] br[216] wl[179] vdd gnd cell_6t
Xbit_r180_c216 bl[216] br[216] wl[180] vdd gnd cell_6t
Xbit_r181_c216 bl[216] br[216] wl[181] vdd gnd cell_6t
Xbit_r182_c216 bl[216] br[216] wl[182] vdd gnd cell_6t
Xbit_r183_c216 bl[216] br[216] wl[183] vdd gnd cell_6t
Xbit_r184_c216 bl[216] br[216] wl[184] vdd gnd cell_6t
Xbit_r185_c216 bl[216] br[216] wl[185] vdd gnd cell_6t
Xbit_r186_c216 bl[216] br[216] wl[186] vdd gnd cell_6t
Xbit_r187_c216 bl[216] br[216] wl[187] vdd gnd cell_6t
Xbit_r188_c216 bl[216] br[216] wl[188] vdd gnd cell_6t
Xbit_r189_c216 bl[216] br[216] wl[189] vdd gnd cell_6t
Xbit_r190_c216 bl[216] br[216] wl[190] vdd gnd cell_6t
Xbit_r191_c216 bl[216] br[216] wl[191] vdd gnd cell_6t
Xbit_r192_c216 bl[216] br[216] wl[192] vdd gnd cell_6t
Xbit_r193_c216 bl[216] br[216] wl[193] vdd gnd cell_6t
Xbit_r194_c216 bl[216] br[216] wl[194] vdd gnd cell_6t
Xbit_r195_c216 bl[216] br[216] wl[195] vdd gnd cell_6t
Xbit_r196_c216 bl[216] br[216] wl[196] vdd gnd cell_6t
Xbit_r197_c216 bl[216] br[216] wl[197] vdd gnd cell_6t
Xbit_r198_c216 bl[216] br[216] wl[198] vdd gnd cell_6t
Xbit_r199_c216 bl[216] br[216] wl[199] vdd gnd cell_6t
Xbit_r200_c216 bl[216] br[216] wl[200] vdd gnd cell_6t
Xbit_r201_c216 bl[216] br[216] wl[201] vdd gnd cell_6t
Xbit_r202_c216 bl[216] br[216] wl[202] vdd gnd cell_6t
Xbit_r203_c216 bl[216] br[216] wl[203] vdd gnd cell_6t
Xbit_r204_c216 bl[216] br[216] wl[204] vdd gnd cell_6t
Xbit_r205_c216 bl[216] br[216] wl[205] vdd gnd cell_6t
Xbit_r206_c216 bl[216] br[216] wl[206] vdd gnd cell_6t
Xbit_r207_c216 bl[216] br[216] wl[207] vdd gnd cell_6t
Xbit_r208_c216 bl[216] br[216] wl[208] vdd gnd cell_6t
Xbit_r209_c216 bl[216] br[216] wl[209] vdd gnd cell_6t
Xbit_r210_c216 bl[216] br[216] wl[210] vdd gnd cell_6t
Xbit_r211_c216 bl[216] br[216] wl[211] vdd gnd cell_6t
Xbit_r212_c216 bl[216] br[216] wl[212] vdd gnd cell_6t
Xbit_r213_c216 bl[216] br[216] wl[213] vdd gnd cell_6t
Xbit_r214_c216 bl[216] br[216] wl[214] vdd gnd cell_6t
Xbit_r215_c216 bl[216] br[216] wl[215] vdd gnd cell_6t
Xbit_r216_c216 bl[216] br[216] wl[216] vdd gnd cell_6t
Xbit_r217_c216 bl[216] br[216] wl[217] vdd gnd cell_6t
Xbit_r218_c216 bl[216] br[216] wl[218] vdd gnd cell_6t
Xbit_r219_c216 bl[216] br[216] wl[219] vdd gnd cell_6t
Xbit_r220_c216 bl[216] br[216] wl[220] vdd gnd cell_6t
Xbit_r221_c216 bl[216] br[216] wl[221] vdd gnd cell_6t
Xbit_r222_c216 bl[216] br[216] wl[222] vdd gnd cell_6t
Xbit_r223_c216 bl[216] br[216] wl[223] vdd gnd cell_6t
Xbit_r224_c216 bl[216] br[216] wl[224] vdd gnd cell_6t
Xbit_r225_c216 bl[216] br[216] wl[225] vdd gnd cell_6t
Xbit_r226_c216 bl[216] br[216] wl[226] vdd gnd cell_6t
Xbit_r227_c216 bl[216] br[216] wl[227] vdd gnd cell_6t
Xbit_r228_c216 bl[216] br[216] wl[228] vdd gnd cell_6t
Xbit_r229_c216 bl[216] br[216] wl[229] vdd gnd cell_6t
Xbit_r230_c216 bl[216] br[216] wl[230] vdd gnd cell_6t
Xbit_r231_c216 bl[216] br[216] wl[231] vdd gnd cell_6t
Xbit_r232_c216 bl[216] br[216] wl[232] vdd gnd cell_6t
Xbit_r233_c216 bl[216] br[216] wl[233] vdd gnd cell_6t
Xbit_r234_c216 bl[216] br[216] wl[234] vdd gnd cell_6t
Xbit_r235_c216 bl[216] br[216] wl[235] vdd gnd cell_6t
Xbit_r236_c216 bl[216] br[216] wl[236] vdd gnd cell_6t
Xbit_r237_c216 bl[216] br[216] wl[237] vdd gnd cell_6t
Xbit_r238_c216 bl[216] br[216] wl[238] vdd gnd cell_6t
Xbit_r239_c216 bl[216] br[216] wl[239] vdd gnd cell_6t
Xbit_r240_c216 bl[216] br[216] wl[240] vdd gnd cell_6t
Xbit_r241_c216 bl[216] br[216] wl[241] vdd gnd cell_6t
Xbit_r242_c216 bl[216] br[216] wl[242] vdd gnd cell_6t
Xbit_r243_c216 bl[216] br[216] wl[243] vdd gnd cell_6t
Xbit_r244_c216 bl[216] br[216] wl[244] vdd gnd cell_6t
Xbit_r245_c216 bl[216] br[216] wl[245] vdd gnd cell_6t
Xbit_r246_c216 bl[216] br[216] wl[246] vdd gnd cell_6t
Xbit_r247_c216 bl[216] br[216] wl[247] vdd gnd cell_6t
Xbit_r248_c216 bl[216] br[216] wl[248] vdd gnd cell_6t
Xbit_r249_c216 bl[216] br[216] wl[249] vdd gnd cell_6t
Xbit_r250_c216 bl[216] br[216] wl[250] vdd gnd cell_6t
Xbit_r251_c216 bl[216] br[216] wl[251] vdd gnd cell_6t
Xbit_r252_c216 bl[216] br[216] wl[252] vdd gnd cell_6t
Xbit_r253_c216 bl[216] br[216] wl[253] vdd gnd cell_6t
Xbit_r254_c216 bl[216] br[216] wl[254] vdd gnd cell_6t
Xbit_r255_c216 bl[216] br[216] wl[255] vdd gnd cell_6t
Xbit_r0_c217 bl[217] br[217] wl[0] vdd gnd cell_6t
Xbit_r1_c217 bl[217] br[217] wl[1] vdd gnd cell_6t
Xbit_r2_c217 bl[217] br[217] wl[2] vdd gnd cell_6t
Xbit_r3_c217 bl[217] br[217] wl[3] vdd gnd cell_6t
Xbit_r4_c217 bl[217] br[217] wl[4] vdd gnd cell_6t
Xbit_r5_c217 bl[217] br[217] wl[5] vdd gnd cell_6t
Xbit_r6_c217 bl[217] br[217] wl[6] vdd gnd cell_6t
Xbit_r7_c217 bl[217] br[217] wl[7] vdd gnd cell_6t
Xbit_r8_c217 bl[217] br[217] wl[8] vdd gnd cell_6t
Xbit_r9_c217 bl[217] br[217] wl[9] vdd gnd cell_6t
Xbit_r10_c217 bl[217] br[217] wl[10] vdd gnd cell_6t
Xbit_r11_c217 bl[217] br[217] wl[11] vdd gnd cell_6t
Xbit_r12_c217 bl[217] br[217] wl[12] vdd gnd cell_6t
Xbit_r13_c217 bl[217] br[217] wl[13] vdd gnd cell_6t
Xbit_r14_c217 bl[217] br[217] wl[14] vdd gnd cell_6t
Xbit_r15_c217 bl[217] br[217] wl[15] vdd gnd cell_6t
Xbit_r16_c217 bl[217] br[217] wl[16] vdd gnd cell_6t
Xbit_r17_c217 bl[217] br[217] wl[17] vdd gnd cell_6t
Xbit_r18_c217 bl[217] br[217] wl[18] vdd gnd cell_6t
Xbit_r19_c217 bl[217] br[217] wl[19] vdd gnd cell_6t
Xbit_r20_c217 bl[217] br[217] wl[20] vdd gnd cell_6t
Xbit_r21_c217 bl[217] br[217] wl[21] vdd gnd cell_6t
Xbit_r22_c217 bl[217] br[217] wl[22] vdd gnd cell_6t
Xbit_r23_c217 bl[217] br[217] wl[23] vdd gnd cell_6t
Xbit_r24_c217 bl[217] br[217] wl[24] vdd gnd cell_6t
Xbit_r25_c217 bl[217] br[217] wl[25] vdd gnd cell_6t
Xbit_r26_c217 bl[217] br[217] wl[26] vdd gnd cell_6t
Xbit_r27_c217 bl[217] br[217] wl[27] vdd gnd cell_6t
Xbit_r28_c217 bl[217] br[217] wl[28] vdd gnd cell_6t
Xbit_r29_c217 bl[217] br[217] wl[29] vdd gnd cell_6t
Xbit_r30_c217 bl[217] br[217] wl[30] vdd gnd cell_6t
Xbit_r31_c217 bl[217] br[217] wl[31] vdd gnd cell_6t
Xbit_r32_c217 bl[217] br[217] wl[32] vdd gnd cell_6t
Xbit_r33_c217 bl[217] br[217] wl[33] vdd gnd cell_6t
Xbit_r34_c217 bl[217] br[217] wl[34] vdd gnd cell_6t
Xbit_r35_c217 bl[217] br[217] wl[35] vdd gnd cell_6t
Xbit_r36_c217 bl[217] br[217] wl[36] vdd gnd cell_6t
Xbit_r37_c217 bl[217] br[217] wl[37] vdd gnd cell_6t
Xbit_r38_c217 bl[217] br[217] wl[38] vdd gnd cell_6t
Xbit_r39_c217 bl[217] br[217] wl[39] vdd gnd cell_6t
Xbit_r40_c217 bl[217] br[217] wl[40] vdd gnd cell_6t
Xbit_r41_c217 bl[217] br[217] wl[41] vdd gnd cell_6t
Xbit_r42_c217 bl[217] br[217] wl[42] vdd gnd cell_6t
Xbit_r43_c217 bl[217] br[217] wl[43] vdd gnd cell_6t
Xbit_r44_c217 bl[217] br[217] wl[44] vdd gnd cell_6t
Xbit_r45_c217 bl[217] br[217] wl[45] vdd gnd cell_6t
Xbit_r46_c217 bl[217] br[217] wl[46] vdd gnd cell_6t
Xbit_r47_c217 bl[217] br[217] wl[47] vdd gnd cell_6t
Xbit_r48_c217 bl[217] br[217] wl[48] vdd gnd cell_6t
Xbit_r49_c217 bl[217] br[217] wl[49] vdd gnd cell_6t
Xbit_r50_c217 bl[217] br[217] wl[50] vdd gnd cell_6t
Xbit_r51_c217 bl[217] br[217] wl[51] vdd gnd cell_6t
Xbit_r52_c217 bl[217] br[217] wl[52] vdd gnd cell_6t
Xbit_r53_c217 bl[217] br[217] wl[53] vdd gnd cell_6t
Xbit_r54_c217 bl[217] br[217] wl[54] vdd gnd cell_6t
Xbit_r55_c217 bl[217] br[217] wl[55] vdd gnd cell_6t
Xbit_r56_c217 bl[217] br[217] wl[56] vdd gnd cell_6t
Xbit_r57_c217 bl[217] br[217] wl[57] vdd gnd cell_6t
Xbit_r58_c217 bl[217] br[217] wl[58] vdd gnd cell_6t
Xbit_r59_c217 bl[217] br[217] wl[59] vdd gnd cell_6t
Xbit_r60_c217 bl[217] br[217] wl[60] vdd gnd cell_6t
Xbit_r61_c217 bl[217] br[217] wl[61] vdd gnd cell_6t
Xbit_r62_c217 bl[217] br[217] wl[62] vdd gnd cell_6t
Xbit_r63_c217 bl[217] br[217] wl[63] vdd gnd cell_6t
Xbit_r64_c217 bl[217] br[217] wl[64] vdd gnd cell_6t
Xbit_r65_c217 bl[217] br[217] wl[65] vdd gnd cell_6t
Xbit_r66_c217 bl[217] br[217] wl[66] vdd gnd cell_6t
Xbit_r67_c217 bl[217] br[217] wl[67] vdd gnd cell_6t
Xbit_r68_c217 bl[217] br[217] wl[68] vdd gnd cell_6t
Xbit_r69_c217 bl[217] br[217] wl[69] vdd gnd cell_6t
Xbit_r70_c217 bl[217] br[217] wl[70] vdd gnd cell_6t
Xbit_r71_c217 bl[217] br[217] wl[71] vdd gnd cell_6t
Xbit_r72_c217 bl[217] br[217] wl[72] vdd gnd cell_6t
Xbit_r73_c217 bl[217] br[217] wl[73] vdd gnd cell_6t
Xbit_r74_c217 bl[217] br[217] wl[74] vdd gnd cell_6t
Xbit_r75_c217 bl[217] br[217] wl[75] vdd gnd cell_6t
Xbit_r76_c217 bl[217] br[217] wl[76] vdd gnd cell_6t
Xbit_r77_c217 bl[217] br[217] wl[77] vdd gnd cell_6t
Xbit_r78_c217 bl[217] br[217] wl[78] vdd gnd cell_6t
Xbit_r79_c217 bl[217] br[217] wl[79] vdd gnd cell_6t
Xbit_r80_c217 bl[217] br[217] wl[80] vdd gnd cell_6t
Xbit_r81_c217 bl[217] br[217] wl[81] vdd gnd cell_6t
Xbit_r82_c217 bl[217] br[217] wl[82] vdd gnd cell_6t
Xbit_r83_c217 bl[217] br[217] wl[83] vdd gnd cell_6t
Xbit_r84_c217 bl[217] br[217] wl[84] vdd gnd cell_6t
Xbit_r85_c217 bl[217] br[217] wl[85] vdd gnd cell_6t
Xbit_r86_c217 bl[217] br[217] wl[86] vdd gnd cell_6t
Xbit_r87_c217 bl[217] br[217] wl[87] vdd gnd cell_6t
Xbit_r88_c217 bl[217] br[217] wl[88] vdd gnd cell_6t
Xbit_r89_c217 bl[217] br[217] wl[89] vdd gnd cell_6t
Xbit_r90_c217 bl[217] br[217] wl[90] vdd gnd cell_6t
Xbit_r91_c217 bl[217] br[217] wl[91] vdd gnd cell_6t
Xbit_r92_c217 bl[217] br[217] wl[92] vdd gnd cell_6t
Xbit_r93_c217 bl[217] br[217] wl[93] vdd gnd cell_6t
Xbit_r94_c217 bl[217] br[217] wl[94] vdd gnd cell_6t
Xbit_r95_c217 bl[217] br[217] wl[95] vdd gnd cell_6t
Xbit_r96_c217 bl[217] br[217] wl[96] vdd gnd cell_6t
Xbit_r97_c217 bl[217] br[217] wl[97] vdd gnd cell_6t
Xbit_r98_c217 bl[217] br[217] wl[98] vdd gnd cell_6t
Xbit_r99_c217 bl[217] br[217] wl[99] vdd gnd cell_6t
Xbit_r100_c217 bl[217] br[217] wl[100] vdd gnd cell_6t
Xbit_r101_c217 bl[217] br[217] wl[101] vdd gnd cell_6t
Xbit_r102_c217 bl[217] br[217] wl[102] vdd gnd cell_6t
Xbit_r103_c217 bl[217] br[217] wl[103] vdd gnd cell_6t
Xbit_r104_c217 bl[217] br[217] wl[104] vdd gnd cell_6t
Xbit_r105_c217 bl[217] br[217] wl[105] vdd gnd cell_6t
Xbit_r106_c217 bl[217] br[217] wl[106] vdd gnd cell_6t
Xbit_r107_c217 bl[217] br[217] wl[107] vdd gnd cell_6t
Xbit_r108_c217 bl[217] br[217] wl[108] vdd gnd cell_6t
Xbit_r109_c217 bl[217] br[217] wl[109] vdd gnd cell_6t
Xbit_r110_c217 bl[217] br[217] wl[110] vdd gnd cell_6t
Xbit_r111_c217 bl[217] br[217] wl[111] vdd gnd cell_6t
Xbit_r112_c217 bl[217] br[217] wl[112] vdd gnd cell_6t
Xbit_r113_c217 bl[217] br[217] wl[113] vdd gnd cell_6t
Xbit_r114_c217 bl[217] br[217] wl[114] vdd gnd cell_6t
Xbit_r115_c217 bl[217] br[217] wl[115] vdd gnd cell_6t
Xbit_r116_c217 bl[217] br[217] wl[116] vdd gnd cell_6t
Xbit_r117_c217 bl[217] br[217] wl[117] vdd gnd cell_6t
Xbit_r118_c217 bl[217] br[217] wl[118] vdd gnd cell_6t
Xbit_r119_c217 bl[217] br[217] wl[119] vdd gnd cell_6t
Xbit_r120_c217 bl[217] br[217] wl[120] vdd gnd cell_6t
Xbit_r121_c217 bl[217] br[217] wl[121] vdd gnd cell_6t
Xbit_r122_c217 bl[217] br[217] wl[122] vdd gnd cell_6t
Xbit_r123_c217 bl[217] br[217] wl[123] vdd gnd cell_6t
Xbit_r124_c217 bl[217] br[217] wl[124] vdd gnd cell_6t
Xbit_r125_c217 bl[217] br[217] wl[125] vdd gnd cell_6t
Xbit_r126_c217 bl[217] br[217] wl[126] vdd gnd cell_6t
Xbit_r127_c217 bl[217] br[217] wl[127] vdd gnd cell_6t
Xbit_r128_c217 bl[217] br[217] wl[128] vdd gnd cell_6t
Xbit_r129_c217 bl[217] br[217] wl[129] vdd gnd cell_6t
Xbit_r130_c217 bl[217] br[217] wl[130] vdd gnd cell_6t
Xbit_r131_c217 bl[217] br[217] wl[131] vdd gnd cell_6t
Xbit_r132_c217 bl[217] br[217] wl[132] vdd gnd cell_6t
Xbit_r133_c217 bl[217] br[217] wl[133] vdd gnd cell_6t
Xbit_r134_c217 bl[217] br[217] wl[134] vdd gnd cell_6t
Xbit_r135_c217 bl[217] br[217] wl[135] vdd gnd cell_6t
Xbit_r136_c217 bl[217] br[217] wl[136] vdd gnd cell_6t
Xbit_r137_c217 bl[217] br[217] wl[137] vdd gnd cell_6t
Xbit_r138_c217 bl[217] br[217] wl[138] vdd gnd cell_6t
Xbit_r139_c217 bl[217] br[217] wl[139] vdd gnd cell_6t
Xbit_r140_c217 bl[217] br[217] wl[140] vdd gnd cell_6t
Xbit_r141_c217 bl[217] br[217] wl[141] vdd gnd cell_6t
Xbit_r142_c217 bl[217] br[217] wl[142] vdd gnd cell_6t
Xbit_r143_c217 bl[217] br[217] wl[143] vdd gnd cell_6t
Xbit_r144_c217 bl[217] br[217] wl[144] vdd gnd cell_6t
Xbit_r145_c217 bl[217] br[217] wl[145] vdd gnd cell_6t
Xbit_r146_c217 bl[217] br[217] wl[146] vdd gnd cell_6t
Xbit_r147_c217 bl[217] br[217] wl[147] vdd gnd cell_6t
Xbit_r148_c217 bl[217] br[217] wl[148] vdd gnd cell_6t
Xbit_r149_c217 bl[217] br[217] wl[149] vdd gnd cell_6t
Xbit_r150_c217 bl[217] br[217] wl[150] vdd gnd cell_6t
Xbit_r151_c217 bl[217] br[217] wl[151] vdd gnd cell_6t
Xbit_r152_c217 bl[217] br[217] wl[152] vdd gnd cell_6t
Xbit_r153_c217 bl[217] br[217] wl[153] vdd gnd cell_6t
Xbit_r154_c217 bl[217] br[217] wl[154] vdd gnd cell_6t
Xbit_r155_c217 bl[217] br[217] wl[155] vdd gnd cell_6t
Xbit_r156_c217 bl[217] br[217] wl[156] vdd gnd cell_6t
Xbit_r157_c217 bl[217] br[217] wl[157] vdd gnd cell_6t
Xbit_r158_c217 bl[217] br[217] wl[158] vdd gnd cell_6t
Xbit_r159_c217 bl[217] br[217] wl[159] vdd gnd cell_6t
Xbit_r160_c217 bl[217] br[217] wl[160] vdd gnd cell_6t
Xbit_r161_c217 bl[217] br[217] wl[161] vdd gnd cell_6t
Xbit_r162_c217 bl[217] br[217] wl[162] vdd gnd cell_6t
Xbit_r163_c217 bl[217] br[217] wl[163] vdd gnd cell_6t
Xbit_r164_c217 bl[217] br[217] wl[164] vdd gnd cell_6t
Xbit_r165_c217 bl[217] br[217] wl[165] vdd gnd cell_6t
Xbit_r166_c217 bl[217] br[217] wl[166] vdd gnd cell_6t
Xbit_r167_c217 bl[217] br[217] wl[167] vdd gnd cell_6t
Xbit_r168_c217 bl[217] br[217] wl[168] vdd gnd cell_6t
Xbit_r169_c217 bl[217] br[217] wl[169] vdd gnd cell_6t
Xbit_r170_c217 bl[217] br[217] wl[170] vdd gnd cell_6t
Xbit_r171_c217 bl[217] br[217] wl[171] vdd gnd cell_6t
Xbit_r172_c217 bl[217] br[217] wl[172] vdd gnd cell_6t
Xbit_r173_c217 bl[217] br[217] wl[173] vdd gnd cell_6t
Xbit_r174_c217 bl[217] br[217] wl[174] vdd gnd cell_6t
Xbit_r175_c217 bl[217] br[217] wl[175] vdd gnd cell_6t
Xbit_r176_c217 bl[217] br[217] wl[176] vdd gnd cell_6t
Xbit_r177_c217 bl[217] br[217] wl[177] vdd gnd cell_6t
Xbit_r178_c217 bl[217] br[217] wl[178] vdd gnd cell_6t
Xbit_r179_c217 bl[217] br[217] wl[179] vdd gnd cell_6t
Xbit_r180_c217 bl[217] br[217] wl[180] vdd gnd cell_6t
Xbit_r181_c217 bl[217] br[217] wl[181] vdd gnd cell_6t
Xbit_r182_c217 bl[217] br[217] wl[182] vdd gnd cell_6t
Xbit_r183_c217 bl[217] br[217] wl[183] vdd gnd cell_6t
Xbit_r184_c217 bl[217] br[217] wl[184] vdd gnd cell_6t
Xbit_r185_c217 bl[217] br[217] wl[185] vdd gnd cell_6t
Xbit_r186_c217 bl[217] br[217] wl[186] vdd gnd cell_6t
Xbit_r187_c217 bl[217] br[217] wl[187] vdd gnd cell_6t
Xbit_r188_c217 bl[217] br[217] wl[188] vdd gnd cell_6t
Xbit_r189_c217 bl[217] br[217] wl[189] vdd gnd cell_6t
Xbit_r190_c217 bl[217] br[217] wl[190] vdd gnd cell_6t
Xbit_r191_c217 bl[217] br[217] wl[191] vdd gnd cell_6t
Xbit_r192_c217 bl[217] br[217] wl[192] vdd gnd cell_6t
Xbit_r193_c217 bl[217] br[217] wl[193] vdd gnd cell_6t
Xbit_r194_c217 bl[217] br[217] wl[194] vdd gnd cell_6t
Xbit_r195_c217 bl[217] br[217] wl[195] vdd gnd cell_6t
Xbit_r196_c217 bl[217] br[217] wl[196] vdd gnd cell_6t
Xbit_r197_c217 bl[217] br[217] wl[197] vdd gnd cell_6t
Xbit_r198_c217 bl[217] br[217] wl[198] vdd gnd cell_6t
Xbit_r199_c217 bl[217] br[217] wl[199] vdd gnd cell_6t
Xbit_r200_c217 bl[217] br[217] wl[200] vdd gnd cell_6t
Xbit_r201_c217 bl[217] br[217] wl[201] vdd gnd cell_6t
Xbit_r202_c217 bl[217] br[217] wl[202] vdd gnd cell_6t
Xbit_r203_c217 bl[217] br[217] wl[203] vdd gnd cell_6t
Xbit_r204_c217 bl[217] br[217] wl[204] vdd gnd cell_6t
Xbit_r205_c217 bl[217] br[217] wl[205] vdd gnd cell_6t
Xbit_r206_c217 bl[217] br[217] wl[206] vdd gnd cell_6t
Xbit_r207_c217 bl[217] br[217] wl[207] vdd gnd cell_6t
Xbit_r208_c217 bl[217] br[217] wl[208] vdd gnd cell_6t
Xbit_r209_c217 bl[217] br[217] wl[209] vdd gnd cell_6t
Xbit_r210_c217 bl[217] br[217] wl[210] vdd gnd cell_6t
Xbit_r211_c217 bl[217] br[217] wl[211] vdd gnd cell_6t
Xbit_r212_c217 bl[217] br[217] wl[212] vdd gnd cell_6t
Xbit_r213_c217 bl[217] br[217] wl[213] vdd gnd cell_6t
Xbit_r214_c217 bl[217] br[217] wl[214] vdd gnd cell_6t
Xbit_r215_c217 bl[217] br[217] wl[215] vdd gnd cell_6t
Xbit_r216_c217 bl[217] br[217] wl[216] vdd gnd cell_6t
Xbit_r217_c217 bl[217] br[217] wl[217] vdd gnd cell_6t
Xbit_r218_c217 bl[217] br[217] wl[218] vdd gnd cell_6t
Xbit_r219_c217 bl[217] br[217] wl[219] vdd gnd cell_6t
Xbit_r220_c217 bl[217] br[217] wl[220] vdd gnd cell_6t
Xbit_r221_c217 bl[217] br[217] wl[221] vdd gnd cell_6t
Xbit_r222_c217 bl[217] br[217] wl[222] vdd gnd cell_6t
Xbit_r223_c217 bl[217] br[217] wl[223] vdd gnd cell_6t
Xbit_r224_c217 bl[217] br[217] wl[224] vdd gnd cell_6t
Xbit_r225_c217 bl[217] br[217] wl[225] vdd gnd cell_6t
Xbit_r226_c217 bl[217] br[217] wl[226] vdd gnd cell_6t
Xbit_r227_c217 bl[217] br[217] wl[227] vdd gnd cell_6t
Xbit_r228_c217 bl[217] br[217] wl[228] vdd gnd cell_6t
Xbit_r229_c217 bl[217] br[217] wl[229] vdd gnd cell_6t
Xbit_r230_c217 bl[217] br[217] wl[230] vdd gnd cell_6t
Xbit_r231_c217 bl[217] br[217] wl[231] vdd gnd cell_6t
Xbit_r232_c217 bl[217] br[217] wl[232] vdd gnd cell_6t
Xbit_r233_c217 bl[217] br[217] wl[233] vdd gnd cell_6t
Xbit_r234_c217 bl[217] br[217] wl[234] vdd gnd cell_6t
Xbit_r235_c217 bl[217] br[217] wl[235] vdd gnd cell_6t
Xbit_r236_c217 bl[217] br[217] wl[236] vdd gnd cell_6t
Xbit_r237_c217 bl[217] br[217] wl[237] vdd gnd cell_6t
Xbit_r238_c217 bl[217] br[217] wl[238] vdd gnd cell_6t
Xbit_r239_c217 bl[217] br[217] wl[239] vdd gnd cell_6t
Xbit_r240_c217 bl[217] br[217] wl[240] vdd gnd cell_6t
Xbit_r241_c217 bl[217] br[217] wl[241] vdd gnd cell_6t
Xbit_r242_c217 bl[217] br[217] wl[242] vdd gnd cell_6t
Xbit_r243_c217 bl[217] br[217] wl[243] vdd gnd cell_6t
Xbit_r244_c217 bl[217] br[217] wl[244] vdd gnd cell_6t
Xbit_r245_c217 bl[217] br[217] wl[245] vdd gnd cell_6t
Xbit_r246_c217 bl[217] br[217] wl[246] vdd gnd cell_6t
Xbit_r247_c217 bl[217] br[217] wl[247] vdd gnd cell_6t
Xbit_r248_c217 bl[217] br[217] wl[248] vdd gnd cell_6t
Xbit_r249_c217 bl[217] br[217] wl[249] vdd gnd cell_6t
Xbit_r250_c217 bl[217] br[217] wl[250] vdd gnd cell_6t
Xbit_r251_c217 bl[217] br[217] wl[251] vdd gnd cell_6t
Xbit_r252_c217 bl[217] br[217] wl[252] vdd gnd cell_6t
Xbit_r253_c217 bl[217] br[217] wl[253] vdd gnd cell_6t
Xbit_r254_c217 bl[217] br[217] wl[254] vdd gnd cell_6t
Xbit_r255_c217 bl[217] br[217] wl[255] vdd gnd cell_6t
Xbit_r0_c218 bl[218] br[218] wl[0] vdd gnd cell_6t
Xbit_r1_c218 bl[218] br[218] wl[1] vdd gnd cell_6t
Xbit_r2_c218 bl[218] br[218] wl[2] vdd gnd cell_6t
Xbit_r3_c218 bl[218] br[218] wl[3] vdd gnd cell_6t
Xbit_r4_c218 bl[218] br[218] wl[4] vdd gnd cell_6t
Xbit_r5_c218 bl[218] br[218] wl[5] vdd gnd cell_6t
Xbit_r6_c218 bl[218] br[218] wl[6] vdd gnd cell_6t
Xbit_r7_c218 bl[218] br[218] wl[7] vdd gnd cell_6t
Xbit_r8_c218 bl[218] br[218] wl[8] vdd gnd cell_6t
Xbit_r9_c218 bl[218] br[218] wl[9] vdd gnd cell_6t
Xbit_r10_c218 bl[218] br[218] wl[10] vdd gnd cell_6t
Xbit_r11_c218 bl[218] br[218] wl[11] vdd gnd cell_6t
Xbit_r12_c218 bl[218] br[218] wl[12] vdd gnd cell_6t
Xbit_r13_c218 bl[218] br[218] wl[13] vdd gnd cell_6t
Xbit_r14_c218 bl[218] br[218] wl[14] vdd gnd cell_6t
Xbit_r15_c218 bl[218] br[218] wl[15] vdd gnd cell_6t
Xbit_r16_c218 bl[218] br[218] wl[16] vdd gnd cell_6t
Xbit_r17_c218 bl[218] br[218] wl[17] vdd gnd cell_6t
Xbit_r18_c218 bl[218] br[218] wl[18] vdd gnd cell_6t
Xbit_r19_c218 bl[218] br[218] wl[19] vdd gnd cell_6t
Xbit_r20_c218 bl[218] br[218] wl[20] vdd gnd cell_6t
Xbit_r21_c218 bl[218] br[218] wl[21] vdd gnd cell_6t
Xbit_r22_c218 bl[218] br[218] wl[22] vdd gnd cell_6t
Xbit_r23_c218 bl[218] br[218] wl[23] vdd gnd cell_6t
Xbit_r24_c218 bl[218] br[218] wl[24] vdd gnd cell_6t
Xbit_r25_c218 bl[218] br[218] wl[25] vdd gnd cell_6t
Xbit_r26_c218 bl[218] br[218] wl[26] vdd gnd cell_6t
Xbit_r27_c218 bl[218] br[218] wl[27] vdd gnd cell_6t
Xbit_r28_c218 bl[218] br[218] wl[28] vdd gnd cell_6t
Xbit_r29_c218 bl[218] br[218] wl[29] vdd gnd cell_6t
Xbit_r30_c218 bl[218] br[218] wl[30] vdd gnd cell_6t
Xbit_r31_c218 bl[218] br[218] wl[31] vdd gnd cell_6t
Xbit_r32_c218 bl[218] br[218] wl[32] vdd gnd cell_6t
Xbit_r33_c218 bl[218] br[218] wl[33] vdd gnd cell_6t
Xbit_r34_c218 bl[218] br[218] wl[34] vdd gnd cell_6t
Xbit_r35_c218 bl[218] br[218] wl[35] vdd gnd cell_6t
Xbit_r36_c218 bl[218] br[218] wl[36] vdd gnd cell_6t
Xbit_r37_c218 bl[218] br[218] wl[37] vdd gnd cell_6t
Xbit_r38_c218 bl[218] br[218] wl[38] vdd gnd cell_6t
Xbit_r39_c218 bl[218] br[218] wl[39] vdd gnd cell_6t
Xbit_r40_c218 bl[218] br[218] wl[40] vdd gnd cell_6t
Xbit_r41_c218 bl[218] br[218] wl[41] vdd gnd cell_6t
Xbit_r42_c218 bl[218] br[218] wl[42] vdd gnd cell_6t
Xbit_r43_c218 bl[218] br[218] wl[43] vdd gnd cell_6t
Xbit_r44_c218 bl[218] br[218] wl[44] vdd gnd cell_6t
Xbit_r45_c218 bl[218] br[218] wl[45] vdd gnd cell_6t
Xbit_r46_c218 bl[218] br[218] wl[46] vdd gnd cell_6t
Xbit_r47_c218 bl[218] br[218] wl[47] vdd gnd cell_6t
Xbit_r48_c218 bl[218] br[218] wl[48] vdd gnd cell_6t
Xbit_r49_c218 bl[218] br[218] wl[49] vdd gnd cell_6t
Xbit_r50_c218 bl[218] br[218] wl[50] vdd gnd cell_6t
Xbit_r51_c218 bl[218] br[218] wl[51] vdd gnd cell_6t
Xbit_r52_c218 bl[218] br[218] wl[52] vdd gnd cell_6t
Xbit_r53_c218 bl[218] br[218] wl[53] vdd gnd cell_6t
Xbit_r54_c218 bl[218] br[218] wl[54] vdd gnd cell_6t
Xbit_r55_c218 bl[218] br[218] wl[55] vdd gnd cell_6t
Xbit_r56_c218 bl[218] br[218] wl[56] vdd gnd cell_6t
Xbit_r57_c218 bl[218] br[218] wl[57] vdd gnd cell_6t
Xbit_r58_c218 bl[218] br[218] wl[58] vdd gnd cell_6t
Xbit_r59_c218 bl[218] br[218] wl[59] vdd gnd cell_6t
Xbit_r60_c218 bl[218] br[218] wl[60] vdd gnd cell_6t
Xbit_r61_c218 bl[218] br[218] wl[61] vdd gnd cell_6t
Xbit_r62_c218 bl[218] br[218] wl[62] vdd gnd cell_6t
Xbit_r63_c218 bl[218] br[218] wl[63] vdd gnd cell_6t
Xbit_r64_c218 bl[218] br[218] wl[64] vdd gnd cell_6t
Xbit_r65_c218 bl[218] br[218] wl[65] vdd gnd cell_6t
Xbit_r66_c218 bl[218] br[218] wl[66] vdd gnd cell_6t
Xbit_r67_c218 bl[218] br[218] wl[67] vdd gnd cell_6t
Xbit_r68_c218 bl[218] br[218] wl[68] vdd gnd cell_6t
Xbit_r69_c218 bl[218] br[218] wl[69] vdd gnd cell_6t
Xbit_r70_c218 bl[218] br[218] wl[70] vdd gnd cell_6t
Xbit_r71_c218 bl[218] br[218] wl[71] vdd gnd cell_6t
Xbit_r72_c218 bl[218] br[218] wl[72] vdd gnd cell_6t
Xbit_r73_c218 bl[218] br[218] wl[73] vdd gnd cell_6t
Xbit_r74_c218 bl[218] br[218] wl[74] vdd gnd cell_6t
Xbit_r75_c218 bl[218] br[218] wl[75] vdd gnd cell_6t
Xbit_r76_c218 bl[218] br[218] wl[76] vdd gnd cell_6t
Xbit_r77_c218 bl[218] br[218] wl[77] vdd gnd cell_6t
Xbit_r78_c218 bl[218] br[218] wl[78] vdd gnd cell_6t
Xbit_r79_c218 bl[218] br[218] wl[79] vdd gnd cell_6t
Xbit_r80_c218 bl[218] br[218] wl[80] vdd gnd cell_6t
Xbit_r81_c218 bl[218] br[218] wl[81] vdd gnd cell_6t
Xbit_r82_c218 bl[218] br[218] wl[82] vdd gnd cell_6t
Xbit_r83_c218 bl[218] br[218] wl[83] vdd gnd cell_6t
Xbit_r84_c218 bl[218] br[218] wl[84] vdd gnd cell_6t
Xbit_r85_c218 bl[218] br[218] wl[85] vdd gnd cell_6t
Xbit_r86_c218 bl[218] br[218] wl[86] vdd gnd cell_6t
Xbit_r87_c218 bl[218] br[218] wl[87] vdd gnd cell_6t
Xbit_r88_c218 bl[218] br[218] wl[88] vdd gnd cell_6t
Xbit_r89_c218 bl[218] br[218] wl[89] vdd gnd cell_6t
Xbit_r90_c218 bl[218] br[218] wl[90] vdd gnd cell_6t
Xbit_r91_c218 bl[218] br[218] wl[91] vdd gnd cell_6t
Xbit_r92_c218 bl[218] br[218] wl[92] vdd gnd cell_6t
Xbit_r93_c218 bl[218] br[218] wl[93] vdd gnd cell_6t
Xbit_r94_c218 bl[218] br[218] wl[94] vdd gnd cell_6t
Xbit_r95_c218 bl[218] br[218] wl[95] vdd gnd cell_6t
Xbit_r96_c218 bl[218] br[218] wl[96] vdd gnd cell_6t
Xbit_r97_c218 bl[218] br[218] wl[97] vdd gnd cell_6t
Xbit_r98_c218 bl[218] br[218] wl[98] vdd gnd cell_6t
Xbit_r99_c218 bl[218] br[218] wl[99] vdd gnd cell_6t
Xbit_r100_c218 bl[218] br[218] wl[100] vdd gnd cell_6t
Xbit_r101_c218 bl[218] br[218] wl[101] vdd gnd cell_6t
Xbit_r102_c218 bl[218] br[218] wl[102] vdd gnd cell_6t
Xbit_r103_c218 bl[218] br[218] wl[103] vdd gnd cell_6t
Xbit_r104_c218 bl[218] br[218] wl[104] vdd gnd cell_6t
Xbit_r105_c218 bl[218] br[218] wl[105] vdd gnd cell_6t
Xbit_r106_c218 bl[218] br[218] wl[106] vdd gnd cell_6t
Xbit_r107_c218 bl[218] br[218] wl[107] vdd gnd cell_6t
Xbit_r108_c218 bl[218] br[218] wl[108] vdd gnd cell_6t
Xbit_r109_c218 bl[218] br[218] wl[109] vdd gnd cell_6t
Xbit_r110_c218 bl[218] br[218] wl[110] vdd gnd cell_6t
Xbit_r111_c218 bl[218] br[218] wl[111] vdd gnd cell_6t
Xbit_r112_c218 bl[218] br[218] wl[112] vdd gnd cell_6t
Xbit_r113_c218 bl[218] br[218] wl[113] vdd gnd cell_6t
Xbit_r114_c218 bl[218] br[218] wl[114] vdd gnd cell_6t
Xbit_r115_c218 bl[218] br[218] wl[115] vdd gnd cell_6t
Xbit_r116_c218 bl[218] br[218] wl[116] vdd gnd cell_6t
Xbit_r117_c218 bl[218] br[218] wl[117] vdd gnd cell_6t
Xbit_r118_c218 bl[218] br[218] wl[118] vdd gnd cell_6t
Xbit_r119_c218 bl[218] br[218] wl[119] vdd gnd cell_6t
Xbit_r120_c218 bl[218] br[218] wl[120] vdd gnd cell_6t
Xbit_r121_c218 bl[218] br[218] wl[121] vdd gnd cell_6t
Xbit_r122_c218 bl[218] br[218] wl[122] vdd gnd cell_6t
Xbit_r123_c218 bl[218] br[218] wl[123] vdd gnd cell_6t
Xbit_r124_c218 bl[218] br[218] wl[124] vdd gnd cell_6t
Xbit_r125_c218 bl[218] br[218] wl[125] vdd gnd cell_6t
Xbit_r126_c218 bl[218] br[218] wl[126] vdd gnd cell_6t
Xbit_r127_c218 bl[218] br[218] wl[127] vdd gnd cell_6t
Xbit_r128_c218 bl[218] br[218] wl[128] vdd gnd cell_6t
Xbit_r129_c218 bl[218] br[218] wl[129] vdd gnd cell_6t
Xbit_r130_c218 bl[218] br[218] wl[130] vdd gnd cell_6t
Xbit_r131_c218 bl[218] br[218] wl[131] vdd gnd cell_6t
Xbit_r132_c218 bl[218] br[218] wl[132] vdd gnd cell_6t
Xbit_r133_c218 bl[218] br[218] wl[133] vdd gnd cell_6t
Xbit_r134_c218 bl[218] br[218] wl[134] vdd gnd cell_6t
Xbit_r135_c218 bl[218] br[218] wl[135] vdd gnd cell_6t
Xbit_r136_c218 bl[218] br[218] wl[136] vdd gnd cell_6t
Xbit_r137_c218 bl[218] br[218] wl[137] vdd gnd cell_6t
Xbit_r138_c218 bl[218] br[218] wl[138] vdd gnd cell_6t
Xbit_r139_c218 bl[218] br[218] wl[139] vdd gnd cell_6t
Xbit_r140_c218 bl[218] br[218] wl[140] vdd gnd cell_6t
Xbit_r141_c218 bl[218] br[218] wl[141] vdd gnd cell_6t
Xbit_r142_c218 bl[218] br[218] wl[142] vdd gnd cell_6t
Xbit_r143_c218 bl[218] br[218] wl[143] vdd gnd cell_6t
Xbit_r144_c218 bl[218] br[218] wl[144] vdd gnd cell_6t
Xbit_r145_c218 bl[218] br[218] wl[145] vdd gnd cell_6t
Xbit_r146_c218 bl[218] br[218] wl[146] vdd gnd cell_6t
Xbit_r147_c218 bl[218] br[218] wl[147] vdd gnd cell_6t
Xbit_r148_c218 bl[218] br[218] wl[148] vdd gnd cell_6t
Xbit_r149_c218 bl[218] br[218] wl[149] vdd gnd cell_6t
Xbit_r150_c218 bl[218] br[218] wl[150] vdd gnd cell_6t
Xbit_r151_c218 bl[218] br[218] wl[151] vdd gnd cell_6t
Xbit_r152_c218 bl[218] br[218] wl[152] vdd gnd cell_6t
Xbit_r153_c218 bl[218] br[218] wl[153] vdd gnd cell_6t
Xbit_r154_c218 bl[218] br[218] wl[154] vdd gnd cell_6t
Xbit_r155_c218 bl[218] br[218] wl[155] vdd gnd cell_6t
Xbit_r156_c218 bl[218] br[218] wl[156] vdd gnd cell_6t
Xbit_r157_c218 bl[218] br[218] wl[157] vdd gnd cell_6t
Xbit_r158_c218 bl[218] br[218] wl[158] vdd gnd cell_6t
Xbit_r159_c218 bl[218] br[218] wl[159] vdd gnd cell_6t
Xbit_r160_c218 bl[218] br[218] wl[160] vdd gnd cell_6t
Xbit_r161_c218 bl[218] br[218] wl[161] vdd gnd cell_6t
Xbit_r162_c218 bl[218] br[218] wl[162] vdd gnd cell_6t
Xbit_r163_c218 bl[218] br[218] wl[163] vdd gnd cell_6t
Xbit_r164_c218 bl[218] br[218] wl[164] vdd gnd cell_6t
Xbit_r165_c218 bl[218] br[218] wl[165] vdd gnd cell_6t
Xbit_r166_c218 bl[218] br[218] wl[166] vdd gnd cell_6t
Xbit_r167_c218 bl[218] br[218] wl[167] vdd gnd cell_6t
Xbit_r168_c218 bl[218] br[218] wl[168] vdd gnd cell_6t
Xbit_r169_c218 bl[218] br[218] wl[169] vdd gnd cell_6t
Xbit_r170_c218 bl[218] br[218] wl[170] vdd gnd cell_6t
Xbit_r171_c218 bl[218] br[218] wl[171] vdd gnd cell_6t
Xbit_r172_c218 bl[218] br[218] wl[172] vdd gnd cell_6t
Xbit_r173_c218 bl[218] br[218] wl[173] vdd gnd cell_6t
Xbit_r174_c218 bl[218] br[218] wl[174] vdd gnd cell_6t
Xbit_r175_c218 bl[218] br[218] wl[175] vdd gnd cell_6t
Xbit_r176_c218 bl[218] br[218] wl[176] vdd gnd cell_6t
Xbit_r177_c218 bl[218] br[218] wl[177] vdd gnd cell_6t
Xbit_r178_c218 bl[218] br[218] wl[178] vdd gnd cell_6t
Xbit_r179_c218 bl[218] br[218] wl[179] vdd gnd cell_6t
Xbit_r180_c218 bl[218] br[218] wl[180] vdd gnd cell_6t
Xbit_r181_c218 bl[218] br[218] wl[181] vdd gnd cell_6t
Xbit_r182_c218 bl[218] br[218] wl[182] vdd gnd cell_6t
Xbit_r183_c218 bl[218] br[218] wl[183] vdd gnd cell_6t
Xbit_r184_c218 bl[218] br[218] wl[184] vdd gnd cell_6t
Xbit_r185_c218 bl[218] br[218] wl[185] vdd gnd cell_6t
Xbit_r186_c218 bl[218] br[218] wl[186] vdd gnd cell_6t
Xbit_r187_c218 bl[218] br[218] wl[187] vdd gnd cell_6t
Xbit_r188_c218 bl[218] br[218] wl[188] vdd gnd cell_6t
Xbit_r189_c218 bl[218] br[218] wl[189] vdd gnd cell_6t
Xbit_r190_c218 bl[218] br[218] wl[190] vdd gnd cell_6t
Xbit_r191_c218 bl[218] br[218] wl[191] vdd gnd cell_6t
Xbit_r192_c218 bl[218] br[218] wl[192] vdd gnd cell_6t
Xbit_r193_c218 bl[218] br[218] wl[193] vdd gnd cell_6t
Xbit_r194_c218 bl[218] br[218] wl[194] vdd gnd cell_6t
Xbit_r195_c218 bl[218] br[218] wl[195] vdd gnd cell_6t
Xbit_r196_c218 bl[218] br[218] wl[196] vdd gnd cell_6t
Xbit_r197_c218 bl[218] br[218] wl[197] vdd gnd cell_6t
Xbit_r198_c218 bl[218] br[218] wl[198] vdd gnd cell_6t
Xbit_r199_c218 bl[218] br[218] wl[199] vdd gnd cell_6t
Xbit_r200_c218 bl[218] br[218] wl[200] vdd gnd cell_6t
Xbit_r201_c218 bl[218] br[218] wl[201] vdd gnd cell_6t
Xbit_r202_c218 bl[218] br[218] wl[202] vdd gnd cell_6t
Xbit_r203_c218 bl[218] br[218] wl[203] vdd gnd cell_6t
Xbit_r204_c218 bl[218] br[218] wl[204] vdd gnd cell_6t
Xbit_r205_c218 bl[218] br[218] wl[205] vdd gnd cell_6t
Xbit_r206_c218 bl[218] br[218] wl[206] vdd gnd cell_6t
Xbit_r207_c218 bl[218] br[218] wl[207] vdd gnd cell_6t
Xbit_r208_c218 bl[218] br[218] wl[208] vdd gnd cell_6t
Xbit_r209_c218 bl[218] br[218] wl[209] vdd gnd cell_6t
Xbit_r210_c218 bl[218] br[218] wl[210] vdd gnd cell_6t
Xbit_r211_c218 bl[218] br[218] wl[211] vdd gnd cell_6t
Xbit_r212_c218 bl[218] br[218] wl[212] vdd gnd cell_6t
Xbit_r213_c218 bl[218] br[218] wl[213] vdd gnd cell_6t
Xbit_r214_c218 bl[218] br[218] wl[214] vdd gnd cell_6t
Xbit_r215_c218 bl[218] br[218] wl[215] vdd gnd cell_6t
Xbit_r216_c218 bl[218] br[218] wl[216] vdd gnd cell_6t
Xbit_r217_c218 bl[218] br[218] wl[217] vdd gnd cell_6t
Xbit_r218_c218 bl[218] br[218] wl[218] vdd gnd cell_6t
Xbit_r219_c218 bl[218] br[218] wl[219] vdd gnd cell_6t
Xbit_r220_c218 bl[218] br[218] wl[220] vdd gnd cell_6t
Xbit_r221_c218 bl[218] br[218] wl[221] vdd gnd cell_6t
Xbit_r222_c218 bl[218] br[218] wl[222] vdd gnd cell_6t
Xbit_r223_c218 bl[218] br[218] wl[223] vdd gnd cell_6t
Xbit_r224_c218 bl[218] br[218] wl[224] vdd gnd cell_6t
Xbit_r225_c218 bl[218] br[218] wl[225] vdd gnd cell_6t
Xbit_r226_c218 bl[218] br[218] wl[226] vdd gnd cell_6t
Xbit_r227_c218 bl[218] br[218] wl[227] vdd gnd cell_6t
Xbit_r228_c218 bl[218] br[218] wl[228] vdd gnd cell_6t
Xbit_r229_c218 bl[218] br[218] wl[229] vdd gnd cell_6t
Xbit_r230_c218 bl[218] br[218] wl[230] vdd gnd cell_6t
Xbit_r231_c218 bl[218] br[218] wl[231] vdd gnd cell_6t
Xbit_r232_c218 bl[218] br[218] wl[232] vdd gnd cell_6t
Xbit_r233_c218 bl[218] br[218] wl[233] vdd gnd cell_6t
Xbit_r234_c218 bl[218] br[218] wl[234] vdd gnd cell_6t
Xbit_r235_c218 bl[218] br[218] wl[235] vdd gnd cell_6t
Xbit_r236_c218 bl[218] br[218] wl[236] vdd gnd cell_6t
Xbit_r237_c218 bl[218] br[218] wl[237] vdd gnd cell_6t
Xbit_r238_c218 bl[218] br[218] wl[238] vdd gnd cell_6t
Xbit_r239_c218 bl[218] br[218] wl[239] vdd gnd cell_6t
Xbit_r240_c218 bl[218] br[218] wl[240] vdd gnd cell_6t
Xbit_r241_c218 bl[218] br[218] wl[241] vdd gnd cell_6t
Xbit_r242_c218 bl[218] br[218] wl[242] vdd gnd cell_6t
Xbit_r243_c218 bl[218] br[218] wl[243] vdd gnd cell_6t
Xbit_r244_c218 bl[218] br[218] wl[244] vdd gnd cell_6t
Xbit_r245_c218 bl[218] br[218] wl[245] vdd gnd cell_6t
Xbit_r246_c218 bl[218] br[218] wl[246] vdd gnd cell_6t
Xbit_r247_c218 bl[218] br[218] wl[247] vdd gnd cell_6t
Xbit_r248_c218 bl[218] br[218] wl[248] vdd gnd cell_6t
Xbit_r249_c218 bl[218] br[218] wl[249] vdd gnd cell_6t
Xbit_r250_c218 bl[218] br[218] wl[250] vdd gnd cell_6t
Xbit_r251_c218 bl[218] br[218] wl[251] vdd gnd cell_6t
Xbit_r252_c218 bl[218] br[218] wl[252] vdd gnd cell_6t
Xbit_r253_c218 bl[218] br[218] wl[253] vdd gnd cell_6t
Xbit_r254_c218 bl[218] br[218] wl[254] vdd gnd cell_6t
Xbit_r255_c218 bl[218] br[218] wl[255] vdd gnd cell_6t
Xbit_r0_c219 bl[219] br[219] wl[0] vdd gnd cell_6t
Xbit_r1_c219 bl[219] br[219] wl[1] vdd gnd cell_6t
Xbit_r2_c219 bl[219] br[219] wl[2] vdd gnd cell_6t
Xbit_r3_c219 bl[219] br[219] wl[3] vdd gnd cell_6t
Xbit_r4_c219 bl[219] br[219] wl[4] vdd gnd cell_6t
Xbit_r5_c219 bl[219] br[219] wl[5] vdd gnd cell_6t
Xbit_r6_c219 bl[219] br[219] wl[6] vdd gnd cell_6t
Xbit_r7_c219 bl[219] br[219] wl[7] vdd gnd cell_6t
Xbit_r8_c219 bl[219] br[219] wl[8] vdd gnd cell_6t
Xbit_r9_c219 bl[219] br[219] wl[9] vdd gnd cell_6t
Xbit_r10_c219 bl[219] br[219] wl[10] vdd gnd cell_6t
Xbit_r11_c219 bl[219] br[219] wl[11] vdd gnd cell_6t
Xbit_r12_c219 bl[219] br[219] wl[12] vdd gnd cell_6t
Xbit_r13_c219 bl[219] br[219] wl[13] vdd gnd cell_6t
Xbit_r14_c219 bl[219] br[219] wl[14] vdd gnd cell_6t
Xbit_r15_c219 bl[219] br[219] wl[15] vdd gnd cell_6t
Xbit_r16_c219 bl[219] br[219] wl[16] vdd gnd cell_6t
Xbit_r17_c219 bl[219] br[219] wl[17] vdd gnd cell_6t
Xbit_r18_c219 bl[219] br[219] wl[18] vdd gnd cell_6t
Xbit_r19_c219 bl[219] br[219] wl[19] vdd gnd cell_6t
Xbit_r20_c219 bl[219] br[219] wl[20] vdd gnd cell_6t
Xbit_r21_c219 bl[219] br[219] wl[21] vdd gnd cell_6t
Xbit_r22_c219 bl[219] br[219] wl[22] vdd gnd cell_6t
Xbit_r23_c219 bl[219] br[219] wl[23] vdd gnd cell_6t
Xbit_r24_c219 bl[219] br[219] wl[24] vdd gnd cell_6t
Xbit_r25_c219 bl[219] br[219] wl[25] vdd gnd cell_6t
Xbit_r26_c219 bl[219] br[219] wl[26] vdd gnd cell_6t
Xbit_r27_c219 bl[219] br[219] wl[27] vdd gnd cell_6t
Xbit_r28_c219 bl[219] br[219] wl[28] vdd gnd cell_6t
Xbit_r29_c219 bl[219] br[219] wl[29] vdd gnd cell_6t
Xbit_r30_c219 bl[219] br[219] wl[30] vdd gnd cell_6t
Xbit_r31_c219 bl[219] br[219] wl[31] vdd gnd cell_6t
Xbit_r32_c219 bl[219] br[219] wl[32] vdd gnd cell_6t
Xbit_r33_c219 bl[219] br[219] wl[33] vdd gnd cell_6t
Xbit_r34_c219 bl[219] br[219] wl[34] vdd gnd cell_6t
Xbit_r35_c219 bl[219] br[219] wl[35] vdd gnd cell_6t
Xbit_r36_c219 bl[219] br[219] wl[36] vdd gnd cell_6t
Xbit_r37_c219 bl[219] br[219] wl[37] vdd gnd cell_6t
Xbit_r38_c219 bl[219] br[219] wl[38] vdd gnd cell_6t
Xbit_r39_c219 bl[219] br[219] wl[39] vdd gnd cell_6t
Xbit_r40_c219 bl[219] br[219] wl[40] vdd gnd cell_6t
Xbit_r41_c219 bl[219] br[219] wl[41] vdd gnd cell_6t
Xbit_r42_c219 bl[219] br[219] wl[42] vdd gnd cell_6t
Xbit_r43_c219 bl[219] br[219] wl[43] vdd gnd cell_6t
Xbit_r44_c219 bl[219] br[219] wl[44] vdd gnd cell_6t
Xbit_r45_c219 bl[219] br[219] wl[45] vdd gnd cell_6t
Xbit_r46_c219 bl[219] br[219] wl[46] vdd gnd cell_6t
Xbit_r47_c219 bl[219] br[219] wl[47] vdd gnd cell_6t
Xbit_r48_c219 bl[219] br[219] wl[48] vdd gnd cell_6t
Xbit_r49_c219 bl[219] br[219] wl[49] vdd gnd cell_6t
Xbit_r50_c219 bl[219] br[219] wl[50] vdd gnd cell_6t
Xbit_r51_c219 bl[219] br[219] wl[51] vdd gnd cell_6t
Xbit_r52_c219 bl[219] br[219] wl[52] vdd gnd cell_6t
Xbit_r53_c219 bl[219] br[219] wl[53] vdd gnd cell_6t
Xbit_r54_c219 bl[219] br[219] wl[54] vdd gnd cell_6t
Xbit_r55_c219 bl[219] br[219] wl[55] vdd gnd cell_6t
Xbit_r56_c219 bl[219] br[219] wl[56] vdd gnd cell_6t
Xbit_r57_c219 bl[219] br[219] wl[57] vdd gnd cell_6t
Xbit_r58_c219 bl[219] br[219] wl[58] vdd gnd cell_6t
Xbit_r59_c219 bl[219] br[219] wl[59] vdd gnd cell_6t
Xbit_r60_c219 bl[219] br[219] wl[60] vdd gnd cell_6t
Xbit_r61_c219 bl[219] br[219] wl[61] vdd gnd cell_6t
Xbit_r62_c219 bl[219] br[219] wl[62] vdd gnd cell_6t
Xbit_r63_c219 bl[219] br[219] wl[63] vdd gnd cell_6t
Xbit_r64_c219 bl[219] br[219] wl[64] vdd gnd cell_6t
Xbit_r65_c219 bl[219] br[219] wl[65] vdd gnd cell_6t
Xbit_r66_c219 bl[219] br[219] wl[66] vdd gnd cell_6t
Xbit_r67_c219 bl[219] br[219] wl[67] vdd gnd cell_6t
Xbit_r68_c219 bl[219] br[219] wl[68] vdd gnd cell_6t
Xbit_r69_c219 bl[219] br[219] wl[69] vdd gnd cell_6t
Xbit_r70_c219 bl[219] br[219] wl[70] vdd gnd cell_6t
Xbit_r71_c219 bl[219] br[219] wl[71] vdd gnd cell_6t
Xbit_r72_c219 bl[219] br[219] wl[72] vdd gnd cell_6t
Xbit_r73_c219 bl[219] br[219] wl[73] vdd gnd cell_6t
Xbit_r74_c219 bl[219] br[219] wl[74] vdd gnd cell_6t
Xbit_r75_c219 bl[219] br[219] wl[75] vdd gnd cell_6t
Xbit_r76_c219 bl[219] br[219] wl[76] vdd gnd cell_6t
Xbit_r77_c219 bl[219] br[219] wl[77] vdd gnd cell_6t
Xbit_r78_c219 bl[219] br[219] wl[78] vdd gnd cell_6t
Xbit_r79_c219 bl[219] br[219] wl[79] vdd gnd cell_6t
Xbit_r80_c219 bl[219] br[219] wl[80] vdd gnd cell_6t
Xbit_r81_c219 bl[219] br[219] wl[81] vdd gnd cell_6t
Xbit_r82_c219 bl[219] br[219] wl[82] vdd gnd cell_6t
Xbit_r83_c219 bl[219] br[219] wl[83] vdd gnd cell_6t
Xbit_r84_c219 bl[219] br[219] wl[84] vdd gnd cell_6t
Xbit_r85_c219 bl[219] br[219] wl[85] vdd gnd cell_6t
Xbit_r86_c219 bl[219] br[219] wl[86] vdd gnd cell_6t
Xbit_r87_c219 bl[219] br[219] wl[87] vdd gnd cell_6t
Xbit_r88_c219 bl[219] br[219] wl[88] vdd gnd cell_6t
Xbit_r89_c219 bl[219] br[219] wl[89] vdd gnd cell_6t
Xbit_r90_c219 bl[219] br[219] wl[90] vdd gnd cell_6t
Xbit_r91_c219 bl[219] br[219] wl[91] vdd gnd cell_6t
Xbit_r92_c219 bl[219] br[219] wl[92] vdd gnd cell_6t
Xbit_r93_c219 bl[219] br[219] wl[93] vdd gnd cell_6t
Xbit_r94_c219 bl[219] br[219] wl[94] vdd gnd cell_6t
Xbit_r95_c219 bl[219] br[219] wl[95] vdd gnd cell_6t
Xbit_r96_c219 bl[219] br[219] wl[96] vdd gnd cell_6t
Xbit_r97_c219 bl[219] br[219] wl[97] vdd gnd cell_6t
Xbit_r98_c219 bl[219] br[219] wl[98] vdd gnd cell_6t
Xbit_r99_c219 bl[219] br[219] wl[99] vdd gnd cell_6t
Xbit_r100_c219 bl[219] br[219] wl[100] vdd gnd cell_6t
Xbit_r101_c219 bl[219] br[219] wl[101] vdd gnd cell_6t
Xbit_r102_c219 bl[219] br[219] wl[102] vdd gnd cell_6t
Xbit_r103_c219 bl[219] br[219] wl[103] vdd gnd cell_6t
Xbit_r104_c219 bl[219] br[219] wl[104] vdd gnd cell_6t
Xbit_r105_c219 bl[219] br[219] wl[105] vdd gnd cell_6t
Xbit_r106_c219 bl[219] br[219] wl[106] vdd gnd cell_6t
Xbit_r107_c219 bl[219] br[219] wl[107] vdd gnd cell_6t
Xbit_r108_c219 bl[219] br[219] wl[108] vdd gnd cell_6t
Xbit_r109_c219 bl[219] br[219] wl[109] vdd gnd cell_6t
Xbit_r110_c219 bl[219] br[219] wl[110] vdd gnd cell_6t
Xbit_r111_c219 bl[219] br[219] wl[111] vdd gnd cell_6t
Xbit_r112_c219 bl[219] br[219] wl[112] vdd gnd cell_6t
Xbit_r113_c219 bl[219] br[219] wl[113] vdd gnd cell_6t
Xbit_r114_c219 bl[219] br[219] wl[114] vdd gnd cell_6t
Xbit_r115_c219 bl[219] br[219] wl[115] vdd gnd cell_6t
Xbit_r116_c219 bl[219] br[219] wl[116] vdd gnd cell_6t
Xbit_r117_c219 bl[219] br[219] wl[117] vdd gnd cell_6t
Xbit_r118_c219 bl[219] br[219] wl[118] vdd gnd cell_6t
Xbit_r119_c219 bl[219] br[219] wl[119] vdd gnd cell_6t
Xbit_r120_c219 bl[219] br[219] wl[120] vdd gnd cell_6t
Xbit_r121_c219 bl[219] br[219] wl[121] vdd gnd cell_6t
Xbit_r122_c219 bl[219] br[219] wl[122] vdd gnd cell_6t
Xbit_r123_c219 bl[219] br[219] wl[123] vdd gnd cell_6t
Xbit_r124_c219 bl[219] br[219] wl[124] vdd gnd cell_6t
Xbit_r125_c219 bl[219] br[219] wl[125] vdd gnd cell_6t
Xbit_r126_c219 bl[219] br[219] wl[126] vdd gnd cell_6t
Xbit_r127_c219 bl[219] br[219] wl[127] vdd gnd cell_6t
Xbit_r128_c219 bl[219] br[219] wl[128] vdd gnd cell_6t
Xbit_r129_c219 bl[219] br[219] wl[129] vdd gnd cell_6t
Xbit_r130_c219 bl[219] br[219] wl[130] vdd gnd cell_6t
Xbit_r131_c219 bl[219] br[219] wl[131] vdd gnd cell_6t
Xbit_r132_c219 bl[219] br[219] wl[132] vdd gnd cell_6t
Xbit_r133_c219 bl[219] br[219] wl[133] vdd gnd cell_6t
Xbit_r134_c219 bl[219] br[219] wl[134] vdd gnd cell_6t
Xbit_r135_c219 bl[219] br[219] wl[135] vdd gnd cell_6t
Xbit_r136_c219 bl[219] br[219] wl[136] vdd gnd cell_6t
Xbit_r137_c219 bl[219] br[219] wl[137] vdd gnd cell_6t
Xbit_r138_c219 bl[219] br[219] wl[138] vdd gnd cell_6t
Xbit_r139_c219 bl[219] br[219] wl[139] vdd gnd cell_6t
Xbit_r140_c219 bl[219] br[219] wl[140] vdd gnd cell_6t
Xbit_r141_c219 bl[219] br[219] wl[141] vdd gnd cell_6t
Xbit_r142_c219 bl[219] br[219] wl[142] vdd gnd cell_6t
Xbit_r143_c219 bl[219] br[219] wl[143] vdd gnd cell_6t
Xbit_r144_c219 bl[219] br[219] wl[144] vdd gnd cell_6t
Xbit_r145_c219 bl[219] br[219] wl[145] vdd gnd cell_6t
Xbit_r146_c219 bl[219] br[219] wl[146] vdd gnd cell_6t
Xbit_r147_c219 bl[219] br[219] wl[147] vdd gnd cell_6t
Xbit_r148_c219 bl[219] br[219] wl[148] vdd gnd cell_6t
Xbit_r149_c219 bl[219] br[219] wl[149] vdd gnd cell_6t
Xbit_r150_c219 bl[219] br[219] wl[150] vdd gnd cell_6t
Xbit_r151_c219 bl[219] br[219] wl[151] vdd gnd cell_6t
Xbit_r152_c219 bl[219] br[219] wl[152] vdd gnd cell_6t
Xbit_r153_c219 bl[219] br[219] wl[153] vdd gnd cell_6t
Xbit_r154_c219 bl[219] br[219] wl[154] vdd gnd cell_6t
Xbit_r155_c219 bl[219] br[219] wl[155] vdd gnd cell_6t
Xbit_r156_c219 bl[219] br[219] wl[156] vdd gnd cell_6t
Xbit_r157_c219 bl[219] br[219] wl[157] vdd gnd cell_6t
Xbit_r158_c219 bl[219] br[219] wl[158] vdd gnd cell_6t
Xbit_r159_c219 bl[219] br[219] wl[159] vdd gnd cell_6t
Xbit_r160_c219 bl[219] br[219] wl[160] vdd gnd cell_6t
Xbit_r161_c219 bl[219] br[219] wl[161] vdd gnd cell_6t
Xbit_r162_c219 bl[219] br[219] wl[162] vdd gnd cell_6t
Xbit_r163_c219 bl[219] br[219] wl[163] vdd gnd cell_6t
Xbit_r164_c219 bl[219] br[219] wl[164] vdd gnd cell_6t
Xbit_r165_c219 bl[219] br[219] wl[165] vdd gnd cell_6t
Xbit_r166_c219 bl[219] br[219] wl[166] vdd gnd cell_6t
Xbit_r167_c219 bl[219] br[219] wl[167] vdd gnd cell_6t
Xbit_r168_c219 bl[219] br[219] wl[168] vdd gnd cell_6t
Xbit_r169_c219 bl[219] br[219] wl[169] vdd gnd cell_6t
Xbit_r170_c219 bl[219] br[219] wl[170] vdd gnd cell_6t
Xbit_r171_c219 bl[219] br[219] wl[171] vdd gnd cell_6t
Xbit_r172_c219 bl[219] br[219] wl[172] vdd gnd cell_6t
Xbit_r173_c219 bl[219] br[219] wl[173] vdd gnd cell_6t
Xbit_r174_c219 bl[219] br[219] wl[174] vdd gnd cell_6t
Xbit_r175_c219 bl[219] br[219] wl[175] vdd gnd cell_6t
Xbit_r176_c219 bl[219] br[219] wl[176] vdd gnd cell_6t
Xbit_r177_c219 bl[219] br[219] wl[177] vdd gnd cell_6t
Xbit_r178_c219 bl[219] br[219] wl[178] vdd gnd cell_6t
Xbit_r179_c219 bl[219] br[219] wl[179] vdd gnd cell_6t
Xbit_r180_c219 bl[219] br[219] wl[180] vdd gnd cell_6t
Xbit_r181_c219 bl[219] br[219] wl[181] vdd gnd cell_6t
Xbit_r182_c219 bl[219] br[219] wl[182] vdd gnd cell_6t
Xbit_r183_c219 bl[219] br[219] wl[183] vdd gnd cell_6t
Xbit_r184_c219 bl[219] br[219] wl[184] vdd gnd cell_6t
Xbit_r185_c219 bl[219] br[219] wl[185] vdd gnd cell_6t
Xbit_r186_c219 bl[219] br[219] wl[186] vdd gnd cell_6t
Xbit_r187_c219 bl[219] br[219] wl[187] vdd gnd cell_6t
Xbit_r188_c219 bl[219] br[219] wl[188] vdd gnd cell_6t
Xbit_r189_c219 bl[219] br[219] wl[189] vdd gnd cell_6t
Xbit_r190_c219 bl[219] br[219] wl[190] vdd gnd cell_6t
Xbit_r191_c219 bl[219] br[219] wl[191] vdd gnd cell_6t
Xbit_r192_c219 bl[219] br[219] wl[192] vdd gnd cell_6t
Xbit_r193_c219 bl[219] br[219] wl[193] vdd gnd cell_6t
Xbit_r194_c219 bl[219] br[219] wl[194] vdd gnd cell_6t
Xbit_r195_c219 bl[219] br[219] wl[195] vdd gnd cell_6t
Xbit_r196_c219 bl[219] br[219] wl[196] vdd gnd cell_6t
Xbit_r197_c219 bl[219] br[219] wl[197] vdd gnd cell_6t
Xbit_r198_c219 bl[219] br[219] wl[198] vdd gnd cell_6t
Xbit_r199_c219 bl[219] br[219] wl[199] vdd gnd cell_6t
Xbit_r200_c219 bl[219] br[219] wl[200] vdd gnd cell_6t
Xbit_r201_c219 bl[219] br[219] wl[201] vdd gnd cell_6t
Xbit_r202_c219 bl[219] br[219] wl[202] vdd gnd cell_6t
Xbit_r203_c219 bl[219] br[219] wl[203] vdd gnd cell_6t
Xbit_r204_c219 bl[219] br[219] wl[204] vdd gnd cell_6t
Xbit_r205_c219 bl[219] br[219] wl[205] vdd gnd cell_6t
Xbit_r206_c219 bl[219] br[219] wl[206] vdd gnd cell_6t
Xbit_r207_c219 bl[219] br[219] wl[207] vdd gnd cell_6t
Xbit_r208_c219 bl[219] br[219] wl[208] vdd gnd cell_6t
Xbit_r209_c219 bl[219] br[219] wl[209] vdd gnd cell_6t
Xbit_r210_c219 bl[219] br[219] wl[210] vdd gnd cell_6t
Xbit_r211_c219 bl[219] br[219] wl[211] vdd gnd cell_6t
Xbit_r212_c219 bl[219] br[219] wl[212] vdd gnd cell_6t
Xbit_r213_c219 bl[219] br[219] wl[213] vdd gnd cell_6t
Xbit_r214_c219 bl[219] br[219] wl[214] vdd gnd cell_6t
Xbit_r215_c219 bl[219] br[219] wl[215] vdd gnd cell_6t
Xbit_r216_c219 bl[219] br[219] wl[216] vdd gnd cell_6t
Xbit_r217_c219 bl[219] br[219] wl[217] vdd gnd cell_6t
Xbit_r218_c219 bl[219] br[219] wl[218] vdd gnd cell_6t
Xbit_r219_c219 bl[219] br[219] wl[219] vdd gnd cell_6t
Xbit_r220_c219 bl[219] br[219] wl[220] vdd gnd cell_6t
Xbit_r221_c219 bl[219] br[219] wl[221] vdd gnd cell_6t
Xbit_r222_c219 bl[219] br[219] wl[222] vdd gnd cell_6t
Xbit_r223_c219 bl[219] br[219] wl[223] vdd gnd cell_6t
Xbit_r224_c219 bl[219] br[219] wl[224] vdd gnd cell_6t
Xbit_r225_c219 bl[219] br[219] wl[225] vdd gnd cell_6t
Xbit_r226_c219 bl[219] br[219] wl[226] vdd gnd cell_6t
Xbit_r227_c219 bl[219] br[219] wl[227] vdd gnd cell_6t
Xbit_r228_c219 bl[219] br[219] wl[228] vdd gnd cell_6t
Xbit_r229_c219 bl[219] br[219] wl[229] vdd gnd cell_6t
Xbit_r230_c219 bl[219] br[219] wl[230] vdd gnd cell_6t
Xbit_r231_c219 bl[219] br[219] wl[231] vdd gnd cell_6t
Xbit_r232_c219 bl[219] br[219] wl[232] vdd gnd cell_6t
Xbit_r233_c219 bl[219] br[219] wl[233] vdd gnd cell_6t
Xbit_r234_c219 bl[219] br[219] wl[234] vdd gnd cell_6t
Xbit_r235_c219 bl[219] br[219] wl[235] vdd gnd cell_6t
Xbit_r236_c219 bl[219] br[219] wl[236] vdd gnd cell_6t
Xbit_r237_c219 bl[219] br[219] wl[237] vdd gnd cell_6t
Xbit_r238_c219 bl[219] br[219] wl[238] vdd gnd cell_6t
Xbit_r239_c219 bl[219] br[219] wl[239] vdd gnd cell_6t
Xbit_r240_c219 bl[219] br[219] wl[240] vdd gnd cell_6t
Xbit_r241_c219 bl[219] br[219] wl[241] vdd gnd cell_6t
Xbit_r242_c219 bl[219] br[219] wl[242] vdd gnd cell_6t
Xbit_r243_c219 bl[219] br[219] wl[243] vdd gnd cell_6t
Xbit_r244_c219 bl[219] br[219] wl[244] vdd gnd cell_6t
Xbit_r245_c219 bl[219] br[219] wl[245] vdd gnd cell_6t
Xbit_r246_c219 bl[219] br[219] wl[246] vdd gnd cell_6t
Xbit_r247_c219 bl[219] br[219] wl[247] vdd gnd cell_6t
Xbit_r248_c219 bl[219] br[219] wl[248] vdd gnd cell_6t
Xbit_r249_c219 bl[219] br[219] wl[249] vdd gnd cell_6t
Xbit_r250_c219 bl[219] br[219] wl[250] vdd gnd cell_6t
Xbit_r251_c219 bl[219] br[219] wl[251] vdd gnd cell_6t
Xbit_r252_c219 bl[219] br[219] wl[252] vdd gnd cell_6t
Xbit_r253_c219 bl[219] br[219] wl[253] vdd gnd cell_6t
Xbit_r254_c219 bl[219] br[219] wl[254] vdd gnd cell_6t
Xbit_r255_c219 bl[219] br[219] wl[255] vdd gnd cell_6t
Xbit_r0_c220 bl[220] br[220] wl[0] vdd gnd cell_6t
Xbit_r1_c220 bl[220] br[220] wl[1] vdd gnd cell_6t
Xbit_r2_c220 bl[220] br[220] wl[2] vdd gnd cell_6t
Xbit_r3_c220 bl[220] br[220] wl[3] vdd gnd cell_6t
Xbit_r4_c220 bl[220] br[220] wl[4] vdd gnd cell_6t
Xbit_r5_c220 bl[220] br[220] wl[5] vdd gnd cell_6t
Xbit_r6_c220 bl[220] br[220] wl[6] vdd gnd cell_6t
Xbit_r7_c220 bl[220] br[220] wl[7] vdd gnd cell_6t
Xbit_r8_c220 bl[220] br[220] wl[8] vdd gnd cell_6t
Xbit_r9_c220 bl[220] br[220] wl[9] vdd gnd cell_6t
Xbit_r10_c220 bl[220] br[220] wl[10] vdd gnd cell_6t
Xbit_r11_c220 bl[220] br[220] wl[11] vdd gnd cell_6t
Xbit_r12_c220 bl[220] br[220] wl[12] vdd gnd cell_6t
Xbit_r13_c220 bl[220] br[220] wl[13] vdd gnd cell_6t
Xbit_r14_c220 bl[220] br[220] wl[14] vdd gnd cell_6t
Xbit_r15_c220 bl[220] br[220] wl[15] vdd gnd cell_6t
Xbit_r16_c220 bl[220] br[220] wl[16] vdd gnd cell_6t
Xbit_r17_c220 bl[220] br[220] wl[17] vdd gnd cell_6t
Xbit_r18_c220 bl[220] br[220] wl[18] vdd gnd cell_6t
Xbit_r19_c220 bl[220] br[220] wl[19] vdd gnd cell_6t
Xbit_r20_c220 bl[220] br[220] wl[20] vdd gnd cell_6t
Xbit_r21_c220 bl[220] br[220] wl[21] vdd gnd cell_6t
Xbit_r22_c220 bl[220] br[220] wl[22] vdd gnd cell_6t
Xbit_r23_c220 bl[220] br[220] wl[23] vdd gnd cell_6t
Xbit_r24_c220 bl[220] br[220] wl[24] vdd gnd cell_6t
Xbit_r25_c220 bl[220] br[220] wl[25] vdd gnd cell_6t
Xbit_r26_c220 bl[220] br[220] wl[26] vdd gnd cell_6t
Xbit_r27_c220 bl[220] br[220] wl[27] vdd gnd cell_6t
Xbit_r28_c220 bl[220] br[220] wl[28] vdd gnd cell_6t
Xbit_r29_c220 bl[220] br[220] wl[29] vdd gnd cell_6t
Xbit_r30_c220 bl[220] br[220] wl[30] vdd gnd cell_6t
Xbit_r31_c220 bl[220] br[220] wl[31] vdd gnd cell_6t
Xbit_r32_c220 bl[220] br[220] wl[32] vdd gnd cell_6t
Xbit_r33_c220 bl[220] br[220] wl[33] vdd gnd cell_6t
Xbit_r34_c220 bl[220] br[220] wl[34] vdd gnd cell_6t
Xbit_r35_c220 bl[220] br[220] wl[35] vdd gnd cell_6t
Xbit_r36_c220 bl[220] br[220] wl[36] vdd gnd cell_6t
Xbit_r37_c220 bl[220] br[220] wl[37] vdd gnd cell_6t
Xbit_r38_c220 bl[220] br[220] wl[38] vdd gnd cell_6t
Xbit_r39_c220 bl[220] br[220] wl[39] vdd gnd cell_6t
Xbit_r40_c220 bl[220] br[220] wl[40] vdd gnd cell_6t
Xbit_r41_c220 bl[220] br[220] wl[41] vdd gnd cell_6t
Xbit_r42_c220 bl[220] br[220] wl[42] vdd gnd cell_6t
Xbit_r43_c220 bl[220] br[220] wl[43] vdd gnd cell_6t
Xbit_r44_c220 bl[220] br[220] wl[44] vdd gnd cell_6t
Xbit_r45_c220 bl[220] br[220] wl[45] vdd gnd cell_6t
Xbit_r46_c220 bl[220] br[220] wl[46] vdd gnd cell_6t
Xbit_r47_c220 bl[220] br[220] wl[47] vdd gnd cell_6t
Xbit_r48_c220 bl[220] br[220] wl[48] vdd gnd cell_6t
Xbit_r49_c220 bl[220] br[220] wl[49] vdd gnd cell_6t
Xbit_r50_c220 bl[220] br[220] wl[50] vdd gnd cell_6t
Xbit_r51_c220 bl[220] br[220] wl[51] vdd gnd cell_6t
Xbit_r52_c220 bl[220] br[220] wl[52] vdd gnd cell_6t
Xbit_r53_c220 bl[220] br[220] wl[53] vdd gnd cell_6t
Xbit_r54_c220 bl[220] br[220] wl[54] vdd gnd cell_6t
Xbit_r55_c220 bl[220] br[220] wl[55] vdd gnd cell_6t
Xbit_r56_c220 bl[220] br[220] wl[56] vdd gnd cell_6t
Xbit_r57_c220 bl[220] br[220] wl[57] vdd gnd cell_6t
Xbit_r58_c220 bl[220] br[220] wl[58] vdd gnd cell_6t
Xbit_r59_c220 bl[220] br[220] wl[59] vdd gnd cell_6t
Xbit_r60_c220 bl[220] br[220] wl[60] vdd gnd cell_6t
Xbit_r61_c220 bl[220] br[220] wl[61] vdd gnd cell_6t
Xbit_r62_c220 bl[220] br[220] wl[62] vdd gnd cell_6t
Xbit_r63_c220 bl[220] br[220] wl[63] vdd gnd cell_6t
Xbit_r64_c220 bl[220] br[220] wl[64] vdd gnd cell_6t
Xbit_r65_c220 bl[220] br[220] wl[65] vdd gnd cell_6t
Xbit_r66_c220 bl[220] br[220] wl[66] vdd gnd cell_6t
Xbit_r67_c220 bl[220] br[220] wl[67] vdd gnd cell_6t
Xbit_r68_c220 bl[220] br[220] wl[68] vdd gnd cell_6t
Xbit_r69_c220 bl[220] br[220] wl[69] vdd gnd cell_6t
Xbit_r70_c220 bl[220] br[220] wl[70] vdd gnd cell_6t
Xbit_r71_c220 bl[220] br[220] wl[71] vdd gnd cell_6t
Xbit_r72_c220 bl[220] br[220] wl[72] vdd gnd cell_6t
Xbit_r73_c220 bl[220] br[220] wl[73] vdd gnd cell_6t
Xbit_r74_c220 bl[220] br[220] wl[74] vdd gnd cell_6t
Xbit_r75_c220 bl[220] br[220] wl[75] vdd gnd cell_6t
Xbit_r76_c220 bl[220] br[220] wl[76] vdd gnd cell_6t
Xbit_r77_c220 bl[220] br[220] wl[77] vdd gnd cell_6t
Xbit_r78_c220 bl[220] br[220] wl[78] vdd gnd cell_6t
Xbit_r79_c220 bl[220] br[220] wl[79] vdd gnd cell_6t
Xbit_r80_c220 bl[220] br[220] wl[80] vdd gnd cell_6t
Xbit_r81_c220 bl[220] br[220] wl[81] vdd gnd cell_6t
Xbit_r82_c220 bl[220] br[220] wl[82] vdd gnd cell_6t
Xbit_r83_c220 bl[220] br[220] wl[83] vdd gnd cell_6t
Xbit_r84_c220 bl[220] br[220] wl[84] vdd gnd cell_6t
Xbit_r85_c220 bl[220] br[220] wl[85] vdd gnd cell_6t
Xbit_r86_c220 bl[220] br[220] wl[86] vdd gnd cell_6t
Xbit_r87_c220 bl[220] br[220] wl[87] vdd gnd cell_6t
Xbit_r88_c220 bl[220] br[220] wl[88] vdd gnd cell_6t
Xbit_r89_c220 bl[220] br[220] wl[89] vdd gnd cell_6t
Xbit_r90_c220 bl[220] br[220] wl[90] vdd gnd cell_6t
Xbit_r91_c220 bl[220] br[220] wl[91] vdd gnd cell_6t
Xbit_r92_c220 bl[220] br[220] wl[92] vdd gnd cell_6t
Xbit_r93_c220 bl[220] br[220] wl[93] vdd gnd cell_6t
Xbit_r94_c220 bl[220] br[220] wl[94] vdd gnd cell_6t
Xbit_r95_c220 bl[220] br[220] wl[95] vdd gnd cell_6t
Xbit_r96_c220 bl[220] br[220] wl[96] vdd gnd cell_6t
Xbit_r97_c220 bl[220] br[220] wl[97] vdd gnd cell_6t
Xbit_r98_c220 bl[220] br[220] wl[98] vdd gnd cell_6t
Xbit_r99_c220 bl[220] br[220] wl[99] vdd gnd cell_6t
Xbit_r100_c220 bl[220] br[220] wl[100] vdd gnd cell_6t
Xbit_r101_c220 bl[220] br[220] wl[101] vdd gnd cell_6t
Xbit_r102_c220 bl[220] br[220] wl[102] vdd gnd cell_6t
Xbit_r103_c220 bl[220] br[220] wl[103] vdd gnd cell_6t
Xbit_r104_c220 bl[220] br[220] wl[104] vdd gnd cell_6t
Xbit_r105_c220 bl[220] br[220] wl[105] vdd gnd cell_6t
Xbit_r106_c220 bl[220] br[220] wl[106] vdd gnd cell_6t
Xbit_r107_c220 bl[220] br[220] wl[107] vdd gnd cell_6t
Xbit_r108_c220 bl[220] br[220] wl[108] vdd gnd cell_6t
Xbit_r109_c220 bl[220] br[220] wl[109] vdd gnd cell_6t
Xbit_r110_c220 bl[220] br[220] wl[110] vdd gnd cell_6t
Xbit_r111_c220 bl[220] br[220] wl[111] vdd gnd cell_6t
Xbit_r112_c220 bl[220] br[220] wl[112] vdd gnd cell_6t
Xbit_r113_c220 bl[220] br[220] wl[113] vdd gnd cell_6t
Xbit_r114_c220 bl[220] br[220] wl[114] vdd gnd cell_6t
Xbit_r115_c220 bl[220] br[220] wl[115] vdd gnd cell_6t
Xbit_r116_c220 bl[220] br[220] wl[116] vdd gnd cell_6t
Xbit_r117_c220 bl[220] br[220] wl[117] vdd gnd cell_6t
Xbit_r118_c220 bl[220] br[220] wl[118] vdd gnd cell_6t
Xbit_r119_c220 bl[220] br[220] wl[119] vdd gnd cell_6t
Xbit_r120_c220 bl[220] br[220] wl[120] vdd gnd cell_6t
Xbit_r121_c220 bl[220] br[220] wl[121] vdd gnd cell_6t
Xbit_r122_c220 bl[220] br[220] wl[122] vdd gnd cell_6t
Xbit_r123_c220 bl[220] br[220] wl[123] vdd gnd cell_6t
Xbit_r124_c220 bl[220] br[220] wl[124] vdd gnd cell_6t
Xbit_r125_c220 bl[220] br[220] wl[125] vdd gnd cell_6t
Xbit_r126_c220 bl[220] br[220] wl[126] vdd gnd cell_6t
Xbit_r127_c220 bl[220] br[220] wl[127] vdd gnd cell_6t
Xbit_r128_c220 bl[220] br[220] wl[128] vdd gnd cell_6t
Xbit_r129_c220 bl[220] br[220] wl[129] vdd gnd cell_6t
Xbit_r130_c220 bl[220] br[220] wl[130] vdd gnd cell_6t
Xbit_r131_c220 bl[220] br[220] wl[131] vdd gnd cell_6t
Xbit_r132_c220 bl[220] br[220] wl[132] vdd gnd cell_6t
Xbit_r133_c220 bl[220] br[220] wl[133] vdd gnd cell_6t
Xbit_r134_c220 bl[220] br[220] wl[134] vdd gnd cell_6t
Xbit_r135_c220 bl[220] br[220] wl[135] vdd gnd cell_6t
Xbit_r136_c220 bl[220] br[220] wl[136] vdd gnd cell_6t
Xbit_r137_c220 bl[220] br[220] wl[137] vdd gnd cell_6t
Xbit_r138_c220 bl[220] br[220] wl[138] vdd gnd cell_6t
Xbit_r139_c220 bl[220] br[220] wl[139] vdd gnd cell_6t
Xbit_r140_c220 bl[220] br[220] wl[140] vdd gnd cell_6t
Xbit_r141_c220 bl[220] br[220] wl[141] vdd gnd cell_6t
Xbit_r142_c220 bl[220] br[220] wl[142] vdd gnd cell_6t
Xbit_r143_c220 bl[220] br[220] wl[143] vdd gnd cell_6t
Xbit_r144_c220 bl[220] br[220] wl[144] vdd gnd cell_6t
Xbit_r145_c220 bl[220] br[220] wl[145] vdd gnd cell_6t
Xbit_r146_c220 bl[220] br[220] wl[146] vdd gnd cell_6t
Xbit_r147_c220 bl[220] br[220] wl[147] vdd gnd cell_6t
Xbit_r148_c220 bl[220] br[220] wl[148] vdd gnd cell_6t
Xbit_r149_c220 bl[220] br[220] wl[149] vdd gnd cell_6t
Xbit_r150_c220 bl[220] br[220] wl[150] vdd gnd cell_6t
Xbit_r151_c220 bl[220] br[220] wl[151] vdd gnd cell_6t
Xbit_r152_c220 bl[220] br[220] wl[152] vdd gnd cell_6t
Xbit_r153_c220 bl[220] br[220] wl[153] vdd gnd cell_6t
Xbit_r154_c220 bl[220] br[220] wl[154] vdd gnd cell_6t
Xbit_r155_c220 bl[220] br[220] wl[155] vdd gnd cell_6t
Xbit_r156_c220 bl[220] br[220] wl[156] vdd gnd cell_6t
Xbit_r157_c220 bl[220] br[220] wl[157] vdd gnd cell_6t
Xbit_r158_c220 bl[220] br[220] wl[158] vdd gnd cell_6t
Xbit_r159_c220 bl[220] br[220] wl[159] vdd gnd cell_6t
Xbit_r160_c220 bl[220] br[220] wl[160] vdd gnd cell_6t
Xbit_r161_c220 bl[220] br[220] wl[161] vdd gnd cell_6t
Xbit_r162_c220 bl[220] br[220] wl[162] vdd gnd cell_6t
Xbit_r163_c220 bl[220] br[220] wl[163] vdd gnd cell_6t
Xbit_r164_c220 bl[220] br[220] wl[164] vdd gnd cell_6t
Xbit_r165_c220 bl[220] br[220] wl[165] vdd gnd cell_6t
Xbit_r166_c220 bl[220] br[220] wl[166] vdd gnd cell_6t
Xbit_r167_c220 bl[220] br[220] wl[167] vdd gnd cell_6t
Xbit_r168_c220 bl[220] br[220] wl[168] vdd gnd cell_6t
Xbit_r169_c220 bl[220] br[220] wl[169] vdd gnd cell_6t
Xbit_r170_c220 bl[220] br[220] wl[170] vdd gnd cell_6t
Xbit_r171_c220 bl[220] br[220] wl[171] vdd gnd cell_6t
Xbit_r172_c220 bl[220] br[220] wl[172] vdd gnd cell_6t
Xbit_r173_c220 bl[220] br[220] wl[173] vdd gnd cell_6t
Xbit_r174_c220 bl[220] br[220] wl[174] vdd gnd cell_6t
Xbit_r175_c220 bl[220] br[220] wl[175] vdd gnd cell_6t
Xbit_r176_c220 bl[220] br[220] wl[176] vdd gnd cell_6t
Xbit_r177_c220 bl[220] br[220] wl[177] vdd gnd cell_6t
Xbit_r178_c220 bl[220] br[220] wl[178] vdd gnd cell_6t
Xbit_r179_c220 bl[220] br[220] wl[179] vdd gnd cell_6t
Xbit_r180_c220 bl[220] br[220] wl[180] vdd gnd cell_6t
Xbit_r181_c220 bl[220] br[220] wl[181] vdd gnd cell_6t
Xbit_r182_c220 bl[220] br[220] wl[182] vdd gnd cell_6t
Xbit_r183_c220 bl[220] br[220] wl[183] vdd gnd cell_6t
Xbit_r184_c220 bl[220] br[220] wl[184] vdd gnd cell_6t
Xbit_r185_c220 bl[220] br[220] wl[185] vdd gnd cell_6t
Xbit_r186_c220 bl[220] br[220] wl[186] vdd gnd cell_6t
Xbit_r187_c220 bl[220] br[220] wl[187] vdd gnd cell_6t
Xbit_r188_c220 bl[220] br[220] wl[188] vdd gnd cell_6t
Xbit_r189_c220 bl[220] br[220] wl[189] vdd gnd cell_6t
Xbit_r190_c220 bl[220] br[220] wl[190] vdd gnd cell_6t
Xbit_r191_c220 bl[220] br[220] wl[191] vdd gnd cell_6t
Xbit_r192_c220 bl[220] br[220] wl[192] vdd gnd cell_6t
Xbit_r193_c220 bl[220] br[220] wl[193] vdd gnd cell_6t
Xbit_r194_c220 bl[220] br[220] wl[194] vdd gnd cell_6t
Xbit_r195_c220 bl[220] br[220] wl[195] vdd gnd cell_6t
Xbit_r196_c220 bl[220] br[220] wl[196] vdd gnd cell_6t
Xbit_r197_c220 bl[220] br[220] wl[197] vdd gnd cell_6t
Xbit_r198_c220 bl[220] br[220] wl[198] vdd gnd cell_6t
Xbit_r199_c220 bl[220] br[220] wl[199] vdd gnd cell_6t
Xbit_r200_c220 bl[220] br[220] wl[200] vdd gnd cell_6t
Xbit_r201_c220 bl[220] br[220] wl[201] vdd gnd cell_6t
Xbit_r202_c220 bl[220] br[220] wl[202] vdd gnd cell_6t
Xbit_r203_c220 bl[220] br[220] wl[203] vdd gnd cell_6t
Xbit_r204_c220 bl[220] br[220] wl[204] vdd gnd cell_6t
Xbit_r205_c220 bl[220] br[220] wl[205] vdd gnd cell_6t
Xbit_r206_c220 bl[220] br[220] wl[206] vdd gnd cell_6t
Xbit_r207_c220 bl[220] br[220] wl[207] vdd gnd cell_6t
Xbit_r208_c220 bl[220] br[220] wl[208] vdd gnd cell_6t
Xbit_r209_c220 bl[220] br[220] wl[209] vdd gnd cell_6t
Xbit_r210_c220 bl[220] br[220] wl[210] vdd gnd cell_6t
Xbit_r211_c220 bl[220] br[220] wl[211] vdd gnd cell_6t
Xbit_r212_c220 bl[220] br[220] wl[212] vdd gnd cell_6t
Xbit_r213_c220 bl[220] br[220] wl[213] vdd gnd cell_6t
Xbit_r214_c220 bl[220] br[220] wl[214] vdd gnd cell_6t
Xbit_r215_c220 bl[220] br[220] wl[215] vdd gnd cell_6t
Xbit_r216_c220 bl[220] br[220] wl[216] vdd gnd cell_6t
Xbit_r217_c220 bl[220] br[220] wl[217] vdd gnd cell_6t
Xbit_r218_c220 bl[220] br[220] wl[218] vdd gnd cell_6t
Xbit_r219_c220 bl[220] br[220] wl[219] vdd gnd cell_6t
Xbit_r220_c220 bl[220] br[220] wl[220] vdd gnd cell_6t
Xbit_r221_c220 bl[220] br[220] wl[221] vdd gnd cell_6t
Xbit_r222_c220 bl[220] br[220] wl[222] vdd gnd cell_6t
Xbit_r223_c220 bl[220] br[220] wl[223] vdd gnd cell_6t
Xbit_r224_c220 bl[220] br[220] wl[224] vdd gnd cell_6t
Xbit_r225_c220 bl[220] br[220] wl[225] vdd gnd cell_6t
Xbit_r226_c220 bl[220] br[220] wl[226] vdd gnd cell_6t
Xbit_r227_c220 bl[220] br[220] wl[227] vdd gnd cell_6t
Xbit_r228_c220 bl[220] br[220] wl[228] vdd gnd cell_6t
Xbit_r229_c220 bl[220] br[220] wl[229] vdd gnd cell_6t
Xbit_r230_c220 bl[220] br[220] wl[230] vdd gnd cell_6t
Xbit_r231_c220 bl[220] br[220] wl[231] vdd gnd cell_6t
Xbit_r232_c220 bl[220] br[220] wl[232] vdd gnd cell_6t
Xbit_r233_c220 bl[220] br[220] wl[233] vdd gnd cell_6t
Xbit_r234_c220 bl[220] br[220] wl[234] vdd gnd cell_6t
Xbit_r235_c220 bl[220] br[220] wl[235] vdd gnd cell_6t
Xbit_r236_c220 bl[220] br[220] wl[236] vdd gnd cell_6t
Xbit_r237_c220 bl[220] br[220] wl[237] vdd gnd cell_6t
Xbit_r238_c220 bl[220] br[220] wl[238] vdd gnd cell_6t
Xbit_r239_c220 bl[220] br[220] wl[239] vdd gnd cell_6t
Xbit_r240_c220 bl[220] br[220] wl[240] vdd gnd cell_6t
Xbit_r241_c220 bl[220] br[220] wl[241] vdd gnd cell_6t
Xbit_r242_c220 bl[220] br[220] wl[242] vdd gnd cell_6t
Xbit_r243_c220 bl[220] br[220] wl[243] vdd gnd cell_6t
Xbit_r244_c220 bl[220] br[220] wl[244] vdd gnd cell_6t
Xbit_r245_c220 bl[220] br[220] wl[245] vdd gnd cell_6t
Xbit_r246_c220 bl[220] br[220] wl[246] vdd gnd cell_6t
Xbit_r247_c220 bl[220] br[220] wl[247] vdd gnd cell_6t
Xbit_r248_c220 bl[220] br[220] wl[248] vdd gnd cell_6t
Xbit_r249_c220 bl[220] br[220] wl[249] vdd gnd cell_6t
Xbit_r250_c220 bl[220] br[220] wl[250] vdd gnd cell_6t
Xbit_r251_c220 bl[220] br[220] wl[251] vdd gnd cell_6t
Xbit_r252_c220 bl[220] br[220] wl[252] vdd gnd cell_6t
Xbit_r253_c220 bl[220] br[220] wl[253] vdd gnd cell_6t
Xbit_r254_c220 bl[220] br[220] wl[254] vdd gnd cell_6t
Xbit_r255_c220 bl[220] br[220] wl[255] vdd gnd cell_6t
Xbit_r0_c221 bl[221] br[221] wl[0] vdd gnd cell_6t
Xbit_r1_c221 bl[221] br[221] wl[1] vdd gnd cell_6t
Xbit_r2_c221 bl[221] br[221] wl[2] vdd gnd cell_6t
Xbit_r3_c221 bl[221] br[221] wl[3] vdd gnd cell_6t
Xbit_r4_c221 bl[221] br[221] wl[4] vdd gnd cell_6t
Xbit_r5_c221 bl[221] br[221] wl[5] vdd gnd cell_6t
Xbit_r6_c221 bl[221] br[221] wl[6] vdd gnd cell_6t
Xbit_r7_c221 bl[221] br[221] wl[7] vdd gnd cell_6t
Xbit_r8_c221 bl[221] br[221] wl[8] vdd gnd cell_6t
Xbit_r9_c221 bl[221] br[221] wl[9] vdd gnd cell_6t
Xbit_r10_c221 bl[221] br[221] wl[10] vdd gnd cell_6t
Xbit_r11_c221 bl[221] br[221] wl[11] vdd gnd cell_6t
Xbit_r12_c221 bl[221] br[221] wl[12] vdd gnd cell_6t
Xbit_r13_c221 bl[221] br[221] wl[13] vdd gnd cell_6t
Xbit_r14_c221 bl[221] br[221] wl[14] vdd gnd cell_6t
Xbit_r15_c221 bl[221] br[221] wl[15] vdd gnd cell_6t
Xbit_r16_c221 bl[221] br[221] wl[16] vdd gnd cell_6t
Xbit_r17_c221 bl[221] br[221] wl[17] vdd gnd cell_6t
Xbit_r18_c221 bl[221] br[221] wl[18] vdd gnd cell_6t
Xbit_r19_c221 bl[221] br[221] wl[19] vdd gnd cell_6t
Xbit_r20_c221 bl[221] br[221] wl[20] vdd gnd cell_6t
Xbit_r21_c221 bl[221] br[221] wl[21] vdd gnd cell_6t
Xbit_r22_c221 bl[221] br[221] wl[22] vdd gnd cell_6t
Xbit_r23_c221 bl[221] br[221] wl[23] vdd gnd cell_6t
Xbit_r24_c221 bl[221] br[221] wl[24] vdd gnd cell_6t
Xbit_r25_c221 bl[221] br[221] wl[25] vdd gnd cell_6t
Xbit_r26_c221 bl[221] br[221] wl[26] vdd gnd cell_6t
Xbit_r27_c221 bl[221] br[221] wl[27] vdd gnd cell_6t
Xbit_r28_c221 bl[221] br[221] wl[28] vdd gnd cell_6t
Xbit_r29_c221 bl[221] br[221] wl[29] vdd gnd cell_6t
Xbit_r30_c221 bl[221] br[221] wl[30] vdd gnd cell_6t
Xbit_r31_c221 bl[221] br[221] wl[31] vdd gnd cell_6t
Xbit_r32_c221 bl[221] br[221] wl[32] vdd gnd cell_6t
Xbit_r33_c221 bl[221] br[221] wl[33] vdd gnd cell_6t
Xbit_r34_c221 bl[221] br[221] wl[34] vdd gnd cell_6t
Xbit_r35_c221 bl[221] br[221] wl[35] vdd gnd cell_6t
Xbit_r36_c221 bl[221] br[221] wl[36] vdd gnd cell_6t
Xbit_r37_c221 bl[221] br[221] wl[37] vdd gnd cell_6t
Xbit_r38_c221 bl[221] br[221] wl[38] vdd gnd cell_6t
Xbit_r39_c221 bl[221] br[221] wl[39] vdd gnd cell_6t
Xbit_r40_c221 bl[221] br[221] wl[40] vdd gnd cell_6t
Xbit_r41_c221 bl[221] br[221] wl[41] vdd gnd cell_6t
Xbit_r42_c221 bl[221] br[221] wl[42] vdd gnd cell_6t
Xbit_r43_c221 bl[221] br[221] wl[43] vdd gnd cell_6t
Xbit_r44_c221 bl[221] br[221] wl[44] vdd gnd cell_6t
Xbit_r45_c221 bl[221] br[221] wl[45] vdd gnd cell_6t
Xbit_r46_c221 bl[221] br[221] wl[46] vdd gnd cell_6t
Xbit_r47_c221 bl[221] br[221] wl[47] vdd gnd cell_6t
Xbit_r48_c221 bl[221] br[221] wl[48] vdd gnd cell_6t
Xbit_r49_c221 bl[221] br[221] wl[49] vdd gnd cell_6t
Xbit_r50_c221 bl[221] br[221] wl[50] vdd gnd cell_6t
Xbit_r51_c221 bl[221] br[221] wl[51] vdd gnd cell_6t
Xbit_r52_c221 bl[221] br[221] wl[52] vdd gnd cell_6t
Xbit_r53_c221 bl[221] br[221] wl[53] vdd gnd cell_6t
Xbit_r54_c221 bl[221] br[221] wl[54] vdd gnd cell_6t
Xbit_r55_c221 bl[221] br[221] wl[55] vdd gnd cell_6t
Xbit_r56_c221 bl[221] br[221] wl[56] vdd gnd cell_6t
Xbit_r57_c221 bl[221] br[221] wl[57] vdd gnd cell_6t
Xbit_r58_c221 bl[221] br[221] wl[58] vdd gnd cell_6t
Xbit_r59_c221 bl[221] br[221] wl[59] vdd gnd cell_6t
Xbit_r60_c221 bl[221] br[221] wl[60] vdd gnd cell_6t
Xbit_r61_c221 bl[221] br[221] wl[61] vdd gnd cell_6t
Xbit_r62_c221 bl[221] br[221] wl[62] vdd gnd cell_6t
Xbit_r63_c221 bl[221] br[221] wl[63] vdd gnd cell_6t
Xbit_r64_c221 bl[221] br[221] wl[64] vdd gnd cell_6t
Xbit_r65_c221 bl[221] br[221] wl[65] vdd gnd cell_6t
Xbit_r66_c221 bl[221] br[221] wl[66] vdd gnd cell_6t
Xbit_r67_c221 bl[221] br[221] wl[67] vdd gnd cell_6t
Xbit_r68_c221 bl[221] br[221] wl[68] vdd gnd cell_6t
Xbit_r69_c221 bl[221] br[221] wl[69] vdd gnd cell_6t
Xbit_r70_c221 bl[221] br[221] wl[70] vdd gnd cell_6t
Xbit_r71_c221 bl[221] br[221] wl[71] vdd gnd cell_6t
Xbit_r72_c221 bl[221] br[221] wl[72] vdd gnd cell_6t
Xbit_r73_c221 bl[221] br[221] wl[73] vdd gnd cell_6t
Xbit_r74_c221 bl[221] br[221] wl[74] vdd gnd cell_6t
Xbit_r75_c221 bl[221] br[221] wl[75] vdd gnd cell_6t
Xbit_r76_c221 bl[221] br[221] wl[76] vdd gnd cell_6t
Xbit_r77_c221 bl[221] br[221] wl[77] vdd gnd cell_6t
Xbit_r78_c221 bl[221] br[221] wl[78] vdd gnd cell_6t
Xbit_r79_c221 bl[221] br[221] wl[79] vdd gnd cell_6t
Xbit_r80_c221 bl[221] br[221] wl[80] vdd gnd cell_6t
Xbit_r81_c221 bl[221] br[221] wl[81] vdd gnd cell_6t
Xbit_r82_c221 bl[221] br[221] wl[82] vdd gnd cell_6t
Xbit_r83_c221 bl[221] br[221] wl[83] vdd gnd cell_6t
Xbit_r84_c221 bl[221] br[221] wl[84] vdd gnd cell_6t
Xbit_r85_c221 bl[221] br[221] wl[85] vdd gnd cell_6t
Xbit_r86_c221 bl[221] br[221] wl[86] vdd gnd cell_6t
Xbit_r87_c221 bl[221] br[221] wl[87] vdd gnd cell_6t
Xbit_r88_c221 bl[221] br[221] wl[88] vdd gnd cell_6t
Xbit_r89_c221 bl[221] br[221] wl[89] vdd gnd cell_6t
Xbit_r90_c221 bl[221] br[221] wl[90] vdd gnd cell_6t
Xbit_r91_c221 bl[221] br[221] wl[91] vdd gnd cell_6t
Xbit_r92_c221 bl[221] br[221] wl[92] vdd gnd cell_6t
Xbit_r93_c221 bl[221] br[221] wl[93] vdd gnd cell_6t
Xbit_r94_c221 bl[221] br[221] wl[94] vdd gnd cell_6t
Xbit_r95_c221 bl[221] br[221] wl[95] vdd gnd cell_6t
Xbit_r96_c221 bl[221] br[221] wl[96] vdd gnd cell_6t
Xbit_r97_c221 bl[221] br[221] wl[97] vdd gnd cell_6t
Xbit_r98_c221 bl[221] br[221] wl[98] vdd gnd cell_6t
Xbit_r99_c221 bl[221] br[221] wl[99] vdd gnd cell_6t
Xbit_r100_c221 bl[221] br[221] wl[100] vdd gnd cell_6t
Xbit_r101_c221 bl[221] br[221] wl[101] vdd gnd cell_6t
Xbit_r102_c221 bl[221] br[221] wl[102] vdd gnd cell_6t
Xbit_r103_c221 bl[221] br[221] wl[103] vdd gnd cell_6t
Xbit_r104_c221 bl[221] br[221] wl[104] vdd gnd cell_6t
Xbit_r105_c221 bl[221] br[221] wl[105] vdd gnd cell_6t
Xbit_r106_c221 bl[221] br[221] wl[106] vdd gnd cell_6t
Xbit_r107_c221 bl[221] br[221] wl[107] vdd gnd cell_6t
Xbit_r108_c221 bl[221] br[221] wl[108] vdd gnd cell_6t
Xbit_r109_c221 bl[221] br[221] wl[109] vdd gnd cell_6t
Xbit_r110_c221 bl[221] br[221] wl[110] vdd gnd cell_6t
Xbit_r111_c221 bl[221] br[221] wl[111] vdd gnd cell_6t
Xbit_r112_c221 bl[221] br[221] wl[112] vdd gnd cell_6t
Xbit_r113_c221 bl[221] br[221] wl[113] vdd gnd cell_6t
Xbit_r114_c221 bl[221] br[221] wl[114] vdd gnd cell_6t
Xbit_r115_c221 bl[221] br[221] wl[115] vdd gnd cell_6t
Xbit_r116_c221 bl[221] br[221] wl[116] vdd gnd cell_6t
Xbit_r117_c221 bl[221] br[221] wl[117] vdd gnd cell_6t
Xbit_r118_c221 bl[221] br[221] wl[118] vdd gnd cell_6t
Xbit_r119_c221 bl[221] br[221] wl[119] vdd gnd cell_6t
Xbit_r120_c221 bl[221] br[221] wl[120] vdd gnd cell_6t
Xbit_r121_c221 bl[221] br[221] wl[121] vdd gnd cell_6t
Xbit_r122_c221 bl[221] br[221] wl[122] vdd gnd cell_6t
Xbit_r123_c221 bl[221] br[221] wl[123] vdd gnd cell_6t
Xbit_r124_c221 bl[221] br[221] wl[124] vdd gnd cell_6t
Xbit_r125_c221 bl[221] br[221] wl[125] vdd gnd cell_6t
Xbit_r126_c221 bl[221] br[221] wl[126] vdd gnd cell_6t
Xbit_r127_c221 bl[221] br[221] wl[127] vdd gnd cell_6t
Xbit_r128_c221 bl[221] br[221] wl[128] vdd gnd cell_6t
Xbit_r129_c221 bl[221] br[221] wl[129] vdd gnd cell_6t
Xbit_r130_c221 bl[221] br[221] wl[130] vdd gnd cell_6t
Xbit_r131_c221 bl[221] br[221] wl[131] vdd gnd cell_6t
Xbit_r132_c221 bl[221] br[221] wl[132] vdd gnd cell_6t
Xbit_r133_c221 bl[221] br[221] wl[133] vdd gnd cell_6t
Xbit_r134_c221 bl[221] br[221] wl[134] vdd gnd cell_6t
Xbit_r135_c221 bl[221] br[221] wl[135] vdd gnd cell_6t
Xbit_r136_c221 bl[221] br[221] wl[136] vdd gnd cell_6t
Xbit_r137_c221 bl[221] br[221] wl[137] vdd gnd cell_6t
Xbit_r138_c221 bl[221] br[221] wl[138] vdd gnd cell_6t
Xbit_r139_c221 bl[221] br[221] wl[139] vdd gnd cell_6t
Xbit_r140_c221 bl[221] br[221] wl[140] vdd gnd cell_6t
Xbit_r141_c221 bl[221] br[221] wl[141] vdd gnd cell_6t
Xbit_r142_c221 bl[221] br[221] wl[142] vdd gnd cell_6t
Xbit_r143_c221 bl[221] br[221] wl[143] vdd gnd cell_6t
Xbit_r144_c221 bl[221] br[221] wl[144] vdd gnd cell_6t
Xbit_r145_c221 bl[221] br[221] wl[145] vdd gnd cell_6t
Xbit_r146_c221 bl[221] br[221] wl[146] vdd gnd cell_6t
Xbit_r147_c221 bl[221] br[221] wl[147] vdd gnd cell_6t
Xbit_r148_c221 bl[221] br[221] wl[148] vdd gnd cell_6t
Xbit_r149_c221 bl[221] br[221] wl[149] vdd gnd cell_6t
Xbit_r150_c221 bl[221] br[221] wl[150] vdd gnd cell_6t
Xbit_r151_c221 bl[221] br[221] wl[151] vdd gnd cell_6t
Xbit_r152_c221 bl[221] br[221] wl[152] vdd gnd cell_6t
Xbit_r153_c221 bl[221] br[221] wl[153] vdd gnd cell_6t
Xbit_r154_c221 bl[221] br[221] wl[154] vdd gnd cell_6t
Xbit_r155_c221 bl[221] br[221] wl[155] vdd gnd cell_6t
Xbit_r156_c221 bl[221] br[221] wl[156] vdd gnd cell_6t
Xbit_r157_c221 bl[221] br[221] wl[157] vdd gnd cell_6t
Xbit_r158_c221 bl[221] br[221] wl[158] vdd gnd cell_6t
Xbit_r159_c221 bl[221] br[221] wl[159] vdd gnd cell_6t
Xbit_r160_c221 bl[221] br[221] wl[160] vdd gnd cell_6t
Xbit_r161_c221 bl[221] br[221] wl[161] vdd gnd cell_6t
Xbit_r162_c221 bl[221] br[221] wl[162] vdd gnd cell_6t
Xbit_r163_c221 bl[221] br[221] wl[163] vdd gnd cell_6t
Xbit_r164_c221 bl[221] br[221] wl[164] vdd gnd cell_6t
Xbit_r165_c221 bl[221] br[221] wl[165] vdd gnd cell_6t
Xbit_r166_c221 bl[221] br[221] wl[166] vdd gnd cell_6t
Xbit_r167_c221 bl[221] br[221] wl[167] vdd gnd cell_6t
Xbit_r168_c221 bl[221] br[221] wl[168] vdd gnd cell_6t
Xbit_r169_c221 bl[221] br[221] wl[169] vdd gnd cell_6t
Xbit_r170_c221 bl[221] br[221] wl[170] vdd gnd cell_6t
Xbit_r171_c221 bl[221] br[221] wl[171] vdd gnd cell_6t
Xbit_r172_c221 bl[221] br[221] wl[172] vdd gnd cell_6t
Xbit_r173_c221 bl[221] br[221] wl[173] vdd gnd cell_6t
Xbit_r174_c221 bl[221] br[221] wl[174] vdd gnd cell_6t
Xbit_r175_c221 bl[221] br[221] wl[175] vdd gnd cell_6t
Xbit_r176_c221 bl[221] br[221] wl[176] vdd gnd cell_6t
Xbit_r177_c221 bl[221] br[221] wl[177] vdd gnd cell_6t
Xbit_r178_c221 bl[221] br[221] wl[178] vdd gnd cell_6t
Xbit_r179_c221 bl[221] br[221] wl[179] vdd gnd cell_6t
Xbit_r180_c221 bl[221] br[221] wl[180] vdd gnd cell_6t
Xbit_r181_c221 bl[221] br[221] wl[181] vdd gnd cell_6t
Xbit_r182_c221 bl[221] br[221] wl[182] vdd gnd cell_6t
Xbit_r183_c221 bl[221] br[221] wl[183] vdd gnd cell_6t
Xbit_r184_c221 bl[221] br[221] wl[184] vdd gnd cell_6t
Xbit_r185_c221 bl[221] br[221] wl[185] vdd gnd cell_6t
Xbit_r186_c221 bl[221] br[221] wl[186] vdd gnd cell_6t
Xbit_r187_c221 bl[221] br[221] wl[187] vdd gnd cell_6t
Xbit_r188_c221 bl[221] br[221] wl[188] vdd gnd cell_6t
Xbit_r189_c221 bl[221] br[221] wl[189] vdd gnd cell_6t
Xbit_r190_c221 bl[221] br[221] wl[190] vdd gnd cell_6t
Xbit_r191_c221 bl[221] br[221] wl[191] vdd gnd cell_6t
Xbit_r192_c221 bl[221] br[221] wl[192] vdd gnd cell_6t
Xbit_r193_c221 bl[221] br[221] wl[193] vdd gnd cell_6t
Xbit_r194_c221 bl[221] br[221] wl[194] vdd gnd cell_6t
Xbit_r195_c221 bl[221] br[221] wl[195] vdd gnd cell_6t
Xbit_r196_c221 bl[221] br[221] wl[196] vdd gnd cell_6t
Xbit_r197_c221 bl[221] br[221] wl[197] vdd gnd cell_6t
Xbit_r198_c221 bl[221] br[221] wl[198] vdd gnd cell_6t
Xbit_r199_c221 bl[221] br[221] wl[199] vdd gnd cell_6t
Xbit_r200_c221 bl[221] br[221] wl[200] vdd gnd cell_6t
Xbit_r201_c221 bl[221] br[221] wl[201] vdd gnd cell_6t
Xbit_r202_c221 bl[221] br[221] wl[202] vdd gnd cell_6t
Xbit_r203_c221 bl[221] br[221] wl[203] vdd gnd cell_6t
Xbit_r204_c221 bl[221] br[221] wl[204] vdd gnd cell_6t
Xbit_r205_c221 bl[221] br[221] wl[205] vdd gnd cell_6t
Xbit_r206_c221 bl[221] br[221] wl[206] vdd gnd cell_6t
Xbit_r207_c221 bl[221] br[221] wl[207] vdd gnd cell_6t
Xbit_r208_c221 bl[221] br[221] wl[208] vdd gnd cell_6t
Xbit_r209_c221 bl[221] br[221] wl[209] vdd gnd cell_6t
Xbit_r210_c221 bl[221] br[221] wl[210] vdd gnd cell_6t
Xbit_r211_c221 bl[221] br[221] wl[211] vdd gnd cell_6t
Xbit_r212_c221 bl[221] br[221] wl[212] vdd gnd cell_6t
Xbit_r213_c221 bl[221] br[221] wl[213] vdd gnd cell_6t
Xbit_r214_c221 bl[221] br[221] wl[214] vdd gnd cell_6t
Xbit_r215_c221 bl[221] br[221] wl[215] vdd gnd cell_6t
Xbit_r216_c221 bl[221] br[221] wl[216] vdd gnd cell_6t
Xbit_r217_c221 bl[221] br[221] wl[217] vdd gnd cell_6t
Xbit_r218_c221 bl[221] br[221] wl[218] vdd gnd cell_6t
Xbit_r219_c221 bl[221] br[221] wl[219] vdd gnd cell_6t
Xbit_r220_c221 bl[221] br[221] wl[220] vdd gnd cell_6t
Xbit_r221_c221 bl[221] br[221] wl[221] vdd gnd cell_6t
Xbit_r222_c221 bl[221] br[221] wl[222] vdd gnd cell_6t
Xbit_r223_c221 bl[221] br[221] wl[223] vdd gnd cell_6t
Xbit_r224_c221 bl[221] br[221] wl[224] vdd gnd cell_6t
Xbit_r225_c221 bl[221] br[221] wl[225] vdd gnd cell_6t
Xbit_r226_c221 bl[221] br[221] wl[226] vdd gnd cell_6t
Xbit_r227_c221 bl[221] br[221] wl[227] vdd gnd cell_6t
Xbit_r228_c221 bl[221] br[221] wl[228] vdd gnd cell_6t
Xbit_r229_c221 bl[221] br[221] wl[229] vdd gnd cell_6t
Xbit_r230_c221 bl[221] br[221] wl[230] vdd gnd cell_6t
Xbit_r231_c221 bl[221] br[221] wl[231] vdd gnd cell_6t
Xbit_r232_c221 bl[221] br[221] wl[232] vdd gnd cell_6t
Xbit_r233_c221 bl[221] br[221] wl[233] vdd gnd cell_6t
Xbit_r234_c221 bl[221] br[221] wl[234] vdd gnd cell_6t
Xbit_r235_c221 bl[221] br[221] wl[235] vdd gnd cell_6t
Xbit_r236_c221 bl[221] br[221] wl[236] vdd gnd cell_6t
Xbit_r237_c221 bl[221] br[221] wl[237] vdd gnd cell_6t
Xbit_r238_c221 bl[221] br[221] wl[238] vdd gnd cell_6t
Xbit_r239_c221 bl[221] br[221] wl[239] vdd gnd cell_6t
Xbit_r240_c221 bl[221] br[221] wl[240] vdd gnd cell_6t
Xbit_r241_c221 bl[221] br[221] wl[241] vdd gnd cell_6t
Xbit_r242_c221 bl[221] br[221] wl[242] vdd gnd cell_6t
Xbit_r243_c221 bl[221] br[221] wl[243] vdd gnd cell_6t
Xbit_r244_c221 bl[221] br[221] wl[244] vdd gnd cell_6t
Xbit_r245_c221 bl[221] br[221] wl[245] vdd gnd cell_6t
Xbit_r246_c221 bl[221] br[221] wl[246] vdd gnd cell_6t
Xbit_r247_c221 bl[221] br[221] wl[247] vdd gnd cell_6t
Xbit_r248_c221 bl[221] br[221] wl[248] vdd gnd cell_6t
Xbit_r249_c221 bl[221] br[221] wl[249] vdd gnd cell_6t
Xbit_r250_c221 bl[221] br[221] wl[250] vdd gnd cell_6t
Xbit_r251_c221 bl[221] br[221] wl[251] vdd gnd cell_6t
Xbit_r252_c221 bl[221] br[221] wl[252] vdd gnd cell_6t
Xbit_r253_c221 bl[221] br[221] wl[253] vdd gnd cell_6t
Xbit_r254_c221 bl[221] br[221] wl[254] vdd gnd cell_6t
Xbit_r255_c221 bl[221] br[221] wl[255] vdd gnd cell_6t
Xbit_r0_c222 bl[222] br[222] wl[0] vdd gnd cell_6t
Xbit_r1_c222 bl[222] br[222] wl[1] vdd gnd cell_6t
Xbit_r2_c222 bl[222] br[222] wl[2] vdd gnd cell_6t
Xbit_r3_c222 bl[222] br[222] wl[3] vdd gnd cell_6t
Xbit_r4_c222 bl[222] br[222] wl[4] vdd gnd cell_6t
Xbit_r5_c222 bl[222] br[222] wl[5] vdd gnd cell_6t
Xbit_r6_c222 bl[222] br[222] wl[6] vdd gnd cell_6t
Xbit_r7_c222 bl[222] br[222] wl[7] vdd gnd cell_6t
Xbit_r8_c222 bl[222] br[222] wl[8] vdd gnd cell_6t
Xbit_r9_c222 bl[222] br[222] wl[9] vdd gnd cell_6t
Xbit_r10_c222 bl[222] br[222] wl[10] vdd gnd cell_6t
Xbit_r11_c222 bl[222] br[222] wl[11] vdd gnd cell_6t
Xbit_r12_c222 bl[222] br[222] wl[12] vdd gnd cell_6t
Xbit_r13_c222 bl[222] br[222] wl[13] vdd gnd cell_6t
Xbit_r14_c222 bl[222] br[222] wl[14] vdd gnd cell_6t
Xbit_r15_c222 bl[222] br[222] wl[15] vdd gnd cell_6t
Xbit_r16_c222 bl[222] br[222] wl[16] vdd gnd cell_6t
Xbit_r17_c222 bl[222] br[222] wl[17] vdd gnd cell_6t
Xbit_r18_c222 bl[222] br[222] wl[18] vdd gnd cell_6t
Xbit_r19_c222 bl[222] br[222] wl[19] vdd gnd cell_6t
Xbit_r20_c222 bl[222] br[222] wl[20] vdd gnd cell_6t
Xbit_r21_c222 bl[222] br[222] wl[21] vdd gnd cell_6t
Xbit_r22_c222 bl[222] br[222] wl[22] vdd gnd cell_6t
Xbit_r23_c222 bl[222] br[222] wl[23] vdd gnd cell_6t
Xbit_r24_c222 bl[222] br[222] wl[24] vdd gnd cell_6t
Xbit_r25_c222 bl[222] br[222] wl[25] vdd gnd cell_6t
Xbit_r26_c222 bl[222] br[222] wl[26] vdd gnd cell_6t
Xbit_r27_c222 bl[222] br[222] wl[27] vdd gnd cell_6t
Xbit_r28_c222 bl[222] br[222] wl[28] vdd gnd cell_6t
Xbit_r29_c222 bl[222] br[222] wl[29] vdd gnd cell_6t
Xbit_r30_c222 bl[222] br[222] wl[30] vdd gnd cell_6t
Xbit_r31_c222 bl[222] br[222] wl[31] vdd gnd cell_6t
Xbit_r32_c222 bl[222] br[222] wl[32] vdd gnd cell_6t
Xbit_r33_c222 bl[222] br[222] wl[33] vdd gnd cell_6t
Xbit_r34_c222 bl[222] br[222] wl[34] vdd gnd cell_6t
Xbit_r35_c222 bl[222] br[222] wl[35] vdd gnd cell_6t
Xbit_r36_c222 bl[222] br[222] wl[36] vdd gnd cell_6t
Xbit_r37_c222 bl[222] br[222] wl[37] vdd gnd cell_6t
Xbit_r38_c222 bl[222] br[222] wl[38] vdd gnd cell_6t
Xbit_r39_c222 bl[222] br[222] wl[39] vdd gnd cell_6t
Xbit_r40_c222 bl[222] br[222] wl[40] vdd gnd cell_6t
Xbit_r41_c222 bl[222] br[222] wl[41] vdd gnd cell_6t
Xbit_r42_c222 bl[222] br[222] wl[42] vdd gnd cell_6t
Xbit_r43_c222 bl[222] br[222] wl[43] vdd gnd cell_6t
Xbit_r44_c222 bl[222] br[222] wl[44] vdd gnd cell_6t
Xbit_r45_c222 bl[222] br[222] wl[45] vdd gnd cell_6t
Xbit_r46_c222 bl[222] br[222] wl[46] vdd gnd cell_6t
Xbit_r47_c222 bl[222] br[222] wl[47] vdd gnd cell_6t
Xbit_r48_c222 bl[222] br[222] wl[48] vdd gnd cell_6t
Xbit_r49_c222 bl[222] br[222] wl[49] vdd gnd cell_6t
Xbit_r50_c222 bl[222] br[222] wl[50] vdd gnd cell_6t
Xbit_r51_c222 bl[222] br[222] wl[51] vdd gnd cell_6t
Xbit_r52_c222 bl[222] br[222] wl[52] vdd gnd cell_6t
Xbit_r53_c222 bl[222] br[222] wl[53] vdd gnd cell_6t
Xbit_r54_c222 bl[222] br[222] wl[54] vdd gnd cell_6t
Xbit_r55_c222 bl[222] br[222] wl[55] vdd gnd cell_6t
Xbit_r56_c222 bl[222] br[222] wl[56] vdd gnd cell_6t
Xbit_r57_c222 bl[222] br[222] wl[57] vdd gnd cell_6t
Xbit_r58_c222 bl[222] br[222] wl[58] vdd gnd cell_6t
Xbit_r59_c222 bl[222] br[222] wl[59] vdd gnd cell_6t
Xbit_r60_c222 bl[222] br[222] wl[60] vdd gnd cell_6t
Xbit_r61_c222 bl[222] br[222] wl[61] vdd gnd cell_6t
Xbit_r62_c222 bl[222] br[222] wl[62] vdd gnd cell_6t
Xbit_r63_c222 bl[222] br[222] wl[63] vdd gnd cell_6t
Xbit_r64_c222 bl[222] br[222] wl[64] vdd gnd cell_6t
Xbit_r65_c222 bl[222] br[222] wl[65] vdd gnd cell_6t
Xbit_r66_c222 bl[222] br[222] wl[66] vdd gnd cell_6t
Xbit_r67_c222 bl[222] br[222] wl[67] vdd gnd cell_6t
Xbit_r68_c222 bl[222] br[222] wl[68] vdd gnd cell_6t
Xbit_r69_c222 bl[222] br[222] wl[69] vdd gnd cell_6t
Xbit_r70_c222 bl[222] br[222] wl[70] vdd gnd cell_6t
Xbit_r71_c222 bl[222] br[222] wl[71] vdd gnd cell_6t
Xbit_r72_c222 bl[222] br[222] wl[72] vdd gnd cell_6t
Xbit_r73_c222 bl[222] br[222] wl[73] vdd gnd cell_6t
Xbit_r74_c222 bl[222] br[222] wl[74] vdd gnd cell_6t
Xbit_r75_c222 bl[222] br[222] wl[75] vdd gnd cell_6t
Xbit_r76_c222 bl[222] br[222] wl[76] vdd gnd cell_6t
Xbit_r77_c222 bl[222] br[222] wl[77] vdd gnd cell_6t
Xbit_r78_c222 bl[222] br[222] wl[78] vdd gnd cell_6t
Xbit_r79_c222 bl[222] br[222] wl[79] vdd gnd cell_6t
Xbit_r80_c222 bl[222] br[222] wl[80] vdd gnd cell_6t
Xbit_r81_c222 bl[222] br[222] wl[81] vdd gnd cell_6t
Xbit_r82_c222 bl[222] br[222] wl[82] vdd gnd cell_6t
Xbit_r83_c222 bl[222] br[222] wl[83] vdd gnd cell_6t
Xbit_r84_c222 bl[222] br[222] wl[84] vdd gnd cell_6t
Xbit_r85_c222 bl[222] br[222] wl[85] vdd gnd cell_6t
Xbit_r86_c222 bl[222] br[222] wl[86] vdd gnd cell_6t
Xbit_r87_c222 bl[222] br[222] wl[87] vdd gnd cell_6t
Xbit_r88_c222 bl[222] br[222] wl[88] vdd gnd cell_6t
Xbit_r89_c222 bl[222] br[222] wl[89] vdd gnd cell_6t
Xbit_r90_c222 bl[222] br[222] wl[90] vdd gnd cell_6t
Xbit_r91_c222 bl[222] br[222] wl[91] vdd gnd cell_6t
Xbit_r92_c222 bl[222] br[222] wl[92] vdd gnd cell_6t
Xbit_r93_c222 bl[222] br[222] wl[93] vdd gnd cell_6t
Xbit_r94_c222 bl[222] br[222] wl[94] vdd gnd cell_6t
Xbit_r95_c222 bl[222] br[222] wl[95] vdd gnd cell_6t
Xbit_r96_c222 bl[222] br[222] wl[96] vdd gnd cell_6t
Xbit_r97_c222 bl[222] br[222] wl[97] vdd gnd cell_6t
Xbit_r98_c222 bl[222] br[222] wl[98] vdd gnd cell_6t
Xbit_r99_c222 bl[222] br[222] wl[99] vdd gnd cell_6t
Xbit_r100_c222 bl[222] br[222] wl[100] vdd gnd cell_6t
Xbit_r101_c222 bl[222] br[222] wl[101] vdd gnd cell_6t
Xbit_r102_c222 bl[222] br[222] wl[102] vdd gnd cell_6t
Xbit_r103_c222 bl[222] br[222] wl[103] vdd gnd cell_6t
Xbit_r104_c222 bl[222] br[222] wl[104] vdd gnd cell_6t
Xbit_r105_c222 bl[222] br[222] wl[105] vdd gnd cell_6t
Xbit_r106_c222 bl[222] br[222] wl[106] vdd gnd cell_6t
Xbit_r107_c222 bl[222] br[222] wl[107] vdd gnd cell_6t
Xbit_r108_c222 bl[222] br[222] wl[108] vdd gnd cell_6t
Xbit_r109_c222 bl[222] br[222] wl[109] vdd gnd cell_6t
Xbit_r110_c222 bl[222] br[222] wl[110] vdd gnd cell_6t
Xbit_r111_c222 bl[222] br[222] wl[111] vdd gnd cell_6t
Xbit_r112_c222 bl[222] br[222] wl[112] vdd gnd cell_6t
Xbit_r113_c222 bl[222] br[222] wl[113] vdd gnd cell_6t
Xbit_r114_c222 bl[222] br[222] wl[114] vdd gnd cell_6t
Xbit_r115_c222 bl[222] br[222] wl[115] vdd gnd cell_6t
Xbit_r116_c222 bl[222] br[222] wl[116] vdd gnd cell_6t
Xbit_r117_c222 bl[222] br[222] wl[117] vdd gnd cell_6t
Xbit_r118_c222 bl[222] br[222] wl[118] vdd gnd cell_6t
Xbit_r119_c222 bl[222] br[222] wl[119] vdd gnd cell_6t
Xbit_r120_c222 bl[222] br[222] wl[120] vdd gnd cell_6t
Xbit_r121_c222 bl[222] br[222] wl[121] vdd gnd cell_6t
Xbit_r122_c222 bl[222] br[222] wl[122] vdd gnd cell_6t
Xbit_r123_c222 bl[222] br[222] wl[123] vdd gnd cell_6t
Xbit_r124_c222 bl[222] br[222] wl[124] vdd gnd cell_6t
Xbit_r125_c222 bl[222] br[222] wl[125] vdd gnd cell_6t
Xbit_r126_c222 bl[222] br[222] wl[126] vdd gnd cell_6t
Xbit_r127_c222 bl[222] br[222] wl[127] vdd gnd cell_6t
Xbit_r128_c222 bl[222] br[222] wl[128] vdd gnd cell_6t
Xbit_r129_c222 bl[222] br[222] wl[129] vdd gnd cell_6t
Xbit_r130_c222 bl[222] br[222] wl[130] vdd gnd cell_6t
Xbit_r131_c222 bl[222] br[222] wl[131] vdd gnd cell_6t
Xbit_r132_c222 bl[222] br[222] wl[132] vdd gnd cell_6t
Xbit_r133_c222 bl[222] br[222] wl[133] vdd gnd cell_6t
Xbit_r134_c222 bl[222] br[222] wl[134] vdd gnd cell_6t
Xbit_r135_c222 bl[222] br[222] wl[135] vdd gnd cell_6t
Xbit_r136_c222 bl[222] br[222] wl[136] vdd gnd cell_6t
Xbit_r137_c222 bl[222] br[222] wl[137] vdd gnd cell_6t
Xbit_r138_c222 bl[222] br[222] wl[138] vdd gnd cell_6t
Xbit_r139_c222 bl[222] br[222] wl[139] vdd gnd cell_6t
Xbit_r140_c222 bl[222] br[222] wl[140] vdd gnd cell_6t
Xbit_r141_c222 bl[222] br[222] wl[141] vdd gnd cell_6t
Xbit_r142_c222 bl[222] br[222] wl[142] vdd gnd cell_6t
Xbit_r143_c222 bl[222] br[222] wl[143] vdd gnd cell_6t
Xbit_r144_c222 bl[222] br[222] wl[144] vdd gnd cell_6t
Xbit_r145_c222 bl[222] br[222] wl[145] vdd gnd cell_6t
Xbit_r146_c222 bl[222] br[222] wl[146] vdd gnd cell_6t
Xbit_r147_c222 bl[222] br[222] wl[147] vdd gnd cell_6t
Xbit_r148_c222 bl[222] br[222] wl[148] vdd gnd cell_6t
Xbit_r149_c222 bl[222] br[222] wl[149] vdd gnd cell_6t
Xbit_r150_c222 bl[222] br[222] wl[150] vdd gnd cell_6t
Xbit_r151_c222 bl[222] br[222] wl[151] vdd gnd cell_6t
Xbit_r152_c222 bl[222] br[222] wl[152] vdd gnd cell_6t
Xbit_r153_c222 bl[222] br[222] wl[153] vdd gnd cell_6t
Xbit_r154_c222 bl[222] br[222] wl[154] vdd gnd cell_6t
Xbit_r155_c222 bl[222] br[222] wl[155] vdd gnd cell_6t
Xbit_r156_c222 bl[222] br[222] wl[156] vdd gnd cell_6t
Xbit_r157_c222 bl[222] br[222] wl[157] vdd gnd cell_6t
Xbit_r158_c222 bl[222] br[222] wl[158] vdd gnd cell_6t
Xbit_r159_c222 bl[222] br[222] wl[159] vdd gnd cell_6t
Xbit_r160_c222 bl[222] br[222] wl[160] vdd gnd cell_6t
Xbit_r161_c222 bl[222] br[222] wl[161] vdd gnd cell_6t
Xbit_r162_c222 bl[222] br[222] wl[162] vdd gnd cell_6t
Xbit_r163_c222 bl[222] br[222] wl[163] vdd gnd cell_6t
Xbit_r164_c222 bl[222] br[222] wl[164] vdd gnd cell_6t
Xbit_r165_c222 bl[222] br[222] wl[165] vdd gnd cell_6t
Xbit_r166_c222 bl[222] br[222] wl[166] vdd gnd cell_6t
Xbit_r167_c222 bl[222] br[222] wl[167] vdd gnd cell_6t
Xbit_r168_c222 bl[222] br[222] wl[168] vdd gnd cell_6t
Xbit_r169_c222 bl[222] br[222] wl[169] vdd gnd cell_6t
Xbit_r170_c222 bl[222] br[222] wl[170] vdd gnd cell_6t
Xbit_r171_c222 bl[222] br[222] wl[171] vdd gnd cell_6t
Xbit_r172_c222 bl[222] br[222] wl[172] vdd gnd cell_6t
Xbit_r173_c222 bl[222] br[222] wl[173] vdd gnd cell_6t
Xbit_r174_c222 bl[222] br[222] wl[174] vdd gnd cell_6t
Xbit_r175_c222 bl[222] br[222] wl[175] vdd gnd cell_6t
Xbit_r176_c222 bl[222] br[222] wl[176] vdd gnd cell_6t
Xbit_r177_c222 bl[222] br[222] wl[177] vdd gnd cell_6t
Xbit_r178_c222 bl[222] br[222] wl[178] vdd gnd cell_6t
Xbit_r179_c222 bl[222] br[222] wl[179] vdd gnd cell_6t
Xbit_r180_c222 bl[222] br[222] wl[180] vdd gnd cell_6t
Xbit_r181_c222 bl[222] br[222] wl[181] vdd gnd cell_6t
Xbit_r182_c222 bl[222] br[222] wl[182] vdd gnd cell_6t
Xbit_r183_c222 bl[222] br[222] wl[183] vdd gnd cell_6t
Xbit_r184_c222 bl[222] br[222] wl[184] vdd gnd cell_6t
Xbit_r185_c222 bl[222] br[222] wl[185] vdd gnd cell_6t
Xbit_r186_c222 bl[222] br[222] wl[186] vdd gnd cell_6t
Xbit_r187_c222 bl[222] br[222] wl[187] vdd gnd cell_6t
Xbit_r188_c222 bl[222] br[222] wl[188] vdd gnd cell_6t
Xbit_r189_c222 bl[222] br[222] wl[189] vdd gnd cell_6t
Xbit_r190_c222 bl[222] br[222] wl[190] vdd gnd cell_6t
Xbit_r191_c222 bl[222] br[222] wl[191] vdd gnd cell_6t
Xbit_r192_c222 bl[222] br[222] wl[192] vdd gnd cell_6t
Xbit_r193_c222 bl[222] br[222] wl[193] vdd gnd cell_6t
Xbit_r194_c222 bl[222] br[222] wl[194] vdd gnd cell_6t
Xbit_r195_c222 bl[222] br[222] wl[195] vdd gnd cell_6t
Xbit_r196_c222 bl[222] br[222] wl[196] vdd gnd cell_6t
Xbit_r197_c222 bl[222] br[222] wl[197] vdd gnd cell_6t
Xbit_r198_c222 bl[222] br[222] wl[198] vdd gnd cell_6t
Xbit_r199_c222 bl[222] br[222] wl[199] vdd gnd cell_6t
Xbit_r200_c222 bl[222] br[222] wl[200] vdd gnd cell_6t
Xbit_r201_c222 bl[222] br[222] wl[201] vdd gnd cell_6t
Xbit_r202_c222 bl[222] br[222] wl[202] vdd gnd cell_6t
Xbit_r203_c222 bl[222] br[222] wl[203] vdd gnd cell_6t
Xbit_r204_c222 bl[222] br[222] wl[204] vdd gnd cell_6t
Xbit_r205_c222 bl[222] br[222] wl[205] vdd gnd cell_6t
Xbit_r206_c222 bl[222] br[222] wl[206] vdd gnd cell_6t
Xbit_r207_c222 bl[222] br[222] wl[207] vdd gnd cell_6t
Xbit_r208_c222 bl[222] br[222] wl[208] vdd gnd cell_6t
Xbit_r209_c222 bl[222] br[222] wl[209] vdd gnd cell_6t
Xbit_r210_c222 bl[222] br[222] wl[210] vdd gnd cell_6t
Xbit_r211_c222 bl[222] br[222] wl[211] vdd gnd cell_6t
Xbit_r212_c222 bl[222] br[222] wl[212] vdd gnd cell_6t
Xbit_r213_c222 bl[222] br[222] wl[213] vdd gnd cell_6t
Xbit_r214_c222 bl[222] br[222] wl[214] vdd gnd cell_6t
Xbit_r215_c222 bl[222] br[222] wl[215] vdd gnd cell_6t
Xbit_r216_c222 bl[222] br[222] wl[216] vdd gnd cell_6t
Xbit_r217_c222 bl[222] br[222] wl[217] vdd gnd cell_6t
Xbit_r218_c222 bl[222] br[222] wl[218] vdd gnd cell_6t
Xbit_r219_c222 bl[222] br[222] wl[219] vdd gnd cell_6t
Xbit_r220_c222 bl[222] br[222] wl[220] vdd gnd cell_6t
Xbit_r221_c222 bl[222] br[222] wl[221] vdd gnd cell_6t
Xbit_r222_c222 bl[222] br[222] wl[222] vdd gnd cell_6t
Xbit_r223_c222 bl[222] br[222] wl[223] vdd gnd cell_6t
Xbit_r224_c222 bl[222] br[222] wl[224] vdd gnd cell_6t
Xbit_r225_c222 bl[222] br[222] wl[225] vdd gnd cell_6t
Xbit_r226_c222 bl[222] br[222] wl[226] vdd gnd cell_6t
Xbit_r227_c222 bl[222] br[222] wl[227] vdd gnd cell_6t
Xbit_r228_c222 bl[222] br[222] wl[228] vdd gnd cell_6t
Xbit_r229_c222 bl[222] br[222] wl[229] vdd gnd cell_6t
Xbit_r230_c222 bl[222] br[222] wl[230] vdd gnd cell_6t
Xbit_r231_c222 bl[222] br[222] wl[231] vdd gnd cell_6t
Xbit_r232_c222 bl[222] br[222] wl[232] vdd gnd cell_6t
Xbit_r233_c222 bl[222] br[222] wl[233] vdd gnd cell_6t
Xbit_r234_c222 bl[222] br[222] wl[234] vdd gnd cell_6t
Xbit_r235_c222 bl[222] br[222] wl[235] vdd gnd cell_6t
Xbit_r236_c222 bl[222] br[222] wl[236] vdd gnd cell_6t
Xbit_r237_c222 bl[222] br[222] wl[237] vdd gnd cell_6t
Xbit_r238_c222 bl[222] br[222] wl[238] vdd gnd cell_6t
Xbit_r239_c222 bl[222] br[222] wl[239] vdd gnd cell_6t
Xbit_r240_c222 bl[222] br[222] wl[240] vdd gnd cell_6t
Xbit_r241_c222 bl[222] br[222] wl[241] vdd gnd cell_6t
Xbit_r242_c222 bl[222] br[222] wl[242] vdd gnd cell_6t
Xbit_r243_c222 bl[222] br[222] wl[243] vdd gnd cell_6t
Xbit_r244_c222 bl[222] br[222] wl[244] vdd gnd cell_6t
Xbit_r245_c222 bl[222] br[222] wl[245] vdd gnd cell_6t
Xbit_r246_c222 bl[222] br[222] wl[246] vdd gnd cell_6t
Xbit_r247_c222 bl[222] br[222] wl[247] vdd gnd cell_6t
Xbit_r248_c222 bl[222] br[222] wl[248] vdd gnd cell_6t
Xbit_r249_c222 bl[222] br[222] wl[249] vdd gnd cell_6t
Xbit_r250_c222 bl[222] br[222] wl[250] vdd gnd cell_6t
Xbit_r251_c222 bl[222] br[222] wl[251] vdd gnd cell_6t
Xbit_r252_c222 bl[222] br[222] wl[252] vdd gnd cell_6t
Xbit_r253_c222 bl[222] br[222] wl[253] vdd gnd cell_6t
Xbit_r254_c222 bl[222] br[222] wl[254] vdd gnd cell_6t
Xbit_r255_c222 bl[222] br[222] wl[255] vdd gnd cell_6t
Xbit_r0_c223 bl[223] br[223] wl[0] vdd gnd cell_6t
Xbit_r1_c223 bl[223] br[223] wl[1] vdd gnd cell_6t
Xbit_r2_c223 bl[223] br[223] wl[2] vdd gnd cell_6t
Xbit_r3_c223 bl[223] br[223] wl[3] vdd gnd cell_6t
Xbit_r4_c223 bl[223] br[223] wl[4] vdd gnd cell_6t
Xbit_r5_c223 bl[223] br[223] wl[5] vdd gnd cell_6t
Xbit_r6_c223 bl[223] br[223] wl[6] vdd gnd cell_6t
Xbit_r7_c223 bl[223] br[223] wl[7] vdd gnd cell_6t
Xbit_r8_c223 bl[223] br[223] wl[8] vdd gnd cell_6t
Xbit_r9_c223 bl[223] br[223] wl[9] vdd gnd cell_6t
Xbit_r10_c223 bl[223] br[223] wl[10] vdd gnd cell_6t
Xbit_r11_c223 bl[223] br[223] wl[11] vdd gnd cell_6t
Xbit_r12_c223 bl[223] br[223] wl[12] vdd gnd cell_6t
Xbit_r13_c223 bl[223] br[223] wl[13] vdd gnd cell_6t
Xbit_r14_c223 bl[223] br[223] wl[14] vdd gnd cell_6t
Xbit_r15_c223 bl[223] br[223] wl[15] vdd gnd cell_6t
Xbit_r16_c223 bl[223] br[223] wl[16] vdd gnd cell_6t
Xbit_r17_c223 bl[223] br[223] wl[17] vdd gnd cell_6t
Xbit_r18_c223 bl[223] br[223] wl[18] vdd gnd cell_6t
Xbit_r19_c223 bl[223] br[223] wl[19] vdd gnd cell_6t
Xbit_r20_c223 bl[223] br[223] wl[20] vdd gnd cell_6t
Xbit_r21_c223 bl[223] br[223] wl[21] vdd gnd cell_6t
Xbit_r22_c223 bl[223] br[223] wl[22] vdd gnd cell_6t
Xbit_r23_c223 bl[223] br[223] wl[23] vdd gnd cell_6t
Xbit_r24_c223 bl[223] br[223] wl[24] vdd gnd cell_6t
Xbit_r25_c223 bl[223] br[223] wl[25] vdd gnd cell_6t
Xbit_r26_c223 bl[223] br[223] wl[26] vdd gnd cell_6t
Xbit_r27_c223 bl[223] br[223] wl[27] vdd gnd cell_6t
Xbit_r28_c223 bl[223] br[223] wl[28] vdd gnd cell_6t
Xbit_r29_c223 bl[223] br[223] wl[29] vdd gnd cell_6t
Xbit_r30_c223 bl[223] br[223] wl[30] vdd gnd cell_6t
Xbit_r31_c223 bl[223] br[223] wl[31] vdd gnd cell_6t
Xbit_r32_c223 bl[223] br[223] wl[32] vdd gnd cell_6t
Xbit_r33_c223 bl[223] br[223] wl[33] vdd gnd cell_6t
Xbit_r34_c223 bl[223] br[223] wl[34] vdd gnd cell_6t
Xbit_r35_c223 bl[223] br[223] wl[35] vdd gnd cell_6t
Xbit_r36_c223 bl[223] br[223] wl[36] vdd gnd cell_6t
Xbit_r37_c223 bl[223] br[223] wl[37] vdd gnd cell_6t
Xbit_r38_c223 bl[223] br[223] wl[38] vdd gnd cell_6t
Xbit_r39_c223 bl[223] br[223] wl[39] vdd gnd cell_6t
Xbit_r40_c223 bl[223] br[223] wl[40] vdd gnd cell_6t
Xbit_r41_c223 bl[223] br[223] wl[41] vdd gnd cell_6t
Xbit_r42_c223 bl[223] br[223] wl[42] vdd gnd cell_6t
Xbit_r43_c223 bl[223] br[223] wl[43] vdd gnd cell_6t
Xbit_r44_c223 bl[223] br[223] wl[44] vdd gnd cell_6t
Xbit_r45_c223 bl[223] br[223] wl[45] vdd gnd cell_6t
Xbit_r46_c223 bl[223] br[223] wl[46] vdd gnd cell_6t
Xbit_r47_c223 bl[223] br[223] wl[47] vdd gnd cell_6t
Xbit_r48_c223 bl[223] br[223] wl[48] vdd gnd cell_6t
Xbit_r49_c223 bl[223] br[223] wl[49] vdd gnd cell_6t
Xbit_r50_c223 bl[223] br[223] wl[50] vdd gnd cell_6t
Xbit_r51_c223 bl[223] br[223] wl[51] vdd gnd cell_6t
Xbit_r52_c223 bl[223] br[223] wl[52] vdd gnd cell_6t
Xbit_r53_c223 bl[223] br[223] wl[53] vdd gnd cell_6t
Xbit_r54_c223 bl[223] br[223] wl[54] vdd gnd cell_6t
Xbit_r55_c223 bl[223] br[223] wl[55] vdd gnd cell_6t
Xbit_r56_c223 bl[223] br[223] wl[56] vdd gnd cell_6t
Xbit_r57_c223 bl[223] br[223] wl[57] vdd gnd cell_6t
Xbit_r58_c223 bl[223] br[223] wl[58] vdd gnd cell_6t
Xbit_r59_c223 bl[223] br[223] wl[59] vdd gnd cell_6t
Xbit_r60_c223 bl[223] br[223] wl[60] vdd gnd cell_6t
Xbit_r61_c223 bl[223] br[223] wl[61] vdd gnd cell_6t
Xbit_r62_c223 bl[223] br[223] wl[62] vdd gnd cell_6t
Xbit_r63_c223 bl[223] br[223] wl[63] vdd gnd cell_6t
Xbit_r64_c223 bl[223] br[223] wl[64] vdd gnd cell_6t
Xbit_r65_c223 bl[223] br[223] wl[65] vdd gnd cell_6t
Xbit_r66_c223 bl[223] br[223] wl[66] vdd gnd cell_6t
Xbit_r67_c223 bl[223] br[223] wl[67] vdd gnd cell_6t
Xbit_r68_c223 bl[223] br[223] wl[68] vdd gnd cell_6t
Xbit_r69_c223 bl[223] br[223] wl[69] vdd gnd cell_6t
Xbit_r70_c223 bl[223] br[223] wl[70] vdd gnd cell_6t
Xbit_r71_c223 bl[223] br[223] wl[71] vdd gnd cell_6t
Xbit_r72_c223 bl[223] br[223] wl[72] vdd gnd cell_6t
Xbit_r73_c223 bl[223] br[223] wl[73] vdd gnd cell_6t
Xbit_r74_c223 bl[223] br[223] wl[74] vdd gnd cell_6t
Xbit_r75_c223 bl[223] br[223] wl[75] vdd gnd cell_6t
Xbit_r76_c223 bl[223] br[223] wl[76] vdd gnd cell_6t
Xbit_r77_c223 bl[223] br[223] wl[77] vdd gnd cell_6t
Xbit_r78_c223 bl[223] br[223] wl[78] vdd gnd cell_6t
Xbit_r79_c223 bl[223] br[223] wl[79] vdd gnd cell_6t
Xbit_r80_c223 bl[223] br[223] wl[80] vdd gnd cell_6t
Xbit_r81_c223 bl[223] br[223] wl[81] vdd gnd cell_6t
Xbit_r82_c223 bl[223] br[223] wl[82] vdd gnd cell_6t
Xbit_r83_c223 bl[223] br[223] wl[83] vdd gnd cell_6t
Xbit_r84_c223 bl[223] br[223] wl[84] vdd gnd cell_6t
Xbit_r85_c223 bl[223] br[223] wl[85] vdd gnd cell_6t
Xbit_r86_c223 bl[223] br[223] wl[86] vdd gnd cell_6t
Xbit_r87_c223 bl[223] br[223] wl[87] vdd gnd cell_6t
Xbit_r88_c223 bl[223] br[223] wl[88] vdd gnd cell_6t
Xbit_r89_c223 bl[223] br[223] wl[89] vdd gnd cell_6t
Xbit_r90_c223 bl[223] br[223] wl[90] vdd gnd cell_6t
Xbit_r91_c223 bl[223] br[223] wl[91] vdd gnd cell_6t
Xbit_r92_c223 bl[223] br[223] wl[92] vdd gnd cell_6t
Xbit_r93_c223 bl[223] br[223] wl[93] vdd gnd cell_6t
Xbit_r94_c223 bl[223] br[223] wl[94] vdd gnd cell_6t
Xbit_r95_c223 bl[223] br[223] wl[95] vdd gnd cell_6t
Xbit_r96_c223 bl[223] br[223] wl[96] vdd gnd cell_6t
Xbit_r97_c223 bl[223] br[223] wl[97] vdd gnd cell_6t
Xbit_r98_c223 bl[223] br[223] wl[98] vdd gnd cell_6t
Xbit_r99_c223 bl[223] br[223] wl[99] vdd gnd cell_6t
Xbit_r100_c223 bl[223] br[223] wl[100] vdd gnd cell_6t
Xbit_r101_c223 bl[223] br[223] wl[101] vdd gnd cell_6t
Xbit_r102_c223 bl[223] br[223] wl[102] vdd gnd cell_6t
Xbit_r103_c223 bl[223] br[223] wl[103] vdd gnd cell_6t
Xbit_r104_c223 bl[223] br[223] wl[104] vdd gnd cell_6t
Xbit_r105_c223 bl[223] br[223] wl[105] vdd gnd cell_6t
Xbit_r106_c223 bl[223] br[223] wl[106] vdd gnd cell_6t
Xbit_r107_c223 bl[223] br[223] wl[107] vdd gnd cell_6t
Xbit_r108_c223 bl[223] br[223] wl[108] vdd gnd cell_6t
Xbit_r109_c223 bl[223] br[223] wl[109] vdd gnd cell_6t
Xbit_r110_c223 bl[223] br[223] wl[110] vdd gnd cell_6t
Xbit_r111_c223 bl[223] br[223] wl[111] vdd gnd cell_6t
Xbit_r112_c223 bl[223] br[223] wl[112] vdd gnd cell_6t
Xbit_r113_c223 bl[223] br[223] wl[113] vdd gnd cell_6t
Xbit_r114_c223 bl[223] br[223] wl[114] vdd gnd cell_6t
Xbit_r115_c223 bl[223] br[223] wl[115] vdd gnd cell_6t
Xbit_r116_c223 bl[223] br[223] wl[116] vdd gnd cell_6t
Xbit_r117_c223 bl[223] br[223] wl[117] vdd gnd cell_6t
Xbit_r118_c223 bl[223] br[223] wl[118] vdd gnd cell_6t
Xbit_r119_c223 bl[223] br[223] wl[119] vdd gnd cell_6t
Xbit_r120_c223 bl[223] br[223] wl[120] vdd gnd cell_6t
Xbit_r121_c223 bl[223] br[223] wl[121] vdd gnd cell_6t
Xbit_r122_c223 bl[223] br[223] wl[122] vdd gnd cell_6t
Xbit_r123_c223 bl[223] br[223] wl[123] vdd gnd cell_6t
Xbit_r124_c223 bl[223] br[223] wl[124] vdd gnd cell_6t
Xbit_r125_c223 bl[223] br[223] wl[125] vdd gnd cell_6t
Xbit_r126_c223 bl[223] br[223] wl[126] vdd gnd cell_6t
Xbit_r127_c223 bl[223] br[223] wl[127] vdd gnd cell_6t
Xbit_r128_c223 bl[223] br[223] wl[128] vdd gnd cell_6t
Xbit_r129_c223 bl[223] br[223] wl[129] vdd gnd cell_6t
Xbit_r130_c223 bl[223] br[223] wl[130] vdd gnd cell_6t
Xbit_r131_c223 bl[223] br[223] wl[131] vdd gnd cell_6t
Xbit_r132_c223 bl[223] br[223] wl[132] vdd gnd cell_6t
Xbit_r133_c223 bl[223] br[223] wl[133] vdd gnd cell_6t
Xbit_r134_c223 bl[223] br[223] wl[134] vdd gnd cell_6t
Xbit_r135_c223 bl[223] br[223] wl[135] vdd gnd cell_6t
Xbit_r136_c223 bl[223] br[223] wl[136] vdd gnd cell_6t
Xbit_r137_c223 bl[223] br[223] wl[137] vdd gnd cell_6t
Xbit_r138_c223 bl[223] br[223] wl[138] vdd gnd cell_6t
Xbit_r139_c223 bl[223] br[223] wl[139] vdd gnd cell_6t
Xbit_r140_c223 bl[223] br[223] wl[140] vdd gnd cell_6t
Xbit_r141_c223 bl[223] br[223] wl[141] vdd gnd cell_6t
Xbit_r142_c223 bl[223] br[223] wl[142] vdd gnd cell_6t
Xbit_r143_c223 bl[223] br[223] wl[143] vdd gnd cell_6t
Xbit_r144_c223 bl[223] br[223] wl[144] vdd gnd cell_6t
Xbit_r145_c223 bl[223] br[223] wl[145] vdd gnd cell_6t
Xbit_r146_c223 bl[223] br[223] wl[146] vdd gnd cell_6t
Xbit_r147_c223 bl[223] br[223] wl[147] vdd gnd cell_6t
Xbit_r148_c223 bl[223] br[223] wl[148] vdd gnd cell_6t
Xbit_r149_c223 bl[223] br[223] wl[149] vdd gnd cell_6t
Xbit_r150_c223 bl[223] br[223] wl[150] vdd gnd cell_6t
Xbit_r151_c223 bl[223] br[223] wl[151] vdd gnd cell_6t
Xbit_r152_c223 bl[223] br[223] wl[152] vdd gnd cell_6t
Xbit_r153_c223 bl[223] br[223] wl[153] vdd gnd cell_6t
Xbit_r154_c223 bl[223] br[223] wl[154] vdd gnd cell_6t
Xbit_r155_c223 bl[223] br[223] wl[155] vdd gnd cell_6t
Xbit_r156_c223 bl[223] br[223] wl[156] vdd gnd cell_6t
Xbit_r157_c223 bl[223] br[223] wl[157] vdd gnd cell_6t
Xbit_r158_c223 bl[223] br[223] wl[158] vdd gnd cell_6t
Xbit_r159_c223 bl[223] br[223] wl[159] vdd gnd cell_6t
Xbit_r160_c223 bl[223] br[223] wl[160] vdd gnd cell_6t
Xbit_r161_c223 bl[223] br[223] wl[161] vdd gnd cell_6t
Xbit_r162_c223 bl[223] br[223] wl[162] vdd gnd cell_6t
Xbit_r163_c223 bl[223] br[223] wl[163] vdd gnd cell_6t
Xbit_r164_c223 bl[223] br[223] wl[164] vdd gnd cell_6t
Xbit_r165_c223 bl[223] br[223] wl[165] vdd gnd cell_6t
Xbit_r166_c223 bl[223] br[223] wl[166] vdd gnd cell_6t
Xbit_r167_c223 bl[223] br[223] wl[167] vdd gnd cell_6t
Xbit_r168_c223 bl[223] br[223] wl[168] vdd gnd cell_6t
Xbit_r169_c223 bl[223] br[223] wl[169] vdd gnd cell_6t
Xbit_r170_c223 bl[223] br[223] wl[170] vdd gnd cell_6t
Xbit_r171_c223 bl[223] br[223] wl[171] vdd gnd cell_6t
Xbit_r172_c223 bl[223] br[223] wl[172] vdd gnd cell_6t
Xbit_r173_c223 bl[223] br[223] wl[173] vdd gnd cell_6t
Xbit_r174_c223 bl[223] br[223] wl[174] vdd gnd cell_6t
Xbit_r175_c223 bl[223] br[223] wl[175] vdd gnd cell_6t
Xbit_r176_c223 bl[223] br[223] wl[176] vdd gnd cell_6t
Xbit_r177_c223 bl[223] br[223] wl[177] vdd gnd cell_6t
Xbit_r178_c223 bl[223] br[223] wl[178] vdd gnd cell_6t
Xbit_r179_c223 bl[223] br[223] wl[179] vdd gnd cell_6t
Xbit_r180_c223 bl[223] br[223] wl[180] vdd gnd cell_6t
Xbit_r181_c223 bl[223] br[223] wl[181] vdd gnd cell_6t
Xbit_r182_c223 bl[223] br[223] wl[182] vdd gnd cell_6t
Xbit_r183_c223 bl[223] br[223] wl[183] vdd gnd cell_6t
Xbit_r184_c223 bl[223] br[223] wl[184] vdd gnd cell_6t
Xbit_r185_c223 bl[223] br[223] wl[185] vdd gnd cell_6t
Xbit_r186_c223 bl[223] br[223] wl[186] vdd gnd cell_6t
Xbit_r187_c223 bl[223] br[223] wl[187] vdd gnd cell_6t
Xbit_r188_c223 bl[223] br[223] wl[188] vdd gnd cell_6t
Xbit_r189_c223 bl[223] br[223] wl[189] vdd gnd cell_6t
Xbit_r190_c223 bl[223] br[223] wl[190] vdd gnd cell_6t
Xbit_r191_c223 bl[223] br[223] wl[191] vdd gnd cell_6t
Xbit_r192_c223 bl[223] br[223] wl[192] vdd gnd cell_6t
Xbit_r193_c223 bl[223] br[223] wl[193] vdd gnd cell_6t
Xbit_r194_c223 bl[223] br[223] wl[194] vdd gnd cell_6t
Xbit_r195_c223 bl[223] br[223] wl[195] vdd gnd cell_6t
Xbit_r196_c223 bl[223] br[223] wl[196] vdd gnd cell_6t
Xbit_r197_c223 bl[223] br[223] wl[197] vdd gnd cell_6t
Xbit_r198_c223 bl[223] br[223] wl[198] vdd gnd cell_6t
Xbit_r199_c223 bl[223] br[223] wl[199] vdd gnd cell_6t
Xbit_r200_c223 bl[223] br[223] wl[200] vdd gnd cell_6t
Xbit_r201_c223 bl[223] br[223] wl[201] vdd gnd cell_6t
Xbit_r202_c223 bl[223] br[223] wl[202] vdd gnd cell_6t
Xbit_r203_c223 bl[223] br[223] wl[203] vdd gnd cell_6t
Xbit_r204_c223 bl[223] br[223] wl[204] vdd gnd cell_6t
Xbit_r205_c223 bl[223] br[223] wl[205] vdd gnd cell_6t
Xbit_r206_c223 bl[223] br[223] wl[206] vdd gnd cell_6t
Xbit_r207_c223 bl[223] br[223] wl[207] vdd gnd cell_6t
Xbit_r208_c223 bl[223] br[223] wl[208] vdd gnd cell_6t
Xbit_r209_c223 bl[223] br[223] wl[209] vdd gnd cell_6t
Xbit_r210_c223 bl[223] br[223] wl[210] vdd gnd cell_6t
Xbit_r211_c223 bl[223] br[223] wl[211] vdd gnd cell_6t
Xbit_r212_c223 bl[223] br[223] wl[212] vdd gnd cell_6t
Xbit_r213_c223 bl[223] br[223] wl[213] vdd gnd cell_6t
Xbit_r214_c223 bl[223] br[223] wl[214] vdd gnd cell_6t
Xbit_r215_c223 bl[223] br[223] wl[215] vdd gnd cell_6t
Xbit_r216_c223 bl[223] br[223] wl[216] vdd gnd cell_6t
Xbit_r217_c223 bl[223] br[223] wl[217] vdd gnd cell_6t
Xbit_r218_c223 bl[223] br[223] wl[218] vdd gnd cell_6t
Xbit_r219_c223 bl[223] br[223] wl[219] vdd gnd cell_6t
Xbit_r220_c223 bl[223] br[223] wl[220] vdd gnd cell_6t
Xbit_r221_c223 bl[223] br[223] wl[221] vdd gnd cell_6t
Xbit_r222_c223 bl[223] br[223] wl[222] vdd gnd cell_6t
Xbit_r223_c223 bl[223] br[223] wl[223] vdd gnd cell_6t
Xbit_r224_c223 bl[223] br[223] wl[224] vdd gnd cell_6t
Xbit_r225_c223 bl[223] br[223] wl[225] vdd gnd cell_6t
Xbit_r226_c223 bl[223] br[223] wl[226] vdd gnd cell_6t
Xbit_r227_c223 bl[223] br[223] wl[227] vdd gnd cell_6t
Xbit_r228_c223 bl[223] br[223] wl[228] vdd gnd cell_6t
Xbit_r229_c223 bl[223] br[223] wl[229] vdd gnd cell_6t
Xbit_r230_c223 bl[223] br[223] wl[230] vdd gnd cell_6t
Xbit_r231_c223 bl[223] br[223] wl[231] vdd gnd cell_6t
Xbit_r232_c223 bl[223] br[223] wl[232] vdd gnd cell_6t
Xbit_r233_c223 bl[223] br[223] wl[233] vdd gnd cell_6t
Xbit_r234_c223 bl[223] br[223] wl[234] vdd gnd cell_6t
Xbit_r235_c223 bl[223] br[223] wl[235] vdd gnd cell_6t
Xbit_r236_c223 bl[223] br[223] wl[236] vdd gnd cell_6t
Xbit_r237_c223 bl[223] br[223] wl[237] vdd gnd cell_6t
Xbit_r238_c223 bl[223] br[223] wl[238] vdd gnd cell_6t
Xbit_r239_c223 bl[223] br[223] wl[239] vdd gnd cell_6t
Xbit_r240_c223 bl[223] br[223] wl[240] vdd gnd cell_6t
Xbit_r241_c223 bl[223] br[223] wl[241] vdd gnd cell_6t
Xbit_r242_c223 bl[223] br[223] wl[242] vdd gnd cell_6t
Xbit_r243_c223 bl[223] br[223] wl[243] vdd gnd cell_6t
Xbit_r244_c223 bl[223] br[223] wl[244] vdd gnd cell_6t
Xbit_r245_c223 bl[223] br[223] wl[245] vdd gnd cell_6t
Xbit_r246_c223 bl[223] br[223] wl[246] vdd gnd cell_6t
Xbit_r247_c223 bl[223] br[223] wl[247] vdd gnd cell_6t
Xbit_r248_c223 bl[223] br[223] wl[248] vdd gnd cell_6t
Xbit_r249_c223 bl[223] br[223] wl[249] vdd gnd cell_6t
Xbit_r250_c223 bl[223] br[223] wl[250] vdd gnd cell_6t
Xbit_r251_c223 bl[223] br[223] wl[251] vdd gnd cell_6t
Xbit_r252_c223 bl[223] br[223] wl[252] vdd gnd cell_6t
Xbit_r253_c223 bl[223] br[223] wl[253] vdd gnd cell_6t
Xbit_r254_c223 bl[223] br[223] wl[254] vdd gnd cell_6t
Xbit_r255_c223 bl[223] br[223] wl[255] vdd gnd cell_6t
Xbit_r0_c224 bl[224] br[224] wl[0] vdd gnd cell_6t
Xbit_r1_c224 bl[224] br[224] wl[1] vdd gnd cell_6t
Xbit_r2_c224 bl[224] br[224] wl[2] vdd gnd cell_6t
Xbit_r3_c224 bl[224] br[224] wl[3] vdd gnd cell_6t
Xbit_r4_c224 bl[224] br[224] wl[4] vdd gnd cell_6t
Xbit_r5_c224 bl[224] br[224] wl[5] vdd gnd cell_6t
Xbit_r6_c224 bl[224] br[224] wl[6] vdd gnd cell_6t
Xbit_r7_c224 bl[224] br[224] wl[7] vdd gnd cell_6t
Xbit_r8_c224 bl[224] br[224] wl[8] vdd gnd cell_6t
Xbit_r9_c224 bl[224] br[224] wl[9] vdd gnd cell_6t
Xbit_r10_c224 bl[224] br[224] wl[10] vdd gnd cell_6t
Xbit_r11_c224 bl[224] br[224] wl[11] vdd gnd cell_6t
Xbit_r12_c224 bl[224] br[224] wl[12] vdd gnd cell_6t
Xbit_r13_c224 bl[224] br[224] wl[13] vdd gnd cell_6t
Xbit_r14_c224 bl[224] br[224] wl[14] vdd gnd cell_6t
Xbit_r15_c224 bl[224] br[224] wl[15] vdd gnd cell_6t
Xbit_r16_c224 bl[224] br[224] wl[16] vdd gnd cell_6t
Xbit_r17_c224 bl[224] br[224] wl[17] vdd gnd cell_6t
Xbit_r18_c224 bl[224] br[224] wl[18] vdd gnd cell_6t
Xbit_r19_c224 bl[224] br[224] wl[19] vdd gnd cell_6t
Xbit_r20_c224 bl[224] br[224] wl[20] vdd gnd cell_6t
Xbit_r21_c224 bl[224] br[224] wl[21] vdd gnd cell_6t
Xbit_r22_c224 bl[224] br[224] wl[22] vdd gnd cell_6t
Xbit_r23_c224 bl[224] br[224] wl[23] vdd gnd cell_6t
Xbit_r24_c224 bl[224] br[224] wl[24] vdd gnd cell_6t
Xbit_r25_c224 bl[224] br[224] wl[25] vdd gnd cell_6t
Xbit_r26_c224 bl[224] br[224] wl[26] vdd gnd cell_6t
Xbit_r27_c224 bl[224] br[224] wl[27] vdd gnd cell_6t
Xbit_r28_c224 bl[224] br[224] wl[28] vdd gnd cell_6t
Xbit_r29_c224 bl[224] br[224] wl[29] vdd gnd cell_6t
Xbit_r30_c224 bl[224] br[224] wl[30] vdd gnd cell_6t
Xbit_r31_c224 bl[224] br[224] wl[31] vdd gnd cell_6t
Xbit_r32_c224 bl[224] br[224] wl[32] vdd gnd cell_6t
Xbit_r33_c224 bl[224] br[224] wl[33] vdd gnd cell_6t
Xbit_r34_c224 bl[224] br[224] wl[34] vdd gnd cell_6t
Xbit_r35_c224 bl[224] br[224] wl[35] vdd gnd cell_6t
Xbit_r36_c224 bl[224] br[224] wl[36] vdd gnd cell_6t
Xbit_r37_c224 bl[224] br[224] wl[37] vdd gnd cell_6t
Xbit_r38_c224 bl[224] br[224] wl[38] vdd gnd cell_6t
Xbit_r39_c224 bl[224] br[224] wl[39] vdd gnd cell_6t
Xbit_r40_c224 bl[224] br[224] wl[40] vdd gnd cell_6t
Xbit_r41_c224 bl[224] br[224] wl[41] vdd gnd cell_6t
Xbit_r42_c224 bl[224] br[224] wl[42] vdd gnd cell_6t
Xbit_r43_c224 bl[224] br[224] wl[43] vdd gnd cell_6t
Xbit_r44_c224 bl[224] br[224] wl[44] vdd gnd cell_6t
Xbit_r45_c224 bl[224] br[224] wl[45] vdd gnd cell_6t
Xbit_r46_c224 bl[224] br[224] wl[46] vdd gnd cell_6t
Xbit_r47_c224 bl[224] br[224] wl[47] vdd gnd cell_6t
Xbit_r48_c224 bl[224] br[224] wl[48] vdd gnd cell_6t
Xbit_r49_c224 bl[224] br[224] wl[49] vdd gnd cell_6t
Xbit_r50_c224 bl[224] br[224] wl[50] vdd gnd cell_6t
Xbit_r51_c224 bl[224] br[224] wl[51] vdd gnd cell_6t
Xbit_r52_c224 bl[224] br[224] wl[52] vdd gnd cell_6t
Xbit_r53_c224 bl[224] br[224] wl[53] vdd gnd cell_6t
Xbit_r54_c224 bl[224] br[224] wl[54] vdd gnd cell_6t
Xbit_r55_c224 bl[224] br[224] wl[55] vdd gnd cell_6t
Xbit_r56_c224 bl[224] br[224] wl[56] vdd gnd cell_6t
Xbit_r57_c224 bl[224] br[224] wl[57] vdd gnd cell_6t
Xbit_r58_c224 bl[224] br[224] wl[58] vdd gnd cell_6t
Xbit_r59_c224 bl[224] br[224] wl[59] vdd gnd cell_6t
Xbit_r60_c224 bl[224] br[224] wl[60] vdd gnd cell_6t
Xbit_r61_c224 bl[224] br[224] wl[61] vdd gnd cell_6t
Xbit_r62_c224 bl[224] br[224] wl[62] vdd gnd cell_6t
Xbit_r63_c224 bl[224] br[224] wl[63] vdd gnd cell_6t
Xbit_r64_c224 bl[224] br[224] wl[64] vdd gnd cell_6t
Xbit_r65_c224 bl[224] br[224] wl[65] vdd gnd cell_6t
Xbit_r66_c224 bl[224] br[224] wl[66] vdd gnd cell_6t
Xbit_r67_c224 bl[224] br[224] wl[67] vdd gnd cell_6t
Xbit_r68_c224 bl[224] br[224] wl[68] vdd gnd cell_6t
Xbit_r69_c224 bl[224] br[224] wl[69] vdd gnd cell_6t
Xbit_r70_c224 bl[224] br[224] wl[70] vdd gnd cell_6t
Xbit_r71_c224 bl[224] br[224] wl[71] vdd gnd cell_6t
Xbit_r72_c224 bl[224] br[224] wl[72] vdd gnd cell_6t
Xbit_r73_c224 bl[224] br[224] wl[73] vdd gnd cell_6t
Xbit_r74_c224 bl[224] br[224] wl[74] vdd gnd cell_6t
Xbit_r75_c224 bl[224] br[224] wl[75] vdd gnd cell_6t
Xbit_r76_c224 bl[224] br[224] wl[76] vdd gnd cell_6t
Xbit_r77_c224 bl[224] br[224] wl[77] vdd gnd cell_6t
Xbit_r78_c224 bl[224] br[224] wl[78] vdd gnd cell_6t
Xbit_r79_c224 bl[224] br[224] wl[79] vdd gnd cell_6t
Xbit_r80_c224 bl[224] br[224] wl[80] vdd gnd cell_6t
Xbit_r81_c224 bl[224] br[224] wl[81] vdd gnd cell_6t
Xbit_r82_c224 bl[224] br[224] wl[82] vdd gnd cell_6t
Xbit_r83_c224 bl[224] br[224] wl[83] vdd gnd cell_6t
Xbit_r84_c224 bl[224] br[224] wl[84] vdd gnd cell_6t
Xbit_r85_c224 bl[224] br[224] wl[85] vdd gnd cell_6t
Xbit_r86_c224 bl[224] br[224] wl[86] vdd gnd cell_6t
Xbit_r87_c224 bl[224] br[224] wl[87] vdd gnd cell_6t
Xbit_r88_c224 bl[224] br[224] wl[88] vdd gnd cell_6t
Xbit_r89_c224 bl[224] br[224] wl[89] vdd gnd cell_6t
Xbit_r90_c224 bl[224] br[224] wl[90] vdd gnd cell_6t
Xbit_r91_c224 bl[224] br[224] wl[91] vdd gnd cell_6t
Xbit_r92_c224 bl[224] br[224] wl[92] vdd gnd cell_6t
Xbit_r93_c224 bl[224] br[224] wl[93] vdd gnd cell_6t
Xbit_r94_c224 bl[224] br[224] wl[94] vdd gnd cell_6t
Xbit_r95_c224 bl[224] br[224] wl[95] vdd gnd cell_6t
Xbit_r96_c224 bl[224] br[224] wl[96] vdd gnd cell_6t
Xbit_r97_c224 bl[224] br[224] wl[97] vdd gnd cell_6t
Xbit_r98_c224 bl[224] br[224] wl[98] vdd gnd cell_6t
Xbit_r99_c224 bl[224] br[224] wl[99] vdd gnd cell_6t
Xbit_r100_c224 bl[224] br[224] wl[100] vdd gnd cell_6t
Xbit_r101_c224 bl[224] br[224] wl[101] vdd gnd cell_6t
Xbit_r102_c224 bl[224] br[224] wl[102] vdd gnd cell_6t
Xbit_r103_c224 bl[224] br[224] wl[103] vdd gnd cell_6t
Xbit_r104_c224 bl[224] br[224] wl[104] vdd gnd cell_6t
Xbit_r105_c224 bl[224] br[224] wl[105] vdd gnd cell_6t
Xbit_r106_c224 bl[224] br[224] wl[106] vdd gnd cell_6t
Xbit_r107_c224 bl[224] br[224] wl[107] vdd gnd cell_6t
Xbit_r108_c224 bl[224] br[224] wl[108] vdd gnd cell_6t
Xbit_r109_c224 bl[224] br[224] wl[109] vdd gnd cell_6t
Xbit_r110_c224 bl[224] br[224] wl[110] vdd gnd cell_6t
Xbit_r111_c224 bl[224] br[224] wl[111] vdd gnd cell_6t
Xbit_r112_c224 bl[224] br[224] wl[112] vdd gnd cell_6t
Xbit_r113_c224 bl[224] br[224] wl[113] vdd gnd cell_6t
Xbit_r114_c224 bl[224] br[224] wl[114] vdd gnd cell_6t
Xbit_r115_c224 bl[224] br[224] wl[115] vdd gnd cell_6t
Xbit_r116_c224 bl[224] br[224] wl[116] vdd gnd cell_6t
Xbit_r117_c224 bl[224] br[224] wl[117] vdd gnd cell_6t
Xbit_r118_c224 bl[224] br[224] wl[118] vdd gnd cell_6t
Xbit_r119_c224 bl[224] br[224] wl[119] vdd gnd cell_6t
Xbit_r120_c224 bl[224] br[224] wl[120] vdd gnd cell_6t
Xbit_r121_c224 bl[224] br[224] wl[121] vdd gnd cell_6t
Xbit_r122_c224 bl[224] br[224] wl[122] vdd gnd cell_6t
Xbit_r123_c224 bl[224] br[224] wl[123] vdd gnd cell_6t
Xbit_r124_c224 bl[224] br[224] wl[124] vdd gnd cell_6t
Xbit_r125_c224 bl[224] br[224] wl[125] vdd gnd cell_6t
Xbit_r126_c224 bl[224] br[224] wl[126] vdd gnd cell_6t
Xbit_r127_c224 bl[224] br[224] wl[127] vdd gnd cell_6t
Xbit_r128_c224 bl[224] br[224] wl[128] vdd gnd cell_6t
Xbit_r129_c224 bl[224] br[224] wl[129] vdd gnd cell_6t
Xbit_r130_c224 bl[224] br[224] wl[130] vdd gnd cell_6t
Xbit_r131_c224 bl[224] br[224] wl[131] vdd gnd cell_6t
Xbit_r132_c224 bl[224] br[224] wl[132] vdd gnd cell_6t
Xbit_r133_c224 bl[224] br[224] wl[133] vdd gnd cell_6t
Xbit_r134_c224 bl[224] br[224] wl[134] vdd gnd cell_6t
Xbit_r135_c224 bl[224] br[224] wl[135] vdd gnd cell_6t
Xbit_r136_c224 bl[224] br[224] wl[136] vdd gnd cell_6t
Xbit_r137_c224 bl[224] br[224] wl[137] vdd gnd cell_6t
Xbit_r138_c224 bl[224] br[224] wl[138] vdd gnd cell_6t
Xbit_r139_c224 bl[224] br[224] wl[139] vdd gnd cell_6t
Xbit_r140_c224 bl[224] br[224] wl[140] vdd gnd cell_6t
Xbit_r141_c224 bl[224] br[224] wl[141] vdd gnd cell_6t
Xbit_r142_c224 bl[224] br[224] wl[142] vdd gnd cell_6t
Xbit_r143_c224 bl[224] br[224] wl[143] vdd gnd cell_6t
Xbit_r144_c224 bl[224] br[224] wl[144] vdd gnd cell_6t
Xbit_r145_c224 bl[224] br[224] wl[145] vdd gnd cell_6t
Xbit_r146_c224 bl[224] br[224] wl[146] vdd gnd cell_6t
Xbit_r147_c224 bl[224] br[224] wl[147] vdd gnd cell_6t
Xbit_r148_c224 bl[224] br[224] wl[148] vdd gnd cell_6t
Xbit_r149_c224 bl[224] br[224] wl[149] vdd gnd cell_6t
Xbit_r150_c224 bl[224] br[224] wl[150] vdd gnd cell_6t
Xbit_r151_c224 bl[224] br[224] wl[151] vdd gnd cell_6t
Xbit_r152_c224 bl[224] br[224] wl[152] vdd gnd cell_6t
Xbit_r153_c224 bl[224] br[224] wl[153] vdd gnd cell_6t
Xbit_r154_c224 bl[224] br[224] wl[154] vdd gnd cell_6t
Xbit_r155_c224 bl[224] br[224] wl[155] vdd gnd cell_6t
Xbit_r156_c224 bl[224] br[224] wl[156] vdd gnd cell_6t
Xbit_r157_c224 bl[224] br[224] wl[157] vdd gnd cell_6t
Xbit_r158_c224 bl[224] br[224] wl[158] vdd gnd cell_6t
Xbit_r159_c224 bl[224] br[224] wl[159] vdd gnd cell_6t
Xbit_r160_c224 bl[224] br[224] wl[160] vdd gnd cell_6t
Xbit_r161_c224 bl[224] br[224] wl[161] vdd gnd cell_6t
Xbit_r162_c224 bl[224] br[224] wl[162] vdd gnd cell_6t
Xbit_r163_c224 bl[224] br[224] wl[163] vdd gnd cell_6t
Xbit_r164_c224 bl[224] br[224] wl[164] vdd gnd cell_6t
Xbit_r165_c224 bl[224] br[224] wl[165] vdd gnd cell_6t
Xbit_r166_c224 bl[224] br[224] wl[166] vdd gnd cell_6t
Xbit_r167_c224 bl[224] br[224] wl[167] vdd gnd cell_6t
Xbit_r168_c224 bl[224] br[224] wl[168] vdd gnd cell_6t
Xbit_r169_c224 bl[224] br[224] wl[169] vdd gnd cell_6t
Xbit_r170_c224 bl[224] br[224] wl[170] vdd gnd cell_6t
Xbit_r171_c224 bl[224] br[224] wl[171] vdd gnd cell_6t
Xbit_r172_c224 bl[224] br[224] wl[172] vdd gnd cell_6t
Xbit_r173_c224 bl[224] br[224] wl[173] vdd gnd cell_6t
Xbit_r174_c224 bl[224] br[224] wl[174] vdd gnd cell_6t
Xbit_r175_c224 bl[224] br[224] wl[175] vdd gnd cell_6t
Xbit_r176_c224 bl[224] br[224] wl[176] vdd gnd cell_6t
Xbit_r177_c224 bl[224] br[224] wl[177] vdd gnd cell_6t
Xbit_r178_c224 bl[224] br[224] wl[178] vdd gnd cell_6t
Xbit_r179_c224 bl[224] br[224] wl[179] vdd gnd cell_6t
Xbit_r180_c224 bl[224] br[224] wl[180] vdd gnd cell_6t
Xbit_r181_c224 bl[224] br[224] wl[181] vdd gnd cell_6t
Xbit_r182_c224 bl[224] br[224] wl[182] vdd gnd cell_6t
Xbit_r183_c224 bl[224] br[224] wl[183] vdd gnd cell_6t
Xbit_r184_c224 bl[224] br[224] wl[184] vdd gnd cell_6t
Xbit_r185_c224 bl[224] br[224] wl[185] vdd gnd cell_6t
Xbit_r186_c224 bl[224] br[224] wl[186] vdd gnd cell_6t
Xbit_r187_c224 bl[224] br[224] wl[187] vdd gnd cell_6t
Xbit_r188_c224 bl[224] br[224] wl[188] vdd gnd cell_6t
Xbit_r189_c224 bl[224] br[224] wl[189] vdd gnd cell_6t
Xbit_r190_c224 bl[224] br[224] wl[190] vdd gnd cell_6t
Xbit_r191_c224 bl[224] br[224] wl[191] vdd gnd cell_6t
Xbit_r192_c224 bl[224] br[224] wl[192] vdd gnd cell_6t
Xbit_r193_c224 bl[224] br[224] wl[193] vdd gnd cell_6t
Xbit_r194_c224 bl[224] br[224] wl[194] vdd gnd cell_6t
Xbit_r195_c224 bl[224] br[224] wl[195] vdd gnd cell_6t
Xbit_r196_c224 bl[224] br[224] wl[196] vdd gnd cell_6t
Xbit_r197_c224 bl[224] br[224] wl[197] vdd gnd cell_6t
Xbit_r198_c224 bl[224] br[224] wl[198] vdd gnd cell_6t
Xbit_r199_c224 bl[224] br[224] wl[199] vdd gnd cell_6t
Xbit_r200_c224 bl[224] br[224] wl[200] vdd gnd cell_6t
Xbit_r201_c224 bl[224] br[224] wl[201] vdd gnd cell_6t
Xbit_r202_c224 bl[224] br[224] wl[202] vdd gnd cell_6t
Xbit_r203_c224 bl[224] br[224] wl[203] vdd gnd cell_6t
Xbit_r204_c224 bl[224] br[224] wl[204] vdd gnd cell_6t
Xbit_r205_c224 bl[224] br[224] wl[205] vdd gnd cell_6t
Xbit_r206_c224 bl[224] br[224] wl[206] vdd gnd cell_6t
Xbit_r207_c224 bl[224] br[224] wl[207] vdd gnd cell_6t
Xbit_r208_c224 bl[224] br[224] wl[208] vdd gnd cell_6t
Xbit_r209_c224 bl[224] br[224] wl[209] vdd gnd cell_6t
Xbit_r210_c224 bl[224] br[224] wl[210] vdd gnd cell_6t
Xbit_r211_c224 bl[224] br[224] wl[211] vdd gnd cell_6t
Xbit_r212_c224 bl[224] br[224] wl[212] vdd gnd cell_6t
Xbit_r213_c224 bl[224] br[224] wl[213] vdd gnd cell_6t
Xbit_r214_c224 bl[224] br[224] wl[214] vdd gnd cell_6t
Xbit_r215_c224 bl[224] br[224] wl[215] vdd gnd cell_6t
Xbit_r216_c224 bl[224] br[224] wl[216] vdd gnd cell_6t
Xbit_r217_c224 bl[224] br[224] wl[217] vdd gnd cell_6t
Xbit_r218_c224 bl[224] br[224] wl[218] vdd gnd cell_6t
Xbit_r219_c224 bl[224] br[224] wl[219] vdd gnd cell_6t
Xbit_r220_c224 bl[224] br[224] wl[220] vdd gnd cell_6t
Xbit_r221_c224 bl[224] br[224] wl[221] vdd gnd cell_6t
Xbit_r222_c224 bl[224] br[224] wl[222] vdd gnd cell_6t
Xbit_r223_c224 bl[224] br[224] wl[223] vdd gnd cell_6t
Xbit_r224_c224 bl[224] br[224] wl[224] vdd gnd cell_6t
Xbit_r225_c224 bl[224] br[224] wl[225] vdd gnd cell_6t
Xbit_r226_c224 bl[224] br[224] wl[226] vdd gnd cell_6t
Xbit_r227_c224 bl[224] br[224] wl[227] vdd gnd cell_6t
Xbit_r228_c224 bl[224] br[224] wl[228] vdd gnd cell_6t
Xbit_r229_c224 bl[224] br[224] wl[229] vdd gnd cell_6t
Xbit_r230_c224 bl[224] br[224] wl[230] vdd gnd cell_6t
Xbit_r231_c224 bl[224] br[224] wl[231] vdd gnd cell_6t
Xbit_r232_c224 bl[224] br[224] wl[232] vdd gnd cell_6t
Xbit_r233_c224 bl[224] br[224] wl[233] vdd gnd cell_6t
Xbit_r234_c224 bl[224] br[224] wl[234] vdd gnd cell_6t
Xbit_r235_c224 bl[224] br[224] wl[235] vdd gnd cell_6t
Xbit_r236_c224 bl[224] br[224] wl[236] vdd gnd cell_6t
Xbit_r237_c224 bl[224] br[224] wl[237] vdd gnd cell_6t
Xbit_r238_c224 bl[224] br[224] wl[238] vdd gnd cell_6t
Xbit_r239_c224 bl[224] br[224] wl[239] vdd gnd cell_6t
Xbit_r240_c224 bl[224] br[224] wl[240] vdd gnd cell_6t
Xbit_r241_c224 bl[224] br[224] wl[241] vdd gnd cell_6t
Xbit_r242_c224 bl[224] br[224] wl[242] vdd gnd cell_6t
Xbit_r243_c224 bl[224] br[224] wl[243] vdd gnd cell_6t
Xbit_r244_c224 bl[224] br[224] wl[244] vdd gnd cell_6t
Xbit_r245_c224 bl[224] br[224] wl[245] vdd gnd cell_6t
Xbit_r246_c224 bl[224] br[224] wl[246] vdd gnd cell_6t
Xbit_r247_c224 bl[224] br[224] wl[247] vdd gnd cell_6t
Xbit_r248_c224 bl[224] br[224] wl[248] vdd gnd cell_6t
Xbit_r249_c224 bl[224] br[224] wl[249] vdd gnd cell_6t
Xbit_r250_c224 bl[224] br[224] wl[250] vdd gnd cell_6t
Xbit_r251_c224 bl[224] br[224] wl[251] vdd gnd cell_6t
Xbit_r252_c224 bl[224] br[224] wl[252] vdd gnd cell_6t
Xbit_r253_c224 bl[224] br[224] wl[253] vdd gnd cell_6t
Xbit_r254_c224 bl[224] br[224] wl[254] vdd gnd cell_6t
Xbit_r255_c224 bl[224] br[224] wl[255] vdd gnd cell_6t
Xbit_r0_c225 bl[225] br[225] wl[0] vdd gnd cell_6t
Xbit_r1_c225 bl[225] br[225] wl[1] vdd gnd cell_6t
Xbit_r2_c225 bl[225] br[225] wl[2] vdd gnd cell_6t
Xbit_r3_c225 bl[225] br[225] wl[3] vdd gnd cell_6t
Xbit_r4_c225 bl[225] br[225] wl[4] vdd gnd cell_6t
Xbit_r5_c225 bl[225] br[225] wl[5] vdd gnd cell_6t
Xbit_r6_c225 bl[225] br[225] wl[6] vdd gnd cell_6t
Xbit_r7_c225 bl[225] br[225] wl[7] vdd gnd cell_6t
Xbit_r8_c225 bl[225] br[225] wl[8] vdd gnd cell_6t
Xbit_r9_c225 bl[225] br[225] wl[9] vdd gnd cell_6t
Xbit_r10_c225 bl[225] br[225] wl[10] vdd gnd cell_6t
Xbit_r11_c225 bl[225] br[225] wl[11] vdd gnd cell_6t
Xbit_r12_c225 bl[225] br[225] wl[12] vdd gnd cell_6t
Xbit_r13_c225 bl[225] br[225] wl[13] vdd gnd cell_6t
Xbit_r14_c225 bl[225] br[225] wl[14] vdd gnd cell_6t
Xbit_r15_c225 bl[225] br[225] wl[15] vdd gnd cell_6t
Xbit_r16_c225 bl[225] br[225] wl[16] vdd gnd cell_6t
Xbit_r17_c225 bl[225] br[225] wl[17] vdd gnd cell_6t
Xbit_r18_c225 bl[225] br[225] wl[18] vdd gnd cell_6t
Xbit_r19_c225 bl[225] br[225] wl[19] vdd gnd cell_6t
Xbit_r20_c225 bl[225] br[225] wl[20] vdd gnd cell_6t
Xbit_r21_c225 bl[225] br[225] wl[21] vdd gnd cell_6t
Xbit_r22_c225 bl[225] br[225] wl[22] vdd gnd cell_6t
Xbit_r23_c225 bl[225] br[225] wl[23] vdd gnd cell_6t
Xbit_r24_c225 bl[225] br[225] wl[24] vdd gnd cell_6t
Xbit_r25_c225 bl[225] br[225] wl[25] vdd gnd cell_6t
Xbit_r26_c225 bl[225] br[225] wl[26] vdd gnd cell_6t
Xbit_r27_c225 bl[225] br[225] wl[27] vdd gnd cell_6t
Xbit_r28_c225 bl[225] br[225] wl[28] vdd gnd cell_6t
Xbit_r29_c225 bl[225] br[225] wl[29] vdd gnd cell_6t
Xbit_r30_c225 bl[225] br[225] wl[30] vdd gnd cell_6t
Xbit_r31_c225 bl[225] br[225] wl[31] vdd gnd cell_6t
Xbit_r32_c225 bl[225] br[225] wl[32] vdd gnd cell_6t
Xbit_r33_c225 bl[225] br[225] wl[33] vdd gnd cell_6t
Xbit_r34_c225 bl[225] br[225] wl[34] vdd gnd cell_6t
Xbit_r35_c225 bl[225] br[225] wl[35] vdd gnd cell_6t
Xbit_r36_c225 bl[225] br[225] wl[36] vdd gnd cell_6t
Xbit_r37_c225 bl[225] br[225] wl[37] vdd gnd cell_6t
Xbit_r38_c225 bl[225] br[225] wl[38] vdd gnd cell_6t
Xbit_r39_c225 bl[225] br[225] wl[39] vdd gnd cell_6t
Xbit_r40_c225 bl[225] br[225] wl[40] vdd gnd cell_6t
Xbit_r41_c225 bl[225] br[225] wl[41] vdd gnd cell_6t
Xbit_r42_c225 bl[225] br[225] wl[42] vdd gnd cell_6t
Xbit_r43_c225 bl[225] br[225] wl[43] vdd gnd cell_6t
Xbit_r44_c225 bl[225] br[225] wl[44] vdd gnd cell_6t
Xbit_r45_c225 bl[225] br[225] wl[45] vdd gnd cell_6t
Xbit_r46_c225 bl[225] br[225] wl[46] vdd gnd cell_6t
Xbit_r47_c225 bl[225] br[225] wl[47] vdd gnd cell_6t
Xbit_r48_c225 bl[225] br[225] wl[48] vdd gnd cell_6t
Xbit_r49_c225 bl[225] br[225] wl[49] vdd gnd cell_6t
Xbit_r50_c225 bl[225] br[225] wl[50] vdd gnd cell_6t
Xbit_r51_c225 bl[225] br[225] wl[51] vdd gnd cell_6t
Xbit_r52_c225 bl[225] br[225] wl[52] vdd gnd cell_6t
Xbit_r53_c225 bl[225] br[225] wl[53] vdd gnd cell_6t
Xbit_r54_c225 bl[225] br[225] wl[54] vdd gnd cell_6t
Xbit_r55_c225 bl[225] br[225] wl[55] vdd gnd cell_6t
Xbit_r56_c225 bl[225] br[225] wl[56] vdd gnd cell_6t
Xbit_r57_c225 bl[225] br[225] wl[57] vdd gnd cell_6t
Xbit_r58_c225 bl[225] br[225] wl[58] vdd gnd cell_6t
Xbit_r59_c225 bl[225] br[225] wl[59] vdd gnd cell_6t
Xbit_r60_c225 bl[225] br[225] wl[60] vdd gnd cell_6t
Xbit_r61_c225 bl[225] br[225] wl[61] vdd gnd cell_6t
Xbit_r62_c225 bl[225] br[225] wl[62] vdd gnd cell_6t
Xbit_r63_c225 bl[225] br[225] wl[63] vdd gnd cell_6t
Xbit_r64_c225 bl[225] br[225] wl[64] vdd gnd cell_6t
Xbit_r65_c225 bl[225] br[225] wl[65] vdd gnd cell_6t
Xbit_r66_c225 bl[225] br[225] wl[66] vdd gnd cell_6t
Xbit_r67_c225 bl[225] br[225] wl[67] vdd gnd cell_6t
Xbit_r68_c225 bl[225] br[225] wl[68] vdd gnd cell_6t
Xbit_r69_c225 bl[225] br[225] wl[69] vdd gnd cell_6t
Xbit_r70_c225 bl[225] br[225] wl[70] vdd gnd cell_6t
Xbit_r71_c225 bl[225] br[225] wl[71] vdd gnd cell_6t
Xbit_r72_c225 bl[225] br[225] wl[72] vdd gnd cell_6t
Xbit_r73_c225 bl[225] br[225] wl[73] vdd gnd cell_6t
Xbit_r74_c225 bl[225] br[225] wl[74] vdd gnd cell_6t
Xbit_r75_c225 bl[225] br[225] wl[75] vdd gnd cell_6t
Xbit_r76_c225 bl[225] br[225] wl[76] vdd gnd cell_6t
Xbit_r77_c225 bl[225] br[225] wl[77] vdd gnd cell_6t
Xbit_r78_c225 bl[225] br[225] wl[78] vdd gnd cell_6t
Xbit_r79_c225 bl[225] br[225] wl[79] vdd gnd cell_6t
Xbit_r80_c225 bl[225] br[225] wl[80] vdd gnd cell_6t
Xbit_r81_c225 bl[225] br[225] wl[81] vdd gnd cell_6t
Xbit_r82_c225 bl[225] br[225] wl[82] vdd gnd cell_6t
Xbit_r83_c225 bl[225] br[225] wl[83] vdd gnd cell_6t
Xbit_r84_c225 bl[225] br[225] wl[84] vdd gnd cell_6t
Xbit_r85_c225 bl[225] br[225] wl[85] vdd gnd cell_6t
Xbit_r86_c225 bl[225] br[225] wl[86] vdd gnd cell_6t
Xbit_r87_c225 bl[225] br[225] wl[87] vdd gnd cell_6t
Xbit_r88_c225 bl[225] br[225] wl[88] vdd gnd cell_6t
Xbit_r89_c225 bl[225] br[225] wl[89] vdd gnd cell_6t
Xbit_r90_c225 bl[225] br[225] wl[90] vdd gnd cell_6t
Xbit_r91_c225 bl[225] br[225] wl[91] vdd gnd cell_6t
Xbit_r92_c225 bl[225] br[225] wl[92] vdd gnd cell_6t
Xbit_r93_c225 bl[225] br[225] wl[93] vdd gnd cell_6t
Xbit_r94_c225 bl[225] br[225] wl[94] vdd gnd cell_6t
Xbit_r95_c225 bl[225] br[225] wl[95] vdd gnd cell_6t
Xbit_r96_c225 bl[225] br[225] wl[96] vdd gnd cell_6t
Xbit_r97_c225 bl[225] br[225] wl[97] vdd gnd cell_6t
Xbit_r98_c225 bl[225] br[225] wl[98] vdd gnd cell_6t
Xbit_r99_c225 bl[225] br[225] wl[99] vdd gnd cell_6t
Xbit_r100_c225 bl[225] br[225] wl[100] vdd gnd cell_6t
Xbit_r101_c225 bl[225] br[225] wl[101] vdd gnd cell_6t
Xbit_r102_c225 bl[225] br[225] wl[102] vdd gnd cell_6t
Xbit_r103_c225 bl[225] br[225] wl[103] vdd gnd cell_6t
Xbit_r104_c225 bl[225] br[225] wl[104] vdd gnd cell_6t
Xbit_r105_c225 bl[225] br[225] wl[105] vdd gnd cell_6t
Xbit_r106_c225 bl[225] br[225] wl[106] vdd gnd cell_6t
Xbit_r107_c225 bl[225] br[225] wl[107] vdd gnd cell_6t
Xbit_r108_c225 bl[225] br[225] wl[108] vdd gnd cell_6t
Xbit_r109_c225 bl[225] br[225] wl[109] vdd gnd cell_6t
Xbit_r110_c225 bl[225] br[225] wl[110] vdd gnd cell_6t
Xbit_r111_c225 bl[225] br[225] wl[111] vdd gnd cell_6t
Xbit_r112_c225 bl[225] br[225] wl[112] vdd gnd cell_6t
Xbit_r113_c225 bl[225] br[225] wl[113] vdd gnd cell_6t
Xbit_r114_c225 bl[225] br[225] wl[114] vdd gnd cell_6t
Xbit_r115_c225 bl[225] br[225] wl[115] vdd gnd cell_6t
Xbit_r116_c225 bl[225] br[225] wl[116] vdd gnd cell_6t
Xbit_r117_c225 bl[225] br[225] wl[117] vdd gnd cell_6t
Xbit_r118_c225 bl[225] br[225] wl[118] vdd gnd cell_6t
Xbit_r119_c225 bl[225] br[225] wl[119] vdd gnd cell_6t
Xbit_r120_c225 bl[225] br[225] wl[120] vdd gnd cell_6t
Xbit_r121_c225 bl[225] br[225] wl[121] vdd gnd cell_6t
Xbit_r122_c225 bl[225] br[225] wl[122] vdd gnd cell_6t
Xbit_r123_c225 bl[225] br[225] wl[123] vdd gnd cell_6t
Xbit_r124_c225 bl[225] br[225] wl[124] vdd gnd cell_6t
Xbit_r125_c225 bl[225] br[225] wl[125] vdd gnd cell_6t
Xbit_r126_c225 bl[225] br[225] wl[126] vdd gnd cell_6t
Xbit_r127_c225 bl[225] br[225] wl[127] vdd gnd cell_6t
Xbit_r128_c225 bl[225] br[225] wl[128] vdd gnd cell_6t
Xbit_r129_c225 bl[225] br[225] wl[129] vdd gnd cell_6t
Xbit_r130_c225 bl[225] br[225] wl[130] vdd gnd cell_6t
Xbit_r131_c225 bl[225] br[225] wl[131] vdd gnd cell_6t
Xbit_r132_c225 bl[225] br[225] wl[132] vdd gnd cell_6t
Xbit_r133_c225 bl[225] br[225] wl[133] vdd gnd cell_6t
Xbit_r134_c225 bl[225] br[225] wl[134] vdd gnd cell_6t
Xbit_r135_c225 bl[225] br[225] wl[135] vdd gnd cell_6t
Xbit_r136_c225 bl[225] br[225] wl[136] vdd gnd cell_6t
Xbit_r137_c225 bl[225] br[225] wl[137] vdd gnd cell_6t
Xbit_r138_c225 bl[225] br[225] wl[138] vdd gnd cell_6t
Xbit_r139_c225 bl[225] br[225] wl[139] vdd gnd cell_6t
Xbit_r140_c225 bl[225] br[225] wl[140] vdd gnd cell_6t
Xbit_r141_c225 bl[225] br[225] wl[141] vdd gnd cell_6t
Xbit_r142_c225 bl[225] br[225] wl[142] vdd gnd cell_6t
Xbit_r143_c225 bl[225] br[225] wl[143] vdd gnd cell_6t
Xbit_r144_c225 bl[225] br[225] wl[144] vdd gnd cell_6t
Xbit_r145_c225 bl[225] br[225] wl[145] vdd gnd cell_6t
Xbit_r146_c225 bl[225] br[225] wl[146] vdd gnd cell_6t
Xbit_r147_c225 bl[225] br[225] wl[147] vdd gnd cell_6t
Xbit_r148_c225 bl[225] br[225] wl[148] vdd gnd cell_6t
Xbit_r149_c225 bl[225] br[225] wl[149] vdd gnd cell_6t
Xbit_r150_c225 bl[225] br[225] wl[150] vdd gnd cell_6t
Xbit_r151_c225 bl[225] br[225] wl[151] vdd gnd cell_6t
Xbit_r152_c225 bl[225] br[225] wl[152] vdd gnd cell_6t
Xbit_r153_c225 bl[225] br[225] wl[153] vdd gnd cell_6t
Xbit_r154_c225 bl[225] br[225] wl[154] vdd gnd cell_6t
Xbit_r155_c225 bl[225] br[225] wl[155] vdd gnd cell_6t
Xbit_r156_c225 bl[225] br[225] wl[156] vdd gnd cell_6t
Xbit_r157_c225 bl[225] br[225] wl[157] vdd gnd cell_6t
Xbit_r158_c225 bl[225] br[225] wl[158] vdd gnd cell_6t
Xbit_r159_c225 bl[225] br[225] wl[159] vdd gnd cell_6t
Xbit_r160_c225 bl[225] br[225] wl[160] vdd gnd cell_6t
Xbit_r161_c225 bl[225] br[225] wl[161] vdd gnd cell_6t
Xbit_r162_c225 bl[225] br[225] wl[162] vdd gnd cell_6t
Xbit_r163_c225 bl[225] br[225] wl[163] vdd gnd cell_6t
Xbit_r164_c225 bl[225] br[225] wl[164] vdd gnd cell_6t
Xbit_r165_c225 bl[225] br[225] wl[165] vdd gnd cell_6t
Xbit_r166_c225 bl[225] br[225] wl[166] vdd gnd cell_6t
Xbit_r167_c225 bl[225] br[225] wl[167] vdd gnd cell_6t
Xbit_r168_c225 bl[225] br[225] wl[168] vdd gnd cell_6t
Xbit_r169_c225 bl[225] br[225] wl[169] vdd gnd cell_6t
Xbit_r170_c225 bl[225] br[225] wl[170] vdd gnd cell_6t
Xbit_r171_c225 bl[225] br[225] wl[171] vdd gnd cell_6t
Xbit_r172_c225 bl[225] br[225] wl[172] vdd gnd cell_6t
Xbit_r173_c225 bl[225] br[225] wl[173] vdd gnd cell_6t
Xbit_r174_c225 bl[225] br[225] wl[174] vdd gnd cell_6t
Xbit_r175_c225 bl[225] br[225] wl[175] vdd gnd cell_6t
Xbit_r176_c225 bl[225] br[225] wl[176] vdd gnd cell_6t
Xbit_r177_c225 bl[225] br[225] wl[177] vdd gnd cell_6t
Xbit_r178_c225 bl[225] br[225] wl[178] vdd gnd cell_6t
Xbit_r179_c225 bl[225] br[225] wl[179] vdd gnd cell_6t
Xbit_r180_c225 bl[225] br[225] wl[180] vdd gnd cell_6t
Xbit_r181_c225 bl[225] br[225] wl[181] vdd gnd cell_6t
Xbit_r182_c225 bl[225] br[225] wl[182] vdd gnd cell_6t
Xbit_r183_c225 bl[225] br[225] wl[183] vdd gnd cell_6t
Xbit_r184_c225 bl[225] br[225] wl[184] vdd gnd cell_6t
Xbit_r185_c225 bl[225] br[225] wl[185] vdd gnd cell_6t
Xbit_r186_c225 bl[225] br[225] wl[186] vdd gnd cell_6t
Xbit_r187_c225 bl[225] br[225] wl[187] vdd gnd cell_6t
Xbit_r188_c225 bl[225] br[225] wl[188] vdd gnd cell_6t
Xbit_r189_c225 bl[225] br[225] wl[189] vdd gnd cell_6t
Xbit_r190_c225 bl[225] br[225] wl[190] vdd gnd cell_6t
Xbit_r191_c225 bl[225] br[225] wl[191] vdd gnd cell_6t
Xbit_r192_c225 bl[225] br[225] wl[192] vdd gnd cell_6t
Xbit_r193_c225 bl[225] br[225] wl[193] vdd gnd cell_6t
Xbit_r194_c225 bl[225] br[225] wl[194] vdd gnd cell_6t
Xbit_r195_c225 bl[225] br[225] wl[195] vdd gnd cell_6t
Xbit_r196_c225 bl[225] br[225] wl[196] vdd gnd cell_6t
Xbit_r197_c225 bl[225] br[225] wl[197] vdd gnd cell_6t
Xbit_r198_c225 bl[225] br[225] wl[198] vdd gnd cell_6t
Xbit_r199_c225 bl[225] br[225] wl[199] vdd gnd cell_6t
Xbit_r200_c225 bl[225] br[225] wl[200] vdd gnd cell_6t
Xbit_r201_c225 bl[225] br[225] wl[201] vdd gnd cell_6t
Xbit_r202_c225 bl[225] br[225] wl[202] vdd gnd cell_6t
Xbit_r203_c225 bl[225] br[225] wl[203] vdd gnd cell_6t
Xbit_r204_c225 bl[225] br[225] wl[204] vdd gnd cell_6t
Xbit_r205_c225 bl[225] br[225] wl[205] vdd gnd cell_6t
Xbit_r206_c225 bl[225] br[225] wl[206] vdd gnd cell_6t
Xbit_r207_c225 bl[225] br[225] wl[207] vdd gnd cell_6t
Xbit_r208_c225 bl[225] br[225] wl[208] vdd gnd cell_6t
Xbit_r209_c225 bl[225] br[225] wl[209] vdd gnd cell_6t
Xbit_r210_c225 bl[225] br[225] wl[210] vdd gnd cell_6t
Xbit_r211_c225 bl[225] br[225] wl[211] vdd gnd cell_6t
Xbit_r212_c225 bl[225] br[225] wl[212] vdd gnd cell_6t
Xbit_r213_c225 bl[225] br[225] wl[213] vdd gnd cell_6t
Xbit_r214_c225 bl[225] br[225] wl[214] vdd gnd cell_6t
Xbit_r215_c225 bl[225] br[225] wl[215] vdd gnd cell_6t
Xbit_r216_c225 bl[225] br[225] wl[216] vdd gnd cell_6t
Xbit_r217_c225 bl[225] br[225] wl[217] vdd gnd cell_6t
Xbit_r218_c225 bl[225] br[225] wl[218] vdd gnd cell_6t
Xbit_r219_c225 bl[225] br[225] wl[219] vdd gnd cell_6t
Xbit_r220_c225 bl[225] br[225] wl[220] vdd gnd cell_6t
Xbit_r221_c225 bl[225] br[225] wl[221] vdd gnd cell_6t
Xbit_r222_c225 bl[225] br[225] wl[222] vdd gnd cell_6t
Xbit_r223_c225 bl[225] br[225] wl[223] vdd gnd cell_6t
Xbit_r224_c225 bl[225] br[225] wl[224] vdd gnd cell_6t
Xbit_r225_c225 bl[225] br[225] wl[225] vdd gnd cell_6t
Xbit_r226_c225 bl[225] br[225] wl[226] vdd gnd cell_6t
Xbit_r227_c225 bl[225] br[225] wl[227] vdd gnd cell_6t
Xbit_r228_c225 bl[225] br[225] wl[228] vdd gnd cell_6t
Xbit_r229_c225 bl[225] br[225] wl[229] vdd gnd cell_6t
Xbit_r230_c225 bl[225] br[225] wl[230] vdd gnd cell_6t
Xbit_r231_c225 bl[225] br[225] wl[231] vdd gnd cell_6t
Xbit_r232_c225 bl[225] br[225] wl[232] vdd gnd cell_6t
Xbit_r233_c225 bl[225] br[225] wl[233] vdd gnd cell_6t
Xbit_r234_c225 bl[225] br[225] wl[234] vdd gnd cell_6t
Xbit_r235_c225 bl[225] br[225] wl[235] vdd gnd cell_6t
Xbit_r236_c225 bl[225] br[225] wl[236] vdd gnd cell_6t
Xbit_r237_c225 bl[225] br[225] wl[237] vdd gnd cell_6t
Xbit_r238_c225 bl[225] br[225] wl[238] vdd gnd cell_6t
Xbit_r239_c225 bl[225] br[225] wl[239] vdd gnd cell_6t
Xbit_r240_c225 bl[225] br[225] wl[240] vdd gnd cell_6t
Xbit_r241_c225 bl[225] br[225] wl[241] vdd gnd cell_6t
Xbit_r242_c225 bl[225] br[225] wl[242] vdd gnd cell_6t
Xbit_r243_c225 bl[225] br[225] wl[243] vdd gnd cell_6t
Xbit_r244_c225 bl[225] br[225] wl[244] vdd gnd cell_6t
Xbit_r245_c225 bl[225] br[225] wl[245] vdd gnd cell_6t
Xbit_r246_c225 bl[225] br[225] wl[246] vdd gnd cell_6t
Xbit_r247_c225 bl[225] br[225] wl[247] vdd gnd cell_6t
Xbit_r248_c225 bl[225] br[225] wl[248] vdd gnd cell_6t
Xbit_r249_c225 bl[225] br[225] wl[249] vdd gnd cell_6t
Xbit_r250_c225 bl[225] br[225] wl[250] vdd gnd cell_6t
Xbit_r251_c225 bl[225] br[225] wl[251] vdd gnd cell_6t
Xbit_r252_c225 bl[225] br[225] wl[252] vdd gnd cell_6t
Xbit_r253_c225 bl[225] br[225] wl[253] vdd gnd cell_6t
Xbit_r254_c225 bl[225] br[225] wl[254] vdd gnd cell_6t
Xbit_r255_c225 bl[225] br[225] wl[255] vdd gnd cell_6t
Xbit_r0_c226 bl[226] br[226] wl[0] vdd gnd cell_6t
Xbit_r1_c226 bl[226] br[226] wl[1] vdd gnd cell_6t
Xbit_r2_c226 bl[226] br[226] wl[2] vdd gnd cell_6t
Xbit_r3_c226 bl[226] br[226] wl[3] vdd gnd cell_6t
Xbit_r4_c226 bl[226] br[226] wl[4] vdd gnd cell_6t
Xbit_r5_c226 bl[226] br[226] wl[5] vdd gnd cell_6t
Xbit_r6_c226 bl[226] br[226] wl[6] vdd gnd cell_6t
Xbit_r7_c226 bl[226] br[226] wl[7] vdd gnd cell_6t
Xbit_r8_c226 bl[226] br[226] wl[8] vdd gnd cell_6t
Xbit_r9_c226 bl[226] br[226] wl[9] vdd gnd cell_6t
Xbit_r10_c226 bl[226] br[226] wl[10] vdd gnd cell_6t
Xbit_r11_c226 bl[226] br[226] wl[11] vdd gnd cell_6t
Xbit_r12_c226 bl[226] br[226] wl[12] vdd gnd cell_6t
Xbit_r13_c226 bl[226] br[226] wl[13] vdd gnd cell_6t
Xbit_r14_c226 bl[226] br[226] wl[14] vdd gnd cell_6t
Xbit_r15_c226 bl[226] br[226] wl[15] vdd gnd cell_6t
Xbit_r16_c226 bl[226] br[226] wl[16] vdd gnd cell_6t
Xbit_r17_c226 bl[226] br[226] wl[17] vdd gnd cell_6t
Xbit_r18_c226 bl[226] br[226] wl[18] vdd gnd cell_6t
Xbit_r19_c226 bl[226] br[226] wl[19] vdd gnd cell_6t
Xbit_r20_c226 bl[226] br[226] wl[20] vdd gnd cell_6t
Xbit_r21_c226 bl[226] br[226] wl[21] vdd gnd cell_6t
Xbit_r22_c226 bl[226] br[226] wl[22] vdd gnd cell_6t
Xbit_r23_c226 bl[226] br[226] wl[23] vdd gnd cell_6t
Xbit_r24_c226 bl[226] br[226] wl[24] vdd gnd cell_6t
Xbit_r25_c226 bl[226] br[226] wl[25] vdd gnd cell_6t
Xbit_r26_c226 bl[226] br[226] wl[26] vdd gnd cell_6t
Xbit_r27_c226 bl[226] br[226] wl[27] vdd gnd cell_6t
Xbit_r28_c226 bl[226] br[226] wl[28] vdd gnd cell_6t
Xbit_r29_c226 bl[226] br[226] wl[29] vdd gnd cell_6t
Xbit_r30_c226 bl[226] br[226] wl[30] vdd gnd cell_6t
Xbit_r31_c226 bl[226] br[226] wl[31] vdd gnd cell_6t
Xbit_r32_c226 bl[226] br[226] wl[32] vdd gnd cell_6t
Xbit_r33_c226 bl[226] br[226] wl[33] vdd gnd cell_6t
Xbit_r34_c226 bl[226] br[226] wl[34] vdd gnd cell_6t
Xbit_r35_c226 bl[226] br[226] wl[35] vdd gnd cell_6t
Xbit_r36_c226 bl[226] br[226] wl[36] vdd gnd cell_6t
Xbit_r37_c226 bl[226] br[226] wl[37] vdd gnd cell_6t
Xbit_r38_c226 bl[226] br[226] wl[38] vdd gnd cell_6t
Xbit_r39_c226 bl[226] br[226] wl[39] vdd gnd cell_6t
Xbit_r40_c226 bl[226] br[226] wl[40] vdd gnd cell_6t
Xbit_r41_c226 bl[226] br[226] wl[41] vdd gnd cell_6t
Xbit_r42_c226 bl[226] br[226] wl[42] vdd gnd cell_6t
Xbit_r43_c226 bl[226] br[226] wl[43] vdd gnd cell_6t
Xbit_r44_c226 bl[226] br[226] wl[44] vdd gnd cell_6t
Xbit_r45_c226 bl[226] br[226] wl[45] vdd gnd cell_6t
Xbit_r46_c226 bl[226] br[226] wl[46] vdd gnd cell_6t
Xbit_r47_c226 bl[226] br[226] wl[47] vdd gnd cell_6t
Xbit_r48_c226 bl[226] br[226] wl[48] vdd gnd cell_6t
Xbit_r49_c226 bl[226] br[226] wl[49] vdd gnd cell_6t
Xbit_r50_c226 bl[226] br[226] wl[50] vdd gnd cell_6t
Xbit_r51_c226 bl[226] br[226] wl[51] vdd gnd cell_6t
Xbit_r52_c226 bl[226] br[226] wl[52] vdd gnd cell_6t
Xbit_r53_c226 bl[226] br[226] wl[53] vdd gnd cell_6t
Xbit_r54_c226 bl[226] br[226] wl[54] vdd gnd cell_6t
Xbit_r55_c226 bl[226] br[226] wl[55] vdd gnd cell_6t
Xbit_r56_c226 bl[226] br[226] wl[56] vdd gnd cell_6t
Xbit_r57_c226 bl[226] br[226] wl[57] vdd gnd cell_6t
Xbit_r58_c226 bl[226] br[226] wl[58] vdd gnd cell_6t
Xbit_r59_c226 bl[226] br[226] wl[59] vdd gnd cell_6t
Xbit_r60_c226 bl[226] br[226] wl[60] vdd gnd cell_6t
Xbit_r61_c226 bl[226] br[226] wl[61] vdd gnd cell_6t
Xbit_r62_c226 bl[226] br[226] wl[62] vdd gnd cell_6t
Xbit_r63_c226 bl[226] br[226] wl[63] vdd gnd cell_6t
Xbit_r64_c226 bl[226] br[226] wl[64] vdd gnd cell_6t
Xbit_r65_c226 bl[226] br[226] wl[65] vdd gnd cell_6t
Xbit_r66_c226 bl[226] br[226] wl[66] vdd gnd cell_6t
Xbit_r67_c226 bl[226] br[226] wl[67] vdd gnd cell_6t
Xbit_r68_c226 bl[226] br[226] wl[68] vdd gnd cell_6t
Xbit_r69_c226 bl[226] br[226] wl[69] vdd gnd cell_6t
Xbit_r70_c226 bl[226] br[226] wl[70] vdd gnd cell_6t
Xbit_r71_c226 bl[226] br[226] wl[71] vdd gnd cell_6t
Xbit_r72_c226 bl[226] br[226] wl[72] vdd gnd cell_6t
Xbit_r73_c226 bl[226] br[226] wl[73] vdd gnd cell_6t
Xbit_r74_c226 bl[226] br[226] wl[74] vdd gnd cell_6t
Xbit_r75_c226 bl[226] br[226] wl[75] vdd gnd cell_6t
Xbit_r76_c226 bl[226] br[226] wl[76] vdd gnd cell_6t
Xbit_r77_c226 bl[226] br[226] wl[77] vdd gnd cell_6t
Xbit_r78_c226 bl[226] br[226] wl[78] vdd gnd cell_6t
Xbit_r79_c226 bl[226] br[226] wl[79] vdd gnd cell_6t
Xbit_r80_c226 bl[226] br[226] wl[80] vdd gnd cell_6t
Xbit_r81_c226 bl[226] br[226] wl[81] vdd gnd cell_6t
Xbit_r82_c226 bl[226] br[226] wl[82] vdd gnd cell_6t
Xbit_r83_c226 bl[226] br[226] wl[83] vdd gnd cell_6t
Xbit_r84_c226 bl[226] br[226] wl[84] vdd gnd cell_6t
Xbit_r85_c226 bl[226] br[226] wl[85] vdd gnd cell_6t
Xbit_r86_c226 bl[226] br[226] wl[86] vdd gnd cell_6t
Xbit_r87_c226 bl[226] br[226] wl[87] vdd gnd cell_6t
Xbit_r88_c226 bl[226] br[226] wl[88] vdd gnd cell_6t
Xbit_r89_c226 bl[226] br[226] wl[89] vdd gnd cell_6t
Xbit_r90_c226 bl[226] br[226] wl[90] vdd gnd cell_6t
Xbit_r91_c226 bl[226] br[226] wl[91] vdd gnd cell_6t
Xbit_r92_c226 bl[226] br[226] wl[92] vdd gnd cell_6t
Xbit_r93_c226 bl[226] br[226] wl[93] vdd gnd cell_6t
Xbit_r94_c226 bl[226] br[226] wl[94] vdd gnd cell_6t
Xbit_r95_c226 bl[226] br[226] wl[95] vdd gnd cell_6t
Xbit_r96_c226 bl[226] br[226] wl[96] vdd gnd cell_6t
Xbit_r97_c226 bl[226] br[226] wl[97] vdd gnd cell_6t
Xbit_r98_c226 bl[226] br[226] wl[98] vdd gnd cell_6t
Xbit_r99_c226 bl[226] br[226] wl[99] vdd gnd cell_6t
Xbit_r100_c226 bl[226] br[226] wl[100] vdd gnd cell_6t
Xbit_r101_c226 bl[226] br[226] wl[101] vdd gnd cell_6t
Xbit_r102_c226 bl[226] br[226] wl[102] vdd gnd cell_6t
Xbit_r103_c226 bl[226] br[226] wl[103] vdd gnd cell_6t
Xbit_r104_c226 bl[226] br[226] wl[104] vdd gnd cell_6t
Xbit_r105_c226 bl[226] br[226] wl[105] vdd gnd cell_6t
Xbit_r106_c226 bl[226] br[226] wl[106] vdd gnd cell_6t
Xbit_r107_c226 bl[226] br[226] wl[107] vdd gnd cell_6t
Xbit_r108_c226 bl[226] br[226] wl[108] vdd gnd cell_6t
Xbit_r109_c226 bl[226] br[226] wl[109] vdd gnd cell_6t
Xbit_r110_c226 bl[226] br[226] wl[110] vdd gnd cell_6t
Xbit_r111_c226 bl[226] br[226] wl[111] vdd gnd cell_6t
Xbit_r112_c226 bl[226] br[226] wl[112] vdd gnd cell_6t
Xbit_r113_c226 bl[226] br[226] wl[113] vdd gnd cell_6t
Xbit_r114_c226 bl[226] br[226] wl[114] vdd gnd cell_6t
Xbit_r115_c226 bl[226] br[226] wl[115] vdd gnd cell_6t
Xbit_r116_c226 bl[226] br[226] wl[116] vdd gnd cell_6t
Xbit_r117_c226 bl[226] br[226] wl[117] vdd gnd cell_6t
Xbit_r118_c226 bl[226] br[226] wl[118] vdd gnd cell_6t
Xbit_r119_c226 bl[226] br[226] wl[119] vdd gnd cell_6t
Xbit_r120_c226 bl[226] br[226] wl[120] vdd gnd cell_6t
Xbit_r121_c226 bl[226] br[226] wl[121] vdd gnd cell_6t
Xbit_r122_c226 bl[226] br[226] wl[122] vdd gnd cell_6t
Xbit_r123_c226 bl[226] br[226] wl[123] vdd gnd cell_6t
Xbit_r124_c226 bl[226] br[226] wl[124] vdd gnd cell_6t
Xbit_r125_c226 bl[226] br[226] wl[125] vdd gnd cell_6t
Xbit_r126_c226 bl[226] br[226] wl[126] vdd gnd cell_6t
Xbit_r127_c226 bl[226] br[226] wl[127] vdd gnd cell_6t
Xbit_r128_c226 bl[226] br[226] wl[128] vdd gnd cell_6t
Xbit_r129_c226 bl[226] br[226] wl[129] vdd gnd cell_6t
Xbit_r130_c226 bl[226] br[226] wl[130] vdd gnd cell_6t
Xbit_r131_c226 bl[226] br[226] wl[131] vdd gnd cell_6t
Xbit_r132_c226 bl[226] br[226] wl[132] vdd gnd cell_6t
Xbit_r133_c226 bl[226] br[226] wl[133] vdd gnd cell_6t
Xbit_r134_c226 bl[226] br[226] wl[134] vdd gnd cell_6t
Xbit_r135_c226 bl[226] br[226] wl[135] vdd gnd cell_6t
Xbit_r136_c226 bl[226] br[226] wl[136] vdd gnd cell_6t
Xbit_r137_c226 bl[226] br[226] wl[137] vdd gnd cell_6t
Xbit_r138_c226 bl[226] br[226] wl[138] vdd gnd cell_6t
Xbit_r139_c226 bl[226] br[226] wl[139] vdd gnd cell_6t
Xbit_r140_c226 bl[226] br[226] wl[140] vdd gnd cell_6t
Xbit_r141_c226 bl[226] br[226] wl[141] vdd gnd cell_6t
Xbit_r142_c226 bl[226] br[226] wl[142] vdd gnd cell_6t
Xbit_r143_c226 bl[226] br[226] wl[143] vdd gnd cell_6t
Xbit_r144_c226 bl[226] br[226] wl[144] vdd gnd cell_6t
Xbit_r145_c226 bl[226] br[226] wl[145] vdd gnd cell_6t
Xbit_r146_c226 bl[226] br[226] wl[146] vdd gnd cell_6t
Xbit_r147_c226 bl[226] br[226] wl[147] vdd gnd cell_6t
Xbit_r148_c226 bl[226] br[226] wl[148] vdd gnd cell_6t
Xbit_r149_c226 bl[226] br[226] wl[149] vdd gnd cell_6t
Xbit_r150_c226 bl[226] br[226] wl[150] vdd gnd cell_6t
Xbit_r151_c226 bl[226] br[226] wl[151] vdd gnd cell_6t
Xbit_r152_c226 bl[226] br[226] wl[152] vdd gnd cell_6t
Xbit_r153_c226 bl[226] br[226] wl[153] vdd gnd cell_6t
Xbit_r154_c226 bl[226] br[226] wl[154] vdd gnd cell_6t
Xbit_r155_c226 bl[226] br[226] wl[155] vdd gnd cell_6t
Xbit_r156_c226 bl[226] br[226] wl[156] vdd gnd cell_6t
Xbit_r157_c226 bl[226] br[226] wl[157] vdd gnd cell_6t
Xbit_r158_c226 bl[226] br[226] wl[158] vdd gnd cell_6t
Xbit_r159_c226 bl[226] br[226] wl[159] vdd gnd cell_6t
Xbit_r160_c226 bl[226] br[226] wl[160] vdd gnd cell_6t
Xbit_r161_c226 bl[226] br[226] wl[161] vdd gnd cell_6t
Xbit_r162_c226 bl[226] br[226] wl[162] vdd gnd cell_6t
Xbit_r163_c226 bl[226] br[226] wl[163] vdd gnd cell_6t
Xbit_r164_c226 bl[226] br[226] wl[164] vdd gnd cell_6t
Xbit_r165_c226 bl[226] br[226] wl[165] vdd gnd cell_6t
Xbit_r166_c226 bl[226] br[226] wl[166] vdd gnd cell_6t
Xbit_r167_c226 bl[226] br[226] wl[167] vdd gnd cell_6t
Xbit_r168_c226 bl[226] br[226] wl[168] vdd gnd cell_6t
Xbit_r169_c226 bl[226] br[226] wl[169] vdd gnd cell_6t
Xbit_r170_c226 bl[226] br[226] wl[170] vdd gnd cell_6t
Xbit_r171_c226 bl[226] br[226] wl[171] vdd gnd cell_6t
Xbit_r172_c226 bl[226] br[226] wl[172] vdd gnd cell_6t
Xbit_r173_c226 bl[226] br[226] wl[173] vdd gnd cell_6t
Xbit_r174_c226 bl[226] br[226] wl[174] vdd gnd cell_6t
Xbit_r175_c226 bl[226] br[226] wl[175] vdd gnd cell_6t
Xbit_r176_c226 bl[226] br[226] wl[176] vdd gnd cell_6t
Xbit_r177_c226 bl[226] br[226] wl[177] vdd gnd cell_6t
Xbit_r178_c226 bl[226] br[226] wl[178] vdd gnd cell_6t
Xbit_r179_c226 bl[226] br[226] wl[179] vdd gnd cell_6t
Xbit_r180_c226 bl[226] br[226] wl[180] vdd gnd cell_6t
Xbit_r181_c226 bl[226] br[226] wl[181] vdd gnd cell_6t
Xbit_r182_c226 bl[226] br[226] wl[182] vdd gnd cell_6t
Xbit_r183_c226 bl[226] br[226] wl[183] vdd gnd cell_6t
Xbit_r184_c226 bl[226] br[226] wl[184] vdd gnd cell_6t
Xbit_r185_c226 bl[226] br[226] wl[185] vdd gnd cell_6t
Xbit_r186_c226 bl[226] br[226] wl[186] vdd gnd cell_6t
Xbit_r187_c226 bl[226] br[226] wl[187] vdd gnd cell_6t
Xbit_r188_c226 bl[226] br[226] wl[188] vdd gnd cell_6t
Xbit_r189_c226 bl[226] br[226] wl[189] vdd gnd cell_6t
Xbit_r190_c226 bl[226] br[226] wl[190] vdd gnd cell_6t
Xbit_r191_c226 bl[226] br[226] wl[191] vdd gnd cell_6t
Xbit_r192_c226 bl[226] br[226] wl[192] vdd gnd cell_6t
Xbit_r193_c226 bl[226] br[226] wl[193] vdd gnd cell_6t
Xbit_r194_c226 bl[226] br[226] wl[194] vdd gnd cell_6t
Xbit_r195_c226 bl[226] br[226] wl[195] vdd gnd cell_6t
Xbit_r196_c226 bl[226] br[226] wl[196] vdd gnd cell_6t
Xbit_r197_c226 bl[226] br[226] wl[197] vdd gnd cell_6t
Xbit_r198_c226 bl[226] br[226] wl[198] vdd gnd cell_6t
Xbit_r199_c226 bl[226] br[226] wl[199] vdd gnd cell_6t
Xbit_r200_c226 bl[226] br[226] wl[200] vdd gnd cell_6t
Xbit_r201_c226 bl[226] br[226] wl[201] vdd gnd cell_6t
Xbit_r202_c226 bl[226] br[226] wl[202] vdd gnd cell_6t
Xbit_r203_c226 bl[226] br[226] wl[203] vdd gnd cell_6t
Xbit_r204_c226 bl[226] br[226] wl[204] vdd gnd cell_6t
Xbit_r205_c226 bl[226] br[226] wl[205] vdd gnd cell_6t
Xbit_r206_c226 bl[226] br[226] wl[206] vdd gnd cell_6t
Xbit_r207_c226 bl[226] br[226] wl[207] vdd gnd cell_6t
Xbit_r208_c226 bl[226] br[226] wl[208] vdd gnd cell_6t
Xbit_r209_c226 bl[226] br[226] wl[209] vdd gnd cell_6t
Xbit_r210_c226 bl[226] br[226] wl[210] vdd gnd cell_6t
Xbit_r211_c226 bl[226] br[226] wl[211] vdd gnd cell_6t
Xbit_r212_c226 bl[226] br[226] wl[212] vdd gnd cell_6t
Xbit_r213_c226 bl[226] br[226] wl[213] vdd gnd cell_6t
Xbit_r214_c226 bl[226] br[226] wl[214] vdd gnd cell_6t
Xbit_r215_c226 bl[226] br[226] wl[215] vdd gnd cell_6t
Xbit_r216_c226 bl[226] br[226] wl[216] vdd gnd cell_6t
Xbit_r217_c226 bl[226] br[226] wl[217] vdd gnd cell_6t
Xbit_r218_c226 bl[226] br[226] wl[218] vdd gnd cell_6t
Xbit_r219_c226 bl[226] br[226] wl[219] vdd gnd cell_6t
Xbit_r220_c226 bl[226] br[226] wl[220] vdd gnd cell_6t
Xbit_r221_c226 bl[226] br[226] wl[221] vdd gnd cell_6t
Xbit_r222_c226 bl[226] br[226] wl[222] vdd gnd cell_6t
Xbit_r223_c226 bl[226] br[226] wl[223] vdd gnd cell_6t
Xbit_r224_c226 bl[226] br[226] wl[224] vdd gnd cell_6t
Xbit_r225_c226 bl[226] br[226] wl[225] vdd gnd cell_6t
Xbit_r226_c226 bl[226] br[226] wl[226] vdd gnd cell_6t
Xbit_r227_c226 bl[226] br[226] wl[227] vdd gnd cell_6t
Xbit_r228_c226 bl[226] br[226] wl[228] vdd gnd cell_6t
Xbit_r229_c226 bl[226] br[226] wl[229] vdd gnd cell_6t
Xbit_r230_c226 bl[226] br[226] wl[230] vdd gnd cell_6t
Xbit_r231_c226 bl[226] br[226] wl[231] vdd gnd cell_6t
Xbit_r232_c226 bl[226] br[226] wl[232] vdd gnd cell_6t
Xbit_r233_c226 bl[226] br[226] wl[233] vdd gnd cell_6t
Xbit_r234_c226 bl[226] br[226] wl[234] vdd gnd cell_6t
Xbit_r235_c226 bl[226] br[226] wl[235] vdd gnd cell_6t
Xbit_r236_c226 bl[226] br[226] wl[236] vdd gnd cell_6t
Xbit_r237_c226 bl[226] br[226] wl[237] vdd gnd cell_6t
Xbit_r238_c226 bl[226] br[226] wl[238] vdd gnd cell_6t
Xbit_r239_c226 bl[226] br[226] wl[239] vdd gnd cell_6t
Xbit_r240_c226 bl[226] br[226] wl[240] vdd gnd cell_6t
Xbit_r241_c226 bl[226] br[226] wl[241] vdd gnd cell_6t
Xbit_r242_c226 bl[226] br[226] wl[242] vdd gnd cell_6t
Xbit_r243_c226 bl[226] br[226] wl[243] vdd gnd cell_6t
Xbit_r244_c226 bl[226] br[226] wl[244] vdd gnd cell_6t
Xbit_r245_c226 bl[226] br[226] wl[245] vdd gnd cell_6t
Xbit_r246_c226 bl[226] br[226] wl[246] vdd gnd cell_6t
Xbit_r247_c226 bl[226] br[226] wl[247] vdd gnd cell_6t
Xbit_r248_c226 bl[226] br[226] wl[248] vdd gnd cell_6t
Xbit_r249_c226 bl[226] br[226] wl[249] vdd gnd cell_6t
Xbit_r250_c226 bl[226] br[226] wl[250] vdd gnd cell_6t
Xbit_r251_c226 bl[226] br[226] wl[251] vdd gnd cell_6t
Xbit_r252_c226 bl[226] br[226] wl[252] vdd gnd cell_6t
Xbit_r253_c226 bl[226] br[226] wl[253] vdd gnd cell_6t
Xbit_r254_c226 bl[226] br[226] wl[254] vdd gnd cell_6t
Xbit_r255_c226 bl[226] br[226] wl[255] vdd gnd cell_6t
Xbit_r0_c227 bl[227] br[227] wl[0] vdd gnd cell_6t
Xbit_r1_c227 bl[227] br[227] wl[1] vdd gnd cell_6t
Xbit_r2_c227 bl[227] br[227] wl[2] vdd gnd cell_6t
Xbit_r3_c227 bl[227] br[227] wl[3] vdd gnd cell_6t
Xbit_r4_c227 bl[227] br[227] wl[4] vdd gnd cell_6t
Xbit_r5_c227 bl[227] br[227] wl[5] vdd gnd cell_6t
Xbit_r6_c227 bl[227] br[227] wl[6] vdd gnd cell_6t
Xbit_r7_c227 bl[227] br[227] wl[7] vdd gnd cell_6t
Xbit_r8_c227 bl[227] br[227] wl[8] vdd gnd cell_6t
Xbit_r9_c227 bl[227] br[227] wl[9] vdd gnd cell_6t
Xbit_r10_c227 bl[227] br[227] wl[10] vdd gnd cell_6t
Xbit_r11_c227 bl[227] br[227] wl[11] vdd gnd cell_6t
Xbit_r12_c227 bl[227] br[227] wl[12] vdd gnd cell_6t
Xbit_r13_c227 bl[227] br[227] wl[13] vdd gnd cell_6t
Xbit_r14_c227 bl[227] br[227] wl[14] vdd gnd cell_6t
Xbit_r15_c227 bl[227] br[227] wl[15] vdd gnd cell_6t
Xbit_r16_c227 bl[227] br[227] wl[16] vdd gnd cell_6t
Xbit_r17_c227 bl[227] br[227] wl[17] vdd gnd cell_6t
Xbit_r18_c227 bl[227] br[227] wl[18] vdd gnd cell_6t
Xbit_r19_c227 bl[227] br[227] wl[19] vdd gnd cell_6t
Xbit_r20_c227 bl[227] br[227] wl[20] vdd gnd cell_6t
Xbit_r21_c227 bl[227] br[227] wl[21] vdd gnd cell_6t
Xbit_r22_c227 bl[227] br[227] wl[22] vdd gnd cell_6t
Xbit_r23_c227 bl[227] br[227] wl[23] vdd gnd cell_6t
Xbit_r24_c227 bl[227] br[227] wl[24] vdd gnd cell_6t
Xbit_r25_c227 bl[227] br[227] wl[25] vdd gnd cell_6t
Xbit_r26_c227 bl[227] br[227] wl[26] vdd gnd cell_6t
Xbit_r27_c227 bl[227] br[227] wl[27] vdd gnd cell_6t
Xbit_r28_c227 bl[227] br[227] wl[28] vdd gnd cell_6t
Xbit_r29_c227 bl[227] br[227] wl[29] vdd gnd cell_6t
Xbit_r30_c227 bl[227] br[227] wl[30] vdd gnd cell_6t
Xbit_r31_c227 bl[227] br[227] wl[31] vdd gnd cell_6t
Xbit_r32_c227 bl[227] br[227] wl[32] vdd gnd cell_6t
Xbit_r33_c227 bl[227] br[227] wl[33] vdd gnd cell_6t
Xbit_r34_c227 bl[227] br[227] wl[34] vdd gnd cell_6t
Xbit_r35_c227 bl[227] br[227] wl[35] vdd gnd cell_6t
Xbit_r36_c227 bl[227] br[227] wl[36] vdd gnd cell_6t
Xbit_r37_c227 bl[227] br[227] wl[37] vdd gnd cell_6t
Xbit_r38_c227 bl[227] br[227] wl[38] vdd gnd cell_6t
Xbit_r39_c227 bl[227] br[227] wl[39] vdd gnd cell_6t
Xbit_r40_c227 bl[227] br[227] wl[40] vdd gnd cell_6t
Xbit_r41_c227 bl[227] br[227] wl[41] vdd gnd cell_6t
Xbit_r42_c227 bl[227] br[227] wl[42] vdd gnd cell_6t
Xbit_r43_c227 bl[227] br[227] wl[43] vdd gnd cell_6t
Xbit_r44_c227 bl[227] br[227] wl[44] vdd gnd cell_6t
Xbit_r45_c227 bl[227] br[227] wl[45] vdd gnd cell_6t
Xbit_r46_c227 bl[227] br[227] wl[46] vdd gnd cell_6t
Xbit_r47_c227 bl[227] br[227] wl[47] vdd gnd cell_6t
Xbit_r48_c227 bl[227] br[227] wl[48] vdd gnd cell_6t
Xbit_r49_c227 bl[227] br[227] wl[49] vdd gnd cell_6t
Xbit_r50_c227 bl[227] br[227] wl[50] vdd gnd cell_6t
Xbit_r51_c227 bl[227] br[227] wl[51] vdd gnd cell_6t
Xbit_r52_c227 bl[227] br[227] wl[52] vdd gnd cell_6t
Xbit_r53_c227 bl[227] br[227] wl[53] vdd gnd cell_6t
Xbit_r54_c227 bl[227] br[227] wl[54] vdd gnd cell_6t
Xbit_r55_c227 bl[227] br[227] wl[55] vdd gnd cell_6t
Xbit_r56_c227 bl[227] br[227] wl[56] vdd gnd cell_6t
Xbit_r57_c227 bl[227] br[227] wl[57] vdd gnd cell_6t
Xbit_r58_c227 bl[227] br[227] wl[58] vdd gnd cell_6t
Xbit_r59_c227 bl[227] br[227] wl[59] vdd gnd cell_6t
Xbit_r60_c227 bl[227] br[227] wl[60] vdd gnd cell_6t
Xbit_r61_c227 bl[227] br[227] wl[61] vdd gnd cell_6t
Xbit_r62_c227 bl[227] br[227] wl[62] vdd gnd cell_6t
Xbit_r63_c227 bl[227] br[227] wl[63] vdd gnd cell_6t
Xbit_r64_c227 bl[227] br[227] wl[64] vdd gnd cell_6t
Xbit_r65_c227 bl[227] br[227] wl[65] vdd gnd cell_6t
Xbit_r66_c227 bl[227] br[227] wl[66] vdd gnd cell_6t
Xbit_r67_c227 bl[227] br[227] wl[67] vdd gnd cell_6t
Xbit_r68_c227 bl[227] br[227] wl[68] vdd gnd cell_6t
Xbit_r69_c227 bl[227] br[227] wl[69] vdd gnd cell_6t
Xbit_r70_c227 bl[227] br[227] wl[70] vdd gnd cell_6t
Xbit_r71_c227 bl[227] br[227] wl[71] vdd gnd cell_6t
Xbit_r72_c227 bl[227] br[227] wl[72] vdd gnd cell_6t
Xbit_r73_c227 bl[227] br[227] wl[73] vdd gnd cell_6t
Xbit_r74_c227 bl[227] br[227] wl[74] vdd gnd cell_6t
Xbit_r75_c227 bl[227] br[227] wl[75] vdd gnd cell_6t
Xbit_r76_c227 bl[227] br[227] wl[76] vdd gnd cell_6t
Xbit_r77_c227 bl[227] br[227] wl[77] vdd gnd cell_6t
Xbit_r78_c227 bl[227] br[227] wl[78] vdd gnd cell_6t
Xbit_r79_c227 bl[227] br[227] wl[79] vdd gnd cell_6t
Xbit_r80_c227 bl[227] br[227] wl[80] vdd gnd cell_6t
Xbit_r81_c227 bl[227] br[227] wl[81] vdd gnd cell_6t
Xbit_r82_c227 bl[227] br[227] wl[82] vdd gnd cell_6t
Xbit_r83_c227 bl[227] br[227] wl[83] vdd gnd cell_6t
Xbit_r84_c227 bl[227] br[227] wl[84] vdd gnd cell_6t
Xbit_r85_c227 bl[227] br[227] wl[85] vdd gnd cell_6t
Xbit_r86_c227 bl[227] br[227] wl[86] vdd gnd cell_6t
Xbit_r87_c227 bl[227] br[227] wl[87] vdd gnd cell_6t
Xbit_r88_c227 bl[227] br[227] wl[88] vdd gnd cell_6t
Xbit_r89_c227 bl[227] br[227] wl[89] vdd gnd cell_6t
Xbit_r90_c227 bl[227] br[227] wl[90] vdd gnd cell_6t
Xbit_r91_c227 bl[227] br[227] wl[91] vdd gnd cell_6t
Xbit_r92_c227 bl[227] br[227] wl[92] vdd gnd cell_6t
Xbit_r93_c227 bl[227] br[227] wl[93] vdd gnd cell_6t
Xbit_r94_c227 bl[227] br[227] wl[94] vdd gnd cell_6t
Xbit_r95_c227 bl[227] br[227] wl[95] vdd gnd cell_6t
Xbit_r96_c227 bl[227] br[227] wl[96] vdd gnd cell_6t
Xbit_r97_c227 bl[227] br[227] wl[97] vdd gnd cell_6t
Xbit_r98_c227 bl[227] br[227] wl[98] vdd gnd cell_6t
Xbit_r99_c227 bl[227] br[227] wl[99] vdd gnd cell_6t
Xbit_r100_c227 bl[227] br[227] wl[100] vdd gnd cell_6t
Xbit_r101_c227 bl[227] br[227] wl[101] vdd gnd cell_6t
Xbit_r102_c227 bl[227] br[227] wl[102] vdd gnd cell_6t
Xbit_r103_c227 bl[227] br[227] wl[103] vdd gnd cell_6t
Xbit_r104_c227 bl[227] br[227] wl[104] vdd gnd cell_6t
Xbit_r105_c227 bl[227] br[227] wl[105] vdd gnd cell_6t
Xbit_r106_c227 bl[227] br[227] wl[106] vdd gnd cell_6t
Xbit_r107_c227 bl[227] br[227] wl[107] vdd gnd cell_6t
Xbit_r108_c227 bl[227] br[227] wl[108] vdd gnd cell_6t
Xbit_r109_c227 bl[227] br[227] wl[109] vdd gnd cell_6t
Xbit_r110_c227 bl[227] br[227] wl[110] vdd gnd cell_6t
Xbit_r111_c227 bl[227] br[227] wl[111] vdd gnd cell_6t
Xbit_r112_c227 bl[227] br[227] wl[112] vdd gnd cell_6t
Xbit_r113_c227 bl[227] br[227] wl[113] vdd gnd cell_6t
Xbit_r114_c227 bl[227] br[227] wl[114] vdd gnd cell_6t
Xbit_r115_c227 bl[227] br[227] wl[115] vdd gnd cell_6t
Xbit_r116_c227 bl[227] br[227] wl[116] vdd gnd cell_6t
Xbit_r117_c227 bl[227] br[227] wl[117] vdd gnd cell_6t
Xbit_r118_c227 bl[227] br[227] wl[118] vdd gnd cell_6t
Xbit_r119_c227 bl[227] br[227] wl[119] vdd gnd cell_6t
Xbit_r120_c227 bl[227] br[227] wl[120] vdd gnd cell_6t
Xbit_r121_c227 bl[227] br[227] wl[121] vdd gnd cell_6t
Xbit_r122_c227 bl[227] br[227] wl[122] vdd gnd cell_6t
Xbit_r123_c227 bl[227] br[227] wl[123] vdd gnd cell_6t
Xbit_r124_c227 bl[227] br[227] wl[124] vdd gnd cell_6t
Xbit_r125_c227 bl[227] br[227] wl[125] vdd gnd cell_6t
Xbit_r126_c227 bl[227] br[227] wl[126] vdd gnd cell_6t
Xbit_r127_c227 bl[227] br[227] wl[127] vdd gnd cell_6t
Xbit_r128_c227 bl[227] br[227] wl[128] vdd gnd cell_6t
Xbit_r129_c227 bl[227] br[227] wl[129] vdd gnd cell_6t
Xbit_r130_c227 bl[227] br[227] wl[130] vdd gnd cell_6t
Xbit_r131_c227 bl[227] br[227] wl[131] vdd gnd cell_6t
Xbit_r132_c227 bl[227] br[227] wl[132] vdd gnd cell_6t
Xbit_r133_c227 bl[227] br[227] wl[133] vdd gnd cell_6t
Xbit_r134_c227 bl[227] br[227] wl[134] vdd gnd cell_6t
Xbit_r135_c227 bl[227] br[227] wl[135] vdd gnd cell_6t
Xbit_r136_c227 bl[227] br[227] wl[136] vdd gnd cell_6t
Xbit_r137_c227 bl[227] br[227] wl[137] vdd gnd cell_6t
Xbit_r138_c227 bl[227] br[227] wl[138] vdd gnd cell_6t
Xbit_r139_c227 bl[227] br[227] wl[139] vdd gnd cell_6t
Xbit_r140_c227 bl[227] br[227] wl[140] vdd gnd cell_6t
Xbit_r141_c227 bl[227] br[227] wl[141] vdd gnd cell_6t
Xbit_r142_c227 bl[227] br[227] wl[142] vdd gnd cell_6t
Xbit_r143_c227 bl[227] br[227] wl[143] vdd gnd cell_6t
Xbit_r144_c227 bl[227] br[227] wl[144] vdd gnd cell_6t
Xbit_r145_c227 bl[227] br[227] wl[145] vdd gnd cell_6t
Xbit_r146_c227 bl[227] br[227] wl[146] vdd gnd cell_6t
Xbit_r147_c227 bl[227] br[227] wl[147] vdd gnd cell_6t
Xbit_r148_c227 bl[227] br[227] wl[148] vdd gnd cell_6t
Xbit_r149_c227 bl[227] br[227] wl[149] vdd gnd cell_6t
Xbit_r150_c227 bl[227] br[227] wl[150] vdd gnd cell_6t
Xbit_r151_c227 bl[227] br[227] wl[151] vdd gnd cell_6t
Xbit_r152_c227 bl[227] br[227] wl[152] vdd gnd cell_6t
Xbit_r153_c227 bl[227] br[227] wl[153] vdd gnd cell_6t
Xbit_r154_c227 bl[227] br[227] wl[154] vdd gnd cell_6t
Xbit_r155_c227 bl[227] br[227] wl[155] vdd gnd cell_6t
Xbit_r156_c227 bl[227] br[227] wl[156] vdd gnd cell_6t
Xbit_r157_c227 bl[227] br[227] wl[157] vdd gnd cell_6t
Xbit_r158_c227 bl[227] br[227] wl[158] vdd gnd cell_6t
Xbit_r159_c227 bl[227] br[227] wl[159] vdd gnd cell_6t
Xbit_r160_c227 bl[227] br[227] wl[160] vdd gnd cell_6t
Xbit_r161_c227 bl[227] br[227] wl[161] vdd gnd cell_6t
Xbit_r162_c227 bl[227] br[227] wl[162] vdd gnd cell_6t
Xbit_r163_c227 bl[227] br[227] wl[163] vdd gnd cell_6t
Xbit_r164_c227 bl[227] br[227] wl[164] vdd gnd cell_6t
Xbit_r165_c227 bl[227] br[227] wl[165] vdd gnd cell_6t
Xbit_r166_c227 bl[227] br[227] wl[166] vdd gnd cell_6t
Xbit_r167_c227 bl[227] br[227] wl[167] vdd gnd cell_6t
Xbit_r168_c227 bl[227] br[227] wl[168] vdd gnd cell_6t
Xbit_r169_c227 bl[227] br[227] wl[169] vdd gnd cell_6t
Xbit_r170_c227 bl[227] br[227] wl[170] vdd gnd cell_6t
Xbit_r171_c227 bl[227] br[227] wl[171] vdd gnd cell_6t
Xbit_r172_c227 bl[227] br[227] wl[172] vdd gnd cell_6t
Xbit_r173_c227 bl[227] br[227] wl[173] vdd gnd cell_6t
Xbit_r174_c227 bl[227] br[227] wl[174] vdd gnd cell_6t
Xbit_r175_c227 bl[227] br[227] wl[175] vdd gnd cell_6t
Xbit_r176_c227 bl[227] br[227] wl[176] vdd gnd cell_6t
Xbit_r177_c227 bl[227] br[227] wl[177] vdd gnd cell_6t
Xbit_r178_c227 bl[227] br[227] wl[178] vdd gnd cell_6t
Xbit_r179_c227 bl[227] br[227] wl[179] vdd gnd cell_6t
Xbit_r180_c227 bl[227] br[227] wl[180] vdd gnd cell_6t
Xbit_r181_c227 bl[227] br[227] wl[181] vdd gnd cell_6t
Xbit_r182_c227 bl[227] br[227] wl[182] vdd gnd cell_6t
Xbit_r183_c227 bl[227] br[227] wl[183] vdd gnd cell_6t
Xbit_r184_c227 bl[227] br[227] wl[184] vdd gnd cell_6t
Xbit_r185_c227 bl[227] br[227] wl[185] vdd gnd cell_6t
Xbit_r186_c227 bl[227] br[227] wl[186] vdd gnd cell_6t
Xbit_r187_c227 bl[227] br[227] wl[187] vdd gnd cell_6t
Xbit_r188_c227 bl[227] br[227] wl[188] vdd gnd cell_6t
Xbit_r189_c227 bl[227] br[227] wl[189] vdd gnd cell_6t
Xbit_r190_c227 bl[227] br[227] wl[190] vdd gnd cell_6t
Xbit_r191_c227 bl[227] br[227] wl[191] vdd gnd cell_6t
Xbit_r192_c227 bl[227] br[227] wl[192] vdd gnd cell_6t
Xbit_r193_c227 bl[227] br[227] wl[193] vdd gnd cell_6t
Xbit_r194_c227 bl[227] br[227] wl[194] vdd gnd cell_6t
Xbit_r195_c227 bl[227] br[227] wl[195] vdd gnd cell_6t
Xbit_r196_c227 bl[227] br[227] wl[196] vdd gnd cell_6t
Xbit_r197_c227 bl[227] br[227] wl[197] vdd gnd cell_6t
Xbit_r198_c227 bl[227] br[227] wl[198] vdd gnd cell_6t
Xbit_r199_c227 bl[227] br[227] wl[199] vdd gnd cell_6t
Xbit_r200_c227 bl[227] br[227] wl[200] vdd gnd cell_6t
Xbit_r201_c227 bl[227] br[227] wl[201] vdd gnd cell_6t
Xbit_r202_c227 bl[227] br[227] wl[202] vdd gnd cell_6t
Xbit_r203_c227 bl[227] br[227] wl[203] vdd gnd cell_6t
Xbit_r204_c227 bl[227] br[227] wl[204] vdd gnd cell_6t
Xbit_r205_c227 bl[227] br[227] wl[205] vdd gnd cell_6t
Xbit_r206_c227 bl[227] br[227] wl[206] vdd gnd cell_6t
Xbit_r207_c227 bl[227] br[227] wl[207] vdd gnd cell_6t
Xbit_r208_c227 bl[227] br[227] wl[208] vdd gnd cell_6t
Xbit_r209_c227 bl[227] br[227] wl[209] vdd gnd cell_6t
Xbit_r210_c227 bl[227] br[227] wl[210] vdd gnd cell_6t
Xbit_r211_c227 bl[227] br[227] wl[211] vdd gnd cell_6t
Xbit_r212_c227 bl[227] br[227] wl[212] vdd gnd cell_6t
Xbit_r213_c227 bl[227] br[227] wl[213] vdd gnd cell_6t
Xbit_r214_c227 bl[227] br[227] wl[214] vdd gnd cell_6t
Xbit_r215_c227 bl[227] br[227] wl[215] vdd gnd cell_6t
Xbit_r216_c227 bl[227] br[227] wl[216] vdd gnd cell_6t
Xbit_r217_c227 bl[227] br[227] wl[217] vdd gnd cell_6t
Xbit_r218_c227 bl[227] br[227] wl[218] vdd gnd cell_6t
Xbit_r219_c227 bl[227] br[227] wl[219] vdd gnd cell_6t
Xbit_r220_c227 bl[227] br[227] wl[220] vdd gnd cell_6t
Xbit_r221_c227 bl[227] br[227] wl[221] vdd gnd cell_6t
Xbit_r222_c227 bl[227] br[227] wl[222] vdd gnd cell_6t
Xbit_r223_c227 bl[227] br[227] wl[223] vdd gnd cell_6t
Xbit_r224_c227 bl[227] br[227] wl[224] vdd gnd cell_6t
Xbit_r225_c227 bl[227] br[227] wl[225] vdd gnd cell_6t
Xbit_r226_c227 bl[227] br[227] wl[226] vdd gnd cell_6t
Xbit_r227_c227 bl[227] br[227] wl[227] vdd gnd cell_6t
Xbit_r228_c227 bl[227] br[227] wl[228] vdd gnd cell_6t
Xbit_r229_c227 bl[227] br[227] wl[229] vdd gnd cell_6t
Xbit_r230_c227 bl[227] br[227] wl[230] vdd gnd cell_6t
Xbit_r231_c227 bl[227] br[227] wl[231] vdd gnd cell_6t
Xbit_r232_c227 bl[227] br[227] wl[232] vdd gnd cell_6t
Xbit_r233_c227 bl[227] br[227] wl[233] vdd gnd cell_6t
Xbit_r234_c227 bl[227] br[227] wl[234] vdd gnd cell_6t
Xbit_r235_c227 bl[227] br[227] wl[235] vdd gnd cell_6t
Xbit_r236_c227 bl[227] br[227] wl[236] vdd gnd cell_6t
Xbit_r237_c227 bl[227] br[227] wl[237] vdd gnd cell_6t
Xbit_r238_c227 bl[227] br[227] wl[238] vdd gnd cell_6t
Xbit_r239_c227 bl[227] br[227] wl[239] vdd gnd cell_6t
Xbit_r240_c227 bl[227] br[227] wl[240] vdd gnd cell_6t
Xbit_r241_c227 bl[227] br[227] wl[241] vdd gnd cell_6t
Xbit_r242_c227 bl[227] br[227] wl[242] vdd gnd cell_6t
Xbit_r243_c227 bl[227] br[227] wl[243] vdd gnd cell_6t
Xbit_r244_c227 bl[227] br[227] wl[244] vdd gnd cell_6t
Xbit_r245_c227 bl[227] br[227] wl[245] vdd gnd cell_6t
Xbit_r246_c227 bl[227] br[227] wl[246] vdd gnd cell_6t
Xbit_r247_c227 bl[227] br[227] wl[247] vdd gnd cell_6t
Xbit_r248_c227 bl[227] br[227] wl[248] vdd gnd cell_6t
Xbit_r249_c227 bl[227] br[227] wl[249] vdd gnd cell_6t
Xbit_r250_c227 bl[227] br[227] wl[250] vdd gnd cell_6t
Xbit_r251_c227 bl[227] br[227] wl[251] vdd gnd cell_6t
Xbit_r252_c227 bl[227] br[227] wl[252] vdd gnd cell_6t
Xbit_r253_c227 bl[227] br[227] wl[253] vdd gnd cell_6t
Xbit_r254_c227 bl[227] br[227] wl[254] vdd gnd cell_6t
Xbit_r255_c227 bl[227] br[227] wl[255] vdd gnd cell_6t
Xbit_r0_c228 bl[228] br[228] wl[0] vdd gnd cell_6t
Xbit_r1_c228 bl[228] br[228] wl[1] vdd gnd cell_6t
Xbit_r2_c228 bl[228] br[228] wl[2] vdd gnd cell_6t
Xbit_r3_c228 bl[228] br[228] wl[3] vdd gnd cell_6t
Xbit_r4_c228 bl[228] br[228] wl[4] vdd gnd cell_6t
Xbit_r5_c228 bl[228] br[228] wl[5] vdd gnd cell_6t
Xbit_r6_c228 bl[228] br[228] wl[6] vdd gnd cell_6t
Xbit_r7_c228 bl[228] br[228] wl[7] vdd gnd cell_6t
Xbit_r8_c228 bl[228] br[228] wl[8] vdd gnd cell_6t
Xbit_r9_c228 bl[228] br[228] wl[9] vdd gnd cell_6t
Xbit_r10_c228 bl[228] br[228] wl[10] vdd gnd cell_6t
Xbit_r11_c228 bl[228] br[228] wl[11] vdd gnd cell_6t
Xbit_r12_c228 bl[228] br[228] wl[12] vdd gnd cell_6t
Xbit_r13_c228 bl[228] br[228] wl[13] vdd gnd cell_6t
Xbit_r14_c228 bl[228] br[228] wl[14] vdd gnd cell_6t
Xbit_r15_c228 bl[228] br[228] wl[15] vdd gnd cell_6t
Xbit_r16_c228 bl[228] br[228] wl[16] vdd gnd cell_6t
Xbit_r17_c228 bl[228] br[228] wl[17] vdd gnd cell_6t
Xbit_r18_c228 bl[228] br[228] wl[18] vdd gnd cell_6t
Xbit_r19_c228 bl[228] br[228] wl[19] vdd gnd cell_6t
Xbit_r20_c228 bl[228] br[228] wl[20] vdd gnd cell_6t
Xbit_r21_c228 bl[228] br[228] wl[21] vdd gnd cell_6t
Xbit_r22_c228 bl[228] br[228] wl[22] vdd gnd cell_6t
Xbit_r23_c228 bl[228] br[228] wl[23] vdd gnd cell_6t
Xbit_r24_c228 bl[228] br[228] wl[24] vdd gnd cell_6t
Xbit_r25_c228 bl[228] br[228] wl[25] vdd gnd cell_6t
Xbit_r26_c228 bl[228] br[228] wl[26] vdd gnd cell_6t
Xbit_r27_c228 bl[228] br[228] wl[27] vdd gnd cell_6t
Xbit_r28_c228 bl[228] br[228] wl[28] vdd gnd cell_6t
Xbit_r29_c228 bl[228] br[228] wl[29] vdd gnd cell_6t
Xbit_r30_c228 bl[228] br[228] wl[30] vdd gnd cell_6t
Xbit_r31_c228 bl[228] br[228] wl[31] vdd gnd cell_6t
Xbit_r32_c228 bl[228] br[228] wl[32] vdd gnd cell_6t
Xbit_r33_c228 bl[228] br[228] wl[33] vdd gnd cell_6t
Xbit_r34_c228 bl[228] br[228] wl[34] vdd gnd cell_6t
Xbit_r35_c228 bl[228] br[228] wl[35] vdd gnd cell_6t
Xbit_r36_c228 bl[228] br[228] wl[36] vdd gnd cell_6t
Xbit_r37_c228 bl[228] br[228] wl[37] vdd gnd cell_6t
Xbit_r38_c228 bl[228] br[228] wl[38] vdd gnd cell_6t
Xbit_r39_c228 bl[228] br[228] wl[39] vdd gnd cell_6t
Xbit_r40_c228 bl[228] br[228] wl[40] vdd gnd cell_6t
Xbit_r41_c228 bl[228] br[228] wl[41] vdd gnd cell_6t
Xbit_r42_c228 bl[228] br[228] wl[42] vdd gnd cell_6t
Xbit_r43_c228 bl[228] br[228] wl[43] vdd gnd cell_6t
Xbit_r44_c228 bl[228] br[228] wl[44] vdd gnd cell_6t
Xbit_r45_c228 bl[228] br[228] wl[45] vdd gnd cell_6t
Xbit_r46_c228 bl[228] br[228] wl[46] vdd gnd cell_6t
Xbit_r47_c228 bl[228] br[228] wl[47] vdd gnd cell_6t
Xbit_r48_c228 bl[228] br[228] wl[48] vdd gnd cell_6t
Xbit_r49_c228 bl[228] br[228] wl[49] vdd gnd cell_6t
Xbit_r50_c228 bl[228] br[228] wl[50] vdd gnd cell_6t
Xbit_r51_c228 bl[228] br[228] wl[51] vdd gnd cell_6t
Xbit_r52_c228 bl[228] br[228] wl[52] vdd gnd cell_6t
Xbit_r53_c228 bl[228] br[228] wl[53] vdd gnd cell_6t
Xbit_r54_c228 bl[228] br[228] wl[54] vdd gnd cell_6t
Xbit_r55_c228 bl[228] br[228] wl[55] vdd gnd cell_6t
Xbit_r56_c228 bl[228] br[228] wl[56] vdd gnd cell_6t
Xbit_r57_c228 bl[228] br[228] wl[57] vdd gnd cell_6t
Xbit_r58_c228 bl[228] br[228] wl[58] vdd gnd cell_6t
Xbit_r59_c228 bl[228] br[228] wl[59] vdd gnd cell_6t
Xbit_r60_c228 bl[228] br[228] wl[60] vdd gnd cell_6t
Xbit_r61_c228 bl[228] br[228] wl[61] vdd gnd cell_6t
Xbit_r62_c228 bl[228] br[228] wl[62] vdd gnd cell_6t
Xbit_r63_c228 bl[228] br[228] wl[63] vdd gnd cell_6t
Xbit_r64_c228 bl[228] br[228] wl[64] vdd gnd cell_6t
Xbit_r65_c228 bl[228] br[228] wl[65] vdd gnd cell_6t
Xbit_r66_c228 bl[228] br[228] wl[66] vdd gnd cell_6t
Xbit_r67_c228 bl[228] br[228] wl[67] vdd gnd cell_6t
Xbit_r68_c228 bl[228] br[228] wl[68] vdd gnd cell_6t
Xbit_r69_c228 bl[228] br[228] wl[69] vdd gnd cell_6t
Xbit_r70_c228 bl[228] br[228] wl[70] vdd gnd cell_6t
Xbit_r71_c228 bl[228] br[228] wl[71] vdd gnd cell_6t
Xbit_r72_c228 bl[228] br[228] wl[72] vdd gnd cell_6t
Xbit_r73_c228 bl[228] br[228] wl[73] vdd gnd cell_6t
Xbit_r74_c228 bl[228] br[228] wl[74] vdd gnd cell_6t
Xbit_r75_c228 bl[228] br[228] wl[75] vdd gnd cell_6t
Xbit_r76_c228 bl[228] br[228] wl[76] vdd gnd cell_6t
Xbit_r77_c228 bl[228] br[228] wl[77] vdd gnd cell_6t
Xbit_r78_c228 bl[228] br[228] wl[78] vdd gnd cell_6t
Xbit_r79_c228 bl[228] br[228] wl[79] vdd gnd cell_6t
Xbit_r80_c228 bl[228] br[228] wl[80] vdd gnd cell_6t
Xbit_r81_c228 bl[228] br[228] wl[81] vdd gnd cell_6t
Xbit_r82_c228 bl[228] br[228] wl[82] vdd gnd cell_6t
Xbit_r83_c228 bl[228] br[228] wl[83] vdd gnd cell_6t
Xbit_r84_c228 bl[228] br[228] wl[84] vdd gnd cell_6t
Xbit_r85_c228 bl[228] br[228] wl[85] vdd gnd cell_6t
Xbit_r86_c228 bl[228] br[228] wl[86] vdd gnd cell_6t
Xbit_r87_c228 bl[228] br[228] wl[87] vdd gnd cell_6t
Xbit_r88_c228 bl[228] br[228] wl[88] vdd gnd cell_6t
Xbit_r89_c228 bl[228] br[228] wl[89] vdd gnd cell_6t
Xbit_r90_c228 bl[228] br[228] wl[90] vdd gnd cell_6t
Xbit_r91_c228 bl[228] br[228] wl[91] vdd gnd cell_6t
Xbit_r92_c228 bl[228] br[228] wl[92] vdd gnd cell_6t
Xbit_r93_c228 bl[228] br[228] wl[93] vdd gnd cell_6t
Xbit_r94_c228 bl[228] br[228] wl[94] vdd gnd cell_6t
Xbit_r95_c228 bl[228] br[228] wl[95] vdd gnd cell_6t
Xbit_r96_c228 bl[228] br[228] wl[96] vdd gnd cell_6t
Xbit_r97_c228 bl[228] br[228] wl[97] vdd gnd cell_6t
Xbit_r98_c228 bl[228] br[228] wl[98] vdd gnd cell_6t
Xbit_r99_c228 bl[228] br[228] wl[99] vdd gnd cell_6t
Xbit_r100_c228 bl[228] br[228] wl[100] vdd gnd cell_6t
Xbit_r101_c228 bl[228] br[228] wl[101] vdd gnd cell_6t
Xbit_r102_c228 bl[228] br[228] wl[102] vdd gnd cell_6t
Xbit_r103_c228 bl[228] br[228] wl[103] vdd gnd cell_6t
Xbit_r104_c228 bl[228] br[228] wl[104] vdd gnd cell_6t
Xbit_r105_c228 bl[228] br[228] wl[105] vdd gnd cell_6t
Xbit_r106_c228 bl[228] br[228] wl[106] vdd gnd cell_6t
Xbit_r107_c228 bl[228] br[228] wl[107] vdd gnd cell_6t
Xbit_r108_c228 bl[228] br[228] wl[108] vdd gnd cell_6t
Xbit_r109_c228 bl[228] br[228] wl[109] vdd gnd cell_6t
Xbit_r110_c228 bl[228] br[228] wl[110] vdd gnd cell_6t
Xbit_r111_c228 bl[228] br[228] wl[111] vdd gnd cell_6t
Xbit_r112_c228 bl[228] br[228] wl[112] vdd gnd cell_6t
Xbit_r113_c228 bl[228] br[228] wl[113] vdd gnd cell_6t
Xbit_r114_c228 bl[228] br[228] wl[114] vdd gnd cell_6t
Xbit_r115_c228 bl[228] br[228] wl[115] vdd gnd cell_6t
Xbit_r116_c228 bl[228] br[228] wl[116] vdd gnd cell_6t
Xbit_r117_c228 bl[228] br[228] wl[117] vdd gnd cell_6t
Xbit_r118_c228 bl[228] br[228] wl[118] vdd gnd cell_6t
Xbit_r119_c228 bl[228] br[228] wl[119] vdd gnd cell_6t
Xbit_r120_c228 bl[228] br[228] wl[120] vdd gnd cell_6t
Xbit_r121_c228 bl[228] br[228] wl[121] vdd gnd cell_6t
Xbit_r122_c228 bl[228] br[228] wl[122] vdd gnd cell_6t
Xbit_r123_c228 bl[228] br[228] wl[123] vdd gnd cell_6t
Xbit_r124_c228 bl[228] br[228] wl[124] vdd gnd cell_6t
Xbit_r125_c228 bl[228] br[228] wl[125] vdd gnd cell_6t
Xbit_r126_c228 bl[228] br[228] wl[126] vdd gnd cell_6t
Xbit_r127_c228 bl[228] br[228] wl[127] vdd gnd cell_6t
Xbit_r128_c228 bl[228] br[228] wl[128] vdd gnd cell_6t
Xbit_r129_c228 bl[228] br[228] wl[129] vdd gnd cell_6t
Xbit_r130_c228 bl[228] br[228] wl[130] vdd gnd cell_6t
Xbit_r131_c228 bl[228] br[228] wl[131] vdd gnd cell_6t
Xbit_r132_c228 bl[228] br[228] wl[132] vdd gnd cell_6t
Xbit_r133_c228 bl[228] br[228] wl[133] vdd gnd cell_6t
Xbit_r134_c228 bl[228] br[228] wl[134] vdd gnd cell_6t
Xbit_r135_c228 bl[228] br[228] wl[135] vdd gnd cell_6t
Xbit_r136_c228 bl[228] br[228] wl[136] vdd gnd cell_6t
Xbit_r137_c228 bl[228] br[228] wl[137] vdd gnd cell_6t
Xbit_r138_c228 bl[228] br[228] wl[138] vdd gnd cell_6t
Xbit_r139_c228 bl[228] br[228] wl[139] vdd gnd cell_6t
Xbit_r140_c228 bl[228] br[228] wl[140] vdd gnd cell_6t
Xbit_r141_c228 bl[228] br[228] wl[141] vdd gnd cell_6t
Xbit_r142_c228 bl[228] br[228] wl[142] vdd gnd cell_6t
Xbit_r143_c228 bl[228] br[228] wl[143] vdd gnd cell_6t
Xbit_r144_c228 bl[228] br[228] wl[144] vdd gnd cell_6t
Xbit_r145_c228 bl[228] br[228] wl[145] vdd gnd cell_6t
Xbit_r146_c228 bl[228] br[228] wl[146] vdd gnd cell_6t
Xbit_r147_c228 bl[228] br[228] wl[147] vdd gnd cell_6t
Xbit_r148_c228 bl[228] br[228] wl[148] vdd gnd cell_6t
Xbit_r149_c228 bl[228] br[228] wl[149] vdd gnd cell_6t
Xbit_r150_c228 bl[228] br[228] wl[150] vdd gnd cell_6t
Xbit_r151_c228 bl[228] br[228] wl[151] vdd gnd cell_6t
Xbit_r152_c228 bl[228] br[228] wl[152] vdd gnd cell_6t
Xbit_r153_c228 bl[228] br[228] wl[153] vdd gnd cell_6t
Xbit_r154_c228 bl[228] br[228] wl[154] vdd gnd cell_6t
Xbit_r155_c228 bl[228] br[228] wl[155] vdd gnd cell_6t
Xbit_r156_c228 bl[228] br[228] wl[156] vdd gnd cell_6t
Xbit_r157_c228 bl[228] br[228] wl[157] vdd gnd cell_6t
Xbit_r158_c228 bl[228] br[228] wl[158] vdd gnd cell_6t
Xbit_r159_c228 bl[228] br[228] wl[159] vdd gnd cell_6t
Xbit_r160_c228 bl[228] br[228] wl[160] vdd gnd cell_6t
Xbit_r161_c228 bl[228] br[228] wl[161] vdd gnd cell_6t
Xbit_r162_c228 bl[228] br[228] wl[162] vdd gnd cell_6t
Xbit_r163_c228 bl[228] br[228] wl[163] vdd gnd cell_6t
Xbit_r164_c228 bl[228] br[228] wl[164] vdd gnd cell_6t
Xbit_r165_c228 bl[228] br[228] wl[165] vdd gnd cell_6t
Xbit_r166_c228 bl[228] br[228] wl[166] vdd gnd cell_6t
Xbit_r167_c228 bl[228] br[228] wl[167] vdd gnd cell_6t
Xbit_r168_c228 bl[228] br[228] wl[168] vdd gnd cell_6t
Xbit_r169_c228 bl[228] br[228] wl[169] vdd gnd cell_6t
Xbit_r170_c228 bl[228] br[228] wl[170] vdd gnd cell_6t
Xbit_r171_c228 bl[228] br[228] wl[171] vdd gnd cell_6t
Xbit_r172_c228 bl[228] br[228] wl[172] vdd gnd cell_6t
Xbit_r173_c228 bl[228] br[228] wl[173] vdd gnd cell_6t
Xbit_r174_c228 bl[228] br[228] wl[174] vdd gnd cell_6t
Xbit_r175_c228 bl[228] br[228] wl[175] vdd gnd cell_6t
Xbit_r176_c228 bl[228] br[228] wl[176] vdd gnd cell_6t
Xbit_r177_c228 bl[228] br[228] wl[177] vdd gnd cell_6t
Xbit_r178_c228 bl[228] br[228] wl[178] vdd gnd cell_6t
Xbit_r179_c228 bl[228] br[228] wl[179] vdd gnd cell_6t
Xbit_r180_c228 bl[228] br[228] wl[180] vdd gnd cell_6t
Xbit_r181_c228 bl[228] br[228] wl[181] vdd gnd cell_6t
Xbit_r182_c228 bl[228] br[228] wl[182] vdd gnd cell_6t
Xbit_r183_c228 bl[228] br[228] wl[183] vdd gnd cell_6t
Xbit_r184_c228 bl[228] br[228] wl[184] vdd gnd cell_6t
Xbit_r185_c228 bl[228] br[228] wl[185] vdd gnd cell_6t
Xbit_r186_c228 bl[228] br[228] wl[186] vdd gnd cell_6t
Xbit_r187_c228 bl[228] br[228] wl[187] vdd gnd cell_6t
Xbit_r188_c228 bl[228] br[228] wl[188] vdd gnd cell_6t
Xbit_r189_c228 bl[228] br[228] wl[189] vdd gnd cell_6t
Xbit_r190_c228 bl[228] br[228] wl[190] vdd gnd cell_6t
Xbit_r191_c228 bl[228] br[228] wl[191] vdd gnd cell_6t
Xbit_r192_c228 bl[228] br[228] wl[192] vdd gnd cell_6t
Xbit_r193_c228 bl[228] br[228] wl[193] vdd gnd cell_6t
Xbit_r194_c228 bl[228] br[228] wl[194] vdd gnd cell_6t
Xbit_r195_c228 bl[228] br[228] wl[195] vdd gnd cell_6t
Xbit_r196_c228 bl[228] br[228] wl[196] vdd gnd cell_6t
Xbit_r197_c228 bl[228] br[228] wl[197] vdd gnd cell_6t
Xbit_r198_c228 bl[228] br[228] wl[198] vdd gnd cell_6t
Xbit_r199_c228 bl[228] br[228] wl[199] vdd gnd cell_6t
Xbit_r200_c228 bl[228] br[228] wl[200] vdd gnd cell_6t
Xbit_r201_c228 bl[228] br[228] wl[201] vdd gnd cell_6t
Xbit_r202_c228 bl[228] br[228] wl[202] vdd gnd cell_6t
Xbit_r203_c228 bl[228] br[228] wl[203] vdd gnd cell_6t
Xbit_r204_c228 bl[228] br[228] wl[204] vdd gnd cell_6t
Xbit_r205_c228 bl[228] br[228] wl[205] vdd gnd cell_6t
Xbit_r206_c228 bl[228] br[228] wl[206] vdd gnd cell_6t
Xbit_r207_c228 bl[228] br[228] wl[207] vdd gnd cell_6t
Xbit_r208_c228 bl[228] br[228] wl[208] vdd gnd cell_6t
Xbit_r209_c228 bl[228] br[228] wl[209] vdd gnd cell_6t
Xbit_r210_c228 bl[228] br[228] wl[210] vdd gnd cell_6t
Xbit_r211_c228 bl[228] br[228] wl[211] vdd gnd cell_6t
Xbit_r212_c228 bl[228] br[228] wl[212] vdd gnd cell_6t
Xbit_r213_c228 bl[228] br[228] wl[213] vdd gnd cell_6t
Xbit_r214_c228 bl[228] br[228] wl[214] vdd gnd cell_6t
Xbit_r215_c228 bl[228] br[228] wl[215] vdd gnd cell_6t
Xbit_r216_c228 bl[228] br[228] wl[216] vdd gnd cell_6t
Xbit_r217_c228 bl[228] br[228] wl[217] vdd gnd cell_6t
Xbit_r218_c228 bl[228] br[228] wl[218] vdd gnd cell_6t
Xbit_r219_c228 bl[228] br[228] wl[219] vdd gnd cell_6t
Xbit_r220_c228 bl[228] br[228] wl[220] vdd gnd cell_6t
Xbit_r221_c228 bl[228] br[228] wl[221] vdd gnd cell_6t
Xbit_r222_c228 bl[228] br[228] wl[222] vdd gnd cell_6t
Xbit_r223_c228 bl[228] br[228] wl[223] vdd gnd cell_6t
Xbit_r224_c228 bl[228] br[228] wl[224] vdd gnd cell_6t
Xbit_r225_c228 bl[228] br[228] wl[225] vdd gnd cell_6t
Xbit_r226_c228 bl[228] br[228] wl[226] vdd gnd cell_6t
Xbit_r227_c228 bl[228] br[228] wl[227] vdd gnd cell_6t
Xbit_r228_c228 bl[228] br[228] wl[228] vdd gnd cell_6t
Xbit_r229_c228 bl[228] br[228] wl[229] vdd gnd cell_6t
Xbit_r230_c228 bl[228] br[228] wl[230] vdd gnd cell_6t
Xbit_r231_c228 bl[228] br[228] wl[231] vdd gnd cell_6t
Xbit_r232_c228 bl[228] br[228] wl[232] vdd gnd cell_6t
Xbit_r233_c228 bl[228] br[228] wl[233] vdd gnd cell_6t
Xbit_r234_c228 bl[228] br[228] wl[234] vdd gnd cell_6t
Xbit_r235_c228 bl[228] br[228] wl[235] vdd gnd cell_6t
Xbit_r236_c228 bl[228] br[228] wl[236] vdd gnd cell_6t
Xbit_r237_c228 bl[228] br[228] wl[237] vdd gnd cell_6t
Xbit_r238_c228 bl[228] br[228] wl[238] vdd gnd cell_6t
Xbit_r239_c228 bl[228] br[228] wl[239] vdd gnd cell_6t
Xbit_r240_c228 bl[228] br[228] wl[240] vdd gnd cell_6t
Xbit_r241_c228 bl[228] br[228] wl[241] vdd gnd cell_6t
Xbit_r242_c228 bl[228] br[228] wl[242] vdd gnd cell_6t
Xbit_r243_c228 bl[228] br[228] wl[243] vdd gnd cell_6t
Xbit_r244_c228 bl[228] br[228] wl[244] vdd gnd cell_6t
Xbit_r245_c228 bl[228] br[228] wl[245] vdd gnd cell_6t
Xbit_r246_c228 bl[228] br[228] wl[246] vdd gnd cell_6t
Xbit_r247_c228 bl[228] br[228] wl[247] vdd gnd cell_6t
Xbit_r248_c228 bl[228] br[228] wl[248] vdd gnd cell_6t
Xbit_r249_c228 bl[228] br[228] wl[249] vdd gnd cell_6t
Xbit_r250_c228 bl[228] br[228] wl[250] vdd gnd cell_6t
Xbit_r251_c228 bl[228] br[228] wl[251] vdd gnd cell_6t
Xbit_r252_c228 bl[228] br[228] wl[252] vdd gnd cell_6t
Xbit_r253_c228 bl[228] br[228] wl[253] vdd gnd cell_6t
Xbit_r254_c228 bl[228] br[228] wl[254] vdd gnd cell_6t
Xbit_r255_c228 bl[228] br[228] wl[255] vdd gnd cell_6t
Xbit_r0_c229 bl[229] br[229] wl[0] vdd gnd cell_6t
Xbit_r1_c229 bl[229] br[229] wl[1] vdd gnd cell_6t
Xbit_r2_c229 bl[229] br[229] wl[2] vdd gnd cell_6t
Xbit_r3_c229 bl[229] br[229] wl[3] vdd gnd cell_6t
Xbit_r4_c229 bl[229] br[229] wl[4] vdd gnd cell_6t
Xbit_r5_c229 bl[229] br[229] wl[5] vdd gnd cell_6t
Xbit_r6_c229 bl[229] br[229] wl[6] vdd gnd cell_6t
Xbit_r7_c229 bl[229] br[229] wl[7] vdd gnd cell_6t
Xbit_r8_c229 bl[229] br[229] wl[8] vdd gnd cell_6t
Xbit_r9_c229 bl[229] br[229] wl[9] vdd gnd cell_6t
Xbit_r10_c229 bl[229] br[229] wl[10] vdd gnd cell_6t
Xbit_r11_c229 bl[229] br[229] wl[11] vdd gnd cell_6t
Xbit_r12_c229 bl[229] br[229] wl[12] vdd gnd cell_6t
Xbit_r13_c229 bl[229] br[229] wl[13] vdd gnd cell_6t
Xbit_r14_c229 bl[229] br[229] wl[14] vdd gnd cell_6t
Xbit_r15_c229 bl[229] br[229] wl[15] vdd gnd cell_6t
Xbit_r16_c229 bl[229] br[229] wl[16] vdd gnd cell_6t
Xbit_r17_c229 bl[229] br[229] wl[17] vdd gnd cell_6t
Xbit_r18_c229 bl[229] br[229] wl[18] vdd gnd cell_6t
Xbit_r19_c229 bl[229] br[229] wl[19] vdd gnd cell_6t
Xbit_r20_c229 bl[229] br[229] wl[20] vdd gnd cell_6t
Xbit_r21_c229 bl[229] br[229] wl[21] vdd gnd cell_6t
Xbit_r22_c229 bl[229] br[229] wl[22] vdd gnd cell_6t
Xbit_r23_c229 bl[229] br[229] wl[23] vdd gnd cell_6t
Xbit_r24_c229 bl[229] br[229] wl[24] vdd gnd cell_6t
Xbit_r25_c229 bl[229] br[229] wl[25] vdd gnd cell_6t
Xbit_r26_c229 bl[229] br[229] wl[26] vdd gnd cell_6t
Xbit_r27_c229 bl[229] br[229] wl[27] vdd gnd cell_6t
Xbit_r28_c229 bl[229] br[229] wl[28] vdd gnd cell_6t
Xbit_r29_c229 bl[229] br[229] wl[29] vdd gnd cell_6t
Xbit_r30_c229 bl[229] br[229] wl[30] vdd gnd cell_6t
Xbit_r31_c229 bl[229] br[229] wl[31] vdd gnd cell_6t
Xbit_r32_c229 bl[229] br[229] wl[32] vdd gnd cell_6t
Xbit_r33_c229 bl[229] br[229] wl[33] vdd gnd cell_6t
Xbit_r34_c229 bl[229] br[229] wl[34] vdd gnd cell_6t
Xbit_r35_c229 bl[229] br[229] wl[35] vdd gnd cell_6t
Xbit_r36_c229 bl[229] br[229] wl[36] vdd gnd cell_6t
Xbit_r37_c229 bl[229] br[229] wl[37] vdd gnd cell_6t
Xbit_r38_c229 bl[229] br[229] wl[38] vdd gnd cell_6t
Xbit_r39_c229 bl[229] br[229] wl[39] vdd gnd cell_6t
Xbit_r40_c229 bl[229] br[229] wl[40] vdd gnd cell_6t
Xbit_r41_c229 bl[229] br[229] wl[41] vdd gnd cell_6t
Xbit_r42_c229 bl[229] br[229] wl[42] vdd gnd cell_6t
Xbit_r43_c229 bl[229] br[229] wl[43] vdd gnd cell_6t
Xbit_r44_c229 bl[229] br[229] wl[44] vdd gnd cell_6t
Xbit_r45_c229 bl[229] br[229] wl[45] vdd gnd cell_6t
Xbit_r46_c229 bl[229] br[229] wl[46] vdd gnd cell_6t
Xbit_r47_c229 bl[229] br[229] wl[47] vdd gnd cell_6t
Xbit_r48_c229 bl[229] br[229] wl[48] vdd gnd cell_6t
Xbit_r49_c229 bl[229] br[229] wl[49] vdd gnd cell_6t
Xbit_r50_c229 bl[229] br[229] wl[50] vdd gnd cell_6t
Xbit_r51_c229 bl[229] br[229] wl[51] vdd gnd cell_6t
Xbit_r52_c229 bl[229] br[229] wl[52] vdd gnd cell_6t
Xbit_r53_c229 bl[229] br[229] wl[53] vdd gnd cell_6t
Xbit_r54_c229 bl[229] br[229] wl[54] vdd gnd cell_6t
Xbit_r55_c229 bl[229] br[229] wl[55] vdd gnd cell_6t
Xbit_r56_c229 bl[229] br[229] wl[56] vdd gnd cell_6t
Xbit_r57_c229 bl[229] br[229] wl[57] vdd gnd cell_6t
Xbit_r58_c229 bl[229] br[229] wl[58] vdd gnd cell_6t
Xbit_r59_c229 bl[229] br[229] wl[59] vdd gnd cell_6t
Xbit_r60_c229 bl[229] br[229] wl[60] vdd gnd cell_6t
Xbit_r61_c229 bl[229] br[229] wl[61] vdd gnd cell_6t
Xbit_r62_c229 bl[229] br[229] wl[62] vdd gnd cell_6t
Xbit_r63_c229 bl[229] br[229] wl[63] vdd gnd cell_6t
Xbit_r64_c229 bl[229] br[229] wl[64] vdd gnd cell_6t
Xbit_r65_c229 bl[229] br[229] wl[65] vdd gnd cell_6t
Xbit_r66_c229 bl[229] br[229] wl[66] vdd gnd cell_6t
Xbit_r67_c229 bl[229] br[229] wl[67] vdd gnd cell_6t
Xbit_r68_c229 bl[229] br[229] wl[68] vdd gnd cell_6t
Xbit_r69_c229 bl[229] br[229] wl[69] vdd gnd cell_6t
Xbit_r70_c229 bl[229] br[229] wl[70] vdd gnd cell_6t
Xbit_r71_c229 bl[229] br[229] wl[71] vdd gnd cell_6t
Xbit_r72_c229 bl[229] br[229] wl[72] vdd gnd cell_6t
Xbit_r73_c229 bl[229] br[229] wl[73] vdd gnd cell_6t
Xbit_r74_c229 bl[229] br[229] wl[74] vdd gnd cell_6t
Xbit_r75_c229 bl[229] br[229] wl[75] vdd gnd cell_6t
Xbit_r76_c229 bl[229] br[229] wl[76] vdd gnd cell_6t
Xbit_r77_c229 bl[229] br[229] wl[77] vdd gnd cell_6t
Xbit_r78_c229 bl[229] br[229] wl[78] vdd gnd cell_6t
Xbit_r79_c229 bl[229] br[229] wl[79] vdd gnd cell_6t
Xbit_r80_c229 bl[229] br[229] wl[80] vdd gnd cell_6t
Xbit_r81_c229 bl[229] br[229] wl[81] vdd gnd cell_6t
Xbit_r82_c229 bl[229] br[229] wl[82] vdd gnd cell_6t
Xbit_r83_c229 bl[229] br[229] wl[83] vdd gnd cell_6t
Xbit_r84_c229 bl[229] br[229] wl[84] vdd gnd cell_6t
Xbit_r85_c229 bl[229] br[229] wl[85] vdd gnd cell_6t
Xbit_r86_c229 bl[229] br[229] wl[86] vdd gnd cell_6t
Xbit_r87_c229 bl[229] br[229] wl[87] vdd gnd cell_6t
Xbit_r88_c229 bl[229] br[229] wl[88] vdd gnd cell_6t
Xbit_r89_c229 bl[229] br[229] wl[89] vdd gnd cell_6t
Xbit_r90_c229 bl[229] br[229] wl[90] vdd gnd cell_6t
Xbit_r91_c229 bl[229] br[229] wl[91] vdd gnd cell_6t
Xbit_r92_c229 bl[229] br[229] wl[92] vdd gnd cell_6t
Xbit_r93_c229 bl[229] br[229] wl[93] vdd gnd cell_6t
Xbit_r94_c229 bl[229] br[229] wl[94] vdd gnd cell_6t
Xbit_r95_c229 bl[229] br[229] wl[95] vdd gnd cell_6t
Xbit_r96_c229 bl[229] br[229] wl[96] vdd gnd cell_6t
Xbit_r97_c229 bl[229] br[229] wl[97] vdd gnd cell_6t
Xbit_r98_c229 bl[229] br[229] wl[98] vdd gnd cell_6t
Xbit_r99_c229 bl[229] br[229] wl[99] vdd gnd cell_6t
Xbit_r100_c229 bl[229] br[229] wl[100] vdd gnd cell_6t
Xbit_r101_c229 bl[229] br[229] wl[101] vdd gnd cell_6t
Xbit_r102_c229 bl[229] br[229] wl[102] vdd gnd cell_6t
Xbit_r103_c229 bl[229] br[229] wl[103] vdd gnd cell_6t
Xbit_r104_c229 bl[229] br[229] wl[104] vdd gnd cell_6t
Xbit_r105_c229 bl[229] br[229] wl[105] vdd gnd cell_6t
Xbit_r106_c229 bl[229] br[229] wl[106] vdd gnd cell_6t
Xbit_r107_c229 bl[229] br[229] wl[107] vdd gnd cell_6t
Xbit_r108_c229 bl[229] br[229] wl[108] vdd gnd cell_6t
Xbit_r109_c229 bl[229] br[229] wl[109] vdd gnd cell_6t
Xbit_r110_c229 bl[229] br[229] wl[110] vdd gnd cell_6t
Xbit_r111_c229 bl[229] br[229] wl[111] vdd gnd cell_6t
Xbit_r112_c229 bl[229] br[229] wl[112] vdd gnd cell_6t
Xbit_r113_c229 bl[229] br[229] wl[113] vdd gnd cell_6t
Xbit_r114_c229 bl[229] br[229] wl[114] vdd gnd cell_6t
Xbit_r115_c229 bl[229] br[229] wl[115] vdd gnd cell_6t
Xbit_r116_c229 bl[229] br[229] wl[116] vdd gnd cell_6t
Xbit_r117_c229 bl[229] br[229] wl[117] vdd gnd cell_6t
Xbit_r118_c229 bl[229] br[229] wl[118] vdd gnd cell_6t
Xbit_r119_c229 bl[229] br[229] wl[119] vdd gnd cell_6t
Xbit_r120_c229 bl[229] br[229] wl[120] vdd gnd cell_6t
Xbit_r121_c229 bl[229] br[229] wl[121] vdd gnd cell_6t
Xbit_r122_c229 bl[229] br[229] wl[122] vdd gnd cell_6t
Xbit_r123_c229 bl[229] br[229] wl[123] vdd gnd cell_6t
Xbit_r124_c229 bl[229] br[229] wl[124] vdd gnd cell_6t
Xbit_r125_c229 bl[229] br[229] wl[125] vdd gnd cell_6t
Xbit_r126_c229 bl[229] br[229] wl[126] vdd gnd cell_6t
Xbit_r127_c229 bl[229] br[229] wl[127] vdd gnd cell_6t
Xbit_r128_c229 bl[229] br[229] wl[128] vdd gnd cell_6t
Xbit_r129_c229 bl[229] br[229] wl[129] vdd gnd cell_6t
Xbit_r130_c229 bl[229] br[229] wl[130] vdd gnd cell_6t
Xbit_r131_c229 bl[229] br[229] wl[131] vdd gnd cell_6t
Xbit_r132_c229 bl[229] br[229] wl[132] vdd gnd cell_6t
Xbit_r133_c229 bl[229] br[229] wl[133] vdd gnd cell_6t
Xbit_r134_c229 bl[229] br[229] wl[134] vdd gnd cell_6t
Xbit_r135_c229 bl[229] br[229] wl[135] vdd gnd cell_6t
Xbit_r136_c229 bl[229] br[229] wl[136] vdd gnd cell_6t
Xbit_r137_c229 bl[229] br[229] wl[137] vdd gnd cell_6t
Xbit_r138_c229 bl[229] br[229] wl[138] vdd gnd cell_6t
Xbit_r139_c229 bl[229] br[229] wl[139] vdd gnd cell_6t
Xbit_r140_c229 bl[229] br[229] wl[140] vdd gnd cell_6t
Xbit_r141_c229 bl[229] br[229] wl[141] vdd gnd cell_6t
Xbit_r142_c229 bl[229] br[229] wl[142] vdd gnd cell_6t
Xbit_r143_c229 bl[229] br[229] wl[143] vdd gnd cell_6t
Xbit_r144_c229 bl[229] br[229] wl[144] vdd gnd cell_6t
Xbit_r145_c229 bl[229] br[229] wl[145] vdd gnd cell_6t
Xbit_r146_c229 bl[229] br[229] wl[146] vdd gnd cell_6t
Xbit_r147_c229 bl[229] br[229] wl[147] vdd gnd cell_6t
Xbit_r148_c229 bl[229] br[229] wl[148] vdd gnd cell_6t
Xbit_r149_c229 bl[229] br[229] wl[149] vdd gnd cell_6t
Xbit_r150_c229 bl[229] br[229] wl[150] vdd gnd cell_6t
Xbit_r151_c229 bl[229] br[229] wl[151] vdd gnd cell_6t
Xbit_r152_c229 bl[229] br[229] wl[152] vdd gnd cell_6t
Xbit_r153_c229 bl[229] br[229] wl[153] vdd gnd cell_6t
Xbit_r154_c229 bl[229] br[229] wl[154] vdd gnd cell_6t
Xbit_r155_c229 bl[229] br[229] wl[155] vdd gnd cell_6t
Xbit_r156_c229 bl[229] br[229] wl[156] vdd gnd cell_6t
Xbit_r157_c229 bl[229] br[229] wl[157] vdd gnd cell_6t
Xbit_r158_c229 bl[229] br[229] wl[158] vdd gnd cell_6t
Xbit_r159_c229 bl[229] br[229] wl[159] vdd gnd cell_6t
Xbit_r160_c229 bl[229] br[229] wl[160] vdd gnd cell_6t
Xbit_r161_c229 bl[229] br[229] wl[161] vdd gnd cell_6t
Xbit_r162_c229 bl[229] br[229] wl[162] vdd gnd cell_6t
Xbit_r163_c229 bl[229] br[229] wl[163] vdd gnd cell_6t
Xbit_r164_c229 bl[229] br[229] wl[164] vdd gnd cell_6t
Xbit_r165_c229 bl[229] br[229] wl[165] vdd gnd cell_6t
Xbit_r166_c229 bl[229] br[229] wl[166] vdd gnd cell_6t
Xbit_r167_c229 bl[229] br[229] wl[167] vdd gnd cell_6t
Xbit_r168_c229 bl[229] br[229] wl[168] vdd gnd cell_6t
Xbit_r169_c229 bl[229] br[229] wl[169] vdd gnd cell_6t
Xbit_r170_c229 bl[229] br[229] wl[170] vdd gnd cell_6t
Xbit_r171_c229 bl[229] br[229] wl[171] vdd gnd cell_6t
Xbit_r172_c229 bl[229] br[229] wl[172] vdd gnd cell_6t
Xbit_r173_c229 bl[229] br[229] wl[173] vdd gnd cell_6t
Xbit_r174_c229 bl[229] br[229] wl[174] vdd gnd cell_6t
Xbit_r175_c229 bl[229] br[229] wl[175] vdd gnd cell_6t
Xbit_r176_c229 bl[229] br[229] wl[176] vdd gnd cell_6t
Xbit_r177_c229 bl[229] br[229] wl[177] vdd gnd cell_6t
Xbit_r178_c229 bl[229] br[229] wl[178] vdd gnd cell_6t
Xbit_r179_c229 bl[229] br[229] wl[179] vdd gnd cell_6t
Xbit_r180_c229 bl[229] br[229] wl[180] vdd gnd cell_6t
Xbit_r181_c229 bl[229] br[229] wl[181] vdd gnd cell_6t
Xbit_r182_c229 bl[229] br[229] wl[182] vdd gnd cell_6t
Xbit_r183_c229 bl[229] br[229] wl[183] vdd gnd cell_6t
Xbit_r184_c229 bl[229] br[229] wl[184] vdd gnd cell_6t
Xbit_r185_c229 bl[229] br[229] wl[185] vdd gnd cell_6t
Xbit_r186_c229 bl[229] br[229] wl[186] vdd gnd cell_6t
Xbit_r187_c229 bl[229] br[229] wl[187] vdd gnd cell_6t
Xbit_r188_c229 bl[229] br[229] wl[188] vdd gnd cell_6t
Xbit_r189_c229 bl[229] br[229] wl[189] vdd gnd cell_6t
Xbit_r190_c229 bl[229] br[229] wl[190] vdd gnd cell_6t
Xbit_r191_c229 bl[229] br[229] wl[191] vdd gnd cell_6t
Xbit_r192_c229 bl[229] br[229] wl[192] vdd gnd cell_6t
Xbit_r193_c229 bl[229] br[229] wl[193] vdd gnd cell_6t
Xbit_r194_c229 bl[229] br[229] wl[194] vdd gnd cell_6t
Xbit_r195_c229 bl[229] br[229] wl[195] vdd gnd cell_6t
Xbit_r196_c229 bl[229] br[229] wl[196] vdd gnd cell_6t
Xbit_r197_c229 bl[229] br[229] wl[197] vdd gnd cell_6t
Xbit_r198_c229 bl[229] br[229] wl[198] vdd gnd cell_6t
Xbit_r199_c229 bl[229] br[229] wl[199] vdd gnd cell_6t
Xbit_r200_c229 bl[229] br[229] wl[200] vdd gnd cell_6t
Xbit_r201_c229 bl[229] br[229] wl[201] vdd gnd cell_6t
Xbit_r202_c229 bl[229] br[229] wl[202] vdd gnd cell_6t
Xbit_r203_c229 bl[229] br[229] wl[203] vdd gnd cell_6t
Xbit_r204_c229 bl[229] br[229] wl[204] vdd gnd cell_6t
Xbit_r205_c229 bl[229] br[229] wl[205] vdd gnd cell_6t
Xbit_r206_c229 bl[229] br[229] wl[206] vdd gnd cell_6t
Xbit_r207_c229 bl[229] br[229] wl[207] vdd gnd cell_6t
Xbit_r208_c229 bl[229] br[229] wl[208] vdd gnd cell_6t
Xbit_r209_c229 bl[229] br[229] wl[209] vdd gnd cell_6t
Xbit_r210_c229 bl[229] br[229] wl[210] vdd gnd cell_6t
Xbit_r211_c229 bl[229] br[229] wl[211] vdd gnd cell_6t
Xbit_r212_c229 bl[229] br[229] wl[212] vdd gnd cell_6t
Xbit_r213_c229 bl[229] br[229] wl[213] vdd gnd cell_6t
Xbit_r214_c229 bl[229] br[229] wl[214] vdd gnd cell_6t
Xbit_r215_c229 bl[229] br[229] wl[215] vdd gnd cell_6t
Xbit_r216_c229 bl[229] br[229] wl[216] vdd gnd cell_6t
Xbit_r217_c229 bl[229] br[229] wl[217] vdd gnd cell_6t
Xbit_r218_c229 bl[229] br[229] wl[218] vdd gnd cell_6t
Xbit_r219_c229 bl[229] br[229] wl[219] vdd gnd cell_6t
Xbit_r220_c229 bl[229] br[229] wl[220] vdd gnd cell_6t
Xbit_r221_c229 bl[229] br[229] wl[221] vdd gnd cell_6t
Xbit_r222_c229 bl[229] br[229] wl[222] vdd gnd cell_6t
Xbit_r223_c229 bl[229] br[229] wl[223] vdd gnd cell_6t
Xbit_r224_c229 bl[229] br[229] wl[224] vdd gnd cell_6t
Xbit_r225_c229 bl[229] br[229] wl[225] vdd gnd cell_6t
Xbit_r226_c229 bl[229] br[229] wl[226] vdd gnd cell_6t
Xbit_r227_c229 bl[229] br[229] wl[227] vdd gnd cell_6t
Xbit_r228_c229 bl[229] br[229] wl[228] vdd gnd cell_6t
Xbit_r229_c229 bl[229] br[229] wl[229] vdd gnd cell_6t
Xbit_r230_c229 bl[229] br[229] wl[230] vdd gnd cell_6t
Xbit_r231_c229 bl[229] br[229] wl[231] vdd gnd cell_6t
Xbit_r232_c229 bl[229] br[229] wl[232] vdd gnd cell_6t
Xbit_r233_c229 bl[229] br[229] wl[233] vdd gnd cell_6t
Xbit_r234_c229 bl[229] br[229] wl[234] vdd gnd cell_6t
Xbit_r235_c229 bl[229] br[229] wl[235] vdd gnd cell_6t
Xbit_r236_c229 bl[229] br[229] wl[236] vdd gnd cell_6t
Xbit_r237_c229 bl[229] br[229] wl[237] vdd gnd cell_6t
Xbit_r238_c229 bl[229] br[229] wl[238] vdd gnd cell_6t
Xbit_r239_c229 bl[229] br[229] wl[239] vdd gnd cell_6t
Xbit_r240_c229 bl[229] br[229] wl[240] vdd gnd cell_6t
Xbit_r241_c229 bl[229] br[229] wl[241] vdd gnd cell_6t
Xbit_r242_c229 bl[229] br[229] wl[242] vdd gnd cell_6t
Xbit_r243_c229 bl[229] br[229] wl[243] vdd gnd cell_6t
Xbit_r244_c229 bl[229] br[229] wl[244] vdd gnd cell_6t
Xbit_r245_c229 bl[229] br[229] wl[245] vdd gnd cell_6t
Xbit_r246_c229 bl[229] br[229] wl[246] vdd gnd cell_6t
Xbit_r247_c229 bl[229] br[229] wl[247] vdd gnd cell_6t
Xbit_r248_c229 bl[229] br[229] wl[248] vdd gnd cell_6t
Xbit_r249_c229 bl[229] br[229] wl[249] vdd gnd cell_6t
Xbit_r250_c229 bl[229] br[229] wl[250] vdd gnd cell_6t
Xbit_r251_c229 bl[229] br[229] wl[251] vdd gnd cell_6t
Xbit_r252_c229 bl[229] br[229] wl[252] vdd gnd cell_6t
Xbit_r253_c229 bl[229] br[229] wl[253] vdd gnd cell_6t
Xbit_r254_c229 bl[229] br[229] wl[254] vdd gnd cell_6t
Xbit_r255_c229 bl[229] br[229] wl[255] vdd gnd cell_6t
Xbit_r0_c230 bl[230] br[230] wl[0] vdd gnd cell_6t
Xbit_r1_c230 bl[230] br[230] wl[1] vdd gnd cell_6t
Xbit_r2_c230 bl[230] br[230] wl[2] vdd gnd cell_6t
Xbit_r3_c230 bl[230] br[230] wl[3] vdd gnd cell_6t
Xbit_r4_c230 bl[230] br[230] wl[4] vdd gnd cell_6t
Xbit_r5_c230 bl[230] br[230] wl[5] vdd gnd cell_6t
Xbit_r6_c230 bl[230] br[230] wl[6] vdd gnd cell_6t
Xbit_r7_c230 bl[230] br[230] wl[7] vdd gnd cell_6t
Xbit_r8_c230 bl[230] br[230] wl[8] vdd gnd cell_6t
Xbit_r9_c230 bl[230] br[230] wl[9] vdd gnd cell_6t
Xbit_r10_c230 bl[230] br[230] wl[10] vdd gnd cell_6t
Xbit_r11_c230 bl[230] br[230] wl[11] vdd gnd cell_6t
Xbit_r12_c230 bl[230] br[230] wl[12] vdd gnd cell_6t
Xbit_r13_c230 bl[230] br[230] wl[13] vdd gnd cell_6t
Xbit_r14_c230 bl[230] br[230] wl[14] vdd gnd cell_6t
Xbit_r15_c230 bl[230] br[230] wl[15] vdd gnd cell_6t
Xbit_r16_c230 bl[230] br[230] wl[16] vdd gnd cell_6t
Xbit_r17_c230 bl[230] br[230] wl[17] vdd gnd cell_6t
Xbit_r18_c230 bl[230] br[230] wl[18] vdd gnd cell_6t
Xbit_r19_c230 bl[230] br[230] wl[19] vdd gnd cell_6t
Xbit_r20_c230 bl[230] br[230] wl[20] vdd gnd cell_6t
Xbit_r21_c230 bl[230] br[230] wl[21] vdd gnd cell_6t
Xbit_r22_c230 bl[230] br[230] wl[22] vdd gnd cell_6t
Xbit_r23_c230 bl[230] br[230] wl[23] vdd gnd cell_6t
Xbit_r24_c230 bl[230] br[230] wl[24] vdd gnd cell_6t
Xbit_r25_c230 bl[230] br[230] wl[25] vdd gnd cell_6t
Xbit_r26_c230 bl[230] br[230] wl[26] vdd gnd cell_6t
Xbit_r27_c230 bl[230] br[230] wl[27] vdd gnd cell_6t
Xbit_r28_c230 bl[230] br[230] wl[28] vdd gnd cell_6t
Xbit_r29_c230 bl[230] br[230] wl[29] vdd gnd cell_6t
Xbit_r30_c230 bl[230] br[230] wl[30] vdd gnd cell_6t
Xbit_r31_c230 bl[230] br[230] wl[31] vdd gnd cell_6t
Xbit_r32_c230 bl[230] br[230] wl[32] vdd gnd cell_6t
Xbit_r33_c230 bl[230] br[230] wl[33] vdd gnd cell_6t
Xbit_r34_c230 bl[230] br[230] wl[34] vdd gnd cell_6t
Xbit_r35_c230 bl[230] br[230] wl[35] vdd gnd cell_6t
Xbit_r36_c230 bl[230] br[230] wl[36] vdd gnd cell_6t
Xbit_r37_c230 bl[230] br[230] wl[37] vdd gnd cell_6t
Xbit_r38_c230 bl[230] br[230] wl[38] vdd gnd cell_6t
Xbit_r39_c230 bl[230] br[230] wl[39] vdd gnd cell_6t
Xbit_r40_c230 bl[230] br[230] wl[40] vdd gnd cell_6t
Xbit_r41_c230 bl[230] br[230] wl[41] vdd gnd cell_6t
Xbit_r42_c230 bl[230] br[230] wl[42] vdd gnd cell_6t
Xbit_r43_c230 bl[230] br[230] wl[43] vdd gnd cell_6t
Xbit_r44_c230 bl[230] br[230] wl[44] vdd gnd cell_6t
Xbit_r45_c230 bl[230] br[230] wl[45] vdd gnd cell_6t
Xbit_r46_c230 bl[230] br[230] wl[46] vdd gnd cell_6t
Xbit_r47_c230 bl[230] br[230] wl[47] vdd gnd cell_6t
Xbit_r48_c230 bl[230] br[230] wl[48] vdd gnd cell_6t
Xbit_r49_c230 bl[230] br[230] wl[49] vdd gnd cell_6t
Xbit_r50_c230 bl[230] br[230] wl[50] vdd gnd cell_6t
Xbit_r51_c230 bl[230] br[230] wl[51] vdd gnd cell_6t
Xbit_r52_c230 bl[230] br[230] wl[52] vdd gnd cell_6t
Xbit_r53_c230 bl[230] br[230] wl[53] vdd gnd cell_6t
Xbit_r54_c230 bl[230] br[230] wl[54] vdd gnd cell_6t
Xbit_r55_c230 bl[230] br[230] wl[55] vdd gnd cell_6t
Xbit_r56_c230 bl[230] br[230] wl[56] vdd gnd cell_6t
Xbit_r57_c230 bl[230] br[230] wl[57] vdd gnd cell_6t
Xbit_r58_c230 bl[230] br[230] wl[58] vdd gnd cell_6t
Xbit_r59_c230 bl[230] br[230] wl[59] vdd gnd cell_6t
Xbit_r60_c230 bl[230] br[230] wl[60] vdd gnd cell_6t
Xbit_r61_c230 bl[230] br[230] wl[61] vdd gnd cell_6t
Xbit_r62_c230 bl[230] br[230] wl[62] vdd gnd cell_6t
Xbit_r63_c230 bl[230] br[230] wl[63] vdd gnd cell_6t
Xbit_r64_c230 bl[230] br[230] wl[64] vdd gnd cell_6t
Xbit_r65_c230 bl[230] br[230] wl[65] vdd gnd cell_6t
Xbit_r66_c230 bl[230] br[230] wl[66] vdd gnd cell_6t
Xbit_r67_c230 bl[230] br[230] wl[67] vdd gnd cell_6t
Xbit_r68_c230 bl[230] br[230] wl[68] vdd gnd cell_6t
Xbit_r69_c230 bl[230] br[230] wl[69] vdd gnd cell_6t
Xbit_r70_c230 bl[230] br[230] wl[70] vdd gnd cell_6t
Xbit_r71_c230 bl[230] br[230] wl[71] vdd gnd cell_6t
Xbit_r72_c230 bl[230] br[230] wl[72] vdd gnd cell_6t
Xbit_r73_c230 bl[230] br[230] wl[73] vdd gnd cell_6t
Xbit_r74_c230 bl[230] br[230] wl[74] vdd gnd cell_6t
Xbit_r75_c230 bl[230] br[230] wl[75] vdd gnd cell_6t
Xbit_r76_c230 bl[230] br[230] wl[76] vdd gnd cell_6t
Xbit_r77_c230 bl[230] br[230] wl[77] vdd gnd cell_6t
Xbit_r78_c230 bl[230] br[230] wl[78] vdd gnd cell_6t
Xbit_r79_c230 bl[230] br[230] wl[79] vdd gnd cell_6t
Xbit_r80_c230 bl[230] br[230] wl[80] vdd gnd cell_6t
Xbit_r81_c230 bl[230] br[230] wl[81] vdd gnd cell_6t
Xbit_r82_c230 bl[230] br[230] wl[82] vdd gnd cell_6t
Xbit_r83_c230 bl[230] br[230] wl[83] vdd gnd cell_6t
Xbit_r84_c230 bl[230] br[230] wl[84] vdd gnd cell_6t
Xbit_r85_c230 bl[230] br[230] wl[85] vdd gnd cell_6t
Xbit_r86_c230 bl[230] br[230] wl[86] vdd gnd cell_6t
Xbit_r87_c230 bl[230] br[230] wl[87] vdd gnd cell_6t
Xbit_r88_c230 bl[230] br[230] wl[88] vdd gnd cell_6t
Xbit_r89_c230 bl[230] br[230] wl[89] vdd gnd cell_6t
Xbit_r90_c230 bl[230] br[230] wl[90] vdd gnd cell_6t
Xbit_r91_c230 bl[230] br[230] wl[91] vdd gnd cell_6t
Xbit_r92_c230 bl[230] br[230] wl[92] vdd gnd cell_6t
Xbit_r93_c230 bl[230] br[230] wl[93] vdd gnd cell_6t
Xbit_r94_c230 bl[230] br[230] wl[94] vdd gnd cell_6t
Xbit_r95_c230 bl[230] br[230] wl[95] vdd gnd cell_6t
Xbit_r96_c230 bl[230] br[230] wl[96] vdd gnd cell_6t
Xbit_r97_c230 bl[230] br[230] wl[97] vdd gnd cell_6t
Xbit_r98_c230 bl[230] br[230] wl[98] vdd gnd cell_6t
Xbit_r99_c230 bl[230] br[230] wl[99] vdd gnd cell_6t
Xbit_r100_c230 bl[230] br[230] wl[100] vdd gnd cell_6t
Xbit_r101_c230 bl[230] br[230] wl[101] vdd gnd cell_6t
Xbit_r102_c230 bl[230] br[230] wl[102] vdd gnd cell_6t
Xbit_r103_c230 bl[230] br[230] wl[103] vdd gnd cell_6t
Xbit_r104_c230 bl[230] br[230] wl[104] vdd gnd cell_6t
Xbit_r105_c230 bl[230] br[230] wl[105] vdd gnd cell_6t
Xbit_r106_c230 bl[230] br[230] wl[106] vdd gnd cell_6t
Xbit_r107_c230 bl[230] br[230] wl[107] vdd gnd cell_6t
Xbit_r108_c230 bl[230] br[230] wl[108] vdd gnd cell_6t
Xbit_r109_c230 bl[230] br[230] wl[109] vdd gnd cell_6t
Xbit_r110_c230 bl[230] br[230] wl[110] vdd gnd cell_6t
Xbit_r111_c230 bl[230] br[230] wl[111] vdd gnd cell_6t
Xbit_r112_c230 bl[230] br[230] wl[112] vdd gnd cell_6t
Xbit_r113_c230 bl[230] br[230] wl[113] vdd gnd cell_6t
Xbit_r114_c230 bl[230] br[230] wl[114] vdd gnd cell_6t
Xbit_r115_c230 bl[230] br[230] wl[115] vdd gnd cell_6t
Xbit_r116_c230 bl[230] br[230] wl[116] vdd gnd cell_6t
Xbit_r117_c230 bl[230] br[230] wl[117] vdd gnd cell_6t
Xbit_r118_c230 bl[230] br[230] wl[118] vdd gnd cell_6t
Xbit_r119_c230 bl[230] br[230] wl[119] vdd gnd cell_6t
Xbit_r120_c230 bl[230] br[230] wl[120] vdd gnd cell_6t
Xbit_r121_c230 bl[230] br[230] wl[121] vdd gnd cell_6t
Xbit_r122_c230 bl[230] br[230] wl[122] vdd gnd cell_6t
Xbit_r123_c230 bl[230] br[230] wl[123] vdd gnd cell_6t
Xbit_r124_c230 bl[230] br[230] wl[124] vdd gnd cell_6t
Xbit_r125_c230 bl[230] br[230] wl[125] vdd gnd cell_6t
Xbit_r126_c230 bl[230] br[230] wl[126] vdd gnd cell_6t
Xbit_r127_c230 bl[230] br[230] wl[127] vdd gnd cell_6t
Xbit_r128_c230 bl[230] br[230] wl[128] vdd gnd cell_6t
Xbit_r129_c230 bl[230] br[230] wl[129] vdd gnd cell_6t
Xbit_r130_c230 bl[230] br[230] wl[130] vdd gnd cell_6t
Xbit_r131_c230 bl[230] br[230] wl[131] vdd gnd cell_6t
Xbit_r132_c230 bl[230] br[230] wl[132] vdd gnd cell_6t
Xbit_r133_c230 bl[230] br[230] wl[133] vdd gnd cell_6t
Xbit_r134_c230 bl[230] br[230] wl[134] vdd gnd cell_6t
Xbit_r135_c230 bl[230] br[230] wl[135] vdd gnd cell_6t
Xbit_r136_c230 bl[230] br[230] wl[136] vdd gnd cell_6t
Xbit_r137_c230 bl[230] br[230] wl[137] vdd gnd cell_6t
Xbit_r138_c230 bl[230] br[230] wl[138] vdd gnd cell_6t
Xbit_r139_c230 bl[230] br[230] wl[139] vdd gnd cell_6t
Xbit_r140_c230 bl[230] br[230] wl[140] vdd gnd cell_6t
Xbit_r141_c230 bl[230] br[230] wl[141] vdd gnd cell_6t
Xbit_r142_c230 bl[230] br[230] wl[142] vdd gnd cell_6t
Xbit_r143_c230 bl[230] br[230] wl[143] vdd gnd cell_6t
Xbit_r144_c230 bl[230] br[230] wl[144] vdd gnd cell_6t
Xbit_r145_c230 bl[230] br[230] wl[145] vdd gnd cell_6t
Xbit_r146_c230 bl[230] br[230] wl[146] vdd gnd cell_6t
Xbit_r147_c230 bl[230] br[230] wl[147] vdd gnd cell_6t
Xbit_r148_c230 bl[230] br[230] wl[148] vdd gnd cell_6t
Xbit_r149_c230 bl[230] br[230] wl[149] vdd gnd cell_6t
Xbit_r150_c230 bl[230] br[230] wl[150] vdd gnd cell_6t
Xbit_r151_c230 bl[230] br[230] wl[151] vdd gnd cell_6t
Xbit_r152_c230 bl[230] br[230] wl[152] vdd gnd cell_6t
Xbit_r153_c230 bl[230] br[230] wl[153] vdd gnd cell_6t
Xbit_r154_c230 bl[230] br[230] wl[154] vdd gnd cell_6t
Xbit_r155_c230 bl[230] br[230] wl[155] vdd gnd cell_6t
Xbit_r156_c230 bl[230] br[230] wl[156] vdd gnd cell_6t
Xbit_r157_c230 bl[230] br[230] wl[157] vdd gnd cell_6t
Xbit_r158_c230 bl[230] br[230] wl[158] vdd gnd cell_6t
Xbit_r159_c230 bl[230] br[230] wl[159] vdd gnd cell_6t
Xbit_r160_c230 bl[230] br[230] wl[160] vdd gnd cell_6t
Xbit_r161_c230 bl[230] br[230] wl[161] vdd gnd cell_6t
Xbit_r162_c230 bl[230] br[230] wl[162] vdd gnd cell_6t
Xbit_r163_c230 bl[230] br[230] wl[163] vdd gnd cell_6t
Xbit_r164_c230 bl[230] br[230] wl[164] vdd gnd cell_6t
Xbit_r165_c230 bl[230] br[230] wl[165] vdd gnd cell_6t
Xbit_r166_c230 bl[230] br[230] wl[166] vdd gnd cell_6t
Xbit_r167_c230 bl[230] br[230] wl[167] vdd gnd cell_6t
Xbit_r168_c230 bl[230] br[230] wl[168] vdd gnd cell_6t
Xbit_r169_c230 bl[230] br[230] wl[169] vdd gnd cell_6t
Xbit_r170_c230 bl[230] br[230] wl[170] vdd gnd cell_6t
Xbit_r171_c230 bl[230] br[230] wl[171] vdd gnd cell_6t
Xbit_r172_c230 bl[230] br[230] wl[172] vdd gnd cell_6t
Xbit_r173_c230 bl[230] br[230] wl[173] vdd gnd cell_6t
Xbit_r174_c230 bl[230] br[230] wl[174] vdd gnd cell_6t
Xbit_r175_c230 bl[230] br[230] wl[175] vdd gnd cell_6t
Xbit_r176_c230 bl[230] br[230] wl[176] vdd gnd cell_6t
Xbit_r177_c230 bl[230] br[230] wl[177] vdd gnd cell_6t
Xbit_r178_c230 bl[230] br[230] wl[178] vdd gnd cell_6t
Xbit_r179_c230 bl[230] br[230] wl[179] vdd gnd cell_6t
Xbit_r180_c230 bl[230] br[230] wl[180] vdd gnd cell_6t
Xbit_r181_c230 bl[230] br[230] wl[181] vdd gnd cell_6t
Xbit_r182_c230 bl[230] br[230] wl[182] vdd gnd cell_6t
Xbit_r183_c230 bl[230] br[230] wl[183] vdd gnd cell_6t
Xbit_r184_c230 bl[230] br[230] wl[184] vdd gnd cell_6t
Xbit_r185_c230 bl[230] br[230] wl[185] vdd gnd cell_6t
Xbit_r186_c230 bl[230] br[230] wl[186] vdd gnd cell_6t
Xbit_r187_c230 bl[230] br[230] wl[187] vdd gnd cell_6t
Xbit_r188_c230 bl[230] br[230] wl[188] vdd gnd cell_6t
Xbit_r189_c230 bl[230] br[230] wl[189] vdd gnd cell_6t
Xbit_r190_c230 bl[230] br[230] wl[190] vdd gnd cell_6t
Xbit_r191_c230 bl[230] br[230] wl[191] vdd gnd cell_6t
Xbit_r192_c230 bl[230] br[230] wl[192] vdd gnd cell_6t
Xbit_r193_c230 bl[230] br[230] wl[193] vdd gnd cell_6t
Xbit_r194_c230 bl[230] br[230] wl[194] vdd gnd cell_6t
Xbit_r195_c230 bl[230] br[230] wl[195] vdd gnd cell_6t
Xbit_r196_c230 bl[230] br[230] wl[196] vdd gnd cell_6t
Xbit_r197_c230 bl[230] br[230] wl[197] vdd gnd cell_6t
Xbit_r198_c230 bl[230] br[230] wl[198] vdd gnd cell_6t
Xbit_r199_c230 bl[230] br[230] wl[199] vdd gnd cell_6t
Xbit_r200_c230 bl[230] br[230] wl[200] vdd gnd cell_6t
Xbit_r201_c230 bl[230] br[230] wl[201] vdd gnd cell_6t
Xbit_r202_c230 bl[230] br[230] wl[202] vdd gnd cell_6t
Xbit_r203_c230 bl[230] br[230] wl[203] vdd gnd cell_6t
Xbit_r204_c230 bl[230] br[230] wl[204] vdd gnd cell_6t
Xbit_r205_c230 bl[230] br[230] wl[205] vdd gnd cell_6t
Xbit_r206_c230 bl[230] br[230] wl[206] vdd gnd cell_6t
Xbit_r207_c230 bl[230] br[230] wl[207] vdd gnd cell_6t
Xbit_r208_c230 bl[230] br[230] wl[208] vdd gnd cell_6t
Xbit_r209_c230 bl[230] br[230] wl[209] vdd gnd cell_6t
Xbit_r210_c230 bl[230] br[230] wl[210] vdd gnd cell_6t
Xbit_r211_c230 bl[230] br[230] wl[211] vdd gnd cell_6t
Xbit_r212_c230 bl[230] br[230] wl[212] vdd gnd cell_6t
Xbit_r213_c230 bl[230] br[230] wl[213] vdd gnd cell_6t
Xbit_r214_c230 bl[230] br[230] wl[214] vdd gnd cell_6t
Xbit_r215_c230 bl[230] br[230] wl[215] vdd gnd cell_6t
Xbit_r216_c230 bl[230] br[230] wl[216] vdd gnd cell_6t
Xbit_r217_c230 bl[230] br[230] wl[217] vdd gnd cell_6t
Xbit_r218_c230 bl[230] br[230] wl[218] vdd gnd cell_6t
Xbit_r219_c230 bl[230] br[230] wl[219] vdd gnd cell_6t
Xbit_r220_c230 bl[230] br[230] wl[220] vdd gnd cell_6t
Xbit_r221_c230 bl[230] br[230] wl[221] vdd gnd cell_6t
Xbit_r222_c230 bl[230] br[230] wl[222] vdd gnd cell_6t
Xbit_r223_c230 bl[230] br[230] wl[223] vdd gnd cell_6t
Xbit_r224_c230 bl[230] br[230] wl[224] vdd gnd cell_6t
Xbit_r225_c230 bl[230] br[230] wl[225] vdd gnd cell_6t
Xbit_r226_c230 bl[230] br[230] wl[226] vdd gnd cell_6t
Xbit_r227_c230 bl[230] br[230] wl[227] vdd gnd cell_6t
Xbit_r228_c230 bl[230] br[230] wl[228] vdd gnd cell_6t
Xbit_r229_c230 bl[230] br[230] wl[229] vdd gnd cell_6t
Xbit_r230_c230 bl[230] br[230] wl[230] vdd gnd cell_6t
Xbit_r231_c230 bl[230] br[230] wl[231] vdd gnd cell_6t
Xbit_r232_c230 bl[230] br[230] wl[232] vdd gnd cell_6t
Xbit_r233_c230 bl[230] br[230] wl[233] vdd gnd cell_6t
Xbit_r234_c230 bl[230] br[230] wl[234] vdd gnd cell_6t
Xbit_r235_c230 bl[230] br[230] wl[235] vdd gnd cell_6t
Xbit_r236_c230 bl[230] br[230] wl[236] vdd gnd cell_6t
Xbit_r237_c230 bl[230] br[230] wl[237] vdd gnd cell_6t
Xbit_r238_c230 bl[230] br[230] wl[238] vdd gnd cell_6t
Xbit_r239_c230 bl[230] br[230] wl[239] vdd gnd cell_6t
Xbit_r240_c230 bl[230] br[230] wl[240] vdd gnd cell_6t
Xbit_r241_c230 bl[230] br[230] wl[241] vdd gnd cell_6t
Xbit_r242_c230 bl[230] br[230] wl[242] vdd gnd cell_6t
Xbit_r243_c230 bl[230] br[230] wl[243] vdd gnd cell_6t
Xbit_r244_c230 bl[230] br[230] wl[244] vdd gnd cell_6t
Xbit_r245_c230 bl[230] br[230] wl[245] vdd gnd cell_6t
Xbit_r246_c230 bl[230] br[230] wl[246] vdd gnd cell_6t
Xbit_r247_c230 bl[230] br[230] wl[247] vdd gnd cell_6t
Xbit_r248_c230 bl[230] br[230] wl[248] vdd gnd cell_6t
Xbit_r249_c230 bl[230] br[230] wl[249] vdd gnd cell_6t
Xbit_r250_c230 bl[230] br[230] wl[250] vdd gnd cell_6t
Xbit_r251_c230 bl[230] br[230] wl[251] vdd gnd cell_6t
Xbit_r252_c230 bl[230] br[230] wl[252] vdd gnd cell_6t
Xbit_r253_c230 bl[230] br[230] wl[253] vdd gnd cell_6t
Xbit_r254_c230 bl[230] br[230] wl[254] vdd gnd cell_6t
Xbit_r255_c230 bl[230] br[230] wl[255] vdd gnd cell_6t
Xbit_r0_c231 bl[231] br[231] wl[0] vdd gnd cell_6t
Xbit_r1_c231 bl[231] br[231] wl[1] vdd gnd cell_6t
Xbit_r2_c231 bl[231] br[231] wl[2] vdd gnd cell_6t
Xbit_r3_c231 bl[231] br[231] wl[3] vdd gnd cell_6t
Xbit_r4_c231 bl[231] br[231] wl[4] vdd gnd cell_6t
Xbit_r5_c231 bl[231] br[231] wl[5] vdd gnd cell_6t
Xbit_r6_c231 bl[231] br[231] wl[6] vdd gnd cell_6t
Xbit_r7_c231 bl[231] br[231] wl[7] vdd gnd cell_6t
Xbit_r8_c231 bl[231] br[231] wl[8] vdd gnd cell_6t
Xbit_r9_c231 bl[231] br[231] wl[9] vdd gnd cell_6t
Xbit_r10_c231 bl[231] br[231] wl[10] vdd gnd cell_6t
Xbit_r11_c231 bl[231] br[231] wl[11] vdd gnd cell_6t
Xbit_r12_c231 bl[231] br[231] wl[12] vdd gnd cell_6t
Xbit_r13_c231 bl[231] br[231] wl[13] vdd gnd cell_6t
Xbit_r14_c231 bl[231] br[231] wl[14] vdd gnd cell_6t
Xbit_r15_c231 bl[231] br[231] wl[15] vdd gnd cell_6t
Xbit_r16_c231 bl[231] br[231] wl[16] vdd gnd cell_6t
Xbit_r17_c231 bl[231] br[231] wl[17] vdd gnd cell_6t
Xbit_r18_c231 bl[231] br[231] wl[18] vdd gnd cell_6t
Xbit_r19_c231 bl[231] br[231] wl[19] vdd gnd cell_6t
Xbit_r20_c231 bl[231] br[231] wl[20] vdd gnd cell_6t
Xbit_r21_c231 bl[231] br[231] wl[21] vdd gnd cell_6t
Xbit_r22_c231 bl[231] br[231] wl[22] vdd gnd cell_6t
Xbit_r23_c231 bl[231] br[231] wl[23] vdd gnd cell_6t
Xbit_r24_c231 bl[231] br[231] wl[24] vdd gnd cell_6t
Xbit_r25_c231 bl[231] br[231] wl[25] vdd gnd cell_6t
Xbit_r26_c231 bl[231] br[231] wl[26] vdd gnd cell_6t
Xbit_r27_c231 bl[231] br[231] wl[27] vdd gnd cell_6t
Xbit_r28_c231 bl[231] br[231] wl[28] vdd gnd cell_6t
Xbit_r29_c231 bl[231] br[231] wl[29] vdd gnd cell_6t
Xbit_r30_c231 bl[231] br[231] wl[30] vdd gnd cell_6t
Xbit_r31_c231 bl[231] br[231] wl[31] vdd gnd cell_6t
Xbit_r32_c231 bl[231] br[231] wl[32] vdd gnd cell_6t
Xbit_r33_c231 bl[231] br[231] wl[33] vdd gnd cell_6t
Xbit_r34_c231 bl[231] br[231] wl[34] vdd gnd cell_6t
Xbit_r35_c231 bl[231] br[231] wl[35] vdd gnd cell_6t
Xbit_r36_c231 bl[231] br[231] wl[36] vdd gnd cell_6t
Xbit_r37_c231 bl[231] br[231] wl[37] vdd gnd cell_6t
Xbit_r38_c231 bl[231] br[231] wl[38] vdd gnd cell_6t
Xbit_r39_c231 bl[231] br[231] wl[39] vdd gnd cell_6t
Xbit_r40_c231 bl[231] br[231] wl[40] vdd gnd cell_6t
Xbit_r41_c231 bl[231] br[231] wl[41] vdd gnd cell_6t
Xbit_r42_c231 bl[231] br[231] wl[42] vdd gnd cell_6t
Xbit_r43_c231 bl[231] br[231] wl[43] vdd gnd cell_6t
Xbit_r44_c231 bl[231] br[231] wl[44] vdd gnd cell_6t
Xbit_r45_c231 bl[231] br[231] wl[45] vdd gnd cell_6t
Xbit_r46_c231 bl[231] br[231] wl[46] vdd gnd cell_6t
Xbit_r47_c231 bl[231] br[231] wl[47] vdd gnd cell_6t
Xbit_r48_c231 bl[231] br[231] wl[48] vdd gnd cell_6t
Xbit_r49_c231 bl[231] br[231] wl[49] vdd gnd cell_6t
Xbit_r50_c231 bl[231] br[231] wl[50] vdd gnd cell_6t
Xbit_r51_c231 bl[231] br[231] wl[51] vdd gnd cell_6t
Xbit_r52_c231 bl[231] br[231] wl[52] vdd gnd cell_6t
Xbit_r53_c231 bl[231] br[231] wl[53] vdd gnd cell_6t
Xbit_r54_c231 bl[231] br[231] wl[54] vdd gnd cell_6t
Xbit_r55_c231 bl[231] br[231] wl[55] vdd gnd cell_6t
Xbit_r56_c231 bl[231] br[231] wl[56] vdd gnd cell_6t
Xbit_r57_c231 bl[231] br[231] wl[57] vdd gnd cell_6t
Xbit_r58_c231 bl[231] br[231] wl[58] vdd gnd cell_6t
Xbit_r59_c231 bl[231] br[231] wl[59] vdd gnd cell_6t
Xbit_r60_c231 bl[231] br[231] wl[60] vdd gnd cell_6t
Xbit_r61_c231 bl[231] br[231] wl[61] vdd gnd cell_6t
Xbit_r62_c231 bl[231] br[231] wl[62] vdd gnd cell_6t
Xbit_r63_c231 bl[231] br[231] wl[63] vdd gnd cell_6t
Xbit_r64_c231 bl[231] br[231] wl[64] vdd gnd cell_6t
Xbit_r65_c231 bl[231] br[231] wl[65] vdd gnd cell_6t
Xbit_r66_c231 bl[231] br[231] wl[66] vdd gnd cell_6t
Xbit_r67_c231 bl[231] br[231] wl[67] vdd gnd cell_6t
Xbit_r68_c231 bl[231] br[231] wl[68] vdd gnd cell_6t
Xbit_r69_c231 bl[231] br[231] wl[69] vdd gnd cell_6t
Xbit_r70_c231 bl[231] br[231] wl[70] vdd gnd cell_6t
Xbit_r71_c231 bl[231] br[231] wl[71] vdd gnd cell_6t
Xbit_r72_c231 bl[231] br[231] wl[72] vdd gnd cell_6t
Xbit_r73_c231 bl[231] br[231] wl[73] vdd gnd cell_6t
Xbit_r74_c231 bl[231] br[231] wl[74] vdd gnd cell_6t
Xbit_r75_c231 bl[231] br[231] wl[75] vdd gnd cell_6t
Xbit_r76_c231 bl[231] br[231] wl[76] vdd gnd cell_6t
Xbit_r77_c231 bl[231] br[231] wl[77] vdd gnd cell_6t
Xbit_r78_c231 bl[231] br[231] wl[78] vdd gnd cell_6t
Xbit_r79_c231 bl[231] br[231] wl[79] vdd gnd cell_6t
Xbit_r80_c231 bl[231] br[231] wl[80] vdd gnd cell_6t
Xbit_r81_c231 bl[231] br[231] wl[81] vdd gnd cell_6t
Xbit_r82_c231 bl[231] br[231] wl[82] vdd gnd cell_6t
Xbit_r83_c231 bl[231] br[231] wl[83] vdd gnd cell_6t
Xbit_r84_c231 bl[231] br[231] wl[84] vdd gnd cell_6t
Xbit_r85_c231 bl[231] br[231] wl[85] vdd gnd cell_6t
Xbit_r86_c231 bl[231] br[231] wl[86] vdd gnd cell_6t
Xbit_r87_c231 bl[231] br[231] wl[87] vdd gnd cell_6t
Xbit_r88_c231 bl[231] br[231] wl[88] vdd gnd cell_6t
Xbit_r89_c231 bl[231] br[231] wl[89] vdd gnd cell_6t
Xbit_r90_c231 bl[231] br[231] wl[90] vdd gnd cell_6t
Xbit_r91_c231 bl[231] br[231] wl[91] vdd gnd cell_6t
Xbit_r92_c231 bl[231] br[231] wl[92] vdd gnd cell_6t
Xbit_r93_c231 bl[231] br[231] wl[93] vdd gnd cell_6t
Xbit_r94_c231 bl[231] br[231] wl[94] vdd gnd cell_6t
Xbit_r95_c231 bl[231] br[231] wl[95] vdd gnd cell_6t
Xbit_r96_c231 bl[231] br[231] wl[96] vdd gnd cell_6t
Xbit_r97_c231 bl[231] br[231] wl[97] vdd gnd cell_6t
Xbit_r98_c231 bl[231] br[231] wl[98] vdd gnd cell_6t
Xbit_r99_c231 bl[231] br[231] wl[99] vdd gnd cell_6t
Xbit_r100_c231 bl[231] br[231] wl[100] vdd gnd cell_6t
Xbit_r101_c231 bl[231] br[231] wl[101] vdd gnd cell_6t
Xbit_r102_c231 bl[231] br[231] wl[102] vdd gnd cell_6t
Xbit_r103_c231 bl[231] br[231] wl[103] vdd gnd cell_6t
Xbit_r104_c231 bl[231] br[231] wl[104] vdd gnd cell_6t
Xbit_r105_c231 bl[231] br[231] wl[105] vdd gnd cell_6t
Xbit_r106_c231 bl[231] br[231] wl[106] vdd gnd cell_6t
Xbit_r107_c231 bl[231] br[231] wl[107] vdd gnd cell_6t
Xbit_r108_c231 bl[231] br[231] wl[108] vdd gnd cell_6t
Xbit_r109_c231 bl[231] br[231] wl[109] vdd gnd cell_6t
Xbit_r110_c231 bl[231] br[231] wl[110] vdd gnd cell_6t
Xbit_r111_c231 bl[231] br[231] wl[111] vdd gnd cell_6t
Xbit_r112_c231 bl[231] br[231] wl[112] vdd gnd cell_6t
Xbit_r113_c231 bl[231] br[231] wl[113] vdd gnd cell_6t
Xbit_r114_c231 bl[231] br[231] wl[114] vdd gnd cell_6t
Xbit_r115_c231 bl[231] br[231] wl[115] vdd gnd cell_6t
Xbit_r116_c231 bl[231] br[231] wl[116] vdd gnd cell_6t
Xbit_r117_c231 bl[231] br[231] wl[117] vdd gnd cell_6t
Xbit_r118_c231 bl[231] br[231] wl[118] vdd gnd cell_6t
Xbit_r119_c231 bl[231] br[231] wl[119] vdd gnd cell_6t
Xbit_r120_c231 bl[231] br[231] wl[120] vdd gnd cell_6t
Xbit_r121_c231 bl[231] br[231] wl[121] vdd gnd cell_6t
Xbit_r122_c231 bl[231] br[231] wl[122] vdd gnd cell_6t
Xbit_r123_c231 bl[231] br[231] wl[123] vdd gnd cell_6t
Xbit_r124_c231 bl[231] br[231] wl[124] vdd gnd cell_6t
Xbit_r125_c231 bl[231] br[231] wl[125] vdd gnd cell_6t
Xbit_r126_c231 bl[231] br[231] wl[126] vdd gnd cell_6t
Xbit_r127_c231 bl[231] br[231] wl[127] vdd gnd cell_6t
Xbit_r128_c231 bl[231] br[231] wl[128] vdd gnd cell_6t
Xbit_r129_c231 bl[231] br[231] wl[129] vdd gnd cell_6t
Xbit_r130_c231 bl[231] br[231] wl[130] vdd gnd cell_6t
Xbit_r131_c231 bl[231] br[231] wl[131] vdd gnd cell_6t
Xbit_r132_c231 bl[231] br[231] wl[132] vdd gnd cell_6t
Xbit_r133_c231 bl[231] br[231] wl[133] vdd gnd cell_6t
Xbit_r134_c231 bl[231] br[231] wl[134] vdd gnd cell_6t
Xbit_r135_c231 bl[231] br[231] wl[135] vdd gnd cell_6t
Xbit_r136_c231 bl[231] br[231] wl[136] vdd gnd cell_6t
Xbit_r137_c231 bl[231] br[231] wl[137] vdd gnd cell_6t
Xbit_r138_c231 bl[231] br[231] wl[138] vdd gnd cell_6t
Xbit_r139_c231 bl[231] br[231] wl[139] vdd gnd cell_6t
Xbit_r140_c231 bl[231] br[231] wl[140] vdd gnd cell_6t
Xbit_r141_c231 bl[231] br[231] wl[141] vdd gnd cell_6t
Xbit_r142_c231 bl[231] br[231] wl[142] vdd gnd cell_6t
Xbit_r143_c231 bl[231] br[231] wl[143] vdd gnd cell_6t
Xbit_r144_c231 bl[231] br[231] wl[144] vdd gnd cell_6t
Xbit_r145_c231 bl[231] br[231] wl[145] vdd gnd cell_6t
Xbit_r146_c231 bl[231] br[231] wl[146] vdd gnd cell_6t
Xbit_r147_c231 bl[231] br[231] wl[147] vdd gnd cell_6t
Xbit_r148_c231 bl[231] br[231] wl[148] vdd gnd cell_6t
Xbit_r149_c231 bl[231] br[231] wl[149] vdd gnd cell_6t
Xbit_r150_c231 bl[231] br[231] wl[150] vdd gnd cell_6t
Xbit_r151_c231 bl[231] br[231] wl[151] vdd gnd cell_6t
Xbit_r152_c231 bl[231] br[231] wl[152] vdd gnd cell_6t
Xbit_r153_c231 bl[231] br[231] wl[153] vdd gnd cell_6t
Xbit_r154_c231 bl[231] br[231] wl[154] vdd gnd cell_6t
Xbit_r155_c231 bl[231] br[231] wl[155] vdd gnd cell_6t
Xbit_r156_c231 bl[231] br[231] wl[156] vdd gnd cell_6t
Xbit_r157_c231 bl[231] br[231] wl[157] vdd gnd cell_6t
Xbit_r158_c231 bl[231] br[231] wl[158] vdd gnd cell_6t
Xbit_r159_c231 bl[231] br[231] wl[159] vdd gnd cell_6t
Xbit_r160_c231 bl[231] br[231] wl[160] vdd gnd cell_6t
Xbit_r161_c231 bl[231] br[231] wl[161] vdd gnd cell_6t
Xbit_r162_c231 bl[231] br[231] wl[162] vdd gnd cell_6t
Xbit_r163_c231 bl[231] br[231] wl[163] vdd gnd cell_6t
Xbit_r164_c231 bl[231] br[231] wl[164] vdd gnd cell_6t
Xbit_r165_c231 bl[231] br[231] wl[165] vdd gnd cell_6t
Xbit_r166_c231 bl[231] br[231] wl[166] vdd gnd cell_6t
Xbit_r167_c231 bl[231] br[231] wl[167] vdd gnd cell_6t
Xbit_r168_c231 bl[231] br[231] wl[168] vdd gnd cell_6t
Xbit_r169_c231 bl[231] br[231] wl[169] vdd gnd cell_6t
Xbit_r170_c231 bl[231] br[231] wl[170] vdd gnd cell_6t
Xbit_r171_c231 bl[231] br[231] wl[171] vdd gnd cell_6t
Xbit_r172_c231 bl[231] br[231] wl[172] vdd gnd cell_6t
Xbit_r173_c231 bl[231] br[231] wl[173] vdd gnd cell_6t
Xbit_r174_c231 bl[231] br[231] wl[174] vdd gnd cell_6t
Xbit_r175_c231 bl[231] br[231] wl[175] vdd gnd cell_6t
Xbit_r176_c231 bl[231] br[231] wl[176] vdd gnd cell_6t
Xbit_r177_c231 bl[231] br[231] wl[177] vdd gnd cell_6t
Xbit_r178_c231 bl[231] br[231] wl[178] vdd gnd cell_6t
Xbit_r179_c231 bl[231] br[231] wl[179] vdd gnd cell_6t
Xbit_r180_c231 bl[231] br[231] wl[180] vdd gnd cell_6t
Xbit_r181_c231 bl[231] br[231] wl[181] vdd gnd cell_6t
Xbit_r182_c231 bl[231] br[231] wl[182] vdd gnd cell_6t
Xbit_r183_c231 bl[231] br[231] wl[183] vdd gnd cell_6t
Xbit_r184_c231 bl[231] br[231] wl[184] vdd gnd cell_6t
Xbit_r185_c231 bl[231] br[231] wl[185] vdd gnd cell_6t
Xbit_r186_c231 bl[231] br[231] wl[186] vdd gnd cell_6t
Xbit_r187_c231 bl[231] br[231] wl[187] vdd gnd cell_6t
Xbit_r188_c231 bl[231] br[231] wl[188] vdd gnd cell_6t
Xbit_r189_c231 bl[231] br[231] wl[189] vdd gnd cell_6t
Xbit_r190_c231 bl[231] br[231] wl[190] vdd gnd cell_6t
Xbit_r191_c231 bl[231] br[231] wl[191] vdd gnd cell_6t
Xbit_r192_c231 bl[231] br[231] wl[192] vdd gnd cell_6t
Xbit_r193_c231 bl[231] br[231] wl[193] vdd gnd cell_6t
Xbit_r194_c231 bl[231] br[231] wl[194] vdd gnd cell_6t
Xbit_r195_c231 bl[231] br[231] wl[195] vdd gnd cell_6t
Xbit_r196_c231 bl[231] br[231] wl[196] vdd gnd cell_6t
Xbit_r197_c231 bl[231] br[231] wl[197] vdd gnd cell_6t
Xbit_r198_c231 bl[231] br[231] wl[198] vdd gnd cell_6t
Xbit_r199_c231 bl[231] br[231] wl[199] vdd gnd cell_6t
Xbit_r200_c231 bl[231] br[231] wl[200] vdd gnd cell_6t
Xbit_r201_c231 bl[231] br[231] wl[201] vdd gnd cell_6t
Xbit_r202_c231 bl[231] br[231] wl[202] vdd gnd cell_6t
Xbit_r203_c231 bl[231] br[231] wl[203] vdd gnd cell_6t
Xbit_r204_c231 bl[231] br[231] wl[204] vdd gnd cell_6t
Xbit_r205_c231 bl[231] br[231] wl[205] vdd gnd cell_6t
Xbit_r206_c231 bl[231] br[231] wl[206] vdd gnd cell_6t
Xbit_r207_c231 bl[231] br[231] wl[207] vdd gnd cell_6t
Xbit_r208_c231 bl[231] br[231] wl[208] vdd gnd cell_6t
Xbit_r209_c231 bl[231] br[231] wl[209] vdd gnd cell_6t
Xbit_r210_c231 bl[231] br[231] wl[210] vdd gnd cell_6t
Xbit_r211_c231 bl[231] br[231] wl[211] vdd gnd cell_6t
Xbit_r212_c231 bl[231] br[231] wl[212] vdd gnd cell_6t
Xbit_r213_c231 bl[231] br[231] wl[213] vdd gnd cell_6t
Xbit_r214_c231 bl[231] br[231] wl[214] vdd gnd cell_6t
Xbit_r215_c231 bl[231] br[231] wl[215] vdd gnd cell_6t
Xbit_r216_c231 bl[231] br[231] wl[216] vdd gnd cell_6t
Xbit_r217_c231 bl[231] br[231] wl[217] vdd gnd cell_6t
Xbit_r218_c231 bl[231] br[231] wl[218] vdd gnd cell_6t
Xbit_r219_c231 bl[231] br[231] wl[219] vdd gnd cell_6t
Xbit_r220_c231 bl[231] br[231] wl[220] vdd gnd cell_6t
Xbit_r221_c231 bl[231] br[231] wl[221] vdd gnd cell_6t
Xbit_r222_c231 bl[231] br[231] wl[222] vdd gnd cell_6t
Xbit_r223_c231 bl[231] br[231] wl[223] vdd gnd cell_6t
Xbit_r224_c231 bl[231] br[231] wl[224] vdd gnd cell_6t
Xbit_r225_c231 bl[231] br[231] wl[225] vdd gnd cell_6t
Xbit_r226_c231 bl[231] br[231] wl[226] vdd gnd cell_6t
Xbit_r227_c231 bl[231] br[231] wl[227] vdd gnd cell_6t
Xbit_r228_c231 bl[231] br[231] wl[228] vdd gnd cell_6t
Xbit_r229_c231 bl[231] br[231] wl[229] vdd gnd cell_6t
Xbit_r230_c231 bl[231] br[231] wl[230] vdd gnd cell_6t
Xbit_r231_c231 bl[231] br[231] wl[231] vdd gnd cell_6t
Xbit_r232_c231 bl[231] br[231] wl[232] vdd gnd cell_6t
Xbit_r233_c231 bl[231] br[231] wl[233] vdd gnd cell_6t
Xbit_r234_c231 bl[231] br[231] wl[234] vdd gnd cell_6t
Xbit_r235_c231 bl[231] br[231] wl[235] vdd gnd cell_6t
Xbit_r236_c231 bl[231] br[231] wl[236] vdd gnd cell_6t
Xbit_r237_c231 bl[231] br[231] wl[237] vdd gnd cell_6t
Xbit_r238_c231 bl[231] br[231] wl[238] vdd gnd cell_6t
Xbit_r239_c231 bl[231] br[231] wl[239] vdd gnd cell_6t
Xbit_r240_c231 bl[231] br[231] wl[240] vdd gnd cell_6t
Xbit_r241_c231 bl[231] br[231] wl[241] vdd gnd cell_6t
Xbit_r242_c231 bl[231] br[231] wl[242] vdd gnd cell_6t
Xbit_r243_c231 bl[231] br[231] wl[243] vdd gnd cell_6t
Xbit_r244_c231 bl[231] br[231] wl[244] vdd gnd cell_6t
Xbit_r245_c231 bl[231] br[231] wl[245] vdd gnd cell_6t
Xbit_r246_c231 bl[231] br[231] wl[246] vdd gnd cell_6t
Xbit_r247_c231 bl[231] br[231] wl[247] vdd gnd cell_6t
Xbit_r248_c231 bl[231] br[231] wl[248] vdd gnd cell_6t
Xbit_r249_c231 bl[231] br[231] wl[249] vdd gnd cell_6t
Xbit_r250_c231 bl[231] br[231] wl[250] vdd gnd cell_6t
Xbit_r251_c231 bl[231] br[231] wl[251] vdd gnd cell_6t
Xbit_r252_c231 bl[231] br[231] wl[252] vdd gnd cell_6t
Xbit_r253_c231 bl[231] br[231] wl[253] vdd gnd cell_6t
Xbit_r254_c231 bl[231] br[231] wl[254] vdd gnd cell_6t
Xbit_r255_c231 bl[231] br[231] wl[255] vdd gnd cell_6t
Xbit_r0_c232 bl[232] br[232] wl[0] vdd gnd cell_6t
Xbit_r1_c232 bl[232] br[232] wl[1] vdd gnd cell_6t
Xbit_r2_c232 bl[232] br[232] wl[2] vdd gnd cell_6t
Xbit_r3_c232 bl[232] br[232] wl[3] vdd gnd cell_6t
Xbit_r4_c232 bl[232] br[232] wl[4] vdd gnd cell_6t
Xbit_r5_c232 bl[232] br[232] wl[5] vdd gnd cell_6t
Xbit_r6_c232 bl[232] br[232] wl[6] vdd gnd cell_6t
Xbit_r7_c232 bl[232] br[232] wl[7] vdd gnd cell_6t
Xbit_r8_c232 bl[232] br[232] wl[8] vdd gnd cell_6t
Xbit_r9_c232 bl[232] br[232] wl[9] vdd gnd cell_6t
Xbit_r10_c232 bl[232] br[232] wl[10] vdd gnd cell_6t
Xbit_r11_c232 bl[232] br[232] wl[11] vdd gnd cell_6t
Xbit_r12_c232 bl[232] br[232] wl[12] vdd gnd cell_6t
Xbit_r13_c232 bl[232] br[232] wl[13] vdd gnd cell_6t
Xbit_r14_c232 bl[232] br[232] wl[14] vdd gnd cell_6t
Xbit_r15_c232 bl[232] br[232] wl[15] vdd gnd cell_6t
Xbit_r16_c232 bl[232] br[232] wl[16] vdd gnd cell_6t
Xbit_r17_c232 bl[232] br[232] wl[17] vdd gnd cell_6t
Xbit_r18_c232 bl[232] br[232] wl[18] vdd gnd cell_6t
Xbit_r19_c232 bl[232] br[232] wl[19] vdd gnd cell_6t
Xbit_r20_c232 bl[232] br[232] wl[20] vdd gnd cell_6t
Xbit_r21_c232 bl[232] br[232] wl[21] vdd gnd cell_6t
Xbit_r22_c232 bl[232] br[232] wl[22] vdd gnd cell_6t
Xbit_r23_c232 bl[232] br[232] wl[23] vdd gnd cell_6t
Xbit_r24_c232 bl[232] br[232] wl[24] vdd gnd cell_6t
Xbit_r25_c232 bl[232] br[232] wl[25] vdd gnd cell_6t
Xbit_r26_c232 bl[232] br[232] wl[26] vdd gnd cell_6t
Xbit_r27_c232 bl[232] br[232] wl[27] vdd gnd cell_6t
Xbit_r28_c232 bl[232] br[232] wl[28] vdd gnd cell_6t
Xbit_r29_c232 bl[232] br[232] wl[29] vdd gnd cell_6t
Xbit_r30_c232 bl[232] br[232] wl[30] vdd gnd cell_6t
Xbit_r31_c232 bl[232] br[232] wl[31] vdd gnd cell_6t
Xbit_r32_c232 bl[232] br[232] wl[32] vdd gnd cell_6t
Xbit_r33_c232 bl[232] br[232] wl[33] vdd gnd cell_6t
Xbit_r34_c232 bl[232] br[232] wl[34] vdd gnd cell_6t
Xbit_r35_c232 bl[232] br[232] wl[35] vdd gnd cell_6t
Xbit_r36_c232 bl[232] br[232] wl[36] vdd gnd cell_6t
Xbit_r37_c232 bl[232] br[232] wl[37] vdd gnd cell_6t
Xbit_r38_c232 bl[232] br[232] wl[38] vdd gnd cell_6t
Xbit_r39_c232 bl[232] br[232] wl[39] vdd gnd cell_6t
Xbit_r40_c232 bl[232] br[232] wl[40] vdd gnd cell_6t
Xbit_r41_c232 bl[232] br[232] wl[41] vdd gnd cell_6t
Xbit_r42_c232 bl[232] br[232] wl[42] vdd gnd cell_6t
Xbit_r43_c232 bl[232] br[232] wl[43] vdd gnd cell_6t
Xbit_r44_c232 bl[232] br[232] wl[44] vdd gnd cell_6t
Xbit_r45_c232 bl[232] br[232] wl[45] vdd gnd cell_6t
Xbit_r46_c232 bl[232] br[232] wl[46] vdd gnd cell_6t
Xbit_r47_c232 bl[232] br[232] wl[47] vdd gnd cell_6t
Xbit_r48_c232 bl[232] br[232] wl[48] vdd gnd cell_6t
Xbit_r49_c232 bl[232] br[232] wl[49] vdd gnd cell_6t
Xbit_r50_c232 bl[232] br[232] wl[50] vdd gnd cell_6t
Xbit_r51_c232 bl[232] br[232] wl[51] vdd gnd cell_6t
Xbit_r52_c232 bl[232] br[232] wl[52] vdd gnd cell_6t
Xbit_r53_c232 bl[232] br[232] wl[53] vdd gnd cell_6t
Xbit_r54_c232 bl[232] br[232] wl[54] vdd gnd cell_6t
Xbit_r55_c232 bl[232] br[232] wl[55] vdd gnd cell_6t
Xbit_r56_c232 bl[232] br[232] wl[56] vdd gnd cell_6t
Xbit_r57_c232 bl[232] br[232] wl[57] vdd gnd cell_6t
Xbit_r58_c232 bl[232] br[232] wl[58] vdd gnd cell_6t
Xbit_r59_c232 bl[232] br[232] wl[59] vdd gnd cell_6t
Xbit_r60_c232 bl[232] br[232] wl[60] vdd gnd cell_6t
Xbit_r61_c232 bl[232] br[232] wl[61] vdd gnd cell_6t
Xbit_r62_c232 bl[232] br[232] wl[62] vdd gnd cell_6t
Xbit_r63_c232 bl[232] br[232] wl[63] vdd gnd cell_6t
Xbit_r64_c232 bl[232] br[232] wl[64] vdd gnd cell_6t
Xbit_r65_c232 bl[232] br[232] wl[65] vdd gnd cell_6t
Xbit_r66_c232 bl[232] br[232] wl[66] vdd gnd cell_6t
Xbit_r67_c232 bl[232] br[232] wl[67] vdd gnd cell_6t
Xbit_r68_c232 bl[232] br[232] wl[68] vdd gnd cell_6t
Xbit_r69_c232 bl[232] br[232] wl[69] vdd gnd cell_6t
Xbit_r70_c232 bl[232] br[232] wl[70] vdd gnd cell_6t
Xbit_r71_c232 bl[232] br[232] wl[71] vdd gnd cell_6t
Xbit_r72_c232 bl[232] br[232] wl[72] vdd gnd cell_6t
Xbit_r73_c232 bl[232] br[232] wl[73] vdd gnd cell_6t
Xbit_r74_c232 bl[232] br[232] wl[74] vdd gnd cell_6t
Xbit_r75_c232 bl[232] br[232] wl[75] vdd gnd cell_6t
Xbit_r76_c232 bl[232] br[232] wl[76] vdd gnd cell_6t
Xbit_r77_c232 bl[232] br[232] wl[77] vdd gnd cell_6t
Xbit_r78_c232 bl[232] br[232] wl[78] vdd gnd cell_6t
Xbit_r79_c232 bl[232] br[232] wl[79] vdd gnd cell_6t
Xbit_r80_c232 bl[232] br[232] wl[80] vdd gnd cell_6t
Xbit_r81_c232 bl[232] br[232] wl[81] vdd gnd cell_6t
Xbit_r82_c232 bl[232] br[232] wl[82] vdd gnd cell_6t
Xbit_r83_c232 bl[232] br[232] wl[83] vdd gnd cell_6t
Xbit_r84_c232 bl[232] br[232] wl[84] vdd gnd cell_6t
Xbit_r85_c232 bl[232] br[232] wl[85] vdd gnd cell_6t
Xbit_r86_c232 bl[232] br[232] wl[86] vdd gnd cell_6t
Xbit_r87_c232 bl[232] br[232] wl[87] vdd gnd cell_6t
Xbit_r88_c232 bl[232] br[232] wl[88] vdd gnd cell_6t
Xbit_r89_c232 bl[232] br[232] wl[89] vdd gnd cell_6t
Xbit_r90_c232 bl[232] br[232] wl[90] vdd gnd cell_6t
Xbit_r91_c232 bl[232] br[232] wl[91] vdd gnd cell_6t
Xbit_r92_c232 bl[232] br[232] wl[92] vdd gnd cell_6t
Xbit_r93_c232 bl[232] br[232] wl[93] vdd gnd cell_6t
Xbit_r94_c232 bl[232] br[232] wl[94] vdd gnd cell_6t
Xbit_r95_c232 bl[232] br[232] wl[95] vdd gnd cell_6t
Xbit_r96_c232 bl[232] br[232] wl[96] vdd gnd cell_6t
Xbit_r97_c232 bl[232] br[232] wl[97] vdd gnd cell_6t
Xbit_r98_c232 bl[232] br[232] wl[98] vdd gnd cell_6t
Xbit_r99_c232 bl[232] br[232] wl[99] vdd gnd cell_6t
Xbit_r100_c232 bl[232] br[232] wl[100] vdd gnd cell_6t
Xbit_r101_c232 bl[232] br[232] wl[101] vdd gnd cell_6t
Xbit_r102_c232 bl[232] br[232] wl[102] vdd gnd cell_6t
Xbit_r103_c232 bl[232] br[232] wl[103] vdd gnd cell_6t
Xbit_r104_c232 bl[232] br[232] wl[104] vdd gnd cell_6t
Xbit_r105_c232 bl[232] br[232] wl[105] vdd gnd cell_6t
Xbit_r106_c232 bl[232] br[232] wl[106] vdd gnd cell_6t
Xbit_r107_c232 bl[232] br[232] wl[107] vdd gnd cell_6t
Xbit_r108_c232 bl[232] br[232] wl[108] vdd gnd cell_6t
Xbit_r109_c232 bl[232] br[232] wl[109] vdd gnd cell_6t
Xbit_r110_c232 bl[232] br[232] wl[110] vdd gnd cell_6t
Xbit_r111_c232 bl[232] br[232] wl[111] vdd gnd cell_6t
Xbit_r112_c232 bl[232] br[232] wl[112] vdd gnd cell_6t
Xbit_r113_c232 bl[232] br[232] wl[113] vdd gnd cell_6t
Xbit_r114_c232 bl[232] br[232] wl[114] vdd gnd cell_6t
Xbit_r115_c232 bl[232] br[232] wl[115] vdd gnd cell_6t
Xbit_r116_c232 bl[232] br[232] wl[116] vdd gnd cell_6t
Xbit_r117_c232 bl[232] br[232] wl[117] vdd gnd cell_6t
Xbit_r118_c232 bl[232] br[232] wl[118] vdd gnd cell_6t
Xbit_r119_c232 bl[232] br[232] wl[119] vdd gnd cell_6t
Xbit_r120_c232 bl[232] br[232] wl[120] vdd gnd cell_6t
Xbit_r121_c232 bl[232] br[232] wl[121] vdd gnd cell_6t
Xbit_r122_c232 bl[232] br[232] wl[122] vdd gnd cell_6t
Xbit_r123_c232 bl[232] br[232] wl[123] vdd gnd cell_6t
Xbit_r124_c232 bl[232] br[232] wl[124] vdd gnd cell_6t
Xbit_r125_c232 bl[232] br[232] wl[125] vdd gnd cell_6t
Xbit_r126_c232 bl[232] br[232] wl[126] vdd gnd cell_6t
Xbit_r127_c232 bl[232] br[232] wl[127] vdd gnd cell_6t
Xbit_r128_c232 bl[232] br[232] wl[128] vdd gnd cell_6t
Xbit_r129_c232 bl[232] br[232] wl[129] vdd gnd cell_6t
Xbit_r130_c232 bl[232] br[232] wl[130] vdd gnd cell_6t
Xbit_r131_c232 bl[232] br[232] wl[131] vdd gnd cell_6t
Xbit_r132_c232 bl[232] br[232] wl[132] vdd gnd cell_6t
Xbit_r133_c232 bl[232] br[232] wl[133] vdd gnd cell_6t
Xbit_r134_c232 bl[232] br[232] wl[134] vdd gnd cell_6t
Xbit_r135_c232 bl[232] br[232] wl[135] vdd gnd cell_6t
Xbit_r136_c232 bl[232] br[232] wl[136] vdd gnd cell_6t
Xbit_r137_c232 bl[232] br[232] wl[137] vdd gnd cell_6t
Xbit_r138_c232 bl[232] br[232] wl[138] vdd gnd cell_6t
Xbit_r139_c232 bl[232] br[232] wl[139] vdd gnd cell_6t
Xbit_r140_c232 bl[232] br[232] wl[140] vdd gnd cell_6t
Xbit_r141_c232 bl[232] br[232] wl[141] vdd gnd cell_6t
Xbit_r142_c232 bl[232] br[232] wl[142] vdd gnd cell_6t
Xbit_r143_c232 bl[232] br[232] wl[143] vdd gnd cell_6t
Xbit_r144_c232 bl[232] br[232] wl[144] vdd gnd cell_6t
Xbit_r145_c232 bl[232] br[232] wl[145] vdd gnd cell_6t
Xbit_r146_c232 bl[232] br[232] wl[146] vdd gnd cell_6t
Xbit_r147_c232 bl[232] br[232] wl[147] vdd gnd cell_6t
Xbit_r148_c232 bl[232] br[232] wl[148] vdd gnd cell_6t
Xbit_r149_c232 bl[232] br[232] wl[149] vdd gnd cell_6t
Xbit_r150_c232 bl[232] br[232] wl[150] vdd gnd cell_6t
Xbit_r151_c232 bl[232] br[232] wl[151] vdd gnd cell_6t
Xbit_r152_c232 bl[232] br[232] wl[152] vdd gnd cell_6t
Xbit_r153_c232 bl[232] br[232] wl[153] vdd gnd cell_6t
Xbit_r154_c232 bl[232] br[232] wl[154] vdd gnd cell_6t
Xbit_r155_c232 bl[232] br[232] wl[155] vdd gnd cell_6t
Xbit_r156_c232 bl[232] br[232] wl[156] vdd gnd cell_6t
Xbit_r157_c232 bl[232] br[232] wl[157] vdd gnd cell_6t
Xbit_r158_c232 bl[232] br[232] wl[158] vdd gnd cell_6t
Xbit_r159_c232 bl[232] br[232] wl[159] vdd gnd cell_6t
Xbit_r160_c232 bl[232] br[232] wl[160] vdd gnd cell_6t
Xbit_r161_c232 bl[232] br[232] wl[161] vdd gnd cell_6t
Xbit_r162_c232 bl[232] br[232] wl[162] vdd gnd cell_6t
Xbit_r163_c232 bl[232] br[232] wl[163] vdd gnd cell_6t
Xbit_r164_c232 bl[232] br[232] wl[164] vdd gnd cell_6t
Xbit_r165_c232 bl[232] br[232] wl[165] vdd gnd cell_6t
Xbit_r166_c232 bl[232] br[232] wl[166] vdd gnd cell_6t
Xbit_r167_c232 bl[232] br[232] wl[167] vdd gnd cell_6t
Xbit_r168_c232 bl[232] br[232] wl[168] vdd gnd cell_6t
Xbit_r169_c232 bl[232] br[232] wl[169] vdd gnd cell_6t
Xbit_r170_c232 bl[232] br[232] wl[170] vdd gnd cell_6t
Xbit_r171_c232 bl[232] br[232] wl[171] vdd gnd cell_6t
Xbit_r172_c232 bl[232] br[232] wl[172] vdd gnd cell_6t
Xbit_r173_c232 bl[232] br[232] wl[173] vdd gnd cell_6t
Xbit_r174_c232 bl[232] br[232] wl[174] vdd gnd cell_6t
Xbit_r175_c232 bl[232] br[232] wl[175] vdd gnd cell_6t
Xbit_r176_c232 bl[232] br[232] wl[176] vdd gnd cell_6t
Xbit_r177_c232 bl[232] br[232] wl[177] vdd gnd cell_6t
Xbit_r178_c232 bl[232] br[232] wl[178] vdd gnd cell_6t
Xbit_r179_c232 bl[232] br[232] wl[179] vdd gnd cell_6t
Xbit_r180_c232 bl[232] br[232] wl[180] vdd gnd cell_6t
Xbit_r181_c232 bl[232] br[232] wl[181] vdd gnd cell_6t
Xbit_r182_c232 bl[232] br[232] wl[182] vdd gnd cell_6t
Xbit_r183_c232 bl[232] br[232] wl[183] vdd gnd cell_6t
Xbit_r184_c232 bl[232] br[232] wl[184] vdd gnd cell_6t
Xbit_r185_c232 bl[232] br[232] wl[185] vdd gnd cell_6t
Xbit_r186_c232 bl[232] br[232] wl[186] vdd gnd cell_6t
Xbit_r187_c232 bl[232] br[232] wl[187] vdd gnd cell_6t
Xbit_r188_c232 bl[232] br[232] wl[188] vdd gnd cell_6t
Xbit_r189_c232 bl[232] br[232] wl[189] vdd gnd cell_6t
Xbit_r190_c232 bl[232] br[232] wl[190] vdd gnd cell_6t
Xbit_r191_c232 bl[232] br[232] wl[191] vdd gnd cell_6t
Xbit_r192_c232 bl[232] br[232] wl[192] vdd gnd cell_6t
Xbit_r193_c232 bl[232] br[232] wl[193] vdd gnd cell_6t
Xbit_r194_c232 bl[232] br[232] wl[194] vdd gnd cell_6t
Xbit_r195_c232 bl[232] br[232] wl[195] vdd gnd cell_6t
Xbit_r196_c232 bl[232] br[232] wl[196] vdd gnd cell_6t
Xbit_r197_c232 bl[232] br[232] wl[197] vdd gnd cell_6t
Xbit_r198_c232 bl[232] br[232] wl[198] vdd gnd cell_6t
Xbit_r199_c232 bl[232] br[232] wl[199] vdd gnd cell_6t
Xbit_r200_c232 bl[232] br[232] wl[200] vdd gnd cell_6t
Xbit_r201_c232 bl[232] br[232] wl[201] vdd gnd cell_6t
Xbit_r202_c232 bl[232] br[232] wl[202] vdd gnd cell_6t
Xbit_r203_c232 bl[232] br[232] wl[203] vdd gnd cell_6t
Xbit_r204_c232 bl[232] br[232] wl[204] vdd gnd cell_6t
Xbit_r205_c232 bl[232] br[232] wl[205] vdd gnd cell_6t
Xbit_r206_c232 bl[232] br[232] wl[206] vdd gnd cell_6t
Xbit_r207_c232 bl[232] br[232] wl[207] vdd gnd cell_6t
Xbit_r208_c232 bl[232] br[232] wl[208] vdd gnd cell_6t
Xbit_r209_c232 bl[232] br[232] wl[209] vdd gnd cell_6t
Xbit_r210_c232 bl[232] br[232] wl[210] vdd gnd cell_6t
Xbit_r211_c232 bl[232] br[232] wl[211] vdd gnd cell_6t
Xbit_r212_c232 bl[232] br[232] wl[212] vdd gnd cell_6t
Xbit_r213_c232 bl[232] br[232] wl[213] vdd gnd cell_6t
Xbit_r214_c232 bl[232] br[232] wl[214] vdd gnd cell_6t
Xbit_r215_c232 bl[232] br[232] wl[215] vdd gnd cell_6t
Xbit_r216_c232 bl[232] br[232] wl[216] vdd gnd cell_6t
Xbit_r217_c232 bl[232] br[232] wl[217] vdd gnd cell_6t
Xbit_r218_c232 bl[232] br[232] wl[218] vdd gnd cell_6t
Xbit_r219_c232 bl[232] br[232] wl[219] vdd gnd cell_6t
Xbit_r220_c232 bl[232] br[232] wl[220] vdd gnd cell_6t
Xbit_r221_c232 bl[232] br[232] wl[221] vdd gnd cell_6t
Xbit_r222_c232 bl[232] br[232] wl[222] vdd gnd cell_6t
Xbit_r223_c232 bl[232] br[232] wl[223] vdd gnd cell_6t
Xbit_r224_c232 bl[232] br[232] wl[224] vdd gnd cell_6t
Xbit_r225_c232 bl[232] br[232] wl[225] vdd gnd cell_6t
Xbit_r226_c232 bl[232] br[232] wl[226] vdd gnd cell_6t
Xbit_r227_c232 bl[232] br[232] wl[227] vdd gnd cell_6t
Xbit_r228_c232 bl[232] br[232] wl[228] vdd gnd cell_6t
Xbit_r229_c232 bl[232] br[232] wl[229] vdd gnd cell_6t
Xbit_r230_c232 bl[232] br[232] wl[230] vdd gnd cell_6t
Xbit_r231_c232 bl[232] br[232] wl[231] vdd gnd cell_6t
Xbit_r232_c232 bl[232] br[232] wl[232] vdd gnd cell_6t
Xbit_r233_c232 bl[232] br[232] wl[233] vdd gnd cell_6t
Xbit_r234_c232 bl[232] br[232] wl[234] vdd gnd cell_6t
Xbit_r235_c232 bl[232] br[232] wl[235] vdd gnd cell_6t
Xbit_r236_c232 bl[232] br[232] wl[236] vdd gnd cell_6t
Xbit_r237_c232 bl[232] br[232] wl[237] vdd gnd cell_6t
Xbit_r238_c232 bl[232] br[232] wl[238] vdd gnd cell_6t
Xbit_r239_c232 bl[232] br[232] wl[239] vdd gnd cell_6t
Xbit_r240_c232 bl[232] br[232] wl[240] vdd gnd cell_6t
Xbit_r241_c232 bl[232] br[232] wl[241] vdd gnd cell_6t
Xbit_r242_c232 bl[232] br[232] wl[242] vdd gnd cell_6t
Xbit_r243_c232 bl[232] br[232] wl[243] vdd gnd cell_6t
Xbit_r244_c232 bl[232] br[232] wl[244] vdd gnd cell_6t
Xbit_r245_c232 bl[232] br[232] wl[245] vdd gnd cell_6t
Xbit_r246_c232 bl[232] br[232] wl[246] vdd gnd cell_6t
Xbit_r247_c232 bl[232] br[232] wl[247] vdd gnd cell_6t
Xbit_r248_c232 bl[232] br[232] wl[248] vdd gnd cell_6t
Xbit_r249_c232 bl[232] br[232] wl[249] vdd gnd cell_6t
Xbit_r250_c232 bl[232] br[232] wl[250] vdd gnd cell_6t
Xbit_r251_c232 bl[232] br[232] wl[251] vdd gnd cell_6t
Xbit_r252_c232 bl[232] br[232] wl[252] vdd gnd cell_6t
Xbit_r253_c232 bl[232] br[232] wl[253] vdd gnd cell_6t
Xbit_r254_c232 bl[232] br[232] wl[254] vdd gnd cell_6t
Xbit_r255_c232 bl[232] br[232] wl[255] vdd gnd cell_6t
Xbit_r0_c233 bl[233] br[233] wl[0] vdd gnd cell_6t
Xbit_r1_c233 bl[233] br[233] wl[1] vdd gnd cell_6t
Xbit_r2_c233 bl[233] br[233] wl[2] vdd gnd cell_6t
Xbit_r3_c233 bl[233] br[233] wl[3] vdd gnd cell_6t
Xbit_r4_c233 bl[233] br[233] wl[4] vdd gnd cell_6t
Xbit_r5_c233 bl[233] br[233] wl[5] vdd gnd cell_6t
Xbit_r6_c233 bl[233] br[233] wl[6] vdd gnd cell_6t
Xbit_r7_c233 bl[233] br[233] wl[7] vdd gnd cell_6t
Xbit_r8_c233 bl[233] br[233] wl[8] vdd gnd cell_6t
Xbit_r9_c233 bl[233] br[233] wl[9] vdd gnd cell_6t
Xbit_r10_c233 bl[233] br[233] wl[10] vdd gnd cell_6t
Xbit_r11_c233 bl[233] br[233] wl[11] vdd gnd cell_6t
Xbit_r12_c233 bl[233] br[233] wl[12] vdd gnd cell_6t
Xbit_r13_c233 bl[233] br[233] wl[13] vdd gnd cell_6t
Xbit_r14_c233 bl[233] br[233] wl[14] vdd gnd cell_6t
Xbit_r15_c233 bl[233] br[233] wl[15] vdd gnd cell_6t
Xbit_r16_c233 bl[233] br[233] wl[16] vdd gnd cell_6t
Xbit_r17_c233 bl[233] br[233] wl[17] vdd gnd cell_6t
Xbit_r18_c233 bl[233] br[233] wl[18] vdd gnd cell_6t
Xbit_r19_c233 bl[233] br[233] wl[19] vdd gnd cell_6t
Xbit_r20_c233 bl[233] br[233] wl[20] vdd gnd cell_6t
Xbit_r21_c233 bl[233] br[233] wl[21] vdd gnd cell_6t
Xbit_r22_c233 bl[233] br[233] wl[22] vdd gnd cell_6t
Xbit_r23_c233 bl[233] br[233] wl[23] vdd gnd cell_6t
Xbit_r24_c233 bl[233] br[233] wl[24] vdd gnd cell_6t
Xbit_r25_c233 bl[233] br[233] wl[25] vdd gnd cell_6t
Xbit_r26_c233 bl[233] br[233] wl[26] vdd gnd cell_6t
Xbit_r27_c233 bl[233] br[233] wl[27] vdd gnd cell_6t
Xbit_r28_c233 bl[233] br[233] wl[28] vdd gnd cell_6t
Xbit_r29_c233 bl[233] br[233] wl[29] vdd gnd cell_6t
Xbit_r30_c233 bl[233] br[233] wl[30] vdd gnd cell_6t
Xbit_r31_c233 bl[233] br[233] wl[31] vdd gnd cell_6t
Xbit_r32_c233 bl[233] br[233] wl[32] vdd gnd cell_6t
Xbit_r33_c233 bl[233] br[233] wl[33] vdd gnd cell_6t
Xbit_r34_c233 bl[233] br[233] wl[34] vdd gnd cell_6t
Xbit_r35_c233 bl[233] br[233] wl[35] vdd gnd cell_6t
Xbit_r36_c233 bl[233] br[233] wl[36] vdd gnd cell_6t
Xbit_r37_c233 bl[233] br[233] wl[37] vdd gnd cell_6t
Xbit_r38_c233 bl[233] br[233] wl[38] vdd gnd cell_6t
Xbit_r39_c233 bl[233] br[233] wl[39] vdd gnd cell_6t
Xbit_r40_c233 bl[233] br[233] wl[40] vdd gnd cell_6t
Xbit_r41_c233 bl[233] br[233] wl[41] vdd gnd cell_6t
Xbit_r42_c233 bl[233] br[233] wl[42] vdd gnd cell_6t
Xbit_r43_c233 bl[233] br[233] wl[43] vdd gnd cell_6t
Xbit_r44_c233 bl[233] br[233] wl[44] vdd gnd cell_6t
Xbit_r45_c233 bl[233] br[233] wl[45] vdd gnd cell_6t
Xbit_r46_c233 bl[233] br[233] wl[46] vdd gnd cell_6t
Xbit_r47_c233 bl[233] br[233] wl[47] vdd gnd cell_6t
Xbit_r48_c233 bl[233] br[233] wl[48] vdd gnd cell_6t
Xbit_r49_c233 bl[233] br[233] wl[49] vdd gnd cell_6t
Xbit_r50_c233 bl[233] br[233] wl[50] vdd gnd cell_6t
Xbit_r51_c233 bl[233] br[233] wl[51] vdd gnd cell_6t
Xbit_r52_c233 bl[233] br[233] wl[52] vdd gnd cell_6t
Xbit_r53_c233 bl[233] br[233] wl[53] vdd gnd cell_6t
Xbit_r54_c233 bl[233] br[233] wl[54] vdd gnd cell_6t
Xbit_r55_c233 bl[233] br[233] wl[55] vdd gnd cell_6t
Xbit_r56_c233 bl[233] br[233] wl[56] vdd gnd cell_6t
Xbit_r57_c233 bl[233] br[233] wl[57] vdd gnd cell_6t
Xbit_r58_c233 bl[233] br[233] wl[58] vdd gnd cell_6t
Xbit_r59_c233 bl[233] br[233] wl[59] vdd gnd cell_6t
Xbit_r60_c233 bl[233] br[233] wl[60] vdd gnd cell_6t
Xbit_r61_c233 bl[233] br[233] wl[61] vdd gnd cell_6t
Xbit_r62_c233 bl[233] br[233] wl[62] vdd gnd cell_6t
Xbit_r63_c233 bl[233] br[233] wl[63] vdd gnd cell_6t
Xbit_r64_c233 bl[233] br[233] wl[64] vdd gnd cell_6t
Xbit_r65_c233 bl[233] br[233] wl[65] vdd gnd cell_6t
Xbit_r66_c233 bl[233] br[233] wl[66] vdd gnd cell_6t
Xbit_r67_c233 bl[233] br[233] wl[67] vdd gnd cell_6t
Xbit_r68_c233 bl[233] br[233] wl[68] vdd gnd cell_6t
Xbit_r69_c233 bl[233] br[233] wl[69] vdd gnd cell_6t
Xbit_r70_c233 bl[233] br[233] wl[70] vdd gnd cell_6t
Xbit_r71_c233 bl[233] br[233] wl[71] vdd gnd cell_6t
Xbit_r72_c233 bl[233] br[233] wl[72] vdd gnd cell_6t
Xbit_r73_c233 bl[233] br[233] wl[73] vdd gnd cell_6t
Xbit_r74_c233 bl[233] br[233] wl[74] vdd gnd cell_6t
Xbit_r75_c233 bl[233] br[233] wl[75] vdd gnd cell_6t
Xbit_r76_c233 bl[233] br[233] wl[76] vdd gnd cell_6t
Xbit_r77_c233 bl[233] br[233] wl[77] vdd gnd cell_6t
Xbit_r78_c233 bl[233] br[233] wl[78] vdd gnd cell_6t
Xbit_r79_c233 bl[233] br[233] wl[79] vdd gnd cell_6t
Xbit_r80_c233 bl[233] br[233] wl[80] vdd gnd cell_6t
Xbit_r81_c233 bl[233] br[233] wl[81] vdd gnd cell_6t
Xbit_r82_c233 bl[233] br[233] wl[82] vdd gnd cell_6t
Xbit_r83_c233 bl[233] br[233] wl[83] vdd gnd cell_6t
Xbit_r84_c233 bl[233] br[233] wl[84] vdd gnd cell_6t
Xbit_r85_c233 bl[233] br[233] wl[85] vdd gnd cell_6t
Xbit_r86_c233 bl[233] br[233] wl[86] vdd gnd cell_6t
Xbit_r87_c233 bl[233] br[233] wl[87] vdd gnd cell_6t
Xbit_r88_c233 bl[233] br[233] wl[88] vdd gnd cell_6t
Xbit_r89_c233 bl[233] br[233] wl[89] vdd gnd cell_6t
Xbit_r90_c233 bl[233] br[233] wl[90] vdd gnd cell_6t
Xbit_r91_c233 bl[233] br[233] wl[91] vdd gnd cell_6t
Xbit_r92_c233 bl[233] br[233] wl[92] vdd gnd cell_6t
Xbit_r93_c233 bl[233] br[233] wl[93] vdd gnd cell_6t
Xbit_r94_c233 bl[233] br[233] wl[94] vdd gnd cell_6t
Xbit_r95_c233 bl[233] br[233] wl[95] vdd gnd cell_6t
Xbit_r96_c233 bl[233] br[233] wl[96] vdd gnd cell_6t
Xbit_r97_c233 bl[233] br[233] wl[97] vdd gnd cell_6t
Xbit_r98_c233 bl[233] br[233] wl[98] vdd gnd cell_6t
Xbit_r99_c233 bl[233] br[233] wl[99] vdd gnd cell_6t
Xbit_r100_c233 bl[233] br[233] wl[100] vdd gnd cell_6t
Xbit_r101_c233 bl[233] br[233] wl[101] vdd gnd cell_6t
Xbit_r102_c233 bl[233] br[233] wl[102] vdd gnd cell_6t
Xbit_r103_c233 bl[233] br[233] wl[103] vdd gnd cell_6t
Xbit_r104_c233 bl[233] br[233] wl[104] vdd gnd cell_6t
Xbit_r105_c233 bl[233] br[233] wl[105] vdd gnd cell_6t
Xbit_r106_c233 bl[233] br[233] wl[106] vdd gnd cell_6t
Xbit_r107_c233 bl[233] br[233] wl[107] vdd gnd cell_6t
Xbit_r108_c233 bl[233] br[233] wl[108] vdd gnd cell_6t
Xbit_r109_c233 bl[233] br[233] wl[109] vdd gnd cell_6t
Xbit_r110_c233 bl[233] br[233] wl[110] vdd gnd cell_6t
Xbit_r111_c233 bl[233] br[233] wl[111] vdd gnd cell_6t
Xbit_r112_c233 bl[233] br[233] wl[112] vdd gnd cell_6t
Xbit_r113_c233 bl[233] br[233] wl[113] vdd gnd cell_6t
Xbit_r114_c233 bl[233] br[233] wl[114] vdd gnd cell_6t
Xbit_r115_c233 bl[233] br[233] wl[115] vdd gnd cell_6t
Xbit_r116_c233 bl[233] br[233] wl[116] vdd gnd cell_6t
Xbit_r117_c233 bl[233] br[233] wl[117] vdd gnd cell_6t
Xbit_r118_c233 bl[233] br[233] wl[118] vdd gnd cell_6t
Xbit_r119_c233 bl[233] br[233] wl[119] vdd gnd cell_6t
Xbit_r120_c233 bl[233] br[233] wl[120] vdd gnd cell_6t
Xbit_r121_c233 bl[233] br[233] wl[121] vdd gnd cell_6t
Xbit_r122_c233 bl[233] br[233] wl[122] vdd gnd cell_6t
Xbit_r123_c233 bl[233] br[233] wl[123] vdd gnd cell_6t
Xbit_r124_c233 bl[233] br[233] wl[124] vdd gnd cell_6t
Xbit_r125_c233 bl[233] br[233] wl[125] vdd gnd cell_6t
Xbit_r126_c233 bl[233] br[233] wl[126] vdd gnd cell_6t
Xbit_r127_c233 bl[233] br[233] wl[127] vdd gnd cell_6t
Xbit_r128_c233 bl[233] br[233] wl[128] vdd gnd cell_6t
Xbit_r129_c233 bl[233] br[233] wl[129] vdd gnd cell_6t
Xbit_r130_c233 bl[233] br[233] wl[130] vdd gnd cell_6t
Xbit_r131_c233 bl[233] br[233] wl[131] vdd gnd cell_6t
Xbit_r132_c233 bl[233] br[233] wl[132] vdd gnd cell_6t
Xbit_r133_c233 bl[233] br[233] wl[133] vdd gnd cell_6t
Xbit_r134_c233 bl[233] br[233] wl[134] vdd gnd cell_6t
Xbit_r135_c233 bl[233] br[233] wl[135] vdd gnd cell_6t
Xbit_r136_c233 bl[233] br[233] wl[136] vdd gnd cell_6t
Xbit_r137_c233 bl[233] br[233] wl[137] vdd gnd cell_6t
Xbit_r138_c233 bl[233] br[233] wl[138] vdd gnd cell_6t
Xbit_r139_c233 bl[233] br[233] wl[139] vdd gnd cell_6t
Xbit_r140_c233 bl[233] br[233] wl[140] vdd gnd cell_6t
Xbit_r141_c233 bl[233] br[233] wl[141] vdd gnd cell_6t
Xbit_r142_c233 bl[233] br[233] wl[142] vdd gnd cell_6t
Xbit_r143_c233 bl[233] br[233] wl[143] vdd gnd cell_6t
Xbit_r144_c233 bl[233] br[233] wl[144] vdd gnd cell_6t
Xbit_r145_c233 bl[233] br[233] wl[145] vdd gnd cell_6t
Xbit_r146_c233 bl[233] br[233] wl[146] vdd gnd cell_6t
Xbit_r147_c233 bl[233] br[233] wl[147] vdd gnd cell_6t
Xbit_r148_c233 bl[233] br[233] wl[148] vdd gnd cell_6t
Xbit_r149_c233 bl[233] br[233] wl[149] vdd gnd cell_6t
Xbit_r150_c233 bl[233] br[233] wl[150] vdd gnd cell_6t
Xbit_r151_c233 bl[233] br[233] wl[151] vdd gnd cell_6t
Xbit_r152_c233 bl[233] br[233] wl[152] vdd gnd cell_6t
Xbit_r153_c233 bl[233] br[233] wl[153] vdd gnd cell_6t
Xbit_r154_c233 bl[233] br[233] wl[154] vdd gnd cell_6t
Xbit_r155_c233 bl[233] br[233] wl[155] vdd gnd cell_6t
Xbit_r156_c233 bl[233] br[233] wl[156] vdd gnd cell_6t
Xbit_r157_c233 bl[233] br[233] wl[157] vdd gnd cell_6t
Xbit_r158_c233 bl[233] br[233] wl[158] vdd gnd cell_6t
Xbit_r159_c233 bl[233] br[233] wl[159] vdd gnd cell_6t
Xbit_r160_c233 bl[233] br[233] wl[160] vdd gnd cell_6t
Xbit_r161_c233 bl[233] br[233] wl[161] vdd gnd cell_6t
Xbit_r162_c233 bl[233] br[233] wl[162] vdd gnd cell_6t
Xbit_r163_c233 bl[233] br[233] wl[163] vdd gnd cell_6t
Xbit_r164_c233 bl[233] br[233] wl[164] vdd gnd cell_6t
Xbit_r165_c233 bl[233] br[233] wl[165] vdd gnd cell_6t
Xbit_r166_c233 bl[233] br[233] wl[166] vdd gnd cell_6t
Xbit_r167_c233 bl[233] br[233] wl[167] vdd gnd cell_6t
Xbit_r168_c233 bl[233] br[233] wl[168] vdd gnd cell_6t
Xbit_r169_c233 bl[233] br[233] wl[169] vdd gnd cell_6t
Xbit_r170_c233 bl[233] br[233] wl[170] vdd gnd cell_6t
Xbit_r171_c233 bl[233] br[233] wl[171] vdd gnd cell_6t
Xbit_r172_c233 bl[233] br[233] wl[172] vdd gnd cell_6t
Xbit_r173_c233 bl[233] br[233] wl[173] vdd gnd cell_6t
Xbit_r174_c233 bl[233] br[233] wl[174] vdd gnd cell_6t
Xbit_r175_c233 bl[233] br[233] wl[175] vdd gnd cell_6t
Xbit_r176_c233 bl[233] br[233] wl[176] vdd gnd cell_6t
Xbit_r177_c233 bl[233] br[233] wl[177] vdd gnd cell_6t
Xbit_r178_c233 bl[233] br[233] wl[178] vdd gnd cell_6t
Xbit_r179_c233 bl[233] br[233] wl[179] vdd gnd cell_6t
Xbit_r180_c233 bl[233] br[233] wl[180] vdd gnd cell_6t
Xbit_r181_c233 bl[233] br[233] wl[181] vdd gnd cell_6t
Xbit_r182_c233 bl[233] br[233] wl[182] vdd gnd cell_6t
Xbit_r183_c233 bl[233] br[233] wl[183] vdd gnd cell_6t
Xbit_r184_c233 bl[233] br[233] wl[184] vdd gnd cell_6t
Xbit_r185_c233 bl[233] br[233] wl[185] vdd gnd cell_6t
Xbit_r186_c233 bl[233] br[233] wl[186] vdd gnd cell_6t
Xbit_r187_c233 bl[233] br[233] wl[187] vdd gnd cell_6t
Xbit_r188_c233 bl[233] br[233] wl[188] vdd gnd cell_6t
Xbit_r189_c233 bl[233] br[233] wl[189] vdd gnd cell_6t
Xbit_r190_c233 bl[233] br[233] wl[190] vdd gnd cell_6t
Xbit_r191_c233 bl[233] br[233] wl[191] vdd gnd cell_6t
Xbit_r192_c233 bl[233] br[233] wl[192] vdd gnd cell_6t
Xbit_r193_c233 bl[233] br[233] wl[193] vdd gnd cell_6t
Xbit_r194_c233 bl[233] br[233] wl[194] vdd gnd cell_6t
Xbit_r195_c233 bl[233] br[233] wl[195] vdd gnd cell_6t
Xbit_r196_c233 bl[233] br[233] wl[196] vdd gnd cell_6t
Xbit_r197_c233 bl[233] br[233] wl[197] vdd gnd cell_6t
Xbit_r198_c233 bl[233] br[233] wl[198] vdd gnd cell_6t
Xbit_r199_c233 bl[233] br[233] wl[199] vdd gnd cell_6t
Xbit_r200_c233 bl[233] br[233] wl[200] vdd gnd cell_6t
Xbit_r201_c233 bl[233] br[233] wl[201] vdd gnd cell_6t
Xbit_r202_c233 bl[233] br[233] wl[202] vdd gnd cell_6t
Xbit_r203_c233 bl[233] br[233] wl[203] vdd gnd cell_6t
Xbit_r204_c233 bl[233] br[233] wl[204] vdd gnd cell_6t
Xbit_r205_c233 bl[233] br[233] wl[205] vdd gnd cell_6t
Xbit_r206_c233 bl[233] br[233] wl[206] vdd gnd cell_6t
Xbit_r207_c233 bl[233] br[233] wl[207] vdd gnd cell_6t
Xbit_r208_c233 bl[233] br[233] wl[208] vdd gnd cell_6t
Xbit_r209_c233 bl[233] br[233] wl[209] vdd gnd cell_6t
Xbit_r210_c233 bl[233] br[233] wl[210] vdd gnd cell_6t
Xbit_r211_c233 bl[233] br[233] wl[211] vdd gnd cell_6t
Xbit_r212_c233 bl[233] br[233] wl[212] vdd gnd cell_6t
Xbit_r213_c233 bl[233] br[233] wl[213] vdd gnd cell_6t
Xbit_r214_c233 bl[233] br[233] wl[214] vdd gnd cell_6t
Xbit_r215_c233 bl[233] br[233] wl[215] vdd gnd cell_6t
Xbit_r216_c233 bl[233] br[233] wl[216] vdd gnd cell_6t
Xbit_r217_c233 bl[233] br[233] wl[217] vdd gnd cell_6t
Xbit_r218_c233 bl[233] br[233] wl[218] vdd gnd cell_6t
Xbit_r219_c233 bl[233] br[233] wl[219] vdd gnd cell_6t
Xbit_r220_c233 bl[233] br[233] wl[220] vdd gnd cell_6t
Xbit_r221_c233 bl[233] br[233] wl[221] vdd gnd cell_6t
Xbit_r222_c233 bl[233] br[233] wl[222] vdd gnd cell_6t
Xbit_r223_c233 bl[233] br[233] wl[223] vdd gnd cell_6t
Xbit_r224_c233 bl[233] br[233] wl[224] vdd gnd cell_6t
Xbit_r225_c233 bl[233] br[233] wl[225] vdd gnd cell_6t
Xbit_r226_c233 bl[233] br[233] wl[226] vdd gnd cell_6t
Xbit_r227_c233 bl[233] br[233] wl[227] vdd gnd cell_6t
Xbit_r228_c233 bl[233] br[233] wl[228] vdd gnd cell_6t
Xbit_r229_c233 bl[233] br[233] wl[229] vdd gnd cell_6t
Xbit_r230_c233 bl[233] br[233] wl[230] vdd gnd cell_6t
Xbit_r231_c233 bl[233] br[233] wl[231] vdd gnd cell_6t
Xbit_r232_c233 bl[233] br[233] wl[232] vdd gnd cell_6t
Xbit_r233_c233 bl[233] br[233] wl[233] vdd gnd cell_6t
Xbit_r234_c233 bl[233] br[233] wl[234] vdd gnd cell_6t
Xbit_r235_c233 bl[233] br[233] wl[235] vdd gnd cell_6t
Xbit_r236_c233 bl[233] br[233] wl[236] vdd gnd cell_6t
Xbit_r237_c233 bl[233] br[233] wl[237] vdd gnd cell_6t
Xbit_r238_c233 bl[233] br[233] wl[238] vdd gnd cell_6t
Xbit_r239_c233 bl[233] br[233] wl[239] vdd gnd cell_6t
Xbit_r240_c233 bl[233] br[233] wl[240] vdd gnd cell_6t
Xbit_r241_c233 bl[233] br[233] wl[241] vdd gnd cell_6t
Xbit_r242_c233 bl[233] br[233] wl[242] vdd gnd cell_6t
Xbit_r243_c233 bl[233] br[233] wl[243] vdd gnd cell_6t
Xbit_r244_c233 bl[233] br[233] wl[244] vdd gnd cell_6t
Xbit_r245_c233 bl[233] br[233] wl[245] vdd gnd cell_6t
Xbit_r246_c233 bl[233] br[233] wl[246] vdd gnd cell_6t
Xbit_r247_c233 bl[233] br[233] wl[247] vdd gnd cell_6t
Xbit_r248_c233 bl[233] br[233] wl[248] vdd gnd cell_6t
Xbit_r249_c233 bl[233] br[233] wl[249] vdd gnd cell_6t
Xbit_r250_c233 bl[233] br[233] wl[250] vdd gnd cell_6t
Xbit_r251_c233 bl[233] br[233] wl[251] vdd gnd cell_6t
Xbit_r252_c233 bl[233] br[233] wl[252] vdd gnd cell_6t
Xbit_r253_c233 bl[233] br[233] wl[253] vdd gnd cell_6t
Xbit_r254_c233 bl[233] br[233] wl[254] vdd gnd cell_6t
Xbit_r255_c233 bl[233] br[233] wl[255] vdd gnd cell_6t
Xbit_r0_c234 bl[234] br[234] wl[0] vdd gnd cell_6t
Xbit_r1_c234 bl[234] br[234] wl[1] vdd gnd cell_6t
Xbit_r2_c234 bl[234] br[234] wl[2] vdd gnd cell_6t
Xbit_r3_c234 bl[234] br[234] wl[3] vdd gnd cell_6t
Xbit_r4_c234 bl[234] br[234] wl[4] vdd gnd cell_6t
Xbit_r5_c234 bl[234] br[234] wl[5] vdd gnd cell_6t
Xbit_r6_c234 bl[234] br[234] wl[6] vdd gnd cell_6t
Xbit_r7_c234 bl[234] br[234] wl[7] vdd gnd cell_6t
Xbit_r8_c234 bl[234] br[234] wl[8] vdd gnd cell_6t
Xbit_r9_c234 bl[234] br[234] wl[9] vdd gnd cell_6t
Xbit_r10_c234 bl[234] br[234] wl[10] vdd gnd cell_6t
Xbit_r11_c234 bl[234] br[234] wl[11] vdd gnd cell_6t
Xbit_r12_c234 bl[234] br[234] wl[12] vdd gnd cell_6t
Xbit_r13_c234 bl[234] br[234] wl[13] vdd gnd cell_6t
Xbit_r14_c234 bl[234] br[234] wl[14] vdd gnd cell_6t
Xbit_r15_c234 bl[234] br[234] wl[15] vdd gnd cell_6t
Xbit_r16_c234 bl[234] br[234] wl[16] vdd gnd cell_6t
Xbit_r17_c234 bl[234] br[234] wl[17] vdd gnd cell_6t
Xbit_r18_c234 bl[234] br[234] wl[18] vdd gnd cell_6t
Xbit_r19_c234 bl[234] br[234] wl[19] vdd gnd cell_6t
Xbit_r20_c234 bl[234] br[234] wl[20] vdd gnd cell_6t
Xbit_r21_c234 bl[234] br[234] wl[21] vdd gnd cell_6t
Xbit_r22_c234 bl[234] br[234] wl[22] vdd gnd cell_6t
Xbit_r23_c234 bl[234] br[234] wl[23] vdd gnd cell_6t
Xbit_r24_c234 bl[234] br[234] wl[24] vdd gnd cell_6t
Xbit_r25_c234 bl[234] br[234] wl[25] vdd gnd cell_6t
Xbit_r26_c234 bl[234] br[234] wl[26] vdd gnd cell_6t
Xbit_r27_c234 bl[234] br[234] wl[27] vdd gnd cell_6t
Xbit_r28_c234 bl[234] br[234] wl[28] vdd gnd cell_6t
Xbit_r29_c234 bl[234] br[234] wl[29] vdd gnd cell_6t
Xbit_r30_c234 bl[234] br[234] wl[30] vdd gnd cell_6t
Xbit_r31_c234 bl[234] br[234] wl[31] vdd gnd cell_6t
Xbit_r32_c234 bl[234] br[234] wl[32] vdd gnd cell_6t
Xbit_r33_c234 bl[234] br[234] wl[33] vdd gnd cell_6t
Xbit_r34_c234 bl[234] br[234] wl[34] vdd gnd cell_6t
Xbit_r35_c234 bl[234] br[234] wl[35] vdd gnd cell_6t
Xbit_r36_c234 bl[234] br[234] wl[36] vdd gnd cell_6t
Xbit_r37_c234 bl[234] br[234] wl[37] vdd gnd cell_6t
Xbit_r38_c234 bl[234] br[234] wl[38] vdd gnd cell_6t
Xbit_r39_c234 bl[234] br[234] wl[39] vdd gnd cell_6t
Xbit_r40_c234 bl[234] br[234] wl[40] vdd gnd cell_6t
Xbit_r41_c234 bl[234] br[234] wl[41] vdd gnd cell_6t
Xbit_r42_c234 bl[234] br[234] wl[42] vdd gnd cell_6t
Xbit_r43_c234 bl[234] br[234] wl[43] vdd gnd cell_6t
Xbit_r44_c234 bl[234] br[234] wl[44] vdd gnd cell_6t
Xbit_r45_c234 bl[234] br[234] wl[45] vdd gnd cell_6t
Xbit_r46_c234 bl[234] br[234] wl[46] vdd gnd cell_6t
Xbit_r47_c234 bl[234] br[234] wl[47] vdd gnd cell_6t
Xbit_r48_c234 bl[234] br[234] wl[48] vdd gnd cell_6t
Xbit_r49_c234 bl[234] br[234] wl[49] vdd gnd cell_6t
Xbit_r50_c234 bl[234] br[234] wl[50] vdd gnd cell_6t
Xbit_r51_c234 bl[234] br[234] wl[51] vdd gnd cell_6t
Xbit_r52_c234 bl[234] br[234] wl[52] vdd gnd cell_6t
Xbit_r53_c234 bl[234] br[234] wl[53] vdd gnd cell_6t
Xbit_r54_c234 bl[234] br[234] wl[54] vdd gnd cell_6t
Xbit_r55_c234 bl[234] br[234] wl[55] vdd gnd cell_6t
Xbit_r56_c234 bl[234] br[234] wl[56] vdd gnd cell_6t
Xbit_r57_c234 bl[234] br[234] wl[57] vdd gnd cell_6t
Xbit_r58_c234 bl[234] br[234] wl[58] vdd gnd cell_6t
Xbit_r59_c234 bl[234] br[234] wl[59] vdd gnd cell_6t
Xbit_r60_c234 bl[234] br[234] wl[60] vdd gnd cell_6t
Xbit_r61_c234 bl[234] br[234] wl[61] vdd gnd cell_6t
Xbit_r62_c234 bl[234] br[234] wl[62] vdd gnd cell_6t
Xbit_r63_c234 bl[234] br[234] wl[63] vdd gnd cell_6t
Xbit_r64_c234 bl[234] br[234] wl[64] vdd gnd cell_6t
Xbit_r65_c234 bl[234] br[234] wl[65] vdd gnd cell_6t
Xbit_r66_c234 bl[234] br[234] wl[66] vdd gnd cell_6t
Xbit_r67_c234 bl[234] br[234] wl[67] vdd gnd cell_6t
Xbit_r68_c234 bl[234] br[234] wl[68] vdd gnd cell_6t
Xbit_r69_c234 bl[234] br[234] wl[69] vdd gnd cell_6t
Xbit_r70_c234 bl[234] br[234] wl[70] vdd gnd cell_6t
Xbit_r71_c234 bl[234] br[234] wl[71] vdd gnd cell_6t
Xbit_r72_c234 bl[234] br[234] wl[72] vdd gnd cell_6t
Xbit_r73_c234 bl[234] br[234] wl[73] vdd gnd cell_6t
Xbit_r74_c234 bl[234] br[234] wl[74] vdd gnd cell_6t
Xbit_r75_c234 bl[234] br[234] wl[75] vdd gnd cell_6t
Xbit_r76_c234 bl[234] br[234] wl[76] vdd gnd cell_6t
Xbit_r77_c234 bl[234] br[234] wl[77] vdd gnd cell_6t
Xbit_r78_c234 bl[234] br[234] wl[78] vdd gnd cell_6t
Xbit_r79_c234 bl[234] br[234] wl[79] vdd gnd cell_6t
Xbit_r80_c234 bl[234] br[234] wl[80] vdd gnd cell_6t
Xbit_r81_c234 bl[234] br[234] wl[81] vdd gnd cell_6t
Xbit_r82_c234 bl[234] br[234] wl[82] vdd gnd cell_6t
Xbit_r83_c234 bl[234] br[234] wl[83] vdd gnd cell_6t
Xbit_r84_c234 bl[234] br[234] wl[84] vdd gnd cell_6t
Xbit_r85_c234 bl[234] br[234] wl[85] vdd gnd cell_6t
Xbit_r86_c234 bl[234] br[234] wl[86] vdd gnd cell_6t
Xbit_r87_c234 bl[234] br[234] wl[87] vdd gnd cell_6t
Xbit_r88_c234 bl[234] br[234] wl[88] vdd gnd cell_6t
Xbit_r89_c234 bl[234] br[234] wl[89] vdd gnd cell_6t
Xbit_r90_c234 bl[234] br[234] wl[90] vdd gnd cell_6t
Xbit_r91_c234 bl[234] br[234] wl[91] vdd gnd cell_6t
Xbit_r92_c234 bl[234] br[234] wl[92] vdd gnd cell_6t
Xbit_r93_c234 bl[234] br[234] wl[93] vdd gnd cell_6t
Xbit_r94_c234 bl[234] br[234] wl[94] vdd gnd cell_6t
Xbit_r95_c234 bl[234] br[234] wl[95] vdd gnd cell_6t
Xbit_r96_c234 bl[234] br[234] wl[96] vdd gnd cell_6t
Xbit_r97_c234 bl[234] br[234] wl[97] vdd gnd cell_6t
Xbit_r98_c234 bl[234] br[234] wl[98] vdd gnd cell_6t
Xbit_r99_c234 bl[234] br[234] wl[99] vdd gnd cell_6t
Xbit_r100_c234 bl[234] br[234] wl[100] vdd gnd cell_6t
Xbit_r101_c234 bl[234] br[234] wl[101] vdd gnd cell_6t
Xbit_r102_c234 bl[234] br[234] wl[102] vdd gnd cell_6t
Xbit_r103_c234 bl[234] br[234] wl[103] vdd gnd cell_6t
Xbit_r104_c234 bl[234] br[234] wl[104] vdd gnd cell_6t
Xbit_r105_c234 bl[234] br[234] wl[105] vdd gnd cell_6t
Xbit_r106_c234 bl[234] br[234] wl[106] vdd gnd cell_6t
Xbit_r107_c234 bl[234] br[234] wl[107] vdd gnd cell_6t
Xbit_r108_c234 bl[234] br[234] wl[108] vdd gnd cell_6t
Xbit_r109_c234 bl[234] br[234] wl[109] vdd gnd cell_6t
Xbit_r110_c234 bl[234] br[234] wl[110] vdd gnd cell_6t
Xbit_r111_c234 bl[234] br[234] wl[111] vdd gnd cell_6t
Xbit_r112_c234 bl[234] br[234] wl[112] vdd gnd cell_6t
Xbit_r113_c234 bl[234] br[234] wl[113] vdd gnd cell_6t
Xbit_r114_c234 bl[234] br[234] wl[114] vdd gnd cell_6t
Xbit_r115_c234 bl[234] br[234] wl[115] vdd gnd cell_6t
Xbit_r116_c234 bl[234] br[234] wl[116] vdd gnd cell_6t
Xbit_r117_c234 bl[234] br[234] wl[117] vdd gnd cell_6t
Xbit_r118_c234 bl[234] br[234] wl[118] vdd gnd cell_6t
Xbit_r119_c234 bl[234] br[234] wl[119] vdd gnd cell_6t
Xbit_r120_c234 bl[234] br[234] wl[120] vdd gnd cell_6t
Xbit_r121_c234 bl[234] br[234] wl[121] vdd gnd cell_6t
Xbit_r122_c234 bl[234] br[234] wl[122] vdd gnd cell_6t
Xbit_r123_c234 bl[234] br[234] wl[123] vdd gnd cell_6t
Xbit_r124_c234 bl[234] br[234] wl[124] vdd gnd cell_6t
Xbit_r125_c234 bl[234] br[234] wl[125] vdd gnd cell_6t
Xbit_r126_c234 bl[234] br[234] wl[126] vdd gnd cell_6t
Xbit_r127_c234 bl[234] br[234] wl[127] vdd gnd cell_6t
Xbit_r128_c234 bl[234] br[234] wl[128] vdd gnd cell_6t
Xbit_r129_c234 bl[234] br[234] wl[129] vdd gnd cell_6t
Xbit_r130_c234 bl[234] br[234] wl[130] vdd gnd cell_6t
Xbit_r131_c234 bl[234] br[234] wl[131] vdd gnd cell_6t
Xbit_r132_c234 bl[234] br[234] wl[132] vdd gnd cell_6t
Xbit_r133_c234 bl[234] br[234] wl[133] vdd gnd cell_6t
Xbit_r134_c234 bl[234] br[234] wl[134] vdd gnd cell_6t
Xbit_r135_c234 bl[234] br[234] wl[135] vdd gnd cell_6t
Xbit_r136_c234 bl[234] br[234] wl[136] vdd gnd cell_6t
Xbit_r137_c234 bl[234] br[234] wl[137] vdd gnd cell_6t
Xbit_r138_c234 bl[234] br[234] wl[138] vdd gnd cell_6t
Xbit_r139_c234 bl[234] br[234] wl[139] vdd gnd cell_6t
Xbit_r140_c234 bl[234] br[234] wl[140] vdd gnd cell_6t
Xbit_r141_c234 bl[234] br[234] wl[141] vdd gnd cell_6t
Xbit_r142_c234 bl[234] br[234] wl[142] vdd gnd cell_6t
Xbit_r143_c234 bl[234] br[234] wl[143] vdd gnd cell_6t
Xbit_r144_c234 bl[234] br[234] wl[144] vdd gnd cell_6t
Xbit_r145_c234 bl[234] br[234] wl[145] vdd gnd cell_6t
Xbit_r146_c234 bl[234] br[234] wl[146] vdd gnd cell_6t
Xbit_r147_c234 bl[234] br[234] wl[147] vdd gnd cell_6t
Xbit_r148_c234 bl[234] br[234] wl[148] vdd gnd cell_6t
Xbit_r149_c234 bl[234] br[234] wl[149] vdd gnd cell_6t
Xbit_r150_c234 bl[234] br[234] wl[150] vdd gnd cell_6t
Xbit_r151_c234 bl[234] br[234] wl[151] vdd gnd cell_6t
Xbit_r152_c234 bl[234] br[234] wl[152] vdd gnd cell_6t
Xbit_r153_c234 bl[234] br[234] wl[153] vdd gnd cell_6t
Xbit_r154_c234 bl[234] br[234] wl[154] vdd gnd cell_6t
Xbit_r155_c234 bl[234] br[234] wl[155] vdd gnd cell_6t
Xbit_r156_c234 bl[234] br[234] wl[156] vdd gnd cell_6t
Xbit_r157_c234 bl[234] br[234] wl[157] vdd gnd cell_6t
Xbit_r158_c234 bl[234] br[234] wl[158] vdd gnd cell_6t
Xbit_r159_c234 bl[234] br[234] wl[159] vdd gnd cell_6t
Xbit_r160_c234 bl[234] br[234] wl[160] vdd gnd cell_6t
Xbit_r161_c234 bl[234] br[234] wl[161] vdd gnd cell_6t
Xbit_r162_c234 bl[234] br[234] wl[162] vdd gnd cell_6t
Xbit_r163_c234 bl[234] br[234] wl[163] vdd gnd cell_6t
Xbit_r164_c234 bl[234] br[234] wl[164] vdd gnd cell_6t
Xbit_r165_c234 bl[234] br[234] wl[165] vdd gnd cell_6t
Xbit_r166_c234 bl[234] br[234] wl[166] vdd gnd cell_6t
Xbit_r167_c234 bl[234] br[234] wl[167] vdd gnd cell_6t
Xbit_r168_c234 bl[234] br[234] wl[168] vdd gnd cell_6t
Xbit_r169_c234 bl[234] br[234] wl[169] vdd gnd cell_6t
Xbit_r170_c234 bl[234] br[234] wl[170] vdd gnd cell_6t
Xbit_r171_c234 bl[234] br[234] wl[171] vdd gnd cell_6t
Xbit_r172_c234 bl[234] br[234] wl[172] vdd gnd cell_6t
Xbit_r173_c234 bl[234] br[234] wl[173] vdd gnd cell_6t
Xbit_r174_c234 bl[234] br[234] wl[174] vdd gnd cell_6t
Xbit_r175_c234 bl[234] br[234] wl[175] vdd gnd cell_6t
Xbit_r176_c234 bl[234] br[234] wl[176] vdd gnd cell_6t
Xbit_r177_c234 bl[234] br[234] wl[177] vdd gnd cell_6t
Xbit_r178_c234 bl[234] br[234] wl[178] vdd gnd cell_6t
Xbit_r179_c234 bl[234] br[234] wl[179] vdd gnd cell_6t
Xbit_r180_c234 bl[234] br[234] wl[180] vdd gnd cell_6t
Xbit_r181_c234 bl[234] br[234] wl[181] vdd gnd cell_6t
Xbit_r182_c234 bl[234] br[234] wl[182] vdd gnd cell_6t
Xbit_r183_c234 bl[234] br[234] wl[183] vdd gnd cell_6t
Xbit_r184_c234 bl[234] br[234] wl[184] vdd gnd cell_6t
Xbit_r185_c234 bl[234] br[234] wl[185] vdd gnd cell_6t
Xbit_r186_c234 bl[234] br[234] wl[186] vdd gnd cell_6t
Xbit_r187_c234 bl[234] br[234] wl[187] vdd gnd cell_6t
Xbit_r188_c234 bl[234] br[234] wl[188] vdd gnd cell_6t
Xbit_r189_c234 bl[234] br[234] wl[189] vdd gnd cell_6t
Xbit_r190_c234 bl[234] br[234] wl[190] vdd gnd cell_6t
Xbit_r191_c234 bl[234] br[234] wl[191] vdd gnd cell_6t
Xbit_r192_c234 bl[234] br[234] wl[192] vdd gnd cell_6t
Xbit_r193_c234 bl[234] br[234] wl[193] vdd gnd cell_6t
Xbit_r194_c234 bl[234] br[234] wl[194] vdd gnd cell_6t
Xbit_r195_c234 bl[234] br[234] wl[195] vdd gnd cell_6t
Xbit_r196_c234 bl[234] br[234] wl[196] vdd gnd cell_6t
Xbit_r197_c234 bl[234] br[234] wl[197] vdd gnd cell_6t
Xbit_r198_c234 bl[234] br[234] wl[198] vdd gnd cell_6t
Xbit_r199_c234 bl[234] br[234] wl[199] vdd gnd cell_6t
Xbit_r200_c234 bl[234] br[234] wl[200] vdd gnd cell_6t
Xbit_r201_c234 bl[234] br[234] wl[201] vdd gnd cell_6t
Xbit_r202_c234 bl[234] br[234] wl[202] vdd gnd cell_6t
Xbit_r203_c234 bl[234] br[234] wl[203] vdd gnd cell_6t
Xbit_r204_c234 bl[234] br[234] wl[204] vdd gnd cell_6t
Xbit_r205_c234 bl[234] br[234] wl[205] vdd gnd cell_6t
Xbit_r206_c234 bl[234] br[234] wl[206] vdd gnd cell_6t
Xbit_r207_c234 bl[234] br[234] wl[207] vdd gnd cell_6t
Xbit_r208_c234 bl[234] br[234] wl[208] vdd gnd cell_6t
Xbit_r209_c234 bl[234] br[234] wl[209] vdd gnd cell_6t
Xbit_r210_c234 bl[234] br[234] wl[210] vdd gnd cell_6t
Xbit_r211_c234 bl[234] br[234] wl[211] vdd gnd cell_6t
Xbit_r212_c234 bl[234] br[234] wl[212] vdd gnd cell_6t
Xbit_r213_c234 bl[234] br[234] wl[213] vdd gnd cell_6t
Xbit_r214_c234 bl[234] br[234] wl[214] vdd gnd cell_6t
Xbit_r215_c234 bl[234] br[234] wl[215] vdd gnd cell_6t
Xbit_r216_c234 bl[234] br[234] wl[216] vdd gnd cell_6t
Xbit_r217_c234 bl[234] br[234] wl[217] vdd gnd cell_6t
Xbit_r218_c234 bl[234] br[234] wl[218] vdd gnd cell_6t
Xbit_r219_c234 bl[234] br[234] wl[219] vdd gnd cell_6t
Xbit_r220_c234 bl[234] br[234] wl[220] vdd gnd cell_6t
Xbit_r221_c234 bl[234] br[234] wl[221] vdd gnd cell_6t
Xbit_r222_c234 bl[234] br[234] wl[222] vdd gnd cell_6t
Xbit_r223_c234 bl[234] br[234] wl[223] vdd gnd cell_6t
Xbit_r224_c234 bl[234] br[234] wl[224] vdd gnd cell_6t
Xbit_r225_c234 bl[234] br[234] wl[225] vdd gnd cell_6t
Xbit_r226_c234 bl[234] br[234] wl[226] vdd gnd cell_6t
Xbit_r227_c234 bl[234] br[234] wl[227] vdd gnd cell_6t
Xbit_r228_c234 bl[234] br[234] wl[228] vdd gnd cell_6t
Xbit_r229_c234 bl[234] br[234] wl[229] vdd gnd cell_6t
Xbit_r230_c234 bl[234] br[234] wl[230] vdd gnd cell_6t
Xbit_r231_c234 bl[234] br[234] wl[231] vdd gnd cell_6t
Xbit_r232_c234 bl[234] br[234] wl[232] vdd gnd cell_6t
Xbit_r233_c234 bl[234] br[234] wl[233] vdd gnd cell_6t
Xbit_r234_c234 bl[234] br[234] wl[234] vdd gnd cell_6t
Xbit_r235_c234 bl[234] br[234] wl[235] vdd gnd cell_6t
Xbit_r236_c234 bl[234] br[234] wl[236] vdd gnd cell_6t
Xbit_r237_c234 bl[234] br[234] wl[237] vdd gnd cell_6t
Xbit_r238_c234 bl[234] br[234] wl[238] vdd gnd cell_6t
Xbit_r239_c234 bl[234] br[234] wl[239] vdd gnd cell_6t
Xbit_r240_c234 bl[234] br[234] wl[240] vdd gnd cell_6t
Xbit_r241_c234 bl[234] br[234] wl[241] vdd gnd cell_6t
Xbit_r242_c234 bl[234] br[234] wl[242] vdd gnd cell_6t
Xbit_r243_c234 bl[234] br[234] wl[243] vdd gnd cell_6t
Xbit_r244_c234 bl[234] br[234] wl[244] vdd gnd cell_6t
Xbit_r245_c234 bl[234] br[234] wl[245] vdd gnd cell_6t
Xbit_r246_c234 bl[234] br[234] wl[246] vdd gnd cell_6t
Xbit_r247_c234 bl[234] br[234] wl[247] vdd gnd cell_6t
Xbit_r248_c234 bl[234] br[234] wl[248] vdd gnd cell_6t
Xbit_r249_c234 bl[234] br[234] wl[249] vdd gnd cell_6t
Xbit_r250_c234 bl[234] br[234] wl[250] vdd gnd cell_6t
Xbit_r251_c234 bl[234] br[234] wl[251] vdd gnd cell_6t
Xbit_r252_c234 bl[234] br[234] wl[252] vdd gnd cell_6t
Xbit_r253_c234 bl[234] br[234] wl[253] vdd gnd cell_6t
Xbit_r254_c234 bl[234] br[234] wl[254] vdd gnd cell_6t
Xbit_r255_c234 bl[234] br[234] wl[255] vdd gnd cell_6t
Xbit_r0_c235 bl[235] br[235] wl[0] vdd gnd cell_6t
Xbit_r1_c235 bl[235] br[235] wl[1] vdd gnd cell_6t
Xbit_r2_c235 bl[235] br[235] wl[2] vdd gnd cell_6t
Xbit_r3_c235 bl[235] br[235] wl[3] vdd gnd cell_6t
Xbit_r4_c235 bl[235] br[235] wl[4] vdd gnd cell_6t
Xbit_r5_c235 bl[235] br[235] wl[5] vdd gnd cell_6t
Xbit_r6_c235 bl[235] br[235] wl[6] vdd gnd cell_6t
Xbit_r7_c235 bl[235] br[235] wl[7] vdd gnd cell_6t
Xbit_r8_c235 bl[235] br[235] wl[8] vdd gnd cell_6t
Xbit_r9_c235 bl[235] br[235] wl[9] vdd gnd cell_6t
Xbit_r10_c235 bl[235] br[235] wl[10] vdd gnd cell_6t
Xbit_r11_c235 bl[235] br[235] wl[11] vdd gnd cell_6t
Xbit_r12_c235 bl[235] br[235] wl[12] vdd gnd cell_6t
Xbit_r13_c235 bl[235] br[235] wl[13] vdd gnd cell_6t
Xbit_r14_c235 bl[235] br[235] wl[14] vdd gnd cell_6t
Xbit_r15_c235 bl[235] br[235] wl[15] vdd gnd cell_6t
Xbit_r16_c235 bl[235] br[235] wl[16] vdd gnd cell_6t
Xbit_r17_c235 bl[235] br[235] wl[17] vdd gnd cell_6t
Xbit_r18_c235 bl[235] br[235] wl[18] vdd gnd cell_6t
Xbit_r19_c235 bl[235] br[235] wl[19] vdd gnd cell_6t
Xbit_r20_c235 bl[235] br[235] wl[20] vdd gnd cell_6t
Xbit_r21_c235 bl[235] br[235] wl[21] vdd gnd cell_6t
Xbit_r22_c235 bl[235] br[235] wl[22] vdd gnd cell_6t
Xbit_r23_c235 bl[235] br[235] wl[23] vdd gnd cell_6t
Xbit_r24_c235 bl[235] br[235] wl[24] vdd gnd cell_6t
Xbit_r25_c235 bl[235] br[235] wl[25] vdd gnd cell_6t
Xbit_r26_c235 bl[235] br[235] wl[26] vdd gnd cell_6t
Xbit_r27_c235 bl[235] br[235] wl[27] vdd gnd cell_6t
Xbit_r28_c235 bl[235] br[235] wl[28] vdd gnd cell_6t
Xbit_r29_c235 bl[235] br[235] wl[29] vdd gnd cell_6t
Xbit_r30_c235 bl[235] br[235] wl[30] vdd gnd cell_6t
Xbit_r31_c235 bl[235] br[235] wl[31] vdd gnd cell_6t
Xbit_r32_c235 bl[235] br[235] wl[32] vdd gnd cell_6t
Xbit_r33_c235 bl[235] br[235] wl[33] vdd gnd cell_6t
Xbit_r34_c235 bl[235] br[235] wl[34] vdd gnd cell_6t
Xbit_r35_c235 bl[235] br[235] wl[35] vdd gnd cell_6t
Xbit_r36_c235 bl[235] br[235] wl[36] vdd gnd cell_6t
Xbit_r37_c235 bl[235] br[235] wl[37] vdd gnd cell_6t
Xbit_r38_c235 bl[235] br[235] wl[38] vdd gnd cell_6t
Xbit_r39_c235 bl[235] br[235] wl[39] vdd gnd cell_6t
Xbit_r40_c235 bl[235] br[235] wl[40] vdd gnd cell_6t
Xbit_r41_c235 bl[235] br[235] wl[41] vdd gnd cell_6t
Xbit_r42_c235 bl[235] br[235] wl[42] vdd gnd cell_6t
Xbit_r43_c235 bl[235] br[235] wl[43] vdd gnd cell_6t
Xbit_r44_c235 bl[235] br[235] wl[44] vdd gnd cell_6t
Xbit_r45_c235 bl[235] br[235] wl[45] vdd gnd cell_6t
Xbit_r46_c235 bl[235] br[235] wl[46] vdd gnd cell_6t
Xbit_r47_c235 bl[235] br[235] wl[47] vdd gnd cell_6t
Xbit_r48_c235 bl[235] br[235] wl[48] vdd gnd cell_6t
Xbit_r49_c235 bl[235] br[235] wl[49] vdd gnd cell_6t
Xbit_r50_c235 bl[235] br[235] wl[50] vdd gnd cell_6t
Xbit_r51_c235 bl[235] br[235] wl[51] vdd gnd cell_6t
Xbit_r52_c235 bl[235] br[235] wl[52] vdd gnd cell_6t
Xbit_r53_c235 bl[235] br[235] wl[53] vdd gnd cell_6t
Xbit_r54_c235 bl[235] br[235] wl[54] vdd gnd cell_6t
Xbit_r55_c235 bl[235] br[235] wl[55] vdd gnd cell_6t
Xbit_r56_c235 bl[235] br[235] wl[56] vdd gnd cell_6t
Xbit_r57_c235 bl[235] br[235] wl[57] vdd gnd cell_6t
Xbit_r58_c235 bl[235] br[235] wl[58] vdd gnd cell_6t
Xbit_r59_c235 bl[235] br[235] wl[59] vdd gnd cell_6t
Xbit_r60_c235 bl[235] br[235] wl[60] vdd gnd cell_6t
Xbit_r61_c235 bl[235] br[235] wl[61] vdd gnd cell_6t
Xbit_r62_c235 bl[235] br[235] wl[62] vdd gnd cell_6t
Xbit_r63_c235 bl[235] br[235] wl[63] vdd gnd cell_6t
Xbit_r64_c235 bl[235] br[235] wl[64] vdd gnd cell_6t
Xbit_r65_c235 bl[235] br[235] wl[65] vdd gnd cell_6t
Xbit_r66_c235 bl[235] br[235] wl[66] vdd gnd cell_6t
Xbit_r67_c235 bl[235] br[235] wl[67] vdd gnd cell_6t
Xbit_r68_c235 bl[235] br[235] wl[68] vdd gnd cell_6t
Xbit_r69_c235 bl[235] br[235] wl[69] vdd gnd cell_6t
Xbit_r70_c235 bl[235] br[235] wl[70] vdd gnd cell_6t
Xbit_r71_c235 bl[235] br[235] wl[71] vdd gnd cell_6t
Xbit_r72_c235 bl[235] br[235] wl[72] vdd gnd cell_6t
Xbit_r73_c235 bl[235] br[235] wl[73] vdd gnd cell_6t
Xbit_r74_c235 bl[235] br[235] wl[74] vdd gnd cell_6t
Xbit_r75_c235 bl[235] br[235] wl[75] vdd gnd cell_6t
Xbit_r76_c235 bl[235] br[235] wl[76] vdd gnd cell_6t
Xbit_r77_c235 bl[235] br[235] wl[77] vdd gnd cell_6t
Xbit_r78_c235 bl[235] br[235] wl[78] vdd gnd cell_6t
Xbit_r79_c235 bl[235] br[235] wl[79] vdd gnd cell_6t
Xbit_r80_c235 bl[235] br[235] wl[80] vdd gnd cell_6t
Xbit_r81_c235 bl[235] br[235] wl[81] vdd gnd cell_6t
Xbit_r82_c235 bl[235] br[235] wl[82] vdd gnd cell_6t
Xbit_r83_c235 bl[235] br[235] wl[83] vdd gnd cell_6t
Xbit_r84_c235 bl[235] br[235] wl[84] vdd gnd cell_6t
Xbit_r85_c235 bl[235] br[235] wl[85] vdd gnd cell_6t
Xbit_r86_c235 bl[235] br[235] wl[86] vdd gnd cell_6t
Xbit_r87_c235 bl[235] br[235] wl[87] vdd gnd cell_6t
Xbit_r88_c235 bl[235] br[235] wl[88] vdd gnd cell_6t
Xbit_r89_c235 bl[235] br[235] wl[89] vdd gnd cell_6t
Xbit_r90_c235 bl[235] br[235] wl[90] vdd gnd cell_6t
Xbit_r91_c235 bl[235] br[235] wl[91] vdd gnd cell_6t
Xbit_r92_c235 bl[235] br[235] wl[92] vdd gnd cell_6t
Xbit_r93_c235 bl[235] br[235] wl[93] vdd gnd cell_6t
Xbit_r94_c235 bl[235] br[235] wl[94] vdd gnd cell_6t
Xbit_r95_c235 bl[235] br[235] wl[95] vdd gnd cell_6t
Xbit_r96_c235 bl[235] br[235] wl[96] vdd gnd cell_6t
Xbit_r97_c235 bl[235] br[235] wl[97] vdd gnd cell_6t
Xbit_r98_c235 bl[235] br[235] wl[98] vdd gnd cell_6t
Xbit_r99_c235 bl[235] br[235] wl[99] vdd gnd cell_6t
Xbit_r100_c235 bl[235] br[235] wl[100] vdd gnd cell_6t
Xbit_r101_c235 bl[235] br[235] wl[101] vdd gnd cell_6t
Xbit_r102_c235 bl[235] br[235] wl[102] vdd gnd cell_6t
Xbit_r103_c235 bl[235] br[235] wl[103] vdd gnd cell_6t
Xbit_r104_c235 bl[235] br[235] wl[104] vdd gnd cell_6t
Xbit_r105_c235 bl[235] br[235] wl[105] vdd gnd cell_6t
Xbit_r106_c235 bl[235] br[235] wl[106] vdd gnd cell_6t
Xbit_r107_c235 bl[235] br[235] wl[107] vdd gnd cell_6t
Xbit_r108_c235 bl[235] br[235] wl[108] vdd gnd cell_6t
Xbit_r109_c235 bl[235] br[235] wl[109] vdd gnd cell_6t
Xbit_r110_c235 bl[235] br[235] wl[110] vdd gnd cell_6t
Xbit_r111_c235 bl[235] br[235] wl[111] vdd gnd cell_6t
Xbit_r112_c235 bl[235] br[235] wl[112] vdd gnd cell_6t
Xbit_r113_c235 bl[235] br[235] wl[113] vdd gnd cell_6t
Xbit_r114_c235 bl[235] br[235] wl[114] vdd gnd cell_6t
Xbit_r115_c235 bl[235] br[235] wl[115] vdd gnd cell_6t
Xbit_r116_c235 bl[235] br[235] wl[116] vdd gnd cell_6t
Xbit_r117_c235 bl[235] br[235] wl[117] vdd gnd cell_6t
Xbit_r118_c235 bl[235] br[235] wl[118] vdd gnd cell_6t
Xbit_r119_c235 bl[235] br[235] wl[119] vdd gnd cell_6t
Xbit_r120_c235 bl[235] br[235] wl[120] vdd gnd cell_6t
Xbit_r121_c235 bl[235] br[235] wl[121] vdd gnd cell_6t
Xbit_r122_c235 bl[235] br[235] wl[122] vdd gnd cell_6t
Xbit_r123_c235 bl[235] br[235] wl[123] vdd gnd cell_6t
Xbit_r124_c235 bl[235] br[235] wl[124] vdd gnd cell_6t
Xbit_r125_c235 bl[235] br[235] wl[125] vdd gnd cell_6t
Xbit_r126_c235 bl[235] br[235] wl[126] vdd gnd cell_6t
Xbit_r127_c235 bl[235] br[235] wl[127] vdd gnd cell_6t
Xbit_r128_c235 bl[235] br[235] wl[128] vdd gnd cell_6t
Xbit_r129_c235 bl[235] br[235] wl[129] vdd gnd cell_6t
Xbit_r130_c235 bl[235] br[235] wl[130] vdd gnd cell_6t
Xbit_r131_c235 bl[235] br[235] wl[131] vdd gnd cell_6t
Xbit_r132_c235 bl[235] br[235] wl[132] vdd gnd cell_6t
Xbit_r133_c235 bl[235] br[235] wl[133] vdd gnd cell_6t
Xbit_r134_c235 bl[235] br[235] wl[134] vdd gnd cell_6t
Xbit_r135_c235 bl[235] br[235] wl[135] vdd gnd cell_6t
Xbit_r136_c235 bl[235] br[235] wl[136] vdd gnd cell_6t
Xbit_r137_c235 bl[235] br[235] wl[137] vdd gnd cell_6t
Xbit_r138_c235 bl[235] br[235] wl[138] vdd gnd cell_6t
Xbit_r139_c235 bl[235] br[235] wl[139] vdd gnd cell_6t
Xbit_r140_c235 bl[235] br[235] wl[140] vdd gnd cell_6t
Xbit_r141_c235 bl[235] br[235] wl[141] vdd gnd cell_6t
Xbit_r142_c235 bl[235] br[235] wl[142] vdd gnd cell_6t
Xbit_r143_c235 bl[235] br[235] wl[143] vdd gnd cell_6t
Xbit_r144_c235 bl[235] br[235] wl[144] vdd gnd cell_6t
Xbit_r145_c235 bl[235] br[235] wl[145] vdd gnd cell_6t
Xbit_r146_c235 bl[235] br[235] wl[146] vdd gnd cell_6t
Xbit_r147_c235 bl[235] br[235] wl[147] vdd gnd cell_6t
Xbit_r148_c235 bl[235] br[235] wl[148] vdd gnd cell_6t
Xbit_r149_c235 bl[235] br[235] wl[149] vdd gnd cell_6t
Xbit_r150_c235 bl[235] br[235] wl[150] vdd gnd cell_6t
Xbit_r151_c235 bl[235] br[235] wl[151] vdd gnd cell_6t
Xbit_r152_c235 bl[235] br[235] wl[152] vdd gnd cell_6t
Xbit_r153_c235 bl[235] br[235] wl[153] vdd gnd cell_6t
Xbit_r154_c235 bl[235] br[235] wl[154] vdd gnd cell_6t
Xbit_r155_c235 bl[235] br[235] wl[155] vdd gnd cell_6t
Xbit_r156_c235 bl[235] br[235] wl[156] vdd gnd cell_6t
Xbit_r157_c235 bl[235] br[235] wl[157] vdd gnd cell_6t
Xbit_r158_c235 bl[235] br[235] wl[158] vdd gnd cell_6t
Xbit_r159_c235 bl[235] br[235] wl[159] vdd gnd cell_6t
Xbit_r160_c235 bl[235] br[235] wl[160] vdd gnd cell_6t
Xbit_r161_c235 bl[235] br[235] wl[161] vdd gnd cell_6t
Xbit_r162_c235 bl[235] br[235] wl[162] vdd gnd cell_6t
Xbit_r163_c235 bl[235] br[235] wl[163] vdd gnd cell_6t
Xbit_r164_c235 bl[235] br[235] wl[164] vdd gnd cell_6t
Xbit_r165_c235 bl[235] br[235] wl[165] vdd gnd cell_6t
Xbit_r166_c235 bl[235] br[235] wl[166] vdd gnd cell_6t
Xbit_r167_c235 bl[235] br[235] wl[167] vdd gnd cell_6t
Xbit_r168_c235 bl[235] br[235] wl[168] vdd gnd cell_6t
Xbit_r169_c235 bl[235] br[235] wl[169] vdd gnd cell_6t
Xbit_r170_c235 bl[235] br[235] wl[170] vdd gnd cell_6t
Xbit_r171_c235 bl[235] br[235] wl[171] vdd gnd cell_6t
Xbit_r172_c235 bl[235] br[235] wl[172] vdd gnd cell_6t
Xbit_r173_c235 bl[235] br[235] wl[173] vdd gnd cell_6t
Xbit_r174_c235 bl[235] br[235] wl[174] vdd gnd cell_6t
Xbit_r175_c235 bl[235] br[235] wl[175] vdd gnd cell_6t
Xbit_r176_c235 bl[235] br[235] wl[176] vdd gnd cell_6t
Xbit_r177_c235 bl[235] br[235] wl[177] vdd gnd cell_6t
Xbit_r178_c235 bl[235] br[235] wl[178] vdd gnd cell_6t
Xbit_r179_c235 bl[235] br[235] wl[179] vdd gnd cell_6t
Xbit_r180_c235 bl[235] br[235] wl[180] vdd gnd cell_6t
Xbit_r181_c235 bl[235] br[235] wl[181] vdd gnd cell_6t
Xbit_r182_c235 bl[235] br[235] wl[182] vdd gnd cell_6t
Xbit_r183_c235 bl[235] br[235] wl[183] vdd gnd cell_6t
Xbit_r184_c235 bl[235] br[235] wl[184] vdd gnd cell_6t
Xbit_r185_c235 bl[235] br[235] wl[185] vdd gnd cell_6t
Xbit_r186_c235 bl[235] br[235] wl[186] vdd gnd cell_6t
Xbit_r187_c235 bl[235] br[235] wl[187] vdd gnd cell_6t
Xbit_r188_c235 bl[235] br[235] wl[188] vdd gnd cell_6t
Xbit_r189_c235 bl[235] br[235] wl[189] vdd gnd cell_6t
Xbit_r190_c235 bl[235] br[235] wl[190] vdd gnd cell_6t
Xbit_r191_c235 bl[235] br[235] wl[191] vdd gnd cell_6t
Xbit_r192_c235 bl[235] br[235] wl[192] vdd gnd cell_6t
Xbit_r193_c235 bl[235] br[235] wl[193] vdd gnd cell_6t
Xbit_r194_c235 bl[235] br[235] wl[194] vdd gnd cell_6t
Xbit_r195_c235 bl[235] br[235] wl[195] vdd gnd cell_6t
Xbit_r196_c235 bl[235] br[235] wl[196] vdd gnd cell_6t
Xbit_r197_c235 bl[235] br[235] wl[197] vdd gnd cell_6t
Xbit_r198_c235 bl[235] br[235] wl[198] vdd gnd cell_6t
Xbit_r199_c235 bl[235] br[235] wl[199] vdd gnd cell_6t
Xbit_r200_c235 bl[235] br[235] wl[200] vdd gnd cell_6t
Xbit_r201_c235 bl[235] br[235] wl[201] vdd gnd cell_6t
Xbit_r202_c235 bl[235] br[235] wl[202] vdd gnd cell_6t
Xbit_r203_c235 bl[235] br[235] wl[203] vdd gnd cell_6t
Xbit_r204_c235 bl[235] br[235] wl[204] vdd gnd cell_6t
Xbit_r205_c235 bl[235] br[235] wl[205] vdd gnd cell_6t
Xbit_r206_c235 bl[235] br[235] wl[206] vdd gnd cell_6t
Xbit_r207_c235 bl[235] br[235] wl[207] vdd gnd cell_6t
Xbit_r208_c235 bl[235] br[235] wl[208] vdd gnd cell_6t
Xbit_r209_c235 bl[235] br[235] wl[209] vdd gnd cell_6t
Xbit_r210_c235 bl[235] br[235] wl[210] vdd gnd cell_6t
Xbit_r211_c235 bl[235] br[235] wl[211] vdd gnd cell_6t
Xbit_r212_c235 bl[235] br[235] wl[212] vdd gnd cell_6t
Xbit_r213_c235 bl[235] br[235] wl[213] vdd gnd cell_6t
Xbit_r214_c235 bl[235] br[235] wl[214] vdd gnd cell_6t
Xbit_r215_c235 bl[235] br[235] wl[215] vdd gnd cell_6t
Xbit_r216_c235 bl[235] br[235] wl[216] vdd gnd cell_6t
Xbit_r217_c235 bl[235] br[235] wl[217] vdd gnd cell_6t
Xbit_r218_c235 bl[235] br[235] wl[218] vdd gnd cell_6t
Xbit_r219_c235 bl[235] br[235] wl[219] vdd gnd cell_6t
Xbit_r220_c235 bl[235] br[235] wl[220] vdd gnd cell_6t
Xbit_r221_c235 bl[235] br[235] wl[221] vdd gnd cell_6t
Xbit_r222_c235 bl[235] br[235] wl[222] vdd gnd cell_6t
Xbit_r223_c235 bl[235] br[235] wl[223] vdd gnd cell_6t
Xbit_r224_c235 bl[235] br[235] wl[224] vdd gnd cell_6t
Xbit_r225_c235 bl[235] br[235] wl[225] vdd gnd cell_6t
Xbit_r226_c235 bl[235] br[235] wl[226] vdd gnd cell_6t
Xbit_r227_c235 bl[235] br[235] wl[227] vdd gnd cell_6t
Xbit_r228_c235 bl[235] br[235] wl[228] vdd gnd cell_6t
Xbit_r229_c235 bl[235] br[235] wl[229] vdd gnd cell_6t
Xbit_r230_c235 bl[235] br[235] wl[230] vdd gnd cell_6t
Xbit_r231_c235 bl[235] br[235] wl[231] vdd gnd cell_6t
Xbit_r232_c235 bl[235] br[235] wl[232] vdd gnd cell_6t
Xbit_r233_c235 bl[235] br[235] wl[233] vdd gnd cell_6t
Xbit_r234_c235 bl[235] br[235] wl[234] vdd gnd cell_6t
Xbit_r235_c235 bl[235] br[235] wl[235] vdd gnd cell_6t
Xbit_r236_c235 bl[235] br[235] wl[236] vdd gnd cell_6t
Xbit_r237_c235 bl[235] br[235] wl[237] vdd gnd cell_6t
Xbit_r238_c235 bl[235] br[235] wl[238] vdd gnd cell_6t
Xbit_r239_c235 bl[235] br[235] wl[239] vdd gnd cell_6t
Xbit_r240_c235 bl[235] br[235] wl[240] vdd gnd cell_6t
Xbit_r241_c235 bl[235] br[235] wl[241] vdd gnd cell_6t
Xbit_r242_c235 bl[235] br[235] wl[242] vdd gnd cell_6t
Xbit_r243_c235 bl[235] br[235] wl[243] vdd gnd cell_6t
Xbit_r244_c235 bl[235] br[235] wl[244] vdd gnd cell_6t
Xbit_r245_c235 bl[235] br[235] wl[245] vdd gnd cell_6t
Xbit_r246_c235 bl[235] br[235] wl[246] vdd gnd cell_6t
Xbit_r247_c235 bl[235] br[235] wl[247] vdd gnd cell_6t
Xbit_r248_c235 bl[235] br[235] wl[248] vdd gnd cell_6t
Xbit_r249_c235 bl[235] br[235] wl[249] vdd gnd cell_6t
Xbit_r250_c235 bl[235] br[235] wl[250] vdd gnd cell_6t
Xbit_r251_c235 bl[235] br[235] wl[251] vdd gnd cell_6t
Xbit_r252_c235 bl[235] br[235] wl[252] vdd gnd cell_6t
Xbit_r253_c235 bl[235] br[235] wl[253] vdd gnd cell_6t
Xbit_r254_c235 bl[235] br[235] wl[254] vdd gnd cell_6t
Xbit_r255_c235 bl[235] br[235] wl[255] vdd gnd cell_6t
Xbit_r0_c236 bl[236] br[236] wl[0] vdd gnd cell_6t
Xbit_r1_c236 bl[236] br[236] wl[1] vdd gnd cell_6t
Xbit_r2_c236 bl[236] br[236] wl[2] vdd gnd cell_6t
Xbit_r3_c236 bl[236] br[236] wl[3] vdd gnd cell_6t
Xbit_r4_c236 bl[236] br[236] wl[4] vdd gnd cell_6t
Xbit_r5_c236 bl[236] br[236] wl[5] vdd gnd cell_6t
Xbit_r6_c236 bl[236] br[236] wl[6] vdd gnd cell_6t
Xbit_r7_c236 bl[236] br[236] wl[7] vdd gnd cell_6t
Xbit_r8_c236 bl[236] br[236] wl[8] vdd gnd cell_6t
Xbit_r9_c236 bl[236] br[236] wl[9] vdd gnd cell_6t
Xbit_r10_c236 bl[236] br[236] wl[10] vdd gnd cell_6t
Xbit_r11_c236 bl[236] br[236] wl[11] vdd gnd cell_6t
Xbit_r12_c236 bl[236] br[236] wl[12] vdd gnd cell_6t
Xbit_r13_c236 bl[236] br[236] wl[13] vdd gnd cell_6t
Xbit_r14_c236 bl[236] br[236] wl[14] vdd gnd cell_6t
Xbit_r15_c236 bl[236] br[236] wl[15] vdd gnd cell_6t
Xbit_r16_c236 bl[236] br[236] wl[16] vdd gnd cell_6t
Xbit_r17_c236 bl[236] br[236] wl[17] vdd gnd cell_6t
Xbit_r18_c236 bl[236] br[236] wl[18] vdd gnd cell_6t
Xbit_r19_c236 bl[236] br[236] wl[19] vdd gnd cell_6t
Xbit_r20_c236 bl[236] br[236] wl[20] vdd gnd cell_6t
Xbit_r21_c236 bl[236] br[236] wl[21] vdd gnd cell_6t
Xbit_r22_c236 bl[236] br[236] wl[22] vdd gnd cell_6t
Xbit_r23_c236 bl[236] br[236] wl[23] vdd gnd cell_6t
Xbit_r24_c236 bl[236] br[236] wl[24] vdd gnd cell_6t
Xbit_r25_c236 bl[236] br[236] wl[25] vdd gnd cell_6t
Xbit_r26_c236 bl[236] br[236] wl[26] vdd gnd cell_6t
Xbit_r27_c236 bl[236] br[236] wl[27] vdd gnd cell_6t
Xbit_r28_c236 bl[236] br[236] wl[28] vdd gnd cell_6t
Xbit_r29_c236 bl[236] br[236] wl[29] vdd gnd cell_6t
Xbit_r30_c236 bl[236] br[236] wl[30] vdd gnd cell_6t
Xbit_r31_c236 bl[236] br[236] wl[31] vdd gnd cell_6t
Xbit_r32_c236 bl[236] br[236] wl[32] vdd gnd cell_6t
Xbit_r33_c236 bl[236] br[236] wl[33] vdd gnd cell_6t
Xbit_r34_c236 bl[236] br[236] wl[34] vdd gnd cell_6t
Xbit_r35_c236 bl[236] br[236] wl[35] vdd gnd cell_6t
Xbit_r36_c236 bl[236] br[236] wl[36] vdd gnd cell_6t
Xbit_r37_c236 bl[236] br[236] wl[37] vdd gnd cell_6t
Xbit_r38_c236 bl[236] br[236] wl[38] vdd gnd cell_6t
Xbit_r39_c236 bl[236] br[236] wl[39] vdd gnd cell_6t
Xbit_r40_c236 bl[236] br[236] wl[40] vdd gnd cell_6t
Xbit_r41_c236 bl[236] br[236] wl[41] vdd gnd cell_6t
Xbit_r42_c236 bl[236] br[236] wl[42] vdd gnd cell_6t
Xbit_r43_c236 bl[236] br[236] wl[43] vdd gnd cell_6t
Xbit_r44_c236 bl[236] br[236] wl[44] vdd gnd cell_6t
Xbit_r45_c236 bl[236] br[236] wl[45] vdd gnd cell_6t
Xbit_r46_c236 bl[236] br[236] wl[46] vdd gnd cell_6t
Xbit_r47_c236 bl[236] br[236] wl[47] vdd gnd cell_6t
Xbit_r48_c236 bl[236] br[236] wl[48] vdd gnd cell_6t
Xbit_r49_c236 bl[236] br[236] wl[49] vdd gnd cell_6t
Xbit_r50_c236 bl[236] br[236] wl[50] vdd gnd cell_6t
Xbit_r51_c236 bl[236] br[236] wl[51] vdd gnd cell_6t
Xbit_r52_c236 bl[236] br[236] wl[52] vdd gnd cell_6t
Xbit_r53_c236 bl[236] br[236] wl[53] vdd gnd cell_6t
Xbit_r54_c236 bl[236] br[236] wl[54] vdd gnd cell_6t
Xbit_r55_c236 bl[236] br[236] wl[55] vdd gnd cell_6t
Xbit_r56_c236 bl[236] br[236] wl[56] vdd gnd cell_6t
Xbit_r57_c236 bl[236] br[236] wl[57] vdd gnd cell_6t
Xbit_r58_c236 bl[236] br[236] wl[58] vdd gnd cell_6t
Xbit_r59_c236 bl[236] br[236] wl[59] vdd gnd cell_6t
Xbit_r60_c236 bl[236] br[236] wl[60] vdd gnd cell_6t
Xbit_r61_c236 bl[236] br[236] wl[61] vdd gnd cell_6t
Xbit_r62_c236 bl[236] br[236] wl[62] vdd gnd cell_6t
Xbit_r63_c236 bl[236] br[236] wl[63] vdd gnd cell_6t
Xbit_r64_c236 bl[236] br[236] wl[64] vdd gnd cell_6t
Xbit_r65_c236 bl[236] br[236] wl[65] vdd gnd cell_6t
Xbit_r66_c236 bl[236] br[236] wl[66] vdd gnd cell_6t
Xbit_r67_c236 bl[236] br[236] wl[67] vdd gnd cell_6t
Xbit_r68_c236 bl[236] br[236] wl[68] vdd gnd cell_6t
Xbit_r69_c236 bl[236] br[236] wl[69] vdd gnd cell_6t
Xbit_r70_c236 bl[236] br[236] wl[70] vdd gnd cell_6t
Xbit_r71_c236 bl[236] br[236] wl[71] vdd gnd cell_6t
Xbit_r72_c236 bl[236] br[236] wl[72] vdd gnd cell_6t
Xbit_r73_c236 bl[236] br[236] wl[73] vdd gnd cell_6t
Xbit_r74_c236 bl[236] br[236] wl[74] vdd gnd cell_6t
Xbit_r75_c236 bl[236] br[236] wl[75] vdd gnd cell_6t
Xbit_r76_c236 bl[236] br[236] wl[76] vdd gnd cell_6t
Xbit_r77_c236 bl[236] br[236] wl[77] vdd gnd cell_6t
Xbit_r78_c236 bl[236] br[236] wl[78] vdd gnd cell_6t
Xbit_r79_c236 bl[236] br[236] wl[79] vdd gnd cell_6t
Xbit_r80_c236 bl[236] br[236] wl[80] vdd gnd cell_6t
Xbit_r81_c236 bl[236] br[236] wl[81] vdd gnd cell_6t
Xbit_r82_c236 bl[236] br[236] wl[82] vdd gnd cell_6t
Xbit_r83_c236 bl[236] br[236] wl[83] vdd gnd cell_6t
Xbit_r84_c236 bl[236] br[236] wl[84] vdd gnd cell_6t
Xbit_r85_c236 bl[236] br[236] wl[85] vdd gnd cell_6t
Xbit_r86_c236 bl[236] br[236] wl[86] vdd gnd cell_6t
Xbit_r87_c236 bl[236] br[236] wl[87] vdd gnd cell_6t
Xbit_r88_c236 bl[236] br[236] wl[88] vdd gnd cell_6t
Xbit_r89_c236 bl[236] br[236] wl[89] vdd gnd cell_6t
Xbit_r90_c236 bl[236] br[236] wl[90] vdd gnd cell_6t
Xbit_r91_c236 bl[236] br[236] wl[91] vdd gnd cell_6t
Xbit_r92_c236 bl[236] br[236] wl[92] vdd gnd cell_6t
Xbit_r93_c236 bl[236] br[236] wl[93] vdd gnd cell_6t
Xbit_r94_c236 bl[236] br[236] wl[94] vdd gnd cell_6t
Xbit_r95_c236 bl[236] br[236] wl[95] vdd gnd cell_6t
Xbit_r96_c236 bl[236] br[236] wl[96] vdd gnd cell_6t
Xbit_r97_c236 bl[236] br[236] wl[97] vdd gnd cell_6t
Xbit_r98_c236 bl[236] br[236] wl[98] vdd gnd cell_6t
Xbit_r99_c236 bl[236] br[236] wl[99] vdd gnd cell_6t
Xbit_r100_c236 bl[236] br[236] wl[100] vdd gnd cell_6t
Xbit_r101_c236 bl[236] br[236] wl[101] vdd gnd cell_6t
Xbit_r102_c236 bl[236] br[236] wl[102] vdd gnd cell_6t
Xbit_r103_c236 bl[236] br[236] wl[103] vdd gnd cell_6t
Xbit_r104_c236 bl[236] br[236] wl[104] vdd gnd cell_6t
Xbit_r105_c236 bl[236] br[236] wl[105] vdd gnd cell_6t
Xbit_r106_c236 bl[236] br[236] wl[106] vdd gnd cell_6t
Xbit_r107_c236 bl[236] br[236] wl[107] vdd gnd cell_6t
Xbit_r108_c236 bl[236] br[236] wl[108] vdd gnd cell_6t
Xbit_r109_c236 bl[236] br[236] wl[109] vdd gnd cell_6t
Xbit_r110_c236 bl[236] br[236] wl[110] vdd gnd cell_6t
Xbit_r111_c236 bl[236] br[236] wl[111] vdd gnd cell_6t
Xbit_r112_c236 bl[236] br[236] wl[112] vdd gnd cell_6t
Xbit_r113_c236 bl[236] br[236] wl[113] vdd gnd cell_6t
Xbit_r114_c236 bl[236] br[236] wl[114] vdd gnd cell_6t
Xbit_r115_c236 bl[236] br[236] wl[115] vdd gnd cell_6t
Xbit_r116_c236 bl[236] br[236] wl[116] vdd gnd cell_6t
Xbit_r117_c236 bl[236] br[236] wl[117] vdd gnd cell_6t
Xbit_r118_c236 bl[236] br[236] wl[118] vdd gnd cell_6t
Xbit_r119_c236 bl[236] br[236] wl[119] vdd gnd cell_6t
Xbit_r120_c236 bl[236] br[236] wl[120] vdd gnd cell_6t
Xbit_r121_c236 bl[236] br[236] wl[121] vdd gnd cell_6t
Xbit_r122_c236 bl[236] br[236] wl[122] vdd gnd cell_6t
Xbit_r123_c236 bl[236] br[236] wl[123] vdd gnd cell_6t
Xbit_r124_c236 bl[236] br[236] wl[124] vdd gnd cell_6t
Xbit_r125_c236 bl[236] br[236] wl[125] vdd gnd cell_6t
Xbit_r126_c236 bl[236] br[236] wl[126] vdd gnd cell_6t
Xbit_r127_c236 bl[236] br[236] wl[127] vdd gnd cell_6t
Xbit_r128_c236 bl[236] br[236] wl[128] vdd gnd cell_6t
Xbit_r129_c236 bl[236] br[236] wl[129] vdd gnd cell_6t
Xbit_r130_c236 bl[236] br[236] wl[130] vdd gnd cell_6t
Xbit_r131_c236 bl[236] br[236] wl[131] vdd gnd cell_6t
Xbit_r132_c236 bl[236] br[236] wl[132] vdd gnd cell_6t
Xbit_r133_c236 bl[236] br[236] wl[133] vdd gnd cell_6t
Xbit_r134_c236 bl[236] br[236] wl[134] vdd gnd cell_6t
Xbit_r135_c236 bl[236] br[236] wl[135] vdd gnd cell_6t
Xbit_r136_c236 bl[236] br[236] wl[136] vdd gnd cell_6t
Xbit_r137_c236 bl[236] br[236] wl[137] vdd gnd cell_6t
Xbit_r138_c236 bl[236] br[236] wl[138] vdd gnd cell_6t
Xbit_r139_c236 bl[236] br[236] wl[139] vdd gnd cell_6t
Xbit_r140_c236 bl[236] br[236] wl[140] vdd gnd cell_6t
Xbit_r141_c236 bl[236] br[236] wl[141] vdd gnd cell_6t
Xbit_r142_c236 bl[236] br[236] wl[142] vdd gnd cell_6t
Xbit_r143_c236 bl[236] br[236] wl[143] vdd gnd cell_6t
Xbit_r144_c236 bl[236] br[236] wl[144] vdd gnd cell_6t
Xbit_r145_c236 bl[236] br[236] wl[145] vdd gnd cell_6t
Xbit_r146_c236 bl[236] br[236] wl[146] vdd gnd cell_6t
Xbit_r147_c236 bl[236] br[236] wl[147] vdd gnd cell_6t
Xbit_r148_c236 bl[236] br[236] wl[148] vdd gnd cell_6t
Xbit_r149_c236 bl[236] br[236] wl[149] vdd gnd cell_6t
Xbit_r150_c236 bl[236] br[236] wl[150] vdd gnd cell_6t
Xbit_r151_c236 bl[236] br[236] wl[151] vdd gnd cell_6t
Xbit_r152_c236 bl[236] br[236] wl[152] vdd gnd cell_6t
Xbit_r153_c236 bl[236] br[236] wl[153] vdd gnd cell_6t
Xbit_r154_c236 bl[236] br[236] wl[154] vdd gnd cell_6t
Xbit_r155_c236 bl[236] br[236] wl[155] vdd gnd cell_6t
Xbit_r156_c236 bl[236] br[236] wl[156] vdd gnd cell_6t
Xbit_r157_c236 bl[236] br[236] wl[157] vdd gnd cell_6t
Xbit_r158_c236 bl[236] br[236] wl[158] vdd gnd cell_6t
Xbit_r159_c236 bl[236] br[236] wl[159] vdd gnd cell_6t
Xbit_r160_c236 bl[236] br[236] wl[160] vdd gnd cell_6t
Xbit_r161_c236 bl[236] br[236] wl[161] vdd gnd cell_6t
Xbit_r162_c236 bl[236] br[236] wl[162] vdd gnd cell_6t
Xbit_r163_c236 bl[236] br[236] wl[163] vdd gnd cell_6t
Xbit_r164_c236 bl[236] br[236] wl[164] vdd gnd cell_6t
Xbit_r165_c236 bl[236] br[236] wl[165] vdd gnd cell_6t
Xbit_r166_c236 bl[236] br[236] wl[166] vdd gnd cell_6t
Xbit_r167_c236 bl[236] br[236] wl[167] vdd gnd cell_6t
Xbit_r168_c236 bl[236] br[236] wl[168] vdd gnd cell_6t
Xbit_r169_c236 bl[236] br[236] wl[169] vdd gnd cell_6t
Xbit_r170_c236 bl[236] br[236] wl[170] vdd gnd cell_6t
Xbit_r171_c236 bl[236] br[236] wl[171] vdd gnd cell_6t
Xbit_r172_c236 bl[236] br[236] wl[172] vdd gnd cell_6t
Xbit_r173_c236 bl[236] br[236] wl[173] vdd gnd cell_6t
Xbit_r174_c236 bl[236] br[236] wl[174] vdd gnd cell_6t
Xbit_r175_c236 bl[236] br[236] wl[175] vdd gnd cell_6t
Xbit_r176_c236 bl[236] br[236] wl[176] vdd gnd cell_6t
Xbit_r177_c236 bl[236] br[236] wl[177] vdd gnd cell_6t
Xbit_r178_c236 bl[236] br[236] wl[178] vdd gnd cell_6t
Xbit_r179_c236 bl[236] br[236] wl[179] vdd gnd cell_6t
Xbit_r180_c236 bl[236] br[236] wl[180] vdd gnd cell_6t
Xbit_r181_c236 bl[236] br[236] wl[181] vdd gnd cell_6t
Xbit_r182_c236 bl[236] br[236] wl[182] vdd gnd cell_6t
Xbit_r183_c236 bl[236] br[236] wl[183] vdd gnd cell_6t
Xbit_r184_c236 bl[236] br[236] wl[184] vdd gnd cell_6t
Xbit_r185_c236 bl[236] br[236] wl[185] vdd gnd cell_6t
Xbit_r186_c236 bl[236] br[236] wl[186] vdd gnd cell_6t
Xbit_r187_c236 bl[236] br[236] wl[187] vdd gnd cell_6t
Xbit_r188_c236 bl[236] br[236] wl[188] vdd gnd cell_6t
Xbit_r189_c236 bl[236] br[236] wl[189] vdd gnd cell_6t
Xbit_r190_c236 bl[236] br[236] wl[190] vdd gnd cell_6t
Xbit_r191_c236 bl[236] br[236] wl[191] vdd gnd cell_6t
Xbit_r192_c236 bl[236] br[236] wl[192] vdd gnd cell_6t
Xbit_r193_c236 bl[236] br[236] wl[193] vdd gnd cell_6t
Xbit_r194_c236 bl[236] br[236] wl[194] vdd gnd cell_6t
Xbit_r195_c236 bl[236] br[236] wl[195] vdd gnd cell_6t
Xbit_r196_c236 bl[236] br[236] wl[196] vdd gnd cell_6t
Xbit_r197_c236 bl[236] br[236] wl[197] vdd gnd cell_6t
Xbit_r198_c236 bl[236] br[236] wl[198] vdd gnd cell_6t
Xbit_r199_c236 bl[236] br[236] wl[199] vdd gnd cell_6t
Xbit_r200_c236 bl[236] br[236] wl[200] vdd gnd cell_6t
Xbit_r201_c236 bl[236] br[236] wl[201] vdd gnd cell_6t
Xbit_r202_c236 bl[236] br[236] wl[202] vdd gnd cell_6t
Xbit_r203_c236 bl[236] br[236] wl[203] vdd gnd cell_6t
Xbit_r204_c236 bl[236] br[236] wl[204] vdd gnd cell_6t
Xbit_r205_c236 bl[236] br[236] wl[205] vdd gnd cell_6t
Xbit_r206_c236 bl[236] br[236] wl[206] vdd gnd cell_6t
Xbit_r207_c236 bl[236] br[236] wl[207] vdd gnd cell_6t
Xbit_r208_c236 bl[236] br[236] wl[208] vdd gnd cell_6t
Xbit_r209_c236 bl[236] br[236] wl[209] vdd gnd cell_6t
Xbit_r210_c236 bl[236] br[236] wl[210] vdd gnd cell_6t
Xbit_r211_c236 bl[236] br[236] wl[211] vdd gnd cell_6t
Xbit_r212_c236 bl[236] br[236] wl[212] vdd gnd cell_6t
Xbit_r213_c236 bl[236] br[236] wl[213] vdd gnd cell_6t
Xbit_r214_c236 bl[236] br[236] wl[214] vdd gnd cell_6t
Xbit_r215_c236 bl[236] br[236] wl[215] vdd gnd cell_6t
Xbit_r216_c236 bl[236] br[236] wl[216] vdd gnd cell_6t
Xbit_r217_c236 bl[236] br[236] wl[217] vdd gnd cell_6t
Xbit_r218_c236 bl[236] br[236] wl[218] vdd gnd cell_6t
Xbit_r219_c236 bl[236] br[236] wl[219] vdd gnd cell_6t
Xbit_r220_c236 bl[236] br[236] wl[220] vdd gnd cell_6t
Xbit_r221_c236 bl[236] br[236] wl[221] vdd gnd cell_6t
Xbit_r222_c236 bl[236] br[236] wl[222] vdd gnd cell_6t
Xbit_r223_c236 bl[236] br[236] wl[223] vdd gnd cell_6t
Xbit_r224_c236 bl[236] br[236] wl[224] vdd gnd cell_6t
Xbit_r225_c236 bl[236] br[236] wl[225] vdd gnd cell_6t
Xbit_r226_c236 bl[236] br[236] wl[226] vdd gnd cell_6t
Xbit_r227_c236 bl[236] br[236] wl[227] vdd gnd cell_6t
Xbit_r228_c236 bl[236] br[236] wl[228] vdd gnd cell_6t
Xbit_r229_c236 bl[236] br[236] wl[229] vdd gnd cell_6t
Xbit_r230_c236 bl[236] br[236] wl[230] vdd gnd cell_6t
Xbit_r231_c236 bl[236] br[236] wl[231] vdd gnd cell_6t
Xbit_r232_c236 bl[236] br[236] wl[232] vdd gnd cell_6t
Xbit_r233_c236 bl[236] br[236] wl[233] vdd gnd cell_6t
Xbit_r234_c236 bl[236] br[236] wl[234] vdd gnd cell_6t
Xbit_r235_c236 bl[236] br[236] wl[235] vdd gnd cell_6t
Xbit_r236_c236 bl[236] br[236] wl[236] vdd gnd cell_6t
Xbit_r237_c236 bl[236] br[236] wl[237] vdd gnd cell_6t
Xbit_r238_c236 bl[236] br[236] wl[238] vdd gnd cell_6t
Xbit_r239_c236 bl[236] br[236] wl[239] vdd gnd cell_6t
Xbit_r240_c236 bl[236] br[236] wl[240] vdd gnd cell_6t
Xbit_r241_c236 bl[236] br[236] wl[241] vdd gnd cell_6t
Xbit_r242_c236 bl[236] br[236] wl[242] vdd gnd cell_6t
Xbit_r243_c236 bl[236] br[236] wl[243] vdd gnd cell_6t
Xbit_r244_c236 bl[236] br[236] wl[244] vdd gnd cell_6t
Xbit_r245_c236 bl[236] br[236] wl[245] vdd gnd cell_6t
Xbit_r246_c236 bl[236] br[236] wl[246] vdd gnd cell_6t
Xbit_r247_c236 bl[236] br[236] wl[247] vdd gnd cell_6t
Xbit_r248_c236 bl[236] br[236] wl[248] vdd gnd cell_6t
Xbit_r249_c236 bl[236] br[236] wl[249] vdd gnd cell_6t
Xbit_r250_c236 bl[236] br[236] wl[250] vdd gnd cell_6t
Xbit_r251_c236 bl[236] br[236] wl[251] vdd gnd cell_6t
Xbit_r252_c236 bl[236] br[236] wl[252] vdd gnd cell_6t
Xbit_r253_c236 bl[236] br[236] wl[253] vdd gnd cell_6t
Xbit_r254_c236 bl[236] br[236] wl[254] vdd gnd cell_6t
Xbit_r255_c236 bl[236] br[236] wl[255] vdd gnd cell_6t
Xbit_r0_c237 bl[237] br[237] wl[0] vdd gnd cell_6t
Xbit_r1_c237 bl[237] br[237] wl[1] vdd gnd cell_6t
Xbit_r2_c237 bl[237] br[237] wl[2] vdd gnd cell_6t
Xbit_r3_c237 bl[237] br[237] wl[3] vdd gnd cell_6t
Xbit_r4_c237 bl[237] br[237] wl[4] vdd gnd cell_6t
Xbit_r5_c237 bl[237] br[237] wl[5] vdd gnd cell_6t
Xbit_r6_c237 bl[237] br[237] wl[6] vdd gnd cell_6t
Xbit_r7_c237 bl[237] br[237] wl[7] vdd gnd cell_6t
Xbit_r8_c237 bl[237] br[237] wl[8] vdd gnd cell_6t
Xbit_r9_c237 bl[237] br[237] wl[9] vdd gnd cell_6t
Xbit_r10_c237 bl[237] br[237] wl[10] vdd gnd cell_6t
Xbit_r11_c237 bl[237] br[237] wl[11] vdd gnd cell_6t
Xbit_r12_c237 bl[237] br[237] wl[12] vdd gnd cell_6t
Xbit_r13_c237 bl[237] br[237] wl[13] vdd gnd cell_6t
Xbit_r14_c237 bl[237] br[237] wl[14] vdd gnd cell_6t
Xbit_r15_c237 bl[237] br[237] wl[15] vdd gnd cell_6t
Xbit_r16_c237 bl[237] br[237] wl[16] vdd gnd cell_6t
Xbit_r17_c237 bl[237] br[237] wl[17] vdd gnd cell_6t
Xbit_r18_c237 bl[237] br[237] wl[18] vdd gnd cell_6t
Xbit_r19_c237 bl[237] br[237] wl[19] vdd gnd cell_6t
Xbit_r20_c237 bl[237] br[237] wl[20] vdd gnd cell_6t
Xbit_r21_c237 bl[237] br[237] wl[21] vdd gnd cell_6t
Xbit_r22_c237 bl[237] br[237] wl[22] vdd gnd cell_6t
Xbit_r23_c237 bl[237] br[237] wl[23] vdd gnd cell_6t
Xbit_r24_c237 bl[237] br[237] wl[24] vdd gnd cell_6t
Xbit_r25_c237 bl[237] br[237] wl[25] vdd gnd cell_6t
Xbit_r26_c237 bl[237] br[237] wl[26] vdd gnd cell_6t
Xbit_r27_c237 bl[237] br[237] wl[27] vdd gnd cell_6t
Xbit_r28_c237 bl[237] br[237] wl[28] vdd gnd cell_6t
Xbit_r29_c237 bl[237] br[237] wl[29] vdd gnd cell_6t
Xbit_r30_c237 bl[237] br[237] wl[30] vdd gnd cell_6t
Xbit_r31_c237 bl[237] br[237] wl[31] vdd gnd cell_6t
Xbit_r32_c237 bl[237] br[237] wl[32] vdd gnd cell_6t
Xbit_r33_c237 bl[237] br[237] wl[33] vdd gnd cell_6t
Xbit_r34_c237 bl[237] br[237] wl[34] vdd gnd cell_6t
Xbit_r35_c237 bl[237] br[237] wl[35] vdd gnd cell_6t
Xbit_r36_c237 bl[237] br[237] wl[36] vdd gnd cell_6t
Xbit_r37_c237 bl[237] br[237] wl[37] vdd gnd cell_6t
Xbit_r38_c237 bl[237] br[237] wl[38] vdd gnd cell_6t
Xbit_r39_c237 bl[237] br[237] wl[39] vdd gnd cell_6t
Xbit_r40_c237 bl[237] br[237] wl[40] vdd gnd cell_6t
Xbit_r41_c237 bl[237] br[237] wl[41] vdd gnd cell_6t
Xbit_r42_c237 bl[237] br[237] wl[42] vdd gnd cell_6t
Xbit_r43_c237 bl[237] br[237] wl[43] vdd gnd cell_6t
Xbit_r44_c237 bl[237] br[237] wl[44] vdd gnd cell_6t
Xbit_r45_c237 bl[237] br[237] wl[45] vdd gnd cell_6t
Xbit_r46_c237 bl[237] br[237] wl[46] vdd gnd cell_6t
Xbit_r47_c237 bl[237] br[237] wl[47] vdd gnd cell_6t
Xbit_r48_c237 bl[237] br[237] wl[48] vdd gnd cell_6t
Xbit_r49_c237 bl[237] br[237] wl[49] vdd gnd cell_6t
Xbit_r50_c237 bl[237] br[237] wl[50] vdd gnd cell_6t
Xbit_r51_c237 bl[237] br[237] wl[51] vdd gnd cell_6t
Xbit_r52_c237 bl[237] br[237] wl[52] vdd gnd cell_6t
Xbit_r53_c237 bl[237] br[237] wl[53] vdd gnd cell_6t
Xbit_r54_c237 bl[237] br[237] wl[54] vdd gnd cell_6t
Xbit_r55_c237 bl[237] br[237] wl[55] vdd gnd cell_6t
Xbit_r56_c237 bl[237] br[237] wl[56] vdd gnd cell_6t
Xbit_r57_c237 bl[237] br[237] wl[57] vdd gnd cell_6t
Xbit_r58_c237 bl[237] br[237] wl[58] vdd gnd cell_6t
Xbit_r59_c237 bl[237] br[237] wl[59] vdd gnd cell_6t
Xbit_r60_c237 bl[237] br[237] wl[60] vdd gnd cell_6t
Xbit_r61_c237 bl[237] br[237] wl[61] vdd gnd cell_6t
Xbit_r62_c237 bl[237] br[237] wl[62] vdd gnd cell_6t
Xbit_r63_c237 bl[237] br[237] wl[63] vdd gnd cell_6t
Xbit_r64_c237 bl[237] br[237] wl[64] vdd gnd cell_6t
Xbit_r65_c237 bl[237] br[237] wl[65] vdd gnd cell_6t
Xbit_r66_c237 bl[237] br[237] wl[66] vdd gnd cell_6t
Xbit_r67_c237 bl[237] br[237] wl[67] vdd gnd cell_6t
Xbit_r68_c237 bl[237] br[237] wl[68] vdd gnd cell_6t
Xbit_r69_c237 bl[237] br[237] wl[69] vdd gnd cell_6t
Xbit_r70_c237 bl[237] br[237] wl[70] vdd gnd cell_6t
Xbit_r71_c237 bl[237] br[237] wl[71] vdd gnd cell_6t
Xbit_r72_c237 bl[237] br[237] wl[72] vdd gnd cell_6t
Xbit_r73_c237 bl[237] br[237] wl[73] vdd gnd cell_6t
Xbit_r74_c237 bl[237] br[237] wl[74] vdd gnd cell_6t
Xbit_r75_c237 bl[237] br[237] wl[75] vdd gnd cell_6t
Xbit_r76_c237 bl[237] br[237] wl[76] vdd gnd cell_6t
Xbit_r77_c237 bl[237] br[237] wl[77] vdd gnd cell_6t
Xbit_r78_c237 bl[237] br[237] wl[78] vdd gnd cell_6t
Xbit_r79_c237 bl[237] br[237] wl[79] vdd gnd cell_6t
Xbit_r80_c237 bl[237] br[237] wl[80] vdd gnd cell_6t
Xbit_r81_c237 bl[237] br[237] wl[81] vdd gnd cell_6t
Xbit_r82_c237 bl[237] br[237] wl[82] vdd gnd cell_6t
Xbit_r83_c237 bl[237] br[237] wl[83] vdd gnd cell_6t
Xbit_r84_c237 bl[237] br[237] wl[84] vdd gnd cell_6t
Xbit_r85_c237 bl[237] br[237] wl[85] vdd gnd cell_6t
Xbit_r86_c237 bl[237] br[237] wl[86] vdd gnd cell_6t
Xbit_r87_c237 bl[237] br[237] wl[87] vdd gnd cell_6t
Xbit_r88_c237 bl[237] br[237] wl[88] vdd gnd cell_6t
Xbit_r89_c237 bl[237] br[237] wl[89] vdd gnd cell_6t
Xbit_r90_c237 bl[237] br[237] wl[90] vdd gnd cell_6t
Xbit_r91_c237 bl[237] br[237] wl[91] vdd gnd cell_6t
Xbit_r92_c237 bl[237] br[237] wl[92] vdd gnd cell_6t
Xbit_r93_c237 bl[237] br[237] wl[93] vdd gnd cell_6t
Xbit_r94_c237 bl[237] br[237] wl[94] vdd gnd cell_6t
Xbit_r95_c237 bl[237] br[237] wl[95] vdd gnd cell_6t
Xbit_r96_c237 bl[237] br[237] wl[96] vdd gnd cell_6t
Xbit_r97_c237 bl[237] br[237] wl[97] vdd gnd cell_6t
Xbit_r98_c237 bl[237] br[237] wl[98] vdd gnd cell_6t
Xbit_r99_c237 bl[237] br[237] wl[99] vdd gnd cell_6t
Xbit_r100_c237 bl[237] br[237] wl[100] vdd gnd cell_6t
Xbit_r101_c237 bl[237] br[237] wl[101] vdd gnd cell_6t
Xbit_r102_c237 bl[237] br[237] wl[102] vdd gnd cell_6t
Xbit_r103_c237 bl[237] br[237] wl[103] vdd gnd cell_6t
Xbit_r104_c237 bl[237] br[237] wl[104] vdd gnd cell_6t
Xbit_r105_c237 bl[237] br[237] wl[105] vdd gnd cell_6t
Xbit_r106_c237 bl[237] br[237] wl[106] vdd gnd cell_6t
Xbit_r107_c237 bl[237] br[237] wl[107] vdd gnd cell_6t
Xbit_r108_c237 bl[237] br[237] wl[108] vdd gnd cell_6t
Xbit_r109_c237 bl[237] br[237] wl[109] vdd gnd cell_6t
Xbit_r110_c237 bl[237] br[237] wl[110] vdd gnd cell_6t
Xbit_r111_c237 bl[237] br[237] wl[111] vdd gnd cell_6t
Xbit_r112_c237 bl[237] br[237] wl[112] vdd gnd cell_6t
Xbit_r113_c237 bl[237] br[237] wl[113] vdd gnd cell_6t
Xbit_r114_c237 bl[237] br[237] wl[114] vdd gnd cell_6t
Xbit_r115_c237 bl[237] br[237] wl[115] vdd gnd cell_6t
Xbit_r116_c237 bl[237] br[237] wl[116] vdd gnd cell_6t
Xbit_r117_c237 bl[237] br[237] wl[117] vdd gnd cell_6t
Xbit_r118_c237 bl[237] br[237] wl[118] vdd gnd cell_6t
Xbit_r119_c237 bl[237] br[237] wl[119] vdd gnd cell_6t
Xbit_r120_c237 bl[237] br[237] wl[120] vdd gnd cell_6t
Xbit_r121_c237 bl[237] br[237] wl[121] vdd gnd cell_6t
Xbit_r122_c237 bl[237] br[237] wl[122] vdd gnd cell_6t
Xbit_r123_c237 bl[237] br[237] wl[123] vdd gnd cell_6t
Xbit_r124_c237 bl[237] br[237] wl[124] vdd gnd cell_6t
Xbit_r125_c237 bl[237] br[237] wl[125] vdd gnd cell_6t
Xbit_r126_c237 bl[237] br[237] wl[126] vdd gnd cell_6t
Xbit_r127_c237 bl[237] br[237] wl[127] vdd gnd cell_6t
Xbit_r128_c237 bl[237] br[237] wl[128] vdd gnd cell_6t
Xbit_r129_c237 bl[237] br[237] wl[129] vdd gnd cell_6t
Xbit_r130_c237 bl[237] br[237] wl[130] vdd gnd cell_6t
Xbit_r131_c237 bl[237] br[237] wl[131] vdd gnd cell_6t
Xbit_r132_c237 bl[237] br[237] wl[132] vdd gnd cell_6t
Xbit_r133_c237 bl[237] br[237] wl[133] vdd gnd cell_6t
Xbit_r134_c237 bl[237] br[237] wl[134] vdd gnd cell_6t
Xbit_r135_c237 bl[237] br[237] wl[135] vdd gnd cell_6t
Xbit_r136_c237 bl[237] br[237] wl[136] vdd gnd cell_6t
Xbit_r137_c237 bl[237] br[237] wl[137] vdd gnd cell_6t
Xbit_r138_c237 bl[237] br[237] wl[138] vdd gnd cell_6t
Xbit_r139_c237 bl[237] br[237] wl[139] vdd gnd cell_6t
Xbit_r140_c237 bl[237] br[237] wl[140] vdd gnd cell_6t
Xbit_r141_c237 bl[237] br[237] wl[141] vdd gnd cell_6t
Xbit_r142_c237 bl[237] br[237] wl[142] vdd gnd cell_6t
Xbit_r143_c237 bl[237] br[237] wl[143] vdd gnd cell_6t
Xbit_r144_c237 bl[237] br[237] wl[144] vdd gnd cell_6t
Xbit_r145_c237 bl[237] br[237] wl[145] vdd gnd cell_6t
Xbit_r146_c237 bl[237] br[237] wl[146] vdd gnd cell_6t
Xbit_r147_c237 bl[237] br[237] wl[147] vdd gnd cell_6t
Xbit_r148_c237 bl[237] br[237] wl[148] vdd gnd cell_6t
Xbit_r149_c237 bl[237] br[237] wl[149] vdd gnd cell_6t
Xbit_r150_c237 bl[237] br[237] wl[150] vdd gnd cell_6t
Xbit_r151_c237 bl[237] br[237] wl[151] vdd gnd cell_6t
Xbit_r152_c237 bl[237] br[237] wl[152] vdd gnd cell_6t
Xbit_r153_c237 bl[237] br[237] wl[153] vdd gnd cell_6t
Xbit_r154_c237 bl[237] br[237] wl[154] vdd gnd cell_6t
Xbit_r155_c237 bl[237] br[237] wl[155] vdd gnd cell_6t
Xbit_r156_c237 bl[237] br[237] wl[156] vdd gnd cell_6t
Xbit_r157_c237 bl[237] br[237] wl[157] vdd gnd cell_6t
Xbit_r158_c237 bl[237] br[237] wl[158] vdd gnd cell_6t
Xbit_r159_c237 bl[237] br[237] wl[159] vdd gnd cell_6t
Xbit_r160_c237 bl[237] br[237] wl[160] vdd gnd cell_6t
Xbit_r161_c237 bl[237] br[237] wl[161] vdd gnd cell_6t
Xbit_r162_c237 bl[237] br[237] wl[162] vdd gnd cell_6t
Xbit_r163_c237 bl[237] br[237] wl[163] vdd gnd cell_6t
Xbit_r164_c237 bl[237] br[237] wl[164] vdd gnd cell_6t
Xbit_r165_c237 bl[237] br[237] wl[165] vdd gnd cell_6t
Xbit_r166_c237 bl[237] br[237] wl[166] vdd gnd cell_6t
Xbit_r167_c237 bl[237] br[237] wl[167] vdd gnd cell_6t
Xbit_r168_c237 bl[237] br[237] wl[168] vdd gnd cell_6t
Xbit_r169_c237 bl[237] br[237] wl[169] vdd gnd cell_6t
Xbit_r170_c237 bl[237] br[237] wl[170] vdd gnd cell_6t
Xbit_r171_c237 bl[237] br[237] wl[171] vdd gnd cell_6t
Xbit_r172_c237 bl[237] br[237] wl[172] vdd gnd cell_6t
Xbit_r173_c237 bl[237] br[237] wl[173] vdd gnd cell_6t
Xbit_r174_c237 bl[237] br[237] wl[174] vdd gnd cell_6t
Xbit_r175_c237 bl[237] br[237] wl[175] vdd gnd cell_6t
Xbit_r176_c237 bl[237] br[237] wl[176] vdd gnd cell_6t
Xbit_r177_c237 bl[237] br[237] wl[177] vdd gnd cell_6t
Xbit_r178_c237 bl[237] br[237] wl[178] vdd gnd cell_6t
Xbit_r179_c237 bl[237] br[237] wl[179] vdd gnd cell_6t
Xbit_r180_c237 bl[237] br[237] wl[180] vdd gnd cell_6t
Xbit_r181_c237 bl[237] br[237] wl[181] vdd gnd cell_6t
Xbit_r182_c237 bl[237] br[237] wl[182] vdd gnd cell_6t
Xbit_r183_c237 bl[237] br[237] wl[183] vdd gnd cell_6t
Xbit_r184_c237 bl[237] br[237] wl[184] vdd gnd cell_6t
Xbit_r185_c237 bl[237] br[237] wl[185] vdd gnd cell_6t
Xbit_r186_c237 bl[237] br[237] wl[186] vdd gnd cell_6t
Xbit_r187_c237 bl[237] br[237] wl[187] vdd gnd cell_6t
Xbit_r188_c237 bl[237] br[237] wl[188] vdd gnd cell_6t
Xbit_r189_c237 bl[237] br[237] wl[189] vdd gnd cell_6t
Xbit_r190_c237 bl[237] br[237] wl[190] vdd gnd cell_6t
Xbit_r191_c237 bl[237] br[237] wl[191] vdd gnd cell_6t
Xbit_r192_c237 bl[237] br[237] wl[192] vdd gnd cell_6t
Xbit_r193_c237 bl[237] br[237] wl[193] vdd gnd cell_6t
Xbit_r194_c237 bl[237] br[237] wl[194] vdd gnd cell_6t
Xbit_r195_c237 bl[237] br[237] wl[195] vdd gnd cell_6t
Xbit_r196_c237 bl[237] br[237] wl[196] vdd gnd cell_6t
Xbit_r197_c237 bl[237] br[237] wl[197] vdd gnd cell_6t
Xbit_r198_c237 bl[237] br[237] wl[198] vdd gnd cell_6t
Xbit_r199_c237 bl[237] br[237] wl[199] vdd gnd cell_6t
Xbit_r200_c237 bl[237] br[237] wl[200] vdd gnd cell_6t
Xbit_r201_c237 bl[237] br[237] wl[201] vdd gnd cell_6t
Xbit_r202_c237 bl[237] br[237] wl[202] vdd gnd cell_6t
Xbit_r203_c237 bl[237] br[237] wl[203] vdd gnd cell_6t
Xbit_r204_c237 bl[237] br[237] wl[204] vdd gnd cell_6t
Xbit_r205_c237 bl[237] br[237] wl[205] vdd gnd cell_6t
Xbit_r206_c237 bl[237] br[237] wl[206] vdd gnd cell_6t
Xbit_r207_c237 bl[237] br[237] wl[207] vdd gnd cell_6t
Xbit_r208_c237 bl[237] br[237] wl[208] vdd gnd cell_6t
Xbit_r209_c237 bl[237] br[237] wl[209] vdd gnd cell_6t
Xbit_r210_c237 bl[237] br[237] wl[210] vdd gnd cell_6t
Xbit_r211_c237 bl[237] br[237] wl[211] vdd gnd cell_6t
Xbit_r212_c237 bl[237] br[237] wl[212] vdd gnd cell_6t
Xbit_r213_c237 bl[237] br[237] wl[213] vdd gnd cell_6t
Xbit_r214_c237 bl[237] br[237] wl[214] vdd gnd cell_6t
Xbit_r215_c237 bl[237] br[237] wl[215] vdd gnd cell_6t
Xbit_r216_c237 bl[237] br[237] wl[216] vdd gnd cell_6t
Xbit_r217_c237 bl[237] br[237] wl[217] vdd gnd cell_6t
Xbit_r218_c237 bl[237] br[237] wl[218] vdd gnd cell_6t
Xbit_r219_c237 bl[237] br[237] wl[219] vdd gnd cell_6t
Xbit_r220_c237 bl[237] br[237] wl[220] vdd gnd cell_6t
Xbit_r221_c237 bl[237] br[237] wl[221] vdd gnd cell_6t
Xbit_r222_c237 bl[237] br[237] wl[222] vdd gnd cell_6t
Xbit_r223_c237 bl[237] br[237] wl[223] vdd gnd cell_6t
Xbit_r224_c237 bl[237] br[237] wl[224] vdd gnd cell_6t
Xbit_r225_c237 bl[237] br[237] wl[225] vdd gnd cell_6t
Xbit_r226_c237 bl[237] br[237] wl[226] vdd gnd cell_6t
Xbit_r227_c237 bl[237] br[237] wl[227] vdd gnd cell_6t
Xbit_r228_c237 bl[237] br[237] wl[228] vdd gnd cell_6t
Xbit_r229_c237 bl[237] br[237] wl[229] vdd gnd cell_6t
Xbit_r230_c237 bl[237] br[237] wl[230] vdd gnd cell_6t
Xbit_r231_c237 bl[237] br[237] wl[231] vdd gnd cell_6t
Xbit_r232_c237 bl[237] br[237] wl[232] vdd gnd cell_6t
Xbit_r233_c237 bl[237] br[237] wl[233] vdd gnd cell_6t
Xbit_r234_c237 bl[237] br[237] wl[234] vdd gnd cell_6t
Xbit_r235_c237 bl[237] br[237] wl[235] vdd gnd cell_6t
Xbit_r236_c237 bl[237] br[237] wl[236] vdd gnd cell_6t
Xbit_r237_c237 bl[237] br[237] wl[237] vdd gnd cell_6t
Xbit_r238_c237 bl[237] br[237] wl[238] vdd gnd cell_6t
Xbit_r239_c237 bl[237] br[237] wl[239] vdd gnd cell_6t
Xbit_r240_c237 bl[237] br[237] wl[240] vdd gnd cell_6t
Xbit_r241_c237 bl[237] br[237] wl[241] vdd gnd cell_6t
Xbit_r242_c237 bl[237] br[237] wl[242] vdd gnd cell_6t
Xbit_r243_c237 bl[237] br[237] wl[243] vdd gnd cell_6t
Xbit_r244_c237 bl[237] br[237] wl[244] vdd gnd cell_6t
Xbit_r245_c237 bl[237] br[237] wl[245] vdd gnd cell_6t
Xbit_r246_c237 bl[237] br[237] wl[246] vdd gnd cell_6t
Xbit_r247_c237 bl[237] br[237] wl[247] vdd gnd cell_6t
Xbit_r248_c237 bl[237] br[237] wl[248] vdd gnd cell_6t
Xbit_r249_c237 bl[237] br[237] wl[249] vdd gnd cell_6t
Xbit_r250_c237 bl[237] br[237] wl[250] vdd gnd cell_6t
Xbit_r251_c237 bl[237] br[237] wl[251] vdd gnd cell_6t
Xbit_r252_c237 bl[237] br[237] wl[252] vdd gnd cell_6t
Xbit_r253_c237 bl[237] br[237] wl[253] vdd gnd cell_6t
Xbit_r254_c237 bl[237] br[237] wl[254] vdd gnd cell_6t
Xbit_r255_c237 bl[237] br[237] wl[255] vdd gnd cell_6t
Xbit_r0_c238 bl[238] br[238] wl[0] vdd gnd cell_6t
Xbit_r1_c238 bl[238] br[238] wl[1] vdd gnd cell_6t
Xbit_r2_c238 bl[238] br[238] wl[2] vdd gnd cell_6t
Xbit_r3_c238 bl[238] br[238] wl[3] vdd gnd cell_6t
Xbit_r4_c238 bl[238] br[238] wl[4] vdd gnd cell_6t
Xbit_r5_c238 bl[238] br[238] wl[5] vdd gnd cell_6t
Xbit_r6_c238 bl[238] br[238] wl[6] vdd gnd cell_6t
Xbit_r7_c238 bl[238] br[238] wl[7] vdd gnd cell_6t
Xbit_r8_c238 bl[238] br[238] wl[8] vdd gnd cell_6t
Xbit_r9_c238 bl[238] br[238] wl[9] vdd gnd cell_6t
Xbit_r10_c238 bl[238] br[238] wl[10] vdd gnd cell_6t
Xbit_r11_c238 bl[238] br[238] wl[11] vdd gnd cell_6t
Xbit_r12_c238 bl[238] br[238] wl[12] vdd gnd cell_6t
Xbit_r13_c238 bl[238] br[238] wl[13] vdd gnd cell_6t
Xbit_r14_c238 bl[238] br[238] wl[14] vdd gnd cell_6t
Xbit_r15_c238 bl[238] br[238] wl[15] vdd gnd cell_6t
Xbit_r16_c238 bl[238] br[238] wl[16] vdd gnd cell_6t
Xbit_r17_c238 bl[238] br[238] wl[17] vdd gnd cell_6t
Xbit_r18_c238 bl[238] br[238] wl[18] vdd gnd cell_6t
Xbit_r19_c238 bl[238] br[238] wl[19] vdd gnd cell_6t
Xbit_r20_c238 bl[238] br[238] wl[20] vdd gnd cell_6t
Xbit_r21_c238 bl[238] br[238] wl[21] vdd gnd cell_6t
Xbit_r22_c238 bl[238] br[238] wl[22] vdd gnd cell_6t
Xbit_r23_c238 bl[238] br[238] wl[23] vdd gnd cell_6t
Xbit_r24_c238 bl[238] br[238] wl[24] vdd gnd cell_6t
Xbit_r25_c238 bl[238] br[238] wl[25] vdd gnd cell_6t
Xbit_r26_c238 bl[238] br[238] wl[26] vdd gnd cell_6t
Xbit_r27_c238 bl[238] br[238] wl[27] vdd gnd cell_6t
Xbit_r28_c238 bl[238] br[238] wl[28] vdd gnd cell_6t
Xbit_r29_c238 bl[238] br[238] wl[29] vdd gnd cell_6t
Xbit_r30_c238 bl[238] br[238] wl[30] vdd gnd cell_6t
Xbit_r31_c238 bl[238] br[238] wl[31] vdd gnd cell_6t
Xbit_r32_c238 bl[238] br[238] wl[32] vdd gnd cell_6t
Xbit_r33_c238 bl[238] br[238] wl[33] vdd gnd cell_6t
Xbit_r34_c238 bl[238] br[238] wl[34] vdd gnd cell_6t
Xbit_r35_c238 bl[238] br[238] wl[35] vdd gnd cell_6t
Xbit_r36_c238 bl[238] br[238] wl[36] vdd gnd cell_6t
Xbit_r37_c238 bl[238] br[238] wl[37] vdd gnd cell_6t
Xbit_r38_c238 bl[238] br[238] wl[38] vdd gnd cell_6t
Xbit_r39_c238 bl[238] br[238] wl[39] vdd gnd cell_6t
Xbit_r40_c238 bl[238] br[238] wl[40] vdd gnd cell_6t
Xbit_r41_c238 bl[238] br[238] wl[41] vdd gnd cell_6t
Xbit_r42_c238 bl[238] br[238] wl[42] vdd gnd cell_6t
Xbit_r43_c238 bl[238] br[238] wl[43] vdd gnd cell_6t
Xbit_r44_c238 bl[238] br[238] wl[44] vdd gnd cell_6t
Xbit_r45_c238 bl[238] br[238] wl[45] vdd gnd cell_6t
Xbit_r46_c238 bl[238] br[238] wl[46] vdd gnd cell_6t
Xbit_r47_c238 bl[238] br[238] wl[47] vdd gnd cell_6t
Xbit_r48_c238 bl[238] br[238] wl[48] vdd gnd cell_6t
Xbit_r49_c238 bl[238] br[238] wl[49] vdd gnd cell_6t
Xbit_r50_c238 bl[238] br[238] wl[50] vdd gnd cell_6t
Xbit_r51_c238 bl[238] br[238] wl[51] vdd gnd cell_6t
Xbit_r52_c238 bl[238] br[238] wl[52] vdd gnd cell_6t
Xbit_r53_c238 bl[238] br[238] wl[53] vdd gnd cell_6t
Xbit_r54_c238 bl[238] br[238] wl[54] vdd gnd cell_6t
Xbit_r55_c238 bl[238] br[238] wl[55] vdd gnd cell_6t
Xbit_r56_c238 bl[238] br[238] wl[56] vdd gnd cell_6t
Xbit_r57_c238 bl[238] br[238] wl[57] vdd gnd cell_6t
Xbit_r58_c238 bl[238] br[238] wl[58] vdd gnd cell_6t
Xbit_r59_c238 bl[238] br[238] wl[59] vdd gnd cell_6t
Xbit_r60_c238 bl[238] br[238] wl[60] vdd gnd cell_6t
Xbit_r61_c238 bl[238] br[238] wl[61] vdd gnd cell_6t
Xbit_r62_c238 bl[238] br[238] wl[62] vdd gnd cell_6t
Xbit_r63_c238 bl[238] br[238] wl[63] vdd gnd cell_6t
Xbit_r64_c238 bl[238] br[238] wl[64] vdd gnd cell_6t
Xbit_r65_c238 bl[238] br[238] wl[65] vdd gnd cell_6t
Xbit_r66_c238 bl[238] br[238] wl[66] vdd gnd cell_6t
Xbit_r67_c238 bl[238] br[238] wl[67] vdd gnd cell_6t
Xbit_r68_c238 bl[238] br[238] wl[68] vdd gnd cell_6t
Xbit_r69_c238 bl[238] br[238] wl[69] vdd gnd cell_6t
Xbit_r70_c238 bl[238] br[238] wl[70] vdd gnd cell_6t
Xbit_r71_c238 bl[238] br[238] wl[71] vdd gnd cell_6t
Xbit_r72_c238 bl[238] br[238] wl[72] vdd gnd cell_6t
Xbit_r73_c238 bl[238] br[238] wl[73] vdd gnd cell_6t
Xbit_r74_c238 bl[238] br[238] wl[74] vdd gnd cell_6t
Xbit_r75_c238 bl[238] br[238] wl[75] vdd gnd cell_6t
Xbit_r76_c238 bl[238] br[238] wl[76] vdd gnd cell_6t
Xbit_r77_c238 bl[238] br[238] wl[77] vdd gnd cell_6t
Xbit_r78_c238 bl[238] br[238] wl[78] vdd gnd cell_6t
Xbit_r79_c238 bl[238] br[238] wl[79] vdd gnd cell_6t
Xbit_r80_c238 bl[238] br[238] wl[80] vdd gnd cell_6t
Xbit_r81_c238 bl[238] br[238] wl[81] vdd gnd cell_6t
Xbit_r82_c238 bl[238] br[238] wl[82] vdd gnd cell_6t
Xbit_r83_c238 bl[238] br[238] wl[83] vdd gnd cell_6t
Xbit_r84_c238 bl[238] br[238] wl[84] vdd gnd cell_6t
Xbit_r85_c238 bl[238] br[238] wl[85] vdd gnd cell_6t
Xbit_r86_c238 bl[238] br[238] wl[86] vdd gnd cell_6t
Xbit_r87_c238 bl[238] br[238] wl[87] vdd gnd cell_6t
Xbit_r88_c238 bl[238] br[238] wl[88] vdd gnd cell_6t
Xbit_r89_c238 bl[238] br[238] wl[89] vdd gnd cell_6t
Xbit_r90_c238 bl[238] br[238] wl[90] vdd gnd cell_6t
Xbit_r91_c238 bl[238] br[238] wl[91] vdd gnd cell_6t
Xbit_r92_c238 bl[238] br[238] wl[92] vdd gnd cell_6t
Xbit_r93_c238 bl[238] br[238] wl[93] vdd gnd cell_6t
Xbit_r94_c238 bl[238] br[238] wl[94] vdd gnd cell_6t
Xbit_r95_c238 bl[238] br[238] wl[95] vdd gnd cell_6t
Xbit_r96_c238 bl[238] br[238] wl[96] vdd gnd cell_6t
Xbit_r97_c238 bl[238] br[238] wl[97] vdd gnd cell_6t
Xbit_r98_c238 bl[238] br[238] wl[98] vdd gnd cell_6t
Xbit_r99_c238 bl[238] br[238] wl[99] vdd gnd cell_6t
Xbit_r100_c238 bl[238] br[238] wl[100] vdd gnd cell_6t
Xbit_r101_c238 bl[238] br[238] wl[101] vdd gnd cell_6t
Xbit_r102_c238 bl[238] br[238] wl[102] vdd gnd cell_6t
Xbit_r103_c238 bl[238] br[238] wl[103] vdd gnd cell_6t
Xbit_r104_c238 bl[238] br[238] wl[104] vdd gnd cell_6t
Xbit_r105_c238 bl[238] br[238] wl[105] vdd gnd cell_6t
Xbit_r106_c238 bl[238] br[238] wl[106] vdd gnd cell_6t
Xbit_r107_c238 bl[238] br[238] wl[107] vdd gnd cell_6t
Xbit_r108_c238 bl[238] br[238] wl[108] vdd gnd cell_6t
Xbit_r109_c238 bl[238] br[238] wl[109] vdd gnd cell_6t
Xbit_r110_c238 bl[238] br[238] wl[110] vdd gnd cell_6t
Xbit_r111_c238 bl[238] br[238] wl[111] vdd gnd cell_6t
Xbit_r112_c238 bl[238] br[238] wl[112] vdd gnd cell_6t
Xbit_r113_c238 bl[238] br[238] wl[113] vdd gnd cell_6t
Xbit_r114_c238 bl[238] br[238] wl[114] vdd gnd cell_6t
Xbit_r115_c238 bl[238] br[238] wl[115] vdd gnd cell_6t
Xbit_r116_c238 bl[238] br[238] wl[116] vdd gnd cell_6t
Xbit_r117_c238 bl[238] br[238] wl[117] vdd gnd cell_6t
Xbit_r118_c238 bl[238] br[238] wl[118] vdd gnd cell_6t
Xbit_r119_c238 bl[238] br[238] wl[119] vdd gnd cell_6t
Xbit_r120_c238 bl[238] br[238] wl[120] vdd gnd cell_6t
Xbit_r121_c238 bl[238] br[238] wl[121] vdd gnd cell_6t
Xbit_r122_c238 bl[238] br[238] wl[122] vdd gnd cell_6t
Xbit_r123_c238 bl[238] br[238] wl[123] vdd gnd cell_6t
Xbit_r124_c238 bl[238] br[238] wl[124] vdd gnd cell_6t
Xbit_r125_c238 bl[238] br[238] wl[125] vdd gnd cell_6t
Xbit_r126_c238 bl[238] br[238] wl[126] vdd gnd cell_6t
Xbit_r127_c238 bl[238] br[238] wl[127] vdd gnd cell_6t
Xbit_r128_c238 bl[238] br[238] wl[128] vdd gnd cell_6t
Xbit_r129_c238 bl[238] br[238] wl[129] vdd gnd cell_6t
Xbit_r130_c238 bl[238] br[238] wl[130] vdd gnd cell_6t
Xbit_r131_c238 bl[238] br[238] wl[131] vdd gnd cell_6t
Xbit_r132_c238 bl[238] br[238] wl[132] vdd gnd cell_6t
Xbit_r133_c238 bl[238] br[238] wl[133] vdd gnd cell_6t
Xbit_r134_c238 bl[238] br[238] wl[134] vdd gnd cell_6t
Xbit_r135_c238 bl[238] br[238] wl[135] vdd gnd cell_6t
Xbit_r136_c238 bl[238] br[238] wl[136] vdd gnd cell_6t
Xbit_r137_c238 bl[238] br[238] wl[137] vdd gnd cell_6t
Xbit_r138_c238 bl[238] br[238] wl[138] vdd gnd cell_6t
Xbit_r139_c238 bl[238] br[238] wl[139] vdd gnd cell_6t
Xbit_r140_c238 bl[238] br[238] wl[140] vdd gnd cell_6t
Xbit_r141_c238 bl[238] br[238] wl[141] vdd gnd cell_6t
Xbit_r142_c238 bl[238] br[238] wl[142] vdd gnd cell_6t
Xbit_r143_c238 bl[238] br[238] wl[143] vdd gnd cell_6t
Xbit_r144_c238 bl[238] br[238] wl[144] vdd gnd cell_6t
Xbit_r145_c238 bl[238] br[238] wl[145] vdd gnd cell_6t
Xbit_r146_c238 bl[238] br[238] wl[146] vdd gnd cell_6t
Xbit_r147_c238 bl[238] br[238] wl[147] vdd gnd cell_6t
Xbit_r148_c238 bl[238] br[238] wl[148] vdd gnd cell_6t
Xbit_r149_c238 bl[238] br[238] wl[149] vdd gnd cell_6t
Xbit_r150_c238 bl[238] br[238] wl[150] vdd gnd cell_6t
Xbit_r151_c238 bl[238] br[238] wl[151] vdd gnd cell_6t
Xbit_r152_c238 bl[238] br[238] wl[152] vdd gnd cell_6t
Xbit_r153_c238 bl[238] br[238] wl[153] vdd gnd cell_6t
Xbit_r154_c238 bl[238] br[238] wl[154] vdd gnd cell_6t
Xbit_r155_c238 bl[238] br[238] wl[155] vdd gnd cell_6t
Xbit_r156_c238 bl[238] br[238] wl[156] vdd gnd cell_6t
Xbit_r157_c238 bl[238] br[238] wl[157] vdd gnd cell_6t
Xbit_r158_c238 bl[238] br[238] wl[158] vdd gnd cell_6t
Xbit_r159_c238 bl[238] br[238] wl[159] vdd gnd cell_6t
Xbit_r160_c238 bl[238] br[238] wl[160] vdd gnd cell_6t
Xbit_r161_c238 bl[238] br[238] wl[161] vdd gnd cell_6t
Xbit_r162_c238 bl[238] br[238] wl[162] vdd gnd cell_6t
Xbit_r163_c238 bl[238] br[238] wl[163] vdd gnd cell_6t
Xbit_r164_c238 bl[238] br[238] wl[164] vdd gnd cell_6t
Xbit_r165_c238 bl[238] br[238] wl[165] vdd gnd cell_6t
Xbit_r166_c238 bl[238] br[238] wl[166] vdd gnd cell_6t
Xbit_r167_c238 bl[238] br[238] wl[167] vdd gnd cell_6t
Xbit_r168_c238 bl[238] br[238] wl[168] vdd gnd cell_6t
Xbit_r169_c238 bl[238] br[238] wl[169] vdd gnd cell_6t
Xbit_r170_c238 bl[238] br[238] wl[170] vdd gnd cell_6t
Xbit_r171_c238 bl[238] br[238] wl[171] vdd gnd cell_6t
Xbit_r172_c238 bl[238] br[238] wl[172] vdd gnd cell_6t
Xbit_r173_c238 bl[238] br[238] wl[173] vdd gnd cell_6t
Xbit_r174_c238 bl[238] br[238] wl[174] vdd gnd cell_6t
Xbit_r175_c238 bl[238] br[238] wl[175] vdd gnd cell_6t
Xbit_r176_c238 bl[238] br[238] wl[176] vdd gnd cell_6t
Xbit_r177_c238 bl[238] br[238] wl[177] vdd gnd cell_6t
Xbit_r178_c238 bl[238] br[238] wl[178] vdd gnd cell_6t
Xbit_r179_c238 bl[238] br[238] wl[179] vdd gnd cell_6t
Xbit_r180_c238 bl[238] br[238] wl[180] vdd gnd cell_6t
Xbit_r181_c238 bl[238] br[238] wl[181] vdd gnd cell_6t
Xbit_r182_c238 bl[238] br[238] wl[182] vdd gnd cell_6t
Xbit_r183_c238 bl[238] br[238] wl[183] vdd gnd cell_6t
Xbit_r184_c238 bl[238] br[238] wl[184] vdd gnd cell_6t
Xbit_r185_c238 bl[238] br[238] wl[185] vdd gnd cell_6t
Xbit_r186_c238 bl[238] br[238] wl[186] vdd gnd cell_6t
Xbit_r187_c238 bl[238] br[238] wl[187] vdd gnd cell_6t
Xbit_r188_c238 bl[238] br[238] wl[188] vdd gnd cell_6t
Xbit_r189_c238 bl[238] br[238] wl[189] vdd gnd cell_6t
Xbit_r190_c238 bl[238] br[238] wl[190] vdd gnd cell_6t
Xbit_r191_c238 bl[238] br[238] wl[191] vdd gnd cell_6t
Xbit_r192_c238 bl[238] br[238] wl[192] vdd gnd cell_6t
Xbit_r193_c238 bl[238] br[238] wl[193] vdd gnd cell_6t
Xbit_r194_c238 bl[238] br[238] wl[194] vdd gnd cell_6t
Xbit_r195_c238 bl[238] br[238] wl[195] vdd gnd cell_6t
Xbit_r196_c238 bl[238] br[238] wl[196] vdd gnd cell_6t
Xbit_r197_c238 bl[238] br[238] wl[197] vdd gnd cell_6t
Xbit_r198_c238 bl[238] br[238] wl[198] vdd gnd cell_6t
Xbit_r199_c238 bl[238] br[238] wl[199] vdd gnd cell_6t
Xbit_r200_c238 bl[238] br[238] wl[200] vdd gnd cell_6t
Xbit_r201_c238 bl[238] br[238] wl[201] vdd gnd cell_6t
Xbit_r202_c238 bl[238] br[238] wl[202] vdd gnd cell_6t
Xbit_r203_c238 bl[238] br[238] wl[203] vdd gnd cell_6t
Xbit_r204_c238 bl[238] br[238] wl[204] vdd gnd cell_6t
Xbit_r205_c238 bl[238] br[238] wl[205] vdd gnd cell_6t
Xbit_r206_c238 bl[238] br[238] wl[206] vdd gnd cell_6t
Xbit_r207_c238 bl[238] br[238] wl[207] vdd gnd cell_6t
Xbit_r208_c238 bl[238] br[238] wl[208] vdd gnd cell_6t
Xbit_r209_c238 bl[238] br[238] wl[209] vdd gnd cell_6t
Xbit_r210_c238 bl[238] br[238] wl[210] vdd gnd cell_6t
Xbit_r211_c238 bl[238] br[238] wl[211] vdd gnd cell_6t
Xbit_r212_c238 bl[238] br[238] wl[212] vdd gnd cell_6t
Xbit_r213_c238 bl[238] br[238] wl[213] vdd gnd cell_6t
Xbit_r214_c238 bl[238] br[238] wl[214] vdd gnd cell_6t
Xbit_r215_c238 bl[238] br[238] wl[215] vdd gnd cell_6t
Xbit_r216_c238 bl[238] br[238] wl[216] vdd gnd cell_6t
Xbit_r217_c238 bl[238] br[238] wl[217] vdd gnd cell_6t
Xbit_r218_c238 bl[238] br[238] wl[218] vdd gnd cell_6t
Xbit_r219_c238 bl[238] br[238] wl[219] vdd gnd cell_6t
Xbit_r220_c238 bl[238] br[238] wl[220] vdd gnd cell_6t
Xbit_r221_c238 bl[238] br[238] wl[221] vdd gnd cell_6t
Xbit_r222_c238 bl[238] br[238] wl[222] vdd gnd cell_6t
Xbit_r223_c238 bl[238] br[238] wl[223] vdd gnd cell_6t
Xbit_r224_c238 bl[238] br[238] wl[224] vdd gnd cell_6t
Xbit_r225_c238 bl[238] br[238] wl[225] vdd gnd cell_6t
Xbit_r226_c238 bl[238] br[238] wl[226] vdd gnd cell_6t
Xbit_r227_c238 bl[238] br[238] wl[227] vdd gnd cell_6t
Xbit_r228_c238 bl[238] br[238] wl[228] vdd gnd cell_6t
Xbit_r229_c238 bl[238] br[238] wl[229] vdd gnd cell_6t
Xbit_r230_c238 bl[238] br[238] wl[230] vdd gnd cell_6t
Xbit_r231_c238 bl[238] br[238] wl[231] vdd gnd cell_6t
Xbit_r232_c238 bl[238] br[238] wl[232] vdd gnd cell_6t
Xbit_r233_c238 bl[238] br[238] wl[233] vdd gnd cell_6t
Xbit_r234_c238 bl[238] br[238] wl[234] vdd gnd cell_6t
Xbit_r235_c238 bl[238] br[238] wl[235] vdd gnd cell_6t
Xbit_r236_c238 bl[238] br[238] wl[236] vdd gnd cell_6t
Xbit_r237_c238 bl[238] br[238] wl[237] vdd gnd cell_6t
Xbit_r238_c238 bl[238] br[238] wl[238] vdd gnd cell_6t
Xbit_r239_c238 bl[238] br[238] wl[239] vdd gnd cell_6t
Xbit_r240_c238 bl[238] br[238] wl[240] vdd gnd cell_6t
Xbit_r241_c238 bl[238] br[238] wl[241] vdd gnd cell_6t
Xbit_r242_c238 bl[238] br[238] wl[242] vdd gnd cell_6t
Xbit_r243_c238 bl[238] br[238] wl[243] vdd gnd cell_6t
Xbit_r244_c238 bl[238] br[238] wl[244] vdd gnd cell_6t
Xbit_r245_c238 bl[238] br[238] wl[245] vdd gnd cell_6t
Xbit_r246_c238 bl[238] br[238] wl[246] vdd gnd cell_6t
Xbit_r247_c238 bl[238] br[238] wl[247] vdd gnd cell_6t
Xbit_r248_c238 bl[238] br[238] wl[248] vdd gnd cell_6t
Xbit_r249_c238 bl[238] br[238] wl[249] vdd gnd cell_6t
Xbit_r250_c238 bl[238] br[238] wl[250] vdd gnd cell_6t
Xbit_r251_c238 bl[238] br[238] wl[251] vdd gnd cell_6t
Xbit_r252_c238 bl[238] br[238] wl[252] vdd gnd cell_6t
Xbit_r253_c238 bl[238] br[238] wl[253] vdd gnd cell_6t
Xbit_r254_c238 bl[238] br[238] wl[254] vdd gnd cell_6t
Xbit_r255_c238 bl[238] br[238] wl[255] vdd gnd cell_6t
Xbit_r0_c239 bl[239] br[239] wl[0] vdd gnd cell_6t
Xbit_r1_c239 bl[239] br[239] wl[1] vdd gnd cell_6t
Xbit_r2_c239 bl[239] br[239] wl[2] vdd gnd cell_6t
Xbit_r3_c239 bl[239] br[239] wl[3] vdd gnd cell_6t
Xbit_r4_c239 bl[239] br[239] wl[4] vdd gnd cell_6t
Xbit_r5_c239 bl[239] br[239] wl[5] vdd gnd cell_6t
Xbit_r6_c239 bl[239] br[239] wl[6] vdd gnd cell_6t
Xbit_r7_c239 bl[239] br[239] wl[7] vdd gnd cell_6t
Xbit_r8_c239 bl[239] br[239] wl[8] vdd gnd cell_6t
Xbit_r9_c239 bl[239] br[239] wl[9] vdd gnd cell_6t
Xbit_r10_c239 bl[239] br[239] wl[10] vdd gnd cell_6t
Xbit_r11_c239 bl[239] br[239] wl[11] vdd gnd cell_6t
Xbit_r12_c239 bl[239] br[239] wl[12] vdd gnd cell_6t
Xbit_r13_c239 bl[239] br[239] wl[13] vdd gnd cell_6t
Xbit_r14_c239 bl[239] br[239] wl[14] vdd gnd cell_6t
Xbit_r15_c239 bl[239] br[239] wl[15] vdd gnd cell_6t
Xbit_r16_c239 bl[239] br[239] wl[16] vdd gnd cell_6t
Xbit_r17_c239 bl[239] br[239] wl[17] vdd gnd cell_6t
Xbit_r18_c239 bl[239] br[239] wl[18] vdd gnd cell_6t
Xbit_r19_c239 bl[239] br[239] wl[19] vdd gnd cell_6t
Xbit_r20_c239 bl[239] br[239] wl[20] vdd gnd cell_6t
Xbit_r21_c239 bl[239] br[239] wl[21] vdd gnd cell_6t
Xbit_r22_c239 bl[239] br[239] wl[22] vdd gnd cell_6t
Xbit_r23_c239 bl[239] br[239] wl[23] vdd gnd cell_6t
Xbit_r24_c239 bl[239] br[239] wl[24] vdd gnd cell_6t
Xbit_r25_c239 bl[239] br[239] wl[25] vdd gnd cell_6t
Xbit_r26_c239 bl[239] br[239] wl[26] vdd gnd cell_6t
Xbit_r27_c239 bl[239] br[239] wl[27] vdd gnd cell_6t
Xbit_r28_c239 bl[239] br[239] wl[28] vdd gnd cell_6t
Xbit_r29_c239 bl[239] br[239] wl[29] vdd gnd cell_6t
Xbit_r30_c239 bl[239] br[239] wl[30] vdd gnd cell_6t
Xbit_r31_c239 bl[239] br[239] wl[31] vdd gnd cell_6t
Xbit_r32_c239 bl[239] br[239] wl[32] vdd gnd cell_6t
Xbit_r33_c239 bl[239] br[239] wl[33] vdd gnd cell_6t
Xbit_r34_c239 bl[239] br[239] wl[34] vdd gnd cell_6t
Xbit_r35_c239 bl[239] br[239] wl[35] vdd gnd cell_6t
Xbit_r36_c239 bl[239] br[239] wl[36] vdd gnd cell_6t
Xbit_r37_c239 bl[239] br[239] wl[37] vdd gnd cell_6t
Xbit_r38_c239 bl[239] br[239] wl[38] vdd gnd cell_6t
Xbit_r39_c239 bl[239] br[239] wl[39] vdd gnd cell_6t
Xbit_r40_c239 bl[239] br[239] wl[40] vdd gnd cell_6t
Xbit_r41_c239 bl[239] br[239] wl[41] vdd gnd cell_6t
Xbit_r42_c239 bl[239] br[239] wl[42] vdd gnd cell_6t
Xbit_r43_c239 bl[239] br[239] wl[43] vdd gnd cell_6t
Xbit_r44_c239 bl[239] br[239] wl[44] vdd gnd cell_6t
Xbit_r45_c239 bl[239] br[239] wl[45] vdd gnd cell_6t
Xbit_r46_c239 bl[239] br[239] wl[46] vdd gnd cell_6t
Xbit_r47_c239 bl[239] br[239] wl[47] vdd gnd cell_6t
Xbit_r48_c239 bl[239] br[239] wl[48] vdd gnd cell_6t
Xbit_r49_c239 bl[239] br[239] wl[49] vdd gnd cell_6t
Xbit_r50_c239 bl[239] br[239] wl[50] vdd gnd cell_6t
Xbit_r51_c239 bl[239] br[239] wl[51] vdd gnd cell_6t
Xbit_r52_c239 bl[239] br[239] wl[52] vdd gnd cell_6t
Xbit_r53_c239 bl[239] br[239] wl[53] vdd gnd cell_6t
Xbit_r54_c239 bl[239] br[239] wl[54] vdd gnd cell_6t
Xbit_r55_c239 bl[239] br[239] wl[55] vdd gnd cell_6t
Xbit_r56_c239 bl[239] br[239] wl[56] vdd gnd cell_6t
Xbit_r57_c239 bl[239] br[239] wl[57] vdd gnd cell_6t
Xbit_r58_c239 bl[239] br[239] wl[58] vdd gnd cell_6t
Xbit_r59_c239 bl[239] br[239] wl[59] vdd gnd cell_6t
Xbit_r60_c239 bl[239] br[239] wl[60] vdd gnd cell_6t
Xbit_r61_c239 bl[239] br[239] wl[61] vdd gnd cell_6t
Xbit_r62_c239 bl[239] br[239] wl[62] vdd gnd cell_6t
Xbit_r63_c239 bl[239] br[239] wl[63] vdd gnd cell_6t
Xbit_r64_c239 bl[239] br[239] wl[64] vdd gnd cell_6t
Xbit_r65_c239 bl[239] br[239] wl[65] vdd gnd cell_6t
Xbit_r66_c239 bl[239] br[239] wl[66] vdd gnd cell_6t
Xbit_r67_c239 bl[239] br[239] wl[67] vdd gnd cell_6t
Xbit_r68_c239 bl[239] br[239] wl[68] vdd gnd cell_6t
Xbit_r69_c239 bl[239] br[239] wl[69] vdd gnd cell_6t
Xbit_r70_c239 bl[239] br[239] wl[70] vdd gnd cell_6t
Xbit_r71_c239 bl[239] br[239] wl[71] vdd gnd cell_6t
Xbit_r72_c239 bl[239] br[239] wl[72] vdd gnd cell_6t
Xbit_r73_c239 bl[239] br[239] wl[73] vdd gnd cell_6t
Xbit_r74_c239 bl[239] br[239] wl[74] vdd gnd cell_6t
Xbit_r75_c239 bl[239] br[239] wl[75] vdd gnd cell_6t
Xbit_r76_c239 bl[239] br[239] wl[76] vdd gnd cell_6t
Xbit_r77_c239 bl[239] br[239] wl[77] vdd gnd cell_6t
Xbit_r78_c239 bl[239] br[239] wl[78] vdd gnd cell_6t
Xbit_r79_c239 bl[239] br[239] wl[79] vdd gnd cell_6t
Xbit_r80_c239 bl[239] br[239] wl[80] vdd gnd cell_6t
Xbit_r81_c239 bl[239] br[239] wl[81] vdd gnd cell_6t
Xbit_r82_c239 bl[239] br[239] wl[82] vdd gnd cell_6t
Xbit_r83_c239 bl[239] br[239] wl[83] vdd gnd cell_6t
Xbit_r84_c239 bl[239] br[239] wl[84] vdd gnd cell_6t
Xbit_r85_c239 bl[239] br[239] wl[85] vdd gnd cell_6t
Xbit_r86_c239 bl[239] br[239] wl[86] vdd gnd cell_6t
Xbit_r87_c239 bl[239] br[239] wl[87] vdd gnd cell_6t
Xbit_r88_c239 bl[239] br[239] wl[88] vdd gnd cell_6t
Xbit_r89_c239 bl[239] br[239] wl[89] vdd gnd cell_6t
Xbit_r90_c239 bl[239] br[239] wl[90] vdd gnd cell_6t
Xbit_r91_c239 bl[239] br[239] wl[91] vdd gnd cell_6t
Xbit_r92_c239 bl[239] br[239] wl[92] vdd gnd cell_6t
Xbit_r93_c239 bl[239] br[239] wl[93] vdd gnd cell_6t
Xbit_r94_c239 bl[239] br[239] wl[94] vdd gnd cell_6t
Xbit_r95_c239 bl[239] br[239] wl[95] vdd gnd cell_6t
Xbit_r96_c239 bl[239] br[239] wl[96] vdd gnd cell_6t
Xbit_r97_c239 bl[239] br[239] wl[97] vdd gnd cell_6t
Xbit_r98_c239 bl[239] br[239] wl[98] vdd gnd cell_6t
Xbit_r99_c239 bl[239] br[239] wl[99] vdd gnd cell_6t
Xbit_r100_c239 bl[239] br[239] wl[100] vdd gnd cell_6t
Xbit_r101_c239 bl[239] br[239] wl[101] vdd gnd cell_6t
Xbit_r102_c239 bl[239] br[239] wl[102] vdd gnd cell_6t
Xbit_r103_c239 bl[239] br[239] wl[103] vdd gnd cell_6t
Xbit_r104_c239 bl[239] br[239] wl[104] vdd gnd cell_6t
Xbit_r105_c239 bl[239] br[239] wl[105] vdd gnd cell_6t
Xbit_r106_c239 bl[239] br[239] wl[106] vdd gnd cell_6t
Xbit_r107_c239 bl[239] br[239] wl[107] vdd gnd cell_6t
Xbit_r108_c239 bl[239] br[239] wl[108] vdd gnd cell_6t
Xbit_r109_c239 bl[239] br[239] wl[109] vdd gnd cell_6t
Xbit_r110_c239 bl[239] br[239] wl[110] vdd gnd cell_6t
Xbit_r111_c239 bl[239] br[239] wl[111] vdd gnd cell_6t
Xbit_r112_c239 bl[239] br[239] wl[112] vdd gnd cell_6t
Xbit_r113_c239 bl[239] br[239] wl[113] vdd gnd cell_6t
Xbit_r114_c239 bl[239] br[239] wl[114] vdd gnd cell_6t
Xbit_r115_c239 bl[239] br[239] wl[115] vdd gnd cell_6t
Xbit_r116_c239 bl[239] br[239] wl[116] vdd gnd cell_6t
Xbit_r117_c239 bl[239] br[239] wl[117] vdd gnd cell_6t
Xbit_r118_c239 bl[239] br[239] wl[118] vdd gnd cell_6t
Xbit_r119_c239 bl[239] br[239] wl[119] vdd gnd cell_6t
Xbit_r120_c239 bl[239] br[239] wl[120] vdd gnd cell_6t
Xbit_r121_c239 bl[239] br[239] wl[121] vdd gnd cell_6t
Xbit_r122_c239 bl[239] br[239] wl[122] vdd gnd cell_6t
Xbit_r123_c239 bl[239] br[239] wl[123] vdd gnd cell_6t
Xbit_r124_c239 bl[239] br[239] wl[124] vdd gnd cell_6t
Xbit_r125_c239 bl[239] br[239] wl[125] vdd gnd cell_6t
Xbit_r126_c239 bl[239] br[239] wl[126] vdd gnd cell_6t
Xbit_r127_c239 bl[239] br[239] wl[127] vdd gnd cell_6t
Xbit_r128_c239 bl[239] br[239] wl[128] vdd gnd cell_6t
Xbit_r129_c239 bl[239] br[239] wl[129] vdd gnd cell_6t
Xbit_r130_c239 bl[239] br[239] wl[130] vdd gnd cell_6t
Xbit_r131_c239 bl[239] br[239] wl[131] vdd gnd cell_6t
Xbit_r132_c239 bl[239] br[239] wl[132] vdd gnd cell_6t
Xbit_r133_c239 bl[239] br[239] wl[133] vdd gnd cell_6t
Xbit_r134_c239 bl[239] br[239] wl[134] vdd gnd cell_6t
Xbit_r135_c239 bl[239] br[239] wl[135] vdd gnd cell_6t
Xbit_r136_c239 bl[239] br[239] wl[136] vdd gnd cell_6t
Xbit_r137_c239 bl[239] br[239] wl[137] vdd gnd cell_6t
Xbit_r138_c239 bl[239] br[239] wl[138] vdd gnd cell_6t
Xbit_r139_c239 bl[239] br[239] wl[139] vdd gnd cell_6t
Xbit_r140_c239 bl[239] br[239] wl[140] vdd gnd cell_6t
Xbit_r141_c239 bl[239] br[239] wl[141] vdd gnd cell_6t
Xbit_r142_c239 bl[239] br[239] wl[142] vdd gnd cell_6t
Xbit_r143_c239 bl[239] br[239] wl[143] vdd gnd cell_6t
Xbit_r144_c239 bl[239] br[239] wl[144] vdd gnd cell_6t
Xbit_r145_c239 bl[239] br[239] wl[145] vdd gnd cell_6t
Xbit_r146_c239 bl[239] br[239] wl[146] vdd gnd cell_6t
Xbit_r147_c239 bl[239] br[239] wl[147] vdd gnd cell_6t
Xbit_r148_c239 bl[239] br[239] wl[148] vdd gnd cell_6t
Xbit_r149_c239 bl[239] br[239] wl[149] vdd gnd cell_6t
Xbit_r150_c239 bl[239] br[239] wl[150] vdd gnd cell_6t
Xbit_r151_c239 bl[239] br[239] wl[151] vdd gnd cell_6t
Xbit_r152_c239 bl[239] br[239] wl[152] vdd gnd cell_6t
Xbit_r153_c239 bl[239] br[239] wl[153] vdd gnd cell_6t
Xbit_r154_c239 bl[239] br[239] wl[154] vdd gnd cell_6t
Xbit_r155_c239 bl[239] br[239] wl[155] vdd gnd cell_6t
Xbit_r156_c239 bl[239] br[239] wl[156] vdd gnd cell_6t
Xbit_r157_c239 bl[239] br[239] wl[157] vdd gnd cell_6t
Xbit_r158_c239 bl[239] br[239] wl[158] vdd gnd cell_6t
Xbit_r159_c239 bl[239] br[239] wl[159] vdd gnd cell_6t
Xbit_r160_c239 bl[239] br[239] wl[160] vdd gnd cell_6t
Xbit_r161_c239 bl[239] br[239] wl[161] vdd gnd cell_6t
Xbit_r162_c239 bl[239] br[239] wl[162] vdd gnd cell_6t
Xbit_r163_c239 bl[239] br[239] wl[163] vdd gnd cell_6t
Xbit_r164_c239 bl[239] br[239] wl[164] vdd gnd cell_6t
Xbit_r165_c239 bl[239] br[239] wl[165] vdd gnd cell_6t
Xbit_r166_c239 bl[239] br[239] wl[166] vdd gnd cell_6t
Xbit_r167_c239 bl[239] br[239] wl[167] vdd gnd cell_6t
Xbit_r168_c239 bl[239] br[239] wl[168] vdd gnd cell_6t
Xbit_r169_c239 bl[239] br[239] wl[169] vdd gnd cell_6t
Xbit_r170_c239 bl[239] br[239] wl[170] vdd gnd cell_6t
Xbit_r171_c239 bl[239] br[239] wl[171] vdd gnd cell_6t
Xbit_r172_c239 bl[239] br[239] wl[172] vdd gnd cell_6t
Xbit_r173_c239 bl[239] br[239] wl[173] vdd gnd cell_6t
Xbit_r174_c239 bl[239] br[239] wl[174] vdd gnd cell_6t
Xbit_r175_c239 bl[239] br[239] wl[175] vdd gnd cell_6t
Xbit_r176_c239 bl[239] br[239] wl[176] vdd gnd cell_6t
Xbit_r177_c239 bl[239] br[239] wl[177] vdd gnd cell_6t
Xbit_r178_c239 bl[239] br[239] wl[178] vdd gnd cell_6t
Xbit_r179_c239 bl[239] br[239] wl[179] vdd gnd cell_6t
Xbit_r180_c239 bl[239] br[239] wl[180] vdd gnd cell_6t
Xbit_r181_c239 bl[239] br[239] wl[181] vdd gnd cell_6t
Xbit_r182_c239 bl[239] br[239] wl[182] vdd gnd cell_6t
Xbit_r183_c239 bl[239] br[239] wl[183] vdd gnd cell_6t
Xbit_r184_c239 bl[239] br[239] wl[184] vdd gnd cell_6t
Xbit_r185_c239 bl[239] br[239] wl[185] vdd gnd cell_6t
Xbit_r186_c239 bl[239] br[239] wl[186] vdd gnd cell_6t
Xbit_r187_c239 bl[239] br[239] wl[187] vdd gnd cell_6t
Xbit_r188_c239 bl[239] br[239] wl[188] vdd gnd cell_6t
Xbit_r189_c239 bl[239] br[239] wl[189] vdd gnd cell_6t
Xbit_r190_c239 bl[239] br[239] wl[190] vdd gnd cell_6t
Xbit_r191_c239 bl[239] br[239] wl[191] vdd gnd cell_6t
Xbit_r192_c239 bl[239] br[239] wl[192] vdd gnd cell_6t
Xbit_r193_c239 bl[239] br[239] wl[193] vdd gnd cell_6t
Xbit_r194_c239 bl[239] br[239] wl[194] vdd gnd cell_6t
Xbit_r195_c239 bl[239] br[239] wl[195] vdd gnd cell_6t
Xbit_r196_c239 bl[239] br[239] wl[196] vdd gnd cell_6t
Xbit_r197_c239 bl[239] br[239] wl[197] vdd gnd cell_6t
Xbit_r198_c239 bl[239] br[239] wl[198] vdd gnd cell_6t
Xbit_r199_c239 bl[239] br[239] wl[199] vdd gnd cell_6t
Xbit_r200_c239 bl[239] br[239] wl[200] vdd gnd cell_6t
Xbit_r201_c239 bl[239] br[239] wl[201] vdd gnd cell_6t
Xbit_r202_c239 bl[239] br[239] wl[202] vdd gnd cell_6t
Xbit_r203_c239 bl[239] br[239] wl[203] vdd gnd cell_6t
Xbit_r204_c239 bl[239] br[239] wl[204] vdd gnd cell_6t
Xbit_r205_c239 bl[239] br[239] wl[205] vdd gnd cell_6t
Xbit_r206_c239 bl[239] br[239] wl[206] vdd gnd cell_6t
Xbit_r207_c239 bl[239] br[239] wl[207] vdd gnd cell_6t
Xbit_r208_c239 bl[239] br[239] wl[208] vdd gnd cell_6t
Xbit_r209_c239 bl[239] br[239] wl[209] vdd gnd cell_6t
Xbit_r210_c239 bl[239] br[239] wl[210] vdd gnd cell_6t
Xbit_r211_c239 bl[239] br[239] wl[211] vdd gnd cell_6t
Xbit_r212_c239 bl[239] br[239] wl[212] vdd gnd cell_6t
Xbit_r213_c239 bl[239] br[239] wl[213] vdd gnd cell_6t
Xbit_r214_c239 bl[239] br[239] wl[214] vdd gnd cell_6t
Xbit_r215_c239 bl[239] br[239] wl[215] vdd gnd cell_6t
Xbit_r216_c239 bl[239] br[239] wl[216] vdd gnd cell_6t
Xbit_r217_c239 bl[239] br[239] wl[217] vdd gnd cell_6t
Xbit_r218_c239 bl[239] br[239] wl[218] vdd gnd cell_6t
Xbit_r219_c239 bl[239] br[239] wl[219] vdd gnd cell_6t
Xbit_r220_c239 bl[239] br[239] wl[220] vdd gnd cell_6t
Xbit_r221_c239 bl[239] br[239] wl[221] vdd gnd cell_6t
Xbit_r222_c239 bl[239] br[239] wl[222] vdd gnd cell_6t
Xbit_r223_c239 bl[239] br[239] wl[223] vdd gnd cell_6t
Xbit_r224_c239 bl[239] br[239] wl[224] vdd gnd cell_6t
Xbit_r225_c239 bl[239] br[239] wl[225] vdd gnd cell_6t
Xbit_r226_c239 bl[239] br[239] wl[226] vdd gnd cell_6t
Xbit_r227_c239 bl[239] br[239] wl[227] vdd gnd cell_6t
Xbit_r228_c239 bl[239] br[239] wl[228] vdd gnd cell_6t
Xbit_r229_c239 bl[239] br[239] wl[229] vdd gnd cell_6t
Xbit_r230_c239 bl[239] br[239] wl[230] vdd gnd cell_6t
Xbit_r231_c239 bl[239] br[239] wl[231] vdd gnd cell_6t
Xbit_r232_c239 bl[239] br[239] wl[232] vdd gnd cell_6t
Xbit_r233_c239 bl[239] br[239] wl[233] vdd gnd cell_6t
Xbit_r234_c239 bl[239] br[239] wl[234] vdd gnd cell_6t
Xbit_r235_c239 bl[239] br[239] wl[235] vdd gnd cell_6t
Xbit_r236_c239 bl[239] br[239] wl[236] vdd gnd cell_6t
Xbit_r237_c239 bl[239] br[239] wl[237] vdd gnd cell_6t
Xbit_r238_c239 bl[239] br[239] wl[238] vdd gnd cell_6t
Xbit_r239_c239 bl[239] br[239] wl[239] vdd gnd cell_6t
Xbit_r240_c239 bl[239] br[239] wl[240] vdd gnd cell_6t
Xbit_r241_c239 bl[239] br[239] wl[241] vdd gnd cell_6t
Xbit_r242_c239 bl[239] br[239] wl[242] vdd gnd cell_6t
Xbit_r243_c239 bl[239] br[239] wl[243] vdd gnd cell_6t
Xbit_r244_c239 bl[239] br[239] wl[244] vdd gnd cell_6t
Xbit_r245_c239 bl[239] br[239] wl[245] vdd gnd cell_6t
Xbit_r246_c239 bl[239] br[239] wl[246] vdd gnd cell_6t
Xbit_r247_c239 bl[239] br[239] wl[247] vdd gnd cell_6t
Xbit_r248_c239 bl[239] br[239] wl[248] vdd gnd cell_6t
Xbit_r249_c239 bl[239] br[239] wl[249] vdd gnd cell_6t
Xbit_r250_c239 bl[239] br[239] wl[250] vdd gnd cell_6t
Xbit_r251_c239 bl[239] br[239] wl[251] vdd gnd cell_6t
Xbit_r252_c239 bl[239] br[239] wl[252] vdd gnd cell_6t
Xbit_r253_c239 bl[239] br[239] wl[253] vdd gnd cell_6t
Xbit_r254_c239 bl[239] br[239] wl[254] vdd gnd cell_6t
Xbit_r255_c239 bl[239] br[239] wl[255] vdd gnd cell_6t
Xbit_r0_c240 bl[240] br[240] wl[0] vdd gnd cell_6t
Xbit_r1_c240 bl[240] br[240] wl[1] vdd gnd cell_6t
Xbit_r2_c240 bl[240] br[240] wl[2] vdd gnd cell_6t
Xbit_r3_c240 bl[240] br[240] wl[3] vdd gnd cell_6t
Xbit_r4_c240 bl[240] br[240] wl[4] vdd gnd cell_6t
Xbit_r5_c240 bl[240] br[240] wl[5] vdd gnd cell_6t
Xbit_r6_c240 bl[240] br[240] wl[6] vdd gnd cell_6t
Xbit_r7_c240 bl[240] br[240] wl[7] vdd gnd cell_6t
Xbit_r8_c240 bl[240] br[240] wl[8] vdd gnd cell_6t
Xbit_r9_c240 bl[240] br[240] wl[9] vdd gnd cell_6t
Xbit_r10_c240 bl[240] br[240] wl[10] vdd gnd cell_6t
Xbit_r11_c240 bl[240] br[240] wl[11] vdd gnd cell_6t
Xbit_r12_c240 bl[240] br[240] wl[12] vdd gnd cell_6t
Xbit_r13_c240 bl[240] br[240] wl[13] vdd gnd cell_6t
Xbit_r14_c240 bl[240] br[240] wl[14] vdd gnd cell_6t
Xbit_r15_c240 bl[240] br[240] wl[15] vdd gnd cell_6t
Xbit_r16_c240 bl[240] br[240] wl[16] vdd gnd cell_6t
Xbit_r17_c240 bl[240] br[240] wl[17] vdd gnd cell_6t
Xbit_r18_c240 bl[240] br[240] wl[18] vdd gnd cell_6t
Xbit_r19_c240 bl[240] br[240] wl[19] vdd gnd cell_6t
Xbit_r20_c240 bl[240] br[240] wl[20] vdd gnd cell_6t
Xbit_r21_c240 bl[240] br[240] wl[21] vdd gnd cell_6t
Xbit_r22_c240 bl[240] br[240] wl[22] vdd gnd cell_6t
Xbit_r23_c240 bl[240] br[240] wl[23] vdd gnd cell_6t
Xbit_r24_c240 bl[240] br[240] wl[24] vdd gnd cell_6t
Xbit_r25_c240 bl[240] br[240] wl[25] vdd gnd cell_6t
Xbit_r26_c240 bl[240] br[240] wl[26] vdd gnd cell_6t
Xbit_r27_c240 bl[240] br[240] wl[27] vdd gnd cell_6t
Xbit_r28_c240 bl[240] br[240] wl[28] vdd gnd cell_6t
Xbit_r29_c240 bl[240] br[240] wl[29] vdd gnd cell_6t
Xbit_r30_c240 bl[240] br[240] wl[30] vdd gnd cell_6t
Xbit_r31_c240 bl[240] br[240] wl[31] vdd gnd cell_6t
Xbit_r32_c240 bl[240] br[240] wl[32] vdd gnd cell_6t
Xbit_r33_c240 bl[240] br[240] wl[33] vdd gnd cell_6t
Xbit_r34_c240 bl[240] br[240] wl[34] vdd gnd cell_6t
Xbit_r35_c240 bl[240] br[240] wl[35] vdd gnd cell_6t
Xbit_r36_c240 bl[240] br[240] wl[36] vdd gnd cell_6t
Xbit_r37_c240 bl[240] br[240] wl[37] vdd gnd cell_6t
Xbit_r38_c240 bl[240] br[240] wl[38] vdd gnd cell_6t
Xbit_r39_c240 bl[240] br[240] wl[39] vdd gnd cell_6t
Xbit_r40_c240 bl[240] br[240] wl[40] vdd gnd cell_6t
Xbit_r41_c240 bl[240] br[240] wl[41] vdd gnd cell_6t
Xbit_r42_c240 bl[240] br[240] wl[42] vdd gnd cell_6t
Xbit_r43_c240 bl[240] br[240] wl[43] vdd gnd cell_6t
Xbit_r44_c240 bl[240] br[240] wl[44] vdd gnd cell_6t
Xbit_r45_c240 bl[240] br[240] wl[45] vdd gnd cell_6t
Xbit_r46_c240 bl[240] br[240] wl[46] vdd gnd cell_6t
Xbit_r47_c240 bl[240] br[240] wl[47] vdd gnd cell_6t
Xbit_r48_c240 bl[240] br[240] wl[48] vdd gnd cell_6t
Xbit_r49_c240 bl[240] br[240] wl[49] vdd gnd cell_6t
Xbit_r50_c240 bl[240] br[240] wl[50] vdd gnd cell_6t
Xbit_r51_c240 bl[240] br[240] wl[51] vdd gnd cell_6t
Xbit_r52_c240 bl[240] br[240] wl[52] vdd gnd cell_6t
Xbit_r53_c240 bl[240] br[240] wl[53] vdd gnd cell_6t
Xbit_r54_c240 bl[240] br[240] wl[54] vdd gnd cell_6t
Xbit_r55_c240 bl[240] br[240] wl[55] vdd gnd cell_6t
Xbit_r56_c240 bl[240] br[240] wl[56] vdd gnd cell_6t
Xbit_r57_c240 bl[240] br[240] wl[57] vdd gnd cell_6t
Xbit_r58_c240 bl[240] br[240] wl[58] vdd gnd cell_6t
Xbit_r59_c240 bl[240] br[240] wl[59] vdd gnd cell_6t
Xbit_r60_c240 bl[240] br[240] wl[60] vdd gnd cell_6t
Xbit_r61_c240 bl[240] br[240] wl[61] vdd gnd cell_6t
Xbit_r62_c240 bl[240] br[240] wl[62] vdd gnd cell_6t
Xbit_r63_c240 bl[240] br[240] wl[63] vdd gnd cell_6t
Xbit_r64_c240 bl[240] br[240] wl[64] vdd gnd cell_6t
Xbit_r65_c240 bl[240] br[240] wl[65] vdd gnd cell_6t
Xbit_r66_c240 bl[240] br[240] wl[66] vdd gnd cell_6t
Xbit_r67_c240 bl[240] br[240] wl[67] vdd gnd cell_6t
Xbit_r68_c240 bl[240] br[240] wl[68] vdd gnd cell_6t
Xbit_r69_c240 bl[240] br[240] wl[69] vdd gnd cell_6t
Xbit_r70_c240 bl[240] br[240] wl[70] vdd gnd cell_6t
Xbit_r71_c240 bl[240] br[240] wl[71] vdd gnd cell_6t
Xbit_r72_c240 bl[240] br[240] wl[72] vdd gnd cell_6t
Xbit_r73_c240 bl[240] br[240] wl[73] vdd gnd cell_6t
Xbit_r74_c240 bl[240] br[240] wl[74] vdd gnd cell_6t
Xbit_r75_c240 bl[240] br[240] wl[75] vdd gnd cell_6t
Xbit_r76_c240 bl[240] br[240] wl[76] vdd gnd cell_6t
Xbit_r77_c240 bl[240] br[240] wl[77] vdd gnd cell_6t
Xbit_r78_c240 bl[240] br[240] wl[78] vdd gnd cell_6t
Xbit_r79_c240 bl[240] br[240] wl[79] vdd gnd cell_6t
Xbit_r80_c240 bl[240] br[240] wl[80] vdd gnd cell_6t
Xbit_r81_c240 bl[240] br[240] wl[81] vdd gnd cell_6t
Xbit_r82_c240 bl[240] br[240] wl[82] vdd gnd cell_6t
Xbit_r83_c240 bl[240] br[240] wl[83] vdd gnd cell_6t
Xbit_r84_c240 bl[240] br[240] wl[84] vdd gnd cell_6t
Xbit_r85_c240 bl[240] br[240] wl[85] vdd gnd cell_6t
Xbit_r86_c240 bl[240] br[240] wl[86] vdd gnd cell_6t
Xbit_r87_c240 bl[240] br[240] wl[87] vdd gnd cell_6t
Xbit_r88_c240 bl[240] br[240] wl[88] vdd gnd cell_6t
Xbit_r89_c240 bl[240] br[240] wl[89] vdd gnd cell_6t
Xbit_r90_c240 bl[240] br[240] wl[90] vdd gnd cell_6t
Xbit_r91_c240 bl[240] br[240] wl[91] vdd gnd cell_6t
Xbit_r92_c240 bl[240] br[240] wl[92] vdd gnd cell_6t
Xbit_r93_c240 bl[240] br[240] wl[93] vdd gnd cell_6t
Xbit_r94_c240 bl[240] br[240] wl[94] vdd gnd cell_6t
Xbit_r95_c240 bl[240] br[240] wl[95] vdd gnd cell_6t
Xbit_r96_c240 bl[240] br[240] wl[96] vdd gnd cell_6t
Xbit_r97_c240 bl[240] br[240] wl[97] vdd gnd cell_6t
Xbit_r98_c240 bl[240] br[240] wl[98] vdd gnd cell_6t
Xbit_r99_c240 bl[240] br[240] wl[99] vdd gnd cell_6t
Xbit_r100_c240 bl[240] br[240] wl[100] vdd gnd cell_6t
Xbit_r101_c240 bl[240] br[240] wl[101] vdd gnd cell_6t
Xbit_r102_c240 bl[240] br[240] wl[102] vdd gnd cell_6t
Xbit_r103_c240 bl[240] br[240] wl[103] vdd gnd cell_6t
Xbit_r104_c240 bl[240] br[240] wl[104] vdd gnd cell_6t
Xbit_r105_c240 bl[240] br[240] wl[105] vdd gnd cell_6t
Xbit_r106_c240 bl[240] br[240] wl[106] vdd gnd cell_6t
Xbit_r107_c240 bl[240] br[240] wl[107] vdd gnd cell_6t
Xbit_r108_c240 bl[240] br[240] wl[108] vdd gnd cell_6t
Xbit_r109_c240 bl[240] br[240] wl[109] vdd gnd cell_6t
Xbit_r110_c240 bl[240] br[240] wl[110] vdd gnd cell_6t
Xbit_r111_c240 bl[240] br[240] wl[111] vdd gnd cell_6t
Xbit_r112_c240 bl[240] br[240] wl[112] vdd gnd cell_6t
Xbit_r113_c240 bl[240] br[240] wl[113] vdd gnd cell_6t
Xbit_r114_c240 bl[240] br[240] wl[114] vdd gnd cell_6t
Xbit_r115_c240 bl[240] br[240] wl[115] vdd gnd cell_6t
Xbit_r116_c240 bl[240] br[240] wl[116] vdd gnd cell_6t
Xbit_r117_c240 bl[240] br[240] wl[117] vdd gnd cell_6t
Xbit_r118_c240 bl[240] br[240] wl[118] vdd gnd cell_6t
Xbit_r119_c240 bl[240] br[240] wl[119] vdd gnd cell_6t
Xbit_r120_c240 bl[240] br[240] wl[120] vdd gnd cell_6t
Xbit_r121_c240 bl[240] br[240] wl[121] vdd gnd cell_6t
Xbit_r122_c240 bl[240] br[240] wl[122] vdd gnd cell_6t
Xbit_r123_c240 bl[240] br[240] wl[123] vdd gnd cell_6t
Xbit_r124_c240 bl[240] br[240] wl[124] vdd gnd cell_6t
Xbit_r125_c240 bl[240] br[240] wl[125] vdd gnd cell_6t
Xbit_r126_c240 bl[240] br[240] wl[126] vdd gnd cell_6t
Xbit_r127_c240 bl[240] br[240] wl[127] vdd gnd cell_6t
Xbit_r128_c240 bl[240] br[240] wl[128] vdd gnd cell_6t
Xbit_r129_c240 bl[240] br[240] wl[129] vdd gnd cell_6t
Xbit_r130_c240 bl[240] br[240] wl[130] vdd gnd cell_6t
Xbit_r131_c240 bl[240] br[240] wl[131] vdd gnd cell_6t
Xbit_r132_c240 bl[240] br[240] wl[132] vdd gnd cell_6t
Xbit_r133_c240 bl[240] br[240] wl[133] vdd gnd cell_6t
Xbit_r134_c240 bl[240] br[240] wl[134] vdd gnd cell_6t
Xbit_r135_c240 bl[240] br[240] wl[135] vdd gnd cell_6t
Xbit_r136_c240 bl[240] br[240] wl[136] vdd gnd cell_6t
Xbit_r137_c240 bl[240] br[240] wl[137] vdd gnd cell_6t
Xbit_r138_c240 bl[240] br[240] wl[138] vdd gnd cell_6t
Xbit_r139_c240 bl[240] br[240] wl[139] vdd gnd cell_6t
Xbit_r140_c240 bl[240] br[240] wl[140] vdd gnd cell_6t
Xbit_r141_c240 bl[240] br[240] wl[141] vdd gnd cell_6t
Xbit_r142_c240 bl[240] br[240] wl[142] vdd gnd cell_6t
Xbit_r143_c240 bl[240] br[240] wl[143] vdd gnd cell_6t
Xbit_r144_c240 bl[240] br[240] wl[144] vdd gnd cell_6t
Xbit_r145_c240 bl[240] br[240] wl[145] vdd gnd cell_6t
Xbit_r146_c240 bl[240] br[240] wl[146] vdd gnd cell_6t
Xbit_r147_c240 bl[240] br[240] wl[147] vdd gnd cell_6t
Xbit_r148_c240 bl[240] br[240] wl[148] vdd gnd cell_6t
Xbit_r149_c240 bl[240] br[240] wl[149] vdd gnd cell_6t
Xbit_r150_c240 bl[240] br[240] wl[150] vdd gnd cell_6t
Xbit_r151_c240 bl[240] br[240] wl[151] vdd gnd cell_6t
Xbit_r152_c240 bl[240] br[240] wl[152] vdd gnd cell_6t
Xbit_r153_c240 bl[240] br[240] wl[153] vdd gnd cell_6t
Xbit_r154_c240 bl[240] br[240] wl[154] vdd gnd cell_6t
Xbit_r155_c240 bl[240] br[240] wl[155] vdd gnd cell_6t
Xbit_r156_c240 bl[240] br[240] wl[156] vdd gnd cell_6t
Xbit_r157_c240 bl[240] br[240] wl[157] vdd gnd cell_6t
Xbit_r158_c240 bl[240] br[240] wl[158] vdd gnd cell_6t
Xbit_r159_c240 bl[240] br[240] wl[159] vdd gnd cell_6t
Xbit_r160_c240 bl[240] br[240] wl[160] vdd gnd cell_6t
Xbit_r161_c240 bl[240] br[240] wl[161] vdd gnd cell_6t
Xbit_r162_c240 bl[240] br[240] wl[162] vdd gnd cell_6t
Xbit_r163_c240 bl[240] br[240] wl[163] vdd gnd cell_6t
Xbit_r164_c240 bl[240] br[240] wl[164] vdd gnd cell_6t
Xbit_r165_c240 bl[240] br[240] wl[165] vdd gnd cell_6t
Xbit_r166_c240 bl[240] br[240] wl[166] vdd gnd cell_6t
Xbit_r167_c240 bl[240] br[240] wl[167] vdd gnd cell_6t
Xbit_r168_c240 bl[240] br[240] wl[168] vdd gnd cell_6t
Xbit_r169_c240 bl[240] br[240] wl[169] vdd gnd cell_6t
Xbit_r170_c240 bl[240] br[240] wl[170] vdd gnd cell_6t
Xbit_r171_c240 bl[240] br[240] wl[171] vdd gnd cell_6t
Xbit_r172_c240 bl[240] br[240] wl[172] vdd gnd cell_6t
Xbit_r173_c240 bl[240] br[240] wl[173] vdd gnd cell_6t
Xbit_r174_c240 bl[240] br[240] wl[174] vdd gnd cell_6t
Xbit_r175_c240 bl[240] br[240] wl[175] vdd gnd cell_6t
Xbit_r176_c240 bl[240] br[240] wl[176] vdd gnd cell_6t
Xbit_r177_c240 bl[240] br[240] wl[177] vdd gnd cell_6t
Xbit_r178_c240 bl[240] br[240] wl[178] vdd gnd cell_6t
Xbit_r179_c240 bl[240] br[240] wl[179] vdd gnd cell_6t
Xbit_r180_c240 bl[240] br[240] wl[180] vdd gnd cell_6t
Xbit_r181_c240 bl[240] br[240] wl[181] vdd gnd cell_6t
Xbit_r182_c240 bl[240] br[240] wl[182] vdd gnd cell_6t
Xbit_r183_c240 bl[240] br[240] wl[183] vdd gnd cell_6t
Xbit_r184_c240 bl[240] br[240] wl[184] vdd gnd cell_6t
Xbit_r185_c240 bl[240] br[240] wl[185] vdd gnd cell_6t
Xbit_r186_c240 bl[240] br[240] wl[186] vdd gnd cell_6t
Xbit_r187_c240 bl[240] br[240] wl[187] vdd gnd cell_6t
Xbit_r188_c240 bl[240] br[240] wl[188] vdd gnd cell_6t
Xbit_r189_c240 bl[240] br[240] wl[189] vdd gnd cell_6t
Xbit_r190_c240 bl[240] br[240] wl[190] vdd gnd cell_6t
Xbit_r191_c240 bl[240] br[240] wl[191] vdd gnd cell_6t
Xbit_r192_c240 bl[240] br[240] wl[192] vdd gnd cell_6t
Xbit_r193_c240 bl[240] br[240] wl[193] vdd gnd cell_6t
Xbit_r194_c240 bl[240] br[240] wl[194] vdd gnd cell_6t
Xbit_r195_c240 bl[240] br[240] wl[195] vdd gnd cell_6t
Xbit_r196_c240 bl[240] br[240] wl[196] vdd gnd cell_6t
Xbit_r197_c240 bl[240] br[240] wl[197] vdd gnd cell_6t
Xbit_r198_c240 bl[240] br[240] wl[198] vdd gnd cell_6t
Xbit_r199_c240 bl[240] br[240] wl[199] vdd gnd cell_6t
Xbit_r200_c240 bl[240] br[240] wl[200] vdd gnd cell_6t
Xbit_r201_c240 bl[240] br[240] wl[201] vdd gnd cell_6t
Xbit_r202_c240 bl[240] br[240] wl[202] vdd gnd cell_6t
Xbit_r203_c240 bl[240] br[240] wl[203] vdd gnd cell_6t
Xbit_r204_c240 bl[240] br[240] wl[204] vdd gnd cell_6t
Xbit_r205_c240 bl[240] br[240] wl[205] vdd gnd cell_6t
Xbit_r206_c240 bl[240] br[240] wl[206] vdd gnd cell_6t
Xbit_r207_c240 bl[240] br[240] wl[207] vdd gnd cell_6t
Xbit_r208_c240 bl[240] br[240] wl[208] vdd gnd cell_6t
Xbit_r209_c240 bl[240] br[240] wl[209] vdd gnd cell_6t
Xbit_r210_c240 bl[240] br[240] wl[210] vdd gnd cell_6t
Xbit_r211_c240 bl[240] br[240] wl[211] vdd gnd cell_6t
Xbit_r212_c240 bl[240] br[240] wl[212] vdd gnd cell_6t
Xbit_r213_c240 bl[240] br[240] wl[213] vdd gnd cell_6t
Xbit_r214_c240 bl[240] br[240] wl[214] vdd gnd cell_6t
Xbit_r215_c240 bl[240] br[240] wl[215] vdd gnd cell_6t
Xbit_r216_c240 bl[240] br[240] wl[216] vdd gnd cell_6t
Xbit_r217_c240 bl[240] br[240] wl[217] vdd gnd cell_6t
Xbit_r218_c240 bl[240] br[240] wl[218] vdd gnd cell_6t
Xbit_r219_c240 bl[240] br[240] wl[219] vdd gnd cell_6t
Xbit_r220_c240 bl[240] br[240] wl[220] vdd gnd cell_6t
Xbit_r221_c240 bl[240] br[240] wl[221] vdd gnd cell_6t
Xbit_r222_c240 bl[240] br[240] wl[222] vdd gnd cell_6t
Xbit_r223_c240 bl[240] br[240] wl[223] vdd gnd cell_6t
Xbit_r224_c240 bl[240] br[240] wl[224] vdd gnd cell_6t
Xbit_r225_c240 bl[240] br[240] wl[225] vdd gnd cell_6t
Xbit_r226_c240 bl[240] br[240] wl[226] vdd gnd cell_6t
Xbit_r227_c240 bl[240] br[240] wl[227] vdd gnd cell_6t
Xbit_r228_c240 bl[240] br[240] wl[228] vdd gnd cell_6t
Xbit_r229_c240 bl[240] br[240] wl[229] vdd gnd cell_6t
Xbit_r230_c240 bl[240] br[240] wl[230] vdd gnd cell_6t
Xbit_r231_c240 bl[240] br[240] wl[231] vdd gnd cell_6t
Xbit_r232_c240 bl[240] br[240] wl[232] vdd gnd cell_6t
Xbit_r233_c240 bl[240] br[240] wl[233] vdd gnd cell_6t
Xbit_r234_c240 bl[240] br[240] wl[234] vdd gnd cell_6t
Xbit_r235_c240 bl[240] br[240] wl[235] vdd gnd cell_6t
Xbit_r236_c240 bl[240] br[240] wl[236] vdd gnd cell_6t
Xbit_r237_c240 bl[240] br[240] wl[237] vdd gnd cell_6t
Xbit_r238_c240 bl[240] br[240] wl[238] vdd gnd cell_6t
Xbit_r239_c240 bl[240] br[240] wl[239] vdd gnd cell_6t
Xbit_r240_c240 bl[240] br[240] wl[240] vdd gnd cell_6t
Xbit_r241_c240 bl[240] br[240] wl[241] vdd gnd cell_6t
Xbit_r242_c240 bl[240] br[240] wl[242] vdd gnd cell_6t
Xbit_r243_c240 bl[240] br[240] wl[243] vdd gnd cell_6t
Xbit_r244_c240 bl[240] br[240] wl[244] vdd gnd cell_6t
Xbit_r245_c240 bl[240] br[240] wl[245] vdd gnd cell_6t
Xbit_r246_c240 bl[240] br[240] wl[246] vdd gnd cell_6t
Xbit_r247_c240 bl[240] br[240] wl[247] vdd gnd cell_6t
Xbit_r248_c240 bl[240] br[240] wl[248] vdd gnd cell_6t
Xbit_r249_c240 bl[240] br[240] wl[249] vdd gnd cell_6t
Xbit_r250_c240 bl[240] br[240] wl[250] vdd gnd cell_6t
Xbit_r251_c240 bl[240] br[240] wl[251] vdd gnd cell_6t
Xbit_r252_c240 bl[240] br[240] wl[252] vdd gnd cell_6t
Xbit_r253_c240 bl[240] br[240] wl[253] vdd gnd cell_6t
Xbit_r254_c240 bl[240] br[240] wl[254] vdd gnd cell_6t
Xbit_r255_c240 bl[240] br[240] wl[255] vdd gnd cell_6t
Xbit_r0_c241 bl[241] br[241] wl[0] vdd gnd cell_6t
Xbit_r1_c241 bl[241] br[241] wl[1] vdd gnd cell_6t
Xbit_r2_c241 bl[241] br[241] wl[2] vdd gnd cell_6t
Xbit_r3_c241 bl[241] br[241] wl[3] vdd gnd cell_6t
Xbit_r4_c241 bl[241] br[241] wl[4] vdd gnd cell_6t
Xbit_r5_c241 bl[241] br[241] wl[5] vdd gnd cell_6t
Xbit_r6_c241 bl[241] br[241] wl[6] vdd gnd cell_6t
Xbit_r7_c241 bl[241] br[241] wl[7] vdd gnd cell_6t
Xbit_r8_c241 bl[241] br[241] wl[8] vdd gnd cell_6t
Xbit_r9_c241 bl[241] br[241] wl[9] vdd gnd cell_6t
Xbit_r10_c241 bl[241] br[241] wl[10] vdd gnd cell_6t
Xbit_r11_c241 bl[241] br[241] wl[11] vdd gnd cell_6t
Xbit_r12_c241 bl[241] br[241] wl[12] vdd gnd cell_6t
Xbit_r13_c241 bl[241] br[241] wl[13] vdd gnd cell_6t
Xbit_r14_c241 bl[241] br[241] wl[14] vdd gnd cell_6t
Xbit_r15_c241 bl[241] br[241] wl[15] vdd gnd cell_6t
Xbit_r16_c241 bl[241] br[241] wl[16] vdd gnd cell_6t
Xbit_r17_c241 bl[241] br[241] wl[17] vdd gnd cell_6t
Xbit_r18_c241 bl[241] br[241] wl[18] vdd gnd cell_6t
Xbit_r19_c241 bl[241] br[241] wl[19] vdd gnd cell_6t
Xbit_r20_c241 bl[241] br[241] wl[20] vdd gnd cell_6t
Xbit_r21_c241 bl[241] br[241] wl[21] vdd gnd cell_6t
Xbit_r22_c241 bl[241] br[241] wl[22] vdd gnd cell_6t
Xbit_r23_c241 bl[241] br[241] wl[23] vdd gnd cell_6t
Xbit_r24_c241 bl[241] br[241] wl[24] vdd gnd cell_6t
Xbit_r25_c241 bl[241] br[241] wl[25] vdd gnd cell_6t
Xbit_r26_c241 bl[241] br[241] wl[26] vdd gnd cell_6t
Xbit_r27_c241 bl[241] br[241] wl[27] vdd gnd cell_6t
Xbit_r28_c241 bl[241] br[241] wl[28] vdd gnd cell_6t
Xbit_r29_c241 bl[241] br[241] wl[29] vdd gnd cell_6t
Xbit_r30_c241 bl[241] br[241] wl[30] vdd gnd cell_6t
Xbit_r31_c241 bl[241] br[241] wl[31] vdd gnd cell_6t
Xbit_r32_c241 bl[241] br[241] wl[32] vdd gnd cell_6t
Xbit_r33_c241 bl[241] br[241] wl[33] vdd gnd cell_6t
Xbit_r34_c241 bl[241] br[241] wl[34] vdd gnd cell_6t
Xbit_r35_c241 bl[241] br[241] wl[35] vdd gnd cell_6t
Xbit_r36_c241 bl[241] br[241] wl[36] vdd gnd cell_6t
Xbit_r37_c241 bl[241] br[241] wl[37] vdd gnd cell_6t
Xbit_r38_c241 bl[241] br[241] wl[38] vdd gnd cell_6t
Xbit_r39_c241 bl[241] br[241] wl[39] vdd gnd cell_6t
Xbit_r40_c241 bl[241] br[241] wl[40] vdd gnd cell_6t
Xbit_r41_c241 bl[241] br[241] wl[41] vdd gnd cell_6t
Xbit_r42_c241 bl[241] br[241] wl[42] vdd gnd cell_6t
Xbit_r43_c241 bl[241] br[241] wl[43] vdd gnd cell_6t
Xbit_r44_c241 bl[241] br[241] wl[44] vdd gnd cell_6t
Xbit_r45_c241 bl[241] br[241] wl[45] vdd gnd cell_6t
Xbit_r46_c241 bl[241] br[241] wl[46] vdd gnd cell_6t
Xbit_r47_c241 bl[241] br[241] wl[47] vdd gnd cell_6t
Xbit_r48_c241 bl[241] br[241] wl[48] vdd gnd cell_6t
Xbit_r49_c241 bl[241] br[241] wl[49] vdd gnd cell_6t
Xbit_r50_c241 bl[241] br[241] wl[50] vdd gnd cell_6t
Xbit_r51_c241 bl[241] br[241] wl[51] vdd gnd cell_6t
Xbit_r52_c241 bl[241] br[241] wl[52] vdd gnd cell_6t
Xbit_r53_c241 bl[241] br[241] wl[53] vdd gnd cell_6t
Xbit_r54_c241 bl[241] br[241] wl[54] vdd gnd cell_6t
Xbit_r55_c241 bl[241] br[241] wl[55] vdd gnd cell_6t
Xbit_r56_c241 bl[241] br[241] wl[56] vdd gnd cell_6t
Xbit_r57_c241 bl[241] br[241] wl[57] vdd gnd cell_6t
Xbit_r58_c241 bl[241] br[241] wl[58] vdd gnd cell_6t
Xbit_r59_c241 bl[241] br[241] wl[59] vdd gnd cell_6t
Xbit_r60_c241 bl[241] br[241] wl[60] vdd gnd cell_6t
Xbit_r61_c241 bl[241] br[241] wl[61] vdd gnd cell_6t
Xbit_r62_c241 bl[241] br[241] wl[62] vdd gnd cell_6t
Xbit_r63_c241 bl[241] br[241] wl[63] vdd gnd cell_6t
Xbit_r64_c241 bl[241] br[241] wl[64] vdd gnd cell_6t
Xbit_r65_c241 bl[241] br[241] wl[65] vdd gnd cell_6t
Xbit_r66_c241 bl[241] br[241] wl[66] vdd gnd cell_6t
Xbit_r67_c241 bl[241] br[241] wl[67] vdd gnd cell_6t
Xbit_r68_c241 bl[241] br[241] wl[68] vdd gnd cell_6t
Xbit_r69_c241 bl[241] br[241] wl[69] vdd gnd cell_6t
Xbit_r70_c241 bl[241] br[241] wl[70] vdd gnd cell_6t
Xbit_r71_c241 bl[241] br[241] wl[71] vdd gnd cell_6t
Xbit_r72_c241 bl[241] br[241] wl[72] vdd gnd cell_6t
Xbit_r73_c241 bl[241] br[241] wl[73] vdd gnd cell_6t
Xbit_r74_c241 bl[241] br[241] wl[74] vdd gnd cell_6t
Xbit_r75_c241 bl[241] br[241] wl[75] vdd gnd cell_6t
Xbit_r76_c241 bl[241] br[241] wl[76] vdd gnd cell_6t
Xbit_r77_c241 bl[241] br[241] wl[77] vdd gnd cell_6t
Xbit_r78_c241 bl[241] br[241] wl[78] vdd gnd cell_6t
Xbit_r79_c241 bl[241] br[241] wl[79] vdd gnd cell_6t
Xbit_r80_c241 bl[241] br[241] wl[80] vdd gnd cell_6t
Xbit_r81_c241 bl[241] br[241] wl[81] vdd gnd cell_6t
Xbit_r82_c241 bl[241] br[241] wl[82] vdd gnd cell_6t
Xbit_r83_c241 bl[241] br[241] wl[83] vdd gnd cell_6t
Xbit_r84_c241 bl[241] br[241] wl[84] vdd gnd cell_6t
Xbit_r85_c241 bl[241] br[241] wl[85] vdd gnd cell_6t
Xbit_r86_c241 bl[241] br[241] wl[86] vdd gnd cell_6t
Xbit_r87_c241 bl[241] br[241] wl[87] vdd gnd cell_6t
Xbit_r88_c241 bl[241] br[241] wl[88] vdd gnd cell_6t
Xbit_r89_c241 bl[241] br[241] wl[89] vdd gnd cell_6t
Xbit_r90_c241 bl[241] br[241] wl[90] vdd gnd cell_6t
Xbit_r91_c241 bl[241] br[241] wl[91] vdd gnd cell_6t
Xbit_r92_c241 bl[241] br[241] wl[92] vdd gnd cell_6t
Xbit_r93_c241 bl[241] br[241] wl[93] vdd gnd cell_6t
Xbit_r94_c241 bl[241] br[241] wl[94] vdd gnd cell_6t
Xbit_r95_c241 bl[241] br[241] wl[95] vdd gnd cell_6t
Xbit_r96_c241 bl[241] br[241] wl[96] vdd gnd cell_6t
Xbit_r97_c241 bl[241] br[241] wl[97] vdd gnd cell_6t
Xbit_r98_c241 bl[241] br[241] wl[98] vdd gnd cell_6t
Xbit_r99_c241 bl[241] br[241] wl[99] vdd gnd cell_6t
Xbit_r100_c241 bl[241] br[241] wl[100] vdd gnd cell_6t
Xbit_r101_c241 bl[241] br[241] wl[101] vdd gnd cell_6t
Xbit_r102_c241 bl[241] br[241] wl[102] vdd gnd cell_6t
Xbit_r103_c241 bl[241] br[241] wl[103] vdd gnd cell_6t
Xbit_r104_c241 bl[241] br[241] wl[104] vdd gnd cell_6t
Xbit_r105_c241 bl[241] br[241] wl[105] vdd gnd cell_6t
Xbit_r106_c241 bl[241] br[241] wl[106] vdd gnd cell_6t
Xbit_r107_c241 bl[241] br[241] wl[107] vdd gnd cell_6t
Xbit_r108_c241 bl[241] br[241] wl[108] vdd gnd cell_6t
Xbit_r109_c241 bl[241] br[241] wl[109] vdd gnd cell_6t
Xbit_r110_c241 bl[241] br[241] wl[110] vdd gnd cell_6t
Xbit_r111_c241 bl[241] br[241] wl[111] vdd gnd cell_6t
Xbit_r112_c241 bl[241] br[241] wl[112] vdd gnd cell_6t
Xbit_r113_c241 bl[241] br[241] wl[113] vdd gnd cell_6t
Xbit_r114_c241 bl[241] br[241] wl[114] vdd gnd cell_6t
Xbit_r115_c241 bl[241] br[241] wl[115] vdd gnd cell_6t
Xbit_r116_c241 bl[241] br[241] wl[116] vdd gnd cell_6t
Xbit_r117_c241 bl[241] br[241] wl[117] vdd gnd cell_6t
Xbit_r118_c241 bl[241] br[241] wl[118] vdd gnd cell_6t
Xbit_r119_c241 bl[241] br[241] wl[119] vdd gnd cell_6t
Xbit_r120_c241 bl[241] br[241] wl[120] vdd gnd cell_6t
Xbit_r121_c241 bl[241] br[241] wl[121] vdd gnd cell_6t
Xbit_r122_c241 bl[241] br[241] wl[122] vdd gnd cell_6t
Xbit_r123_c241 bl[241] br[241] wl[123] vdd gnd cell_6t
Xbit_r124_c241 bl[241] br[241] wl[124] vdd gnd cell_6t
Xbit_r125_c241 bl[241] br[241] wl[125] vdd gnd cell_6t
Xbit_r126_c241 bl[241] br[241] wl[126] vdd gnd cell_6t
Xbit_r127_c241 bl[241] br[241] wl[127] vdd gnd cell_6t
Xbit_r128_c241 bl[241] br[241] wl[128] vdd gnd cell_6t
Xbit_r129_c241 bl[241] br[241] wl[129] vdd gnd cell_6t
Xbit_r130_c241 bl[241] br[241] wl[130] vdd gnd cell_6t
Xbit_r131_c241 bl[241] br[241] wl[131] vdd gnd cell_6t
Xbit_r132_c241 bl[241] br[241] wl[132] vdd gnd cell_6t
Xbit_r133_c241 bl[241] br[241] wl[133] vdd gnd cell_6t
Xbit_r134_c241 bl[241] br[241] wl[134] vdd gnd cell_6t
Xbit_r135_c241 bl[241] br[241] wl[135] vdd gnd cell_6t
Xbit_r136_c241 bl[241] br[241] wl[136] vdd gnd cell_6t
Xbit_r137_c241 bl[241] br[241] wl[137] vdd gnd cell_6t
Xbit_r138_c241 bl[241] br[241] wl[138] vdd gnd cell_6t
Xbit_r139_c241 bl[241] br[241] wl[139] vdd gnd cell_6t
Xbit_r140_c241 bl[241] br[241] wl[140] vdd gnd cell_6t
Xbit_r141_c241 bl[241] br[241] wl[141] vdd gnd cell_6t
Xbit_r142_c241 bl[241] br[241] wl[142] vdd gnd cell_6t
Xbit_r143_c241 bl[241] br[241] wl[143] vdd gnd cell_6t
Xbit_r144_c241 bl[241] br[241] wl[144] vdd gnd cell_6t
Xbit_r145_c241 bl[241] br[241] wl[145] vdd gnd cell_6t
Xbit_r146_c241 bl[241] br[241] wl[146] vdd gnd cell_6t
Xbit_r147_c241 bl[241] br[241] wl[147] vdd gnd cell_6t
Xbit_r148_c241 bl[241] br[241] wl[148] vdd gnd cell_6t
Xbit_r149_c241 bl[241] br[241] wl[149] vdd gnd cell_6t
Xbit_r150_c241 bl[241] br[241] wl[150] vdd gnd cell_6t
Xbit_r151_c241 bl[241] br[241] wl[151] vdd gnd cell_6t
Xbit_r152_c241 bl[241] br[241] wl[152] vdd gnd cell_6t
Xbit_r153_c241 bl[241] br[241] wl[153] vdd gnd cell_6t
Xbit_r154_c241 bl[241] br[241] wl[154] vdd gnd cell_6t
Xbit_r155_c241 bl[241] br[241] wl[155] vdd gnd cell_6t
Xbit_r156_c241 bl[241] br[241] wl[156] vdd gnd cell_6t
Xbit_r157_c241 bl[241] br[241] wl[157] vdd gnd cell_6t
Xbit_r158_c241 bl[241] br[241] wl[158] vdd gnd cell_6t
Xbit_r159_c241 bl[241] br[241] wl[159] vdd gnd cell_6t
Xbit_r160_c241 bl[241] br[241] wl[160] vdd gnd cell_6t
Xbit_r161_c241 bl[241] br[241] wl[161] vdd gnd cell_6t
Xbit_r162_c241 bl[241] br[241] wl[162] vdd gnd cell_6t
Xbit_r163_c241 bl[241] br[241] wl[163] vdd gnd cell_6t
Xbit_r164_c241 bl[241] br[241] wl[164] vdd gnd cell_6t
Xbit_r165_c241 bl[241] br[241] wl[165] vdd gnd cell_6t
Xbit_r166_c241 bl[241] br[241] wl[166] vdd gnd cell_6t
Xbit_r167_c241 bl[241] br[241] wl[167] vdd gnd cell_6t
Xbit_r168_c241 bl[241] br[241] wl[168] vdd gnd cell_6t
Xbit_r169_c241 bl[241] br[241] wl[169] vdd gnd cell_6t
Xbit_r170_c241 bl[241] br[241] wl[170] vdd gnd cell_6t
Xbit_r171_c241 bl[241] br[241] wl[171] vdd gnd cell_6t
Xbit_r172_c241 bl[241] br[241] wl[172] vdd gnd cell_6t
Xbit_r173_c241 bl[241] br[241] wl[173] vdd gnd cell_6t
Xbit_r174_c241 bl[241] br[241] wl[174] vdd gnd cell_6t
Xbit_r175_c241 bl[241] br[241] wl[175] vdd gnd cell_6t
Xbit_r176_c241 bl[241] br[241] wl[176] vdd gnd cell_6t
Xbit_r177_c241 bl[241] br[241] wl[177] vdd gnd cell_6t
Xbit_r178_c241 bl[241] br[241] wl[178] vdd gnd cell_6t
Xbit_r179_c241 bl[241] br[241] wl[179] vdd gnd cell_6t
Xbit_r180_c241 bl[241] br[241] wl[180] vdd gnd cell_6t
Xbit_r181_c241 bl[241] br[241] wl[181] vdd gnd cell_6t
Xbit_r182_c241 bl[241] br[241] wl[182] vdd gnd cell_6t
Xbit_r183_c241 bl[241] br[241] wl[183] vdd gnd cell_6t
Xbit_r184_c241 bl[241] br[241] wl[184] vdd gnd cell_6t
Xbit_r185_c241 bl[241] br[241] wl[185] vdd gnd cell_6t
Xbit_r186_c241 bl[241] br[241] wl[186] vdd gnd cell_6t
Xbit_r187_c241 bl[241] br[241] wl[187] vdd gnd cell_6t
Xbit_r188_c241 bl[241] br[241] wl[188] vdd gnd cell_6t
Xbit_r189_c241 bl[241] br[241] wl[189] vdd gnd cell_6t
Xbit_r190_c241 bl[241] br[241] wl[190] vdd gnd cell_6t
Xbit_r191_c241 bl[241] br[241] wl[191] vdd gnd cell_6t
Xbit_r192_c241 bl[241] br[241] wl[192] vdd gnd cell_6t
Xbit_r193_c241 bl[241] br[241] wl[193] vdd gnd cell_6t
Xbit_r194_c241 bl[241] br[241] wl[194] vdd gnd cell_6t
Xbit_r195_c241 bl[241] br[241] wl[195] vdd gnd cell_6t
Xbit_r196_c241 bl[241] br[241] wl[196] vdd gnd cell_6t
Xbit_r197_c241 bl[241] br[241] wl[197] vdd gnd cell_6t
Xbit_r198_c241 bl[241] br[241] wl[198] vdd gnd cell_6t
Xbit_r199_c241 bl[241] br[241] wl[199] vdd gnd cell_6t
Xbit_r200_c241 bl[241] br[241] wl[200] vdd gnd cell_6t
Xbit_r201_c241 bl[241] br[241] wl[201] vdd gnd cell_6t
Xbit_r202_c241 bl[241] br[241] wl[202] vdd gnd cell_6t
Xbit_r203_c241 bl[241] br[241] wl[203] vdd gnd cell_6t
Xbit_r204_c241 bl[241] br[241] wl[204] vdd gnd cell_6t
Xbit_r205_c241 bl[241] br[241] wl[205] vdd gnd cell_6t
Xbit_r206_c241 bl[241] br[241] wl[206] vdd gnd cell_6t
Xbit_r207_c241 bl[241] br[241] wl[207] vdd gnd cell_6t
Xbit_r208_c241 bl[241] br[241] wl[208] vdd gnd cell_6t
Xbit_r209_c241 bl[241] br[241] wl[209] vdd gnd cell_6t
Xbit_r210_c241 bl[241] br[241] wl[210] vdd gnd cell_6t
Xbit_r211_c241 bl[241] br[241] wl[211] vdd gnd cell_6t
Xbit_r212_c241 bl[241] br[241] wl[212] vdd gnd cell_6t
Xbit_r213_c241 bl[241] br[241] wl[213] vdd gnd cell_6t
Xbit_r214_c241 bl[241] br[241] wl[214] vdd gnd cell_6t
Xbit_r215_c241 bl[241] br[241] wl[215] vdd gnd cell_6t
Xbit_r216_c241 bl[241] br[241] wl[216] vdd gnd cell_6t
Xbit_r217_c241 bl[241] br[241] wl[217] vdd gnd cell_6t
Xbit_r218_c241 bl[241] br[241] wl[218] vdd gnd cell_6t
Xbit_r219_c241 bl[241] br[241] wl[219] vdd gnd cell_6t
Xbit_r220_c241 bl[241] br[241] wl[220] vdd gnd cell_6t
Xbit_r221_c241 bl[241] br[241] wl[221] vdd gnd cell_6t
Xbit_r222_c241 bl[241] br[241] wl[222] vdd gnd cell_6t
Xbit_r223_c241 bl[241] br[241] wl[223] vdd gnd cell_6t
Xbit_r224_c241 bl[241] br[241] wl[224] vdd gnd cell_6t
Xbit_r225_c241 bl[241] br[241] wl[225] vdd gnd cell_6t
Xbit_r226_c241 bl[241] br[241] wl[226] vdd gnd cell_6t
Xbit_r227_c241 bl[241] br[241] wl[227] vdd gnd cell_6t
Xbit_r228_c241 bl[241] br[241] wl[228] vdd gnd cell_6t
Xbit_r229_c241 bl[241] br[241] wl[229] vdd gnd cell_6t
Xbit_r230_c241 bl[241] br[241] wl[230] vdd gnd cell_6t
Xbit_r231_c241 bl[241] br[241] wl[231] vdd gnd cell_6t
Xbit_r232_c241 bl[241] br[241] wl[232] vdd gnd cell_6t
Xbit_r233_c241 bl[241] br[241] wl[233] vdd gnd cell_6t
Xbit_r234_c241 bl[241] br[241] wl[234] vdd gnd cell_6t
Xbit_r235_c241 bl[241] br[241] wl[235] vdd gnd cell_6t
Xbit_r236_c241 bl[241] br[241] wl[236] vdd gnd cell_6t
Xbit_r237_c241 bl[241] br[241] wl[237] vdd gnd cell_6t
Xbit_r238_c241 bl[241] br[241] wl[238] vdd gnd cell_6t
Xbit_r239_c241 bl[241] br[241] wl[239] vdd gnd cell_6t
Xbit_r240_c241 bl[241] br[241] wl[240] vdd gnd cell_6t
Xbit_r241_c241 bl[241] br[241] wl[241] vdd gnd cell_6t
Xbit_r242_c241 bl[241] br[241] wl[242] vdd gnd cell_6t
Xbit_r243_c241 bl[241] br[241] wl[243] vdd gnd cell_6t
Xbit_r244_c241 bl[241] br[241] wl[244] vdd gnd cell_6t
Xbit_r245_c241 bl[241] br[241] wl[245] vdd gnd cell_6t
Xbit_r246_c241 bl[241] br[241] wl[246] vdd gnd cell_6t
Xbit_r247_c241 bl[241] br[241] wl[247] vdd gnd cell_6t
Xbit_r248_c241 bl[241] br[241] wl[248] vdd gnd cell_6t
Xbit_r249_c241 bl[241] br[241] wl[249] vdd gnd cell_6t
Xbit_r250_c241 bl[241] br[241] wl[250] vdd gnd cell_6t
Xbit_r251_c241 bl[241] br[241] wl[251] vdd gnd cell_6t
Xbit_r252_c241 bl[241] br[241] wl[252] vdd gnd cell_6t
Xbit_r253_c241 bl[241] br[241] wl[253] vdd gnd cell_6t
Xbit_r254_c241 bl[241] br[241] wl[254] vdd gnd cell_6t
Xbit_r255_c241 bl[241] br[241] wl[255] vdd gnd cell_6t
Xbit_r0_c242 bl[242] br[242] wl[0] vdd gnd cell_6t
Xbit_r1_c242 bl[242] br[242] wl[1] vdd gnd cell_6t
Xbit_r2_c242 bl[242] br[242] wl[2] vdd gnd cell_6t
Xbit_r3_c242 bl[242] br[242] wl[3] vdd gnd cell_6t
Xbit_r4_c242 bl[242] br[242] wl[4] vdd gnd cell_6t
Xbit_r5_c242 bl[242] br[242] wl[5] vdd gnd cell_6t
Xbit_r6_c242 bl[242] br[242] wl[6] vdd gnd cell_6t
Xbit_r7_c242 bl[242] br[242] wl[7] vdd gnd cell_6t
Xbit_r8_c242 bl[242] br[242] wl[8] vdd gnd cell_6t
Xbit_r9_c242 bl[242] br[242] wl[9] vdd gnd cell_6t
Xbit_r10_c242 bl[242] br[242] wl[10] vdd gnd cell_6t
Xbit_r11_c242 bl[242] br[242] wl[11] vdd gnd cell_6t
Xbit_r12_c242 bl[242] br[242] wl[12] vdd gnd cell_6t
Xbit_r13_c242 bl[242] br[242] wl[13] vdd gnd cell_6t
Xbit_r14_c242 bl[242] br[242] wl[14] vdd gnd cell_6t
Xbit_r15_c242 bl[242] br[242] wl[15] vdd gnd cell_6t
Xbit_r16_c242 bl[242] br[242] wl[16] vdd gnd cell_6t
Xbit_r17_c242 bl[242] br[242] wl[17] vdd gnd cell_6t
Xbit_r18_c242 bl[242] br[242] wl[18] vdd gnd cell_6t
Xbit_r19_c242 bl[242] br[242] wl[19] vdd gnd cell_6t
Xbit_r20_c242 bl[242] br[242] wl[20] vdd gnd cell_6t
Xbit_r21_c242 bl[242] br[242] wl[21] vdd gnd cell_6t
Xbit_r22_c242 bl[242] br[242] wl[22] vdd gnd cell_6t
Xbit_r23_c242 bl[242] br[242] wl[23] vdd gnd cell_6t
Xbit_r24_c242 bl[242] br[242] wl[24] vdd gnd cell_6t
Xbit_r25_c242 bl[242] br[242] wl[25] vdd gnd cell_6t
Xbit_r26_c242 bl[242] br[242] wl[26] vdd gnd cell_6t
Xbit_r27_c242 bl[242] br[242] wl[27] vdd gnd cell_6t
Xbit_r28_c242 bl[242] br[242] wl[28] vdd gnd cell_6t
Xbit_r29_c242 bl[242] br[242] wl[29] vdd gnd cell_6t
Xbit_r30_c242 bl[242] br[242] wl[30] vdd gnd cell_6t
Xbit_r31_c242 bl[242] br[242] wl[31] vdd gnd cell_6t
Xbit_r32_c242 bl[242] br[242] wl[32] vdd gnd cell_6t
Xbit_r33_c242 bl[242] br[242] wl[33] vdd gnd cell_6t
Xbit_r34_c242 bl[242] br[242] wl[34] vdd gnd cell_6t
Xbit_r35_c242 bl[242] br[242] wl[35] vdd gnd cell_6t
Xbit_r36_c242 bl[242] br[242] wl[36] vdd gnd cell_6t
Xbit_r37_c242 bl[242] br[242] wl[37] vdd gnd cell_6t
Xbit_r38_c242 bl[242] br[242] wl[38] vdd gnd cell_6t
Xbit_r39_c242 bl[242] br[242] wl[39] vdd gnd cell_6t
Xbit_r40_c242 bl[242] br[242] wl[40] vdd gnd cell_6t
Xbit_r41_c242 bl[242] br[242] wl[41] vdd gnd cell_6t
Xbit_r42_c242 bl[242] br[242] wl[42] vdd gnd cell_6t
Xbit_r43_c242 bl[242] br[242] wl[43] vdd gnd cell_6t
Xbit_r44_c242 bl[242] br[242] wl[44] vdd gnd cell_6t
Xbit_r45_c242 bl[242] br[242] wl[45] vdd gnd cell_6t
Xbit_r46_c242 bl[242] br[242] wl[46] vdd gnd cell_6t
Xbit_r47_c242 bl[242] br[242] wl[47] vdd gnd cell_6t
Xbit_r48_c242 bl[242] br[242] wl[48] vdd gnd cell_6t
Xbit_r49_c242 bl[242] br[242] wl[49] vdd gnd cell_6t
Xbit_r50_c242 bl[242] br[242] wl[50] vdd gnd cell_6t
Xbit_r51_c242 bl[242] br[242] wl[51] vdd gnd cell_6t
Xbit_r52_c242 bl[242] br[242] wl[52] vdd gnd cell_6t
Xbit_r53_c242 bl[242] br[242] wl[53] vdd gnd cell_6t
Xbit_r54_c242 bl[242] br[242] wl[54] vdd gnd cell_6t
Xbit_r55_c242 bl[242] br[242] wl[55] vdd gnd cell_6t
Xbit_r56_c242 bl[242] br[242] wl[56] vdd gnd cell_6t
Xbit_r57_c242 bl[242] br[242] wl[57] vdd gnd cell_6t
Xbit_r58_c242 bl[242] br[242] wl[58] vdd gnd cell_6t
Xbit_r59_c242 bl[242] br[242] wl[59] vdd gnd cell_6t
Xbit_r60_c242 bl[242] br[242] wl[60] vdd gnd cell_6t
Xbit_r61_c242 bl[242] br[242] wl[61] vdd gnd cell_6t
Xbit_r62_c242 bl[242] br[242] wl[62] vdd gnd cell_6t
Xbit_r63_c242 bl[242] br[242] wl[63] vdd gnd cell_6t
Xbit_r64_c242 bl[242] br[242] wl[64] vdd gnd cell_6t
Xbit_r65_c242 bl[242] br[242] wl[65] vdd gnd cell_6t
Xbit_r66_c242 bl[242] br[242] wl[66] vdd gnd cell_6t
Xbit_r67_c242 bl[242] br[242] wl[67] vdd gnd cell_6t
Xbit_r68_c242 bl[242] br[242] wl[68] vdd gnd cell_6t
Xbit_r69_c242 bl[242] br[242] wl[69] vdd gnd cell_6t
Xbit_r70_c242 bl[242] br[242] wl[70] vdd gnd cell_6t
Xbit_r71_c242 bl[242] br[242] wl[71] vdd gnd cell_6t
Xbit_r72_c242 bl[242] br[242] wl[72] vdd gnd cell_6t
Xbit_r73_c242 bl[242] br[242] wl[73] vdd gnd cell_6t
Xbit_r74_c242 bl[242] br[242] wl[74] vdd gnd cell_6t
Xbit_r75_c242 bl[242] br[242] wl[75] vdd gnd cell_6t
Xbit_r76_c242 bl[242] br[242] wl[76] vdd gnd cell_6t
Xbit_r77_c242 bl[242] br[242] wl[77] vdd gnd cell_6t
Xbit_r78_c242 bl[242] br[242] wl[78] vdd gnd cell_6t
Xbit_r79_c242 bl[242] br[242] wl[79] vdd gnd cell_6t
Xbit_r80_c242 bl[242] br[242] wl[80] vdd gnd cell_6t
Xbit_r81_c242 bl[242] br[242] wl[81] vdd gnd cell_6t
Xbit_r82_c242 bl[242] br[242] wl[82] vdd gnd cell_6t
Xbit_r83_c242 bl[242] br[242] wl[83] vdd gnd cell_6t
Xbit_r84_c242 bl[242] br[242] wl[84] vdd gnd cell_6t
Xbit_r85_c242 bl[242] br[242] wl[85] vdd gnd cell_6t
Xbit_r86_c242 bl[242] br[242] wl[86] vdd gnd cell_6t
Xbit_r87_c242 bl[242] br[242] wl[87] vdd gnd cell_6t
Xbit_r88_c242 bl[242] br[242] wl[88] vdd gnd cell_6t
Xbit_r89_c242 bl[242] br[242] wl[89] vdd gnd cell_6t
Xbit_r90_c242 bl[242] br[242] wl[90] vdd gnd cell_6t
Xbit_r91_c242 bl[242] br[242] wl[91] vdd gnd cell_6t
Xbit_r92_c242 bl[242] br[242] wl[92] vdd gnd cell_6t
Xbit_r93_c242 bl[242] br[242] wl[93] vdd gnd cell_6t
Xbit_r94_c242 bl[242] br[242] wl[94] vdd gnd cell_6t
Xbit_r95_c242 bl[242] br[242] wl[95] vdd gnd cell_6t
Xbit_r96_c242 bl[242] br[242] wl[96] vdd gnd cell_6t
Xbit_r97_c242 bl[242] br[242] wl[97] vdd gnd cell_6t
Xbit_r98_c242 bl[242] br[242] wl[98] vdd gnd cell_6t
Xbit_r99_c242 bl[242] br[242] wl[99] vdd gnd cell_6t
Xbit_r100_c242 bl[242] br[242] wl[100] vdd gnd cell_6t
Xbit_r101_c242 bl[242] br[242] wl[101] vdd gnd cell_6t
Xbit_r102_c242 bl[242] br[242] wl[102] vdd gnd cell_6t
Xbit_r103_c242 bl[242] br[242] wl[103] vdd gnd cell_6t
Xbit_r104_c242 bl[242] br[242] wl[104] vdd gnd cell_6t
Xbit_r105_c242 bl[242] br[242] wl[105] vdd gnd cell_6t
Xbit_r106_c242 bl[242] br[242] wl[106] vdd gnd cell_6t
Xbit_r107_c242 bl[242] br[242] wl[107] vdd gnd cell_6t
Xbit_r108_c242 bl[242] br[242] wl[108] vdd gnd cell_6t
Xbit_r109_c242 bl[242] br[242] wl[109] vdd gnd cell_6t
Xbit_r110_c242 bl[242] br[242] wl[110] vdd gnd cell_6t
Xbit_r111_c242 bl[242] br[242] wl[111] vdd gnd cell_6t
Xbit_r112_c242 bl[242] br[242] wl[112] vdd gnd cell_6t
Xbit_r113_c242 bl[242] br[242] wl[113] vdd gnd cell_6t
Xbit_r114_c242 bl[242] br[242] wl[114] vdd gnd cell_6t
Xbit_r115_c242 bl[242] br[242] wl[115] vdd gnd cell_6t
Xbit_r116_c242 bl[242] br[242] wl[116] vdd gnd cell_6t
Xbit_r117_c242 bl[242] br[242] wl[117] vdd gnd cell_6t
Xbit_r118_c242 bl[242] br[242] wl[118] vdd gnd cell_6t
Xbit_r119_c242 bl[242] br[242] wl[119] vdd gnd cell_6t
Xbit_r120_c242 bl[242] br[242] wl[120] vdd gnd cell_6t
Xbit_r121_c242 bl[242] br[242] wl[121] vdd gnd cell_6t
Xbit_r122_c242 bl[242] br[242] wl[122] vdd gnd cell_6t
Xbit_r123_c242 bl[242] br[242] wl[123] vdd gnd cell_6t
Xbit_r124_c242 bl[242] br[242] wl[124] vdd gnd cell_6t
Xbit_r125_c242 bl[242] br[242] wl[125] vdd gnd cell_6t
Xbit_r126_c242 bl[242] br[242] wl[126] vdd gnd cell_6t
Xbit_r127_c242 bl[242] br[242] wl[127] vdd gnd cell_6t
Xbit_r128_c242 bl[242] br[242] wl[128] vdd gnd cell_6t
Xbit_r129_c242 bl[242] br[242] wl[129] vdd gnd cell_6t
Xbit_r130_c242 bl[242] br[242] wl[130] vdd gnd cell_6t
Xbit_r131_c242 bl[242] br[242] wl[131] vdd gnd cell_6t
Xbit_r132_c242 bl[242] br[242] wl[132] vdd gnd cell_6t
Xbit_r133_c242 bl[242] br[242] wl[133] vdd gnd cell_6t
Xbit_r134_c242 bl[242] br[242] wl[134] vdd gnd cell_6t
Xbit_r135_c242 bl[242] br[242] wl[135] vdd gnd cell_6t
Xbit_r136_c242 bl[242] br[242] wl[136] vdd gnd cell_6t
Xbit_r137_c242 bl[242] br[242] wl[137] vdd gnd cell_6t
Xbit_r138_c242 bl[242] br[242] wl[138] vdd gnd cell_6t
Xbit_r139_c242 bl[242] br[242] wl[139] vdd gnd cell_6t
Xbit_r140_c242 bl[242] br[242] wl[140] vdd gnd cell_6t
Xbit_r141_c242 bl[242] br[242] wl[141] vdd gnd cell_6t
Xbit_r142_c242 bl[242] br[242] wl[142] vdd gnd cell_6t
Xbit_r143_c242 bl[242] br[242] wl[143] vdd gnd cell_6t
Xbit_r144_c242 bl[242] br[242] wl[144] vdd gnd cell_6t
Xbit_r145_c242 bl[242] br[242] wl[145] vdd gnd cell_6t
Xbit_r146_c242 bl[242] br[242] wl[146] vdd gnd cell_6t
Xbit_r147_c242 bl[242] br[242] wl[147] vdd gnd cell_6t
Xbit_r148_c242 bl[242] br[242] wl[148] vdd gnd cell_6t
Xbit_r149_c242 bl[242] br[242] wl[149] vdd gnd cell_6t
Xbit_r150_c242 bl[242] br[242] wl[150] vdd gnd cell_6t
Xbit_r151_c242 bl[242] br[242] wl[151] vdd gnd cell_6t
Xbit_r152_c242 bl[242] br[242] wl[152] vdd gnd cell_6t
Xbit_r153_c242 bl[242] br[242] wl[153] vdd gnd cell_6t
Xbit_r154_c242 bl[242] br[242] wl[154] vdd gnd cell_6t
Xbit_r155_c242 bl[242] br[242] wl[155] vdd gnd cell_6t
Xbit_r156_c242 bl[242] br[242] wl[156] vdd gnd cell_6t
Xbit_r157_c242 bl[242] br[242] wl[157] vdd gnd cell_6t
Xbit_r158_c242 bl[242] br[242] wl[158] vdd gnd cell_6t
Xbit_r159_c242 bl[242] br[242] wl[159] vdd gnd cell_6t
Xbit_r160_c242 bl[242] br[242] wl[160] vdd gnd cell_6t
Xbit_r161_c242 bl[242] br[242] wl[161] vdd gnd cell_6t
Xbit_r162_c242 bl[242] br[242] wl[162] vdd gnd cell_6t
Xbit_r163_c242 bl[242] br[242] wl[163] vdd gnd cell_6t
Xbit_r164_c242 bl[242] br[242] wl[164] vdd gnd cell_6t
Xbit_r165_c242 bl[242] br[242] wl[165] vdd gnd cell_6t
Xbit_r166_c242 bl[242] br[242] wl[166] vdd gnd cell_6t
Xbit_r167_c242 bl[242] br[242] wl[167] vdd gnd cell_6t
Xbit_r168_c242 bl[242] br[242] wl[168] vdd gnd cell_6t
Xbit_r169_c242 bl[242] br[242] wl[169] vdd gnd cell_6t
Xbit_r170_c242 bl[242] br[242] wl[170] vdd gnd cell_6t
Xbit_r171_c242 bl[242] br[242] wl[171] vdd gnd cell_6t
Xbit_r172_c242 bl[242] br[242] wl[172] vdd gnd cell_6t
Xbit_r173_c242 bl[242] br[242] wl[173] vdd gnd cell_6t
Xbit_r174_c242 bl[242] br[242] wl[174] vdd gnd cell_6t
Xbit_r175_c242 bl[242] br[242] wl[175] vdd gnd cell_6t
Xbit_r176_c242 bl[242] br[242] wl[176] vdd gnd cell_6t
Xbit_r177_c242 bl[242] br[242] wl[177] vdd gnd cell_6t
Xbit_r178_c242 bl[242] br[242] wl[178] vdd gnd cell_6t
Xbit_r179_c242 bl[242] br[242] wl[179] vdd gnd cell_6t
Xbit_r180_c242 bl[242] br[242] wl[180] vdd gnd cell_6t
Xbit_r181_c242 bl[242] br[242] wl[181] vdd gnd cell_6t
Xbit_r182_c242 bl[242] br[242] wl[182] vdd gnd cell_6t
Xbit_r183_c242 bl[242] br[242] wl[183] vdd gnd cell_6t
Xbit_r184_c242 bl[242] br[242] wl[184] vdd gnd cell_6t
Xbit_r185_c242 bl[242] br[242] wl[185] vdd gnd cell_6t
Xbit_r186_c242 bl[242] br[242] wl[186] vdd gnd cell_6t
Xbit_r187_c242 bl[242] br[242] wl[187] vdd gnd cell_6t
Xbit_r188_c242 bl[242] br[242] wl[188] vdd gnd cell_6t
Xbit_r189_c242 bl[242] br[242] wl[189] vdd gnd cell_6t
Xbit_r190_c242 bl[242] br[242] wl[190] vdd gnd cell_6t
Xbit_r191_c242 bl[242] br[242] wl[191] vdd gnd cell_6t
Xbit_r192_c242 bl[242] br[242] wl[192] vdd gnd cell_6t
Xbit_r193_c242 bl[242] br[242] wl[193] vdd gnd cell_6t
Xbit_r194_c242 bl[242] br[242] wl[194] vdd gnd cell_6t
Xbit_r195_c242 bl[242] br[242] wl[195] vdd gnd cell_6t
Xbit_r196_c242 bl[242] br[242] wl[196] vdd gnd cell_6t
Xbit_r197_c242 bl[242] br[242] wl[197] vdd gnd cell_6t
Xbit_r198_c242 bl[242] br[242] wl[198] vdd gnd cell_6t
Xbit_r199_c242 bl[242] br[242] wl[199] vdd gnd cell_6t
Xbit_r200_c242 bl[242] br[242] wl[200] vdd gnd cell_6t
Xbit_r201_c242 bl[242] br[242] wl[201] vdd gnd cell_6t
Xbit_r202_c242 bl[242] br[242] wl[202] vdd gnd cell_6t
Xbit_r203_c242 bl[242] br[242] wl[203] vdd gnd cell_6t
Xbit_r204_c242 bl[242] br[242] wl[204] vdd gnd cell_6t
Xbit_r205_c242 bl[242] br[242] wl[205] vdd gnd cell_6t
Xbit_r206_c242 bl[242] br[242] wl[206] vdd gnd cell_6t
Xbit_r207_c242 bl[242] br[242] wl[207] vdd gnd cell_6t
Xbit_r208_c242 bl[242] br[242] wl[208] vdd gnd cell_6t
Xbit_r209_c242 bl[242] br[242] wl[209] vdd gnd cell_6t
Xbit_r210_c242 bl[242] br[242] wl[210] vdd gnd cell_6t
Xbit_r211_c242 bl[242] br[242] wl[211] vdd gnd cell_6t
Xbit_r212_c242 bl[242] br[242] wl[212] vdd gnd cell_6t
Xbit_r213_c242 bl[242] br[242] wl[213] vdd gnd cell_6t
Xbit_r214_c242 bl[242] br[242] wl[214] vdd gnd cell_6t
Xbit_r215_c242 bl[242] br[242] wl[215] vdd gnd cell_6t
Xbit_r216_c242 bl[242] br[242] wl[216] vdd gnd cell_6t
Xbit_r217_c242 bl[242] br[242] wl[217] vdd gnd cell_6t
Xbit_r218_c242 bl[242] br[242] wl[218] vdd gnd cell_6t
Xbit_r219_c242 bl[242] br[242] wl[219] vdd gnd cell_6t
Xbit_r220_c242 bl[242] br[242] wl[220] vdd gnd cell_6t
Xbit_r221_c242 bl[242] br[242] wl[221] vdd gnd cell_6t
Xbit_r222_c242 bl[242] br[242] wl[222] vdd gnd cell_6t
Xbit_r223_c242 bl[242] br[242] wl[223] vdd gnd cell_6t
Xbit_r224_c242 bl[242] br[242] wl[224] vdd gnd cell_6t
Xbit_r225_c242 bl[242] br[242] wl[225] vdd gnd cell_6t
Xbit_r226_c242 bl[242] br[242] wl[226] vdd gnd cell_6t
Xbit_r227_c242 bl[242] br[242] wl[227] vdd gnd cell_6t
Xbit_r228_c242 bl[242] br[242] wl[228] vdd gnd cell_6t
Xbit_r229_c242 bl[242] br[242] wl[229] vdd gnd cell_6t
Xbit_r230_c242 bl[242] br[242] wl[230] vdd gnd cell_6t
Xbit_r231_c242 bl[242] br[242] wl[231] vdd gnd cell_6t
Xbit_r232_c242 bl[242] br[242] wl[232] vdd gnd cell_6t
Xbit_r233_c242 bl[242] br[242] wl[233] vdd gnd cell_6t
Xbit_r234_c242 bl[242] br[242] wl[234] vdd gnd cell_6t
Xbit_r235_c242 bl[242] br[242] wl[235] vdd gnd cell_6t
Xbit_r236_c242 bl[242] br[242] wl[236] vdd gnd cell_6t
Xbit_r237_c242 bl[242] br[242] wl[237] vdd gnd cell_6t
Xbit_r238_c242 bl[242] br[242] wl[238] vdd gnd cell_6t
Xbit_r239_c242 bl[242] br[242] wl[239] vdd gnd cell_6t
Xbit_r240_c242 bl[242] br[242] wl[240] vdd gnd cell_6t
Xbit_r241_c242 bl[242] br[242] wl[241] vdd gnd cell_6t
Xbit_r242_c242 bl[242] br[242] wl[242] vdd gnd cell_6t
Xbit_r243_c242 bl[242] br[242] wl[243] vdd gnd cell_6t
Xbit_r244_c242 bl[242] br[242] wl[244] vdd gnd cell_6t
Xbit_r245_c242 bl[242] br[242] wl[245] vdd gnd cell_6t
Xbit_r246_c242 bl[242] br[242] wl[246] vdd gnd cell_6t
Xbit_r247_c242 bl[242] br[242] wl[247] vdd gnd cell_6t
Xbit_r248_c242 bl[242] br[242] wl[248] vdd gnd cell_6t
Xbit_r249_c242 bl[242] br[242] wl[249] vdd gnd cell_6t
Xbit_r250_c242 bl[242] br[242] wl[250] vdd gnd cell_6t
Xbit_r251_c242 bl[242] br[242] wl[251] vdd gnd cell_6t
Xbit_r252_c242 bl[242] br[242] wl[252] vdd gnd cell_6t
Xbit_r253_c242 bl[242] br[242] wl[253] vdd gnd cell_6t
Xbit_r254_c242 bl[242] br[242] wl[254] vdd gnd cell_6t
Xbit_r255_c242 bl[242] br[242] wl[255] vdd gnd cell_6t
Xbit_r0_c243 bl[243] br[243] wl[0] vdd gnd cell_6t
Xbit_r1_c243 bl[243] br[243] wl[1] vdd gnd cell_6t
Xbit_r2_c243 bl[243] br[243] wl[2] vdd gnd cell_6t
Xbit_r3_c243 bl[243] br[243] wl[3] vdd gnd cell_6t
Xbit_r4_c243 bl[243] br[243] wl[4] vdd gnd cell_6t
Xbit_r5_c243 bl[243] br[243] wl[5] vdd gnd cell_6t
Xbit_r6_c243 bl[243] br[243] wl[6] vdd gnd cell_6t
Xbit_r7_c243 bl[243] br[243] wl[7] vdd gnd cell_6t
Xbit_r8_c243 bl[243] br[243] wl[8] vdd gnd cell_6t
Xbit_r9_c243 bl[243] br[243] wl[9] vdd gnd cell_6t
Xbit_r10_c243 bl[243] br[243] wl[10] vdd gnd cell_6t
Xbit_r11_c243 bl[243] br[243] wl[11] vdd gnd cell_6t
Xbit_r12_c243 bl[243] br[243] wl[12] vdd gnd cell_6t
Xbit_r13_c243 bl[243] br[243] wl[13] vdd gnd cell_6t
Xbit_r14_c243 bl[243] br[243] wl[14] vdd gnd cell_6t
Xbit_r15_c243 bl[243] br[243] wl[15] vdd gnd cell_6t
Xbit_r16_c243 bl[243] br[243] wl[16] vdd gnd cell_6t
Xbit_r17_c243 bl[243] br[243] wl[17] vdd gnd cell_6t
Xbit_r18_c243 bl[243] br[243] wl[18] vdd gnd cell_6t
Xbit_r19_c243 bl[243] br[243] wl[19] vdd gnd cell_6t
Xbit_r20_c243 bl[243] br[243] wl[20] vdd gnd cell_6t
Xbit_r21_c243 bl[243] br[243] wl[21] vdd gnd cell_6t
Xbit_r22_c243 bl[243] br[243] wl[22] vdd gnd cell_6t
Xbit_r23_c243 bl[243] br[243] wl[23] vdd gnd cell_6t
Xbit_r24_c243 bl[243] br[243] wl[24] vdd gnd cell_6t
Xbit_r25_c243 bl[243] br[243] wl[25] vdd gnd cell_6t
Xbit_r26_c243 bl[243] br[243] wl[26] vdd gnd cell_6t
Xbit_r27_c243 bl[243] br[243] wl[27] vdd gnd cell_6t
Xbit_r28_c243 bl[243] br[243] wl[28] vdd gnd cell_6t
Xbit_r29_c243 bl[243] br[243] wl[29] vdd gnd cell_6t
Xbit_r30_c243 bl[243] br[243] wl[30] vdd gnd cell_6t
Xbit_r31_c243 bl[243] br[243] wl[31] vdd gnd cell_6t
Xbit_r32_c243 bl[243] br[243] wl[32] vdd gnd cell_6t
Xbit_r33_c243 bl[243] br[243] wl[33] vdd gnd cell_6t
Xbit_r34_c243 bl[243] br[243] wl[34] vdd gnd cell_6t
Xbit_r35_c243 bl[243] br[243] wl[35] vdd gnd cell_6t
Xbit_r36_c243 bl[243] br[243] wl[36] vdd gnd cell_6t
Xbit_r37_c243 bl[243] br[243] wl[37] vdd gnd cell_6t
Xbit_r38_c243 bl[243] br[243] wl[38] vdd gnd cell_6t
Xbit_r39_c243 bl[243] br[243] wl[39] vdd gnd cell_6t
Xbit_r40_c243 bl[243] br[243] wl[40] vdd gnd cell_6t
Xbit_r41_c243 bl[243] br[243] wl[41] vdd gnd cell_6t
Xbit_r42_c243 bl[243] br[243] wl[42] vdd gnd cell_6t
Xbit_r43_c243 bl[243] br[243] wl[43] vdd gnd cell_6t
Xbit_r44_c243 bl[243] br[243] wl[44] vdd gnd cell_6t
Xbit_r45_c243 bl[243] br[243] wl[45] vdd gnd cell_6t
Xbit_r46_c243 bl[243] br[243] wl[46] vdd gnd cell_6t
Xbit_r47_c243 bl[243] br[243] wl[47] vdd gnd cell_6t
Xbit_r48_c243 bl[243] br[243] wl[48] vdd gnd cell_6t
Xbit_r49_c243 bl[243] br[243] wl[49] vdd gnd cell_6t
Xbit_r50_c243 bl[243] br[243] wl[50] vdd gnd cell_6t
Xbit_r51_c243 bl[243] br[243] wl[51] vdd gnd cell_6t
Xbit_r52_c243 bl[243] br[243] wl[52] vdd gnd cell_6t
Xbit_r53_c243 bl[243] br[243] wl[53] vdd gnd cell_6t
Xbit_r54_c243 bl[243] br[243] wl[54] vdd gnd cell_6t
Xbit_r55_c243 bl[243] br[243] wl[55] vdd gnd cell_6t
Xbit_r56_c243 bl[243] br[243] wl[56] vdd gnd cell_6t
Xbit_r57_c243 bl[243] br[243] wl[57] vdd gnd cell_6t
Xbit_r58_c243 bl[243] br[243] wl[58] vdd gnd cell_6t
Xbit_r59_c243 bl[243] br[243] wl[59] vdd gnd cell_6t
Xbit_r60_c243 bl[243] br[243] wl[60] vdd gnd cell_6t
Xbit_r61_c243 bl[243] br[243] wl[61] vdd gnd cell_6t
Xbit_r62_c243 bl[243] br[243] wl[62] vdd gnd cell_6t
Xbit_r63_c243 bl[243] br[243] wl[63] vdd gnd cell_6t
Xbit_r64_c243 bl[243] br[243] wl[64] vdd gnd cell_6t
Xbit_r65_c243 bl[243] br[243] wl[65] vdd gnd cell_6t
Xbit_r66_c243 bl[243] br[243] wl[66] vdd gnd cell_6t
Xbit_r67_c243 bl[243] br[243] wl[67] vdd gnd cell_6t
Xbit_r68_c243 bl[243] br[243] wl[68] vdd gnd cell_6t
Xbit_r69_c243 bl[243] br[243] wl[69] vdd gnd cell_6t
Xbit_r70_c243 bl[243] br[243] wl[70] vdd gnd cell_6t
Xbit_r71_c243 bl[243] br[243] wl[71] vdd gnd cell_6t
Xbit_r72_c243 bl[243] br[243] wl[72] vdd gnd cell_6t
Xbit_r73_c243 bl[243] br[243] wl[73] vdd gnd cell_6t
Xbit_r74_c243 bl[243] br[243] wl[74] vdd gnd cell_6t
Xbit_r75_c243 bl[243] br[243] wl[75] vdd gnd cell_6t
Xbit_r76_c243 bl[243] br[243] wl[76] vdd gnd cell_6t
Xbit_r77_c243 bl[243] br[243] wl[77] vdd gnd cell_6t
Xbit_r78_c243 bl[243] br[243] wl[78] vdd gnd cell_6t
Xbit_r79_c243 bl[243] br[243] wl[79] vdd gnd cell_6t
Xbit_r80_c243 bl[243] br[243] wl[80] vdd gnd cell_6t
Xbit_r81_c243 bl[243] br[243] wl[81] vdd gnd cell_6t
Xbit_r82_c243 bl[243] br[243] wl[82] vdd gnd cell_6t
Xbit_r83_c243 bl[243] br[243] wl[83] vdd gnd cell_6t
Xbit_r84_c243 bl[243] br[243] wl[84] vdd gnd cell_6t
Xbit_r85_c243 bl[243] br[243] wl[85] vdd gnd cell_6t
Xbit_r86_c243 bl[243] br[243] wl[86] vdd gnd cell_6t
Xbit_r87_c243 bl[243] br[243] wl[87] vdd gnd cell_6t
Xbit_r88_c243 bl[243] br[243] wl[88] vdd gnd cell_6t
Xbit_r89_c243 bl[243] br[243] wl[89] vdd gnd cell_6t
Xbit_r90_c243 bl[243] br[243] wl[90] vdd gnd cell_6t
Xbit_r91_c243 bl[243] br[243] wl[91] vdd gnd cell_6t
Xbit_r92_c243 bl[243] br[243] wl[92] vdd gnd cell_6t
Xbit_r93_c243 bl[243] br[243] wl[93] vdd gnd cell_6t
Xbit_r94_c243 bl[243] br[243] wl[94] vdd gnd cell_6t
Xbit_r95_c243 bl[243] br[243] wl[95] vdd gnd cell_6t
Xbit_r96_c243 bl[243] br[243] wl[96] vdd gnd cell_6t
Xbit_r97_c243 bl[243] br[243] wl[97] vdd gnd cell_6t
Xbit_r98_c243 bl[243] br[243] wl[98] vdd gnd cell_6t
Xbit_r99_c243 bl[243] br[243] wl[99] vdd gnd cell_6t
Xbit_r100_c243 bl[243] br[243] wl[100] vdd gnd cell_6t
Xbit_r101_c243 bl[243] br[243] wl[101] vdd gnd cell_6t
Xbit_r102_c243 bl[243] br[243] wl[102] vdd gnd cell_6t
Xbit_r103_c243 bl[243] br[243] wl[103] vdd gnd cell_6t
Xbit_r104_c243 bl[243] br[243] wl[104] vdd gnd cell_6t
Xbit_r105_c243 bl[243] br[243] wl[105] vdd gnd cell_6t
Xbit_r106_c243 bl[243] br[243] wl[106] vdd gnd cell_6t
Xbit_r107_c243 bl[243] br[243] wl[107] vdd gnd cell_6t
Xbit_r108_c243 bl[243] br[243] wl[108] vdd gnd cell_6t
Xbit_r109_c243 bl[243] br[243] wl[109] vdd gnd cell_6t
Xbit_r110_c243 bl[243] br[243] wl[110] vdd gnd cell_6t
Xbit_r111_c243 bl[243] br[243] wl[111] vdd gnd cell_6t
Xbit_r112_c243 bl[243] br[243] wl[112] vdd gnd cell_6t
Xbit_r113_c243 bl[243] br[243] wl[113] vdd gnd cell_6t
Xbit_r114_c243 bl[243] br[243] wl[114] vdd gnd cell_6t
Xbit_r115_c243 bl[243] br[243] wl[115] vdd gnd cell_6t
Xbit_r116_c243 bl[243] br[243] wl[116] vdd gnd cell_6t
Xbit_r117_c243 bl[243] br[243] wl[117] vdd gnd cell_6t
Xbit_r118_c243 bl[243] br[243] wl[118] vdd gnd cell_6t
Xbit_r119_c243 bl[243] br[243] wl[119] vdd gnd cell_6t
Xbit_r120_c243 bl[243] br[243] wl[120] vdd gnd cell_6t
Xbit_r121_c243 bl[243] br[243] wl[121] vdd gnd cell_6t
Xbit_r122_c243 bl[243] br[243] wl[122] vdd gnd cell_6t
Xbit_r123_c243 bl[243] br[243] wl[123] vdd gnd cell_6t
Xbit_r124_c243 bl[243] br[243] wl[124] vdd gnd cell_6t
Xbit_r125_c243 bl[243] br[243] wl[125] vdd gnd cell_6t
Xbit_r126_c243 bl[243] br[243] wl[126] vdd gnd cell_6t
Xbit_r127_c243 bl[243] br[243] wl[127] vdd gnd cell_6t
Xbit_r128_c243 bl[243] br[243] wl[128] vdd gnd cell_6t
Xbit_r129_c243 bl[243] br[243] wl[129] vdd gnd cell_6t
Xbit_r130_c243 bl[243] br[243] wl[130] vdd gnd cell_6t
Xbit_r131_c243 bl[243] br[243] wl[131] vdd gnd cell_6t
Xbit_r132_c243 bl[243] br[243] wl[132] vdd gnd cell_6t
Xbit_r133_c243 bl[243] br[243] wl[133] vdd gnd cell_6t
Xbit_r134_c243 bl[243] br[243] wl[134] vdd gnd cell_6t
Xbit_r135_c243 bl[243] br[243] wl[135] vdd gnd cell_6t
Xbit_r136_c243 bl[243] br[243] wl[136] vdd gnd cell_6t
Xbit_r137_c243 bl[243] br[243] wl[137] vdd gnd cell_6t
Xbit_r138_c243 bl[243] br[243] wl[138] vdd gnd cell_6t
Xbit_r139_c243 bl[243] br[243] wl[139] vdd gnd cell_6t
Xbit_r140_c243 bl[243] br[243] wl[140] vdd gnd cell_6t
Xbit_r141_c243 bl[243] br[243] wl[141] vdd gnd cell_6t
Xbit_r142_c243 bl[243] br[243] wl[142] vdd gnd cell_6t
Xbit_r143_c243 bl[243] br[243] wl[143] vdd gnd cell_6t
Xbit_r144_c243 bl[243] br[243] wl[144] vdd gnd cell_6t
Xbit_r145_c243 bl[243] br[243] wl[145] vdd gnd cell_6t
Xbit_r146_c243 bl[243] br[243] wl[146] vdd gnd cell_6t
Xbit_r147_c243 bl[243] br[243] wl[147] vdd gnd cell_6t
Xbit_r148_c243 bl[243] br[243] wl[148] vdd gnd cell_6t
Xbit_r149_c243 bl[243] br[243] wl[149] vdd gnd cell_6t
Xbit_r150_c243 bl[243] br[243] wl[150] vdd gnd cell_6t
Xbit_r151_c243 bl[243] br[243] wl[151] vdd gnd cell_6t
Xbit_r152_c243 bl[243] br[243] wl[152] vdd gnd cell_6t
Xbit_r153_c243 bl[243] br[243] wl[153] vdd gnd cell_6t
Xbit_r154_c243 bl[243] br[243] wl[154] vdd gnd cell_6t
Xbit_r155_c243 bl[243] br[243] wl[155] vdd gnd cell_6t
Xbit_r156_c243 bl[243] br[243] wl[156] vdd gnd cell_6t
Xbit_r157_c243 bl[243] br[243] wl[157] vdd gnd cell_6t
Xbit_r158_c243 bl[243] br[243] wl[158] vdd gnd cell_6t
Xbit_r159_c243 bl[243] br[243] wl[159] vdd gnd cell_6t
Xbit_r160_c243 bl[243] br[243] wl[160] vdd gnd cell_6t
Xbit_r161_c243 bl[243] br[243] wl[161] vdd gnd cell_6t
Xbit_r162_c243 bl[243] br[243] wl[162] vdd gnd cell_6t
Xbit_r163_c243 bl[243] br[243] wl[163] vdd gnd cell_6t
Xbit_r164_c243 bl[243] br[243] wl[164] vdd gnd cell_6t
Xbit_r165_c243 bl[243] br[243] wl[165] vdd gnd cell_6t
Xbit_r166_c243 bl[243] br[243] wl[166] vdd gnd cell_6t
Xbit_r167_c243 bl[243] br[243] wl[167] vdd gnd cell_6t
Xbit_r168_c243 bl[243] br[243] wl[168] vdd gnd cell_6t
Xbit_r169_c243 bl[243] br[243] wl[169] vdd gnd cell_6t
Xbit_r170_c243 bl[243] br[243] wl[170] vdd gnd cell_6t
Xbit_r171_c243 bl[243] br[243] wl[171] vdd gnd cell_6t
Xbit_r172_c243 bl[243] br[243] wl[172] vdd gnd cell_6t
Xbit_r173_c243 bl[243] br[243] wl[173] vdd gnd cell_6t
Xbit_r174_c243 bl[243] br[243] wl[174] vdd gnd cell_6t
Xbit_r175_c243 bl[243] br[243] wl[175] vdd gnd cell_6t
Xbit_r176_c243 bl[243] br[243] wl[176] vdd gnd cell_6t
Xbit_r177_c243 bl[243] br[243] wl[177] vdd gnd cell_6t
Xbit_r178_c243 bl[243] br[243] wl[178] vdd gnd cell_6t
Xbit_r179_c243 bl[243] br[243] wl[179] vdd gnd cell_6t
Xbit_r180_c243 bl[243] br[243] wl[180] vdd gnd cell_6t
Xbit_r181_c243 bl[243] br[243] wl[181] vdd gnd cell_6t
Xbit_r182_c243 bl[243] br[243] wl[182] vdd gnd cell_6t
Xbit_r183_c243 bl[243] br[243] wl[183] vdd gnd cell_6t
Xbit_r184_c243 bl[243] br[243] wl[184] vdd gnd cell_6t
Xbit_r185_c243 bl[243] br[243] wl[185] vdd gnd cell_6t
Xbit_r186_c243 bl[243] br[243] wl[186] vdd gnd cell_6t
Xbit_r187_c243 bl[243] br[243] wl[187] vdd gnd cell_6t
Xbit_r188_c243 bl[243] br[243] wl[188] vdd gnd cell_6t
Xbit_r189_c243 bl[243] br[243] wl[189] vdd gnd cell_6t
Xbit_r190_c243 bl[243] br[243] wl[190] vdd gnd cell_6t
Xbit_r191_c243 bl[243] br[243] wl[191] vdd gnd cell_6t
Xbit_r192_c243 bl[243] br[243] wl[192] vdd gnd cell_6t
Xbit_r193_c243 bl[243] br[243] wl[193] vdd gnd cell_6t
Xbit_r194_c243 bl[243] br[243] wl[194] vdd gnd cell_6t
Xbit_r195_c243 bl[243] br[243] wl[195] vdd gnd cell_6t
Xbit_r196_c243 bl[243] br[243] wl[196] vdd gnd cell_6t
Xbit_r197_c243 bl[243] br[243] wl[197] vdd gnd cell_6t
Xbit_r198_c243 bl[243] br[243] wl[198] vdd gnd cell_6t
Xbit_r199_c243 bl[243] br[243] wl[199] vdd gnd cell_6t
Xbit_r200_c243 bl[243] br[243] wl[200] vdd gnd cell_6t
Xbit_r201_c243 bl[243] br[243] wl[201] vdd gnd cell_6t
Xbit_r202_c243 bl[243] br[243] wl[202] vdd gnd cell_6t
Xbit_r203_c243 bl[243] br[243] wl[203] vdd gnd cell_6t
Xbit_r204_c243 bl[243] br[243] wl[204] vdd gnd cell_6t
Xbit_r205_c243 bl[243] br[243] wl[205] vdd gnd cell_6t
Xbit_r206_c243 bl[243] br[243] wl[206] vdd gnd cell_6t
Xbit_r207_c243 bl[243] br[243] wl[207] vdd gnd cell_6t
Xbit_r208_c243 bl[243] br[243] wl[208] vdd gnd cell_6t
Xbit_r209_c243 bl[243] br[243] wl[209] vdd gnd cell_6t
Xbit_r210_c243 bl[243] br[243] wl[210] vdd gnd cell_6t
Xbit_r211_c243 bl[243] br[243] wl[211] vdd gnd cell_6t
Xbit_r212_c243 bl[243] br[243] wl[212] vdd gnd cell_6t
Xbit_r213_c243 bl[243] br[243] wl[213] vdd gnd cell_6t
Xbit_r214_c243 bl[243] br[243] wl[214] vdd gnd cell_6t
Xbit_r215_c243 bl[243] br[243] wl[215] vdd gnd cell_6t
Xbit_r216_c243 bl[243] br[243] wl[216] vdd gnd cell_6t
Xbit_r217_c243 bl[243] br[243] wl[217] vdd gnd cell_6t
Xbit_r218_c243 bl[243] br[243] wl[218] vdd gnd cell_6t
Xbit_r219_c243 bl[243] br[243] wl[219] vdd gnd cell_6t
Xbit_r220_c243 bl[243] br[243] wl[220] vdd gnd cell_6t
Xbit_r221_c243 bl[243] br[243] wl[221] vdd gnd cell_6t
Xbit_r222_c243 bl[243] br[243] wl[222] vdd gnd cell_6t
Xbit_r223_c243 bl[243] br[243] wl[223] vdd gnd cell_6t
Xbit_r224_c243 bl[243] br[243] wl[224] vdd gnd cell_6t
Xbit_r225_c243 bl[243] br[243] wl[225] vdd gnd cell_6t
Xbit_r226_c243 bl[243] br[243] wl[226] vdd gnd cell_6t
Xbit_r227_c243 bl[243] br[243] wl[227] vdd gnd cell_6t
Xbit_r228_c243 bl[243] br[243] wl[228] vdd gnd cell_6t
Xbit_r229_c243 bl[243] br[243] wl[229] vdd gnd cell_6t
Xbit_r230_c243 bl[243] br[243] wl[230] vdd gnd cell_6t
Xbit_r231_c243 bl[243] br[243] wl[231] vdd gnd cell_6t
Xbit_r232_c243 bl[243] br[243] wl[232] vdd gnd cell_6t
Xbit_r233_c243 bl[243] br[243] wl[233] vdd gnd cell_6t
Xbit_r234_c243 bl[243] br[243] wl[234] vdd gnd cell_6t
Xbit_r235_c243 bl[243] br[243] wl[235] vdd gnd cell_6t
Xbit_r236_c243 bl[243] br[243] wl[236] vdd gnd cell_6t
Xbit_r237_c243 bl[243] br[243] wl[237] vdd gnd cell_6t
Xbit_r238_c243 bl[243] br[243] wl[238] vdd gnd cell_6t
Xbit_r239_c243 bl[243] br[243] wl[239] vdd gnd cell_6t
Xbit_r240_c243 bl[243] br[243] wl[240] vdd gnd cell_6t
Xbit_r241_c243 bl[243] br[243] wl[241] vdd gnd cell_6t
Xbit_r242_c243 bl[243] br[243] wl[242] vdd gnd cell_6t
Xbit_r243_c243 bl[243] br[243] wl[243] vdd gnd cell_6t
Xbit_r244_c243 bl[243] br[243] wl[244] vdd gnd cell_6t
Xbit_r245_c243 bl[243] br[243] wl[245] vdd gnd cell_6t
Xbit_r246_c243 bl[243] br[243] wl[246] vdd gnd cell_6t
Xbit_r247_c243 bl[243] br[243] wl[247] vdd gnd cell_6t
Xbit_r248_c243 bl[243] br[243] wl[248] vdd gnd cell_6t
Xbit_r249_c243 bl[243] br[243] wl[249] vdd gnd cell_6t
Xbit_r250_c243 bl[243] br[243] wl[250] vdd gnd cell_6t
Xbit_r251_c243 bl[243] br[243] wl[251] vdd gnd cell_6t
Xbit_r252_c243 bl[243] br[243] wl[252] vdd gnd cell_6t
Xbit_r253_c243 bl[243] br[243] wl[253] vdd gnd cell_6t
Xbit_r254_c243 bl[243] br[243] wl[254] vdd gnd cell_6t
Xbit_r255_c243 bl[243] br[243] wl[255] vdd gnd cell_6t
Xbit_r0_c244 bl[244] br[244] wl[0] vdd gnd cell_6t
Xbit_r1_c244 bl[244] br[244] wl[1] vdd gnd cell_6t
Xbit_r2_c244 bl[244] br[244] wl[2] vdd gnd cell_6t
Xbit_r3_c244 bl[244] br[244] wl[3] vdd gnd cell_6t
Xbit_r4_c244 bl[244] br[244] wl[4] vdd gnd cell_6t
Xbit_r5_c244 bl[244] br[244] wl[5] vdd gnd cell_6t
Xbit_r6_c244 bl[244] br[244] wl[6] vdd gnd cell_6t
Xbit_r7_c244 bl[244] br[244] wl[7] vdd gnd cell_6t
Xbit_r8_c244 bl[244] br[244] wl[8] vdd gnd cell_6t
Xbit_r9_c244 bl[244] br[244] wl[9] vdd gnd cell_6t
Xbit_r10_c244 bl[244] br[244] wl[10] vdd gnd cell_6t
Xbit_r11_c244 bl[244] br[244] wl[11] vdd gnd cell_6t
Xbit_r12_c244 bl[244] br[244] wl[12] vdd gnd cell_6t
Xbit_r13_c244 bl[244] br[244] wl[13] vdd gnd cell_6t
Xbit_r14_c244 bl[244] br[244] wl[14] vdd gnd cell_6t
Xbit_r15_c244 bl[244] br[244] wl[15] vdd gnd cell_6t
Xbit_r16_c244 bl[244] br[244] wl[16] vdd gnd cell_6t
Xbit_r17_c244 bl[244] br[244] wl[17] vdd gnd cell_6t
Xbit_r18_c244 bl[244] br[244] wl[18] vdd gnd cell_6t
Xbit_r19_c244 bl[244] br[244] wl[19] vdd gnd cell_6t
Xbit_r20_c244 bl[244] br[244] wl[20] vdd gnd cell_6t
Xbit_r21_c244 bl[244] br[244] wl[21] vdd gnd cell_6t
Xbit_r22_c244 bl[244] br[244] wl[22] vdd gnd cell_6t
Xbit_r23_c244 bl[244] br[244] wl[23] vdd gnd cell_6t
Xbit_r24_c244 bl[244] br[244] wl[24] vdd gnd cell_6t
Xbit_r25_c244 bl[244] br[244] wl[25] vdd gnd cell_6t
Xbit_r26_c244 bl[244] br[244] wl[26] vdd gnd cell_6t
Xbit_r27_c244 bl[244] br[244] wl[27] vdd gnd cell_6t
Xbit_r28_c244 bl[244] br[244] wl[28] vdd gnd cell_6t
Xbit_r29_c244 bl[244] br[244] wl[29] vdd gnd cell_6t
Xbit_r30_c244 bl[244] br[244] wl[30] vdd gnd cell_6t
Xbit_r31_c244 bl[244] br[244] wl[31] vdd gnd cell_6t
Xbit_r32_c244 bl[244] br[244] wl[32] vdd gnd cell_6t
Xbit_r33_c244 bl[244] br[244] wl[33] vdd gnd cell_6t
Xbit_r34_c244 bl[244] br[244] wl[34] vdd gnd cell_6t
Xbit_r35_c244 bl[244] br[244] wl[35] vdd gnd cell_6t
Xbit_r36_c244 bl[244] br[244] wl[36] vdd gnd cell_6t
Xbit_r37_c244 bl[244] br[244] wl[37] vdd gnd cell_6t
Xbit_r38_c244 bl[244] br[244] wl[38] vdd gnd cell_6t
Xbit_r39_c244 bl[244] br[244] wl[39] vdd gnd cell_6t
Xbit_r40_c244 bl[244] br[244] wl[40] vdd gnd cell_6t
Xbit_r41_c244 bl[244] br[244] wl[41] vdd gnd cell_6t
Xbit_r42_c244 bl[244] br[244] wl[42] vdd gnd cell_6t
Xbit_r43_c244 bl[244] br[244] wl[43] vdd gnd cell_6t
Xbit_r44_c244 bl[244] br[244] wl[44] vdd gnd cell_6t
Xbit_r45_c244 bl[244] br[244] wl[45] vdd gnd cell_6t
Xbit_r46_c244 bl[244] br[244] wl[46] vdd gnd cell_6t
Xbit_r47_c244 bl[244] br[244] wl[47] vdd gnd cell_6t
Xbit_r48_c244 bl[244] br[244] wl[48] vdd gnd cell_6t
Xbit_r49_c244 bl[244] br[244] wl[49] vdd gnd cell_6t
Xbit_r50_c244 bl[244] br[244] wl[50] vdd gnd cell_6t
Xbit_r51_c244 bl[244] br[244] wl[51] vdd gnd cell_6t
Xbit_r52_c244 bl[244] br[244] wl[52] vdd gnd cell_6t
Xbit_r53_c244 bl[244] br[244] wl[53] vdd gnd cell_6t
Xbit_r54_c244 bl[244] br[244] wl[54] vdd gnd cell_6t
Xbit_r55_c244 bl[244] br[244] wl[55] vdd gnd cell_6t
Xbit_r56_c244 bl[244] br[244] wl[56] vdd gnd cell_6t
Xbit_r57_c244 bl[244] br[244] wl[57] vdd gnd cell_6t
Xbit_r58_c244 bl[244] br[244] wl[58] vdd gnd cell_6t
Xbit_r59_c244 bl[244] br[244] wl[59] vdd gnd cell_6t
Xbit_r60_c244 bl[244] br[244] wl[60] vdd gnd cell_6t
Xbit_r61_c244 bl[244] br[244] wl[61] vdd gnd cell_6t
Xbit_r62_c244 bl[244] br[244] wl[62] vdd gnd cell_6t
Xbit_r63_c244 bl[244] br[244] wl[63] vdd gnd cell_6t
Xbit_r64_c244 bl[244] br[244] wl[64] vdd gnd cell_6t
Xbit_r65_c244 bl[244] br[244] wl[65] vdd gnd cell_6t
Xbit_r66_c244 bl[244] br[244] wl[66] vdd gnd cell_6t
Xbit_r67_c244 bl[244] br[244] wl[67] vdd gnd cell_6t
Xbit_r68_c244 bl[244] br[244] wl[68] vdd gnd cell_6t
Xbit_r69_c244 bl[244] br[244] wl[69] vdd gnd cell_6t
Xbit_r70_c244 bl[244] br[244] wl[70] vdd gnd cell_6t
Xbit_r71_c244 bl[244] br[244] wl[71] vdd gnd cell_6t
Xbit_r72_c244 bl[244] br[244] wl[72] vdd gnd cell_6t
Xbit_r73_c244 bl[244] br[244] wl[73] vdd gnd cell_6t
Xbit_r74_c244 bl[244] br[244] wl[74] vdd gnd cell_6t
Xbit_r75_c244 bl[244] br[244] wl[75] vdd gnd cell_6t
Xbit_r76_c244 bl[244] br[244] wl[76] vdd gnd cell_6t
Xbit_r77_c244 bl[244] br[244] wl[77] vdd gnd cell_6t
Xbit_r78_c244 bl[244] br[244] wl[78] vdd gnd cell_6t
Xbit_r79_c244 bl[244] br[244] wl[79] vdd gnd cell_6t
Xbit_r80_c244 bl[244] br[244] wl[80] vdd gnd cell_6t
Xbit_r81_c244 bl[244] br[244] wl[81] vdd gnd cell_6t
Xbit_r82_c244 bl[244] br[244] wl[82] vdd gnd cell_6t
Xbit_r83_c244 bl[244] br[244] wl[83] vdd gnd cell_6t
Xbit_r84_c244 bl[244] br[244] wl[84] vdd gnd cell_6t
Xbit_r85_c244 bl[244] br[244] wl[85] vdd gnd cell_6t
Xbit_r86_c244 bl[244] br[244] wl[86] vdd gnd cell_6t
Xbit_r87_c244 bl[244] br[244] wl[87] vdd gnd cell_6t
Xbit_r88_c244 bl[244] br[244] wl[88] vdd gnd cell_6t
Xbit_r89_c244 bl[244] br[244] wl[89] vdd gnd cell_6t
Xbit_r90_c244 bl[244] br[244] wl[90] vdd gnd cell_6t
Xbit_r91_c244 bl[244] br[244] wl[91] vdd gnd cell_6t
Xbit_r92_c244 bl[244] br[244] wl[92] vdd gnd cell_6t
Xbit_r93_c244 bl[244] br[244] wl[93] vdd gnd cell_6t
Xbit_r94_c244 bl[244] br[244] wl[94] vdd gnd cell_6t
Xbit_r95_c244 bl[244] br[244] wl[95] vdd gnd cell_6t
Xbit_r96_c244 bl[244] br[244] wl[96] vdd gnd cell_6t
Xbit_r97_c244 bl[244] br[244] wl[97] vdd gnd cell_6t
Xbit_r98_c244 bl[244] br[244] wl[98] vdd gnd cell_6t
Xbit_r99_c244 bl[244] br[244] wl[99] vdd gnd cell_6t
Xbit_r100_c244 bl[244] br[244] wl[100] vdd gnd cell_6t
Xbit_r101_c244 bl[244] br[244] wl[101] vdd gnd cell_6t
Xbit_r102_c244 bl[244] br[244] wl[102] vdd gnd cell_6t
Xbit_r103_c244 bl[244] br[244] wl[103] vdd gnd cell_6t
Xbit_r104_c244 bl[244] br[244] wl[104] vdd gnd cell_6t
Xbit_r105_c244 bl[244] br[244] wl[105] vdd gnd cell_6t
Xbit_r106_c244 bl[244] br[244] wl[106] vdd gnd cell_6t
Xbit_r107_c244 bl[244] br[244] wl[107] vdd gnd cell_6t
Xbit_r108_c244 bl[244] br[244] wl[108] vdd gnd cell_6t
Xbit_r109_c244 bl[244] br[244] wl[109] vdd gnd cell_6t
Xbit_r110_c244 bl[244] br[244] wl[110] vdd gnd cell_6t
Xbit_r111_c244 bl[244] br[244] wl[111] vdd gnd cell_6t
Xbit_r112_c244 bl[244] br[244] wl[112] vdd gnd cell_6t
Xbit_r113_c244 bl[244] br[244] wl[113] vdd gnd cell_6t
Xbit_r114_c244 bl[244] br[244] wl[114] vdd gnd cell_6t
Xbit_r115_c244 bl[244] br[244] wl[115] vdd gnd cell_6t
Xbit_r116_c244 bl[244] br[244] wl[116] vdd gnd cell_6t
Xbit_r117_c244 bl[244] br[244] wl[117] vdd gnd cell_6t
Xbit_r118_c244 bl[244] br[244] wl[118] vdd gnd cell_6t
Xbit_r119_c244 bl[244] br[244] wl[119] vdd gnd cell_6t
Xbit_r120_c244 bl[244] br[244] wl[120] vdd gnd cell_6t
Xbit_r121_c244 bl[244] br[244] wl[121] vdd gnd cell_6t
Xbit_r122_c244 bl[244] br[244] wl[122] vdd gnd cell_6t
Xbit_r123_c244 bl[244] br[244] wl[123] vdd gnd cell_6t
Xbit_r124_c244 bl[244] br[244] wl[124] vdd gnd cell_6t
Xbit_r125_c244 bl[244] br[244] wl[125] vdd gnd cell_6t
Xbit_r126_c244 bl[244] br[244] wl[126] vdd gnd cell_6t
Xbit_r127_c244 bl[244] br[244] wl[127] vdd gnd cell_6t
Xbit_r128_c244 bl[244] br[244] wl[128] vdd gnd cell_6t
Xbit_r129_c244 bl[244] br[244] wl[129] vdd gnd cell_6t
Xbit_r130_c244 bl[244] br[244] wl[130] vdd gnd cell_6t
Xbit_r131_c244 bl[244] br[244] wl[131] vdd gnd cell_6t
Xbit_r132_c244 bl[244] br[244] wl[132] vdd gnd cell_6t
Xbit_r133_c244 bl[244] br[244] wl[133] vdd gnd cell_6t
Xbit_r134_c244 bl[244] br[244] wl[134] vdd gnd cell_6t
Xbit_r135_c244 bl[244] br[244] wl[135] vdd gnd cell_6t
Xbit_r136_c244 bl[244] br[244] wl[136] vdd gnd cell_6t
Xbit_r137_c244 bl[244] br[244] wl[137] vdd gnd cell_6t
Xbit_r138_c244 bl[244] br[244] wl[138] vdd gnd cell_6t
Xbit_r139_c244 bl[244] br[244] wl[139] vdd gnd cell_6t
Xbit_r140_c244 bl[244] br[244] wl[140] vdd gnd cell_6t
Xbit_r141_c244 bl[244] br[244] wl[141] vdd gnd cell_6t
Xbit_r142_c244 bl[244] br[244] wl[142] vdd gnd cell_6t
Xbit_r143_c244 bl[244] br[244] wl[143] vdd gnd cell_6t
Xbit_r144_c244 bl[244] br[244] wl[144] vdd gnd cell_6t
Xbit_r145_c244 bl[244] br[244] wl[145] vdd gnd cell_6t
Xbit_r146_c244 bl[244] br[244] wl[146] vdd gnd cell_6t
Xbit_r147_c244 bl[244] br[244] wl[147] vdd gnd cell_6t
Xbit_r148_c244 bl[244] br[244] wl[148] vdd gnd cell_6t
Xbit_r149_c244 bl[244] br[244] wl[149] vdd gnd cell_6t
Xbit_r150_c244 bl[244] br[244] wl[150] vdd gnd cell_6t
Xbit_r151_c244 bl[244] br[244] wl[151] vdd gnd cell_6t
Xbit_r152_c244 bl[244] br[244] wl[152] vdd gnd cell_6t
Xbit_r153_c244 bl[244] br[244] wl[153] vdd gnd cell_6t
Xbit_r154_c244 bl[244] br[244] wl[154] vdd gnd cell_6t
Xbit_r155_c244 bl[244] br[244] wl[155] vdd gnd cell_6t
Xbit_r156_c244 bl[244] br[244] wl[156] vdd gnd cell_6t
Xbit_r157_c244 bl[244] br[244] wl[157] vdd gnd cell_6t
Xbit_r158_c244 bl[244] br[244] wl[158] vdd gnd cell_6t
Xbit_r159_c244 bl[244] br[244] wl[159] vdd gnd cell_6t
Xbit_r160_c244 bl[244] br[244] wl[160] vdd gnd cell_6t
Xbit_r161_c244 bl[244] br[244] wl[161] vdd gnd cell_6t
Xbit_r162_c244 bl[244] br[244] wl[162] vdd gnd cell_6t
Xbit_r163_c244 bl[244] br[244] wl[163] vdd gnd cell_6t
Xbit_r164_c244 bl[244] br[244] wl[164] vdd gnd cell_6t
Xbit_r165_c244 bl[244] br[244] wl[165] vdd gnd cell_6t
Xbit_r166_c244 bl[244] br[244] wl[166] vdd gnd cell_6t
Xbit_r167_c244 bl[244] br[244] wl[167] vdd gnd cell_6t
Xbit_r168_c244 bl[244] br[244] wl[168] vdd gnd cell_6t
Xbit_r169_c244 bl[244] br[244] wl[169] vdd gnd cell_6t
Xbit_r170_c244 bl[244] br[244] wl[170] vdd gnd cell_6t
Xbit_r171_c244 bl[244] br[244] wl[171] vdd gnd cell_6t
Xbit_r172_c244 bl[244] br[244] wl[172] vdd gnd cell_6t
Xbit_r173_c244 bl[244] br[244] wl[173] vdd gnd cell_6t
Xbit_r174_c244 bl[244] br[244] wl[174] vdd gnd cell_6t
Xbit_r175_c244 bl[244] br[244] wl[175] vdd gnd cell_6t
Xbit_r176_c244 bl[244] br[244] wl[176] vdd gnd cell_6t
Xbit_r177_c244 bl[244] br[244] wl[177] vdd gnd cell_6t
Xbit_r178_c244 bl[244] br[244] wl[178] vdd gnd cell_6t
Xbit_r179_c244 bl[244] br[244] wl[179] vdd gnd cell_6t
Xbit_r180_c244 bl[244] br[244] wl[180] vdd gnd cell_6t
Xbit_r181_c244 bl[244] br[244] wl[181] vdd gnd cell_6t
Xbit_r182_c244 bl[244] br[244] wl[182] vdd gnd cell_6t
Xbit_r183_c244 bl[244] br[244] wl[183] vdd gnd cell_6t
Xbit_r184_c244 bl[244] br[244] wl[184] vdd gnd cell_6t
Xbit_r185_c244 bl[244] br[244] wl[185] vdd gnd cell_6t
Xbit_r186_c244 bl[244] br[244] wl[186] vdd gnd cell_6t
Xbit_r187_c244 bl[244] br[244] wl[187] vdd gnd cell_6t
Xbit_r188_c244 bl[244] br[244] wl[188] vdd gnd cell_6t
Xbit_r189_c244 bl[244] br[244] wl[189] vdd gnd cell_6t
Xbit_r190_c244 bl[244] br[244] wl[190] vdd gnd cell_6t
Xbit_r191_c244 bl[244] br[244] wl[191] vdd gnd cell_6t
Xbit_r192_c244 bl[244] br[244] wl[192] vdd gnd cell_6t
Xbit_r193_c244 bl[244] br[244] wl[193] vdd gnd cell_6t
Xbit_r194_c244 bl[244] br[244] wl[194] vdd gnd cell_6t
Xbit_r195_c244 bl[244] br[244] wl[195] vdd gnd cell_6t
Xbit_r196_c244 bl[244] br[244] wl[196] vdd gnd cell_6t
Xbit_r197_c244 bl[244] br[244] wl[197] vdd gnd cell_6t
Xbit_r198_c244 bl[244] br[244] wl[198] vdd gnd cell_6t
Xbit_r199_c244 bl[244] br[244] wl[199] vdd gnd cell_6t
Xbit_r200_c244 bl[244] br[244] wl[200] vdd gnd cell_6t
Xbit_r201_c244 bl[244] br[244] wl[201] vdd gnd cell_6t
Xbit_r202_c244 bl[244] br[244] wl[202] vdd gnd cell_6t
Xbit_r203_c244 bl[244] br[244] wl[203] vdd gnd cell_6t
Xbit_r204_c244 bl[244] br[244] wl[204] vdd gnd cell_6t
Xbit_r205_c244 bl[244] br[244] wl[205] vdd gnd cell_6t
Xbit_r206_c244 bl[244] br[244] wl[206] vdd gnd cell_6t
Xbit_r207_c244 bl[244] br[244] wl[207] vdd gnd cell_6t
Xbit_r208_c244 bl[244] br[244] wl[208] vdd gnd cell_6t
Xbit_r209_c244 bl[244] br[244] wl[209] vdd gnd cell_6t
Xbit_r210_c244 bl[244] br[244] wl[210] vdd gnd cell_6t
Xbit_r211_c244 bl[244] br[244] wl[211] vdd gnd cell_6t
Xbit_r212_c244 bl[244] br[244] wl[212] vdd gnd cell_6t
Xbit_r213_c244 bl[244] br[244] wl[213] vdd gnd cell_6t
Xbit_r214_c244 bl[244] br[244] wl[214] vdd gnd cell_6t
Xbit_r215_c244 bl[244] br[244] wl[215] vdd gnd cell_6t
Xbit_r216_c244 bl[244] br[244] wl[216] vdd gnd cell_6t
Xbit_r217_c244 bl[244] br[244] wl[217] vdd gnd cell_6t
Xbit_r218_c244 bl[244] br[244] wl[218] vdd gnd cell_6t
Xbit_r219_c244 bl[244] br[244] wl[219] vdd gnd cell_6t
Xbit_r220_c244 bl[244] br[244] wl[220] vdd gnd cell_6t
Xbit_r221_c244 bl[244] br[244] wl[221] vdd gnd cell_6t
Xbit_r222_c244 bl[244] br[244] wl[222] vdd gnd cell_6t
Xbit_r223_c244 bl[244] br[244] wl[223] vdd gnd cell_6t
Xbit_r224_c244 bl[244] br[244] wl[224] vdd gnd cell_6t
Xbit_r225_c244 bl[244] br[244] wl[225] vdd gnd cell_6t
Xbit_r226_c244 bl[244] br[244] wl[226] vdd gnd cell_6t
Xbit_r227_c244 bl[244] br[244] wl[227] vdd gnd cell_6t
Xbit_r228_c244 bl[244] br[244] wl[228] vdd gnd cell_6t
Xbit_r229_c244 bl[244] br[244] wl[229] vdd gnd cell_6t
Xbit_r230_c244 bl[244] br[244] wl[230] vdd gnd cell_6t
Xbit_r231_c244 bl[244] br[244] wl[231] vdd gnd cell_6t
Xbit_r232_c244 bl[244] br[244] wl[232] vdd gnd cell_6t
Xbit_r233_c244 bl[244] br[244] wl[233] vdd gnd cell_6t
Xbit_r234_c244 bl[244] br[244] wl[234] vdd gnd cell_6t
Xbit_r235_c244 bl[244] br[244] wl[235] vdd gnd cell_6t
Xbit_r236_c244 bl[244] br[244] wl[236] vdd gnd cell_6t
Xbit_r237_c244 bl[244] br[244] wl[237] vdd gnd cell_6t
Xbit_r238_c244 bl[244] br[244] wl[238] vdd gnd cell_6t
Xbit_r239_c244 bl[244] br[244] wl[239] vdd gnd cell_6t
Xbit_r240_c244 bl[244] br[244] wl[240] vdd gnd cell_6t
Xbit_r241_c244 bl[244] br[244] wl[241] vdd gnd cell_6t
Xbit_r242_c244 bl[244] br[244] wl[242] vdd gnd cell_6t
Xbit_r243_c244 bl[244] br[244] wl[243] vdd gnd cell_6t
Xbit_r244_c244 bl[244] br[244] wl[244] vdd gnd cell_6t
Xbit_r245_c244 bl[244] br[244] wl[245] vdd gnd cell_6t
Xbit_r246_c244 bl[244] br[244] wl[246] vdd gnd cell_6t
Xbit_r247_c244 bl[244] br[244] wl[247] vdd gnd cell_6t
Xbit_r248_c244 bl[244] br[244] wl[248] vdd gnd cell_6t
Xbit_r249_c244 bl[244] br[244] wl[249] vdd gnd cell_6t
Xbit_r250_c244 bl[244] br[244] wl[250] vdd gnd cell_6t
Xbit_r251_c244 bl[244] br[244] wl[251] vdd gnd cell_6t
Xbit_r252_c244 bl[244] br[244] wl[252] vdd gnd cell_6t
Xbit_r253_c244 bl[244] br[244] wl[253] vdd gnd cell_6t
Xbit_r254_c244 bl[244] br[244] wl[254] vdd gnd cell_6t
Xbit_r255_c244 bl[244] br[244] wl[255] vdd gnd cell_6t
Xbit_r0_c245 bl[245] br[245] wl[0] vdd gnd cell_6t
Xbit_r1_c245 bl[245] br[245] wl[1] vdd gnd cell_6t
Xbit_r2_c245 bl[245] br[245] wl[2] vdd gnd cell_6t
Xbit_r3_c245 bl[245] br[245] wl[3] vdd gnd cell_6t
Xbit_r4_c245 bl[245] br[245] wl[4] vdd gnd cell_6t
Xbit_r5_c245 bl[245] br[245] wl[5] vdd gnd cell_6t
Xbit_r6_c245 bl[245] br[245] wl[6] vdd gnd cell_6t
Xbit_r7_c245 bl[245] br[245] wl[7] vdd gnd cell_6t
Xbit_r8_c245 bl[245] br[245] wl[8] vdd gnd cell_6t
Xbit_r9_c245 bl[245] br[245] wl[9] vdd gnd cell_6t
Xbit_r10_c245 bl[245] br[245] wl[10] vdd gnd cell_6t
Xbit_r11_c245 bl[245] br[245] wl[11] vdd gnd cell_6t
Xbit_r12_c245 bl[245] br[245] wl[12] vdd gnd cell_6t
Xbit_r13_c245 bl[245] br[245] wl[13] vdd gnd cell_6t
Xbit_r14_c245 bl[245] br[245] wl[14] vdd gnd cell_6t
Xbit_r15_c245 bl[245] br[245] wl[15] vdd gnd cell_6t
Xbit_r16_c245 bl[245] br[245] wl[16] vdd gnd cell_6t
Xbit_r17_c245 bl[245] br[245] wl[17] vdd gnd cell_6t
Xbit_r18_c245 bl[245] br[245] wl[18] vdd gnd cell_6t
Xbit_r19_c245 bl[245] br[245] wl[19] vdd gnd cell_6t
Xbit_r20_c245 bl[245] br[245] wl[20] vdd gnd cell_6t
Xbit_r21_c245 bl[245] br[245] wl[21] vdd gnd cell_6t
Xbit_r22_c245 bl[245] br[245] wl[22] vdd gnd cell_6t
Xbit_r23_c245 bl[245] br[245] wl[23] vdd gnd cell_6t
Xbit_r24_c245 bl[245] br[245] wl[24] vdd gnd cell_6t
Xbit_r25_c245 bl[245] br[245] wl[25] vdd gnd cell_6t
Xbit_r26_c245 bl[245] br[245] wl[26] vdd gnd cell_6t
Xbit_r27_c245 bl[245] br[245] wl[27] vdd gnd cell_6t
Xbit_r28_c245 bl[245] br[245] wl[28] vdd gnd cell_6t
Xbit_r29_c245 bl[245] br[245] wl[29] vdd gnd cell_6t
Xbit_r30_c245 bl[245] br[245] wl[30] vdd gnd cell_6t
Xbit_r31_c245 bl[245] br[245] wl[31] vdd gnd cell_6t
Xbit_r32_c245 bl[245] br[245] wl[32] vdd gnd cell_6t
Xbit_r33_c245 bl[245] br[245] wl[33] vdd gnd cell_6t
Xbit_r34_c245 bl[245] br[245] wl[34] vdd gnd cell_6t
Xbit_r35_c245 bl[245] br[245] wl[35] vdd gnd cell_6t
Xbit_r36_c245 bl[245] br[245] wl[36] vdd gnd cell_6t
Xbit_r37_c245 bl[245] br[245] wl[37] vdd gnd cell_6t
Xbit_r38_c245 bl[245] br[245] wl[38] vdd gnd cell_6t
Xbit_r39_c245 bl[245] br[245] wl[39] vdd gnd cell_6t
Xbit_r40_c245 bl[245] br[245] wl[40] vdd gnd cell_6t
Xbit_r41_c245 bl[245] br[245] wl[41] vdd gnd cell_6t
Xbit_r42_c245 bl[245] br[245] wl[42] vdd gnd cell_6t
Xbit_r43_c245 bl[245] br[245] wl[43] vdd gnd cell_6t
Xbit_r44_c245 bl[245] br[245] wl[44] vdd gnd cell_6t
Xbit_r45_c245 bl[245] br[245] wl[45] vdd gnd cell_6t
Xbit_r46_c245 bl[245] br[245] wl[46] vdd gnd cell_6t
Xbit_r47_c245 bl[245] br[245] wl[47] vdd gnd cell_6t
Xbit_r48_c245 bl[245] br[245] wl[48] vdd gnd cell_6t
Xbit_r49_c245 bl[245] br[245] wl[49] vdd gnd cell_6t
Xbit_r50_c245 bl[245] br[245] wl[50] vdd gnd cell_6t
Xbit_r51_c245 bl[245] br[245] wl[51] vdd gnd cell_6t
Xbit_r52_c245 bl[245] br[245] wl[52] vdd gnd cell_6t
Xbit_r53_c245 bl[245] br[245] wl[53] vdd gnd cell_6t
Xbit_r54_c245 bl[245] br[245] wl[54] vdd gnd cell_6t
Xbit_r55_c245 bl[245] br[245] wl[55] vdd gnd cell_6t
Xbit_r56_c245 bl[245] br[245] wl[56] vdd gnd cell_6t
Xbit_r57_c245 bl[245] br[245] wl[57] vdd gnd cell_6t
Xbit_r58_c245 bl[245] br[245] wl[58] vdd gnd cell_6t
Xbit_r59_c245 bl[245] br[245] wl[59] vdd gnd cell_6t
Xbit_r60_c245 bl[245] br[245] wl[60] vdd gnd cell_6t
Xbit_r61_c245 bl[245] br[245] wl[61] vdd gnd cell_6t
Xbit_r62_c245 bl[245] br[245] wl[62] vdd gnd cell_6t
Xbit_r63_c245 bl[245] br[245] wl[63] vdd gnd cell_6t
Xbit_r64_c245 bl[245] br[245] wl[64] vdd gnd cell_6t
Xbit_r65_c245 bl[245] br[245] wl[65] vdd gnd cell_6t
Xbit_r66_c245 bl[245] br[245] wl[66] vdd gnd cell_6t
Xbit_r67_c245 bl[245] br[245] wl[67] vdd gnd cell_6t
Xbit_r68_c245 bl[245] br[245] wl[68] vdd gnd cell_6t
Xbit_r69_c245 bl[245] br[245] wl[69] vdd gnd cell_6t
Xbit_r70_c245 bl[245] br[245] wl[70] vdd gnd cell_6t
Xbit_r71_c245 bl[245] br[245] wl[71] vdd gnd cell_6t
Xbit_r72_c245 bl[245] br[245] wl[72] vdd gnd cell_6t
Xbit_r73_c245 bl[245] br[245] wl[73] vdd gnd cell_6t
Xbit_r74_c245 bl[245] br[245] wl[74] vdd gnd cell_6t
Xbit_r75_c245 bl[245] br[245] wl[75] vdd gnd cell_6t
Xbit_r76_c245 bl[245] br[245] wl[76] vdd gnd cell_6t
Xbit_r77_c245 bl[245] br[245] wl[77] vdd gnd cell_6t
Xbit_r78_c245 bl[245] br[245] wl[78] vdd gnd cell_6t
Xbit_r79_c245 bl[245] br[245] wl[79] vdd gnd cell_6t
Xbit_r80_c245 bl[245] br[245] wl[80] vdd gnd cell_6t
Xbit_r81_c245 bl[245] br[245] wl[81] vdd gnd cell_6t
Xbit_r82_c245 bl[245] br[245] wl[82] vdd gnd cell_6t
Xbit_r83_c245 bl[245] br[245] wl[83] vdd gnd cell_6t
Xbit_r84_c245 bl[245] br[245] wl[84] vdd gnd cell_6t
Xbit_r85_c245 bl[245] br[245] wl[85] vdd gnd cell_6t
Xbit_r86_c245 bl[245] br[245] wl[86] vdd gnd cell_6t
Xbit_r87_c245 bl[245] br[245] wl[87] vdd gnd cell_6t
Xbit_r88_c245 bl[245] br[245] wl[88] vdd gnd cell_6t
Xbit_r89_c245 bl[245] br[245] wl[89] vdd gnd cell_6t
Xbit_r90_c245 bl[245] br[245] wl[90] vdd gnd cell_6t
Xbit_r91_c245 bl[245] br[245] wl[91] vdd gnd cell_6t
Xbit_r92_c245 bl[245] br[245] wl[92] vdd gnd cell_6t
Xbit_r93_c245 bl[245] br[245] wl[93] vdd gnd cell_6t
Xbit_r94_c245 bl[245] br[245] wl[94] vdd gnd cell_6t
Xbit_r95_c245 bl[245] br[245] wl[95] vdd gnd cell_6t
Xbit_r96_c245 bl[245] br[245] wl[96] vdd gnd cell_6t
Xbit_r97_c245 bl[245] br[245] wl[97] vdd gnd cell_6t
Xbit_r98_c245 bl[245] br[245] wl[98] vdd gnd cell_6t
Xbit_r99_c245 bl[245] br[245] wl[99] vdd gnd cell_6t
Xbit_r100_c245 bl[245] br[245] wl[100] vdd gnd cell_6t
Xbit_r101_c245 bl[245] br[245] wl[101] vdd gnd cell_6t
Xbit_r102_c245 bl[245] br[245] wl[102] vdd gnd cell_6t
Xbit_r103_c245 bl[245] br[245] wl[103] vdd gnd cell_6t
Xbit_r104_c245 bl[245] br[245] wl[104] vdd gnd cell_6t
Xbit_r105_c245 bl[245] br[245] wl[105] vdd gnd cell_6t
Xbit_r106_c245 bl[245] br[245] wl[106] vdd gnd cell_6t
Xbit_r107_c245 bl[245] br[245] wl[107] vdd gnd cell_6t
Xbit_r108_c245 bl[245] br[245] wl[108] vdd gnd cell_6t
Xbit_r109_c245 bl[245] br[245] wl[109] vdd gnd cell_6t
Xbit_r110_c245 bl[245] br[245] wl[110] vdd gnd cell_6t
Xbit_r111_c245 bl[245] br[245] wl[111] vdd gnd cell_6t
Xbit_r112_c245 bl[245] br[245] wl[112] vdd gnd cell_6t
Xbit_r113_c245 bl[245] br[245] wl[113] vdd gnd cell_6t
Xbit_r114_c245 bl[245] br[245] wl[114] vdd gnd cell_6t
Xbit_r115_c245 bl[245] br[245] wl[115] vdd gnd cell_6t
Xbit_r116_c245 bl[245] br[245] wl[116] vdd gnd cell_6t
Xbit_r117_c245 bl[245] br[245] wl[117] vdd gnd cell_6t
Xbit_r118_c245 bl[245] br[245] wl[118] vdd gnd cell_6t
Xbit_r119_c245 bl[245] br[245] wl[119] vdd gnd cell_6t
Xbit_r120_c245 bl[245] br[245] wl[120] vdd gnd cell_6t
Xbit_r121_c245 bl[245] br[245] wl[121] vdd gnd cell_6t
Xbit_r122_c245 bl[245] br[245] wl[122] vdd gnd cell_6t
Xbit_r123_c245 bl[245] br[245] wl[123] vdd gnd cell_6t
Xbit_r124_c245 bl[245] br[245] wl[124] vdd gnd cell_6t
Xbit_r125_c245 bl[245] br[245] wl[125] vdd gnd cell_6t
Xbit_r126_c245 bl[245] br[245] wl[126] vdd gnd cell_6t
Xbit_r127_c245 bl[245] br[245] wl[127] vdd gnd cell_6t
Xbit_r128_c245 bl[245] br[245] wl[128] vdd gnd cell_6t
Xbit_r129_c245 bl[245] br[245] wl[129] vdd gnd cell_6t
Xbit_r130_c245 bl[245] br[245] wl[130] vdd gnd cell_6t
Xbit_r131_c245 bl[245] br[245] wl[131] vdd gnd cell_6t
Xbit_r132_c245 bl[245] br[245] wl[132] vdd gnd cell_6t
Xbit_r133_c245 bl[245] br[245] wl[133] vdd gnd cell_6t
Xbit_r134_c245 bl[245] br[245] wl[134] vdd gnd cell_6t
Xbit_r135_c245 bl[245] br[245] wl[135] vdd gnd cell_6t
Xbit_r136_c245 bl[245] br[245] wl[136] vdd gnd cell_6t
Xbit_r137_c245 bl[245] br[245] wl[137] vdd gnd cell_6t
Xbit_r138_c245 bl[245] br[245] wl[138] vdd gnd cell_6t
Xbit_r139_c245 bl[245] br[245] wl[139] vdd gnd cell_6t
Xbit_r140_c245 bl[245] br[245] wl[140] vdd gnd cell_6t
Xbit_r141_c245 bl[245] br[245] wl[141] vdd gnd cell_6t
Xbit_r142_c245 bl[245] br[245] wl[142] vdd gnd cell_6t
Xbit_r143_c245 bl[245] br[245] wl[143] vdd gnd cell_6t
Xbit_r144_c245 bl[245] br[245] wl[144] vdd gnd cell_6t
Xbit_r145_c245 bl[245] br[245] wl[145] vdd gnd cell_6t
Xbit_r146_c245 bl[245] br[245] wl[146] vdd gnd cell_6t
Xbit_r147_c245 bl[245] br[245] wl[147] vdd gnd cell_6t
Xbit_r148_c245 bl[245] br[245] wl[148] vdd gnd cell_6t
Xbit_r149_c245 bl[245] br[245] wl[149] vdd gnd cell_6t
Xbit_r150_c245 bl[245] br[245] wl[150] vdd gnd cell_6t
Xbit_r151_c245 bl[245] br[245] wl[151] vdd gnd cell_6t
Xbit_r152_c245 bl[245] br[245] wl[152] vdd gnd cell_6t
Xbit_r153_c245 bl[245] br[245] wl[153] vdd gnd cell_6t
Xbit_r154_c245 bl[245] br[245] wl[154] vdd gnd cell_6t
Xbit_r155_c245 bl[245] br[245] wl[155] vdd gnd cell_6t
Xbit_r156_c245 bl[245] br[245] wl[156] vdd gnd cell_6t
Xbit_r157_c245 bl[245] br[245] wl[157] vdd gnd cell_6t
Xbit_r158_c245 bl[245] br[245] wl[158] vdd gnd cell_6t
Xbit_r159_c245 bl[245] br[245] wl[159] vdd gnd cell_6t
Xbit_r160_c245 bl[245] br[245] wl[160] vdd gnd cell_6t
Xbit_r161_c245 bl[245] br[245] wl[161] vdd gnd cell_6t
Xbit_r162_c245 bl[245] br[245] wl[162] vdd gnd cell_6t
Xbit_r163_c245 bl[245] br[245] wl[163] vdd gnd cell_6t
Xbit_r164_c245 bl[245] br[245] wl[164] vdd gnd cell_6t
Xbit_r165_c245 bl[245] br[245] wl[165] vdd gnd cell_6t
Xbit_r166_c245 bl[245] br[245] wl[166] vdd gnd cell_6t
Xbit_r167_c245 bl[245] br[245] wl[167] vdd gnd cell_6t
Xbit_r168_c245 bl[245] br[245] wl[168] vdd gnd cell_6t
Xbit_r169_c245 bl[245] br[245] wl[169] vdd gnd cell_6t
Xbit_r170_c245 bl[245] br[245] wl[170] vdd gnd cell_6t
Xbit_r171_c245 bl[245] br[245] wl[171] vdd gnd cell_6t
Xbit_r172_c245 bl[245] br[245] wl[172] vdd gnd cell_6t
Xbit_r173_c245 bl[245] br[245] wl[173] vdd gnd cell_6t
Xbit_r174_c245 bl[245] br[245] wl[174] vdd gnd cell_6t
Xbit_r175_c245 bl[245] br[245] wl[175] vdd gnd cell_6t
Xbit_r176_c245 bl[245] br[245] wl[176] vdd gnd cell_6t
Xbit_r177_c245 bl[245] br[245] wl[177] vdd gnd cell_6t
Xbit_r178_c245 bl[245] br[245] wl[178] vdd gnd cell_6t
Xbit_r179_c245 bl[245] br[245] wl[179] vdd gnd cell_6t
Xbit_r180_c245 bl[245] br[245] wl[180] vdd gnd cell_6t
Xbit_r181_c245 bl[245] br[245] wl[181] vdd gnd cell_6t
Xbit_r182_c245 bl[245] br[245] wl[182] vdd gnd cell_6t
Xbit_r183_c245 bl[245] br[245] wl[183] vdd gnd cell_6t
Xbit_r184_c245 bl[245] br[245] wl[184] vdd gnd cell_6t
Xbit_r185_c245 bl[245] br[245] wl[185] vdd gnd cell_6t
Xbit_r186_c245 bl[245] br[245] wl[186] vdd gnd cell_6t
Xbit_r187_c245 bl[245] br[245] wl[187] vdd gnd cell_6t
Xbit_r188_c245 bl[245] br[245] wl[188] vdd gnd cell_6t
Xbit_r189_c245 bl[245] br[245] wl[189] vdd gnd cell_6t
Xbit_r190_c245 bl[245] br[245] wl[190] vdd gnd cell_6t
Xbit_r191_c245 bl[245] br[245] wl[191] vdd gnd cell_6t
Xbit_r192_c245 bl[245] br[245] wl[192] vdd gnd cell_6t
Xbit_r193_c245 bl[245] br[245] wl[193] vdd gnd cell_6t
Xbit_r194_c245 bl[245] br[245] wl[194] vdd gnd cell_6t
Xbit_r195_c245 bl[245] br[245] wl[195] vdd gnd cell_6t
Xbit_r196_c245 bl[245] br[245] wl[196] vdd gnd cell_6t
Xbit_r197_c245 bl[245] br[245] wl[197] vdd gnd cell_6t
Xbit_r198_c245 bl[245] br[245] wl[198] vdd gnd cell_6t
Xbit_r199_c245 bl[245] br[245] wl[199] vdd gnd cell_6t
Xbit_r200_c245 bl[245] br[245] wl[200] vdd gnd cell_6t
Xbit_r201_c245 bl[245] br[245] wl[201] vdd gnd cell_6t
Xbit_r202_c245 bl[245] br[245] wl[202] vdd gnd cell_6t
Xbit_r203_c245 bl[245] br[245] wl[203] vdd gnd cell_6t
Xbit_r204_c245 bl[245] br[245] wl[204] vdd gnd cell_6t
Xbit_r205_c245 bl[245] br[245] wl[205] vdd gnd cell_6t
Xbit_r206_c245 bl[245] br[245] wl[206] vdd gnd cell_6t
Xbit_r207_c245 bl[245] br[245] wl[207] vdd gnd cell_6t
Xbit_r208_c245 bl[245] br[245] wl[208] vdd gnd cell_6t
Xbit_r209_c245 bl[245] br[245] wl[209] vdd gnd cell_6t
Xbit_r210_c245 bl[245] br[245] wl[210] vdd gnd cell_6t
Xbit_r211_c245 bl[245] br[245] wl[211] vdd gnd cell_6t
Xbit_r212_c245 bl[245] br[245] wl[212] vdd gnd cell_6t
Xbit_r213_c245 bl[245] br[245] wl[213] vdd gnd cell_6t
Xbit_r214_c245 bl[245] br[245] wl[214] vdd gnd cell_6t
Xbit_r215_c245 bl[245] br[245] wl[215] vdd gnd cell_6t
Xbit_r216_c245 bl[245] br[245] wl[216] vdd gnd cell_6t
Xbit_r217_c245 bl[245] br[245] wl[217] vdd gnd cell_6t
Xbit_r218_c245 bl[245] br[245] wl[218] vdd gnd cell_6t
Xbit_r219_c245 bl[245] br[245] wl[219] vdd gnd cell_6t
Xbit_r220_c245 bl[245] br[245] wl[220] vdd gnd cell_6t
Xbit_r221_c245 bl[245] br[245] wl[221] vdd gnd cell_6t
Xbit_r222_c245 bl[245] br[245] wl[222] vdd gnd cell_6t
Xbit_r223_c245 bl[245] br[245] wl[223] vdd gnd cell_6t
Xbit_r224_c245 bl[245] br[245] wl[224] vdd gnd cell_6t
Xbit_r225_c245 bl[245] br[245] wl[225] vdd gnd cell_6t
Xbit_r226_c245 bl[245] br[245] wl[226] vdd gnd cell_6t
Xbit_r227_c245 bl[245] br[245] wl[227] vdd gnd cell_6t
Xbit_r228_c245 bl[245] br[245] wl[228] vdd gnd cell_6t
Xbit_r229_c245 bl[245] br[245] wl[229] vdd gnd cell_6t
Xbit_r230_c245 bl[245] br[245] wl[230] vdd gnd cell_6t
Xbit_r231_c245 bl[245] br[245] wl[231] vdd gnd cell_6t
Xbit_r232_c245 bl[245] br[245] wl[232] vdd gnd cell_6t
Xbit_r233_c245 bl[245] br[245] wl[233] vdd gnd cell_6t
Xbit_r234_c245 bl[245] br[245] wl[234] vdd gnd cell_6t
Xbit_r235_c245 bl[245] br[245] wl[235] vdd gnd cell_6t
Xbit_r236_c245 bl[245] br[245] wl[236] vdd gnd cell_6t
Xbit_r237_c245 bl[245] br[245] wl[237] vdd gnd cell_6t
Xbit_r238_c245 bl[245] br[245] wl[238] vdd gnd cell_6t
Xbit_r239_c245 bl[245] br[245] wl[239] vdd gnd cell_6t
Xbit_r240_c245 bl[245] br[245] wl[240] vdd gnd cell_6t
Xbit_r241_c245 bl[245] br[245] wl[241] vdd gnd cell_6t
Xbit_r242_c245 bl[245] br[245] wl[242] vdd gnd cell_6t
Xbit_r243_c245 bl[245] br[245] wl[243] vdd gnd cell_6t
Xbit_r244_c245 bl[245] br[245] wl[244] vdd gnd cell_6t
Xbit_r245_c245 bl[245] br[245] wl[245] vdd gnd cell_6t
Xbit_r246_c245 bl[245] br[245] wl[246] vdd gnd cell_6t
Xbit_r247_c245 bl[245] br[245] wl[247] vdd gnd cell_6t
Xbit_r248_c245 bl[245] br[245] wl[248] vdd gnd cell_6t
Xbit_r249_c245 bl[245] br[245] wl[249] vdd gnd cell_6t
Xbit_r250_c245 bl[245] br[245] wl[250] vdd gnd cell_6t
Xbit_r251_c245 bl[245] br[245] wl[251] vdd gnd cell_6t
Xbit_r252_c245 bl[245] br[245] wl[252] vdd gnd cell_6t
Xbit_r253_c245 bl[245] br[245] wl[253] vdd gnd cell_6t
Xbit_r254_c245 bl[245] br[245] wl[254] vdd gnd cell_6t
Xbit_r255_c245 bl[245] br[245] wl[255] vdd gnd cell_6t
Xbit_r0_c246 bl[246] br[246] wl[0] vdd gnd cell_6t
Xbit_r1_c246 bl[246] br[246] wl[1] vdd gnd cell_6t
Xbit_r2_c246 bl[246] br[246] wl[2] vdd gnd cell_6t
Xbit_r3_c246 bl[246] br[246] wl[3] vdd gnd cell_6t
Xbit_r4_c246 bl[246] br[246] wl[4] vdd gnd cell_6t
Xbit_r5_c246 bl[246] br[246] wl[5] vdd gnd cell_6t
Xbit_r6_c246 bl[246] br[246] wl[6] vdd gnd cell_6t
Xbit_r7_c246 bl[246] br[246] wl[7] vdd gnd cell_6t
Xbit_r8_c246 bl[246] br[246] wl[8] vdd gnd cell_6t
Xbit_r9_c246 bl[246] br[246] wl[9] vdd gnd cell_6t
Xbit_r10_c246 bl[246] br[246] wl[10] vdd gnd cell_6t
Xbit_r11_c246 bl[246] br[246] wl[11] vdd gnd cell_6t
Xbit_r12_c246 bl[246] br[246] wl[12] vdd gnd cell_6t
Xbit_r13_c246 bl[246] br[246] wl[13] vdd gnd cell_6t
Xbit_r14_c246 bl[246] br[246] wl[14] vdd gnd cell_6t
Xbit_r15_c246 bl[246] br[246] wl[15] vdd gnd cell_6t
Xbit_r16_c246 bl[246] br[246] wl[16] vdd gnd cell_6t
Xbit_r17_c246 bl[246] br[246] wl[17] vdd gnd cell_6t
Xbit_r18_c246 bl[246] br[246] wl[18] vdd gnd cell_6t
Xbit_r19_c246 bl[246] br[246] wl[19] vdd gnd cell_6t
Xbit_r20_c246 bl[246] br[246] wl[20] vdd gnd cell_6t
Xbit_r21_c246 bl[246] br[246] wl[21] vdd gnd cell_6t
Xbit_r22_c246 bl[246] br[246] wl[22] vdd gnd cell_6t
Xbit_r23_c246 bl[246] br[246] wl[23] vdd gnd cell_6t
Xbit_r24_c246 bl[246] br[246] wl[24] vdd gnd cell_6t
Xbit_r25_c246 bl[246] br[246] wl[25] vdd gnd cell_6t
Xbit_r26_c246 bl[246] br[246] wl[26] vdd gnd cell_6t
Xbit_r27_c246 bl[246] br[246] wl[27] vdd gnd cell_6t
Xbit_r28_c246 bl[246] br[246] wl[28] vdd gnd cell_6t
Xbit_r29_c246 bl[246] br[246] wl[29] vdd gnd cell_6t
Xbit_r30_c246 bl[246] br[246] wl[30] vdd gnd cell_6t
Xbit_r31_c246 bl[246] br[246] wl[31] vdd gnd cell_6t
Xbit_r32_c246 bl[246] br[246] wl[32] vdd gnd cell_6t
Xbit_r33_c246 bl[246] br[246] wl[33] vdd gnd cell_6t
Xbit_r34_c246 bl[246] br[246] wl[34] vdd gnd cell_6t
Xbit_r35_c246 bl[246] br[246] wl[35] vdd gnd cell_6t
Xbit_r36_c246 bl[246] br[246] wl[36] vdd gnd cell_6t
Xbit_r37_c246 bl[246] br[246] wl[37] vdd gnd cell_6t
Xbit_r38_c246 bl[246] br[246] wl[38] vdd gnd cell_6t
Xbit_r39_c246 bl[246] br[246] wl[39] vdd gnd cell_6t
Xbit_r40_c246 bl[246] br[246] wl[40] vdd gnd cell_6t
Xbit_r41_c246 bl[246] br[246] wl[41] vdd gnd cell_6t
Xbit_r42_c246 bl[246] br[246] wl[42] vdd gnd cell_6t
Xbit_r43_c246 bl[246] br[246] wl[43] vdd gnd cell_6t
Xbit_r44_c246 bl[246] br[246] wl[44] vdd gnd cell_6t
Xbit_r45_c246 bl[246] br[246] wl[45] vdd gnd cell_6t
Xbit_r46_c246 bl[246] br[246] wl[46] vdd gnd cell_6t
Xbit_r47_c246 bl[246] br[246] wl[47] vdd gnd cell_6t
Xbit_r48_c246 bl[246] br[246] wl[48] vdd gnd cell_6t
Xbit_r49_c246 bl[246] br[246] wl[49] vdd gnd cell_6t
Xbit_r50_c246 bl[246] br[246] wl[50] vdd gnd cell_6t
Xbit_r51_c246 bl[246] br[246] wl[51] vdd gnd cell_6t
Xbit_r52_c246 bl[246] br[246] wl[52] vdd gnd cell_6t
Xbit_r53_c246 bl[246] br[246] wl[53] vdd gnd cell_6t
Xbit_r54_c246 bl[246] br[246] wl[54] vdd gnd cell_6t
Xbit_r55_c246 bl[246] br[246] wl[55] vdd gnd cell_6t
Xbit_r56_c246 bl[246] br[246] wl[56] vdd gnd cell_6t
Xbit_r57_c246 bl[246] br[246] wl[57] vdd gnd cell_6t
Xbit_r58_c246 bl[246] br[246] wl[58] vdd gnd cell_6t
Xbit_r59_c246 bl[246] br[246] wl[59] vdd gnd cell_6t
Xbit_r60_c246 bl[246] br[246] wl[60] vdd gnd cell_6t
Xbit_r61_c246 bl[246] br[246] wl[61] vdd gnd cell_6t
Xbit_r62_c246 bl[246] br[246] wl[62] vdd gnd cell_6t
Xbit_r63_c246 bl[246] br[246] wl[63] vdd gnd cell_6t
Xbit_r64_c246 bl[246] br[246] wl[64] vdd gnd cell_6t
Xbit_r65_c246 bl[246] br[246] wl[65] vdd gnd cell_6t
Xbit_r66_c246 bl[246] br[246] wl[66] vdd gnd cell_6t
Xbit_r67_c246 bl[246] br[246] wl[67] vdd gnd cell_6t
Xbit_r68_c246 bl[246] br[246] wl[68] vdd gnd cell_6t
Xbit_r69_c246 bl[246] br[246] wl[69] vdd gnd cell_6t
Xbit_r70_c246 bl[246] br[246] wl[70] vdd gnd cell_6t
Xbit_r71_c246 bl[246] br[246] wl[71] vdd gnd cell_6t
Xbit_r72_c246 bl[246] br[246] wl[72] vdd gnd cell_6t
Xbit_r73_c246 bl[246] br[246] wl[73] vdd gnd cell_6t
Xbit_r74_c246 bl[246] br[246] wl[74] vdd gnd cell_6t
Xbit_r75_c246 bl[246] br[246] wl[75] vdd gnd cell_6t
Xbit_r76_c246 bl[246] br[246] wl[76] vdd gnd cell_6t
Xbit_r77_c246 bl[246] br[246] wl[77] vdd gnd cell_6t
Xbit_r78_c246 bl[246] br[246] wl[78] vdd gnd cell_6t
Xbit_r79_c246 bl[246] br[246] wl[79] vdd gnd cell_6t
Xbit_r80_c246 bl[246] br[246] wl[80] vdd gnd cell_6t
Xbit_r81_c246 bl[246] br[246] wl[81] vdd gnd cell_6t
Xbit_r82_c246 bl[246] br[246] wl[82] vdd gnd cell_6t
Xbit_r83_c246 bl[246] br[246] wl[83] vdd gnd cell_6t
Xbit_r84_c246 bl[246] br[246] wl[84] vdd gnd cell_6t
Xbit_r85_c246 bl[246] br[246] wl[85] vdd gnd cell_6t
Xbit_r86_c246 bl[246] br[246] wl[86] vdd gnd cell_6t
Xbit_r87_c246 bl[246] br[246] wl[87] vdd gnd cell_6t
Xbit_r88_c246 bl[246] br[246] wl[88] vdd gnd cell_6t
Xbit_r89_c246 bl[246] br[246] wl[89] vdd gnd cell_6t
Xbit_r90_c246 bl[246] br[246] wl[90] vdd gnd cell_6t
Xbit_r91_c246 bl[246] br[246] wl[91] vdd gnd cell_6t
Xbit_r92_c246 bl[246] br[246] wl[92] vdd gnd cell_6t
Xbit_r93_c246 bl[246] br[246] wl[93] vdd gnd cell_6t
Xbit_r94_c246 bl[246] br[246] wl[94] vdd gnd cell_6t
Xbit_r95_c246 bl[246] br[246] wl[95] vdd gnd cell_6t
Xbit_r96_c246 bl[246] br[246] wl[96] vdd gnd cell_6t
Xbit_r97_c246 bl[246] br[246] wl[97] vdd gnd cell_6t
Xbit_r98_c246 bl[246] br[246] wl[98] vdd gnd cell_6t
Xbit_r99_c246 bl[246] br[246] wl[99] vdd gnd cell_6t
Xbit_r100_c246 bl[246] br[246] wl[100] vdd gnd cell_6t
Xbit_r101_c246 bl[246] br[246] wl[101] vdd gnd cell_6t
Xbit_r102_c246 bl[246] br[246] wl[102] vdd gnd cell_6t
Xbit_r103_c246 bl[246] br[246] wl[103] vdd gnd cell_6t
Xbit_r104_c246 bl[246] br[246] wl[104] vdd gnd cell_6t
Xbit_r105_c246 bl[246] br[246] wl[105] vdd gnd cell_6t
Xbit_r106_c246 bl[246] br[246] wl[106] vdd gnd cell_6t
Xbit_r107_c246 bl[246] br[246] wl[107] vdd gnd cell_6t
Xbit_r108_c246 bl[246] br[246] wl[108] vdd gnd cell_6t
Xbit_r109_c246 bl[246] br[246] wl[109] vdd gnd cell_6t
Xbit_r110_c246 bl[246] br[246] wl[110] vdd gnd cell_6t
Xbit_r111_c246 bl[246] br[246] wl[111] vdd gnd cell_6t
Xbit_r112_c246 bl[246] br[246] wl[112] vdd gnd cell_6t
Xbit_r113_c246 bl[246] br[246] wl[113] vdd gnd cell_6t
Xbit_r114_c246 bl[246] br[246] wl[114] vdd gnd cell_6t
Xbit_r115_c246 bl[246] br[246] wl[115] vdd gnd cell_6t
Xbit_r116_c246 bl[246] br[246] wl[116] vdd gnd cell_6t
Xbit_r117_c246 bl[246] br[246] wl[117] vdd gnd cell_6t
Xbit_r118_c246 bl[246] br[246] wl[118] vdd gnd cell_6t
Xbit_r119_c246 bl[246] br[246] wl[119] vdd gnd cell_6t
Xbit_r120_c246 bl[246] br[246] wl[120] vdd gnd cell_6t
Xbit_r121_c246 bl[246] br[246] wl[121] vdd gnd cell_6t
Xbit_r122_c246 bl[246] br[246] wl[122] vdd gnd cell_6t
Xbit_r123_c246 bl[246] br[246] wl[123] vdd gnd cell_6t
Xbit_r124_c246 bl[246] br[246] wl[124] vdd gnd cell_6t
Xbit_r125_c246 bl[246] br[246] wl[125] vdd gnd cell_6t
Xbit_r126_c246 bl[246] br[246] wl[126] vdd gnd cell_6t
Xbit_r127_c246 bl[246] br[246] wl[127] vdd gnd cell_6t
Xbit_r128_c246 bl[246] br[246] wl[128] vdd gnd cell_6t
Xbit_r129_c246 bl[246] br[246] wl[129] vdd gnd cell_6t
Xbit_r130_c246 bl[246] br[246] wl[130] vdd gnd cell_6t
Xbit_r131_c246 bl[246] br[246] wl[131] vdd gnd cell_6t
Xbit_r132_c246 bl[246] br[246] wl[132] vdd gnd cell_6t
Xbit_r133_c246 bl[246] br[246] wl[133] vdd gnd cell_6t
Xbit_r134_c246 bl[246] br[246] wl[134] vdd gnd cell_6t
Xbit_r135_c246 bl[246] br[246] wl[135] vdd gnd cell_6t
Xbit_r136_c246 bl[246] br[246] wl[136] vdd gnd cell_6t
Xbit_r137_c246 bl[246] br[246] wl[137] vdd gnd cell_6t
Xbit_r138_c246 bl[246] br[246] wl[138] vdd gnd cell_6t
Xbit_r139_c246 bl[246] br[246] wl[139] vdd gnd cell_6t
Xbit_r140_c246 bl[246] br[246] wl[140] vdd gnd cell_6t
Xbit_r141_c246 bl[246] br[246] wl[141] vdd gnd cell_6t
Xbit_r142_c246 bl[246] br[246] wl[142] vdd gnd cell_6t
Xbit_r143_c246 bl[246] br[246] wl[143] vdd gnd cell_6t
Xbit_r144_c246 bl[246] br[246] wl[144] vdd gnd cell_6t
Xbit_r145_c246 bl[246] br[246] wl[145] vdd gnd cell_6t
Xbit_r146_c246 bl[246] br[246] wl[146] vdd gnd cell_6t
Xbit_r147_c246 bl[246] br[246] wl[147] vdd gnd cell_6t
Xbit_r148_c246 bl[246] br[246] wl[148] vdd gnd cell_6t
Xbit_r149_c246 bl[246] br[246] wl[149] vdd gnd cell_6t
Xbit_r150_c246 bl[246] br[246] wl[150] vdd gnd cell_6t
Xbit_r151_c246 bl[246] br[246] wl[151] vdd gnd cell_6t
Xbit_r152_c246 bl[246] br[246] wl[152] vdd gnd cell_6t
Xbit_r153_c246 bl[246] br[246] wl[153] vdd gnd cell_6t
Xbit_r154_c246 bl[246] br[246] wl[154] vdd gnd cell_6t
Xbit_r155_c246 bl[246] br[246] wl[155] vdd gnd cell_6t
Xbit_r156_c246 bl[246] br[246] wl[156] vdd gnd cell_6t
Xbit_r157_c246 bl[246] br[246] wl[157] vdd gnd cell_6t
Xbit_r158_c246 bl[246] br[246] wl[158] vdd gnd cell_6t
Xbit_r159_c246 bl[246] br[246] wl[159] vdd gnd cell_6t
Xbit_r160_c246 bl[246] br[246] wl[160] vdd gnd cell_6t
Xbit_r161_c246 bl[246] br[246] wl[161] vdd gnd cell_6t
Xbit_r162_c246 bl[246] br[246] wl[162] vdd gnd cell_6t
Xbit_r163_c246 bl[246] br[246] wl[163] vdd gnd cell_6t
Xbit_r164_c246 bl[246] br[246] wl[164] vdd gnd cell_6t
Xbit_r165_c246 bl[246] br[246] wl[165] vdd gnd cell_6t
Xbit_r166_c246 bl[246] br[246] wl[166] vdd gnd cell_6t
Xbit_r167_c246 bl[246] br[246] wl[167] vdd gnd cell_6t
Xbit_r168_c246 bl[246] br[246] wl[168] vdd gnd cell_6t
Xbit_r169_c246 bl[246] br[246] wl[169] vdd gnd cell_6t
Xbit_r170_c246 bl[246] br[246] wl[170] vdd gnd cell_6t
Xbit_r171_c246 bl[246] br[246] wl[171] vdd gnd cell_6t
Xbit_r172_c246 bl[246] br[246] wl[172] vdd gnd cell_6t
Xbit_r173_c246 bl[246] br[246] wl[173] vdd gnd cell_6t
Xbit_r174_c246 bl[246] br[246] wl[174] vdd gnd cell_6t
Xbit_r175_c246 bl[246] br[246] wl[175] vdd gnd cell_6t
Xbit_r176_c246 bl[246] br[246] wl[176] vdd gnd cell_6t
Xbit_r177_c246 bl[246] br[246] wl[177] vdd gnd cell_6t
Xbit_r178_c246 bl[246] br[246] wl[178] vdd gnd cell_6t
Xbit_r179_c246 bl[246] br[246] wl[179] vdd gnd cell_6t
Xbit_r180_c246 bl[246] br[246] wl[180] vdd gnd cell_6t
Xbit_r181_c246 bl[246] br[246] wl[181] vdd gnd cell_6t
Xbit_r182_c246 bl[246] br[246] wl[182] vdd gnd cell_6t
Xbit_r183_c246 bl[246] br[246] wl[183] vdd gnd cell_6t
Xbit_r184_c246 bl[246] br[246] wl[184] vdd gnd cell_6t
Xbit_r185_c246 bl[246] br[246] wl[185] vdd gnd cell_6t
Xbit_r186_c246 bl[246] br[246] wl[186] vdd gnd cell_6t
Xbit_r187_c246 bl[246] br[246] wl[187] vdd gnd cell_6t
Xbit_r188_c246 bl[246] br[246] wl[188] vdd gnd cell_6t
Xbit_r189_c246 bl[246] br[246] wl[189] vdd gnd cell_6t
Xbit_r190_c246 bl[246] br[246] wl[190] vdd gnd cell_6t
Xbit_r191_c246 bl[246] br[246] wl[191] vdd gnd cell_6t
Xbit_r192_c246 bl[246] br[246] wl[192] vdd gnd cell_6t
Xbit_r193_c246 bl[246] br[246] wl[193] vdd gnd cell_6t
Xbit_r194_c246 bl[246] br[246] wl[194] vdd gnd cell_6t
Xbit_r195_c246 bl[246] br[246] wl[195] vdd gnd cell_6t
Xbit_r196_c246 bl[246] br[246] wl[196] vdd gnd cell_6t
Xbit_r197_c246 bl[246] br[246] wl[197] vdd gnd cell_6t
Xbit_r198_c246 bl[246] br[246] wl[198] vdd gnd cell_6t
Xbit_r199_c246 bl[246] br[246] wl[199] vdd gnd cell_6t
Xbit_r200_c246 bl[246] br[246] wl[200] vdd gnd cell_6t
Xbit_r201_c246 bl[246] br[246] wl[201] vdd gnd cell_6t
Xbit_r202_c246 bl[246] br[246] wl[202] vdd gnd cell_6t
Xbit_r203_c246 bl[246] br[246] wl[203] vdd gnd cell_6t
Xbit_r204_c246 bl[246] br[246] wl[204] vdd gnd cell_6t
Xbit_r205_c246 bl[246] br[246] wl[205] vdd gnd cell_6t
Xbit_r206_c246 bl[246] br[246] wl[206] vdd gnd cell_6t
Xbit_r207_c246 bl[246] br[246] wl[207] vdd gnd cell_6t
Xbit_r208_c246 bl[246] br[246] wl[208] vdd gnd cell_6t
Xbit_r209_c246 bl[246] br[246] wl[209] vdd gnd cell_6t
Xbit_r210_c246 bl[246] br[246] wl[210] vdd gnd cell_6t
Xbit_r211_c246 bl[246] br[246] wl[211] vdd gnd cell_6t
Xbit_r212_c246 bl[246] br[246] wl[212] vdd gnd cell_6t
Xbit_r213_c246 bl[246] br[246] wl[213] vdd gnd cell_6t
Xbit_r214_c246 bl[246] br[246] wl[214] vdd gnd cell_6t
Xbit_r215_c246 bl[246] br[246] wl[215] vdd gnd cell_6t
Xbit_r216_c246 bl[246] br[246] wl[216] vdd gnd cell_6t
Xbit_r217_c246 bl[246] br[246] wl[217] vdd gnd cell_6t
Xbit_r218_c246 bl[246] br[246] wl[218] vdd gnd cell_6t
Xbit_r219_c246 bl[246] br[246] wl[219] vdd gnd cell_6t
Xbit_r220_c246 bl[246] br[246] wl[220] vdd gnd cell_6t
Xbit_r221_c246 bl[246] br[246] wl[221] vdd gnd cell_6t
Xbit_r222_c246 bl[246] br[246] wl[222] vdd gnd cell_6t
Xbit_r223_c246 bl[246] br[246] wl[223] vdd gnd cell_6t
Xbit_r224_c246 bl[246] br[246] wl[224] vdd gnd cell_6t
Xbit_r225_c246 bl[246] br[246] wl[225] vdd gnd cell_6t
Xbit_r226_c246 bl[246] br[246] wl[226] vdd gnd cell_6t
Xbit_r227_c246 bl[246] br[246] wl[227] vdd gnd cell_6t
Xbit_r228_c246 bl[246] br[246] wl[228] vdd gnd cell_6t
Xbit_r229_c246 bl[246] br[246] wl[229] vdd gnd cell_6t
Xbit_r230_c246 bl[246] br[246] wl[230] vdd gnd cell_6t
Xbit_r231_c246 bl[246] br[246] wl[231] vdd gnd cell_6t
Xbit_r232_c246 bl[246] br[246] wl[232] vdd gnd cell_6t
Xbit_r233_c246 bl[246] br[246] wl[233] vdd gnd cell_6t
Xbit_r234_c246 bl[246] br[246] wl[234] vdd gnd cell_6t
Xbit_r235_c246 bl[246] br[246] wl[235] vdd gnd cell_6t
Xbit_r236_c246 bl[246] br[246] wl[236] vdd gnd cell_6t
Xbit_r237_c246 bl[246] br[246] wl[237] vdd gnd cell_6t
Xbit_r238_c246 bl[246] br[246] wl[238] vdd gnd cell_6t
Xbit_r239_c246 bl[246] br[246] wl[239] vdd gnd cell_6t
Xbit_r240_c246 bl[246] br[246] wl[240] vdd gnd cell_6t
Xbit_r241_c246 bl[246] br[246] wl[241] vdd gnd cell_6t
Xbit_r242_c246 bl[246] br[246] wl[242] vdd gnd cell_6t
Xbit_r243_c246 bl[246] br[246] wl[243] vdd gnd cell_6t
Xbit_r244_c246 bl[246] br[246] wl[244] vdd gnd cell_6t
Xbit_r245_c246 bl[246] br[246] wl[245] vdd gnd cell_6t
Xbit_r246_c246 bl[246] br[246] wl[246] vdd gnd cell_6t
Xbit_r247_c246 bl[246] br[246] wl[247] vdd gnd cell_6t
Xbit_r248_c246 bl[246] br[246] wl[248] vdd gnd cell_6t
Xbit_r249_c246 bl[246] br[246] wl[249] vdd gnd cell_6t
Xbit_r250_c246 bl[246] br[246] wl[250] vdd gnd cell_6t
Xbit_r251_c246 bl[246] br[246] wl[251] vdd gnd cell_6t
Xbit_r252_c246 bl[246] br[246] wl[252] vdd gnd cell_6t
Xbit_r253_c246 bl[246] br[246] wl[253] vdd gnd cell_6t
Xbit_r254_c246 bl[246] br[246] wl[254] vdd gnd cell_6t
Xbit_r255_c246 bl[246] br[246] wl[255] vdd gnd cell_6t
Xbit_r0_c247 bl[247] br[247] wl[0] vdd gnd cell_6t
Xbit_r1_c247 bl[247] br[247] wl[1] vdd gnd cell_6t
Xbit_r2_c247 bl[247] br[247] wl[2] vdd gnd cell_6t
Xbit_r3_c247 bl[247] br[247] wl[3] vdd gnd cell_6t
Xbit_r4_c247 bl[247] br[247] wl[4] vdd gnd cell_6t
Xbit_r5_c247 bl[247] br[247] wl[5] vdd gnd cell_6t
Xbit_r6_c247 bl[247] br[247] wl[6] vdd gnd cell_6t
Xbit_r7_c247 bl[247] br[247] wl[7] vdd gnd cell_6t
Xbit_r8_c247 bl[247] br[247] wl[8] vdd gnd cell_6t
Xbit_r9_c247 bl[247] br[247] wl[9] vdd gnd cell_6t
Xbit_r10_c247 bl[247] br[247] wl[10] vdd gnd cell_6t
Xbit_r11_c247 bl[247] br[247] wl[11] vdd gnd cell_6t
Xbit_r12_c247 bl[247] br[247] wl[12] vdd gnd cell_6t
Xbit_r13_c247 bl[247] br[247] wl[13] vdd gnd cell_6t
Xbit_r14_c247 bl[247] br[247] wl[14] vdd gnd cell_6t
Xbit_r15_c247 bl[247] br[247] wl[15] vdd gnd cell_6t
Xbit_r16_c247 bl[247] br[247] wl[16] vdd gnd cell_6t
Xbit_r17_c247 bl[247] br[247] wl[17] vdd gnd cell_6t
Xbit_r18_c247 bl[247] br[247] wl[18] vdd gnd cell_6t
Xbit_r19_c247 bl[247] br[247] wl[19] vdd gnd cell_6t
Xbit_r20_c247 bl[247] br[247] wl[20] vdd gnd cell_6t
Xbit_r21_c247 bl[247] br[247] wl[21] vdd gnd cell_6t
Xbit_r22_c247 bl[247] br[247] wl[22] vdd gnd cell_6t
Xbit_r23_c247 bl[247] br[247] wl[23] vdd gnd cell_6t
Xbit_r24_c247 bl[247] br[247] wl[24] vdd gnd cell_6t
Xbit_r25_c247 bl[247] br[247] wl[25] vdd gnd cell_6t
Xbit_r26_c247 bl[247] br[247] wl[26] vdd gnd cell_6t
Xbit_r27_c247 bl[247] br[247] wl[27] vdd gnd cell_6t
Xbit_r28_c247 bl[247] br[247] wl[28] vdd gnd cell_6t
Xbit_r29_c247 bl[247] br[247] wl[29] vdd gnd cell_6t
Xbit_r30_c247 bl[247] br[247] wl[30] vdd gnd cell_6t
Xbit_r31_c247 bl[247] br[247] wl[31] vdd gnd cell_6t
Xbit_r32_c247 bl[247] br[247] wl[32] vdd gnd cell_6t
Xbit_r33_c247 bl[247] br[247] wl[33] vdd gnd cell_6t
Xbit_r34_c247 bl[247] br[247] wl[34] vdd gnd cell_6t
Xbit_r35_c247 bl[247] br[247] wl[35] vdd gnd cell_6t
Xbit_r36_c247 bl[247] br[247] wl[36] vdd gnd cell_6t
Xbit_r37_c247 bl[247] br[247] wl[37] vdd gnd cell_6t
Xbit_r38_c247 bl[247] br[247] wl[38] vdd gnd cell_6t
Xbit_r39_c247 bl[247] br[247] wl[39] vdd gnd cell_6t
Xbit_r40_c247 bl[247] br[247] wl[40] vdd gnd cell_6t
Xbit_r41_c247 bl[247] br[247] wl[41] vdd gnd cell_6t
Xbit_r42_c247 bl[247] br[247] wl[42] vdd gnd cell_6t
Xbit_r43_c247 bl[247] br[247] wl[43] vdd gnd cell_6t
Xbit_r44_c247 bl[247] br[247] wl[44] vdd gnd cell_6t
Xbit_r45_c247 bl[247] br[247] wl[45] vdd gnd cell_6t
Xbit_r46_c247 bl[247] br[247] wl[46] vdd gnd cell_6t
Xbit_r47_c247 bl[247] br[247] wl[47] vdd gnd cell_6t
Xbit_r48_c247 bl[247] br[247] wl[48] vdd gnd cell_6t
Xbit_r49_c247 bl[247] br[247] wl[49] vdd gnd cell_6t
Xbit_r50_c247 bl[247] br[247] wl[50] vdd gnd cell_6t
Xbit_r51_c247 bl[247] br[247] wl[51] vdd gnd cell_6t
Xbit_r52_c247 bl[247] br[247] wl[52] vdd gnd cell_6t
Xbit_r53_c247 bl[247] br[247] wl[53] vdd gnd cell_6t
Xbit_r54_c247 bl[247] br[247] wl[54] vdd gnd cell_6t
Xbit_r55_c247 bl[247] br[247] wl[55] vdd gnd cell_6t
Xbit_r56_c247 bl[247] br[247] wl[56] vdd gnd cell_6t
Xbit_r57_c247 bl[247] br[247] wl[57] vdd gnd cell_6t
Xbit_r58_c247 bl[247] br[247] wl[58] vdd gnd cell_6t
Xbit_r59_c247 bl[247] br[247] wl[59] vdd gnd cell_6t
Xbit_r60_c247 bl[247] br[247] wl[60] vdd gnd cell_6t
Xbit_r61_c247 bl[247] br[247] wl[61] vdd gnd cell_6t
Xbit_r62_c247 bl[247] br[247] wl[62] vdd gnd cell_6t
Xbit_r63_c247 bl[247] br[247] wl[63] vdd gnd cell_6t
Xbit_r64_c247 bl[247] br[247] wl[64] vdd gnd cell_6t
Xbit_r65_c247 bl[247] br[247] wl[65] vdd gnd cell_6t
Xbit_r66_c247 bl[247] br[247] wl[66] vdd gnd cell_6t
Xbit_r67_c247 bl[247] br[247] wl[67] vdd gnd cell_6t
Xbit_r68_c247 bl[247] br[247] wl[68] vdd gnd cell_6t
Xbit_r69_c247 bl[247] br[247] wl[69] vdd gnd cell_6t
Xbit_r70_c247 bl[247] br[247] wl[70] vdd gnd cell_6t
Xbit_r71_c247 bl[247] br[247] wl[71] vdd gnd cell_6t
Xbit_r72_c247 bl[247] br[247] wl[72] vdd gnd cell_6t
Xbit_r73_c247 bl[247] br[247] wl[73] vdd gnd cell_6t
Xbit_r74_c247 bl[247] br[247] wl[74] vdd gnd cell_6t
Xbit_r75_c247 bl[247] br[247] wl[75] vdd gnd cell_6t
Xbit_r76_c247 bl[247] br[247] wl[76] vdd gnd cell_6t
Xbit_r77_c247 bl[247] br[247] wl[77] vdd gnd cell_6t
Xbit_r78_c247 bl[247] br[247] wl[78] vdd gnd cell_6t
Xbit_r79_c247 bl[247] br[247] wl[79] vdd gnd cell_6t
Xbit_r80_c247 bl[247] br[247] wl[80] vdd gnd cell_6t
Xbit_r81_c247 bl[247] br[247] wl[81] vdd gnd cell_6t
Xbit_r82_c247 bl[247] br[247] wl[82] vdd gnd cell_6t
Xbit_r83_c247 bl[247] br[247] wl[83] vdd gnd cell_6t
Xbit_r84_c247 bl[247] br[247] wl[84] vdd gnd cell_6t
Xbit_r85_c247 bl[247] br[247] wl[85] vdd gnd cell_6t
Xbit_r86_c247 bl[247] br[247] wl[86] vdd gnd cell_6t
Xbit_r87_c247 bl[247] br[247] wl[87] vdd gnd cell_6t
Xbit_r88_c247 bl[247] br[247] wl[88] vdd gnd cell_6t
Xbit_r89_c247 bl[247] br[247] wl[89] vdd gnd cell_6t
Xbit_r90_c247 bl[247] br[247] wl[90] vdd gnd cell_6t
Xbit_r91_c247 bl[247] br[247] wl[91] vdd gnd cell_6t
Xbit_r92_c247 bl[247] br[247] wl[92] vdd gnd cell_6t
Xbit_r93_c247 bl[247] br[247] wl[93] vdd gnd cell_6t
Xbit_r94_c247 bl[247] br[247] wl[94] vdd gnd cell_6t
Xbit_r95_c247 bl[247] br[247] wl[95] vdd gnd cell_6t
Xbit_r96_c247 bl[247] br[247] wl[96] vdd gnd cell_6t
Xbit_r97_c247 bl[247] br[247] wl[97] vdd gnd cell_6t
Xbit_r98_c247 bl[247] br[247] wl[98] vdd gnd cell_6t
Xbit_r99_c247 bl[247] br[247] wl[99] vdd gnd cell_6t
Xbit_r100_c247 bl[247] br[247] wl[100] vdd gnd cell_6t
Xbit_r101_c247 bl[247] br[247] wl[101] vdd gnd cell_6t
Xbit_r102_c247 bl[247] br[247] wl[102] vdd gnd cell_6t
Xbit_r103_c247 bl[247] br[247] wl[103] vdd gnd cell_6t
Xbit_r104_c247 bl[247] br[247] wl[104] vdd gnd cell_6t
Xbit_r105_c247 bl[247] br[247] wl[105] vdd gnd cell_6t
Xbit_r106_c247 bl[247] br[247] wl[106] vdd gnd cell_6t
Xbit_r107_c247 bl[247] br[247] wl[107] vdd gnd cell_6t
Xbit_r108_c247 bl[247] br[247] wl[108] vdd gnd cell_6t
Xbit_r109_c247 bl[247] br[247] wl[109] vdd gnd cell_6t
Xbit_r110_c247 bl[247] br[247] wl[110] vdd gnd cell_6t
Xbit_r111_c247 bl[247] br[247] wl[111] vdd gnd cell_6t
Xbit_r112_c247 bl[247] br[247] wl[112] vdd gnd cell_6t
Xbit_r113_c247 bl[247] br[247] wl[113] vdd gnd cell_6t
Xbit_r114_c247 bl[247] br[247] wl[114] vdd gnd cell_6t
Xbit_r115_c247 bl[247] br[247] wl[115] vdd gnd cell_6t
Xbit_r116_c247 bl[247] br[247] wl[116] vdd gnd cell_6t
Xbit_r117_c247 bl[247] br[247] wl[117] vdd gnd cell_6t
Xbit_r118_c247 bl[247] br[247] wl[118] vdd gnd cell_6t
Xbit_r119_c247 bl[247] br[247] wl[119] vdd gnd cell_6t
Xbit_r120_c247 bl[247] br[247] wl[120] vdd gnd cell_6t
Xbit_r121_c247 bl[247] br[247] wl[121] vdd gnd cell_6t
Xbit_r122_c247 bl[247] br[247] wl[122] vdd gnd cell_6t
Xbit_r123_c247 bl[247] br[247] wl[123] vdd gnd cell_6t
Xbit_r124_c247 bl[247] br[247] wl[124] vdd gnd cell_6t
Xbit_r125_c247 bl[247] br[247] wl[125] vdd gnd cell_6t
Xbit_r126_c247 bl[247] br[247] wl[126] vdd gnd cell_6t
Xbit_r127_c247 bl[247] br[247] wl[127] vdd gnd cell_6t
Xbit_r128_c247 bl[247] br[247] wl[128] vdd gnd cell_6t
Xbit_r129_c247 bl[247] br[247] wl[129] vdd gnd cell_6t
Xbit_r130_c247 bl[247] br[247] wl[130] vdd gnd cell_6t
Xbit_r131_c247 bl[247] br[247] wl[131] vdd gnd cell_6t
Xbit_r132_c247 bl[247] br[247] wl[132] vdd gnd cell_6t
Xbit_r133_c247 bl[247] br[247] wl[133] vdd gnd cell_6t
Xbit_r134_c247 bl[247] br[247] wl[134] vdd gnd cell_6t
Xbit_r135_c247 bl[247] br[247] wl[135] vdd gnd cell_6t
Xbit_r136_c247 bl[247] br[247] wl[136] vdd gnd cell_6t
Xbit_r137_c247 bl[247] br[247] wl[137] vdd gnd cell_6t
Xbit_r138_c247 bl[247] br[247] wl[138] vdd gnd cell_6t
Xbit_r139_c247 bl[247] br[247] wl[139] vdd gnd cell_6t
Xbit_r140_c247 bl[247] br[247] wl[140] vdd gnd cell_6t
Xbit_r141_c247 bl[247] br[247] wl[141] vdd gnd cell_6t
Xbit_r142_c247 bl[247] br[247] wl[142] vdd gnd cell_6t
Xbit_r143_c247 bl[247] br[247] wl[143] vdd gnd cell_6t
Xbit_r144_c247 bl[247] br[247] wl[144] vdd gnd cell_6t
Xbit_r145_c247 bl[247] br[247] wl[145] vdd gnd cell_6t
Xbit_r146_c247 bl[247] br[247] wl[146] vdd gnd cell_6t
Xbit_r147_c247 bl[247] br[247] wl[147] vdd gnd cell_6t
Xbit_r148_c247 bl[247] br[247] wl[148] vdd gnd cell_6t
Xbit_r149_c247 bl[247] br[247] wl[149] vdd gnd cell_6t
Xbit_r150_c247 bl[247] br[247] wl[150] vdd gnd cell_6t
Xbit_r151_c247 bl[247] br[247] wl[151] vdd gnd cell_6t
Xbit_r152_c247 bl[247] br[247] wl[152] vdd gnd cell_6t
Xbit_r153_c247 bl[247] br[247] wl[153] vdd gnd cell_6t
Xbit_r154_c247 bl[247] br[247] wl[154] vdd gnd cell_6t
Xbit_r155_c247 bl[247] br[247] wl[155] vdd gnd cell_6t
Xbit_r156_c247 bl[247] br[247] wl[156] vdd gnd cell_6t
Xbit_r157_c247 bl[247] br[247] wl[157] vdd gnd cell_6t
Xbit_r158_c247 bl[247] br[247] wl[158] vdd gnd cell_6t
Xbit_r159_c247 bl[247] br[247] wl[159] vdd gnd cell_6t
Xbit_r160_c247 bl[247] br[247] wl[160] vdd gnd cell_6t
Xbit_r161_c247 bl[247] br[247] wl[161] vdd gnd cell_6t
Xbit_r162_c247 bl[247] br[247] wl[162] vdd gnd cell_6t
Xbit_r163_c247 bl[247] br[247] wl[163] vdd gnd cell_6t
Xbit_r164_c247 bl[247] br[247] wl[164] vdd gnd cell_6t
Xbit_r165_c247 bl[247] br[247] wl[165] vdd gnd cell_6t
Xbit_r166_c247 bl[247] br[247] wl[166] vdd gnd cell_6t
Xbit_r167_c247 bl[247] br[247] wl[167] vdd gnd cell_6t
Xbit_r168_c247 bl[247] br[247] wl[168] vdd gnd cell_6t
Xbit_r169_c247 bl[247] br[247] wl[169] vdd gnd cell_6t
Xbit_r170_c247 bl[247] br[247] wl[170] vdd gnd cell_6t
Xbit_r171_c247 bl[247] br[247] wl[171] vdd gnd cell_6t
Xbit_r172_c247 bl[247] br[247] wl[172] vdd gnd cell_6t
Xbit_r173_c247 bl[247] br[247] wl[173] vdd gnd cell_6t
Xbit_r174_c247 bl[247] br[247] wl[174] vdd gnd cell_6t
Xbit_r175_c247 bl[247] br[247] wl[175] vdd gnd cell_6t
Xbit_r176_c247 bl[247] br[247] wl[176] vdd gnd cell_6t
Xbit_r177_c247 bl[247] br[247] wl[177] vdd gnd cell_6t
Xbit_r178_c247 bl[247] br[247] wl[178] vdd gnd cell_6t
Xbit_r179_c247 bl[247] br[247] wl[179] vdd gnd cell_6t
Xbit_r180_c247 bl[247] br[247] wl[180] vdd gnd cell_6t
Xbit_r181_c247 bl[247] br[247] wl[181] vdd gnd cell_6t
Xbit_r182_c247 bl[247] br[247] wl[182] vdd gnd cell_6t
Xbit_r183_c247 bl[247] br[247] wl[183] vdd gnd cell_6t
Xbit_r184_c247 bl[247] br[247] wl[184] vdd gnd cell_6t
Xbit_r185_c247 bl[247] br[247] wl[185] vdd gnd cell_6t
Xbit_r186_c247 bl[247] br[247] wl[186] vdd gnd cell_6t
Xbit_r187_c247 bl[247] br[247] wl[187] vdd gnd cell_6t
Xbit_r188_c247 bl[247] br[247] wl[188] vdd gnd cell_6t
Xbit_r189_c247 bl[247] br[247] wl[189] vdd gnd cell_6t
Xbit_r190_c247 bl[247] br[247] wl[190] vdd gnd cell_6t
Xbit_r191_c247 bl[247] br[247] wl[191] vdd gnd cell_6t
Xbit_r192_c247 bl[247] br[247] wl[192] vdd gnd cell_6t
Xbit_r193_c247 bl[247] br[247] wl[193] vdd gnd cell_6t
Xbit_r194_c247 bl[247] br[247] wl[194] vdd gnd cell_6t
Xbit_r195_c247 bl[247] br[247] wl[195] vdd gnd cell_6t
Xbit_r196_c247 bl[247] br[247] wl[196] vdd gnd cell_6t
Xbit_r197_c247 bl[247] br[247] wl[197] vdd gnd cell_6t
Xbit_r198_c247 bl[247] br[247] wl[198] vdd gnd cell_6t
Xbit_r199_c247 bl[247] br[247] wl[199] vdd gnd cell_6t
Xbit_r200_c247 bl[247] br[247] wl[200] vdd gnd cell_6t
Xbit_r201_c247 bl[247] br[247] wl[201] vdd gnd cell_6t
Xbit_r202_c247 bl[247] br[247] wl[202] vdd gnd cell_6t
Xbit_r203_c247 bl[247] br[247] wl[203] vdd gnd cell_6t
Xbit_r204_c247 bl[247] br[247] wl[204] vdd gnd cell_6t
Xbit_r205_c247 bl[247] br[247] wl[205] vdd gnd cell_6t
Xbit_r206_c247 bl[247] br[247] wl[206] vdd gnd cell_6t
Xbit_r207_c247 bl[247] br[247] wl[207] vdd gnd cell_6t
Xbit_r208_c247 bl[247] br[247] wl[208] vdd gnd cell_6t
Xbit_r209_c247 bl[247] br[247] wl[209] vdd gnd cell_6t
Xbit_r210_c247 bl[247] br[247] wl[210] vdd gnd cell_6t
Xbit_r211_c247 bl[247] br[247] wl[211] vdd gnd cell_6t
Xbit_r212_c247 bl[247] br[247] wl[212] vdd gnd cell_6t
Xbit_r213_c247 bl[247] br[247] wl[213] vdd gnd cell_6t
Xbit_r214_c247 bl[247] br[247] wl[214] vdd gnd cell_6t
Xbit_r215_c247 bl[247] br[247] wl[215] vdd gnd cell_6t
Xbit_r216_c247 bl[247] br[247] wl[216] vdd gnd cell_6t
Xbit_r217_c247 bl[247] br[247] wl[217] vdd gnd cell_6t
Xbit_r218_c247 bl[247] br[247] wl[218] vdd gnd cell_6t
Xbit_r219_c247 bl[247] br[247] wl[219] vdd gnd cell_6t
Xbit_r220_c247 bl[247] br[247] wl[220] vdd gnd cell_6t
Xbit_r221_c247 bl[247] br[247] wl[221] vdd gnd cell_6t
Xbit_r222_c247 bl[247] br[247] wl[222] vdd gnd cell_6t
Xbit_r223_c247 bl[247] br[247] wl[223] vdd gnd cell_6t
Xbit_r224_c247 bl[247] br[247] wl[224] vdd gnd cell_6t
Xbit_r225_c247 bl[247] br[247] wl[225] vdd gnd cell_6t
Xbit_r226_c247 bl[247] br[247] wl[226] vdd gnd cell_6t
Xbit_r227_c247 bl[247] br[247] wl[227] vdd gnd cell_6t
Xbit_r228_c247 bl[247] br[247] wl[228] vdd gnd cell_6t
Xbit_r229_c247 bl[247] br[247] wl[229] vdd gnd cell_6t
Xbit_r230_c247 bl[247] br[247] wl[230] vdd gnd cell_6t
Xbit_r231_c247 bl[247] br[247] wl[231] vdd gnd cell_6t
Xbit_r232_c247 bl[247] br[247] wl[232] vdd gnd cell_6t
Xbit_r233_c247 bl[247] br[247] wl[233] vdd gnd cell_6t
Xbit_r234_c247 bl[247] br[247] wl[234] vdd gnd cell_6t
Xbit_r235_c247 bl[247] br[247] wl[235] vdd gnd cell_6t
Xbit_r236_c247 bl[247] br[247] wl[236] vdd gnd cell_6t
Xbit_r237_c247 bl[247] br[247] wl[237] vdd gnd cell_6t
Xbit_r238_c247 bl[247] br[247] wl[238] vdd gnd cell_6t
Xbit_r239_c247 bl[247] br[247] wl[239] vdd gnd cell_6t
Xbit_r240_c247 bl[247] br[247] wl[240] vdd gnd cell_6t
Xbit_r241_c247 bl[247] br[247] wl[241] vdd gnd cell_6t
Xbit_r242_c247 bl[247] br[247] wl[242] vdd gnd cell_6t
Xbit_r243_c247 bl[247] br[247] wl[243] vdd gnd cell_6t
Xbit_r244_c247 bl[247] br[247] wl[244] vdd gnd cell_6t
Xbit_r245_c247 bl[247] br[247] wl[245] vdd gnd cell_6t
Xbit_r246_c247 bl[247] br[247] wl[246] vdd gnd cell_6t
Xbit_r247_c247 bl[247] br[247] wl[247] vdd gnd cell_6t
Xbit_r248_c247 bl[247] br[247] wl[248] vdd gnd cell_6t
Xbit_r249_c247 bl[247] br[247] wl[249] vdd gnd cell_6t
Xbit_r250_c247 bl[247] br[247] wl[250] vdd gnd cell_6t
Xbit_r251_c247 bl[247] br[247] wl[251] vdd gnd cell_6t
Xbit_r252_c247 bl[247] br[247] wl[252] vdd gnd cell_6t
Xbit_r253_c247 bl[247] br[247] wl[253] vdd gnd cell_6t
Xbit_r254_c247 bl[247] br[247] wl[254] vdd gnd cell_6t
Xbit_r255_c247 bl[247] br[247] wl[255] vdd gnd cell_6t
Xbit_r0_c248 bl[248] br[248] wl[0] vdd gnd cell_6t
Xbit_r1_c248 bl[248] br[248] wl[1] vdd gnd cell_6t
Xbit_r2_c248 bl[248] br[248] wl[2] vdd gnd cell_6t
Xbit_r3_c248 bl[248] br[248] wl[3] vdd gnd cell_6t
Xbit_r4_c248 bl[248] br[248] wl[4] vdd gnd cell_6t
Xbit_r5_c248 bl[248] br[248] wl[5] vdd gnd cell_6t
Xbit_r6_c248 bl[248] br[248] wl[6] vdd gnd cell_6t
Xbit_r7_c248 bl[248] br[248] wl[7] vdd gnd cell_6t
Xbit_r8_c248 bl[248] br[248] wl[8] vdd gnd cell_6t
Xbit_r9_c248 bl[248] br[248] wl[9] vdd gnd cell_6t
Xbit_r10_c248 bl[248] br[248] wl[10] vdd gnd cell_6t
Xbit_r11_c248 bl[248] br[248] wl[11] vdd gnd cell_6t
Xbit_r12_c248 bl[248] br[248] wl[12] vdd gnd cell_6t
Xbit_r13_c248 bl[248] br[248] wl[13] vdd gnd cell_6t
Xbit_r14_c248 bl[248] br[248] wl[14] vdd gnd cell_6t
Xbit_r15_c248 bl[248] br[248] wl[15] vdd gnd cell_6t
Xbit_r16_c248 bl[248] br[248] wl[16] vdd gnd cell_6t
Xbit_r17_c248 bl[248] br[248] wl[17] vdd gnd cell_6t
Xbit_r18_c248 bl[248] br[248] wl[18] vdd gnd cell_6t
Xbit_r19_c248 bl[248] br[248] wl[19] vdd gnd cell_6t
Xbit_r20_c248 bl[248] br[248] wl[20] vdd gnd cell_6t
Xbit_r21_c248 bl[248] br[248] wl[21] vdd gnd cell_6t
Xbit_r22_c248 bl[248] br[248] wl[22] vdd gnd cell_6t
Xbit_r23_c248 bl[248] br[248] wl[23] vdd gnd cell_6t
Xbit_r24_c248 bl[248] br[248] wl[24] vdd gnd cell_6t
Xbit_r25_c248 bl[248] br[248] wl[25] vdd gnd cell_6t
Xbit_r26_c248 bl[248] br[248] wl[26] vdd gnd cell_6t
Xbit_r27_c248 bl[248] br[248] wl[27] vdd gnd cell_6t
Xbit_r28_c248 bl[248] br[248] wl[28] vdd gnd cell_6t
Xbit_r29_c248 bl[248] br[248] wl[29] vdd gnd cell_6t
Xbit_r30_c248 bl[248] br[248] wl[30] vdd gnd cell_6t
Xbit_r31_c248 bl[248] br[248] wl[31] vdd gnd cell_6t
Xbit_r32_c248 bl[248] br[248] wl[32] vdd gnd cell_6t
Xbit_r33_c248 bl[248] br[248] wl[33] vdd gnd cell_6t
Xbit_r34_c248 bl[248] br[248] wl[34] vdd gnd cell_6t
Xbit_r35_c248 bl[248] br[248] wl[35] vdd gnd cell_6t
Xbit_r36_c248 bl[248] br[248] wl[36] vdd gnd cell_6t
Xbit_r37_c248 bl[248] br[248] wl[37] vdd gnd cell_6t
Xbit_r38_c248 bl[248] br[248] wl[38] vdd gnd cell_6t
Xbit_r39_c248 bl[248] br[248] wl[39] vdd gnd cell_6t
Xbit_r40_c248 bl[248] br[248] wl[40] vdd gnd cell_6t
Xbit_r41_c248 bl[248] br[248] wl[41] vdd gnd cell_6t
Xbit_r42_c248 bl[248] br[248] wl[42] vdd gnd cell_6t
Xbit_r43_c248 bl[248] br[248] wl[43] vdd gnd cell_6t
Xbit_r44_c248 bl[248] br[248] wl[44] vdd gnd cell_6t
Xbit_r45_c248 bl[248] br[248] wl[45] vdd gnd cell_6t
Xbit_r46_c248 bl[248] br[248] wl[46] vdd gnd cell_6t
Xbit_r47_c248 bl[248] br[248] wl[47] vdd gnd cell_6t
Xbit_r48_c248 bl[248] br[248] wl[48] vdd gnd cell_6t
Xbit_r49_c248 bl[248] br[248] wl[49] vdd gnd cell_6t
Xbit_r50_c248 bl[248] br[248] wl[50] vdd gnd cell_6t
Xbit_r51_c248 bl[248] br[248] wl[51] vdd gnd cell_6t
Xbit_r52_c248 bl[248] br[248] wl[52] vdd gnd cell_6t
Xbit_r53_c248 bl[248] br[248] wl[53] vdd gnd cell_6t
Xbit_r54_c248 bl[248] br[248] wl[54] vdd gnd cell_6t
Xbit_r55_c248 bl[248] br[248] wl[55] vdd gnd cell_6t
Xbit_r56_c248 bl[248] br[248] wl[56] vdd gnd cell_6t
Xbit_r57_c248 bl[248] br[248] wl[57] vdd gnd cell_6t
Xbit_r58_c248 bl[248] br[248] wl[58] vdd gnd cell_6t
Xbit_r59_c248 bl[248] br[248] wl[59] vdd gnd cell_6t
Xbit_r60_c248 bl[248] br[248] wl[60] vdd gnd cell_6t
Xbit_r61_c248 bl[248] br[248] wl[61] vdd gnd cell_6t
Xbit_r62_c248 bl[248] br[248] wl[62] vdd gnd cell_6t
Xbit_r63_c248 bl[248] br[248] wl[63] vdd gnd cell_6t
Xbit_r64_c248 bl[248] br[248] wl[64] vdd gnd cell_6t
Xbit_r65_c248 bl[248] br[248] wl[65] vdd gnd cell_6t
Xbit_r66_c248 bl[248] br[248] wl[66] vdd gnd cell_6t
Xbit_r67_c248 bl[248] br[248] wl[67] vdd gnd cell_6t
Xbit_r68_c248 bl[248] br[248] wl[68] vdd gnd cell_6t
Xbit_r69_c248 bl[248] br[248] wl[69] vdd gnd cell_6t
Xbit_r70_c248 bl[248] br[248] wl[70] vdd gnd cell_6t
Xbit_r71_c248 bl[248] br[248] wl[71] vdd gnd cell_6t
Xbit_r72_c248 bl[248] br[248] wl[72] vdd gnd cell_6t
Xbit_r73_c248 bl[248] br[248] wl[73] vdd gnd cell_6t
Xbit_r74_c248 bl[248] br[248] wl[74] vdd gnd cell_6t
Xbit_r75_c248 bl[248] br[248] wl[75] vdd gnd cell_6t
Xbit_r76_c248 bl[248] br[248] wl[76] vdd gnd cell_6t
Xbit_r77_c248 bl[248] br[248] wl[77] vdd gnd cell_6t
Xbit_r78_c248 bl[248] br[248] wl[78] vdd gnd cell_6t
Xbit_r79_c248 bl[248] br[248] wl[79] vdd gnd cell_6t
Xbit_r80_c248 bl[248] br[248] wl[80] vdd gnd cell_6t
Xbit_r81_c248 bl[248] br[248] wl[81] vdd gnd cell_6t
Xbit_r82_c248 bl[248] br[248] wl[82] vdd gnd cell_6t
Xbit_r83_c248 bl[248] br[248] wl[83] vdd gnd cell_6t
Xbit_r84_c248 bl[248] br[248] wl[84] vdd gnd cell_6t
Xbit_r85_c248 bl[248] br[248] wl[85] vdd gnd cell_6t
Xbit_r86_c248 bl[248] br[248] wl[86] vdd gnd cell_6t
Xbit_r87_c248 bl[248] br[248] wl[87] vdd gnd cell_6t
Xbit_r88_c248 bl[248] br[248] wl[88] vdd gnd cell_6t
Xbit_r89_c248 bl[248] br[248] wl[89] vdd gnd cell_6t
Xbit_r90_c248 bl[248] br[248] wl[90] vdd gnd cell_6t
Xbit_r91_c248 bl[248] br[248] wl[91] vdd gnd cell_6t
Xbit_r92_c248 bl[248] br[248] wl[92] vdd gnd cell_6t
Xbit_r93_c248 bl[248] br[248] wl[93] vdd gnd cell_6t
Xbit_r94_c248 bl[248] br[248] wl[94] vdd gnd cell_6t
Xbit_r95_c248 bl[248] br[248] wl[95] vdd gnd cell_6t
Xbit_r96_c248 bl[248] br[248] wl[96] vdd gnd cell_6t
Xbit_r97_c248 bl[248] br[248] wl[97] vdd gnd cell_6t
Xbit_r98_c248 bl[248] br[248] wl[98] vdd gnd cell_6t
Xbit_r99_c248 bl[248] br[248] wl[99] vdd gnd cell_6t
Xbit_r100_c248 bl[248] br[248] wl[100] vdd gnd cell_6t
Xbit_r101_c248 bl[248] br[248] wl[101] vdd gnd cell_6t
Xbit_r102_c248 bl[248] br[248] wl[102] vdd gnd cell_6t
Xbit_r103_c248 bl[248] br[248] wl[103] vdd gnd cell_6t
Xbit_r104_c248 bl[248] br[248] wl[104] vdd gnd cell_6t
Xbit_r105_c248 bl[248] br[248] wl[105] vdd gnd cell_6t
Xbit_r106_c248 bl[248] br[248] wl[106] vdd gnd cell_6t
Xbit_r107_c248 bl[248] br[248] wl[107] vdd gnd cell_6t
Xbit_r108_c248 bl[248] br[248] wl[108] vdd gnd cell_6t
Xbit_r109_c248 bl[248] br[248] wl[109] vdd gnd cell_6t
Xbit_r110_c248 bl[248] br[248] wl[110] vdd gnd cell_6t
Xbit_r111_c248 bl[248] br[248] wl[111] vdd gnd cell_6t
Xbit_r112_c248 bl[248] br[248] wl[112] vdd gnd cell_6t
Xbit_r113_c248 bl[248] br[248] wl[113] vdd gnd cell_6t
Xbit_r114_c248 bl[248] br[248] wl[114] vdd gnd cell_6t
Xbit_r115_c248 bl[248] br[248] wl[115] vdd gnd cell_6t
Xbit_r116_c248 bl[248] br[248] wl[116] vdd gnd cell_6t
Xbit_r117_c248 bl[248] br[248] wl[117] vdd gnd cell_6t
Xbit_r118_c248 bl[248] br[248] wl[118] vdd gnd cell_6t
Xbit_r119_c248 bl[248] br[248] wl[119] vdd gnd cell_6t
Xbit_r120_c248 bl[248] br[248] wl[120] vdd gnd cell_6t
Xbit_r121_c248 bl[248] br[248] wl[121] vdd gnd cell_6t
Xbit_r122_c248 bl[248] br[248] wl[122] vdd gnd cell_6t
Xbit_r123_c248 bl[248] br[248] wl[123] vdd gnd cell_6t
Xbit_r124_c248 bl[248] br[248] wl[124] vdd gnd cell_6t
Xbit_r125_c248 bl[248] br[248] wl[125] vdd gnd cell_6t
Xbit_r126_c248 bl[248] br[248] wl[126] vdd gnd cell_6t
Xbit_r127_c248 bl[248] br[248] wl[127] vdd gnd cell_6t
Xbit_r128_c248 bl[248] br[248] wl[128] vdd gnd cell_6t
Xbit_r129_c248 bl[248] br[248] wl[129] vdd gnd cell_6t
Xbit_r130_c248 bl[248] br[248] wl[130] vdd gnd cell_6t
Xbit_r131_c248 bl[248] br[248] wl[131] vdd gnd cell_6t
Xbit_r132_c248 bl[248] br[248] wl[132] vdd gnd cell_6t
Xbit_r133_c248 bl[248] br[248] wl[133] vdd gnd cell_6t
Xbit_r134_c248 bl[248] br[248] wl[134] vdd gnd cell_6t
Xbit_r135_c248 bl[248] br[248] wl[135] vdd gnd cell_6t
Xbit_r136_c248 bl[248] br[248] wl[136] vdd gnd cell_6t
Xbit_r137_c248 bl[248] br[248] wl[137] vdd gnd cell_6t
Xbit_r138_c248 bl[248] br[248] wl[138] vdd gnd cell_6t
Xbit_r139_c248 bl[248] br[248] wl[139] vdd gnd cell_6t
Xbit_r140_c248 bl[248] br[248] wl[140] vdd gnd cell_6t
Xbit_r141_c248 bl[248] br[248] wl[141] vdd gnd cell_6t
Xbit_r142_c248 bl[248] br[248] wl[142] vdd gnd cell_6t
Xbit_r143_c248 bl[248] br[248] wl[143] vdd gnd cell_6t
Xbit_r144_c248 bl[248] br[248] wl[144] vdd gnd cell_6t
Xbit_r145_c248 bl[248] br[248] wl[145] vdd gnd cell_6t
Xbit_r146_c248 bl[248] br[248] wl[146] vdd gnd cell_6t
Xbit_r147_c248 bl[248] br[248] wl[147] vdd gnd cell_6t
Xbit_r148_c248 bl[248] br[248] wl[148] vdd gnd cell_6t
Xbit_r149_c248 bl[248] br[248] wl[149] vdd gnd cell_6t
Xbit_r150_c248 bl[248] br[248] wl[150] vdd gnd cell_6t
Xbit_r151_c248 bl[248] br[248] wl[151] vdd gnd cell_6t
Xbit_r152_c248 bl[248] br[248] wl[152] vdd gnd cell_6t
Xbit_r153_c248 bl[248] br[248] wl[153] vdd gnd cell_6t
Xbit_r154_c248 bl[248] br[248] wl[154] vdd gnd cell_6t
Xbit_r155_c248 bl[248] br[248] wl[155] vdd gnd cell_6t
Xbit_r156_c248 bl[248] br[248] wl[156] vdd gnd cell_6t
Xbit_r157_c248 bl[248] br[248] wl[157] vdd gnd cell_6t
Xbit_r158_c248 bl[248] br[248] wl[158] vdd gnd cell_6t
Xbit_r159_c248 bl[248] br[248] wl[159] vdd gnd cell_6t
Xbit_r160_c248 bl[248] br[248] wl[160] vdd gnd cell_6t
Xbit_r161_c248 bl[248] br[248] wl[161] vdd gnd cell_6t
Xbit_r162_c248 bl[248] br[248] wl[162] vdd gnd cell_6t
Xbit_r163_c248 bl[248] br[248] wl[163] vdd gnd cell_6t
Xbit_r164_c248 bl[248] br[248] wl[164] vdd gnd cell_6t
Xbit_r165_c248 bl[248] br[248] wl[165] vdd gnd cell_6t
Xbit_r166_c248 bl[248] br[248] wl[166] vdd gnd cell_6t
Xbit_r167_c248 bl[248] br[248] wl[167] vdd gnd cell_6t
Xbit_r168_c248 bl[248] br[248] wl[168] vdd gnd cell_6t
Xbit_r169_c248 bl[248] br[248] wl[169] vdd gnd cell_6t
Xbit_r170_c248 bl[248] br[248] wl[170] vdd gnd cell_6t
Xbit_r171_c248 bl[248] br[248] wl[171] vdd gnd cell_6t
Xbit_r172_c248 bl[248] br[248] wl[172] vdd gnd cell_6t
Xbit_r173_c248 bl[248] br[248] wl[173] vdd gnd cell_6t
Xbit_r174_c248 bl[248] br[248] wl[174] vdd gnd cell_6t
Xbit_r175_c248 bl[248] br[248] wl[175] vdd gnd cell_6t
Xbit_r176_c248 bl[248] br[248] wl[176] vdd gnd cell_6t
Xbit_r177_c248 bl[248] br[248] wl[177] vdd gnd cell_6t
Xbit_r178_c248 bl[248] br[248] wl[178] vdd gnd cell_6t
Xbit_r179_c248 bl[248] br[248] wl[179] vdd gnd cell_6t
Xbit_r180_c248 bl[248] br[248] wl[180] vdd gnd cell_6t
Xbit_r181_c248 bl[248] br[248] wl[181] vdd gnd cell_6t
Xbit_r182_c248 bl[248] br[248] wl[182] vdd gnd cell_6t
Xbit_r183_c248 bl[248] br[248] wl[183] vdd gnd cell_6t
Xbit_r184_c248 bl[248] br[248] wl[184] vdd gnd cell_6t
Xbit_r185_c248 bl[248] br[248] wl[185] vdd gnd cell_6t
Xbit_r186_c248 bl[248] br[248] wl[186] vdd gnd cell_6t
Xbit_r187_c248 bl[248] br[248] wl[187] vdd gnd cell_6t
Xbit_r188_c248 bl[248] br[248] wl[188] vdd gnd cell_6t
Xbit_r189_c248 bl[248] br[248] wl[189] vdd gnd cell_6t
Xbit_r190_c248 bl[248] br[248] wl[190] vdd gnd cell_6t
Xbit_r191_c248 bl[248] br[248] wl[191] vdd gnd cell_6t
Xbit_r192_c248 bl[248] br[248] wl[192] vdd gnd cell_6t
Xbit_r193_c248 bl[248] br[248] wl[193] vdd gnd cell_6t
Xbit_r194_c248 bl[248] br[248] wl[194] vdd gnd cell_6t
Xbit_r195_c248 bl[248] br[248] wl[195] vdd gnd cell_6t
Xbit_r196_c248 bl[248] br[248] wl[196] vdd gnd cell_6t
Xbit_r197_c248 bl[248] br[248] wl[197] vdd gnd cell_6t
Xbit_r198_c248 bl[248] br[248] wl[198] vdd gnd cell_6t
Xbit_r199_c248 bl[248] br[248] wl[199] vdd gnd cell_6t
Xbit_r200_c248 bl[248] br[248] wl[200] vdd gnd cell_6t
Xbit_r201_c248 bl[248] br[248] wl[201] vdd gnd cell_6t
Xbit_r202_c248 bl[248] br[248] wl[202] vdd gnd cell_6t
Xbit_r203_c248 bl[248] br[248] wl[203] vdd gnd cell_6t
Xbit_r204_c248 bl[248] br[248] wl[204] vdd gnd cell_6t
Xbit_r205_c248 bl[248] br[248] wl[205] vdd gnd cell_6t
Xbit_r206_c248 bl[248] br[248] wl[206] vdd gnd cell_6t
Xbit_r207_c248 bl[248] br[248] wl[207] vdd gnd cell_6t
Xbit_r208_c248 bl[248] br[248] wl[208] vdd gnd cell_6t
Xbit_r209_c248 bl[248] br[248] wl[209] vdd gnd cell_6t
Xbit_r210_c248 bl[248] br[248] wl[210] vdd gnd cell_6t
Xbit_r211_c248 bl[248] br[248] wl[211] vdd gnd cell_6t
Xbit_r212_c248 bl[248] br[248] wl[212] vdd gnd cell_6t
Xbit_r213_c248 bl[248] br[248] wl[213] vdd gnd cell_6t
Xbit_r214_c248 bl[248] br[248] wl[214] vdd gnd cell_6t
Xbit_r215_c248 bl[248] br[248] wl[215] vdd gnd cell_6t
Xbit_r216_c248 bl[248] br[248] wl[216] vdd gnd cell_6t
Xbit_r217_c248 bl[248] br[248] wl[217] vdd gnd cell_6t
Xbit_r218_c248 bl[248] br[248] wl[218] vdd gnd cell_6t
Xbit_r219_c248 bl[248] br[248] wl[219] vdd gnd cell_6t
Xbit_r220_c248 bl[248] br[248] wl[220] vdd gnd cell_6t
Xbit_r221_c248 bl[248] br[248] wl[221] vdd gnd cell_6t
Xbit_r222_c248 bl[248] br[248] wl[222] vdd gnd cell_6t
Xbit_r223_c248 bl[248] br[248] wl[223] vdd gnd cell_6t
Xbit_r224_c248 bl[248] br[248] wl[224] vdd gnd cell_6t
Xbit_r225_c248 bl[248] br[248] wl[225] vdd gnd cell_6t
Xbit_r226_c248 bl[248] br[248] wl[226] vdd gnd cell_6t
Xbit_r227_c248 bl[248] br[248] wl[227] vdd gnd cell_6t
Xbit_r228_c248 bl[248] br[248] wl[228] vdd gnd cell_6t
Xbit_r229_c248 bl[248] br[248] wl[229] vdd gnd cell_6t
Xbit_r230_c248 bl[248] br[248] wl[230] vdd gnd cell_6t
Xbit_r231_c248 bl[248] br[248] wl[231] vdd gnd cell_6t
Xbit_r232_c248 bl[248] br[248] wl[232] vdd gnd cell_6t
Xbit_r233_c248 bl[248] br[248] wl[233] vdd gnd cell_6t
Xbit_r234_c248 bl[248] br[248] wl[234] vdd gnd cell_6t
Xbit_r235_c248 bl[248] br[248] wl[235] vdd gnd cell_6t
Xbit_r236_c248 bl[248] br[248] wl[236] vdd gnd cell_6t
Xbit_r237_c248 bl[248] br[248] wl[237] vdd gnd cell_6t
Xbit_r238_c248 bl[248] br[248] wl[238] vdd gnd cell_6t
Xbit_r239_c248 bl[248] br[248] wl[239] vdd gnd cell_6t
Xbit_r240_c248 bl[248] br[248] wl[240] vdd gnd cell_6t
Xbit_r241_c248 bl[248] br[248] wl[241] vdd gnd cell_6t
Xbit_r242_c248 bl[248] br[248] wl[242] vdd gnd cell_6t
Xbit_r243_c248 bl[248] br[248] wl[243] vdd gnd cell_6t
Xbit_r244_c248 bl[248] br[248] wl[244] vdd gnd cell_6t
Xbit_r245_c248 bl[248] br[248] wl[245] vdd gnd cell_6t
Xbit_r246_c248 bl[248] br[248] wl[246] vdd gnd cell_6t
Xbit_r247_c248 bl[248] br[248] wl[247] vdd gnd cell_6t
Xbit_r248_c248 bl[248] br[248] wl[248] vdd gnd cell_6t
Xbit_r249_c248 bl[248] br[248] wl[249] vdd gnd cell_6t
Xbit_r250_c248 bl[248] br[248] wl[250] vdd gnd cell_6t
Xbit_r251_c248 bl[248] br[248] wl[251] vdd gnd cell_6t
Xbit_r252_c248 bl[248] br[248] wl[252] vdd gnd cell_6t
Xbit_r253_c248 bl[248] br[248] wl[253] vdd gnd cell_6t
Xbit_r254_c248 bl[248] br[248] wl[254] vdd gnd cell_6t
Xbit_r255_c248 bl[248] br[248] wl[255] vdd gnd cell_6t
Xbit_r0_c249 bl[249] br[249] wl[0] vdd gnd cell_6t
Xbit_r1_c249 bl[249] br[249] wl[1] vdd gnd cell_6t
Xbit_r2_c249 bl[249] br[249] wl[2] vdd gnd cell_6t
Xbit_r3_c249 bl[249] br[249] wl[3] vdd gnd cell_6t
Xbit_r4_c249 bl[249] br[249] wl[4] vdd gnd cell_6t
Xbit_r5_c249 bl[249] br[249] wl[5] vdd gnd cell_6t
Xbit_r6_c249 bl[249] br[249] wl[6] vdd gnd cell_6t
Xbit_r7_c249 bl[249] br[249] wl[7] vdd gnd cell_6t
Xbit_r8_c249 bl[249] br[249] wl[8] vdd gnd cell_6t
Xbit_r9_c249 bl[249] br[249] wl[9] vdd gnd cell_6t
Xbit_r10_c249 bl[249] br[249] wl[10] vdd gnd cell_6t
Xbit_r11_c249 bl[249] br[249] wl[11] vdd gnd cell_6t
Xbit_r12_c249 bl[249] br[249] wl[12] vdd gnd cell_6t
Xbit_r13_c249 bl[249] br[249] wl[13] vdd gnd cell_6t
Xbit_r14_c249 bl[249] br[249] wl[14] vdd gnd cell_6t
Xbit_r15_c249 bl[249] br[249] wl[15] vdd gnd cell_6t
Xbit_r16_c249 bl[249] br[249] wl[16] vdd gnd cell_6t
Xbit_r17_c249 bl[249] br[249] wl[17] vdd gnd cell_6t
Xbit_r18_c249 bl[249] br[249] wl[18] vdd gnd cell_6t
Xbit_r19_c249 bl[249] br[249] wl[19] vdd gnd cell_6t
Xbit_r20_c249 bl[249] br[249] wl[20] vdd gnd cell_6t
Xbit_r21_c249 bl[249] br[249] wl[21] vdd gnd cell_6t
Xbit_r22_c249 bl[249] br[249] wl[22] vdd gnd cell_6t
Xbit_r23_c249 bl[249] br[249] wl[23] vdd gnd cell_6t
Xbit_r24_c249 bl[249] br[249] wl[24] vdd gnd cell_6t
Xbit_r25_c249 bl[249] br[249] wl[25] vdd gnd cell_6t
Xbit_r26_c249 bl[249] br[249] wl[26] vdd gnd cell_6t
Xbit_r27_c249 bl[249] br[249] wl[27] vdd gnd cell_6t
Xbit_r28_c249 bl[249] br[249] wl[28] vdd gnd cell_6t
Xbit_r29_c249 bl[249] br[249] wl[29] vdd gnd cell_6t
Xbit_r30_c249 bl[249] br[249] wl[30] vdd gnd cell_6t
Xbit_r31_c249 bl[249] br[249] wl[31] vdd gnd cell_6t
Xbit_r32_c249 bl[249] br[249] wl[32] vdd gnd cell_6t
Xbit_r33_c249 bl[249] br[249] wl[33] vdd gnd cell_6t
Xbit_r34_c249 bl[249] br[249] wl[34] vdd gnd cell_6t
Xbit_r35_c249 bl[249] br[249] wl[35] vdd gnd cell_6t
Xbit_r36_c249 bl[249] br[249] wl[36] vdd gnd cell_6t
Xbit_r37_c249 bl[249] br[249] wl[37] vdd gnd cell_6t
Xbit_r38_c249 bl[249] br[249] wl[38] vdd gnd cell_6t
Xbit_r39_c249 bl[249] br[249] wl[39] vdd gnd cell_6t
Xbit_r40_c249 bl[249] br[249] wl[40] vdd gnd cell_6t
Xbit_r41_c249 bl[249] br[249] wl[41] vdd gnd cell_6t
Xbit_r42_c249 bl[249] br[249] wl[42] vdd gnd cell_6t
Xbit_r43_c249 bl[249] br[249] wl[43] vdd gnd cell_6t
Xbit_r44_c249 bl[249] br[249] wl[44] vdd gnd cell_6t
Xbit_r45_c249 bl[249] br[249] wl[45] vdd gnd cell_6t
Xbit_r46_c249 bl[249] br[249] wl[46] vdd gnd cell_6t
Xbit_r47_c249 bl[249] br[249] wl[47] vdd gnd cell_6t
Xbit_r48_c249 bl[249] br[249] wl[48] vdd gnd cell_6t
Xbit_r49_c249 bl[249] br[249] wl[49] vdd gnd cell_6t
Xbit_r50_c249 bl[249] br[249] wl[50] vdd gnd cell_6t
Xbit_r51_c249 bl[249] br[249] wl[51] vdd gnd cell_6t
Xbit_r52_c249 bl[249] br[249] wl[52] vdd gnd cell_6t
Xbit_r53_c249 bl[249] br[249] wl[53] vdd gnd cell_6t
Xbit_r54_c249 bl[249] br[249] wl[54] vdd gnd cell_6t
Xbit_r55_c249 bl[249] br[249] wl[55] vdd gnd cell_6t
Xbit_r56_c249 bl[249] br[249] wl[56] vdd gnd cell_6t
Xbit_r57_c249 bl[249] br[249] wl[57] vdd gnd cell_6t
Xbit_r58_c249 bl[249] br[249] wl[58] vdd gnd cell_6t
Xbit_r59_c249 bl[249] br[249] wl[59] vdd gnd cell_6t
Xbit_r60_c249 bl[249] br[249] wl[60] vdd gnd cell_6t
Xbit_r61_c249 bl[249] br[249] wl[61] vdd gnd cell_6t
Xbit_r62_c249 bl[249] br[249] wl[62] vdd gnd cell_6t
Xbit_r63_c249 bl[249] br[249] wl[63] vdd gnd cell_6t
Xbit_r64_c249 bl[249] br[249] wl[64] vdd gnd cell_6t
Xbit_r65_c249 bl[249] br[249] wl[65] vdd gnd cell_6t
Xbit_r66_c249 bl[249] br[249] wl[66] vdd gnd cell_6t
Xbit_r67_c249 bl[249] br[249] wl[67] vdd gnd cell_6t
Xbit_r68_c249 bl[249] br[249] wl[68] vdd gnd cell_6t
Xbit_r69_c249 bl[249] br[249] wl[69] vdd gnd cell_6t
Xbit_r70_c249 bl[249] br[249] wl[70] vdd gnd cell_6t
Xbit_r71_c249 bl[249] br[249] wl[71] vdd gnd cell_6t
Xbit_r72_c249 bl[249] br[249] wl[72] vdd gnd cell_6t
Xbit_r73_c249 bl[249] br[249] wl[73] vdd gnd cell_6t
Xbit_r74_c249 bl[249] br[249] wl[74] vdd gnd cell_6t
Xbit_r75_c249 bl[249] br[249] wl[75] vdd gnd cell_6t
Xbit_r76_c249 bl[249] br[249] wl[76] vdd gnd cell_6t
Xbit_r77_c249 bl[249] br[249] wl[77] vdd gnd cell_6t
Xbit_r78_c249 bl[249] br[249] wl[78] vdd gnd cell_6t
Xbit_r79_c249 bl[249] br[249] wl[79] vdd gnd cell_6t
Xbit_r80_c249 bl[249] br[249] wl[80] vdd gnd cell_6t
Xbit_r81_c249 bl[249] br[249] wl[81] vdd gnd cell_6t
Xbit_r82_c249 bl[249] br[249] wl[82] vdd gnd cell_6t
Xbit_r83_c249 bl[249] br[249] wl[83] vdd gnd cell_6t
Xbit_r84_c249 bl[249] br[249] wl[84] vdd gnd cell_6t
Xbit_r85_c249 bl[249] br[249] wl[85] vdd gnd cell_6t
Xbit_r86_c249 bl[249] br[249] wl[86] vdd gnd cell_6t
Xbit_r87_c249 bl[249] br[249] wl[87] vdd gnd cell_6t
Xbit_r88_c249 bl[249] br[249] wl[88] vdd gnd cell_6t
Xbit_r89_c249 bl[249] br[249] wl[89] vdd gnd cell_6t
Xbit_r90_c249 bl[249] br[249] wl[90] vdd gnd cell_6t
Xbit_r91_c249 bl[249] br[249] wl[91] vdd gnd cell_6t
Xbit_r92_c249 bl[249] br[249] wl[92] vdd gnd cell_6t
Xbit_r93_c249 bl[249] br[249] wl[93] vdd gnd cell_6t
Xbit_r94_c249 bl[249] br[249] wl[94] vdd gnd cell_6t
Xbit_r95_c249 bl[249] br[249] wl[95] vdd gnd cell_6t
Xbit_r96_c249 bl[249] br[249] wl[96] vdd gnd cell_6t
Xbit_r97_c249 bl[249] br[249] wl[97] vdd gnd cell_6t
Xbit_r98_c249 bl[249] br[249] wl[98] vdd gnd cell_6t
Xbit_r99_c249 bl[249] br[249] wl[99] vdd gnd cell_6t
Xbit_r100_c249 bl[249] br[249] wl[100] vdd gnd cell_6t
Xbit_r101_c249 bl[249] br[249] wl[101] vdd gnd cell_6t
Xbit_r102_c249 bl[249] br[249] wl[102] vdd gnd cell_6t
Xbit_r103_c249 bl[249] br[249] wl[103] vdd gnd cell_6t
Xbit_r104_c249 bl[249] br[249] wl[104] vdd gnd cell_6t
Xbit_r105_c249 bl[249] br[249] wl[105] vdd gnd cell_6t
Xbit_r106_c249 bl[249] br[249] wl[106] vdd gnd cell_6t
Xbit_r107_c249 bl[249] br[249] wl[107] vdd gnd cell_6t
Xbit_r108_c249 bl[249] br[249] wl[108] vdd gnd cell_6t
Xbit_r109_c249 bl[249] br[249] wl[109] vdd gnd cell_6t
Xbit_r110_c249 bl[249] br[249] wl[110] vdd gnd cell_6t
Xbit_r111_c249 bl[249] br[249] wl[111] vdd gnd cell_6t
Xbit_r112_c249 bl[249] br[249] wl[112] vdd gnd cell_6t
Xbit_r113_c249 bl[249] br[249] wl[113] vdd gnd cell_6t
Xbit_r114_c249 bl[249] br[249] wl[114] vdd gnd cell_6t
Xbit_r115_c249 bl[249] br[249] wl[115] vdd gnd cell_6t
Xbit_r116_c249 bl[249] br[249] wl[116] vdd gnd cell_6t
Xbit_r117_c249 bl[249] br[249] wl[117] vdd gnd cell_6t
Xbit_r118_c249 bl[249] br[249] wl[118] vdd gnd cell_6t
Xbit_r119_c249 bl[249] br[249] wl[119] vdd gnd cell_6t
Xbit_r120_c249 bl[249] br[249] wl[120] vdd gnd cell_6t
Xbit_r121_c249 bl[249] br[249] wl[121] vdd gnd cell_6t
Xbit_r122_c249 bl[249] br[249] wl[122] vdd gnd cell_6t
Xbit_r123_c249 bl[249] br[249] wl[123] vdd gnd cell_6t
Xbit_r124_c249 bl[249] br[249] wl[124] vdd gnd cell_6t
Xbit_r125_c249 bl[249] br[249] wl[125] vdd gnd cell_6t
Xbit_r126_c249 bl[249] br[249] wl[126] vdd gnd cell_6t
Xbit_r127_c249 bl[249] br[249] wl[127] vdd gnd cell_6t
Xbit_r128_c249 bl[249] br[249] wl[128] vdd gnd cell_6t
Xbit_r129_c249 bl[249] br[249] wl[129] vdd gnd cell_6t
Xbit_r130_c249 bl[249] br[249] wl[130] vdd gnd cell_6t
Xbit_r131_c249 bl[249] br[249] wl[131] vdd gnd cell_6t
Xbit_r132_c249 bl[249] br[249] wl[132] vdd gnd cell_6t
Xbit_r133_c249 bl[249] br[249] wl[133] vdd gnd cell_6t
Xbit_r134_c249 bl[249] br[249] wl[134] vdd gnd cell_6t
Xbit_r135_c249 bl[249] br[249] wl[135] vdd gnd cell_6t
Xbit_r136_c249 bl[249] br[249] wl[136] vdd gnd cell_6t
Xbit_r137_c249 bl[249] br[249] wl[137] vdd gnd cell_6t
Xbit_r138_c249 bl[249] br[249] wl[138] vdd gnd cell_6t
Xbit_r139_c249 bl[249] br[249] wl[139] vdd gnd cell_6t
Xbit_r140_c249 bl[249] br[249] wl[140] vdd gnd cell_6t
Xbit_r141_c249 bl[249] br[249] wl[141] vdd gnd cell_6t
Xbit_r142_c249 bl[249] br[249] wl[142] vdd gnd cell_6t
Xbit_r143_c249 bl[249] br[249] wl[143] vdd gnd cell_6t
Xbit_r144_c249 bl[249] br[249] wl[144] vdd gnd cell_6t
Xbit_r145_c249 bl[249] br[249] wl[145] vdd gnd cell_6t
Xbit_r146_c249 bl[249] br[249] wl[146] vdd gnd cell_6t
Xbit_r147_c249 bl[249] br[249] wl[147] vdd gnd cell_6t
Xbit_r148_c249 bl[249] br[249] wl[148] vdd gnd cell_6t
Xbit_r149_c249 bl[249] br[249] wl[149] vdd gnd cell_6t
Xbit_r150_c249 bl[249] br[249] wl[150] vdd gnd cell_6t
Xbit_r151_c249 bl[249] br[249] wl[151] vdd gnd cell_6t
Xbit_r152_c249 bl[249] br[249] wl[152] vdd gnd cell_6t
Xbit_r153_c249 bl[249] br[249] wl[153] vdd gnd cell_6t
Xbit_r154_c249 bl[249] br[249] wl[154] vdd gnd cell_6t
Xbit_r155_c249 bl[249] br[249] wl[155] vdd gnd cell_6t
Xbit_r156_c249 bl[249] br[249] wl[156] vdd gnd cell_6t
Xbit_r157_c249 bl[249] br[249] wl[157] vdd gnd cell_6t
Xbit_r158_c249 bl[249] br[249] wl[158] vdd gnd cell_6t
Xbit_r159_c249 bl[249] br[249] wl[159] vdd gnd cell_6t
Xbit_r160_c249 bl[249] br[249] wl[160] vdd gnd cell_6t
Xbit_r161_c249 bl[249] br[249] wl[161] vdd gnd cell_6t
Xbit_r162_c249 bl[249] br[249] wl[162] vdd gnd cell_6t
Xbit_r163_c249 bl[249] br[249] wl[163] vdd gnd cell_6t
Xbit_r164_c249 bl[249] br[249] wl[164] vdd gnd cell_6t
Xbit_r165_c249 bl[249] br[249] wl[165] vdd gnd cell_6t
Xbit_r166_c249 bl[249] br[249] wl[166] vdd gnd cell_6t
Xbit_r167_c249 bl[249] br[249] wl[167] vdd gnd cell_6t
Xbit_r168_c249 bl[249] br[249] wl[168] vdd gnd cell_6t
Xbit_r169_c249 bl[249] br[249] wl[169] vdd gnd cell_6t
Xbit_r170_c249 bl[249] br[249] wl[170] vdd gnd cell_6t
Xbit_r171_c249 bl[249] br[249] wl[171] vdd gnd cell_6t
Xbit_r172_c249 bl[249] br[249] wl[172] vdd gnd cell_6t
Xbit_r173_c249 bl[249] br[249] wl[173] vdd gnd cell_6t
Xbit_r174_c249 bl[249] br[249] wl[174] vdd gnd cell_6t
Xbit_r175_c249 bl[249] br[249] wl[175] vdd gnd cell_6t
Xbit_r176_c249 bl[249] br[249] wl[176] vdd gnd cell_6t
Xbit_r177_c249 bl[249] br[249] wl[177] vdd gnd cell_6t
Xbit_r178_c249 bl[249] br[249] wl[178] vdd gnd cell_6t
Xbit_r179_c249 bl[249] br[249] wl[179] vdd gnd cell_6t
Xbit_r180_c249 bl[249] br[249] wl[180] vdd gnd cell_6t
Xbit_r181_c249 bl[249] br[249] wl[181] vdd gnd cell_6t
Xbit_r182_c249 bl[249] br[249] wl[182] vdd gnd cell_6t
Xbit_r183_c249 bl[249] br[249] wl[183] vdd gnd cell_6t
Xbit_r184_c249 bl[249] br[249] wl[184] vdd gnd cell_6t
Xbit_r185_c249 bl[249] br[249] wl[185] vdd gnd cell_6t
Xbit_r186_c249 bl[249] br[249] wl[186] vdd gnd cell_6t
Xbit_r187_c249 bl[249] br[249] wl[187] vdd gnd cell_6t
Xbit_r188_c249 bl[249] br[249] wl[188] vdd gnd cell_6t
Xbit_r189_c249 bl[249] br[249] wl[189] vdd gnd cell_6t
Xbit_r190_c249 bl[249] br[249] wl[190] vdd gnd cell_6t
Xbit_r191_c249 bl[249] br[249] wl[191] vdd gnd cell_6t
Xbit_r192_c249 bl[249] br[249] wl[192] vdd gnd cell_6t
Xbit_r193_c249 bl[249] br[249] wl[193] vdd gnd cell_6t
Xbit_r194_c249 bl[249] br[249] wl[194] vdd gnd cell_6t
Xbit_r195_c249 bl[249] br[249] wl[195] vdd gnd cell_6t
Xbit_r196_c249 bl[249] br[249] wl[196] vdd gnd cell_6t
Xbit_r197_c249 bl[249] br[249] wl[197] vdd gnd cell_6t
Xbit_r198_c249 bl[249] br[249] wl[198] vdd gnd cell_6t
Xbit_r199_c249 bl[249] br[249] wl[199] vdd gnd cell_6t
Xbit_r200_c249 bl[249] br[249] wl[200] vdd gnd cell_6t
Xbit_r201_c249 bl[249] br[249] wl[201] vdd gnd cell_6t
Xbit_r202_c249 bl[249] br[249] wl[202] vdd gnd cell_6t
Xbit_r203_c249 bl[249] br[249] wl[203] vdd gnd cell_6t
Xbit_r204_c249 bl[249] br[249] wl[204] vdd gnd cell_6t
Xbit_r205_c249 bl[249] br[249] wl[205] vdd gnd cell_6t
Xbit_r206_c249 bl[249] br[249] wl[206] vdd gnd cell_6t
Xbit_r207_c249 bl[249] br[249] wl[207] vdd gnd cell_6t
Xbit_r208_c249 bl[249] br[249] wl[208] vdd gnd cell_6t
Xbit_r209_c249 bl[249] br[249] wl[209] vdd gnd cell_6t
Xbit_r210_c249 bl[249] br[249] wl[210] vdd gnd cell_6t
Xbit_r211_c249 bl[249] br[249] wl[211] vdd gnd cell_6t
Xbit_r212_c249 bl[249] br[249] wl[212] vdd gnd cell_6t
Xbit_r213_c249 bl[249] br[249] wl[213] vdd gnd cell_6t
Xbit_r214_c249 bl[249] br[249] wl[214] vdd gnd cell_6t
Xbit_r215_c249 bl[249] br[249] wl[215] vdd gnd cell_6t
Xbit_r216_c249 bl[249] br[249] wl[216] vdd gnd cell_6t
Xbit_r217_c249 bl[249] br[249] wl[217] vdd gnd cell_6t
Xbit_r218_c249 bl[249] br[249] wl[218] vdd gnd cell_6t
Xbit_r219_c249 bl[249] br[249] wl[219] vdd gnd cell_6t
Xbit_r220_c249 bl[249] br[249] wl[220] vdd gnd cell_6t
Xbit_r221_c249 bl[249] br[249] wl[221] vdd gnd cell_6t
Xbit_r222_c249 bl[249] br[249] wl[222] vdd gnd cell_6t
Xbit_r223_c249 bl[249] br[249] wl[223] vdd gnd cell_6t
Xbit_r224_c249 bl[249] br[249] wl[224] vdd gnd cell_6t
Xbit_r225_c249 bl[249] br[249] wl[225] vdd gnd cell_6t
Xbit_r226_c249 bl[249] br[249] wl[226] vdd gnd cell_6t
Xbit_r227_c249 bl[249] br[249] wl[227] vdd gnd cell_6t
Xbit_r228_c249 bl[249] br[249] wl[228] vdd gnd cell_6t
Xbit_r229_c249 bl[249] br[249] wl[229] vdd gnd cell_6t
Xbit_r230_c249 bl[249] br[249] wl[230] vdd gnd cell_6t
Xbit_r231_c249 bl[249] br[249] wl[231] vdd gnd cell_6t
Xbit_r232_c249 bl[249] br[249] wl[232] vdd gnd cell_6t
Xbit_r233_c249 bl[249] br[249] wl[233] vdd gnd cell_6t
Xbit_r234_c249 bl[249] br[249] wl[234] vdd gnd cell_6t
Xbit_r235_c249 bl[249] br[249] wl[235] vdd gnd cell_6t
Xbit_r236_c249 bl[249] br[249] wl[236] vdd gnd cell_6t
Xbit_r237_c249 bl[249] br[249] wl[237] vdd gnd cell_6t
Xbit_r238_c249 bl[249] br[249] wl[238] vdd gnd cell_6t
Xbit_r239_c249 bl[249] br[249] wl[239] vdd gnd cell_6t
Xbit_r240_c249 bl[249] br[249] wl[240] vdd gnd cell_6t
Xbit_r241_c249 bl[249] br[249] wl[241] vdd gnd cell_6t
Xbit_r242_c249 bl[249] br[249] wl[242] vdd gnd cell_6t
Xbit_r243_c249 bl[249] br[249] wl[243] vdd gnd cell_6t
Xbit_r244_c249 bl[249] br[249] wl[244] vdd gnd cell_6t
Xbit_r245_c249 bl[249] br[249] wl[245] vdd gnd cell_6t
Xbit_r246_c249 bl[249] br[249] wl[246] vdd gnd cell_6t
Xbit_r247_c249 bl[249] br[249] wl[247] vdd gnd cell_6t
Xbit_r248_c249 bl[249] br[249] wl[248] vdd gnd cell_6t
Xbit_r249_c249 bl[249] br[249] wl[249] vdd gnd cell_6t
Xbit_r250_c249 bl[249] br[249] wl[250] vdd gnd cell_6t
Xbit_r251_c249 bl[249] br[249] wl[251] vdd gnd cell_6t
Xbit_r252_c249 bl[249] br[249] wl[252] vdd gnd cell_6t
Xbit_r253_c249 bl[249] br[249] wl[253] vdd gnd cell_6t
Xbit_r254_c249 bl[249] br[249] wl[254] vdd gnd cell_6t
Xbit_r255_c249 bl[249] br[249] wl[255] vdd gnd cell_6t
Xbit_r0_c250 bl[250] br[250] wl[0] vdd gnd cell_6t
Xbit_r1_c250 bl[250] br[250] wl[1] vdd gnd cell_6t
Xbit_r2_c250 bl[250] br[250] wl[2] vdd gnd cell_6t
Xbit_r3_c250 bl[250] br[250] wl[3] vdd gnd cell_6t
Xbit_r4_c250 bl[250] br[250] wl[4] vdd gnd cell_6t
Xbit_r5_c250 bl[250] br[250] wl[5] vdd gnd cell_6t
Xbit_r6_c250 bl[250] br[250] wl[6] vdd gnd cell_6t
Xbit_r7_c250 bl[250] br[250] wl[7] vdd gnd cell_6t
Xbit_r8_c250 bl[250] br[250] wl[8] vdd gnd cell_6t
Xbit_r9_c250 bl[250] br[250] wl[9] vdd gnd cell_6t
Xbit_r10_c250 bl[250] br[250] wl[10] vdd gnd cell_6t
Xbit_r11_c250 bl[250] br[250] wl[11] vdd gnd cell_6t
Xbit_r12_c250 bl[250] br[250] wl[12] vdd gnd cell_6t
Xbit_r13_c250 bl[250] br[250] wl[13] vdd gnd cell_6t
Xbit_r14_c250 bl[250] br[250] wl[14] vdd gnd cell_6t
Xbit_r15_c250 bl[250] br[250] wl[15] vdd gnd cell_6t
Xbit_r16_c250 bl[250] br[250] wl[16] vdd gnd cell_6t
Xbit_r17_c250 bl[250] br[250] wl[17] vdd gnd cell_6t
Xbit_r18_c250 bl[250] br[250] wl[18] vdd gnd cell_6t
Xbit_r19_c250 bl[250] br[250] wl[19] vdd gnd cell_6t
Xbit_r20_c250 bl[250] br[250] wl[20] vdd gnd cell_6t
Xbit_r21_c250 bl[250] br[250] wl[21] vdd gnd cell_6t
Xbit_r22_c250 bl[250] br[250] wl[22] vdd gnd cell_6t
Xbit_r23_c250 bl[250] br[250] wl[23] vdd gnd cell_6t
Xbit_r24_c250 bl[250] br[250] wl[24] vdd gnd cell_6t
Xbit_r25_c250 bl[250] br[250] wl[25] vdd gnd cell_6t
Xbit_r26_c250 bl[250] br[250] wl[26] vdd gnd cell_6t
Xbit_r27_c250 bl[250] br[250] wl[27] vdd gnd cell_6t
Xbit_r28_c250 bl[250] br[250] wl[28] vdd gnd cell_6t
Xbit_r29_c250 bl[250] br[250] wl[29] vdd gnd cell_6t
Xbit_r30_c250 bl[250] br[250] wl[30] vdd gnd cell_6t
Xbit_r31_c250 bl[250] br[250] wl[31] vdd gnd cell_6t
Xbit_r32_c250 bl[250] br[250] wl[32] vdd gnd cell_6t
Xbit_r33_c250 bl[250] br[250] wl[33] vdd gnd cell_6t
Xbit_r34_c250 bl[250] br[250] wl[34] vdd gnd cell_6t
Xbit_r35_c250 bl[250] br[250] wl[35] vdd gnd cell_6t
Xbit_r36_c250 bl[250] br[250] wl[36] vdd gnd cell_6t
Xbit_r37_c250 bl[250] br[250] wl[37] vdd gnd cell_6t
Xbit_r38_c250 bl[250] br[250] wl[38] vdd gnd cell_6t
Xbit_r39_c250 bl[250] br[250] wl[39] vdd gnd cell_6t
Xbit_r40_c250 bl[250] br[250] wl[40] vdd gnd cell_6t
Xbit_r41_c250 bl[250] br[250] wl[41] vdd gnd cell_6t
Xbit_r42_c250 bl[250] br[250] wl[42] vdd gnd cell_6t
Xbit_r43_c250 bl[250] br[250] wl[43] vdd gnd cell_6t
Xbit_r44_c250 bl[250] br[250] wl[44] vdd gnd cell_6t
Xbit_r45_c250 bl[250] br[250] wl[45] vdd gnd cell_6t
Xbit_r46_c250 bl[250] br[250] wl[46] vdd gnd cell_6t
Xbit_r47_c250 bl[250] br[250] wl[47] vdd gnd cell_6t
Xbit_r48_c250 bl[250] br[250] wl[48] vdd gnd cell_6t
Xbit_r49_c250 bl[250] br[250] wl[49] vdd gnd cell_6t
Xbit_r50_c250 bl[250] br[250] wl[50] vdd gnd cell_6t
Xbit_r51_c250 bl[250] br[250] wl[51] vdd gnd cell_6t
Xbit_r52_c250 bl[250] br[250] wl[52] vdd gnd cell_6t
Xbit_r53_c250 bl[250] br[250] wl[53] vdd gnd cell_6t
Xbit_r54_c250 bl[250] br[250] wl[54] vdd gnd cell_6t
Xbit_r55_c250 bl[250] br[250] wl[55] vdd gnd cell_6t
Xbit_r56_c250 bl[250] br[250] wl[56] vdd gnd cell_6t
Xbit_r57_c250 bl[250] br[250] wl[57] vdd gnd cell_6t
Xbit_r58_c250 bl[250] br[250] wl[58] vdd gnd cell_6t
Xbit_r59_c250 bl[250] br[250] wl[59] vdd gnd cell_6t
Xbit_r60_c250 bl[250] br[250] wl[60] vdd gnd cell_6t
Xbit_r61_c250 bl[250] br[250] wl[61] vdd gnd cell_6t
Xbit_r62_c250 bl[250] br[250] wl[62] vdd gnd cell_6t
Xbit_r63_c250 bl[250] br[250] wl[63] vdd gnd cell_6t
Xbit_r64_c250 bl[250] br[250] wl[64] vdd gnd cell_6t
Xbit_r65_c250 bl[250] br[250] wl[65] vdd gnd cell_6t
Xbit_r66_c250 bl[250] br[250] wl[66] vdd gnd cell_6t
Xbit_r67_c250 bl[250] br[250] wl[67] vdd gnd cell_6t
Xbit_r68_c250 bl[250] br[250] wl[68] vdd gnd cell_6t
Xbit_r69_c250 bl[250] br[250] wl[69] vdd gnd cell_6t
Xbit_r70_c250 bl[250] br[250] wl[70] vdd gnd cell_6t
Xbit_r71_c250 bl[250] br[250] wl[71] vdd gnd cell_6t
Xbit_r72_c250 bl[250] br[250] wl[72] vdd gnd cell_6t
Xbit_r73_c250 bl[250] br[250] wl[73] vdd gnd cell_6t
Xbit_r74_c250 bl[250] br[250] wl[74] vdd gnd cell_6t
Xbit_r75_c250 bl[250] br[250] wl[75] vdd gnd cell_6t
Xbit_r76_c250 bl[250] br[250] wl[76] vdd gnd cell_6t
Xbit_r77_c250 bl[250] br[250] wl[77] vdd gnd cell_6t
Xbit_r78_c250 bl[250] br[250] wl[78] vdd gnd cell_6t
Xbit_r79_c250 bl[250] br[250] wl[79] vdd gnd cell_6t
Xbit_r80_c250 bl[250] br[250] wl[80] vdd gnd cell_6t
Xbit_r81_c250 bl[250] br[250] wl[81] vdd gnd cell_6t
Xbit_r82_c250 bl[250] br[250] wl[82] vdd gnd cell_6t
Xbit_r83_c250 bl[250] br[250] wl[83] vdd gnd cell_6t
Xbit_r84_c250 bl[250] br[250] wl[84] vdd gnd cell_6t
Xbit_r85_c250 bl[250] br[250] wl[85] vdd gnd cell_6t
Xbit_r86_c250 bl[250] br[250] wl[86] vdd gnd cell_6t
Xbit_r87_c250 bl[250] br[250] wl[87] vdd gnd cell_6t
Xbit_r88_c250 bl[250] br[250] wl[88] vdd gnd cell_6t
Xbit_r89_c250 bl[250] br[250] wl[89] vdd gnd cell_6t
Xbit_r90_c250 bl[250] br[250] wl[90] vdd gnd cell_6t
Xbit_r91_c250 bl[250] br[250] wl[91] vdd gnd cell_6t
Xbit_r92_c250 bl[250] br[250] wl[92] vdd gnd cell_6t
Xbit_r93_c250 bl[250] br[250] wl[93] vdd gnd cell_6t
Xbit_r94_c250 bl[250] br[250] wl[94] vdd gnd cell_6t
Xbit_r95_c250 bl[250] br[250] wl[95] vdd gnd cell_6t
Xbit_r96_c250 bl[250] br[250] wl[96] vdd gnd cell_6t
Xbit_r97_c250 bl[250] br[250] wl[97] vdd gnd cell_6t
Xbit_r98_c250 bl[250] br[250] wl[98] vdd gnd cell_6t
Xbit_r99_c250 bl[250] br[250] wl[99] vdd gnd cell_6t
Xbit_r100_c250 bl[250] br[250] wl[100] vdd gnd cell_6t
Xbit_r101_c250 bl[250] br[250] wl[101] vdd gnd cell_6t
Xbit_r102_c250 bl[250] br[250] wl[102] vdd gnd cell_6t
Xbit_r103_c250 bl[250] br[250] wl[103] vdd gnd cell_6t
Xbit_r104_c250 bl[250] br[250] wl[104] vdd gnd cell_6t
Xbit_r105_c250 bl[250] br[250] wl[105] vdd gnd cell_6t
Xbit_r106_c250 bl[250] br[250] wl[106] vdd gnd cell_6t
Xbit_r107_c250 bl[250] br[250] wl[107] vdd gnd cell_6t
Xbit_r108_c250 bl[250] br[250] wl[108] vdd gnd cell_6t
Xbit_r109_c250 bl[250] br[250] wl[109] vdd gnd cell_6t
Xbit_r110_c250 bl[250] br[250] wl[110] vdd gnd cell_6t
Xbit_r111_c250 bl[250] br[250] wl[111] vdd gnd cell_6t
Xbit_r112_c250 bl[250] br[250] wl[112] vdd gnd cell_6t
Xbit_r113_c250 bl[250] br[250] wl[113] vdd gnd cell_6t
Xbit_r114_c250 bl[250] br[250] wl[114] vdd gnd cell_6t
Xbit_r115_c250 bl[250] br[250] wl[115] vdd gnd cell_6t
Xbit_r116_c250 bl[250] br[250] wl[116] vdd gnd cell_6t
Xbit_r117_c250 bl[250] br[250] wl[117] vdd gnd cell_6t
Xbit_r118_c250 bl[250] br[250] wl[118] vdd gnd cell_6t
Xbit_r119_c250 bl[250] br[250] wl[119] vdd gnd cell_6t
Xbit_r120_c250 bl[250] br[250] wl[120] vdd gnd cell_6t
Xbit_r121_c250 bl[250] br[250] wl[121] vdd gnd cell_6t
Xbit_r122_c250 bl[250] br[250] wl[122] vdd gnd cell_6t
Xbit_r123_c250 bl[250] br[250] wl[123] vdd gnd cell_6t
Xbit_r124_c250 bl[250] br[250] wl[124] vdd gnd cell_6t
Xbit_r125_c250 bl[250] br[250] wl[125] vdd gnd cell_6t
Xbit_r126_c250 bl[250] br[250] wl[126] vdd gnd cell_6t
Xbit_r127_c250 bl[250] br[250] wl[127] vdd gnd cell_6t
Xbit_r128_c250 bl[250] br[250] wl[128] vdd gnd cell_6t
Xbit_r129_c250 bl[250] br[250] wl[129] vdd gnd cell_6t
Xbit_r130_c250 bl[250] br[250] wl[130] vdd gnd cell_6t
Xbit_r131_c250 bl[250] br[250] wl[131] vdd gnd cell_6t
Xbit_r132_c250 bl[250] br[250] wl[132] vdd gnd cell_6t
Xbit_r133_c250 bl[250] br[250] wl[133] vdd gnd cell_6t
Xbit_r134_c250 bl[250] br[250] wl[134] vdd gnd cell_6t
Xbit_r135_c250 bl[250] br[250] wl[135] vdd gnd cell_6t
Xbit_r136_c250 bl[250] br[250] wl[136] vdd gnd cell_6t
Xbit_r137_c250 bl[250] br[250] wl[137] vdd gnd cell_6t
Xbit_r138_c250 bl[250] br[250] wl[138] vdd gnd cell_6t
Xbit_r139_c250 bl[250] br[250] wl[139] vdd gnd cell_6t
Xbit_r140_c250 bl[250] br[250] wl[140] vdd gnd cell_6t
Xbit_r141_c250 bl[250] br[250] wl[141] vdd gnd cell_6t
Xbit_r142_c250 bl[250] br[250] wl[142] vdd gnd cell_6t
Xbit_r143_c250 bl[250] br[250] wl[143] vdd gnd cell_6t
Xbit_r144_c250 bl[250] br[250] wl[144] vdd gnd cell_6t
Xbit_r145_c250 bl[250] br[250] wl[145] vdd gnd cell_6t
Xbit_r146_c250 bl[250] br[250] wl[146] vdd gnd cell_6t
Xbit_r147_c250 bl[250] br[250] wl[147] vdd gnd cell_6t
Xbit_r148_c250 bl[250] br[250] wl[148] vdd gnd cell_6t
Xbit_r149_c250 bl[250] br[250] wl[149] vdd gnd cell_6t
Xbit_r150_c250 bl[250] br[250] wl[150] vdd gnd cell_6t
Xbit_r151_c250 bl[250] br[250] wl[151] vdd gnd cell_6t
Xbit_r152_c250 bl[250] br[250] wl[152] vdd gnd cell_6t
Xbit_r153_c250 bl[250] br[250] wl[153] vdd gnd cell_6t
Xbit_r154_c250 bl[250] br[250] wl[154] vdd gnd cell_6t
Xbit_r155_c250 bl[250] br[250] wl[155] vdd gnd cell_6t
Xbit_r156_c250 bl[250] br[250] wl[156] vdd gnd cell_6t
Xbit_r157_c250 bl[250] br[250] wl[157] vdd gnd cell_6t
Xbit_r158_c250 bl[250] br[250] wl[158] vdd gnd cell_6t
Xbit_r159_c250 bl[250] br[250] wl[159] vdd gnd cell_6t
Xbit_r160_c250 bl[250] br[250] wl[160] vdd gnd cell_6t
Xbit_r161_c250 bl[250] br[250] wl[161] vdd gnd cell_6t
Xbit_r162_c250 bl[250] br[250] wl[162] vdd gnd cell_6t
Xbit_r163_c250 bl[250] br[250] wl[163] vdd gnd cell_6t
Xbit_r164_c250 bl[250] br[250] wl[164] vdd gnd cell_6t
Xbit_r165_c250 bl[250] br[250] wl[165] vdd gnd cell_6t
Xbit_r166_c250 bl[250] br[250] wl[166] vdd gnd cell_6t
Xbit_r167_c250 bl[250] br[250] wl[167] vdd gnd cell_6t
Xbit_r168_c250 bl[250] br[250] wl[168] vdd gnd cell_6t
Xbit_r169_c250 bl[250] br[250] wl[169] vdd gnd cell_6t
Xbit_r170_c250 bl[250] br[250] wl[170] vdd gnd cell_6t
Xbit_r171_c250 bl[250] br[250] wl[171] vdd gnd cell_6t
Xbit_r172_c250 bl[250] br[250] wl[172] vdd gnd cell_6t
Xbit_r173_c250 bl[250] br[250] wl[173] vdd gnd cell_6t
Xbit_r174_c250 bl[250] br[250] wl[174] vdd gnd cell_6t
Xbit_r175_c250 bl[250] br[250] wl[175] vdd gnd cell_6t
Xbit_r176_c250 bl[250] br[250] wl[176] vdd gnd cell_6t
Xbit_r177_c250 bl[250] br[250] wl[177] vdd gnd cell_6t
Xbit_r178_c250 bl[250] br[250] wl[178] vdd gnd cell_6t
Xbit_r179_c250 bl[250] br[250] wl[179] vdd gnd cell_6t
Xbit_r180_c250 bl[250] br[250] wl[180] vdd gnd cell_6t
Xbit_r181_c250 bl[250] br[250] wl[181] vdd gnd cell_6t
Xbit_r182_c250 bl[250] br[250] wl[182] vdd gnd cell_6t
Xbit_r183_c250 bl[250] br[250] wl[183] vdd gnd cell_6t
Xbit_r184_c250 bl[250] br[250] wl[184] vdd gnd cell_6t
Xbit_r185_c250 bl[250] br[250] wl[185] vdd gnd cell_6t
Xbit_r186_c250 bl[250] br[250] wl[186] vdd gnd cell_6t
Xbit_r187_c250 bl[250] br[250] wl[187] vdd gnd cell_6t
Xbit_r188_c250 bl[250] br[250] wl[188] vdd gnd cell_6t
Xbit_r189_c250 bl[250] br[250] wl[189] vdd gnd cell_6t
Xbit_r190_c250 bl[250] br[250] wl[190] vdd gnd cell_6t
Xbit_r191_c250 bl[250] br[250] wl[191] vdd gnd cell_6t
Xbit_r192_c250 bl[250] br[250] wl[192] vdd gnd cell_6t
Xbit_r193_c250 bl[250] br[250] wl[193] vdd gnd cell_6t
Xbit_r194_c250 bl[250] br[250] wl[194] vdd gnd cell_6t
Xbit_r195_c250 bl[250] br[250] wl[195] vdd gnd cell_6t
Xbit_r196_c250 bl[250] br[250] wl[196] vdd gnd cell_6t
Xbit_r197_c250 bl[250] br[250] wl[197] vdd gnd cell_6t
Xbit_r198_c250 bl[250] br[250] wl[198] vdd gnd cell_6t
Xbit_r199_c250 bl[250] br[250] wl[199] vdd gnd cell_6t
Xbit_r200_c250 bl[250] br[250] wl[200] vdd gnd cell_6t
Xbit_r201_c250 bl[250] br[250] wl[201] vdd gnd cell_6t
Xbit_r202_c250 bl[250] br[250] wl[202] vdd gnd cell_6t
Xbit_r203_c250 bl[250] br[250] wl[203] vdd gnd cell_6t
Xbit_r204_c250 bl[250] br[250] wl[204] vdd gnd cell_6t
Xbit_r205_c250 bl[250] br[250] wl[205] vdd gnd cell_6t
Xbit_r206_c250 bl[250] br[250] wl[206] vdd gnd cell_6t
Xbit_r207_c250 bl[250] br[250] wl[207] vdd gnd cell_6t
Xbit_r208_c250 bl[250] br[250] wl[208] vdd gnd cell_6t
Xbit_r209_c250 bl[250] br[250] wl[209] vdd gnd cell_6t
Xbit_r210_c250 bl[250] br[250] wl[210] vdd gnd cell_6t
Xbit_r211_c250 bl[250] br[250] wl[211] vdd gnd cell_6t
Xbit_r212_c250 bl[250] br[250] wl[212] vdd gnd cell_6t
Xbit_r213_c250 bl[250] br[250] wl[213] vdd gnd cell_6t
Xbit_r214_c250 bl[250] br[250] wl[214] vdd gnd cell_6t
Xbit_r215_c250 bl[250] br[250] wl[215] vdd gnd cell_6t
Xbit_r216_c250 bl[250] br[250] wl[216] vdd gnd cell_6t
Xbit_r217_c250 bl[250] br[250] wl[217] vdd gnd cell_6t
Xbit_r218_c250 bl[250] br[250] wl[218] vdd gnd cell_6t
Xbit_r219_c250 bl[250] br[250] wl[219] vdd gnd cell_6t
Xbit_r220_c250 bl[250] br[250] wl[220] vdd gnd cell_6t
Xbit_r221_c250 bl[250] br[250] wl[221] vdd gnd cell_6t
Xbit_r222_c250 bl[250] br[250] wl[222] vdd gnd cell_6t
Xbit_r223_c250 bl[250] br[250] wl[223] vdd gnd cell_6t
Xbit_r224_c250 bl[250] br[250] wl[224] vdd gnd cell_6t
Xbit_r225_c250 bl[250] br[250] wl[225] vdd gnd cell_6t
Xbit_r226_c250 bl[250] br[250] wl[226] vdd gnd cell_6t
Xbit_r227_c250 bl[250] br[250] wl[227] vdd gnd cell_6t
Xbit_r228_c250 bl[250] br[250] wl[228] vdd gnd cell_6t
Xbit_r229_c250 bl[250] br[250] wl[229] vdd gnd cell_6t
Xbit_r230_c250 bl[250] br[250] wl[230] vdd gnd cell_6t
Xbit_r231_c250 bl[250] br[250] wl[231] vdd gnd cell_6t
Xbit_r232_c250 bl[250] br[250] wl[232] vdd gnd cell_6t
Xbit_r233_c250 bl[250] br[250] wl[233] vdd gnd cell_6t
Xbit_r234_c250 bl[250] br[250] wl[234] vdd gnd cell_6t
Xbit_r235_c250 bl[250] br[250] wl[235] vdd gnd cell_6t
Xbit_r236_c250 bl[250] br[250] wl[236] vdd gnd cell_6t
Xbit_r237_c250 bl[250] br[250] wl[237] vdd gnd cell_6t
Xbit_r238_c250 bl[250] br[250] wl[238] vdd gnd cell_6t
Xbit_r239_c250 bl[250] br[250] wl[239] vdd gnd cell_6t
Xbit_r240_c250 bl[250] br[250] wl[240] vdd gnd cell_6t
Xbit_r241_c250 bl[250] br[250] wl[241] vdd gnd cell_6t
Xbit_r242_c250 bl[250] br[250] wl[242] vdd gnd cell_6t
Xbit_r243_c250 bl[250] br[250] wl[243] vdd gnd cell_6t
Xbit_r244_c250 bl[250] br[250] wl[244] vdd gnd cell_6t
Xbit_r245_c250 bl[250] br[250] wl[245] vdd gnd cell_6t
Xbit_r246_c250 bl[250] br[250] wl[246] vdd gnd cell_6t
Xbit_r247_c250 bl[250] br[250] wl[247] vdd gnd cell_6t
Xbit_r248_c250 bl[250] br[250] wl[248] vdd gnd cell_6t
Xbit_r249_c250 bl[250] br[250] wl[249] vdd gnd cell_6t
Xbit_r250_c250 bl[250] br[250] wl[250] vdd gnd cell_6t
Xbit_r251_c250 bl[250] br[250] wl[251] vdd gnd cell_6t
Xbit_r252_c250 bl[250] br[250] wl[252] vdd gnd cell_6t
Xbit_r253_c250 bl[250] br[250] wl[253] vdd gnd cell_6t
Xbit_r254_c250 bl[250] br[250] wl[254] vdd gnd cell_6t
Xbit_r255_c250 bl[250] br[250] wl[255] vdd gnd cell_6t
Xbit_r0_c251 bl[251] br[251] wl[0] vdd gnd cell_6t
Xbit_r1_c251 bl[251] br[251] wl[1] vdd gnd cell_6t
Xbit_r2_c251 bl[251] br[251] wl[2] vdd gnd cell_6t
Xbit_r3_c251 bl[251] br[251] wl[3] vdd gnd cell_6t
Xbit_r4_c251 bl[251] br[251] wl[4] vdd gnd cell_6t
Xbit_r5_c251 bl[251] br[251] wl[5] vdd gnd cell_6t
Xbit_r6_c251 bl[251] br[251] wl[6] vdd gnd cell_6t
Xbit_r7_c251 bl[251] br[251] wl[7] vdd gnd cell_6t
Xbit_r8_c251 bl[251] br[251] wl[8] vdd gnd cell_6t
Xbit_r9_c251 bl[251] br[251] wl[9] vdd gnd cell_6t
Xbit_r10_c251 bl[251] br[251] wl[10] vdd gnd cell_6t
Xbit_r11_c251 bl[251] br[251] wl[11] vdd gnd cell_6t
Xbit_r12_c251 bl[251] br[251] wl[12] vdd gnd cell_6t
Xbit_r13_c251 bl[251] br[251] wl[13] vdd gnd cell_6t
Xbit_r14_c251 bl[251] br[251] wl[14] vdd gnd cell_6t
Xbit_r15_c251 bl[251] br[251] wl[15] vdd gnd cell_6t
Xbit_r16_c251 bl[251] br[251] wl[16] vdd gnd cell_6t
Xbit_r17_c251 bl[251] br[251] wl[17] vdd gnd cell_6t
Xbit_r18_c251 bl[251] br[251] wl[18] vdd gnd cell_6t
Xbit_r19_c251 bl[251] br[251] wl[19] vdd gnd cell_6t
Xbit_r20_c251 bl[251] br[251] wl[20] vdd gnd cell_6t
Xbit_r21_c251 bl[251] br[251] wl[21] vdd gnd cell_6t
Xbit_r22_c251 bl[251] br[251] wl[22] vdd gnd cell_6t
Xbit_r23_c251 bl[251] br[251] wl[23] vdd gnd cell_6t
Xbit_r24_c251 bl[251] br[251] wl[24] vdd gnd cell_6t
Xbit_r25_c251 bl[251] br[251] wl[25] vdd gnd cell_6t
Xbit_r26_c251 bl[251] br[251] wl[26] vdd gnd cell_6t
Xbit_r27_c251 bl[251] br[251] wl[27] vdd gnd cell_6t
Xbit_r28_c251 bl[251] br[251] wl[28] vdd gnd cell_6t
Xbit_r29_c251 bl[251] br[251] wl[29] vdd gnd cell_6t
Xbit_r30_c251 bl[251] br[251] wl[30] vdd gnd cell_6t
Xbit_r31_c251 bl[251] br[251] wl[31] vdd gnd cell_6t
Xbit_r32_c251 bl[251] br[251] wl[32] vdd gnd cell_6t
Xbit_r33_c251 bl[251] br[251] wl[33] vdd gnd cell_6t
Xbit_r34_c251 bl[251] br[251] wl[34] vdd gnd cell_6t
Xbit_r35_c251 bl[251] br[251] wl[35] vdd gnd cell_6t
Xbit_r36_c251 bl[251] br[251] wl[36] vdd gnd cell_6t
Xbit_r37_c251 bl[251] br[251] wl[37] vdd gnd cell_6t
Xbit_r38_c251 bl[251] br[251] wl[38] vdd gnd cell_6t
Xbit_r39_c251 bl[251] br[251] wl[39] vdd gnd cell_6t
Xbit_r40_c251 bl[251] br[251] wl[40] vdd gnd cell_6t
Xbit_r41_c251 bl[251] br[251] wl[41] vdd gnd cell_6t
Xbit_r42_c251 bl[251] br[251] wl[42] vdd gnd cell_6t
Xbit_r43_c251 bl[251] br[251] wl[43] vdd gnd cell_6t
Xbit_r44_c251 bl[251] br[251] wl[44] vdd gnd cell_6t
Xbit_r45_c251 bl[251] br[251] wl[45] vdd gnd cell_6t
Xbit_r46_c251 bl[251] br[251] wl[46] vdd gnd cell_6t
Xbit_r47_c251 bl[251] br[251] wl[47] vdd gnd cell_6t
Xbit_r48_c251 bl[251] br[251] wl[48] vdd gnd cell_6t
Xbit_r49_c251 bl[251] br[251] wl[49] vdd gnd cell_6t
Xbit_r50_c251 bl[251] br[251] wl[50] vdd gnd cell_6t
Xbit_r51_c251 bl[251] br[251] wl[51] vdd gnd cell_6t
Xbit_r52_c251 bl[251] br[251] wl[52] vdd gnd cell_6t
Xbit_r53_c251 bl[251] br[251] wl[53] vdd gnd cell_6t
Xbit_r54_c251 bl[251] br[251] wl[54] vdd gnd cell_6t
Xbit_r55_c251 bl[251] br[251] wl[55] vdd gnd cell_6t
Xbit_r56_c251 bl[251] br[251] wl[56] vdd gnd cell_6t
Xbit_r57_c251 bl[251] br[251] wl[57] vdd gnd cell_6t
Xbit_r58_c251 bl[251] br[251] wl[58] vdd gnd cell_6t
Xbit_r59_c251 bl[251] br[251] wl[59] vdd gnd cell_6t
Xbit_r60_c251 bl[251] br[251] wl[60] vdd gnd cell_6t
Xbit_r61_c251 bl[251] br[251] wl[61] vdd gnd cell_6t
Xbit_r62_c251 bl[251] br[251] wl[62] vdd gnd cell_6t
Xbit_r63_c251 bl[251] br[251] wl[63] vdd gnd cell_6t
Xbit_r64_c251 bl[251] br[251] wl[64] vdd gnd cell_6t
Xbit_r65_c251 bl[251] br[251] wl[65] vdd gnd cell_6t
Xbit_r66_c251 bl[251] br[251] wl[66] vdd gnd cell_6t
Xbit_r67_c251 bl[251] br[251] wl[67] vdd gnd cell_6t
Xbit_r68_c251 bl[251] br[251] wl[68] vdd gnd cell_6t
Xbit_r69_c251 bl[251] br[251] wl[69] vdd gnd cell_6t
Xbit_r70_c251 bl[251] br[251] wl[70] vdd gnd cell_6t
Xbit_r71_c251 bl[251] br[251] wl[71] vdd gnd cell_6t
Xbit_r72_c251 bl[251] br[251] wl[72] vdd gnd cell_6t
Xbit_r73_c251 bl[251] br[251] wl[73] vdd gnd cell_6t
Xbit_r74_c251 bl[251] br[251] wl[74] vdd gnd cell_6t
Xbit_r75_c251 bl[251] br[251] wl[75] vdd gnd cell_6t
Xbit_r76_c251 bl[251] br[251] wl[76] vdd gnd cell_6t
Xbit_r77_c251 bl[251] br[251] wl[77] vdd gnd cell_6t
Xbit_r78_c251 bl[251] br[251] wl[78] vdd gnd cell_6t
Xbit_r79_c251 bl[251] br[251] wl[79] vdd gnd cell_6t
Xbit_r80_c251 bl[251] br[251] wl[80] vdd gnd cell_6t
Xbit_r81_c251 bl[251] br[251] wl[81] vdd gnd cell_6t
Xbit_r82_c251 bl[251] br[251] wl[82] vdd gnd cell_6t
Xbit_r83_c251 bl[251] br[251] wl[83] vdd gnd cell_6t
Xbit_r84_c251 bl[251] br[251] wl[84] vdd gnd cell_6t
Xbit_r85_c251 bl[251] br[251] wl[85] vdd gnd cell_6t
Xbit_r86_c251 bl[251] br[251] wl[86] vdd gnd cell_6t
Xbit_r87_c251 bl[251] br[251] wl[87] vdd gnd cell_6t
Xbit_r88_c251 bl[251] br[251] wl[88] vdd gnd cell_6t
Xbit_r89_c251 bl[251] br[251] wl[89] vdd gnd cell_6t
Xbit_r90_c251 bl[251] br[251] wl[90] vdd gnd cell_6t
Xbit_r91_c251 bl[251] br[251] wl[91] vdd gnd cell_6t
Xbit_r92_c251 bl[251] br[251] wl[92] vdd gnd cell_6t
Xbit_r93_c251 bl[251] br[251] wl[93] vdd gnd cell_6t
Xbit_r94_c251 bl[251] br[251] wl[94] vdd gnd cell_6t
Xbit_r95_c251 bl[251] br[251] wl[95] vdd gnd cell_6t
Xbit_r96_c251 bl[251] br[251] wl[96] vdd gnd cell_6t
Xbit_r97_c251 bl[251] br[251] wl[97] vdd gnd cell_6t
Xbit_r98_c251 bl[251] br[251] wl[98] vdd gnd cell_6t
Xbit_r99_c251 bl[251] br[251] wl[99] vdd gnd cell_6t
Xbit_r100_c251 bl[251] br[251] wl[100] vdd gnd cell_6t
Xbit_r101_c251 bl[251] br[251] wl[101] vdd gnd cell_6t
Xbit_r102_c251 bl[251] br[251] wl[102] vdd gnd cell_6t
Xbit_r103_c251 bl[251] br[251] wl[103] vdd gnd cell_6t
Xbit_r104_c251 bl[251] br[251] wl[104] vdd gnd cell_6t
Xbit_r105_c251 bl[251] br[251] wl[105] vdd gnd cell_6t
Xbit_r106_c251 bl[251] br[251] wl[106] vdd gnd cell_6t
Xbit_r107_c251 bl[251] br[251] wl[107] vdd gnd cell_6t
Xbit_r108_c251 bl[251] br[251] wl[108] vdd gnd cell_6t
Xbit_r109_c251 bl[251] br[251] wl[109] vdd gnd cell_6t
Xbit_r110_c251 bl[251] br[251] wl[110] vdd gnd cell_6t
Xbit_r111_c251 bl[251] br[251] wl[111] vdd gnd cell_6t
Xbit_r112_c251 bl[251] br[251] wl[112] vdd gnd cell_6t
Xbit_r113_c251 bl[251] br[251] wl[113] vdd gnd cell_6t
Xbit_r114_c251 bl[251] br[251] wl[114] vdd gnd cell_6t
Xbit_r115_c251 bl[251] br[251] wl[115] vdd gnd cell_6t
Xbit_r116_c251 bl[251] br[251] wl[116] vdd gnd cell_6t
Xbit_r117_c251 bl[251] br[251] wl[117] vdd gnd cell_6t
Xbit_r118_c251 bl[251] br[251] wl[118] vdd gnd cell_6t
Xbit_r119_c251 bl[251] br[251] wl[119] vdd gnd cell_6t
Xbit_r120_c251 bl[251] br[251] wl[120] vdd gnd cell_6t
Xbit_r121_c251 bl[251] br[251] wl[121] vdd gnd cell_6t
Xbit_r122_c251 bl[251] br[251] wl[122] vdd gnd cell_6t
Xbit_r123_c251 bl[251] br[251] wl[123] vdd gnd cell_6t
Xbit_r124_c251 bl[251] br[251] wl[124] vdd gnd cell_6t
Xbit_r125_c251 bl[251] br[251] wl[125] vdd gnd cell_6t
Xbit_r126_c251 bl[251] br[251] wl[126] vdd gnd cell_6t
Xbit_r127_c251 bl[251] br[251] wl[127] vdd gnd cell_6t
Xbit_r128_c251 bl[251] br[251] wl[128] vdd gnd cell_6t
Xbit_r129_c251 bl[251] br[251] wl[129] vdd gnd cell_6t
Xbit_r130_c251 bl[251] br[251] wl[130] vdd gnd cell_6t
Xbit_r131_c251 bl[251] br[251] wl[131] vdd gnd cell_6t
Xbit_r132_c251 bl[251] br[251] wl[132] vdd gnd cell_6t
Xbit_r133_c251 bl[251] br[251] wl[133] vdd gnd cell_6t
Xbit_r134_c251 bl[251] br[251] wl[134] vdd gnd cell_6t
Xbit_r135_c251 bl[251] br[251] wl[135] vdd gnd cell_6t
Xbit_r136_c251 bl[251] br[251] wl[136] vdd gnd cell_6t
Xbit_r137_c251 bl[251] br[251] wl[137] vdd gnd cell_6t
Xbit_r138_c251 bl[251] br[251] wl[138] vdd gnd cell_6t
Xbit_r139_c251 bl[251] br[251] wl[139] vdd gnd cell_6t
Xbit_r140_c251 bl[251] br[251] wl[140] vdd gnd cell_6t
Xbit_r141_c251 bl[251] br[251] wl[141] vdd gnd cell_6t
Xbit_r142_c251 bl[251] br[251] wl[142] vdd gnd cell_6t
Xbit_r143_c251 bl[251] br[251] wl[143] vdd gnd cell_6t
Xbit_r144_c251 bl[251] br[251] wl[144] vdd gnd cell_6t
Xbit_r145_c251 bl[251] br[251] wl[145] vdd gnd cell_6t
Xbit_r146_c251 bl[251] br[251] wl[146] vdd gnd cell_6t
Xbit_r147_c251 bl[251] br[251] wl[147] vdd gnd cell_6t
Xbit_r148_c251 bl[251] br[251] wl[148] vdd gnd cell_6t
Xbit_r149_c251 bl[251] br[251] wl[149] vdd gnd cell_6t
Xbit_r150_c251 bl[251] br[251] wl[150] vdd gnd cell_6t
Xbit_r151_c251 bl[251] br[251] wl[151] vdd gnd cell_6t
Xbit_r152_c251 bl[251] br[251] wl[152] vdd gnd cell_6t
Xbit_r153_c251 bl[251] br[251] wl[153] vdd gnd cell_6t
Xbit_r154_c251 bl[251] br[251] wl[154] vdd gnd cell_6t
Xbit_r155_c251 bl[251] br[251] wl[155] vdd gnd cell_6t
Xbit_r156_c251 bl[251] br[251] wl[156] vdd gnd cell_6t
Xbit_r157_c251 bl[251] br[251] wl[157] vdd gnd cell_6t
Xbit_r158_c251 bl[251] br[251] wl[158] vdd gnd cell_6t
Xbit_r159_c251 bl[251] br[251] wl[159] vdd gnd cell_6t
Xbit_r160_c251 bl[251] br[251] wl[160] vdd gnd cell_6t
Xbit_r161_c251 bl[251] br[251] wl[161] vdd gnd cell_6t
Xbit_r162_c251 bl[251] br[251] wl[162] vdd gnd cell_6t
Xbit_r163_c251 bl[251] br[251] wl[163] vdd gnd cell_6t
Xbit_r164_c251 bl[251] br[251] wl[164] vdd gnd cell_6t
Xbit_r165_c251 bl[251] br[251] wl[165] vdd gnd cell_6t
Xbit_r166_c251 bl[251] br[251] wl[166] vdd gnd cell_6t
Xbit_r167_c251 bl[251] br[251] wl[167] vdd gnd cell_6t
Xbit_r168_c251 bl[251] br[251] wl[168] vdd gnd cell_6t
Xbit_r169_c251 bl[251] br[251] wl[169] vdd gnd cell_6t
Xbit_r170_c251 bl[251] br[251] wl[170] vdd gnd cell_6t
Xbit_r171_c251 bl[251] br[251] wl[171] vdd gnd cell_6t
Xbit_r172_c251 bl[251] br[251] wl[172] vdd gnd cell_6t
Xbit_r173_c251 bl[251] br[251] wl[173] vdd gnd cell_6t
Xbit_r174_c251 bl[251] br[251] wl[174] vdd gnd cell_6t
Xbit_r175_c251 bl[251] br[251] wl[175] vdd gnd cell_6t
Xbit_r176_c251 bl[251] br[251] wl[176] vdd gnd cell_6t
Xbit_r177_c251 bl[251] br[251] wl[177] vdd gnd cell_6t
Xbit_r178_c251 bl[251] br[251] wl[178] vdd gnd cell_6t
Xbit_r179_c251 bl[251] br[251] wl[179] vdd gnd cell_6t
Xbit_r180_c251 bl[251] br[251] wl[180] vdd gnd cell_6t
Xbit_r181_c251 bl[251] br[251] wl[181] vdd gnd cell_6t
Xbit_r182_c251 bl[251] br[251] wl[182] vdd gnd cell_6t
Xbit_r183_c251 bl[251] br[251] wl[183] vdd gnd cell_6t
Xbit_r184_c251 bl[251] br[251] wl[184] vdd gnd cell_6t
Xbit_r185_c251 bl[251] br[251] wl[185] vdd gnd cell_6t
Xbit_r186_c251 bl[251] br[251] wl[186] vdd gnd cell_6t
Xbit_r187_c251 bl[251] br[251] wl[187] vdd gnd cell_6t
Xbit_r188_c251 bl[251] br[251] wl[188] vdd gnd cell_6t
Xbit_r189_c251 bl[251] br[251] wl[189] vdd gnd cell_6t
Xbit_r190_c251 bl[251] br[251] wl[190] vdd gnd cell_6t
Xbit_r191_c251 bl[251] br[251] wl[191] vdd gnd cell_6t
Xbit_r192_c251 bl[251] br[251] wl[192] vdd gnd cell_6t
Xbit_r193_c251 bl[251] br[251] wl[193] vdd gnd cell_6t
Xbit_r194_c251 bl[251] br[251] wl[194] vdd gnd cell_6t
Xbit_r195_c251 bl[251] br[251] wl[195] vdd gnd cell_6t
Xbit_r196_c251 bl[251] br[251] wl[196] vdd gnd cell_6t
Xbit_r197_c251 bl[251] br[251] wl[197] vdd gnd cell_6t
Xbit_r198_c251 bl[251] br[251] wl[198] vdd gnd cell_6t
Xbit_r199_c251 bl[251] br[251] wl[199] vdd gnd cell_6t
Xbit_r200_c251 bl[251] br[251] wl[200] vdd gnd cell_6t
Xbit_r201_c251 bl[251] br[251] wl[201] vdd gnd cell_6t
Xbit_r202_c251 bl[251] br[251] wl[202] vdd gnd cell_6t
Xbit_r203_c251 bl[251] br[251] wl[203] vdd gnd cell_6t
Xbit_r204_c251 bl[251] br[251] wl[204] vdd gnd cell_6t
Xbit_r205_c251 bl[251] br[251] wl[205] vdd gnd cell_6t
Xbit_r206_c251 bl[251] br[251] wl[206] vdd gnd cell_6t
Xbit_r207_c251 bl[251] br[251] wl[207] vdd gnd cell_6t
Xbit_r208_c251 bl[251] br[251] wl[208] vdd gnd cell_6t
Xbit_r209_c251 bl[251] br[251] wl[209] vdd gnd cell_6t
Xbit_r210_c251 bl[251] br[251] wl[210] vdd gnd cell_6t
Xbit_r211_c251 bl[251] br[251] wl[211] vdd gnd cell_6t
Xbit_r212_c251 bl[251] br[251] wl[212] vdd gnd cell_6t
Xbit_r213_c251 bl[251] br[251] wl[213] vdd gnd cell_6t
Xbit_r214_c251 bl[251] br[251] wl[214] vdd gnd cell_6t
Xbit_r215_c251 bl[251] br[251] wl[215] vdd gnd cell_6t
Xbit_r216_c251 bl[251] br[251] wl[216] vdd gnd cell_6t
Xbit_r217_c251 bl[251] br[251] wl[217] vdd gnd cell_6t
Xbit_r218_c251 bl[251] br[251] wl[218] vdd gnd cell_6t
Xbit_r219_c251 bl[251] br[251] wl[219] vdd gnd cell_6t
Xbit_r220_c251 bl[251] br[251] wl[220] vdd gnd cell_6t
Xbit_r221_c251 bl[251] br[251] wl[221] vdd gnd cell_6t
Xbit_r222_c251 bl[251] br[251] wl[222] vdd gnd cell_6t
Xbit_r223_c251 bl[251] br[251] wl[223] vdd gnd cell_6t
Xbit_r224_c251 bl[251] br[251] wl[224] vdd gnd cell_6t
Xbit_r225_c251 bl[251] br[251] wl[225] vdd gnd cell_6t
Xbit_r226_c251 bl[251] br[251] wl[226] vdd gnd cell_6t
Xbit_r227_c251 bl[251] br[251] wl[227] vdd gnd cell_6t
Xbit_r228_c251 bl[251] br[251] wl[228] vdd gnd cell_6t
Xbit_r229_c251 bl[251] br[251] wl[229] vdd gnd cell_6t
Xbit_r230_c251 bl[251] br[251] wl[230] vdd gnd cell_6t
Xbit_r231_c251 bl[251] br[251] wl[231] vdd gnd cell_6t
Xbit_r232_c251 bl[251] br[251] wl[232] vdd gnd cell_6t
Xbit_r233_c251 bl[251] br[251] wl[233] vdd gnd cell_6t
Xbit_r234_c251 bl[251] br[251] wl[234] vdd gnd cell_6t
Xbit_r235_c251 bl[251] br[251] wl[235] vdd gnd cell_6t
Xbit_r236_c251 bl[251] br[251] wl[236] vdd gnd cell_6t
Xbit_r237_c251 bl[251] br[251] wl[237] vdd gnd cell_6t
Xbit_r238_c251 bl[251] br[251] wl[238] vdd gnd cell_6t
Xbit_r239_c251 bl[251] br[251] wl[239] vdd gnd cell_6t
Xbit_r240_c251 bl[251] br[251] wl[240] vdd gnd cell_6t
Xbit_r241_c251 bl[251] br[251] wl[241] vdd gnd cell_6t
Xbit_r242_c251 bl[251] br[251] wl[242] vdd gnd cell_6t
Xbit_r243_c251 bl[251] br[251] wl[243] vdd gnd cell_6t
Xbit_r244_c251 bl[251] br[251] wl[244] vdd gnd cell_6t
Xbit_r245_c251 bl[251] br[251] wl[245] vdd gnd cell_6t
Xbit_r246_c251 bl[251] br[251] wl[246] vdd gnd cell_6t
Xbit_r247_c251 bl[251] br[251] wl[247] vdd gnd cell_6t
Xbit_r248_c251 bl[251] br[251] wl[248] vdd gnd cell_6t
Xbit_r249_c251 bl[251] br[251] wl[249] vdd gnd cell_6t
Xbit_r250_c251 bl[251] br[251] wl[250] vdd gnd cell_6t
Xbit_r251_c251 bl[251] br[251] wl[251] vdd gnd cell_6t
Xbit_r252_c251 bl[251] br[251] wl[252] vdd gnd cell_6t
Xbit_r253_c251 bl[251] br[251] wl[253] vdd gnd cell_6t
Xbit_r254_c251 bl[251] br[251] wl[254] vdd gnd cell_6t
Xbit_r255_c251 bl[251] br[251] wl[255] vdd gnd cell_6t
Xbit_r0_c252 bl[252] br[252] wl[0] vdd gnd cell_6t
Xbit_r1_c252 bl[252] br[252] wl[1] vdd gnd cell_6t
Xbit_r2_c252 bl[252] br[252] wl[2] vdd gnd cell_6t
Xbit_r3_c252 bl[252] br[252] wl[3] vdd gnd cell_6t
Xbit_r4_c252 bl[252] br[252] wl[4] vdd gnd cell_6t
Xbit_r5_c252 bl[252] br[252] wl[5] vdd gnd cell_6t
Xbit_r6_c252 bl[252] br[252] wl[6] vdd gnd cell_6t
Xbit_r7_c252 bl[252] br[252] wl[7] vdd gnd cell_6t
Xbit_r8_c252 bl[252] br[252] wl[8] vdd gnd cell_6t
Xbit_r9_c252 bl[252] br[252] wl[9] vdd gnd cell_6t
Xbit_r10_c252 bl[252] br[252] wl[10] vdd gnd cell_6t
Xbit_r11_c252 bl[252] br[252] wl[11] vdd gnd cell_6t
Xbit_r12_c252 bl[252] br[252] wl[12] vdd gnd cell_6t
Xbit_r13_c252 bl[252] br[252] wl[13] vdd gnd cell_6t
Xbit_r14_c252 bl[252] br[252] wl[14] vdd gnd cell_6t
Xbit_r15_c252 bl[252] br[252] wl[15] vdd gnd cell_6t
Xbit_r16_c252 bl[252] br[252] wl[16] vdd gnd cell_6t
Xbit_r17_c252 bl[252] br[252] wl[17] vdd gnd cell_6t
Xbit_r18_c252 bl[252] br[252] wl[18] vdd gnd cell_6t
Xbit_r19_c252 bl[252] br[252] wl[19] vdd gnd cell_6t
Xbit_r20_c252 bl[252] br[252] wl[20] vdd gnd cell_6t
Xbit_r21_c252 bl[252] br[252] wl[21] vdd gnd cell_6t
Xbit_r22_c252 bl[252] br[252] wl[22] vdd gnd cell_6t
Xbit_r23_c252 bl[252] br[252] wl[23] vdd gnd cell_6t
Xbit_r24_c252 bl[252] br[252] wl[24] vdd gnd cell_6t
Xbit_r25_c252 bl[252] br[252] wl[25] vdd gnd cell_6t
Xbit_r26_c252 bl[252] br[252] wl[26] vdd gnd cell_6t
Xbit_r27_c252 bl[252] br[252] wl[27] vdd gnd cell_6t
Xbit_r28_c252 bl[252] br[252] wl[28] vdd gnd cell_6t
Xbit_r29_c252 bl[252] br[252] wl[29] vdd gnd cell_6t
Xbit_r30_c252 bl[252] br[252] wl[30] vdd gnd cell_6t
Xbit_r31_c252 bl[252] br[252] wl[31] vdd gnd cell_6t
Xbit_r32_c252 bl[252] br[252] wl[32] vdd gnd cell_6t
Xbit_r33_c252 bl[252] br[252] wl[33] vdd gnd cell_6t
Xbit_r34_c252 bl[252] br[252] wl[34] vdd gnd cell_6t
Xbit_r35_c252 bl[252] br[252] wl[35] vdd gnd cell_6t
Xbit_r36_c252 bl[252] br[252] wl[36] vdd gnd cell_6t
Xbit_r37_c252 bl[252] br[252] wl[37] vdd gnd cell_6t
Xbit_r38_c252 bl[252] br[252] wl[38] vdd gnd cell_6t
Xbit_r39_c252 bl[252] br[252] wl[39] vdd gnd cell_6t
Xbit_r40_c252 bl[252] br[252] wl[40] vdd gnd cell_6t
Xbit_r41_c252 bl[252] br[252] wl[41] vdd gnd cell_6t
Xbit_r42_c252 bl[252] br[252] wl[42] vdd gnd cell_6t
Xbit_r43_c252 bl[252] br[252] wl[43] vdd gnd cell_6t
Xbit_r44_c252 bl[252] br[252] wl[44] vdd gnd cell_6t
Xbit_r45_c252 bl[252] br[252] wl[45] vdd gnd cell_6t
Xbit_r46_c252 bl[252] br[252] wl[46] vdd gnd cell_6t
Xbit_r47_c252 bl[252] br[252] wl[47] vdd gnd cell_6t
Xbit_r48_c252 bl[252] br[252] wl[48] vdd gnd cell_6t
Xbit_r49_c252 bl[252] br[252] wl[49] vdd gnd cell_6t
Xbit_r50_c252 bl[252] br[252] wl[50] vdd gnd cell_6t
Xbit_r51_c252 bl[252] br[252] wl[51] vdd gnd cell_6t
Xbit_r52_c252 bl[252] br[252] wl[52] vdd gnd cell_6t
Xbit_r53_c252 bl[252] br[252] wl[53] vdd gnd cell_6t
Xbit_r54_c252 bl[252] br[252] wl[54] vdd gnd cell_6t
Xbit_r55_c252 bl[252] br[252] wl[55] vdd gnd cell_6t
Xbit_r56_c252 bl[252] br[252] wl[56] vdd gnd cell_6t
Xbit_r57_c252 bl[252] br[252] wl[57] vdd gnd cell_6t
Xbit_r58_c252 bl[252] br[252] wl[58] vdd gnd cell_6t
Xbit_r59_c252 bl[252] br[252] wl[59] vdd gnd cell_6t
Xbit_r60_c252 bl[252] br[252] wl[60] vdd gnd cell_6t
Xbit_r61_c252 bl[252] br[252] wl[61] vdd gnd cell_6t
Xbit_r62_c252 bl[252] br[252] wl[62] vdd gnd cell_6t
Xbit_r63_c252 bl[252] br[252] wl[63] vdd gnd cell_6t
Xbit_r64_c252 bl[252] br[252] wl[64] vdd gnd cell_6t
Xbit_r65_c252 bl[252] br[252] wl[65] vdd gnd cell_6t
Xbit_r66_c252 bl[252] br[252] wl[66] vdd gnd cell_6t
Xbit_r67_c252 bl[252] br[252] wl[67] vdd gnd cell_6t
Xbit_r68_c252 bl[252] br[252] wl[68] vdd gnd cell_6t
Xbit_r69_c252 bl[252] br[252] wl[69] vdd gnd cell_6t
Xbit_r70_c252 bl[252] br[252] wl[70] vdd gnd cell_6t
Xbit_r71_c252 bl[252] br[252] wl[71] vdd gnd cell_6t
Xbit_r72_c252 bl[252] br[252] wl[72] vdd gnd cell_6t
Xbit_r73_c252 bl[252] br[252] wl[73] vdd gnd cell_6t
Xbit_r74_c252 bl[252] br[252] wl[74] vdd gnd cell_6t
Xbit_r75_c252 bl[252] br[252] wl[75] vdd gnd cell_6t
Xbit_r76_c252 bl[252] br[252] wl[76] vdd gnd cell_6t
Xbit_r77_c252 bl[252] br[252] wl[77] vdd gnd cell_6t
Xbit_r78_c252 bl[252] br[252] wl[78] vdd gnd cell_6t
Xbit_r79_c252 bl[252] br[252] wl[79] vdd gnd cell_6t
Xbit_r80_c252 bl[252] br[252] wl[80] vdd gnd cell_6t
Xbit_r81_c252 bl[252] br[252] wl[81] vdd gnd cell_6t
Xbit_r82_c252 bl[252] br[252] wl[82] vdd gnd cell_6t
Xbit_r83_c252 bl[252] br[252] wl[83] vdd gnd cell_6t
Xbit_r84_c252 bl[252] br[252] wl[84] vdd gnd cell_6t
Xbit_r85_c252 bl[252] br[252] wl[85] vdd gnd cell_6t
Xbit_r86_c252 bl[252] br[252] wl[86] vdd gnd cell_6t
Xbit_r87_c252 bl[252] br[252] wl[87] vdd gnd cell_6t
Xbit_r88_c252 bl[252] br[252] wl[88] vdd gnd cell_6t
Xbit_r89_c252 bl[252] br[252] wl[89] vdd gnd cell_6t
Xbit_r90_c252 bl[252] br[252] wl[90] vdd gnd cell_6t
Xbit_r91_c252 bl[252] br[252] wl[91] vdd gnd cell_6t
Xbit_r92_c252 bl[252] br[252] wl[92] vdd gnd cell_6t
Xbit_r93_c252 bl[252] br[252] wl[93] vdd gnd cell_6t
Xbit_r94_c252 bl[252] br[252] wl[94] vdd gnd cell_6t
Xbit_r95_c252 bl[252] br[252] wl[95] vdd gnd cell_6t
Xbit_r96_c252 bl[252] br[252] wl[96] vdd gnd cell_6t
Xbit_r97_c252 bl[252] br[252] wl[97] vdd gnd cell_6t
Xbit_r98_c252 bl[252] br[252] wl[98] vdd gnd cell_6t
Xbit_r99_c252 bl[252] br[252] wl[99] vdd gnd cell_6t
Xbit_r100_c252 bl[252] br[252] wl[100] vdd gnd cell_6t
Xbit_r101_c252 bl[252] br[252] wl[101] vdd gnd cell_6t
Xbit_r102_c252 bl[252] br[252] wl[102] vdd gnd cell_6t
Xbit_r103_c252 bl[252] br[252] wl[103] vdd gnd cell_6t
Xbit_r104_c252 bl[252] br[252] wl[104] vdd gnd cell_6t
Xbit_r105_c252 bl[252] br[252] wl[105] vdd gnd cell_6t
Xbit_r106_c252 bl[252] br[252] wl[106] vdd gnd cell_6t
Xbit_r107_c252 bl[252] br[252] wl[107] vdd gnd cell_6t
Xbit_r108_c252 bl[252] br[252] wl[108] vdd gnd cell_6t
Xbit_r109_c252 bl[252] br[252] wl[109] vdd gnd cell_6t
Xbit_r110_c252 bl[252] br[252] wl[110] vdd gnd cell_6t
Xbit_r111_c252 bl[252] br[252] wl[111] vdd gnd cell_6t
Xbit_r112_c252 bl[252] br[252] wl[112] vdd gnd cell_6t
Xbit_r113_c252 bl[252] br[252] wl[113] vdd gnd cell_6t
Xbit_r114_c252 bl[252] br[252] wl[114] vdd gnd cell_6t
Xbit_r115_c252 bl[252] br[252] wl[115] vdd gnd cell_6t
Xbit_r116_c252 bl[252] br[252] wl[116] vdd gnd cell_6t
Xbit_r117_c252 bl[252] br[252] wl[117] vdd gnd cell_6t
Xbit_r118_c252 bl[252] br[252] wl[118] vdd gnd cell_6t
Xbit_r119_c252 bl[252] br[252] wl[119] vdd gnd cell_6t
Xbit_r120_c252 bl[252] br[252] wl[120] vdd gnd cell_6t
Xbit_r121_c252 bl[252] br[252] wl[121] vdd gnd cell_6t
Xbit_r122_c252 bl[252] br[252] wl[122] vdd gnd cell_6t
Xbit_r123_c252 bl[252] br[252] wl[123] vdd gnd cell_6t
Xbit_r124_c252 bl[252] br[252] wl[124] vdd gnd cell_6t
Xbit_r125_c252 bl[252] br[252] wl[125] vdd gnd cell_6t
Xbit_r126_c252 bl[252] br[252] wl[126] vdd gnd cell_6t
Xbit_r127_c252 bl[252] br[252] wl[127] vdd gnd cell_6t
Xbit_r128_c252 bl[252] br[252] wl[128] vdd gnd cell_6t
Xbit_r129_c252 bl[252] br[252] wl[129] vdd gnd cell_6t
Xbit_r130_c252 bl[252] br[252] wl[130] vdd gnd cell_6t
Xbit_r131_c252 bl[252] br[252] wl[131] vdd gnd cell_6t
Xbit_r132_c252 bl[252] br[252] wl[132] vdd gnd cell_6t
Xbit_r133_c252 bl[252] br[252] wl[133] vdd gnd cell_6t
Xbit_r134_c252 bl[252] br[252] wl[134] vdd gnd cell_6t
Xbit_r135_c252 bl[252] br[252] wl[135] vdd gnd cell_6t
Xbit_r136_c252 bl[252] br[252] wl[136] vdd gnd cell_6t
Xbit_r137_c252 bl[252] br[252] wl[137] vdd gnd cell_6t
Xbit_r138_c252 bl[252] br[252] wl[138] vdd gnd cell_6t
Xbit_r139_c252 bl[252] br[252] wl[139] vdd gnd cell_6t
Xbit_r140_c252 bl[252] br[252] wl[140] vdd gnd cell_6t
Xbit_r141_c252 bl[252] br[252] wl[141] vdd gnd cell_6t
Xbit_r142_c252 bl[252] br[252] wl[142] vdd gnd cell_6t
Xbit_r143_c252 bl[252] br[252] wl[143] vdd gnd cell_6t
Xbit_r144_c252 bl[252] br[252] wl[144] vdd gnd cell_6t
Xbit_r145_c252 bl[252] br[252] wl[145] vdd gnd cell_6t
Xbit_r146_c252 bl[252] br[252] wl[146] vdd gnd cell_6t
Xbit_r147_c252 bl[252] br[252] wl[147] vdd gnd cell_6t
Xbit_r148_c252 bl[252] br[252] wl[148] vdd gnd cell_6t
Xbit_r149_c252 bl[252] br[252] wl[149] vdd gnd cell_6t
Xbit_r150_c252 bl[252] br[252] wl[150] vdd gnd cell_6t
Xbit_r151_c252 bl[252] br[252] wl[151] vdd gnd cell_6t
Xbit_r152_c252 bl[252] br[252] wl[152] vdd gnd cell_6t
Xbit_r153_c252 bl[252] br[252] wl[153] vdd gnd cell_6t
Xbit_r154_c252 bl[252] br[252] wl[154] vdd gnd cell_6t
Xbit_r155_c252 bl[252] br[252] wl[155] vdd gnd cell_6t
Xbit_r156_c252 bl[252] br[252] wl[156] vdd gnd cell_6t
Xbit_r157_c252 bl[252] br[252] wl[157] vdd gnd cell_6t
Xbit_r158_c252 bl[252] br[252] wl[158] vdd gnd cell_6t
Xbit_r159_c252 bl[252] br[252] wl[159] vdd gnd cell_6t
Xbit_r160_c252 bl[252] br[252] wl[160] vdd gnd cell_6t
Xbit_r161_c252 bl[252] br[252] wl[161] vdd gnd cell_6t
Xbit_r162_c252 bl[252] br[252] wl[162] vdd gnd cell_6t
Xbit_r163_c252 bl[252] br[252] wl[163] vdd gnd cell_6t
Xbit_r164_c252 bl[252] br[252] wl[164] vdd gnd cell_6t
Xbit_r165_c252 bl[252] br[252] wl[165] vdd gnd cell_6t
Xbit_r166_c252 bl[252] br[252] wl[166] vdd gnd cell_6t
Xbit_r167_c252 bl[252] br[252] wl[167] vdd gnd cell_6t
Xbit_r168_c252 bl[252] br[252] wl[168] vdd gnd cell_6t
Xbit_r169_c252 bl[252] br[252] wl[169] vdd gnd cell_6t
Xbit_r170_c252 bl[252] br[252] wl[170] vdd gnd cell_6t
Xbit_r171_c252 bl[252] br[252] wl[171] vdd gnd cell_6t
Xbit_r172_c252 bl[252] br[252] wl[172] vdd gnd cell_6t
Xbit_r173_c252 bl[252] br[252] wl[173] vdd gnd cell_6t
Xbit_r174_c252 bl[252] br[252] wl[174] vdd gnd cell_6t
Xbit_r175_c252 bl[252] br[252] wl[175] vdd gnd cell_6t
Xbit_r176_c252 bl[252] br[252] wl[176] vdd gnd cell_6t
Xbit_r177_c252 bl[252] br[252] wl[177] vdd gnd cell_6t
Xbit_r178_c252 bl[252] br[252] wl[178] vdd gnd cell_6t
Xbit_r179_c252 bl[252] br[252] wl[179] vdd gnd cell_6t
Xbit_r180_c252 bl[252] br[252] wl[180] vdd gnd cell_6t
Xbit_r181_c252 bl[252] br[252] wl[181] vdd gnd cell_6t
Xbit_r182_c252 bl[252] br[252] wl[182] vdd gnd cell_6t
Xbit_r183_c252 bl[252] br[252] wl[183] vdd gnd cell_6t
Xbit_r184_c252 bl[252] br[252] wl[184] vdd gnd cell_6t
Xbit_r185_c252 bl[252] br[252] wl[185] vdd gnd cell_6t
Xbit_r186_c252 bl[252] br[252] wl[186] vdd gnd cell_6t
Xbit_r187_c252 bl[252] br[252] wl[187] vdd gnd cell_6t
Xbit_r188_c252 bl[252] br[252] wl[188] vdd gnd cell_6t
Xbit_r189_c252 bl[252] br[252] wl[189] vdd gnd cell_6t
Xbit_r190_c252 bl[252] br[252] wl[190] vdd gnd cell_6t
Xbit_r191_c252 bl[252] br[252] wl[191] vdd gnd cell_6t
Xbit_r192_c252 bl[252] br[252] wl[192] vdd gnd cell_6t
Xbit_r193_c252 bl[252] br[252] wl[193] vdd gnd cell_6t
Xbit_r194_c252 bl[252] br[252] wl[194] vdd gnd cell_6t
Xbit_r195_c252 bl[252] br[252] wl[195] vdd gnd cell_6t
Xbit_r196_c252 bl[252] br[252] wl[196] vdd gnd cell_6t
Xbit_r197_c252 bl[252] br[252] wl[197] vdd gnd cell_6t
Xbit_r198_c252 bl[252] br[252] wl[198] vdd gnd cell_6t
Xbit_r199_c252 bl[252] br[252] wl[199] vdd gnd cell_6t
Xbit_r200_c252 bl[252] br[252] wl[200] vdd gnd cell_6t
Xbit_r201_c252 bl[252] br[252] wl[201] vdd gnd cell_6t
Xbit_r202_c252 bl[252] br[252] wl[202] vdd gnd cell_6t
Xbit_r203_c252 bl[252] br[252] wl[203] vdd gnd cell_6t
Xbit_r204_c252 bl[252] br[252] wl[204] vdd gnd cell_6t
Xbit_r205_c252 bl[252] br[252] wl[205] vdd gnd cell_6t
Xbit_r206_c252 bl[252] br[252] wl[206] vdd gnd cell_6t
Xbit_r207_c252 bl[252] br[252] wl[207] vdd gnd cell_6t
Xbit_r208_c252 bl[252] br[252] wl[208] vdd gnd cell_6t
Xbit_r209_c252 bl[252] br[252] wl[209] vdd gnd cell_6t
Xbit_r210_c252 bl[252] br[252] wl[210] vdd gnd cell_6t
Xbit_r211_c252 bl[252] br[252] wl[211] vdd gnd cell_6t
Xbit_r212_c252 bl[252] br[252] wl[212] vdd gnd cell_6t
Xbit_r213_c252 bl[252] br[252] wl[213] vdd gnd cell_6t
Xbit_r214_c252 bl[252] br[252] wl[214] vdd gnd cell_6t
Xbit_r215_c252 bl[252] br[252] wl[215] vdd gnd cell_6t
Xbit_r216_c252 bl[252] br[252] wl[216] vdd gnd cell_6t
Xbit_r217_c252 bl[252] br[252] wl[217] vdd gnd cell_6t
Xbit_r218_c252 bl[252] br[252] wl[218] vdd gnd cell_6t
Xbit_r219_c252 bl[252] br[252] wl[219] vdd gnd cell_6t
Xbit_r220_c252 bl[252] br[252] wl[220] vdd gnd cell_6t
Xbit_r221_c252 bl[252] br[252] wl[221] vdd gnd cell_6t
Xbit_r222_c252 bl[252] br[252] wl[222] vdd gnd cell_6t
Xbit_r223_c252 bl[252] br[252] wl[223] vdd gnd cell_6t
Xbit_r224_c252 bl[252] br[252] wl[224] vdd gnd cell_6t
Xbit_r225_c252 bl[252] br[252] wl[225] vdd gnd cell_6t
Xbit_r226_c252 bl[252] br[252] wl[226] vdd gnd cell_6t
Xbit_r227_c252 bl[252] br[252] wl[227] vdd gnd cell_6t
Xbit_r228_c252 bl[252] br[252] wl[228] vdd gnd cell_6t
Xbit_r229_c252 bl[252] br[252] wl[229] vdd gnd cell_6t
Xbit_r230_c252 bl[252] br[252] wl[230] vdd gnd cell_6t
Xbit_r231_c252 bl[252] br[252] wl[231] vdd gnd cell_6t
Xbit_r232_c252 bl[252] br[252] wl[232] vdd gnd cell_6t
Xbit_r233_c252 bl[252] br[252] wl[233] vdd gnd cell_6t
Xbit_r234_c252 bl[252] br[252] wl[234] vdd gnd cell_6t
Xbit_r235_c252 bl[252] br[252] wl[235] vdd gnd cell_6t
Xbit_r236_c252 bl[252] br[252] wl[236] vdd gnd cell_6t
Xbit_r237_c252 bl[252] br[252] wl[237] vdd gnd cell_6t
Xbit_r238_c252 bl[252] br[252] wl[238] vdd gnd cell_6t
Xbit_r239_c252 bl[252] br[252] wl[239] vdd gnd cell_6t
Xbit_r240_c252 bl[252] br[252] wl[240] vdd gnd cell_6t
Xbit_r241_c252 bl[252] br[252] wl[241] vdd gnd cell_6t
Xbit_r242_c252 bl[252] br[252] wl[242] vdd gnd cell_6t
Xbit_r243_c252 bl[252] br[252] wl[243] vdd gnd cell_6t
Xbit_r244_c252 bl[252] br[252] wl[244] vdd gnd cell_6t
Xbit_r245_c252 bl[252] br[252] wl[245] vdd gnd cell_6t
Xbit_r246_c252 bl[252] br[252] wl[246] vdd gnd cell_6t
Xbit_r247_c252 bl[252] br[252] wl[247] vdd gnd cell_6t
Xbit_r248_c252 bl[252] br[252] wl[248] vdd gnd cell_6t
Xbit_r249_c252 bl[252] br[252] wl[249] vdd gnd cell_6t
Xbit_r250_c252 bl[252] br[252] wl[250] vdd gnd cell_6t
Xbit_r251_c252 bl[252] br[252] wl[251] vdd gnd cell_6t
Xbit_r252_c252 bl[252] br[252] wl[252] vdd gnd cell_6t
Xbit_r253_c252 bl[252] br[252] wl[253] vdd gnd cell_6t
Xbit_r254_c252 bl[252] br[252] wl[254] vdd gnd cell_6t
Xbit_r255_c252 bl[252] br[252] wl[255] vdd gnd cell_6t
Xbit_r0_c253 bl[253] br[253] wl[0] vdd gnd cell_6t
Xbit_r1_c253 bl[253] br[253] wl[1] vdd gnd cell_6t
Xbit_r2_c253 bl[253] br[253] wl[2] vdd gnd cell_6t
Xbit_r3_c253 bl[253] br[253] wl[3] vdd gnd cell_6t
Xbit_r4_c253 bl[253] br[253] wl[4] vdd gnd cell_6t
Xbit_r5_c253 bl[253] br[253] wl[5] vdd gnd cell_6t
Xbit_r6_c253 bl[253] br[253] wl[6] vdd gnd cell_6t
Xbit_r7_c253 bl[253] br[253] wl[7] vdd gnd cell_6t
Xbit_r8_c253 bl[253] br[253] wl[8] vdd gnd cell_6t
Xbit_r9_c253 bl[253] br[253] wl[9] vdd gnd cell_6t
Xbit_r10_c253 bl[253] br[253] wl[10] vdd gnd cell_6t
Xbit_r11_c253 bl[253] br[253] wl[11] vdd gnd cell_6t
Xbit_r12_c253 bl[253] br[253] wl[12] vdd gnd cell_6t
Xbit_r13_c253 bl[253] br[253] wl[13] vdd gnd cell_6t
Xbit_r14_c253 bl[253] br[253] wl[14] vdd gnd cell_6t
Xbit_r15_c253 bl[253] br[253] wl[15] vdd gnd cell_6t
Xbit_r16_c253 bl[253] br[253] wl[16] vdd gnd cell_6t
Xbit_r17_c253 bl[253] br[253] wl[17] vdd gnd cell_6t
Xbit_r18_c253 bl[253] br[253] wl[18] vdd gnd cell_6t
Xbit_r19_c253 bl[253] br[253] wl[19] vdd gnd cell_6t
Xbit_r20_c253 bl[253] br[253] wl[20] vdd gnd cell_6t
Xbit_r21_c253 bl[253] br[253] wl[21] vdd gnd cell_6t
Xbit_r22_c253 bl[253] br[253] wl[22] vdd gnd cell_6t
Xbit_r23_c253 bl[253] br[253] wl[23] vdd gnd cell_6t
Xbit_r24_c253 bl[253] br[253] wl[24] vdd gnd cell_6t
Xbit_r25_c253 bl[253] br[253] wl[25] vdd gnd cell_6t
Xbit_r26_c253 bl[253] br[253] wl[26] vdd gnd cell_6t
Xbit_r27_c253 bl[253] br[253] wl[27] vdd gnd cell_6t
Xbit_r28_c253 bl[253] br[253] wl[28] vdd gnd cell_6t
Xbit_r29_c253 bl[253] br[253] wl[29] vdd gnd cell_6t
Xbit_r30_c253 bl[253] br[253] wl[30] vdd gnd cell_6t
Xbit_r31_c253 bl[253] br[253] wl[31] vdd gnd cell_6t
Xbit_r32_c253 bl[253] br[253] wl[32] vdd gnd cell_6t
Xbit_r33_c253 bl[253] br[253] wl[33] vdd gnd cell_6t
Xbit_r34_c253 bl[253] br[253] wl[34] vdd gnd cell_6t
Xbit_r35_c253 bl[253] br[253] wl[35] vdd gnd cell_6t
Xbit_r36_c253 bl[253] br[253] wl[36] vdd gnd cell_6t
Xbit_r37_c253 bl[253] br[253] wl[37] vdd gnd cell_6t
Xbit_r38_c253 bl[253] br[253] wl[38] vdd gnd cell_6t
Xbit_r39_c253 bl[253] br[253] wl[39] vdd gnd cell_6t
Xbit_r40_c253 bl[253] br[253] wl[40] vdd gnd cell_6t
Xbit_r41_c253 bl[253] br[253] wl[41] vdd gnd cell_6t
Xbit_r42_c253 bl[253] br[253] wl[42] vdd gnd cell_6t
Xbit_r43_c253 bl[253] br[253] wl[43] vdd gnd cell_6t
Xbit_r44_c253 bl[253] br[253] wl[44] vdd gnd cell_6t
Xbit_r45_c253 bl[253] br[253] wl[45] vdd gnd cell_6t
Xbit_r46_c253 bl[253] br[253] wl[46] vdd gnd cell_6t
Xbit_r47_c253 bl[253] br[253] wl[47] vdd gnd cell_6t
Xbit_r48_c253 bl[253] br[253] wl[48] vdd gnd cell_6t
Xbit_r49_c253 bl[253] br[253] wl[49] vdd gnd cell_6t
Xbit_r50_c253 bl[253] br[253] wl[50] vdd gnd cell_6t
Xbit_r51_c253 bl[253] br[253] wl[51] vdd gnd cell_6t
Xbit_r52_c253 bl[253] br[253] wl[52] vdd gnd cell_6t
Xbit_r53_c253 bl[253] br[253] wl[53] vdd gnd cell_6t
Xbit_r54_c253 bl[253] br[253] wl[54] vdd gnd cell_6t
Xbit_r55_c253 bl[253] br[253] wl[55] vdd gnd cell_6t
Xbit_r56_c253 bl[253] br[253] wl[56] vdd gnd cell_6t
Xbit_r57_c253 bl[253] br[253] wl[57] vdd gnd cell_6t
Xbit_r58_c253 bl[253] br[253] wl[58] vdd gnd cell_6t
Xbit_r59_c253 bl[253] br[253] wl[59] vdd gnd cell_6t
Xbit_r60_c253 bl[253] br[253] wl[60] vdd gnd cell_6t
Xbit_r61_c253 bl[253] br[253] wl[61] vdd gnd cell_6t
Xbit_r62_c253 bl[253] br[253] wl[62] vdd gnd cell_6t
Xbit_r63_c253 bl[253] br[253] wl[63] vdd gnd cell_6t
Xbit_r64_c253 bl[253] br[253] wl[64] vdd gnd cell_6t
Xbit_r65_c253 bl[253] br[253] wl[65] vdd gnd cell_6t
Xbit_r66_c253 bl[253] br[253] wl[66] vdd gnd cell_6t
Xbit_r67_c253 bl[253] br[253] wl[67] vdd gnd cell_6t
Xbit_r68_c253 bl[253] br[253] wl[68] vdd gnd cell_6t
Xbit_r69_c253 bl[253] br[253] wl[69] vdd gnd cell_6t
Xbit_r70_c253 bl[253] br[253] wl[70] vdd gnd cell_6t
Xbit_r71_c253 bl[253] br[253] wl[71] vdd gnd cell_6t
Xbit_r72_c253 bl[253] br[253] wl[72] vdd gnd cell_6t
Xbit_r73_c253 bl[253] br[253] wl[73] vdd gnd cell_6t
Xbit_r74_c253 bl[253] br[253] wl[74] vdd gnd cell_6t
Xbit_r75_c253 bl[253] br[253] wl[75] vdd gnd cell_6t
Xbit_r76_c253 bl[253] br[253] wl[76] vdd gnd cell_6t
Xbit_r77_c253 bl[253] br[253] wl[77] vdd gnd cell_6t
Xbit_r78_c253 bl[253] br[253] wl[78] vdd gnd cell_6t
Xbit_r79_c253 bl[253] br[253] wl[79] vdd gnd cell_6t
Xbit_r80_c253 bl[253] br[253] wl[80] vdd gnd cell_6t
Xbit_r81_c253 bl[253] br[253] wl[81] vdd gnd cell_6t
Xbit_r82_c253 bl[253] br[253] wl[82] vdd gnd cell_6t
Xbit_r83_c253 bl[253] br[253] wl[83] vdd gnd cell_6t
Xbit_r84_c253 bl[253] br[253] wl[84] vdd gnd cell_6t
Xbit_r85_c253 bl[253] br[253] wl[85] vdd gnd cell_6t
Xbit_r86_c253 bl[253] br[253] wl[86] vdd gnd cell_6t
Xbit_r87_c253 bl[253] br[253] wl[87] vdd gnd cell_6t
Xbit_r88_c253 bl[253] br[253] wl[88] vdd gnd cell_6t
Xbit_r89_c253 bl[253] br[253] wl[89] vdd gnd cell_6t
Xbit_r90_c253 bl[253] br[253] wl[90] vdd gnd cell_6t
Xbit_r91_c253 bl[253] br[253] wl[91] vdd gnd cell_6t
Xbit_r92_c253 bl[253] br[253] wl[92] vdd gnd cell_6t
Xbit_r93_c253 bl[253] br[253] wl[93] vdd gnd cell_6t
Xbit_r94_c253 bl[253] br[253] wl[94] vdd gnd cell_6t
Xbit_r95_c253 bl[253] br[253] wl[95] vdd gnd cell_6t
Xbit_r96_c253 bl[253] br[253] wl[96] vdd gnd cell_6t
Xbit_r97_c253 bl[253] br[253] wl[97] vdd gnd cell_6t
Xbit_r98_c253 bl[253] br[253] wl[98] vdd gnd cell_6t
Xbit_r99_c253 bl[253] br[253] wl[99] vdd gnd cell_6t
Xbit_r100_c253 bl[253] br[253] wl[100] vdd gnd cell_6t
Xbit_r101_c253 bl[253] br[253] wl[101] vdd gnd cell_6t
Xbit_r102_c253 bl[253] br[253] wl[102] vdd gnd cell_6t
Xbit_r103_c253 bl[253] br[253] wl[103] vdd gnd cell_6t
Xbit_r104_c253 bl[253] br[253] wl[104] vdd gnd cell_6t
Xbit_r105_c253 bl[253] br[253] wl[105] vdd gnd cell_6t
Xbit_r106_c253 bl[253] br[253] wl[106] vdd gnd cell_6t
Xbit_r107_c253 bl[253] br[253] wl[107] vdd gnd cell_6t
Xbit_r108_c253 bl[253] br[253] wl[108] vdd gnd cell_6t
Xbit_r109_c253 bl[253] br[253] wl[109] vdd gnd cell_6t
Xbit_r110_c253 bl[253] br[253] wl[110] vdd gnd cell_6t
Xbit_r111_c253 bl[253] br[253] wl[111] vdd gnd cell_6t
Xbit_r112_c253 bl[253] br[253] wl[112] vdd gnd cell_6t
Xbit_r113_c253 bl[253] br[253] wl[113] vdd gnd cell_6t
Xbit_r114_c253 bl[253] br[253] wl[114] vdd gnd cell_6t
Xbit_r115_c253 bl[253] br[253] wl[115] vdd gnd cell_6t
Xbit_r116_c253 bl[253] br[253] wl[116] vdd gnd cell_6t
Xbit_r117_c253 bl[253] br[253] wl[117] vdd gnd cell_6t
Xbit_r118_c253 bl[253] br[253] wl[118] vdd gnd cell_6t
Xbit_r119_c253 bl[253] br[253] wl[119] vdd gnd cell_6t
Xbit_r120_c253 bl[253] br[253] wl[120] vdd gnd cell_6t
Xbit_r121_c253 bl[253] br[253] wl[121] vdd gnd cell_6t
Xbit_r122_c253 bl[253] br[253] wl[122] vdd gnd cell_6t
Xbit_r123_c253 bl[253] br[253] wl[123] vdd gnd cell_6t
Xbit_r124_c253 bl[253] br[253] wl[124] vdd gnd cell_6t
Xbit_r125_c253 bl[253] br[253] wl[125] vdd gnd cell_6t
Xbit_r126_c253 bl[253] br[253] wl[126] vdd gnd cell_6t
Xbit_r127_c253 bl[253] br[253] wl[127] vdd gnd cell_6t
Xbit_r128_c253 bl[253] br[253] wl[128] vdd gnd cell_6t
Xbit_r129_c253 bl[253] br[253] wl[129] vdd gnd cell_6t
Xbit_r130_c253 bl[253] br[253] wl[130] vdd gnd cell_6t
Xbit_r131_c253 bl[253] br[253] wl[131] vdd gnd cell_6t
Xbit_r132_c253 bl[253] br[253] wl[132] vdd gnd cell_6t
Xbit_r133_c253 bl[253] br[253] wl[133] vdd gnd cell_6t
Xbit_r134_c253 bl[253] br[253] wl[134] vdd gnd cell_6t
Xbit_r135_c253 bl[253] br[253] wl[135] vdd gnd cell_6t
Xbit_r136_c253 bl[253] br[253] wl[136] vdd gnd cell_6t
Xbit_r137_c253 bl[253] br[253] wl[137] vdd gnd cell_6t
Xbit_r138_c253 bl[253] br[253] wl[138] vdd gnd cell_6t
Xbit_r139_c253 bl[253] br[253] wl[139] vdd gnd cell_6t
Xbit_r140_c253 bl[253] br[253] wl[140] vdd gnd cell_6t
Xbit_r141_c253 bl[253] br[253] wl[141] vdd gnd cell_6t
Xbit_r142_c253 bl[253] br[253] wl[142] vdd gnd cell_6t
Xbit_r143_c253 bl[253] br[253] wl[143] vdd gnd cell_6t
Xbit_r144_c253 bl[253] br[253] wl[144] vdd gnd cell_6t
Xbit_r145_c253 bl[253] br[253] wl[145] vdd gnd cell_6t
Xbit_r146_c253 bl[253] br[253] wl[146] vdd gnd cell_6t
Xbit_r147_c253 bl[253] br[253] wl[147] vdd gnd cell_6t
Xbit_r148_c253 bl[253] br[253] wl[148] vdd gnd cell_6t
Xbit_r149_c253 bl[253] br[253] wl[149] vdd gnd cell_6t
Xbit_r150_c253 bl[253] br[253] wl[150] vdd gnd cell_6t
Xbit_r151_c253 bl[253] br[253] wl[151] vdd gnd cell_6t
Xbit_r152_c253 bl[253] br[253] wl[152] vdd gnd cell_6t
Xbit_r153_c253 bl[253] br[253] wl[153] vdd gnd cell_6t
Xbit_r154_c253 bl[253] br[253] wl[154] vdd gnd cell_6t
Xbit_r155_c253 bl[253] br[253] wl[155] vdd gnd cell_6t
Xbit_r156_c253 bl[253] br[253] wl[156] vdd gnd cell_6t
Xbit_r157_c253 bl[253] br[253] wl[157] vdd gnd cell_6t
Xbit_r158_c253 bl[253] br[253] wl[158] vdd gnd cell_6t
Xbit_r159_c253 bl[253] br[253] wl[159] vdd gnd cell_6t
Xbit_r160_c253 bl[253] br[253] wl[160] vdd gnd cell_6t
Xbit_r161_c253 bl[253] br[253] wl[161] vdd gnd cell_6t
Xbit_r162_c253 bl[253] br[253] wl[162] vdd gnd cell_6t
Xbit_r163_c253 bl[253] br[253] wl[163] vdd gnd cell_6t
Xbit_r164_c253 bl[253] br[253] wl[164] vdd gnd cell_6t
Xbit_r165_c253 bl[253] br[253] wl[165] vdd gnd cell_6t
Xbit_r166_c253 bl[253] br[253] wl[166] vdd gnd cell_6t
Xbit_r167_c253 bl[253] br[253] wl[167] vdd gnd cell_6t
Xbit_r168_c253 bl[253] br[253] wl[168] vdd gnd cell_6t
Xbit_r169_c253 bl[253] br[253] wl[169] vdd gnd cell_6t
Xbit_r170_c253 bl[253] br[253] wl[170] vdd gnd cell_6t
Xbit_r171_c253 bl[253] br[253] wl[171] vdd gnd cell_6t
Xbit_r172_c253 bl[253] br[253] wl[172] vdd gnd cell_6t
Xbit_r173_c253 bl[253] br[253] wl[173] vdd gnd cell_6t
Xbit_r174_c253 bl[253] br[253] wl[174] vdd gnd cell_6t
Xbit_r175_c253 bl[253] br[253] wl[175] vdd gnd cell_6t
Xbit_r176_c253 bl[253] br[253] wl[176] vdd gnd cell_6t
Xbit_r177_c253 bl[253] br[253] wl[177] vdd gnd cell_6t
Xbit_r178_c253 bl[253] br[253] wl[178] vdd gnd cell_6t
Xbit_r179_c253 bl[253] br[253] wl[179] vdd gnd cell_6t
Xbit_r180_c253 bl[253] br[253] wl[180] vdd gnd cell_6t
Xbit_r181_c253 bl[253] br[253] wl[181] vdd gnd cell_6t
Xbit_r182_c253 bl[253] br[253] wl[182] vdd gnd cell_6t
Xbit_r183_c253 bl[253] br[253] wl[183] vdd gnd cell_6t
Xbit_r184_c253 bl[253] br[253] wl[184] vdd gnd cell_6t
Xbit_r185_c253 bl[253] br[253] wl[185] vdd gnd cell_6t
Xbit_r186_c253 bl[253] br[253] wl[186] vdd gnd cell_6t
Xbit_r187_c253 bl[253] br[253] wl[187] vdd gnd cell_6t
Xbit_r188_c253 bl[253] br[253] wl[188] vdd gnd cell_6t
Xbit_r189_c253 bl[253] br[253] wl[189] vdd gnd cell_6t
Xbit_r190_c253 bl[253] br[253] wl[190] vdd gnd cell_6t
Xbit_r191_c253 bl[253] br[253] wl[191] vdd gnd cell_6t
Xbit_r192_c253 bl[253] br[253] wl[192] vdd gnd cell_6t
Xbit_r193_c253 bl[253] br[253] wl[193] vdd gnd cell_6t
Xbit_r194_c253 bl[253] br[253] wl[194] vdd gnd cell_6t
Xbit_r195_c253 bl[253] br[253] wl[195] vdd gnd cell_6t
Xbit_r196_c253 bl[253] br[253] wl[196] vdd gnd cell_6t
Xbit_r197_c253 bl[253] br[253] wl[197] vdd gnd cell_6t
Xbit_r198_c253 bl[253] br[253] wl[198] vdd gnd cell_6t
Xbit_r199_c253 bl[253] br[253] wl[199] vdd gnd cell_6t
Xbit_r200_c253 bl[253] br[253] wl[200] vdd gnd cell_6t
Xbit_r201_c253 bl[253] br[253] wl[201] vdd gnd cell_6t
Xbit_r202_c253 bl[253] br[253] wl[202] vdd gnd cell_6t
Xbit_r203_c253 bl[253] br[253] wl[203] vdd gnd cell_6t
Xbit_r204_c253 bl[253] br[253] wl[204] vdd gnd cell_6t
Xbit_r205_c253 bl[253] br[253] wl[205] vdd gnd cell_6t
Xbit_r206_c253 bl[253] br[253] wl[206] vdd gnd cell_6t
Xbit_r207_c253 bl[253] br[253] wl[207] vdd gnd cell_6t
Xbit_r208_c253 bl[253] br[253] wl[208] vdd gnd cell_6t
Xbit_r209_c253 bl[253] br[253] wl[209] vdd gnd cell_6t
Xbit_r210_c253 bl[253] br[253] wl[210] vdd gnd cell_6t
Xbit_r211_c253 bl[253] br[253] wl[211] vdd gnd cell_6t
Xbit_r212_c253 bl[253] br[253] wl[212] vdd gnd cell_6t
Xbit_r213_c253 bl[253] br[253] wl[213] vdd gnd cell_6t
Xbit_r214_c253 bl[253] br[253] wl[214] vdd gnd cell_6t
Xbit_r215_c253 bl[253] br[253] wl[215] vdd gnd cell_6t
Xbit_r216_c253 bl[253] br[253] wl[216] vdd gnd cell_6t
Xbit_r217_c253 bl[253] br[253] wl[217] vdd gnd cell_6t
Xbit_r218_c253 bl[253] br[253] wl[218] vdd gnd cell_6t
Xbit_r219_c253 bl[253] br[253] wl[219] vdd gnd cell_6t
Xbit_r220_c253 bl[253] br[253] wl[220] vdd gnd cell_6t
Xbit_r221_c253 bl[253] br[253] wl[221] vdd gnd cell_6t
Xbit_r222_c253 bl[253] br[253] wl[222] vdd gnd cell_6t
Xbit_r223_c253 bl[253] br[253] wl[223] vdd gnd cell_6t
Xbit_r224_c253 bl[253] br[253] wl[224] vdd gnd cell_6t
Xbit_r225_c253 bl[253] br[253] wl[225] vdd gnd cell_6t
Xbit_r226_c253 bl[253] br[253] wl[226] vdd gnd cell_6t
Xbit_r227_c253 bl[253] br[253] wl[227] vdd gnd cell_6t
Xbit_r228_c253 bl[253] br[253] wl[228] vdd gnd cell_6t
Xbit_r229_c253 bl[253] br[253] wl[229] vdd gnd cell_6t
Xbit_r230_c253 bl[253] br[253] wl[230] vdd gnd cell_6t
Xbit_r231_c253 bl[253] br[253] wl[231] vdd gnd cell_6t
Xbit_r232_c253 bl[253] br[253] wl[232] vdd gnd cell_6t
Xbit_r233_c253 bl[253] br[253] wl[233] vdd gnd cell_6t
Xbit_r234_c253 bl[253] br[253] wl[234] vdd gnd cell_6t
Xbit_r235_c253 bl[253] br[253] wl[235] vdd gnd cell_6t
Xbit_r236_c253 bl[253] br[253] wl[236] vdd gnd cell_6t
Xbit_r237_c253 bl[253] br[253] wl[237] vdd gnd cell_6t
Xbit_r238_c253 bl[253] br[253] wl[238] vdd gnd cell_6t
Xbit_r239_c253 bl[253] br[253] wl[239] vdd gnd cell_6t
Xbit_r240_c253 bl[253] br[253] wl[240] vdd gnd cell_6t
Xbit_r241_c253 bl[253] br[253] wl[241] vdd gnd cell_6t
Xbit_r242_c253 bl[253] br[253] wl[242] vdd gnd cell_6t
Xbit_r243_c253 bl[253] br[253] wl[243] vdd gnd cell_6t
Xbit_r244_c253 bl[253] br[253] wl[244] vdd gnd cell_6t
Xbit_r245_c253 bl[253] br[253] wl[245] vdd gnd cell_6t
Xbit_r246_c253 bl[253] br[253] wl[246] vdd gnd cell_6t
Xbit_r247_c253 bl[253] br[253] wl[247] vdd gnd cell_6t
Xbit_r248_c253 bl[253] br[253] wl[248] vdd gnd cell_6t
Xbit_r249_c253 bl[253] br[253] wl[249] vdd gnd cell_6t
Xbit_r250_c253 bl[253] br[253] wl[250] vdd gnd cell_6t
Xbit_r251_c253 bl[253] br[253] wl[251] vdd gnd cell_6t
Xbit_r252_c253 bl[253] br[253] wl[252] vdd gnd cell_6t
Xbit_r253_c253 bl[253] br[253] wl[253] vdd gnd cell_6t
Xbit_r254_c253 bl[253] br[253] wl[254] vdd gnd cell_6t
Xbit_r255_c253 bl[253] br[253] wl[255] vdd gnd cell_6t
Xbit_r0_c254 bl[254] br[254] wl[0] vdd gnd cell_6t
Xbit_r1_c254 bl[254] br[254] wl[1] vdd gnd cell_6t
Xbit_r2_c254 bl[254] br[254] wl[2] vdd gnd cell_6t
Xbit_r3_c254 bl[254] br[254] wl[3] vdd gnd cell_6t
Xbit_r4_c254 bl[254] br[254] wl[4] vdd gnd cell_6t
Xbit_r5_c254 bl[254] br[254] wl[5] vdd gnd cell_6t
Xbit_r6_c254 bl[254] br[254] wl[6] vdd gnd cell_6t
Xbit_r7_c254 bl[254] br[254] wl[7] vdd gnd cell_6t
Xbit_r8_c254 bl[254] br[254] wl[8] vdd gnd cell_6t
Xbit_r9_c254 bl[254] br[254] wl[9] vdd gnd cell_6t
Xbit_r10_c254 bl[254] br[254] wl[10] vdd gnd cell_6t
Xbit_r11_c254 bl[254] br[254] wl[11] vdd gnd cell_6t
Xbit_r12_c254 bl[254] br[254] wl[12] vdd gnd cell_6t
Xbit_r13_c254 bl[254] br[254] wl[13] vdd gnd cell_6t
Xbit_r14_c254 bl[254] br[254] wl[14] vdd gnd cell_6t
Xbit_r15_c254 bl[254] br[254] wl[15] vdd gnd cell_6t
Xbit_r16_c254 bl[254] br[254] wl[16] vdd gnd cell_6t
Xbit_r17_c254 bl[254] br[254] wl[17] vdd gnd cell_6t
Xbit_r18_c254 bl[254] br[254] wl[18] vdd gnd cell_6t
Xbit_r19_c254 bl[254] br[254] wl[19] vdd gnd cell_6t
Xbit_r20_c254 bl[254] br[254] wl[20] vdd gnd cell_6t
Xbit_r21_c254 bl[254] br[254] wl[21] vdd gnd cell_6t
Xbit_r22_c254 bl[254] br[254] wl[22] vdd gnd cell_6t
Xbit_r23_c254 bl[254] br[254] wl[23] vdd gnd cell_6t
Xbit_r24_c254 bl[254] br[254] wl[24] vdd gnd cell_6t
Xbit_r25_c254 bl[254] br[254] wl[25] vdd gnd cell_6t
Xbit_r26_c254 bl[254] br[254] wl[26] vdd gnd cell_6t
Xbit_r27_c254 bl[254] br[254] wl[27] vdd gnd cell_6t
Xbit_r28_c254 bl[254] br[254] wl[28] vdd gnd cell_6t
Xbit_r29_c254 bl[254] br[254] wl[29] vdd gnd cell_6t
Xbit_r30_c254 bl[254] br[254] wl[30] vdd gnd cell_6t
Xbit_r31_c254 bl[254] br[254] wl[31] vdd gnd cell_6t
Xbit_r32_c254 bl[254] br[254] wl[32] vdd gnd cell_6t
Xbit_r33_c254 bl[254] br[254] wl[33] vdd gnd cell_6t
Xbit_r34_c254 bl[254] br[254] wl[34] vdd gnd cell_6t
Xbit_r35_c254 bl[254] br[254] wl[35] vdd gnd cell_6t
Xbit_r36_c254 bl[254] br[254] wl[36] vdd gnd cell_6t
Xbit_r37_c254 bl[254] br[254] wl[37] vdd gnd cell_6t
Xbit_r38_c254 bl[254] br[254] wl[38] vdd gnd cell_6t
Xbit_r39_c254 bl[254] br[254] wl[39] vdd gnd cell_6t
Xbit_r40_c254 bl[254] br[254] wl[40] vdd gnd cell_6t
Xbit_r41_c254 bl[254] br[254] wl[41] vdd gnd cell_6t
Xbit_r42_c254 bl[254] br[254] wl[42] vdd gnd cell_6t
Xbit_r43_c254 bl[254] br[254] wl[43] vdd gnd cell_6t
Xbit_r44_c254 bl[254] br[254] wl[44] vdd gnd cell_6t
Xbit_r45_c254 bl[254] br[254] wl[45] vdd gnd cell_6t
Xbit_r46_c254 bl[254] br[254] wl[46] vdd gnd cell_6t
Xbit_r47_c254 bl[254] br[254] wl[47] vdd gnd cell_6t
Xbit_r48_c254 bl[254] br[254] wl[48] vdd gnd cell_6t
Xbit_r49_c254 bl[254] br[254] wl[49] vdd gnd cell_6t
Xbit_r50_c254 bl[254] br[254] wl[50] vdd gnd cell_6t
Xbit_r51_c254 bl[254] br[254] wl[51] vdd gnd cell_6t
Xbit_r52_c254 bl[254] br[254] wl[52] vdd gnd cell_6t
Xbit_r53_c254 bl[254] br[254] wl[53] vdd gnd cell_6t
Xbit_r54_c254 bl[254] br[254] wl[54] vdd gnd cell_6t
Xbit_r55_c254 bl[254] br[254] wl[55] vdd gnd cell_6t
Xbit_r56_c254 bl[254] br[254] wl[56] vdd gnd cell_6t
Xbit_r57_c254 bl[254] br[254] wl[57] vdd gnd cell_6t
Xbit_r58_c254 bl[254] br[254] wl[58] vdd gnd cell_6t
Xbit_r59_c254 bl[254] br[254] wl[59] vdd gnd cell_6t
Xbit_r60_c254 bl[254] br[254] wl[60] vdd gnd cell_6t
Xbit_r61_c254 bl[254] br[254] wl[61] vdd gnd cell_6t
Xbit_r62_c254 bl[254] br[254] wl[62] vdd gnd cell_6t
Xbit_r63_c254 bl[254] br[254] wl[63] vdd gnd cell_6t
Xbit_r64_c254 bl[254] br[254] wl[64] vdd gnd cell_6t
Xbit_r65_c254 bl[254] br[254] wl[65] vdd gnd cell_6t
Xbit_r66_c254 bl[254] br[254] wl[66] vdd gnd cell_6t
Xbit_r67_c254 bl[254] br[254] wl[67] vdd gnd cell_6t
Xbit_r68_c254 bl[254] br[254] wl[68] vdd gnd cell_6t
Xbit_r69_c254 bl[254] br[254] wl[69] vdd gnd cell_6t
Xbit_r70_c254 bl[254] br[254] wl[70] vdd gnd cell_6t
Xbit_r71_c254 bl[254] br[254] wl[71] vdd gnd cell_6t
Xbit_r72_c254 bl[254] br[254] wl[72] vdd gnd cell_6t
Xbit_r73_c254 bl[254] br[254] wl[73] vdd gnd cell_6t
Xbit_r74_c254 bl[254] br[254] wl[74] vdd gnd cell_6t
Xbit_r75_c254 bl[254] br[254] wl[75] vdd gnd cell_6t
Xbit_r76_c254 bl[254] br[254] wl[76] vdd gnd cell_6t
Xbit_r77_c254 bl[254] br[254] wl[77] vdd gnd cell_6t
Xbit_r78_c254 bl[254] br[254] wl[78] vdd gnd cell_6t
Xbit_r79_c254 bl[254] br[254] wl[79] vdd gnd cell_6t
Xbit_r80_c254 bl[254] br[254] wl[80] vdd gnd cell_6t
Xbit_r81_c254 bl[254] br[254] wl[81] vdd gnd cell_6t
Xbit_r82_c254 bl[254] br[254] wl[82] vdd gnd cell_6t
Xbit_r83_c254 bl[254] br[254] wl[83] vdd gnd cell_6t
Xbit_r84_c254 bl[254] br[254] wl[84] vdd gnd cell_6t
Xbit_r85_c254 bl[254] br[254] wl[85] vdd gnd cell_6t
Xbit_r86_c254 bl[254] br[254] wl[86] vdd gnd cell_6t
Xbit_r87_c254 bl[254] br[254] wl[87] vdd gnd cell_6t
Xbit_r88_c254 bl[254] br[254] wl[88] vdd gnd cell_6t
Xbit_r89_c254 bl[254] br[254] wl[89] vdd gnd cell_6t
Xbit_r90_c254 bl[254] br[254] wl[90] vdd gnd cell_6t
Xbit_r91_c254 bl[254] br[254] wl[91] vdd gnd cell_6t
Xbit_r92_c254 bl[254] br[254] wl[92] vdd gnd cell_6t
Xbit_r93_c254 bl[254] br[254] wl[93] vdd gnd cell_6t
Xbit_r94_c254 bl[254] br[254] wl[94] vdd gnd cell_6t
Xbit_r95_c254 bl[254] br[254] wl[95] vdd gnd cell_6t
Xbit_r96_c254 bl[254] br[254] wl[96] vdd gnd cell_6t
Xbit_r97_c254 bl[254] br[254] wl[97] vdd gnd cell_6t
Xbit_r98_c254 bl[254] br[254] wl[98] vdd gnd cell_6t
Xbit_r99_c254 bl[254] br[254] wl[99] vdd gnd cell_6t
Xbit_r100_c254 bl[254] br[254] wl[100] vdd gnd cell_6t
Xbit_r101_c254 bl[254] br[254] wl[101] vdd gnd cell_6t
Xbit_r102_c254 bl[254] br[254] wl[102] vdd gnd cell_6t
Xbit_r103_c254 bl[254] br[254] wl[103] vdd gnd cell_6t
Xbit_r104_c254 bl[254] br[254] wl[104] vdd gnd cell_6t
Xbit_r105_c254 bl[254] br[254] wl[105] vdd gnd cell_6t
Xbit_r106_c254 bl[254] br[254] wl[106] vdd gnd cell_6t
Xbit_r107_c254 bl[254] br[254] wl[107] vdd gnd cell_6t
Xbit_r108_c254 bl[254] br[254] wl[108] vdd gnd cell_6t
Xbit_r109_c254 bl[254] br[254] wl[109] vdd gnd cell_6t
Xbit_r110_c254 bl[254] br[254] wl[110] vdd gnd cell_6t
Xbit_r111_c254 bl[254] br[254] wl[111] vdd gnd cell_6t
Xbit_r112_c254 bl[254] br[254] wl[112] vdd gnd cell_6t
Xbit_r113_c254 bl[254] br[254] wl[113] vdd gnd cell_6t
Xbit_r114_c254 bl[254] br[254] wl[114] vdd gnd cell_6t
Xbit_r115_c254 bl[254] br[254] wl[115] vdd gnd cell_6t
Xbit_r116_c254 bl[254] br[254] wl[116] vdd gnd cell_6t
Xbit_r117_c254 bl[254] br[254] wl[117] vdd gnd cell_6t
Xbit_r118_c254 bl[254] br[254] wl[118] vdd gnd cell_6t
Xbit_r119_c254 bl[254] br[254] wl[119] vdd gnd cell_6t
Xbit_r120_c254 bl[254] br[254] wl[120] vdd gnd cell_6t
Xbit_r121_c254 bl[254] br[254] wl[121] vdd gnd cell_6t
Xbit_r122_c254 bl[254] br[254] wl[122] vdd gnd cell_6t
Xbit_r123_c254 bl[254] br[254] wl[123] vdd gnd cell_6t
Xbit_r124_c254 bl[254] br[254] wl[124] vdd gnd cell_6t
Xbit_r125_c254 bl[254] br[254] wl[125] vdd gnd cell_6t
Xbit_r126_c254 bl[254] br[254] wl[126] vdd gnd cell_6t
Xbit_r127_c254 bl[254] br[254] wl[127] vdd gnd cell_6t
Xbit_r128_c254 bl[254] br[254] wl[128] vdd gnd cell_6t
Xbit_r129_c254 bl[254] br[254] wl[129] vdd gnd cell_6t
Xbit_r130_c254 bl[254] br[254] wl[130] vdd gnd cell_6t
Xbit_r131_c254 bl[254] br[254] wl[131] vdd gnd cell_6t
Xbit_r132_c254 bl[254] br[254] wl[132] vdd gnd cell_6t
Xbit_r133_c254 bl[254] br[254] wl[133] vdd gnd cell_6t
Xbit_r134_c254 bl[254] br[254] wl[134] vdd gnd cell_6t
Xbit_r135_c254 bl[254] br[254] wl[135] vdd gnd cell_6t
Xbit_r136_c254 bl[254] br[254] wl[136] vdd gnd cell_6t
Xbit_r137_c254 bl[254] br[254] wl[137] vdd gnd cell_6t
Xbit_r138_c254 bl[254] br[254] wl[138] vdd gnd cell_6t
Xbit_r139_c254 bl[254] br[254] wl[139] vdd gnd cell_6t
Xbit_r140_c254 bl[254] br[254] wl[140] vdd gnd cell_6t
Xbit_r141_c254 bl[254] br[254] wl[141] vdd gnd cell_6t
Xbit_r142_c254 bl[254] br[254] wl[142] vdd gnd cell_6t
Xbit_r143_c254 bl[254] br[254] wl[143] vdd gnd cell_6t
Xbit_r144_c254 bl[254] br[254] wl[144] vdd gnd cell_6t
Xbit_r145_c254 bl[254] br[254] wl[145] vdd gnd cell_6t
Xbit_r146_c254 bl[254] br[254] wl[146] vdd gnd cell_6t
Xbit_r147_c254 bl[254] br[254] wl[147] vdd gnd cell_6t
Xbit_r148_c254 bl[254] br[254] wl[148] vdd gnd cell_6t
Xbit_r149_c254 bl[254] br[254] wl[149] vdd gnd cell_6t
Xbit_r150_c254 bl[254] br[254] wl[150] vdd gnd cell_6t
Xbit_r151_c254 bl[254] br[254] wl[151] vdd gnd cell_6t
Xbit_r152_c254 bl[254] br[254] wl[152] vdd gnd cell_6t
Xbit_r153_c254 bl[254] br[254] wl[153] vdd gnd cell_6t
Xbit_r154_c254 bl[254] br[254] wl[154] vdd gnd cell_6t
Xbit_r155_c254 bl[254] br[254] wl[155] vdd gnd cell_6t
Xbit_r156_c254 bl[254] br[254] wl[156] vdd gnd cell_6t
Xbit_r157_c254 bl[254] br[254] wl[157] vdd gnd cell_6t
Xbit_r158_c254 bl[254] br[254] wl[158] vdd gnd cell_6t
Xbit_r159_c254 bl[254] br[254] wl[159] vdd gnd cell_6t
Xbit_r160_c254 bl[254] br[254] wl[160] vdd gnd cell_6t
Xbit_r161_c254 bl[254] br[254] wl[161] vdd gnd cell_6t
Xbit_r162_c254 bl[254] br[254] wl[162] vdd gnd cell_6t
Xbit_r163_c254 bl[254] br[254] wl[163] vdd gnd cell_6t
Xbit_r164_c254 bl[254] br[254] wl[164] vdd gnd cell_6t
Xbit_r165_c254 bl[254] br[254] wl[165] vdd gnd cell_6t
Xbit_r166_c254 bl[254] br[254] wl[166] vdd gnd cell_6t
Xbit_r167_c254 bl[254] br[254] wl[167] vdd gnd cell_6t
Xbit_r168_c254 bl[254] br[254] wl[168] vdd gnd cell_6t
Xbit_r169_c254 bl[254] br[254] wl[169] vdd gnd cell_6t
Xbit_r170_c254 bl[254] br[254] wl[170] vdd gnd cell_6t
Xbit_r171_c254 bl[254] br[254] wl[171] vdd gnd cell_6t
Xbit_r172_c254 bl[254] br[254] wl[172] vdd gnd cell_6t
Xbit_r173_c254 bl[254] br[254] wl[173] vdd gnd cell_6t
Xbit_r174_c254 bl[254] br[254] wl[174] vdd gnd cell_6t
Xbit_r175_c254 bl[254] br[254] wl[175] vdd gnd cell_6t
Xbit_r176_c254 bl[254] br[254] wl[176] vdd gnd cell_6t
Xbit_r177_c254 bl[254] br[254] wl[177] vdd gnd cell_6t
Xbit_r178_c254 bl[254] br[254] wl[178] vdd gnd cell_6t
Xbit_r179_c254 bl[254] br[254] wl[179] vdd gnd cell_6t
Xbit_r180_c254 bl[254] br[254] wl[180] vdd gnd cell_6t
Xbit_r181_c254 bl[254] br[254] wl[181] vdd gnd cell_6t
Xbit_r182_c254 bl[254] br[254] wl[182] vdd gnd cell_6t
Xbit_r183_c254 bl[254] br[254] wl[183] vdd gnd cell_6t
Xbit_r184_c254 bl[254] br[254] wl[184] vdd gnd cell_6t
Xbit_r185_c254 bl[254] br[254] wl[185] vdd gnd cell_6t
Xbit_r186_c254 bl[254] br[254] wl[186] vdd gnd cell_6t
Xbit_r187_c254 bl[254] br[254] wl[187] vdd gnd cell_6t
Xbit_r188_c254 bl[254] br[254] wl[188] vdd gnd cell_6t
Xbit_r189_c254 bl[254] br[254] wl[189] vdd gnd cell_6t
Xbit_r190_c254 bl[254] br[254] wl[190] vdd gnd cell_6t
Xbit_r191_c254 bl[254] br[254] wl[191] vdd gnd cell_6t
Xbit_r192_c254 bl[254] br[254] wl[192] vdd gnd cell_6t
Xbit_r193_c254 bl[254] br[254] wl[193] vdd gnd cell_6t
Xbit_r194_c254 bl[254] br[254] wl[194] vdd gnd cell_6t
Xbit_r195_c254 bl[254] br[254] wl[195] vdd gnd cell_6t
Xbit_r196_c254 bl[254] br[254] wl[196] vdd gnd cell_6t
Xbit_r197_c254 bl[254] br[254] wl[197] vdd gnd cell_6t
Xbit_r198_c254 bl[254] br[254] wl[198] vdd gnd cell_6t
Xbit_r199_c254 bl[254] br[254] wl[199] vdd gnd cell_6t
Xbit_r200_c254 bl[254] br[254] wl[200] vdd gnd cell_6t
Xbit_r201_c254 bl[254] br[254] wl[201] vdd gnd cell_6t
Xbit_r202_c254 bl[254] br[254] wl[202] vdd gnd cell_6t
Xbit_r203_c254 bl[254] br[254] wl[203] vdd gnd cell_6t
Xbit_r204_c254 bl[254] br[254] wl[204] vdd gnd cell_6t
Xbit_r205_c254 bl[254] br[254] wl[205] vdd gnd cell_6t
Xbit_r206_c254 bl[254] br[254] wl[206] vdd gnd cell_6t
Xbit_r207_c254 bl[254] br[254] wl[207] vdd gnd cell_6t
Xbit_r208_c254 bl[254] br[254] wl[208] vdd gnd cell_6t
Xbit_r209_c254 bl[254] br[254] wl[209] vdd gnd cell_6t
Xbit_r210_c254 bl[254] br[254] wl[210] vdd gnd cell_6t
Xbit_r211_c254 bl[254] br[254] wl[211] vdd gnd cell_6t
Xbit_r212_c254 bl[254] br[254] wl[212] vdd gnd cell_6t
Xbit_r213_c254 bl[254] br[254] wl[213] vdd gnd cell_6t
Xbit_r214_c254 bl[254] br[254] wl[214] vdd gnd cell_6t
Xbit_r215_c254 bl[254] br[254] wl[215] vdd gnd cell_6t
Xbit_r216_c254 bl[254] br[254] wl[216] vdd gnd cell_6t
Xbit_r217_c254 bl[254] br[254] wl[217] vdd gnd cell_6t
Xbit_r218_c254 bl[254] br[254] wl[218] vdd gnd cell_6t
Xbit_r219_c254 bl[254] br[254] wl[219] vdd gnd cell_6t
Xbit_r220_c254 bl[254] br[254] wl[220] vdd gnd cell_6t
Xbit_r221_c254 bl[254] br[254] wl[221] vdd gnd cell_6t
Xbit_r222_c254 bl[254] br[254] wl[222] vdd gnd cell_6t
Xbit_r223_c254 bl[254] br[254] wl[223] vdd gnd cell_6t
Xbit_r224_c254 bl[254] br[254] wl[224] vdd gnd cell_6t
Xbit_r225_c254 bl[254] br[254] wl[225] vdd gnd cell_6t
Xbit_r226_c254 bl[254] br[254] wl[226] vdd gnd cell_6t
Xbit_r227_c254 bl[254] br[254] wl[227] vdd gnd cell_6t
Xbit_r228_c254 bl[254] br[254] wl[228] vdd gnd cell_6t
Xbit_r229_c254 bl[254] br[254] wl[229] vdd gnd cell_6t
Xbit_r230_c254 bl[254] br[254] wl[230] vdd gnd cell_6t
Xbit_r231_c254 bl[254] br[254] wl[231] vdd gnd cell_6t
Xbit_r232_c254 bl[254] br[254] wl[232] vdd gnd cell_6t
Xbit_r233_c254 bl[254] br[254] wl[233] vdd gnd cell_6t
Xbit_r234_c254 bl[254] br[254] wl[234] vdd gnd cell_6t
Xbit_r235_c254 bl[254] br[254] wl[235] vdd gnd cell_6t
Xbit_r236_c254 bl[254] br[254] wl[236] vdd gnd cell_6t
Xbit_r237_c254 bl[254] br[254] wl[237] vdd gnd cell_6t
Xbit_r238_c254 bl[254] br[254] wl[238] vdd gnd cell_6t
Xbit_r239_c254 bl[254] br[254] wl[239] vdd gnd cell_6t
Xbit_r240_c254 bl[254] br[254] wl[240] vdd gnd cell_6t
Xbit_r241_c254 bl[254] br[254] wl[241] vdd gnd cell_6t
Xbit_r242_c254 bl[254] br[254] wl[242] vdd gnd cell_6t
Xbit_r243_c254 bl[254] br[254] wl[243] vdd gnd cell_6t
Xbit_r244_c254 bl[254] br[254] wl[244] vdd gnd cell_6t
Xbit_r245_c254 bl[254] br[254] wl[245] vdd gnd cell_6t
Xbit_r246_c254 bl[254] br[254] wl[246] vdd gnd cell_6t
Xbit_r247_c254 bl[254] br[254] wl[247] vdd gnd cell_6t
Xbit_r248_c254 bl[254] br[254] wl[248] vdd gnd cell_6t
Xbit_r249_c254 bl[254] br[254] wl[249] vdd gnd cell_6t
Xbit_r250_c254 bl[254] br[254] wl[250] vdd gnd cell_6t
Xbit_r251_c254 bl[254] br[254] wl[251] vdd gnd cell_6t
Xbit_r252_c254 bl[254] br[254] wl[252] vdd gnd cell_6t
Xbit_r253_c254 bl[254] br[254] wl[253] vdd gnd cell_6t
Xbit_r254_c254 bl[254] br[254] wl[254] vdd gnd cell_6t
Xbit_r255_c254 bl[254] br[254] wl[255] vdd gnd cell_6t
Xbit_r0_c255 bl[255] br[255] wl[0] vdd gnd cell_6t
Xbit_r1_c255 bl[255] br[255] wl[1] vdd gnd cell_6t
Xbit_r2_c255 bl[255] br[255] wl[2] vdd gnd cell_6t
Xbit_r3_c255 bl[255] br[255] wl[3] vdd gnd cell_6t
Xbit_r4_c255 bl[255] br[255] wl[4] vdd gnd cell_6t
Xbit_r5_c255 bl[255] br[255] wl[5] vdd gnd cell_6t
Xbit_r6_c255 bl[255] br[255] wl[6] vdd gnd cell_6t
Xbit_r7_c255 bl[255] br[255] wl[7] vdd gnd cell_6t
Xbit_r8_c255 bl[255] br[255] wl[8] vdd gnd cell_6t
Xbit_r9_c255 bl[255] br[255] wl[9] vdd gnd cell_6t
Xbit_r10_c255 bl[255] br[255] wl[10] vdd gnd cell_6t
Xbit_r11_c255 bl[255] br[255] wl[11] vdd gnd cell_6t
Xbit_r12_c255 bl[255] br[255] wl[12] vdd gnd cell_6t
Xbit_r13_c255 bl[255] br[255] wl[13] vdd gnd cell_6t
Xbit_r14_c255 bl[255] br[255] wl[14] vdd gnd cell_6t
Xbit_r15_c255 bl[255] br[255] wl[15] vdd gnd cell_6t
Xbit_r16_c255 bl[255] br[255] wl[16] vdd gnd cell_6t
Xbit_r17_c255 bl[255] br[255] wl[17] vdd gnd cell_6t
Xbit_r18_c255 bl[255] br[255] wl[18] vdd gnd cell_6t
Xbit_r19_c255 bl[255] br[255] wl[19] vdd gnd cell_6t
Xbit_r20_c255 bl[255] br[255] wl[20] vdd gnd cell_6t
Xbit_r21_c255 bl[255] br[255] wl[21] vdd gnd cell_6t
Xbit_r22_c255 bl[255] br[255] wl[22] vdd gnd cell_6t
Xbit_r23_c255 bl[255] br[255] wl[23] vdd gnd cell_6t
Xbit_r24_c255 bl[255] br[255] wl[24] vdd gnd cell_6t
Xbit_r25_c255 bl[255] br[255] wl[25] vdd gnd cell_6t
Xbit_r26_c255 bl[255] br[255] wl[26] vdd gnd cell_6t
Xbit_r27_c255 bl[255] br[255] wl[27] vdd gnd cell_6t
Xbit_r28_c255 bl[255] br[255] wl[28] vdd gnd cell_6t
Xbit_r29_c255 bl[255] br[255] wl[29] vdd gnd cell_6t
Xbit_r30_c255 bl[255] br[255] wl[30] vdd gnd cell_6t
Xbit_r31_c255 bl[255] br[255] wl[31] vdd gnd cell_6t
Xbit_r32_c255 bl[255] br[255] wl[32] vdd gnd cell_6t
Xbit_r33_c255 bl[255] br[255] wl[33] vdd gnd cell_6t
Xbit_r34_c255 bl[255] br[255] wl[34] vdd gnd cell_6t
Xbit_r35_c255 bl[255] br[255] wl[35] vdd gnd cell_6t
Xbit_r36_c255 bl[255] br[255] wl[36] vdd gnd cell_6t
Xbit_r37_c255 bl[255] br[255] wl[37] vdd gnd cell_6t
Xbit_r38_c255 bl[255] br[255] wl[38] vdd gnd cell_6t
Xbit_r39_c255 bl[255] br[255] wl[39] vdd gnd cell_6t
Xbit_r40_c255 bl[255] br[255] wl[40] vdd gnd cell_6t
Xbit_r41_c255 bl[255] br[255] wl[41] vdd gnd cell_6t
Xbit_r42_c255 bl[255] br[255] wl[42] vdd gnd cell_6t
Xbit_r43_c255 bl[255] br[255] wl[43] vdd gnd cell_6t
Xbit_r44_c255 bl[255] br[255] wl[44] vdd gnd cell_6t
Xbit_r45_c255 bl[255] br[255] wl[45] vdd gnd cell_6t
Xbit_r46_c255 bl[255] br[255] wl[46] vdd gnd cell_6t
Xbit_r47_c255 bl[255] br[255] wl[47] vdd gnd cell_6t
Xbit_r48_c255 bl[255] br[255] wl[48] vdd gnd cell_6t
Xbit_r49_c255 bl[255] br[255] wl[49] vdd gnd cell_6t
Xbit_r50_c255 bl[255] br[255] wl[50] vdd gnd cell_6t
Xbit_r51_c255 bl[255] br[255] wl[51] vdd gnd cell_6t
Xbit_r52_c255 bl[255] br[255] wl[52] vdd gnd cell_6t
Xbit_r53_c255 bl[255] br[255] wl[53] vdd gnd cell_6t
Xbit_r54_c255 bl[255] br[255] wl[54] vdd gnd cell_6t
Xbit_r55_c255 bl[255] br[255] wl[55] vdd gnd cell_6t
Xbit_r56_c255 bl[255] br[255] wl[56] vdd gnd cell_6t
Xbit_r57_c255 bl[255] br[255] wl[57] vdd gnd cell_6t
Xbit_r58_c255 bl[255] br[255] wl[58] vdd gnd cell_6t
Xbit_r59_c255 bl[255] br[255] wl[59] vdd gnd cell_6t
Xbit_r60_c255 bl[255] br[255] wl[60] vdd gnd cell_6t
Xbit_r61_c255 bl[255] br[255] wl[61] vdd gnd cell_6t
Xbit_r62_c255 bl[255] br[255] wl[62] vdd gnd cell_6t
Xbit_r63_c255 bl[255] br[255] wl[63] vdd gnd cell_6t
Xbit_r64_c255 bl[255] br[255] wl[64] vdd gnd cell_6t
Xbit_r65_c255 bl[255] br[255] wl[65] vdd gnd cell_6t
Xbit_r66_c255 bl[255] br[255] wl[66] vdd gnd cell_6t
Xbit_r67_c255 bl[255] br[255] wl[67] vdd gnd cell_6t
Xbit_r68_c255 bl[255] br[255] wl[68] vdd gnd cell_6t
Xbit_r69_c255 bl[255] br[255] wl[69] vdd gnd cell_6t
Xbit_r70_c255 bl[255] br[255] wl[70] vdd gnd cell_6t
Xbit_r71_c255 bl[255] br[255] wl[71] vdd gnd cell_6t
Xbit_r72_c255 bl[255] br[255] wl[72] vdd gnd cell_6t
Xbit_r73_c255 bl[255] br[255] wl[73] vdd gnd cell_6t
Xbit_r74_c255 bl[255] br[255] wl[74] vdd gnd cell_6t
Xbit_r75_c255 bl[255] br[255] wl[75] vdd gnd cell_6t
Xbit_r76_c255 bl[255] br[255] wl[76] vdd gnd cell_6t
Xbit_r77_c255 bl[255] br[255] wl[77] vdd gnd cell_6t
Xbit_r78_c255 bl[255] br[255] wl[78] vdd gnd cell_6t
Xbit_r79_c255 bl[255] br[255] wl[79] vdd gnd cell_6t
Xbit_r80_c255 bl[255] br[255] wl[80] vdd gnd cell_6t
Xbit_r81_c255 bl[255] br[255] wl[81] vdd gnd cell_6t
Xbit_r82_c255 bl[255] br[255] wl[82] vdd gnd cell_6t
Xbit_r83_c255 bl[255] br[255] wl[83] vdd gnd cell_6t
Xbit_r84_c255 bl[255] br[255] wl[84] vdd gnd cell_6t
Xbit_r85_c255 bl[255] br[255] wl[85] vdd gnd cell_6t
Xbit_r86_c255 bl[255] br[255] wl[86] vdd gnd cell_6t
Xbit_r87_c255 bl[255] br[255] wl[87] vdd gnd cell_6t
Xbit_r88_c255 bl[255] br[255] wl[88] vdd gnd cell_6t
Xbit_r89_c255 bl[255] br[255] wl[89] vdd gnd cell_6t
Xbit_r90_c255 bl[255] br[255] wl[90] vdd gnd cell_6t
Xbit_r91_c255 bl[255] br[255] wl[91] vdd gnd cell_6t
Xbit_r92_c255 bl[255] br[255] wl[92] vdd gnd cell_6t
Xbit_r93_c255 bl[255] br[255] wl[93] vdd gnd cell_6t
Xbit_r94_c255 bl[255] br[255] wl[94] vdd gnd cell_6t
Xbit_r95_c255 bl[255] br[255] wl[95] vdd gnd cell_6t
Xbit_r96_c255 bl[255] br[255] wl[96] vdd gnd cell_6t
Xbit_r97_c255 bl[255] br[255] wl[97] vdd gnd cell_6t
Xbit_r98_c255 bl[255] br[255] wl[98] vdd gnd cell_6t
Xbit_r99_c255 bl[255] br[255] wl[99] vdd gnd cell_6t
Xbit_r100_c255 bl[255] br[255] wl[100] vdd gnd cell_6t
Xbit_r101_c255 bl[255] br[255] wl[101] vdd gnd cell_6t
Xbit_r102_c255 bl[255] br[255] wl[102] vdd gnd cell_6t
Xbit_r103_c255 bl[255] br[255] wl[103] vdd gnd cell_6t
Xbit_r104_c255 bl[255] br[255] wl[104] vdd gnd cell_6t
Xbit_r105_c255 bl[255] br[255] wl[105] vdd gnd cell_6t
Xbit_r106_c255 bl[255] br[255] wl[106] vdd gnd cell_6t
Xbit_r107_c255 bl[255] br[255] wl[107] vdd gnd cell_6t
Xbit_r108_c255 bl[255] br[255] wl[108] vdd gnd cell_6t
Xbit_r109_c255 bl[255] br[255] wl[109] vdd gnd cell_6t
Xbit_r110_c255 bl[255] br[255] wl[110] vdd gnd cell_6t
Xbit_r111_c255 bl[255] br[255] wl[111] vdd gnd cell_6t
Xbit_r112_c255 bl[255] br[255] wl[112] vdd gnd cell_6t
Xbit_r113_c255 bl[255] br[255] wl[113] vdd gnd cell_6t
Xbit_r114_c255 bl[255] br[255] wl[114] vdd gnd cell_6t
Xbit_r115_c255 bl[255] br[255] wl[115] vdd gnd cell_6t
Xbit_r116_c255 bl[255] br[255] wl[116] vdd gnd cell_6t
Xbit_r117_c255 bl[255] br[255] wl[117] vdd gnd cell_6t
Xbit_r118_c255 bl[255] br[255] wl[118] vdd gnd cell_6t
Xbit_r119_c255 bl[255] br[255] wl[119] vdd gnd cell_6t
Xbit_r120_c255 bl[255] br[255] wl[120] vdd gnd cell_6t
Xbit_r121_c255 bl[255] br[255] wl[121] vdd gnd cell_6t
Xbit_r122_c255 bl[255] br[255] wl[122] vdd gnd cell_6t
Xbit_r123_c255 bl[255] br[255] wl[123] vdd gnd cell_6t
Xbit_r124_c255 bl[255] br[255] wl[124] vdd gnd cell_6t
Xbit_r125_c255 bl[255] br[255] wl[125] vdd gnd cell_6t
Xbit_r126_c255 bl[255] br[255] wl[126] vdd gnd cell_6t
Xbit_r127_c255 bl[255] br[255] wl[127] vdd gnd cell_6t
Xbit_r128_c255 bl[255] br[255] wl[128] vdd gnd cell_6t
Xbit_r129_c255 bl[255] br[255] wl[129] vdd gnd cell_6t
Xbit_r130_c255 bl[255] br[255] wl[130] vdd gnd cell_6t
Xbit_r131_c255 bl[255] br[255] wl[131] vdd gnd cell_6t
Xbit_r132_c255 bl[255] br[255] wl[132] vdd gnd cell_6t
Xbit_r133_c255 bl[255] br[255] wl[133] vdd gnd cell_6t
Xbit_r134_c255 bl[255] br[255] wl[134] vdd gnd cell_6t
Xbit_r135_c255 bl[255] br[255] wl[135] vdd gnd cell_6t
Xbit_r136_c255 bl[255] br[255] wl[136] vdd gnd cell_6t
Xbit_r137_c255 bl[255] br[255] wl[137] vdd gnd cell_6t
Xbit_r138_c255 bl[255] br[255] wl[138] vdd gnd cell_6t
Xbit_r139_c255 bl[255] br[255] wl[139] vdd gnd cell_6t
Xbit_r140_c255 bl[255] br[255] wl[140] vdd gnd cell_6t
Xbit_r141_c255 bl[255] br[255] wl[141] vdd gnd cell_6t
Xbit_r142_c255 bl[255] br[255] wl[142] vdd gnd cell_6t
Xbit_r143_c255 bl[255] br[255] wl[143] vdd gnd cell_6t
Xbit_r144_c255 bl[255] br[255] wl[144] vdd gnd cell_6t
Xbit_r145_c255 bl[255] br[255] wl[145] vdd gnd cell_6t
Xbit_r146_c255 bl[255] br[255] wl[146] vdd gnd cell_6t
Xbit_r147_c255 bl[255] br[255] wl[147] vdd gnd cell_6t
Xbit_r148_c255 bl[255] br[255] wl[148] vdd gnd cell_6t
Xbit_r149_c255 bl[255] br[255] wl[149] vdd gnd cell_6t
Xbit_r150_c255 bl[255] br[255] wl[150] vdd gnd cell_6t
Xbit_r151_c255 bl[255] br[255] wl[151] vdd gnd cell_6t
Xbit_r152_c255 bl[255] br[255] wl[152] vdd gnd cell_6t
Xbit_r153_c255 bl[255] br[255] wl[153] vdd gnd cell_6t
Xbit_r154_c255 bl[255] br[255] wl[154] vdd gnd cell_6t
Xbit_r155_c255 bl[255] br[255] wl[155] vdd gnd cell_6t
Xbit_r156_c255 bl[255] br[255] wl[156] vdd gnd cell_6t
Xbit_r157_c255 bl[255] br[255] wl[157] vdd gnd cell_6t
Xbit_r158_c255 bl[255] br[255] wl[158] vdd gnd cell_6t
Xbit_r159_c255 bl[255] br[255] wl[159] vdd gnd cell_6t
Xbit_r160_c255 bl[255] br[255] wl[160] vdd gnd cell_6t
Xbit_r161_c255 bl[255] br[255] wl[161] vdd gnd cell_6t
Xbit_r162_c255 bl[255] br[255] wl[162] vdd gnd cell_6t
Xbit_r163_c255 bl[255] br[255] wl[163] vdd gnd cell_6t
Xbit_r164_c255 bl[255] br[255] wl[164] vdd gnd cell_6t
Xbit_r165_c255 bl[255] br[255] wl[165] vdd gnd cell_6t
Xbit_r166_c255 bl[255] br[255] wl[166] vdd gnd cell_6t
Xbit_r167_c255 bl[255] br[255] wl[167] vdd gnd cell_6t
Xbit_r168_c255 bl[255] br[255] wl[168] vdd gnd cell_6t
Xbit_r169_c255 bl[255] br[255] wl[169] vdd gnd cell_6t
Xbit_r170_c255 bl[255] br[255] wl[170] vdd gnd cell_6t
Xbit_r171_c255 bl[255] br[255] wl[171] vdd gnd cell_6t
Xbit_r172_c255 bl[255] br[255] wl[172] vdd gnd cell_6t
Xbit_r173_c255 bl[255] br[255] wl[173] vdd gnd cell_6t
Xbit_r174_c255 bl[255] br[255] wl[174] vdd gnd cell_6t
Xbit_r175_c255 bl[255] br[255] wl[175] vdd gnd cell_6t
Xbit_r176_c255 bl[255] br[255] wl[176] vdd gnd cell_6t
Xbit_r177_c255 bl[255] br[255] wl[177] vdd gnd cell_6t
Xbit_r178_c255 bl[255] br[255] wl[178] vdd gnd cell_6t
Xbit_r179_c255 bl[255] br[255] wl[179] vdd gnd cell_6t
Xbit_r180_c255 bl[255] br[255] wl[180] vdd gnd cell_6t
Xbit_r181_c255 bl[255] br[255] wl[181] vdd gnd cell_6t
Xbit_r182_c255 bl[255] br[255] wl[182] vdd gnd cell_6t
Xbit_r183_c255 bl[255] br[255] wl[183] vdd gnd cell_6t
Xbit_r184_c255 bl[255] br[255] wl[184] vdd gnd cell_6t
Xbit_r185_c255 bl[255] br[255] wl[185] vdd gnd cell_6t
Xbit_r186_c255 bl[255] br[255] wl[186] vdd gnd cell_6t
Xbit_r187_c255 bl[255] br[255] wl[187] vdd gnd cell_6t
Xbit_r188_c255 bl[255] br[255] wl[188] vdd gnd cell_6t
Xbit_r189_c255 bl[255] br[255] wl[189] vdd gnd cell_6t
Xbit_r190_c255 bl[255] br[255] wl[190] vdd gnd cell_6t
Xbit_r191_c255 bl[255] br[255] wl[191] vdd gnd cell_6t
Xbit_r192_c255 bl[255] br[255] wl[192] vdd gnd cell_6t
Xbit_r193_c255 bl[255] br[255] wl[193] vdd gnd cell_6t
Xbit_r194_c255 bl[255] br[255] wl[194] vdd gnd cell_6t
Xbit_r195_c255 bl[255] br[255] wl[195] vdd gnd cell_6t
Xbit_r196_c255 bl[255] br[255] wl[196] vdd gnd cell_6t
Xbit_r197_c255 bl[255] br[255] wl[197] vdd gnd cell_6t
Xbit_r198_c255 bl[255] br[255] wl[198] vdd gnd cell_6t
Xbit_r199_c255 bl[255] br[255] wl[199] vdd gnd cell_6t
Xbit_r200_c255 bl[255] br[255] wl[200] vdd gnd cell_6t
Xbit_r201_c255 bl[255] br[255] wl[201] vdd gnd cell_6t
Xbit_r202_c255 bl[255] br[255] wl[202] vdd gnd cell_6t
Xbit_r203_c255 bl[255] br[255] wl[203] vdd gnd cell_6t
Xbit_r204_c255 bl[255] br[255] wl[204] vdd gnd cell_6t
Xbit_r205_c255 bl[255] br[255] wl[205] vdd gnd cell_6t
Xbit_r206_c255 bl[255] br[255] wl[206] vdd gnd cell_6t
Xbit_r207_c255 bl[255] br[255] wl[207] vdd gnd cell_6t
Xbit_r208_c255 bl[255] br[255] wl[208] vdd gnd cell_6t
Xbit_r209_c255 bl[255] br[255] wl[209] vdd gnd cell_6t
Xbit_r210_c255 bl[255] br[255] wl[210] vdd gnd cell_6t
Xbit_r211_c255 bl[255] br[255] wl[211] vdd gnd cell_6t
Xbit_r212_c255 bl[255] br[255] wl[212] vdd gnd cell_6t
Xbit_r213_c255 bl[255] br[255] wl[213] vdd gnd cell_6t
Xbit_r214_c255 bl[255] br[255] wl[214] vdd gnd cell_6t
Xbit_r215_c255 bl[255] br[255] wl[215] vdd gnd cell_6t
Xbit_r216_c255 bl[255] br[255] wl[216] vdd gnd cell_6t
Xbit_r217_c255 bl[255] br[255] wl[217] vdd gnd cell_6t
Xbit_r218_c255 bl[255] br[255] wl[218] vdd gnd cell_6t
Xbit_r219_c255 bl[255] br[255] wl[219] vdd gnd cell_6t
Xbit_r220_c255 bl[255] br[255] wl[220] vdd gnd cell_6t
Xbit_r221_c255 bl[255] br[255] wl[221] vdd gnd cell_6t
Xbit_r222_c255 bl[255] br[255] wl[222] vdd gnd cell_6t
Xbit_r223_c255 bl[255] br[255] wl[223] vdd gnd cell_6t
Xbit_r224_c255 bl[255] br[255] wl[224] vdd gnd cell_6t
Xbit_r225_c255 bl[255] br[255] wl[225] vdd gnd cell_6t
Xbit_r226_c255 bl[255] br[255] wl[226] vdd gnd cell_6t
Xbit_r227_c255 bl[255] br[255] wl[227] vdd gnd cell_6t
Xbit_r228_c255 bl[255] br[255] wl[228] vdd gnd cell_6t
Xbit_r229_c255 bl[255] br[255] wl[229] vdd gnd cell_6t
Xbit_r230_c255 bl[255] br[255] wl[230] vdd gnd cell_6t
Xbit_r231_c255 bl[255] br[255] wl[231] vdd gnd cell_6t
Xbit_r232_c255 bl[255] br[255] wl[232] vdd gnd cell_6t
Xbit_r233_c255 bl[255] br[255] wl[233] vdd gnd cell_6t
Xbit_r234_c255 bl[255] br[255] wl[234] vdd gnd cell_6t
Xbit_r235_c255 bl[255] br[255] wl[235] vdd gnd cell_6t
Xbit_r236_c255 bl[255] br[255] wl[236] vdd gnd cell_6t
Xbit_r237_c255 bl[255] br[255] wl[237] vdd gnd cell_6t
Xbit_r238_c255 bl[255] br[255] wl[238] vdd gnd cell_6t
Xbit_r239_c255 bl[255] br[255] wl[239] vdd gnd cell_6t
Xbit_r240_c255 bl[255] br[255] wl[240] vdd gnd cell_6t
Xbit_r241_c255 bl[255] br[255] wl[241] vdd gnd cell_6t
Xbit_r242_c255 bl[255] br[255] wl[242] vdd gnd cell_6t
Xbit_r243_c255 bl[255] br[255] wl[243] vdd gnd cell_6t
Xbit_r244_c255 bl[255] br[255] wl[244] vdd gnd cell_6t
Xbit_r245_c255 bl[255] br[255] wl[245] vdd gnd cell_6t
Xbit_r246_c255 bl[255] br[255] wl[246] vdd gnd cell_6t
Xbit_r247_c255 bl[255] br[255] wl[247] vdd gnd cell_6t
Xbit_r248_c255 bl[255] br[255] wl[248] vdd gnd cell_6t
Xbit_r249_c255 bl[255] br[255] wl[249] vdd gnd cell_6t
Xbit_r250_c255 bl[255] br[255] wl[250] vdd gnd cell_6t
Xbit_r251_c255 bl[255] br[255] wl[251] vdd gnd cell_6t
Xbit_r252_c255 bl[255] br[255] wl[252] vdd gnd cell_6t
Xbit_r253_c255 bl[255] br[255] wl[253] vdd gnd cell_6t
Xbit_r254_c255 bl[255] br[255] wl[254] vdd gnd cell_6t
Xbit_r255_c255 bl[255] br[255] wl[255] vdd gnd cell_6t
.ENDS bitcell_array

* ptx M{0} {1} p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p

.SUBCKT precharge bl br en vdd
Mlower_pmos bl en BR vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mupper_pmos1 bl en vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mupper_pmos2 br en vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
.ENDS precharge

.SUBCKT precharge_array bl[0] br[0] bl[1] br[1] bl[2] br[2] bl[3] br[3] bl[4] br[4] bl[5] br[5] bl[6] br[6] bl[7] br[7] bl[8] br[8] bl[9] br[9] bl[10] br[10] bl[11] br[11] bl[12] br[12] bl[13] br[13] bl[14] br[14] bl[15] br[15] bl[16] br[16] bl[17] br[17] bl[18] br[18] bl[19] br[19] bl[20] br[20] bl[21] br[21] bl[22] br[22] bl[23] br[23] bl[24] br[24] bl[25] br[25] bl[26] br[26] bl[27] br[27] bl[28] br[28] bl[29] br[29] bl[30] br[30] bl[31] br[31] bl[32] br[32] bl[33] br[33] bl[34] br[34] bl[35] br[35] bl[36] br[36] bl[37] br[37] bl[38] br[38] bl[39] br[39] bl[40] br[40] bl[41] br[41] bl[42] br[42] bl[43] br[43] bl[44] br[44] bl[45] br[45] bl[46] br[46] bl[47] br[47] bl[48] br[48] bl[49] br[49] bl[50] br[50] bl[51] br[51] bl[52] br[52] bl[53] br[53] bl[54] br[54] bl[55] br[55] bl[56] br[56] bl[57] br[57] bl[58] br[58] bl[59] br[59] bl[60] br[60] bl[61] br[61] bl[62] br[62] bl[63] br[63] bl[64] br[64] bl[65] br[65] bl[66] br[66] bl[67] br[67] bl[68] br[68] bl[69] br[69] bl[70] br[70] bl[71] br[71] bl[72] br[72] bl[73] br[73] bl[74] br[74] bl[75] br[75] bl[76] br[76] bl[77] br[77] bl[78] br[78] bl[79] br[79] bl[80] br[80] bl[81] br[81] bl[82] br[82] bl[83] br[83] bl[84] br[84] bl[85] br[85] bl[86] br[86] bl[87] br[87] bl[88] br[88] bl[89] br[89] bl[90] br[90] bl[91] br[91] bl[92] br[92] bl[93] br[93] bl[94] br[94] bl[95] br[95] bl[96] br[96] bl[97] br[97] bl[98] br[98] bl[99] br[99] bl[100] br[100] bl[101] br[101] bl[102] br[102] bl[103] br[103] bl[104] br[104] bl[105] br[105] bl[106] br[106] bl[107] br[107] bl[108] br[108] bl[109] br[109] bl[110] br[110] bl[111] br[111] bl[112] br[112] bl[113] br[113] bl[114] br[114] bl[115] br[115] bl[116] br[116] bl[117] br[117] bl[118] br[118] bl[119] br[119] bl[120] br[120] bl[121] br[121] bl[122] br[122] bl[123] br[123] bl[124] br[124] bl[125] br[125] bl[126] br[126] bl[127] br[127] bl[128] br[128] bl[129] br[129] bl[130] br[130] bl[131] br[131] bl[132] br[132] bl[133] br[133] bl[134] br[134] bl[135] br[135] bl[136] br[136] bl[137] br[137] bl[138] br[138] bl[139] br[139] bl[140] br[140] bl[141] br[141] bl[142] br[142] bl[143] br[143] bl[144] br[144] bl[145] br[145] bl[146] br[146] bl[147] br[147] bl[148] br[148] bl[149] br[149] bl[150] br[150] bl[151] br[151] bl[152] br[152] bl[153] br[153] bl[154] br[154] bl[155] br[155] bl[156] br[156] bl[157] br[157] bl[158] br[158] bl[159] br[159] bl[160] br[160] bl[161] br[161] bl[162] br[162] bl[163] br[163] bl[164] br[164] bl[165] br[165] bl[166] br[166] bl[167] br[167] bl[168] br[168] bl[169] br[169] bl[170] br[170] bl[171] br[171] bl[172] br[172] bl[173] br[173] bl[174] br[174] bl[175] br[175] bl[176] br[176] bl[177] br[177] bl[178] br[178] bl[179] br[179] bl[180] br[180] bl[181] br[181] bl[182] br[182] bl[183] br[183] bl[184] br[184] bl[185] br[185] bl[186] br[186] bl[187] br[187] bl[188] br[188] bl[189] br[189] bl[190] br[190] bl[191] br[191] bl[192] br[192] bl[193] br[193] bl[194] br[194] bl[195] br[195] bl[196] br[196] bl[197] br[197] bl[198] br[198] bl[199] br[199] bl[200] br[200] bl[201] br[201] bl[202] br[202] bl[203] br[203] bl[204] br[204] bl[205] br[205] bl[206] br[206] bl[207] br[207] bl[208] br[208] bl[209] br[209] bl[210] br[210] bl[211] br[211] bl[212] br[212] bl[213] br[213] bl[214] br[214] bl[215] br[215] bl[216] br[216] bl[217] br[217] bl[218] br[218] bl[219] br[219] bl[220] br[220] bl[221] br[221] bl[222] br[222] bl[223] br[223] bl[224] br[224] bl[225] br[225] bl[226] br[226] bl[227] br[227] bl[228] br[228] bl[229] br[229] bl[230] br[230] bl[231] br[231] bl[232] br[232] bl[233] br[233] bl[234] br[234] bl[235] br[235] bl[236] br[236] bl[237] br[237] bl[238] br[238] bl[239] br[239] bl[240] br[240] bl[241] br[241] bl[242] br[242] bl[243] br[243] bl[244] br[244] bl[245] br[245] bl[246] br[246] bl[247] br[247] bl[248] br[248] bl[249] br[249] bl[250] br[250] bl[251] br[251] bl[252] br[252] bl[253] br[253] bl[254] br[254] bl[255] br[255] en vdd
Xpre_column_0 bl[0] br[0] en vdd precharge
Xpre_column_1 bl[1] br[1] en vdd precharge
Xpre_column_2 bl[2] br[2] en vdd precharge
Xpre_column_3 bl[3] br[3] en vdd precharge
Xpre_column_4 bl[4] br[4] en vdd precharge
Xpre_column_5 bl[5] br[5] en vdd precharge
Xpre_column_6 bl[6] br[6] en vdd precharge
Xpre_column_7 bl[7] br[7] en vdd precharge
Xpre_column_8 bl[8] br[8] en vdd precharge
Xpre_column_9 bl[9] br[9] en vdd precharge
Xpre_column_10 bl[10] br[10] en vdd precharge
Xpre_column_11 bl[11] br[11] en vdd precharge
Xpre_column_12 bl[12] br[12] en vdd precharge
Xpre_column_13 bl[13] br[13] en vdd precharge
Xpre_column_14 bl[14] br[14] en vdd precharge
Xpre_column_15 bl[15] br[15] en vdd precharge
Xpre_column_16 bl[16] br[16] en vdd precharge
Xpre_column_17 bl[17] br[17] en vdd precharge
Xpre_column_18 bl[18] br[18] en vdd precharge
Xpre_column_19 bl[19] br[19] en vdd precharge
Xpre_column_20 bl[20] br[20] en vdd precharge
Xpre_column_21 bl[21] br[21] en vdd precharge
Xpre_column_22 bl[22] br[22] en vdd precharge
Xpre_column_23 bl[23] br[23] en vdd precharge
Xpre_column_24 bl[24] br[24] en vdd precharge
Xpre_column_25 bl[25] br[25] en vdd precharge
Xpre_column_26 bl[26] br[26] en vdd precharge
Xpre_column_27 bl[27] br[27] en vdd precharge
Xpre_column_28 bl[28] br[28] en vdd precharge
Xpre_column_29 bl[29] br[29] en vdd precharge
Xpre_column_30 bl[30] br[30] en vdd precharge
Xpre_column_31 bl[31] br[31] en vdd precharge
Xpre_column_32 bl[32] br[32] en vdd precharge
Xpre_column_33 bl[33] br[33] en vdd precharge
Xpre_column_34 bl[34] br[34] en vdd precharge
Xpre_column_35 bl[35] br[35] en vdd precharge
Xpre_column_36 bl[36] br[36] en vdd precharge
Xpre_column_37 bl[37] br[37] en vdd precharge
Xpre_column_38 bl[38] br[38] en vdd precharge
Xpre_column_39 bl[39] br[39] en vdd precharge
Xpre_column_40 bl[40] br[40] en vdd precharge
Xpre_column_41 bl[41] br[41] en vdd precharge
Xpre_column_42 bl[42] br[42] en vdd precharge
Xpre_column_43 bl[43] br[43] en vdd precharge
Xpre_column_44 bl[44] br[44] en vdd precharge
Xpre_column_45 bl[45] br[45] en vdd precharge
Xpre_column_46 bl[46] br[46] en vdd precharge
Xpre_column_47 bl[47] br[47] en vdd precharge
Xpre_column_48 bl[48] br[48] en vdd precharge
Xpre_column_49 bl[49] br[49] en vdd precharge
Xpre_column_50 bl[50] br[50] en vdd precharge
Xpre_column_51 bl[51] br[51] en vdd precharge
Xpre_column_52 bl[52] br[52] en vdd precharge
Xpre_column_53 bl[53] br[53] en vdd precharge
Xpre_column_54 bl[54] br[54] en vdd precharge
Xpre_column_55 bl[55] br[55] en vdd precharge
Xpre_column_56 bl[56] br[56] en vdd precharge
Xpre_column_57 bl[57] br[57] en vdd precharge
Xpre_column_58 bl[58] br[58] en vdd precharge
Xpre_column_59 bl[59] br[59] en vdd precharge
Xpre_column_60 bl[60] br[60] en vdd precharge
Xpre_column_61 bl[61] br[61] en vdd precharge
Xpre_column_62 bl[62] br[62] en vdd precharge
Xpre_column_63 bl[63] br[63] en vdd precharge
Xpre_column_64 bl[64] br[64] en vdd precharge
Xpre_column_65 bl[65] br[65] en vdd precharge
Xpre_column_66 bl[66] br[66] en vdd precharge
Xpre_column_67 bl[67] br[67] en vdd precharge
Xpre_column_68 bl[68] br[68] en vdd precharge
Xpre_column_69 bl[69] br[69] en vdd precharge
Xpre_column_70 bl[70] br[70] en vdd precharge
Xpre_column_71 bl[71] br[71] en vdd precharge
Xpre_column_72 bl[72] br[72] en vdd precharge
Xpre_column_73 bl[73] br[73] en vdd precharge
Xpre_column_74 bl[74] br[74] en vdd precharge
Xpre_column_75 bl[75] br[75] en vdd precharge
Xpre_column_76 bl[76] br[76] en vdd precharge
Xpre_column_77 bl[77] br[77] en vdd precharge
Xpre_column_78 bl[78] br[78] en vdd precharge
Xpre_column_79 bl[79] br[79] en vdd precharge
Xpre_column_80 bl[80] br[80] en vdd precharge
Xpre_column_81 bl[81] br[81] en vdd precharge
Xpre_column_82 bl[82] br[82] en vdd precharge
Xpre_column_83 bl[83] br[83] en vdd precharge
Xpre_column_84 bl[84] br[84] en vdd precharge
Xpre_column_85 bl[85] br[85] en vdd precharge
Xpre_column_86 bl[86] br[86] en vdd precharge
Xpre_column_87 bl[87] br[87] en vdd precharge
Xpre_column_88 bl[88] br[88] en vdd precharge
Xpre_column_89 bl[89] br[89] en vdd precharge
Xpre_column_90 bl[90] br[90] en vdd precharge
Xpre_column_91 bl[91] br[91] en vdd precharge
Xpre_column_92 bl[92] br[92] en vdd precharge
Xpre_column_93 bl[93] br[93] en vdd precharge
Xpre_column_94 bl[94] br[94] en vdd precharge
Xpre_column_95 bl[95] br[95] en vdd precharge
Xpre_column_96 bl[96] br[96] en vdd precharge
Xpre_column_97 bl[97] br[97] en vdd precharge
Xpre_column_98 bl[98] br[98] en vdd precharge
Xpre_column_99 bl[99] br[99] en vdd precharge
Xpre_column_100 bl[100] br[100] en vdd precharge
Xpre_column_101 bl[101] br[101] en vdd precharge
Xpre_column_102 bl[102] br[102] en vdd precharge
Xpre_column_103 bl[103] br[103] en vdd precharge
Xpre_column_104 bl[104] br[104] en vdd precharge
Xpre_column_105 bl[105] br[105] en vdd precharge
Xpre_column_106 bl[106] br[106] en vdd precharge
Xpre_column_107 bl[107] br[107] en vdd precharge
Xpre_column_108 bl[108] br[108] en vdd precharge
Xpre_column_109 bl[109] br[109] en vdd precharge
Xpre_column_110 bl[110] br[110] en vdd precharge
Xpre_column_111 bl[111] br[111] en vdd precharge
Xpre_column_112 bl[112] br[112] en vdd precharge
Xpre_column_113 bl[113] br[113] en vdd precharge
Xpre_column_114 bl[114] br[114] en vdd precharge
Xpre_column_115 bl[115] br[115] en vdd precharge
Xpre_column_116 bl[116] br[116] en vdd precharge
Xpre_column_117 bl[117] br[117] en vdd precharge
Xpre_column_118 bl[118] br[118] en vdd precharge
Xpre_column_119 bl[119] br[119] en vdd precharge
Xpre_column_120 bl[120] br[120] en vdd precharge
Xpre_column_121 bl[121] br[121] en vdd precharge
Xpre_column_122 bl[122] br[122] en vdd precharge
Xpre_column_123 bl[123] br[123] en vdd precharge
Xpre_column_124 bl[124] br[124] en vdd precharge
Xpre_column_125 bl[125] br[125] en vdd precharge
Xpre_column_126 bl[126] br[126] en vdd precharge
Xpre_column_127 bl[127] br[127] en vdd precharge
Xpre_column_128 bl[128] br[128] en vdd precharge
Xpre_column_129 bl[129] br[129] en vdd precharge
Xpre_column_130 bl[130] br[130] en vdd precharge
Xpre_column_131 bl[131] br[131] en vdd precharge
Xpre_column_132 bl[132] br[132] en vdd precharge
Xpre_column_133 bl[133] br[133] en vdd precharge
Xpre_column_134 bl[134] br[134] en vdd precharge
Xpre_column_135 bl[135] br[135] en vdd precharge
Xpre_column_136 bl[136] br[136] en vdd precharge
Xpre_column_137 bl[137] br[137] en vdd precharge
Xpre_column_138 bl[138] br[138] en vdd precharge
Xpre_column_139 bl[139] br[139] en vdd precharge
Xpre_column_140 bl[140] br[140] en vdd precharge
Xpre_column_141 bl[141] br[141] en vdd precharge
Xpre_column_142 bl[142] br[142] en vdd precharge
Xpre_column_143 bl[143] br[143] en vdd precharge
Xpre_column_144 bl[144] br[144] en vdd precharge
Xpre_column_145 bl[145] br[145] en vdd precharge
Xpre_column_146 bl[146] br[146] en vdd precharge
Xpre_column_147 bl[147] br[147] en vdd precharge
Xpre_column_148 bl[148] br[148] en vdd precharge
Xpre_column_149 bl[149] br[149] en vdd precharge
Xpre_column_150 bl[150] br[150] en vdd precharge
Xpre_column_151 bl[151] br[151] en vdd precharge
Xpre_column_152 bl[152] br[152] en vdd precharge
Xpre_column_153 bl[153] br[153] en vdd precharge
Xpre_column_154 bl[154] br[154] en vdd precharge
Xpre_column_155 bl[155] br[155] en vdd precharge
Xpre_column_156 bl[156] br[156] en vdd precharge
Xpre_column_157 bl[157] br[157] en vdd precharge
Xpre_column_158 bl[158] br[158] en vdd precharge
Xpre_column_159 bl[159] br[159] en vdd precharge
Xpre_column_160 bl[160] br[160] en vdd precharge
Xpre_column_161 bl[161] br[161] en vdd precharge
Xpre_column_162 bl[162] br[162] en vdd precharge
Xpre_column_163 bl[163] br[163] en vdd precharge
Xpre_column_164 bl[164] br[164] en vdd precharge
Xpre_column_165 bl[165] br[165] en vdd precharge
Xpre_column_166 bl[166] br[166] en vdd precharge
Xpre_column_167 bl[167] br[167] en vdd precharge
Xpre_column_168 bl[168] br[168] en vdd precharge
Xpre_column_169 bl[169] br[169] en vdd precharge
Xpre_column_170 bl[170] br[170] en vdd precharge
Xpre_column_171 bl[171] br[171] en vdd precharge
Xpre_column_172 bl[172] br[172] en vdd precharge
Xpre_column_173 bl[173] br[173] en vdd precharge
Xpre_column_174 bl[174] br[174] en vdd precharge
Xpre_column_175 bl[175] br[175] en vdd precharge
Xpre_column_176 bl[176] br[176] en vdd precharge
Xpre_column_177 bl[177] br[177] en vdd precharge
Xpre_column_178 bl[178] br[178] en vdd precharge
Xpre_column_179 bl[179] br[179] en vdd precharge
Xpre_column_180 bl[180] br[180] en vdd precharge
Xpre_column_181 bl[181] br[181] en vdd precharge
Xpre_column_182 bl[182] br[182] en vdd precharge
Xpre_column_183 bl[183] br[183] en vdd precharge
Xpre_column_184 bl[184] br[184] en vdd precharge
Xpre_column_185 bl[185] br[185] en vdd precharge
Xpre_column_186 bl[186] br[186] en vdd precharge
Xpre_column_187 bl[187] br[187] en vdd precharge
Xpre_column_188 bl[188] br[188] en vdd precharge
Xpre_column_189 bl[189] br[189] en vdd precharge
Xpre_column_190 bl[190] br[190] en vdd precharge
Xpre_column_191 bl[191] br[191] en vdd precharge
Xpre_column_192 bl[192] br[192] en vdd precharge
Xpre_column_193 bl[193] br[193] en vdd precharge
Xpre_column_194 bl[194] br[194] en vdd precharge
Xpre_column_195 bl[195] br[195] en vdd precharge
Xpre_column_196 bl[196] br[196] en vdd precharge
Xpre_column_197 bl[197] br[197] en vdd precharge
Xpre_column_198 bl[198] br[198] en vdd precharge
Xpre_column_199 bl[199] br[199] en vdd precharge
Xpre_column_200 bl[200] br[200] en vdd precharge
Xpre_column_201 bl[201] br[201] en vdd precharge
Xpre_column_202 bl[202] br[202] en vdd precharge
Xpre_column_203 bl[203] br[203] en vdd precharge
Xpre_column_204 bl[204] br[204] en vdd precharge
Xpre_column_205 bl[205] br[205] en vdd precharge
Xpre_column_206 bl[206] br[206] en vdd precharge
Xpre_column_207 bl[207] br[207] en vdd precharge
Xpre_column_208 bl[208] br[208] en vdd precharge
Xpre_column_209 bl[209] br[209] en vdd precharge
Xpre_column_210 bl[210] br[210] en vdd precharge
Xpre_column_211 bl[211] br[211] en vdd precharge
Xpre_column_212 bl[212] br[212] en vdd precharge
Xpre_column_213 bl[213] br[213] en vdd precharge
Xpre_column_214 bl[214] br[214] en vdd precharge
Xpre_column_215 bl[215] br[215] en vdd precharge
Xpre_column_216 bl[216] br[216] en vdd precharge
Xpre_column_217 bl[217] br[217] en vdd precharge
Xpre_column_218 bl[218] br[218] en vdd precharge
Xpre_column_219 bl[219] br[219] en vdd precharge
Xpre_column_220 bl[220] br[220] en vdd precharge
Xpre_column_221 bl[221] br[221] en vdd precharge
Xpre_column_222 bl[222] br[222] en vdd precharge
Xpre_column_223 bl[223] br[223] en vdd precharge
Xpre_column_224 bl[224] br[224] en vdd precharge
Xpre_column_225 bl[225] br[225] en vdd precharge
Xpre_column_226 bl[226] br[226] en vdd precharge
Xpre_column_227 bl[227] br[227] en vdd precharge
Xpre_column_228 bl[228] br[228] en vdd precharge
Xpre_column_229 bl[229] br[229] en vdd precharge
Xpre_column_230 bl[230] br[230] en vdd precharge
Xpre_column_231 bl[231] br[231] en vdd precharge
Xpre_column_232 bl[232] br[232] en vdd precharge
Xpre_column_233 bl[233] br[233] en vdd precharge
Xpre_column_234 bl[234] br[234] en vdd precharge
Xpre_column_235 bl[235] br[235] en vdd precharge
Xpre_column_236 bl[236] br[236] en vdd precharge
Xpre_column_237 bl[237] br[237] en vdd precharge
Xpre_column_238 bl[238] br[238] en vdd precharge
Xpre_column_239 bl[239] br[239] en vdd precharge
Xpre_column_240 bl[240] br[240] en vdd precharge
Xpre_column_241 bl[241] br[241] en vdd precharge
Xpre_column_242 bl[242] br[242] en vdd precharge
Xpre_column_243 bl[243] br[243] en vdd precharge
Xpre_column_244 bl[244] br[244] en vdd precharge
Xpre_column_245 bl[245] br[245] en vdd precharge
Xpre_column_246 bl[246] br[246] en vdd precharge
Xpre_column_247 bl[247] br[247] en vdd precharge
Xpre_column_248 bl[248] br[248] en vdd precharge
Xpre_column_249 bl[249] br[249] en vdd precharge
Xpre_column_250 bl[250] br[250] en vdd precharge
Xpre_column_251 bl[251] br[251] en vdd precharge
Xpre_column_252 bl[252] br[252] en vdd precharge
Xpre_column_253 bl[253] br[253] en vdd precharge
Xpre_column_254 bl[254] br[254] en vdd precharge
Xpre_column_255 bl[255] br[255] en vdd precharge
.ENDS precharge_array

* ptx M{0} {1} n m=1 w=9.6u l=0.6u pd=20.4u ps=20.4u as=14.4p ad=14.4p

.SUBCKT single_level_column_mux_8 bl br bl_out br_out sel gnd
Mmux_tx1 bl sel bl_out gnd n m=1 w=9.6u l=0.6u pd=20.4u ps=20.4u as=14.4p ad=14.4p
Mmux_tx2 br sel br_out gnd n m=1 w=9.6u l=0.6u pd=20.4u ps=20.4u as=14.4p ad=14.4p
.ENDS single_level_column_mux_8

.SUBCKT columnmux_array bl[0] br[0] bl[1] br[1] bl[2] br[2] bl[3] br[3] bl[4] br[4] bl[5] br[5] bl[6] br[6] bl[7] br[7] bl[8] br[8] bl[9] br[9] bl[10] br[10] bl[11] br[11] bl[12] br[12] bl[13] br[13] bl[14] br[14] bl[15] br[15] bl[16] br[16] bl[17] br[17] bl[18] br[18] bl[19] br[19] bl[20] br[20] bl[21] br[21] bl[22] br[22] bl[23] br[23] bl[24] br[24] bl[25] br[25] bl[26] br[26] bl[27] br[27] bl[28] br[28] bl[29] br[29] bl[30] br[30] bl[31] br[31] bl[32] br[32] bl[33] br[33] bl[34] br[34] bl[35] br[35] bl[36] br[36] bl[37] br[37] bl[38] br[38] bl[39] br[39] bl[40] br[40] bl[41] br[41] bl[42] br[42] bl[43] br[43] bl[44] br[44] bl[45] br[45] bl[46] br[46] bl[47] br[47] bl[48] br[48] bl[49] br[49] bl[50] br[50] bl[51] br[51] bl[52] br[52] bl[53] br[53] bl[54] br[54] bl[55] br[55] bl[56] br[56] bl[57] br[57] bl[58] br[58] bl[59] br[59] bl[60] br[60] bl[61] br[61] bl[62] br[62] bl[63] br[63] bl[64] br[64] bl[65] br[65] bl[66] br[66] bl[67] br[67] bl[68] br[68] bl[69] br[69] bl[70] br[70] bl[71] br[71] bl[72] br[72] bl[73] br[73] bl[74] br[74] bl[75] br[75] bl[76] br[76] bl[77] br[77] bl[78] br[78] bl[79] br[79] bl[80] br[80] bl[81] br[81] bl[82] br[82] bl[83] br[83] bl[84] br[84] bl[85] br[85] bl[86] br[86] bl[87] br[87] bl[88] br[88] bl[89] br[89] bl[90] br[90] bl[91] br[91] bl[92] br[92] bl[93] br[93] bl[94] br[94] bl[95] br[95] bl[96] br[96] bl[97] br[97] bl[98] br[98] bl[99] br[99] bl[100] br[100] bl[101] br[101] bl[102] br[102] bl[103] br[103] bl[104] br[104] bl[105] br[105] bl[106] br[106] bl[107] br[107] bl[108] br[108] bl[109] br[109] bl[110] br[110] bl[111] br[111] bl[112] br[112] bl[113] br[113] bl[114] br[114] bl[115] br[115] bl[116] br[116] bl[117] br[117] bl[118] br[118] bl[119] br[119] bl[120] br[120] bl[121] br[121] bl[122] br[122] bl[123] br[123] bl[124] br[124] bl[125] br[125] bl[126] br[126] bl[127] br[127] bl[128] br[128] bl[129] br[129] bl[130] br[130] bl[131] br[131] bl[132] br[132] bl[133] br[133] bl[134] br[134] bl[135] br[135] bl[136] br[136] bl[137] br[137] bl[138] br[138] bl[139] br[139] bl[140] br[140] bl[141] br[141] bl[142] br[142] bl[143] br[143] bl[144] br[144] bl[145] br[145] bl[146] br[146] bl[147] br[147] bl[148] br[148] bl[149] br[149] bl[150] br[150] bl[151] br[151] bl[152] br[152] bl[153] br[153] bl[154] br[154] bl[155] br[155] bl[156] br[156] bl[157] br[157] bl[158] br[158] bl[159] br[159] bl[160] br[160] bl[161] br[161] bl[162] br[162] bl[163] br[163] bl[164] br[164] bl[165] br[165] bl[166] br[166] bl[167] br[167] bl[168] br[168] bl[169] br[169] bl[170] br[170] bl[171] br[171] bl[172] br[172] bl[173] br[173] bl[174] br[174] bl[175] br[175] bl[176] br[176] bl[177] br[177] bl[178] br[178] bl[179] br[179] bl[180] br[180] bl[181] br[181] bl[182] br[182] bl[183] br[183] bl[184] br[184] bl[185] br[185] bl[186] br[186] bl[187] br[187] bl[188] br[188] bl[189] br[189] bl[190] br[190] bl[191] br[191] bl[192] br[192] bl[193] br[193] bl[194] br[194] bl[195] br[195] bl[196] br[196] bl[197] br[197] bl[198] br[198] bl[199] br[199] bl[200] br[200] bl[201] br[201] bl[202] br[202] bl[203] br[203] bl[204] br[204] bl[205] br[205] bl[206] br[206] bl[207] br[207] bl[208] br[208] bl[209] br[209] bl[210] br[210] bl[211] br[211] bl[212] br[212] bl[213] br[213] bl[214] br[214] bl[215] br[215] bl[216] br[216] bl[217] br[217] bl[218] br[218] bl[219] br[219] bl[220] br[220] bl[221] br[221] bl[222] br[222] bl[223] br[223] bl[224] br[224] bl[225] br[225] bl[226] br[226] bl[227] br[227] bl[228] br[228] bl[229] br[229] bl[230] br[230] bl[231] br[231] bl[232] br[232] bl[233] br[233] bl[234] br[234] bl[235] br[235] bl[236] br[236] bl[237] br[237] bl[238] br[238] bl[239] br[239] bl[240] br[240] bl[241] br[241] bl[242] br[242] bl[243] br[243] bl[244] br[244] bl[245] br[245] bl[246] br[246] bl[247] br[247] bl[248] br[248] bl[249] br[249] bl[250] br[250] bl[251] br[251] bl[252] br[252] bl[253] br[253] bl[254] br[254] bl[255] br[255] sel[0] sel[1] bl_out[0] br_out[0] bl_out[1] br_out[1] bl_out[2] br_out[2] bl_out[3] br_out[3] bl_out[4] br_out[4] bl_out[5] br_out[5] bl_out[6] br_out[6] bl_out[7] br_out[7] bl_out[8] br_out[8] bl_out[9] br_out[9] bl_out[10] br_out[10] bl_out[11] br_out[11] bl_out[12] br_out[12] bl_out[13] br_out[13] bl_out[14] br_out[14] bl_out[15] br_out[15] bl_out[16] br_out[16] bl_out[17] br_out[17] bl_out[18] br_out[18] bl_out[19] br_out[19] bl_out[20] br_out[20] bl_out[21] br_out[21] bl_out[22] br_out[22] bl_out[23] br_out[23] bl_out[24] br_out[24] bl_out[25] br_out[25] bl_out[26] br_out[26] bl_out[27] br_out[27] bl_out[28] br_out[28] bl_out[29] br_out[29] bl_out[30] br_out[30] bl_out[31] br_out[31] bl_out[32] br_out[32] bl_out[33] br_out[33] bl_out[34] br_out[34] bl_out[35] br_out[35] bl_out[36] br_out[36] bl_out[37] br_out[37] bl_out[38] br_out[38] bl_out[39] br_out[39] bl_out[40] br_out[40] bl_out[41] br_out[41] bl_out[42] br_out[42] bl_out[43] br_out[43] bl_out[44] br_out[44] bl_out[45] br_out[45] bl_out[46] br_out[46] bl_out[47] br_out[47] bl_out[48] br_out[48] bl_out[49] br_out[49] bl_out[50] br_out[50] bl_out[51] br_out[51] bl_out[52] br_out[52] bl_out[53] br_out[53] bl_out[54] br_out[54] bl_out[55] br_out[55] bl_out[56] br_out[56] bl_out[57] br_out[57] bl_out[58] br_out[58] bl_out[59] br_out[59] bl_out[60] br_out[60] bl_out[61] br_out[61] bl_out[62] br_out[62] bl_out[63] br_out[63] bl_out[64] br_out[64] bl_out[65] br_out[65] bl_out[66] br_out[66] bl_out[67] br_out[67] bl_out[68] br_out[68] bl_out[69] br_out[69] bl_out[70] br_out[70] bl_out[71] br_out[71] bl_out[72] br_out[72] bl_out[73] br_out[73] bl_out[74] br_out[74] bl_out[75] br_out[75] bl_out[76] br_out[76] bl_out[77] br_out[77] bl_out[78] br_out[78] bl_out[79] br_out[79] bl_out[80] br_out[80] bl_out[81] br_out[81] bl_out[82] br_out[82] bl_out[83] br_out[83] bl_out[84] br_out[84] bl_out[85] br_out[85] bl_out[86] br_out[86] bl_out[87] br_out[87] bl_out[88] br_out[88] bl_out[89] br_out[89] bl_out[90] br_out[90] bl_out[91] br_out[91] bl_out[92] br_out[92] bl_out[93] br_out[93] bl_out[94] br_out[94] bl_out[95] br_out[95] bl_out[96] br_out[96] bl_out[97] br_out[97] bl_out[98] br_out[98] bl_out[99] br_out[99] bl_out[100] br_out[100] bl_out[101] br_out[101] bl_out[102] br_out[102] bl_out[103] br_out[103] bl_out[104] br_out[104] bl_out[105] br_out[105] bl_out[106] br_out[106] bl_out[107] br_out[107] bl_out[108] br_out[108] bl_out[109] br_out[109] bl_out[110] br_out[110] bl_out[111] br_out[111] bl_out[112] br_out[112] bl_out[113] br_out[113] bl_out[114] br_out[114] bl_out[115] br_out[115] bl_out[116] br_out[116] bl_out[117] br_out[117] bl_out[118] br_out[118] bl_out[119] br_out[119] bl_out[120] br_out[120] bl_out[121] br_out[121] bl_out[122] br_out[122] bl_out[123] br_out[123] bl_out[124] br_out[124] bl_out[125] br_out[125] bl_out[126] br_out[126] bl_out[127] br_out[127] gnd
XXMUX0 bl[0] br[0] bl_out[0] br_out[0] sel[0] gnd single_level_column_mux_8
XXMUX1 bl[1] br[1] bl_out[0] br_out[0] sel[1] gnd single_level_column_mux_8
XXMUX2 bl[2] br[2] bl_out[1] br_out[1] sel[0] gnd single_level_column_mux_8
XXMUX3 bl[3] br[3] bl_out[1] br_out[1] sel[1] gnd single_level_column_mux_8
XXMUX4 bl[4] br[4] bl_out[2] br_out[2] sel[0] gnd single_level_column_mux_8
XXMUX5 bl[5] br[5] bl_out[2] br_out[2] sel[1] gnd single_level_column_mux_8
XXMUX6 bl[6] br[6] bl_out[3] br_out[3] sel[0] gnd single_level_column_mux_8
XXMUX7 bl[7] br[7] bl_out[3] br_out[3] sel[1] gnd single_level_column_mux_8
XXMUX8 bl[8] br[8] bl_out[4] br_out[4] sel[0] gnd single_level_column_mux_8
XXMUX9 bl[9] br[9] bl_out[4] br_out[4] sel[1] gnd single_level_column_mux_8
XXMUX10 bl[10] br[10] bl_out[5] br_out[5] sel[0] gnd single_level_column_mux_8
XXMUX11 bl[11] br[11] bl_out[5] br_out[5] sel[1] gnd single_level_column_mux_8
XXMUX12 bl[12] br[12] bl_out[6] br_out[6] sel[0] gnd single_level_column_mux_8
XXMUX13 bl[13] br[13] bl_out[6] br_out[6] sel[1] gnd single_level_column_mux_8
XXMUX14 bl[14] br[14] bl_out[7] br_out[7] sel[0] gnd single_level_column_mux_8
XXMUX15 bl[15] br[15] bl_out[7] br_out[7] sel[1] gnd single_level_column_mux_8
XXMUX16 bl[16] br[16] bl_out[8] br_out[8] sel[0] gnd single_level_column_mux_8
XXMUX17 bl[17] br[17] bl_out[8] br_out[8] sel[1] gnd single_level_column_mux_8
XXMUX18 bl[18] br[18] bl_out[9] br_out[9] sel[0] gnd single_level_column_mux_8
XXMUX19 bl[19] br[19] bl_out[9] br_out[9] sel[1] gnd single_level_column_mux_8
XXMUX20 bl[20] br[20] bl_out[10] br_out[10] sel[0] gnd single_level_column_mux_8
XXMUX21 bl[21] br[21] bl_out[10] br_out[10] sel[1] gnd single_level_column_mux_8
XXMUX22 bl[22] br[22] bl_out[11] br_out[11] sel[0] gnd single_level_column_mux_8
XXMUX23 bl[23] br[23] bl_out[11] br_out[11] sel[1] gnd single_level_column_mux_8
XXMUX24 bl[24] br[24] bl_out[12] br_out[12] sel[0] gnd single_level_column_mux_8
XXMUX25 bl[25] br[25] bl_out[12] br_out[12] sel[1] gnd single_level_column_mux_8
XXMUX26 bl[26] br[26] bl_out[13] br_out[13] sel[0] gnd single_level_column_mux_8
XXMUX27 bl[27] br[27] bl_out[13] br_out[13] sel[1] gnd single_level_column_mux_8
XXMUX28 bl[28] br[28] bl_out[14] br_out[14] sel[0] gnd single_level_column_mux_8
XXMUX29 bl[29] br[29] bl_out[14] br_out[14] sel[1] gnd single_level_column_mux_8
XXMUX30 bl[30] br[30] bl_out[15] br_out[15] sel[0] gnd single_level_column_mux_8
XXMUX31 bl[31] br[31] bl_out[15] br_out[15] sel[1] gnd single_level_column_mux_8
XXMUX32 bl[32] br[32] bl_out[16] br_out[16] sel[0] gnd single_level_column_mux_8
XXMUX33 bl[33] br[33] bl_out[16] br_out[16] sel[1] gnd single_level_column_mux_8
XXMUX34 bl[34] br[34] bl_out[17] br_out[17] sel[0] gnd single_level_column_mux_8
XXMUX35 bl[35] br[35] bl_out[17] br_out[17] sel[1] gnd single_level_column_mux_8
XXMUX36 bl[36] br[36] bl_out[18] br_out[18] sel[0] gnd single_level_column_mux_8
XXMUX37 bl[37] br[37] bl_out[18] br_out[18] sel[1] gnd single_level_column_mux_8
XXMUX38 bl[38] br[38] bl_out[19] br_out[19] sel[0] gnd single_level_column_mux_8
XXMUX39 bl[39] br[39] bl_out[19] br_out[19] sel[1] gnd single_level_column_mux_8
XXMUX40 bl[40] br[40] bl_out[20] br_out[20] sel[0] gnd single_level_column_mux_8
XXMUX41 bl[41] br[41] bl_out[20] br_out[20] sel[1] gnd single_level_column_mux_8
XXMUX42 bl[42] br[42] bl_out[21] br_out[21] sel[0] gnd single_level_column_mux_8
XXMUX43 bl[43] br[43] bl_out[21] br_out[21] sel[1] gnd single_level_column_mux_8
XXMUX44 bl[44] br[44] bl_out[22] br_out[22] sel[0] gnd single_level_column_mux_8
XXMUX45 bl[45] br[45] bl_out[22] br_out[22] sel[1] gnd single_level_column_mux_8
XXMUX46 bl[46] br[46] bl_out[23] br_out[23] sel[0] gnd single_level_column_mux_8
XXMUX47 bl[47] br[47] bl_out[23] br_out[23] sel[1] gnd single_level_column_mux_8
XXMUX48 bl[48] br[48] bl_out[24] br_out[24] sel[0] gnd single_level_column_mux_8
XXMUX49 bl[49] br[49] bl_out[24] br_out[24] sel[1] gnd single_level_column_mux_8
XXMUX50 bl[50] br[50] bl_out[25] br_out[25] sel[0] gnd single_level_column_mux_8
XXMUX51 bl[51] br[51] bl_out[25] br_out[25] sel[1] gnd single_level_column_mux_8
XXMUX52 bl[52] br[52] bl_out[26] br_out[26] sel[0] gnd single_level_column_mux_8
XXMUX53 bl[53] br[53] bl_out[26] br_out[26] sel[1] gnd single_level_column_mux_8
XXMUX54 bl[54] br[54] bl_out[27] br_out[27] sel[0] gnd single_level_column_mux_8
XXMUX55 bl[55] br[55] bl_out[27] br_out[27] sel[1] gnd single_level_column_mux_8
XXMUX56 bl[56] br[56] bl_out[28] br_out[28] sel[0] gnd single_level_column_mux_8
XXMUX57 bl[57] br[57] bl_out[28] br_out[28] sel[1] gnd single_level_column_mux_8
XXMUX58 bl[58] br[58] bl_out[29] br_out[29] sel[0] gnd single_level_column_mux_8
XXMUX59 bl[59] br[59] bl_out[29] br_out[29] sel[1] gnd single_level_column_mux_8
XXMUX60 bl[60] br[60] bl_out[30] br_out[30] sel[0] gnd single_level_column_mux_8
XXMUX61 bl[61] br[61] bl_out[30] br_out[30] sel[1] gnd single_level_column_mux_8
XXMUX62 bl[62] br[62] bl_out[31] br_out[31] sel[0] gnd single_level_column_mux_8
XXMUX63 bl[63] br[63] bl_out[31] br_out[31] sel[1] gnd single_level_column_mux_8
XXMUX64 bl[64] br[64] bl_out[32] br_out[32] sel[0] gnd single_level_column_mux_8
XXMUX65 bl[65] br[65] bl_out[32] br_out[32] sel[1] gnd single_level_column_mux_8
XXMUX66 bl[66] br[66] bl_out[33] br_out[33] sel[0] gnd single_level_column_mux_8
XXMUX67 bl[67] br[67] bl_out[33] br_out[33] sel[1] gnd single_level_column_mux_8
XXMUX68 bl[68] br[68] bl_out[34] br_out[34] sel[0] gnd single_level_column_mux_8
XXMUX69 bl[69] br[69] bl_out[34] br_out[34] sel[1] gnd single_level_column_mux_8
XXMUX70 bl[70] br[70] bl_out[35] br_out[35] sel[0] gnd single_level_column_mux_8
XXMUX71 bl[71] br[71] bl_out[35] br_out[35] sel[1] gnd single_level_column_mux_8
XXMUX72 bl[72] br[72] bl_out[36] br_out[36] sel[0] gnd single_level_column_mux_8
XXMUX73 bl[73] br[73] bl_out[36] br_out[36] sel[1] gnd single_level_column_mux_8
XXMUX74 bl[74] br[74] bl_out[37] br_out[37] sel[0] gnd single_level_column_mux_8
XXMUX75 bl[75] br[75] bl_out[37] br_out[37] sel[1] gnd single_level_column_mux_8
XXMUX76 bl[76] br[76] bl_out[38] br_out[38] sel[0] gnd single_level_column_mux_8
XXMUX77 bl[77] br[77] bl_out[38] br_out[38] sel[1] gnd single_level_column_mux_8
XXMUX78 bl[78] br[78] bl_out[39] br_out[39] sel[0] gnd single_level_column_mux_8
XXMUX79 bl[79] br[79] bl_out[39] br_out[39] sel[1] gnd single_level_column_mux_8
XXMUX80 bl[80] br[80] bl_out[40] br_out[40] sel[0] gnd single_level_column_mux_8
XXMUX81 bl[81] br[81] bl_out[40] br_out[40] sel[1] gnd single_level_column_mux_8
XXMUX82 bl[82] br[82] bl_out[41] br_out[41] sel[0] gnd single_level_column_mux_8
XXMUX83 bl[83] br[83] bl_out[41] br_out[41] sel[1] gnd single_level_column_mux_8
XXMUX84 bl[84] br[84] bl_out[42] br_out[42] sel[0] gnd single_level_column_mux_8
XXMUX85 bl[85] br[85] bl_out[42] br_out[42] sel[1] gnd single_level_column_mux_8
XXMUX86 bl[86] br[86] bl_out[43] br_out[43] sel[0] gnd single_level_column_mux_8
XXMUX87 bl[87] br[87] bl_out[43] br_out[43] sel[1] gnd single_level_column_mux_8
XXMUX88 bl[88] br[88] bl_out[44] br_out[44] sel[0] gnd single_level_column_mux_8
XXMUX89 bl[89] br[89] bl_out[44] br_out[44] sel[1] gnd single_level_column_mux_8
XXMUX90 bl[90] br[90] bl_out[45] br_out[45] sel[0] gnd single_level_column_mux_8
XXMUX91 bl[91] br[91] bl_out[45] br_out[45] sel[1] gnd single_level_column_mux_8
XXMUX92 bl[92] br[92] bl_out[46] br_out[46] sel[0] gnd single_level_column_mux_8
XXMUX93 bl[93] br[93] bl_out[46] br_out[46] sel[1] gnd single_level_column_mux_8
XXMUX94 bl[94] br[94] bl_out[47] br_out[47] sel[0] gnd single_level_column_mux_8
XXMUX95 bl[95] br[95] bl_out[47] br_out[47] sel[1] gnd single_level_column_mux_8
XXMUX96 bl[96] br[96] bl_out[48] br_out[48] sel[0] gnd single_level_column_mux_8
XXMUX97 bl[97] br[97] bl_out[48] br_out[48] sel[1] gnd single_level_column_mux_8
XXMUX98 bl[98] br[98] bl_out[49] br_out[49] sel[0] gnd single_level_column_mux_8
XXMUX99 bl[99] br[99] bl_out[49] br_out[49] sel[1] gnd single_level_column_mux_8
XXMUX100 bl[100] br[100] bl_out[50] br_out[50] sel[0] gnd single_level_column_mux_8
XXMUX101 bl[101] br[101] bl_out[50] br_out[50] sel[1] gnd single_level_column_mux_8
XXMUX102 bl[102] br[102] bl_out[51] br_out[51] sel[0] gnd single_level_column_mux_8
XXMUX103 bl[103] br[103] bl_out[51] br_out[51] sel[1] gnd single_level_column_mux_8
XXMUX104 bl[104] br[104] bl_out[52] br_out[52] sel[0] gnd single_level_column_mux_8
XXMUX105 bl[105] br[105] bl_out[52] br_out[52] sel[1] gnd single_level_column_mux_8
XXMUX106 bl[106] br[106] bl_out[53] br_out[53] sel[0] gnd single_level_column_mux_8
XXMUX107 bl[107] br[107] bl_out[53] br_out[53] sel[1] gnd single_level_column_mux_8
XXMUX108 bl[108] br[108] bl_out[54] br_out[54] sel[0] gnd single_level_column_mux_8
XXMUX109 bl[109] br[109] bl_out[54] br_out[54] sel[1] gnd single_level_column_mux_8
XXMUX110 bl[110] br[110] bl_out[55] br_out[55] sel[0] gnd single_level_column_mux_8
XXMUX111 bl[111] br[111] bl_out[55] br_out[55] sel[1] gnd single_level_column_mux_8
XXMUX112 bl[112] br[112] bl_out[56] br_out[56] sel[0] gnd single_level_column_mux_8
XXMUX113 bl[113] br[113] bl_out[56] br_out[56] sel[1] gnd single_level_column_mux_8
XXMUX114 bl[114] br[114] bl_out[57] br_out[57] sel[0] gnd single_level_column_mux_8
XXMUX115 bl[115] br[115] bl_out[57] br_out[57] sel[1] gnd single_level_column_mux_8
XXMUX116 bl[116] br[116] bl_out[58] br_out[58] sel[0] gnd single_level_column_mux_8
XXMUX117 bl[117] br[117] bl_out[58] br_out[58] sel[1] gnd single_level_column_mux_8
XXMUX118 bl[118] br[118] bl_out[59] br_out[59] sel[0] gnd single_level_column_mux_8
XXMUX119 bl[119] br[119] bl_out[59] br_out[59] sel[1] gnd single_level_column_mux_8
XXMUX120 bl[120] br[120] bl_out[60] br_out[60] sel[0] gnd single_level_column_mux_8
XXMUX121 bl[121] br[121] bl_out[60] br_out[60] sel[1] gnd single_level_column_mux_8
XXMUX122 bl[122] br[122] bl_out[61] br_out[61] sel[0] gnd single_level_column_mux_8
XXMUX123 bl[123] br[123] bl_out[61] br_out[61] sel[1] gnd single_level_column_mux_8
XXMUX124 bl[124] br[124] bl_out[62] br_out[62] sel[0] gnd single_level_column_mux_8
XXMUX125 bl[125] br[125] bl_out[62] br_out[62] sel[1] gnd single_level_column_mux_8
XXMUX126 bl[126] br[126] bl_out[63] br_out[63] sel[0] gnd single_level_column_mux_8
XXMUX127 bl[127] br[127] bl_out[63] br_out[63] sel[1] gnd single_level_column_mux_8
XXMUX128 bl[128] br[128] bl_out[64] br_out[64] sel[0] gnd single_level_column_mux_8
XXMUX129 bl[129] br[129] bl_out[64] br_out[64] sel[1] gnd single_level_column_mux_8
XXMUX130 bl[130] br[130] bl_out[65] br_out[65] sel[0] gnd single_level_column_mux_8
XXMUX131 bl[131] br[131] bl_out[65] br_out[65] sel[1] gnd single_level_column_mux_8
XXMUX132 bl[132] br[132] bl_out[66] br_out[66] sel[0] gnd single_level_column_mux_8
XXMUX133 bl[133] br[133] bl_out[66] br_out[66] sel[1] gnd single_level_column_mux_8
XXMUX134 bl[134] br[134] bl_out[67] br_out[67] sel[0] gnd single_level_column_mux_8
XXMUX135 bl[135] br[135] bl_out[67] br_out[67] sel[1] gnd single_level_column_mux_8
XXMUX136 bl[136] br[136] bl_out[68] br_out[68] sel[0] gnd single_level_column_mux_8
XXMUX137 bl[137] br[137] bl_out[68] br_out[68] sel[1] gnd single_level_column_mux_8
XXMUX138 bl[138] br[138] bl_out[69] br_out[69] sel[0] gnd single_level_column_mux_8
XXMUX139 bl[139] br[139] bl_out[69] br_out[69] sel[1] gnd single_level_column_mux_8
XXMUX140 bl[140] br[140] bl_out[70] br_out[70] sel[0] gnd single_level_column_mux_8
XXMUX141 bl[141] br[141] bl_out[70] br_out[70] sel[1] gnd single_level_column_mux_8
XXMUX142 bl[142] br[142] bl_out[71] br_out[71] sel[0] gnd single_level_column_mux_8
XXMUX143 bl[143] br[143] bl_out[71] br_out[71] sel[1] gnd single_level_column_mux_8
XXMUX144 bl[144] br[144] bl_out[72] br_out[72] sel[0] gnd single_level_column_mux_8
XXMUX145 bl[145] br[145] bl_out[72] br_out[72] sel[1] gnd single_level_column_mux_8
XXMUX146 bl[146] br[146] bl_out[73] br_out[73] sel[0] gnd single_level_column_mux_8
XXMUX147 bl[147] br[147] bl_out[73] br_out[73] sel[1] gnd single_level_column_mux_8
XXMUX148 bl[148] br[148] bl_out[74] br_out[74] sel[0] gnd single_level_column_mux_8
XXMUX149 bl[149] br[149] bl_out[74] br_out[74] sel[1] gnd single_level_column_mux_8
XXMUX150 bl[150] br[150] bl_out[75] br_out[75] sel[0] gnd single_level_column_mux_8
XXMUX151 bl[151] br[151] bl_out[75] br_out[75] sel[1] gnd single_level_column_mux_8
XXMUX152 bl[152] br[152] bl_out[76] br_out[76] sel[0] gnd single_level_column_mux_8
XXMUX153 bl[153] br[153] bl_out[76] br_out[76] sel[1] gnd single_level_column_mux_8
XXMUX154 bl[154] br[154] bl_out[77] br_out[77] sel[0] gnd single_level_column_mux_8
XXMUX155 bl[155] br[155] bl_out[77] br_out[77] sel[1] gnd single_level_column_mux_8
XXMUX156 bl[156] br[156] bl_out[78] br_out[78] sel[0] gnd single_level_column_mux_8
XXMUX157 bl[157] br[157] bl_out[78] br_out[78] sel[1] gnd single_level_column_mux_8
XXMUX158 bl[158] br[158] bl_out[79] br_out[79] sel[0] gnd single_level_column_mux_8
XXMUX159 bl[159] br[159] bl_out[79] br_out[79] sel[1] gnd single_level_column_mux_8
XXMUX160 bl[160] br[160] bl_out[80] br_out[80] sel[0] gnd single_level_column_mux_8
XXMUX161 bl[161] br[161] bl_out[80] br_out[80] sel[1] gnd single_level_column_mux_8
XXMUX162 bl[162] br[162] bl_out[81] br_out[81] sel[0] gnd single_level_column_mux_8
XXMUX163 bl[163] br[163] bl_out[81] br_out[81] sel[1] gnd single_level_column_mux_8
XXMUX164 bl[164] br[164] bl_out[82] br_out[82] sel[0] gnd single_level_column_mux_8
XXMUX165 bl[165] br[165] bl_out[82] br_out[82] sel[1] gnd single_level_column_mux_8
XXMUX166 bl[166] br[166] bl_out[83] br_out[83] sel[0] gnd single_level_column_mux_8
XXMUX167 bl[167] br[167] bl_out[83] br_out[83] sel[1] gnd single_level_column_mux_8
XXMUX168 bl[168] br[168] bl_out[84] br_out[84] sel[0] gnd single_level_column_mux_8
XXMUX169 bl[169] br[169] bl_out[84] br_out[84] sel[1] gnd single_level_column_mux_8
XXMUX170 bl[170] br[170] bl_out[85] br_out[85] sel[0] gnd single_level_column_mux_8
XXMUX171 bl[171] br[171] bl_out[85] br_out[85] sel[1] gnd single_level_column_mux_8
XXMUX172 bl[172] br[172] bl_out[86] br_out[86] sel[0] gnd single_level_column_mux_8
XXMUX173 bl[173] br[173] bl_out[86] br_out[86] sel[1] gnd single_level_column_mux_8
XXMUX174 bl[174] br[174] bl_out[87] br_out[87] sel[0] gnd single_level_column_mux_8
XXMUX175 bl[175] br[175] bl_out[87] br_out[87] sel[1] gnd single_level_column_mux_8
XXMUX176 bl[176] br[176] bl_out[88] br_out[88] sel[0] gnd single_level_column_mux_8
XXMUX177 bl[177] br[177] bl_out[88] br_out[88] sel[1] gnd single_level_column_mux_8
XXMUX178 bl[178] br[178] bl_out[89] br_out[89] sel[0] gnd single_level_column_mux_8
XXMUX179 bl[179] br[179] bl_out[89] br_out[89] sel[1] gnd single_level_column_mux_8
XXMUX180 bl[180] br[180] bl_out[90] br_out[90] sel[0] gnd single_level_column_mux_8
XXMUX181 bl[181] br[181] bl_out[90] br_out[90] sel[1] gnd single_level_column_mux_8
XXMUX182 bl[182] br[182] bl_out[91] br_out[91] sel[0] gnd single_level_column_mux_8
XXMUX183 bl[183] br[183] bl_out[91] br_out[91] sel[1] gnd single_level_column_mux_8
XXMUX184 bl[184] br[184] bl_out[92] br_out[92] sel[0] gnd single_level_column_mux_8
XXMUX185 bl[185] br[185] bl_out[92] br_out[92] sel[1] gnd single_level_column_mux_8
XXMUX186 bl[186] br[186] bl_out[93] br_out[93] sel[0] gnd single_level_column_mux_8
XXMUX187 bl[187] br[187] bl_out[93] br_out[93] sel[1] gnd single_level_column_mux_8
XXMUX188 bl[188] br[188] bl_out[94] br_out[94] sel[0] gnd single_level_column_mux_8
XXMUX189 bl[189] br[189] bl_out[94] br_out[94] sel[1] gnd single_level_column_mux_8
XXMUX190 bl[190] br[190] bl_out[95] br_out[95] sel[0] gnd single_level_column_mux_8
XXMUX191 bl[191] br[191] bl_out[95] br_out[95] sel[1] gnd single_level_column_mux_8
XXMUX192 bl[192] br[192] bl_out[96] br_out[96] sel[0] gnd single_level_column_mux_8
XXMUX193 bl[193] br[193] bl_out[96] br_out[96] sel[1] gnd single_level_column_mux_8
XXMUX194 bl[194] br[194] bl_out[97] br_out[97] sel[0] gnd single_level_column_mux_8
XXMUX195 bl[195] br[195] bl_out[97] br_out[97] sel[1] gnd single_level_column_mux_8
XXMUX196 bl[196] br[196] bl_out[98] br_out[98] sel[0] gnd single_level_column_mux_8
XXMUX197 bl[197] br[197] bl_out[98] br_out[98] sel[1] gnd single_level_column_mux_8
XXMUX198 bl[198] br[198] bl_out[99] br_out[99] sel[0] gnd single_level_column_mux_8
XXMUX199 bl[199] br[199] bl_out[99] br_out[99] sel[1] gnd single_level_column_mux_8
XXMUX200 bl[200] br[200] bl_out[100] br_out[100] sel[0] gnd single_level_column_mux_8
XXMUX201 bl[201] br[201] bl_out[100] br_out[100] sel[1] gnd single_level_column_mux_8
XXMUX202 bl[202] br[202] bl_out[101] br_out[101] sel[0] gnd single_level_column_mux_8
XXMUX203 bl[203] br[203] bl_out[101] br_out[101] sel[1] gnd single_level_column_mux_8
XXMUX204 bl[204] br[204] bl_out[102] br_out[102] sel[0] gnd single_level_column_mux_8
XXMUX205 bl[205] br[205] bl_out[102] br_out[102] sel[1] gnd single_level_column_mux_8
XXMUX206 bl[206] br[206] bl_out[103] br_out[103] sel[0] gnd single_level_column_mux_8
XXMUX207 bl[207] br[207] bl_out[103] br_out[103] sel[1] gnd single_level_column_mux_8
XXMUX208 bl[208] br[208] bl_out[104] br_out[104] sel[0] gnd single_level_column_mux_8
XXMUX209 bl[209] br[209] bl_out[104] br_out[104] sel[1] gnd single_level_column_mux_8
XXMUX210 bl[210] br[210] bl_out[105] br_out[105] sel[0] gnd single_level_column_mux_8
XXMUX211 bl[211] br[211] bl_out[105] br_out[105] sel[1] gnd single_level_column_mux_8
XXMUX212 bl[212] br[212] bl_out[106] br_out[106] sel[0] gnd single_level_column_mux_8
XXMUX213 bl[213] br[213] bl_out[106] br_out[106] sel[1] gnd single_level_column_mux_8
XXMUX214 bl[214] br[214] bl_out[107] br_out[107] sel[0] gnd single_level_column_mux_8
XXMUX215 bl[215] br[215] bl_out[107] br_out[107] sel[1] gnd single_level_column_mux_8
XXMUX216 bl[216] br[216] bl_out[108] br_out[108] sel[0] gnd single_level_column_mux_8
XXMUX217 bl[217] br[217] bl_out[108] br_out[108] sel[1] gnd single_level_column_mux_8
XXMUX218 bl[218] br[218] bl_out[109] br_out[109] sel[0] gnd single_level_column_mux_8
XXMUX219 bl[219] br[219] bl_out[109] br_out[109] sel[1] gnd single_level_column_mux_8
XXMUX220 bl[220] br[220] bl_out[110] br_out[110] sel[0] gnd single_level_column_mux_8
XXMUX221 bl[221] br[221] bl_out[110] br_out[110] sel[1] gnd single_level_column_mux_8
XXMUX222 bl[222] br[222] bl_out[111] br_out[111] sel[0] gnd single_level_column_mux_8
XXMUX223 bl[223] br[223] bl_out[111] br_out[111] sel[1] gnd single_level_column_mux_8
XXMUX224 bl[224] br[224] bl_out[112] br_out[112] sel[0] gnd single_level_column_mux_8
XXMUX225 bl[225] br[225] bl_out[112] br_out[112] sel[1] gnd single_level_column_mux_8
XXMUX226 bl[226] br[226] bl_out[113] br_out[113] sel[0] gnd single_level_column_mux_8
XXMUX227 bl[227] br[227] bl_out[113] br_out[113] sel[1] gnd single_level_column_mux_8
XXMUX228 bl[228] br[228] bl_out[114] br_out[114] sel[0] gnd single_level_column_mux_8
XXMUX229 bl[229] br[229] bl_out[114] br_out[114] sel[1] gnd single_level_column_mux_8
XXMUX230 bl[230] br[230] bl_out[115] br_out[115] sel[0] gnd single_level_column_mux_8
XXMUX231 bl[231] br[231] bl_out[115] br_out[115] sel[1] gnd single_level_column_mux_8
XXMUX232 bl[232] br[232] bl_out[116] br_out[116] sel[0] gnd single_level_column_mux_8
XXMUX233 bl[233] br[233] bl_out[116] br_out[116] sel[1] gnd single_level_column_mux_8
XXMUX234 bl[234] br[234] bl_out[117] br_out[117] sel[0] gnd single_level_column_mux_8
XXMUX235 bl[235] br[235] bl_out[117] br_out[117] sel[1] gnd single_level_column_mux_8
XXMUX236 bl[236] br[236] bl_out[118] br_out[118] sel[0] gnd single_level_column_mux_8
XXMUX237 bl[237] br[237] bl_out[118] br_out[118] sel[1] gnd single_level_column_mux_8
XXMUX238 bl[238] br[238] bl_out[119] br_out[119] sel[0] gnd single_level_column_mux_8
XXMUX239 bl[239] br[239] bl_out[119] br_out[119] sel[1] gnd single_level_column_mux_8
XXMUX240 bl[240] br[240] bl_out[120] br_out[120] sel[0] gnd single_level_column_mux_8
XXMUX241 bl[241] br[241] bl_out[120] br_out[120] sel[1] gnd single_level_column_mux_8
XXMUX242 bl[242] br[242] bl_out[121] br_out[121] sel[0] gnd single_level_column_mux_8
XXMUX243 bl[243] br[243] bl_out[121] br_out[121] sel[1] gnd single_level_column_mux_8
XXMUX244 bl[244] br[244] bl_out[122] br_out[122] sel[0] gnd single_level_column_mux_8
XXMUX245 bl[245] br[245] bl_out[122] br_out[122] sel[1] gnd single_level_column_mux_8
XXMUX246 bl[246] br[246] bl_out[123] br_out[123] sel[0] gnd single_level_column_mux_8
XXMUX247 bl[247] br[247] bl_out[123] br_out[123] sel[1] gnd single_level_column_mux_8
XXMUX248 bl[248] br[248] bl_out[124] br_out[124] sel[0] gnd single_level_column_mux_8
XXMUX249 bl[249] br[249] bl_out[124] br_out[124] sel[1] gnd single_level_column_mux_8
XXMUX250 bl[250] br[250] bl_out[125] br_out[125] sel[0] gnd single_level_column_mux_8
XXMUX251 bl[251] br[251] bl_out[125] br_out[125] sel[1] gnd single_level_column_mux_8
XXMUX252 bl[252] br[252] bl_out[126] br_out[126] sel[0] gnd single_level_column_mux_8
XXMUX253 bl[253] br[253] bl_out[126] br_out[126] sel[1] gnd single_level_column_mux_8
XXMUX254 bl[254] br[254] bl_out[127] br_out[127] sel[0] gnd single_level_column_mux_8
XXMUX255 bl[255] br[255] bl_out[127] br_out[127] sel[1] gnd single_level_column_mux_8
.ENDS columnmux_array
*********************** "sense_amp" ******************************

.SUBCKT sense_amp bl br dout en vdd gnd
M_1 dout net_1 vdd vdd p W='5.4*1u' L=0.6u
M_2 dout net_1 net_2 gnd n W='2.7*1u' L=0.6u
M_3 net_1 dout vdd vdd p W='5.4*1u' L=0.6u
M_4 net_1 dout net_2 gnd n W='2.7*1u' L=0.6u
M_5 bl en dout vdd p W='7.2*1u' L=0.6u
M_6 br en net_1 vdd p W='7.2*1u' L=0.6u
M_7 net_2 en gnd gnd n W='2.7*1u' L=0.6u
.ENDS	 sense_amp


.SUBCKT sense_amp_array data[0] bl[0] br[0] data[1] bl[2] br[2] data[2] bl[4] br[4] data[3] bl[6] br[6] data[4] bl[8] br[8] data[5] bl[10] br[10] data[6] bl[12] br[12] data[7] bl[14] br[14] data[8] bl[16] br[16] data[9] bl[18] br[18] data[10] bl[20] br[20] data[11] bl[22] br[22] data[12] bl[24] br[24] data[13] bl[26] br[26] data[14] bl[28] br[28] data[15] bl[30] br[30] data[16] bl[32] br[32] data[17] bl[34] br[34] data[18] bl[36] br[36] data[19] bl[38] br[38] data[20] bl[40] br[40] data[21] bl[42] br[42] data[22] bl[44] br[44] data[23] bl[46] br[46] data[24] bl[48] br[48] data[25] bl[50] br[50] data[26] bl[52] br[52] data[27] bl[54] br[54] data[28] bl[56] br[56] data[29] bl[58] br[58] data[30] bl[60] br[60] data[31] bl[62] br[62] data[32] bl[64] br[64] data[33] bl[66] br[66] data[34] bl[68] br[68] data[35] bl[70] br[70] data[36] bl[72] br[72] data[37] bl[74] br[74] data[38] bl[76] br[76] data[39] bl[78] br[78] data[40] bl[80] br[80] data[41] bl[82] br[82] data[42] bl[84] br[84] data[43] bl[86] br[86] data[44] bl[88] br[88] data[45] bl[90] br[90] data[46] bl[92] br[92] data[47] bl[94] br[94] data[48] bl[96] br[96] data[49] bl[98] br[98] data[50] bl[100] br[100] data[51] bl[102] br[102] data[52] bl[104] br[104] data[53] bl[106] br[106] data[54] bl[108] br[108] data[55] bl[110] br[110] data[56] bl[112] br[112] data[57] bl[114] br[114] data[58] bl[116] br[116] data[59] bl[118] br[118] data[60] bl[120] br[120] data[61] bl[122] br[122] data[62] bl[124] br[124] data[63] bl[126] br[126] data[64] bl[128] br[128] data[65] bl[130] br[130] data[66] bl[132] br[132] data[67] bl[134] br[134] data[68] bl[136] br[136] data[69] bl[138] br[138] data[70] bl[140] br[140] data[71] bl[142] br[142] data[72] bl[144] br[144] data[73] bl[146] br[146] data[74] bl[148] br[148] data[75] bl[150] br[150] data[76] bl[152] br[152] data[77] bl[154] br[154] data[78] bl[156] br[156] data[79] bl[158] br[158] data[80] bl[160] br[160] data[81] bl[162] br[162] data[82] bl[164] br[164] data[83] bl[166] br[166] data[84] bl[168] br[168] data[85] bl[170] br[170] data[86] bl[172] br[172] data[87] bl[174] br[174] data[88] bl[176] br[176] data[89] bl[178] br[178] data[90] bl[180] br[180] data[91] bl[182] br[182] data[92] bl[184] br[184] data[93] bl[186] br[186] data[94] bl[188] br[188] data[95] bl[190] br[190] data[96] bl[192] br[192] data[97] bl[194] br[194] data[98] bl[196] br[196] data[99] bl[198] br[198] data[100] bl[200] br[200] data[101] bl[202] br[202] data[102] bl[204] br[204] data[103] bl[206] br[206] data[104] bl[208] br[208] data[105] bl[210] br[210] data[106] bl[212] br[212] data[107] bl[214] br[214] data[108] bl[216] br[216] data[109] bl[218] br[218] data[110] bl[220] br[220] data[111] bl[222] br[222] data[112] bl[224] br[224] data[113] bl[226] br[226] data[114] bl[228] br[228] data[115] bl[230] br[230] data[116] bl[232] br[232] data[117] bl[234] br[234] data[118] bl[236] br[236] data[119] bl[238] br[238] data[120] bl[240] br[240] data[121] bl[242] br[242] data[122] bl[244] br[244] data[123] bl[246] br[246] data[124] bl[248] br[248] data[125] bl[250] br[250] data[126] bl[252] br[252] data[127] bl[254] br[254] en vdd gnd
Xsa_d0 bl[0] br[0] data[0] en vdd gnd sense_amp
Xsa_d2 bl[2] br[2] data[1] en vdd gnd sense_amp
Xsa_d4 bl[4] br[4] data[2] en vdd gnd sense_amp
Xsa_d6 bl[6] br[6] data[3] en vdd gnd sense_amp
Xsa_d8 bl[8] br[8] data[4] en vdd gnd sense_amp
Xsa_d10 bl[10] br[10] data[5] en vdd gnd sense_amp
Xsa_d12 bl[12] br[12] data[6] en vdd gnd sense_amp
Xsa_d14 bl[14] br[14] data[7] en vdd gnd sense_amp
Xsa_d16 bl[16] br[16] data[8] en vdd gnd sense_amp
Xsa_d18 bl[18] br[18] data[9] en vdd gnd sense_amp
Xsa_d20 bl[20] br[20] data[10] en vdd gnd sense_amp
Xsa_d22 bl[22] br[22] data[11] en vdd gnd sense_amp
Xsa_d24 bl[24] br[24] data[12] en vdd gnd sense_amp
Xsa_d26 bl[26] br[26] data[13] en vdd gnd sense_amp
Xsa_d28 bl[28] br[28] data[14] en vdd gnd sense_amp
Xsa_d30 bl[30] br[30] data[15] en vdd gnd sense_amp
Xsa_d32 bl[32] br[32] data[16] en vdd gnd sense_amp
Xsa_d34 bl[34] br[34] data[17] en vdd gnd sense_amp
Xsa_d36 bl[36] br[36] data[18] en vdd gnd sense_amp
Xsa_d38 bl[38] br[38] data[19] en vdd gnd sense_amp
Xsa_d40 bl[40] br[40] data[20] en vdd gnd sense_amp
Xsa_d42 bl[42] br[42] data[21] en vdd gnd sense_amp
Xsa_d44 bl[44] br[44] data[22] en vdd gnd sense_amp
Xsa_d46 bl[46] br[46] data[23] en vdd gnd sense_amp
Xsa_d48 bl[48] br[48] data[24] en vdd gnd sense_amp
Xsa_d50 bl[50] br[50] data[25] en vdd gnd sense_amp
Xsa_d52 bl[52] br[52] data[26] en vdd gnd sense_amp
Xsa_d54 bl[54] br[54] data[27] en vdd gnd sense_amp
Xsa_d56 bl[56] br[56] data[28] en vdd gnd sense_amp
Xsa_d58 bl[58] br[58] data[29] en vdd gnd sense_amp
Xsa_d60 bl[60] br[60] data[30] en vdd gnd sense_amp
Xsa_d62 bl[62] br[62] data[31] en vdd gnd sense_amp
Xsa_d64 bl[64] br[64] data[32] en vdd gnd sense_amp
Xsa_d66 bl[66] br[66] data[33] en vdd gnd sense_amp
Xsa_d68 bl[68] br[68] data[34] en vdd gnd sense_amp
Xsa_d70 bl[70] br[70] data[35] en vdd gnd sense_amp
Xsa_d72 bl[72] br[72] data[36] en vdd gnd sense_amp
Xsa_d74 bl[74] br[74] data[37] en vdd gnd sense_amp
Xsa_d76 bl[76] br[76] data[38] en vdd gnd sense_amp
Xsa_d78 bl[78] br[78] data[39] en vdd gnd sense_amp
Xsa_d80 bl[80] br[80] data[40] en vdd gnd sense_amp
Xsa_d82 bl[82] br[82] data[41] en vdd gnd sense_amp
Xsa_d84 bl[84] br[84] data[42] en vdd gnd sense_amp
Xsa_d86 bl[86] br[86] data[43] en vdd gnd sense_amp
Xsa_d88 bl[88] br[88] data[44] en vdd gnd sense_amp
Xsa_d90 bl[90] br[90] data[45] en vdd gnd sense_amp
Xsa_d92 bl[92] br[92] data[46] en vdd gnd sense_amp
Xsa_d94 bl[94] br[94] data[47] en vdd gnd sense_amp
Xsa_d96 bl[96] br[96] data[48] en vdd gnd sense_amp
Xsa_d98 bl[98] br[98] data[49] en vdd gnd sense_amp
Xsa_d100 bl[100] br[100] data[50] en vdd gnd sense_amp
Xsa_d102 bl[102] br[102] data[51] en vdd gnd sense_amp
Xsa_d104 bl[104] br[104] data[52] en vdd gnd sense_amp
Xsa_d106 bl[106] br[106] data[53] en vdd gnd sense_amp
Xsa_d108 bl[108] br[108] data[54] en vdd gnd sense_amp
Xsa_d110 bl[110] br[110] data[55] en vdd gnd sense_amp
Xsa_d112 bl[112] br[112] data[56] en vdd gnd sense_amp
Xsa_d114 bl[114] br[114] data[57] en vdd gnd sense_amp
Xsa_d116 bl[116] br[116] data[58] en vdd gnd sense_amp
Xsa_d118 bl[118] br[118] data[59] en vdd gnd sense_amp
Xsa_d120 bl[120] br[120] data[60] en vdd gnd sense_amp
Xsa_d122 bl[122] br[122] data[61] en vdd gnd sense_amp
Xsa_d124 bl[124] br[124] data[62] en vdd gnd sense_amp
Xsa_d126 bl[126] br[126] data[63] en vdd gnd sense_amp
Xsa_d128 bl[128] br[128] data[64] en vdd gnd sense_amp
Xsa_d130 bl[130] br[130] data[65] en vdd gnd sense_amp
Xsa_d132 bl[132] br[132] data[66] en vdd gnd sense_amp
Xsa_d134 bl[134] br[134] data[67] en vdd gnd sense_amp
Xsa_d136 bl[136] br[136] data[68] en vdd gnd sense_amp
Xsa_d138 bl[138] br[138] data[69] en vdd gnd sense_amp
Xsa_d140 bl[140] br[140] data[70] en vdd gnd sense_amp
Xsa_d142 bl[142] br[142] data[71] en vdd gnd sense_amp
Xsa_d144 bl[144] br[144] data[72] en vdd gnd sense_amp
Xsa_d146 bl[146] br[146] data[73] en vdd gnd sense_amp
Xsa_d148 bl[148] br[148] data[74] en vdd gnd sense_amp
Xsa_d150 bl[150] br[150] data[75] en vdd gnd sense_amp
Xsa_d152 bl[152] br[152] data[76] en vdd gnd sense_amp
Xsa_d154 bl[154] br[154] data[77] en vdd gnd sense_amp
Xsa_d156 bl[156] br[156] data[78] en vdd gnd sense_amp
Xsa_d158 bl[158] br[158] data[79] en vdd gnd sense_amp
Xsa_d160 bl[160] br[160] data[80] en vdd gnd sense_amp
Xsa_d162 bl[162] br[162] data[81] en vdd gnd sense_amp
Xsa_d164 bl[164] br[164] data[82] en vdd gnd sense_amp
Xsa_d166 bl[166] br[166] data[83] en vdd gnd sense_amp
Xsa_d168 bl[168] br[168] data[84] en vdd gnd sense_amp
Xsa_d170 bl[170] br[170] data[85] en vdd gnd sense_amp
Xsa_d172 bl[172] br[172] data[86] en vdd gnd sense_amp
Xsa_d174 bl[174] br[174] data[87] en vdd gnd sense_amp
Xsa_d176 bl[176] br[176] data[88] en vdd gnd sense_amp
Xsa_d178 bl[178] br[178] data[89] en vdd gnd sense_amp
Xsa_d180 bl[180] br[180] data[90] en vdd gnd sense_amp
Xsa_d182 bl[182] br[182] data[91] en vdd gnd sense_amp
Xsa_d184 bl[184] br[184] data[92] en vdd gnd sense_amp
Xsa_d186 bl[186] br[186] data[93] en vdd gnd sense_amp
Xsa_d188 bl[188] br[188] data[94] en vdd gnd sense_amp
Xsa_d190 bl[190] br[190] data[95] en vdd gnd sense_amp
Xsa_d192 bl[192] br[192] data[96] en vdd gnd sense_amp
Xsa_d194 bl[194] br[194] data[97] en vdd gnd sense_amp
Xsa_d196 bl[196] br[196] data[98] en vdd gnd sense_amp
Xsa_d198 bl[198] br[198] data[99] en vdd gnd sense_amp
Xsa_d200 bl[200] br[200] data[100] en vdd gnd sense_amp
Xsa_d202 bl[202] br[202] data[101] en vdd gnd sense_amp
Xsa_d204 bl[204] br[204] data[102] en vdd gnd sense_amp
Xsa_d206 bl[206] br[206] data[103] en vdd gnd sense_amp
Xsa_d208 bl[208] br[208] data[104] en vdd gnd sense_amp
Xsa_d210 bl[210] br[210] data[105] en vdd gnd sense_amp
Xsa_d212 bl[212] br[212] data[106] en vdd gnd sense_amp
Xsa_d214 bl[214] br[214] data[107] en vdd gnd sense_amp
Xsa_d216 bl[216] br[216] data[108] en vdd gnd sense_amp
Xsa_d218 bl[218] br[218] data[109] en vdd gnd sense_amp
Xsa_d220 bl[220] br[220] data[110] en vdd gnd sense_amp
Xsa_d222 bl[222] br[222] data[111] en vdd gnd sense_amp
Xsa_d224 bl[224] br[224] data[112] en vdd gnd sense_amp
Xsa_d226 bl[226] br[226] data[113] en vdd gnd sense_amp
Xsa_d228 bl[228] br[228] data[114] en vdd gnd sense_amp
Xsa_d230 bl[230] br[230] data[115] en vdd gnd sense_amp
Xsa_d232 bl[232] br[232] data[116] en vdd gnd sense_amp
Xsa_d234 bl[234] br[234] data[117] en vdd gnd sense_amp
Xsa_d236 bl[236] br[236] data[118] en vdd gnd sense_amp
Xsa_d238 bl[238] br[238] data[119] en vdd gnd sense_amp
Xsa_d240 bl[240] br[240] data[120] en vdd gnd sense_amp
Xsa_d242 bl[242] br[242] data[121] en vdd gnd sense_amp
Xsa_d244 bl[244] br[244] data[122] en vdd gnd sense_amp
Xsa_d246 bl[246] br[246] data[123] en vdd gnd sense_amp
Xsa_d248 bl[248] br[248] data[124] en vdd gnd sense_amp
Xsa_d250 bl[250] br[250] data[125] en vdd gnd sense_amp
Xsa_d252 bl[252] br[252] data[126] en vdd gnd sense_amp
Xsa_d254 bl[254] br[254] data[127] en vdd gnd sense_amp
.ENDS sense_amp_array
*********************** Write_Driver ******************************
.SUBCKT write_driver din bl br en vdd gnd

**** Inverter to conver Data_in to data_in_bar ******
M_1 net_3 din gnd gnd n W='1.2*1u' L=0.6u
M_2 net_3 din vdd vdd p W='2.1*1u' L=0.6u

**** 2input nand gate follwed by inverter to drive BL ******
M_3 net_2 en net_7 gnd n W='2.1*1u' L=0.6u
M_4 net_7 din gnd gnd n W='2.1*1u' L=0.6u
M_5 net_2 en vdd vdd p W='2.1*1u' L=0.6u
M_6 net_2 din vdd vdd p W='2.1*1u' L=0.6u


M_7 net_1 net_2 vdd vdd p W='2.1*1u' L=0.6u
M_8 net_1 net_2 gnd gnd n W='1.2*1u' L=0.6u

**** 2input nand gate follwed by inverter to drive BR******

M_9 net_4 en vdd vdd p W='2.1*1u' L=0.6u
M_10 net_4 en net_8 gnd n W='2.1*1u' L=0.6u
M_11 net_8 net_3 gnd gnd n W='2.1*1u' L=0.6u
M_12 net_4 net_3 vdd vdd p W='2.1*1u' L=0.6u

M_13 net_6 net_4 vdd vdd p W='2.1*1u' L=0.6u
M_14 net_6 net_4 gnd gnd n W='1.2*1u' L=0.6u

************************************************

M_15 bl net_6 net_5 gnd n W='3.6*1u' L=0.6u
M_16 br net_1 net_5 gnd n W='3.6*1u' L=0.6u
M_17 net_5 en gnd gnd n W='3.6*1u' L=0.6u



.ENDS	$ write_driver


.SUBCKT write_driver_array data[0] data[1] data[2] data[3] data[4] data[5] data[6] data[7] data[8] data[9] data[10] data[11] data[12] data[13] data[14] data[15] data[16] data[17] data[18] data[19] data[20] data[21] data[22] data[23] data[24] data[25] data[26] data[27] data[28] data[29] data[30] data[31] data[32] data[33] data[34] data[35] data[36] data[37] data[38] data[39] data[40] data[41] data[42] data[43] data[44] data[45] data[46] data[47] data[48] data[49] data[50] data[51] data[52] data[53] data[54] data[55] data[56] data[57] data[58] data[59] data[60] data[61] data[62] data[63] data[64] data[65] data[66] data[67] data[68] data[69] data[70] data[71] data[72] data[73] data[74] data[75] data[76] data[77] data[78] data[79] data[80] data[81] data[82] data[83] data[84] data[85] data[86] data[87] data[88] data[89] data[90] data[91] data[92] data[93] data[94] data[95] data[96] data[97] data[98] data[99] data[100] data[101] data[102] data[103] data[104] data[105] data[106] data[107] data[108] data[109] data[110] data[111] data[112] data[113] data[114] data[115] data[116] data[117] data[118] data[119] data[120] data[121] data[122] data[123] data[124] data[125] data[126] data[127] bl[0] br[0] bl[1] br[1] bl[2] br[2] bl[3] br[3] bl[4] br[4] bl[5] br[5] bl[6] br[6] bl[7] br[7] bl[8] br[8] bl[9] br[9] bl[10] br[10] bl[11] br[11] bl[12] br[12] bl[13] br[13] bl[14] br[14] bl[15] br[15] bl[16] br[16] bl[17] br[17] bl[18] br[18] bl[19] br[19] bl[20] br[20] bl[21] br[21] bl[22] br[22] bl[23] br[23] bl[24] br[24] bl[25] br[25] bl[26] br[26] bl[27] br[27] bl[28] br[28] bl[29] br[29] bl[30] br[30] bl[31] br[31] bl[32] br[32] bl[33] br[33] bl[34] br[34] bl[35] br[35] bl[36] br[36] bl[37] br[37] bl[38] br[38] bl[39] br[39] bl[40] br[40] bl[41] br[41] bl[42] br[42] bl[43] br[43] bl[44] br[44] bl[45] br[45] bl[46] br[46] bl[47] br[47] bl[48] br[48] bl[49] br[49] bl[50] br[50] bl[51] br[51] bl[52] br[52] bl[53] br[53] bl[54] br[54] bl[55] br[55] bl[56] br[56] bl[57] br[57] bl[58] br[58] bl[59] br[59] bl[60] br[60] bl[61] br[61] bl[62] br[62] bl[63] br[63] bl[64] br[64] bl[65] br[65] bl[66] br[66] bl[67] br[67] bl[68] br[68] bl[69] br[69] bl[70] br[70] bl[71] br[71] bl[72] br[72] bl[73] br[73] bl[74] br[74] bl[75] br[75] bl[76] br[76] bl[77] br[77] bl[78] br[78] bl[79] br[79] bl[80] br[80] bl[81] br[81] bl[82] br[82] bl[83] br[83] bl[84] br[84] bl[85] br[85] bl[86] br[86] bl[87] br[87] bl[88] br[88] bl[89] br[89] bl[90] br[90] bl[91] br[91] bl[92] br[92] bl[93] br[93] bl[94] br[94] bl[95] br[95] bl[96] br[96] bl[97] br[97] bl[98] br[98] bl[99] br[99] bl[100] br[100] bl[101] br[101] bl[102] br[102] bl[103] br[103] bl[104] br[104] bl[105] br[105] bl[106] br[106] bl[107] br[107] bl[108] br[108] bl[109] br[109] bl[110] br[110] bl[111] br[111] bl[112] br[112] bl[113] br[113] bl[114] br[114] bl[115] br[115] bl[116] br[116] bl[117] br[117] bl[118] br[118] bl[119] br[119] bl[120] br[120] bl[121] br[121] bl[122] br[122] bl[123] br[123] bl[124] br[124] bl[125] br[125] bl[126] br[126] bl[127] br[127] en vdd gnd
XXwrite_driver0 data[0] bl[0] br[0] en vdd gnd write_driver
XXwrite_driver2 data[1] bl[1] br[1] en vdd gnd write_driver
XXwrite_driver4 data[2] bl[2] br[2] en vdd gnd write_driver
XXwrite_driver6 data[3] bl[3] br[3] en vdd gnd write_driver
XXwrite_driver8 data[4] bl[4] br[4] en vdd gnd write_driver
XXwrite_driver10 data[5] bl[5] br[5] en vdd gnd write_driver
XXwrite_driver12 data[6] bl[6] br[6] en vdd gnd write_driver
XXwrite_driver14 data[7] bl[7] br[7] en vdd gnd write_driver
XXwrite_driver16 data[8] bl[8] br[8] en vdd gnd write_driver
XXwrite_driver18 data[9] bl[9] br[9] en vdd gnd write_driver
XXwrite_driver20 data[10] bl[10] br[10] en vdd gnd write_driver
XXwrite_driver22 data[11] bl[11] br[11] en vdd gnd write_driver
XXwrite_driver24 data[12] bl[12] br[12] en vdd gnd write_driver
XXwrite_driver26 data[13] bl[13] br[13] en vdd gnd write_driver
XXwrite_driver28 data[14] bl[14] br[14] en vdd gnd write_driver
XXwrite_driver30 data[15] bl[15] br[15] en vdd gnd write_driver
XXwrite_driver32 data[16] bl[16] br[16] en vdd gnd write_driver
XXwrite_driver34 data[17] bl[17] br[17] en vdd gnd write_driver
XXwrite_driver36 data[18] bl[18] br[18] en vdd gnd write_driver
XXwrite_driver38 data[19] bl[19] br[19] en vdd gnd write_driver
XXwrite_driver40 data[20] bl[20] br[20] en vdd gnd write_driver
XXwrite_driver42 data[21] bl[21] br[21] en vdd gnd write_driver
XXwrite_driver44 data[22] bl[22] br[22] en vdd gnd write_driver
XXwrite_driver46 data[23] bl[23] br[23] en vdd gnd write_driver
XXwrite_driver48 data[24] bl[24] br[24] en vdd gnd write_driver
XXwrite_driver50 data[25] bl[25] br[25] en vdd gnd write_driver
XXwrite_driver52 data[26] bl[26] br[26] en vdd gnd write_driver
XXwrite_driver54 data[27] bl[27] br[27] en vdd gnd write_driver
XXwrite_driver56 data[28] bl[28] br[28] en vdd gnd write_driver
XXwrite_driver58 data[29] bl[29] br[29] en vdd gnd write_driver
XXwrite_driver60 data[30] bl[30] br[30] en vdd gnd write_driver
XXwrite_driver62 data[31] bl[31] br[31] en vdd gnd write_driver
XXwrite_driver64 data[32] bl[32] br[32] en vdd gnd write_driver
XXwrite_driver66 data[33] bl[33] br[33] en vdd gnd write_driver
XXwrite_driver68 data[34] bl[34] br[34] en vdd gnd write_driver
XXwrite_driver70 data[35] bl[35] br[35] en vdd gnd write_driver
XXwrite_driver72 data[36] bl[36] br[36] en vdd gnd write_driver
XXwrite_driver74 data[37] bl[37] br[37] en vdd gnd write_driver
XXwrite_driver76 data[38] bl[38] br[38] en vdd gnd write_driver
XXwrite_driver78 data[39] bl[39] br[39] en vdd gnd write_driver
XXwrite_driver80 data[40] bl[40] br[40] en vdd gnd write_driver
XXwrite_driver82 data[41] bl[41] br[41] en vdd gnd write_driver
XXwrite_driver84 data[42] bl[42] br[42] en vdd gnd write_driver
XXwrite_driver86 data[43] bl[43] br[43] en vdd gnd write_driver
XXwrite_driver88 data[44] bl[44] br[44] en vdd gnd write_driver
XXwrite_driver90 data[45] bl[45] br[45] en vdd gnd write_driver
XXwrite_driver92 data[46] bl[46] br[46] en vdd gnd write_driver
XXwrite_driver94 data[47] bl[47] br[47] en vdd gnd write_driver
XXwrite_driver96 data[48] bl[48] br[48] en vdd gnd write_driver
XXwrite_driver98 data[49] bl[49] br[49] en vdd gnd write_driver
XXwrite_driver100 data[50] bl[50] br[50] en vdd gnd write_driver
XXwrite_driver102 data[51] bl[51] br[51] en vdd gnd write_driver
XXwrite_driver104 data[52] bl[52] br[52] en vdd gnd write_driver
XXwrite_driver106 data[53] bl[53] br[53] en vdd gnd write_driver
XXwrite_driver108 data[54] bl[54] br[54] en vdd gnd write_driver
XXwrite_driver110 data[55] bl[55] br[55] en vdd gnd write_driver
XXwrite_driver112 data[56] bl[56] br[56] en vdd gnd write_driver
XXwrite_driver114 data[57] bl[57] br[57] en vdd gnd write_driver
XXwrite_driver116 data[58] bl[58] br[58] en vdd gnd write_driver
XXwrite_driver118 data[59] bl[59] br[59] en vdd gnd write_driver
XXwrite_driver120 data[60] bl[60] br[60] en vdd gnd write_driver
XXwrite_driver122 data[61] bl[61] br[61] en vdd gnd write_driver
XXwrite_driver124 data[62] bl[62] br[62] en vdd gnd write_driver
XXwrite_driver126 data[63] bl[63] br[63] en vdd gnd write_driver
XXwrite_driver128 data[64] bl[64] br[64] en vdd gnd write_driver
XXwrite_driver130 data[65] bl[65] br[65] en vdd gnd write_driver
XXwrite_driver132 data[66] bl[66] br[66] en vdd gnd write_driver
XXwrite_driver134 data[67] bl[67] br[67] en vdd gnd write_driver
XXwrite_driver136 data[68] bl[68] br[68] en vdd gnd write_driver
XXwrite_driver138 data[69] bl[69] br[69] en vdd gnd write_driver
XXwrite_driver140 data[70] bl[70] br[70] en vdd gnd write_driver
XXwrite_driver142 data[71] bl[71] br[71] en vdd gnd write_driver
XXwrite_driver144 data[72] bl[72] br[72] en vdd gnd write_driver
XXwrite_driver146 data[73] bl[73] br[73] en vdd gnd write_driver
XXwrite_driver148 data[74] bl[74] br[74] en vdd gnd write_driver
XXwrite_driver150 data[75] bl[75] br[75] en vdd gnd write_driver
XXwrite_driver152 data[76] bl[76] br[76] en vdd gnd write_driver
XXwrite_driver154 data[77] bl[77] br[77] en vdd gnd write_driver
XXwrite_driver156 data[78] bl[78] br[78] en vdd gnd write_driver
XXwrite_driver158 data[79] bl[79] br[79] en vdd gnd write_driver
XXwrite_driver160 data[80] bl[80] br[80] en vdd gnd write_driver
XXwrite_driver162 data[81] bl[81] br[81] en vdd gnd write_driver
XXwrite_driver164 data[82] bl[82] br[82] en vdd gnd write_driver
XXwrite_driver166 data[83] bl[83] br[83] en vdd gnd write_driver
XXwrite_driver168 data[84] bl[84] br[84] en vdd gnd write_driver
XXwrite_driver170 data[85] bl[85] br[85] en vdd gnd write_driver
XXwrite_driver172 data[86] bl[86] br[86] en vdd gnd write_driver
XXwrite_driver174 data[87] bl[87] br[87] en vdd gnd write_driver
XXwrite_driver176 data[88] bl[88] br[88] en vdd gnd write_driver
XXwrite_driver178 data[89] bl[89] br[89] en vdd gnd write_driver
XXwrite_driver180 data[90] bl[90] br[90] en vdd gnd write_driver
XXwrite_driver182 data[91] bl[91] br[91] en vdd gnd write_driver
XXwrite_driver184 data[92] bl[92] br[92] en vdd gnd write_driver
XXwrite_driver186 data[93] bl[93] br[93] en vdd gnd write_driver
XXwrite_driver188 data[94] bl[94] br[94] en vdd gnd write_driver
XXwrite_driver190 data[95] bl[95] br[95] en vdd gnd write_driver
XXwrite_driver192 data[96] bl[96] br[96] en vdd gnd write_driver
XXwrite_driver194 data[97] bl[97] br[97] en vdd gnd write_driver
XXwrite_driver196 data[98] bl[98] br[98] en vdd gnd write_driver
XXwrite_driver198 data[99] bl[99] br[99] en vdd gnd write_driver
XXwrite_driver200 data[100] bl[100] br[100] en vdd gnd write_driver
XXwrite_driver202 data[101] bl[101] br[101] en vdd gnd write_driver
XXwrite_driver204 data[102] bl[102] br[102] en vdd gnd write_driver
XXwrite_driver206 data[103] bl[103] br[103] en vdd gnd write_driver
XXwrite_driver208 data[104] bl[104] br[104] en vdd gnd write_driver
XXwrite_driver210 data[105] bl[105] br[105] en vdd gnd write_driver
XXwrite_driver212 data[106] bl[106] br[106] en vdd gnd write_driver
XXwrite_driver214 data[107] bl[107] br[107] en vdd gnd write_driver
XXwrite_driver216 data[108] bl[108] br[108] en vdd gnd write_driver
XXwrite_driver218 data[109] bl[109] br[109] en vdd gnd write_driver
XXwrite_driver220 data[110] bl[110] br[110] en vdd gnd write_driver
XXwrite_driver222 data[111] bl[111] br[111] en vdd gnd write_driver
XXwrite_driver224 data[112] bl[112] br[112] en vdd gnd write_driver
XXwrite_driver226 data[113] bl[113] br[113] en vdd gnd write_driver
XXwrite_driver228 data[114] bl[114] br[114] en vdd gnd write_driver
XXwrite_driver230 data[115] bl[115] br[115] en vdd gnd write_driver
XXwrite_driver232 data[116] bl[116] br[116] en vdd gnd write_driver
XXwrite_driver234 data[117] bl[117] br[117] en vdd gnd write_driver
XXwrite_driver236 data[118] bl[118] br[118] en vdd gnd write_driver
XXwrite_driver238 data[119] bl[119] br[119] en vdd gnd write_driver
XXwrite_driver240 data[120] bl[120] br[120] en vdd gnd write_driver
XXwrite_driver242 data[121] bl[121] br[121] en vdd gnd write_driver
XXwrite_driver244 data[122] bl[122] br[122] en vdd gnd write_driver
XXwrite_driver246 data[123] bl[123] br[123] en vdd gnd write_driver
XXwrite_driver248 data[124] bl[124] br[124] en vdd gnd write_driver
XXwrite_driver250 data[125] bl[125] br[125] en vdd gnd write_driver
XXwrite_driver252 data[126] bl[126] br[126] en vdd gnd write_driver
XXwrite_driver254 data[127] bl[127] br[127] en vdd gnd write_driver
.ENDS write_driver_array

.SUBCKT pinv_8 A Z vdd gnd
Mpinv_pmos Z A vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpinv_nmos Z A gnd gnd n m=1 w=1.2u l=0.6u pd=3.6u ps=3.6u as=1.8p ad=1.8p
.ENDS pinv_8

.SUBCKT pnand2_2 A B Z vdd gnd
Mpnand2_pmos1 vdd A Z vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand2_pmos2 Z B vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand2_nmos1 Z B net1 gnd n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand2_nmos2 net1 A gnd gnd n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
.ENDS pnand2_2

.SUBCKT pnand3_2 A B C Z vdd gnd
Mpnand3_pmos1 vdd A Z vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand3_pmos2 Z B vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand3_pmos3 Z C vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand3_nmos1 Z C net1 gnd n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand3_nmos2 net1 B net2 gnd n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand3_nmos3 net2 A gnd gnd n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
.ENDS pnand3_2

.SUBCKT pinv_9 A Z vdd gnd
Mpinv_pmos Z A vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpinv_nmos Z A gnd gnd n m=1 w=1.2u l=0.6u pd=3.6u ps=3.6u as=1.8p ad=1.8p
.ENDS pinv_9

.SUBCKT pnand2_3 A B Z vdd gnd
Mpnand2_pmos1 vdd A Z vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand2_pmos2 Z B vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand2_nmos1 Z B net1 gnd n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand2_nmos2 net1 A gnd gnd n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
.ENDS pnand2_3

.SUBCKT pre2x4 in[0] in[1] out[0] out[1] out[2] out[3] vdd gnd
XXpre_inv[0] in[0] inbar[0] vdd gnd pinv_9
XXpre_inv[1] in[1] inbar[1] vdd gnd pinv_9
XXpre_nand_inv[0] Z[0] out[0] vdd gnd pinv_9
XXpre_nand_inv[1] Z[1] out[1] vdd gnd pinv_9
XXpre_nand_inv[2] Z[2] out[2] vdd gnd pinv_9
XXpre_nand_inv[3] Z[3] out[3] vdd gnd pinv_9
XXpre2x4_nand[0] inbar[0] inbar[1] Z[0] vdd gnd pnand2_3
XXpre2x4_nand[1] in[0] inbar[1] Z[1] vdd gnd pnand2_3
XXpre2x4_nand[2] inbar[0] in[1] Z[2] vdd gnd pnand2_3
XXpre2x4_nand[3] in[0] in[1] Z[3] vdd gnd pnand2_3
.ENDS pre2x4

.SUBCKT pinv_10 A Z vdd gnd
Mpinv_pmos Z A vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpinv_nmos Z A gnd gnd n m=1 w=1.2u l=0.6u pd=3.6u ps=3.6u as=1.8p ad=1.8p
.ENDS pinv_10

.SUBCKT pnand3_3 A B C Z vdd gnd
Mpnand3_pmos1 vdd A Z vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand3_pmos2 Z B vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand3_pmos3 Z C vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand3_nmos1 Z C net1 gnd n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand3_nmos2 net1 B net2 gnd n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand3_nmos3 net2 A gnd gnd n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
.ENDS pnand3_3

.SUBCKT pre3x8 in[0] in[1] in[2] out[0] out[1] out[2] out[3] out[4] out[5] out[6] out[7] vdd gnd
XXpre_inv[0] in[0] inbar[0] vdd gnd pinv_10
XXpre_inv[1] in[1] inbar[1] vdd gnd pinv_10
XXpre_inv[2] in[2] inbar[2] vdd gnd pinv_10
XXpre_nand_inv[0] Z[0] out[0] vdd gnd pinv_10
XXpre_nand_inv[1] Z[1] out[1] vdd gnd pinv_10
XXpre_nand_inv[2] Z[2] out[2] vdd gnd pinv_10
XXpre_nand_inv[3] Z[3] out[3] vdd gnd pinv_10
XXpre_nand_inv[4] Z[4] out[4] vdd gnd pinv_10
XXpre_nand_inv[5] Z[5] out[5] vdd gnd pinv_10
XXpre_nand_inv[6] Z[6] out[6] vdd gnd pinv_10
XXpre_nand_inv[7] Z[7] out[7] vdd gnd pinv_10
XXpre3x8_nand[0] inbar[0] inbar[1] inbar[2] Z[0] vdd gnd pnand3_3
XXpre3x8_nand[1] in[0] inbar[1] inbar[2] Z[1] vdd gnd pnand3_3
XXpre3x8_nand[2] inbar[0] in[1] inbar[2] Z[2] vdd gnd pnand3_3
XXpre3x8_nand[3] in[0] in[1] inbar[2] Z[3] vdd gnd pnand3_3
XXpre3x8_nand[4] inbar[0] inbar[1] in[2] Z[4] vdd gnd pnand3_3
XXpre3x8_nand[5] in[0] inbar[1] in[2] Z[5] vdd gnd pnand3_3
XXpre3x8_nand[6] inbar[0] in[1] in[2] Z[6] vdd gnd pnand3_3
XXpre3x8_nand[7] in[0] in[1] in[2] Z[7] vdd gnd pnand3_3
.ENDS pre3x8

.SUBCKT hierarchical_decoder_256rows A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7] decode[0] decode[1] decode[2] decode[3] decode[4] decode[5] decode[6] decode[7] decode[8] decode[9] decode[10] decode[11] decode[12] decode[13] decode[14] decode[15] decode[16] decode[17] decode[18] decode[19] decode[20] decode[21] decode[22] decode[23] decode[24] decode[25] decode[26] decode[27] decode[28] decode[29] decode[30] decode[31] decode[32] decode[33] decode[34] decode[35] decode[36] decode[37] decode[38] decode[39] decode[40] decode[41] decode[42] decode[43] decode[44] decode[45] decode[46] decode[47] decode[48] decode[49] decode[50] decode[51] decode[52] decode[53] decode[54] decode[55] decode[56] decode[57] decode[58] decode[59] decode[60] decode[61] decode[62] decode[63] decode[64] decode[65] decode[66] decode[67] decode[68] decode[69] decode[70] decode[71] decode[72] decode[73] decode[74] decode[75] decode[76] decode[77] decode[78] decode[79] decode[80] decode[81] decode[82] decode[83] decode[84] decode[85] decode[86] decode[87] decode[88] decode[89] decode[90] decode[91] decode[92] decode[93] decode[94] decode[95] decode[96] decode[97] decode[98] decode[99] decode[100] decode[101] decode[102] decode[103] decode[104] decode[105] decode[106] decode[107] decode[108] decode[109] decode[110] decode[111] decode[112] decode[113] decode[114] decode[115] decode[116] decode[117] decode[118] decode[119] decode[120] decode[121] decode[122] decode[123] decode[124] decode[125] decode[126] decode[127] decode[128] decode[129] decode[130] decode[131] decode[132] decode[133] decode[134] decode[135] decode[136] decode[137] decode[138] decode[139] decode[140] decode[141] decode[142] decode[143] decode[144] decode[145] decode[146] decode[147] decode[148] decode[149] decode[150] decode[151] decode[152] decode[153] decode[154] decode[155] decode[156] decode[157] decode[158] decode[159] decode[160] decode[161] decode[162] decode[163] decode[164] decode[165] decode[166] decode[167] decode[168] decode[169] decode[170] decode[171] decode[172] decode[173] decode[174] decode[175] decode[176] decode[177] decode[178] decode[179] decode[180] decode[181] decode[182] decode[183] decode[184] decode[185] decode[186] decode[187] decode[188] decode[189] decode[190] decode[191] decode[192] decode[193] decode[194] decode[195] decode[196] decode[197] decode[198] decode[199] decode[200] decode[201] decode[202] decode[203] decode[204] decode[205] decode[206] decode[207] decode[208] decode[209] decode[210] decode[211] decode[212] decode[213] decode[214] decode[215] decode[216] decode[217] decode[218] decode[219] decode[220] decode[221] decode[222] decode[223] decode[224] decode[225] decode[226] decode[227] decode[228] decode[229] decode[230] decode[231] decode[232] decode[233] decode[234] decode[235] decode[236] decode[237] decode[238] decode[239] decode[240] decode[241] decode[242] decode[243] decode[244] decode[245] decode[246] decode[247] decode[248] decode[249] decode[250] decode[251] decode[252] decode[253] decode[254] decode[255] vdd gnd
Xpre[0] A[0] A[1] out[0] out[1] out[2] out[3] vdd gnd pre2x4
Xpre3x8[0] A[2] A[3] A[4] out[4] out[5] out[6] out[7] out[8] out[9] out[10] out[11] vdd gnd pre3x8
Xpre3x8[1] A[5] A[6] A[7] out[12] out[13] out[14] out[15] out[16] out[17] out[18] out[19] vdd gnd pre3x8
XDEC_NAND[0] out[0] out[4] out[12] Z[0] vdd gnd pnand3_2
XDEC_NAND[1] out[0] out[4] out[13] Z[1] vdd gnd pnand3_2
XDEC_NAND[2] out[0] out[4] out[14] Z[2] vdd gnd pnand3_2
XDEC_NAND[3] out[0] out[4] out[15] Z[3] vdd gnd pnand3_2
XDEC_NAND[4] out[0] out[4] out[16] Z[4] vdd gnd pnand3_2
XDEC_NAND[5] out[0] out[4] out[17] Z[5] vdd gnd pnand3_2
XDEC_NAND[6] out[0] out[4] out[18] Z[6] vdd gnd pnand3_2
XDEC_NAND[7] out[0] out[4] out[19] Z[7] vdd gnd pnand3_2
XDEC_NAND[8] out[0] out[5] out[12] Z[8] vdd gnd pnand3_2
XDEC_NAND[9] out[0] out[5] out[13] Z[9] vdd gnd pnand3_2
XDEC_NAND[10] out[0] out[5] out[14] Z[10] vdd gnd pnand3_2
XDEC_NAND[11] out[0] out[5] out[15] Z[11] vdd gnd pnand3_2
XDEC_NAND[12] out[0] out[5] out[16] Z[12] vdd gnd pnand3_2
XDEC_NAND[13] out[0] out[5] out[17] Z[13] vdd gnd pnand3_2
XDEC_NAND[14] out[0] out[5] out[18] Z[14] vdd gnd pnand3_2
XDEC_NAND[15] out[0] out[5] out[19] Z[15] vdd gnd pnand3_2
XDEC_NAND[16] out[0] out[6] out[12] Z[16] vdd gnd pnand3_2
XDEC_NAND[17] out[0] out[6] out[13] Z[17] vdd gnd pnand3_2
XDEC_NAND[18] out[0] out[6] out[14] Z[18] vdd gnd pnand3_2
XDEC_NAND[19] out[0] out[6] out[15] Z[19] vdd gnd pnand3_2
XDEC_NAND[20] out[0] out[6] out[16] Z[20] vdd gnd pnand3_2
XDEC_NAND[21] out[0] out[6] out[17] Z[21] vdd gnd pnand3_2
XDEC_NAND[22] out[0] out[6] out[18] Z[22] vdd gnd pnand3_2
XDEC_NAND[23] out[0] out[6] out[19] Z[23] vdd gnd pnand3_2
XDEC_NAND[24] out[0] out[7] out[12] Z[24] vdd gnd pnand3_2
XDEC_NAND[25] out[0] out[7] out[13] Z[25] vdd gnd pnand3_2
XDEC_NAND[26] out[0] out[7] out[14] Z[26] vdd gnd pnand3_2
XDEC_NAND[27] out[0] out[7] out[15] Z[27] vdd gnd pnand3_2
XDEC_NAND[28] out[0] out[7] out[16] Z[28] vdd gnd pnand3_2
XDEC_NAND[29] out[0] out[7] out[17] Z[29] vdd gnd pnand3_2
XDEC_NAND[30] out[0] out[7] out[18] Z[30] vdd gnd pnand3_2
XDEC_NAND[31] out[0] out[7] out[19] Z[31] vdd gnd pnand3_2
XDEC_NAND[32] out[0] out[8] out[12] Z[32] vdd gnd pnand3_2
XDEC_NAND[33] out[0] out[8] out[13] Z[33] vdd gnd pnand3_2
XDEC_NAND[34] out[0] out[8] out[14] Z[34] vdd gnd pnand3_2
XDEC_NAND[35] out[0] out[8] out[15] Z[35] vdd gnd pnand3_2
XDEC_NAND[36] out[0] out[8] out[16] Z[36] vdd gnd pnand3_2
XDEC_NAND[37] out[0] out[8] out[17] Z[37] vdd gnd pnand3_2
XDEC_NAND[38] out[0] out[8] out[18] Z[38] vdd gnd pnand3_2
XDEC_NAND[39] out[0] out[8] out[19] Z[39] vdd gnd pnand3_2
XDEC_NAND[40] out[0] out[9] out[12] Z[40] vdd gnd pnand3_2
XDEC_NAND[41] out[0] out[9] out[13] Z[41] vdd gnd pnand3_2
XDEC_NAND[42] out[0] out[9] out[14] Z[42] vdd gnd pnand3_2
XDEC_NAND[43] out[0] out[9] out[15] Z[43] vdd gnd pnand3_2
XDEC_NAND[44] out[0] out[9] out[16] Z[44] vdd gnd pnand3_2
XDEC_NAND[45] out[0] out[9] out[17] Z[45] vdd gnd pnand3_2
XDEC_NAND[46] out[0] out[9] out[18] Z[46] vdd gnd pnand3_2
XDEC_NAND[47] out[0] out[9] out[19] Z[47] vdd gnd pnand3_2
XDEC_NAND[48] out[0] out[10] out[12] Z[48] vdd gnd pnand3_2
XDEC_NAND[49] out[0] out[10] out[13] Z[49] vdd gnd pnand3_2
XDEC_NAND[50] out[0] out[10] out[14] Z[50] vdd gnd pnand3_2
XDEC_NAND[51] out[0] out[10] out[15] Z[51] vdd gnd pnand3_2
XDEC_NAND[52] out[0] out[10] out[16] Z[52] vdd gnd pnand3_2
XDEC_NAND[53] out[0] out[10] out[17] Z[53] vdd gnd pnand3_2
XDEC_NAND[54] out[0] out[10] out[18] Z[54] vdd gnd pnand3_2
XDEC_NAND[55] out[0] out[10] out[19] Z[55] vdd gnd pnand3_2
XDEC_NAND[56] out[0] out[11] out[12] Z[56] vdd gnd pnand3_2
XDEC_NAND[57] out[0] out[11] out[13] Z[57] vdd gnd pnand3_2
XDEC_NAND[58] out[0] out[11] out[14] Z[58] vdd gnd pnand3_2
XDEC_NAND[59] out[0] out[11] out[15] Z[59] vdd gnd pnand3_2
XDEC_NAND[60] out[0] out[11] out[16] Z[60] vdd gnd pnand3_2
XDEC_NAND[61] out[0] out[11] out[17] Z[61] vdd gnd pnand3_2
XDEC_NAND[62] out[0] out[11] out[18] Z[62] vdd gnd pnand3_2
XDEC_NAND[63] out[0] out[11] out[19] Z[63] vdd gnd pnand3_2
XDEC_NAND[64] out[1] out[4] out[12] Z[64] vdd gnd pnand3_2
XDEC_NAND[65] out[1] out[4] out[13] Z[65] vdd gnd pnand3_2
XDEC_NAND[66] out[1] out[4] out[14] Z[66] vdd gnd pnand3_2
XDEC_NAND[67] out[1] out[4] out[15] Z[67] vdd gnd pnand3_2
XDEC_NAND[68] out[1] out[4] out[16] Z[68] vdd gnd pnand3_2
XDEC_NAND[69] out[1] out[4] out[17] Z[69] vdd gnd pnand3_2
XDEC_NAND[70] out[1] out[4] out[18] Z[70] vdd gnd pnand3_2
XDEC_NAND[71] out[1] out[4] out[19] Z[71] vdd gnd pnand3_2
XDEC_NAND[72] out[1] out[5] out[12] Z[72] vdd gnd pnand3_2
XDEC_NAND[73] out[1] out[5] out[13] Z[73] vdd gnd pnand3_2
XDEC_NAND[74] out[1] out[5] out[14] Z[74] vdd gnd pnand3_2
XDEC_NAND[75] out[1] out[5] out[15] Z[75] vdd gnd pnand3_2
XDEC_NAND[76] out[1] out[5] out[16] Z[76] vdd gnd pnand3_2
XDEC_NAND[77] out[1] out[5] out[17] Z[77] vdd gnd pnand3_2
XDEC_NAND[78] out[1] out[5] out[18] Z[78] vdd gnd pnand3_2
XDEC_NAND[79] out[1] out[5] out[19] Z[79] vdd gnd pnand3_2
XDEC_NAND[80] out[1] out[6] out[12] Z[80] vdd gnd pnand3_2
XDEC_NAND[81] out[1] out[6] out[13] Z[81] vdd gnd pnand3_2
XDEC_NAND[82] out[1] out[6] out[14] Z[82] vdd gnd pnand3_2
XDEC_NAND[83] out[1] out[6] out[15] Z[83] vdd gnd pnand3_2
XDEC_NAND[84] out[1] out[6] out[16] Z[84] vdd gnd pnand3_2
XDEC_NAND[85] out[1] out[6] out[17] Z[85] vdd gnd pnand3_2
XDEC_NAND[86] out[1] out[6] out[18] Z[86] vdd gnd pnand3_2
XDEC_NAND[87] out[1] out[6] out[19] Z[87] vdd gnd pnand3_2
XDEC_NAND[88] out[1] out[7] out[12] Z[88] vdd gnd pnand3_2
XDEC_NAND[89] out[1] out[7] out[13] Z[89] vdd gnd pnand3_2
XDEC_NAND[90] out[1] out[7] out[14] Z[90] vdd gnd pnand3_2
XDEC_NAND[91] out[1] out[7] out[15] Z[91] vdd gnd pnand3_2
XDEC_NAND[92] out[1] out[7] out[16] Z[92] vdd gnd pnand3_2
XDEC_NAND[93] out[1] out[7] out[17] Z[93] vdd gnd pnand3_2
XDEC_NAND[94] out[1] out[7] out[18] Z[94] vdd gnd pnand3_2
XDEC_NAND[95] out[1] out[7] out[19] Z[95] vdd gnd pnand3_2
XDEC_NAND[96] out[1] out[8] out[12] Z[96] vdd gnd pnand3_2
XDEC_NAND[97] out[1] out[8] out[13] Z[97] vdd gnd pnand3_2
XDEC_NAND[98] out[1] out[8] out[14] Z[98] vdd gnd pnand3_2
XDEC_NAND[99] out[1] out[8] out[15] Z[99] vdd gnd pnand3_2
XDEC_NAND[100] out[1] out[8] out[16] Z[100] vdd gnd pnand3_2
XDEC_NAND[101] out[1] out[8] out[17] Z[101] vdd gnd pnand3_2
XDEC_NAND[102] out[1] out[8] out[18] Z[102] vdd gnd pnand3_2
XDEC_NAND[103] out[1] out[8] out[19] Z[103] vdd gnd pnand3_2
XDEC_NAND[104] out[1] out[9] out[12] Z[104] vdd gnd pnand3_2
XDEC_NAND[105] out[1] out[9] out[13] Z[105] vdd gnd pnand3_2
XDEC_NAND[106] out[1] out[9] out[14] Z[106] vdd gnd pnand3_2
XDEC_NAND[107] out[1] out[9] out[15] Z[107] vdd gnd pnand3_2
XDEC_NAND[108] out[1] out[9] out[16] Z[108] vdd gnd pnand3_2
XDEC_NAND[109] out[1] out[9] out[17] Z[109] vdd gnd pnand3_2
XDEC_NAND[110] out[1] out[9] out[18] Z[110] vdd gnd pnand3_2
XDEC_NAND[111] out[1] out[9] out[19] Z[111] vdd gnd pnand3_2
XDEC_NAND[112] out[1] out[10] out[12] Z[112] vdd gnd pnand3_2
XDEC_NAND[113] out[1] out[10] out[13] Z[113] vdd gnd pnand3_2
XDEC_NAND[114] out[1] out[10] out[14] Z[114] vdd gnd pnand3_2
XDEC_NAND[115] out[1] out[10] out[15] Z[115] vdd gnd pnand3_2
XDEC_NAND[116] out[1] out[10] out[16] Z[116] vdd gnd pnand3_2
XDEC_NAND[117] out[1] out[10] out[17] Z[117] vdd gnd pnand3_2
XDEC_NAND[118] out[1] out[10] out[18] Z[118] vdd gnd pnand3_2
XDEC_NAND[119] out[1] out[10] out[19] Z[119] vdd gnd pnand3_2
XDEC_NAND[120] out[1] out[11] out[12] Z[120] vdd gnd pnand3_2
XDEC_NAND[121] out[1] out[11] out[13] Z[121] vdd gnd pnand3_2
XDEC_NAND[122] out[1] out[11] out[14] Z[122] vdd gnd pnand3_2
XDEC_NAND[123] out[1] out[11] out[15] Z[123] vdd gnd pnand3_2
XDEC_NAND[124] out[1] out[11] out[16] Z[124] vdd gnd pnand3_2
XDEC_NAND[125] out[1] out[11] out[17] Z[125] vdd gnd pnand3_2
XDEC_NAND[126] out[1] out[11] out[18] Z[126] vdd gnd pnand3_2
XDEC_NAND[127] out[1] out[11] out[19] Z[127] vdd gnd pnand3_2
XDEC_NAND[128] out[2] out[4] out[12] Z[128] vdd gnd pnand3_2
XDEC_NAND[129] out[2] out[4] out[13] Z[129] vdd gnd pnand3_2
XDEC_NAND[130] out[2] out[4] out[14] Z[130] vdd gnd pnand3_2
XDEC_NAND[131] out[2] out[4] out[15] Z[131] vdd gnd pnand3_2
XDEC_NAND[132] out[2] out[4] out[16] Z[132] vdd gnd pnand3_2
XDEC_NAND[133] out[2] out[4] out[17] Z[133] vdd gnd pnand3_2
XDEC_NAND[134] out[2] out[4] out[18] Z[134] vdd gnd pnand3_2
XDEC_NAND[135] out[2] out[4] out[19] Z[135] vdd gnd pnand3_2
XDEC_NAND[136] out[2] out[5] out[12] Z[136] vdd gnd pnand3_2
XDEC_NAND[137] out[2] out[5] out[13] Z[137] vdd gnd pnand3_2
XDEC_NAND[138] out[2] out[5] out[14] Z[138] vdd gnd pnand3_2
XDEC_NAND[139] out[2] out[5] out[15] Z[139] vdd gnd pnand3_2
XDEC_NAND[140] out[2] out[5] out[16] Z[140] vdd gnd pnand3_2
XDEC_NAND[141] out[2] out[5] out[17] Z[141] vdd gnd pnand3_2
XDEC_NAND[142] out[2] out[5] out[18] Z[142] vdd gnd pnand3_2
XDEC_NAND[143] out[2] out[5] out[19] Z[143] vdd gnd pnand3_2
XDEC_NAND[144] out[2] out[6] out[12] Z[144] vdd gnd pnand3_2
XDEC_NAND[145] out[2] out[6] out[13] Z[145] vdd gnd pnand3_2
XDEC_NAND[146] out[2] out[6] out[14] Z[146] vdd gnd pnand3_2
XDEC_NAND[147] out[2] out[6] out[15] Z[147] vdd gnd pnand3_2
XDEC_NAND[148] out[2] out[6] out[16] Z[148] vdd gnd pnand3_2
XDEC_NAND[149] out[2] out[6] out[17] Z[149] vdd gnd pnand3_2
XDEC_NAND[150] out[2] out[6] out[18] Z[150] vdd gnd pnand3_2
XDEC_NAND[151] out[2] out[6] out[19] Z[151] vdd gnd pnand3_2
XDEC_NAND[152] out[2] out[7] out[12] Z[152] vdd gnd pnand3_2
XDEC_NAND[153] out[2] out[7] out[13] Z[153] vdd gnd pnand3_2
XDEC_NAND[154] out[2] out[7] out[14] Z[154] vdd gnd pnand3_2
XDEC_NAND[155] out[2] out[7] out[15] Z[155] vdd gnd pnand3_2
XDEC_NAND[156] out[2] out[7] out[16] Z[156] vdd gnd pnand3_2
XDEC_NAND[157] out[2] out[7] out[17] Z[157] vdd gnd pnand3_2
XDEC_NAND[158] out[2] out[7] out[18] Z[158] vdd gnd pnand3_2
XDEC_NAND[159] out[2] out[7] out[19] Z[159] vdd gnd pnand3_2
XDEC_NAND[160] out[2] out[8] out[12] Z[160] vdd gnd pnand3_2
XDEC_NAND[161] out[2] out[8] out[13] Z[161] vdd gnd pnand3_2
XDEC_NAND[162] out[2] out[8] out[14] Z[162] vdd gnd pnand3_2
XDEC_NAND[163] out[2] out[8] out[15] Z[163] vdd gnd pnand3_2
XDEC_NAND[164] out[2] out[8] out[16] Z[164] vdd gnd pnand3_2
XDEC_NAND[165] out[2] out[8] out[17] Z[165] vdd gnd pnand3_2
XDEC_NAND[166] out[2] out[8] out[18] Z[166] vdd gnd pnand3_2
XDEC_NAND[167] out[2] out[8] out[19] Z[167] vdd gnd pnand3_2
XDEC_NAND[168] out[2] out[9] out[12] Z[168] vdd gnd pnand3_2
XDEC_NAND[169] out[2] out[9] out[13] Z[169] vdd gnd pnand3_2
XDEC_NAND[170] out[2] out[9] out[14] Z[170] vdd gnd pnand3_2
XDEC_NAND[171] out[2] out[9] out[15] Z[171] vdd gnd pnand3_2
XDEC_NAND[172] out[2] out[9] out[16] Z[172] vdd gnd pnand3_2
XDEC_NAND[173] out[2] out[9] out[17] Z[173] vdd gnd pnand3_2
XDEC_NAND[174] out[2] out[9] out[18] Z[174] vdd gnd pnand3_2
XDEC_NAND[175] out[2] out[9] out[19] Z[175] vdd gnd pnand3_2
XDEC_NAND[176] out[2] out[10] out[12] Z[176] vdd gnd pnand3_2
XDEC_NAND[177] out[2] out[10] out[13] Z[177] vdd gnd pnand3_2
XDEC_NAND[178] out[2] out[10] out[14] Z[178] vdd gnd pnand3_2
XDEC_NAND[179] out[2] out[10] out[15] Z[179] vdd gnd pnand3_2
XDEC_NAND[180] out[2] out[10] out[16] Z[180] vdd gnd pnand3_2
XDEC_NAND[181] out[2] out[10] out[17] Z[181] vdd gnd pnand3_2
XDEC_NAND[182] out[2] out[10] out[18] Z[182] vdd gnd pnand3_2
XDEC_NAND[183] out[2] out[10] out[19] Z[183] vdd gnd pnand3_2
XDEC_NAND[184] out[2] out[11] out[12] Z[184] vdd gnd pnand3_2
XDEC_NAND[185] out[2] out[11] out[13] Z[185] vdd gnd pnand3_2
XDEC_NAND[186] out[2] out[11] out[14] Z[186] vdd gnd pnand3_2
XDEC_NAND[187] out[2] out[11] out[15] Z[187] vdd gnd pnand3_2
XDEC_NAND[188] out[2] out[11] out[16] Z[188] vdd gnd pnand3_2
XDEC_NAND[189] out[2] out[11] out[17] Z[189] vdd gnd pnand3_2
XDEC_NAND[190] out[2] out[11] out[18] Z[190] vdd gnd pnand3_2
XDEC_NAND[191] out[2] out[11] out[19] Z[191] vdd gnd pnand3_2
XDEC_NAND[192] out[3] out[4] out[12] Z[192] vdd gnd pnand3_2
XDEC_NAND[193] out[3] out[4] out[13] Z[193] vdd gnd pnand3_2
XDEC_NAND[194] out[3] out[4] out[14] Z[194] vdd gnd pnand3_2
XDEC_NAND[195] out[3] out[4] out[15] Z[195] vdd gnd pnand3_2
XDEC_NAND[196] out[3] out[4] out[16] Z[196] vdd gnd pnand3_2
XDEC_NAND[197] out[3] out[4] out[17] Z[197] vdd gnd pnand3_2
XDEC_NAND[198] out[3] out[4] out[18] Z[198] vdd gnd pnand3_2
XDEC_NAND[199] out[3] out[4] out[19] Z[199] vdd gnd pnand3_2
XDEC_NAND[200] out[3] out[5] out[12] Z[200] vdd gnd pnand3_2
XDEC_NAND[201] out[3] out[5] out[13] Z[201] vdd gnd pnand3_2
XDEC_NAND[202] out[3] out[5] out[14] Z[202] vdd gnd pnand3_2
XDEC_NAND[203] out[3] out[5] out[15] Z[203] vdd gnd pnand3_2
XDEC_NAND[204] out[3] out[5] out[16] Z[204] vdd gnd pnand3_2
XDEC_NAND[205] out[3] out[5] out[17] Z[205] vdd gnd pnand3_2
XDEC_NAND[206] out[3] out[5] out[18] Z[206] vdd gnd pnand3_2
XDEC_NAND[207] out[3] out[5] out[19] Z[207] vdd gnd pnand3_2
XDEC_NAND[208] out[3] out[6] out[12] Z[208] vdd gnd pnand3_2
XDEC_NAND[209] out[3] out[6] out[13] Z[209] vdd gnd pnand3_2
XDEC_NAND[210] out[3] out[6] out[14] Z[210] vdd gnd pnand3_2
XDEC_NAND[211] out[3] out[6] out[15] Z[211] vdd gnd pnand3_2
XDEC_NAND[212] out[3] out[6] out[16] Z[212] vdd gnd pnand3_2
XDEC_NAND[213] out[3] out[6] out[17] Z[213] vdd gnd pnand3_2
XDEC_NAND[214] out[3] out[6] out[18] Z[214] vdd gnd pnand3_2
XDEC_NAND[215] out[3] out[6] out[19] Z[215] vdd gnd pnand3_2
XDEC_NAND[216] out[3] out[7] out[12] Z[216] vdd gnd pnand3_2
XDEC_NAND[217] out[3] out[7] out[13] Z[217] vdd gnd pnand3_2
XDEC_NAND[218] out[3] out[7] out[14] Z[218] vdd gnd pnand3_2
XDEC_NAND[219] out[3] out[7] out[15] Z[219] vdd gnd pnand3_2
XDEC_NAND[220] out[3] out[7] out[16] Z[220] vdd gnd pnand3_2
XDEC_NAND[221] out[3] out[7] out[17] Z[221] vdd gnd pnand3_2
XDEC_NAND[222] out[3] out[7] out[18] Z[222] vdd gnd pnand3_2
XDEC_NAND[223] out[3] out[7] out[19] Z[223] vdd gnd pnand3_2
XDEC_NAND[224] out[3] out[8] out[12] Z[224] vdd gnd pnand3_2
XDEC_NAND[225] out[3] out[8] out[13] Z[225] vdd gnd pnand3_2
XDEC_NAND[226] out[3] out[8] out[14] Z[226] vdd gnd pnand3_2
XDEC_NAND[227] out[3] out[8] out[15] Z[227] vdd gnd pnand3_2
XDEC_NAND[228] out[3] out[8] out[16] Z[228] vdd gnd pnand3_2
XDEC_NAND[229] out[3] out[8] out[17] Z[229] vdd gnd pnand3_2
XDEC_NAND[230] out[3] out[8] out[18] Z[230] vdd gnd pnand3_2
XDEC_NAND[231] out[3] out[8] out[19] Z[231] vdd gnd pnand3_2
XDEC_NAND[232] out[3] out[9] out[12] Z[232] vdd gnd pnand3_2
XDEC_NAND[233] out[3] out[9] out[13] Z[233] vdd gnd pnand3_2
XDEC_NAND[234] out[3] out[9] out[14] Z[234] vdd gnd pnand3_2
XDEC_NAND[235] out[3] out[9] out[15] Z[235] vdd gnd pnand3_2
XDEC_NAND[236] out[3] out[9] out[16] Z[236] vdd gnd pnand3_2
XDEC_NAND[237] out[3] out[9] out[17] Z[237] vdd gnd pnand3_2
XDEC_NAND[238] out[3] out[9] out[18] Z[238] vdd gnd pnand3_2
XDEC_NAND[239] out[3] out[9] out[19] Z[239] vdd gnd pnand3_2
XDEC_NAND[240] out[3] out[10] out[12] Z[240] vdd gnd pnand3_2
XDEC_NAND[241] out[3] out[10] out[13] Z[241] vdd gnd pnand3_2
XDEC_NAND[242] out[3] out[10] out[14] Z[242] vdd gnd pnand3_2
XDEC_NAND[243] out[3] out[10] out[15] Z[243] vdd gnd pnand3_2
XDEC_NAND[244] out[3] out[10] out[16] Z[244] vdd gnd pnand3_2
XDEC_NAND[245] out[3] out[10] out[17] Z[245] vdd gnd pnand3_2
XDEC_NAND[246] out[3] out[10] out[18] Z[246] vdd gnd pnand3_2
XDEC_NAND[247] out[3] out[10] out[19] Z[247] vdd gnd pnand3_2
XDEC_NAND[248] out[3] out[11] out[12] Z[248] vdd gnd pnand3_2
XDEC_NAND[249] out[3] out[11] out[13] Z[249] vdd gnd pnand3_2
XDEC_NAND[250] out[3] out[11] out[14] Z[250] vdd gnd pnand3_2
XDEC_NAND[251] out[3] out[11] out[15] Z[251] vdd gnd pnand3_2
XDEC_NAND[252] out[3] out[11] out[16] Z[252] vdd gnd pnand3_2
XDEC_NAND[253] out[3] out[11] out[17] Z[253] vdd gnd pnand3_2
XDEC_NAND[254] out[3] out[11] out[18] Z[254] vdd gnd pnand3_2
XDEC_NAND[255] out[3] out[11] out[19] Z[255] vdd gnd pnand3_2
XDEC_INV_[0] Z[0] decode[0] vdd gnd pinv_8
XDEC_INV_[1] Z[1] decode[1] vdd gnd pinv_8
XDEC_INV_[2] Z[2] decode[2] vdd gnd pinv_8
XDEC_INV_[3] Z[3] decode[3] vdd gnd pinv_8
XDEC_INV_[4] Z[4] decode[4] vdd gnd pinv_8
XDEC_INV_[5] Z[5] decode[5] vdd gnd pinv_8
XDEC_INV_[6] Z[6] decode[6] vdd gnd pinv_8
XDEC_INV_[7] Z[7] decode[7] vdd gnd pinv_8
XDEC_INV_[8] Z[8] decode[8] vdd gnd pinv_8
XDEC_INV_[9] Z[9] decode[9] vdd gnd pinv_8
XDEC_INV_[10] Z[10] decode[10] vdd gnd pinv_8
XDEC_INV_[11] Z[11] decode[11] vdd gnd pinv_8
XDEC_INV_[12] Z[12] decode[12] vdd gnd pinv_8
XDEC_INV_[13] Z[13] decode[13] vdd gnd pinv_8
XDEC_INV_[14] Z[14] decode[14] vdd gnd pinv_8
XDEC_INV_[15] Z[15] decode[15] vdd gnd pinv_8
XDEC_INV_[16] Z[16] decode[16] vdd gnd pinv_8
XDEC_INV_[17] Z[17] decode[17] vdd gnd pinv_8
XDEC_INV_[18] Z[18] decode[18] vdd gnd pinv_8
XDEC_INV_[19] Z[19] decode[19] vdd gnd pinv_8
XDEC_INV_[20] Z[20] decode[20] vdd gnd pinv_8
XDEC_INV_[21] Z[21] decode[21] vdd gnd pinv_8
XDEC_INV_[22] Z[22] decode[22] vdd gnd pinv_8
XDEC_INV_[23] Z[23] decode[23] vdd gnd pinv_8
XDEC_INV_[24] Z[24] decode[24] vdd gnd pinv_8
XDEC_INV_[25] Z[25] decode[25] vdd gnd pinv_8
XDEC_INV_[26] Z[26] decode[26] vdd gnd pinv_8
XDEC_INV_[27] Z[27] decode[27] vdd gnd pinv_8
XDEC_INV_[28] Z[28] decode[28] vdd gnd pinv_8
XDEC_INV_[29] Z[29] decode[29] vdd gnd pinv_8
XDEC_INV_[30] Z[30] decode[30] vdd gnd pinv_8
XDEC_INV_[31] Z[31] decode[31] vdd gnd pinv_8
XDEC_INV_[32] Z[32] decode[32] vdd gnd pinv_8
XDEC_INV_[33] Z[33] decode[33] vdd gnd pinv_8
XDEC_INV_[34] Z[34] decode[34] vdd gnd pinv_8
XDEC_INV_[35] Z[35] decode[35] vdd gnd pinv_8
XDEC_INV_[36] Z[36] decode[36] vdd gnd pinv_8
XDEC_INV_[37] Z[37] decode[37] vdd gnd pinv_8
XDEC_INV_[38] Z[38] decode[38] vdd gnd pinv_8
XDEC_INV_[39] Z[39] decode[39] vdd gnd pinv_8
XDEC_INV_[40] Z[40] decode[40] vdd gnd pinv_8
XDEC_INV_[41] Z[41] decode[41] vdd gnd pinv_8
XDEC_INV_[42] Z[42] decode[42] vdd gnd pinv_8
XDEC_INV_[43] Z[43] decode[43] vdd gnd pinv_8
XDEC_INV_[44] Z[44] decode[44] vdd gnd pinv_8
XDEC_INV_[45] Z[45] decode[45] vdd gnd pinv_8
XDEC_INV_[46] Z[46] decode[46] vdd gnd pinv_8
XDEC_INV_[47] Z[47] decode[47] vdd gnd pinv_8
XDEC_INV_[48] Z[48] decode[48] vdd gnd pinv_8
XDEC_INV_[49] Z[49] decode[49] vdd gnd pinv_8
XDEC_INV_[50] Z[50] decode[50] vdd gnd pinv_8
XDEC_INV_[51] Z[51] decode[51] vdd gnd pinv_8
XDEC_INV_[52] Z[52] decode[52] vdd gnd pinv_8
XDEC_INV_[53] Z[53] decode[53] vdd gnd pinv_8
XDEC_INV_[54] Z[54] decode[54] vdd gnd pinv_8
XDEC_INV_[55] Z[55] decode[55] vdd gnd pinv_8
XDEC_INV_[56] Z[56] decode[56] vdd gnd pinv_8
XDEC_INV_[57] Z[57] decode[57] vdd gnd pinv_8
XDEC_INV_[58] Z[58] decode[58] vdd gnd pinv_8
XDEC_INV_[59] Z[59] decode[59] vdd gnd pinv_8
XDEC_INV_[60] Z[60] decode[60] vdd gnd pinv_8
XDEC_INV_[61] Z[61] decode[61] vdd gnd pinv_8
XDEC_INV_[62] Z[62] decode[62] vdd gnd pinv_8
XDEC_INV_[63] Z[63] decode[63] vdd gnd pinv_8
XDEC_INV_[64] Z[64] decode[64] vdd gnd pinv_8
XDEC_INV_[65] Z[65] decode[65] vdd gnd pinv_8
XDEC_INV_[66] Z[66] decode[66] vdd gnd pinv_8
XDEC_INV_[67] Z[67] decode[67] vdd gnd pinv_8
XDEC_INV_[68] Z[68] decode[68] vdd gnd pinv_8
XDEC_INV_[69] Z[69] decode[69] vdd gnd pinv_8
XDEC_INV_[70] Z[70] decode[70] vdd gnd pinv_8
XDEC_INV_[71] Z[71] decode[71] vdd gnd pinv_8
XDEC_INV_[72] Z[72] decode[72] vdd gnd pinv_8
XDEC_INV_[73] Z[73] decode[73] vdd gnd pinv_8
XDEC_INV_[74] Z[74] decode[74] vdd gnd pinv_8
XDEC_INV_[75] Z[75] decode[75] vdd gnd pinv_8
XDEC_INV_[76] Z[76] decode[76] vdd gnd pinv_8
XDEC_INV_[77] Z[77] decode[77] vdd gnd pinv_8
XDEC_INV_[78] Z[78] decode[78] vdd gnd pinv_8
XDEC_INV_[79] Z[79] decode[79] vdd gnd pinv_8
XDEC_INV_[80] Z[80] decode[80] vdd gnd pinv_8
XDEC_INV_[81] Z[81] decode[81] vdd gnd pinv_8
XDEC_INV_[82] Z[82] decode[82] vdd gnd pinv_8
XDEC_INV_[83] Z[83] decode[83] vdd gnd pinv_8
XDEC_INV_[84] Z[84] decode[84] vdd gnd pinv_8
XDEC_INV_[85] Z[85] decode[85] vdd gnd pinv_8
XDEC_INV_[86] Z[86] decode[86] vdd gnd pinv_8
XDEC_INV_[87] Z[87] decode[87] vdd gnd pinv_8
XDEC_INV_[88] Z[88] decode[88] vdd gnd pinv_8
XDEC_INV_[89] Z[89] decode[89] vdd gnd pinv_8
XDEC_INV_[90] Z[90] decode[90] vdd gnd pinv_8
XDEC_INV_[91] Z[91] decode[91] vdd gnd pinv_8
XDEC_INV_[92] Z[92] decode[92] vdd gnd pinv_8
XDEC_INV_[93] Z[93] decode[93] vdd gnd pinv_8
XDEC_INV_[94] Z[94] decode[94] vdd gnd pinv_8
XDEC_INV_[95] Z[95] decode[95] vdd gnd pinv_8
XDEC_INV_[96] Z[96] decode[96] vdd gnd pinv_8
XDEC_INV_[97] Z[97] decode[97] vdd gnd pinv_8
XDEC_INV_[98] Z[98] decode[98] vdd gnd pinv_8
XDEC_INV_[99] Z[99] decode[99] vdd gnd pinv_8
XDEC_INV_[100] Z[100] decode[100] vdd gnd pinv_8
XDEC_INV_[101] Z[101] decode[101] vdd gnd pinv_8
XDEC_INV_[102] Z[102] decode[102] vdd gnd pinv_8
XDEC_INV_[103] Z[103] decode[103] vdd gnd pinv_8
XDEC_INV_[104] Z[104] decode[104] vdd gnd pinv_8
XDEC_INV_[105] Z[105] decode[105] vdd gnd pinv_8
XDEC_INV_[106] Z[106] decode[106] vdd gnd pinv_8
XDEC_INV_[107] Z[107] decode[107] vdd gnd pinv_8
XDEC_INV_[108] Z[108] decode[108] vdd gnd pinv_8
XDEC_INV_[109] Z[109] decode[109] vdd gnd pinv_8
XDEC_INV_[110] Z[110] decode[110] vdd gnd pinv_8
XDEC_INV_[111] Z[111] decode[111] vdd gnd pinv_8
XDEC_INV_[112] Z[112] decode[112] vdd gnd pinv_8
XDEC_INV_[113] Z[113] decode[113] vdd gnd pinv_8
XDEC_INV_[114] Z[114] decode[114] vdd gnd pinv_8
XDEC_INV_[115] Z[115] decode[115] vdd gnd pinv_8
XDEC_INV_[116] Z[116] decode[116] vdd gnd pinv_8
XDEC_INV_[117] Z[117] decode[117] vdd gnd pinv_8
XDEC_INV_[118] Z[118] decode[118] vdd gnd pinv_8
XDEC_INV_[119] Z[119] decode[119] vdd gnd pinv_8
XDEC_INV_[120] Z[120] decode[120] vdd gnd pinv_8
XDEC_INV_[121] Z[121] decode[121] vdd gnd pinv_8
XDEC_INV_[122] Z[122] decode[122] vdd gnd pinv_8
XDEC_INV_[123] Z[123] decode[123] vdd gnd pinv_8
XDEC_INV_[124] Z[124] decode[124] vdd gnd pinv_8
XDEC_INV_[125] Z[125] decode[125] vdd gnd pinv_8
XDEC_INV_[126] Z[126] decode[126] vdd gnd pinv_8
XDEC_INV_[127] Z[127] decode[127] vdd gnd pinv_8
XDEC_INV_[128] Z[128] decode[128] vdd gnd pinv_8
XDEC_INV_[129] Z[129] decode[129] vdd gnd pinv_8
XDEC_INV_[130] Z[130] decode[130] vdd gnd pinv_8
XDEC_INV_[131] Z[131] decode[131] vdd gnd pinv_8
XDEC_INV_[132] Z[132] decode[132] vdd gnd pinv_8
XDEC_INV_[133] Z[133] decode[133] vdd gnd pinv_8
XDEC_INV_[134] Z[134] decode[134] vdd gnd pinv_8
XDEC_INV_[135] Z[135] decode[135] vdd gnd pinv_8
XDEC_INV_[136] Z[136] decode[136] vdd gnd pinv_8
XDEC_INV_[137] Z[137] decode[137] vdd gnd pinv_8
XDEC_INV_[138] Z[138] decode[138] vdd gnd pinv_8
XDEC_INV_[139] Z[139] decode[139] vdd gnd pinv_8
XDEC_INV_[140] Z[140] decode[140] vdd gnd pinv_8
XDEC_INV_[141] Z[141] decode[141] vdd gnd pinv_8
XDEC_INV_[142] Z[142] decode[142] vdd gnd pinv_8
XDEC_INV_[143] Z[143] decode[143] vdd gnd pinv_8
XDEC_INV_[144] Z[144] decode[144] vdd gnd pinv_8
XDEC_INV_[145] Z[145] decode[145] vdd gnd pinv_8
XDEC_INV_[146] Z[146] decode[146] vdd gnd pinv_8
XDEC_INV_[147] Z[147] decode[147] vdd gnd pinv_8
XDEC_INV_[148] Z[148] decode[148] vdd gnd pinv_8
XDEC_INV_[149] Z[149] decode[149] vdd gnd pinv_8
XDEC_INV_[150] Z[150] decode[150] vdd gnd pinv_8
XDEC_INV_[151] Z[151] decode[151] vdd gnd pinv_8
XDEC_INV_[152] Z[152] decode[152] vdd gnd pinv_8
XDEC_INV_[153] Z[153] decode[153] vdd gnd pinv_8
XDEC_INV_[154] Z[154] decode[154] vdd gnd pinv_8
XDEC_INV_[155] Z[155] decode[155] vdd gnd pinv_8
XDEC_INV_[156] Z[156] decode[156] vdd gnd pinv_8
XDEC_INV_[157] Z[157] decode[157] vdd gnd pinv_8
XDEC_INV_[158] Z[158] decode[158] vdd gnd pinv_8
XDEC_INV_[159] Z[159] decode[159] vdd gnd pinv_8
XDEC_INV_[160] Z[160] decode[160] vdd gnd pinv_8
XDEC_INV_[161] Z[161] decode[161] vdd gnd pinv_8
XDEC_INV_[162] Z[162] decode[162] vdd gnd pinv_8
XDEC_INV_[163] Z[163] decode[163] vdd gnd pinv_8
XDEC_INV_[164] Z[164] decode[164] vdd gnd pinv_8
XDEC_INV_[165] Z[165] decode[165] vdd gnd pinv_8
XDEC_INV_[166] Z[166] decode[166] vdd gnd pinv_8
XDEC_INV_[167] Z[167] decode[167] vdd gnd pinv_8
XDEC_INV_[168] Z[168] decode[168] vdd gnd pinv_8
XDEC_INV_[169] Z[169] decode[169] vdd gnd pinv_8
XDEC_INV_[170] Z[170] decode[170] vdd gnd pinv_8
XDEC_INV_[171] Z[171] decode[171] vdd gnd pinv_8
XDEC_INV_[172] Z[172] decode[172] vdd gnd pinv_8
XDEC_INV_[173] Z[173] decode[173] vdd gnd pinv_8
XDEC_INV_[174] Z[174] decode[174] vdd gnd pinv_8
XDEC_INV_[175] Z[175] decode[175] vdd gnd pinv_8
XDEC_INV_[176] Z[176] decode[176] vdd gnd pinv_8
XDEC_INV_[177] Z[177] decode[177] vdd gnd pinv_8
XDEC_INV_[178] Z[178] decode[178] vdd gnd pinv_8
XDEC_INV_[179] Z[179] decode[179] vdd gnd pinv_8
XDEC_INV_[180] Z[180] decode[180] vdd gnd pinv_8
XDEC_INV_[181] Z[181] decode[181] vdd gnd pinv_8
XDEC_INV_[182] Z[182] decode[182] vdd gnd pinv_8
XDEC_INV_[183] Z[183] decode[183] vdd gnd pinv_8
XDEC_INV_[184] Z[184] decode[184] vdd gnd pinv_8
XDEC_INV_[185] Z[185] decode[185] vdd gnd pinv_8
XDEC_INV_[186] Z[186] decode[186] vdd gnd pinv_8
XDEC_INV_[187] Z[187] decode[187] vdd gnd pinv_8
XDEC_INV_[188] Z[188] decode[188] vdd gnd pinv_8
XDEC_INV_[189] Z[189] decode[189] vdd gnd pinv_8
XDEC_INV_[190] Z[190] decode[190] vdd gnd pinv_8
XDEC_INV_[191] Z[191] decode[191] vdd gnd pinv_8
XDEC_INV_[192] Z[192] decode[192] vdd gnd pinv_8
XDEC_INV_[193] Z[193] decode[193] vdd gnd pinv_8
XDEC_INV_[194] Z[194] decode[194] vdd gnd pinv_8
XDEC_INV_[195] Z[195] decode[195] vdd gnd pinv_8
XDEC_INV_[196] Z[196] decode[196] vdd gnd pinv_8
XDEC_INV_[197] Z[197] decode[197] vdd gnd pinv_8
XDEC_INV_[198] Z[198] decode[198] vdd gnd pinv_8
XDEC_INV_[199] Z[199] decode[199] vdd gnd pinv_8
XDEC_INV_[200] Z[200] decode[200] vdd gnd pinv_8
XDEC_INV_[201] Z[201] decode[201] vdd gnd pinv_8
XDEC_INV_[202] Z[202] decode[202] vdd gnd pinv_8
XDEC_INV_[203] Z[203] decode[203] vdd gnd pinv_8
XDEC_INV_[204] Z[204] decode[204] vdd gnd pinv_8
XDEC_INV_[205] Z[205] decode[205] vdd gnd pinv_8
XDEC_INV_[206] Z[206] decode[206] vdd gnd pinv_8
XDEC_INV_[207] Z[207] decode[207] vdd gnd pinv_8
XDEC_INV_[208] Z[208] decode[208] vdd gnd pinv_8
XDEC_INV_[209] Z[209] decode[209] vdd gnd pinv_8
XDEC_INV_[210] Z[210] decode[210] vdd gnd pinv_8
XDEC_INV_[211] Z[211] decode[211] vdd gnd pinv_8
XDEC_INV_[212] Z[212] decode[212] vdd gnd pinv_8
XDEC_INV_[213] Z[213] decode[213] vdd gnd pinv_8
XDEC_INV_[214] Z[214] decode[214] vdd gnd pinv_8
XDEC_INV_[215] Z[215] decode[215] vdd gnd pinv_8
XDEC_INV_[216] Z[216] decode[216] vdd gnd pinv_8
XDEC_INV_[217] Z[217] decode[217] vdd gnd pinv_8
XDEC_INV_[218] Z[218] decode[218] vdd gnd pinv_8
XDEC_INV_[219] Z[219] decode[219] vdd gnd pinv_8
XDEC_INV_[220] Z[220] decode[220] vdd gnd pinv_8
XDEC_INV_[221] Z[221] decode[221] vdd gnd pinv_8
XDEC_INV_[222] Z[222] decode[222] vdd gnd pinv_8
XDEC_INV_[223] Z[223] decode[223] vdd gnd pinv_8
XDEC_INV_[224] Z[224] decode[224] vdd gnd pinv_8
XDEC_INV_[225] Z[225] decode[225] vdd gnd pinv_8
XDEC_INV_[226] Z[226] decode[226] vdd gnd pinv_8
XDEC_INV_[227] Z[227] decode[227] vdd gnd pinv_8
XDEC_INV_[228] Z[228] decode[228] vdd gnd pinv_8
XDEC_INV_[229] Z[229] decode[229] vdd gnd pinv_8
XDEC_INV_[230] Z[230] decode[230] vdd gnd pinv_8
XDEC_INV_[231] Z[231] decode[231] vdd gnd pinv_8
XDEC_INV_[232] Z[232] decode[232] vdd gnd pinv_8
XDEC_INV_[233] Z[233] decode[233] vdd gnd pinv_8
XDEC_INV_[234] Z[234] decode[234] vdd gnd pinv_8
XDEC_INV_[235] Z[235] decode[235] vdd gnd pinv_8
XDEC_INV_[236] Z[236] decode[236] vdd gnd pinv_8
XDEC_INV_[237] Z[237] decode[237] vdd gnd pinv_8
XDEC_INV_[238] Z[238] decode[238] vdd gnd pinv_8
XDEC_INV_[239] Z[239] decode[239] vdd gnd pinv_8
XDEC_INV_[240] Z[240] decode[240] vdd gnd pinv_8
XDEC_INV_[241] Z[241] decode[241] vdd gnd pinv_8
XDEC_INV_[242] Z[242] decode[242] vdd gnd pinv_8
XDEC_INV_[243] Z[243] decode[243] vdd gnd pinv_8
XDEC_INV_[244] Z[244] decode[244] vdd gnd pinv_8
XDEC_INV_[245] Z[245] decode[245] vdd gnd pinv_8
XDEC_INV_[246] Z[246] decode[246] vdd gnd pinv_8
XDEC_INV_[247] Z[247] decode[247] vdd gnd pinv_8
XDEC_INV_[248] Z[248] decode[248] vdd gnd pinv_8
XDEC_INV_[249] Z[249] decode[249] vdd gnd pinv_8
XDEC_INV_[250] Z[250] decode[250] vdd gnd pinv_8
XDEC_INV_[251] Z[251] decode[251] vdd gnd pinv_8
XDEC_INV_[252] Z[252] decode[252] vdd gnd pinv_8
XDEC_INV_[253] Z[253] decode[253] vdd gnd pinv_8
XDEC_INV_[254] Z[254] decode[254] vdd gnd pinv_8
XDEC_INV_[255] Z[255] decode[255] vdd gnd pinv_8
.ENDS hierarchical_decoder_256rows

.SUBCKT msf_address din[0] din[1] din[2] din[3] din[4] din[5] din[6] din[7] din[8] dout[0] dout_bar[0] dout[1] dout_bar[1] dout[2] dout_bar[2] dout[3] dout_bar[3] dout[4] dout_bar[4] dout[5] dout_bar[5] dout[6] dout_bar[6] dout[7] dout_bar[7] dout[8] dout_bar[8] clk vdd gnd
XXdff0 din[0] dout[0] dout_bar[0] clk vdd gnd ms_flop
XXdff1 din[1] dout[1] dout_bar[1] clk vdd gnd ms_flop
XXdff2 din[2] dout[2] dout_bar[2] clk vdd gnd ms_flop
XXdff3 din[3] dout[3] dout_bar[3] clk vdd gnd ms_flop
XXdff4 din[4] dout[4] dout_bar[4] clk vdd gnd ms_flop
XXdff5 din[5] dout[5] dout_bar[5] clk vdd gnd ms_flop
XXdff6 din[6] dout[6] dout_bar[6] clk vdd gnd ms_flop
XXdff7 din[7] dout[7] dout_bar[7] clk vdd gnd ms_flop
XXdff8 din[8] dout[8] dout_bar[8] clk vdd gnd ms_flop
.ENDS msf_address

.SUBCKT msf_data_in din[0] din[1] din[2] din[3] din[4] din[5] din[6] din[7] din[8] din[9] din[10] din[11] din[12] din[13] din[14] din[15] din[16] din[17] din[18] din[19] din[20] din[21] din[22] din[23] din[24] din[25] din[26] din[27] din[28] din[29] din[30] din[31] din[32] din[33] din[34] din[35] din[36] din[37] din[38] din[39] din[40] din[41] din[42] din[43] din[44] din[45] din[46] din[47] din[48] din[49] din[50] din[51] din[52] din[53] din[54] din[55] din[56] din[57] din[58] din[59] din[60] din[61] din[62] din[63] din[64] din[65] din[66] din[67] din[68] din[69] din[70] din[71] din[72] din[73] din[74] din[75] din[76] din[77] din[78] din[79] din[80] din[81] din[82] din[83] din[84] din[85] din[86] din[87] din[88] din[89] din[90] din[91] din[92] din[93] din[94] din[95] din[96] din[97] din[98] din[99] din[100] din[101] din[102] din[103] din[104] din[105] din[106] din[107] din[108] din[109] din[110] din[111] din[112] din[113] din[114] din[115] din[116] din[117] din[118] din[119] din[120] din[121] din[122] din[123] din[124] din[125] din[126] din[127] dout[0] dout_bar[0] dout[1] dout_bar[1] dout[2] dout_bar[2] dout[3] dout_bar[3] dout[4] dout_bar[4] dout[5] dout_bar[5] dout[6] dout_bar[6] dout[7] dout_bar[7] dout[8] dout_bar[8] dout[9] dout_bar[9] dout[10] dout_bar[10] dout[11] dout_bar[11] dout[12] dout_bar[12] dout[13] dout_bar[13] dout[14] dout_bar[14] dout[15] dout_bar[15] dout[16] dout_bar[16] dout[17] dout_bar[17] dout[18] dout_bar[18] dout[19] dout_bar[19] dout[20] dout_bar[20] dout[21] dout_bar[21] dout[22] dout_bar[22] dout[23] dout_bar[23] dout[24] dout_bar[24] dout[25] dout_bar[25] dout[26] dout_bar[26] dout[27] dout_bar[27] dout[28] dout_bar[28] dout[29] dout_bar[29] dout[30] dout_bar[30] dout[31] dout_bar[31] dout[32] dout_bar[32] dout[33] dout_bar[33] dout[34] dout_bar[34] dout[35] dout_bar[35] dout[36] dout_bar[36] dout[37] dout_bar[37] dout[38] dout_bar[38] dout[39] dout_bar[39] dout[40] dout_bar[40] dout[41] dout_bar[41] dout[42] dout_bar[42] dout[43] dout_bar[43] dout[44] dout_bar[44] dout[45] dout_bar[45] dout[46] dout_bar[46] dout[47] dout_bar[47] dout[48] dout_bar[48] dout[49] dout_bar[49] dout[50] dout_bar[50] dout[51] dout_bar[51] dout[52] dout_bar[52] dout[53] dout_bar[53] dout[54] dout_bar[54] dout[55] dout_bar[55] dout[56] dout_bar[56] dout[57] dout_bar[57] dout[58] dout_bar[58] dout[59] dout_bar[59] dout[60] dout_bar[60] dout[61] dout_bar[61] dout[62] dout_bar[62] dout[63] dout_bar[63] dout[64] dout_bar[64] dout[65] dout_bar[65] dout[66] dout_bar[66] dout[67] dout_bar[67] dout[68] dout_bar[68] dout[69] dout_bar[69] dout[70] dout_bar[70] dout[71] dout_bar[71] dout[72] dout_bar[72] dout[73] dout_bar[73] dout[74] dout_bar[74] dout[75] dout_bar[75] dout[76] dout_bar[76] dout[77] dout_bar[77] dout[78] dout_bar[78] dout[79] dout_bar[79] dout[80] dout_bar[80] dout[81] dout_bar[81] dout[82] dout_bar[82] dout[83] dout_bar[83] dout[84] dout_bar[84] dout[85] dout_bar[85] dout[86] dout_bar[86] dout[87] dout_bar[87] dout[88] dout_bar[88] dout[89] dout_bar[89] dout[90] dout_bar[90] dout[91] dout_bar[91] dout[92] dout_bar[92] dout[93] dout_bar[93] dout[94] dout_bar[94] dout[95] dout_bar[95] dout[96] dout_bar[96] dout[97] dout_bar[97] dout[98] dout_bar[98] dout[99] dout_bar[99] dout[100] dout_bar[100] dout[101] dout_bar[101] dout[102] dout_bar[102] dout[103] dout_bar[103] dout[104] dout_bar[104] dout[105] dout_bar[105] dout[106] dout_bar[106] dout[107] dout_bar[107] dout[108] dout_bar[108] dout[109] dout_bar[109] dout[110] dout_bar[110] dout[111] dout_bar[111] dout[112] dout_bar[112] dout[113] dout_bar[113] dout[114] dout_bar[114] dout[115] dout_bar[115] dout[116] dout_bar[116] dout[117] dout_bar[117] dout[118] dout_bar[118] dout[119] dout_bar[119] dout[120] dout_bar[120] dout[121] dout_bar[121] dout[122] dout_bar[122] dout[123] dout_bar[123] dout[124] dout_bar[124] dout[125] dout_bar[125] dout[126] dout_bar[126] dout[127] dout_bar[127] clk vdd gnd
XXdff0 din[0] dout[0] dout_bar[0] clk vdd gnd ms_flop
XXdff2 din[1] dout[1] dout_bar[1] clk vdd gnd ms_flop
XXdff4 din[2] dout[2] dout_bar[2] clk vdd gnd ms_flop
XXdff6 din[3] dout[3] dout_bar[3] clk vdd gnd ms_flop
XXdff8 din[4] dout[4] dout_bar[4] clk vdd gnd ms_flop
XXdff10 din[5] dout[5] dout_bar[5] clk vdd gnd ms_flop
XXdff12 din[6] dout[6] dout_bar[6] clk vdd gnd ms_flop
XXdff14 din[7] dout[7] dout_bar[7] clk vdd gnd ms_flop
XXdff16 din[8] dout[8] dout_bar[8] clk vdd gnd ms_flop
XXdff18 din[9] dout[9] dout_bar[9] clk vdd gnd ms_flop
XXdff20 din[10] dout[10] dout_bar[10] clk vdd gnd ms_flop
XXdff22 din[11] dout[11] dout_bar[11] clk vdd gnd ms_flop
XXdff24 din[12] dout[12] dout_bar[12] clk vdd gnd ms_flop
XXdff26 din[13] dout[13] dout_bar[13] clk vdd gnd ms_flop
XXdff28 din[14] dout[14] dout_bar[14] clk vdd gnd ms_flop
XXdff30 din[15] dout[15] dout_bar[15] clk vdd gnd ms_flop
XXdff32 din[16] dout[16] dout_bar[16] clk vdd gnd ms_flop
XXdff34 din[17] dout[17] dout_bar[17] clk vdd gnd ms_flop
XXdff36 din[18] dout[18] dout_bar[18] clk vdd gnd ms_flop
XXdff38 din[19] dout[19] dout_bar[19] clk vdd gnd ms_flop
XXdff40 din[20] dout[20] dout_bar[20] clk vdd gnd ms_flop
XXdff42 din[21] dout[21] dout_bar[21] clk vdd gnd ms_flop
XXdff44 din[22] dout[22] dout_bar[22] clk vdd gnd ms_flop
XXdff46 din[23] dout[23] dout_bar[23] clk vdd gnd ms_flop
XXdff48 din[24] dout[24] dout_bar[24] clk vdd gnd ms_flop
XXdff50 din[25] dout[25] dout_bar[25] clk vdd gnd ms_flop
XXdff52 din[26] dout[26] dout_bar[26] clk vdd gnd ms_flop
XXdff54 din[27] dout[27] dout_bar[27] clk vdd gnd ms_flop
XXdff56 din[28] dout[28] dout_bar[28] clk vdd gnd ms_flop
XXdff58 din[29] dout[29] dout_bar[29] clk vdd gnd ms_flop
XXdff60 din[30] dout[30] dout_bar[30] clk vdd gnd ms_flop
XXdff62 din[31] dout[31] dout_bar[31] clk vdd gnd ms_flop
XXdff64 din[32] dout[32] dout_bar[32] clk vdd gnd ms_flop
XXdff66 din[33] dout[33] dout_bar[33] clk vdd gnd ms_flop
XXdff68 din[34] dout[34] dout_bar[34] clk vdd gnd ms_flop
XXdff70 din[35] dout[35] dout_bar[35] clk vdd gnd ms_flop
XXdff72 din[36] dout[36] dout_bar[36] clk vdd gnd ms_flop
XXdff74 din[37] dout[37] dout_bar[37] clk vdd gnd ms_flop
XXdff76 din[38] dout[38] dout_bar[38] clk vdd gnd ms_flop
XXdff78 din[39] dout[39] dout_bar[39] clk vdd gnd ms_flop
XXdff80 din[40] dout[40] dout_bar[40] clk vdd gnd ms_flop
XXdff82 din[41] dout[41] dout_bar[41] clk vdd gnd ms_flop
XXdff84 din[42] dout[42] dout_bar[42] clk vdd gnd ms_flop
XXdff86 din[43] dout[43] dout_bar[43] clk vdd gnd ms_flop
XXdff88 din[44] dout[44] dout_bar[44] clk vdd gnd ms_flop
XXdff90 din[45] dout[45] dout_bar[45] clk vdd gnd ms_flop
XXdff92 din[46] dout[46] dout_bar[46] clk vdd gnd ms_flop
XXdff94 din[47] dout[47] dout_bar[47] clk vdd gnd ms_flop
XXdff96 din[48] dout[48] dout_bar[48] clk vdd gnd ms_flop
XXdff98 din[49] dout[49] dout_bar[49] clk vdd gnd ms_flop
XXdff100 din[50] dout[50] dout_bar[50] clk vdd gnd ms_flop
XXdff102 din[51] dout[51] dout_bar[51] clk vdd gnd ms_flop
XXdff104 din[52] dout[52] dout_bar[52] clk vdd gnd ms_flop
XXdff106 din[53] dout[53] dout_bar[53] clk vdd gnd ms_flop
XXdff108 din[54] dout[54] dout_bar[54] clk vdd gnd ms_flop
XXdff110 din[55] dout[55] dout_bar[55] clk vdd gnd ms_flop
XXdff112 din[56] dout[56] dout_bar[56] clk vdd gnd ms_flop
XXdff114 din[57] dout[57] dout_bar[57] clk vdd gnd ms_flop
XXdff116 din[58] dout[58] dout_bar[58] clk vdd gnd ms_flop
XXdff118 din[59] dout[59] dout_bar[59] clk vdd gnd ms_flop
XXdff120 din[60] dout[60] dout_bar[60] clk vdd gnd ms_flop
XXdff122 din[61] dout[61] dout_bar[61] clk vdd gnd ms_flop
XXdff124 din[62] dout[62] dout_bar[62] clk vdd gnd ms_flop
XXdff126 din[63] dout[63] dout_bar[63] clk vdd gnd ms_flop
XXdff128 din[64] dout[64] dout_bar[64] clk vdd gnd ms_flop
XXdff130 din[65] dout[65] dout_bar[65] clk vdd gnd ms_flop
XXdff132 din[66] dout[66] dout_bar[66] clk vdd gnd ms_flop
XXdff134 din[67] dout[67] dout_bar[67] clk vdd gnd ms_flop
XXdff136 din[68] dout[68] dout_bar[68] clk vdd gnd ms_flop
XXdff138 din[69] dout[69] dout_bar[69] clk vdd gnd ms_flop
XXdff140 din[70] dout[70] dout_bar[70] clk vdd gnd ms_flop
XXdff142 din[71] dout[71] dout_bar[71] clk vdd gnd ms_flop
XXdff144 din[72] dout[72] dout_bar[72] clk vdd gnd ms_flop
XXdff146 din[73] dout[73] dout_bar[73] clk vdd gnd ms_flop
XXdff148 din[74] dout[74] dout_bar[74] clk vdd gnd ms_flop
XXdff150 din[75] dout[75] dout_bar[75] clk vdd gnd ms_flop
XXdff152 din[76] dout[76] dout_bar[76] clk vdd gnd ms_flop
XXdff154 din[77] dout[77] dout_bar[77] clk vdd gnd ms_flop
XXdff156 din[78] dout[78] dout_bar[78] clk vdd gnd ms_flop
XXdff158 din[79] dout[79] dout_bar[79] clk vdd gnd ms_flop
XXdff160 din[80] dout[80] dout_bar[80] clk vdd gnd ms_flop
XXdff162 din[81] dout[81] dout_bar[81] clk vdd gnd ms_flop
XXdff164 din[82] dout[82] dout_bar[82] clk vdd gnd ms_flop
XXdff166 din[83] dout[83] dout_bar[83] clk vdd gnd ms_flop
XXdff168 din[84] dout[84] dout_bar[84] clk vdd gnd ms_flop
XXdff170 din[85] dout[85] dout_bar[85] clk vdd gnd ms_flop
XXdff172 din[86] dout[86] dout_bar[86] clk vdd gnd ms_flop
XXdff174 din[87] dout[87] dout_bar[87] clk vdd gnd ms_flop
XXdff176 din[88] dout[88] dout_bar[88] clk vdd gnd ms_flop
XXdff178 din[89] dout[89] dout_bar[89] clk vdd gnd ms_flop
XXdff180 din[90] dout[90] dout_bar[90] clk vdd gnd ms_flop
XXdff182 din[91] dout[91] dout_bar[91] clk vdd gnd ms_flop
XXdff184 din[92] dout[92] dout_bar[92] clk vdd gnd ms_flop
XXdff186 din[93] dout[93] dout_bar[93] clk vdd gnd ms_flop
XXdff188 din[94] dout[94] dout_bar[94] clk vdd gnd ms_flop
XXdff190 din[95] dout[95] dout_bar[95] clk vdd gnd ms_flop
XXdff192 din[96] dout[96] dout_bar[96] clk vdd gnd ms_flop
XXdff194 din[97] dout[97] dout_bar[97] clk vdd gnd ms_flop
XXdff196 din[98] dout[98] dout_bar[98] clk vdd gnd ms_flop
XXdff198 din[99] dout[99] dout_bar[99] clk vdd gnd ms_flop
XXdff200 din[100] dout[100] dout_bar[100] clk vdd gnd ms_flop
XXdff202 din[101] dout[101] dout_bar[101] clk vdd gnd ms_flop
XXdff204 din[102] dout[102] dout_bar[102] clk vdd gnd ms_flop
XXdff206 din[103] dout[103] dout_bar[103] clk vdd gnd ms_flop
XXdff208 din[104] dout[104] dout_bar[104] clk vdd gnd ms_flop
XXdff210 din[105] dout[105] dout_bar[105] clk vdd gnd ms_flop
XXdff212 din[106] dout[106] dout_bar[106] clk vdd gnd ms_flop
XXdff214 din[107] dout[107] dout_bar[107] clk vdd gnd ms_flop
XXdff216 din[108] dout[108] dout_bar[108] clk vdd gnd ms_flop
XXdff218 din[109] dout[109] dout_bar[109] clk vdd gnd ms_flop
XXdff220 din[110] dout[110] dout_bar[110] clk vdd gnd ms_flop
XXdff222 din[111] dout[111] dout_bar[111] clk vdd gnd ms_flop
XXdff224 din[112] dout[112] dout_bar[112] clk vdd gnd ms_flop
XXdff226 din[113] dout[113] dout_bar[113] clk vdd gnd ms_flop
XXdff228 din[114] dout[114] dout_bar[114] clk vdd gnd ms_flop
XXdff230 din[115] dout[115] dout_bar[115] clk vdd gnd ms_flop
XXdff232 din[116] dout[116] dout_bar[116] clk vdd gnd ms_flop
XXdff234 din[117] dout[117] dout_bar[117] clk vdd gnd ms_flop
XXdff236 din[118] dout[118] dout_bar[118] clk vdd gnd ms_flop
XXdff238 din[119] dout[119] dout_bar[119] clk vdd gnd ms_flop
XXdff240 din[120] dout[120] dout_bar[120] clk vdd gnd ms_flop
XXdff242 din[121] dout[121] dout_bar[121] clk vdd gnd ms_flop
XXdff244 din[122] dout[122] dout_bar[122] clk vdd gnd ms_flop
XXdff246 din[123] dout[123] dout_bar[123] clk vdd gnd ms_flop
XXdff248 din[124] dout[124] dout_bar[124] clk vdd gnd ms_flop
XXdff250 din[125] dout[125] dout_bar[125] clk vdd gnd ms_flop
XXdff252 din[126] dout[126] dout_bar[126] clk vdd gnd ms_flop
XXdff254 din[127] dout[127] dout_bar[127] clk vdd gnd ms_flop
.ENDS msf_data_in
*********************** tri_gate ******************************

.SUBCKT tri_gate in out en en_bar vdd gnd

M_1 net_2 in_inv gnd gnd n W='1.2*1u' L=0.6u
M_2 net_3 in_inv vdd vdd p W='2.4*1u' L=0.6u
M_3 out en_bar net_3 vdd p W='2.4*1u' L=0.6u
M_4 out en net_2 gnd n W='1.2*1u' L=0.6u
M_5 in_inv in vdd vdd p W='2.4*1u' L=0.6u
M_6 in_inv in gnd gnd n W='1.2*1u' L=0.6u


.ENDS	

.SUBCKT tri_gate_array in[0] in[1] in[2] in[3] in[4] in[5] in[6] in[7] in[8] in[9] in[10] in[11] in[12] in[13] in[14] in[15] in[16] in[17] in[18] in[19] in[20] in[21] in[22] in[23] in[24] in[25] in[26] in[27] in[28] in[29] in[30] in[31] in[32] in[33] in[34] in[35] in[36] in[37] in[38] in[39] in[40] in[41] in[42] in[43] in[44] in[45] in[46] in[47] in[48] in[49] in[50] in[51] in[52] in[53] in[54] in[55] in[56] in[57] in[58] in[59] in[60] in[61] in[62] in[63] in[64] in[65] in[66] in[67] in[68] in[69] in[70] in[71] in[72] in[73] in[74] in[75] in[76] in[77] in[78] in[79] in[80] in[81] in[82] in[83] in[84] in[85] in[86] in[87] in[88] in[89] in[90] in[91] in[92] in[93] in[94] in[95] in[96] in[97] in[98] in[99] in[100] in[101] in[102] in[103] in[104] in[105] in[106] in[107] in[108] in[109] in[110] in[111] in[112] in[113] in[114] in[115] in[116] in[117] in[118] in[119] in[120] in[121] in[122] in[123] in[124] in[125] in[126] in[127] out[0] out[1] out[2] out[3] out[4] out[5] out[6] out[7] out[8] out[9] out[10] out[11] out[12] out[13] out[14] out[15] out[16] out[17] out[18] out[19] out[20] out[21] out[22] out[23] out[24] out[25] out[26] out[27] out[28] out[29] out[30] out[31] out[32] out[33] out[34] out[35] out[36] out[37] out[38] out[39] out[40] out[41] out[42] out[43] out[44] out[45] out[46] out[47] out[48] out[49] out[50] out[51] out[52] out[53] out[54] out[55] out[56] out[57] out[58] out[59] out[60] out[61] out[62] out[63] out[64] out[65] out[66] out[67] out[68] out[69] out[70] out[71] out[72] out[73] out[74] out[75] out[76] out[77] out[78] out[79] out[80] out[81] out[82] out[83] out[84] out[85] out[86] out[87] out[88] out[89] out[90] out[91] out[92] out[93] out[94] out[95] out[96] out[97] out[98] out[99] out[100] out[101] out[102] out[103] out[104] out[105] out[106] out[107] out[108] out[109] out[110] out[111] out[112] out[113] out[114] out[115] out[116] out[117] out[118] out[119] out[120] out[121] out[122] out[123] out[124] out[125] out[126] out[127] en en_bar vdd gnd
XXtri_gate0 in[0] out[0] en en_bar vdd gnd tri_gate
XXtri_gate2 in[1] out[1] en en_bar vdd gnd tri_gate
XXtri_gate4 in[2] out[2] en en_bar vdd gnd tri_gate
XXtri_gate6 in[3] out[3] en en_bar vdd gnd tri_gate
XXtri_gate8 in[4] out[4] en en_bar vdd gnd tri_gate
XXtri_gate10 in[5] out[5] en en_bar vdd gnd tri_gate
XXtri_gate12 in[6] out[6] en en_bar vdd gnd tri_gate
XXtri_gate14 in[7] out[7] en en_bar vdd gnd tri_gate
XXtri_gate16 in[8] out[8] en en_bar vdd gnd tri_gate
XXtri_gate18 in[9] out[9] en en_bar vdd gnd tri_gate
XXtri_gate20 in[10] out[10] en en_bar vdd gnd tri_gate
XXtri_gate22 in[11] out[11] en en_bar vdd gnd tri_gate
XXtri_gate24 in[12] out[12] en en_bar vdd gnd tri_gate
XXtri_gate26 in[13] out[13] en en_bar vdd gnd tri_gate
XXtri_gate28 in[14] out[14] en en_bar vdd gnd tri_gate
XXtri_gate30 in[15] out[15] en en_bar vdd gnd tri_gate
XXtri_gate32 in[16] out[16] en en_bar vdd gnd tri_gate
XXtri_gate34 in[17] out[17] en en_bar vdd gnd tri_gate
XXtri_gate36 in[18] out[18] en en_bar vdd gnd tri_gate
XXtri_gate38 in[19] out[19] en en_bar vdd gnd tri_gate
XXtri_gate40 in[20] out[20] en en_bar vdd gnd tri_gate
XXtri_gate42 in[21] out[21] en en_bar vdd gnd tri_gate
XXtri_gate44 in[22] out[22] en en_bar vdd gnd tri_gate
XXtri_gate46 in[23] out[23] en en_bar vdd gnd tri_gate
XXtri_gate48 in[24] out[24] en en_bar vdd gnd tri_gate
XXtri_gate50 in[25] out[25] en en_bar vdd gnd tri_gate
XXtri_gate52 in[26] out[26] en en_bar vdd gnd tri_gate
XXtri_gate54 in[27] out[27] en en_bar vdd gnd tri_gate
XXtri_gate56 in[28] out[28] en en_bar vdd gnd tri_gate
XXtri_gate58 in[29] out[29] en en_bar vdd gnd tri_gate
XXtri_gate60 in[30] out[30] en en_bar vdd gnd tri_gate
XXtri_gate62 in[31] out[31] en en_bar vdd gnd tri_gate
XXtri_gate64 in[32] out[32] en en_bar vdd gnd tri_gate
XXtri_gate66 in[33] out[33] en en_bar vdd gnd tri_gate
XXtri_gate68 in[34] out[34] en en_bar vdd gnd tri_gate
XXtri_gate70 in[35] out[35] en en_bar vdd gnd tri_gate
XXtri_gate72 in[36] out[36] en en_bar vdd gnd tri_gate
XXtri_gate74 in[37] out[37] en en_bar vdd gnd tri_gate
XXtri_gate76 in[38] out[38] en en_bar vdd gnd tri_gate
XXtri_gate78 in[39] out[39] en en_bar vdd gnd tri_gate
XXtri_gate80 in[40] out[40] en en_bar vdd gnd tri_gate
XXtri_gate82 in[41] out[41] en en_bar vdd gnd tri_gate
XXtri_gate84 in[42] out[42] en en_bar vdd gnd tri_gate
XXtri_gate86 in[43] out[43] en en_bar vdd gnd tri_gate
XXtri_gate88 in[44] out[44] en en_bar vdd gnd tri_gate
XXtri_gate90 in[45] out[45] en en_bar vdd gnd tri_gate
XXtri_gate92 in[46] out[46] en en_bar vdd gnd tri_gate
XXtri_gate94 in[47] out[47] en en_bar vdd gnd tri_gate
XXtri_gate96 in[48] out[48] en en_bar vdd gnd tri_gate
XXtri_gate98 in[49] out[49] en en_bar vdd gnd tri_gate
XXtri_gate100 in[50] out[50] en en_bar vdd gnd tri_gate
XXtri_gate102 in[51] out[51] en en_bar vdd gnd tri_gate
XXtri_gate104 in[52] out[52] en en_bar vdd gnd tri_gate
XXtri_gate106 in[53] out[53] en en_bar vdd gnd tri_gate
XXtri_gate108 in[54] out[54] en en_bar vdd gnd tri_gate
XXtri_gate110 in[55] out[55] en en_bar vdd gnd tri_gate
XXtri_gate112 in[56] out[56] en en_bar vdd gnd tri_gate
XXtri_gate114 in[57] out[57] en en_bar vdd gnd tri_gate
XXtri_gate116 in[58] out[58] en en_bar vdd gnd tri_gate
XXtri_gate118 in[59] out[59] en en_bar vdd gnd tri_gate
XXtri_gate120 in[60] out[60] en en_bar vdd gnd tri_gate
XXtri_gate122 in[61] out[61] en en_bar vdd gnd tri_gate
XXtri_gate124 in[62] out[62] en en_bar vdd gnd tri_gate
XXtri_gate126 in[63] out[63] en en_bar vdd gnd tri_gate
XXtri_gate128 in[64] out[64] en en_bar vdd gnd tri_gate
XXtri_gate130 in[65] out[65] en en_bar vdd gnd tri_gate
XXtri_gate132 in[66] out[66] en en_bar vdd gnd tri_gate
XXtri_gate134 in[67] out[67] en en_bar vdd gnd tri_gate
XXtri_gate136 in[68] out[68] en en_bar vdd gnd tri_gate
XXtri_gate138 in[69] out[69] en en_bar vdd gnd tri_gate
XXtri_gate140 in[70] out[70] en en_bar vdd gnd tri_gate
XXtri_gate142 in[71] out[71] en en_bar vdd gnd tri_gate
XXtri_gate144 in[72] out[72] en en_bar vdd gnd tri_gate
XXtri_gate146 in[73] out[73] en en_bar vdd gnd tri_gate
XXtri_gate148 in[74] out[74] en en_bar vdd gnd tri_gate
XXtri_gate150 in[75] out[75] en en_bar vdd gnd tri_gate
XXtri_gate152 in[76] out[76] en en_bar vdd gnd tri_gate
XXtri_gate154 in[77] out[77] en en_bar vdd gnd tri_gate
XXtri_gate156 in[78] out[78] en en_bar vdd gnd tri_gate
XXtri_gate158 in[79] out[79] en en_bar vdd gnd tri_gate
XXtri_gate160 in[80] out[80] en en_bar vdd gnd tri_gate
XXtri_gate162 in[81] out[81] en en_bar vdd gnd tri_gate
XXtri_gate164 in[82] out[82] en en_bar vdd gnd tri_gate
XXtri_gate166 in[83] out[83] en en_bar vdd gnd tri_gate
XXtri_gate168 in[84] out[84] en en_bar vdd gnd tri_gate
XXtri_gate170 in[85] out[85] en en_bar vdd gnd tri_gate
XXtri_gate172 in[86] out[86] en en_bar vdd gnd tri_gate
XXtri_gate174 in[87] out[87] en en_bar vdd gnd tri_gate
XXtri_gate176 in[88] out[88] en en_bar vdd gnd tri_gate
XXtri_gate178 in[89] out[89] en en_bar vdd gnd tri_gate
XXtri_gate180 in[90] out[90] en en_bar vdd gnd tri_gate
XXtri_gate182 in[91] out[91] en en_bar vdd gnd tri_gate
XXtri_gate184 in[92] out[92] en en_bar vdd gnd tri_gate
XXtri_gate186 in[93] out[93] en en_bar vdd gnd tri_gate
XXtri_gate188 in[94] out[94] en en_bar vdd gnd tri_gate
XXtri_gate190 in[95] out[95] en en_bar vdd gnd tri_gate
XXtri_gate192 in[96] out[96] en en_bar vdd gnd tri_gate
XXtri_gate194 in[97] out[97] en en_bar vdd gnd tri_gate
XXtri_gate196 in[98] out[98] en en_bar vdd gnd tri_gate
XXtri_gate198 in[99] out[99] en en_bar vdd gnd tri_gate
XXtri_gate200 in[100] out[100] en en_bar vdd gnd tri_gate
XXtri_gate202 in[101] out[101] en en_bar vdd gnd tri_gate
XXtri_gate204 in[102] out[102] en en_bar vdd gnd tri_gate
XXtri_gate206 in[103] out[103] en en_bar vdd gnd tri_gate
XXtri_gate208 in[104] out[104] en en_bar vdd gnd tri_gate
XXtri_gate210 in[105] out[105] en en_bar vdd gnd tri_gate
XXtri_gate212 in[106] out[106] en en_bar vdd gnd tri_gate
XXtri_gate214 in[107] out[107] en en_bar vdd gnd tri_gate
XXtri_gate216 in[108] out[108] en en_bar vdd gnd tri_gate
XXtri_gate218 in[109] out[109] en en_bar vdd gnd tri_gate
XXtri_gate220 in[110] out[110] en en_bar vdd gnd tri_gate
XXtri_gate222 in[111] out[111] en en_bar vdd gnd tri_gate
XXtri_gate224 in[112] out[112] en en_bar vdd gnd tri_gate
XXtri_gate226 in[113] out[113] en en_bar vdd gnd tri_gate
XXtri_gate228 in[114] out[114] en en_bar vdd gnd tri_gate
XXtri_gate230 in[115] out[115] en en_bar vdd gnd tri_gate
XXtri_gate232 in[116] out[116] en en_bar vdd gnd tri_gate
XXtri_gate234 in[117] out[117] en en_bar vdd gnd tri_gate
XXtri_gate236 in[118] out[118] en en_bar vdd gnd tri_gate
XXtri_gate238 in[119] out[119] en en_bar vdd gnd tri_gate
XXtri_gate240 in[120] out[120] en en_bar vdd gnd tri_gate
XXtri_gate242 in[121] out[121] en en_bar vdd gnd tri_gate
XXtri_gate244 in[122] out[122] en en_bar vdd gnd tri_gate
XXtri_gate246 in[123] out[123] en en_bar vdd gnd tri_gate
XXtri_gate248 in[124] out[124] en en_bar vdd gnd tri_gate
XXtri_gate250 in[125] out[125] en en_bar vdd gnd tri_gate
XXtri_gate252 in[126] out[126] en en_bar vdd gnd tri_gate
XXtri_gate254 in[127] out[127] en en_bar vdd gnd tri_gate
.ENDS tri_gate_array

.SUBCKT pinv_11 A Z vdd gnd
Mpinv_pmos Z A vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpinv_nmos Z A gnd gnd n m=1 w=1.2u l=0.6u pd=3.6u ps=3.6u as=1.8p ad=1.8p
.ENDS pinv_11

.SUBCKT pinv_12 A Z vdd gnd
Mpinv_pmos Z A vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpinv_nmos Z A gnd gnd n m=1 w=1.2u l=0.6u pd=3.6u ps=3.6u as=1.8p ad=1.8p
.ENDS pinv_12

.SUBCKT pnand2_4 A B Z vdd gnd
Mpnand2_pmos1 vdd A Z vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand2_pmos2 Z B vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand2_nmos1 Z B net1 gnd n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand2_nmos2 net1 A gnd gnd n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
.ENDS pnand2_4

.SUBCKT wordline_driver in[0] in[1] in[2] in[3] in[4] in[5] in[6] in[7] in[8] in[9] in[10] in[11] in[12] in[13] in[14] in[15] in[16] in[17] in[18] in[19] in[20] in[21] in[22] in[23] in[24] in[25] in[26] in[27] in[28] in[29] in[30] in[31] in[32] in[33] in[34] in[35] in[36] in[37] in[38] in[39] in[40] in[41] in[42] in[43] in[44] in[45] in[46] in[47] in[48] in[49] in[50] in[51] in[52] in[53] in[54] in[55] in[56] in[57] in[58] in[59] in[60] in[61] in[62] in[63] in[64] in[65] in[66] in[67] in[68] in[69] in[70] in[71] in[72] in[73] in[74] in[75] in[76] in[77] in[78] in[79] in[80] in[81] in[82] in[83] in[84] in[85] in[86] in[87] in[88] in[89] in[90] in[91] in[92] in[93] in[94] in[95] in[96] in[97] in[98] in[99] in[100] in[101] in[102] in[103] in[104] in[105] in[106] in[107] in[108] in[109] in[110] in[111] in[112] in[113] in[114] in[115] in[116] in[117] in[118] in[119] in[120] in[121] in[122] in[123] in[124] in[125] in[126] in[127] in[128] in[129] in[130] in[131] in[132] in[133] in[134] in[135] in[136] in[137] in[138] in[139] in[140] in[141] in[142] in[143] in[144] in[145] in[146] in[147] in[148] in[149] in[150] in[151] in[152] in[153] in[154] in[155] in[156] in[157] in[158] in[159] in[160] in[161] in[162] in[163] in[164] in[165] in[166] in[167] in[168] in[169] in[170] in[171] in[172] in[173] in[174] in[175] in[176] in[177] in[178] in[179] in[180] in[181] in[182] in[183] in[184] in[185] in[186] in[187] in[188] in[189] in[190] in[191] in[192] in[193] in[194] in[195] in[196] in[197] in[198] in[199] in[200] in[201] in[202] in[203] in[204] in[205] in[206] in[207] in[208] in[209] in[210] in[211] in[212] in[213] in[214] in[215] in[216] in[217] in[218] in[219] in[220] in[221] in[222] in[223] in[224] in[225] in[226] in[227] in[228] in[229] in[230] in[231] in[232] in[233] in[234] in[235] in[236] in[237] in[238] in[239] in[240] in[241] in[242] in[243] in[244] in[245] in[246] in[247] in[248] in[249] in[250] in[251] in[252] in[253] in[254] in[255] wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] wl[128] wl[129] wl[130] wl[131] wl[132] wl[133] wl[134] wl[135] wl[136] wl[137] wl[138] wl[139] wl[140] wl[141] wl[142] wl[143] wl[144] wl[145] wl[146] wl[147] wl[148] wl[149] wl[150] wl[151] wl[152] wl[153] wl[154] wl[155] wl[156] wl[157] wl[158] wl[159] wl[160] wl[161] wl[162] wl[163] wl[164] wl[165] wl[166] wl[167] wl[168] wl[169] wl[170] wl[171] wl[172] wl[173] wl[174] wl[175] wl[176] wl[177] wl[178] wl[179] wl[180] wl[181] wl[182] wl[183] wl[184] wl[185] wl[186] wl[187] wl[188] wl[189] wl[190] wl[191] wl[192] wl[193] wl[194] wl[195] wl[196] wl[197] wl[198] wl[199] wl[200] wl[201] wl[202] wl[203] wl[204] wl[205] wl[206] wl[207] wl[208] wl[209] wl[210] wl[211] wl[212] wl[213] wl[214] wl[215] wl[216] wl[217] wl[218] wl[219] wl[220] wl[221] wl[222] wl[223] wl[224] wl[225] wl[226] wl[227] wl[228] wl[229] wl[230] wl[231] wl[232] wl[233] wl[234] wl[235] wl[236] wl[237] wl[238] wl[239] wl[240] wl[241] wl[242] wl[243] wl[244] wl[245] wl[246] wl[247] wl[248] wl[249] wl[250] wl[251] wl[252] wl[253] wl[254] wl[255] en vdd gnd
Xwl_driver_inv_en0 en en_bar[0] vdd gnd pinv_12
Xwl_driver_nand0 en_bar[0] in[0] net[0] vdd gnd pnand2_4
Xwl_driver_inv0 net[0] wl[0] vdd gnd pinv_11
Xwl_driver_inv_en1 en en_bar[1] vdd gnd pinv_12
Xwl_driver_nand1 en_bar[1] in[1] net[1] vdd gnd pnand2_4
Xwl_driver_inv1 net[1] wl[1] vdd gnd pinv_11
Xwl_driver_inv_en2 en en_bar[2] vdd gnd pinv_12
Xwl_driver_nand2 en_bar[2] in[2] net[2] vdd gnd pnand2_4
Xwl_driver_inv2 net[2] wl[2] vdd gnd pinv_11
Xwl_driver_inv_en3 en en_bar[3] vdd gnd pinv_12
Xwl_driver_nand3 en_bar[3] in[3] net[3] vdd gnd pnand2_4
Xwl_driver_inv3 net[3] wl[3] vdd gnd pinv_11
Xwl_driver_inv_en4 en en_bar[4] vdd gnd pinv_12
Xwl_driver_nand4 en_bar[4] in[4] net[4] vdd gnd pnand2_4
Xwl_driver_inv4 net[4] wl[4] vdd gnd pinv_11
Xwl_driver_inv_en5 en en_bar[5] vdd gnd pinv_12
Xwl_driver_nand5 en_bar[5] in[5] net[5] vdd gnd pnand2_4
Xwl_driver_inv5 net[5] wl[5] vdd gnd pinv_11
Xwl_driver_inv_en6 en en_bar[6] vdd gnd pinv_12
Xwl_driver_nand6 en_bar[6] in[6] net[6] vdd gnd pnand2_4
Xwl_driver_inv6 net[6] wl[6] vdd gnd pinv_11
Xwl_driver_inv_en7 en en_bar[7] vdd gnd pinv_12
Xwl_driver_nand7 en_bar[7] in[7] net[7] vdd gnd pnand2_4
Xwl_driver_inv7 net[7] wl[7] vdd gnd pinv_11
Xwl_driver_inv_en8 en en_bar[8] vdd gnd pinv_12
Xwl_driver_nand8 en_bar[8] in[8] net[8] vdd gnd pnand2_4
Xwl_driver_inv8 net[8] wl[8] vdd gnd pinv_11
Xwl_driver_inv_en9 en en_bar[9] vdd gnd pinv_12
Xwl_driver_nand9 en_bar[9] in[9] net[9] vdd gnd pnand2_4
Xwl_driver_inv9 net[9] wl[9] vdd gnd pinv_11
Xwl_driver_inv_en10 en en_bar[10] vdd gnd pinv_12
Xwl_driver_nand10 en_bar[10] in[10] net[10] vdd gnd pnand2_4
Xwl_driver_inv10 net[10] wl[10] vdd gnd pinv_11
Xwl_driver_inv_en11 en en_bar[11] vdd gnd pinv_12
Xwl_driver_nand11 en_bar[11] in[11] net[11] vdd gnd pnand2_4
Xwl_driver_inv11 net[11] wl[11] vdd gnd pinv_11
Xwl_driver_inv_en12 en en_bar[12] vdd gnd pinv_12
Xwl_driver_nand12 en_bar[12] in[12] net[12] vdd gnd pnand2_4
Xwl_driver_inv12 net[12] wl[12] vdd gnd pinv_11
Xwl_driver_inv_en13 en en_bar[13] vdd gnd pinv_12
Xwl_driver_nand13 en_bar[13] in[13] net[13] vdd gnd pnand2_4
Xwl_driver_inv13 net[13] wl[13] vdd gnd pinv_11
Xwl_driver_inv_en14 en en_bar[14] vdd gnd pinv_12
Xwl_driver_nand14 en_bar[14] in[14] net[14] vdd gnd pnand2_4
Xwl_driver_inv14 net[14] wl[14] vdd gnd pinv_11
Xwl_driver_inv_en15 en en_bar[15] vdd gnd pinv_12
Xwl_driver_nand15 en_bar[15] in[15] net[15] vdd gnd pnand2_4
Xwl_driver_inv15 net[15] wl[15] vdd gnd pinv_11
Xwl_driver_inv_en16 en en_bar[16] vdd gnd pinv_12
Xwl_driver_nand16 en_bar[16] in[16] net[16] vdd gnd pnand2_4
Xwl_driver_inv16 net[16] wl[16] vdd gnd pinv_11
Xwl_driver_inv_en17 en en_bar[17] vdd gnd pinv_12
Xwl_driver_nand17 en_bar[17] in[17] net[17] vdd gnd pnand2_4
Xwl_driver_inv17 net[17] wl[17] vdd gnd pinv_11
Xwl_driver_inv_en18 en en_bar[18] vdd gnd pinv_12
Xwl_driver_nand18 en_bar[18] in[18] net[18] vdd gnd pnand2_4
Xwl_driver_inv18 net[18] wl[18] vdd gnd pinv_11
Xwl_driver_inv_en19 en en_bar[19] vdd gnd pinv_12
Xwl_driver_nand19 en_bar[19] in[19] net[19] vdd gnd pnand2_4
Xwl_driver_inv19 net[19] wl[19] vdd gnd pinv_11
Xwl_driver_inv_en20 en en_bar[20] vdd gnd pinv_12
Xwl_driver_nand20 en_bar[20] in[20] net[20] vdd gnd pnand2_4
Xwl_driver_inv20 net[20] wl[20] vdd gnd pinv_11
Xwl_driver_inv_en21 en en_bar[21] vdd gnd pinv_12
Xwl_driver_nand21 en_bar[21] in[21] net[21] vdd gnd pnand2_4
Xwl_driver_inv21 net[21] wl[21] vdd gnd pinv_11
Xwl_driver_inv_en22 en en_bar[22] vdd gnd pinv_12
Xwl_driver_nand22 en_bar[22] in[22] net[22] vdd gnd pnand2_4
Xwl_driver_inv22 net[22] wl[22] vdd gnd pinv_11
Xwl_driver_inv_en23 en en_bar[23] vdd gnd pinv_12
Xwl_driver_nand23 en_bar[23] in[23] net[23] vdd gnd pnand2_4
Xwl_driver_inv23 net[23] wl[23] vdd gnd pinv_11
Xwl_driver_inv_en24 en en_bar[24] vdd gnd pinv_12
Xwl_driver_nand24 en_bar[24] in[24] net[24] vdd gnd pnand2_4
Xwl_driver_inv24 net[24] wl[24] vdd gnd pinv_11
Xwl_driver_inv_en25 en en_bar[25] vdd gnd pinv_12
Xwl_driver_nand25 en_bar[25] in[25] net[25] vdd gnd pnand2_4
Xwl_driver_inv25 net[25] wl[25] vdd gnd pinv_11
Xwl_driver_inv_en26 en en_bar[26] vdd gnd pinv_12
Xwl_driver_nand26 en_bar[26] in[26] net[26] vdd gnd pnand2_4
Xwl_driver_inv26 net[26] wl[26] vdd gnd pinv_11
Xwl_driver_inv_en27 en en_bar[27] vdd gnd pinv_12
Xwl_driver_nand27 en_bar[27] in[27] net[27] vdd gnd pnand2_4
Xwl_driver_inv27 net[27] wl[27] vdd gnd pinv_11
Xwl_driver_inv_en28 en en_bar[28] vdd gnd pinv_12
Xwl_driver_nand28 en_bar[28] in[28] net[28] vdd gnd pnand2_4
Xwl_driver_inv28 net[28] wl[28] vdd gnd pinv_11
Xwl_driver_inv_en29 en en_bar[29] vdd gnd pinv_12
Xwl_driver_nand29 en_bar[29] in[29] net[29] vdd gnd pnand2_4
Xwl_driver_inv29 net[29] wl[29] vdd gnd pinv_11
Xwl_driver_inv_en30 en en_bar[30] vdd gnd pinv_12
Xwl_driver_nand30 en_bar[30] in[30] net[30] vdd gnd pnand2_4
Xwl_driver_inv30 net[30] wl[30] vdd gnd pinv_11
Xwl_driver_inv_en31 en en_bar[31] vdd gnd pinv_12
Xwl_driver_nand31 en_bar[31] in[31] net[31] vdd gnd pnand2_4
Xwl_driver_inv31 net[31] wl[31] vdd gnd pinv_11
Xwl_driver_inv_en32 en en_bar[32] vdd gnd pinv_12
Xwl_driver_nand32 en_bar[32] in[32] net[32] vdd gnd pnand2_4
Xwl_driver_inv32 net[32] wl[32] vdd gnd pinv_11
Xwl_driver_inv_en33 en en_bar[33] vdd gnd pinv_12
Xwl_driver_nand33 en_bar[33] in[33] net[33] vdd gnd pnand2_4
Xwl_driver_inv33 net[33] wl[33] vdd gnd pinv_11
Xwl_driver_inv_en34 en en_bar[34] vdd gnd pinv_12
Xwl_driver_nand34 en_bar[34] in[34] net[34] vdd gnd pnand2_4
Xwl_driver_inv34 net[34] wl[34] vdd gnd pinv_11
Xwl_driver_inv_en35 en en_bar[35] vdd gnd pinv_12
Xwl_driver_nand35 en_bar[35] in[35] net[35] vdd gnd pnand2_4
Xwl_driver_inv35 net[35] wl[35] vdd gnd pinv_11
Xwl_driver_inv_en36 en en_bar[36] vdd gnd pinv_12
Xwl_driver_nand36 en_bar[36] in[36] net[36] vdd gnd pnand2_4
Xwl_driver_inv36 net[36] wl[36] vdd gnd pinv_11
Xwl_driver_inv_en37 en en_bar[37] vdd gnd pinv_12
Xwl_driver_nand37 en_bar[37] in[37] net[37] vdd gnd pnand2_4
Xwl_driver_inv37 net[37] wl[37] vdd gnd pinv_11
Xwl_driver_inv_en38 en en_bar[38] vdd gnd pinv_12
Xwl_driver_nand38 en_bar[38] in[38] net[38] vdd gnd pnand2_4
Xwl_driver_inv38 net[38] wl[38] vdd gnd pinv_11
Xwl_driver_inv_en39 en en_bar[39] vdd gnd pinv_12
Xwl_driver_nand39 en_bar[39] in[39] net[39] vdd gnd pnand2_4
Xwl_driver_inv39 net[39] wl[39] vdd gnd pinv_11
Xwl_driver_inv_en40 en en_bar[40] vdd gnd pinv_12
Xwl_driver_nand40 en_bar[40] in[40] net[40] vdd gnd pnand2_4
Xwl_driver_inv40 net[40] wl[40] vdd gnd pinv_11
Xwl_driver_inv_en41 en en_bar[41] vdd gnd pinv_12
Xwl_driver_nand41 en_bar[41] in[41] net[41] vdd gnd pnand2_4
Xwl_driver_inv41 net[41] wl[41] vdd gnd pinv_11
Xwl_driver_inv_en42 en en_bar[42] vdd gnd pinv_12
Xwl_driver_nand42 en_bar[42] in[42] net[42] vdd gnd pnand2_4
Xwl_driver_inv42 net[42] wl[42] vdd gnd pinv_11
Xwl_driver_inv_en43 en en_bar[43] vdd gnd pinv_12
Xwl_driver_nand43 en_bar[43] in[43] net[43] vdd gnd pnand2_4
Xwl_driver_inv43 net[43] wl[43] vdd gnd pinv_11
Xwl_driver_inv_en44 en en_bar[44] vdd gnd pinv_12
Xwl_driver_nand44 en_bar[44] in[44] net[44] vdd gnd pnand2_4
Xwl_driver_inv44 net[44] wl[44] vdd gnd pinv_11
Xwl_driver_inv_en45 en en_bar[45] vdd gnd pinv_12
Xwl_driver_nand45 en_bar[45] in[45] net[45] vdd gnd pnand2_4
Xwl_driver_inv45 net[45] wl[45] vdd gnd pinv_11
Xwl_driver_inv_en46 en en_bar[46] vdd gnd pinv_12
Xwl_driver_nand46 en_bar[46] in[46] net[46] vdd gnd pnand2_4
Xwl_driver_inv46 net[46] wl[46] vdd gnd pinv_11
Xwl_driver_inv_en47 en en_bar[47] vdd gnd pinv_12
Xwl_driver_nand47 en_bar[47] in[47] net[47] vdd gnd pnand2_4
Xwl_driver_inv47 net[47] wl[47] vdd gnd pinv_11
Xwl_driver_inv_en48 en en_bar[48] vdd gnd pinv_12
Xwl_driver_nand48 en_bar[48] in[48] net[48] vdd gnd pnand2_4
Xwl_driver_inv48 net[48] wl[48] vdd gnd pinv_11
Xwl_driver_inv_en49 en en_bar[49] vdd gnd pinv_12
Xwl_driver_nand49 en_bar[49] in[49] net[49] vdd gnd pnand2_4
Xwl_driver_inv49 net[49] wl[49] vdd gnd pinv_11
Xwl_driver_inv_en50 en en_bar[50] vdd gnd pinv_12
Xwl_driver_nand50 en_bar[50] in[50] net[50] vdd gnd pnand2_4
Xwl_driver_inv50 net[50] wl[50] vdd gnd pinv_11
Xwl_driver_inv_en51 en en_bar[51] vdd gnd pinv_12
Xwl_driver_nand51 en_bar[51] in[51] net[51] vdd gnd pnand2_4
Xwl_driver_inv51 net[51] wl[51] vdd gnd pinv_11
Xwl_driver_inv_en52 en en_bar[52] vdd gnd pinv_12
Xwl_driver_nand52 en_bar[52] in[52] net[52] vdd gnd pnand2_4
Xwl_driver_inv52 net[52] wl[52] vdd gnd pinv_11
Xwl_driver_inv_en53 en en_bar[53] vdd gnd pinv_12
Xwl_driver_nand53 en_bar[53] in[53] net[53] vdd gnd pnand2_4
Xwl_driver_inv53 net[53] wl[53] vdd gnd pinv_11
Xwl_driver_inv_en54 en en_bar[54] vdd gnd pinv_12
Xwl_driver_nand54 en_bar[54] in[54] net[54] vdd gnd pnand2_4
Xwl_driver_inv54 net[54] wl[54] vdd gnd pinv_11
Xwl_driver_inv_en55 en en_bar[55] vdd gnd pinv_12
Xwl_driver_nand55 en_bar[55] in[55] net[55] vdd gnd pnand2_4
Xwl_driver_inv55 net[55] wl[55] vdd gnd pinv_11
Xwl_driver_inv_en56 en en_bar[56] vdd gnd pinv_12
Xwl_driver_nand56 en_bar[56] in[56] net[56] vdd gnd pnand2_4
Xwl_driver_inv56 net[56] wl[56] vdd gnd pinv_11
Xwl_driver_inv_en57 en en_bar[57] vdd gnd pinv_12
Xwl_driver_nand57 en_bar[57] in[57] net[57] vdd gnd pnand2_4
Xwl_driver_inv57 net[57] wl[57] vdd gnd pinv_11
Xwl_driver_inv_en58 en en_bar[58] vdd gnd pinv_12
Xwl_driver_nand58 en_bar[58] in[58] net[58] vdd gnd pnand2_4
Xwl_driver_inv58 net[58] wl[58] vdd gnd pinv_11
Xwl_driver_inv_en59 en en_bar[59] vdd gnd pinv_12
Xwl_driver_nand59 en_bar[59] in[59] net[59] vdd gnd pnand2_4
Xwl_driver_inv59 net[59] wl[59] vdd gnd pinv_11
Xwl_driver_inv_en60 en en_bar[60] vdd gnd pinv_12
Xwl_driver_nand60 en_bar[60] in[60] net[60] vdd gnd pnand2_4
Xwl_driver_inv60 net[60] wl[60] vdd gnd pinv_11
Xwl_driver_inv_en61 en en_bar[61] vdd gnd pinv_12
Xwl_driver_nand61 en_bar[61] in[61] net[61] vdd gnd pnand2_4
Xwl_driver_inv61 net[61] wl[61] vdd gnd pinv_11
Xwl_driver_inv_en62 en en_bar[62] vdd gnd pinv_12
Xwl_driver_nand62 en_bar[62] in[62] net[62] vdd gnd pnand2_4
Xwl_driver_inv62 net[62] wl[62] vdd gnd pinv_11
Xwl_driver_inv_en63 en en_bar[63] vdd gnd pinv_12
Xwl_driver_nand63 en_bar[63] in[63] net[63] vdd gnd pnand2_4
Xwl_driver_inv63 net[63] wl[63] vdd gnd pinv_11
Xwl_driver_inv_en64 en en_bar[64] vdd gnd pinv_12
Xwl_driver_nand64 en_bar[64] in[64] net[64] vdd gnd pnand2_4
Xwl_driver_inv64 net[64] wl[64] vdd gnd pinv_11
Xwl_driver_inv_en65 en en_bar[65] vdd gnd pinv_12
Xwl_driver_nand65 en_bar[65] in[65] net[65] vdd gnd pnand2_4
Xwl_driver_inv65 net[65] wl[65] vdd gnd pinv_11
Xwl_driver_inv_en66 en en_bar[66] vdd gnd pinv_12
Xwl_driver_nand66 en_bar[66] in[66] net[66] vdd gnd pnand2_4
Xwl_driver_inv66 net[66] wl[66] vdd gnd pinv_11
Xwl_driver_inv_en67 en en_bar[67] vdd gnd pinv_12
Xwl_driver_nand67 en_bar[67] in[67] net[67] vdd gnd pnand2_4
Xwl_driver_inv67 net[67] wl[67] vdd gnd pinv_11
Xwl_driver_inv_en68 en en_bar[68] vdd gnd pinv_12
Xwl_driver_nand68 en_bar[68] in[68] net[68] vdd gnd pnand2_4
Xwl_driver_inv68 net[68] wl[68] vdd gnd pinv_11
Xwl_driver_inv_en69 en en_bar[69] vdd gnd pinv_12
Xwl_driver_nand69 en_bar[69] in[69] net[69] vdd gnd pnand2_4
Xwl_driver_inv69 net[69] wl[69] vdd gnd pinv_11
Xwl_driver_inv_en70 en en_bar[70] vdd gnd pinv_12
Xwl_driver_nand70 en_bar[70] in[70] net[70] vdd gnd pnand2_4
Xwl_driver_inv70 net[70] wl[70] vdd gnd pinv_11
Xwl_driver_inv_en71 en en_bar[71] vdd gnd pinv_12
Xwl_driver_nand71 en_bar[71] in[71] net[71] vdd gnd pnand2_4
Xwl_driver_inv71 net[71] wl[71] vdd gnd pinv_11
Xwl_driver_inv_en72 en en_bar[72] vdd gnd pinv_12
Xwl_driver_nand72 en_bar[72] in[72] net[72] vdd gnd pnand2_4
Xwl_driver_inv72 net[72] wl[72] vdd gnd pinv_11
Xwl_driver_inv_en73 en en_bar[73] vdd gnd pinv_12
Xwl_driver_nand73 en_bar[73] in[73] net[73] vdd gnd pnand2_4
Xwl_driver_inv73 net[73] wl[73] vdd gnd pinv_11
Xwl_driver_inv_en74 en en_bar[74] vdd gnd pinv_12
Xwl_driver_nand74 en_bar[74] in[74] net[74] vdd gnd pnand2_4
Xwl_driver_inv74 net[74] wl[74] vdd gnd pinv_11
Xwl_driver_inv_en75 en en_bar[75] vdd gnd pinv_12
Xwl_driver_nand75 en_bar[75] in[75] net[75] vdd gnd pnand2_4
Xwl_driver_inv75 net[75] wl[75] vdd gnd pinv_11
Xwl_driver_inv_en76 en en_bar[76] vdd gnd pinv_12
Xwl_driver_nand76 en_bar[76] in[76] net[76] vdd gnd pnand2_4
Xwl_driver_inv76 net[76] wl[76] vdd gnd pinv_11
Xwl_driver_inv_en77 en en_bar[77] vdd gnd pinv_12
Xwl_driver_nand77 en_bar[77] in[77] net[77] vdd gnd pnand2_4
Xwl_driver_inv77 net[77] wl[77] vdd gnd pinv_11
Xwl_driver_inv_en78 en en_bar[78] vdd gnd pinv_12
Xwl_driver_nand78 en_bar[78] in[78] net[78] vdd gnd pnand2_4
Xwl_driver_inv78 net[78] wl[78] vdd gnd pinv_11
Xwl_driver_inv_en79 en en_bar[79] vdd gnd pinv_12
Xwl_driver_nand79 en_bar[79] in[79] net[79] vdd gnd pnand2_4
Xwl_driver_inv79 net[79] wl[79] vdd gnd pinv_11
Xwl_driver_inv_en80 en en_bar[80] vdd gnd pinv_12
Xwl_driver_nand80 en_bar[80] in[80] net[80] vdd gnd pnand2_4
Xwl_driver_inv80 net[80] wl[80] vdd gnd pinv_11
Xwl_driver_inv_en81 en en_bar[81] vdd gnd pinv_12
Xwl_driver_nand81 en_bar[81] in[81] net[81] vdd gnd pnand2_4
Xwl_driver_inv81 net[81] wl[81] vdd gnd pinv_11
Xwl_driver_inv_en82 en en_bar[82] vdd gnd pinv_12
Xwl_driver_nand82 en_bar[82] in[82] net[82] vdd gnd pnand2_4
Xwl_driver_inv82 net[82] wl[82] vdd gnd pinv_11
Xwl_driver_inv_en83 en en_bar[83] vdd gnd pinv_12
Xwl_driver_nand83 en_bar[83] in[83] net[83] vdd gnd pnand2_4
Xwl_driver_inv83 net[83] wl[83] vdd gnd pinv_11
Xwl_driver_inv_en84 en en_bar[84] vdd gnd pinv_12
Xwl_driver_nand84 en_bar[84] in[84] net[84] vdd gnd pnand2_4
Xwl_driver_inv84 net[84] wl[84] vdd gnd pinv_11
Xwl_driver_inv_en85 en en_bar[85] vdd gnd pinv_12
Xwl_driver_nand85 en_bar[85] in[85] net[85] vdd gnd pnand2_4
Xwl_driver_inv85 net[85] wl[85] vdd gnd pinv_11
Xwl_driver_inv_en86 en en_bar[86] vdd gnd pinv_12
Xwl_driver_nand86 en_bar[86] in[86] net[86] vdd gnd pnand2_4
Xwl_driver_inv86 net[86] wl[86] vdd gnd pinv_11
Xwl_driver_inv_en87 en en_bar[87] vdd gnd pinv_12
Xwl_driver_nand87 en_bar[87] in[87] net[87] vdd gnd pnand2_4
Xwl_driver_inv87 net[87] wl[87] vdd gnd pinv_11
Xwl_driver_inv_en88 en en_bar[88] vdd gnd pinv_12
Xwl_driver_nand88 en_bar[88] in[88] net[88] vdd gnd pnand2_4
Xwl_driver_inv88 net[88] wl[88] vdd gnd pinv_11
Xwl_driver_inv_en89 en en_bar[89] vdd gnd pinv_12
Xwl_driver_nand89 en_bar[89] in[89] net[89] vdd gnd pnand2_4
Xwl_driver_inv89 net[89] wl[89] vdd gnd pinv_11
Xwl_driver_inv_en90 en en_bar[90] vdd gnd pinv_12
Xwl_driver_nand90 en_bar[90] in[90] net[90] vdd gnd pnand2_4
Xwl_driver_inv90 net[90] wl[90] vdd gnd pinv_11
Xwl_driver_inv_en91 en en_bar[91] vdd gnd pinv_12
Xwl_driver_nand91 en_bar[91] in[91] net[91] vdd gnd pnand2_4
Xwl_driver_inv91 net[91] wl[91] vdd gnd pinv_11
Xwl_driver_inv_en92 en en_bar[92] vdd gnd pinv_12
Xwl_driver_nand92 en_bar[92] in[92] net[92] vdd gnd pnand2_4
Xwl_driver_inv92 net[92] wl[92] vdd gnd pinv_11
Xwl_driver_inv_en93 en en_bar[93] vdd gnd pinv_12
Xwl_driver_nand93 en_bar[93] in[93] net[93] vdd gnd pnand2_4
Xwl_driver_inv93 net[93] wl[93] vdd gnd pinv_11
Xwl_driver_inv_en94 en en_bar[94] vdd gnd pinv_12
Xwl_driver_nand94 en_bar[94] in[94] net[94] vdd gnd pnand2_4
Xwl_driver_inv94 net[94] wl[94] vdd gnd pinv_11
Xwl_driver_inv_en95 en en_bar[95] vdd gnd pinv_12
Xwl_driver_nand95 en_bar[95] in[95] net[95] vdd gnd pnand2_4
Xwl_driver_inv95 net[95] wl[95] vdd gnd pinv_11
Xwl_driver_inv_en96 en en_bar[96] vdd gnd pinv_12
Xwl_driver_nand96 en_bar[96] in[96] net[96] vdd gnd pnand2_4
Xwl_driver_inv96 net[96] wl[96] vdd gnd pinv_11
Xwl_driver_inv_en97 en en_bar[97] vdd gnd pinv_12
Xwl_driver_nand97 en_bar[97] in[97] net[97] vdd gnd pnand2_4
Xwl_driver_inv97 net[97] wl[97] vdd gnd pinv_11
Xwl_driver_inv_en98 en en_bar[98] vdd gnd pinv_12
Xwl_driver_nand98 en_bar[98] in[98] net[98] vdd gnd pnand2_4
Xwl_driver_inv98 net[98] wl[98] vdd gnd pinv_11
Xwl_driver_inv_en99 en en_bar[99] vdd gnd pinv_12
Xwl_driver_nand99 en_bar[99] in[99] net[99] vdd gnd pnand2_4
Xwl_driver_inv99 net[99] wl[99] vdd gnd pinv_11
Xwl_driver_inv_en100 en en_bar[100] vdd gnd pinv_12
Xwl_driver_nand100 en_bar[100] in[100] net[100] vdd gnd pnand2_4
Xwl_driver_inv100 net[100] wl[100] vdd gnd pinv_11
Xwl_driver_inv_en101 en en_bar[101] vdd gnd pinv_12
Xwl_driver_nand101 en_bar[101] in[101] net[101] vdd gnd pnand2_4
Xwl_driver_inv101 net[101] wl[101] vdd gnd pinv_11
Xwl_driver_inv_en102 en en_bar[102] vdd gnd pinv_12
Xwl_driver_nand102 en_bar[102] in[102] net[102] vdd gnd pnand2_4
Xwl_driver_inv102 net[102] wl[102] vdd gnd pinv_11
Xwl_driver_inv_en103 en en_bar[103] vdd gnd pinv_12
Xwl_driver_nand103 en_bar[103] in[103] net[103] vdd gnd pnand2_4
Xwl_driver_inv103 net[103] wl[103] vdd gnd pinv_11
Xwl_driver_inv_en104 en en_bar[104] vdd gnd pinv_12
Xwl_driver_nand104 en_bar[104] in[104] net[104] vdd gnd pnand2_4
Xwl_driver_inv104 net[104] wl[104] vdd gnd pinv_11
Xwl_driver_inv_en105 en en_bar[105] vdd gnd pinv_12
Xwl_driver_nand105 en_bar[105] in[105] net[105] vdd gnd pnand2_4
Xwl_driver_inv105 net[105] wl[105] vdd gnd pinv_11
Xwl_driver_inv_en106 en en_bar[106] vdd gnd pinv_12
Xwl_driver_nand106 en_bar[106] in[106] net[106] vdd gnd pnand2_4
Xwl_driver_inv106 net[106] wl[106] vdd gnd pinv_11
Xwl_driver_inv_en107 en en_bar[107] vdd gnd pinv_12
Xwl_driver_nand107 en_bar[107] in[107] net[107] vdd gnd pnand2_4
Xwl_driver_inv107 net[107] wl[107] vdd gnd pinv_11
Xwl_driver_inv_en108 en en_bar[108] vdd gnd pinv_12
Xwl_driver_nand108 en_bar[108] in[108] net[108] vdd gnd pnand2_4
Xwl_driver_inv108 net[108] wl[108] vdd gnd pinv_11
Xwl_driver_inv_en109 en en_bar[109] vdd gnd pinv_12
Xwl_driver_nand109 en_bar[109] in[109] net[109] vdd gnd pnand2_4
Xwl_driver_inv109 net[109] wl[109] vdd gnd pinv_11
Xwl_driver_inv_en110 en en_bar[110] vdd gnd pinv_12
Xwl_driver_nand110 en_bar[110] in[110] net[110] vdd gnd pnand2_4
Xwl_driver_inv110 net[110] wl[110] vdd gnd pinv_11
Xwl_driver_inv_en111 en en_bar[111] vdd gnd pinv_12
Xwl_driver_nand111 en_bar[111] in[111] net[111] vdd gnd pnand2_4
Xwl_driver_inv111 net[111] wl[111] vdd gnd pinv_11
Xwl_driver_inv_en112 en en_bar[112] vdd gnd pinv_12
Xwl_driver_nand112 en_bar[112] in[112] net[112] vdd gnd pnand2_4
Xwl_driver_inv112 net[112] wl[112] vdd gnd pinv_11
Xwl_driver_inv_en113 en en_bar[113] vdd gnd pinv_12
Xwl_driver_nand113 en_bar[113] in[113] net[113] vdd gnd pnand2_4
Xwl_driver_inv113 net[113] wl[113] vdd gnd pinv_11
Xwl_driver_inv_en114 en en_bar[114] vdd gnd pinv_12
Xwl_driver_nand114 en_bar[114] in[114] net[114] vdd gnd pnand2_4
Xwl_driver_inv114 net[114] wl[114] vdd gnd pinv_11
Xwl_driver_inv_en115 en en_bar[115] vdd gnd pinv_12
Xwl_driver_nand115 en_bar[115] in[115] net[115] vdd gnd pnand2_4
Xwl_driver_inv115 net[115] wl[115] vdd gnd pinv_11
Xwl_driver_inv_en116 en en_bar[116] vdd gnd pinv_12
Xwl_driver_nand116 en_bar[116] in[116] net[116] vdd gnd pnand2_4
Xwl_driver_inv116 net[116] wl[116] vdd gnd pinv_11
Xwl_driver_inv_en117 en en_bar[117] vdd gnd pinv_12
Xwl_driver_nand117 en_bar[117] in[117] net[117] vdd gnd pnand2_4
Xwl_driver_inv117 net[117] wl[117] vdd gnd pinv_11
Xwl_driver_inv_en118 en en_bar[118] vdd gnd pinv_12
Xwl_driver_nand118 en_bar[118] in[118] net[118] vdd gnd pnand2_4
Xwl_driver_inv118 net[118] wl[118] vdd gnd pinv_11
Xwl_driver_inv_en119 en en_bar[119] vdd gnd pinv_12
Xwl_driver_nand119 en_bar[119] in[119] net[119] vdd gnd pnand2_4
Xwl_driver_inv119 net[119] wl[119] vdd gnd pinv_11
Xwl_driver_inv_en120 en en_bar[120] vdd gnd pinv_12
Xwl_driver_nand120 en_bar[120] in[120] net[120] vdd gnd pnand2_4
Xwl_driver_inv120 net[120] wl[120] vdd gnd pinv_11
Xwl_driver_inv_en121 en en_bar[121] vdd gnd pinv_12
Xwl_driver_nand121 en_bar[121] in[121] net[121] vdd gnd pnand2_4
Xwl_driver_inv121 net[121] wl[121] vdd gnd pinv_11
Xwl_driver_inv_en122 en en_bar[122] vdd gnd pinv_12
Xwl_driver_nand122 en_bar[122] in[122] net[122] vdd gnd pnand2_4
Xwl_driver_inv122 net[122] wl[122] vdd gnd pinv_11
Xwl_driver_inv_en123 en en_bar[123] vdd gnd pinv_12
Xwl_driver_nand123 en_bar[123] in[123] net[123] vdd gnd pnand2_4
Xwl_driver_inv123 net[123] wl[123] vdd gnd pinv_11
Xwl_driver_inv_en124 en en_bar[124] vdd gnd pinv_12
Xwl_driver_nand124 en_bar[124] in[124] net[124] vdd gnd pnand2_4
Xwl_driver_inv124 net[124] wl[124] vdd gnd pinv_11
Xwl_driver_inv_en125 en en_bar[125] vdd gnd pinv_12
Xwl_driver_nand125 en_bar[125] in[125] net[125] vdd gnd pnand2_4
Xwl_driver_inv125 net[125] wl[125] vdd gnd pinv_11
Xwl_driver_inv_en126 en en_bar[126] vdd gnd pinv_12
Xwl_driver_nand126 en_bar[126] in[126] net[126] vdd gnd pnand2_4
Xwl_driver_inv126 net[126] wl[126] vdd gnd pinv_11
Xwl_driver_inv_en127 en en_bar[127] vdd gnd pinv_12
Xwl_driver_nand127 en_bar[127] in[127] net[127] vdd gnd pnand2_4
Xwl_driver_inv127 net[127] wl[127] vdd gnd pinv_11
Xwl_driver_inv_en128 en en_bar[128] vdd gnd pinv_12
Xwl_driver_nand128 en_bar[128] in[128] net[128] vdd gnd pnand2_4
Xwl_driver_inv128 net[128] wl[128] vdd gnd pinv_11
Xwl_driver_inv_en129 en en_bar[129] vdd gnd pinv_12
Xwl_driver_nand129 en_bar[129] in[129] net[129] vdd gnd pnand2_4
Xwl_driver_inv129 net[129] wl[129] vdd gnd pinv_11
Xwl_driver_inv_en130 en en_bar[130] vdd gnd pinv_12
Xwl_driver_nand130 en_bar[130] in[130] net[130] vdd gnd pnand2_4
Xwl_driver_inv130 net[130] wl[130] vdd gnd pinv_11
Xwl_driver_inv_en131 en en_bar[131] vdd gnd pinv_12
Xwl_driver_nand131 en_bar[131] in[131] net[131] vdd gnd pnand2_4
Xwl_driver_inv131 net[131] wl[131] vdd gnd pinv_11
Xwl_driver_inv_en132 en en_bar[132] vdd gnd pinv_12
Xwl_driver_nand132 en_bar[132] in[132] net[132] vdd gnd pnand2_4
Xwl_driver_inv132 net[132] wl[132] vdd gnd pinv_11
Xwl_driver_inv_en133 en en_bar[133] vdd gnd pinv_12
Xwl_driver_nand133 en_bar[133] in[133] net[133] vdd gnd pnand2_4
Xwl_driver_inv133 net[133] wl[133] vdd gnd pinv_11
Xwl_driver_inv_en134 en en_bar[134] vdd gnd pinv_12
Xwl_driver_nand134 en_bar[134] in[134] net[134] vdd gnd pnand2_4
Xwl_driver_inv134 net[134] wl[134] vdd gnd pinv_11
Xwl_driver_inv_en135 en en_bar[135] vdd gnd pinv_12
Xwl_driver_nand135 en_bar[135] in[135] net[135] vdd gnd pnand2_4
Xwl_driver_inv135 net[135] wl[135] vdd gnd pinv_11
Xwl_driver_inv_en136 en en_bar[136] vdd gnd pinv_12
Xwl_driver_nand136 en_bar[136] in[136] net[136] vdd gnd pnand2_4
Xwl_driver_inv136 net[136] wl[136] vdd gnd pinv_11
Xwl_driver_inv_en137 en en_bar[137] vdd gnd pinv_12
Xwl_driver_nand137 en_bar[137] in[137] net[137] vdd gnd pnand2_4
Xwl_driver_inv137 net[137] wl[137] vdd gnd pinv_11
Xwl_driver_inv_en138 en en_bar[138] vdd gnd pinv_12
Xwl_driver_nand138 en_bar[138] in[138] net[138] vdd gnd pnand2_4
Xwl_driver_inv138 net[138] wl[138] vdd gnd pinv_11
Xwl_driver_inv_en139 en en_bar[139] vdd gnd pinv_12
Xwl_driver_nand139 en_bar[139] in[139] net[139] vdd gnd pnand2_4
Xwl_driver_inv139 net[139] wl[139] vdd gnd pinv_11
Xwl_driver_inv_en140 en en_bar[140] vdd gnd pinv_12
Xwl_driver_nand140 en_bar[140] in[140] net[140] vdd gnd pnand2_4
Xwl_driver_inv140 net[140] wl[140] vdd gnd pinv_11
Xwl_driver_inv_en141 en en_bar[141] vdd gnd pinv_12
Xwl_driver_nand141 en_bar[141] in[141] net[141] vdd gnd pnand2_4
Xwl_driver_inv141 net[141] wl[141] vdd gnd pinv_11
Xwl_driver_inv_en142 en en_bar[142] vdd gnd pinv_12
Xwl_driver_nand142 en_bar[142] in[142] net[142] vdd gnd pnand2_4
Xwl_driver_inv142 net[142] wl[142] vdd gnd pinv_11
Xwl_driver_inv_en143 en en_bar[143] vdd gnd pinv_12
Xwl_driver_nand143 en_bar[143] in[143] net[143] vdd gnd pnand2_4
Xwl_driver_inv143 net[143] wl[143] vdd gnd pinv_11
Xwl_driver_inv_en144 en en_bar[144] vdd gnd pinv_12
Xwl_driver_nand144 en_bar[144] in[144] net[144] vdd gnd pnand2_4
Xwl_driver_inv144 net[144] wl[144] vdd gnd pinv_11
Xwl_driver_inv_en145 en en_bar[145] vdd gnd pinv_12
Xwl_driver_nand145 en_bar[145] in[145] net[145] vdd gnd pnand2_4
Xwl_driver_inv145 net[145] wl[145] vdd gnd pinv_11
Xwl_driver_inv_en146 en en_bar[146] vdd gnd pinv_12
Xwl_driver_nand146 en_bar[146] in[146] net[146] vdd gnd pnand2_4
Xwl_driver_inv146 net[146] wl[146] vdd gnd pinv_11
Xwl_driver_inv_en147 en en_bar[147] vdd gnd pinv_12
Xwl_driver_nand147 en_bar[147] in[147] net[147] vdd gnd pnand2_4
Xwl_driver_inv147 net[147] wl[147] vdd gnd pinv_11
Xwl_driver_inv_en148 en en_bar[148] vdd gnd pinv_12
Xwl_driver_nand148 en_bar[148] in[148] net[148] vdd gnd pnand2_4
Xwl_driver_inv148 net[148] wl[148] vdd gnd pinv_11
Xwl_driver_inv_en149 en en_bar[149] vdd gnd pinv_12
Xwl_driver_nand149 en_bar[149] in[149] net[149] vdd gnd pnand2_4
Xwl_driver_inv149 net[149] wl[149] vdd gnd pinv_11
Xwl_driver_inv_en150 en en_bar[150] vdd gnd pinv_12
Xwl_driver_nand150 en_bar[150] in[150] net[150] vdd gnd pnand2_4
Xwl_driver_inv150 net[150] wl[150] vdd gnd pinv_11
Xwl_driver_inv_en151 en en_bar[151] vdd gnd pinv_12
Xwl_driver_nand151 en_bar[151] in[151] net[151] vdd gnd pnand2_4
Xwl_driver_inv151 net[151] wl[151] vdd gnd pinv_11
Xwl_driver_inv_en152 en en_bar[152] vdd gnd pinv_12
Xwl_driver_nand152 en_bar[152] in[152] net[152] vdd gnd pnand2_4
Xwl_driver_inv152 net[152] wl[152] vdd gnd pinv_11
Xwl_driver_inv_en153 en en_bar[153] vdd gnd pinv_12
Xwl_driver_nand153 en_bar[153] in[153] net[153] vdd gnd pnand2_4
Xwl_driver_inv153 net[153] wl[153] vdd gnd pinv_11
Xwl_driver_inv_en154 en en_bar[154] vdd gnd pinv_12
Xwl_driver_nand154 en_bar[154] in[154] net[154] vdd gnd pnand2_4
Xwl_driver_inv154 net[154] wl[154] vdd gnd pinv_11
Xwl_driver_inv_en155 en en_bar[155] vdd gnd pinv_12
Xwl_driver_nand155 en_bar[155] in[155] net[155] vdd gnd pnand2_4
Xwl_driver_inv155 net[155] wl[155] vdd gnd pinv_11
Xwl_driver_inv_en156 en en_bar[156] vdd gnd pinv_12
Xwl_driver_nand156 en_bar[156] in[156] net[156] vdd gnd pnand2_4
Xwl_driver_inv156 net[156] wl[156] vdd gnd pinv_11
Xwl_driver_inv_en157 en en_bar[157] vdd gnd pinv_12
Xwl_driver_nand157 en_bar[157] in[157] net[157] vdd gnd pnand2_4
Xwl_driver_inv157 net[157] wl[157] vdd gnd pinv_11
Xwl_driver_inv_en158 en en_bar[158] vdd gnd pinv_12
Xwl_driver_nand158 en_bar[158] in[158] net[158] vdd gnd pnand2_4
Xwl_driver_inv158 net[158] wl[158] vdd gnd pinv_11
Xwl_driver_inv_en159 en en_bar[159] vdd gnd pinv_12
Xwl_driver_nand159 en_bar[159] in[159] net[159] vdd gnd pnand2_4
Xwl_driver_inv159 net[159] wl[159] vdd gnd pinv_11
Xwl_driver_inv_en160 en en_bar[160] vdd gnd pinv_12
Xwl_driver_nand160 en_bar[160] in[160] net[160] vdd gnd pnand2_4
Xwl_driver_inv160 net[160] wl[160] vdd gnd pinv_11
Xwl_driver_inv_en161 en en_bar[161] vdd gnd pinv_12
Xwl_driver_nand161 en_bar[161] in[161] net[161] vdd gnd pnand2_4
Xwl_driver_inv161 net[161] wl[161] vdd gnd pinv_11
Xwl_driver_inv_en162 en en_bar[162] vdd gnd pinv_12
Xwl_driver_nand162 en_bar[162] in[162] net[162] vdd gnd pnand2_4
Xwl_driver_inv162 net[162] wl[162] vdd gnd pinv_11
Xwl_driver_inv_en163 en en_bar[163] vdd gnd pinv_12
Xwl_driver_nand163 en_bar[163] in[163] net[163] vdd gnd pnand2_4
Xwl_driver_inv163 net[163] wl[163] vdd gnd pinv_11
Xwl_driver_inv_en164 en en_bar[164] vdd gnd pinv_12
Xwl_driver_nand164 en_bar[164] in[164] net[164] vdd gnd pnand2_4
Xwl_driver_inv164 net[164] wl[164] vdd gnd pinv_11
Xwl_driver_inv_en165 en en_bar[165] vdd gnd pinv_12
Xwl_driver_nand165 en_bar[165] in[165] net[165] vdd gnd pnand2_4
Xwl_driver_inv165 net[165] wl[165] vdd gnd pinv_11
Xwl_driver_inv_en166 en en_bar[166] vdd gnd pinv_12
Xwl_driver_nand166 en_bar[166] in[166] net[166] vdd gnd pnand2_4
Xwl_driver_inv166 net[166] wl[166] vdd gnd pinv_11
Xwl_driver_inv_en167 en en_bar[167] vdd gnd pinv_12
Xwl_driver_nand167 en_bar[167] in[167] net[167] vdd gnd pnand2_4
Xwl_driver_inv167 net[167] wl[167] vdd gnd pinv_11
Xwl_driver_inv_en168 en en_bar[168] vdd gnd pinv_12
Xwl_driver_nand168 en_bar[168] in[168] net[168] vdd gnd pnand2_4
Xwl_driver_inv168 net[168] wl[168] vdd gnd pinv_11
Xwl_driver_inv_en169 en en_bar[169] vdd gnd pinv_12
Xwl_driver_nand169 en_bar[169] in[169] net[169] vdd gnd pnand2_4
Xwl_driver_inv169 net[169] wl[169] vdd gnd pinv_11
Xwl_driver_inv_en170 en en_bar[170] vdd gnd pinv_12
Xwl_driver_nand170 en_bar[170] in[170] net[170] vdd gnd pnand2_4
Xwl_driver_inv170 net[170] wl[170] vdd gnd pinv_11
Xwl_driver_inv_en171 en en_bar[171] vdd gnd pinv_12
Xwl_driver_nand171 en_bar[171] in[171] net[171] vdd gnd pnand2_4
Xwl_driver_inv171 net[171] wl[171] vdd gnd pinv_11
Xwl_driver_inv_en172 en en_bar[172] vdd gnd pinv_12
Xwl_driver_nand172 en_bar[172] in[172] net[172] vdd gnd pnand2_4
Xwl_driver_inv172 net[172] wl[172] vdd gnd pinv_11
Xwl_driver_inv_en173 en en_bar[173] vdd gnd pinv_12
Xwl_driver_nand173 en_bar[173] in[173] net[173] vdd gnd pnand2_4
Xwl_driver_inv173 net[173] wl[173] vdd gnd pinv_11
Xwl_driver_inv_en174 en en_bar[174] vdd gnd pinv_12
Xwl_driver_nand174 en_bar[174] in[174] net[174] vdd gnd pnand2_4
Xwl_driver_inv174 net[174] wl[174] vdd gnd pinv_11
Xwl_driver_inv_en175 en en_bar[175] vdd gnd pinv_12
Xwl_driver_nand175 en_bar[175] in[175] net[175] vdd gnd pnand2_4
Xwl_driver_inv175 net[175] wl[175] vdd gnd pinv_11
Xwl_driver_inv_en176 en en_bar[176] vdd gnd pinv_12
Xwl_driver_nand176 en_bar[176] in[176] net[176] vdd gnd pnand2_4
Xwl_driver_inv176 net[176] wl[176] vdd gnd pinv_11
Xwl_driver_inv_en177 en en_bar[177] vdd gnd pinv_12
Xwl_driver_nand177 en_bar[177] in[177] net[177] vdd gnd pnand2_4
Xwl_driver_inv177 net[177] wl[177] vdd gnd pinv_11
Xwl_driver_inv_en178 en en_bar[178] vdd gnd pinv_12
Xwl_driver_nand178 en_bar[178] in[178] net[178] vdd gnd pnand2_4
Xwl_driver_inv178 net[178] wl[178] vdd gnd pinv_11
Xwl_driver_inv_en179 en en_bar[179] vdd gnd pinv_12
Xwl_driver_nand179 en_bar[179] in[179] net[179] vdd gnd pnand2_4
Xwl_driver_inv179 net[179] wl[179] vdd gnd pinv_11
Xwl_driver_inv_en180 en en_bar[180] vdd gnd pinv_12
Xwl_driver_nand180 en_bar[180] in[180] net[180] vdd gnd pnand2_4
Xwl_driver_inv180 net[180] wl[180] vdd gnd pinv_11
Xwl_driver_inv_en181 en en_bar[181] vdd gnd pinv_12
Xwl_driver_nand181 en_bar[181] in[181] net[181] vdd gnd pnand2_4
Xwl_driver_inv181 net[181] wl[181] vdd gnd pinv_11
Xwl_driver_inv_en182 en en_bar[182] vdd gnd pinv_12
Xwl_driver_nand182 en_bar[182] in[182] net[182] vdd gnd pnand2_4
Xwl_driver_inv182 net[182] wl[182] vdd gnd pinv_11
Xwl_driver_inv_en183 en en_bar[183] vdd gnd pinv_12
Xwl_driver_nand183 en_bar[183] in[183] net[183] vdd gnd pnand2_4
Xwl_driver_inv183 net[183] wl[183] vdd gnd pinv_11
Xwl_driver_inv_en184 en en_bar[184] vdd gnd pinv_12
Xwl_driver_nand184 en_bar[184] in[184] net[184] vdd gnd pnand2_4
Xwl_driver_inv184 net[184] wl[184] vdd gnd pinv_11
Xwl_driver_inv_en185 en en_bar[185] vdd gnd pinv_12
Xwl_driver_nand185 en_bar[185] in[185] net[185] vdd gnd pnand2_4
Xwl_driver_inv185 net[185] wl[185] vdd gnd pinv_11
Xwl_driver_inv_en186 en en_bar[186] vdd gnd pinv_12
Xwl_driver_nand186 en_bar[186] in[186] net[186] vdd gnd pnand2_4
Xwl_driver_inv186 net[186] wl[186] vdd gnd pinv_11
Xwl_driver_inv_en187 en en_bar[187] vdd gnd pinv_12
Xwl_driver_nand187 en_bar[187] in[187] net[187] vdd gnd pnand2_4
Xwl_driver_inv187 net[187] wl[187] vdd gnd pinv_11
Xwl_driver_inv_en188 en en_bar[188] vdd gnd pinv_12
Xwl_driver_nand188 en_bar[188] in[188] net[188] vdd gnd pnand2_4
Xwl_driver_inv188 net[188] wl[188] vdd gnd pinv_11
Xwl_driver_inv_en189 en en_bar[189] vdd gnd pinv_12
Xwl_driver_nand189 en_bar[189] in[189] net[189] vdd gnd pnand2_4
Xwl_driver_inv189 net[189] wl[189] vdd gnd pinv_11
Xwl_driver_inv_en190 en en_bar[190] vdd gnd pinv_12
Xwl_driver_nand190 en_bar[190] in[190] net[190] vdd gnd pnand2_4
Xwl_driver_inv190 net[190] wl[190] vdd gnd pinv_11
Xwl_driver_inv_en191 en en_bar[191] vdd gnd pinv_12
Xwl_driver_nand191 en_bar[191] in[191] net[191] vdd gnd pnand2_4
Xwl_driver_inv191 net[191] wl[191] vdd gnd pinv_11
Xwl_driver_inv_en192 en en_bar[192] vdd gnd pinv_12
Xwl_driver_nand192 en_bar[192] in[192] net[192] vdd gnd pnand2_4
Xwl_driver_inv192 net[192] wl[192] vdd gnd pinv_11
Xwl_driver_inv_en193 en en_bar[193] vdd gnd pinv_12
Xwl_driver_nand193 en_bar[193] in[193] net[193] vdd gnd pnand2_4
Xwl_driver_inv193 net[193] wl[193] vdd gnd pinv_11
Xwl_driver_inv_en194 en en_bar[194] vdd gnd pinv_12
Xwl_driver_nand194 en_bar[194] in[194] net[194] vdd gnd pnand2_4
Xwl_driver_inv194 net[194] wl[194] vdd gnd pinv_11
Xwl_driver_inv_en195 en en_bar[195] vdd gnd pinv_12
Xwl_driver_nand195 en_bar[195] in[195] net[195] vdd gnd pnand2_4
Xwl_driver_inv195 net[195] wl[195] vdd gnd pinv_11
Xwl_driver_inv_en196 en en_bar[196] vdd gnd pinv_12
Xwl_driver_nand196 en_bar[196] in[196] net[196] vdd gnd pnand2_4
Xwl_driver_inv196 net[196] wl[196] vdd gnd pinv_11
Xwl_driver_inv_en197 en en_bar[197] vdd gnd pinv_12
Xwl_driver_nand197 en_bar[197] in[197] net[197] vdd gnd pnand2_4
Xwl_driver_inv197 net[197] wl[197] vdd gnd pinv_11
Xwl_driver_inv_en198 en en_bar[198] vdd gnd pinv_12
Xwl_driver_nand198 en_bar[198] in[198] net[198] vdd gnd pnand2_4
Xwl_driver_inv198 net[198] wl[198] vdd gnd pinv_11
Xwl_driver_inv_en199 en en_bar[199] vdd gnd pinv_12
Xwl_driver_nand199 en_bar[199] in[199] net[199] vdd gnd pnand2_4
Xwl_driver_inv199 net[199] wl[199] vdd gnd pinv_11
Xwl_driver_inv_en200 en en_bar[200] vdd gnd pinv_12
Xwl_driver_nand200 en_bar[200] in[200] net[200] vdd gnd pnand2_4
Xwl_driver_inv200 net[200] wl[200] vdd gnd pinv_11
Xwl_driver_inv_en201 en en_bar[201] vdd gnd pinv_12
Xwl_driver_nand201 en_bar[201] in[201] net[201] vdd gnd pnand2_4
Xwl_driver_inv201 net[201] wl[201] vdd gnd pinv_11
Xwl_driver_inv_en202 en en_bar[202] vdd gnd pinv_12
Xwl_driver_nand202 en_bar[202] in[202] net[202] vdd gnd pnand2_4
Xwl_driver_inv202 net[202] wl[202] vdd gnd pinv_11
Xwl_driver_inv_en203 en en_bar[203] vdd gnd pinv_12
Xwl_driver_nand203 en_bar[203] in[203] net[203] vdd gnd pnand2_4
Xwl_driver_inv203 net[203] wl[203] vdd gnd pinv_11
Xwl_driver_inv_en204 en en_bar[204] vdd gnd pinv_12
Xwl_driver_nand204 en_bar[204] in[204] net[204] vdd gnd pnand2_4
Xwl_driver_inv204 net[204] wl[204] vdd gnd pinv_11
Xwl_driver_inv_en205 en en_bar[205] vdd gnd pinv_12
Xwl_driver_nand205 en_bar[205] in[205] net[205] vdd gnd pnand2_4
Xwl_driver_inv205 net[205] wl[205] vdd gnd pinv_11
Xwl_driver_inv_en206 en en_bar[206] vdd gnd pinv_12
Xwl_driver_nand206 en_bar[206] in[206] net[206] vdd gnd pnand2_4
Xwl_driver_inv206 net[206] wl[206] vdd gnd pinv_11
Xwl_driver_inv_en207 en en_bar[207] vdd gnd pinv_12
Xwl_driver_nand207 en_bar[207] in[207] net[207] vdd gnd pnand2_4
Xwl_driver_inv207 net[207] wl[207] vdd gnd pinv_11
Xwl_driver_inv_en208 en en_bar[208] vdd gnd pinv_12
Xwl_driver_nand208 en_bar[208] in[208] net[208] vdd gnd pnand2_4
Xwl_driver_inv208 net[208] wl[208] vdd gnd pinv_11
Xwl_driver_inv_en209 en en_bar[209] vdd gnd pinv_12
Xwl_driver_nand209 en_bar[209] in[209] net[209] vdd gnd pnand2_4
Xwl_driver_inv209 net[209] wl[209] vdd gnd pinv_11
Xwl_driver_inv_en210 en en_bar[210] vdd gnd pinv_12
Xwl_driver_nand210 en_bar[210] in[210] net[210] vdd gnd pnand2_4
Xwl_driver_inv210 net[210] wl[210] vdd gnd pinv_11
Xwl_driver_inv_en211 en en_bar[211] vdd gnd pinv_12
Xwl_driver_nand211 en_bar[211] in[211] net[211] vdd gnd pnand2_4
Xwl_driver_inv211 net[211] wl[211] vdd gnd pinv_11
Xwl_driver_inv_en212 en en_bar[212] vdd gnd pinv_12
Xwl_driver_nand212 en_bar[212] in[212] net[212] vdd gnd pnand2_4
Xwl_driver_inv212 net[212] wl[212] vdd gnd pinv_11
Xwl_driver_inv_en213 en en_bar[213] vdd gnd pinv_12
Xwl_driver_nand213 en_bar[213] in[213] net[213] vdd gnd pnand2_4
Xwl_driver_inv213 net[213] wl[213] vdd gnd pinv_11
Xwl_driver_inv_en214 en en_bar[214] vdd gnd pinv_12
Xwl_driver_nand214 en_bar[214] in[214] net[214] vdd gnd pnand2_4
Xwl_driver_inv214 net[214] wl[214] vdd gnd pinv_11
Xwl_driver_inv_en215 en en_bar[215] vdd gnd pinv_12
Xwl_driver_nand215 en_bar[215] in[215] net[215] vdd gnd pnand2_4
Xwl_driver_inv215 net[215] wl[215] vdd gnd pinv_11
Xwl_driver_inv_en216 en en_bar[216] vdd gnd pinv_12
Xwl_driver_nand216 en_bar[216] in[216] net[216] vdd gnd pnand2_4
Xwl_driver_inv216 net[216] wl[216] vdd gnd pinv_11
Xwl_driver_inv_en217 en en_bar[217] vdd gnd pinv_12
Xwl_driver_nand217 en_bar[217] in[217] net[217] vdd gnd pnand2_4
Xwl_driver_inv217 net[217] wl[217] vdd gnd pinv_11
Xwl_driver_inv_en218 en en_bar[218] vdd gnd pinv_12
Xwl_driver_nand218 en_bar[218] in[218] net[218] vdd gnd pnand2_4
Xwl_driver_inv218 net[218] wl[218] vdd gnd pinv_11
Xwl_driver_inv_en219 en en_bar[219] vdd gnd pinv_12
Xwl_driver_nand219 en_bar[219] in[219] net[219] vdd gnd pnand2_4
Xwl_driver_inv219 net[219] wl[219] vdd gnd pinv_11
Xwl_driver_inv_en220 en en_bar[220] vdd gnd pinv_12
Xwl_driver_nand220 en_bar[220] in[220] net[220] vdd gnd pnand2_4
Xwl_driver_inv220 net[220] wl[220] vdd gnd pinv_11
Xwl_driver_inv_en221 en en_bar[221] vdd gnd pinv_12
Xwl_driver_nand221 en_bar[221] in[221] net[221] vdd gnd pnand2_4
Xwl_driver_inv221 net[221] wl[221] vdd gnd pinv_11
Xwl_driver_inv_en222 en en_bar[222] vdd gnd pinv_12
Xwl_driver_nand222 en_bar[222] in[222] net[222] vdd gnd pnand2_4
Xwl_driver_inv222 net[222] wl[222] vdd gnd pinv_11
Xwl_driver_inv_en223 en en_bar[223] vdd gnd pinv_12
Xwl_driver_nand223 en_bar[223] in[223] net[223] vdd gnd pnand2_4
Xwl_driver_inv223 net[223] wl[223] vdd gnd pinv_11
Xwl_driver_inv_en224 en en_bar[224] vdd gnd pinv_12
Xwl_driver_nand224 en_bar[224] in[224] net[224] vdd gnd pnand2_4
Xwl_driver_inv224 net[224] wl[224] vdd gnd pinv_11
Xwl_driver_inv_en225 en en_bar[225] vdd gnd pinv_12
Xwl_driver_nand225 en_bar[225] in[225] net[225] vdd gnd pnand2_4
Xwl_driver_inv225 net[225] wl[225] vdd gnd pinv_11
Xwl_driver_inv_en226 en en_bar[226] vdd gnd pinv_12
Xwl_driver_nand226 en_bar[226] in[226] net[226] vdd gnd pnand2_4
Xwl_driver_inv226 net[226] wl[226] vdd gnd pinv_11
Xwl_driver_inv_en227 en en_bar[227] vdd gnd pinv_12
Xwl_driver_nand227 en_bar[227] in[227] net[227] vdd gnd pnand2_4
Xwl_driver_inv227 net[227] wl[227] vdd gnd pinv_11
Xwl_driver_inv_en228 en en_bar[228] vdd gnd pinv_12
Xwl_driver_nand228 en_bar[228] in[228] net[228] vdd gnd pnand2_4
Xwl_driver_inv228 net[228] wl[228] vdd gnd pinv_11
Xwl_driver_inv_en229 en en_bar[229] vdd gnd pinv_12
Xwl_driver_nand229 en_bar[229] in[229] net[229] vdd gnd pnand2_4
Xwl_driver_inv229 net[229] wl[229] vdd gnd pinv_11
Xwl_driver_inv_en230 en en_bar[230] vdd gnd pinv_12
Xwl_driver_nand230 en_bar[230] in[230] net[230] vdd gnd pnand2_4
Xwl_driver_inv230 net[230] wl[230] vdd gnd pinv_11
Xwl_driver_inv_en231 en en_bar[231] vdd gnd pinv_12
Xwl_driver_nand231 en_bar[231] in[231] net[231] vdd gnd pnand2_4
Xwl_driver_inv231 net[231] wl[231] vdd gnd pinv_11
Xwl_driver_inv_en232 en en_bar[232] vdd gnd pinv_12
Xwl_driver_nand232 en_bar[232] in[232] net[232] vdd gnd pnand2_4
Xwl_driver_inv232 net[232] wl[232] vdd gnd pinv_11
Xwl_driver_inv_en233 en en_bar[233] vdd gnd pinv_12
Xwl_driver_nand233 en_bar[233] in[233] net[233] vdd gnd pnand2_4
Xwl_driver_inv233 net[233] wl[233] vdd gnd pinv_11
Xwl_driver_inv_en234 en en_bar[234] vdd gnd pinv_12
Xwl_driver_nand234 en_bar[234] in[234] net[234] vdd gnd pnand2_4
Xwl_driver_inv234 net[234] wl[234] vdd gnd pinv_11
Xwl_driver_inv_en235 en en_bar[235] vdd gnd pinv_12
Xwl_driver_nand235 en_bar[235] in[235] net[235] vdd gnd pnand2_4
Xwl_driver_inv235 net[235] wl[235] vdd gnd pinv_11
Xwl_driver_inv_en236 en en_bar[236] vdd gnd pinv_12
Xwl_driver_nand236 en_bar[236] in[236] net[236] vdd gnd pnand2_4
Xwl_driver_inv236 net[236] wl[236] vdd gnd pinv_11
Xwl_driver_inv_en237 en en_bar[237] vdd gnd pinv_12
Xwl_driver_nand237 en_bar[237] in[237] net[237] vdd gnd pnand2_4
Xwl_driver_inv237 net[237] wl[237] vdd gnd pinv_11
Xwl_driver_inv_en238 en en_bar[238] vdd gnd pinv_12
Xwl_driver_nand238 en_bar[238] in[238] net[238] vdd gnd pnand2_4
Xwl_driver_inv238 net[238] wl[238] vdd gnd pinv_11
Xwl_driver_inv_en239 en en_bar[239] vdd gnd pinv_12
Xwl_driver_nand239 en_bar[239] in[239] net[239] vdd gnd pnand2_4
Xwl_driver_inv239 net[239] wl[239] vdd gnd pinv_11
Xwl_driver_inv_en240 en en_bar[240] vdd gnd pinv_12
Xwl_driver_nand240 en_bar[240] in[240] net[240] vdd gnd pnand2_4
Xwl_driver_inv240 net[240] wl[240] vdd gnd pinv_11
Xwl_driver_inv_en241 en en_bar[241] vdd gnd pinv_12
Xwl_driver_nand241 en_bar[241] in[241] net[241] vdd gnd pnand2_4
Xwl_driver_inv241 net[241] wl[241] vdd gnd pinv_11
Xwl_driver_inv_en242 en en_bar[242] vdd gnd pinv_12
Xwl_driver_nand242 en_bar[242] in[242] net[242] vdd gnd pnand2_4
Xwl_driver_inv242 net[242] wl[242] vdd gnd pinv_11
Xwl_driver_inv_en243 en en_bar[243] vdd gnd pinv_12
Xwl_driver_nand243 en_bar[243] in[243] net[243] vdd gnd pnand2_4
Xwl_driver_inv243 net[243] wl[243] vdd gnd pinv_11
Xwl_driver_inv_en244 en en_bar[244] vdd gnd pinv_12
Xwl_driver_nand244 en_bar[244] in[244] net[244] vdd gnd pnand2_4
Xwl_driver_inv244 net[244] wl[244] vdd gnd pinv_11
Xwl_driver_inv_en245 en en_bar[245] vdd gnd pinv_12
Xwl_driver_nand245 en_bar[245] in[245] net[245] vdd gnd pnand2_4
Xwl_driver_inv245 net[245] wl[245] vdd gnd pinv_11
Xwl_driver_inv_en246 en en_bar[246] vdd gnd pinv_12
Xwl_driver_nand246 en_bar[246] in[246] net[246] vdd gnd pnand2_4
Xwl_driver_inv246 net[246] wl[246] vdd gnd pinv_11
Xwl_driver_inv_en247 en en_bar[247] vdd gnd pinv_12
Xwl_driver_nand247 en_bar[247] in[247] net[247] vdd gnd pnand2_4
Xwl_driver_inv247 net[247] wl[247] vdd gnd pinv_11
Xwl_driver_inv_en248 en en_bar[248] vdd gnd pinv_12
Xwl_driver_nand248 en_bar[248] in[248] net[248] vdd gnd pnand2_4
Xwl_driver_inv248 net[248] wl[248] vdd gnd pinv_11
Xwl_driver_inv_en249 en en_bar[249] vdd gnd pinv_12
Xwl_driver_nand249 en_bar[249] in[249] net[249] vdd gnd pnand2_4
Xwl_driver_inv249 net[249] wl[249] vdd gnd pinv_11
Xwl_driver_inv_en250 en en_bar[250] vdd gnd pinv_12
Xwl_driver_nand250 en_bar[250] in[250] net[250] vdd gnd pnand2_4
Xwl_driver_inv250 net[250] wl[250] vdd gnd pinv_11
Xwl_driver_inv_en251 en en_bar[251] vdd gnd pinv_12
Xwl_driver_nand251 en_bar[251] in[251] net[251] vdd gnd pnand2_4
Xwl_driver_inv251 net[251] wl[251] vdd gnd pinv_11
Xwl_driver_inv_en252 en en_bar[252] vdd gnd pinv_12
Xwl_driver_nand252 en_bar[252] in[252] net[252] vdd gnd pnand2_4
Xwl_driver_inv252 net[252] wl[252] vdd gnd pinv_11
Xwl_driver_inv_en253 en en_bar[253] vdd gnd pinv_12
Xwl_driver_nand253 en_bar[253] in[253] net[253] vdd gnd pnand2_4
Xwl_driver_inv253 net[253] wl[253] vdd gnd pinv_11
Xwl_driver_inv_en254 en en_bar[254] vdd gnd pinv_12
Xwl_driver_nand254 en_bar[254] in[254] net[254] vdd gnd pnand2_4
Xwl_driver_inv254 net[254] wl[254] vdd gnd pinv_11
Xwl_driver_inv_en255 en en_bar[255] vdd gnd pinv_12
Xwl_driver_nand255 en_bar[255] in[255] net[255] vdd gnd pnand2_4
Xwl_driver_inv255 net[255] wl[255] vdd gnd pinv_11
.ENDS wordline_driver

.SUBCKT pinv_13 A Z vdd gnd
Mpinv_pmos Z A vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpinv_nmos Z A gnd gnd n m=1 w=1.2u l=0.6u pd=3.6u ps=3.6u as=1.8p ad=1.8p
.ENDS pinv_13

.SUBCKT pinv_14 A Z vdd gnd
Mpinv_pmos Z A vdd vdd p m=3 w=3.15u l=0.6u pd=7.5u ps=7.5u as=4.725p ad=4.725p
Mpinv_nmos Z A gnd gnd n m=3 w=1.65u l=0.6u pd=4.5u ps=4.5u as=2.475p ad=2.475p
.ENDS pinv_14

.SUBCKT pnor2_2 A B Z vdd gnd
Mpnor2_pmos1 vdd A net1 vdd p m=1 w=3.6u l=0.6u pd=8.4u ps=8.4u as=5.4p ad=5.4p
Mpnor2_pmos2 net1 B Z vdd p m=1 w=3.6u l=0.6u pd=8.4u ps=8.4u as=5.4p ad=5.4p
Mpnor2_nmos1 Z A gnd gnd n m=1 w=1.2u l=0.6u pd=3.6u ps=3.6u as=1.8p ad=1.8p
Mpnor2_nmos2 Z B gnd gnd n m=1 w=1.2u l=0.6u pd=3.6u ps=3.6u as=1.8p ad=1.8p
.ENDS pnor2_2

.SUBCKT pnand2_5 A B Z vdd gnd
Mpnand2_pmos1 vdd A Z vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand2_pmos2 Z B vdd vdd p m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand2_nmos1 Z B net1 gnd n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
Mpnand2_nmos2 net1 A gnd gnd n m=1 w=2.4u l=0.6u pd=6.0u ps=6.0u as=3.6p ad=3.6p
.ENDS pnand2_5

.SUBCKT bank DATA[0] DATA[1] DATA[2] DATA[3] DATA[4] DATA[5] DATA[6] DATA[7] DATA[8] DATA[9] DATA[10] DATA[11] DATA[12] DATA[13] DATA[14] DATA[15] DATA[16] DATA[17] DATA[18] DATA[19] DATA[20] DATA[21] DATA[22] DATA[23] DATA[24] DATA[25] DATA[26] DATA[27] DATA[28] DATA[29] DATA[30] DATA[31] DATA[32] DATA[33] DATA[34] DATA[35] DATA[36] DATA[37] DATA[38] DATA[39] DATA[40] DATA[41] DATA[42] DATA[43] DATA[44] DATA[45] DATA[46] DATA[47] DATA[48] DATA[49] DATA[50] DATA[51] DATA[52] DATA[53] DATA[54] DATA[55] DATA[56] DATA[57] DATA[58] DATA[59] DATA[60] DATA[61] DATA[62] DATA[63] DATA[64] DATA[65] DATA[66] DATA[67] DATA[68] DATA[69] DATA[70] DATA[71] DATA[72] DATA[73] DATA[74] DATA[75] DATA[76] DATA[77] DATA[78] DATA[79] DATA[80] DATA[81] DATA[82] DATA[83] DATA[84] DATA[85] DATA[86] DATA[87] DATA[88] DATA[89] DATA[90] DATA[91] DATA[92] DATA[93] DATA[94] DATA[95] DATA[96] DATA[97] DATA[98] DATA[99] DATA[100] DATA[101] DATA[102] DATA[103] DATA[104] DATA[105] DATA[106] DATA[107] DATA[108] DATA[109] DATA[110] DATA[111] DATA[112] DATA[113] DATA[114] DATA[115] DATA[116] DATA[117] DATA[118] DATA[119] DATA[120] DATA[121] DATA[122] DATA[123] DATA[124] DATA[125] DATA[126] DATA[127] ADDR[0] ADDR[1] ADDR[2] ADDR[3] ADDR[4] ADDR[5] ADDR[6] ADDR[7] ADDR[8] bank_sel s_en w_en tri_en_bar tri_en clk_bar clk_buf vdd gnd
Xbitcell_array bl[0] br[0] bl[1] br[1] bl[2] br[2] bl[3] br[3] bl[4] br[4] bl[5] br[5] bl[6] br[6] bl[7] br[7] bl[8] br[8] bl[9] br[9] bl[10] br[10] bl[11] br[11] bl[12] br[12] bl[13] br[13] bl[14] br[14] bl[15] br[15] bl[16] br[16] bl[17] br[17] bl[18] br[18] bl[19] br[19] bl[20] br[20] bl[21] br[21] bl[22] br[22] bl[23] br[23] bl[24] br[24] bl[25] br[25] bl[26] br[26] bl[27] br[27] bl[28] br[28] bl[29] br[29] bl[30] br[30] bl[31] br[31] bl[32] br[32] bl[33] br[33] bl[34] br[34] bl[35] br[35] bl[36] br[36] bl[37] br[37] bl[38] br[38] bl[39] br[39] bl[40] br[40] bl[41] br[41] bl[42] br[42] bl[43] br[43] bl[44] br[44] bl[45] br[45] bl[46] br[46] bl[47] br[47] bl[48] br[48] bl[49] br[49] bl[50] br[50] bl[51] br[51] bl[52] br[52] bl[53] br[53] bl[54] br[54] bl[55] br[55] bl[56] br[56] bl[57] br[57] bl[58] br[58] bl[59] br[59] bl[60] br[60] bl[61] br[61] bl[62] br[62] bl[63] br[63] bl[64] br[64] bl[65] br[65] bl[66] br[66] bl[67] br[67] bl[68] br[68] bl[69] br[69] bl[70] br[70] bl[71] br[71] bl[72] br[72] bl[73] br[73] bl[74] br[74] bl[75] br[75] bl[76] br[76] bl[77] br[77] bl[78] br[78] bl[79] br[79] bl[80] br[80] bl[81] br[81] bl[82] br[82] bl[83] br[83] bl[84] br[84] bl[85] br[85] bl[86] br[86] bl[87] br[87] bl[88] br[88] bl[89] br[89] bl[90] br[90] bl[91] br[91] bl[92] br[92] bl[93] br[93] bl[94] br[94] bl[95] br[95] bl[96] br[96] bl[97] br[97] bl[98] br[98] bl[99] br[99] bl[100] br[100] bl[101] br[101] bl[102] br[102] bl[103] br[103] bl[104] br[104] bl[105] br[105] bl[106] br[106] bl[107] br[107] bl[108] br[108] bl[109] br[109] bl[110] br[110] bl[111] br[111] bl[112] br[112] bl[113] br[113] bl[114] br[114] bl[115] br[115] bl[116] br[116] bl[117] br[117] bl[118] br[118] bl[119] br[119] bl[120] br[120] bl[121] br[121] bl[122] br[122] bl[123] br[123] bl[124] br[124] bl[125] br[125] bl[126] br[126] bl[127] br[127] bl[128] br[128] bl[129] br[129] bl[130] br[130] bl[131] br[131] bl[132] br[132] bl[133] br[133] bl[134] br[134] bl[135] br[135] bl[136] br[136] bl[137] br[137] bl[138] br[138] bl[139] br[139] bl[140] br[140] bl[141] br[141] bl[142] br[142] bl[143] br[143] bl[144] br[144] bl[145] br[145] bl[146] br[146] bl[147] br[147] bl[148] br[148] bl[149] br[149] bl[150] br[150] bl[151] br[151] bl[152] br[152] bl[153] br[153] bl[154] br[154] bl[155] br[155] bl[156] br[156] bl[157] br[157] bl[158] br[158] bl[159] br[159] bl[160] br[160] bl[161] br[161] bl[162] br[162] bl[163] br[163] bl[164] br[164] bl[165] br[165] bl[166] br[166] bl[167] br[167] bl[168] br[168] bl[169] br[169] bl[170] br[170] bl[171] br[171] bl[172] br[172] bl[173] br[173] bl[174] br[174] bl[175] br[175] bl[176] br[176] bl[177] br[177] bl[178] br[178] bl[179] br[179] bl[180] br[180] bl[181] br[181] bl[182] br[182] bl[183] br[183] bl[184] br[184] bl[185] br[185] bl[186] br[186] bl[187] br[187] bl[188] br[188] bl[189] br[189] bl[190] br[190] bl[191] br[191] bl[192] br[192] bl[193] br[193] bl[194] br[194] bl[195] br[195] bl[196] br[196] bl[197] br[197] bl[198] br[198] bl[199] br[199] bl[200] br[200] bl[201] br[201] bl[202] br[202] bl[203] br[203] bl[204] br[204] bl[205] br[205] bl[206] br[206] bl[207] br[207] bl[208] br[208] bl[209] br[209] bl[210] br[210] bl[211] br[211] bl[212] br[212] bl[213] br[213] bl[214] br[214] bl[215] br[215] bl[216] br[216] bl[217] br[217] bl[218] br[218] bl[219] br[219] bl[220] br[220] bl[221] br[221] bl[222] br[222] bl[223] br[223] bl[224] br[224] bl[225] br[225] bl[226] br[226] bl[227] br[227] bl[228] br[228] bl[229] br[229] bl[230] br[230] bl[231] br[231] bl[232] br[232] bl[233] br[233] bl[234] br[234] bl[235] br[235] bl[236] br[236] bl[237] br[237] bl[238] br[238] bl[239] br[239] bl[240] br[240] bl[241] br[241] bl[242] br[242] bl[243] br[243] bl[244] br[244] bl[245] br[245] bl[246] br[246] bl[247] br[247] bl[248] br[248] bl[249] br[249] bl[250] br[250] bl[251] br[251] bl[252] br[252] bl[253] br[253] bl[254] br[254] bl[255] br[255] wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] wl[128] wl[129] wl[130] wl[131] wl[132] wl[133] wl[134] wl[135] wl[136] wl[137] wl[138] wl[139] wl[140] wl[141] wl[142] wl[143] wl[144] wl[145] wl[146] wl[147] wl[148] wl[149] wl[150] wl[151] wl[152] wl[153] wl[154] wl[155] wl[156] wl[157] wl[158] wl[159] wl[160] wl[161] wl[162] wl[163] wl[164] wl[165] wl[166] wl[167] wl[168] wl[169] wl[170] wl[171] wl[172] wl[173] wl[174] wl[175] wl[176] wl[177] wl[178] wl[179] wl[180] wl[181] wl[182] wl[183] wl[184] wl[185] wl[186] wl[187] wl[188] wl[189] wl[190] wl[191] wl[192] wl[193] wl[194] wl[195] wl[196] wl[197] wl[198] wl[199] wl[200] wl[201] wl[202] wl[203] wl[204] wl[205] wl[206] wl[207] wl[208] wl[209] wl[210] wl[211] wl[212] wl[213] wl[214] wl[215] wl[216] wl[217] wl[218] wl[219] wl[220] wl[221] wl[222] wl[223] wl[224] wl[225] wl[226] wl[227] wl[228] wl[229] wl[230] wl[231] wl[232] wl[233] wl[234] wl[235] wl[236] wl[237] wl[238] wl[239] wl[240] wl[241] wl[242] wl[243] wl[244] wl[245] wl[246] wl[247] wl[248] wl[249] wl[250] wl[251] wl[252] wl[253] wl[254] wl[255] vdd gnd bitcell_array
Xprecharge_array bl[0] br[0] bl[1] br[1] bl[2] br[2] bl[3] br[3] bl[4] br[4] bl[5] br[5] bl[6] br[6] bl[7] br[7] bl[8] br[8] bl[9] br[9] bl[10] br[10] bl[11] br[11] bl[12] br[12] bl[13] br[13] bl[14] br[14] bl[15] br[15] bl[16] br[16] bl[17] br[17] bl[18] br[18] bl[19] br[19] bl[20] br[20] bl[21] br[21] bl[22] br[22] bl[23] br[23] bl[24] br[24] bl[25] br[25] bl[26] br[26] bl[27] br[27] bl[28] br[28] bl[29] br[29] bl[30] br[30] bl[31] br[31] bl[32] br[32] bl[33] br[33] bl[34] br[34] bl[35] br[35] bl[36] br[36] bl[37] br[37] bl[38] br[38] bl[39] br[39] bl[40] br[40] bl[41] br[41] bl[42] br[42] bl[43] br[43] bl[44] br[44] bl[45] br[45] bl[46] br[46] bl[47] br[47] bl[48] br[48] bl[49] br[49] bl[50] br[50] bl[51] br[51] bl[52] br[52] bl[53] br[53] bl[54] br[54] bl[55] br[55] bl[56] br[56] bl[57] br[57] bl[58] br[58] bl[59] br[59] bl[60] br[60] bl[61] br[61] bl[62] br[62] bl[63] br[63] bl[64] br[64] bl[65] br[65] bl[66] br[66] bl[67] br[67] bl[68] br[68] bl[69] br[69] bl[70] br[70] bl[71] br[71] bl[72] br[72] bl[73] br[73] bl[74] br[74] bl[75] br[75] bl[76] br[76] bl[77] br[77] bl[78] br[78] bl[79] br[79] bl[80] br[80] bl[81] br[81] bl[82] br[82] bl[83] br[83] bl[84] br[84] bl[85] br[85] bl[86] br[86] bl[87] br[87] bl[88] br[88] bl[89] br[89] bl[90] br[90] bl[91] br[91] bl[92] br[92] bl[93] br[93] bl[94] br[94] bl[95] br[95] bl[96] br[96] bl[97] br[97] bl[98] br[98] bl[99] br[99] bl[100] br[100] bl[101] br[101] bl[102] br[102] bl[103] br[103] bl[104] br[104] bl[105] br[105] bl[106] br[106] bl[107] br[107] bl[108] br[108] bl[109] br[109] bl[110] br[110] bl[111] br[111] bl[112] br[112] bl[113] br[113] bl[114] br[114] bl[115] br[115] bl[116] br[116] bl[117] br[117] bl[118] br[118] bl[119] br[119] bl[120] br[120] bl[121] br[121] bl[122] br[122] bl[123] br[123] bl[124] br[124] bl[125] br[125] bl[126] br[126] bl[127] br[127] bl[128] br[128] bl[129] br[129] bl[130] br[130] bl[131] br[131] bl[132] br[132] bl[133] br[133] bl[134] br[134] bl[135] br[135] bl[136] br[136] bl[137] br[137] bl[138] br[138] bl[139] br[139] bl[140] br[140] bl[141] br[141] bl[142] br[142] bl[143] br[143] bl[144] br[144] bl[145] br[145] bl[146] br[146] bl[147] br[147] bl[148] br[148] bl[149] br[149] bl[150] br[150] bl[151] br[151] bl[152] br[152] bl[153] br[153] bl[154] br[154] bl[155] br[155] bl[156] br[156] bl[157] br[157] bl[158] br[158] bl[159] br[159] bl[160] br[160] bl[161] br[161] bl[162] br[162] bl[163] br[163] bl[164] br[164] bl[165] br[165] bl[166] br[166] bl[167] br[167] bl[168] br[168] bl[169] br[169] bl[170] br[170] bl[171] br[171] bl[172] br[172] bl[173] br[173] bl[174] br[174] bl[175] br[175] bl[176] br[176] bl[177] br[177] bl[178] br[178] bl[179] br[179] bl[180] br[180] bl[181] br[181] bl[182] br[182] bl[183] br[183] bl[184] br[184] bl[185] br[185] bl[186] br[186] bl[187] br[187] bl[188] br[188] bl[189] br[189] bl[190] br[190] bl[191] br[191] bl[192] br[192] bl[193] br[193] bl[194] br[194] bl[195] br[195] bl[196] br[196] bl[197] br[197] bl[198] br[198] bl[199] br[199] bl[200] br[200] bl[201] br[201] bl[202] br[202] bl[203] br[203] bl[204] br[204] bl[205] br[205] bl[206] br[206] bl[207] br[207] bl[208] br[208] bl[209] br[209] bl[210] br[210] bl[211] br[211] bl[212] br[212] bl[213] br[213] bl[214] br[214] bl[215] br[215] bl[216] br[216] bl[217] br[217] bl[218] br[218] bl[219] br[219] bl[220] br[220] bl[221] br[221] bl[222] br[222] bl[223] br[223] bl[224] br[224] bl[225] br[225] bl[226] br[226] bl[227] br[227] bl[228] br[228] bl[229] br[229] bl[230] br[230] bl[231] br[231] bl[232] br[232] bl[233] br[233] bl[234] br[234] bl[235] br[235] bl[236] br[236] bl[237] br[237] bl[238] br[238] bl[239] br[239] bl[240] br[240] bl[241] br[241] bl[242] br[242] bl[243] br[243] bl[244] br[244] bl[245] br[245] bl[246] br[246] bl[247] br[247] bl[248] br[248] bl[249] br[249] bl[250] br[250] bl[251] br[251] bl[252] br[252] bl[253] br[253] bl[254] br[254] bl[255] br[255] gated_clk_bar vdd precharge_array
Xcolumn_mux_array bl[0] br[0] bl[1] br[1] bl[2] br[2] bl[3] br[3] bl[4] br[4] bl[5] br[5] bl[6] br[6] bl[7] br[7] bl[8] br[8] bl[9] br[9] bl[10] br[10] bl[11] br[11] bl[12] br[12] bl[13] br[13] bl[14] br[14] bl[15] br[15] bl[16] br[16] bl[17] br[17] bl[18] br[18] bl[19] br[19] bl[20] br[20] bl[21] br[21] bl[22] br[22] bl[23] br[23] bl[24] br[24] bl[25] br[25] bl[26] br[26] bl[27] br[27] bl[28] br[28] bl[29] br[29] bl[30] br[30] bl[31] br[31] bl[32] br[32] bl[33] br[33] bl[34] br[34] bl[35] br[35] bl[36] br[36] bl[37] br[37] bl[38] br[38] bl[39] br[39] bl[40] br[40] bl[41] br[41] bl[42] br[42] bl[43] br[43] bl[44] br[44] bl[45] br[45] bl[46] br[46] bl[47] br[47] bl[48] br[48] bl[49] br[49] bl[50] br[50] bl[51] br[51] bl[52] br[52] bl[53] br[53] bl[54] br[54] bl[55] br[55] bl[56] br[56] bl[57] br[57] bl[58] br[58] bl[59] br[59] bl[60] br[60] bl[61] br[61] bl[62] br[62] bl[63] br[63] bl[64] br[64] bl[65] br[65] bl[66] br[66] bl[67] br[67] bl[68] br[68] bl[69] br[69] bl[70] br[70] bl[71] br[71] bl[72] br[72] bl[73] br[73] bl[74] br[74] bl[75] br[75] bl[76] br[76] bl[77] br[77] bl[78] br[78] bl[79] br[79] bl[80] br[80] bl[81] br[81] bl[82] br[82] bl[83] br[83] bl[84] br[84] bl[85] br[85] bl[86] br[86] bl[87] br[87] bl[88] br[88] bl[89] br[89] bl[90] br[90] bl[91] br[91] bl[92] br[92] bl[93] br[93] bl[94] br[94] bl[95] br[95] bl[96] br[96] bl[97] br[97] bl[98] br[98] bl[99] br[99] bl[100] br[100] bl[101] br[101] bl[102] br[102] bl[103] br[103] bl[104] br[104] bl[105] br[105] bl[106] br[106] bl[107] br[107] bl[108] br[108] bl[109] br[109] bl[110] br[110] bl[111] br[111] bl[112] br[112] bl[113] br[113] bl[114] br[114] bl[115] br[115] bl[116] br[116] bl[117] br[117] bl[118] br[118] bl[119] br[119] bl[120] br[120] bl[121] br[121] bl[122] br[122] bl[123] br[123] bl[124] br[124] bl[125] br[125] bl[126] br[126] bl[127] br[127] bl[128] br[128] bl[129] br[129] bl[130] br[130] bl[131] br[131] bl[132] br[132] bl[133] br[133] bl[134] br[134] bl[135] br[135] bl[136] br[136] bl[137] br[137] bl[138] br[138] bl[139] br[139] bl[140] br[140] bl[141] br[141] bl[142] br[142] bl[143] br[143] bl[144] br[144] bl[145] br[145] bl[146] br[146] bl[147] br[147] bl[148] br[148] bl[149] br[149] bl[150] br[150] bl[151] br[151] bl[152] br[152] bl[153] br[153] bl[154] br[154] bl[155] br[155] bl[156] br[156] bl[157] br[157] bl[158] br[158] bl[159] br[159] bl[160] br[160] bl[161] br[161] bl[162] br[162] bl[163] br[163] bl[164] br[164] bl[165] br[165] bl[166] br[166] bl[167] br[167] bl[168] br[168] bl[169] br[169] bl[170] br[170] bl[171] br[171] bl[172] br[172] bl[173] br[173] bl[174] br[174] bl[175] br[175] bl[176] br[176] bl[177] br[177] bl[178] br[178] bl[179] br[179] bl[180] br[180] bl[181] br[181] bl[182] br[182] bl[183] br[183] bl[184] br[184] bl[185] br[185] bl[186] br[186] bl[187] br[187] bl[188] br[188] bl[189] br[189] bl[190] br[190] bl[191] br[191] bl[192] br[192] bl[193] br[193] bl[194] br[194] bl[195] br[195] bl[196] br[196] bl[197] br[197] bl[198] br[198] bl[199] br[199] bl[200] br[200] bl[201] br[201] bl[202] br[202] bl[203] br[203] bl[204] br[204] bl[205] br[205] bl[206] br[206] bl[207] br[207] bl[208] br[208] bl[209] br[209] bl[210] br[210] bl[211] br[211] bl[212] br[212] bl[213] br[213] bl[214] br[214] bl[215] br[215] bl[216] br[216] bl[217] br[217] bl[218] br[218] bl[219] br[219] bl[220] br[220] bl[221] br[221] bl[222] br[222] bl[223] br[223] bl[224] br[224] bl[225] br[225] bl[226] br[226] bl[227] br[227] bl[228] br[228] bl[229] br[229] bl[230] br[230] bl[231] br[231] bl[232] br[232] bl[233] br[233] bl[234] br[234] bl[235] br[235] bl[236] br[236] bl[237] br[237] bl[238] br[238] bl[239] br[239] bl[240] br[240] bl[241] br[241] bl[242] br[242] bl[243] br[243] bl[244] br[244] bl[245] br[245] bl[246] br[246] bl[247] br[247] bl[248] br[248] bl[249] br[249] bl[250] br[250] bl[251] br[251] bl[252] br[252] bl[253] br[253] bl[254] br[254] bl[255] br[255] sel[0] sel[1] bl_out[0] br_out[0] bl_out[1] br_out[1] bl_out[2] br_out[2] bl_out[3] br_out[3] bl_out[4] br_out[4] bl_out[5] br_out[5] bl_out[6] br_out[6] bl_out[7] br_out[7] bl_out[8] br_out[8] bl_out[9] br_out[9] bl_out[10] br_out[10] bl_out[11] br_out[11] bl_out[12] br_out[12] bl_out[13] br_out[13] bl_out[14] br_out[14] bl_out[15] br_out[15] bl_out[16] br_out[16] bl_out[17] br_out[17] bl_out[18] br_out[18] bl_out[19] br_out[19] bl_out[20] br_out[20] bl_out[21] br_out[21] bl_out[22] br_out[22] bl_out[23] br_out[23] bl_out[24] br_out[24] bl_out[25] br_out[25] bl_out[26] br_out[26] bl_out[27] br_out[27] bl_out[28] br_out[28] bl_out[29] br_out[29] bl_out[30] br_out[30] bl_out[31] br_out[31] bl_out[32] br_out[32] bl_out[33] br_out[33] bl_out[34] br_out[34] bl_out[35] br_out[35] bl_out[36] br_out[36] bl_out[37] br_out[37] bl_out[38] br_out[38] bl_out[39] br_out[39] bl_out[40] br_out[40] bl_out[41] br_out[41] bl_out[42] br_out[42] bl_out[43] br_out[43] bl_out[44] br_out[44] bl_out[45] br_out[45] bl_out[46] br_out[46] bl_out[47] br_out[47] bl_out[48] br_out[48] bl_out[49] br_out[49] bl_out[50] br_out[50] bl_out[51] br_out[51] bl_out[52] br_out[52] bl_out[53] br_out[53] bl_out[54] br_out[54] bl_out[55] br_out[55] bl_out[56] br_out[56] bl_out[57] br_out[57] bl_out[58] br_out[58] bl_out[59] br_out[59] bl_out[60] br_out[60] bl_out[61] br_out[61] bl_out[62] br_out[62] bl_out[63] br_out[63] bl_out[64] br_out[64] bl_out[65] br_out[65] bl_out[66] br_out[66] bl_out[67] br_out[67] bl_out[68] br_out[68] bl_out[69] br_out[69] bl_out[70] br_out[70] bl_out[71] br_out[71] bl_out[72] br_out[72] bl_out[73] br_out[73] bl_out[74] br_out[74] bl_out[75] br_out[75] bl_out[76] br_out[76] bl_out[77] br_out[77] bl_out[78] br_out[78] bl_out[79] br_out[79] bl_out[80] br_out[80] bl_out[81] br_out[81] bl_out[82] br_out[82] bl_out[83] br_out[83] bl_out[84] br_out[84] bl_out[85] br_out[85] bl_out[86] br_out[86] bl_out[87] br_out[87] bl_out[88] br_out[88] bl_out[89] br_out[89] bl_out[90] br_out[90] bl_out[91] br_out[91] bl_out[92] br_out[92] bl_out[93] br_out[93] bl_out[94] br_out[94] bl_out[95] br_out[95] bl_out[96] br_out[96] bl_out[97] br_out[97] bl_out[98] br_out[98] bl_out[99] br_out[99] bl_out[100] br_out[100] bl_out[101] br_out[101] bl_out[102] br_out[102] bl_out[103] br_out[103] bl_out[104] br_out[104] bl_out[105] br_out[105] bl_out[106] br_out[106] bl_out[107] br_out[107] bl_out[108] br_out[108] bl_out[109] br_out[109] bl_out[110] br_out[110] bl_out[111] br_out[111] bl_out[112] br_out[112] bl_out[113] br_out[113] bl_out[114] br_out[114] bl_out[115] br_out[115] bl_out[116] br_out[116] bl_out[117] br_out[117] bl_out[118] br_out[118] bl_out[119] br_out[119] bl_out[120] br_out[120] bl_out[121] br_out[121] bl_out[122] br_out[122] bl_out[123] br_out[123] bl_out[124] br_out[124] bl_out[125] br_out[125] bl_out[126] br_out[126] bl_out[127] br_out[127] gnd columnmux_array
Xsense_amp_array data_out[0] bl_out[0] br_out[0] data_out[1] bl_out[1] br_out[1] data_out[2] bl_out[2] br_out[2] data_out[3] bl_out[3] br_out[3] data_out[4] bl_out[4] br_out[4] data_out[5] bl_out[5] br_out[5] data_out[6] bl_out[6] br_out[6] data_out[7] bl_out[7] br_out[7] data_out[8] bl_out[8] br_out[8] data_out[9] bl_out[9] br_out[9] data_out[10] bl_out[10] br_out[10] data_out[11] bl_out[11] br_out[11] data_out[12] bl_out[12] br_out[12] data_out[13] bl_out[13] br_out[13] data_out[14] bl_out[14] br_out[14] data_out[15] bl_out[15] br_out[15] data_out[16] bl_out[16] br_out[16] data_out[17] bl_out[17] br_out[17] data_out[18] bl_out[18] br_out[18] data_out[19] bl_out[19] br_out[19] data_out[20] bl_out[20] br_out[20] data_out[21] bl_out[21] br_out[21] data_out[22] bl_out[22] br_out[22] data_out[23] bl_out[23] br_out[23] data_out[24] bl_out[24] br_out[24] data_out[25] bl_out[25] br_out[25] data_out[26] bl_out[26] br_out[26] data_out[27] bl_out[27] br_out[27] data_out[28] bl_out[28] br_out[28] data_out[29] bl_out[29] br_out[29] data_out[30] bl_out[30] br_out[30] data_out[31] bl_out[31] br_out[31] data_out[32] bl_out[32] br_out[32] data_out[33] bl_out[33] br_out[33] data_out[34] bl_out[34] br_out[34] data_out[35] bl_out[35] br_out[35] data_out[36] bl_out[36] br_out[36] data_out[37] bl_out[37] br_out[37] data_out[38] bl_out[38] br_out[38] data_out[39] bl_out[39] br_out[39] data_out[40] bl_out[40] br_out[40] data_out[41] bl_out[41] br_out[41] data_out[42] bl_out[42] br_out[42] data_out[43] bl_out[43] br_out[43] data_out[44] bl_out[44] br_out[44] data_out[45] bl_out[45] br_out[45] data_out[46] bl_out[46] br_out[46] data_out[47] bl_out[47] br_out[47] data_out[48] bl_out[48] br_out[48] data_out[49] bl_out[49] br_out[49] data_out[50] bl_out[50] br_out[50] data_out[51] bl_out[51] br_out[51] data_out[52] bl_out[52] br_out[52] data_out[53] bl_out[53] br_out[53] data_out[54] bl_out[54] br_out[54] data_out[55] bl_out[55] br_out[55] data_out[56] bl_out[56] br_out[56] data_out[57] bl_out[57] br_out[57] data_out[58] bl_out[58] br_out[58] data_out[59] bl_out[59] br_out[59] data_out[60] bl_out[60] br_out[60] data_out[61] bl_out[61] br_out[61] data_out[62] bl_out[62] br_out[62] data_out[63] bl_out[63] br_out[63] data_out[64] bl_out[64] br_out[64] data_out[65] bl_out[65] br_out[65] data_out[66] bl_out[66] br_out[66] data_out[67] bl_out[67] br_out[67] data_out[68] bl_out[68] br_out[68] data_out[69] bl_out[69] br_out[69] data_out[70] bl_out[70] br_out[70] data_out[71] bl_out[71] br_out[71] data_out[72] bl_out[72] br_out[72] data_out[73] bl_out[73] br_out[73] data_out[74] bl_out[74] br_out[74] data_out[75] bl_out[75] br_out[75] data_out[76] bl_out[76] br_out[76] data_out[77] bl_out[77] br_out[77] data_out[78] bl_out[78] br_out[78] data_out[79] bl_out[79] br_out[79] data_out[80] bl_out[80] br_out[80] data_out[81] bl_out[81] br_out[81] data_out[82] bl_out[82] br_out[82] data_out[83] bl_out[83] br_out[83] data_out[84] bl_out[84] br_out[84] data_out[85] bl_out[85] br_out[85] data_out[86] bl_out[86] br_out[86] data_out[87] bl_out[87] br_out[87] data_out[88] bl_out[88] br_out[88] data_out[89] bl_out[89] br_out[89] data_out[90] bl_out[90] br_out[90] data_out[91] bl_out[91] br_out[91] data_out[92] bl_out[92] br_out[92] data_out[93] bl_out[93] br_out[93] data_out[94] bl_out[94] br_out[94] data_out[95] bl_out[95] br_out[95] data_out[96] bl_out[96] br_out[96] data_out[97] bl_out[97] br_out[97] data_out[98] bl_out[98] br_out[98] data_out[99] bl_out[99] br_out[99] data_out[100] bl_out[100] br_out[100] data_out[101] bl_out[101] br_out[101] data_out[102] bl_out[102] br_out[102] data_out[103] bl_out[103] br_out[103] data_out[104] bl_out[104] br_out[104] data_out[105] bl_out[105] br_out[105] data_out[106] bl_out[106] br_out[106] data_out[107] bl_out[107] br_out[107] data_out[108] bl_out[108] br_out[108] data_out[109] bl_out[109] br_out[109] data_out[110] bl_out[110] br_out[110] data_out[111] bl_out[111] br_out[111] data_out[112] bl_out[112] br_out[112] data_out[113] bl_out[113] br_out[113] data_out[114] bl_out[114] br_out[114] data_out[115] bl_out[115] br_out[115] data_out[116] bl_out[116] br_out[116] data_out[117] bl_out[117] br_out[117] data_out[118] bl_out[118] br_out[118] data_out[119] bl_out[119] br_out[119] data_out[120] bl_out[120] br_out[120] data_out[121] bl_out[121] br_out[121] data_out[122] bl_out[122] br_out[122] data_out[123] bl_out[123] br_out[123] data_out[124] bl_out[124] br_out[124] data_out[125] bl_out[125] br_out[125] data_out[126] bl_out[126] br_out[126] data_out[127] bl_out[127] br_out[127] gated_s_en vdd gnd sense_amp_array
Xwrite_driver_array data_in[0] data_in[1] data_in[2] data_in[3] data_in[4] data_in[5] data_in[6] data_in[7] data_in[8] data_in[9] data_in[10] data_in[11] data_in[12] data_in[13] data_in[14] data_in[15] data_in[16] data_in[17] data_in[18] data_in[19] data_in[20] data_in[21] data_in[22] data_in[23] data_in[24] data_in[25] data_in[26] data_in[27] data_in[28] data_in[29] data_in[30] data_in[31] data_in[32] data_in[33] data_in[34] data_in[35] data_in[36] data_in[37] data_in[38] data_in[39] data_in[40] data_in[41] data_in[42] data_in[43] data_in[44] data_in[45] data_in[46] data_in[47] data_in[48] data_in[49] data_in[50] data_in[51] data_in[52] data_in[53] data_in[54] data_in[55] data_in[56] data_in[57] data_in[58] data_in[59] data_in[60] data_in[61] data_in[62] data_in[63] data_in[64] data_in[65] data_in[66] data_in[67] data_in[68] data_in[69] data_in[70] data_in[71] data_in[72] data_in[73] data_in[74] data_in[75] data_in[76] data_in[77] data_in[78] data_in[79] data_in[80] data_in[81] data_in[82] data_in[83] data_in[84] data_in[85] data_in[86] data_in[87] data_in[88] data_in[89] data_in[90] data_in[91] data_in[92] data_in[93] data_in[94] data_in[95] data_in[96] data_in[97] data_in[98] data_in[99] data_in[100] data_in[101] data_in[102] data_in[103] data_in[104] data_in[105] data_in[106] data_in[107] data_in[108] data_in[109] data_in[110] data_in[111] data_in[112] data_in[113] data_in[114] data_in[115] data_in[116] data_in[117] data_in[118] data_in[119] data_in[120] data_in[121] data_in[122] data_in[123] data_in[124] data_in[125] data_in[126] data_in[127] bl_out[0] br_out[0] bl_out[1] br_out[1] bl_out[2] br_out[2] bl_out[3] br_out[3] bl_out[4] br_out[4] bl_out[5] br_out[5] bl_out[6] br_out[6] bl_out[7] br_out[7] bl_out[8] br_out[8] bl_out[9] br_out[9] bl_out[10] br_out[10] bl_out[11] br_out[11] bl_out[12] br_out[12] bl_out[13] br_out[13] bl_out[14] br_out[14] bl_out[15] br_out[15] bl_out[16] br_out[16] bl_out[17] br_out[17] bl_out[18] br_out[18] bl_out[19] br_out[19] bl_out[20] br_out[20] bl_out[21] br_out[21] bl_out[22] br_out[22] bl_out[23] br_out[23] bl_out[24] br_out[24] bl_out[25] br_out[25] bl_out[26] br_out[26] bl_out[27] br_out[27] bl_out[28] br_out[28] bl_out[29] br_out[29] bl_out[30] br_out[30] bl_out[31] br_out[31] bl_out[32] br_out[32] bl_out[33] br_out[33] bl_out[34] br_out[34] bl_out[35] br_out[35] bl_out[36] br_out[36] bl_out[37] br_out[37] bl_out[38] br_out[38] bl_out[39] br_out[39] bl_out[40] br_out[40] bl_out[41] br_out[41] bl_out[42] br_out[42] bl_out[43] br_out[43] bl_out[44] br_out[44] bl_out[45] br_out[45] bl_out[46] br_out[46] bl_out[47] br_out[47] bl_out[48] br_out[48] bl_out[49] br_out[49] bl_out[50] br_out[50] bl_out[51] br_out[51] bl_out[52] br_out[52] bl_out[53] br_out[53] bl_out[54] br_out[54] bl_out[55] br_out[55] bl_out[56] br_out[56] bl_out[57] br_out[57] bl_out[58] br_out[58] bl_out[59] br_out[59] bl_out[60] br_out[60] bl_out[61] br_out[61] bl_out[62] br_out[62] bl_out[63] br_out[63] bl_out[64] br_out[64] bl_out[65] br_out[65] bl_out[66] br_out[66] bl_out[67] br_out[67] bl_out[68] br_out[68] bl_out[69] br_out[69] bl_out[70] br_out[70] bl_out[71] br_out[71] bl_out[72] br_out[72] bl_out[73] br_out[73] bl_out[74] br_out[74] bl_out[75] br_out[75] bl_out[76] br_out[76] bl_out[77] br_out[77] bl_out[78] br_out[78] bl_out[79] br_out[79] bl_out[80] br_out[80] bl_out[81] br_out[81] bl_out[82] br_out[82] bl_out[83] br_out[83] bl_out[84] br_out[84] bl_out[85] br_out[85] bl_out[86] br_out[86] bl_out[87] br_out[87] bl_out[88] br_out[88] bl_out[89] br_out[89] bl_out[90] br_out[90] bl_out[91] br_out[91] bl_out[92] br_out[92] bl_out[93] br_out[93] bl_out[94] br_out[94] bl_out[95] br_out[95] bl_out[96] br_out[96] bl_out[97] br_out[97] bl_out[98] br_out[98] bl_out[99] br_out[99] bl_out[100] br_out[100] bl_out[101] br_out[101] bl_out[102] br_out[102] bl_out[103] br_out[103] bl_out[104] br_out[104] bl_out[105] br_out[105] bl_out[106] br_out[106] bl_out[107] br_out[107] bl_out[108] br_out[108] bl_out[109] br_out[109] bl_out[110] br_out[110] bl_out[111] br_out[111] bl_out[112] br_out[112] bl_out[113] br_out[113] bl_out[114] br_out[114] bl_out[115] br_out[115] bl_out[116] br_out[116] bl_out[117] br_out[117] bl_out[118] br_out[118] bl_out[119] br_out[119] bl_out[120] br_out[120] bl_out[121] br_out[121] bl_out[122] br_out[122] bl_out[123] br_out[123] bl_out[124] br_out[124] bl_out[125] br_out[125] bl_out[126] br_out[126] bl_out[127] br_out[127] gated_w_en vdd gnd write_driver_array
Xdata_in_flop_array DATA[0] DATA[1] DATA[2] DATA[3] DATA[4] DATA[5] DATA[6] DATA[7] DATA[8] DATA[9] DATA[10] DATA[11] DATA[12] DATA[13] DATA[14] DATA[15] DATA[16] DATA[17] DATA[18] DATA[19] DATA[20] DATA[21] DATA[22] DATA[23] DATA[24] DATA[25] DATA[26] DATA[27] DATA[28] DATA[29] DATA[30] DATA[31] DATA[32] DATA[33] DATA[34] DATA[35] DATA[36] DATA[37] DATA[38] DATA[39] DATA[40] DATA[41] DATA[42] DATA[43] DATA[44] DATA[45] DATA[46] DATA[47] DATA[48] DATA[49] DATA[50] DATA[51] DATA[52] DATA[53] DATA[54] DATA[55] DATA[56] DATA[57] DATA[58] DATA[59] DATA[60] DATA[61] DATA[62] DATA[63] DATA[64] DATA[65] DATA[66] DATA[67] DATA[68] DATA[69] DATA[70] DATA[71] DATA[72] DATA[73] DATA[74] DATA[75] DATA[76] DATA[77] DATA[78] DATA[79] DATA[80] DATA[81] DATA[82] DATA[83] DATA[84] DATA[85] DATA[86] DATA[87] DATA[88] DATA[89] DATA[90] DATA[91] DATA[92] DATA[93] DATA[94] DATA[95] DATA[96] DATA[97] DATA[98] DATA[99] DATA[100] DATA[101] DATA[102] DATA[103] DATA[104] DATA[105] DATA[106] DATA[107] DATA[108] DATA[109] DATA[110] DATA[111] DATA[112] DATA[113] DATA[114] DATA[115] DATA[116] DATA[117] DATA[118] DATA[119] DATA[120] DATA[121] DATA[122] DATA[123] DATA[124] DATA[125] DATA[126] DATA[127] data_in[0] data_in_bar[0] data_in[1] data_in_bar[1] data_in[2] data_in_bar[2] data_in[3] data_in_bar[3] data_in[4] data_in_bar[4] data_in[5] data_in_bar[5] data_in[6] data_in_bar[6] data_in[7] data_in_bar[7] data_in[8] data_in_bar[8] data_in[9] data_in_bar[9] data_in[10] data_in_bar[10] data_in[11] data_in_bar[11] data_in[12] data_in_bar[12] data_in[13] data_in_bar[13] data_in[14] data_in_bar[14] data_in[15] data_in_bar[15] data_in[16] data_in_bar[16] data_in[17] data_in_bar[17] data_in[18] data_in_bar[18] data_in[19] data_in_bar[19] data_in[20] data_in_bar[20] data_in[21] data_in_bar[21] data_in[22] data_in_bar[22] data_in[23] data_in_bar[23] data_in[24] data_in_bar[24] data_in[25] data_in_bar[25] data_in[26] data_in_bar[26] data_in[27] data_in_bar[27] data_in[28] data_in_bar[28] data_in[29] data_in_bar[29] data_in[30] data_in_bar[30] data_in[31] data_in_bar[31] data_in[32] data_in_bar[32] data_in[33] data_in_bar[33] data_in[34] data_in_bar[34] data_in[35] data_in_bar[35] data_in[36] data_in_bar[36] data_in[37] data_in_bar[37] data_in[38] data_in_bar[38] data_in[39] data_in_bar[39] data_in[40] data_in_bar[40] data_in[41] data_in_bar[41] data_in[42] data_in_bar[42] data_in[43] data_in_bar[43] data_in[44] data_in_bar[44] data_in[45] data_in_bar[45] data_in[46] data_in_bar[46] data_in[47] data_in_bar[47] data_in[48] data_in_bar[48] data_in[49] data_in_bar[49] data_in[50] data_in_bar[50] data_in[51] data_in_bar[51] data_in[52] data_in_bar[52] data_in[53] data_in_bar[53] data_in[54] data_in_bar[54] data_in[55] data_in_bar[55] data_in[56] data_in_bar[56] data_in[57] data_in_bar[57] data_in[58] data_in_bar[58] data_in[59] data_in_bar[59] data_in[60] data_in_bar[60] data_in[61] data_in_bar[61] data_in[62] data_in_bar[62] data_in[63] data_in_bar[63] data_in[64] data_in_bar[64] data_in[65] data_in_bar[65] data_in[66] data_in_bar[66] data_in[67] data_in_bar[67] data_in[68] data_in_bar[68] data_in[69] data_in_bar[69] data_in[70] data_in_bar[70] data_in[71] data_in_bar[71] data_in[72] data_in_bar[72] data_in[73] data_in_bar[73] data_in[74] data_in_bar[74] data_in[75] data_in_bar[75] data_in[76] data_in_bar[76] data_in[77] data_in_bar[77] data_in[78] data_in_bar[78] data_in[79] data_in_bar[79] data_in[80] data_in_bar[80] data_in[81] data_in_bar[81] data_in[82] data_in_bar[82] data_in[83] data_in_bar[83] data_in[84] data_in_bar[84] data_in[85] data_in_bar[85] data_in[86] data_in_bar[86] data_in[87] data_in_bar[87] data_in[88] data_in_bar[88] data_in[89] data_in_bar[89] data_in[90] data_in_bar[90] data_in[91] data_in_bar[91] data_in[92] data_in_bar[92] data_in[93] data_in_bar[93] data_in[94] data_in_bar[94] data_in[95] data_in_bar[95] data_in[96] data_in_bar[96] data_in[97] data_in_bar[97] data_in[98] data_in_bar[98] data_in[99] data_in_bar[99] data_in[100] data_in_bar[100] data_in[101] data_in_bar[101] data_in[102] data_in_bar[102] data_in[103] data_in_bar[103] data_in[104] data_in_bar[104] data_in[105] data_in_bar[105] data_in[106] data_in_bar[106] data_in[107] data_in_bar[107] data_in[108] data_in_bar[108] data_in[109] data_in_bar[109] data_in[110] data_in_bar[110] data_in[111] data_in_bar[111] data_in[112] data_in_bar[112] data_in[113] data_in_bar[113] data_in[114] data_in_bar[114] data_in[115] data_in_bar[115] data_in[116] data_in_bar[116] data_in[117] data_in_bar[117] data_in[118] data_in_bar[118] data_in[119] data_in_bar[119] data_in[120] data_in_bar[120] data_in[121] data_in_bar[121] data_in[122] data_in_bar[122] data_in[123] data_in_bar[123] data_in[124] data_in_bar[124] data_in[125] data_in_bar[125] data_in[126] data_in_bar[126] data_in[127] data_in_bar[127] gated_clk_bar vdd gnd msf_data_in
Xtri_gate_array data_out[0] data_out[1] data_out[2] data_out[3] data_out[4] data_out[5] data_out[6] data_out[7] data_out[8] data_out[9] data_out[10] data_out[11] data_out[12] data_out[13] data_out[14] data_out[15] data_out[16] data_out[17] data_out[18] data_out[19] data_out[20] data_out[21] data_out[22] data_out[23] data_out[24] data_out[25] data_out[26] data_out[27] data_out[28] data_out[29] data_out[30] data_out[31] data_out[32] data_out[33] data_out[34] data_out[35] data_out[36] data_out[37] data_out[38] data_out[39] data_out[40] data_out[41] data_out[42] data_out[43] data_out[44] data_out[45] data_out[46] data_out[47] data_out[48] data_out[49] data_out[50] data_out[51] data_out[52] data_out[53] data_out[54] data_out[55] data_out[56] data_out[57] data_out[58] data_out[59] data_out[60] data_out[61] data_out[62] data_out[63] data_out[64] data_out[65] data_out[66] data_out[67] data_out[68] data_out[69] data_out[70] data_out[71] data_out[72] data_out[73] data_out[74] data_out[75] data_out[76] data_out[77] data_out[78] data_out[79] data_out[80] data_out[81] data_out[82] data_out[83] data_out[84] data_out[85] data_out[86] data_out[87] data_out[88] data_out[89] data_out[90] data_out[91] data_out[92] data_out[93] data_out[94] data_out[95] data_out[96] data_out[97] data_out[98] data_out[99] data_out[100] data_out[101] data_out[102] data_out[103] data_out[104] data_out[105] data_out[106] data_out[107] data_out[108] data_out[109] data_out[110] data_out[111] data_out[112] data_out[113] data_out[114] data_out[115] data_out[116] data_out[117] data_out[118] data_out[119] data_out[120] data_out[121] data_out[122] data_out[123] data_out[124] data_out[125] data_out[126] data_out[127] DATA[0] DATA[1] DATA[2] DATA[3] DATA[4] DATA[5] DATA[6] DATA[7] DATA[8] DATA[9] DATA[10] DATA[11] DATA[12] DATA[13] DATA[14] DATA[15] DATA[16] DATA[17] DATA[18] DATA[19] DATA[20] DATA[21] DATA[22] DATA[23] DATA[24] DATA[25] DATA[26] DATA[27] DATA[28] DATA[29] DATA[30] DATA[31] DATA[32] DATA[33] DATA[34] DATA[35] DATA[36] DATA[37] DATA[38] DATA[39] DATA[40] DATA[41] DATA[42] DATA[43] DATA[44] DATA[45] DATA[46] DATA[47] DATA[48] DATA[49] DATA[50] DATA[51] DATA[52] DATA[53] DATA[54] DATA[55] DATA[56] DATA[57] DATA[58] DATA[59] DATA[60] DATA[61] DATA[62] DATA[63] DATA[64] DATA[65] DATA[66] DATA[67] DATA[68] DATA[69] DATA[70] DATA[71] DATA[72] DATA[73] DATA[74] DATA[75] DATA[76] DATA[77] DATA[78] DATA[79] DATA[80] DATA[81] DATA[82] DATA[83] DATA[84] DATA[85] DATA[86] DATA[87] DATA[88] DATA[89] DATA[90] DATA[91] DATA[92] DATA[93] DATA[94] DATA[95] DATA[96] DATA[97] DATA[98] DATA[99] DATA[100] DATA[101] DATA[102] DATA[103] DATA[104] DATA[105] DATA[106] DATA[107] DATA[108] DATA[109] DATA[110] DATA[111] DATA[112] DATA[113] DATA[114] DATA[115] DATA[116] DATA[117] DATA[118] DATA[119] DATA[120] DATA[121] DATA[122] DATA[123] DATA[124] DATA[125] DATA[126] DATA[127] gated_tri_en gated_tri_en_bar vdd gnd tri_gate_array
Xrow_decoder A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7] dec_out[0] dec_out[1] dec_out[2] dec_out[3] dec_out[4] dec_out[5] dec_out[6] dec_out[7] dec_out[8] dec_out[9] dec_out[10] dec_out[11] dec_out[12] dec_out[13] dec_out[14] dec_out[15] dec_out[16] dec_out[17] dec_out[18] dec_out[19] dec_out[20] dec_out[21] dec_out[22] dec_out[23] dec_out[24] dec_out[25] dec_out[26] dec_out[27] dec_out[28] dec_out[29] dec_out[30] dec_out[31] dec_out[32] dec_out[33] dec_out[34] dec_out[35] dec_out[36] dec_out[37] dec_out[38] dec_out[39] dec_out[40] dec_out[41] dec_out[42] dec_out[43] dec_out[44] dec_out[45] dec_out[46] dec_out[47] dec_out[48] dec_out[49] dec_out[50] dec_out[51] dec_out[52] dec_out[53] dec_out[54] dec_out[55] dec_out[56] dec_out[57] dec_out[58] dec_out[59] dec_out[60] dec_out[61] dec_out[62] dec_out[63] dec_out[64] dec_out[65] dec_out[66] dec_out[67] dec_out[68] dec_out[69] dec_out[70] dec_out[71] dec_out[72] dec_out[73] dec_out[74] dec_out[75] dec_out[76] dec_out[77] dec_out[78] dec_out[79] dec_out[80] dec_out[81] dec_out[82] dec_out[83] dec_out[84] dec_out[85] dec_out[86] dec_out[87] dec_out[88] dec_out[89] dec_out[90] dec_out[91] dec_out[92] dec_out[93] dec_out[94] dec_out[95] dec_out[96] dec_out[97] dec_out[98] dec_out[99] dec_out[100] dec_out[101] dec_out[102] dec_out[103] dec_out[104] dec_out[105] dec_out[106] dec_out[107] dec_out[108] dec_out[109] dec_out[110] dec_out[111] dec_out[112] dec_out[113] dec_out[114] dec_out[115] dec_out[116] dec_out[117] dec_out[118] dec_out[119] dec_out[120] dec_out[121] dec_out[122] dec_out[123] dec_out[124] dec_out[125] dec_out[126] dec_out[127] dec_out[128] dec_out[129] dec_out[130] dec_out[131] dec_out[132] dec_out[133] dec_out[134] dec_out[135] dec_out[136] dec_out[137] dec_out[138] dec_out[139] dec_out[140] dec_out[141] dec_out[142] dec_out[143] dec_out[144] dec_out[145] dec_out[146] dec_out[147] dec_out[148] dec_out[149] dec_out[150] dec_out[151] dec_out[152] dec_out[153] dec_out[154] dec_out[155] dec_out[156] dec_out[157] dec_out[158] dec_out[159] dec_out[160] dec_out[161] dec_out[162] dec_out[163] dec_out[164] dec_out[165] dec_out[166] dec_out[167] dec_out[168] dec_out[169] dec_out[170] dec_out[171] dec_out[172] dec_out[173] dec_out[174] dec_out[175] dec_out[176] dec_out[177] dec_out[178] dec_out[179] dec_out[180] dec_out[181] dec_out[182] dec_out[183] dec_out[184] dec_out[185] dec_out[186] dec_out[187] dec_out[188] dec_out[189] dec_out[190] dec_out[191] dec_out[192] dec_out[193] dec_out[194] dec_out[195] dec_out[196] dec_out[197] dec_out[198] dec_out[199] dec_out[200] dec_out[201] dec_out[202] dec_out[203] dec_out[204] dec_out[205] dec_out[206] dec_out[207] dec_out[208] dec_out[209] dec_out[210] dec_out[211] dec_out[212] dec_out[213] dec_out[214] dec_out[215] dec_out[216] dec_out[217] dec_out[218] dec_out[219] dec_out[220] dec_out[221] dec_out[222] dec_out[223] dec_out[224] dec_out[225] dec_out[226] dec_out[227] dec_out[228] dec_out[229] dec_out[230] dec_out[231] dec_out[232] dec_out[233] dec_out[234] dec_out[235] dec_out[236] dec_out[237] dec_out[238] dec_out[239] dec_out[240] dec_out[241] dec_out[242] dec_out[243] dec_out[244] dec_out[245] dec_out[246] dec_out[247] dec_out[248] dec_out[249] dec_out[250] dec_out[251] dec_out[252] dec_out[253] dec_out[254] dec_out[255] vdd gnd hierarchical_decoder_256rows
Xwordline_driver dec_out[0] dec_out[1] dec_out[2] dec_out[3] dec_out[4] dec_out[5] dec_out[6] dec_out[7] dec_out[8] dec_out[9] dec_out[10] dec_out[11] dec_out[12] dec_out[13] dec_out[14] dec_out[15] dec_out[16] dec_out[17] dec_out[18] dec_out[19] dec_out[20] dec_out[21] dec_out[22] dec_out[23] dec_out[24] dec_out[25] dec_out[26] dec_out[27] dec_out[28] dec_out[29] dec_out[30] dec_out[31] dec_out[32] dec_out[33] dec_out[34] dec_out[35] dec_out[36] dec_out[37] dec_out[38] dec_out[39] dec_out[40] dec_out[41] dec_out[42] dec_out[43] dec_out[44] dec_out[45] dec_out[46] dec_out[47] dec_out[48] dec_out[49] dec_out[50] dec_out[51] dec_out[52] dec_out[53] dec_out[54] dec_out[55] dec_out[56] dec_out[57] dec_out[58] dec_out[59] dec_out[60] dec_out[61] dec_out[62] dec_out[63] dec_out[64] dec_out[65] dec_out[66] dec_out[67] dec_out[68] dec_out[69] dec_out[70] dec_out[71] dec_out[72] dec_out[73] dec_out[74] dec_out[75] dec_out[76] dec_out[77] dec_out[78] dec_out[79] dec_out[80] dec_out[81] dec_out[82] dec_out[83] dec_out[84] dec_out[85] dec_out[86] dec_out[87] dec_out[88] dec_out[89] dec_out[90] dec_out[91] dec_out[92] dec_out[93] dec_out[94] dec_out[95] dec_out[96] dec_out[97] dec_out[98] dec_out[99] dec_out[100] dec_out[101] dec_out[102] dec_out[103] dec_out[104] dec_out[105] dec_out[106] dec_out[107] dec_out[108] dec_out[109] dec_out[110] dec_out[111] dec_out[112] dec_out[113] dec_out[114] dec_out[115] dec_out[116] dec_out[117] dec_out[118] dec_out[119] dec_out[120] dec_out[121] dec_out[122] dec_out[123] dec_out[124] dec_out[125] dec_out[126] dec_out[127] dec_out[128] dec_out[129] dec_out[130] dec_out[131] dec_out[132] dec_out[133] dec_out[134] dec_out[135] dec_out[136] dec_out[137] dec_out[138] dec_out[139] dec_out[140] dec_out[141] dec_out[142] dec_out[143] dec_out[144] dec_out[145] dec_out[146] dec_out[147] dec_out[148] dec_out[149] dec_out[150] dec_out[151] dec_out[152] dec_out[153] dec_out[154] dec_out[155] dec_out[156] dec_out[157] dec_out[158] dec_out[159] dec_out[160] dec_out[161] dec_out[162] dec_out[163] dec_out[164] dec_out[165] dec_out[166] dec_out[167] dec_out[168] dec_out[169] dec_out[170] dec_out[171] dec_out[172] dec_out[173] dec_out[174] dec_out[175] dec_out[176] dec_out[177] dec_out[178] dec_out[179] dec_out[180] dec_out[181] dec_out[182] dec_out[183] dec_out[184] dec_out[185] dec_out[186] dec_out[187] dec_out[188] dec_out[189] dec_out[190] dec_out[191] dec_out[192] dec_out[193] dec_out[194] dec_out[195] dec_out[196] dec_out[197] dec_out[198] dec_out[199] dec_out[200] dec_out[201] dec_out[202] dec_out[203] dec_out[204] dec_out[205] dec_out[206] dec_out[207] dec_out[208] dec_out[209] dec_out[210] dec_out[211] dec_out[212] dec_out[213] dec_out[214] dec_out[215] dec_out[216] dec_out[217] dec_out[218] dec_out[219] dec_out[220] dec_out[221] dec_out[222] dec_out[223] dec_out[224] dec_out[225] dec_out[226] dec_out[227] dec_out[228] dec_out[229] dec_out[230] dec_out[231] dec_out[232] dec_out[233] dec_out[234] dec_out[235] dec_out[236] dec_out[237] dec_out[238] dec_out[239] dec_out[240] dec_out[241] dec_out[242] dec_out[243] dec_out[244] dec_out[245] dec_out[246] dec_out[247] dec_out[248] dec_out[249] dec_out[250] dec_out[251] dec_out[252] dec_out[253] dec_out[254] dec_out[255] wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] wl[128] wl[129] wl[130] wl[131] wl[132] wl[133] wl[134] wl[135] wl[136] wl[137] wl[138] wl[139] wl[140] wl[141] wl[142] wl[143] wl[144] wl[145] wl[146] wl[147] wl[148] wl[149] wl[150] wl[151] wl[152] wl[153] wl[154] wl[155] wl[156] wl[157] wl[158] wl[159] wl[160] wl[161] wl[162] wl[163] wl[164] wl[165] wl[166] wl[167] wl[168] wl[169] wl[170] wl[171] wl[172] wl[173] wl[174] wl[175] wl[176] wl[177] wl[178] wl[179] wl[180] wl[181] wl[182] wl[183] wl[184] wl[185] wl[186] wl[187] wl[188] wl[189] wl[190] wl[191] wl[192] wl[193] wl[194] wl[195] wl[196] wl[197] wl[198] wl[199] wl[200] wl[201] wl[202] wl[203] wl[204] wl[205] wl[206] wl[207] wl[208] wl[209] wl[210] wl[211] wl[212] wl[213] wl[214] wl[215] wl[216] wl[217] wl[218] wl[219] wl[220] wl[221] wl[222] wl[223] wl[224] wl[225] wl[226] wl[227] wl[228] wl[229] wl[230] wl[231] wl[232] wl[233] wl[234] wl[235] wl[236] wl[237] wl[238] wl[239] wl[240] wl[241] wl[242] wl[243] wl[244] wl[245] wl[246] wl[247] wl[248] wl[249] wl[250] wl[251] wl[252] wl[253] wl[254] wl[255] gated_clk_buf vdd gnd wordline_driver
Xaddress_flop_array ADDR[0] ADDR[1] ADDR[2] ADDR[3] ADDR[4] ADDR[5] ADDR[6] ADDR[7] ADDR[8] A[0] A_bar[0] A[1] A_bar[1] A[2] A_bar[2] A[3] A_bar[3] A[4] A_bar[4] A[5] A_bar[5] A[6] A_bar[6] A[7] A_bar[7] sel[1] sel[0] gated_clk_buf vdd gnd msf_address
Xbank_sel_inv bank_sel bank_sel_bar vdd gnd pinv_13
Xnor_clk_buf clk_buf bank_sel_bar gated_clk_buf_temp_bar vdd gnd pnor2_2
Xinv_clk_buf gated_clk_buf_temp_bar gated_clk_buf vdd gnd pinv_14
Xnor_tri_en_bar tri_en_bar bank_sel_bar gated_tri_en_bar_temp_bar vdd gnd pnor2_2
Xinv_tri_en_bar gated_tri_en_bar_temp_bar gated_tri_en_bar vdd gnd pinv_14
Xnand_tri_en tri_en bank_sel gated_tri_en_temp_bar vdd gnd pnand2_5
Xinv_tri_en gated_tri_en_temp_bar gated_tri_en vdd gnd pinv_14
Xnand_clk_bar clk_bar bank_sel gated_clk_bar_temp_bar vdd gnd pnand2_5
Xinv_clk_bar gated_clk_bar_temp_bar gated_clk_bar vdd gnd pinv_14
Xnand_w_en w_en bank_sel gated_w_en_temp_bar vdd gnd pnand2_5
Xinv_w_en gated_w_en_temp_bar gated_w_en vdd gnd pinv_14
Xnand_s_en s_en bank_sel gated_s_en_temp_bar vdd gnd pnand2_5
Xinv_s_en gated_s_en_temp_bar gated_s_en vdd gnd pinv_14
.ENDS bank

.SUBCKT msb_address din[0] dout[0] dout_bar[0] clk vdd gnd
XXdff0 din[0] dout[0] dout_bar[0] clk vdd gnd ms_flop
.ENDS msb_address

.SUBCKT sram_1rw_128b_1024w_2bank_scn3me_subm DATA[0] DATA[1] DATA[2] DATA[3] DATA[4] DATA[5] DATA[6] DATA[7] DATA[8] DATA[9] DATA[10] DATA[11] DATA[12] DATA[13] DATA[14] DATA[15] DATA[16] DATA[17] DATA[18] DATA[19] DATA[20] DATA[21] DATA[22] DATA[23] DATA[24] DATA[25] DATA[26] DATA[27] DATA[28] DATA[29] DATA[30] DATA[31] DATA[32] DATA[33] DATA[34] DATA[35] DATA[36] DATA[37] DATA[38] DATA[39] DATA[40] DATA[41] DATA[42] DATA[43] DATA[44] DATA[45] DATA[46] DATA[47] DATA[48] DATA[49] DATA[50] DATA[51] DATA[52] DATA[53] DATA[54] DATA[55] DATA[56] DATA[57] DATA[58] DATA[59] DATA[60] DATA[61] DATA[62] DATA[63] DATA[64] DATA[65] DATA[66] DATA[67] DATA[68] DATA[69] DATA[70] DATA[71] DATA[72] DATA[73] DATA[74] DATA[75] DATA[76] DATA[77] DATA[78] DATA[79] DATA[80] DATA[81] DATA[82] DATA[83] DATA[84] DATA[85] DATA[86] DATA[87] DATA[88] DATA[89] DATA[90] DATA[91] DATA[92] DATA[93] DATA[94] DATA[95] DATA[96] DATA[97] DATA[98] DATA[99] DATA[100] DATA[101] DATA[102] DATA[103] DATA[104] DATA[105] DATA[106] DATA[107] DATA[108] DATA[109] DATA[110] DATA[111] DATA[112] DATA[113] DATA[114] DATA[115] DATA[116] DATA[117] DATA[118] DATA[119] DATA[120] DATA[121] DATA[122] DATA[123] DATA[124] DATA[125] DATA[126] DATA[127] ADDR[0] ADDR[1] ADDR[2] ADDR[3] ADDR[4] ADDR[5] ADDR[6] ADDR[7] ADDR[8] ADDR[9] CSb WEb OEb clk vdd gnd
Xbank0 DATA[0] DATA[1] DATA[2] DATA[3] DATA[4] DATA[5] DATA[6] DATA[7] DATA[8] DATA[9] DATA[10] DATA[11] DATA[12] DATA[13] DATA[14] DATA[15] DATA[16] DATA[17] DATA[18] DATA[19] DATA[20] DATA[21] DATA[22] DATA[23] DATA[24] DATA[25] DATA[26] DATA[27] DATA[28] DATA[29] DATA[30] DATA[31] DATA[32] DATA[33] DATA[34] DATA[35] DATA[36] DATA[37] DATA[38] DATA[39] DATA[40] DATA[41] DATA[42] DATA[43] DATA[44] DATA[45] DATA[46] DATA[47] DATA[48] DATA[49] DATA[50] DATA[51] DATA[52] DATA[53] DATA[54] DATA[55] DATA[56] DATA[57] DATA[58] DATA[59] DATA[60] DATA[61] DATA[62] DATA[63] DATA[64] DATA[65] DATA[66] DATA[67] DATA[68] DATA[69] DATA[70] DATA[71] DATA[72] DATA[73] DATA[74] DATA[75] DATA[76] DATA[77] DATA[78] DATA[79] DATA[80] DATA[81] DATA[82] DATA[83] DATA[84] DATA[85] DATA[86] DATA[87] DATA[88] DATA[89] DATA[90] DATA[91] DATA[92] DATA[93] DATA[94] DATA[95] DATA[96] DATA[97] DATA[98] DATA[99] DATA[100] DATA[101] DATA[102] DATA[103] DATA[104] DATA[105] DATA[106] DATA[107] DATA[108] DATA[109] DATA[110] DATA[111] DATA[112] DATA[113] DATA[114] DATA[115] DATA[116] DATA[117] DATA[118] DATA[119] DATA[120] DATA[121] DATA[122] DATA[123] DATA[124] DATA[125] DATA[126] DATA[127] ADDR[0] ADDR[1] ADDR[2] ADDR[3] ADDR[4] ADDR[5] ADDR[6] ADDR[7] ADDR[8] bank_sel[0] s_en w_en tri_en_bar tri_en clk_bar clk_buf vdd gnd bank
Xbank1 DATA[0] DATA[1] DATA[2] DATA[3] DATA[4] DATA[5] DATA[6] DATA[7] DATA[8] DATA[9] DATA[10] DATA[11] DATA[12] DATA[13] DATA[14] DATA[15] DATA[16] DATA[17] DATA[18] DATA[19] DATA[20] DATA[21] DATA[22] DATA[23] DATA[24] DATA[25] DATA[26] DATA[27] DATA[28] DATA[29] DATA[30] DATA[31] DATA[32] DATA[33] DATA[34] DATA[35] DATA[36] DATA[37] DATA[38] DATA[39] DATA[40] DATA[41] DATA[42] DATA[43] DATA[44] DATA[45] DATA[46] DATA[47] DATA[48] DATA[49] DATA[50] DATA[51] DATA[52] DATA[53] DATA[54] DATA[55] DATA[56] DATA[57] DATA[58] DATA[59] DATA[60] DATA[61] DATA[62] DATA[63] DATA[64] DATA[65] DATA[66] DATA[67] DATA[68] DATA[69] DATA[70] DATA[71] DATA[72] DATA[73] DATA[74] DATA[75] DATA[76] DATA[77] DATA[78] DATA[79] DATA[80] DATA[81] DATA[82] DATA[83] DATA[84] DATA[85] DATA[86] DATA[87] DATA[88] DATA[89] DATA[90] DATA[91] DATA[92] DATA[93] DATA[94] DATA[95] DATA[96] DATA[97] DATA[98] DATA[99] DATA[100] DATA[101] DATA[102] DATA[103] DATA[104] DATA[105] DATA[106] DATA[107] DATA[108] DATA[109] DATA[110] DATA[111] DATA[112] DATA[113] DATA[114] DATA[115] DATA[116] DATA[117] DATA[118] DATA[119] DATA[120] DATA[121] DATA[122] DATA[123] DATA[124] DATA[125] DATA[126] DATA[127] ADDR[0] ADDR[1] ADDR[2] ADDR[3] ADDR[4] ADDR[5] ADDR[6] ADDR[7] ADDR[8] bank_sel[1] s_en w_en tri_en_bar tri_en clk_bar clk_buf vdd gnd bank
Xcontrol CSb WEb OEb clk s_en w_en tri_en tri_en_bar clk_bar clk_buf vdd gnd control_logic
Xmsb_address ADDR[9] bank_sel[1] bank_sel[0] clk_buf vdd gnd msb_address
.ENDS sram_1rw_128b_1024w_2bank_scn3me_subm
