magic
tech sky130A
magscale 1 2
timestamp 1595931502
<< checkpaint >>
rect -1296 -1277 2690 2731
<< locali >>
rect 0 1397 1394 1431
rect 330 708 364 1151
rect 330 674 459 708
rect 883 674 917 708
rect 212 485 246 551
rect 112 237 146 303
rect 0 -17 1394 17
use pnand2  pnand2_0
timestamp 1595931502
transform 1 0 0 0 1 0
box -36 -17 414 1471
use pdriver  pdriver_0
timestamp 1595931502
transform 1 0 378 0 1 0
box -36 -17 1052 1471
<< labels >>
rlabel corelocali s 697 0 697 0 4 gnd
rlabel corelocali s 229 518 229 518 4 B
rlabel corelocali s 900 691 900 691 4 Z
rlabel corelocali s 697 1414 697 1414 4 vdd
rlabel corelocali s 129 270 129 270 4 A
<< properties >>
string FIXED_BBOX 0 0 1394 1414
<< end >>
