magic
tech sky130A
magscale 1 2
timestamp 1595931502
<< checkpaint >>
rect -1296 -1277 1922 2731
<< nwell >>
rect -36 679 662 1471
<< locali >>
rect 0 1397 626 1431
rect 64 636 98 702
rect 196 652 449 686
rect 547 652 581 686
rect 0 -17 626 17
use pinv_7  pinv_7_0
timestamp 1595931502
transform 1 0 368 0 1 0
box -36 -17 294 1471
use pinv_4  pinv_4_0
timestamp 1595931502
transform 1 0 0 0 1 0
box -36 -17 404 1471
<< labels >>
rlabel corelocali s 313 0 313 0 4 gnd
rlabel corelocali s 564 669 564 669 4 Z
rlabel corelocali s 313 1414 313 1414 4 vdd
rlabel corelocali s 81 669 81 669 4 A
<< properties >>
string FIXED_BBOX 0 0 626 1414
<< end >>
