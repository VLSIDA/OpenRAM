magic
tech sky130A
magscale 1 2
timestamp 1595931502
<< checkpaint >>
rect -1190 -1316 2148 1736
<< nwell >>
rect 412 -56 888 476
<< nmos >>
rect 196 266 344 296
rect 196 194 344 224
<< pmos >>
rect 582 272 806 302
rect 582 182 806 212
<< ndiff >>
rect 196 348 344 356
rect 196 314 257 348
rect 291 314 344 348
rect 196 296 344 314
rect 196 224 344 266
rect 196 176 344 194
rect 196 142 259 176
rect 293 142 344 176
rect 196 108 344 142
<< pdiff >>
rect 582 348 806 356
rect 582 314 677 348
rect 711 314 806 348
rect 582 302 806 314
rect 582 260 806 272
rect 582 226 677 260
rect 711 226 806 260
rect 582 212 806 226
rect 582 170 806 182
rect 582 136 677 170
rect 711 136 806 170
rect 582 128 806 136
<< ndiffc >>
rect 257 314 291 348
rect 259 142 293 176
<< pdiffc >>
rect 677 314 711 348
rect 677 226 711 260
rect 677 136 711 170
<< psubdiff >>
rect 228 17 312 18
rect 228 -17 253 17
rect 287 -17 312 17
rect 228 -18 312 -17
<< nsubdiff >>
rect 654 17 738 19
rect 654 -17 679 17
rect 713 -17 738 17
rect 654 -19 738 -17
<< psubdiffcont >>
rect 253 -17 287 17
<< nsubdiffcont >>
rect 679 -17 713 17
<< poly >>
rect 76 316 130 332
rect 76 282 86 316
rect 120 296 130 316
rect 460 296 582 302
rect 120 282 196 296
rect 76 266 196 282
rect 344 272 582 296
rect 806 272 832 302
rect 344 266 478 272
rect 76 208 196 224
rect 76 174 86 208
rect 120 194 196 208
rect 344 212 490 224
rect 344 194 582 212
rect 120 174 130 194
rect 76 158 130 174
rect 458 182 582 194
rect 806 182 832 212
<< polycont >>
rect 86 282 120 316
rect 86 174 120 208
<< locali >>
rect 70 282 86 316
rect 120 282 136 316
rect 210 314 257 348
rect 291 314 677 348
rect 711 314 888 348
rect 70 174 86 208
rect 120 174 136 208
rect 208 142 254 176
rect 293 142 340 176
rect 509 170 543 314
rect 660 226 677 260
rect 711 226 727 260
rect 509 169 598 170
rect 660 169 677 170
rect 509 136 677 169
rect 711 136 728 170
rect 509 135 685 136
rect 509 134 572 135
rect 236 17 312 18
rect 236 -17 253 17
rect 287 -17 312 17
rect 236 -18 312 -17
rect 660 17 730 19
rect 660 -17 679 17
rect 713 -17 730 17
rect 660 -19 730 -17
<< viali >>
rect 254 142 259 176
rect 259 142 288 176
rect 677 226 711 260
rect 253 -17 287 17
rect 679 -17 713 17
<< metal1 >>
rect 246 176 294 402
rect 246 142 254 176
rect 288 142 294 176
rect 246 17 294 142
rect 246 -17 253 17
rect 287 -17 294 17
rect 246 -30 294 -17
rect 670 260 720 402
rect 670 226 677 260
rect 711 226 720 260
rect 670 17 720 226
rect 670 -17 679 17
rect 713 -17 720 17
rect 670 -32 720 -17
<< labels >>
rlabel corelocali s 103 191 103 191 4 B
rlabel corelocali s 103 299 103 299 4 A
rlabel corelocali s 854 331 854 331 4 Z
rlabel metal1 s 696 94 696 94 4 vdd
rlabel metal1 s 268 82 268 82 4 gnd
rlabel metal1 s 270 186 270 186 4 gnd
rlabel corelocali s 103 191 103 191 4 B
rlabel corelocali s 549 331 549 331 4 Z
rlabel metal1 s 695 185 695 185 4 vdd
rlabel corelocali s 103 299 103 299 4 A
<< properties >>
string FIXED_BBOX 0 0 876 395
<< end >>
