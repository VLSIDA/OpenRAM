magic
tech sky130A
magscale 1 2
timestamp 1595931502
<< checkpaint >>
rect -1302 -841 1884 8741
<< metal2 >>
rect 0 7433 624 7481
rect 0 7213 624 7261
rect 0 6959 624 7007
rect 0 6739 624 6787
rect 0 6643 624 6691
rect 0 6423 624 6471
rect 0 6169 624 6217
rect 0 5949 624 5997
rect 0 5853 624 5901
rect 0 5633 624 5681
rect 0 5379 624 5427
rect 0 5159 624 5207
rect 0 5063 624 5111
rect 0 4843 624 4891
rect 0 4589 624 4637
rect 0 4369 624 4417
rect 0 4273 624 4321
rect 0 4053 624 4101
rect 0 3799 624 3847
rect 0 3579 624 3627
rect 0 3483 624 3531
rect 0 3263 624 3311
rect 0 3009 624 3057
rect 0 2789 624 2837
rect 0 2693 624 2741
rect 0 2473 624 2521
rect 0 2219 624 2267
rect 0 1999 624 2047
rect 0 1903 624 1951
rect 0 1683 624 1731
rect 0 1429 624 1477
rect 0 1209 624 1257
rect 0 1113 624 1161
rect 0 893 624 941
rect 0 639 624 687
rect 0 419 624 467
<< metal3 >>
rect 191 7298 289 7396
rect 191 7061 289 7159
rect 191 6824 289 6922
rect 191 6508 289 6606
rect 191 6271 289 6369
rect 191 6034 289 6132
rect 191 5718 289 5816
rect 191 5481 289 5579
rect 191 5244 289 5342
rect 191 4928 289 5026
rect 191 4691 289 4789
rect 191 4454 289 4552
rect 191 4138 289 4236
rect 191 3901 289 3999
rect 191 3664 289 3762
rect 191 3348 289 3446
rect 191 3111 289 3209
rect 191 2874 289 2972
rect 191 2558 289 2656
rect 191 2321 289 2419
rect 191 2084 289 2182
rect 191 1768 289 1866
rect 191 1531 289 1629
rect 191 1294 289 1392
rect 191 978 289 1076
rect 191 741 289 839
rect 191 504 289 602
use contact_9  contact_9_35
timestamp 1595931502
transform 1 0 207 0 1 516
box 0 0 66 74
use contact_9  contact_9_34
timestamp 1595931502
transform 1 0 207 0 1 753
box 0 0 66 74
use contact_9  contact_9_33
timestamp 1595931502
transform 1 0 207 0 1 990
box 0 0 66 74
use contact_9  contact_9_32
timestamp 1595931502
transform 1 0 207 0 1 753
box 0 0 66 74
use contact_9  contact_9_31
timestamp 1595931502
transform 1 0 207 0 1 1306
box 0 0 66 74
use contact_9  contact_9_30
timestamp 1595931502
transform 1 0 207 0 1 1543
box 0 0 66 74
use contact_9  contact_9_29
timestamp 1595931502
transform 1 0 207 0 1 1780
box 0 0 66 74
use contact_9  contact_9_28
timestamp 1595931502
transform 1 0 207 0 1 1543
box 0 0 66 74
use contact_9  contact_9_27
timestamp 1595931502
transform 1 0 207 0 1 2096
box 0 0 66 74
use contact_9  contact_9_26
timestamp 1595931502
transform 1 0 207 0 1 2333
box 0 0 66 74
use contact_9  contact_9_25
timestamp 1595931502
transform 1 0 207 0 1 2570
box 0 0 66 74
use contact_9  contact_9_24
timestamp 1595931502
transform 1 0 207 0 1 2333
box 0 0 66 74
use contact_9  contact_9_23
timestamp 1595931502
transform 1 0 207 0 1 2886
box 0 0 66 74
use contact_9  contact_9_22
timestamp 1595931502
transform 1 0 207 0 1 3123
box 0 0 66 74
use contact_9  contact_9_21
timestamp 1595931502
transform 1 0 207 0 1 3360
box 0 0 66 74
use contact_9  contact_9_20
timestamp 1595931502
transform 1 0 207 0 1 3123
box 0 0 66 74
use contact_9  contact_9_19
timestamp 1595931502
transform 1 0 207 0 1 3676
box 0 0 66 74
use contact_9  contact_9_18
timestamp 1595931502
transform 1 0 207 0 1 3913
box 0 0 66 74
use contact_9  contact_9_17
timestamp 1595931502
transform 1 0 207 0 1 4150
box 0 0 66 74
use contact_9  contact_9_16
timestamp 1595931502
transform 1 0 207 0 1 3913
box 0 0 66 74
use contact_9  contact_9_15
timestamp 1595931502
transform 1 0 207 0 1 4466
box 0 0 66 74
use contact_9  contact_9_14
timestamp 1595931502
transform 1 0 207 0 1 4703
box 0 0 66 74
use contact_9  contact_9_13
timestamp 1595931502
transform 1 0 207 0 1 4940
box 0 0 66 74
use contact_9  contact_9_12
timestamp 1595931502
transform 1 0 207 0 1 4703
box 0 0 66 74
use contact_9  contact_9_11
timestamp 1595931502
transform 1 0 207 0 1 5256
box 0 0 66 74
use contact_9  contact_9_10
timestamp 1595931502
transform 1 0 207 0 1 5493
box 0 0 66 74
use contact_9  contact_9_9
timestamp 1595931502
transform 1 0 207 0 1 5730
box 0 0 66 74
use contact_9  contact_9_8
timestamp 1595931502
transform 1 0 207 0 1 5493
box 0 0 66 74
use contact_9  contact_9_7
timestamp 1595931502
transform 1 0 207 0 1 6046
box 0 0 66 74
use contact_9  contact_9_6
timestamp 1595931502
transform 1 0 207 0 1 6283
box 0 0 66 74
use contact_9  contact_9_5
timestamp 1595931502
transform 1 0 207 0 1 6520
box 0 0 66 74
use contact_9  contact_9_4
timestamp 1595931502
transform 1 0 207 0 1 6283
box 0 0 66 74
use contact_9  contact_9_3
timestamp 1595931502
transform 1 0 207 0 1 6836
box 0 0 66 74
use contact_9  contact_9_2
timestamp 1595931502
transform 1 0 207 0 1 7073
box 0 0 66 74
use contact_9  contact_9_1
timestamp 1595931502
transform 1 0 207 0 1 7310
box 0 0 66 74
use contact_9  contact_9_0
timestamp 1595931502
transform 1 0 207 0 1 7073
box 0 0 66 74
use row_cap_cell_1rw_1r  row_cap_cell_1rw_1r_17
timestamp 1595931502
transform 1 0 0 0 -1 790
box -42 -55 624 371
use row_cap_cell_1rw_1r  row_cap_cell_1rw_1r_16
timestamp 1595931502
transform 1 0 0 0 1 790
box -42 -55 624 371
use row_cap_cell_1rw_1r  row_cap_cell_1rw_1r_15
timestamp 1595931502
transform 1 0 0 0 -1 1580
box -42 -55 624 371
use row_cap_cell_1rw_1r  row_cap_cell_1rw_1r_14
timestamp 1595931502
transform 1 0 0 0 1 1580
box -42 -55 624 371
use row_cap_cell_1rw_1r  row_cap_cell_1rw_1r_13
timestamp 1595931502
transform 1 0 0 0 -1 2370
box -42 -55 624 371
use row_cap_cell_1rw_1r  row_cap_cell_1rw_1r_12
timestamp 1595931502
transform 1 0 0 0 1 2370
box -42 -55 624 371
use row_cap_cell_1rw_1r  row_cap_cell_1rw_1r_11
timestamp 1595931502
transform 1 0 0 0 -1 3160
box -42 -55 624 371
use row_cap_cell_1rw_1r  row_cap_cell_1rw_1r_10
timestamp 1595931502
transform 1 0 0 0 1 3160
box -42 -55 624 371
use row_cap_cell_1rw_1r  row_cap_cell_1rw_1r_9
timestamp 1595931502
transform 1 0 0 0 -1 3950
box -42 -55 624 371
use row_cap_cell_1rw_1r  row_cap_cell_1rw_1r_8
timestamp 1595931502
transform 1 0 0 0 1 3950
box -42 -55 624 371
use row_cap_cell_1rw_1r  row_cap_cell_1rw_1r_7
timestamp 1595931502
transform 1 0 0 0 -1 4740
box -42 -55 624 371
use row_cap_cell_1rw_1r  row_cap_cell_1rw_1r_6
timestamp 1595931502
transform 1 0 0 0 1 4740
box -42 -55 624 371
use row_cap_cell_1rw_1r  row_cap_cell_1rw_1r_5
timestamp 1595931502
transform 1 0 0 0 -1 5530
box -42 -55 624 371
use row_cap_cell_1rw_1r  row_cap_cell_1rw_1r_4
timestamp 1595931502
transform 1 0 0 0 1 5530
box -42 -55 624 371
use row_cap_cell_1rw_1r  row_cap_cell_1rw_1r_3
timestamp 1595931502
transform 1 0 0 0 -1 6320
box -42 -55 624 371
use row_cap_cell_1rw_1r  row_cap_cell_1rw_1r_2
timestamp 1595931502
transform 1 0 0 0 1 6320
box -42 -55 624 371
use row_cap_cell_1rw_1r  row_cap_cell_1rw_1r_1
timestamp 1595931502
transform 1 0 0 0 -1 7110
box -42 -55 624 371
use row_cap_cell_1rw_1r  row_cap_cell_1rw_1r_0
timestamp 1595931502
transform 1 0 0 0 1 7110
box -42 -55 624 371
<< labels >>
rlabel metal2 s 312 4613 312 4613 4 wl1_11
rlabel metal2 s 312 6193 312 6193 4 wl1_15
rlabel metal2 s 312 1927 312 1927 4 wl0_4
rlabel metal2 s 312 917 312 917 4 wl1_2
rlabel metal2 s 312 5403 312 5403 4 wl1_13
rlabel metal2 s 312 6667 312 6667 4 wl0_16
rlabel metal2 s 312 3823 312 3823 4 wl1_9
rlabel metal2 s 312 663 312 663 4 wl1_1
rlabel metal2 s 312 1453 312 1453 4 wl1_3
rlabel metal2 s 312 3033 312 3033 4 wl1_7
rlabel metal2 s 312 7237 312 7237 4 wl1_18
rlabel metal2 s 312 5657 312 5657 4 wl1_14
rlabel metal2 s 312 4393 312 4393 4 wl0_11
rlabel metal2 s 312 7457 312 7457 4 wl0_18
rlabel metal2 s 312 6447 312 6447 4 wl1_16
rlabel metal2 s 312 4077 312 4077 4 wl1_10
rlabel metal2 s 312 1707 312 1707 4 wl1_4
rlabel metal2 s 312 1233 312 1233 4 wl0_3
rlabel metal3 s 240 3713 240 3713 4 gnd
rlabel metal3 s 240 5530 240 5530 4 gnd
rlabel metal3 s 240 6557 240 6557 4 gnd
rlabel metal3 s 240 790 240 790 4 gnd
rlabel metal3 s 240 3397 240 3397 4 gnd
rlabel metal3 s 240 4977 240 4977 4 gnd
rlabel metal3 s 240 2133 240 2133 4 gnd
rlabel metal3 s 240 5767 240 5767 4 gnd
rlabel metal3 s 240 1817 240 1817 4 gnd
rlabel metal3 s 240 1580 240 1580 4 gnd
rlabel metal3 s 240 7110 240 7110 4 gnd
rlabel metal3 s 240 4187 240 4187 4 gnd
rlabel metal3 s 240 1027 240 1027 4 gnd
rlabel metal3 s 240 4503 240 4503 4 gnd
rlabel metal3 s 240 3160 240 3160 4 gnd
rlabel metal3 s 240 3950 240 3950 4 gnd
rlabel metal3 s 240 5293 240 5293 4 gnd
rlabel metal3 s 240 2370 240 2370 4 gnd
rlabel metal3 s 240 6320 240 6320 4 gnd
rlabel metal3 s 240 2607 240 2607 4 gnd
rlabel metal3 s 240 4740 240 4740 4 gnd
rlabel metal3 s 240 553 240 553 4 gnd
rlabel metal3 s 240 6873 240 6873 4 gnd
rlabel metal3 s 240 1343 240 1343 4 gnd
rlabel metal3 s 240 7347 240 7347 4 gnd
rlabel metal3 s 240 2923 240 2923 4 gnd
rlabel metal3 s 240 6083 240 6083 4 gnd
rlabel metal2 s 312 2497 312 2497 4 wl1_6
rlabel metal2 s 312 2717 312 2717 4 wl0_6
rlabel metal2 s 312 6763 312 6763 4 wl0_17
rlabel metal2 s 312 3603 312 3603 4 wl0_9
rlabel metal2 s 312 2813 312 2813 4 wl0_7
rlabel metal2 s 312 5973 312 5973 4 wl0_15
rlabel metal2 s 312 3287 312 3287 4 wl1_8
rlabel metal2 s 312 5087 312 5087 4 wl0_12
rlabel metal2 s 312 4867 312 4867 4 wl1_12
rlabel metal2 s 312 5877 312 5877 4 wl0_14
rlabel metal2 s 312 2243 312 2243 4 wl1_5
rlabel metal2 s 312 6983 312 6983 4 wl1_17
rlabel metal2 s 312 2023 312 2023 4 wl0_5
rlabel metal2 s 312 5183 312 5183 4 wl0_13
rlabel metal2 s 312 443 312 443 4 wl0_1
rlabel metal2 s 312 1137 312 1137 4 wl0_2
rlabel metal2 s 312 4297 312 4297 4 wl0_10
rlabel metal2 s 312 3507 312 3507 4 wl0_8
<< properties >>
string FIXED_BBOX 0 0 624 7900
<< end >>
