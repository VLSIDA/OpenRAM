magic
tech sky130A
magscale 1 2
timestamp 1595931502
<< checkpaint >>
rect -780 -965 1791 1637
<< metal1 >>
rect 480 311 531 377
rect 480 295 515 311
tri 515 295 531 311 nw
<< end >>
