magic
tech sky130A
magscale 1 2
timestamp 1595931502
<< checkpaint >>
rect -1260 -1286 2058 1652
<< scnmos >>
rect 60 0 90 336
rect 168 0 198 336
rect 276 0 306 336
rect 384 0 414 336
rect 492 0 522 336
rect 600 0 630 336
rect 708 0 738 336
<< ndiff >>
rect 0 0 60 336
rect 90 0 168 336
rect 198 0 276 336
rect 306 0 384 336
rect 414 0 492 336
rect 522 0 600 336
rect 630 0 708 336
rect 738 0 798 336
<< poly >>
rect 60 362 738 392
rect 60 336 90 362
rect 168 336 198 362
rect 276 336 306 362
rect 384 336 414 362
rect 492 336 522 362
rect 600 336 630 362
rect 708 336 738 362
rect 60 -26 90 0
rect 168 -26 198 0
rect 276 -26 306 0
rect 384 -26 414 0
rect 492 -26 522 0
rect 600 -26 630 0
rect 708 -26 738 0
<< locali >>
rect 112 235 790 269
rect 8 135 42 201
rect 112 168 146 235
rect 220 135 254 201
rect 328 168 362 235
rect 436 135 470 201
rect 544 168 578 235
rect 652 135 686 201
rect 756 168 790 235
use contact_17  contact_17_0
timestamp 1595931502
transform 1 0 748 0 1 135
box 0 0 50 66
use contact_17  contact_17_1
timestamp 1595931502
transform 1 0 644 0 1 135
box 0 0 50 66
use contact_17  contact_17_2
timestamp 1595931502
transform 1 0 536 0 1 135
box 0 0 50 66
use contact_17  contact_17_3
timestamp 1595931502
transform 1 0 428 0 1 135
box 0 0 50 66
use contact_17  contact_17_4
timestamp 1595931502
transform 1 0 320 0 1 135
box 0 0 50 66
use contact_17  contact_17_5
timestamp 1595931502
transform 1 0 212 0 1 135
box 0 0 50 66
use contact_17  contact_17_6
timestamp 1595931502
transform 1 0 104 0 1 135
box 0 0 50 66
use contact_17  contact_17_7
timestamp 1595931502
transform 1 0 0 0 1 135
box 0 0 50 66
<< labels >>
rlabel poly s 399 377 399 377 4 G
rlabel corelocali s 669 168 669 168 4 S
rlabel corelocali s 453 168 453 168 4 S
rlabel corelocali s 237 168 237 168 4 S
rlabel corelocali s 25 168 25 168 4 S
rlabel corelocali s 451 252 451 252 4 D
<< properties >>
string FIXED_BBOX -25 -26 823 362
<< end >>
