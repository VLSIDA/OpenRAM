VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS
SITE  MacroSite
   CLASS Core ;
   SIZE 231500.0 by 299900.00000000006 ;
END  MacroSite
MACRO sram_2_16_scn4m_subm
   CLASS BLOCK ;
   SIZE 231500.0 BY 299900.00000000006 ;
   SYMMETRY X Y R90 ;
   SITE MacroSite ;
   PIN DIN0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  186200.0 8600.000000000002 187000.0 9400.000000000002 ;
      END
   END DIN0[0]
   PIN DIN0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  208000.0 8600.000000000002 208800.0 9400.000000000002 ;
      END
   END DIN0[1]
   PIN ADDR0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  56800.0 220500.0 57599.99999999999 221300.0 ;
      END
   END ADDR0[0]
   PIN ADDR0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  56800.0 242500.0 57599.99999999999 243300.0 ;
      END
   END ADDR0[1]
   PIN ADDR0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  56800.0 260500.0 57599.99999999999 261300.0 ;
      END
   END ADDR0[2]
   PIN ADDR0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  56800.0 282500.0 57599.99999999999 283300.0 ;
      END
   END ADDR0[3]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  7599.9999999999945 28200.000000000004 8399.99999999999 29000.000000000004 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  7599.9999999999945 50200.0 8399.99999999999 51000.0 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  36900.0 19600.0 37499.99999999999 29100.0 ;
      END
   END clk0
   PIN DOUT0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal2 ;
         RECT  179200.0 68800.00000000001 180000.0 71800.00000000001 ;
      END
   END DOUT0[0]
   PIN DOUT0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal2 ;
         RECT  186000.0 68800.00000000001 186800.0 71800.00000000001 ;
      END
   END DOUT0[1]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  181700.00000000003 131300.0 182300.0 131900.0 ;
         LAYER metal3 ;
         RECT  188500.0 131300.0 189100.00000000003 131900.0 ;
         LAYER metal3 ;
         RECT  181700.00000000003 149700.00000000003 182300.0 150300.0 ;
         LAYER metal3 ;
         RECT  188500.0 149700.00000000003 189100.00000000003 150300.0 ;
         LAYER metal3 ;
         RECT  181700.00000000003 168100.00000000003 182300.0 168700.00000000003 ;
         LAYER metal3 ;
         RECT  188500.0 168100.00000000003 189100.00000000003 168700.00000000003 ;
         LAYER metal3 ;
         RECT  181700.00000000003 186500.0 182300.0 187100.00000000003 ;
         LAYER metal3 ;
         RECT  188500.0 186500.0 189100.00000000003 187100.00000000003 ;
         LAYER metal3 ;
         RECT  181700.00000000003 204900.0 182300.0 205500.0 ;
         LAYER metal3 ;
         RECT  188500.0 204900.0 189100.00000000003 205500.0 ;
         LAYER metal3 ;
         RECT  181700.00000000003 223300.0 182300.0 223900.0 ;
         LAYER metal3 ;
         RECT  188500.0 223300.0 189100.00000000003 223900.0 ;
         LAYER metal3 ;
         RECT  181700.00000000003 241700.00000000003 182300.0 242300.0 ;
         LAYER metal3 ;
         RECT  188500.0 241700.00000000003 189100.00000000003 242300.0 ;
         LAYER metal3 ;
         RECT  181700.00000000003 260100.00000000003 182300.0 260700.0 ;
         LAYER metal3 ;
         RECT  188500.0 260100.00000000003 189100.00000000003 260700.0 ;
         LAYER metal3 ;
         RECT  181400.0 112000.0 182200.00000000003 112800.00000000001 ;
         LAYER metal3 ;
         RECT  188200.00000000003 112000.0 189000.0 112800.00000000001 ;
         LAYER metal3 ;
         RECT  184100.00000000003 81700.0 184700.00000000003 82300.00000000001 ;
         LAYER metal3 ;
         RECT  190900.0 81700.0 191500.0 82300.00000000001 ;
         LAYER metal3 ;
         RECT  182500.0 30500.0 183100.00000000003 31100.0 ;
         LAYER metal3 ;
         RECT  181900.0 47900.00000000001 182500.0 48500.0 ;
         LAYER metal3 ;
         RECT  189300.0 30500.0 189900.0 31100.0 ;
         LAYER metal3 ;
         RECT  188700.00000000003 47900.00000000001 189300.0 48500.0 ;
         LAYER metal3 ;
         RECT  130100.0 131600.0 130900.0 132400.0 ;
         LAYER metal3 ;
         RECT  130100.0 150000.0 130900.0 150800.0 ;
         LAYER metal3 ;
         RECT  130100.0 168400.0 130900.0 169200.00000000003 ;
         LAYER metal3 ;
         RECT  130100.0 186800.0 130900.0 187600.00000000003 ;
         LAYER metal3 ;
         RECT  130100.0 205200.00000000003 130900.0 206000.0 ;
         LAYER metal3 ;
         RECT  130100.0 223600.00000000003 130900.0 224400.0 ;
         LAYER metal3 ;
         RECT  130100.0 242000.0 130900.0 242800.0 ;
         LAYER metal3 ;
         RECT  130100.0 260400.00000000003 130900.0 261200.0 ;
         LAYER metal3 ;
         RECT  89700.0 131600.0 90500.0 132400.0 ;
         LAYER metal3 ;
         RECT  107700.0 131600.0 108500.0 132400.0 ;
         LAYER metal3 ;
         RECT  89700.0 150000.0 90500.0 150800.0 ;
         LAYER metal3 ;
         RECT  107700.0 150000.0 108500.0 150800.0 ;
         LAYER metal3 ;
         RECT  89700.0 168400.0 90500.0 169200.00000000003 ;
         LAYER metal3 ;
         RECT  107700.0 168400.0 108500.0 169200.00000000003 ;
         LAYER metal3 ;
         RECT  89700.0 186800.0 90500.0 187600.00000000003 ;
         LAYER metal3 ;
         RECT  107700.0 186800.0 108500.0 187600.00000000003 ;
         LAYER metal3 ;
         RECT  154400.0 131700.00000000003 155000.0 132300.0 ;
         LAYER metal3 ;
         RECT  164000.0 131700.00000000003 164600.00000000003 132300.0 ;
         LAYER metal3 ;
         RECT  154400.0 150100.0 155000.0 150700.00000000003 ;
         LAYER metal3 ;
         RECT  164000.0 150100.0 164600.00000000003 150700.00000000003 ;
         LAYER metal3 ;
         RECT  154400.0 168500.0 155000.0 169100.00000000003 ;
         LAYER metal3 ;
         RECT  164000.0 168500.0 164600.00000000003 169100.00000000003 ;
         LAYER metal3 ;
         RECT  154400.0 186900.0 155000.0 187500.0 ;
         LAYER metal3 ;
         RECT  164000.0 186900.0 164600.00000000003 187500.0 ;
         LAYER metal3 ;
         RECT  154400.0 205300.0 155000.0 205900.0 ;
         LAYER metal3 ;
         RECT  164000.0 205300.0 164600.00000000003 205900.0 ;
         LAYER metal3 ;
         RECT  154400.0 223700.00000000003 155000.0 224300.0 ;
         LAYER metal3 ;
         RECT  164000.0 223700.00000000003 164600.00000000003 224300.0 ;
         LAYER metal3 ;
         RECT  154400.0 242100.00000000003 155000.0 242700.00000000003 ;
         LAYER metal3 ;
         RECT  164000.0 242100.00000000003 164600.00000000003 242700.00000000003 ;
         LAYER metal3 ;
         RECT  154400.0 260500.0 155000.0 261100.00000000003 ;
         LAYER metal3 ;
         RECT  164000.0 260500.0 164600.00000000003 261100.00000000003 ;
         LAYER metal3 ;
         RECT  69200.0 39200.0 70000.0 40000.0 ;
         LAYER metal3 ;
         RECT  69200.0 79200.0 70000.0 80000.0 ;
         LAYER metal3 ;
         RECT  69200.0 119200.0 70000.0 120000.0 ;
         LAYER metal3 ;
         RECT  31500.0 142600.0 32100.0 143200.00000000003 ;
         LAYER metal3 ;
         RECT  31500.0 161000.0 32100.0 161600.00000000003 ;
         LAYER metal3 ;
         RECT  31500.0 179400.0 32100.0 180000.0 ;
         LAYER metal3 ;
         RECT  31500.0 197800.0 32100.0 198400.0 ;
         LAYER metal3 ;
         RECT  12400.0 142500.0 13200.000000000002 143300.0 ;
         LAYER metal3 ;
         RECT  18800.0 142500.0 19600.0 143300.0 ;
         LAYER metal3 ;
         RECT  12400.0 160900.0 13200.000000000002 161700.00000000003 ;
         LAYER metal3 ;
         RECT  18800.0 160900.0 19600.0 161700.00000000003 ;
         LAYER metal3 ;
         RECT  6000.0 124100.00000000001 6800.000000000001 124900.0 ;
         LAYER metal3 ;
         RECT  31400.000000000004 122700.0 32200.000000000004 123500.0 ;
         LAYER metal3 ;
         RECT  17200.0 129100.0 18000.0 129900.0 ;
         LAYER metal3 ;
         RECT  -400.0 39200.0 400.0 40000.0 ;
         LAYER metal3 ;
         RECT  59700.0 231500.0 60500.0 232300.0 ;
         LAYER metal3 ;
         RECT  59700.0 271500.0 60500.0 272300.0 ;
         LAYER metal3 ;
         RECT  189100.00000000003 19600.0 189900.0 20400.000000000004 ;
         LAYER metal3 ;
         RECT  210900.0 19600.0 211700.00000000003 20400.000000000004 ;
         LAYER metal3 ;
         RECT  0.0 3900.0000000000005 168000.0 8100.0 ;
         LAYER metal3 ;
         RECT  0.0 13500.0 232800.0 17700.0 ;
         LAYER metal3 ;
         RECT  0.0 23100.0 232800.0 27300.0 ;
         LAYER metal3 ;
         RECT  0.0 32700.000000000004 177600.00000000003 36900.0 ;
         LAYER metal3 ;
         RECT  194400.0 32700.000000000004 232800.0 36900.0 ;
         LAYER metal3 ;
         RECT  0.0 42300.00000000001 177600.00000000003 46500.0 ;
         LAYER metal3 ;
         RECT  196800.0 42300.00000000001 232800.0 46500.0 ;
         LAYER metal3 ;
         RECT  0.0 51900.00000000001 177600.00000000003 56100.0 ;
         LAYER metal3 ;
         RECT  196800.0 51900.00000000001 232800.0 56100.0 ;
         LAYER metal3 ;
         RECT  0.0 61500.0 232800.0 65700.0 ;
         LAYER metal3 ;
         RECT  0.0 71100.00000000001 232800.0 75300.0 ;
         LAYER metal3 ;
         RECT  0.0 80700.0 232800.0 84900.0 ;
         LAYER metal3 ;
         RECT  52800.00000000001 90300.00000000001 180000.0 94500.0 ;
         LAYER metal3 ;
         RECT  196800.0 90300.00000000001 232800.0 94500.0 ;
         LAYER metal3 ;
         RECT  0.0 99900.0 64800.0 104100.00000000001 ;
         LAYER metal3 ;
         RECT  74400.0 99900.0 232800.0 104100.00000000001 ;
         LAYER metal3 ;
         RECT  0.0 109500.0 64800.0 113700.0 ;
         LAYER metal3 ;
         RECT  182400.0 109500.0 232800.0 113700.0 ;
         LAYER metal3 ;
         RECT  0.0 119100.00000000001 84000.0 123300.00000000001 ;
         LAYER metal3 ;
         RECT  170400.0 119100.00000000001 232800.0 123300.00000000001 ;
         LAYER metal3 ;
         RECT  40800.00000000001 128700.00000000001 69600.00000000001 132900.0 ;
         LAYER metal3 ;
         RECT  86400.0 128700.00000000001 105600.00000000001 132900.0 ;
         LAYER metal3 ;
         RECT  120000.0 128700.00000000001 232800.0 132900.0 ;
         LAYER metal3 ;
         RECT  40800.00000000001 138300.0 69600.00000000001 142500.0 ;
         LAYER metal3 ;
         RECT  170400.0 138300.0 232800.0 142500.0 ;
         LAYER metal3 ;
         RECT  43200.0 147900.0 105600.00000000001 152100.0 ;
         LAYER metal3 ;
         RECT  122400.0 147900.0 232800.0 152100.0 ;
         LAYER metal3 ;
         RECT  40800.00000000001 157500.0 84000.0 161700.00000000003 ;
         LAYER metal3 ;
         RECT  170400.0 157500.0 232800.0 161700.00000000003 ;
         LAYER metal3 ;
         RECT  43200.0 167100.00000000003 72000.0 171300.0 ;
         LAYER metal3 ;
         RECT  86400.0 167100.00000000003 105600.00000000001 171300.0 ;
         LAYER metal3 ;
         RECT  127200.0 167100.00000000003 232800.0 171300.0 ;
         LAYER metal3 ;
         RECT  0.0 176700.00000000003 72000.0 180900.0 ;
         LAYER metal3 ;
         RECT  170400.0 176700.00000000003 232800.0 180900.0 ;
         LAYER metal3 ;
         RECT  0.0 186300.0 31200.000000000004 190500.0 ;
         LAYER metal3 ;
         RECT  43200.0 186300.0 105600.00000000001 190500.0 ;
         LAYER metal3 ;
         RECT  129600.0 186300.0 172800.0 190500.0 ;
         LAYER metal3 ;
         RECT  196800.0 186300.0 232800.0 190500.0 ;
         LAYER metal3 ;
         RECT  0.0 195900.0 84000.0 200100.00000000003 ;
         LAYER metal3 ;
         RECT  196800.0 195900.0 232800.0 200100.00000000003 ;
         LAYER metal3 ;
         RECT  0.0 205500.0 31200.000000000004 209700.00000000003 ;
         LAYER metal3 ;
         RECT  43200.0 205500.0 172800.0 209700.00000000003 ;
         LAYER metal3 ;
         RECT  196800.0 205500.0 232800.0 209700.00000000003 ;
         LAYER metal3 ;
         RECT  0.0 215100.00000000003 43200.0 219300.0 ;
         LAYER metal3 ;
         RECT  76800.00000000001 215100.00000000003 124800.00000000001 219300.0 ;
         LAYER metal3 ;
         RECT  196800.0 215100.00000000003 232800.0 219300.0 ;
         LAYER metal3 ;
         RECT  0.0 224700.00000000003 172800.0 228900.0 ;
         LAYER metal3 ;
         RECT  196800.0 224700.00000000003 232800.0 228900.0 ;
         LAYER metal3 ;
         RECT  0.0 234300.0 172800.0 238500.0 ;
         LAYER metal3 ;
         RECT  196800.0 234300.0 232800.0 238500.0 ;
         LAYER metal3 ;
         RECT  0.0 243900.0 172800.0 248100.00000000003 ;
         LAYER metal3 ;
         RECT  196800.0 243900.0 232800.0 248100.00000000003 ;
         LAYER metal3 ;
         RECT  0.0 253500.0 172800.0 257700.0 ;
         LAYER metal3 ;
         RECT  196800.0 253500.0 232800.0 257700.0 ;
         LAYER metal3 ;
         RECT  0.0 263100.0 172800.0 267300.0 ;
         LAYER metal3 ;
         RECT  196800.0 263100.0 232800.0 267300.0 ;
         LAYER metal3 ;
         RECT  0.0 272700.0 232800.0 276900.00000000006 ;
         LAYER metal3 ;
         RECT  0.0 282300.0 62400.00000000001 286500.0 ;
         LAYER metal3 ;
         RECT  84000.0 282300.0 232800.0 286500.0 ;
         LAYER metal3 ;
         RECT  0.0 291900.00000000006 55200.0 296100.0 ;
         LAYER metal3 ;
         RECT  64800.0 291900.00000000006 232800.0 296100.0 ;
         LAYER metal4 ;
         RECT  4200.0 0.0 7800.000000000001 302400.00000000006 ;
         LAYER metal4 ;
         RECT  13800.0 0.0 17400.000000000004 302400.00000000006 ;
         LAYER metal4 ;
         RECT  23400.000000000004 0.0 27000.0 302400.00000000006 ;
         LAYER metal4 ;
         RECT  33000.0 0.0 36600.0 302400.00000000006 ;
         LAYER metal4 ;
         RECT  42600.0 0.0 46200.0 302400.00000000006 ;
         LAYER metal4 ;
         RECT  52200.0 0.0 55800.00000000001 302400.00000000006 ;
         LAYER metal4 ;
         RECT  61800.00000000001 0.0 65400.00000000001 302400.00000000006 ;
         LAYER metal4 ;
         RECT  71400.0 0.0 75000.0 302400.00000000006 ;
         LAYER metal4 ;
         RECT  81000.0 0.0 84600.00000000001 302400.00000000006 ;
         LAYER metal4 ;
         RECT  90600.00000000001 0.0 94200.0 302400.00000000006 ;
         LAYER metal4 ;
         RECT  100200.0 0.0 103800.00000000001 302400.00000000006 ;
         LAYER metal4 ;
         RECT  109800.00000000001 0.0 113400.0 302400.00000000006 ;
         LAYER metal4 ;
         RECT  119400.0 0.0 123000.0 302400.00000000006 ;
         LAYER metal4 ;
         RECT  129000.0 0.0 132600.0 302400.00000000006 ;
         LAYER metal4 ;
         RECT  138600.0 0.0 142200.00000000003 302400.00000000006 ;
         LAYER metal4 ;
         RECT  148200.00000000003 0.0 151800.0 302400.00000000006 ;
         LAYER metal4 ;
         RECT  157800.0 0.0 161400.0 302400.00000000006 ;
         LAYER metal4 ;
         RECT  167400.0 0.0 171000.0 302400.00000000006 ;
         LAYER metal4 ;
         RECT  177000.0 0.0 180600.00000000003 302400.00000000006 ;
         LAYER metal4 ;
         RECT  186600.00000000003 0.0 190200.00000000003 302400.00000000006 ;
         LAYER metal4 ;
         RECT  196200.00000000003 0.0 199800.0 302400.00000000006 ;
         LAYER metal4 ;
         RECT  205800.0 0.0 209400.0 302400.00000000006 ;
         LAYER metal4 ;
         RECT  215400.0 0.0 219000.0 302400.00000000006 ;
         LAYER metal4 ;
         RECT  225000.0 0.0 228600.00000000003 302400.00000000006 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  178300.0 126700.0 178900.0 127300.00000000001 ;
         LAYER metal3 ;
         RECT  185100.00000000003 126700.0 185700.00000000003 127300.00000000001 ;
         LAYER metal3 ;
         RECT  191900.0 126700.0 192500.0 127300.00000000001 ;
         LAYER metal3 ;
         RECT  178300.0 135900.0 178900.0 136500.0 ;
         LAYER metal3 ;
         RECT  185100.00000000003 135900.0 185700.00000000003 136500.0 ;
         LAYER metal3 ;
         RECT  191900.0 135900.0 192500.0 136500.0 ;
         LAYER metal3 ;
         RECT  178300.0 145100.0 178900.0 145700.00000000003 ;
         LAYER metal3 ;
         RECT  185100.00000000003 145100.0 185700.00000000003 145700.00000000003 ;
         LAYER metal3 ;
         RECT  191900.0 145100.0 192500.0 145700.00000000003 ;
         LAYER metal3 ;
         RECT  178300.0 154300.0 178900.0 154900.0 ;
         LAYER metal3 ;
         RECT  185100.00000000003 154300.0 185700.00000000003 154900.0 ;
         LAYER metal3 ;
         RECT  191900.0 154300.0 192500.0 154900.0 ;
         LAYER metal3 ;
         RECT  178300.0 163500.0 178900.0 164100.00000000003 ;
         LAYER metal3 ;
         RECT  185100.00000000003 163500.0 185700.00000000003 164100.00000000003 ;
         LAYER metal3 ;
         RECT  191900.0 163500.0 192500.0 164100.00000000003 ;
         LAYER metal3 ;
         RECT  178300.0 172700.00000000003 178900.0 173300.0 ;
         LAYER metal3 ;
         RECT  185100.00000000003 172700.00000000003 185700.00000000003 173300.0 ;
         LAYER metal3 ;
         RECT  191900.0 172700.00000000003 192500.0 173300.0 ;
         LAYER metal3 ;
         RECT  178300.0 181900.0 178900.0 182500.0 ;
         LAYER metal3 ;
         RECT  185100.00000000003 181900.0 185700.00000000003 182500.0 ;
         LAYER metal3 ;
         RECT  191900.0 181900.0 192500.0 182500.0 ;
         LAYER metal3 ;
         RECT  178300.0 191100.00000000003 178900.0 191700.00000000003 ;
         LAYER metal3 ;
         RECT  185100.00000000003 191100.00000000003 185700.00000000003 191700.00000000003 ;
         LAYER metal3 ;
         RECT  191900.0 191100.00000000003 192500.0 191700.00000000003 ;
         LAYER metal3 ;
         RECT  178300.0 200300.0 178900.0 200900.0 ;
         LAYER metal3 ;
         RECT  185100.00000000003 200300.0 185700.00000000003 200900.0 ;
         LAYER metal3 ;
         RECT  191900.0 200300.0 192500.0 200900.0 ;
         LAYER metal3 ;
         RECT  178300.0 209500.0 178900.0 210100.00000000003 ;
         LAYER metal3 ;
         RECT  185100.00000000003 209500.0 185700.00000000003 210100.00000000003 ;
         LAYER metal3 ;
         RECT  191900.0 209500.0 192500.0 210100.00000000003 ;
         LAYER metal3 ;
         RECT  178300.0 218700.00000000003 178900.0 219300.0 ;
         LAYER metal3 ;
         RECT  185100.00000000003 218700.00000000003 185700.00000000003 219300.0 ;
         LAYER metal3 ;
         RECT  191900.0 218700.00000000003 192500.0 219300.0 ;
         LAYER metal3 ;
         RECT  178300.0 227900.0 178900.0 228500.0 ;
         LAYER metal3 ;
         RECT  185100.00000000003 227900.0 185700.00000000003 228500.0 ;
         LAYER metal3 ;
         RECT  191900.0 227900.0 192500.0 228500.0 ;
         LAYER metal3 ;
         RECT  178300.0 237100.00000000003 178900.0 237700.00000000003 ;
         LAYER metal3 ;
         RECT  185100.00000000003 237100.00000000003 185700.00000000003 237700.00000000003 ;
         LAYER metal3 ;
         RECT  191900.0 237100.00000000003 192500.0 237700.00000000003 ;
         LAYER metal3 ;
         RECT  178300.0 246300.0 178900.0 246900.0 ;
         LAYER metal3 ;
         RECT  185100.00000000003 246300.0 185700.00000000003 246900.0 ;
         LAYER metal3 ;
         RECT  191900.0 246300.0 192500.0 246900.0 ;
         LAYER metal3 ;
         RECT  178300.0 255500.0 178900.0 256100.00000000003 ;
         LAYER metal3 ;
         RECT  185100.00000000003 255500.0 185700.00000000003 256100.00000000003 ;
         LAYER metal3 ;
         RECT  191900.0 255500.0 192500.0 256100.00000000003 ;
         LAYER metal3 ;
         RECT  178300.0 264700.0 178900.0 265300.0 ;
         LAYER metal3 ;
         RECT  185100.00000000003 264700.0 185700.00000000003 265300.0 ;
         LAYER metal3 ;
         RECT  191900.0 264700.0 192500.0 265300.0 ;
         LAYER metal3 ;
         RECT  185100.00000000003 95100.00000000001 185700.00000000003 95700.0 ;
         LAYER metal3 ;
         RECT  191900.0 95100.00000000001 192500.0 95700.0 ;
         LAYER metal3 ;
         RECT  182500.0 37100.0 183100.00000000003 37700.0 ;
         LAYER metal3 ;
         RECT  183900.0 41500.0 184500.0 42100.0 ;
         LAYER metal3 ;
         RECT  183300.0 54900.00000000001 183900.0 55500.0 ;
         LAYER metal3 ;
         RECT  189300.0 37100.0 189900.0 37700.0 ;
         LAYER metal3 ;
         RECT  190700.00000000003 41500.0 191300.0 42100.0 ;
         LAYER metal3 ;
         RECT  190100.00000000003 54900.00000000001 190700.00000000003 55500.0 ;
         LAYER metal3 ;
         RECT  130100.0 122400.0 130900.0 123200.0 ;
         LAYER metal3 ;
         RECT  130100.0 140800.0 130900.0 141600.0 ;
         LAYER metal3 ;
         RECT  130100.0 159200.00000000003 130900.0 160000.0 ;
         LAYER metal3 ;
         RECT  130100.0 177600.00000000003 130900.0 178400.0 ;
         LAYER metal3 ;
         RECT  130100.0 196000.0 130900.0 196800.0 ;
         LAYER metal3 ;
         RECT  130100.0 214400.0 130900.0 215200.00000000003 ;
         LAYER metal3 ;
         RECT  130100.0 232800.0 130900.0 233600.00000000003 ;
         LAYER metal3 ;
         RECT  130100.0 251200.00000000003 130900.0 252000.0 ;
         LAYER metal3 ;
         RECT  130100.0 269600.0 130900.0 270400.00000000006 ;
         LAYER metal3 ;
         RECT  89700.0 122400.0 90500.0 123200.0 ;
         LAYER metal3 ;
         RECT  107700.0 122400.0 108500.0 123200.0 ;
         LAYER metal3 ;
         RECT  89700.0 140800.0 90500.0 141600.0 ;
         LAYER metal3 ;
         RECT  107700.0 140800.0 108500.0 141600.0 ;
         LAYER metal3 ;
         RECT  89700.0 159200.00000000003 90500.0 160000.0 ;
         LAYER metal3 ;
         RECT  107700.0 159200.00000000003 108500.0 160000.0 ;
         LAYER metal3 ;
         RECT  89700.0 177600.00000000003 90500.0 178400.0 ;
         LAYER metal3 ;
         RECT  107700.0 177600.00000000003 108500.0 178400.0 ;
         LAYER metal3 ;
         RECT  89700.0 196000.0 90500.0 196800.0 ;
         LAYER metal3 ;
         RECT  107700.0 196000.0 108500.0 196800.0 ;
         LAYER metal3 ;
         RECT  154400.0 122500.0 155000.0 123100.00000000001 ;
         LAYER metal3 ;
         RECT  164000.0 122500.0 164600.00000000003 123100.00000000001 ;
         LAYER metal3 ;
         RECT  154400.0 140900.0 155000.0 141500.0 ;
         LAYER metal3 ;
         RECT  164000.0 140900.0 164600.00000000003 141500.0 ;
         LAYER metal3 ;
         RECT  154400.0 159300.0 155000.0 159900.0 ;
         LAYER metal3 ;
         RECT  164000.0 159300.0 164600.00000000003 159900.0 ;
         LAYER metal3 ;
         RECT  154400.0 177700.00000000003 155000.0 178300.0 ;
         LAYER metal3 ;
         RECT  164000.0 177700.00000000003 164600.00000000003 178300.0 ;
         LAYER metal3 ;
         RECT  154400.0 196100.00000000003 155000.0 196700.00000000003 ;
         LAYER metal3 ;
         RECT  164000.0 196100.00000000003 164600.00000000003 196700.00000000003 ;
         LAYER metal3 ;
         RECT  154400.0 214500.0 155000.0 215100.00000000003 ;
         LAYER metal3 ;
         RECT  164000.0 214500.0 164600.00000000003 215100.00000000003 ;
         LAYER metal3 ;
         RECT  154400.0 232900.0 155000.0 233500.0 ;
         LAYER metal3 ;
         RECT  164000.0 232900.0 164600.00000000003 233500.0 ;
         LAYER metal3 ;
         RECT  154400.0 251300.0 155000.0 251900.0 ;
         LAYER metal3 ;
         RECT  164000.0 251300.0 164600.00000000003 251900.0 ;
         LAYER metal3 ;
         RECT  154400.0 269700.0 155000.0 270300.0 ;
         LAYER metal3 ;
         RECT  164000.0 269700.0 164600.00000000003 270300.0 ;
         LAYER metal3 ;
         RECT  69200.0 59200.0 70000.0 60000.0 ;
         LAYER metal3 ;
         RECT  69200.0 19200.000000000004 70000.0 20000.0 ;
         LAYER metal3 ;
         RECT  69200.0 99200.0 70000.0 100000.0 ;
         LAYER metal3 ;
         RECT  28100.0 138000.0 28700.000000000004 138600.0 ;
         LAYER metal3 ;
         RECT  34900.0 138000.0 35500.0 138600.0 ;
         LAYER metal3 ;
         RECT  28100.0 147200.00000000003 28700.000000000004 147800.0 ;
         LAYER metal3 ;
         RECT  34900.0 147200.00000000003 35500.0 147800.0 ;
         LAYER metal3 ;
         RECT  28100.0 156400.0 28700.000000000004 157000.0 ;
         LAYER metal3 ;
         RECT  34900.0 156400.0 35500.0 157000.0 ;
         LAYER metal3 ;
         RECT  28100.0 165600.00000000003 28700.000000000004 166200.00000000003 ;
         LAYER metal3 ;
         RECT  34900.0 165600.00000000003 35500.0 166200.00000000003 ;
         LAYER metal3 ;
         RECT  28100.0 174800.0 28700.000000000004 175400.0 ;
         LAYER metal3 ;
         RECT  34900.0 174800.0 35500.0 175400.0 ;
         LAYER metal3 ;
         RECT  28100.0 184000.0 28700.000000000004 184600.00000000003 ;
         LAYER metal3 ;
         RECT  34900.0 184000.0 35500.0 184600.00000000003 ;
         LAYER metal3 ;
         RECT  28100.0 193200.00000000003 28700.000000000004 193800.0 ;
         LAYER metal3 ;
         RECT  34900.0 193200.00000000003 35500.0 193800.0 ;
         LAYER metal3 ;
         RECT  28100.0 202400.0 28700.000000000004 203000.0 ;
         LAYER metal3 ;
         RECT  34900.0 202400.0 35500.0 203000.0 ;
         LAYER metal3 ;
         RECT  12400.0 133300.0 13200.000000000002 134100.0 ;
         LAYER metal3 ;
         RECT  18800.0 133300.0 19600.0 134100.0 ;
         LAYER metal3 ;
         RECT  12400.0 151700.00000000003 13200.000000000002 152500.0 ;
         LAYER metal3 ;
         RECT  18800.0 151700.00000000003 19600.0 152500.0 ;
         LAYER metal3 ;
         RECT  12400.0 170100.00000000003 13200.000000000002 170900.0 ;
         LAYER metal3 ;
         RECT  18800.0 170100.00000000003 19600.0 170900.0 ;
         LAYER metal3 ;
         RECT  28000.0 128700.00000000001 28800.0 129500.0 ;
         LAYER metal3 ;
         RECT  34800.00000000001 128700.00000000001 35600.0 129500.0 ;
         LAYER metal3 ;
         RECT  36400.0 134700.00000000003 37200.0 135500.0 ;
         LAYER metal3 ;
         RECT  36400.0 150300.0 37200.0 151100.0 ;
         LAYER metal3 ;
         RECT  36400.0 153100.0 37200.0 153900.0 ;
         LAYER metal3 ;
         RECT  36400.0 168700.00000000003 37200.0 169500.0 ;
         LAYER metal3 ;
         RECT  36400.0 171500.0 37200.0 172300.0 ;
         LAYER metal3 ;
         RECT  36400.0 187100.00000000003 37200.0 187900.0 ;
         LAYER metal3 ;
         RECT  36400.0 189900.0 37200.0 190700.00000000003 ;
         LAYER metal3 ;
         RECT  36400.0 205500.0 37200.0 206300.0 ;
         LAYER metal3 ;
         RECT  -400.0 19200.000000000004 400.0 20000.0 ;
         LAYER metal3 ;
         RECT  -400.0 59200.0 400.0 60000.0 ;
         LAYER metal3 ;
         RECT  59700.0 211500.0 60500.0 212300.0 ;
         LAYER metal3 ;
         RECT  59700.0 251500.0 60500.0 252300.0 ;
         LAYER metal3 ;
         RECT  59700.0 291500.0 60500.0 292300.0 ;
         LAYER metal3 ;
         RECT  189100.00000000003 -400.0 189900.0 400.0 ;
         LAYER metal3 ;
         RECT  210900.0 -400.0 211700.00000000003 400.0 ;
         LAYER metal3 ;
         RECT  0.0 -900.0 168000.0 3300.0000000000005 ;
         LAYER metal3 ;
         RECT  0.0 8700.000000000002 232800.0 12900.0 ;
         LAYER metal3 ;
         RECT  0.0 18300.0 184800.0 22500.0 ;
         LAYER metal3 ;
         RECT  216000.0 18300.0 232800.0 22500.0 ;
         LAYER metal3 ;
         RECT  194400.0 27900.000000000004 232800.0 32100.0 ;
         LAYER metal3 ;
         RECT  4800.000000000001 37500.0 64800.0 41700.0 ;
         LAYER metal3 ;
         RECT  74400.0 37500.0 232800.0 41700.0 ;
         LAYER metal3 ;
         RECT  194400.0 47100.0 232800.0 51300.00000000001 ;
         LAYER metal3 ;
         RECT  0.0 56700.0 232800.0 60900.00000000001 ;
         LAYER metal3 ;
         RECT  0.0 66300.0 64800.0 70500.0 ;
         LAYER metal3 ;
         RECT  180000.0 66300.0 232800.0 70500.0 ;
         LAYER metal3 ;
         RECT  0.0 75900.0 64800.0 80100.00000000001 ;
         LAYER metal3 ;
         RECT  74400.0 75900.0 232800.0 80100.00000000001 ;
         LAYER metal3 ;
         RECT  52800.00000000001 85500.0 232800.0 89700.0 ;
         LAYER metal3 ;
         RECT  0.0 95100.00000000001 232800.0 99300.00000000001 ;
         LAYER metal3 ;
         RECT  0.0 104700.0 64800.0 108900.0 ;
         LAYER metal3 ;
         RECT  182400.0 104700.0 232800.0 108900.0 ;
         LAYER metal3 ;
         RECT  0.0 114300.00000000001 232800.0 118500.0 ;
         LAYER metal3 ;
         RECT  38400.00000000001 123900.0 232800.0 128100.0 ;
         LAYER metal3 ;
         RECT  26400.000000000004 133500.0 69600.00000000001 137700.00000000003 ;
         LAYER metal3 ;
         RECT  86400.0 133500.0 232800.0 137700.00000000003 ;
         LAYER metal3 ;
         RECT  38400.00000000001 143100.0 69600.00000000001 147300.0 ;
         LAYER metal3 ;
         RECT  88800.00000000001 143100.0 232800.0 147300.0 ;
         LAYER metal3 ;
         RECT  26400.000000000004 152700.00000000003 232800.0 156900.0 ;
         LAYER metal3 ;
         RECT  38400.00000000001 162300.0 232800.0 166500.0 ;
         LAYER metal3 ;
         RECT  0.0 171900.0 232800.0 176100.00000000003 ;
         LAYER metal3 ;
         RECT  0.0 181500.0 232800.0 185700.00000000003 ;
         LAYER metal3 ;
         RECT  0.0 191100.00000000003 232800.0 195300.0 ;
         LAYER metal3 ;
         RECT  0.0 200700.00000000003 124800.00000000001 204900.0 ;
         LAYER metal3 ;
         RECT  194400.0 200700.00000000003 232800.0 204900.0 ;
         LAYER metal3 ;
         RECT  0.0 210300.0 43200.0 214500.0 ;
         LAYER metal3 ;
         RECT  76800.00000000001 210300.0 232800.0 214500.0 ;
         LAYER metal3 ;
         RECT  0.0 219900.0 62400.00000000001 224100.00000000003 ;
         LAYER metal3 ;
         RECT  79200.0 219900.0 124800.00000000001 224100.00000000003 ;
         LAYER metal3 ;
         RECT  194400.0 219900.0 232800.0 224100.00000000003 ;
         LAYER metal3 ;
         RECT  0.0 229500.0 55200.0 233700.00000000003 ;
         LAYER metal3 ;
         RECT  64800.0 229500.0 232800.0 233700.00000000003 ;
         LAYER metal3 ;
         RECT  0.0 239100.00000000003 62400.00000000001 243300.0 ;
         LAYER metal3 ;
         RECT  81600.00000000001 239100.00000000003 124800.00000000001 243300.0 ;
         LAYER metal3 ;
         RECT  194400.0 239100.00000000003 232800.0 243300.0 ;
         LAYER metal3 ;
         RECT  0.0 248700.00000000003 232800.0 252900.0 ;
         LAYER metal3 ;
         RECT  0.0 258300.0 62400.00000000001 262500.0 ;
         LAYER metal3 ;
         RECT  81600.00000000001 258300.0 124800.00000000001 262500.0 ;
         LAYER metal3 ;
         RECT  194400.0 258300.0 232800.0 262500.0 ;
         LAYER metal3 ;
         RECT  0.0 267900.00000000006 55200.0 272100.0 ;
         LAYER metal3 ;
         RECT  64800.0 267900.00000000006 232800.0 272100.0 ;
         LAYER metal3 ;
         RECT  0.0 277500.0 62400.00000000001 281700.0 ;
         LAYER metal3 ;
         RECT  84000.0 277500.0 232800.0 281700.0 ;
         LAYER metal3 ;
         RECT  0.0 287100.0 232800.0 291300.0 ;
         LAYER metal3 ;
         RECT  0.0 296700.0 232800.0 300900.00000000006 ;
         LAYER metal4 ;
         RECT  -600.0000000000001 0.0 3000.0 302400.00000000006 ;
         LAYER metal4 ;
         RECT  9000.0 0.0 12600.000000000002 302400.00000000006 ;
         LAYER metal4 ;
         RECT  18600.0 0.0 22200.000000000004 302400.00000000006 ;
         LAYER metal4 ;
         RECT  28200.000000000004 0.0 31800.0 302400.00000000006 ;
         LAYER metal4 ;
         RECT  37800.00000000001 0.0 41400.00000000001 302400.00000000006 ;
         LAYER metal4 ;
         RECT  47400.00000000001 0.0 51000.0 302400.00000000006 ;
         LAYER metal4 ;
         RECT  57000.0 0.0 60600.0 302400.00000000006 ;
         LAYER metal4 ;
         RECT  66600.00000000001 0.0 70200.0 302400.00000000006 ;
         LAYER metal4 ;
         RECT  76200.0 0.0 79800.00000000001 302400.00000000006 ;
         LAYER metal4 ;
         RECT  85800.00000000001 0.0 89400.0 302400.00000000006 ;
         LAYER metal4 ;
         RECT  95400.0 0.0 99000.0 302400.00000000006 ;
         LAYER metal4 ;
         RECT  105000.0 0.0 108600.00000000001 302400.00000000006 ;
         LAYER metal4 ;
         RECT  114600.00000000001 0.0 118200.0 302400.00000000006 ;
         LAYER metal4 ;
         RECT  124200.0 0.0 127800.00000000001 302400.00000000006 ;
         LAYER metal4 ;
         RECT  133800.0 0.0 137400.0 302400.00000000006 ;
         LAYER metal4 ;
         RECT  143400.0 0.0 147000.0 302400.00000000006 ;
         LAYER metal4 ;
         RECT  153000.0 0.0 156600.00000000003 302400.00000000006 ;
         LAYER metal4 ;
         RECT  162600.00000000003 0.0 166200.00000000003 302400.00000000006 ;
         LAYER metal4 ;
         RECT  172200.00000000003 0.0 175800.0 302400.00000000006 ;
         LAYER metal4 ;
         RECT  181800.0 0.0 185400.0 302400.00000000006 ;
         LAYER metal4 ;
         RECT  191400.0 0.0 195000.0 302400.00000000006 ;
         LAYER metal4 ;
         RECT  201000.0 0.0 204600.00000000003 302400.00000000006 ;
         LAYER metal4 ;
         RECT  210600.00000000003 0.0 214200.00000000003 302400.00000000006 ;
         LAYER metal4 ;
         RECT  220200.00000000003 0.0 223800.0 302400.00000000006 ;
         LAYER metal4 ;
         RECT  229800.0 0.0 233400.0 302400.00000000006 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  182000.0 22500.000000000004 197800.0 23100.000000000004 ;
      RECT  182000.0 22500.000000000004 189900.0 23100.000000000004 ;
      RECT  189900.0 22500.000000000004 197800.0 23100.000000000004 ;
      RECT  188800.0 23900.000000000004 219600.00000000003 24500.000000000004 ;
      RECT  188800.0 23900.000000000004 204200.00000000003 24500.000000000004 ;
      RECT  204200.0 23900.000000000004 219600.0 24500.000000000004 ;
      RECT  141300.0 126900.0 141899.99999999997 127500.0 ;
      RECT  141300.0 125300.00000000001 141899.99999999997 125900.0 ;
      RECT  139200.0 126900.0 141600.00000000003 127500.0 ;
      RECT  141300.0 125600.00000000001 141899.99999999997 127200.0 ;
      RECT  141600.00000000003 125300.00000000001 144100.00000000003 125900.0 ;
      RECT  172900.0 126900.0 173500.0 127500.0 ;
      RECT  172900.0 123500.0 173500.0 124100.0 ;
      RECT  168200.0 126900.0 173200.0 127500.0 ;
      RECT  172900.0 123800.00000000001 173500.0 127200.00000000001 ;
      RECT  173200.0 123500.0 178200.0 124100.0 ;
      RECT  141300.0 136500.0 141899.99999999997 137100.00000000003 ;
      RECT  141300.0 138100.00000000003 141899.99999999997 138700.0 ;
      RECT  139200.0 136500.0 141600.00000000003 137100.00000000003 ;
      RECT  141300.0 136800.0 141899.99999999997 138400.0 ;
      RECT  141600.00000000003 138100.00000000003 144100.00000000003 138700.0 ;
      RECT  172900.0 136500.0 173500.0 137100.00000000003 ;
      RECT  172900.0 139100.00000000003 173500.0 139700.0 ;
      RECT  168200.0 136500.0 173200.0 137100.00000000003 ;
      RECT  172900.0 136800.0 173500.0 139400.0 ;
      RECT  173200.0 139100.00000000003 178200.0 139700.0 ;
      RECT  141300.0 145300.0 141899.99999999997 145900.0 ;
      RECT  141300.0 143700.0 141899.99999999997 144300.0 ;
      RECT  139200.0 145300.0 141600.00000000003 145900.0 ;
      RECT  141300.0 144000.0 141899.99999999997 145600.00000000003 ;
      RECT  141600.00000000003 143700.0 144100.00000000003 144300.0 ;
      RECT  172900.0 145300.0 173500.0 145900.0 ;
      RECT  172900.0 141900.0 173500.0 142500.0 ;
      RECT  168200.0 145300.0 173200.0 145900.0 ;
      RECT  172900.0 142200.0 173500.0 145600.00000000003 ;
      RECT  173200.0 141900.0 178200.0 142500.0 ;
      RECT  141300.0 154899.99999999997 141899.99999999997 155500.0 ;
      RECT  141300.0 156500.0 141899.99999999997 157100.00000000003 ;
      RECT  139200.0 154899.99999999997 141600.00000000003 155500.0 ;
      RECT  141300.0 155200.0 141899.99999999997 156800.0 ;
      RECT  141600.00000000003 156500.0 144100.00000000003 157100.00000000003 ;
      RECT  172900.0 154899.99999999997 173500.0 155500.0 ;
      RECT  172900.0 157500.0 173500.0 158100.00000000003 ;
      RECT  168200.0 154899.99999999997 173200.0 155500.0 ;
      RECT  172900.0 155200.0 173500.0 157800.0 ;
      RECT  173200.0 157500.0 178200.0 158100.00000000003 ;
      RECT  141300.0 163700.0 141899.99999999997 164300.0 ;
      RECT  141300.0 162100.00000000003 141899.99999999997 162700.0 ;
      RECT  139200.0 163700.0 141600.00000000003 164300.0 ;
      RECT  141300.0 162399.99999999997 141899.99999999997 164000.0 ;
      RECT  141600.00000000003 162100.00000000003 144100.00000000003 162700.0 ;
      RECT  172900.0 163700.0 173500.0 164300.0 ;
      RECT  172900.0 160300.0 173500.0 160899.99999999997 ;
      RECT  168200.0 163700.0 173200.0 164300.0 ;
      RECT  172900.0 160600.00000000003 173500.0 164000.0 ;
      RECT  173200.0 160300.0 178200.0 160899.99999999997 ;
      RECT  141300.0 173300.0 141899.99999999997 173900.00000000003 ;
      RECT  141300.0 174899.99999999997 141899.99999999997 175500.0 ;
      RECT  139200.0 173300.0 141600.00000000003 173900.00000000003 ;
      RECT  141300.0 173600.00000000003 141899.99999999997 175200.0 ;
      RECT  141600.00000000003 174899.99999999997 144100.00000000003 175500.0 ;
      RECT  172900.0 173300.0 173500.0 173900.00000000003 ;
      RECT  172900.0 175899.99999999997 173500.0 176500.0 ;
      RECT  168200.0 173300.0 173200.0 173900.00000000003 ;
      RECT  172900.0 173600.00000000003 173500.0 176200.0 ;
      RECT  173200.0 175899.99999999997 178200.0 176500.0 ;
      RECT  141300.0 182100.00000000003 141899.99999999997 182700.0 ;
      RECT  141300.0 180500.0 141899.99999999997 181100.00000000003 ;
      RECT  139200.0 182100.00000000003 141600.00000000003 182700.0 ;
      RECT  141300.0 180800.0 141899.99999999997 182400.00000000003 ;
      RECT  141600.00000000003 180500.0 144100.00000000003 181100.00000000003 ;
      RECT  172900.0 182100.00000000003 173500.0 182700.0 ;
      RECT  172900.0 178700.0 173500.0 179300.0 ;
      RECT  168200.0 182100.00000000003 173200.0 182700.0 ;
      RECT  172900.0 179000.0 173500.0 182400.00000000003 ;
      RECT  173200.0 178700.0 178200.0 179300.0 ;
      RECT  141300.0 191700.0 141899.99999999997 192300.0 ;
      RECT  141300.0 193300.0 141899.99999999997 193900.00000000003 ;
      RECT  139200.0 191700.0 141600.00000000003 192300.0 ;
      RECT  141300.0 192000.0 141899.99999999997 193600.00000000003 ;
      RECT  141600.00000000003 193300.0 144100.00000000003 193900.00000000003 ;
      RECT  172900.0 191700.0 173500.0 192300.0 ;
      RECT  172900.0 194300.0 173500.0 194900.00000000003 ;
      RECT  168200.0 191700.0 173200.0 192300.0 ;
      RECT  172900.0 192000.0 173500.0 194600.00000000003 ;
      RECT  173200.0 194300.0 178200.0 194900.00000000003 ;
      RECT  141300.0 200500.0 141899.99999999997 201100.00000000003 ;
      RECT  141300.0 198899.99999999997 141899.99999999997 199500.0 ;
      RECT  139200.0 200500.0 141600.00000000003 201100.00000000003 ;
      RECT  141300.0 199200.0 141899.99999999997 200800.0 ;
      RECT  141600.00000000003 198899.99999999997 144100.00000000003 199500.0 ;
      RECT  172900.0 200500.0 173500.0 201100.00000000003 ;
      RECT  172900.0 197100.00000000003 173500.0 197700.0 ;
      RECT  168200.0 200500.0 173200.0 201100.00000000003 ;
      RECT  172900.0 197399.99999999997 173500.0 200800.0 ;
      RECT  173200.0 197100.00000000003 178200.0 197700.0 ;
      RECT  141300.0 210100.00000000003 141899.99999999997 210700.0 ;
      RECT  141300.0 211700.0 141899.99999999997 212300.0 ;
      RECT  139200.0 210100.00000000003 141600.00000000003 210700.0 ;
      RECT  141300.0 210399.99999999997 141899.99999999997 212000.0 ;
      RECT  141600.00000000003 211700.0 144100.00000000003 212300.0 ;
      RECT  172900.0 210100.00000000003 173500.0 210700.0 ;
      RECT  172900.0 212700.0 173500.0 213300.0 ;
      RECT  168200.0 210100.00000000003 173200.0 210700.0 ;
      RECT  172900.0 210399.99999999997 173500.0 213000.0 ;
      RECT  173200.0 212700.0 178200.0 213300.0 ;
      RECT  141300.0 218899.99999999997 141899.99999999997 219500.0 ;
      RECT  141300.0 217300.0 141899.99999999997 217900.00000000003 ;
      RECT  139200.0 218899.99999999997 141600.00000000003 219500.0 ;
      RECT  141300.0 217600.00000000003 141899.99999999997 219200.0 ;
      RECT  141600.00000000003 217300.0 144100.00000000003 217900.00000000003 ;
      RECT  172900.0 218899.99999999997 173500.0 219500.0 ;
      RECT  172900.0 215500.0 173500.0 216100.00000000003 ;
      RECT  168200.0 218899.99999999997 173200.0 219500.0 ;
      RECT  172900.0 215800.0 173500.0 219200.00000000006 ;
      RECT  173200.0 215500.0 178200.0 216100.00000000003 ;
      RECT  141300.0 228500.0 141899.99999999997 229100.00000000003 ;
      RECT  141300.0 230100.00000000003 141899.99999999997 230700.0 ;
      RECT  139200.0 228500.0 141600.00000000003 229100.00000000003 ;
      RECT  141300.0 228800.0 141899.99999999997 230400.00000000003 ;
      RECT  141600.00000000003 230100.00000000003 144100.00000000003 230700.0 ;
      RECT  172900.0 228500.0 173500.0 229100.00000000003 ;
      RECT  172900.0 231100.00000000003 173500.0 231700.0 ;
      RECT  168200.0 228500.0 173200.0 229100.00000000003 ;
      RECT  172900.0 228800.0 173500.0 231400.00000000003 ;
      RECT  173200.0 231100.00000000003 178200.0 231700.0 ;
      RECT  141300.0 237300.0 141899.99999999997 237900.00000000003 ;
      RECT  141300.0 235700.0 141899.99999999997 236300.0 ;
      RECT  139200.0 237300.0 141600.00000000003 237900.00000000003 ;
      RECT  141300.0 236000.0 141899.99999999997 237600.00000000003 ;
      RECT  141600.00000000003 235700.0 144100.00000000003 236300.0 ;
      RECT  172900.0 237300.0 173500.0 237900.00000000003 ;
      RECT  172900.0 233899.99999999997 173500.0 234500.0 ;
      RECT  168200.0 237300.0 173200.0 237900.00000000003 ;
      RECT  172900.0 234200.0 173500.0 237600.00000000003 ;
      RECT  173200.0 233899.99999999997 178200.0 234500.0 ;
      RECT  141300.0 246899.99999999997 141899.99999999997 247500.0 ;
      RECT  141300.0 248500.0 141899.99999999997 249100.00000000003 ;
      RECT  139200.0 246899.99999999997 141600.00000000003 247500.0 ;
      RECT  141300.0 247200.0 141899.99999999997 248800.0 ;
      RECT  141600.00000000003 248500.0 144100.00000000003 249100.00000000003 ;
      RECT  172900.0 246899.99999999997 173500.0 247500.0 ;
      RECT  172900.0 249500.0 173500.0 250100.00000000003 ;
      RECT  168200.0 246899.99999999997 173200.0 247500.0 ;
      RECT  172900.0 247200.0 173500.0 249800.0 ;
      RECT  173200.0 249500.0 178200.0 250100.00000000003 ;
      RECT  141300.0 255700.0 141899.99999999997 256300.0 ;
      RECT  141300.0 254100.00000000003 141899.99999999997 254700.00000000006 ;
      RECT  139200.0 255700.0 141600.00000000003 256300.0 ;
      RECT  141300.0 254399.99999999997 141899.99999999997 256000.0 ;
      RECT  141600.00000000003 254100.00000000003 144100.00000000003 254700.00000000006 ;
      RECT  172900.0 255700.0 173500.0 256300.0 ;
      RECT  172900.0 252300.0 173500.0 252900.00000000003 ;
      RECT  168200.0 255700.0 173200.0 256300.0 ;
      RECT  172900.0 252600.00000000003 173500.0 256000.00000000006 ;
      RECT  173200.0 252300.0 178200.0 252900.00000000003 ;
      RECT  141300.0 265300.0 141899.99999999997 265900.00000000006 ;
      RECT  141300.0 266900.0 141899.99999999997 267500.0 ;
      RECT  139200.0 265300.0 141600.00000000003 265900.00000000006 ;
      RECT  141300.0 265600.0 141899.99999999997 267200.00000000006 ;
      RECT  141600.00000000003 266900.0 144100.00000000003 267500.0 ;
      RECT  172900.0 265300.0 173500.0 265900.00000000006 ;
      RECT  172900.0 267900.0 173500.0 268500.0 ;
      RECT  168200.0 265300.0 173200.0 265900.00000000006 ;
      RECT  172900.0 265600.0 173500.0 268200.00000000006 ;
      RECT  173200.0 267900.0 178200.0 268500.0 ;
      RECT  174100.00000000003 108800.0 178600.00000000003 109399.99999999999 ;
      RECT  175500.0 29000.0 178600.00000000003 29600.0 ;
      RECT  176900.0 98600.00000000001 178600.00000000003 99200.0 ;
      RECT  146200.0 271100.0 172700.0 271700.00000000006 ;
      RECT  178600.00000000003 122400.0 185400.0 131600.00000000003 ;
      RECT  178600.00000000003 140800.0 185400.0 131600.00000000003 ;
      RECT  178600.00000000003 140800.0 185400.0 150000.0 ;
      RECT  178600.00000000003 159200.0 185400.0 150000.0 ;
      RECT  178600.00000000003 159200.0 185400.0 168400.00000000003 ;
      RECT  178600.00000000003 177600.00000000003 185400.0 168399.99999999997 ;
      RECT  178600.00000000003 177600.00000000003 185400.0 186800.0 ;
      RECT  178600.00000000003 196000.0 185400.0 186800.0 ;
      RECT  178600.00000000003 196000.0 185400.0 205200.0 ;
      RECT  178600.00000000003 214399.99999999997 185400.0 205200.0 ;
      RECT  178600.00000000003 214399.99999999997 185400.0 223600.00000000003 ;
      RECT  178600.00000000003 232800.0 185400.0 223600.00000000003 ;
      RECT  178600.00000000003 232800.0 185400.0 242000.0 ;
      RECT  178600.00000000003 251200.0 185400.0 242000.0 ;
      RECT  178600.00000000003 251200.0 185400.0 260399.99999999997 ;
      RECT  178600.00000000003 269600.0 185400.0 260400.00000000003 ;
      RECT  185400.0 122400.0 192200.0 131600.00000000003 ;
      RECT  185400.0 140800.0 192200.0 131600.00000000003 ;
      RECT  185400.0 140800.0 192200.0 150000.0 ;
      RECT  185400.0 159200.0 192200.0 150000.0 ;
      RECT  185400.0 159200.0 192200.0 168400.00000000003 ;
      RECT  185400.0 177600.00000000003 192200.0 168399.99999999997 ;
      RECT  185400.0 177600.00000000003 192200.0 186800.0 ;
      RECT  185400.0 196000.0 192200.0 186800.0 ;
      RECT  185400.0 196000.0 192200.0 205200.0 ;
      RECT  185400.0 214399.99999999997 192200.0 205200.0 ;
      RECT  185400.0 214399.99999999997 192200.0 223600.00000000003 ;
      RECT  185400.0 232800.0 192200.0 223600.00000000003 ;
      RECT  185400.0 232800.0 192200.0 242000.0 ;
      RECT  185400.0 251200.0 192200.0 242000.0 ;
      RECT  185400.0 251200.0 192200.0 260399.99999999997 ;
      RECT  185400.0 269600.0 192200.0 260400.00000000003 ;
      RECT  178200.0 123400.0 192400.0 124200.0 ;
      RECT  178200.0 139000.0 192400.0 139800.0 ;
      RECT  178200.0 141800.0 192400.0 142600.00000000003 ;
      RECT  178200.0 157399.99999999997 192400.0 158200.0 ;
      RECT  178200.0 160200.0 192400.0 161000.0 ;
      RECT  178200.0 175800.0 192400.0 176600.00000000003 ;
      RECT  178200.0 178600.00000000003 192400.0 179399.99999999997 ;
      RECT  178200.0 194200.0 192400.0 195000.0 ;
      RECT  178200.0 197000.0 192400.0 197800.0 ;
      RECT  178200.0 212600.00000000003 192400.0 213399.99999999997 ;
      RECT  178200.0 215399.99999999997 192400.0 216200.0 ;
      RECT  178200.0 231000.0 192400.0 231800.0 ;
      RECT  178200.0 233800.0 192400.0 234600.00000000003 ;
      RECT  178200.0 249399.99999999997 192400.0 250200.0 ;
      RECT  178200.0 252200.0 192400.0 253000.0 ;
      RECT  178200.0 267800.0 192400.0 268600.0 ;
      RECT  178600.00000000003 117900.0 185400.0 118500.00000000001 ;
      RECT  181500.0 112800.00000000001 182100.00000000003 118200.0 ;
      RECT  181800.0 107300.00000000001 183800.0 107900.0 ;
      RECT  183400.0 112100.00000000001 183800.0 112700.0 ;
      RECT  179800.0 107200.0 180600.00000000003 108000.00000000001 ;
      RECT  181400.0 107200.0 182200.0 108000.00000000001 ;
      RECT  181400.0 107200.0 182200.0 108000.00000000001 ;
      RECT  179800.0 107200.0 180600.00000000003 108000.00000000001 ;
      RECT  179800.0 112000.00000000001 180600.00000000003 112800.00000000001 ;
      RECT  181400.0 112000.00000000001 182200.0 112800.00000000001 ;
      RECT  181400.0 112000.00000000001 182200.0 112800.00000000001 ;
      RECT  179800.0 112000.00000000001 180600.00000000003 112800.00000000001 ;
      RECT  181400.0 112000.00000000001 182200.0 112800.00000000001 ;
      RECT  183000.0 112000.00000000001 183800.0 112800.00000000001 ;
      RECT  183000.0 112000.00000000001 183800.0 112800.00000000001 ;
      RECT  181400.0 112000.00000000001 182200.0 112800.00000000001 ;
      RECT  181200.0 108700.0 180400.0 109500.00000000001 ;
      RECT  181400.0 115600.00000000001 182200.0 116400.0 ;
      RECT  181400.0 112000.00000000001 182200.0 112800.00000000001 ;
      RECT  179800.0 112000.00000000001 180600.00000000003 112800.00000000001 ;
      RECT  179800.0 107200.0 180600.00000000003 108000.00000000001 ;
      RECT  183400.0 112000.00000000001 184200.0 112800.00000000001 ;
      RECT  183400.0 107200.0 184200.0 108000.00000000001 ;
      RECT  178600.00000000003 108800.00000000001 185400.0 109400.0 ;
      RECT  185400.0 117900.0 192200.0 118500.00000000001 ;
      RECT  188300.0 112800.00000000001 188900.0 118200.0 ;
      RECT  188600.00000000003 107300.00000000001 190600.00000000003 107900.0 ;
      RECT  190200.0 112100.00000000001 190600.00000000003 112700.0 ;
      RECT  186600.00000000003 107200.0 187400.0 108000.00000000001 ;
      RECT  188200.0 107200.0 189000.0 108000.00000000001 ;
      RECT  188200.0 107200.0 189000.0 108000.00000000001 ;
      RECT  186600.00000000003 107200.0 187400.0 108000.00000000001 ;
      RECT  186600.00000000003 112000.00000000001 187400.0 112800.00000000001 ;
      RECT  188200.0 112000.00000000001 189000.0 112800.00000000001 ;
      RECT  188200.0 112000.00000000001 189000.0 112800.00000000001 ;
      RECT  186600.00000000003 112000.00000000001 187400.0 112800.00000000001 ;
      RECT  188200.0 112000.00000000001 189000.0 112800.00000000001 ;
      RECT  189800.0 112000.00000000001 190600.00000000003 112800.00000000001 ;
      RECT  189800.0 112000.00000000001 190600.00000000003 112800.00000000001 ;
      RECT  188200.0 112000.00000000001 189000.0 112800.00000000001 ;
      RECT  188000.0 108700.0 187200.0 109500.00000000001 ;
      RECT  188200.0 115600.00000000001 189000.0 116400.0 ;
      RECT  188200.0 112000.00000000001 189000.0 112800.00000000001 ;
      RECT  186600.00000000003 112000.00000000001 187400.0 112800.00000000001 ;
      RECT  186600.00000000003 107200.0 187400.0 108000.00000000001 ;
      RECT  190200.0 112000.00000000001 191000.0 112800.00000000001 ;
      RECT  190200.0 107200.0 191000.0 108000.00000000001 ;
      RECT  185400.0 108800.00000000001 192200.0 109400.0 ;
      RECT  178600.00000000003 108800.00000000001 192200.0 109400.0 ;
      RECT  178600.00000000003 68800.00000000001 185400.0 101400.0 ;
      RECT  185400.0 68800.00000000001 192200.0 101400.0 ;
      RECT  178600.00000000003 98600.00000000001 192200.0 99200.0 ;
      RECT  178600.00000000003 24200.000000000004 185400.0 64599.99999999999 ;
      RECT  185400.0 24200.000000000004 192200.0 64599.99999999999 ;
      RECT  178600.00000000003 29000.000000000004 192200.0 29600.0 ;
      RECT  133600.0 127300.00000000001 134200.0 127900.0 ;
      RECT  133600.0 126900.0 134200.0 127500.00000000001 ;
      RECT  130900.0 127300.00000000001 133900.0 127900.0 ;
      RECT  133600.0 127200.0 134200.0 127600.00000000001 ;
      RECT  133900.0 126900.0 136900.0 127500.00000000001 ;
      RECT  133600.0 136100.00000000003 134200.0 136700.0 ;
      RECT  133600.0 136500.0 134200.0 137100.00000000003 ;
      RECT  130900.0 136100.00000000003 133900.0 136700.0 ;
      RECT  133600.0 136400.0 134200.0 136800.0 ;
      RECT  133900.0 136500.0 136900.0 137100.00000000003 ;
      RECT  133600.0 145700.0 134200.0 146300.0 ;
      RECT  133600.0 145300.0 134200.0 145900.0 ;
      RECT  130900.0 145700.0 133900.0 146300.0 ;
      RECT  133600.0 145600.00000000003 134200.0 146000.0 ;
      RECT  133900.0 145300.0 136900.0 145900.0 ;
      RECT  133600.0 154500.0 134200.0 155100.00000000003 ;
      RECT  133600.0 154899.99999999997 134200.0 155500.0 ;
      RECT  130900.0 154500.0 133900.0 155100.00000000003 ;
      RECT  133600.0 154800.0 134200.0 155200.0 ;
      RECT  133900.0 154899.99999999997 136900.0 155500.0 ;
      RECT  133600.0 164100.00000000003 134200.0 164700.0 ;
      RECT  133600.0 163700.0 134200.0 164300.0 ;
      RECT  130900.0 164100.00000000003 133900.0 164700.0 ;
      RECT  133600.0 164000.0 134200.0 164399.99999999997 ;
      RECT  133900.0 163700.0 136900.0 164300.0 ;
      RECT  133600.0 172899.99999999997 134200.0 173500.0 ;
      RECT  133600.0 173300.0 134200.0 173899.99999999997 ;
      RECT  130900.0 172899.99999999997 133900.0 173500.0 ;
      RECT  133600.0 173200.0 134200.0 173600.00000000003 ;
      RECT  133900.0 173300.0 136900.0 173899.99999999997 ;
      RECT  133600.0 182500.0 134200.0 183100.00000000003 ;
      RECT  133600.0 182100.00000000003 134200.0 182700.0 ;
      RECT  130900.0 182500.0 133900.0 183100.00000000003 ;
      RECT  133600.0 182399.99999999997 134200.0 182800.0 ;
      RECT  133900.0 182100.00000000003 136900.0 182700.0 ;
      RECT  133600.0 191300.0 134200.0 191899.99999999997 ;
      RECT  133600.0 191700.0 134200.0 192300.0 ;
      RECT  130900.0 191300.0 133900.0 191899.99999999997 ;
      RECT  133600.0 191600.00000000003 134200.0 192000.0 ;
      RECT  133900.0 191700.0 136900.0 192300.0 ;
      RECT  133600.0 200900.00000000003 134200.0 201500.0 ;
      RECT  133600.0 200500.0 134200.0 201100.00000000003 ;
      RECT  130900.0 200900.00000000003 133900.0 201500.0 ;
      RECT  133600.0 200800.0 134200.0 201200.0 ;
      RECT  133900.0 200500.0 136900.0 201100.00000000003 ;
      RECT  133600.0 209700.0 134200.0 210300.0 ;
      RECT  133600.0 210100.00000000003 134200.0 210700.0 ;
      RECT  130900.0 209700.0 133900.0 210300.0 ;
      RECT  133600.0 210000.0 134200.0 210400.00000000003 ;
      RECT  133900.0 210100.00000000003 136900.0 210700.0 ;
      RECT  133600.0 219300.0 134200.0 219899.99999999997 ;
      RECT  133600.0 218900.00000000003 134200.0 219500.0 ;
      RECT  130900.0 219300.0 133900.0 219899.99999999997 ;
      RECT  133600.0 219200.0 134200.0 219600.00000000003 ;
      RECT  133900.0 218900.00000000003 136900.0 219500.0 ;
      RECT  133600.0 228100.00000000003 134200.0 228700.0 ;
      RECT  133600.0 228500.0 134200.0 229100.00000000003 ;
      RECT  130900.0 228100.00000000003 133900.0 228700.0 ;
      RECT  133600.0 228400.00000000003 134200.0 228800.0 ;
      RECT  133900.0 228500.0 136900.0 229100.00000000003 ;
      RECT  133600.0 237700.0 134200.0 238300.0 ;
      RECT  133600.0 237300.0 134200.0 237899.99999999997 ;
      RECT  130900.0 237700.0 133900.0 238300.0 ;
      RECT  133600.0 237600.00000000003 134200.0 238000.0 ;
      RECT  133900.0 237300.0 136900.0 237899.99999999997 ;
      RECT  133600.0 246500.0 134200.0 247100.00000000003 ;
      RECT  133600.0 246900.00000000003 134200.0 247500.0 ;
      RECT  130900.0 246500.0 133900.0 247100.00000000003 ;
      RECT  133600.0 246800.0 134200.0 247200.0 ;
      RECT  133900.0 246900.00000000003 136900.0 247500.0 ;
      RECT  133600.0 256100.00000000003 134200.0 256700.0 ;
      RECT  133600.0 255700.0 134200.0 256300.0 ;
      RECT  130900.0 256100.00000000003 133900.0 256700.0 ;
      RECT  133600.0 256000.0 134200.0 256400.00000000003 ;
      RECT  133900.0 255700.0 136900.0 256300.0 ;
      RECT  133600.0 264900.0 134200.0 265500.0 ;
      RECT  133600.0 265300.0 134200.0 265900.0 ;
      RECT  130900.0 264900.0 133900.0 265500.0 ;
      RECT  133600.0 265200.0 134200.0 265600.0 ;
      RECT  133900.0 265300.0 136900.0 265900.0 ;
      RECT  115100.0 127300.00000000001 127300.00000000001 127900.0 ;
      RECT  120700.0 125900.0 129300.00000000001 126500.0 ;
      RECT  115100.0 136100.00000000003 127300.00000000001 136700.0 ;
      RECT  122100.0 137500.0 129300.00000000001 138100.00000000003 ;
      RECT  115100.0 145700.0 127300.00000000001 146300.0 ;
      RECT  123500.0 144300.0 129300.00000000001 144900.0 ;
      RECT  115100.0 154500.0 127300.00000000001 155100.00000000003 ;
      RECT  124900.0 155899.99999999997 129300.00000000001 156500.0 ;
      RECT  116500.0 164100.00000000003 127300.0 164700.0 ;
      RECT  120700.0 162700.0 129300.00000000001 163300.0 ;
      RECT  116500.0 172899.99999999997 127300.0 173500.0 ;
      RECT  122100.0 174300.0 129300.00000000001 174899.99999999997 ;
      RECT  116500.0 182500.0 127300.0 183100.00000000003 ;
      RECT  123500.0 181100.00000000003 129300.00000000001 181700.0 ;
      RECT  116500.0 191300.0 127300.0 191899.99999999997 ;
      RECT  124900.0 192700.0 129300.00000000001 193300.0 ;
      RECT  117900.0 200900.00000000003 127300.0 201500.0 ;
      RECT  120700.0 199500.0 129300.00000000001 200100.00000000003 ;
      RECT  117900.0 209700.0 127300.0 210300.0 ;
      RECT  122100.0 211100.00000000003 129300.00000000001 211700.0 ;
      RECT  117900.0 219300.0 127300.0 219899.99999999997 ;
      RECT  123500.0 217900.00000000003 129300.00000000001 218500.0 ;
      RECT  117900.0 228100.00000000003 127300.0 228700.0 ;
      RECT  124900.0 229500.0 129300.00000000001 230100.00000000003 ;
      RECT  119300.0 237700.0 127300.0 238300.0 ;
      RECT  120700.0 236300.0 129300.00000000001 236899.99999999997 ;
      RECT  119300.0 246500.0 127300.0 247100.00000000003 ;
      RECT  122100.0 247900.00000000003 129300.00000000001 248500.0 ;
      RECT  119300.0 256100.00000000003 127300.0 256700.0 ;
      RECT  123500.0 254700.0 129300.00000000001 255300.0 ;
      RECT  119300.0 264900.0 127300.0 265500.0 ;
      RECT  124900.0 266300.0 129300.00000000001 266900.0 ;
      RECT  125700.0 131700.0 141700.0 132300.0 ;
      RECT  125700.0 122500.0 141700.0 123100.00000000001 ;
      RECT  125700.0 150100.00000000003 141700.0 150700.0 ;
      RECT  125700.0 140900.0 141700.0 141500.0 ;
      RECT  125700.0 168500.0 141700.0 169100.00000000003 ;
      RECT  125700.0 159300.0 141700.0 159899.99999999997 ;
      RECT  125700.0 186900.00000000003 141700.0 187500.0 ;
      RECT  125700.0 177700.0 141700.0 178300.0 ;
      RECT  125700.0 205300.0 141700.0 205899.99999999997 ;
      RECT  125700.0 196100.00000000003 141700.0 196700.0 ;
      RECT  125700.0 223700.0 141700.0 224300.0 ;
      RECT  125700.0 214500.0 141700.0 215100.00000000003 ;
      RECT  125700.0 242100.00000000003 141700.0 242700.0 ;
      RECT  125700.0 232900.00000000003 141700.0 233500.0 ;
      RECT  125700.0 260500.0 141700.0 261100.00000000003 ;
      RECT  125700.0 251300.0 141700.0 251899.99999999997 ;
      RECT  90400.0 126900.0 91000.0 127500.00000000001 ;
      RECT  90400.0 129900.0 91000.0 130500.0 ;
      RECT  87600.0 126900.0 90700.0 127500.00000000001 ;
      RECT  90400.0 127200.0 91000.0 130199.99999999999 ;
      RECT  90700.0 129900.0 93200.0 130500.0 ;
      RECT  81500.0 126900.0 85300.0 127500.00000000001 ;
      RECT  90400.0 136500.0 91000.0 137100.00000000003 ;
      RECT  90400.0 139100.00000000003 91000.0 139700.0 ;
      RECT  87600.0 136500.0 90700.0 137100.00000000003 ;
      RECT  90400.0 136800.0 91000.0 139400.0 ;
      RECT  90700.0 139100.00000000003 94600.0 139700.0 ;
      RECT  82900.0 136500.0 85300.0 137100.00000000003 ;
      RECT  81500.0 142300.0 96000.0 142900.0 ;
      RECT  82900.0 151500.0 97400.0 152100.00000000003 ;
      RECT  93200.0 127300.00000000001 100100.0 127900.0 ;
      RECT  94600.0 125900.0 102100.0 126500.0 ;
      RECT  96000.0 136100.00000000003 100100.0 136700.0 ;
      RECT  94600.0 137500.0 102100.0 138100.00000000003 ;
      RECT  93200.0 145700.0 100100.0 146300.0 ;
      RECT  97400.0 144300.0 102100.0 144900.0 ;
      RECT  96000.0 154500.0 100100.0 155100.00000000003 ;
      RECT  97400.0 155899.99999999997 102100.0 156500.0 ;
      RECT  106400.0 127300.00000000001 107000.0 127900.0 ;
      RECT  106400.0 126900.0 107000.0 127500.00000000001 ;
      RECT  103700.0 127300.00000000001 106700.0 127900.0 ;
      RECT  106400.0 127200.0 107000.0 127600.00000000001 ;
      RECT  106700.0 126900.0 109700.0 127500.00000000001 ;
      RECT  106400.0 136100.00000000003 107000.0 136700.0 ;
      RECT  106400.0 136500.0 107000.0 137100.00000000003 ;
      RECT  103700.0 136100.00000000003 106700.0 136700.0 ;
      RECT  106400.0 136400.0 107000.0 136800.0 ;
      RECT  106700.0 136500.0 109700.0 137100.00000000003 ;
      RECT  106400.0 145700.0 107000.0 146300.0 ;
      RECT  106400.0 145300.0 107000.0 145900.0 ;
      RECT  103700.0 145700.0 106700.0 146300.0 ;
      RECT  106400.0 145600.00000000003 107000.0 146000.0 ;
      RECT  106700.0 145300.0 109700.0 145900.0 ;
      RECT  106400.0 154500.0 107000.0 155100.00000000003 ;
      RECT  106400.0 154899.99999999997 107000.0 155500.0 ;
      RECT  103700.0 154500.0 106700.0 155100.00000000003 ;
      RECT  106400.0 154800.0 107000.0 155200.0 ;
      RECT  106700.0 154899.99999999997 109700.0 155500.0 ;
      RECT  80900.0 131700.0 114500.0 132300.0 ;
      RECT  80900.0 122500.0 114500.0 123100.00000000001 ;
      RECT  80900.0 131700.0 114500.0 132300.0 ;
      RECT  80900.0 140900.0 114500.0 141500.0 ;
      RECT  80900.0 150100.00000000003 114500.0 150700.0 ;
      RECT  80900.0 140900.0 114500.0 141500.0 ;
      RECT  80900.0 150100.00000000003 114500.0 150700.0 ;
      RECT  80900.0 159300.0 114500.0 159899.99999999997 ;
      RECT  88100.0 130699.99999999999 88900.0 132000.0 ;
      RECT  88100.0 122800.00000000001 88900.0 124100.00000000001 ;
      RECT  84900.0 123700.0 85700.0 122500.0 ;
      RECT  84900.0 129900.0 85700.0 132300.0 ;
      RECT  86700.0 123700.0 87300.0 129900.0 ;
      RECT  84900.0 129900.0 85700.0 130699.99999999999 ;
      RECT  86500.0 129900.0 87300.0 130699.99999999999 ;
      RECT  86500.0 129900.0 87300.0 130699.99999999999 ;
      RECT  84900.0 129900.0 85700.0 130699.99999999999 ;
      RECT  84900.0 123700.0 85700.0 124500.0 ;
      RECT  86500.0 123700.0 87300.0 124500.0 ;
      RECT  86500.0 123700.0 87300.0 124500.0 ;
      RECT  84900.0 123700.0 85700.0 124500.0 ;
      RECT  88100.0 130300.00000000001 88900.0 131100.00000000003 ;
      RECT  88100.0 123700.0 88900.0 124500.0 ;
      RECT  85300.0 126800.00000000001 86100.0 127600.00000000001 ;
      RECT  85300.0 126800.00000000001 86100.0 127600.00000000001 ;
      RECT  87000.0 126900.0 87600.0 127500.0 ;
      RECT  83700.0 131700.0 90100.0 132300.0 ;
      RECT  83700.0 122500.0 90100.0 123100.00000000001 ;
      RECT  88100.0 133300.0 88900.0 132000.0 ;
      RECT  88100.0 141200.0 88900.0 139900.0 ;
      RECT  84900.0 140300.0 85700.0 141500.0 ;
      RECT  84900.0 134100.00000000003 85700.0 131700.0 ;
      RECT  86700.0 140300.0 87300.0 134100.00000000003 ;
      RECT  84900.0 134100.00000000003 85700.0 133300.0 ;
      RECT  86500.0 134100.00000000003 87300.0 133300.0 ;
      RECT  86500.0 134100.00000000003 87300.0 133300.0 ;
      RECT  84900.0 134100.00000000003 85700.0 133300.0 ;
      RECT  84900.0 140300.0 85700.0 139500.0 ;
      RECT  86500.0 140300.0 87300.0 139500.0 ;
      RECT  86500.0 140300.0 87300.0 139500.0 ;
      RECT  84900.0 140300.0 85700.0 139500.0 ;
      RECT  88100.0 133700.0 88900.0 132900.0 ;
      RECT  88100.0 140300.0 88900.0 139500.0 ;
      RECT  85300.0 137200.0 86100.0 136400.0 ;
      RECT  85300.0 137200.0 86100.0 136400.0 ;
      RECT  87000.0 137100.00000000003 87600.0 136500.0 ;
      RECT  83700.0 132300.0 90100.0 131700.0 ;
      RECT  83700.0 141500.0 90100.0 140900.0 ;
      RECT  112500.0 130699.99999999999 113300.00000000001 132000.0 ;
      RECT  112500.0 122800.00000000001 113300.00000000001 124100.00000000001 ;
      RECT  109300.0 123700.0 110100.0 122500.0 ;
      RECT  109300.0 129900.0 110100.0 132300.0 ;
      RECT  111100.0 123700.0 111700.0 129900.0 ;
      RECT  109300.0 129900.0 110100.0 130699.99999999999 ;
      RECT  110900.0 129900.0 111700.0 130699.99999999999 ;
      RECT  110900.0 129900.0 111700.0 130699.99999999999 ;
      RECT  109300.0 129900.0 110100.0 130699.99999999999 ;
      RECT  109300.0 123700.0 110100.0 124500.0 ;
      RECT  110900.0 123700.0 111700.0 124500.0 ;
      RECT  110900.0 123700.0 111700.0 124500.0 ;
      RECT  109300.0 123700.0 110100.0 124500.0 ;
      RECT  112500.0 130300.00000000001 113300.00000000001 131100.00000000003 ;
      RECT  112500.0 123700.0 113300.00000000001 124500.0 ;
      RECT  109700.0 126800.00000000001 110500.0 127600.00000000001 ;
      RECT  109700.0 126800.00000000001 110500.0 127600.00000000001 ;
      RECT  111400.0 126900.0 112000.0 127500.0 ;
      RECT  108100.0 131700.0 114500.0 132300.0 ;
      RECT  108100.0 122500.0 114500.0 123100.00000000001 ;
      RECT  112500.0 133300.0 113300.00000000001 132000.0 ;
      RECT  112500.0 141200.0 113300.00000000001 139900.0 ;
      RECT  109300.0 140300.0 110100.0 141500.0 ;
      RECT  109300.0 134100.00000000003 110100.0 131700.0 ;
      RECT  111100.0 140300.0 111700.0 134100.00000000003 ;
      RECT  109300.0 134100.00000000003 110100.0 133300.0 ;
      RECT  110900.0 134100.00000000003 111700.0 133300.0 ;
      RECT  110900.0 134100.00000000003 111700.0 133300.0 ;
      RECT  109300.0 134100.00000000003 110100.0 133300.0 ;
      RECT  109300.0 140300.0 110100.0 139500.0 ;
      RECT  110900.0 140300.0 111700.0 139500.0 ;
      RECT  110900.0 140300.0 111700.0 139500.0 ;
      RECT  109300.0 140300.0 110100.0 139500.0 ;
      RECT  112500.0 133700.0 113300.00000000001 132900.0 ;
      RECT  112500.0 140300.0 113300.00000000001 139500.0 ;
      RECT  109700.0 137200.0 110500.0 136400.0 ;
      RECT  109700.0 137200.0 110500.0 136400.0 ;
      RECT  111400.0 137100.00000000003 112000.0 136500.0 ;
      RECT  108100.0 132300.0 114500.0 131700.0 ;
      RECT  108100.0 141500.0 114500.0 140900.0 ;
      RECT  112500.0 149100.00000000003 113300.00000000001 150400.0 ;
      RECT  112500.0 141200.0 113300.00000000001 142500.0 ;
      RECT  109300.0 142100.00000000003 110100.0 140900.0 ;
      RECT  109300.0 148300.0 110100.0 150700.0 ;
      RECT  111100.0 142100.00000000003 111700.0 148300.0 ;
      RECT  109300.0 148300.0 110100.0 149100.00000000003 ;
      RECT  110900.0 148300.0 111700.0 149100.00000000003 ;
      RECT  110900.0 148300.0 111700.0 149100.00000000003 ;
      RECT  109300.0 148300.0 110100.0 149100.00000000003 ;
      RECT  109300.0 142100.00000000003 110100.0 142900.0 ;
      RECT  110900.0 142100.00000000003 111700.0 142900.0 ;
      RECT  110900.0 142100.00000000003 111700.0 142900.0 ;
      RECT  109300.0 142100.00000000003 110100.0 142900.0 ;
      RECT  112500.0 148700.0 113300.00000000001 149500.0 ;
      RECT  112500.0 142100.00000000003 113300.00000000001 142900.0 ;
      RECT  109700.0 145200.0 110500.0 146000.0 ;
      RECT  109700.0 145200.0 110500.0 146000.0 ;
      RECT  111400.0 145300.0 112000.0 145900.0 ;
      RECT  108100.0 150100.00000000003 114500.0 150700.0 ;
      RECT  108100.0 140900.0 114500.0 141500.0 ;
      RECT  112500.0 151700.0 113300.00000000001 150400.0 ;
      RECT  112500.0 159600.00000000003 113300.00000000001 158300.0 ;
      RECT  109300.0 158700.0 110100.0 159899.99999999997 ;
      RECT  109300.0 152500.0 110100.0 150100.00000000003 ;
      RECT  111100.0 158700.0 111700.0 152500.0 ;
      RECT  109300.0 152500.0 110100.0 151700.0 ;
      RECT  110900.0 152500.0 111700.0 151700.0 ;
      RECT  110900.0 152500.0 111700.0 151700.0 ;
      RECT  109300.0 152500.0 110100.0 151700.0 ;
      RECT  109300.0 158700.0 110100.0 157899.99999999997 ;
      RECT  110900.0 158700.0 111700.0 157899.99999999997 ;
      RECT  110900.0 158700.0 111700.0 157899.99999999997 ;
      RECT  109300.0 158700.0 110100.0 157899.99999999997 ;
      RECT  112500.0 152100.00000000003 113300.00000000001 151300.0 ;
      RECT  112500.0 158700.0 113300.00000000001 157899.99999999997 ;
      RECT  109700.0 155600.00000000003 110500.0 154800.0 ;
      RECT  109700.0 155600.00000000003 110500.0 154800.0 ;
      RECT  111400.0 155500.0 112000.0 154899.99999999997 ;
      RECT  108100.0 150700.0 114500.0 150100.00000000003 ;
      RECT  108100.0 159899.99999999997 114500.0 159300.0 ;
      RECT  99700.0 124100.00000000001 100500.0 122500.0 ;
      RECT  99700.0 129900.0 100500.0 132300.0 ;
      RECT  102900.0 129900.0 103700.0 132300.0 ;
      RECT  104500.0 130699.99999999999 105300.0 132000.0 ;
      RECT  104500.0 122800.00000000001 105300.0 124100.00000000001 ;
      RECT  99700.0 129900.0 100500.0 130699.99999999999 ;
      RECT  101300.0 129900.0 102100.0 130699.99999999999 ;
      RECT  101300.0 129900.0 102100.0 130699.99999999999 ;
      RECT  99700.0 129900.0 100500.0 130699.99999999999 ;
      RECT  101300.0 129900.0 102100.0 130699.99999999999 ;
      RECT  102900.0 129900.0 103700.0 130699.99999999999 ;
      RECT  102900.0 129900.0 103700.0 130699.99999999999 ;
      RECT  101300.0 129900.0 102100.0 130699.99999999999 ;
      RECT  99700.0 124100.00000000001 100500.0 124900.0 ;
      RECT  101300.0 124100.00000000001 102100.0 124900.0 ;
      RECT  101300.0 124100.00000000001 102100.0 124900.0 ;
      RECT  99700.0 124100.00000000001 100500.0 124900.0 ;
      RECT  101300.0 124100.00000000001 102100.0 124900.0 ;
      RECT  102900.0 124100.00000000001 103700.0 124900.0 ;
      RECT  102900.0 124100.00000000001 103700.0 124900.0 ;
      RECT  101300.0 124100.00000000001 102100.0 124900.0 ;
      RECT  104500.0 130300.00000000001 105300.0 131100.00000000003 ;
      RECT  104500.0 123700.0 105300.0 124500.0 ;
      RECT  102900.0 125800.00000000001 102100.0 126600.00000000001 ;
      RECT  100900.0 127200.0 100100.0 128000.0 ;
      RECT  101300.0 129900.0 102100.0 130699.99999999999 ;
      RECT  102900.0 124100.00000000001 103700.0 124900.0 ;
      RECT  103700.0 127200.0 102900.0 128000.0 ;
      RECT  100100.0 127200.0 100900.0 128000.0 ;
      RECT  102100.0 125800.00000000001 102900.0 126600.00000000001 ;
      RECT  102900.0 127200.0 103700.0 128000.0 ;
      RECT  98500.0 131700.0 108100.0 132300.0 ;
      RECT  98500.0 122500.0 108100.0 123100.00000000001 ;
      RECT  99700.0 139900.0 100500.0 141500.0 ;
      RECT  99700.0 134100.00000000003 100500.0 131700.0 ;
      RECT  102900.0 134100.00000000003 103700.0 131700.0 ;
      RECT  104500.0 133300.0 105300.0 132000.0 ;
      RECT  104500.0 141200.0 105300.0 139900.0 ;
      RECT  99700.0 134100.00000000003 100500.0 133300.0 ;
      RECT  101300.0 134100.00000000003 102100.0 133300.0 ;
      RECT  101300.0 134100.00000000003 102100.0 133300.0 ;
      RECT  99700.0 134100.00000000003 100500.0 133300.0 ;
      RECT  101300.0 134100.00000000003 102100.0 133300.0 ;
      RECT  102900.0 134100.00000000003 103700.0 133300.0 ;
      RECT  102900.0 134100.00000000003 103700.0 133300.0 ;
      RECT  101300.0 134100.00000000003 102100.0 133300.0 ;
      RECT  99700.0 139900.0 100500.0 139100.00000000003 ;
      RECT  101300.0 139900.0 102100.0 139100.00000000003 ;
      RECT  101300.0 139900.0 102100.0 139100.00000000003 ;
      RECT  99700.0 139900.0 100500.0 139100.00000000003 ;
      RECT  101300.0 139900.0 102100.0 139100.00000000003 ;
      RECT  102900.0 139900.0 103700.0 139100.00000000003 ;
      RECT  102900.0 139900.0 103700.0 139100.00000000003 ;
      RECT  101300.0 139900.0 102100.0 139100.00000000003 ;
      RECT  104500.0 133700.0 105300.0 132900.0 ;
      RECT  104500.0 140300.0 105300.0 139500.0 ;
      RECT  102900.0 138200.0 102100.0 137400.0 ;
      RECT  100900.0 136800.0 100100.0 136000.0 ;
      RECT  101300.0 134100.00000000003 102100.0 133300.0 ;
      RECT  102900.0 139900.0 103700.0 139100.00000000003 ;
      RECT  103700.0 136800.0 102900.0 136000.0 ;
      RECT  100100.0 136800.0 100900.0 136000.0 ;
      RECT  102100.0 138200.0 102900.0 137400.0 ;
      RECT  102900.0 136800.0 103700.0 136000.0 ;
      RECT  98500.0 132300.0 108100.0 131700.0 ;
      RECT  98500.0 141500.0 108100.0 140900.0 ;
      RECT  99700.0 142500.0 100500.0 140900.0 ;
      RECT  99700.0 148300.0 100500.0 150700.0 ;
      RECT  102900.0 148300.0 103700.0 150700.0 ;
      RECT  104500.0 149100.00000000003 105300.0 150400.0 ;
      RECT  104500.0 141200.0 105300.0 142500.0 ;
      RECT  99700.0 148300.0 100500.0 149100.00000000003 ;
      RECT  101300.0 148300.0 102100.0 149100.00000000003 ;
      RECT  101300.0 148300.0 102100.0 149100.00000000003 ;
      RECT  99700.0 148300.0 100500.0 149100.00000000003 ;
      RECT  101300.0 148300.0 102100.0 149100.00000000003 ;
      RECT  102900.0 148300.0 103700.0 149100.00000000003 ;
      RECT  102900.0 148300.0 103700.0 149100.00000000003 ;
      RECT  101300.0 148300.0 102100.0 149100.00000000003 ;
      RECT  99700.0 142500.0 100500.0 143300.0 ;
      RECT  101300.0 142500.0 102100.0 143300.0 ;
      RECT  101300.0 142500.0 102100.0 143300.0 ;
      RECT  99700.0 142500.0 100500.0 143300.0 ;
      RECT  101300.0 142500.0 102100.0 143300.0 ;
      RECT  102900.0 142500.0 103700.0 143300.0 ;
      RECT  102900.0 142500.0 103700.0 143300.0 ;
      RECT  101300.0 142500.0 102100.0 143300.0 ;
      RECT  104500.0 148700.0 105300.0 149500.0 ;
      RECT  104500.0 142100.00000000003 105300.0 142900.0 ;
      RECT  102900.0 144200.0 102100.0 145000.0 ;
      RECT  100900.0 145600.00000000003 100100.0 146400.0 ;
      RECT  101300.0 148300.0 102100.0 149100.00000000003 ;
      RECT  102900.0 142500.0 103700.0 143300.0 ;
      RECT  103700.0 145600.00000000003 102900.0 146400.0 ;
      RECT  100100.0 145600.00000000003 100900.0 146400.0 ;
      RECT  102100.0 144200.0 102900.0 145000.0 ;
      RECT  102900.0 145600.00000000003 103700.0 146400.0 ;
      RECT  98500.0 150100.00000000003 108100.0 150700.0 ;
      RECT  98500.0 140900.0 108100.0 141500.0 ;
      RECT  99700.0 158300.0 100500.0 159899.99999999997 ;
      RECT  99700.0 152500.0 100500.0 150100.00000000003 ;
      RECT  102900.0 152500.0 103700.0 150100.00000000003 ;
      RECT  104500.0 151700.0 105300.0 150400.0 ;
      RECT  104500.0 159600.00000000003 105300.0 158300.0 ;
      RECT  99700.0 152500.0 100500.0 151700.0 ;
      RECT  101300.0 152500.0 102100.0 151700.0 ;
      RECT  101300.0 152500.0 102100.0 151700.0 ;
      RECT  99700.0 152500.0 100500.0 151700.0 ;
      RECT  101300.0 152500.0 102100.0 151700.0 ;
      RECT  102900.0 152500.0 103700.0 151700.0 ;
      RECT  102900.0 152500.0 103700.0 151700.0 ;
      RECT  101300.0 152500.0 102100.0 151700.0 ;
      RECT  99700.0 158300.0 100500.0 157500.0 ;
      RECT  101300.0 158300.0 102100.0 157500.0 ;
      RECT  101300.0 158300.0 102100.0 157500.0 ;
      RECT  99700.0 158300.0 100500.0 157500.0 ;
      RECT  101300.0 158300.0 102100.0 157500.0 ;
      RECT  102900.0 158300.0 103700.0 157500.0 ;
      RECT  102900.0 158300.0 103700.0 157500.0 ;
      RECT  101300.0 158300.0 102100.0 157500.0 ;
      RECT  104500.0 152100.00000000003 105300.0 151300.0 ;
      RECT  104500.0 158700.0 105300.0 157899.99999999997 ;
      RECT  102900.0 156600.00000000003 102100.0 155800.0 ;
      RECT  100900.0 155200.0 100100.0 154400.00000000003 ;
      RECT  101300.0 152500.0 102100.0 151700.0 ;
      RECT  102900.0 158300.0 103700.0 157500.0 ;
      RECT  103700.0 155200.0 102900.0 154400.00000000003 ;
      RECT  100100.0 155200.0 100900.0 154400.00000000003 ;
      RECT  102100.0 156600.00000000003 102900.0 155800.0 ;
      RECT  102900.0 155200.0 103700.0 154400.00000000003 ;
      RECT  98500.0 150700.0 108100.0 150100.00000000003 ;
      RECT  98500.0 159899.99999999997 108100.0 159300.0 ;
      RECT  93600.0 129800.00000000001 92800.0 130600.00000000003 ;
      RECT  81900.0 126800.00000000001 81100.0 127600.00000000001 ;
      RECT  95000.0 139000.0 94200.0 139800.0 ;
      RECT  83300.0 136400.0 82500.0 137200.0 ;
      RECT  81900.0 142200.0 81100.0 143000.0 ;
      RECT  96400.0 142200.0 95600.0 143000.0 ;
      RECT  83300.0 151400.0 82500.0 152200.0 ;
      RECT  97800.0 151400.0 97000.0 152200.0 ;
      RECT  93600.0 127200.0 92800.0 128000.0 ;
      RECT  95000.0 125800.00000000001 94200.0 126600.00000000001 ;
      RECT  96400.0 136000.0 95600.0 136800.0 ;
      RECT  95000.0 137400.0 94200.0 138200.0 ;
      RECT  93600.0 145600.00000000003 92800.0 146400.0 ;
      RECT  97800.0 144200.0 97000.0 145000.0 ;
      RECT  96400.0 154399.99999999997 95600.0 155200.0 ;
      RECT  97800.0 155800.0 97000.0 156600.00000000003 ;
      RECT  90500.0 131600.00000000003 89700.0 132400.0 ;
      RECT  108500.0 131600.00000000003 107700.0 132400.0 ;
      RECT  90500.0 122400.0 89700.0 123200.0 ;
      RECT  108500.0 122400.0 107700.0 123200.0 ;
      RECT  90500.0 131600.00000000003 89700.0 132400.0 ;
      RECT  108500.0 131600.00000000003 107700.0 132400.0 ;
      RECT  90500.0 140800.0 89700.0 141600.00000000003 ;
      RECT  108500.0 140800.0 107700.0 141600.00000000003 ;
      RECT  90500.0 150000.0 89700.0 150800.0 ;
      RECT  108500.0 150000.0 107700.0 150800.0 ;
      RECT  90500.0 140800.0 89700.0 141600.00000000003 ;
      RECT  108500.0 140800.0 107700.0 141600.00000000003 ;
      RECT  90500.0 150000.0 89700.0 150800.0 ;
      RECT  108500.0 150000.0 107700.0 150800.0 ;
      RECT  90500.0 159200.0 89700.0 160000.0 ;
      RECT  108500.0 159200.0 107700.0 160000.0 ;
      RECT  111400.0 126900.0 112000.0 127500.0 ;
      RECT  111400.0 136500.0 112000.0 137100.00000000003 ;
      RECT  111400.0 145300.0 112000.0 145900.0 ;
      RECT  111400.0 154899.99999999997 112000.0 155500.0 ;
      RECT  90400.0 163700.0 91000.0 164300.0 ;
      RECT  90400.0 166700.0 91000.0 167300.0 ;
      RECT  87600.0 163700.0 90700.0 164300.0 ;
      RECT  90400.0 164000.0 91000.0 167000.0 ;
      RECT  90700.0 166700.0 93200.0 167300.0 ;
      RECT  81500.0 163700.0 85300.0 164300.0 ;
      RECT  90400.0 173300.0 91000.0 173899.99999999997 ;
      RECT  90400.0 175899.99999999997 91000.0 176500.0 ;
      RECT  87600.0 173300.0 90700.0 173899.99999999997 ;
      RECT  90400.0 173600.00000000003 91000.0 176200.0 ;
      RECT  90700.0 175899.99999999997 94600.0 176500.0 ;
      RECT  82900.0 173300.0 85300.0 173899.99999999997 ;
      RECT  81500.0 179100.00000000003 96000.0 179700.0 ;
      RECT  82900.0 188300.0 97400.0 188899.99999999997 ;
      RECT  93200.0 164100.00000000003 100100.0 164700.0 ;
      RECT  94600.0 162700.0 102100.0 163300.0 ;
      RECT  96000.0 172899.99999999997 100100.0 173500.0 ;
      RECT  94600.0 174300.0 102100.0 174899.99999999997 ;
      RECT  93200.0 182500.0 100100.0 183100.00000000003 ;
      RECT  97400.0 181100.00000000003 102100.0 181700.0 ;
      RECT  96000.0 191300.0 100100.0 191899.99999999997 ;
      RECT  97400.0 192700.0 102100.0 193300.0 ;
      RECT  106400.0 164100.00000000003 107000.0 164700.0 ;
      RECT  106400.0 163700.0 107000.0 164300.0 ;
      RECT  103700.0 164100.00000000003 106700.0 164700.0 ;
      RECT  106400.0 164000.0 107000.0 164399.99999999997 ;
      RECT  106700.0 163700.0 109700.0 164300.0 ;
      RECT  106400.0 172899.99999999997 107000.0 173500.0 ;
      RECT  106400.0 173300.0 107000.0 173899.99999999997 ;
      RECT  103700.0 172899.99999999997 106700.0 173500.0 ;
      RECT  106400.0 173200.0 107000.0 173600.00000000003 ;
      RECT  106700.0 173300.0 109700.0 173899.99999999997 ;
      RECT  106400.0 182500.0 107000.0 183100.00000000003 ;
      RECT  106400.0 182100.00000000003 107000.0 182700.0 ;
      RECT  103700.0 182500.0 106700.0 183100.00000000003 ;
      RECT  106400.0 182399.99999999997 107000.0 182800.0 ;
      RECT  106700.0 182100.00000000003 109700.0 182700.0 ;
      RECT  106400.0 191300.0 107000.0 191899.99999999997 ;
      RECT  106400.0 191700.0 107000.0 192300.0 ;
      RECT  103700.0 191300.0 106700.0 191899.99999999997 ;
      RECT  106400.0 191600.00000000003 107000.0 192000.0 ;
      RECT  106700.0 191700.0 109700.0 192300.0 ;
      RECT  80900.0 168500.0 114500.0 169100.00000000003 ;
      RECT  80900.0 159300.0 114500.0 159899.99999999997 ;
      RECT  80900.0 168500.0 114500.0 169100.00000000003 ;
      RECT  80900.0 177700.0 114500.0 178300.0 ;
      RECT  80900.0 186899.99999999997 114500.0 187500.0 ;
      RECT  80900.0 177700.0 114500.0 178300.0 ;
      RECT  80900.0 186899.99999999997 114500.0 187500.0 ;
      RECT  80900.0 196100.00000000003 114500.0 196700.0 ;
      RECT  88100.0 167500.0 88900.0 168800.0 ;
      RECT  88100.0 159600.00000000003 88900.0 160899.99999999997 ;
      RECT  84900.0 160500.0 85700.0 159300.0 ;
      RECT  84900.0 166700.0 85700.0 169100.00000000003 ;
      RECT  86700.0 160500.0 87300.0 166700.0 ;
      RECT  84900.0 166700.0 85700.0 167500.0 ;
      RECT  86500.0 166700.0 87300.0 167500.0 ;
      RECT  86500.0 166700.0 87300.0 167500.0 ;
      RECT  84900.0 166700.0 85700.0 167500.0 ;
      RECT  84900.0 160500.0 85700.0 161300.0 ;
      RECT  86500.0 160500.0 87300.0 161300.0 ;
      RECT  86500.0 160500.0 87300.0 161300.0 ;
      RECT  84900.0 160500.0 85700.0 161300.0 ;
      RECT  88100.0 167100.00000000003 88900.0 167899.99999999997 ;
      RECT  88100.0 160500.0 88900.0 161300.0 ;
      RECT  85300.0 163600.00000000003 86100.0 164399.99999999997 ;
      RECT  85300.0 163600.00000000003 86100.0 164399.99999999997 ;
      RECT  87000.0 163700.0 87600.0 164300.0 ;
      RECT  83700.0 168500.0 90100.0 169100.00000000003 ;
      RECT  83700.0 159300.0 90100.0 159899.99999999997 ;
      RECT  88100.0 170100.00000000003 88900.0 168800.0 ;
      RECT  88100.0 178000.0 88900.0 176700.0 ;
      RECT  84900.0 177100.00000000003 85700.0 178300.0 ;
      RECT  84900.0 170899.99999999997 85700.0 168500.0 ;
      RECT  86700.0 177100.00000000003 87300.0 170899.99999999997 ;
      RECT  84900.0 170900.00000000003 85700.0 170100.00000000003 ;
      RECT  86500.0 170900.00000000003 87300.0 170100.00000000003 ;
      RECT  86500.0 170900.00000000003 87300.0 170100.00000000003 ;
      RECT  84900.0 170900.00000000003 85700.0 170100.00000000003 ;
      RECT  84900.0 177100.00000000003 85700.0 176300.0 ;
      RECT  86500.0 177100.00000000003 87300.0 176300.0 ;
      RECT  86500.0 177100.00000000003 87300.0 176300.0 ;
      RECT  84900.0 177100.00000000003 85700.0 176300.0 ;
      RECT  88100.0 170500.0 88900.0 169700.0 ;
      RECT  88100.0 177100.00000000003 88900.0 176300.0 ;
      RECT  85300.0 174000.0 86100.0 173200.0 ;
      RECT  85300.0 174000.0 86100.0 173200.0 ;
      RECT  87000.0 173899.99999999997 87600.0 173300.0 ;
      RECT  83700.0 169100.00000000003 90100.0 168500.0 ;
      RECT  83700.0 178300.0 90100.0 177700.0 ;
      RECT  112500.0 167500.0 113300.00000000001 168800.0 ;
      RECT  112500.0 159600.00000000003 113300.00000000001 160899.99999999997 ;
      RECT  109300.0 160500.0 110100.0 159300.0 ;
      RECT  109300.0 166700.0 110100.0 169100.00000000003 ;
      RECT  111100.0 160500.0 111700.0 166700.0 ;
      RECT  109300.0 166700.0 110100.0 167500.0 ;
      RECT  110900.0 166700.0 111700.0 167500.0 ;
      RECT  110900.0 166700.0 111700.0 167500.0 ;
      RECT  109300.0 166700.0 110100.0 167500.0 ;
      RECT  109300.0 160500.0 110100.0 161300.0 ;
      RECT  110900.0 160500.0 111700.0 161300.0 ;
      RECT  110900.0 160500.0 111700.0 161300.0 ;
      RECT  109300.0 160500.0 110100.0 161300.0 ;
      RECT  112500.0 167100.00000000003 113300.00000000001 167899.99999999997 ;
      RECT  112500.0 160500.0 113300.00000000001 161300.0 ;
      RECT  109700.0 163600.00000000003 110500.0 164399.99999999997 ;
      RECT  109700.0 163600.00000000003 110500.0 164399.99999999997 ;
      RECT  111400.0 163700.0 112000.0 164300.0 ;
      RECT  108100.0 168500.0 114500.0 169100.00000000003 ;
      RECT  108100.0 159300.0 114500.0 159899.99999999997 ;
      RECT  112500.0 170100.00000000003 113300.00000000001 168800.0 ;
      RECT  112500.0 178000.0 113300.00000000001 176700.0 ;
      RECT  109300.0 177100.00000000003 110100.0 178300.0 ;
      RECT  109300.0 170899.99999999997 110100.0 168500.0 ;
      RECT  111100.0 177100.00000000003 111700.0 170899.99999999997 ;
      RECT  109300.0 170900.00000000003 110100.0 170100.00000000003 ;
      RECT  110900.0 170900.00000000003 111700.0 170100.00000000003 ;
      RECT  110900.0 170900.00000000003 111700.0 170100.00000000003 ;
      RECT  109300.0 170900.00000000003 110100.0 170100.00000000003 ;
      RECT  109300.0 177100.00000000003 110100.0 176300.0 ;
      RECT  110900.0 177100.00000000003 111700.0 176300.0 ;
      RECT  110900.0 177100.00000000003 111700.0 176300.0 ;
      RECT  109300.0 177100.00000000003 110100.0 176300.0 ;
      RECT  112500.0 170500.0 113300.00000000001 169700.0 ;
      RECT  112500.0 177100.00000000003 113300.00000000001 176300.0 ;
      RECT  109700.0 174000.0 110500.0 173200.0 ;
      RECT  109700.0 174000.0 110500.0 173200.0 ;
      RECT  111400.0 173899.99999999997 112000.0 173300.0 ;
      RECT  108100.0 169100.00000000003 114500.0 168500.0 ;
      RECT  108100.0 178300.0 114500.0 177700.0 ;
      RECT  112500.0 185900.00000000003 113300.00000000001 187200.0 ;
      RECT  112500.0 178000.0 113300.00000000001 179300.0 ;
      RECT  109300.0 178899.99999999997 110100.0 177700.0 ;
      RECT  109300.0 185100.00000000003 110100.0 187500.0 ;
      RECT  111100.0 178899.99999999997 111700.0 185100.00000000003 ;
      RECT  109300.0 185100.00000000003 110100.0 185900.00000000003 ;
      RECT  110900.0 185100.00000000003 111700.0 185900.00000000003 ;
      RECT  110900.0 185100.00000000003 111700.0 185900.00000000003 ;
      RECT  109300.0 185100.00000000003 110100.0 185900.00000000003 ;
      RECT  109300.0 178899.99999999997 110100.0 179700.0 ;
      RECT  110900.0 178899.99999999997 111700.0 179700.0 ;
      RECT  110900.0 178899.99999999997 111700.0 179700.0 ;
      RECT  109300.0 178899.99999999997 110100.0 179700.0 ;
      RECT  112500.0 185500.0 113300.00000000001 186300.0 ;
      RECT  112500.0 178899.99999999997 113300.00000000001 179700.0 ;
      RECT  109700.0 182000.0 110500.0 182800.0 ;
      RECT  109700.0 182000.0 110500.0 182800.0 ;
      RECT  111400.0 182100.00000000003 112000.0 182700.0 ;
      RECT  108100.0 186899.99999999997 114500.0 187500.0 ;
      RECT  108100.0 177700.0 114500.0 178300.0 ;
      RECT  112500.0 188500.0 113300.00000000001 187200.0 ;
      RECT  112500.0 196399.99999999997 113300.00000000001 195100.00000000003 ;
      RECT  109300.0 195500.0 110100.0 196700.0 ;
      RECT  109300.0 189300.0 110100.0 186899.99999999997 ;
      RECT  111100.0 195500.0 111700.0 189300.0 ;
      RECT  109300.0 189300.0 110100.0 188500.0 ;
      RECT  110900.0 189300.0 111700.0 188500.0 ;
      RECT  110900.0 189300.0 111700.0 188500.0 ;
      RECT  109300.0 189300.0 110100.0 188500.0 ;
      RECT  109300.0 195500.0 110100.0 194700.0 ;
      RECT  110900.0 195500.0 111700.0 194700.0 ;
      RECT  110900.0 195500.0 111700.0 194700.0 ;
      RECT  109300.0 195500.0 110100.0 194700.0 ;
      RECT  112500.0 188899.99999999997 113300.00000000001 188100.00000000003 ;
      RECT  112500.0 195500.0 113300.00000000001 194700.0 ;
      RECT  109700.0 192399.99999999997 110500.0 191600.00000000003 ;
      RECT  109700.0 192399.99999999997 110500.0 191600.00000000003 ;
      RECT  111400.0 192300.0 112000.0 191700.0 ;
      RECT  108100.0 187500.0 114500.0 186899.99999999997 ;
      RECT  108100.0 196700.0 114500.0 196100.00000000003 ;
      RECT  99700.0 160899.99999999997 100500.0 159300.0 ;
      RECT  99700.0 166700.0 100500.0 169100.00000000003 ;
      RECT  102900.0 166700.0 103700.0 169100.00000000003 ;
      RECT  104500.0 167500.0 105300.0 168800.0 ;
      RECT  104500.0 159600.00000000003 105300.0 160899.99999999997 ;
      RECT  99700.0 166700.0 100500.0 167500.0 ;
      RECT  101300.0 166700.0 102100.0 167500.0 ;
      RECT  101300.0 166700.0 102100.0 167500.0 ;
      RECT  99700.0 166700.0 100500.0 167500.0 ;
      RECT  101300.0 166700.0 102100.0 167500.0 ;
      RECT  102900.0 166700.0 103700.0 167500.0 ;
      RECT  102900.0 166700.0 103700.0 167500.0 ;
      RECT  101300.0 166700.0 102100.0 167500.0 ;
      RECT  99700.0 160899.99999999997 100500.0 161700.0 ;
      RECT  101300.0 160899.99999999997 102100.0 161700.0 ;
      RECT  101300.0 160899.99999999997 102100.0 161700.0 ;
      RECT  99700.0 160899.99999999997 100500.0 161700.0 ;
      RECT  101300.0 160899.99999999997 102100.0 161700.0 ;
      RECT  102900.0 160899.99999999997 103700.0 161700.0 ;
      RECT  102900.0 160899.99999999997 103700.0 161700.0 ;
      RECT  101300.0 160899.99999999997 102100.0 161700.0 ;
      RECT  104500.0 167100.00000000003 105300.0 167899.99999999997 ;
      RECT  104500.0 160500.0 105300.0 161300.0 ;
      RECT  102900.0 162600.00000000003 102100.0 163399.99999999997 ;
      RECT  100900.0 164000.0 100100.0 164800.0 ;
      RECT  101300.0 166700.0 102100.0 167500.0 ;
      RECT  102900.0 160899.99999999997 103700.0 161700.0 ;
      RECT  103700.0 164000.0 102900.0 164800.0 ;
      RECT  100100.0 164000.0 100900.0 164800.0 ;
      RECT  102100.0 162600.00000000003 102900.0 163399.99999999997 ;
      RECT  102900.0 164000.0 103700.0 164800.0 ;
      RECT  98500.0 168500.0 108100.0 169100.00000000003 ;
      RECT  98500.0 159300.0 108100.0 159899.99999999997 ;
      RECT  99700.0 176700.0 100500.0 178300.0 ;
      RECT  99700.0 170899.99999999997 100500.0 168500.0 ;
      RECT  102900.0 170899.99999999997 103700.0 168500.0 ;
      RECT  104500.0 170100.00000000003 105300.0 168800.0 ;
      RECT  104500.0 178000.0 105300.0 176700.0 ;
      RECT  99700.0 170900.00000000003 100500.0 170100.00000000003 ;
      RECT  101300.0 170900.00000000003 102100.0 170100.00000000003 ;
      RECT  101300.0 170900.00000000003 102100.0 170100.00000000003 ;
      RECT  99700.0 170900.00000000003 100500.0 170100.00000000003 ;
      RECT  101300.0 170900.00000000003 102100.0 170100.00000000003 ;
      RECT  102900.0 170900.00000000003 103700.0 170100.00000000003 ;
      RECT  102900.0 170900.00000000003 103700.0 170100.00000000003 ;
      RECT  101300.0 170900.00000000003 102100.0 170100.00000000003 ;
      RECT  99700.0 176700.0 100500.0 175899.99999999997 ;
      RECT  101300.0 176700.0 102100.0 175899.99999999997 ;
      RECT  101300.0 176700.0 102100.0 175899.99999999997 ;
      RECT  99700.0 176700.0 100500.0 175899.99999999997 ;
      RECT  101300.0 176700.0 102100.0 175899.99999999997 ;
      RECT  102900.0 176700.0 103700.0 175899.99999999997 ;
      RECT  102900.0 176700.0 103700.0 175899.99999999997 ;
      RECT  101300.0 176700.0 102100.0 175899.99999999997 ;
      RECT  104500.0 170500.0 105300.0 169700.0 ;
      RECT  104500.0 177100.00000000003 105300.0 176300.0 ;
      RECT  102900.0 175000.0 102100.0 174200.0 ;
      RECT  100900.0 173600.00000000003 100100.0 172800.0 ;
      RECT  101300.0 170899.99999999997 102100.0 170100.00000000003 ;
      RECT  102900.0 176700.0 103700.0 175899.99999999997 ;
      RECT  103700.0 173600.00000000003 102900.0 172800.0 ;
      RECT  100100.0 173600.00000000003 100900.0 172800.0 ;
      RECT  102100.0 175000.0 102900.0 174200.0 ;
      RECT  102900.0 173600.00000000003 103700.0 172800.0 ;
      RECT  98500.0 169100.00000000003 108100.0 168500.0 ;
      RECT  98500.0 178300.0 108100.0 177700.0 ;
      RECT  99700.0 179300.0 100500.0 177700.0 ;
      RECT  99700.0 185100.00000000003 100500.0 187500.0 ;
      RECT  102900.0 185100.00000000003 103700.0 187500.0 ;
      RECT  104500.0 185900.00000000003 105300.0 187200.0 ;
      RECT  104500.0 178000.0 105300.0 179300.0 ;
      RECT  99700.0 185100.00000000003 100500.0 185900.00000000003 ;
      RECT  101300.0 185100.00000000003 102100.0 185900.00000000003 ;
      RECT  101300.0 185100.00000000003 102100.0 185900.00000000003 ;
      RECT  99700.0 185100.00000000003 100500.0 185900.00000000003 ;
      RECT  101300.0 185100.00000000003 102100.0 185900.00000000003 ;
      RECT  102900.0 185100.00000000003 103700.0 185900.00000000003 ;
      RECT  102900.0 185100.00000000003 103700.0 185900.00000000003 ;
      RECT  101300.0 185100.00000000003 102100.0 185900.00000000003 ;
      RECT  99700.0 179300.0 100500.0 180100.00000000003 ;
      RECT  101300.0 179300.0 102100.0 180100.00000000003 ;
      RECT  101300.0 179300.0 102100.0 180100.00000000003 ;
      RECT  99700.0 179300.0 100500.0 180100.00000000003 ;
      RECT  101300.0 179300.0 102100.0 180100.00000000003 ;
      RECT  102900.0 179300.0 103700.0 180100.00000000003 ;
      RECT  102900.0 179300.0 103700.0 180100.00000000003 ;
      RECT  101300.0 179300.0 102100.0 180100.00000000003 ;
      RECT  104500.0 185500.0 105300.0 186300.0 ;
      RECT  104500.0 178899.99999999997 105300.0 179700.0 ;
      RECT  102900.0 181000.0 102100.0 181800.0 ;
      RECT  100900.0 182400.00000000003 100100.0 183200.0 ;
      RECT  101300.0 185100.00000000003 102100.0 185900.00000000003 ;
      RECT  102900.0 179300.0 103700.0 180100.00000000003 ;
      RECT  103700.0 182400.00000000003 102900.0 183200.0 ;
      RECT  100100.0 182400.00000000003 100900.0 183200.0 ;
      RECT  102100.0 181000.0 102900.0 181800.0 ;
      RECT  102900.0 182400.00000000003 103700.0 183200.0 ;
      RECT  98500.0 186899.99999999997 108100.0 187500.0 ;
      RECT  98500.0 177700.0 108100.0 178300.0 ;
      RECT  99700.0 195100.00000000003 100500.0 196700.0 ;
      RECT  99700.0 189300.0 100500.0 186899.99999999997 ;
      RECT  102900.0 189300.0 103700.0 186899.99999999997 ;
      RECT  104500.0 188500.0 105300.0 187200.0 ;
      RECT  104500.0 196399.99999999997 105300.0 195100.00000000003 ;
      RECT  99700.0 189300.0 100500.0 188500.0 ;
      RECT  101300.0 189300.0 102100.0 188500.0 ;
      RECT  101300.0 189300.0 102100.0 188500.0 ;
      RECT  99700.0 189300.0 100500.0 188500.0 ;
      RECT  101300.0 189300.0 102100.0 188500.0 ;
      RECT  102900.0 189300.0 103700.0 188500.0 ;
      RECT  102900.0 189300.0 103700.0 188500.0 ;
      RECT  101300.0 189300.0 102100.0 188500.0 ;
      RECT  99700.0 195100.00000000003 100500.0 194300.0 ;
      RECT  101300.0 195100.00000000003 102100.0 194300.0 ;
      RECT  101300.0 195100.00000000003 102100.0 194300.0 ;
      RECT  99700.0 195100.00000000003 100500.0 194300.0 ;
      RECT  101300.0 195100.00000000003 102100.0 194300.0 ;
      RECT  102900.0 195100.00000000003 103700.0 194300.0 ;
      RECT  102900.0 195100.00000000003 103700.0 194300.0 ;
      RECT  101300.0 195100.00000000003 102100.0 194300.0 ;
      RECT  104500.0 188899.99999999997 105300.0 188100.00000000003 ;
      RECT  104500.0 195500.0 105300.0 194700.0 ;
      RECT  102900.0 193399.99999999997 102100.0 192600.00000000003 ;
      RECT  100900.0 192000.0 100100.0 191200.0 ;
      RECT  101300.0 189300.0 102100.0 188500.0 ;
      RECT  102900.0 195100.00000000003 103700.0 194300.0 ;
      RECT  103700.0 192000.0 102900.0 191200.0 ;
      RECT  100100.0 192000.0 100900.0 191200.0 ;
      RECT  102100.0 193399.99999999997 102900.0 192600.00000000003 ;
      RECT  102900.0 192000.0 103700.0 191200.0 ;
      RECT  98500.0 187500.0 108100.0 186899.99999999997 ;
      RECT  98500.0 196700.0 108100.0 196100.00000000003 ;
      RECT  93600.0 166600.00000000003 92800.0 167399.99999999997 ;
      RECT  81900.0 163600.00000000003 81100.0 164399.99999999997 ;
      RECT  95000.0 175800.0 94200.0 176600.00000000003 ;
      RECT  83300.0 173200.0 82500.0 174000.0 ;
      RECT  81900.0 179000.0 81100.0 179800.0 ;
      RECT  96400.0 179000.0 95600.0 179800.0 ;
      RECT  83300.0 188200.0 82500.0 189000.0 ;
      RECT  97800.0 188200.0 97000.0 189000.0 ;
      RECT  93600.0 164000.0 92800.0 164800.0 ;
      RECT  95000.0 162600.00000000003 94200.0 163399.99999999997 ;
      RECT  96400.0 172800.0 95600.0 173600.00000000003 ;
      RECT  95000.0 174200.0 94200.0 175000.0 ;
      RECT  93600.0 182399.99999999997 92800.0 183200.0 ;
      RECT  97800.0 181000.0 97000.0 181800.0 ;
      RECT  96400.0 191200.0 95600.0 192000.0 ;
      RECT  97800.0 192600.00000000003 97000.0 193399.99999999997 ;
      RECT  90500.0 168399.99999999997 89700.0 169200.0 ;
      RECT  108500.0 168399.99999999997 107700.0 169200.0 ;
      RECT  90500.0 159200.0 89700.0 160000.0 ;
      RECT  108500.0 159200.0 107700.0 160000.0 ;
      RECT  90500.0 168399.99999999997 89700.0 169200.0 ;
      RECT  108500.0 168399.99999999997 107700.0 169200.0 ;
      RECT  90500.0 177600.00000000003 89700.0 178399.99999999997 ;
      RECT  108500.0 177600.00000000003 107700.0 178399.99999999997 ;
      RECT  90500.0 186800.0 89700.0 187600.00000000003 ;
      RECT  108500.0 186800.0 107700.0 187600.00000000003 ;
      RECT  90500.0 177600.00000000003 89700.0 178399.99999999997 ;
      RECT  108500.0 177600.00000000003 107700.0 178399.99999999997 ;
      RECT  90500.0 186800.0 89700.0 187600.00000000003 ;
      RECT  108500.0 186800.0 107700.0 187600.00000000003 ;
      RECT  90500.0 196000.0 89700.0 196800.0 ;
      RECT  108500.0 196000.0 107700.0 196800.0 ;
      RECT  111400.0 163700.0 112000.0 164300.0 ;
      RECT  111400.0 173300.0 112000.0 173899.99999999997 ;
      RECT  111400.0 182100.00000000003 112000.0 182700.0 ;
      RECT  111400.0 191700.0 112000.0 192300.0 ;
      RECT  126900.0 124100.00000000001 127700.0 122500.0 ;
      RECT  126900.0 129900.0 127700.0 132300.0 ;
      RECT  130100.0 129900.0 130900.0 132300.0 ;
      RECT  131700.0 130699.99999999999 132500.0 132000.0 ;
      RECT  131700.0 122800.00000000001 132500.0 124100.00000000001 ;
      RECT  126900.0 129900.0 127700.0 130699.99999999999 ;
      RECT  128500.0 129900.0 129300.00000000001 130699.99999999999 ;
      RECT  128500.0 129900.0 129300.00000000001 130699.99999999999 ;
      RECT  126900.0 129900.0 127700.0 130699.99999999999 ;
      RECT  128500.0 129900.0 129300.00000000001 130699.99999999999 ;
      RECT  130100.0 129900.0 130900.0 130699.99999999999 ;
      RECT  130100.0 129900.0 130900.0 130699.99999999999 ;
      RECT  128500.0 129900.0 129300.00000000001 130699.99999999999 ;
      RECT  126900.0 124100.00000000001 127700.0 124900.0 ;
      RECT  128500.0 124100.00000000001 129300.00000000001 124900.0 ;
      RECT  128500.0 124100.00000000001 129300.00000000001 124900.0 ;
      RECT  126900.0 124100.00000000001 127700.0 124900.0 ;
      RECT  128500.0 124100.00000000001 129300.00000000001 124900.0 ;
      RECT  130100.0 124100.00000000001 130900.0 124900.0 ;
      RECT  130100.0 124100.00000000001 130900.0 124900.0 ;
      RECT  128500.0 124100.00000000001 129300.00000000001 124900.0 ;
      RECT  131700.0 130300.00000000001 132500.0 131100.00000000003 ;
      RECT  131700.0 123700.0 132500.0 124500.0 ;
      RECT  130100.0 125800.00000000001 129300.00000000001 126600.00000000001 ;
      RECT  128100.0 127200.0 127300.00000000001 128000.0 ;
      RECT  128500.0 129900.0 129300.00000000001 130699.99999999999 ;
      RECT  130100.0 124100.00000000001 130900.0 124900.0 ;
      RECT  130900.0 127200.0 130100.0 128000.0 ;
      RECT  127300.00000000001 127200.0 128100.0 128000.0 ;
      RECT  129300.00000000001 125800.00000000001 130100.0 126600.00000000001 ;
      RECT  130100.0 127200.0 130900.0 128000.0 ;
      RECT  125700.0 131700.0 135300.0 132300.0 ;
      RECT  125700.0 122500.0 135300.0 123100.00000000001 ;
      RECT  126900.0 139900.0 127700.0 141500.0 ;
      RECT  126900.0 134100.00000000003 127700.0 131700.0 ;
      RECT  130100.0 134100.00000000003 130900.0 131700.0 ;
      RECT  131700.0 133300.0 132500.0 132000.0 ;
      RECT  131700.0 141200.0 132500.0 139900.0 ;
      RECT  126900.0 134100.00000000003 127700.0 133300.0 ;
      RECT  128500.0 134100.00000000003 129300.00000000001 133300.0 ;
      RECT  128500.0 134100.00000000003 129300.00000000001 133300.0 ;
      RECT  126900.0 134100.00000000003 127700.0 133300.0 ;
      RECT  128500.0 134100.00000000003 129300.00000000001 133300.0 ;
      RECT  130100.0 134100.00000000003 130900.0 133300.0 ;
      RECT  130100.0 134100.00000000003 130900.0 133300.0 ;
      RECT  128500.0 134100.00000000003 129300.00000000001 133300.0 ;
      RECT  126900.0 139900.0 127700.0 139100.00000000003 ;
      RECT  128500.0 139900.0 129300.00000000001 139100.00000000003 ;
      RECT  128500.0 139900.0 129300.00000000001 139100.00000000003 ;
      RECT  126900.0 139900.0 127700.0 139100.00000000003 ;
      RECT  128500.0 139900.0 129300.00000000001 139100.00000000003 ;
      RECT  130100.0 139900.0 130900.0 139100.00000000003 ;
      RECT  130100.0 139900.0 130900.0 139100.00000000003 ;
      RECT  128500.0 139900.0 129300.00000000001 139100.00000000003 ;
      RECT  131700.0 133700.0 132500.0 132900.0 ;
      RECT  131700.0 140300.0 132500.0 139500.0 ;
      RECT  130100.0 138200.0 129300.00000000001 137400.0 ;
      RECT  128100.0 136800.0 127300.00000000001 136000.0 ;
      RECT  128500.0 134100.00000000003 129300.00000000001 133300.0 ;
      RECT  130100.0 139900.0 130900.0 139100.00000000003 ;
      RECT  130900.0 136800.0 130100.0 136000.0 ;
      RECT  127300.00000000001 136800.0 128100.0 136000.0 ;
      RECT  129300.00000000001 138200.0 130100.0 137400.0 ;
      RECT  130100.0 136800.0 130900.0 136000.0 ;
      RECT  125700.0 132300.0 135300.0 131700.0 ;
      RECT  125700.0 141500.0 135300.0 140900.0 ;
      RECT  126900.0 142500.0 127700.0 140900.0 ;
      RECT  126900.0 148300.0 127700.0 150700.0 ;
      RECT  130100.0 148300.0 130900.0 150700.0 ;
      RECT  131700.0 149100.00000000003 132500.0 150400.0 ;
      RECT  131700.0 141200.0 132500.0 142500.0 ;
      RECT  126900.0 148300.0 127700.0 149100.00000000003 ;
      RECT  128500.0 148300.0 129300.00000000001 149100.00000000003 ;
      RECT  128500.0 148300.0 129300.00000000001 149100.00000000003 ;
      RECT  126900.0 148300.0 127700.0 149100.00000000003 ;
      RECT  128500.0 148300.0 129300.00000000001 149100.00000000003 ;
      RECT  130100.0 148300.0 130900.0 149100.00000000003 ;
      RECT  130100.0 148300.0 130900.0 149100.00000000003 ;
      RECT  128500.0 148300.0 129300.00000000001 149100.00000000003 ;
      RECT  126900.0 142500.0 127700.0 143300.0 ;
      RECT  128500.0 142500.0 129300.00000000001 143300.0 ;
      RECT  128500.0 142500.0 129300.00000000001 143300.0 ;
      RECT  126900.0 142500.0 127700.0 143300.0 ;
      RECT  128500.0 142500.0 129300.00000000001 143300.0 ;
      RECT  130100.0 142500.0 130900.0 143300.0 ;
      RECT  130100.0 142500.0 130900.0 143300.0 ;
      RECT  128500.0 142500.0 129300.00000000001 143300.0 ;
      RECT  131700.0 148700.0 132500.0 149500.0 ;
      RECT  131700.0 142100.00000000003 132500.0 142900.0 ;
      RECT  130100.0 144200.0 129300.00000000001 145000.0 ;
      RECT  128100.0 145600.00000000003 127300.00000000001 146400.0 ;
      RECT  128500.0 148300.0 129300.00000000001 149100.00000000003 ;
      RECT  130100.0 142500.0 130900.0 143300.0 ;
      RECT  130900.0 145600.00000000003 130100.0 146400.0 ;
      RECT  127300.00000000001 145600.00000000003 128100.0 146400.0 ;
      RECT  129300.00000000001 144200.0 130100.0 145000.0 ;
      RECT  130100.0 145600.00000000003 130900.0 146400.0 ;
      RECT  125700.0 150100.00000000003 135300.0 150700.0 ;
      RECT  125700.0 140900.0 135300.0 141500.0 ;
      RECT  126900.0 158300.0 127700.0 159899.99999999997 ;
      RECT  126900.0 152500.0 127700.0 150100.00000000003 ;
      RECT  130100.0 152500.0 130900.0 150100.00000000003 ;
      RECT  131700.0 151700.0 132500.0 150400.0 ;
      RECT  131700.0 159600.00000000003 132500.0 158300.0 ;
      RECT  126900.0 152500.0 127700.0 151700.0 ;
      RECT  128500.0 152500.0 129300.00000000001 151700.0 ;
      RECT  128500.0 152500.0 129300.00000000001 151700.0 ;
      RECT  126900.0 152500.0 127700.0 151700.0 ;
      RECT  128500.0 152500.0 129300.00000000001 151700.0 ;
      RECT  130100.0 152500.0 130900.0 151700.0 ;
      RECT  130100.0 152500.0 130900.0 151700.0 ;
      RECT  128500.0 152500.0 129300.00000000001 151700.0 ;
      RECT  126900.0 158300.0 127700.0 157500.0 ;
      RECT  128500.0 158300.0 129300.00000000001 157500.0 ;
      RECT  128500.0 158300.0 129300.00000000001 157500.0 ;
      RECT  126900.0 158300.0 127700.0 157500.0 ;
      RECT  128500.0 158300.0 129300.00000000001 157500.0 ;
      RECT  130100.0 158300.0 130900.0 157500.0 ;
      RECT  130100.0 158300.0 130900.0 157500.0 ;
      RECT  128500.0 158300.0 129300.00000000001 157500.0 ;
      RECT  131700.0 152100.00000000003 132500.0 151300.0 ;
      RECT  131700.0 158700.0 132500.0 157899.99999999997 ;
      RECT  130100.0 156600.00000000003 129300.00000000001 155800.0 ;
      RECT  128100.0 155200.0 127300.00000000001 154399.99999999997 ;
      RECT  128500.0 152500.0 129300.00000000001 151700.0 ;
      RECT  130100.0 158300.0 130900.0 157500.0 ;
      RECT  130900.0 155200.0 130100.0 154399.99999999997 ;
      RECT  127300.00000000001 155200.0 128100.0 154399.99999999997 ;
      RECT  129300.00000000001 156600.00000000003 130100.0 155800.0 ;
      RECT  130100.0 155200.0 130900.0 154399.99999999997 ;
      RECT  125700.0 150700.0 135300.0 150100.00000000003 ;
      RECT  125700.0 159899.99999999997 135300.0 159300.0 ;
      RECT  126900.0 160899.99999999997 127700.0 159300.0 ;
      RECT  126900.0 166700.0 127700.0 169100.00000000003 ;
      RECT  130100.0 166700.0 130900.0 169100.00000000003 ;
      RECT  131700.0 167500.0 132500.0 168800.0 ;
      RECT  131700.0 159600.00000000003 132500.0 160899.99999999997 ;
      RECT  126900.0 166700.0 127700.0 167500.0 ;
      RECT  128500.0 166700.0 129300.00000000001 167500.0 ;
      RECT  128500.0 166700.0 129300.00000000001 167500.0 ;
      RECT  126900.0 166700.0 127700.0 167500.0 ;
      RECT  128500.0 166700.0 129300.00000000001 167500.0 ;
      RECT  130100.0 166700.0 130900.0 167500.0 ;
      RECT  130100.0 166700.0 130900.0 167500.0 ;
      RECT  128500.0 166700.0 129300.00000000001 167500.0 ;
      RECT  126900.0 160899.99999999997 127700.0 161700.0 ;
      RECT  128500.0 160899.99999999997 129300.00000000001 161700.0 ;
      RECT  128500.0 160899.99999999997 129300.00000000001 161700.0 ;
      RECT  126900.0 160899.99999999997 127700.0 161700.0 ;
      RECT  128500.0 160899.99999999997 129300.00000000001 161700.0 ;
      RECT  130100.0 160899.99999999997 130900.0 161700.0 ;
      RECT  130100.0 160899.99999999997 130900.0 161700.0 ;
      RECT  128500.0 160899.99999999997 129300.00000000001 161700.0 ;
      RECT  131700.0 167100.00000000003 132500.0 167899.99999999997 ;
      RECT  131700.0 160500.0 132500.0 161300.0 ;
      RECT  130100.0 162600.00000000003 129300.00000000001 163399.99999999997 ;
      RECT  128100.0 164000.0 127300.00000000001 164800.0 ;
      RECT  128500.0 166700.0 129300.00000000001 167500.0 ;
      RECT  130100.0 160899.99999999997 130900.0 161700.0 ;
      RECT  130900.0 164000.0 130100.0 164800.0 ;
      RECT  127300.00000000001 164000.0 128100.0 164800.0 ;
      RECT  129300.00000000001 162600.00000000003 130100.0 163399.99999999997 ;
      RECT  130100.0 164000.0 130900.0 164800.0 ;
      RECT  125700.0 168500.0 135300.0 169100.00000000003 ;
      RECT  125700.0 159300.0 135300.0 159899.99999999997 ;
      RECT  126900.0 176700.0 127700.0 178300.0 ;
      RECT  126900.0 170899.99999999997 127700.0 168500.0 ;
      RECT  130100.0 170899.99999999997 130900.0 168500.0 ;
      RECT  131700.0 170100.00000000003 132500.0 168800.0 ;
      RECT  131700.0 178000.0 132500.0 176700.0 ;
      RECT  126900.0 170899.99999999997 127700.0 170100.00000000003 ;
      RECT  128500.0 170899.99999999997 129300.00000000001 170100.00000000003 ;
      RECT  128500.0 170899.99999999997 129300.00000000001 170100.00000000003 ;
      RECT  126900.0 170899.99999999997 127700.0 170100.00000000003 ;
      RECT  128500.0 170899.99999999997 129300.00000000001 170100.00000000003 ;
      RECT  130100.0 170899.99999999997 130900.0 170100.00000000003 ;
      RECT  130100.0 170899.99999999997 130900.0 170100.00000000003 ;
      RECT  128500.0 170899.99999999997 129300.00000000001 170100.00000000003 ;
      RECT  126900.0 176700.0 127700.0 175899.99999999997 ;
      RECT  128500.0 176700.0 129300.00000000001 175899.99999999997 ;
      RECT  128500.0 176700.0 129300.00000000001 175899.99999999997 ;
      RECT  126900.0 176700.0 127700.0 175899.99999999997 ;
      RECT  128500.0 176700.0 129300.00000000001 175899.99999999997 ;
      RECT  130100.0 176700.0 130900.0 175899.99999999997 ;
      RECT  130100.0 176700.0 130900.0 175899.99999999997 ;
      RECT  128500.0 176700.0 129300.00000000001 175899.99999999997 ;
      RECT  131700.0 170500.0 132500.0 169700.0 ;
      RECT  131700.0 177100.00000000003 132500.0 176300.0 ;
      RECT  130100.0 175000.0 129300.00000000001 174200.0 ;
      RECT  128100.0 173600.00000000003 127300.00000000001 172800.0 ;
      RECT  128500.0 170899.99999999997 129300.00000000001 170100.00000000003 ;
      RECT  130100.0 176700.0 130900.0 175899.99999999997 ;
      RECT  130900.0 173600.00000000003 130100.0 172800.0 ;
      RECT  127300.00000000001 173600.00000000003 128100.0 172800.0 ;
      RECT  129300.00000000001 175000.0 130100.0 174200.0 ;
      RECT  130100.0 173600.00000000003 130900.0 172800.0 ;
      RECT  125700.0 169100.00000000003 135300.0 168500.0 ;
      RECT  125700.0 178300.0 135300.0 177700.0 ;
      RECT  126900.0 179300.0 127700.0 177700.0 ;
      RECT  126900.0 185100.00000000003 127700.0 187500.0 ;
      RECT  130100.0 185100.00000000003 130900.0 187500.0 ;
      RECT  131700.0 185899.99999999997 132500.0 187200.0 ;
      RECT  131700.0 178000.0 132500.0 179300.0 ;
      RECT  126900.0 185100.00000000003 127700.0 185899.99999999997 ;
      RECT  128500.0 185100.00000000003 129300.00000000001 185899.99999999997 ;
      RECT  128500.0 185100.00000000003 129300.00000000001 185899.99999999997 ;
      RECT  126900.0 185100.00000000003 127700.0 185899.99999999997 ;
      RECT  128500.0 185100.00000000003 129300.00000000001 185899.99999999997 ;
      RECT  130100.0 185100.00000000003 130900.0 185899.99999999997 ;
      RECT  130100.0 185100.00000000003 130900.0 185899.99999999997 ;
      RECT  128500.0 185100.00000000003 129300.00000000001 185899.99999999997 ;
      RECT  126900.0 179300.0 127700.0 180100.00000000003 ;
      RECT  128500.0 179300.0 129300.00000000001 180100.00000000003 ;
      RECT  128500.0 179300.0 129300.00000000001 180100.00000000003 ;
      RECT  126900.0 179300.0 127700.0 180100.00000000003 ;
      RECT  128500.0 179300.0 129300.00000000001 180100.00000000003 ;
      RECT  130100.0 179300.0 130900.0 180100.00000000003 ;
      RECT  130100.0 179300.0 130900.0 180100.00000000003 ;
      RECT  128500.0 179300.0 129300.00000000001 180100.00000000003 ;
      RECT  131700.0 185500.0 132500.0 186300.0 ;
      RECT  131700.0 178899.99999999997 132500.0 179700.0 ;
      RECT  130100.0 181000.0 129300.00000000001 181800.0 ;
      RECT  128100.0 182399.99999999997 127300.00000000001 183200.0 ;
      RECT  128500.0 185100.00000000003 129300.00000000001 185899.99999999997 ;
      RECT  130100.0 179300.0 130900.0 180100.00000000003 ;
      RECT  130900.0 182399.99999999997 130100.0 183200.0 ;
      RECT  127300.00000000001 182399.99999999997 128100.0 183200.0 ;
      RECT  129300.00000000001 181000.0 130100.0 181800.0 ;
      RECT  130100.0 182399.99999999997 130900.0 183200.0 ;
      RECT  125700.0 186899.99999999997 135300.0 187500.0 ;
      RECT  125700.0 177700.0 135300.0 178300.0 ;
      RECT  126900.0 195100.00000000003 127700.0 196700.0 ;
      RECT  126900.0 189300.0 127700.0 186900.00000000003 ;
      RECT  130100.0 189300.0 130900.0 186900.00000000003 ;
      RECT  131700.0 188500.0 132500.0 187200.0 ;
      RECT  131700.0 196400.00000000003 132500.0 195100.00000000003 ;
      RECT  126900.0 189300.0 127700.0 188500.0 ;
      RECT  128500.0 189300.0 129300.00000000001 188500.0 ;
      RECT  128500.0 189300.0 129300.00000000001 188500.0 ;
      RECT  126900.0 189300.0 127700.0 188500.0 ;
      RECT  128500.0 189300.0 129300.00000000001 188500.0 ;
      RECT  130100.0 189300.0 130900.0 188500.0 ;
      RECT  130100.0 189300.0 130900.0 188500.0 ;
      RECT  128500.0 189300.0 129300.00000000001 188500.0 ;
      RECT  126900.0 195100.00000000003 127700.0 194300.0 ;
      RECT  128500.0 195100.00000000003 129300.00000000001 194300.0 ;
      RECT  128500.0 195100.00000000003 129300.00000000001 194300.0 ;
      RECT  126900.0 195100.00000000003 127700.0 194300.0 ;
      RECT  128500.0 195100.00000000003 129300.00000000001 194300.0 ;
      RECT  130100.0 195100.00000000003 130900.0 194300.0 ;
      RECT  130100.0 195100.00000000003 130900.0 194300.0 ;
      RECT  128500.0 195100.00000000003 129300.00000000001 194300.0 ;
      RECT  131700.0 188900.00000000003 132500.0 188100.00000000003 ;
      RECT  131700.0 195500.0 132500.0 194700.0 ;
      RECT  130100.0 193400.00000000003 129300.00000000001 192600.00000000003 ;
      RECT  128100.0 192000.0 127300.00000000001 191200.0 ;
      RECT  128500.0 189300.0 129300.00000000001 188500.0 ;
      RECT  130100.0 195100.00000000003 130900.0 194300.0 ;
      RECT  130900.0 192000.0 130100.0 191200.0 ;
      RECT  127300.00000000001 192000.0 128100.0 191200.0 ;
      RECT  129300.00000000001 193400.00000000003 130100.0 192600.00000000003 ;
      RECT  130100.0 192000.0 130900.0 191200.0 ;
      RECT  125700.0 187500.0 135300.0 186900.00000000003 ;
      RECT  125700.0 196700.0 135300.0 196100.00000000003 ;
      RECT  126900.0 197700.0 127700.0 196100.00000000003 ;
      RECT  126900.0 203500.0 127700.0 205900.00000000003 ;
      RECT  130100.0 203500.0 130900.0 205900.00000000003 ;
      RECT  131700.0 204300.0 132500.0 205600.00000000003 ;
      RECT  131700.0 196400.00000000003 132500.0 197700.0 ;
      RECT  126900.0 203500.0 127700.0 204300.0 ;
      RECT  128500.0 203500.0 129300.00000000001 204300.0 ;
      RECT  128500.0 203500.0 129300.00000000001 204300.0 ;
      RECT  126900.0 203500.0 127700.0 204300.0 ;
      RECT  128500.0 203500.0 129300.00000000001 204300.0 ;
      RECT  130100.0 203500.0 130900.0 204300.0 ;
      RECT  130100.0 203500.0 130900.0 204300.0 ;
      RECT  128500.0 203500.0 129300.00000000001 204300.0 ;
      RECT  126900.0 197700.0 127700.0 198500.0 ;
      RECT  128500.0 197700.0 129300.00000000001 198500.0 ;
      RECT  128500.0 197700.0 129300.00000000001 198500.0 ;
      RECT  126900.0 197700.0 127700.0 198500.0 ;
      RECT  128500.0 197700.0 129300.00000000001 198500.0 ;
      RECT  130100.0 197700.0 130900.0 198500.0 ;
      RECT  130100.0 197700.0 130900.0 198500.0 ;
      RECT  128500.0 197700.0 129300.00000000001 198500.0 ;
      RECT  131700.0 203900.00000000003 132500.0 204700.0 ;
      RECT  131700.0 197300.0 132500.0 198100.00000000003 ;
      RECT  130100.0 199400.00000000003 129300.00000000001 200200.0 ;
      RECT  128100.0 200800.0 127300.00000000001 201600.00000000003 ;
      RECT  128500.0 203500.0 129300.00000000001 204300.0 ;
      RECT  130100.0 197700.0 130900.0 198500.0 ;
      RECT  130900.0 200800.0 130100.0 201600.00000000003 ;
      RECT  127300.00000000001 200800.0 128100.0 201600.00000000003 ;
      RECT  129300.00000000001 199400.00000000003 130100.0 200200.0 ;
      RECT  130100.0 200800.0 130900.0 201600.00000000003 ;
      RECT  125700.0 205300.0 135300.0 205900.00000000003 ;
      RECT  125700.0 196100.00000000003 135300.0 196700.0 ;
      RECT  126900.0 213500.0 127700.0 215100.00000000003 ;
      RECT  126900.0 207700.0 127700.0 205300.0 ;
      RECT  130100.0 207700.0 130900.0 205300.0 ;
      RECT  131700.0 206899.99999999997 132500.0 205600.00000000003 ;
      RECT  131700.0 214800.0 132500.0 213500.0 ;
      RECT  126900.0 207700.0 127700.0 206899.99999999997 ;
      RECT  128500.0 207700.0 129300.00000000001 206899.99999999997 ;
      RECT  128500.0 207700.0 129300.00000000001 206899.99999999997 ;
      RECT  126900.0 207700.0 127700.0 206899.99999999997 ;
      RECT  128500.0 207700.0 129300.00000000001 206899.99999999997 ;
      RECT  130100.0 207700.0 130900.0 206899.99999999997 ;
      RECT  130100.0 207700.0 130900.0 206899.99999999997 ;
      RECT  128500.0 207700.0 129300.00000000001 206899.99999999997 ;
      RECT  126900.0 213500.0 127700.0 212700.0 ;
      RECT  128500.0 213500.0 129300.00000000001 212700.0 ;
      RECT  128500.0 213500.0 129300.00000000001 212700.0 ;
      RECT  126900.0 213500.0 127700.0 212700.0 ;
      RECT  128500.0 213500.0 129300.00000000001 212700.0 ;
      RECT  130100.0 213500.0 130900.0 212700.0 ;
      RECT  130100.0 213500.0 130900.0 212700.0 ;
      RECT  128500.0 213500.0 129300.00000000001 212700.0 ;
      RECT  131700.0 207300.0 132500.0 206500.0 ;
      RECT  131700.0 213899.99999999997 132500.0 213100.00000000003 ;
      RECT  130100.0 211800.0 129300.00000000001 211000.0 ;
      RECT  128100.0 210399.99999999997 127300.00000000001 209600.00000000003 ;
      RECT  128500.0 207700.0 129300.00000000001 206899.99999999997 ;
      RECT  130100.0 213500.0 130900.0 212700.0 ;
      RECT  130900.0 210399.99999999997 130100.0 209600.00000000003 ;
      RECT  127300.00000000001 210399.99999999997 128100.0 209600.00000000003 ;
      RECT  129300.00000000001 211800.0 130100.0 211000.0 ;
      RECT  130100.0 210399.99999999997 130900.0 209600.00000000003 ;
      RECT  125700.0 205899.99999999997 135300.0 205300.0 ;
      RECT  125700.0 215100.00000000003 135300.0 214500.0 ;
      RECT  126900.0 216100.00000000003 127700.0 214500.0 ;
      RECT  126900.0 221899.99999999997 127700.0 224300.0 ;
      RECT  130100.0 221899.99999999997 130900.0 224300.0 ;
      RECT  131700.0 222700.0 132500.0 224000.0 ;
      RECT  131700.0 214800.0 132500.0 216100.00000000003 ;
      RECT  126900.0 221899.99999999997 127700.0 222700.0 ;
      RECT  128500.0 221899.99999999997 129300.00000000001 222700.0 ;
      RECT  128500.0 221899.99999999997 129300.00000000001 222700.0 ;
      RECT  126900.0 221899.99999999997 127700.0 222700.0 ;
      RECT  128500.0 221899.99999999997 129300.00000000001 222700.0 ;
      RECT  130100.0 221899.99999999997 130900.0 222700.0 ;
      RECT  130100.0 221899.99999999997 130900.0 222700.0 ;
      RECT  128500.0 221899.99999999997 129300.00000000001 222700.0 ;
      RECT  126900.0 216100.00000000003 127700.0 216899.99999999997 ;
      RECT  128500.0 216100.00000000003 129300.00000000001 216899.99999999997 ;
      RECT  128500.0 216100.00000000003 129300.00000000001 216899.99999999997 ;
      RECT  126900.0 216100.00000000003 127700.0 216899.99999999997 ;
      RECT  128500.0 216100.00000000003 129300.00000000001 216899.99999999997 ;
      RECT  130100.0 216100.00000000003 130900.0 216899.99999999997 ;
      RECT  130100.0 216100.00000000003 130900.0 216899.99999999997 ;
      RECT  128500.0 216100.00000000003 129300.00000000001 216899.99999999997 ;
      RECT  131700.0 222300.0 132500.0 223100.00000000003 ;
      RECT  131700.0 215700.0 132500.0 216500.0 ;
      RECT  130100.0 217800.0 129300.00000000001 218600.00000000003 ;
      RECT  128100.0 219200.0 127300.00000000001 220000.0 ;
      RECT  128500.0 221899.99999999997 129300.00000000001 222700.0 ;
      RECT  130100.0 216100.00000000003 130900.0 216899.99999999997 ;
      RECT  130900.0 219200.0 130100.0 220000.0 ;
      RECT  127300.00000000001 219200.0 128100.0 220000.0 ;
      RECT  129300.00000000001 217800.0 130100.0 218600.00000000003 ;
      RECT  130100.0 219200.0 130900.0 220000.0 ;
      RECT  125700.0 223700.0 135300.0 224300.0 ;
      RECT  125700.0 214500.0 135300.0 215100.00000000003 ;
      RECT  126900.0 231900.00000000003 127700.0 233500.0 ;
      RECT  126900.0 226100.00000000003 127700.0 223700.0 ;
      RECT  130100.0 226100.00000000003 130900.0 223700.0 ;
      RECT  131700.0 225300.0 132500.0 224000.0 ;
      RECT  131700.0 233200.0 132500.0 231900.00000000003 ;
      RECT  126900.0 226100.00000000003 127700.0 225300.0 ;
      RECT  128500.0 226100.00000000003 129300.00000000001 225300.0 ;
      RECT  128500.0 226100.00000000003 129300.00000000001 225300.0 ;
      RECT  126900.0 226100.00000000003 127700.0 225300.0 ;
      RECT  128500.0 226100.00000000003 129300.00000000001 225300.0 ;
      RECT  130100.0 226100.00000000003 130900.0 225300.0 ;
      RECT  130100.0 226100.00000000003 130900.0 225300.0 ;
      RECT  128500.0 226100.00000000003 129300.00000000001 225300.0 ;
      RECT  126900.0 231900.00000000003 127700.0 231100.00000000003 ;
      RECT  128500.0 231900.00000000003 129300.00000000001 231100.00000000003 ;
      RECT  128500.0 231900.00000000003 129300.00000000001 231100.00000000003 ;
      RECT  126900.0 231900.00000000003 127700.0 231100.00000000003 ;
      RECT  128500.0 231900.00000000003 129300.00000000001 231100.00000000003 ;
      RECT  130100.0 231900.00000000003 130900.0 231100.00000000003 ;
      RECT  130100.0 231900.00000000003 130900.0 231100.00000000003 ;
      RECT  128500.0 231900.00000000003 129300.00000000001 231100.00000000003 ;
      RECT  131700.0 225700.0 132500.0 224900.00000000003 ;
      RECT  131700.0 232300.0 132500.0 231500.0 ;
      RECT  130100.0 230200.0 129300.00000000001 229400.00000000003 ;
      RECT  128100.0 228800.0 127300.00000000001 228000.0 ;
      RECT  128500.0 226100.00000000003 129300.00000000001 225300.0 ;
      RECT  130100.0 231900.00000000003 130900.0 231100.00000000003 ;
      RECT  130900.0 228800.0 130100.0 228000.0 ;
      RECT  127300.00000000001 228800.0 128100.0 228000.0 ;
      RECT  129300.00000000001 230200.0 130100.0 229400.00000000003 ;
      RECT  130100.0 228800.0 130900.0 228000.0 ;
      RECT  125700.0 224300.0 135300.0 223700.0 ;
      RECT  125700.0 233500.0 135300.0 232900.00000000003 ;
      RECT  126900.0 234500.0 127700.0 232900.00000000003 ;
      RECT  126900.0 240300.0 127700.0 242700.0 ;
      RECT  130100.0 240300.0 130900.0 242700.0 ;
      RECT  131700.0 241100.00000000003 132500.0 242400.00000000003 ;
      RECT  131700.0 233200.0 132500.0 234500.0 ;
      RECT  126900.0 240300.0 127700.0 241100.00000000003 ;
      RECT  128500.0 240300.0 129300.00000000001 241100.00000000003 ;
      RECT  128500.0 240300.0 129300.00000000001 241100.00000000003 ;
      RECT  126900.0 240300.0 127700.0 241100.00000000003 ;
      RECT  128500.0 240300.0 129300.00000000001 241100.00000000003 ;
      RECT  130100.0 240300.0 130900.0 241100.00000000003 ;
      RECT  130100.0 240300.0 130900.0 241100.00000000003 ;
      RECT  128500.0 240300.0 129300.00000000001 241100.00000000003 ;
      RECT  126900.0 234500.0 127700.0 235300.0 ;
      RECT  128500.0 234500.0 129300.00000000001 235300.0 ;
      RECT  128500.0 234500.0 129300.00000000001 235300.0 ;
      RECT  126900.0 234500.0 127700.0 235300.0 ;
      RECT  128500.0 234500.0 129300.00000000001 235300.0 ;
      RECT  130100.0 234500.0 130900.0 235300.0 ;
      RECT  130100.0 234500.0 130900.0 235300.0 ;
      RECT  128500.0 234500.0 129300.00000000001 235300.0 ;
      RECT  131700.0 240700.0 132500.0 241500.0 ;
      RECT  131700.0 234100.00000000003 132500.0 234900.00000000003 ;
      RECT  130100.0 236200.0 129300.00000000001 237000.0 ;
      RECT  128100.0 237600.00000000003 127300.00000000001 238400.00000000003 ;
      RECT  128500.0 240300.0 129300.00000000001 241100.00000000003 ;
      RECT  130100.0 234500.0 130900.0 235300.0 ;
      RECT  130900.0 237600.00000000003 130100.0 238400.00000000003 ;
      RECT  127300.00000000001 237600.00000000003 128100.0 238400.00000000003 ;
      RECT  129300.00000000001 236200.0 130100.0 237000.0 ;
      RECT  130100.0 237600.00000000003 130900.0 238400.00000000003 ;
      RECT  125700.0 242100.00000000003 135300.0 242700.0 ;
      RECT  125700.0 232900.00000000003 135300.0 233500.0 ;
      RECT  126900.0 250300.0 127700.0 251900.00000000003 ;
      RECT  126900.0 244500.0 127700.0 242100.00000000003 ;
      RECT  130100.0 244500.0 130900.0 242100.00000000003 ;
      RECT  131700.0 243700.0 132500.0 242400.00000000003 ;
      RECT  131700.0 251600.00000000003 132500.0 250300.0 ;
      RECT  126900.0 244500.0 127700.0 243700.0 ;
      RECT  128500.0 244500.0 129300.00000000001 243700.0 ;
      RECT  128500.0 244500.0 129300.00000000001 243700.0 ;
      RECT  126900.0 244500.0 127700.0 243700.0 ;
      RECT  128500.0 244500.0 129300.00000000001 243700.0 ;
      RECT  130100.0 244500.0 130900.0 243700.0 ;
      RECT  130100.0 244500.0 130900.0 243700.0 ;
      RECT  128500.0 244500.0 129300.00000000001 243700.0 ;
      RECT  126900.0 250300.0 127700.0 249500.0 ;
      RECT  128500.0 250300.0 129300.00000000001 249500.0 ;
      RECT  128500.0 250300.0 129300.00000000001 249500.0 ;
      RECT  126900.0 250300.0 127700.0 249500.0 ;
      RECT  128500.0 250300.0 129300.00000000001 249500.0 ;
      RECT  130100.0 250300.0 130900.0 249500.0 ;
      RECT  130100.0 250300.0 130900.0 249500.0 ;
      RECT  128500.0 250300.0 129300.00000000001 249500.0 ;
      RECT  131700.0 244100.00000000003 132500.0 243300.0 ;
      RECT  131700.0 250700.0 132500.0 249900.00000000003 ;
      RECT  130100.0 248600.00000000003 129300.00000000001 247800.0 ;
      RECT  128100.0 247200.0 127300.00000000001 246400.00000000003 ;
      RECT  128500.0 244500.0 129300.00000000001 243700.0 ;
      RECT  130100.0 250300.0 130900.0 249500.0 ;
      RECT  130900.0 247200.0 130100.0 246400.00000000003 ;
      RECT  127300.00000000001 247200.0 128100.0 246400.00000000003 ;
      RECT  129300.00000000001 248600.00000000003 130100.0 247800.0 ;
      RECT  130100.0 247200.0 130900.0 246400.00000000003 ;
      RECT  125700.0 242700.0 135300.0 242100.00000000003 ;
      RECT  125700.0 251900.00000000003 135300.0 251300.0 ;
      RECT  126900.0 252900.00000000003 127700.0 251300.0 ;
      RECT  126900.0 258700.0 127700.0 261100.00000000003 ;
      RECT  130100.0 258700.0 130900.0 261100.00000000003 ;
      RECT  131700.0 259500.0 132500.0 260800.0 ;
      RECT  131700.0 251600.00000000003 132500.0 252900.00000000003 ;
      RECT  126900.0 258700.0 127700.0 259500.0 ;
      RECT  128500.0 258700.0 129300.00000000001 259500.0 ;
      RECT  128500.0 258700.0 129300.00000000001 259500.0 ;
      RECT  126900.0 258700.0 127700.0 259500.0 ;
      RECT  128500.0 258700.0 129300.00000000001 259500.0 ;
      RECT  130100.0 258700.0 130900.0 259500.0 ;
      RECT  130100.0 258700.0 130900.0 259500.0 ;
      RECT  128500.0 258700.0 129300.00000000001 259500.0 ;
      RECT  126900.0 252900.00000000003 127700.0 253700.0 ;
      RECT  128500.0 252900.00000000003 129300.00000000001 253700.0 ;
      RECT  128500.0 252900.00000000003 129300.00000000001 253700.0 ;
      RECT  126900.0 252900.00000000003 127700.0 253700.0 ;
      RECT  128500.0 252900.00000000003 129300.00000000001 253700.0 ;
      RECT  130100.0 252900.00000000003 130900.0 253700.0 ;
      RECT  130100.0 252900.00000000003 130900.0 253700.0 ;
      RECT  128500.0 252900.00000000003 129300.00000000001 253700.0 ;
      RECT  131700.0 259100.00000000003 132500.0 259900.00000000003 ;
      RECT  131700.0 252500.0 132500.0 253300.0 ;
      RECT  130100.0 254600.00000000003 129300.00000000001 255400.00000000003 ;
      RECT  128100.0 256000.0 127300.00000000001 256800.0 ;
      RECT  128500.0 258700.0 129300.00000000001 259500.0 ;
      RECT  130100.0 252900.00000000003 130900.0 253700.0 ;
      RECT  130900.0 256000.0 130100.0 256800.0 ;
      RECT  127300.00000000001 256000.0 128100.0 256800.0 ;
      RECT  129300.00000000001 254600.00000000003 130100.0 255400.00000000003 ;
      RECT  130100.0 256000.0 130900.0 256800.0 ;
      RECT  125700.0 260500.0 135300.0 261100.00000000003 ;
      RECT  125700.0 251300.0 135300.0 251900.00000000003 ;
      RECT  126900.0 268700.0 127700.0 270300.0 ;
      RECT  126900.0 262900.00000000006 127700.0 260500.0 ;
      RECT  130100.0 262900.00000000006 130900.0 260500.0 ;
      RECT  131700.0 262100.00000000003 132500.0 260800.0 ;
      RECT  131700.0 270000.0 132500.0 268700.0 ;
      RECT  126900.0 262900.00000000006 127700.0 262100.00000000003 ;
      RECT  128500.0 262900.00000000006 129300.00000000001 262100.00000000003 ;
      RECT  128500.0 262900.00000000006 129300.00000000001 262100.00000000003 ;
      RECT  126900.0 262900.00000000006 127700.0 262100.00000000003 ;
      RECT  128500.0 262900.00000000006 129300.00000000001 262100.00000000003 ;
      RECT  130100.0 262900.00000000006 130900.0 262100.00000000003 ;
      RECT  130100.0 262900.00000000006 130900.0 262100.00000000003 ;
      RECT  128500.0 262900.00000000006 129300.00000000001 262100.00000000003 ;
      RECT  126900.0 268700.0 127700.0 267900.00000000006 ;
      RECT  128500.0 268700.0 129300.00000000001 267900.00000000006 ;
      RECT  128500.0 268700.0 129300.00000000001 267900.00000000006 ;
      RECT  126900.0 268700.0 127700.0 267900.00000000006 ;
      RECT  128500.0 268700.0 129300.00000000001 267900.00000000006 ;
      RECT  130100.0 268700.0 130900.0 267900.00000000006 ;
      RECT  130100.0 268700.0 130900.0 267900.00000000006 ;
      RECT  128500.0 268700.0 129300.00000000001 267900.00000000006 ;
      RECT  131700.0 262500.0 132500.0 261700.0 ;
      RECT  131700.0 269100.0 132500.0 268300.0 ;
      RECT  130100.0 267000.0 129300.00000000001 266200.0 ;
      RECT  128100.0 265600.0 127300.00000000001 264800.0 ;
      RECT  128500.0 262900.00000000006 129300.00000000001 262100.00000000003 ;
      RECT  130100.0 268700.0 130900.0 267900.00000000006 ;
      RECT  130900.0 265600.0 130100.0 264800.0 ;
      RECT  127300.00000000001 265600.0 128100.0 264800.0 ;
      RECT  129300.00000000001 267000.0 130100.0 266200.0 ;
      RECT  130100.0 265600.0 130900.0 264800.0 ;
      RECT  125700.0 261100.00000000003 135300.0 260500.0 ;
      RECT  125700.0 270300.0 135300.0 269700.0 ;
      RECT  139700.0 130699.99999999999 140500.0 132000.0 ;
      RECT  139700.0 122800.00000000001 140500.0 124100.00000000001 ;
      RECT  136500.0 123700.0 137300.0 122500.0 ;
      RECT  136500.0 129900.0 137300.0 132300.0 ;
      RECT  138300.0 123700.0 138899.99999999997 129900.0 ;
      RECT  136500.0 129900.0 137300.0 130699.99999999999 ;
      RECT  138100.0 129900.0 138899.99999999997 130699.99999999999 ;
      RECT  138100.0 129900.0 138899.99999999997 130699.99999999999 ;
      RECT  136500.0 129900.0 137300.0 130699.99999999999 ;
      RECT  136500.0 123700.0 137300.0 124500.0 ;
      RECT  138100.0 123700.0 138899.99999999997 124500.0 ;
      RECT  138100.0 123700.0 138899.99999999997 124500.0 ;
      RECT  136500.0 123700.0 137300.0 124500.0 ;
      RECT  139700.0 130300.00000000001 140500.0 131100.00000000003 ;
      RECT  139700.0 123700.0 140500.0 124500.0 ;
      RECT  136900.0 126800.00000000001 137700.0 127600.00000000001 ;
      RECT  136900.0 126800.00000000001 137700.0 127600.00000000001 ;
      RECT  138600.0 126900.0 139200.0 127500.0 ;
      RECT  135300.0 131700.0 141700.0 132300.0 ;
      RECT  135300.0 122500.0 141700.0 123100.00000000001 ;
      RECT  139700.0 133300.0 140500.0 132000.0 ;
      RECT  139700.0 141200.0 140500.0 139900.0 ;
      RECT  136500.0 140300.0 137300.0 141500.0 ;
      RECT  136500.0 134100.00000000003 137300.0 131700.0 ;
      RECT  138300.0 140300.0 138899.99999999997 134100.00000000003 ;
      RECT  136500.0 134100.00000000003 137300.0 133300.0 ;
      RECT  138100.0 134100.00000000003 138899.99999999997 133300.0 ;
      RECT  138100.0 134100.00000000003 138899.99999999997 133300.0 ;
      RECT  136500.0 134100.00000000003 137300.0 133300.0 ;
      RECT  136500.0 140300.0 137300.0 139500.0 ;
      RECT  138100.0 140300.0 138899.99999999997 139500.0 ;
      RECT  138100.0 140300.0 138899.99999999997 139500.0 ;
      RECT  136500.0 140300.0 137300.0 139500.0 ;
      RECT  139700.0 133700.0 140500.0 132900.0 ;
      RECT  139700.0 140300.0 140500.0 139500.0 ;
      RECT  136900.0 137200.0 137700.0 136400.0 ;
      RECT  136900.0 137200.0 137700.0 136400.0 ;
      RECT  138600.0 137100.00000000003 139200.0 136500.0 ;
      RECT  135300.0 132300.0 141700.0 131700.0 ;
      RECT  135300.0 141500.0 141700.0 140900.0 ;
      RECT  139700.0 149100.00000000003 140500.0 150400.0 ;
      RECT  139700.0 141200.0 140500.0 142500.0 ;
      RECT  136500.0 142100.00000000003 137300.0 140900.0 ;
      RECT  136500.0 148300.0 137300.0 150700.0 ;
      RECT  138300.0 142100.00000000003 138899.99999999997 148300.0 ;
      RECT  136500.0 148300.0 137300.0 149100.00000000003 ;
      RECT  138100.0 148300.0 138899.99999999997 149100.00000000003 ;
      RECT  138100.0 148300.0 138899.99999999997 149100.00000000003 ;
      RECT  136500.0 148300.0 137300.0 149100.00000000003 ;
      RECT  136500.0 142100.00000000003 137300.0 142900.0 ;
      RECT  138100.0 142100.00000000003 138899.99999999997 142900.0 ;
      RECT  138100.0 142100.00000000003 138899.99999999997 142900.0 ;
      RECT  136500.0 142100.00000000003 137300.0 142900.0 ;
      RECT  139700.0 148700.0 140500.0 149500.0 ;
      RECT  139700.0 142100.00000000003 140500.0 142900.0 ;
      RECT  136900.0 145200.0 137700.0 146000.0 ;
      RECT  136900.0 145200.0 137700.0 146000.0 ;
      RECT  138600.0 145300.0 139200.0 145900.0 ;
      RECT  135300.0 150100.00000000003 141700.0 150700.0 ;
      RECT  135300.0 140900.0 141700.0 141500.0 ;
      RECT  139700.0 151700.0 140500.0 150400.0 ;
      RECT  139700.0 159600.00000000003 140500.0 158300.0 ;
      RECT  136500.0 158700.0 137300.0 159899.99999999997 ;
      RECT  136500.0 152500.0 137300.0 150100.00000000003 ;
      RECT  138300.0 158700.0 138899.99999999997 152500.0 ;
      RECT  136500.0 152500.0 137300.0 151700.0 ;
      RECT  138100.0 152500.0 138899.99999999997 151700.0 ;
      RECT  138100.0 152500.0 138899.99999999997 151700.0 ;
      RECT  136500.0 152500.0 137300.0 151700.0 ;
      RECT  136500.0 158700.0 137300.0 157899.99999999997 ;
      RECT  138100.0 158700.0 138899.99999999997 157899.99999999997 ;
      RECT  138100.0 158700.0 138899.99999999997 157899.99999999997 ;
      RECT  136500.0 158700.0 137300.0 157899.99999999997 ;
      RECT  139700.0 152100.00000000003 140500.0 151300.0 ;
      RECT  139700.0 158700.0 140500.0 157899.99999999997 ;
      RECT  136900.0 155600.00000000003 137700.0 154800.0 ;
      RECT  136900.0 155600.00000000003 137700.0 154800.0 ;
      RECT  138600.0 155500.0 139200.0 154899.99999999997 ;
      RECT  135300.0 150700.0 141700.0 150100.00000000003 ;
      RECT  135300.0 159899.99999999997 141700.0 159300.0 ;
      RECT  139700.0 167500.0 140500.0 168800.0 ;
      RECT  139700.0 159600.00000000003 140500.0 160899.99999999997 ;
      RECT  136500.0 160500.0 137300.0 159300.0 ;
      RECT  136500.0 166700.0 137300.0 169100.00000000003 ;
      RECT  138300.0 160500.0 138899.99999999997 166700.0 ;
      RECT  136500.0 166700.0 137300.0 167500.0 ;
      RECT  138100.0 166700.0 138899.99999999997 167500.0 ;
      RECT  138100.0 166700.0 138899.99999999997 167500.0 ;
      RECT  136500.0 166700.0 137300.0 167500.0 ;
      RECT  136500.0 160500.0 137300.0 161300.0 ;
      RECT  138100.0 160500.0 138899.99999999997 161300.0 ;
      RECT  138100.0 160500.0 138899.99999999997 161300.0 ;
      RECT  136500.0 160500.0 137300.0 161300.0 ;
      RECT  139700.0 167100.00000000003 140500.0 167899.99999999997 ;
      RECT  139700.0 160500.0 140500.0 161300.0 ;
      RECT  136900.0 163600.00000000003 137700.0 164399.99999999997 ;
      RECT  136900.0 163600.00000000003 137700.0 164399.99999999997 ;
      RECT  138600.0 163700.0 139200.0 164300.0 ;
      RECT  135300.0 168500.0 141700.0 169100.00000000003 ;
      RECT  135300.0 159300.0 141700.0 159899.99999999997 ;
      RECT  139700.0 170100.00000000003 140500.0 168800.0 ;
      RECT  139700.0 178000.0 140500.0 176700.0 ;
      RECT  136500.0 177100.00000000003 137300.0 178300.0 ;
      RECT  136500.0 170899.99999999997 137300.0 168500.0 ;
      RECT  138300.0 177100.00000000003 138899.99999999997 170899.99999999997 ;
      RECT  136500.0 170899.99999999997 137300.0 170100.00000000003 ;
      RECT  138100.0 170899.99999999997 138899.99999999997 170100.00000000003 ;
      RECT  138100.0 170899.99999999997 138899.99999999997 170100.00000000003 ;
      RECT  136500.0 170899.99999999997 137300.0 170100.00000000003 ;
      RECT  136500.0 177100.00000000003 137300.0 176300.0 ;
      RECT  138100.0 177100.00000000003 138899.99999999997 176300.0 ;
      RECT  138100.0 177100.00000000003 138899.99999999997 176300.0 ;
      RECT  136500.0 177100.00000000003 137300.0 176300.0 ;
      RECT  139700.0 170500.0 140500.0 169700.0 ;
      RECT  139700.0 177100.00000000003 140500.0 176300.0 ;
      RECT  136900.0 174000.0 137700.0 173200.0 ;
      RECT  136900.0 174000.0 137700.0 173200.0 ;
      RECT  138600.0 173899.99999999997 139200.0 173300.0 ;
      RECT  135300.0 169100.00000000003 141700.0 168500.0 ;
      RECT  135300.0 178300.0 141700.0 177700.0 ;
      RECT  139700.0 185899.99999999997 140500.0 187200.0 ;
      RECT  139700.0 178000.0 140500.0 179300.0 ;
      RECT  136500.0 178899.99999999997 137300.0 177700.0 ;
      RECT  136500.0 185100.00000000003 137300.0 187500.0 ;
      RECT  138300.0 178899.99999999997 138899.99999999997 185100.00000000003 ;
      RECT  136500.0 185100.00000000003 137300.0 185899.99999999997 ;
      RECT  138100.0 185100.00000000003 138899.99999999997 185899.99999999997 ;
      RECT  138100.0 185100.00000000003 138899.99999999997 185899.99999999997 ;
      RECT  136500.0 185100.00000000003 137300.0 185899.99999999997 ;
      RECT  136500.0 178899.99999999997 137300.0 179700.0 ;
      RECT  138100.0 178899.99999999997 138899.99999999997 179700.0 ;
      RECT  138100.0 178899.99999999997 138899.99999999997 179700.0 ;
      RECT  136500.0 178899.99999999997 137300.0 179700.0 ;
      RECT  139700.0 185500.0 140500.0 186300.0 ;
      RECT  139700.0 178899.99999999997 140500.0 179700.0 ;
      RECT  136900.0 182000.0 137700.0 182800.0 ;
      RECT  136900.0 182000.0 137700.0 182800.0 ;
      RECT  138600.0 182100.00000000003 139200.0 182700.0 ;
      RECT  135300.0 186899.99999999997 141700.0 187500.0 ;
      RECT  135300.0 177700.0 141700.0 178300.0 ;
      RECT  139700.0 188500.0 140500.0 187200.0 ;
      RECT  139700.0 196400.00000000003 140500.0 195100.00000000003 ;
      RECT  136500.0 195500.0 137300.0 196700.0 ;
      RECT  136500.0 189300.0 137300.0 186900.00000000003 ;
      RECT  138300.0 195500.0 138899.99999999997 189300.0 ;
      RECT  136500.0 189300.0 137300.0 188500.0 ;
      RECT  138100.0 189300.0 138899.99999999997 188500.0 ;
      RECT  138100.0 189300.0 138899.99999999997 188500.0 ;
      RECT  136500.0 189300.0 137300.0 188500.0 ;
      RECT  136500.0 195500.0 137300.0 194700.0 ;
      RECT  138100.0 195500.0 138899.99999999997 194700.0 ;
      RECT  138100.0 195500.0 138899.99999999997 194700.0 ;
      RECT  136500.0 195500.0 137300.0 194700.0 ;
      RECT  139700.0 188900.00000000003 140500.0 188100.00000000003 ;
      RECT  139700.0 195500.0 140500.0 194700.0 ;
      RECT  136900.0 192400.00000000003 137700.0 191600.00000000003 ;
      RECT  136900.0 192400.00000000003 137700.0 191600.00000000003 ;
      RECT  138600.0 192300.0 139200.0 191700.0 ;
      RECT  135300.0 187500.0 141700.0 186900.00000000003 ;
      RECT  135300.0 196700.0 141700.0 196100.00000000003 ;
      RECT  139700.0 204300.0 140500.0 205600.00000000003 ;
      RECT  139700.0 196400.00000000003 140500.0 197700.0 ;
      RECT  136500.0 197300.0 137300.0 196100.00000000003 ;
      RECT  136500.0 203500.0 137300.0 205900.00000000003 ;
      RECT  138300.0 197300.0 138899.99999999997 203500.0 ;
      RECT  136500.0 203500.0 137300.0 204300.0 ;
      RECT  138100.0 203500.0 138899.99999999997 204300.0 ;
      RECT  138100.0 203500.0 138899.99999999997 204300.0 ;
      RECT  136500.0 203500.0 137300.0 204300.0 ;
      RECT  136500.0 197300.0 137300.0 198100.00000000003 ;
      RECT  138100.0 197300.0 138899.99999999997 198100.00000000003 ;
      RECT  138100.0 197300.0 138899.99999999997 198100.00000000003 ;
      RECT  136500.0 197300.0 137300.0 198100.00000000003 ;
      RECT  139700.0 203900.00000000003 140500.0 204700.0 ;
      RECT  139700.0 197300.0 140500.0 198100.00000000003 ;
      RECT  136900.0 200400.00000000003 137700.0 201200.0 ;
      RECT  136900.0 200400.00000000003 137700.0 201200.0 ;
      RECT  138600.0 200500.0 139200.0 201100.00000000003 ;
      RECT  135300.0 205300.0 141700.0 205900.00000000003 ;
      RECT  135300.0 196100.00000000003 141700.0 196700.0 ;
      RECT  139700.0 206899.99999999997 140500.0 205600.00000000003 ;
      RECT  139700.0 214800.0 140500.0 213500.0 ;
      RECT  136500.0 213899.99999999997 137300.0 215100.00000000003 ;
      RECT  136500.0 207700.0 137300.0 205300.0 ;
      RECT  138300.0 213899.99999999997 138899.99999999997 207700.0 ;
      RECT  136500.0 207700.0 137300.0 206899.99999999997 ;
      RECT  138100.0 207700.0 138899.99999999997 206899.99999999997 ;
      RECT  138100.0 207700.0 138899.99999999997 206899.99999999997 ;
      RECT  136500.0 207700.0 137300.0 206899.99999999997 ;
      RECT  136500.0 213899.99999999997 137300.0 213100.00000000003 ;
      RECT  138100.0 213899.99999999997 138899.99999999997 213100.00000000003 ;
      RECT  138100.0 213899.99999999997 138899.99999999997 213100.00000000003 ;
      RECT  136500.0 213899.99999999997 137300.0 213100.00000000003 ;
      RECT  139700.0 207300.0 140500.0 206500.0 ;
      RECT  139700.0 213899.99999999997 140500.0 213100.00000000003 ;
      RECT  136900.0 210800.0 137700.0 210000.0 ;
      RECT  136900.0 210800.0 137700.0 210000.0 ;
      RECT  138600.0 210700.0 139200.0 210100.00000000003 ;
      RECT  135300.0 205899.99999999997 141700.0 205300.0 ;
      RECT  135300.0 215100.00000000003 141700.0 214500.0 ;
      RECT  139700.0 222700.0 140500.0 224000.0 ;
      RECT  139700.0 214800.0 140500.0 216100.00000000003 ;
      RECT  136500.0 215700.0 137300.0 214500.0 ;
      RECT  136500.0 221899.99999999997 137300.0 224300.0 ;
      RECT  138300.0 215700.0 138899.99999999997 221899.99999999997 ;
      RECT  136500.0 221899.99999999997 137300.0 222700.0 ;
      RECT  138100.0 221899.99999999997 138899.99999999997 222700.0 ;
      RECT  138100.0 221899.99999999997 138899.99999999997 222700.0 ;
      RECT  136500.0 221899.99999999997 137300.0 222700.0 ;
      RECT  136500.0 215700.0 137300.0 216500.0 ;
      RECT  138100.0 215700.0 138899.99999999997 216500.0 ;
      RECT  138100.0 215700.0 138899.99999999997 216500.0 ;
      RECT  136500.0 215700.0 137300.0 216500.0 ;
      RECT  139700.0 222300.0 140500.0 223100.00000000003 ;
      RECT  139700.0 215700.0 140500.0 216500.0 ;
      RECT  136900.0 218800.0 137700.0 219600.00000000003 ;
      RECT  136900.0 218800.0 137700.0 219600.00000000003 ;
      RECT  138600.0 218899.99999999997 139200.0 219500.0 ;
      RECT  135300.0 223700.0 141700.0 224300.0 ;
      RECT  135300.0 214500.0 141700.0 215100.00000000003 ;
      RECT  139700.0 225300.0 140500.0 224000.0 ;
      RECT  139700.0 233200.0 140500.0 231900.00000000003 ;
      RECT  136500.0 232300.0 137300.0 233500.0 ;
      RECT  136500.0 226100.00000000003 137300.0 223700.0 ;
      RECT  138300.0 232300.0 138899.99999999997 226100.00000000003 ;
      RECT  136500.0 226100.00000000003 137300.0 225300.0 ;
      RECT  138100.0 226100.00000000003 138899.99999999997 225300.0 ;
      RECT  138100.0 226100.00000000003 138899.99999999997 225300.0 ;
      RECT  136500.0 226100.00000000003 137300.0 225300.0 ;
      RECT  136500.0 232300.0 137300.0 231500.0 ;
      RECT  138100.0 232300.0 138899.99999999997 231500.0 ;
      RECT  138100.0 232300.0 138899.99999999997 231500.0 ;
      RECT  136500.0 232300.0 137300.0 231500.0 ;
      RECT  139700.0 225700.0 140500.0 224900.00000000003 ;
      RECT  139700.0 232300.0 140500.0 231500.0 ;
      RECT  136900.0 229200.0 137700.0 228400.00000000003 ;
      RECT  136900.0 229200.0 137700.0 228400.00000000003 ;
      RECT  138600.0 229100.00000000003 139200.0 228500.0 ;
      RECT  135300.0 224300.0 141700.0 223700.0 ;
      RECT  135300.0 233500.0 141700.0 232900.00000000003 ;
      RECT  139700.0 241100.00000000003 140500.0 242400.00000000003 ;
      RECT  139700.0 233200.0 140500.0 234500.0 ;
      RECT  136500.0 234100.00000000003 137300.0 232900.00000000003 ;
      RECT  136500.0 240300.0 137300.0 242700.0 ;
      RECT  138300.0 234100.00000000003 138899.99999999997 240300.0 ;
      RECT  136500.0 240300.0 137300.0 241100.00000000003 ;
      RECT  138100.0 240300.0 138899.99999999997 241100.00000000003 ;
      RECT  138100.0 240300.0 138899.99999999997 241100.00000000003 ;
      RECT  136500.0 240300.0 137300.0 241100.00000000003 ;
      RECT  136500.0 234100.00000000003 137300.0 234900.00000000003 ;
      RECT  138100.0 234100.00000000003 138899.99999999997 234900.00000000003 ;
      RECT  138100.0 234100.00000000003 138899.99999999997 234900.00000000003 ;
      RECT  136500.0 234100.00000000003 137300.0 234900.00000000003 ;
      RECT  139700.0 240700.0 140500.0 241500.0 ;
      RECT  139700.0 234100.00000000003 140500.0 234900.00000000003 ;
      RECT  136900.0 237200.0 137700.0 238000.0 ;
      RECT  136900.0 237200.0 137700.0 238000.0 ;
      RECT  138600.0 237300.0 139200.0 237900.00000000003 ;
      RECT  135300.0 242100.00000000003 141700.0 242700.0 ;
      RECT  135300.0 232900.00000000003 141700.0 233500.0 ;
      RECT  139700.0 243700.0 140500.0 242400.00000000003 ;
      RECT  139700.0 251600.00000000003 140500.0 250300.0 ;
      RECT  136500.0 250700.0 137300.0 251900.00000000003 ;
      RECT  136500.0 244500.0 137300.0 242100.00000000003 ;
      RECT  138300.0 250700.0 138899.99999999997 244500.0 ;
      RECT  136500.0 244500.0 137300.0 243700.0 ;
      RECT  138100.0 244500.0 138899.99999999997 243700.0 ;
      RECT  138100.0 244500.0 138899.99999999997 243700.0 ;
      RECT  136500.0 244500.0 137300.0 243700.0 ;
      RECT  136500.0 250700.0 137300.0 249900.00000000003 ;
      RECT  138100.0 250700.0 138899.99999999997 249900.00000000003 ;
      RECT  138100.0 250700.0 138899.99999999997 249900.00000000003 ;
      RECT  136500.0 250700.0 137300.0 249900.00000000003 ;
      RECT  139700.0 244100.00000000003 140500.0 243300.0 ;
      RECT  139700.0 250700.0 140500.0 249900.00000000003 ;
      RECT  136900.0 247600.00000000003 137700.0 246800.0 ;
      RECT  136900.0 247600.00000000003 137700.0 246800.0 ;
      RECT  138600.0 247500.0 139200.0 246900.00000000003 ;
      RECT  135300.0 242700.0 141700.0 242100.00000000003 ;
      RECT  135300.0 251900.00000000003 141700.0 251300.0 ;
      RECT  139700.0 259500.0 140500.0 260800.0 ;
      RECT  139700.0 251600.00000000003 140500.0 252900.00000000003 ;
      RECT  136500.0 252500.0 137300.0 251300.0 ;
      RECT  136500.0 258700.0 137300.0 261100.00000000003 ;
      RECT  138300.0 252500.0 138899.99999999997 258700.0 ;
      RECT  136500.0 258700.0 137300.0 259500.0 ;
      RECT  138100.0 258700.0 138899.99999999997 259500.0 ;
      RECT  138100.0 258700.0 138899.99999999997 259500.0 ;
      RECT  136500.0 258700.0 137300.0 259500.0 ;
      RECT  136500.0 252500.0 137300.0 253300.0 ;
      RECT  138100.0 252500.0 138899.99999999997 253300.0 ;
      RECT  138100.0 252500.0 138899.99999999997 253300.0 ;
      RECT  136500.0 252500.0 137300.0 253300.0 ;
      RECT  139700.0 259100.00000000003 140500.0 259900.00000000003 ;
      RECT  139700.0 252500.0 140500.0 253300.0 ;
      RECT  136900.0 255600.00000000003 137700.0 256400.00000000003 ;
      RECT  136900.0 255600.00000000003 137700.0 256400.00000000003 ;
      RECT  138600.0 255700.0 139200.0 256300.0 ;
      RECT  135300.0 260500.0 141700.0 261100.00000000003 ;
      RECT  135300.0 251300.0 141700.0 251900.00000000003 ;
      RECT  139700.0 262100.00000000003 140500.0 260800.0 ;
      RECT  139700.0 270000.0 140500.0 268700.0 ;
      RECT  136500.0 269100.0 137300.0 270300.0 ;
      RECT  136500.0 262900.00000000006 137300.0 260500.0 ;
      RECT  138300.0 269100.0 138899.99999999997 262900.00000000006 ;
      RECT  136500.0 262900.00000000006 137300.0 262100.00000000003 ;
      RECT  138100.0 262900.00000000006 138899.99999999997 262100.00000000003 ;
      RECT  138100.0 262900.00000000006 138899.99999999997 262100.00000000003 ;
      RECT  136500.0 262900.00000000006 137300.0 262100.00000000003 ;
      RECT  136500.0 269100.0 137300.0 268300.0 ;
      RECT  138100.0 269100.0 138899.99999999997 268300.0 ;
      RECT  138100.0 269100.0 138899.99999999997 268300.0 ;
      RECT  136500.0 269100.0 137300.0 268300.0 ;
      RECT  139700.0 262500.0 140500.0 261700.0 ;
      RECT  139700.0 269100.0 140500.0 268300.0 ;
      RECT  136900.0 266000.0 137700.0 265200.0 ;
      RECT  136900.0 266000.0 137700.0 265200.0 ;
      RECT  138600.0 265900.00000000006 139200.0 265300.0 ;
      RECT  135300.0 261100.00000000003 141700.0 260500.0 ;
      RECT  135300.0 270300.0 141700.0 269700.0 ;
      RECT  112100.0 126800.00000000001 111300.00000000001 127600.00000000001 ;
      RECT  112100.0 136400.0 111300.00000000001 137200.0 ;
      RECT  112100.0 145200.0 111300.00000000001 146000.0 ;
      RECT  112100.0 154800.0 111300.00000000001 155600.00000000003 ;
      RECT  112100.0 163600.00000000003 111300.00000000001 164399.99999999997 ;
      RECT  112100.0 173200.0 111300.00000000001 174000.0 ;
      RECT  112100.0 182000.0 111300.00000000001 182800.0 ;
      RECT  112100.0 191600.00000000003 111300.00000000001 192399.99999999997 ;
      RECT  115500.0 127200.0 114700.0 128000.0 ;
      RECT  121100.0 125800.00000000001 120300.00000000001 126600.00000000001 ;
      RECT  115500.0 136000.0 114700.0 136800.0 ;
      RECT  122500.0 137400.0 121700.0 138200.0 ;
      RECT  115500.0 145600.00000000003 114700.0 146400.0 ;
      RECT  123900.0 144200.0 123100.0 145000.0 ;
      RECT  115500.0 154399.99999999997 114700.0 155200.0 ;
      RECT  125300.0 155800.0 124500.0 156600.00000000003 ;
      RECT  116900.0 164000.0 116100.0 164800.0 ;
      RECT  121100.0 162600.00000000003 120300.00000000001 163399.99999999997 ;
      RECT  116900.0 172800.0 116100.0 173600.00000000003 ;
      RECT  122500.0 174200.0 121700.0 175000.0 ;
      RECT  116900.0 182399.99999999997 116100.0 183200.0 ;
      RECT  123900.0 181000.0 123100.0 181800.0 ;
      RECT  116900.0 191200.0 116100.0 192000.0 ;
      RECT  125300.0 192600.00000000003 124500.0 193399.99999999997 ;
      RECT  118300.0 200800.0 117500.0 201600.00000000003 ;
      RECT  121100.0 199400.00000000003 120300.00000000001 200200.0 ;
      RECT  118300.0 209600.00000000003 117500.0 210400.00000000003 ;
      RECT  122500.0 211000.0 121700.0 211800.0 ;
      RECT  118300.0 219200.0 117500.0 220000.0 ;
      RECT  123900.0 217800.0 123100.0 218600.00000000003 ;
      RECT  118300.0 228000.0 117500.0 228800.0 ;
      RECT  125300.0 229400.00000000003 124500.0 230200.0 ;
      RECT  119700.0 237600.00000000003 118900.0 238400.00000000003 ;
      RECT  121100.0 236200.0 120300.00000000001 237000.0 ;
      RECT  119700.0 246400.00000000003 118900.0 247200.0 ;
      RECT  122500.0 247800.0 121700.0 248600.00000000003 ;
      RECT  119700.0 256000.0 118900.0 256800.0 ;
      RECT  123900.0 254600.00000000003 123100.0 255400.00000000003 ;
      RECT  119700.0 264800.0 118900.0 265600.0 ;
      RECT  125300.0 266200.0 124500.0 267000.0 ;
      RECT  130900.0 131600.00000000003 130100.00000000003 132400.0 ;
      RECT  130900.0 122400.0 130100.00000000003 123200.0 ;
      RECT  130900.0 131600.00000000003 130100.00000000003 132400.0 ;
      RECT  130900.0 140800.0 130100.00000000003 141600.00000000003 ;
      RECT  130900.0 150000.0 130100.00000000003 150800.0 ;
      RECT  130900.0 140800.0 130100.00000000003 141600.00000000003 ;
      RECT  130900.0 150000.0 130100.00000000003 150800.0 ;
      RECT  130900.0 159200.0 130100.00000000003 160000.0 ;
      RECT  130900.0 168399.99999999997 130100.00000000003 169200.0 ;
      RECT  130900.0 159200.0 130100.00000000003 160000.0 ;
      RECT  130900.0 168399.99999999997 130100.00000000003 169200.0 ;
      RECT  130900.0 177600.00000000003 130100.00000000003 178399.99999999997 ;
      RECT  130900.0 186800.0 130100.00000000003 187600.00000000003 ;
      RECT  130900.0 177600.00000000003 130100.00000000003 178399.99999999997 ;
      RECT  130900.0 186800.0 130100.00000000003 187600.00000000003 ;
      RECT  130900.0 196000.0 130100.00000000003 196800.0 ;
      RECT  130900.0 205200.0 130100.00000000003 206000.0 ;
      RECT  130900.0 196000.0 130100.00000000003 196800.0 ;
      RECT  130900.0 205200.0 130100.00000000003 206000.0 ;
      RECT  130900.0 214400.00000000003 130100.00000000003 215200.0 ;
      RECT  130900.0 223600.00000000003 130100.00000000003 224400.00000000003 ;
      RECT  130900.0 214400.00000000003 130100.00000000003 215200.0 ;
      RECT  130900.0 223600.00000000003 130100.00000000003 224400.00000000003 ;
      RECT  130900.0 232800.0 130100.00000000003 233600.00000000003 ;
      RECT  130900.0 242000.0 130100.00000000003 242800.0 ;
      RECT  130900.0 232800.0 130100.00000000003 233600.00000000003 ;
      RECT  130900.0 242000.0 130100.00000000003 242800.0 ;
      RECT  130900.0 251200.0 130100.00000000003 252000.0 ;
      RECT  130900.0 260399.99999999997 130100.00000000003 261200.0 ;
      RECT  130900.0 251200.0 130100.00000000003 252000.0 ;
      RECT  130900.0 260399.99999999997 130100.00000000003 261200.0 ;
      RECT  130900.0 269600.0 130100.00000000003 270400.00000000006 ;
      RECT  138600.00000000003 126900.0 139200.0 127500.0 ;
      RECT  138600.00000000003 136500.0 139200.0 137100.00000000003 ;
      RECT  138600.00000000003 145300.0 139200.0 145900.0 ;
      RECT  138600.00000000003 154899.99999999997 139200.0 155500.0 ;
      RECT  138600.00000000003 163700.0 139200.0 164300.0 ;
      RECT  138600.00000000003 173300.0 139200.0 173899.99999999997 ;
      RECT  138600.00000000003 182100.00000000003 139200.0 182700.0 ;
      RECT  138600.00000000003 191700.0 139200.0 192300.0 ;
      RECT  138600.00000000003 200500.0 139200.0 201100.00000000003 ;
      RECT  138600.00000000003 210100.00000000003 139200.0 210700.0 ;
      RECT  138600.00000000003 218900.00000000003 139200.0 219500.0 ;
      RECT  138600.00000000003 228500.0 139200.0 229100.00000000003 ;
      RECT  138600.00000000003 237300.0 139200.0 237900.00000000003 ;
      RECT  138600.00000000003 246900.00000000003 139200.0 247500.0 ;
      RECT  138600.00000000003 255700.0 139200.0 256300.0 ;
      RECT  138600.00000000003 265300.0 139200.0 265900.0 ;
      RECT  146200.0 126900.0 149899.99999999997 127500.00000000001 ;
      RECT  151600.0 127300.00000000001 152200.0 127900.0 ;
      RECT  151600.0 126900.0 152200.0 127500.00000000001 ;
      RECT  151600.0 127500.0 152200.0 127600.00000000001 ;
      RECT  151899.99999999997 127300.00000000001 156300.0 127900.0 ;
      RECT  156300.0 127300.00000000001 157100.0 127900.0 ;
      RECT  162600.0 127300.00000000001 163200.0 127900.0 ;
      RECT  162600.0 126900.0 163200.0 127500.00000000001 ;
      RECT  159899.99999999997 127300.00000000001 162899.99999999997 127900.0 ;
      RECT  162600.0 127200.0 163200.0 127600.00000000001 ;
      RECT  162899.99999999997 126900.0 165899.99999999997 127500.00000000001 ;
      RECT  146200.0 136500.0 149899.99999999997 137100.00000000003 ;
      RECT  151600.0 136100.00000000003 152200.0 136700.0 ;
      RECT  151600.0 136500.0 152200.0 137100.00000000003 ;
      RECT  151600.0 136400.0 152200.0 137100.00000000003 ;
      RECT  151899.99999999997 136100.00000000003 156300.0 136700.0 ;
      RECT  156300.0 136100.00000000003 157100.0 136700.0 ;
      RECT  162600.0 136100.00000000003 163200.0 136700.0 ;
      RECT  162600.0 136500.0 163200.0 137100.00000000003 ;
      RECT  159899.99999999997 136100.00000000003 162899.99999999997 136700.0 ;
      RECT  162600.0 136400.0 163200.0 136800.0 ;
      RECT  162899.99999999997 136500.0 165899.99999999997 137100.00000000003 ;
      RECT  146200.0 145300.0 149899.99999999997 145900.0 ;
      RECT  151600.0 145700.0 152200.0 146300.0 ;
      RECT  151600.0 145300.0 152200.0 145900.0 ;
      RECT  151600.0 145900.0 152200.0 146000.0 ;
      RECT  151899.99999999997 145700.0 156300.0 146300.0 ;
      RECT  156300.0 145700.0 157100.0 146300.0 ;
      RECT  162600.0 145700.0 163200.0 146300.0 ;
      RECT  162600.0 145300.0 163200.0 145900.0 ;
      RECT  159899.99999999997 145700.0 162899.99999999997 146300.0 ;
      RECT  162600.0 145600.00000000003 163200.0 146000.0 ;
      RECT  162899.99999999997 145300.0 165899.99999999997 145900.0 ;
      RECT  146200.0 154899.99999999997 149899.99999999997 155500.0 ;
      RECT  151600.0 154500.0 152200.0 155100.00000000003 ;
      RECT  151600.0 154899.99999999997 152200.0 155500.0 ;
      RECT  151600.0 154800.0 152200.0 155500.0 ;
      RECT  151899.99999999997 154500.0 156300.0 155100.00000000003 ;
      RECT  156300.0 154500.0 157100.0 155100.00000000003 ;
      RECT  162600.0 154500.0 163200.0 155100.00000000003 ;
      RECT  162600.0 154899.99999999997 163200.0 155500.0 ;
      RECT  159899.99999999997 154500.0 162899.99999999997 155100.00000000003 ;
      RECT  162600.0 154800.0 163200.0 155200.0 ;
      RECT  162899.99999999997 154899.99999999997 165899.99999999997 155500.0 ;
      RECT  146200.0 163700.0 149899.99999999997 164300.0 ;
      RECT  151600.0 164100.00000000003 152200.0 164700.0 ;
      RECT  151600.0 163700.0 152200.0 164300.0 ;
      RECT  151600.0 164300.0 152200.0 164399.99999999997 ;
      RECT  151899.99999999997 164100.00000000003 156300.0 164700.0 ;
      RECT  156300.0 164100.00000000003 157100.0 164700.0 ;
      RECT  162600.0 164100.00000000003 163200.0 164700.0 ;
      RECT  162600.0 163700.0 163200.0 164300.0 ;
      RECT  159899.99999999997 164100.00000000003 162899.99999999997 164700.0 ;
      RECT  162600.0 164000.0 163200.0 164399.99999999997 ;
      RECT  162899.99999999997 163700.0 165899.99999999997 164300.0 ;
      RECT  146200.0 173300.0 149899.99999999997 173899.99999999997 ;
      RECT  151600.0 172899.99999999997 152200.0 173500.0 ;
      RECT  151600.0 173300.0 152200.0 173899.99999999997 ;
      RECT  151600.0 173200.0 152200.0 173900.00000000003 ;
      RECT  151899.99999999997 172899.99999999997 156300.0 173500.0 ;
      RECT  156300.0 172899.99999999997 157100.0 173500.0 ;
      RECT  162600.0 172899.99999999997 163200.0 173500.0 ;
      RECT  162600.0 173300.0 163200.0 173899.99999999997 ;
      RECT  159899.99999999997 172899.99999999997 162899.99999999997 173500.0 ;
      RECT  162600.0 173200.0 163200.0 173600.00000000003 ;
      RECT  162899.99999999997 173300.0 165899.99999999997 173899.99999999997 ;
      RECT  146200.0 182100.00000000003 149899.99999999997 182700.0 ;
      RECT  151600.0 182500.0 152200.0 183100.00000000003 ;
      RECT  151600.0 182100.00000000003 152200.0 182700.0 ;
      RECT  151600.0 182700.0 152200.0 182800.0 ;
      RECT  151899.99999999997 182500.0 156300.0 183100.00000000003 ;
      RECT  156300.0 182500.0 157100.0 183100.00000000003 ;
      RECT  162600.0 182500.0 163200.0 183100.00000000003 ;
      RECT  162600.0 182100.00000000003 163200.0 182700.0 ;
      RECT  159899.99999999997 182500.0 162899.99999999997 183100.00000000003 ;
      RECT  162600.0 182399.99999999997 163200.0 182800.0 ;
      RECT  162899.99999999997 182100.00000000003 165899.99999999997 182700.0 ;
      RECT  146200.0 191700.0 149899.99999999997 192300.0 ;
      RECT  151600.0 191300.0 152200.0 191899.99999999997 ;
      RECT  151600.0 191700.0 152200.0 192300.0 ;
      RECT  151600.0 191600.00000000003 152200.0 192300.0 ;
      RECT  151899.99999999997 191300.0 156300.0 191899.99999999997 ;
      RECT  156300.0 191300.0 157100.0 191899.99999999997 ;
      RECT  162600.0 191300.0 163200.0 191899.99999999997 ;
      RECT  162600.0 191700.0 163200.0 192300.0 ;
      RECT  159899.99999999997 191300.0 162899.99999999997 191899.99999999997 ;
      RECT  162600.0 191600.00000000003 163200.0 192000.0 ;
      RECT  162899.99999999997 191700.0 165899.99999999997 192300.0 ;
      RECT  146200.0 200500.0 149899.99999999997 201100.00000000003 ;
      RECT  151600.0 200900.00000000003 152200.0 201500.0 ;
      RECT  151600.0 200500.0 152200.0 201100.00000000003 ;
      RECT  151600.0 201100.00000000003 152200.0 201200.0 ;
      RECT  151899.99999999997 200900.00000000003 156300.0 201500.0 ;
      RECT  156300.0 200900.00000000003 157100.0 201500.0 ;
      RECT  162600.0 200900.00000000003 163200.0 201500.0 ;
      RECT  162600.0 200500.0 163200.0 201100.00000000003 ;
      RECT  159899.99999999997 200900.00000000003 162899.99999999997 201500.0 ;
      RECT  162600.0 200800.0 163200.0 201200.0 ;
      RECT  162899.99999999997 200500.0 165899.99999999997 201100.00000000003 ;
      RECT  146200.0 210100.00000000003 149899.99999999997 210700.0 ;
      RECT  151600.0 209700.0 152200.0 210300.0 ;
      RECT  151600.0 210100.00000000003 152200.0 210700.0 ;
      RECT  151600.0 210000.0 152200.0 210700.0 ;
      RECT  151899.99999999997 209700.0 156300.0 210300.0 ;
      RECT  156300.0 209700.0 157100.0 210300.0 ;
      RECT  162600.0 209700.0 163200.0 210300.0 ;
      RECT  162600.0 210100.00000000003 163200.0 210700.0 ;
      RECT  159899.99999999997 209700.0 162899.99999999997 210300.0 ;
      RECT  162600.0 210000.0 163200.0 210400.00000000003 ;
      RECT  162899.99999999997 210100.00000000003 165899.99999999997 210700.0 ;
      RECT  146200.0 218900.00000000003 149899.99999999997 219500.0 ;
      RECT  151600.0 219300.0 152200.0 219899.99999999997 ;
      RECT  151600.0 218900.00000000003 152200.0 219500.0 ;
      RECT  151600.0 219500.0 152200.0 219600.00000000003 ;
      RECT  151899.99999999997 219300.0 156300.0 219899.99999999997 ;
      RECT  156300.0 219300.0 157100.0 219899.99999999997 ;
      RECT  162600.0 219300.0 163200.0 219899.99999999997 ;
      RECT  162600.0 218900.00000000003 163200.0 219500.0 ;
      RECT  159899.99999999997 219300.0 162899.99999999997 219899.99999999997 ;
      RECT  162600.0 219200.0 163200.0 219600.00000000003 ;
      RECT  162899.99999999997 218900.00000000003 165899.99999999997 219500.0 ;
      RECT  146200.0 228500.0 149899.99999999997 229100.00000000003 ;
      RECT  151600.0 228100.00000000003 152200.0 228700.0 ;
      RECT  151600.0 228500.0 152200.0 229100.00000000003 ;
      RECT  151600.0 228400.00000000003 152200.0 229100.00000000003 ;
      RECT  151899.99999999997 228100.00000000003 156300.0 228700.0 ;
      RECT  156300.0 228100.00000000003 157100.0 228700.0 ;
      RECT  162600.0 228100.00000000003 163200.0 228700.0 ;
      RECT  162600.0 228500.0 163200.0 229100.00000000003 ;
      RECT  159899.99999999997 228100.00000000003 162899.99999999997 228700.0 ;
      RECT  162600.0 228400.00000000003 163200.0 228800.0 ;
      RECT  162899.99999999997 228500.0 165899.99999999997 229100.00000000003 ;
      RECT  146200.0 237300.0 149899.99999999997 237899.99999999997 ;
      RECT  151600.0 237700.0 152200.0 238300.0 ;
      RECT  151600.0 237300.0 152200.0 237899.99999999997 ;
      RECT  151600.0 237900.00000000003 152200.0 238000.0 ;
      RECT  151899.99999999997 237700.0 156300.0 238300.0 ;
      RECT  156300.0 237700.0 157100.0 238300.0 ;
      RECT  162600.0 237700.0 163200.0 238300.0 ;
      RECT  162600.0 237300.0 163200.0 237899.99999999997 ;
      RECT  159899.99999999997 237700.0 162899.99999999997 238300.0 ;
      RECT  162600.0 237600.00000000003 163200.0 238000.0 ;
      RECT  162899.99999999997 237300.0 165899.99999999997 237899.99999999997 ;
      RECT  146200.0 246900.00000000003 149899.99999999997 247500.0 ;
      RECT  151600.0 246500.0 152200.0 247100.00000000003 ;
      RECT  151600.0 246900.00000000003 152200.0 247500.0 ;
      RECT  151600.0 246800.0 152200.0 247500.0 ;
      RECT  151899.99999999997 246500.0 156300.0 247100.00000000003 ;
      RECT  156300.0 246500.0 157100.0 247100.00000000003 ;
      RECT  162600.0 246500.0 163200.0 247100.00000000003 ;
      RECT  162600.0 246900.00000000003 163200.0 247500.0 ;
      RECT  159899.99999999997 246500.0 162899.99999999997 247100.00000000003 ;
      RECT  162600.0 246800.0 163200.0 247200.0 ;
      RECT  162899.99999999997 246900.00000000003 165899.99999999997 247500.0 ;
      RECT  146200.0 255700.0 149899.99999999997 256300.0 ;
      RECT  151600.0 256100.00000000003 152200.0 256700.0 ;
      RECT  151600.0 255700.0 152200.0 256300.0 ;
      RECT  151600.0 256300.0 152200.0 256399.99999999997 ;
      RECT  151899.99999999997 256100.00000000003 156300.0 256700.0 ;
      RECT  156300.0 256100.00000000003 157100.0 256700.0 ;
      RECT  162600.0 256100.00000000003 163200.0 256700.0 ;
      RECT  162600.0 255700.0 163200.0 256300.0 ;
      RECT  159899.99999999997 256100.00000000003 162899.99999999997 256700.0 ;
      RECT  162600.0 256000.0 163200.0 256400.00000000003 ;
      RECT  162899.99999999997 255700.0 165899.99999999997 256300.0 ;
      RECT  146200.0 265300.0 149899.99999999997 265900.0 ;
      RECT  151600.0 264900.0 152200.0 265500.0 ;
      RECT  151600.0 265300.0 152200.0 265900.0 ;
      RECT  151600.0 265200.0 152200.0 265900.0 ;
      RECT  151899.99999999997 264900.0 156300.0 265500.0 ;
      RECT  156300.0 264900.0 157100.0 265500.0 ;
      RECT  162600.0 264900.0 163200.0 265500.0 ;
      RECT  162600.0 265300.0 163200.0 265900.0 ;
      RECT  159899.99999999997 264900.0 162899.99999999997 265500.0 ;
      RECT  162600.0 265200.0 163200.0 265600.0 ;
      RECT  162899.99999999997 265300.0 165899.99999999997 265900.0 ;
      RECT  152700.0 130699.99999999999 153500.0 132000.0 ;
      RECT  152700.0 122800.00000000001 153500.0 124100.00000000001 ;
      RECT  149500.0 123700.0 150300.0 122500.0 ;
      RECT  149500.0 129900.0 150300.0 132300.0 ;
      RECT  151300.0 123700.0 151899.99999999997 129900.0 ;
      RECT  149500.0 129900.0 150300.0 130699.99999999999 ;
      RECT  151100.0 129900.0 151899.99999999997 130699.99999999999 ;
      RECT  151100.0 129900.0 151899.99999999997 130699.99999999999 ;
      RECT  149500.0 129900.0 150300.0 130699.99999999999 ;
      RECT  149500.0 123700.0 150300.0 124500.0 ;
      RECT  151100.0 123700.0 151899.99999999997 124500.0 ;
      RECT  151100.0 123700.0 151899.99999999997 124500.0 ;
      RECT  149500.0 123700.0 150300.0 124500.0 ;
      RECT  152700.0 130300.00000000001 153500.0 131100.00000000003 ;
      RECT  152700.0 123700.0 153500.0 124500.0 ;
      RECT  149899.99999999997 126800.00000000001 150700.0 127600.00000000001 ;
      RECT  149899.99999999997 126800.00000000001 150700.0 127600.00000000001 ;
      RECT  151600.0 126900.0 152200.0 127500.0 ;
      RECT  148300.0 131700.0 154700.0 132300.0 ;
      RECT  148300.0 122500.0 154700.0 123100.00000000001 ;
      RECT  155899.99999999997 124100.00000000001 156700.0 122500.0 ;
      RECT  155899.99999999997 129900.0 156700.0 132300.0 ;
      RECT  159100.0 129900.0 159899.99999999997 132300.0 ;
      RECT  160700.0 130699.99999999999 161500.0 132000.0 ;
      RECT  160700.0 122800.00000000001 161500.0 124100.00000000001 ;
      RECT  155899.99999999997 129900.0 156700.0 130699.99999999999 ;
      RECT  157500.0 129900.0 158300.0 130699.99999999999 ;
      RECT  157500.0 129900.0 158300.0 130699.99999999999 ;
      RECT  155899.99999999997 129900.0 156700.0 130699.99999999999 ;
      RECT  157500.0 129900.0 158300.0 130699.99999999999 ;
      RECT  159100.0 129900.0 159900.0 130699.99999999999 ;
      RECT  159100.0 129900.0 159899.99999999997 130699.99999999999 ;
      RECT  157500.0 129900.0 158300.0 130699.99999999999 ;
      RECT  155899.99999999997 124100.00000000001 156700.0 124900.0 ;
      RECT  157500.0 124100.00000000001 158300.0 124900.0 ;
      RECT  157500.0 124100.00000000001 158300.0 124900.0 ;
      RECT  155899.99999999997 124100.00000000001 156700.0 124900.0 ;
      RECT  157500.0 124100.00000000001 158300.0 124900.0 ;
      RECT  159100.0 124100.00000000001 159900.0 124900.0 ;
      RECT  159100.0 124100.00000000001 159899.99999999997 124900.0 ;
      RECT  157500.0 124100.00000000001 158300.0 124900.0 ;
      RECT  160700.0 130300.00000000001 161500.0 131100.00000000003 ;
      RECT  160700.0 123700.0 161500.0 124500.0 ;
      RECT  159100.0 125800.00000000001 158300.0 126600.00000000001 ;
      RECT  157100.0 127200.0 156300.0 128000.0 ;
      RECT  157500.0 129900.0 158300.0 130699.99999999999 ;
      RECT  159100.0 124100.00000000001 159899.99999999997 124900.0 ;
      RECT  159899.99999999997 127200.0 159100.0 128000.0 ;
      RECT  156300.0 127200.0 157100.0 128000.0 ;
      RECT  158300.0 125800.00000000001 159100.0 126600.00000000001 ;
      RECT  159100.0 127200.0 159899.99999999997 128000.0 ;
      RECT  154700.0 131700.0 164300.0 132300.0 ;
      RECT  154700.0 122500.0 164300.0 123100.00000000001 ;
      RECT  168700.0 130699.99999999999 169500.0 132000.0 ;
      RECT  168700.0 122800.00000000001 169500.0 124100.00000000001 ;
      RECT  165500.0 123700.0 166300.0 122500.0 ;
      RECT  165500.0 129900.0 166300.0 132300.0 ;
      RECT  167300.0 123700.0 167900.0 129900.0 ;
      RECT  165500.0 129900.0 166300.0 130699.99999999999 ;
      RECT  167100.00000000003 129900.0 167900.0 130699.99999999999 ;
      RECT  167100.00000000003 129900.0 167900.0 130699.99999999999 ;
      RECT  165500.0 129900.0 166300.0 130699.99999999999 ;
      RECT  165500.0 123700.0 166300.0 124500.0 ;
      RECT  167100.00000000003 123700.0 167900.0 124500.0 ;
      RECT  167100.00000000003 123700.0 167900.0 124500.0 ;
      RECT  165500.0 123700.0 166300.0 124500.0 ;
      RECT  168700.0 130300.00000000001 169500.0 131100.00000000003 ;
      RECT  168700.0 123700.0 169500.0 124500.0 ;
      RECT  165900.0 126800.00000000001 166700.0 127600.00000000001 ;
      RECT  165900.0 126800.00000000001 166700.0 127600.00000000001 ;
      RECT  167600.00000000003 126900.0 168200.0 127500.0 ;
      RECT  164300.0 131700.0 170700.0 132300.0 ;
      RECT  164300.0 122500.0 170700.0 123100.00000000001 ;
      RECT  152700.0 133300.0 153500.0 132000.0 ;
      RECT  152700.0 141200.0 153500.0 139900.0 ;
      RECT  149500.0 140300.0 150300.0 141500.0 ;
      RECT  149500.0 134100.00000000003 150300.0 131700.0 ;
      RECT  151300.0 140300.0 151899.99999999997 134100.00000000003 ;
      RECT  149500.0 134100.00000000003 150300.0 133300.0 ;
      RECT  151100.0 134100.00000000003 151899.99999999997 133300.0 ;
      RECT  151100.0 134100.00000000003 151899.99999999997 133300.0 ;
      RECT  149500.0 134100.00000000003 150300.0 133300.0 ;
      RECT  149500.0 140300.0 150300.0 139500.0 ;
      RECT  151100.0 140300.0 151899.99999999997 139500.0 ;
      RECT  151100.0 140300.0 151899.99999999997 139500.0 ;
      RECT  149500.0 140300.0 150300.0 139500.0 ;
      RECT  152700.0 133700.0 153500.0 132900.0 ;
      RECT  152700.0 140300.0 153500.0 139500.0 ;
      RECT  149899.99999999997 137200.0 150700.0 136400.0 ;
      RECT  149899.99999999997 137200.0 150700.0 136400.0 ;
      RECT  151600.0 137100.00000000003 152200.0 136500.0 ;
      RECT  148300.0 132300.0 154700.0 131700.0 ;
      RECT  148300.0 141500.0 154700.0 140900.0 ;
      RECT  155899.99999999997 139900.0 156700.0 141500.0 ;
      RECT  155899.99999999997 134100.00000000003 156700.0 131700.0 ;
      RECT  159100.0 134100.00000000003 159899.99999999997 131700.0 ;
      RECT  160700.0 133300.0 161500.0 132000.0 ;
      RECT  160700.0 141200.0 161500.0 139900.0 ;
      RECT  155899.99999999997 134100.00000000003 156700.0 133300.0 ;
      RECT  157500.0 134100.00000000003 158300.0 133300.0 ;
      RECT  157500.0 134100.00000000003 158300.0 133300.0 ;
      RECT  155899.99999999997 134100.00000000003 156700.0 133300.0 ;
      RECT  157500.0 134100.00000000003 158300.0 133300.0 ;
      RECT  159100.0 134100.00000000003 159900.0 133300.0 ;
      RECT  159100.0 134100.00000000003 159899.99999999997 133300.0 ;
      RECT  157500.0 134100.00000000003 158300.0 133300.0 ;
      RECT  155899.99999999997 139900.0 156700.0 139100.00000000003 ;
      RECT  157500.0 139900.0 158300.0 139100.00000000003 ;
      RECT  157500.0 139900.0 158300.0 139100.00000000003 ;
      RECT  155899.99999999997 139900.0 156700.0 139100.00000000003 ;
      RECT  157500.0 139900.0 158300.0 139100.00000000003 ;
      RECT  159100.0 139900.0 159900.0 139100.00000000003 ;
      RECT  159100.0 139900.0 159899.99999999997 139100.00000000003 ;
      RECT  157500.0 139900.0 158300.0 139100.00000000003 ;
      RECT  160700.0 133700.0 161500.0 132900.0 ;
      RECT  160700.0 140300.0 161500.0 139500.0 ;
      RECT  159100.0 138200.0 158300.0 137400.0 ;
      RECT  157100.0 136800.0 156300.0 136000.0 ;
      RECT  157500.0 134100.00000000003 158300.0 133300.0 ;
      RECT  159100.0 139900.0 159899.99999999997 139100.00000000003 ;
      RECT  159899.99999999997 136800.0 159100.0 136000.0 ;
      RECT  156300.0 136800.0 157100.0 136000.0 ;
      RECT  158300.0 138200.0 159100.0 137400.0 ;
      RECT  159100.0 136800.0 159899.99999999997 136000.0 ;
      RECT  154700.0 132300.0 164300.0 131700.0 ;
      RECT  154700.0 141500.0 164300.0 140900.0 ;
      RECT  168700.0 133300.0 169500.0 132000.0 ;
      RECT  168700.0 141200.0 169500.0 139900.0 ;
      RECT  165500.0 140300.0 166300.0 141500.0 ;
      RECT  165500.0 134100.00000000003 166300.0 131700.0 ;
      RECT  167300.0 140300.0 167900.0 134100.00000000003 ;
      RECT  165500.0 134100.00000000003 166300.0 133300.0 ;
      RECT  167100.00000000003 134100.00000000003 167900.0 133300.0 ;
      RECT  167100.00000000003 134100.00000000003 167900.0 133300.0 ;
      RECT  165500.0 134100.00000000003 166300.0 133300.0 ;
      RECT  165500.0 140300.0 166300.0 139500.0 ;
      RECT  167100.00000000003 140300.0 167900.0 139500.0 ;
      RECT  167100.00000000003 140300.0 167900.0 139500.0 ;
      RECT  165500.0 140300.0 166300.0 139500.0 ;
      RECT  168700.0 133700.0 169500.0 132900.0 ;
      RECT  168700.0 140300.0 169500.0 139500.0 ;
      RECT  165900.0 137200.0 166700.0 136400.0 ;
      RECT  165900.0 137200.0 166700.0 136400.0 ;
      RECT  167600.00000000003 137100.00000000003 168200.0 136500.0 ;
      RECT  164300.0 132300.0 170700.0 131700.0 ;
      RECT  164300.0 141500.0 170700.0 140900.0 ;
      RECT  152700.0 149100.00000000003 153500.0 150400.0 ;
      RECT  152700.0 141200.0 153500.0 142500.0 ;
      RECT  149500.0 142100.00000000003 150300.0 140900.0 ;
      RECT  149500.0 148300.0 150300.0 150700.0 ;
      RECT  151300.0 142100.00000000003 151899.99999999997 148300.0 ;
      RECT  149500.0 148300.0 150300.0 149100.00000000003 ;
      RECT  151100.0 148300.0 151899.99999999997 149100.00000000003 ;
      RECT  151100.0 148300.0 151899.99999999997 149100.00000000003 ;
      RECT  149500.0 148300.0 150300.0 149100.00000000003 ;
      RECT  149500.0 142100.00000000003 150300.0 142900.0 ;
      RECT  151100.0 142100.00000000003 151899.99999999997 142900.0 ;
      RECT  151100.0 142100.00000000003 151899.99999999997 142900.0 ;
      RECT  149500.0 142100.00000000003 150300.0 142900.0 ;
      RECT  152700.0 148700.0 153500.0 149500.0 ;
      RECT  152700.0 142100.00000000003 153500.0 142900.0 ;
      RECT  149899.99999999997 145200.0 150700.0 146000.0 ;
      RECT  149899.99999999997 145200.0 150700.0 146000.0 ;
      RECT  151600.0 145300.0 152200.0 145900.0 ;
      RECT  148300.0 150100.00000000003 154700.0 150700.0 ;
      RECT  148300.0 140900.0 154700.0 141500.0 ;
      RECT  155899.99999999997 142500.0 156700.0 140900.0 ;
      RECT  155899.99999999997 148300.0 156700.0 150700.0 ;
      RECT  159100.0 148300.0 159899.99999999997 150700.0 ;
      RECT  160700.0 149100.00000000003 161500.0 150400.0 ;
      RECT  160700.0 141200.0 161500.0 142500.0 ;
      RECT  155899.99999999997 148300.0 156700.0 149100.00000000003 ;
      RECT  157500.0 148300.0 158300.0 149100.00000000003 ;
      RECT  157500.0 148300.0 158300.0 149100.00000000003 ;
      RECT  155899.99999999997 148300.0 156700.0 149100.00000000003 ;
      RECT  157500.0 148300.0 158300.0 149100.00000000003 ;
      RECT  159100.0 148300.0 159900.0 149100.00000000003 ;
      RECT  159100.0 148300.0 159899.99999999997 149100.00000000003 ;
      RECT  157500.0 148300.0 158300.0 149100.00000000003 ;
      RECT  155899.99999999997 142500.0 156700.0 143300.0 ;
      RECT  157500.0 142500.0 158300.0 143300.0 ;
      RECT  157500.0 142500.0 158300.0 143300.0 ;
      RECT  155899.99999999997 142500.0 156700.0 143300.0 ;
      RECT  157500.0 142500.0 158300.0 143300.0 ;
      RECT  159100.0 142500.0 159900.0 143300.0 ;
      RECT  159100.0 142500.0 159899.99999999997 143300.0 ;
      RECT  157500.0 142500.0 158300.0 143300.0 ;
      RECT  160700.0 148700.0 161500.0 149500.0 ;
      RECT  160700.0 142100.00000000003 161500.0 142900.0 ;
      RECT  159100.0 144200.0 158300.0 145000.0 ;
      RECT  157100.0 145600.00000000003 156300.0 146400.0 ;
      RECT  157500.0 148300.0 158300.0 149100.00000000003 ;
      RECT  159100.0 142500.0 159899.99999999997 143300.0 ;
      RECT  159899.99999999997 145600.00000000003 159100.0 146400.0 ;
      RECT  156300.0 145600.00000000003 157100.0 146400.0 ;
      RECT  158300.0 144200.0 159100.0 145000.0 ;
      RECT  159100.0 145600.00000000003 159899.99999999997 146400.0 ;
      RECT  154700.0 150100.00000000003 164300.0 150700.0 ;
      RECT  154700.0 140900.0 164300.0 141500.0 ;
      RECT  168700.0 149100.00000000003 169500.0 150400.0 ;
      RECT  168700.0 141200.0 169500.0 142500.0 ;
      RECT  165500.0 142100.00000000003 166300.0 140900.0 ;
      RECT  165500.0 148300.0 166300.0 150700.0 ;
      RECT  167300.0 142100.00000000003 167900.0 148300.0 ;
      RECT  165500.0 148300.0 166300.0 149100.00000000003 ;
      RECT  167100.00000000003 148300.0 167900.0 149100.00000000003 ;
      RECT  167100.00000000003 148300.0 167900.0 149100.00000000003 ;
      RECT  165500.0 148300.0 166300.0 149100.00000000003 ;
      RECT  165500.0 142100.00000000003 166300.0 142900.0 ;
      RECT  167100.00000000003 142100.00000000003 167900.0 142900.0 ;
      RECT  167100.00000000003 142100.00000000003 167900.0 142900.0 ;
      RECT  165500.0 142100.00000000003 166300.0 142900.0 ;
      RECT  168700.0 148700.0 169500.0 149500.0 ;
      RECT  168700.0 142100.00000000003 169500.0 142900.0 ;
      RECT  165900.0 145200.0 166700.0 146000.0 ;
      RECT  165900.0 145200.0 166700.0 146000.0 ;
      RECT  167600.00000000003 145300.0 168200.0 145900.0 ;
      RECT  164300.0 150100.00000000003 170700.0 150700.0 ;
      RECT  164300.0 140900.0 170700.0 141500.0 ;
      RECT  152700.0 151700.0 153500.0 150400.0 ;
      RECT  152700.0 159600.00000000003 153500.0 158300.0 ;
      RECT  149500.0 158700.0 150300.0 159899.99999999997 ;
      RECT  149500.0 152500.0 150300.0 150100.00000000003 ;
      RECT  151300.0 158700.0 151899.99999999997 152500.0 ;
      RECT  149500.0 152500.0 150300.0 151700.0 ;
      RECT  151100.0 152500.0 151899.99999999997 151700.0 ;
      RECT  151100.0 152500.0 151899.99999999997 151700.0 ;
      RECT  149500.0 152500.0 150300.0 151700.0 ;
      RECT  149500.0 158700.0 150300.0 157899.99999999997 ;
      RECT  151100.0 158700.0 151899.99999999997 157899.99999999997 ;
      RECT  151100.0 158700.0 151899.99999999997 157899.99999999997 ;
      RECT  149500.0 158700.0 150300.0 157899.99999999997 ;
      RECT  152700.0 152100.00000000003 153500.0 151300.0 ;
      RECT  152700.0 158700.0 153500.0 157899.99999999997 ;
      RECT  149899.99999999997 155600.00000000003 150700.0 154800.0 ;
      RECT  149899.99999999997 155600.00000000003 150700.0 154800.0 ;
      RECT  151600.0 155500.0 152200.0 154899.99999999997 ;
      RECT  148300.0 150700.0 154700.0 150100.00000000003 ;
      RECT  148300.0 159899.99999999997 154700.0 159300.0 ;
      RECT  155899.99999999997 158300.0 156700.0 159899.99999999997 ;
      RECT  155899.99999999997 152500.0 156700.0 150100.00000000003 ;
      RECT  159100.0 152500.0 159899.99999999997 150100.00000000003 ;
      RECT  160700.0 151700.0 161500.0 150400.0 ;
      RECT  160700.0 159600.00000000003 161500.0 158300.0 ;
      RECT  155899.99999999997 152500.0 156700.0 151700.0 ;
      RECT  157500.0 152500.0 158300.0 151700.0 ;
      RECT  157500.0 152500.0 158300.0 151700.0 ;
      RECT  155899.99999999997 152500.0 156700.0 151700.0 ;
      RECT  157500.0 152500.0 158300.0 151700.0 ;
      RECT  159100.0 152500.0 159900.0 151700.0 ;
      RECT  159100.0 152500.0 159899.99999999997 151700.0 ;
      RECT  157500.0 152500.0 158300.0 151700.0 ;
      RECT  155899.99999999997 158300.0 156700.0 157500.0 ;
      RECT  157500.0 158300.0 158300.0 157500.0 ;
      RECT  157500.0 158300.0 158300.0 157500.0 ;
      RECT  155899.99999999997 158300.0 156700.0 157500.0 ;
      RECT  157500.0 158300.0 158300.0 157500.0 ;
      RECT  159100.0 158300.0 159900.0 157500.0 ;
      RECT  159100.0 158300.0 159899.99999999997 157500.0 ;
      RECT  157500.0 158300.0 158300.0 157500.0 ;
      RECT  160700.0 152100.00000000003 161500.0 151300.0 ;
      RECT  160700.0 158700.0 161500.0 157899.99999999997 ;
      RECT  159100.0 156600.00000000003 158300.0 155800.0 ;
      RECT  157100.0 155200.0 156300.0 154399.99999999997 ;
      RECT  157500.0 152500.0 158300.0 151700.0 ;
      RECT  159100.0 158300.0 159899.99999999997 157500.0 ;
      RECT  159899.99999999997 155200.0 159100.0 154399.99999999997 ;
      RECT  156300.0 155200.0 157100.0 154399.99999999997 ;
      RECT  158300.0 156600.00000000003 159100.0 155800.0 ;
      RECT  159100.0 155200.0 159899.99999999997 154399.99999999997 ;
      RECT  154700.0 150700.0 164300.0 150100.00000000003 ;
      RECT  154700.0 159899.99999999997 164300.0 159300.0 ;
      RECT  168700.0 151700.0 169500.0 150400.0 ;
      RECT  168700.0 159600.00000000003 169500.0 158300.0 ;
      RECT  165500.0 158700.0 166300.0 159899.99999999997 ;
      RECT  165500.0 152500.0 166300.0 150100.00000000003 ;
      RECT  167300.0 158700.0 167900.0 152500.0 ;
      RECT  165500.0 152500.0 166300.0 151700.0 ;
      RECT  167100.00000000003 152500.0 167900.0 151700.0 ;
      RECT  167100.00000000003 152500.0 167900.0 151700.0 ;
      RECT  165500.0 152500.0 166300.0 151700.0 ;
      RECT  165500.0 158700.0 166300.0 157899.99999999997 ;
      RECT  167100.00000000003 158700.0 167900.0 157899.99999999997 ;
      RECT  167100.00000000003 158700.0 167900.0 157899.99999999997 ;
      RECT  165500.0 158700.0 166300.0 157899.99999999997 ;
      RECT  168700.0 152100.00000000003 169500.0 151300.0 ;
      RECT  168700.0 158700.0 169500.0 157899.99999999997 ;
      RECT  165900.0 155600.00000000003 166700.0 154800.0 ;
      RECT  165900.0 155600.00000000003 166700.0 154800.0 ;
      RECT  167600.00000000003 155500.0 168200.0 154899.99999999997 ;
      RECT  164300.0 150700.0 170700.0 150100.00000000003 ;
      RECT  164300.0 159899.99999999997 170700.0 159300.0 ;
      RECT  152700.0 167500.0 153500.0 168800.0 ;
      RECT  152700.0 159600.00000000003 153500.0 160899.99999999997 ;
      RECT  149500.0 160500.0 150300.0 159300.0 ;
      RECT  149500.0 166700.0 150300.0 169100.00000000003 ;
      RECT  151300.0 160500.0 151899.99999999997 166700.0 ;
      RECT  149500.0 166700.0 150300.0 167500.0 ;
      RECT  151100.0 166700.0 151899.99999999997 167500.0 ;
      RECT  151100.0 166700.0 151899.99999999997 167500.0 ;
      RECT  149500.0 166700.0 150300.0 167500.0 ;
      RECT  149500.0 160500.0 150300.0 161300.0 ;
      RECT  151100.0 160500.0 151899.99999999997 161300.0 ;
      RECT  151100.0 160500.0 151899.99999999997 161300.0 ;
      RECT  149500.0 160500.0 150300.0 161300.0 ;
      RECT  152700.0 167100.00000000003 153500.0 167899.99999999997 ;
      RECT  152700.0 160500.0 153500.0 161300.0 ;
      RECT  149899.99999999997 163600.00000000003 150700.0 164399.99999999997 ;
      RECT  149899.99999999997 163600.00000000003 150700.0 164399.99999999997 ;
      RECT  151600.0 163700.0 152200.0 164300.0 ;
      RECT  148300.0 168500.0 154700.0 169100.00000000003 ;
      RECT  148300.0 159300.0 154700.0 159899.99999999997 ;
      RECT  155899.99999999997 160899.99999999997 156700.0 159300.0 ;
      RECT  155899.99999999997 166700.0 156700.0 169100.00000000003 ;
      RECT  159100.0 166700.0 159899.99999999997 169100.00000000003 ;
      RECT  160700.0 167500.0 161500.0 168800.0 ;
      RECT  160700.0 159600.00000000003 161500.0 160899.99999999997 ;
      RECT  155899.99999999997 166700.0 156700.0 167500.0 ;
      RECT  157500.0 166700.0 158300.0 167500.0 ;
      RECT  157500.0 166700.0 158300.0 167500.0 ;
      RECT  155899.99999999997 166700.0 156700.0 167500.0 ;
      RECT  157500.0 166700.0 158300.0 167500.0 ;
      RECT  159100.0 166700.0 159900.0 167500.0 ;
      RECT  159100.0 166700.0 159899.99999999997 167500.0 ;
      RECT  157500.0 166700.0 158300.0 167500.0 ;
      RECT  155899.99999999997 160899.99999999997 156700.0 161700.0 ;
      RECT  157500.0 160899.99999999997 158300.0 161700.0 ;
      RECT  157500.0 160899.99999999997 158300.0 161700.0 ;
      RECT  155899.99999999997 160899.99999999997 156700.0 161700.0 ;
      RECT  157500.0 160899.99999999997 158300.0 161700.0 ;
      RECT  159100.0 160899.99999999997 159900.0 161700.0 ;
      RECT  159100.0 160899.99999999997 159899.99999999997 161700.0 ;
      RECT  157500.0 160899.99999999997 158300.0 161700.0 ;
      RECT  160700.0 167100.00000000003 161500.0 167899.99999999997 ;
      RECT  160700.0 160500.0 161500.0 161300.0 ;
      RECT  159100.0 162600.00000000003 158300.0 163399.99999999997 ;
      RECT  157100.0 164000.0 156300.0 164800.0 ;
      RECT  157500.0 166700.0 158300.0 167500.0 ;
      RECT  159100.0 160899.99999999997 159899.99999999997 161700.0 ;
      RECT  159899.99999999997 164000.0 159100.0 164800.0 ;
      RECT  156300.0 164000.0 157100.0 164800.0 ;
      RECT  158300.0 162600.00000000003 159100.0 163399.99999999997 ;
      RECT  159100.0 164000.0 159899.99999999997 164800.0 ;
      RECT  154700.0 168500.0 164300.0 169100.00000000003 ;
      RECT  154700.0 159300.0 164300.0 159899.99999999997 ;
      RECT  168700.0 167500.0 169500.0 168800.0 ;
      RECT  168700.0 159600.00000000003 169500.0 160899.99999999997 ;
      RECT  165500.0 160500.0 166300.0 159300.0 ;
      RECT  165500.0 166700.0 166300.0 169100.00000000003 ;
      RECT  167300.0 160500.0 167900.0 166700.0 ;
      RECT  165500.0 166700.0 166300.0 167500.0 ;
      RECT  167100.00000000003 166700.0 167900.0 167500.0 ;
      RECT  167100.00000000003 166700.0 167900.0 167500.0 ;
      RECT  165500.0 166700.0 166300.0 167500.0 ;
      RECT  165500.0 160500.0 166300.0 161300.0 ;
      RECT  167100.00000000003 160500.0 167900.0 161300.0 ;
      RECT  167100.00000000003 160500.0 167900.0 161300.0 ;
      RECT  165500.0 160500.0 166300.0 161300.0 ;
      RECT  168700.0 167100.00000000003 169500.0 167899.99999999997 ;
      RECT  168700.0 160500.0 169500.0 161300.0 ;
      RECT  165900.0 163600.00000000003 166700.0 164399.99999999997 ;
      RECT  165900.0 163600.00000000003 166700.0 164399.99999999997 ;
      RECT  167600.00000000003 163700.0 168200.0 164300.0 ;
      RECT  164300.0 168500.0 170700.0 169100.00000000003 ;
      RECT  164300.0 159300.0 170700.0 159899.99999999997 ;
      RECT  152700.0 170100.00000000003 153500.0 168800.0 ;
      RECT  152700.0 178000.0 153500.0 176700.0 ;
      RECT  149500.0 177100.00000000003 150300.0 178300.0 ;
      RECT  149500.0 170899.99999999997 150300.0 168500.0 ;
      RECT  151300.0 177100.00000000003 151899.99999999997 170899.99999999997 ;
      RECT  149500.0 170899.99999999997 150300.0 170100.00000000003 ;
      RECT  151100.0 170899.99999999997 151899.99999999997 170100.00000000003 ;
      RECT  151100.0 170899.99999999997 151899.99999999997 170100.00000000003 ;
      RECT  149500.0 170899.99999999997 150300.0 170100.00000000003 ;
      RECT  149500.0 177100.00000000003 150300.0 176300.0 ;
      RECT  151100.0 177100.00000000003 151899.99999999997 176300.0 ;
      RECT  151100.0 177100.00000000003 151899.99999999997 176300.0 ;
      RECT  149500.0 177100.00000000003 150300.0 176300.0 ;
      RECT  152700.0 170500.0 153500.0 169700.0 ;
      RECT  152700.0 177100.00000000003 153500.0 176300.0 ;
      RECT  149899.99999999997 174000.0 150700.0 173200.0 ;
      RECT  149899.99999999997 174000.0 150700.0 173200.0 ;
      RECT  151600.0 173899.99999999997 152200.0 173300.0 ;
      RECT  148300.0 169100.00000000003 154700.0 168500.0 ;
      RECT  148300.0 178300.0 154700.0 177700.0 ;
      RECT  155899.99999999997 176700.0 156700.0 178300.0 ;
      RECT  155899.99999999997 170899.99999999997 156700.0 168500.0 ;
      RECT  159100.0 170899.99999999997 159899.99999999997 168500.0 ;
      RECT  160700.0 170100.00000000003 161500.0 168800.0 ;
      RECT  160700.0 178000.0 161500.0 176700.0 ;
      RECT  155899.99999999997 170899.99999999997 156700.0 170100.00000000003 ;
      RECT  157500.0 170899.99999999997 158300.0 170100.00000000003 ;
      RECT  157500.0 170899.99999999997 158300.0 170100.00000000003 ;
      RECT  155899.99999999997 170899.99999999997 156700.0 170100.00000000003 ;
      RECT  157500.0 170899.99999999997 158300.0 170100.00000000003 ;
      RECT  159100.0 170899.99999999997 159900.0 170100.00000000003 ;
      RECT  159100.0 170899.99999999997 159899.99999999997 170100.00000000003 ;
      RECT  157500.0 170899.99999999997 158300.0 170100.00000000003 ;
      RECT  155899.99999999997 176700.0 156700.0 175899.99999999997 ;
      RECT  157500.0 176700.0 158300.0 175899.99999999997 ;
      RECT  157500.0 176700.0 158300.0 175899.99999999997 ;
      RECT  155899.99999999997 176700.0 156700.0 175899.99999999997 ;
      RECT  157500.0 176700.0 158300.0 175899.99999999997 ;
      RECT  159100.0 176700.0 159900.0 175899.99999999997 ;
      RECT  159100.0 176700.0 159899.99999999997 175899.99999999997 ;
      RECT  157500.0 176700.0 158300.0 175899.99999999997 ;
      RECT  160700.0 170500.0 161500.0 169700.0 ;
      RECT  160700.0 177100.00000000003 161500.0 176300.0 ;
      RECT  159100.0 175000.0 158300.0 174200.0 ;
      RECT  157100.0 173600.00000000003 156300.0 172800.0 ;
      RECT  157500.0 170899.99999999997 158300.0 170100.00000000003 ;
      RECT  159100.0 176700.0 159899.99999999997 175899.99999999997 ;
      RECT  159899.99999999997 173600.00000000003 159100.0 172800.0 ;
      RECT  156300.0 173600.00000000003 157100.0 172800.0 ;
      RECT  158300.0 175000.0 159100.0 174200.0 ;
      RECT  159100.0 173600.00000000003 159899.99999999997 172800.0 ;
      RECT  154700.0 169100.00000000003 164300.0 168500.0 ;
      RECT  154700.0 178300.0 164300.0 177700.0 ;
      RECT  168700.0 170100.00000000003 169500.0 168800.0 ;
      RECT  168700.0 178000.0 169500.0 176700.0 ;
      RECT  165500.0 177100.00000000003 166300.0 178300.0 ;
      RECT  165500.0 170899.99999999997 166300.0 168500.0 ;
      RECT  167300.0 177100.00000000003 167900.0 170899.99999999997 ;
      RECT  165500.0 170899.99999999997 166300.0 170100.00000000003 ;
      RECT  167100.00000000003 170899.99999999997 167900.0 170100.00000000003 ;
      RECT  167100.00000000003 170899.99999999997 167900.0 170100.00000000003 ;
      RECT  165500.0 170899.99999999997 166300.0 170100.00000000003 ;
      RECT  165500.0 177100.00000000003 166300.0 176300.0 ;
      RECT  167100.00000000003 177100.00000000003 167900.0 176300.0 ;
      RECT  167100.00000000003 177100.00000000003 167900.0 176300.0 ;
      RECT  165500.0 177100.00000000003 166300.0 176300.0 ;
      RECT  168700.0 170500.0 169500.0 169700.0 ;
      RECT  168700.0 177100.00000000003 169500.0 176300.0 ;
      RECT  165900.0 174000.0 166700.0 173200.0 ;
      RECT  165900.0 174000.0 166700.0 173200.0 ;
      RECT  167600.00000000003 173899.99999999997 168200.0 173300.0 ;
      RECT  164300.0 169100.00000000003 170700.0 168500.0 ;
      RECT  164300.0 178300.0 170700.0 177700.0 ;
      RECT  152700.0 185899.99999999997 153500.0 187200.0 ;
      RECT  152700.0 178000.0 153500.0 179300.0 ;
      RECT  149500.0 178899.99999999997 150300.0 177700.0 ;
      RECT  149500.0 185100.00000000003 150300.0 187500.0 ;
      RECT  151300.0 178899.99999999997 151899.99999999997 185100.00000000003 ;
      RECT  149500.0 185100.00000000003 150300.0 185899.99999999997 ;
      RECT  151100.0 185100.00000000003 151899.99999999997 185899.99999999997 ;
      RECT  151100.0 185100.00000000003 151899.99999999997 185899.99999999997 ;
      RECT  149500.0 185100.00000000003 150300.0 185899.99999999997 ;
      RECT  149500.0 178899.99999999997 150300.0 179700.0 ;
      RECT  151100.0 178899.99999999997 151899.99999999997 179700.0 ;
      RECT  151100.0 178899.99999999997 151899.99999999997 179700.0 ;
      RECT  149500.0 178899.99999999997 150300.0 179700.0 ;
      RECT  152700.0 185500.0 153500.0 186300.0 ;
      RECT  152700.0 178899.99999999997 153500.0 179700.0 ;
      RECT  149899.99999999997 182000.0 150700.0 182800.0 ;
      RECT  149899.99999999997 182000.0 150700.0 182800.0 ;
      RECT  151600.0 182100.00000000003 152200.0 182700.0 ;
      RECT  148300.0 186899.99999999997 154700.0 187500.0 ;
      RECT  148300.0 177700.0 154700.0 178300.0 ;
      RECT  155899.99999999997 179300.0 156700.0 177700.0 ;
      RECT  155899.99999999997 185100.00000000003 156700.0 187500.0 ;
      RECT  159100.0 185100.00000000003 159899.99999999997 187500.0 ;
      RECT  160700.0 185899.99999999997 161500.0 187200.0 ;
      RECT  160700.0 178000.0 161500.0 179300.0 ;
      RECT  155899.99999999997 185100.00000000003 156700.0 185899.99999999997 ;
      RECT  157500.0 185100.00000000003 158300.0 185899.99999999997 ;
      RECT  157500.0 185100.00000000003 158300.0 185899.99999999997 ;
      RECT  155899.99999999997 185100.00000000003 156700.0 185899.99999999997 ;
      RECT  157500.0 185100.00000000003 158300.0 185899.99999999997 ;
      RECT  159100.0 185100.00000000003 159900.0 185899.99999999997 ;
      RECT  159100.0 185100.00000000003 159899.99999999997 185899.99999999997 ;
      RECT  157500.0 185100.00000000003 158300.0 185899.99999999997 ;
      RECT  155899.99999999997 179300.0 156700.0 180100.00000000003 ;
      RECT  157500.0 179300.0 158300.0 180100.00000000003 ;
      RECT  157500.0 179300.0 158300.0 180100.00000000003 ;
      RECT  155899.99999999997 179300.0 156700.0 180100.00000000003 ;
      RECT  157500.0 179300.0 158300.0 180100.00000000003 ;
      RECT  159100.0 179300.0 159900.0 180100.00000000003 ;
      RECT  159100.0 179300.0 159899.99999999997 180100.00000000003 ;
      RECT  157500.0 179300.0 158300.0 180100.00000000003 ;
      RECT  160700.0 185500.0 161500.0 186300.0 ;
      RECT  160700.0 178899.99999999997 161500.0 179700.0 ;
      RECT  159100.0 181000.0 158300.0 181800.0 ;
      RECT  157100.0 182399.99999999997 156300.0 183200.0 ;
      RECT  157500.0 185100.00000000003 158300.0 185899.99999999997 ;
      RECT  159100.0 179300.0 159899.99999999997 180100.00000000003 ;
      RECT  159899.99999999997 182399.99999999997 159100.0 183200.0 ;
      RECT  156300.0 182399.99999999997 157100.0 183200.0 ;
      RECT  158300.0 181000.0 159100.0 181800.0 ;
      RECT  159100.0 182399.99999999997 159899.99999999997 183200.0 ;
      RECT  154700.0 186899.99999999997 164300.0 187500.0 ;
      RECT  154700.0 177700.0 164300.0 178300.0 ;
      RECT  168700.0 185899.99999999997 169500.0 187200.0 ;
      RECT  168700.0 178000.0 169500.0 179300.0 ;
      RECT  165500.0 178899.99999999997 166300.0 177700.0 ;
      RECT  165500.0 185100.00000000003 166300.0 187500.0 ;
      RECT  167300.0 178899.99999999997 167900.0 185100.00000000003 ;
      RECT  165500.0 185100.00000000003 166300.0 185899.99999999997 ;
      RECT  167100.00000000003 185100.00000000003 167900.0 185899.99999999997 ;
      RECT  167100.00000000003 185100.00000000003 167900.0 185899.99999999997 ;
      RECT  165500.0 185100.00000000003 166300.0 185899.99999999997 ;
      RECT  165500.0 178899.99999999997 166300.0 179700.0 ;
      RECT  167100.00000000003 178899.99999999997 167900.0 179700.0 ;
      RECT  167100.00000000003 178899.99999999997 167900.0 179700.0 ;
      RECT  165500.0 178899.99999999997 166300.0 179700.0 ;
      RECT  168700.0 185500.0 169500.0 186300.0 ;
      RECT  168700.0 178899.99999999997 169500.0 179700.0 ;
      RECT  165900.0 182000.0 166700.0 182800.0 ;
      RECT  165900.0 182000.0 166700.0 182800.0 ;
      RECT  167600.00000000003 182100.00000000003 168200.0 182700.0 ;
      RECT  164300.0 186899.99999999997 170700.0 187500.0 ;
      RECT  164300.0 177700.0 170700.0 178300.0 ;
      RECT  152700.0 188500.0 153500.0 187200.0 ;
      RECT  152700.0 196400.00000000003 153500.0 195100.00000000003 ;
      RECT  149500.0 195500.0 150300.0 196700.0 ;
      RECT  149500.0 189300.0 150300.0 186900.00000000003 ;
      RECT  151300.0 195500.0 151899.99999999997 189300.0 ;
      RECT  149500.0 189300.0 150300.0 188500.0 ;
      RECT  151100.0 189300.0 151899.99999999997 188500.0 ;
      RECT  151100.0 189300.0 151899.99999999997 188500.0 ;
      RECT  149500.0 189300.0 150300.0 188500.0 ;
      RECT  149500.0 195500.0 150300.0 194700.0 ;
      RECT  151100.0 195500.0 151899.99999999997 194700.0 ;
      RECT  151100.0 195500.0 151899.99999999997 194700.0 ;
      RECT  149500.0 195500.0 150300.0 194700.0 ;
      RECT  152700.0 188900.00000000003 153500.0 188100.00000000003 ;
      RECT  152700.0 195500.0 153500.0 194700.0 ;
      RECT  149899.99999999997 192400.00000000003 150700.0 191600.00000000003 ;
      RECT  149899.99999999997 192400.00000000003 150700.0 191600.00000000003 ;
      RECT  151600.0 192300.0 152200.0 191700.0 ;
      RECT  148300.0 187500.0 154700.0 186900.00000000003 ;
      RECT  148300.0 196700.0 154700.0 196100.00000000003 ;
      RECT  155899.99999999997 195100.00000000003 156700.0 196700.0 ;
      RECT  155899.99999999997 189300.0 156700.0 186900.00000000003 ;
      RECT  159100.0 189300.0 159899.99999999997 186900.00000000003 ;
      RECT  160700.0 188500.0 161500.0 187200.0 ;
      RECT  160700.0 196400.00000000003 161500.0 195100.00000000003 ;
      RECT  155899.99999999997 189300.0 156700.0 188500.0 ;
      RECT  157500.0 189300.0 158300.0 188500.0 ;
      RECT  157500.0 189300.0 158300.0 188500.0 ;
      RECT  155899.99999999997 189300.0 156700.0 188500.0 ;
      RECT  157500.0 189300.0 158300.0 188500.0 ;
      RECT  159100.0 189300.0 159900.0 188500.0 ;
      RECT  159100.0 189300.0 159899.99999999997 188500.0 ;
      RECT  157500.0 189300.0 158300.0 188500.0 ;
      RECT  155899.99999999997 195100.00000000003 156700.0 194300.0 ;
      RECT  157500.0 195100.00000000003 158300.0 194300.0 ;
      RECT  157500.0 195100.00000000003 158300.0 194300.0 ;
      RECT  155899.99999999997 195100.00000000003 156700.0 194300.0 ;
      RECT  157500.0 195100.00000000003 158300.0 194300.0 ;
      RECT  159100.0 195100.00000000003 159900.0 194300.0 ;
      RECT  159100.0 195100.00000000003 159899.99999999997 194300.0 ;
      RECT  157500.0 195100.00000000003 158300.0 194300.0 ;
      RECT  160700.0 188900.00000000003 161500.0 188100.00000000003 ;
      RECT  160700.0 195500.0 161500.0 194700.0 ;
      RECT  159100.0 193400.00000000003 158300.0 192600.00000000003 ;
      RECT  157100.0 192000.0 156300.0 191200.0 ;
      RECT  157500.0 189300.0 158300.0 188500.0 ;
      RECT  159100.0 195100.00000000003 159899.99999999997 194300.0 ;
      RECT  159899.99999999997 192000.0 159100.0 191200.0 ;
      RECT  156300.0 192000.0 157100.0 191200.0 ;
      RECT  158300.0 193400.00000000003 159100.0 192600.00000000003 ;
      RECT  159100.0 192000.0 159899.99999999997 191200.0 ;
      RECT  154700.0 187500.0 164300.0 186900.00000000003 ;
      RECT  154700.0 196700.0 164300.0 196100.00000000003 ;
      RECT  168700.0 188500.0 169500.0 187200.0 ;
      RECT  168700.0 196400.00000000003 169500.0 195100.00000000003 ;
      RECT  165500.0 195500.0 166300.0 196700.0 ;
      RECT  165500.0 189300.0 166300.0 186900.00000000003 ;
      RECT  167300.0 195500.0 167900.0 189300.0 ;
      RECT  165500.0 189300.0 166300.0 188500.0 ;
      RECT  167100.00000000003 189300.0 167900.0 188500.0 ;
      RECT  167100.00000000003 189300.0 167900.0 188500.0 ;
      RECT  165500.0 189300.0 166300.0 188500.0 ;
      RECT  165500.0 195500.0 166300.0 194700.0 ;
      RECT  167100.00000000003 195500.0 167900.0 194700.0 ;
      RECT  167100.00000000003 195500.0 167900.0 194700.0 ;
      RECT  165500.0 195500.0 166300.0 194700.0 ;
      RECT  168700.0 188900.00000000003 169500.0 188100.00000000003 ;
      RECT  168700.0 195500.0 169500.0 194700.0 ;
      RECT  165900.0 192400.00000000003 166700.0 191600.00000000003 ;
      RECT  165900.0 192400.00000000003 166700.0 191600.00000000003 ;
      RECT  167600.00000000003 192300.0 168200.0 191700.0 ;
      RECT  164300.0 187500.0 170700.0 186900.00000000003 ;
      RECT  164300.0 196700.0 170700.0 196100.00000000003 ;
      RECT  152700.0 204300.0 153500.0 205600.00000000003 ;
      RECT  152700.0 196400.00000000003 153500.0 197700.0 ;
      RECT  149500.0 197300.0 150300.0 196100.00000000003 ;
      RECT  149500.0 203500.0 150300.0 205900.00000000003 ;
      RECT  151300.0 197300.0 151899.99999999997 203500.0 ;
      RECT  149500.0 203500.0 150300.0 204300.0 ;
      RECT  151100.0 203500.0 151899.99999999997 204300.0 ;
      RECT  151100.0 203500.0 151899.99999999997 204300.0 ;
      RECT  149500.0 203500.0 150300.0 204300.0 ;
      RECT  149500.0 197300.0 150300.0 198100.00000000003 ;
      RECT  151100.0 197300.0 151899.99999999997 198100.00000000003 ;
      RECT  151100.0 197300.0 151899.99999999997 198100.00000000003 ;
      RECT  149500.0 197300.0 150300.0 198100.00000000003 ;
      RECT  152700.0 203900.00000000003 153500.0 204700.0 ;
      RECT  152700.0 197300.0 153500.0 198100.00000000003 ;
      RECT  149899.99999999997 200400.00000000003 150700.0 201200.0 ;
      RECT  149899.99999999997 200400.00000000003 150700.0 201200.0 ;
      RECT  151600.0 200500.0 152200.0 201100.00000000003 ;
      RECT  148300.0 205300.0 154700.0 205900.00000000003 ;
      RECT  148300.0 196100.00000000003 154700.0 196700.0 ;
      RECT  155899.99999999997 197700.0 156700.0 196100.00000000003 ;
      RECT  155899.99999999997 203500.0 156700.0 205900.00000000003 ;
      RECT  159100.0 203500.0 159899.99999999997 205900.00000000003 ;
      RECT  160700.0 204300.0 161500.0 205600.00000000003 ;
      RECT  160700.0 196400.00000000003 161500.0 197700.0 ;
      RECT  155899.99999999997 203500.0 156700.0 204300.0 ;
      RECT  157500.0 203500.0 158300.0 204300.0 ;
      RECT  157500.0 203500.0 158300.0 204300.0 ;
      RECT  155899.99999999997 203500.0 156700.0 204300.0 ;
      RECT  157500.0 203500.0 158300.0 204300.0 ;
      RECT  159100.0 203500.0 159900.0 204300.0 ;
      RECT  159100.0 203500.0 159899.99999999997 204300.0 ;
      RECT  157500.0 203500.0 158300.0 204300.0 ;
      RECT  155899.99999999997 197700.0 156700.0 198500.0 ;
      RECT  157500.0 197700.0 158300.0 198500.0 ;
      RECT  157500.0 197700.0 158300.0 198500.0 ;
      RECT  155899.99999999997 197700.0 156700.0 198500.0 ;
      RECT  157500.0 197700.0 158300.0 198500.0 ;
      RECT  159100.0 197700.0 159900.0 198500.0 ;
      RECT  159100.0 197700.0 159899.99999999997 198500.0 ;
      RECT  157500.0 197700.0 158300.0 198500.0 ;
      RECT  160700.0 203900.00000000003 161500.0 204700.0 ;
      RECT  160700.0 197300.0 161500.0 198100.00000000003 ;
      RECT  159100.0 199400.00000000003 158300.0 200200.0 ;
      RECT  157100.0 200800.0 156300.0 201600.00000000003 ;
      RECT  157500.0 203500.0 158300.0 204300.0 ;
      RECT  159100.0 197700.0 159899.99999999997 198500.0 ;
      RECT  159899.99999999997 200800.0 159100.0 201600.00000000003 ;
      RECT  156300.0 200800.0 157100.0 201600.00000000003 ;
      RECT  158300.0 199400.00000000003 159100.0 200200.0 ;
      RECT  159100.0 200800.0 159899.99999999997 201600.00000000003 ;
      RECT  154700.0 205300.0 164300.0 205900.00000000003 ;
      RECT  154700.0 196100.00000000003 164300.0 196700.0 ;
      RECT  168700.0 204300.0 169500.0 205600.00000000003 ;
      RECT  168700.0 196400.00000000003 169500.0 197700.0 ;
      RECT  165500.0 197300.0 166300.0 196100.00000000003 ;
      RECT  165500.0 203500.0 166300.0 205900.00000000003 ;
      RECT  167300.0 197300.0 167900.0 203500.0 ;
      RECT  165500.0 203500.0 166300.0 204300.0 ;
      RECT  167100.00000000003 203500.0 167900.0 204300.0 ;
      RECT  167100.00000000003 203500.0 167900.0 204300.0 ;
      RECT  165500.0 203500.0 166300.0 204300.0 ;
      RECT  165500.0 197300.0 166300.0 198100.00000000003 ;
      RECT  167100.00000000003 197300.0 167900.0 198100.00000000003 ;
      RECT  167100.00000000003 197300.0 167900.0 198100.00000000003 ;
      RECT  165500.0 197300.0 166300.0 198100.00000000003 ;
      RECT  168700.0 203900.00000000003 169500.0 204700.0 ;
      RECT  168700.0 197300.0 169500.0 198100.00000000003 ;
      RECT  165900.0 200400.00000000003 166700.0 201200.0 ;
      RECT  165900.0 200400.00000000003 166700.0 201200.0 ;
      RECT  167600.00000000003 200500.0 168200.0 201100.00000000003 ;
      RECT  164300.0 205300.0 170700.0 205900.00000000003 ;
      RECT  164300.0 196100.00000000003 170700.0 196700.0 ;
      RECT  152700.0 206899.99999999997 153500.0 205600.00000000003 ;
      RECT  152700.0 214800.0 153500.0 213500.0 ;
      RECT  149500.0 213899.99999999997 150300.0 215100.00000000003 ;
      RECT  149500.0 207700.0 150300.0 205300.0 ;
      RECT  151300.0 213899.99999999997 151899.99999999997 207700.0 ;
      RECT  149500.0 207700.0 150300.0 206899.99999999997 ;
      RECT  151100.0 207700.0 151899.99999999997 206899.99999999997 ;
      RECT  151100.0 207700.0 151899.99999999997 206899.99999999997 ;
      RECT  149500.0 207700.0 150300.0 206899.99999999997 ;
      RECT  149500.0 213899.99999999997 150300.0 213100.00000000003 ;
      RECT  151100.0 213899.99999999997 151899.99999999997 213100.00000000003 ;
      RECT  151100.0 213899.99999999997 151899.99999999997 213100.00000000003 ;
      RECT  149500.0 213899.99999999997 150300.0 213100.00000000003 ;
      RECT  152700.0 207300.0 153500.0 206500.0 ;
      RECT  152700.0 213899.99999999997 153500.0 213100.00000000003 ;
      RECT  149899.99999999997 210800.0 150700.0 210000.0 ;
      RECT  149899.99999999997 210800.0 150700.0 210000.0 ;
      RECT  151600.0 210700.0 152200.0 210100.00000000003 ;
      RECT  148300.0 205899.99999999997 154700.0 205300.0 ;
      RECT  148300.0 215100.00000000003 154700.0 214500.0 ;
      RECT  155899.99999999997 213500.0 156700.0 215100.00000000003 ;
      RECT  155899.99999999997 207700.0 156700.0 205300.0 ;
      RECT  159100.0 207700.0 159899.99999999997 205300.0 ;
      RECT  160700.0 206899.99999999997 161500.0 205600.00000000003 ;
      RECT  160700.0 214800.0 161500.0 213500.0 ;
      RECT  155899.99999999997 207700.0 156700.0 206899.99999999997 ;
      RECT  157500.0 207700.0 158300.0 206899.99999999997 ;
      RECT  157500.0 207700.0 158300.0 206899.99999999997 ;
      RECT  155899.99999999997 207700.0 156700.0 206899.99999999997 ;
      RECT  157500.0 207700.0 158300.0 206899.99999999997 ;
      RECT  159100.0 207700.0 159900.0 206899.99999999997 ;
      RECT  159100.0 207700.0 159899.99999999997 206899.99999999997 ;
      RECT  157500.0 207700.0 158300.0 206899.99999999997 ;
      RECT  155899.99999999997 213500.0 156700.0 212700.0 ;
      RECT  157500.0 213500.0 158300.0 212700.0 ;
      RECT  157500.0 213500.0 158300.0 212700.0 ;
      RECT  155899.99999999997 213500.0 156700.0 212700.0 ;
      RECT  157500.0 213500.0 158300.0 212700.0 ;
      RECT  159100.0 213500.0 159900.0 212700.0 ;
      RECT  159100.0 213500.0 159899.99999999997 212700.0 ;
      RECT  157500.0 213500.0 158300.0 212700.0 ;
      RECT  160700.0 207300.0 161500.0 206500.0 ;
      RECT  160700.0 213899.99999999997 161500.0 213100.00000000003 ;
      RECT  159100.0 211800.0 158300.0 211000.0 ;
      RECT  157100.0 210399.99999999997 156300.0 209600.00000000003 ;
      RECT  157500.0 207700.0 158300.0 206899.99999999997 ;
      RECT  159100.0 213500.0 159899.99999999997 212700.0 ;
      RECT  159899.99999999997 210399.99999999997 159100.0 209600.00000000003 ;
      RECT  156300.0 210399.99999999997 157100.0 209600.00000000003 ;
      RECT  158300.0 211800.0 159100.0 211000.0 ;
      RECT  159100.0 210399.99999999997 159899.99999999997 209600.00000000003 ;
      RECT  154700.0 205899.99999999997 164300.0 205300.0 ;
      RECT  154700.0 215100.00000000003 164300.0 214500.0 ;
      RECT  168700.0 206899.99999999997 169500.0 205600.00000000003 ;
      RECT  168700.0 214800.0 169500.0 213500.0 ;
      RECT  165500.0 213899.99999999997 166300.0 215100.00000000003 ;
      RECT  165500.0 207700.0 166300.0 205300.0 ;
      RECT  167300.0 213899.99999999997 167900.0 207700.0 ;
      RECT  165500.0 207700.0 166300.0 206899.99999999997 ;
      RECT  167100.00000000003 207700.0 167900.0 206899.99999999997 ;
      RECT  167100.00000000003 207700.0 167900.0 206899.99999999997 ;
      RECT  165500.0 207700.0 166300.0 206899.99999999997 ;
      RECT  165500.0 213899.99999999997 166300.0 213100.00000000003 ;
      RECT  167100.00000000003 213899.99999999997 167900.0 213100.00000000003 ;
      RECT  167100.00000000003 213899.99999999997 167900.0 213100.00000000003 ;
      RECT  165500.0 213899.99999999997 166300.0 213100.00000000003 ;
      RECT  168700.0 207300.0 169500.0 206500.0 ;
      RECT  168700.0 213899.99999999997 169500.0 213100.00000000003 ;
      RECT  165900.0 210800.0 166700.0 210000.0 ;
      RECT  165900.0 210800.0 166700.0 210000.0 ;
      RECT  167600.00000000003 210700.0 168200.0 210100.00000000003 ;
      RECT  164300.0 205899.99999999997 170700.0 205300.0 ;
      RECT  164300.0 215100.00000000003 170700.0 214500.0 ;
      RECT  152700.0 222700.0 153500.0 224000.0 ;
      RECT  152700.0 214800.0 153500.0 216100.00000000003 ;
      RECT  149500.0 215700.0 150300.0 214500.0 ;
      RECT  149500.0 221899.99999999997 150300.0 224300.0 ;
      RECT  151300.0 215700.0 151899.99999999997 221899.99999999997 ;
      RECT  149500.0 221899.99999999997 150300.0 222700.0 ;
      RECT  151100.0 221899.99999999997 151899.99999999997 222700.0 ;
      RECT  151100.0 221899.99999999997 151899.99999999997 222700.0 ;
      RECT  149500.0 221899.99999999997 150300.0 222700.0 ;
      RECT  149500.0 215700.0 150300.0 216500.0 ;
      RECT  151100.0 215700.0 151899.99999999997 216500.0 ;
      RECT  151100.0 215700.0 151899.99999999997 216500.0 ;
      RECT  149500.0 215700.0 150300.0 216500.0 ;
      RECT  152700.0 222300.0 153500.0 223100.00000000003 ;
      RECT  152700.0 215700.0 153500.0 216500.0 ;
      RECT  149899.99999999997 218800.0 150700.0 219600.00000000003 ;
      RECT  149899.99999999997 218800.0 150700.0 219600.00000000003 ;
      RECT  151600.0 218899.99999999997 152200.0 219500.0 ;
      RECT  148300.0 223700.0 154700.0 224300.0 ;
      RECT  148300.0 214500.0 154700.0 215100.00000000003 ;
      RECT  155899.99999999997 216100.00000000003 156700.0 214500.0 ;
      RECT  155899.99999999997 221899.99999999997 156700.0 224300.0 ;
      RECT  159100.0 221899.99999999997 159899.99999999997 224300.0 ;
      RECT  160700.0 222700.0 161500.0 224000.0 ;
      RECT  160700.0 214800.0 161500.0 216100.00000000003 ;
      RECT  155899.99999999997 221899.99999999997 156700.0 222700.0 ;
      RECT  157500.0 221899.99999999997 158300.0 222700.0 ;
      RECT  157500.0 221899.99999999997 158300.0 222700.0 ;
      RECT  155899.99999999997 221899.99999999997 156700.0 222700.0 ;
      RECT  157500.0 221899.99999999997 158300.0 222700.0 ;
      RECT  159100.0 221899.99999999997 159900.0 222700.0 ;
      RECT  159100.0 221899.99999999997 159899.99999999997 222700.0 ;
      RECT  157500.0 221899.99999999997 158300.0 222700.0 ;
      RECT  155899.99999999997 216100.00000000003 156700.0 216899.99999999997 ;
      RECT  157500.0 216100.00000000003 158300.0 216899.99999999997 ;
      RECT  157500.0 216100.00000000003 158300.0 216899.99999999997 ;
      RECT  155899.99999999997 216100.00000000003 156700.0 216899.99999999997 ;
      RECT  157500.0 216100.00000000003 158300.0 216899.99999999997 ;
      RECT  159100.0 216100.00000000003 159900.0 216899.99999999997 ;
      RECT  159100.0 216100.00000000003 159899.99999999997 216899.99999999997 ;
      RECT  157500.0 216100.00000000003 158300.0 216899.99999999997 ;
      RECT  160700.0 222300.0 161500.0 223100.00000000003 ;
      RECT  160700.0 215700.0 161500.0 216500.0 ;
      RECT  159100.0 217800.0 158300.0 218600.00000000003 ;
      RECT  157100.0 219200.0 156300.0 220000.0 ;
      RECT  157500.0 221899.99999999997 158300.0 222700.0 ;
      RECT  159100.0 216100.00000000003 159899.99999999997 216899.99999999997 ;
      RECT  159899.99999999997 219200.0 159100.0 220000.0 ;
      RECT  156300.0 219200.0 157100.0 220000.0 ;
      RECT  158300.0 217800.0 159100.0 218600.00000000003 ;
      RECT  159100.0 219200.0 159899.99999999997 220000.0 ;
      RECT  154700.0 223700.0 164300.0 224300.0 ;
      RECT  154700.0 214500.0 164300.0 215100.00000000003 ;
      RECT  168700.0 222700.0 169500.0 224000.0 ;
      RECT  168700.0 214800.0 169500.0 216100.00000000003 ;
      RECT  165500.0 215700.0 166300.0 214500.0 ;
      RECT  165500.0 221899.99999999997 166300.0 224300.0 ;
      RECT  167300.0 215700.0 167900.0 221899.99999999997 ;
      RECT  165500.0 221899.99999999997 166300.0 222700.0 ;
      RECT  167100.00000000003 221899.99999999997 167900.0 222700.0 ;
      RECT  167100.00000000003 221899.99999999997 167900.0 222700.0 ;
      RECT  165500.0 221899.99999999997 166300.0 222700.0 ;
      RECT  165500.0 215700.0 166300.0 216500.0 ;
      RECT  167100.00000000003 215700.0 167900.0 216500.0 ;
      RECT  167100.00000000003 215700.0 167900.0 216500.0 ;
      RECT  165500.0 215700.0 166300.0 216500.0 ;
      RECT  168700.0 222300.0 169500.0 223100.00000000003 ;
      RECT  168700.0 215700.0 169500.0 216500.0 ;
      RECT  165900.0 218800.0 166700.0 219600.00000000003 ;
      RECT  165900.0 218800.0 166700.0 219600.00000000003 ;
      RECT  167600.00000000003 218899.99999999997 168200.0 219500.0 ;
      RECT  164300.0 223700.0 170700.0 224300.0 ;
      RECT  164300.0 214500.0 170700.0 215100.00000000003 ;
      RECT  152700.0 225300.0 153500.0 224000.0 ;
      RECT  152700.0 233200.0 153500.0 231900.00000000003 ;
      RECT  149500.0 232300.0 150300.0 233500.0 ;
      RECT  149500.0 226100.00000000003 150300.0 223700.0 ;
      RECT  151300.0 232300.0 151899.99999999997 226100.00000000003 ;
      RECT  149500.0 226100.00000000003 150300.0 225300.0 ;
      RECT  151100.0 226100.00000000003 151899.99999999997 225300.0 ;
      RECT  151100.0 226100.00000000003 151899.99999999997 225300.0 ;
      RECT  149500.0 226100.00000000003 150300.0 225300.0 ;
      RECT  149500.0 232300.0 150300.0 231500.0 ;
      RECT  151100.0 232300.0 151899.99999999997 231500.0 ;
      RECT  151100.0 232300.0 151899.99999999997 231500.0 ;
      RECT  149500.0 232300.0 150300.0 231500.0 ;
      RECT  152700.0 225700.0 153500.0 224900.00000000003 ;
      RECT  152700.0 232300.0 153500.0 231500.0 ;
      RECT  149899.99999999997 229200.0 150700.0 228400.00000000003 ;
      RECT  149899.99999999997 229200.0 150700.0 228400.00000000003 ;
      RECT  151600.0 229100.00000000003 152200.0 228500.0 ;
      RECT  148300.0 224300.0 154700.0 223700.0 ;
      RECT  148300.0 233500.0 154700.0 232900.00000000003 ;
      RECT  155899.99999999997 231900.00000000003 156700.0 233500.0 ;
      RECT  155899.99999999997 226100.00000000003 156700.0 223700.0 ;
      RECT  159100.0 226100.00000000003 159899.99999999997 223700.0 ;
      RECT  160700.0 225300.0 161500.0 224000.0 ;
      RECT  160700.0 233200.0 161500.0 231900.00000000003 ;
      RECT  155899.99999999997 226100.00000000003 156700.0 225300.0 ;
      RECT  157500.0 226100.00000000003 158300.0 225300.0 ;
      RECT  157500.0 226100.00000000003 158300.0 225300.0 ;
      RECT  155899.99999999997 226100.00000000003 156700.0 225300.0 ;
      RECT  157500.0 226100.00000000003 158300.0 225300.0 ;
      RECT  159100.0 226100.00000000003 159900.0 225300.0 ;
      RECT  159100.0 226100.00000000003 159899.99999999997 225300.0 ;
      RECT  157500.0 226100.00000000003 158300.0 225300.0 ;
      RECT  155899.99999999997 231900.00000000003 156700.0 231100.00000000003 ;
      RECT  157500.0 231900.00000000003 158300.0 231100.00000000003 ;
      RECT  157500.0 231900.00000000003 158300.0 231100.00000000003 ;
      RECT  155899.99999999997 231900.00000000003 156700.0 231100.00000000003 ;
      RECT  157500.0 231900.00000000003 158300.0 231100.00000000003 ;
      RECT  159100.0 231900.00000000003 159900.0 231100.00000000003 ;
      RECT  159100.0 231900.00000000003 159899.99999999997 231100.00000000003 ;
      RECT  157500.0 231900.00000000003 158300.0 231100.00000000003 ;
      RECT  160700.0 225700.0 161500.0 224900.00000000003 ;
      RECT  160700.0 232300.0 161500.0 231500.0 ;
      RECT  159100.0 230200.0 158300.0 229400.00000000003 ;
      RECT  157100.0 228800.0 156300.0 228000.0 ;
      RECT  157500.0 226100.00000000003 158300.0 225300.0 ;
      RECT  159100.0 231900.00000000003 159899.99999999997 231100.00000000003 ;
      RECT  159899.99999999997 228800.0 159100.0 228000.0 ;
      RECT  156300.0 228800.0 157100.0 228000.0 ;
      RECT  158300.0 230200.0 159100.0 229400.00000000003 ;
      RECT  159100.0 228800.0 159899.99999999997 228000.0 ;
      RECT  154700.0 224300.0 164300.0 223700.0 ;
      RECT  154700.0 233500.0 164300.0 232900.00000000003 ;
      RECT  168700.0 225300.0 169500.0 224000.0 ;
      RECT  168700.0 233200.0 169500.0 231900.00000000003 ;
      RECT  165500.0 232300.0 166300.0 233500.0 ;
      RECT  165500.0 226100.00000000003 166300.0 223700.0 ;
      RECT  167300.0 232300.0 167900.0 226100.00000000003 ;
      RECT  165500.0 226100.00000000003 166300.0 225300.0 ;
      RECT  167100.00000000003 226100.00000000003 167900.0 225300.0 ;
      RECT  167100.00000000003 226100.00000000003 167900.0 225300.0 ;
      RECT  165500.0 226100.00000000003 166300.0 225300.0 ;
      RECT  165500.0 232300.0 166300.0 231500.0 ;
      RECT  167100.00000000003 232300.0 167900.0 231500.0 ;
      RECT  167100.00000000003 232300.0 167900.0 231500.0 ;
      RECT  165500.0 232300.0 166300.0 231500.0 ;
      RECT  168700.0 225700.0 169500.0 224900.00000000003 ;
      RECT  168700.0 232300.0 169500.0 231500.0 ;
      RECT  165900.0 229200.0 166700.0 228400.00000000003 ;
      RECT  165900.0 229200.0 166700.0 228400.00000000003 ;
      RECT  167600.00000000003 229100.00000000003 168200.0 228500.0 ;
      RECT  164300.0 224300.0 170700.0 223700.0 ;
      RECT  164300.0 233500.0 170700.0 232900.00000000003 ;
      RECT  152700.0 241100.00000000003 153500.0 242400.00000000003 ;
      RECT  152700.0 233200.0 153500.0 234500.0 ;
      RECT  149500.0 234100.00000000003 150300.0 232900.00000000003 ;
      RECT  149500.0 240300.0 150300.0 242700.0 ;
      RECT  151300.0 234100.00000000003 151899.99999999997 240300.0 ;
      RECT  149500.0 240300.0 150300.0 241100.00000000003 ;
      RECT  151100.0 240300.0 151899.99999999997 241100.00000000003 ;
      RECT  151100.0 240300.0 151899.99999999997 241100.00000000003 ;
      RECT  149500.0 240300.0 150300.0 241100.00000000003 ;
      RECT  149500.0 234100.00000000003 150300.0 234900.00000000003 ;
      RECT  151100.0 234100.00000000003 151899.99999999997 234900.00000000003 ;
      RECT  151100.0 234100.00000000003 151899.99999999997 234900.00000000003 ;
      RECT  149500.0 234100.00000000003 150300.0 234900.00000000003 ;
      RECT  152700.0 240700.0 153500.0 241500.0 ;
      RECT  152700.0 234100.00000000003 153500.0 234900.00000000003 ;
      RECT  149899.99999999997 237200.0 150700.0 238000.0 ;
      RECT  149899.99999999997 237200.0 150700.0 238000.0 ;
      RECT  151600.0 237300.0 152200.0 237900.00000000003 ;
      RECT  148300.0 242100.00000000003 154700.0 242700.0 ;
      RECT  148300.0 232900.00000000003 154700.0 233500.0 ;
      RECT  155899.99999999997 234500.0 156700.0 232900.00000000003 ;
      RECT  155899.99999999997 240300.0 156700.0 242700.0 ;
      RECT  159100.0 240300.0 159899.99999999997 242700.0 ;
      RECT  160700.0 241100.00000000003 161500.0 242400.00000000003 ;
      RECT  160700.0 233200.0 161500.0 234500.0 ;
      RECT  155899.99999999997 240300.0 156700.0 241100.00000000003 ;
      RECT  157500.0 240300.0 158300.0 241100.00000000003 ;
      RECT  157500.0 240300.0 158300.0 241100.00000000003 ;
      RECT  155899.99999999997 240300.0 156700.0 241100.00000000003 ;
      RECT  157500.0 240300.0 158300.0 241100.00000000003 ;
      RECT  159100.0 240300.0 159900.0 241100.00000000003 ;
      RECT  159100.0 240300.0 159899.99999999997 241100.00000000003 ;
      RECT  157500.0 240300.0 158300.0 241100.00000000003 ;
      RECT  155899.99999999997 234500.0 156700.0 235300.0 ;
      RECT  157500.0 234500.0 158300.0 235300.0 ;
      RECT  157500.0 234500.0 158300.0 235300.0 ;
      RECT  155899.99999999997 234500.0 156700.0 235300.0 ;
      RECT  157500.0 234500.0 158300.0 235300.0 ;
      RECT  159100.0 234500.0 159900.0 235300.0 ;
      RECT  159100.0 234500.0 159899.99999999997 235300.0 ;
      RECT  157500.0 234500.0 158300.0 235300.0 ;
      RECT  160700.0 240700.0 161500.0 241500.0 ;
      RECT  160700.0 234100.00000000003 161500.0 234900.00000000003 ;
      RECT  159100.0 236200.0 158300.0 237000.0 ;
      RECT  157100.0 237600.00000000003 156300.0 238400.00000000003 ;
      RECT  157500.0 240300.0 158300.0 241100.00000000003 ;
      RECT  159100.0 234500.0 159899.99999999997 235300.0 ;
      RECT  159899.99999999997 237600.00000000003 159100.0 238400.00000000003 ;
      RECT  156300.0 237600.00000000003 157100.0 238400.00000000003 ;
      RECT  158300.0 236200.0 159100.0 237000.0 ;
      RECT  159100.0 237600.00000000003 159899.99999999997 238400.00000000003 ;
      RECT  154700.0 242100.00000000003 164300.0 242700.0 ;
      RECT  154700.0 232900.00000000003 164300.0 233500.0 ;
      RECT  168700.0 241100.00000000003 169500.0 242400.00000000003 ;
      RECT  168700.0 233200.0 169500.0 234500.0 ;
      RECT  165500.0 234100.00000000003 166300.0 232900.00000000003 ;
      RECT  165500.0 240300.0 166300.0 242700.0 ;
      RECT  167300.0 234100.00000000003 167900.0 240300.0 ;
      RECT  165500.0 240300.0 166300.0 241100.00000000003 ;
      RECT  167100.00000000003 240300.0 167900.0 241100.00000000003 ;
      RECT  167100.00000000003 240300.0 167900.0 241100.00000000003 ;
      RECT  165500.0 240300.0 166300.0 241100.00000000003 ;
      RECT  165500.0 234100.00000000003 166300.0 234900.00000000003 ;
      RECT  167100.00000000003 234100.00000000003 167900.0 234900.00000000003 ;
      RECT  167100.00000000003 234100.00000000003 167900.0 234900.00000000003 ;
      RECT  165500.0 234100.00000000003 166300.0 234900.00000000003 ;
      RECT  168700.0 240700.0 169500.0 241500.0 ;
      RECT  168700.0 234100.00000000003 169500.0 234900.00000000003 ;
      RECT  165900.0 237200.0 166700.0 238000.0 ;
      RECT  165900.0 237200.0 166700.0 238000.0 ;
      RECT  167600.00000000003 237300.0 168200.0 237900.00000000003 ;
      RECT  164300.0 242100.00000000003 170700.0 242700.0 ;
      RECT  164300.0 232900.00000000003 170700.0 233500.0 ;
      RECT  152700.0 243700.0 153500.0 242400.00000000003 ;
      RECT  152700.0 251600.00000000003 153500.0 250300.0 ;
      RECT  149500.0 250700.0 150300.0 251900.00000000003 ;
      RECT  149500.0 244500.0 150300.0 242100.00000000003 ;
      RECT  151300.0 250700.0 151899.99999999997 244500.0 ;
      RECT  149500.0 244500.0 150300.0 243700.0 ;
      RECT  151100.0 244500.0 151899.99999999997 243700.0 ;
      RECT  151100.0 244500.0 151899.99999999997 243700.0 ;
      RECT  149500.0 244500.0 150300.0 243700.0 ;
      RECT  149500.0 250700.0 150300.0 249900.00000000003 ;
      RECT  151100.0 250700.0 151899.99999999997 249900.00000000003 ;
      RECT  151100.0 250700.0 151899.99999999997 249900.00000000003 ;
      RECT  149500.0 250700.0 150300.0 249900.00000000003 ;
      RECT  152700.0 244100.00000000003 153500.0 243300.0 ;
      RECT  152700.0 250700.0 153500.0 249900.00000000003 ;
      RECT  149899.99999999997 247600.00000000003 150700.0 246800.0 ;
      RECT  149899.99999999997 247600.00000000003 150700.0 246800.0 ;
      RECT  151600.0 247500.0 152200.0 246900.00000000003 ;
      RECT  148300.0 242700.0 154700.0 242100.00000000003 ;
      RECT  148300.0 251900.00000000003 154700.0 251300.0 ;
      RECT  155899.99999999997 250300.0 156700.0 251900.00000000003 ;
      RECT  155899.99999999997 244500.0 156700.0 242100.00000000003 ;
      RECT  159100.0 244500.0 159899.99999999997 242100.00000000003 ;
      RECT  160700.0 243700.0 161500.0 242400.00000000003 ;
      RECT  160700.0 251600.00000000003 161500.0 250300.0 ;
      RECT  155899.99999999997 244500.0 156700.0 243700.0 ;
      RECT  157500.0 244500.0 158300.0 243700.0 ;
      RECT  157500.0 244500.0 158300.0 243700.0 ;
      RECT  155899.99999999997 244500.0 156700.0 243700.0 ;
      RECT  157500.0 244500.0 158300.0 243700.0 ;
      RECT  159100.0 244500.0 159900.0 243700.0 ;
      RECT  159100.0 244500.0 159899.99999999997 243700.0 ;
      RECT  157500.0 244500.0 158300.0 243700.0 ;
      RECT  155899.99999999997 250300.0 156700.0 249500.0 ;
      RECT  157500.0 250300.0 158300.0 249500.0 ;
      RECT  157500.0 250300.0 158300.0 249500.0 ;
      RECT  155899.99999999997 250300.0 156700.0 249500.0 ;
      RECT  157500.0 250300.0 158300.0 249500.0 ;
      RECT  159100.0 250300.0 159900.0 249500.0 ;
      RECT  159100.0 250300.0 159899.99999999997 249500.0 ;
      RECT  157500.0 250300.0 158300.0 249500.0 ;
      RECT  160700.0 244100.00000000003 161500.0 243300.0 ;
      RECT  160700.0 250700.0 161500.0 249900.00000000003 ;
      RECT  159100.0 248600.00000000003 158300.0 247800.0 ;
      RECT  157100.0 247200.0 156300.0 246400.00000000003 ;
      RECT  157500.0 244500.0 158300.0 243700.0 ;
      RECT  159100.0 250300.0 159899.99999999997 249500.0 ;
      RECT  159899.99999999997 247200.0 159100.0 246400.00000000003 ;
      RECT  156300.0 247200.0 157100.0 246400.00000000003 ;
      RECT  158300.0 248600.00000000003 159100.0 247800.0 ;
      RECT  159100.0 247200.0 159899.99999999997 246400.00000000003 ;
      RECT  154700.0 242700.0 164300.0 242100.00000000003 ;
      RECT  154700.0 251900.00000000003 164300.0 251300.0 ;
      RECT  168700.0 243700.0 169500.0 242400.00000000003 ;
      RECT  168700.0 251600.00000000003 169500.0 250300.0 ;
      RECT  165500.0 250700.0 166300.0 251900.00000000003 ;
      RECT  165500.0 244500.0 166300.0 242100.00000000003 ;
      RECT  167300.0 250700.0 167900.0 244500.0 ;
      RECT  165500.0 244500.0 166300.0 243700.0 ;
      RECT  167100.00000000003 244500.0 167900.0 243700.0 ;
      RECT  167100.00000000003 244500.0 167900.0 243700.0 ;
      RECT  165500.0 244500.0 166300.0 243700.0 ;
      RECT  165500.0 250700.0 166300.0 249900.00000000003 ;
      RECT  167100.00000000003 250700.0 167900.0 249900.00000000003 ;
      RECT  167100.00000000003 250700.0 167900.0 249900.00000000003 ;
      RECT  165500.0 250700.0 166300.0 249900.00000000003 ;
      RECT  168700.0 244100.00000000003 169500.0 243300.0 ;
      RECT  168700.0 250700.0 169500.0 249900.00000000003 ;
      RECT  165900.0 247600.00000000003 166700.0 246800.0 ;
      RECT  165900.0 247600.00000000003 166700.0 246800.0 ;
      RECT  167600.00000000003 247500.0 168200.0 246900.00000000003 ;
      RECT  164300.0 242700.0 170700.0 242100.00000000003 ;
      RECT  164300.0 251900.00000000003 170700.0 251300.0 ;
      RECT  152700.0 259500.0 153500.0 260800.0 ;
      RECT  152700.0 251600.00000000003 153500.0 252900.00000000003 ;
      RECT  149500.0 252500.0 150300.0 251300.0 ;
      RECT  149500.0 258700.0 150300.0 261100.00000000003 ;
      RECT  151300.0 252500.0 151899.99999999997 258700.0 ;
      RECT  149500.0 258700.0 150300.0 259500.0 ;
      RECT  151100.0 258700.0 151899.99999999997 259500.0 ;
      RECT  151100.0 258700.0 151899.99999999997 259500.0 ;
      RECT  149500.0 258700.0 150300.0 259500.0 ;
      RECT  149500.0 252500.0 150300.0 253300.0 ;
      RECT  151100.0 252500.0 151899.99999999997 253300.0 ;
      RECT  151100.0 252500.0 151899.99999999997 253300.0 ;
      RECT  149500.0 252500.0 150300.0 253300.0 ;
      RECT  152700.0 259100.00000000003 153500.0 259900.00000000003 ;
      RECT  152700.0 252500.0 153500.0 253300.0 ;
      RECT  149899.99999999997 255600.00000000003 150700.0 256400.00000000003 ;
      RECT  149899.99999999997 255600.00000000003 150700.0 256400.00000000003 ;
      RECT  151600.0 255700.0 152200.0 256300.0 ;
      RECT  148300.0 260500.0 154700.0 261100.00000000003 ;
      RECT  148300.0 251300.0 154700.0 251900.00000000003 ;
      RECT  155899.99999999997 252900.00000000003 156700.0 251300.0 ;
      RECT  155899.99999999997 258700.0 156700.0 261100.00000000003 ;
      RECT  159100.0 258700.0 159899.99999999997 261100.00000000003 ;
      RECT  160700.0 259500.0 161500.0 260800.0 ;
      RECT  160700.0 251600.00000000003 161500.0 252900.00000000003 ;
      RECT  155899.99999999997 258700.0 156700.0 259500.0 ;
      RECT  157500.0 258700.0 158300.0 259500.0 ;
      RECT  157500.0 258700.0 158300.0 259500.0 ;
      RECT  155899.99999999997 258700.0 156700.0 259500.0 ;
      RECT  157500.0 258700.0 158300.0 259500.0 ;
      RECT  159100.0 258700.0 159900.0 259500.0 ;
      RECT  159100.0 258700.0 159899.99999999997 259500.0 ;
      RECT  157500.0 258700.0 158300.0 259500.0 ;
      RECT  155899.99999999997 252900.00000000003 156700.0 253700.0 ;
      RECT  157500.0 252900.00000000003 158300.0 253700.0 ;
      RECT  157500.0 252900.00000000003 158300.0 253700.0 ;
      RECT  155899.99999999997 252900.00000000003 156700.0 253700.0 ;
      RECT  157500.0 252900.00000000003 158300.0 253700.0 ;
      RECT  159100.0 252900.00000000003 159900.0 253700.0 ;
      RECT  159100.0 252900.00000000003 159899.99999999997 253700.0 ;
      RECT  157500.0 252900.00000000003 158300.0 253700.0 ;
      RECT  160700.0 259100.00000000003 161500.0 259900.00000000003 ;
      RECT  160700.0 252500.0 161500.0 253300.0 ;
      RECT  159100.0 254600.00000000003 158300.0 255400.00000000003 ;
      RECT  157100.0 256000.0 156300.0 256800.0 ;
      RECT  157500.0 258700.0 158300.0 259500.0 ;
      RECT  159100.0 252900.00000000003 159899.99999999997 253700.0 ;
      RECT  159899.99999999997 256000.0 159100.0 256800.0 ;
      RECT  156300.0 256000.0 157100.0 256800.0 ;
      RECT  158300.0 254600.00000000003 159100.0 255400.00000000003 ;
      RECT  159100.0 256000.0 159899.99999999997 256800.0 ;
      RECT  154700.0 260500.0 164300.0 261100.00000000003 ;
      RECT  154700.0 251300.0 164300.0 251900.00000000003 ;
      RECT  168700.0 259500.0 169500.0 260800.0 ;
      RECT  168700.0 251600.00000000003 169500.0 252900.00000000003 ;
      RECT  165500.0 252500.0 166300.0 251300.0 ;
      RECT  165500.0 258700.0 166300.0 261100.00000000003 ;
      RECT  167300.0 252500.0 167900.0 258700.0 ;
      RECT  165500.0 258700.0 166300.0 259500.0 ;
      RECT  167100.00000000003 258700.0 167900.0 259500.0 ;
      RECT  167100.00000000003 258700.0 167900.0 259500.0 ;
      RECT  165500.0 258700.0 166300.0 259500.0 ;
      RECT  165500.0 252500.0 166300.0 253300.0 ;
      RECT  167100.00000000003 252500.0 167900.0 253300.0 ;
      RECT  167100.00000000003 252500.0 167900.0 253300.0 ;
      RECT  165500.0 252500.0 166300.0 253300.0 ;
      RECT  168700.0 259100.00000000003 169500.0 259900.00000000003 ;
      RECT  168700.0 252500.0 169500.0 253300.0 ;
      RECT  165900.0 255600.00000000003 166700.0 256400.00000000003 ;
      RECT  165900.0 255600.00000000003 166700.0 256400.00000000003 ;
      RECT  167600.00000000003 255700.0 168200.0 256300.0 ;
      RECT  164300.0 260500.0 170700.0 261100.00000000003 ;
      RECT  164300.0 251300.0 170700.0 251900.00000000003 ;
      RECT  152700.0 262100.00000000003 153500.0 260800.0 ;
      RECT  152700.0 270000.0 153500.0 268700.0 ;
      RECT  149500.0 269100.0 150300.0 270300.0 ;
      RECT  149500.0 262900.00000000006 150300.0 260500.0 ;
      RECT  151300.0 269100.0 151899.99999999997 262900.00000000006 ;
      RECT  149500.0 262900.00000000006 150300.0 262100.00000000003 ;
      RECT  151100.0 262900.00000000006 151899.99999999997 262100.00000000003 ;
      RECT  151100.0 262900.00000000006 151899.99999999997 262100.00000000003 ;
      RECT  149500.0 262900.00000000006 150300.0 262100.00000000003 ;
      RECT  149500.0 269100.0 150300.0 268300.0 ;
      RECT  151100.0 269100.0 151899.99999999997 268300.0 ;
      RECT  151100.0 269100.0 151899.99999999997 268300.0 ;
      RECT  149500.0 269100.0 150300.0 268300.0 ;
      RECT  152700.0 262500.0 153500.0 261700.0 ;
      RECT  152700.0 269100.0 153500.0 268300.0 ;
      RECT  149899.99999999997 266000.0 150700.0 265200.0 ;
      RECT  149899.99999999997 266000.0 150700.0 265200.0 ;
      RECT  151600.0 265900.00000000006 152200.0 265300.0 ;
      RECT  148300.0 261100.00000000003 154700.0 260500.0 ;
      RECT  148300.0 270300.0 154700.0 269700.0 ;
      RECT  155899.99999999997 268700.0 156700.0 270300.0 ;
      RECT  155899.99999999997 262900.00000000006 156700.0 260500.0 ;
      RECT  159100.0 262900.00000000006 159899.99999999997 260500.0 ;
      RECT  160700.0 262100.00000000003 161500.0 260800.0 ;
      RECT  160700.0 270000.0 161500.0 268700.0 ;
      RECT  155899.99999999997 262900.00000000006 156700.0 262100.00000000003 ;
      RECT  157500.0 262900.00000000006 158300.0 262100.00000000003 ;
      RECT  157500.0 262900.00000000006 158300.0 262100.00000000003 ;
      RECT  155899.99999999997 262900.00000000006 156700.0 262100.00000000003 ;
      RECT  157500.0 262900.00000000006 158300.0 262100.00000000003 ;
      RECT  159100.0 262900.00000000006 159900.0 262100.00000000003 ;
      RECT  159100.0 262900.00000000006 159899.99999999997 262100.00000000003 ;
      RECT  157500.0 262900.00000000006 158300.0 262100.00000000003 ;
      RECT  155899.99999999997 268700.0 156700.0 267900.00000000006 ;
      RECT  157500.0 268700.0 158300.0 267900.00000000006 ;
      RECT  157500.0 268700.0 158300.0 267900.00000000006 ;
      RECT  155899.99999999997 268700.0 156700.0 267900.00000000006 ;
      RECT  157500.0 268700.0 158300.0 267900.00000000006 ;
      RECT  159100.0 268700.0 159900.0 267900.00000000006 ;
      RECT  159100.0 268700.0 159899.99999999997 267900.00000000006 ;
      RECT  157500.0 268700.0 158300.0 267900.00000000006 ;
      RECT  160700.0 262500.0 161500.0 261700.0 ;
      RECT  160700.0 269100.0 161500.0 268300.0 ;
      RECT  159100.0 267000.0 158300.0 266200.0 ;
      RECT  157100.0 265600.0 156300.0 264800.0 ;
      RECT  157500.0 262900.00000000006 158300.0 262100.00000000003 ;
      RECT  159100.0 268700.0 159899.99999999997 267900.00000000006 ;
      RECT  159899.99999999997 265600.0 159100.0 264800.0 ;
      RECT  156300.0 265600.0 157100.0 264800.0 ;
      RECT  158300.0 267000.0 159100.0 266200.0 ;
      RECT  159100.0 265600.0 159899.99999999997 264800.0 ;
      RECT  154700.0 261100.00000000003 164300.0 260500.0 ;
      RECT  154700.0 270300.0 164300.0 269700.0 ;
      RECT  168700.0 262100.00000000003 169500.0 260800.0 ;
      RECT  168700.0 270000.0 169500.0 268700.0 ;
      RECT  165500.0 269100.0 166300.0 270300.0 ;
      RECT  165500.0 262900.00000000006 166300.0 260500.0 ;
      RECT  167300.0 269100.0 167900.0 262900.00000000006 ;
      RECT  165500.0 262900.00000000006 166300.0 262100.00000000003 ;
      RECT  167100.00000000003 262900.00000000006 167900.0 262100.00000000003 ;
      RECT  167100.00000000003 262900.00000000006 167900.0 262100.00000000003 ;
      RECT  165500.0 262900.00000000006 166300.0 262100.00000000003 ;
      RECT  165500.0 269100.0 166300.0 268300.0 ;
      RECT  167100.00000000003 269100.0 167900.0 268300.0 ;
      RECT  167100.00000000003 269100.0 167900.0 268300.0 ;
      RECT  165500.0 269100.0 166300.0 268300.0 ;
      RECT  168700.0 262500.0 169500.0 261700.0 ;
      RECT  168700.0 269100.0 169500.0 268300.0 ;
      RECT  165900.0 266000.0 166700.0 265200.0 ;
      RECT  165900.0 266000.0 166700.0 265200.0 ;
      RECT  167600.00000000003 265900.00000000006 168200.0 265300.0 ;
      RECT  164300.0 261100.00000000003 170700.0 260500.0 ;
      RECT  164300.0 270300.0 170700.0 269700.0 ;
      RECT  145800.0 126800.00000000001 146600.0 127600.00000000001 ;
      RECT  147100.0 125200.0 147899.99999999997 126000.0 ;
      RECT  158300.0 125800.00000000001 157500.0 126600.00000000001 ;
      RECT  145800.0 136400.0 146600.0 137200.0 ;
      RECT  147100.0 138000.0 147899.99999999997 138800.0 ;
      RECT  158300.0 137400.0 157500.0 138200.0 ;
      RECT  145800.0 145200.0 146600.0 146000.0 ;
      RECT  147100.0 143600.00000000003 147899.99999999997 144400.0 ;
      RECT  158300.0 144200.0 157500.0 145000.0 ;
      RECT  145800.0 154800.0 146600.0 155600.00000000003 ;
      RECT  147100.0 156399.99999999997 147899.99999999997 157200.0 ;
      RECT  158300.0 155800.0 157500.0 156600.00000000003 ;
      RECT  145800.0 163600.00000000003 146600.0 164399.99999999997 ;
      RECT  147100.0 162000.0 147899.99999999997 162800.0 ;
      RECT  158300.0 162600.00000000003 157500.0 163399.99999999997 ;
      RECT  145800.0 173200.0 146600.0 174000.0 ;
      RECT  147100.0 174800.0 147899.99999999997 175600.00000000003 ;
      RECT  158300.0 174200.0 157500.0 175000.0 ;
      RECT  145800.0 182000.0 146600.0 182800.0 ;
      RECT  147100.0 180399.99999999997 147899.99999999997 181200.0 ;
      RECT  158300.0 181000.0 157500.0 181800.0 ;
      RECT  145800.0 191600.00000000003 146600.0 192399.99999999997 ;
      RECT  147100.0 193200.0 147899.99999999997 194000.0 ;
      RECT  158300.0 192600.00000000003 157500.0 193399.99999999997 ;
      RECT  145800.0 200400.00000000003 146600.0 201200.0 ;
      RECT  147100.0 198800.0 147899.99999999997 199600.00000000003 ;
      RECT  158300.0 199400.00000000003 157500.0 200200.0 ;
      RECT  145800.0 210000.0 146600.0 210800.0 ;
      RECT  147100.0 211600.00000000003 147899.99999999997 212400.00000000003 ;
      RECT  158300.0 211000.0 157500.0 211800.0 ;
      RECT  145800.0 218800.0 146600.0 219600.00000000003 ;
      RECT  147100.0 217200.0 147899.99999999997 218000.0 ;
      RECT  158300.0 217800.0 157500.0 218600.00000000003 ;
      RECT  145800.0 228400.00000000003 146600.0 229200.0 ;
      RECT  147100.0 230000.0 147899.99999999997 230800.0 ;
      RECT  158300.0 229400.00000000003 157500.0 230200.0 ;
      RECT  145800.0 237200.0 146600.0 238000.0 ;
      RECT  147100.0 235600.00000000003 147899.99999999997 236400.00000000003 ;
      RECT  158300.0 236200.0 157500.0 237000.0 ;
      RECT  145800.0 246800.0 146600.0 247600.00000000003 ;
      RECT  147100.0 248400.00000000003 147899.99999999997 249200.0 ;
      RECT  158300.0 247800.0 157500.0 248600.00000000003 ;
      RECT  145800.0 255600.00000000003 146600.0 256400.00000000003 ;
      RECT  147100.0 254000.0 147899.99999999997 254800.0 ;
      RECT  158300.0 254600.00000000003 157500.0 255400.00000000003 ;
      RECT  145800.0 265200.0 146600.0 266000.0 ;
      RECT  147100.0 266800.0 147899.99999999997 267600.0 ;
      RECT  158300.0 266200.0 157500.0 267000.0 ;
      RECT  155100.0 131600.00000000003 154300.0 132400.0 ;
      RECT  164700.0 131600.00000000003 163899.99999999997 132400.0 ;
      RECT  155100.0 122400.0 154300.0 123200.0 ;
      RECT  164700.0 122400.0 163899.99999999997 123200.0 ;
      RECT  155100.0 131600.00000000003 154300.0 132400.0 ;
      RECT  164700.0 131600.00000000003 163899.99999999997 132400.0 ;
      RECT  155100.0 140800.0 154300.0 141600.00000000003 ;
      RECT  164700.0 140800.0 163899.99999999997 141600.00000000003 ;
      RECT  155100.0 150000.0 154300.0 150800.0 ;
      RECT  164700.0 150000.0 163899.99999999997 150800.0 ;
      RECT  155100.0 140800.0 154300.0 141600.00000000003 ;
      RECT  164700.0 140800.0 163899.99999999997 141600.00000000003 ;
      RECT  155100.0 150000.0 154300.0 150800.0 ;
      RECT  164700.0 150000.0 163899.99999999997 150800.0 ;
      RECT  155100.0 159200.0 154300.0 160000.0 ;
      RECT  164700.0 159200.0 163899.99999999997 160000.0 ;
      RECT  155100.0 168399.99999999997 154300.0 169200.0 ;
      RECT  164700.0 168399.99999999997 163899.99999999997 169200.0 ;
      RECT  155100.0 159200.0 154300.0 160000.0 ;
      RECT  164700.0 159200.0 163899.99999999997 160000.0 ;
      RECT  155100.0 168399.99999999997 154300.0 169200.0 ;
      RECT  164700.0 168399.99999999997 163899.99999999997 169200.0 ;
      RECT  155100.0 177600.00000000003 154300.0 178399.99999999997 ;
      RECT  164700.0 177600.00000000003 163899.99999999997 178399.99999999997 ;
      RECT  155100.0 186800.0 154300.0 187600.00000000003 ;
      RECT  164700.0 186800.0 163899.99999999997 187600.00000000003 ;
      RECT  155100.0 177600.00000000003 154300.0 178399.99999999997 ;
      RECT  164700.0 177600.00000000003 163899.99999999997 178399.99999999997 ;
      RECT  155100.0 186800.0 154300.0 187600.00000000003 ;
      RECT  164700.0 186800.0 163899.99999999997 187600.00000000003 ;
      RECT  155100.0 196000.0 154300.0 196800.0 ;
      RECT  164700.0 196000.0 163899.99999999997 196800.0 ;
      RECT  155100.0 205200.0 154300.0 206000.0 ;
      RECT  164700.0 205200.0 163899.99999999997 206000.0 ;
      RECT  155100.0 196000.0 154300.0 196800.0 ;
      RECT  164700.0 196000.0 163899.99999999997 196800.0 ;
      RECT  155100.0 205200.0 154300.0 206000.0 ;
      RECT  164700.0 205200.0 163899.99999999997 206000.0 ;
      RECT  155100.0 214400.00000000003 154300.0 215200.0 ;
      RECT  164700.0 214400.00000000003 163899.99999999997 215200.0 ;
      RECT  155100.0 223600.00000000003 154300.0 224400.00000000003 ;
      RECT  164700.0 223600.00000000003 163899.99999999997 224400.00000000003 ;
      RECT  155100.0 214400.00000000003 154300.0 215200.0 ;
      RECT  164700.0 214400.00000000003 163899.99999999997 215200.0 ;
      RECT  155100.0 223600.00000000003 154300.0 224400.00000000003 ;
      RECT  164700.0 223600.00000000003 163899.99999999997 224400.00000000003 ;
      RECT  155100.0 232800.0 154300.0 233600.00000000003 ;
      RECT  164700.0 232800.0 163899.99999999997 233600.00000000003 ;
      RECT  155100.0 242000.0 154300.0 242800.0 ;
      RECT  164700.0 242000.0 163899.99999999997 242800.0 ;
      RECT  155100.0 232800.0 154300.0 233600.00000000003 ;
      RECT  164700.0 232800.0 163899.99999999997 233600.00000000003 ;
      RECT  155100.0 242000.0 154300.0 242800.0 ;
      RECT  164700.0 242000.0 163899.99999999997 242800.0 ;
      RECT  155100.0 251200.0 154300.0 252000.0 ;
      RECT  164700.0 251200.0 163899.99999999997 252000.0 ;
      RECT  155100.0 260399.99999999997 154300.0 261200.0 ;
      RECT  164700.0 260399.99999999997 163899.99999999997 261200.0 ;
      RECT  155100.0 251200.0 154300.0 252000.0 ;
      RECT  164700.0 251200.0 163899.99999999997 252000.0 ;
      RECT  155100.0 260399.99999999997 154300.0 261200.0 ;
      RECT  164700.0 260399.99999999997 163899.99999999997 261200.0 ;
      RECT  155100.0 269600.0 154300.0 270400.00000000006 ;
      RECT  164700.0 269600.0 163899.99999999997 270400.00000000006 ;
      RECT  144100.0 125300.00000000001 147500.0 125900.0 ;
      RECT  144100.0 138100.00000000003 147500.0 138700.0 ;
      RECT  144100.0 143700.0 147500.0 144300.0 ;
      RECT  144100.0 156500.0 147500.0 157100.00000000003 ;
      RECT  144100.0 162100.00000000003 147500.0 162700.0 ;
      RECT  144100.0 174899.99999999997 147500.0 175500.0 ;
      RECT  144100.0 180500.0 147500.0 181100.00000000003 ;
      RECT  144100.0 193300.0 147500.0 193900.00000000003 ;
      RECT  144100.0 198900.00000000003 147500.0 199500.0 ;
      RECT  144100.0 211700.0 147500.0 212300.0 ;
      RECT  144100.0 217300.0 147500.0 217900.00000000003 ;
      RECT  144100.0 230100.00000000003 147500.0 230700.0 ;
      RECT  144100.0 235700.0 147500.0 236300.0 ;
      RECT  144100.0 248500.0 147500.0 249100.00000000003 ;
      RECT  144100.0 254100.00000000003 147500.0 254700.0 ;
      RECT  144100.0 266900.0 147500.0 267500.0 ;
      RECT  167600.0 126900.0 168200.0 127500.0 ;
      RECT  167600.0 136500.0 168200.0 137100.00000000003 ;
      RECT  167600.0 145300.0 168200.0 145900.0 ;
      RECT  167600.0 154899.99999999997 168200.0 155500.0 ;
      RECT  167600.0 163700.0 168200.0 164300.0 ;
      RECT  167600.0 173300.0 168200.0 173899.99999999997 ;
      RECT  167600.0 182100.00000000003 168200.0 182700.0 ;
      RECT  167600.0 191700.0 168200.0 192300.0 ;
      RECT  167600.0 200500.0 168200.0 201100.00000000003 ;
      RECT  167600.0 210100.00000000003 168200.0 210700.0 ;
      RECT  167600.0 218900.00000000003 168200.0 219500.0 ;
      RECT  167600.0 228500.0 168200.0 229100.00000000003 ;
      RECT  167600.0 237300.0 168200.0 237900.00000000003 ;
      RECT  167600.0 246900.00000000003 168200.0 247500.0 ;
      RECT  167600.0 255700.0 168200.0 256300.0 ;
      RECT  167600.0 265300.0 168200.0 265900.0 ;
      RECT  174500.0 108700.0 173700.00000000003 109500.0 ;
      RECT  175900.0 28900.000000000007 175100.00000000003 29700.000000000007 ;
      RECT  177300.0 98500.0 176500.0 99300.0 ;
      RECT  146600.00000000003 271000.0 145800.0 271800.0 ;
      RECT  173100.00000000003 271000.0 172300.0 271800.0 ;
      RECT  25400.000000000004 28900.000000000004 32700.000000000004 29500.0 ;
      RECT  25400.000000000004 49700.0 31300.000000000004 50300.00000000001 ;
      RECT  3100.0 62100.0 28500.000000000004 62700.0 ;
      RECT  29900.000000000004 65000.0 37600.0 65600.00000000001 ;
      RECT  32700.000000000004 63700.0 39200.0 64300.000000000015 ;
      RECT  31300.0 62400.00000000001 40800.0 63000.00000000001 ;
      RECT  47300.00000000001 65000.0 47900.00000000001 65600.00000000001 ;
      RECT  41600.0 65000.0 47600.0 65600.00000000001 ;
      RECT  47300.00000000001 65300.000000000015 47900.00000000001 69400.0 ;
      RECT  48900.00000000001 68500.0 49500.00000000001 69100.00000000001 ;
      RECT  48900.00000000001 68800.00000000001 49500.00000000001 69400.0 ;
      RECT  49200.0 68500.0 54000.0 69100.00000000001 ;
      RECT  55600.0 68500.0 60400.00000000001 69100.00000000001 ;
      RECT  29900.000000000004 94500.0 37200.0 95100.0 ;
      RECT  32700.000000000004 95900.0 39200.0 96500.0 ;
      RECT  46500.0 94500.0 47100.0 95100.0 ;
      RECT  40000.0 94500.0 46800.0 95100.0 ;
      RECT  46500.0 89800.00000000001 47100.0 94800.00000000001 ;
      RECT  9200.000000000002 108500.0 36800.00000000001 109100.0 ;
      RECT  38800.00000000001 108500.0 43600.00000000001 109100.0 ;
      RECT  54400.00000000001 39300.00000000001 69600.00000000001 39900.00000000001 ;
      RECT  54400.00000000001 59300.00000000001 69600.00000000001 59900.00000000001 ;
      RECT  54400.00000000001 19300.0 69600.00000000001 19900.000000000004 ;
      RECT  51200.0 79300.00000000001 69600.00000000001 79900.0 ;
      RECT  51200.0 99300.00000000001 69600.00000000001 99900.0 ;
      RECT  52800.00000000001 119300.00000000001 69600.00000000001 119900.0 ;
      RECT  52800.00000000001 99300.00000000001 69600.00000000001 99900.0 ;
      RECT  0.0 19600.0 21800.0 39600.0 ;
      RECT  26200.000000000004 38300.0 27000.0 39600.0 ;
      RECT  26200.000000000004 19600.0 27000.0 20900.000000000004 ;
      RECT  23000.0 20900.000000000004 23800.0 19300.0 ;
      RECT  23000.0 36700.0 23800.0 39900.00000000001 ;
      RECT  24800.0 20900.000000000004 25400.000000000004 36700.0 ;
      RECT  23000.0 36700.0 23800.0 37500.0 ;
      RECT  24600.0 36700.0 25400.000000000004 37500.0 ;
      RECT  24600.0 36700.0 25400.000000000004 37500.0 ;
      RECT  23000.0 36700.0 23800.0 37500.0 ;
      RECT  23000.0 20900.000000000004 23800.0 21700.000000000004 ;
      RECT  24600.0 20900.000000000004 25400.000000000004 21700.000000000004 ;
      RECT  24600.0 20900.000000000004 25400.000000000004 21700.000000000004 ;
      RECT  23000.0 20900.000000000004 23800.0 21700.000000000004 ;
      RECT  26200.000000000004 37900.00000000001 27000.0 38700.0 ;
      RECT  26200.000000000004 20500.0 27000.0 21300.0 ;
      RECT  23400.000000000004 28800.000000000004 24200.000000000004 29600.0 ;
      RECT  23400.000000000004 28800.000000000004 24200.000000000004 29600.0 ;
      RECT  25100.0 28900.000000000004 25700.000000000004 29500.0 ;
      RECT  21800.0 39300.00000000001 28200.000000000004 39900.00000000001 ;
      RECT  21800.0 19300.0 28200.000000000004 19900.000000000004 ;
      RECT  23400.000000000004 28800.000000000004 24200.000000000004 29600.0 ;
      RECT  25000.0 28800.000000000004 25800.0 29600.0 ;
      RECT  0.0 39000.0 28200.000000000004 40200.0 ;
      RECT  0.0 19000.0 28200.000000000004 20200.000000000004 ;
      RECT  0.0 59600.0 21800.0 39600.0 ;
      RECT  26200.000000000004 40900.00000000001 27000.0 39600.0 ;
      RECT  26200.000000000004 59600.0 27000.0 58300.00000000001 ;
      RECT  23000.0 58300.00000000001 23800.0 59900.0 ;
      RECT  23000.0 42500.0 23800.0 39300.0 ;
      RECT  24800.0 58300.00000000001 25400.000000000004 42500.0 ;
      RECT  23000.0 42500.0 23800.0 41700.0 ;
      RECT  24600.0 42500.0 25400.000000000004 41700.0 ;
      RECT  24600.0 42500.0 25400.000000000004 41700.0 ;
      RECT  23000.0 42500.0 23800.0 41700.0 ;
      RECT  23000.0 58300.00000000001 23800.0 57500.0 ;
      RECT  24600.0 58300.00000000001 25400.000000000004 57500.0 ;
      RECT  24600.0 58300.00000000001 25400.000000000004 57500.0 ;
      RECT  23000.0 58300.00000000001 23800.0 57500.0 ;
      RECT  26200.000000000004 41300.0 27000.0 40500.0 ;
      RECT  26200.000000000004 58700.0 27000.0 57900.0 ;
      RECT  23400.000000000004 50400.0 24200.000000000004 49600.0 ;
      RECT  23400.000000000004 50400.0 24200.000000000004 49600.0 ;
      RECT  25100.0 50300.0 25700.000000000004 49700.0 ;
      RECT  21800.0 39900.0 28200.000000000004 39300.0 ;
      RECT  21800.0 59900.0 28200.000000000004 59300.00000000001 ;
      RECT  23400.000000000004 50400.0 24200.000000000004 49600.0 ;
      RECT  25000.0 50400.0 25800.0 49600.0 ;
      RECT  0.0 40200.0 28200.000000000004 39000.0 ;
      RECT  0.0 60200.0 28200.000000000004 59000.0 ;
      RECT  400.0 39200.0 -400.0 40000.0 ;
      RECT  400.0 19200.000000000004 -400.0 20000.0 ;
      RECT  400.0 39200.0 -400.0 40000.0 ;
      RECT  400.0 59200.0 -400.0 60000.0 ;
      RECT  38500.0 28900.000000000004 39100.0 29500.0 ;
      RECT  38500.0 29200.000000000004 39100.0 29400.000000000004 ;
      RECT  38800.00000000001 28900.000000000004 43600.0 29500.0 ;
      RECT  44900.00000000001 28500.0 45500.0 29100.0 ;
      RECT  44900.00000000001 28800.000000000004 45500.0 29200.000000000004 ;
      RECT  45200.0 28500.0 50000.0 29100.0 ;
      RECT  38800.00000000001 50100.0 50000.0 50700.0 ;
      RECT  39600.0 38300.0 40400.00000000001 39600.0 ;
      RECT  39600.0 19600.0 40400.00000000001 20900.000000000004 ;
      RECT  36400.00000000001 20500.0 37200.0 19300.0 ;
      RECT  36400.00000000001 37500.0 37200.0 39900.00000000001 ;
      RECT  38200.0 20500.0 38800.00000000001 37500.0 ;
      RECT  36400.00000000001 37500.0 37200.0 38300.0 ;
      RECT  38000.0 37500.0 38800.00000000001 38300.0 ;
      RECT  38000.0 37500.0 38800.00000000001 38300.0 ;
      RECT  36400.00000000001 37500.0 37200.0 38300.0 ;
      RECT  36400.00000000001 20500.0 37200.0 21300.0 ;
      RECT  38000.0 20500.0 38800.00000000001 21300.0 ;
      RECT  38000.0 20500.0 38800.00000000001 21300.0 ;
      RECT  36400.00000000001 20500.0 37200.0 21300.0 ;
      RECT  39600.0 37900.00000000001 40400.00000000001 38700.0 ;
      RECT  39600.0 20500.0 40400.00000000001 21300.0 ;
      RECT  36800.00000000001 29000.0 37600.0 29800.000000000004 ;
      RECT  36800.00000000001 29000.0 37600.0 29800.000000000004 ;
      RECT  38500.0 29100.0 39100.0 29700.000000000004 ;
      RECT  35200.0 39300.00000000001 41600.0 39900.00000000001 ;
      RECT  35200.0 19300.0 41600.0 19900.000000000004 ;
      RECT  46000.0 38300.0 46800.00000000001 39600.0 ;
      RECT  46000.0 19600.0 46800.00000000001 20900.000000000004 ;
      RECT  42800.00000000001 20900.000000000004 43600.0 19300.0 ;
      RECT  42800.00000000001 36700.0 43600.0 39900.00000000001 ;
      RECT  44600.0 20900.000000000004 45200.0 36700.0 ;
      RECT  42800.00000000001 36700.0 43600.0 37500.0 ;
      RECT  44400.00000000001 36700.0 45200.0 37500.0 ;
      RECT  44400.00000000001 36700.0 45200.0 37500.0 ;
      RECT  42800.00000000001 36700.0 43600.0 37500.0 ;
      RECT  42800.00000000001 20900.000000000004 43600.0 21700.000000000004 ;
      RECT  44400.00000000001 20900.000000000004 45200.0 21700.000000000004 ;
      RECT  44400.00000000001 20900.000000000004 45200.0 21700.000000000004 ;
      RECT  42800.00000000001 20900.000000000004 43600.0 21700.000000000004 ;
      RECT  46000.0 37900.00000000001 46800.00000000001 38700.0 ;
      RECT  46000.0 20500.0 46800.00000000001 21300.0 ;
      RECT  43200.0 28800.000000000004 44000.0 29600.0 ;
      RECT  43200.0 28800.000000000004 44000.0 29600.0 ;
      RECT  44900.00000000001 28900.000000000004 45500.0 29500.0 ;
      RECT  41600.0 39300.00000000001 48000.0 39900.00000000001 ;
      RECT  41600.0 19300.0 48000.0 19900.000000000004 ;
      RECT  52400.00000000001 38300.0 53200.0 39600.0 ;
      RECT  52400.00000000001 19600.0 53200.0 20900.000000000004 ;
      RECT  49200.0 21700.000000000004 50000.0 19300.0 ;
      RECT  49200.0 35100.0 50000.0 39900.00000000001 ;
      RECT  51000.0 21700.000000000004 51600.00000000001 35100.0 ;
      RECT  49200.0 35100.0 50000.0 35900.00000000001 ;
      RECT  50800.00000000001 35100.0 51600.00000000001 35900.00000000001 ;
      RECT  50800.00000000001 35100.0 51600.00000000001 35900.00000000001 ;
      RECT  49200.0 35100.0 50000.0 35900.00000000001 ;
      RECT  49200.0 21700.000000000004 50000.0 22500.0 ;
      RECT  50800.00000000001 21700.000000000004 51600.00000000001 22500.0 ;
      RECT  50800.00000000001 21700.000000000004 51600.00000000001 22500.0 ;
      RECT  49200.0 21700.000000000004 50000.0 22500.0 ;
      RECT  52400.00000000001 37900.00000000001 53200.0 38700.0 ;
      RECT  52400.00000000001 20500.0 53200.0 21300.0 ;
      RECT  49600.0 28400.000000000004 50400.00000000001 29200.000000000004 ;
      RECT  49600.0 28400.000000000004 50400.00000000001 29200.000000000004 ;
      RECT  51300.00000000001 28500.0 51900.00000000001 29100.0 ;
      RECT  48000.0 39300.00000000001 54400.00000000001 39900.00000000001 ;
      RECT  48000.0 19300.0 54400.00000000001 19900.000000000004 ;
      RECT  52400.00000000001 40900.00000000001 53200.0 39600.0 ;
      RECT  52400.00000000001 59600.0 53200.0 58300.00000000001 ;
      RECT  49200.0 57500.0 50000.0 59900.0 ;
      RECT  49200.0 44100.0 50000.0 39300.0 ;
      RECT  51000.0 57500.0 51600.00000000001 44100.0 ;
      RECT  49200.0 44100.0 50000.0 43300.0 ;
      RECT  50800.00000000001 44100.0 51600.00000000001 43300.0 ;
      RECT  50800.00000000001 44100.0 51600.00000000001 43300.0 ;
      RECT  49200.0 44100.0 50000.0 43300.0 ;
      RECT  49200.0 57500.0 50000.0 56700.0 ;
      RECT  50800.00000000001 57500.0 51600.00000000001 56700.0 ;
      RECT  50800.00000000001 57500.0 51600.00000000001 56700.0 ;
      RECT  49200.0 57500.0 50000.0 56700.0 ;
      RECT  52400.00000000001 41300.0 53200.0 40500.0 ;
      RECT  52400.00000000001 58700.0 53200.0 57900.0 ;
      RECT  49600.0 50800.0 50400.00000000001 50000.0 ;
      RECT  49600.0 50800.0 50400.00000000001 50000.0 ;
      RECT  51300.00000000001 50700.0 51900.00000000001 50100.0 ;
      RECT  48000.0 39900.0 54400.00000000001 39300.0 ;
      RECT  48000.0 59900.0 54400.00000000001 59300.00000000001 ;
      RECT  39200.0 50000.0 38400.00000000001 50800.00000000001 ;
      RECT  38400.00000000001 29000.0 39200.0 29800.000000000004 ;
      RECT  51200.0 50000.0 52000.0 50800.00000000001 ;
      RECT  51200.0 28400.000000000004 52000.0 29200.000000000004 ;
      RECT  36800.00000000001 29000.0 37600.0 29800.000000000004 ;
      RECT  35200.0 39300.00000000001 54400.00000000001 39900.00000000001 ;
      RECT  35200.0 59300.00000000001 54400.00000000001 59900.00000000001 ;
      RECT  35200.0 19300.0 54400.00000000001 19900.000000000004 ;
      RECT  36400.00000000001 60900.0 37200.0 59300.00000000001 ;
      RECT  36400.00000000001 77500.0 37200.0 79900.0 ;
      RECT  39600.0 77500.0 40400.00000000001 79900.0 ;
      RECT  42800.00000000001 78300.00000000001 43600.0 79600.0 ;
      RECT  42800.00000000001 59600.0 43600.0 60900.0 ;
      RECT  36400.00000000001 77500.0 37200.0 78300.00000000001 ;
      RECT  38000.0 77500.0 38800.00000000001 78300.00000000001 ;
      RECT  38000.0 77500.0 38800.00000000001 78300.00000000001 ;
      RECT  36400.00000000001 77500.0 37200.0 78300.00000000001 ;
      RECT  38000.0 77500.0 38800.00000000001 78300.00000000001 ;
      RECT  39600.0 77500.0 40400.00000000001 78300.00000000001 ;
      RECT  39600.0 77500.0 40400.00000000001 78300.00000000001 ;
      RECT  38000.0 77500.0 38800.00000000001 78300.00000000001 ;
      RECT  39600.0 77500.0 40400.00000000001 78300.00000000001 ;
      RECT  41200.0 77500.0 42000.0 78300.00000000001 ;
      RECT  41200.0 77500.0 42000.0 78300.00000000001 ;
      RECT  39600.0 77500.0 40400.00000000001 78300.00000000001 ;
      RECT  36400.00000000001 60900.0 37200.0 61700.0 ;
      RECT  38000.0 60900.0 38800.00000000001 61700.0 ;
      RECT  38000.0 60900.0 38800.00000000001 61700.0 ;
      RECT  36400.00000000001 60900.0 37200.0 61700.0 ;
      RECT  38000.0 60900.0 38800.00000000001 61700.0 ;
      RECT  39600.0 60900.0 40400.00000000001 61700.0 ;
      RECT  39600.0 60900.0 40400.00000000001 61700.0 ;
      RECT  38000.0 60900.0 38800.00000000001 61700.0 ;
      RECT  39600.0 60900.0 40400.00000000001 61700.0 ;
      RECT  41200.0 60900.0 42000.0 61700.0 ;
      RECT  41200.0 60900.0 42000.0 61700.0 ;
      RECT  39600.0 60900.0 40400.00000000001 61700.0 ;
      RECT  42800.00000000001 77900.0 43600.0 78700.0 ;
      RECT  42800.00000000001 60500.0 43600.0 61300.00000000001 ;
      RECT  41200.0 62300.00000000001 40400.00000000001 63100.0 ;
      RECT  39600.0 63600.0 38800.00000000001 64400.00000000001 ;
      RECT  38000.0 64900.00000000001 37200.0 65700.0 ;
      RECT  38000.0 77500.0 38800.00000000001 78300.00000000001 ;
      RECT  41200.0 77500.0 42000.0 78300.00000000001 ;
      RECT  41200.0 60900.0 42000.0 61700.0 ;
      RECT  41200.0 64900.00000000001 42000.0 65700.0 ;
      RECT  37200.0 64900.00000000001 38000.0 65700.0 ;
      RECT  38800.00000000001 63600.0 39600.0 64400.00000000001 ;
      RECT  40400.00000000001 62300.00000000001 41200.0 63100.0 ;
      RECT  41200.0 64900.00000000001 42000.0 65700.0 ;
      RECT  35200.0 79300.00000000001 45600.0 79900.0 ;
      RECT  35200.0 59300.00000000001 45600.0 59900.0 ;
      RECT  50000.0 78300.00000000001 50800.00000000001 79600.0 ;
      RECT  50000.0 59600.0 50800.00000000001 60900.0 ;
      RECT  46800.00000000001 60500.0 47600.0 59300.00000000001 ;
      RECT  46800.00000000001 77500.0 47600.0 79900.0 ;
      RECT  48600.0 60500.0 49200.0 77500.0 ;
      RECT  46800.00000000001 77500.0 47600.0 78300.00000000001 ;
      RECT  48400.0 77500.0 49200.0 78300.00000000001 ;
      RECT  48400.0 77500.0 49200.0 78300.00000000001 ;
      RECT  46800.00000000001 77500.0 47600.0 78300.00000000001 ;
      RECT  46800.00000000001 60500.0 47600.0 61300.00000000001 ;
      RECT  48400.0 60500.0 49200.0 61300.00000000001 ;
      RECT  48400.0 60500.0 49200.0 61300.00000000001 ;
      RECT  46800.00000000001 60500.0 47600.0 61300.00000000001 ;
      RECT  50000.0 77900.0 50800.00000000001 78700.0 ;
      RECT  50000.0 60500.0 50800.00000000001 61300.00000000001 ;
      RECT  47200.0 69000.0 48000.0 69800.00000000001 ;
      RECT  47200.0 69000.0 48000.0 69800.00000000001 ;
      RECT  48900.0 69100.0 49500.0 69700.0 ;
      RECT  45600.0 79300.00000000001 52000.0 79900.0 ;
      RECT  45600.0 59300.00000000001 52000.0 59900.0 ;
      RECT  56400.0 78300.00000000001 57200.0 79600.0 ;
      RECT  56400.0 59600.0 57200.0 60900.0 ;
      RECT  53200.0 61700.0 54000.0 59300.00000000001 ;
      RECT  53200.0 75100.0 54000.0 79900.0 ;
      RECT  55000.0 61700.0 55600.0 75100.0 ;
      RECT  53200.0 75100.0 54000.0 75900.0 ;
      RECT  54800.0 75100.0 55600.0 75900.0 ;
      RECT  54800.0 75100.0 55600.0 75900.0 ;
      RECT  53200.0 75100.0 54000.0 75900.0 ;
      RECT  53200.0 61700.0 54000.0 62500.0 ;
      RECT  54800.0 61700.0 55600.0 62500.0 ;
      RECT  54800.0 61700.0 55600.0 62500.0 ;
      RECT  53200.0 61700.0 54000.0 62500.0 ;
      RECT  56400.0 77900.0 57200.0 78700.0 ;
      RECT  56400.0 60500.0 57200.0 61300.00000000001 ;
      RECT  53600.0 68400.0 54400.0 69200.0 ;
      RECT  53600.0 68400.0 54400.0 69200.0 ;
      RECT  55300.0 68500.0 55900.0 69100.0 ;
      RECT  52000.0 79300.00000000001 58400.0 79900.0 ;
      RECT  52000.0 59300.00000000001 58400.0 59900.0 ;
      RECT  67600.00000000001 78300.00000000001 68400.0 79600.0 ;
      RECT  67600.00000000001 59600.0 68400.0 60900.0 ;
      RECT  59700.0 60500.0 66700.0 59300.00000000001 ;
      RECT  59700.0 76500.0 66700.0 79900.0 ;
      RECT  64500.0 63100.0 65100.00000000001 73900.0 ;
      RECT  59700.0 75500.0 60300.00000000001 76800.00000000001 ;
      RECT  62900.00000000001 75500.0 63500.00000000001 76800.00000000001 ;
      RECT  66100.00000000001 75500.0 66700.0 76800.00000000001 ;
      RECT  61300.00000000001 74200.0 61900.00000000001 75500.0 ;
      RECT  64500.0 74200.0 65100.00000000001 75500.0 ;
      RECT  59600.00000000001 75100.0 60400.00000000001 75900.0 ;
      RECT  62800.00000000001 75100.0 63600.00000000001 75900.0 ;
      RECT  66000.0 75100.0 66800.00000000001 75900.0 ;
      RECT  61200.0 75100.0 62000.00000000001 75900.0 ;
      RECT  64400.00000000001 75100.0 65200.0 75900.0 ;
      RECT  61300.00000000001 73900.0 65100.00000000001 74500.0 ;
      RECT  59700.0 76500.0 66700.0 77100.0 ;
      RECT  59700.0 60800.00000000001 60300.00000000001 62100.0 ;
      RECT  62900.00000000001 60800.00000000001 63500.00000000001 62100.0 ;
      RECT  66100.00000000001 60800.00000000001 66700.0 62100.0 ;
      RECT  61300.00000000001 62100.0 61900.00000000001 63400.0 ;
      RECT  64500.0 62100.0 65100.00000000001 63400.0 ;
      RECT  59600.00000000001 61700.0 60400.00000000001 62500.0 ;
      RECT  62800.00000000001 61700.0 63600.00000000001 62500.0 ;
      RECT  66000.0 61700.0 66800.00000000001 62500.0 ;
      RECT  61200.0 61700.0 62000.00000000001 62500.0 ;
      RECT  64400.00000000001 61700.0 65200.0 62500.0 ;
      RECT  61300.00000000001 63100.0 65100.00000000001 63700.0 ;
      RECT  59700.0 60500.0 66700.0 61100.0 ;
      RECT  67600.00000000001 77900.0 68400.0 78700.0 ;
      RECT  67600.00000000001 60500.0 68400.0 61300.00000000001 ;
      RECT  60000.00000000001 68400.0 60800.00000000001 69200.0 ;
      RECT  60000.00000000001 68400.0 60800.00000000001 69200.0 ;
      RECT  64800.000000000015 68500.0 65400.00000000001 69100.0 ;
      RECT  58400.00000000001 79300.00000000001 69600.00000000001 79900.0 ;
      RECT  58400.00000000001 59300.00000000001 69600.00000000001 59900.0 ;
      RECT  36400.00000000001 98300.00000000001 37200.0 99900.0 ;
      RECT  36400.00000000001 81699.99999999999 37200.0 79300.0 ;
      RECT  39600.0 81699.99999999999 40400.00000000001 79300.0 ;
      RECT  41200.0 80900.0 42000.0 79600.0 ;
      RECT  41200.0 99600.0 42000.0 98300.00000000001 ;
      RECT  36400.00000000001 81700.0 37200.0 80900.0 ;
      RECT  38000.0 81700.0 38800.00000000001 80900.0 ;
      RECT  38000.0 81700.0 38800.00000000001 80900.0 ;
      RECT  36400.00000000001 81700.0 37200.0 80900.0 ;
      RECT  38000.0 81700.0 38800.00000000001 80900.0 ;
      RECT  39600.0 81700.0 40400.00000000001 80900.0 ;
      RECT  39600.0 81700.0 40400.00000000001 80900.0 ;
      RECT  38000.0 81700.0 38800.00000000001 80900.0 ;
      RECT  36400.00000000001 98300.00000000001 37200.0 97500.0 ;
      RECT  38000.0 98300.00000000001 38800.00000000001 97500.0 ;
      RECT  38000.0 98300.00000000001 38800.00000000001 97500.0 ;
      RECT  36400.00000000001 98300.00000000001 37200.0 97500.0 ;
      RECT  38000.0 98300.00000000001 38800.00000000001 97500.0 ;
      RECT  39600.0 98300.00000000001 40400.00000000001 97500.0 ;
      RECT  39600.0 98300.00000000001 40400.00000000001 97500.0 ;
      RECT  38000.0 98300.00000000001 38800.00000000001 97500.0 ;
      RECT  41200.0 81300.00000000001 42000.0 80500.0 ;
      RECT  41200.0 98699.99999999999 42000.0 97900.0 ;
      RECT  39600.0 96600.0 38800.00000000001 95800.00000000001 ;
      RECT  37600.0 95199.99999999999 36800.00000000001 94400.0 ;
      RECT  38000.0 81699.99999999999 38800.00000000001 80900.0 ;
      RECT  39600.0 98300.00000000001 40400.00000000001 97500.0 ;
      RECT  40400.00000000001 95199.99999999999 39600.0 94400.0 ;
      RECT  36800.00000000001 95199.99999999999 37600.0 94400.0 ;
      RECT  38800.00000000001 96600.0 39600.0 95800.00000000001 ;
      RECT  39600.0 95199.99999999999 40400.00000000001 94400.0 ;
      RECT  35200.0 79900.0 44800.00000000001 79300.00000000001 ;
      RECT  35200.0 99900.0 44800.00000000001 99300.00000000001 ;
      RECT  49200.0 80900.0 50000.00000000001 79600.0 ;
      RECT  49200.0 99600.0 50000.00000000001 98300.00000000001 ;
      RECT  46000.00000000001 98699.99999999999 46800.00000000001 99900.0 ;
      RECT  46000.00000000001 81699.99999999999 46800.00000000001 79300.0 ;
      RECT  47800.00000000001 98699.99999999999 48400.00000000001 81700.0 ;
      RECT  46000.00000000001 81700.0 46800.00000000001 80900.0 ;
      RECT  47600.0 81700.0 48400.00000000001 80900.0 ;
      RECT  47600.0 81700.0 48400.00000000001 80900.0 ;
      RECT  46000.00000000001 81700.0 46800.00000000001 80900.0 ;
      RECT  46000.00000000001 98699.99999999999 46800.00000000001 97900.0 ;
      RECT  47600.0 98699.99999999999 48400.00000000001 97900.0 ;
      RECT  47600.0 98699.99999999999 48400.00000000001 97900.0 ;
      RECT  46000.00000000001 98699.99999999999 46800.00000000001 97900.0 ;
      RECT  49200.0 81300.00000000001 50000.00000000001 80500.0 ;
      RECT  49200.0 98699.99999999999 50000.00000000001 97900.0 ;
      RECT  46400.00000000001 90199.99999999999 47200.0 89400.0 ;
      RECT  46400.00000000001 90199.99999999999 47200.0 89400.0 ;
      RECT  48100.0 90100.0 48700.0 89500.0 ;
      RECT  44800.00000000001 79900.0 51200.0 79300.00000000001 ;
      RECT  44800.00000000001 99900.0 51200.0 99300.00000000001 ;
      RECT  39600.0 118300.00000000001 40400.00000000001 119600.0 ;
      RECT  39600.0 99600.0 40400.00000000001 100900.0 ;
      RECT  36400.00000000001 101699.99999999999 37200.0 99300.00000000001 ;
      RECT  36400.00000000001 115100.0 37200.0 119900.0 ;
      RECT  38200.0 101699.99999999999 38800.00000000001 115100.0 ;
      RECT  36400.00000000001 115100.0 37200.0 115900.0 ;
      RECT  38000.0 115100.0 38800.00000000001 115900.0 ;
      RECT  38000.0 115100.0 38800.00000000001 115900.0 ;
      RECT  36400.00000000001 115100.0 37200.0 115900.0 ;
      RECT  36400.00000000001 101699.99999999999 37200.0 102500.0 ;
      RECT  38000.0 101699.99999999999 38800.00000000001 102500.0 ;
      RECT  38000.0 101699.99999999999 38800.00000000001 102500.0 ;
      RECT  36400.00000000001 101699.99999999999 37200.0 102500.0 ;
      RECT  39600.0 117900.0 40400.00000000001 118699.99999999999 ;
      RECT  39600.0 100500.0 40400.00000000001 101300.00000000001 ;
      RECT  36800.00000000001 108400.0 37600.0 109199.99999999999 ;
      RECT  36800.00000000001 108400.0 37600.0 109199.99999999999 ;
      RECT  38500.0 108500.0 39100.0 109100.0 ;
      RECT  35200.0 119300.00000000001 41600.0 119900.0 ;
      RECT  35200.0 99300.00000000001 41600.0 99900.0 ;
      RECT  50800.00000000001 118300.00000000001 51600.0 119600.0 ;
      RECT  50800.00000000001 99600.0 51600.0 100900.0 ;
      RECT  42900.0 100500.0 49900.00000000001 99300.00000000001 ;
      RECT  42900.0 116500.0 49900.00000000001 119900.0 ;
      RECT  47700.0 103100.0 48300.00000000001 113900.0 ;
      RECT  42900.0 115500.0 43500.0 116800.00000000001 ;
      RECT  46100.0 115500.0 46700.0 116800.00000000001 ;
      RECT  49300.00000000001 115500.0 49900.00000000001 116800.00000000001 ;
      RECT  44500.0 114199.99999999999 45100.0 115500.0 ;
      RECT  47700.0 114199.99999999999 48300.00000000001 115500.0 ;
      RECT  42800.00000000001 115100.0 43600.0 115900.0 ;
      RECT  46000.0 115100.0 46800.00000000001 115900.0 ;
      RECT  49200.0 115100.0 50000.0 115900.0 ;
      RECT  44400.0 115100.0 45200.0 115900.0 ;
      RECT  47600.0 115100.0 48400.0 115900.0 ;
      RECT  44500.0 113900.0 48300.00000000001 114500.0 ;
      RECT  42900.0 116500.0 49900.00000000001 117100.0 ;
      RECT  42900.0 100800.00000000001 43500.0 102100.0 ;
      RECT  46100.0 100800.00000000001 46700.0 102100.0 ;
      RECT  49300.00000000001 100800.00000000001 49900.00000000001 102100.0 ;
      RECT  44500.0 102100.0 45100.0 103400.0 ;
      RECT  47700.0 102100.0 48300.00000000001 103400.0 ;
      RECT  42800.00000000001 101699.99999999999 43600.0 102500.0 ;
      RECT  46000.0 101699.99999999999 46800.00000000001 102500.0 ;
      RECT  49200.0 101699.99999999999 50000.0 102500.0 ;
      RECT  44400.0 101699.99999999999 45200.0 102500.0 ;
      RECT  47600.0 101699.99999999999 48400.0 102500.0 ;
      RECT  44500.0 103100.0 48300.00000000001 103699.99999999999 ;
      RECT  42900.0 100500.0 49900.00000000001 101100.0 ;
      RECT  50800.00000000001 117900.0 51600.0 118699.99999999999 ;
      RECT  50800.00000000001 100500.0 51600.0 101300.00000000001 ;
      RECT  43200.0 108400.0 44000.0 109199.99999999999 ;
      RECT  43200.0 108400.0 44000.0 109199.99999999999 ;
      RECT  48000.0 108500.0 48600.0 109100.0 ;
      RECT  41600.0 119300.00000000001 52800.00000000001 119900.0 ;
      RECT  41600.0 99300.00000000001 52800.00000000001 99900.0 ;
      RECT  31500.000000000004 123100.00000000003 32100.0 124500.0 ;
      RECT  35400.00000000001 134700.00000000003 36800.00000000001 135500.0 ;
      RECT  35400.00000000001 150300.0 36800.00000000001 151100.0 ;
      RECT  35400.00000000001 153100.0 36800.00000000001 153900.0 ;
      RECT  35400.00000000001 168700.00000000003 36800.00000000001 169500.0 ;
      RECT  35400.00000000001 171500.0 36800.00000000001 172300.0 ;
      RECT  35400.00000000001 187100.0 36800.00000000001 187900.0 ;
      RECT  35400.00000000001 189900.0 36800.00000000001 190700.00000000003 ;
      RECT  35400.00000000001 205500.0 36800.00000000001 206299.99999999997 ;
      RECT  26800.0 132000.0 27400.000000000004 132600.00000000003 ;
      RECT  26800.0 131400.0 27400.000000000004 132000.0 ;
      RECT  27100.0 132000.0 28000.0 132600.00000000003 ;
      RECT  26800.0 131700.00000000003 27400.000000000004 132300.0 ;
      RECT  16800.0 131400.0 27100.0 132000.0 ;
      RECT  15700.000000000002 129000.0 16300.0 129600.00000000003 ;
      RECT  15700.000000000002 129300.00000000001 16300.0 129500.0 ;
      RECT  10800.0 129000.0 16000.0 129600.00000000003 ;
      RECT  8399.999999999998 125800.00000000001 7600.0 124500.0 ;
      RECT  8400.0 133700.00000000003 7600.000000000001 132400.0 ;
      RECT  11600.000000000002 132800.0 10800.0 134000.0 ;
      RECT  11600.0 126600.00000000003 10799.999999999998 124200.00000000001 ;
      RECT  9800.0 132800.0 9200.0 126600.00000000003 ;
      RECT  11600.0 126600.00000000003 10800.0 125800.00000000001 ;
      RECT  10000.0 126600.00000000003 9200.0 125800.00000000001 ;
      RECT  10000.0 126600.00000000003 9200.0 125800.00000000001 ;
      RECT  11600.0 126600.00000000003 10800.0 125800.00000000001 ;
      RECT  11600.000000000002 132800.0 10800.0 132000.0 ;
      RECT  10000.0 132800.0 9200.0 132000.0 ;
      RECT  10000.0 132800.0 9200.000000000002 132000.0 ;
      RECT  11600.000000000002 132800.0 10800.0 132000.0 ;
      RECT  8399.999999999998 126200.00000000001 7600.0 125400.0 ;
      RECT  8400.0 132800.0 7600.000000000001 132000.0 ;
      RECT  11200.0 129700.00000000001 10400.0 128900.0 ;
      RECT  11200.0 129700.00000000001 10400.0 128900.0 ;
      RECT  9500.0 129600.00000000003 8900.0 129000.0 ;
      RECT  12799.999999999998 124800.00000000001 6399.999999999999 124200.00000000001 ;
      RECT  12800.0 134000.0 6400.0 133400.0 ;
      RECT  15600.000000000002 129100.00000000003 16400.000000000004 129900.0 ;
      RECT  17200.000000000004 129100.00000000003 18000.0 129900.0 ;
      RECT  17200.000000000004 129100.00000000003 18000.0 129900.0 ;
      RECT  15600.000000000002 129100.00000000003 16400.000000000004 129900.0 ;
      RECT  4400.0 141600.00000000003 5200.0 142900.0 ;
      RECT  4400.0 133700.00000000003 5200.0 135000.0 ;
      RECT  1200.0000000000002 134600.00000000003 2000.0 133400.0 ;
      RECT  1200.0000000000002 140800.0 2000.0 143200.00000000003 ;
      RECT  3000.0 134600.00000000003 3600.0 140800.0 ;
      RECT  1200.0000000000002 140800.0 2000.0 141600.00000000003 ;
      RECT  2800.0000000000005 140800.0 3600.0000000000005 141600.00000000003 ;
      RECT  2800.0000000000005 140800.0 3600.0 141600.00000000003 ;
      RECT  1200.0000000000002 140800.0 2000.0 141600.00000000003 ;
      RECT  1200.0000000000002 134600.00000000003 2000.0 135400.0 ;
      RECT  2800.0000000000005 134600.00000000003 3600.0000000000005 135400.0 ;
      RECT  2800.0000000000005 134600.00000000003 3600.0 135400.0 ;
      RECT  1200.0000000000002 134600.00000000003 2000.0 135400.0 ;
      RECT  4400.0 141200.00000000003 5200.0 142000.0 ;
      RECT  4400.0 134600.00000000003 5200.0 135400.0 ;
      RECT  1600.0 137700.00000000003 2400.0000000000005 138500.0 ;
      RECT  1600.0 137700.00000000003 2400.0000000000005 138500.0 ;
      RECT  3300.0000000000005 137800.0 3900.0000000000005 138400.0 ;
      RECT  0.0 142600.00000000003 6400.0 143200.00000000003 ;
      RECT  0.0 133400.0 6400.0 134000.0 ;
      RECT  10800.0 141600.00000000003 11600.000000000002 142900.0 ;
      RECT  10800.0 133700.00000000003 11600.000000000002 135000.0 ;
      RECT  7600.000000000001 134600.00000000003 8400.0 133400.0 ;
      RECT  7600.000000000001 140800.0 8400.0 143200.00000000003 ;
      RECT  9400.0 134600.00000000003 10000.0 140800.0 ;
      RECT  7600.000000000001 140800.0 8400.0 141600.00000000003 ;
      RECT  9200.000000000002 140800.0 10000.0 141600.00000000003 ;
      RECT  9200.000000000002 140800.0 10000.0 141600.00000000003 ;
      RECT  7600.000000000001 140800.0 8400.0 141600.00000000003 ;
      RECT  7600.000000000001 134600.00000000003 8400.0 135400.0 ;
      RECT  9200.000000000002 134600.00000000003 10000.0 135400.0 ;
      RECT  9200.000000000002 134600.00000000003 10000.0 135400.0 ;
      RECT  7600.000000000001 134600.00000000003 8400.0 135400.0 ;
      RECT  10800.0 141200.00000000003 11600.000000000002 142000.0 ;
      RECT  10800.0 134600.00000000003 11600.000000000002 135400.0 ;
      RECT  8000.0 137700.00000000003 8800.0 138500.0 ;
      RECT  8000.0 137700.00000000003 8800.0 138500.0 ;
      RECT  9700.000000000002 137800.0 10300.0 138400.0 ;
      RECT  6400.0 142600.00000000003 12800.0 143200.00000000003 ;
      RECT  6400.0 133400.0 12800.0 134000.0 ;
      RECT  17200.000000000004 141600.00000000003 18000.0 142900.0 ;
      RECT  17200.000000000004 133700.00000000003 18000.0 135000.0 ;
      RECT  14000.0 134600.00000000003 14800.0 133400.0 ;
      RECT  14000.0 140800.0 14800.0 143200.00000000003 ;
      RECT  15800.0 134600.00000000003 16400.000000000004 140800.0 ;
      RECT  14000.0 140800.0 14800.0 141600.00000000003 ;
      RECT  15600.000000000002 140800.0 16400.000000000004 141600.00000000003 ;
      RECT  15600.000000000002 140800.0 16400.000000000004 141600.00000000003 ;
      RECT  14000.0 140800.0 14800.0 141600.00000000003 ;
      RECT  14000.0 134600.00000000003 14800.0 135400.0 ;
      RECT  15600.000000000002 134600.00000000003 16400.000000000004 135400.0 ;
      RECT  15600.000000000002 134600.00000000003 16400.000000000004 135400.0 ;
      RECT  14000.0 134600.00000000003 14800.0 135400.0 ;
      RECT  17200.000000000004 141200.00000000003 18000.0 142000.0 ;
      RECT  17200.000000000004 134600.00000000003 18000.0 135400.0 ;
      RECT  14400.0 137700.00000000003 15200.000000000002 138500.0 ;
      RECT  14400.0 137700.00000000003 15200.000000000002 138500.0 ;
      RECT  16100.000000000002 137800.0 16700.000000000004 138400.0 ;
      RECT  12800.0 142600.00000000003 19200.000000000004 143200.00000000003 ;
      RECT  12800.0 133400.0 19200.000000000004 134000.0 ;
      RECT  23600.0 141600.00000000003 24400.000000000004 142900.0 ;
      RECT  23600.0 133700.00000000003 24400.000000000004 135000.0 ;
      RECT  20400.000000000004 134600.00000000003 21200.000000000004 133400.0 ;
      RECT  20400.000000000004 140800.0 21200.000000000004 143200.00000000003 ;
      RECT  22200.000000000004 134600.00000000003 22800.000000000004 140800.0 ;
      RECT  20400.000000000004 140800.0 21200.000000000004 141600.00000000003 ;
      RECT  22000.000000000004 140800.0 22800.000000000004 141600.00000000003 ;
      RECT  22000.000000000004 140800.0 22800.000000000004 141600.00000000003 ;
      RECT  20400.000000000004 140800.0 21200.000000000004 141600.00000000003 ;
      RECT  20400.000000000004 134600.00000000003 21200.000000000004 135400.0 ;
      RECT  22000.000000000004 134600.00000000003 22800.000000000004 135400.0 ;
      RECT  22000.000000000004 134600.00000000003 22800.000000000004 135400.0 ;
      RECT  20400.000000000004 134600.00000000003 21200.000000000004 135400.0 ;
      RECT  23600.0 141200.00000000003 24400.000000000004 142000.0 ;
      RECT  23600.0 134600.00000000003 24400.000000000004 135400.0 ;
      RECT  20800.000000000004 137700.00000000003 21600.0 138500.0 ;
      RECT  20800.000000000004 137700.00000000003 21600.0 138500.0 ;
      RECT  22500.000000000004 137800.0 23100.0 138400.0 ;
      RECT  19200.000000000004 142600.00000000003 25600.0 143200.00000000003 ;
      RECT  19200.000000000004 133400.0 25600.0 134000.0 ;
      RECT  4400.0 144200.00000000003 5200.0 142900.0 ;
      RECT  4400.0 152100.0 5200.0 150800.0 ;
      RECT  1200.0000000000002 151200.00000000003 2000.0 152400.0 ;
      RECT  1200.0000000000002 145000.0 2000.0 142600.00000000003 ;
      RECT  3000.0 151200.00000000003 3600.0 145000.0 ;
      RECT  1200.0000000000002 145000.0 2000.0 144200.00000000003 ;
      RECT  2800.0000000000005 145000.0 3600.0000000000005 144200.00000000003 ;
      RECT  2800.0000000000005 145000.0 3600.0 144200.00000000003 ;
      RECT  1200.0000000000002 145000.0 2000.0 144200.00000000003 ;
      RECT  1200.0000000000002 151200.00000000003 2000.0 150400.0 ;
      RECT  2800.0000000000005 151200.00000000003 3600.0000000000005 150400.0 ;
      RECT  2800.0000000000005 151200.00000000003 3600.0 150400.0 ;
      RECT  1200.0000000000002 151200.00000000003 2000.0 150400.0 ;
      RECT  4400.0 144600.00000000003 5200.0 143800.0 ;
      RECT  4400.0 151200.00000000003 5200.0 150400.0 ;
      RECT  1600.0 148100.0 2400.0000000000005 147300.0 ;
      RECT  1600.0 148100.0 2400.0000000000005 147300.0 ;
      RECT  3300.0000000000005 148000.0 3900.0000000000005 147400.0 ;
      RECT  0.0 143200.00000000003 6400.0 142600.00000000003 ;
      RECT  0.0 152400.0 6400.0 151800.0 ;
      RECT  10800.0 144200.00000000003 11600.000000000002 142900.0 ;
      RECT  10800.0 152100.0 11600.000000000002 150800.0 ;
      RECT  7600.000000000001 151200.00000000003 8400.0 152400.0 ;
      RECT  7600.000000000001 145000.0 8400.0 142600.00000000003 ;
      RECT  9400.0 151200.00000000003 10000.0 145000.0 ;
      RECT  7600.000000000001 145000.0 8400.0 144200.00000000003 ;
      RECT  9200.000000000002 145000.0 10000.0 144200.00000000003 ;
      RECT  9200.000000000002 145000.0 10000.0 144200.00000000003 ;
      RECT  7600.000000000001 145000.0 8400.0 144200.00000000003 ;
      RECT  7600.000000000001 151200.00000000003 8400.0 150400.0 ;
      RECT  9200.000000000002 151200.00000000003 10000.0 150400.0 ;
      RECT  9200.000000000002 151200.00000000003 10000.0 150400.0 ;
      RECT  7600.000000000001 151200.00000000003 8400.0 150400.0 ;
      RECT  10800.0 144600.00000000003 11600.000000000002 143800.0 ;
      RECT  10800.0 151200.00000000003 11600.000000000002 150400.0 ;
      RECT  8000.0 148100.0 8800.0 147300.0 ;
      RECT  8000.0 148100.0 8800.0 147300.0 ;
      RECT  9700.000000000002 148000.0 10300.0 147400.0 ;
      RECT  6400.0 143200.00000000003 12800.0 142600.00000000003 ;
      RECT  6400.0 152400.0 12800.0 151800.0 ;
      RECT  17200.000000000004 144200.00000000003 18000.0 142900.0 ;
      RECT  17200.000000000004 152100.0 18000.0 150800.0 ;
      RECT  14000.0 151200.00000000003 14800.0 152400.0 ;
      RECT  14000.0 145000.0 14800.0 142600.00000000003 ;
      RECT  15800.0 151200.00000000003 16400.000000000004 145000.0 ;
      RECT  14000.0 145000.0 14800.0 144200.00000000003 ;
      RECT  15600.000000000002 145000.0 16400.000000000004 144200.00000000003 ;
      RECT  15600.000000000002 145000.0 16400.000000000004 144200.00000000003 ;
      RECT  14000.0 145000.0 14800.0 144200.00000000003 ;
      RECT  14000.0 151200.00000000003 14800.0 150400.0 ;
      RECT  15600.000000000002 151200.00000000003 16400.000000000004 150400.0 ;
      RECT  15600.000000000002 151200.00000000003 16400.000000000004 150400.0 ;
      RECT  14000.0 151200.00000000003 14800.0 150400.0 ;
      RECT  17200.000000000004 144600.00000000003 18000.0 143800.0 ;
      RECT  17200.000000000004 151200.00000000003 18000.0 150400.0 ;
      RECT  14400.0 148100.0 15200.000000000002 147300.0 ;
      RECT  14400.0 148100.0 15200.000000000002 147300.0 ;
      RECT  16100.000000000002 148000.0 16700.000000000004 147400.0 ;
      RECT  12800.0 143200.00000000003 19200.000000000004 142600.00000000003 ;
      RECT  12800.0 152400.0 19200.000000000004 151800.0 ;
      RECT  23600.0 144200.00000000003 24400.000000000004 142900.0 ;
      RECT  23600.0 152100.0 24400.000000000004 150800.0 ;
      RECT  20400.000000000004 151200.00000000003 21200.000000000004 152400.0 ;
      RECT  20400.000000000004 145000.0 21200.000000000004 142600.00000000003 ;
      RECT  22200.000000000004 151200.00000000003 22800.000000000004 145000.0 ;
      RECT  20400.000000000004 145000.0 21200.000000000004 144200.00000000003 ;
      RECT  22000.000000000004 145000.0 22800.000000000004 144200.00000000003 ;
      RECT  22000.000000000004 145000.0 22800.000000000004 144200.00000000003 ;
      RECT  20400.000000000004 145000.0 21200.000000000004 144200.00000000003 ;
      RECT  20400.000000000004 151200.00000000003 21200.000000000004 150400.0 ;
      RECT  22000.000000000004 151200.00000000003 22800.000000000004 150400.0 ;
      RECT  22000.000000000004 151200.00000000003 22800.000000000004 150400.0 ;
      RECT  20400.000000000004 151200.00000000003 21200.000000000004 150400.0 ;
      RECT  23600.0 144600.00000000003 24400.000000000004 143800.0 ;
      RECT  23600.0 151200.00000000003 24400.000000000004 150400.0 ;
      RECT  20800.000000000004 148100.0 21600.0 147300.0 ;
      RECT  20800.000000000004 148100.0 21600.0 147300.0 ;
      RECT  22500.000000000004 148000.0 23100.0 147400.0 ;
      RECT  19200.000000000004 143200.00000000003 25600.0 142600.00000000003 ;
      RECT  19200.000000000004 152400.0 25600.0 151800.0 ;
      RECT  4400.0 160000.00000000003 5200.0 161300.0 ;
      RECT  4400.0 152100.0 5200.0 153400.0 ;
      RECT  1200.0000000000002 153000.0 2000.0 151800.0 ;
      RECT  1200.0000000000002 159200.00000000003 2000.0 161600.0 ;
      RECT  3000.0 153000.0 3600.0 159200.00000000003 ;
      RECT  1200.0000000000002 159200.00000000003 2000.0 160000.00000000003 ;
      RECT  2800.0000000000005 159200.00000000003 3600.0000000000005 160000.00000000003 ;
      RECT  2800.0000000000005 159200.00000000003 3600.0 160000.00000000003 ;
      RECT  1200.0000000000002 159200.00000000003 2000.0 160000.00000000003 ;
      RECT  1200.0000000000002 153000.0 2000.0 153800.0 ;
      RECT  2800.0000000000005 153000.0 3600.0000000000005 153800.0 ;
      RECT  2800.0000000000005 153000.0 3600.0 153800.0 ;
      RECT  1200.0000000000002 153000.0 2000.0 153800.0 ;
      RECT  4400.0 159600.0 5200.0 160400.0 ;
      RECT  4400.0 153000.0 5200.0 153800.0 ;
      RECT  1600.0 156100.0 2400.0000000000005 156900.0 ;
      RECT  1600.0 156100.0 2400.0000000000005 156900.0 ;
      RECT  3300.0000000000005 156200.00000000003 3900.0000000000005 156800.0 ;
      RECT  0.0 161000.00000000003 6400.0 161600.0 ;
      RECT  0.0 151800.0 6400.0 152400.0 ;
      RECT  10800.0 160000.00000000003 11600.000000000002 161300.0 ;
      RECT  10800.0 152100.0 11600.000000000002 153400.0 ;
      RECT  7600.000000000001 153000.0 8400.0 151800.0 ;
      RECT  7600.000000000001 159200.00000000003 8400.0 161600.0 ;
      RECT  9400.0 153000.0 10000.0 159200.00000000003 ;
      RECT  7600.000000000001 159200.00000000003 8400.0 160000.00000000003 ;
      RECT  9200.000000000002 159200.00000000003 10000.0 160000.00000000003 ;
      RECT  9200.000000000002 159200.00000000003 10000.0 160000.00000000003 ;
      RECT  7600.000000000001 159200.00000000003 8400.0 160000.00000000003 ;
      RECT  7600.000000000001 153000.0 8400.0 153800.0 ;
      RECT  9200.000000000002 153000.0 10000.0 153800.0 ;
      RECT  9200.000000000002 153000.0 10000.0 153800.0 ;
      RECT  7600.000000000001 153000.0 8400.0 153800.0 ;
      RECT  10800.0 159600.0 11600.000000000002 160400.0 ;
      RECT  10800.0 153000.0 11600.000000000002 153800.0 ;
      RECT  8000.0 156100.0 8800.0 156900.0 ;
      RECT  8000.0 156100.0 8800.0 156900.0 ;
      RECT  9700.000000000002 156200.00000000003 10300.0 156800.0 ;
      RECT  6400.0 161000.00000000003 12800.0 161600.0 ;
      RECT  6400.0 151800.0 12800.0 152400.0 ;
      RECT  17200.000000000004 160000.00000000003 18000.0 161300.0 ;
      RECT  17200.000000000004 152100.0 18000.0 153400.0 ;
      RECT  14000.0 153000.0 14800.0 151800.0 ;
      RECT  14000.0 159200.00000000003 14800.0 161600.0 ;
      RECT  15800.0 153000.0 16400.000000000004 159200.00000000003 ;
      RECT  14000.0 159200.00000000003 14800.0 160000.00000000003 ;
      RECT  15600.000000000002 159200.00000000003 16400.000000000004 160000.00000000003 ;
      RECT  15600.000000000002 159200.00000000003 16400.000000000004 160000.00000000003 ;
      RECT  14000.0 159200.00000000003 14800.0 160000.00000000003 ;
      RECT  14000.0 153000.0 14800.0 153800.0 ;
      RECT  15600.000000000002 153000.0 16400.000000000004 153800.0 ;
      RECT  15600.000000000002 153000.0 16400.000000000004 153800.0 ;
      RECT  14000.0 153000.0 14800.0 153800.0 ;
      RECT  17200.000000000004 159600.0 18000.0 160400.0 ;
      RECT  17200.000000000004 153000.0 18000.0 153800.0 ;
      RECT  14400.0 156100.0 15200.000000000002 156900.0 ;
      RECT  14400.0 156100.0 15200.000000000002 156900.0 ;
      RECT  16100.000000000002 156200.00000000003 16700.000000000004 156800.0 ;
      RECT  12800.0 161000.00000000003 19200.000000000004 161600.0 ;
      RECT  12800.0 151800.0 19200.000000000004 152400.0 ;
      RECT  23600.0 160000.00000000003 24400.000000000004 161300.0 ;
      RECT  23600.0 152100.0 24400.000000000004 153400.0 ;
      RECT  20400.000000000004 153000.0 21200.000000000004 151800.0 ;
      RECT  20400.000000000004 159200.00000000003 21200.000000000004 161600.0 ;
      RECT  22200.000000000004 153000.0 22800.000000000004 159200.00000000003 ;
      RECT  20400.000000000004 159200.00000000003 21200.000000000004 160000.00000000003 ;
      RECT  22000.000000000004 159200.00000000003 22800.000000000004 160000.00000000003 ;
      RECT  22000.000000000004 159200.00000000003 22800.000000000004 160000.00000000003 ;
      RECT  20400.000000000004 159200.00000000003 21200.000000000004 160000.00000000003 ;
      RECT  20400.000000000004 153000.0 21200.000000000004 153800.0 ;
      RECT  22000.000000000004 153000.0 22800.000000000004 153800.0 ;
      RECT  22000.000000000004 153000.0 22800.000000000004 153800.0 ;
      RECT  20400.000000000004 153000.0 21200.000000000004 153800.0 ;
      RECT  23600.0 159600.0 24400.000000000004 160400.0 ;
      RECT  23600.0 153000.0 24400.000000000004 153800.0 ;
      RECT  20800.000000000004 156100.0 21600.0 156900.0 ;
      RECT  20800.000000000004 156100.0 21600.0 156900.0 ;
      RECT  22500.000000000004 156200.00000000003 23100.0 156800.0 ;
      RECT  19200.000000000004 161000.00000000003 25600.0 161600.0 ;
      RECT  19200.000000000004 151800.0 25600.0 152400.0 ;
      RECT  4400.0 162600.0 5200.0 161300.0 ;
      RECT  4400.0 170500.00000000003 5200.0 169200.00000000003 ;
      RECT  1200.0000000000002 169600.0 2000.0 170800.0 ;
      RECT  1200.0000000000002 163400.0 2000.0 161000.00000000003 ;
      RECT  3000.0 169600.0 3600.0 163400.0 ;
      RECT  1200.0000000000002 163400.0 2000.0 162600.0 ;
      RECT  2800.0000000000005 163400.0 3600.0000000000005 162600.0 ;
      RECT  2800.0000000000005 163400.0 3600.0 162600.0 ;
      RECT  1200.0000000000002 163400.0 2000.0 162600.0 ;
      RECT  1200.0000000000002 169600.0 2000.0 168800.0 ;
      RECT  2800.0000000000005 169600.0 3600.0000000000005 168800.0 ;
      RECT  2800.0000000000005 169600.0 3600.0 168800.0 ;
      RECT  1200.0000000000002 169600.0 2000.0 168800.0 ;
      RECT  4400.0 163000.00000000003 5200.0 162200.00000000003 ;
      RECT  4400.0 169600.0 5200.0 168800.0 ;
      RECT  1600.0 166500.00000000003 2400.0000000000005 165700.00000000003 ;
      RECT  1600.0 166500.00000000003 2400.0000000000005 165700.00000000003 ;
      RECT  3300.0000000000005 166400.0 3900.0000000000005 165800.0 ;
      RECT  0.0 161600.0 6400.0 161000.00000000003 ;
      RECT  0.0 170800.0 6400.0 170200.00000000003 ;
      RECT  10800.0 162600.0 11600.000000000002 161300.0 ;
      RECT  10800.0 170500.00000000003 11600.000000000002 169200.00000000003 ;
      RECT  7600.000000000001 169600.0 8400.0 170800.0 ;
      RECT  7600.000000000001 163400.0 8400.0 161000.00000000003 ;
      RECT  9400.0 169600.0 10000.0 163400.0 ;
      RECT  7600.000000000001 163400.0 8400.0 162600.0 ;
      RECT  9200.000000000002 163400.0 10000.0 162600.0 ;
      RECT  9200.000000000002 163400.0 10000.0 162600.0 ;
      RECT  7600.000000000001 163400.0 8400.0 162600.0 ;
      RECT  7600.000000000001 169600.0 8400.0 168800.0 ;
      RECT  9200.000000000002 169600.0 10000.0 168800.0 ;
      RECT  9200.000000000002 169600.0 10000.0 168800.0 ;
      RECT  7600.000000000001 169600.0 8400.0 168800.0 ;
      RECT  10800.0 163000.00000000003 11600.000000000002 162200.00000000003 ;
      RECT  10800.0 169600.0 11600.000000000002 168800.0 ;
      RECT  8000.0 166500.00000000003 8800.0 165700.00000000003 ;
      RECT  8000.0 166500.00000000003 8800.0 165700.00000000003 ;
      RECT  9700.000000000002 166400.0 10300.0 165800.0 ;
      RECT  6400.0 161600.0 12800.0 161000.00000000003 ;
      RECT  6400.0 170800.0 12800.0 170200.00000000003 ;
      RECT  17200.000000000004 162600.0 18000.0 161300.0 ;
      RECT  17200.000000000004 170500.00000000003 18000.0 169200.00000000003 ;
      RECT  14000.0 169600.0 14800.0 170800.0 ;
      RECT  14000.0 163400.0 14800.0 161000.00000000003 ;
      RECT  15800.0 169600.0 16400.000000000004 163400.0 ;
      RECT  14000.0 163400.0 14800.0 162600.0 ;
      RECT  15600.000000000002 163400.0 16400.000000000004 162600.0 ;
      RECT  15600.000000000002 163400.0 16400.000000000004 162600.0 ;
      RECT  14000.0 163400.0 14800.0 162600.0 ;
      RECT  14000.0 169600.0 14800.0 168800.0 ;
      RECT  15600.000000000002 169600.0 16400.000000000004 168800.0 ;
      RECT  15600.000000000002 169600.0 16400.000000000004 168800.0 ;
      RECT  14000.0 169600.0 14800.0 168800.0 ;
      RECT  17200.000000000004 163000.00000000003 18000.0 162200.00000000003 ;
      RECT  17200.000000000004 169600.0 18000.0 168800.0 ;
      RECT  14400.0 166500.00000000003 15200.000000000002 165700.00000000003 ;
      RECT  14400.0 166500.00000000003 15200.000000000002 165700.00000000003 ;
      RECT  16100.000000000002 166400.0 16700.000000000004 165800.0 ;
      RECT  12800.0 161600.0 19200.000000000004 161000.00000000003 ;
      RECT  12800.0 170800.0 19200.000000000004 170200.00000000003 ;
      RECT  23600.0 162600.0 24400.000000000004 161300.0 ;
      RECT  23600.0 170500.00000000003 24400.000000000004 169200.00000000003 ;
      RECT  20400.000000000004 169600.0 21200.000000000004 170800.0 ;
      RECT  20400.000000000004 163400.0 21200.000000000004 161000.00000000003 ;
      RECT  22200.000000000004 169600.0 22800.000000000004 163400.0 ;
      RECT  20400.000000000004 163400.0 21200.000000000004 162600.0 ;
      RECT  22000.000000000004 163400.0 22800.000000000004 162600.0 ;
      RECT  22000.000000000004 163400.0 22800.000000000004 162600.0 ;
      RECT  20400.000000000004 163400.0 21200.000000000004 162600.0 ;
      RECT  20400.000000000004 169600.0 21200.000000000004 168800.0 ;
      RECT  22000.000000000004 169600.0 22800.000000000004 168800.0 ;
      RECT  22000.000000000004 169600.0 22800.000000000004 168800.0 ;
      RECT  20400.000000000004 169600.0 21200.000000000004 168800.0 ;
      RECT  23600.0 163000.00000000003 24400.000000000004 162200.00000000003 ;
      RECT  23600.0 169600.0 24400.000000000004 168800.0 ;
      RECT  20800.000000000004 166500.00000000003 21600.0 165700.00000000003 ;
      RECT  20800.000000000004 166500.00000000003 21600.0 165700.00000000003 ;
      RECT  22500.000000000004 166400.0 23100.0 165800.0 ;
      RECT  19200.000000000004 161600.0 25600.0 161000.00000000003 ;
      RECT  19200.000000000004 170800.0 25600.0 170200.00000000003 ;
      RECT  8000.0 137700.00000000003 8800.0 138500.0 ;
      RECT  14400.0 137700.00000000003 15200.000000000002 138500.0 ;
      RECT  20800.0 137700.00000000003 21600.0 138500.0 ;
      RECT  1600.0 137700.00000000003 2400.0000000000005 138500.0 ;
      RECT  3200.0 137700.00000000003 4000.0 138500.0 ;
      RECT  8000.0 147300.0 8800.0 148100.0 ;
      RECT  14400.0 147300.0 15200.000000000002 148100.0 ;
      RECT  20800.0 147300.0 21600.0 148100.0 ;
      RECT  1600.0 147300.0 2400.0000000000005 148100.0 ;
      RECT  3200.0 147300.0 4000.0 148100.0 ;
      RECT  8000.0 156100.0 8800.0 156900.0 ;
      RECT  14400.0 156100.0 15200.000000000002 156900.0 ;
      RECT  20800.0 156100.0 21600.0 156900.0 ;
      RECT  1600.0 156100.0 2400.0000000000005 156900.0 ;
      RECT  3200.0 156100.0 4000.0 156900.0 ;
      RECT  8000.0 165700.00000000003 8800.0 166500.0 ;
      RECT  14400.0 165700.00000000003 15200.000000000002 166500.0 ;
      RECT  20800.0 165700.00000000003 21600.0 166500.0 ;
      RECT  1600.0 165700.00000000003 2400.0000000000005 166500.0 ;
      RECT  3200.0 165700.00000000003 4000.0 166500.0 ;
      RECT  13200.000000000002 142500.0 12400.0 143300.0 ;
      RECT  13200.000000000002 133300.0 12400.0 134100.00000000003 ;
      RECT  19600.0 142500.0 18800.0 143300.0 ;
      RECT  19600.0 133300.0 18800.0 134100.00000000003 ;
      RECT  13200.000000000002 160900.0 12400.0 161700.00000000003 ;
      RECT  13200.000000000002 151700.00000000003 12400.0 152500.0 ;
      RECT  19600.0 160900.0 18800.0 161700.00000000003 ;
      RECT  19600.0 151700.00000000003 18800.0 152500.0 ;
      RECT  13200.000000000002 170100.0 12400.0 170900.0 ;
      RECT  19600.0 170100.0 18800.0 170900.0 ;
      RECT  1600.0 137700.00000000003 2400.0000000000005 138500.0 ;
      RECT  20800.0 165700.00000000003 21600.0 166500.0 ;
      RECT  28400.000000000004 133700.00000000003 35200.0 124500.0 ;
      RECT  28400.000000000004 133700.00000000003 35200.0 142900.0 ;
      RECT  28400.000000000004 152100.0 35200.0 142900.0 ;
      RECT  28400.000000000004 152100.0 35200.0 161300.0 ;
      RECT  28400.000000000004 170500.00000000003 35200.0 161300.0 ;
      RECT  28400.000000000004 170500.00000000003 35200.0 179700.00000000003 ;
      RECT  28400.000000000004 188900.0 35200.0 179700.00000000003 ;
      RECT  28400.000000000004 188900.0 35200.0 198100.0 ;
      RECT  28400.000000000004 207300.0 35200.0 198100.0 ;
      RECT  28000.000000000004 134700.00000000003 35400.00000000001 135500.0 ;
      RECT  28000.000000000004 150300.0 35400.00000000001 151100.0 ;
      RECT  28000.000000000004 153100.0 35400.00000000001 153900.0 ;
      RECT  28000.000000000004 168700.00000000003 35400.00000000001 169500.00000000003 ;
      RECT  28000.000000000004 171500.00000000003 35400.00000000001 172300.0 ;
      RECT  28000.000000000004 187100.0 35400.00000000001 187900.0 ;
      RECT  28000.000000000004 189900.0 35400.00000000001 190700.00000000003 ;
      RECT  28000.000000000004 205500.0 35400.00000000001 206300.0 ;
      RECT  6800.000000000001 124100.00000000003 6000.000000000001 124900.0 ;
      RECT  31400.000000000004 122700.00000000001 32200.000000000004 123500.0 ;
      RECT  28800.0 128700.00000000001 28000.0 129500.0 ;
      RECT  35600.0 128700.00000000001 34800.00000000001 129500.0 ;
      RECT  37200.0 134700.00000000003 36400.00000000001 135500.0 ;
      RECT  37200.0 150300.0 36400.00000000001 151100.0 ;
      RECT  37200.0 153100.0 36400.00000000001 153900.0 ;
      RECT  37200.0 168700.00000000003 36400.00000000001 169500.0 ;
      RECT  37200.0 171500.0 36400.00000000001 172300.0 ;
      RECT  37200.0 187100.0 36400.00000000001 187900.0 ;
      RECT  37200.0 189900.0 36400.00000000001 190700.00000000003 ;
      RECT  37200.0 205500.0 36400.00000000001 206299.99999999997 ;
      RECT  16400.000000000004 131300.0 17200.000000000004 132100.00000000003 ;
      RECT  16400.000000000004 131300.0 17200.000000000004 132100.00000000003 ;
      RECT  17200.000000000004 129100.00000000003 18000.000000000004 129900.0 ;
      RECT  15600.000000000002 129100.00000000003 16400.000000000004 129900.0 ;
      RECT  8800.0 128900.0 9600.000000000002 129700.00000000001 ;
      RECT  33100.0 28800.000000000004 32300.000000000004 29600.0 ;
      RECT  25000.0 28800.000000000004 25800.0 29600.0 ;
      RECT  31700.000000000004 49600.0 30900.000000000004 50400.00000000001 ;
      RECT  25000.0 49600.0 25800.0 50400.00000000001 ;
      RECT  3500.0 62000.00000000001 2700.0 62800.00000000001 ;
      RECT  28900.000000000004 62000.00000000001 28100.0 62800.00000000001 ;
      RECT  30300.0 64900.00000000001 29500.0 65700.0 ;
      RECT  33100.0 63600.0 32300.000000000004 64400.00000000001 ;
      RECT  31700.000000000004 62300.00000000001 30900.000000000004 63100.0 ;
      RECT  30300.0 94400.0 29500.0 95199.99999999999 ;
      RECT  33100.0 95800.00000000001 32300.000000000004 96600.0 ;
      RECT  48800.00000000001 89400.0 48000.00000000001 90199.99999999999 ;
      RECT  9600.000000000002 108400.0 8800.0 109200.00000000001 ;
      RECT  70000.0 39200.0 69200.0 40000.0 ;
      RECT  70000.0 59200.0 69200.0 60000.0 ;
      RECT  70000.0 19200.000000000004 69200.0 20000.0 ;
      RECT  70000.0 79200.0 69200.0 80000.0 ;
      RECT  70000.0 59200.0 69200.0 60000.0 ;
      RECT  70000.0 79200.0 69200.0 80000.0 ;
      RECT  70000.0 99200.00000000001 69200.0 100000.0 ;
      RECT  70000.0 119200.00000000001 69200.0 120000.0 ;
      RECT  70000.0 99200.00000000001 69200.0 100000.0 ;
      RECT  48300.00000000001 108500.0 71000.0 109100.0 ;
      RECT  65100.00000000001 68500.0 71000.0 69100.0 ;
      RECT  51600.0 28500.0 71000.0 29100.0 ;
      RECT  51600.0 50100.0 71000.0 50700.0 ;
      RECT  49199.99999999999 211900.00000000003 71000.0 231900.00000000003 ;
      RECT  49199.99999999999 251900.00000000003 71000.0 231900.00000000003 ;
      RECT  49199.99999999999 251900.00000000003 71000.0 271900.00000000006 ;
      RECT  49199.99999999999 291900.00000000006 71000.0 271900.00000000006 ;
      RECT  60500.0 231500.00000000003 59699.99999999999 232300.00000000003 ;
      RECT  60500.0 211500.00000000003 59699.99999999999 212300.00000000003 ;
      RECT  60500.0 231500.00000000003 59699.99999999999 232300.00000000003 ;
      RECT  60500.0 251500.00000000003 59699.99999999999 252300.00000000003 ;
      RECT  60500.0 271500.00000000006 59699.99999999999 272300.0 ;
      RECT  60500.0 251500.00000000003 59699.99999999999 252300.00000000003 ;
      RECT  60500.0 271500.00000000006 59699.99999999999 272300.0 ;
      RECT  60500.0 291500.00000000006 59699.99999999999 292300.00000000006 ;
      RECT  178600.00000000003 0.0 200400.00000000003 20000.0 ;
      RECT  200400.00000000003 0.0 222200.00000000003 20000.0 ;
      RECT  189900.00000000003 19600.0 189100.00000000003 20400.000000000004 ;
      RECT  189900.00000000003 -400.0 189100.00000000003 400.0 ;
      RECT  211700.00000000003 19600.0 210900.00000000003 20400.000000000004 ;
      RECT  211700.00000000003 -400.0 210900.00000000003 400.0 ;
      RECT  71399.99999999999 108400.0 70600.0 109200.0 ;
      RECT  71399.99999999999 68400.0 70600.0 69200.0 ;
      RECT  71399.99999999999 28400.000000000004 70600.0 29200.000000000004 ;
      RECT  71399.99999999999 50000.0 70600.0 50800.0 ;
      RECT  182400.0 22400.000000000004 181600.0 23200.000000000004 ;
      RECT  198200.0 22400.000000000004 197399.99999999997 23200.000000000004 ;
      RECT  189200.0 23800.000000000004 188399.99999999997 24600.000000000004 ;
      RECT  220000.0 23800.000000000004 219200.0 24600.000000000004 ;
   LAYER  metal2 ;
      RECT  172400.0 3400.0000000000023 173000.0 148700.00000000003 ;
      RECT  72100.0 50400.00000000001 72699.99999999999 215300.0 ;
      RECT  176600.00000000003 108800.00000000001 177200.00000000003 148700.00000000003 ;
      RECT  175200.0 68800.00000000001 175799.99999999997 148700.00000000003 ;
      RECT  173800.0 28800.000000000004 174400.0 148700.00000000003 ;
      RECT  172400.0 50400.00000000001 173000.0 148700.00000000003 ;
      RECT  73899.99999999999 159600.00000000003 74499.99999999999 221700.00000000003 ;
      RECT  75300.0 159600.00000000003 75899.99999999999 242100.00000000003 ;
      RECT  76700.0 159600.00000000003 77300.0 261700.00000000006 ;
      RECT  78100.0 159600.00000000003 78699.99999999999 282100.0 ;
      RECT  181700.0 22800.000000000004 182299.99999999997 25200.000000000004 ;
      RECT  197500.0 9800.000000000002 198100.0 22800.000000000004 ;
      RECT  188500.0 24200.000000000004 189100.0 25200.000000000004 ;
      RECT  219300.0 9800.000000000002 219900.0 24200.000000000004 ;
      RECT  180700.0 64599.99999999999 181300.0 71500.0 ;
      RECT  180700.0 71500.0 181300.0 78400.0 ;
      RECT  182700.0 64599.99999999999 183300.0 71500.0 ;
      RECT  182700.0 71500.0 183300.0 78400.0 ;
      RECT  187500.0 64599.99999999999 188100.00000000003 71500.0 ;
      RECT  187500.0 71500.0 188100.00000000003 78400.0 ;
      RECT  189500.0 64599.99999999999 190100.00000000003 71500.0 ;
      RECT  189500.0 71500.0 190100.00000000003 78400.0 ;
      RECT  180700.0 103200.0 181300.0 103800.0 ;
      RECT  179900.0 103200.0 180500.0 103800.0 ;
      RECT  180700.0 101400.0 181300.0 103500.0 ;
      RECT  180200.0 103200.0 181000.0 103800.0 ;
      RECT  179900.0 103500.0 180500.0 105600.0 ;
      RECT  182700.0 103200.0 183300.0 103800.0 ;
      RECT  183500.0 103200.0 184100.00000000003 103800.0 ;
      RECT  182700.0 101400.0 183300.0 103500.0 ;
      RECT  183000.0 103200.0 183800.0 103800.0 ;
      RECT  183500.0 103500.0 184100.00000000003 105600.0 ;
      RECT  187500.0 103200.0 188100.00000000003 103800.0 ;
      RECT  186700.0 103200.0 187300.0 103800.0 ;
      RECT  187500.0 101400.0 188100.00000000003 103500.0 ;
      RECT  187000.0 103200.0 187800.0 103800.0 ;
      RECT  186700.0 103500.0 187300.0 105600.0 ;
      RECT  189500.0 103200.0 190100.00000000003 103800.0 ;
      RECT  190300.0 103200.0 190900.0 103800.0 ;
      RECT  189500.0 101400.0 190100.00000000003 103500.0 ;
      RECT  189800.0 103200.0 190600.00000000003 103800.0 ;
      RECT  190300.0 103500.0 190900.0 105600.0 ;
      RECT  179900.0 118200.0 180500.0 120100.00000000001 ;
      RECT  179900.0 120100.00000000001 180500.0 122000.00000000001 ;
      RECT  183500.0 118200.0 184100.00000000003 120100.00000000001 ;
      RECT  183500.0 120100.00000000001 184100.00000000003 122800.00000000001 ;
      RECT  186700.0 118200.0 187300.0 120100.00000000001 ;
      RECT  186700.0 120100.00000000001 187300.0 122000.00000000001 ;
      RECT  190300.0 118200.0 190900.0 120100.00000000001 ;
      RECT  190300.0 120100.00000000001 190900.0 122800.00000000001 ;
      RECT  145900.0 270000.0 146500.0 271400.00000000006 ;
      RECT  178600.00000000003 122400.0 185400.0 131600.00000000003 ;
      RECT  178600.00000000003 140800.0 185400.0 131600.00000000003 ;
      RECT  178600.00000000003 140800.0 185400.0 150000.0 ;
      RECT  178600.00000000003 159200.0 185400.0 150000.0 ;
      RECT  178600.00000000003 159200.0 185400.0 168400.00000000003 ;
      RECT  178600.00000000003 177600.00000000003 185400.0 168399.99999999997 ;
      RECT  178600.00000000003 177600.00000000003 185400.0 186800.0 ;
      RECT  178600.00000000003 196000.0 185400.0 186800.0 ;
      RECT  178600.00000000003 196000.0 185400.0 205200.0 ;
      RECT  178600.00000000003 214399.99999999997 185400.0 205200.0 ;
      RECT  178600.00000000003 214399.99999999997 185400.0 223600.00000000003 ;
      RECT  178600.00000000003 232800.0 185400.0 223600.00000000003 ;
      RECT  178600.00000000003 232800.0 185400.0 242000.0 ;
      RECT  178600.00000000003 251200.0 185400.0 242000.0 ;
      RECT  178600.00000000003 251200.0 185400.0 260399.99999999997 ;
      RECT  178600.00000000003 269600.0 185400.0 260400.00000000003 ;
      RECT  185400.0 122400.0 192200.0 131600.00000000003 ;
      RECT  185400.0 140800.0 192200.0 131600.00000000003 ;
      RECT  185400.0 140800.0 192200.0 150000.0 ;
      RECT  185400.0 159200.0 192200.0 150000.0 ;
      RECT  185400.0 159200.0 192200.0 168400.00000000003 ;
      RECT  185400.0 177600.00000000003 192200.0 168399.99999999997 ;
      RECT  185400.0 177600.00000000003 192200.0 186800.0 ;
      RECT  185400.0 196000.0 192200.0 186800.0 ;
      RECT  185400.0 196000.0 192200.0 205200.0 ;
      RECT  185400.0 214399.99999999997 192200.0 205200.0 ;
      RECT  185400.0 214399.99999999997 192200.0 223600.00000000003 ;
      RECT  185400.0 232800.0 192200.0 223600.00000000003 ;
      RECT  185400.0 232800.0 192200.0 242000.0 ;
      RECT  185400.0 251200.0 192200.0 242000.0 ;
      RECT  185400.0 251200.0 192200.0 260399.99999999997 ;
      RECT  185400.0 269600.0 192200.0 260400.00000000003 ;
      RECT  181600.00000000003 131200.0 182400.0 132000.0 ;
      RECT  188400.0 131200.0 189200.0 132000.0 ;
      RECT  181600.00000000003 131200.0 182400.0 132000.0 ;
      RECT  188400.0 131200.0 189200.0 132000.0 ;
      RECT  181600.00000000003 149600.00000000003 182400.0 150400.0 ;
      RECT  188400.0 149600.00000000003 189200.0 150400.0 ;
      RECT  181600.00000000003 149600.00000000003 182400.0 150400.0 ;
      RECT  188400.0 149600.00000000003 189200.0 150400.0 ;
      RECT  181600.00000000003 168000.0 182400.0 168800.0 ;
      RECT  188400.0 168000.0 189200.0 168800.0 ;
      RECT  181600.00000000003 168000.0 182400.0 168800.0 ;
      RECT  188400.0 168000.0 189200.0 168800.0 ;
      RECT  181600.00000000003 186399.99999999997 182400.0 187200.0 ;
      RECT  188400.0 186399.99999999997 189200.0 187200.0 ;
      RECT  181600.00000000003 186399.99999999997 182400.0 187200.0 ;
      RECT  188400.0 186399.99999999997 189200.0 187200.0 ;
      RECT  181600.00000000003 204800.0 182400.0 205600.00000000003 ;
      RECT  188400.0 204800.0 189200.0 205600.00000000003 ;
      RECT  181600.00000000003 204800.0 182400.0 205600.00000000003 ;
      RECT  188400.0 204800.0 189200.0 205600.00000000003 ;
      RECT  181600.00000000003 223200.0 182400.0 224000.0 ;
      RECT  188400.0 223200.0 189200.0 224000.0 ;
      RECT  181600.00000000003 223200.0 182400.0 224000.0 ;
      RECT  188400.0 223200.0 189200.0 224000.0 ;
      RECT  181600.00000000003 241600.00000000003 182400.0 242399.99999999997 ;
      RECT  188400.0 241600.00000000003 189200.0 242399.99999999997 ;
      RECT  181600.00000000003 241600.00000000003 182400.0 242399.99999999997 ;
      RECT  188400.0 241600.00000000003 189200.0 242399.99999999997 ;
      RECT  181600.00000000003 260000.0 182400.0 260800.0 ;
      RECT  188400.0 260000.0 189200.0 260800.0 ;
      RECT  181600.00000000003 260000.0 182400.0 260800.0 ;
      RECT  188400.0 260000.0 189200.0 260800.0 ;
      RECT  178200.0 126600.00000000001 179000.0 127400.0 ;
      RECT  185000.0 126600.00000000001 185800.0 127400.0 ;
      RECT  185000.0 126600.00000000001 185800.0 127400.0 ;
      RECT  191800.0 126600.00000000001 192600.00000000003 127400.0 ;
      RECT  178200.0 135800.0 179000.0 136600.00000000003 ;
      RECT  185000.0 135800.0 185800.0 136600.00000000003 ;
      RECT  185000.0 135800.0 185800.0 136600.00000000003 ;
      RECT  191800.0 135800.0 192600.00000000003 136600.00000000003 ;
      RECT  178200.0 145000.0 179000.0 145800.0 ;
      RECT  185000.0 145000.0 185800.0 145800.0 ;
      RECT  185000.0 145000.0 185800.0 145800.0 ;
      RECT  191800.0 145000.0 192600.00000000003 145800.0 ;
      RECT  178200.0 154200.0 179000.0 155000.0 ;
      RECT  185000.0 154200.0 185800.0 155000.0 ;
      RECT  185000.0 154200.0 185800.0 155000.0 ;
      RECT  191800.0 154200.0 192600.00000000003 155000.0 ;
      RECT  178200.0 163399.99999999997 179000.0 164200.0 ;
      RECT  185000.0 163399.99999999997 185800.0 164200.0 ;
      RECT  185000.0 163399.99999999997 185800.0 164200.0 ;
      RECT  191800.0 163399.99999999997 192600.00000000003 164200.0 ;
      RECT  178200.0 172600.00000000003 179000.0 173399.99999999997 ;
      RECT  185000.0 172600.00000000003 185800.0 173399.99999999997 ;
      RECT  185000.0 172600.00000000003 185800.0 173399.99999999997 ;
      RECT  191800.0 172600.00000000003 192600.00000000003 173399.99999999997 ;
      RECT  178200.0 181800.0 179000.0 182600.00000000003 ;
      RECT  185000.0 181800.0 185800.0 182600.00000000003 ;
      RECT  185000.0 181800.0 185800.0 182600.00000000003 ;
      RECT  191800.0 181800.0 192600.00000000003 182600.00000000003 ;
      RECT  178200.0 191000.0 179000.0 191800.0 ;
      RECT  185000.0 191000.0 185800.0 191800.0 ;
      RECT  185000.0 191000.0 185800.0 191800.0 ;
      RECT  191800.0 191000.0 192600.00000000003 191800.0 ;
      RECT  178200.0 200200.0 179000.0 201000.0 ;
      RECT  185000.0 200200.0 185800.0 201000.0 ;
      RECT  185000.0 200200.0 185800.0 201000.0 ;
      RECT  191800.0 200200.0 192600.00000000003 201000.0 ;
      RECT  178200.0 209399.99999999997 179000.0 210200.0 ;
      RECT  185000.0 209399.99999999997 185800.0 210200.0 ;
      RECT  185000.0 209399.99999999997 185800.0 210200.0 ;
      RECT  191800.0 209399.99999999997 192600.00000000003 210200.0 ;
      RECT  178200.0 218600.00000000003 179000.0 219399.99999999997 ;
      RECT  185000.0 218600.00000000003 185800.0 219399.99999999997 ;
      RECT  185000.0 218600.00000000003 185800.0 219399.99999999997 ;
      RECT  191800.0 218600.00000000003 192600.00000000003 219399.99999999997 ;
      RECT  178200.0 227800.0 179000.0 228600.00000000003 ;
      RECT  185000.0 227800.0 185800.0 228600.00000000003 ;
      RECT  185000.0 227800.0 185800.0 228600.00000000003 ;
      RECT  191800.0 227800.0 192600.00000000003 228600.00000000003 ;
      RECT  178200.0 237000.0 179000.0 237800.0 ;
      RECT  185000.0 237000.0 185800.0 237800.0 ;
      RECT  185000.0 237000.0 185800.0 237800.0 ;
      RECT  191800.0 237000.0 192600.00000000003 237800.0 ;
      RECT  178200.0 246200.0 179000.0 247000.0 ;
      RECT  185000.0 246200.0 185800.0 247000.0 ;
      RECT  185000.0 246200.0 185800.0 247000.0 ;
      RECT  191800.0 246200.0 192600.00000000003 247000.0 ;
      RECT  178200.0 255399.99999999997 179000.0 256200.0 ;
      RECT  185000.0 255399.99999999997 185800.0 256200.0 ;
      RECT  185000.0 255399.99999999997 185800.0 256200.0 ;
      RECT  191800.0 255399.99999999997 192600.00000000003 256200.0 ;
      RECT  178200.0 264600.0 179000.0 265400.00000000006 ;
      RECT  185000.0 264600.0 185800.0 265400.00000000006 ;
      RECT  185000.0 264600.0 185800.0 265400.00000000006 ;
      RECT  191800.0 264600.0 192600.00000000003 265400.00000000006 ;
      RECT  179800.0 122000.0 180600.00000000003 271000.0 ;
      RECT  183400.0 122800.00000000001 184200.0 271800.0 ;
      RECT  186600.00000000003 122000.0 187400.0 271000.0 ;
      RECT  190200.0 122800.00000000001 191000.0 271800.0 ;
      RECT  181400.0 112000.00000000001 182200.0 112800.00000000001 ;
      RECT  181400.0 112000.00000000001 182200.0 112800.00000000001 ;
      RECT  179800.0 112000.00000000001 180600.00000000003 112800.00000000001 ;
      RECT  179800.0 107200.0 180600.00000000003 108000.00000000001 ;
      RECT  183400.0 112000.00000000001 184200.0 112800.00000000001 ;
      RECT  183400.0 107200.0 184200.0 108000.00000000001 ;
      RECT  179900.0 105600.00000000001 180500.0 118200.0 ;
      RECT  183500.0 105600.00000000001 184100.00000000003 118200.0 ;
      RECT  188200.0 112000.00000000001 189000.0 112800.00000000001 ;
      RECT  188200.0 112000.00000000001 189000.0 112800.00000000001 ;
      RECT  186600.00000000003 112000.00000000001 187400.0 112800.00000000001 ;
      RECT  186600.00000000003 107200.0 187400.0 108000.00000000001 ;
      RECT  190200.0 112000.00000000001 191000.0 112800.00000000001 ;
      RECT  190200.0 107200.0 191000.0 108000.00000000001 ;
      RECT  186700.0 105600.00000000001 187300.0 118200.0 ;
      RECT  190300.0 105600.00000000001 190900.0 118200.0 ;
      RECT  179900.0 105600.00000000001 180500.0 118200.0 ;
      RECT  183500.0 105600.00000000001 184100.00000000003 118200.0 ;
      RECT  186700.0 105600.00000000001 187300.0 118200.0 ;
      RECT  190300.0 105600.00000000001 190900.0 118200.0 ;
      RECT  178600.00000000003 68800.00000000001 185400.0 101400.0 ;
      RECT  185400.0 68800.00000000001 192200.0 101400.0 ;
      RECT  185000.0 95000.00000000001 185800.0 95800.00000000001 ;
      RECT  184000.0 81600.00000000001 184800.0 82400.0 ;
      RECT  191800.0 95000.00000000001 192600.00000000003 95800.00000000001 ;
      RECT  190800.0 81600.00000000001 191600.00000000003 82400.0 ;
      RECT  179200.0 68800.00000000001 180000.0 71800.00000000001 ;
      RECT  180600.00000000003 78400.0 181400.0 101400.0 ;
      RECT  182600.00000000003 78400.0 183400.0 101400.0 ;
      RECT  186000.0 68800.00000000001 186800.0 71800.00000000001 ;
      RECT  187400.0 78400.0 188200.0 101400.0 ;
      RECT  189400.0 78400.0 190200.0 101400.0 ;
      RECT  178600.00000000003 24200.000000000004 185400.0 64599.99999999999 ;
      RECT  185400.0 24200.000000000004 192200.0 64599.99999999999 ;
      RECT  182400.0 30400.000000000004 183200.0 31200.000000000004 ;
      RECT  181800.0 47800.00000000001 182600.00000000003 48600.00000000001 ;
      RECT  182400.0 37000.0 183200.0 37800.00000000001 ;
      RECT  183800.0 41400.00000000001 184600.00000000003 42200.0 ;
      RECT  183200.0 54800.00000000001 184000.0 55600.00000000001 ;
      RECT  189200.0 30400.000000000004 190000.0 31200.000000000004 ;
      RECT  188600.00000000003 47800.00000000001 189400.0 48600.00000000001 ;
      RECT  189200.0 37000.0 190000.0 37800.00000000001 ;
      RECT  190600.00000000003 41400.00000000001 191400.0 42200.0 ;
      RECT  190000.0 54800.00000000001 190800.0 55600.00000000001 ;
      RECT  181600.00000000003 24200.000000000004 182400.0 26200.000000000004 ;
      RECT  188400.0 24200.000000000004 189200.0 26200.000000000004 ;
      RECT  180600.00000000003 62600.00000000001 181400.0 64600.00000000001 ;
      RECT  182600.00000000003 59600.0 183400.0 64600.00000000001 ;
      RECT  187400.0 62600.00000000001 188200.0 64600.00000000001 ;
      RECT  189400.0 59600.0 190200.0 64600.00000000001 ;
      RECT  111400.0 127500.0 112000.0 131800.0 ;
      RECT  111400.0 137100.00000000003 112000.0 141400.0 ;
      RECT  111400.0 145900.0 112000.0 150200.0 ;
      RECT  111400.0 155500.0 112000.0 159800.0 ;
      RECT  111400.0 164300.0 112000.0 168600.00000000003 ;
      RECT  111400.0 173899.99999999997 112000.0 178200.0 ;
      RECT  111400.0 182700.0 112000.0 187000.0 ;
      RECT  111400.0 192300.0 112000.0 196600.00000000003 ;
      RECT  92900.0 124000.0 93500.0 159600.00000000003 ;
      RECT  94300.0 124000.0 94900.0 159600.00000000003 ;
      RECT  95700.0 124000.0 96300.0 159600.00000000003 ;
      RECT  97100.0 124000.0 97700.0 159600.00000000003 ;
      RECT  101400.0 127300.00000000001 102000.0 127900.0 ;
      RECT  103000.0 127300.00000000001 103600.0 127900.0 ;
      RECT  101400.0 127600.00000000001 102000.0 129900.0 ;
      RECT  101700.0 127300.00000000001 103300.0 127900.0 ;
      RECT  103000.0 124900.0 103600.0 127600.00000000001 ;
      RECT  101300.0 129900.0 102100.0 130699.99999999999 ;
      RECT  102900.0 124100.00000000001 103700.0 124900.0 ;
      RECT  103700.0 127200.0 102900.0 128000.0 ;
      RECT  101400.0 136700.0 102000.0 136100.00000000003 ;
      RECT  103000.0 136700.0 103600.0 136100.00000000003 ;
      RECT  101400.0 136400.0 102000.0 134100.00000000003 ;
      RECT  101700.0 136700.0 103300.0 136100.00000000003 ;
      RECT  103000.0 139100.00000000003 103600.0 136400.0 ;
      RECT  101300.0 134100.00000000003 102100.0 133300.0 ;
      RECT  102900.0 139900.0 103700.0 139100.00000000003 ;
      RECT  103700.0 136800.0 102900.0 136000.0 ;
      RECT  101400.0 145700.0 102000.0 146300.0 ;
      RECT  103000.0 145700.0 103600.0 146300.0 ;
      RECT  101400.0 146000.0 102000.0 148300.0 ;
      RECT  101700.0 145700.0 103300.0 146300.0 ;
      RECT  103000.0 143300.0 103600.0 146000.0 ;
      RECT  101300.0 148300.0 102100.0 149100.00000000003 ;
      RECT  102900.0 142500.0 103700.0 143300.0 ;
      RECT  103700.0 145600.00000000003 102900.0 146400.0 ;
      RECT  101400.0 155100.00000000003 102000.0 154500.0 ;
      RECT  103000.0 155100.00000000003 103600.0 154500.0 ;
      RECT  101400.0 154800.0 102000.0 152500.0 ;
      RECT  101700.0 155100.00000000003 103300.0 154500.0 ;
      RECT  103000.0 157500.0 103600.0 154800.0 ;
      RECT  101300.0 152500.0 102100.0 151700.0 ;
      RECT  102900.0 158300.0 103700.0 157500.0 ;
      RECT  103700.0 155200.0 102900.0 154400.00000000003 ;
      RECT  93600.0 129800.00000000001 92800.0 130600.00000000003 ;
      RECT  81900.0 126800.00000000001 81100.0 127600.00000000001 ;
      RECT  95000.0 139000.0 94200.0 139800.0 ;
      RECT  83300.0 136400.0 82500.0 137200.0 ;
      RECT  81900.0 142200.0 81100.0 143000.0 ;
      RECT  96400.0 142200.0 95600.0 143000.0 ;
      RECT  83300.0 151400.0 82500.0 152200.0 ;
      RECT  97800.0 151400.0 97000.0 152200.0 ;
      RECT  93600.0 127200.0 92800.0 128000.0 ;
      RECT  95000.0 125800.00000000001 94200.0 126600.00000000001 ;
      RECT  96400.0 136000.0 95600.0 136800.0 ;
      RECT  95000.0 137400.0 94200.0 138200.0 ;
      RECT  93600.0 145600.00000000003 92800.0 146400.0 ;
      RECT  97800.0 144200.0 97000.0 145000.0 ;
      RECT  96400.0 154399.99999999997 95600.0 155200.0 ;
      RECT  97800.0 155800.0 97000.0 156600.00000000003 ;
      RECT  90500.0 131600.00000000003 89700.0 132400.0 ;
      RECT  90500.0 131600.00000000003 89700.0 132400.0 ;
      RECT  108500.0 131600.00000000003 107700.0 132400.0 ;
      RECT  108500.0 131600.00000000003 107700.0 132400.0 ;
      RECT  90500.0 122400.0 89700.0 123200.0 ;
      RECT  90500.0 122400.0 89700.0 123200.0 ;
      RECT  108500.0 122400.0 107700.0 123200.0 ;
      RECT  108500.0 122400.0 107700.0 123200.0 ;
      RECT  90500.0 131600.00000000003 89700.0 132400.0 ;
      RECT  90500.0 131600.00000000003 89700.0 132400.0 ;
      RECT  108500.0 131600.00000000003 107700.0 132400.0 ;
      RECT  108500.0 131600.00000000003 107700.0 132400.0 ;
      RECT  90500.0 140800.0 89700.0 141600.00000000003 ;
      RECT  90500.0 140800.0 89700.0 141600.00000000003 ;
      RECT  108500.0 140800.0 107700.0 141600.00000000003 ;
      RECT  108500.0 140800.0 107700.0 141600.00000000003 ;
      RECT  90500.0 150000.0 89700.0 150800.0 ;
      RECT  90500.0 150000.0 89700.0 150800.0 ;
      RECT  108500.0 150000.0 107700.0 150800.0 ;
      RECT  108500.0 150000.0 107700.0 150800.0 ;
      RECT  90500.0 140800.0 89700.0 141600.00000000003 ;
      RECT  90500.0 140800.0 89700.0 141600.00000000003 ;
      RECT  108500.0 140800.0 107700.0 141600.00000000003 ;
      RECT  108500.0 140800.0 107700.0 141600.00000000003 ;
      RECT  90500.0 150000.0 89700.0 150800.0 ;
      RECT  90500.0 150000.0 89700.0 150800.0 ;
      RECT  108500.0 150000.0 107700.0 150800.0 ;
      RECT  108500.0 150000.0 107700.0 150800.0 ;
      RECT  90500.0 159200.0 89700.0 160000.0 ;
      RECT  90500.0 159200.0 89700.0 160000.0 ;
      RECT  108500.0 159200.0 107700.0 160000.0 ;
      RECT  108500.0 159200.0 107700.0 160000.0 ;
      RECT  81200.0 124000.0 81800.0 159600.00000000003 ;
      RECT  82600.0 124000.0 83200.0 159600.00000000003 ;
      RECT  92900.0 160800.0 93500.0 196399.99999999997 ;
      RECT  94300.0 160800.0 94900.0 196399.99999999997 ;
      RECT  95700.0 160800.0 96300.0 196399.99999999997 ;
      RECT  97100.0 160800.0 97700.0 196399.99999999997 ;
      RECT  101400.0 164100.00000000003 102000.0 164700.0 ;
      RECT  103000.0 164100.00000000003 103600.0 164700.0 ;
      RECT  101400.0 164399.99999999997 102000.0 166700.0 ;
      RECT  101700.0 164100.00000000003 103300.0 164700.0 ;
      RECT  103000.0 161700.0 103600.0 164399.99999999997 ;
      RECT  101300.0 166700.0 102100.0 167500.0 ;
      RECT  102900.0 160899.99999999997 103700.0 161700.0 ;
      RECT  103700.0 164000.0 102900.0 164800.0 ;
      RECT  101400.0 173500.0 102000.0 172900.00000000003 ;
      RECT  103000.0 173500.0 103600.0 172900.00000000003 ;
      RECT  101400.0 173200.0 102000.0 170899.99999999997 ;
      RECT  101700.0 173500.0 103300.0 172900.00000000003 ;
      RECT  103000.0 175899.99999999997 103600.0 173200.0 ;
      RECT  101300.0 170899.99999999997 102100.0 170100.00000000003 ;
      RECT  102900.0 176700.0 103700.0 175899.99999999997 ;
      RECT  103700.0 173600.00000000003 102900.0 172800.0 ;
      RECT  101400.0 182500.0 102000.0 183100.00000000003 ;
      RECT  103000.0 182500.0 103600.0 183100.00000000003 ;
      RECT  101400.0 182800.0 102000.0 185100.00000000003 ;
      RECT  101700.0 182500.0 103300.0 183100.00000000003 ;
      RECT  103000.0 180100.00000000003 103600.0 182800.0 ;
      RECT  101300.0 185100.00000000003 102100.0 185900.00000000003 ;
      RECT  102900.0 179300.0 103700.0 180100.00000000003 ;
      RECT  103700.0 182400.00000000003 102900.0 183200.0 ;
      RECT  101400.0 191899.99999999997 102000.0 191300.0 ;
      RECT  103000.0 191899.99999999997 103600.0 191300.0 ;
      RECT  101400.0 191600.00000000003 102000.0 189300.0 ;
      RECT  101700.0 191899.99999999997 103300.0 191300.0 ;
      RECT  103000.0 194300.0 103600.0 191600.00000000003 ;
      RECT  101300.0 189300.0 102100.0 188500.0 ;
      RECT  102900.0 195100.00000000003 103700.0 194300.0 ;
      RECT  103700.0 192000.0 102900.0 191200.0 ;
      RECT  93600.0 166600.00000000003 92800.0 167399.99999999997 ;
      RECT  81900.0 163600.00000000003 81100.0 164399.99999999997 ;
      RECT  95000.0 175800.0 94200.0 176600.00000000003 ;
      RECT  83300.0 173200.0 82500.0 174000.0 ;
      RECT  81900.0 179000.0 81100.0 179800.0 ;
      RECT  96400.0 179000.0 95600.0 179800.0 ;
      RECT  83300.0 188200.0 82500.0 189000.0 ;
      RECT  97800.0 188200.0 97000.0 189000.0 ;
      RECT  93600.0 164000.0 92800.0 164800.0 ;
      RECT  95000.0 162600.00000000003 94200.0 163399.99999999997 ;
      RECT  96400.0 172800.0 95600.0 173600.00000000003 ;
      RECT  95000.0 174200.0 94200.0 175000.0 ;
      RECT  93600.0 182399.99999999997 92800.0 183200.0 ;
      RECT  97800.0 181000.0 97000.0 181800.0 ;
      RECT  96400.0 191200.0 95600.0 192000.0 ;
      RECT  97800.0 192600.00000000003 97000.0 193399.99999999997 ;
      RECT  90500.0 168399.99999999997 89700.0 169200.0 ;
      RECT  90500.0 168399.99999999997 89700.0 169200.0 ;
      RECT  108500.0 168399.99999999997 107700.0 169200.0 ;
      RECT  108500.0 168399.99999999997 107700.0 169200.0 ;
      RECT  90500.0 159200.0 89700.0 160000.0 ;
      RECT  90500.0 159200.0 89700.0 160000.0 ;
      RECT  108500.0 159200.0 107700.0 160000.0 ;
      RECT  108500.0 159200.0 107700.0 160000.0 ;
      RECT  90500.0 168399.99999999997 89700.0 169200.0 ;
      RECT  90500.0 168399.99999999997 89700.0 169200.0 ;
      RECT  108500.0 168399.99999999997 107700.0 169200.0 ;
      RECT  108500.0 168399.99999999997 107700.0 169200.0 ;
      RECT  90500.0 177600.00000000003 89700.0 178399.99999999997 ;
      RECT  90500.0 177600.00000000003 89700.0 178399.99999999997 ;
      RECT  108500.0 177600.00000000003 107700.0 178399.99999999997 ;
      RECT  108500.0 177600.00000000003 107700.0 178399.99999999997 ;
      RECT  90500.0 186800.0 89700.0 187600.00000000003 ;
      RECT  90500.0 186800.0 89700.0 187600.00000000003 ;
      RECT  108500.0 186800.0 107700.0 187600.00000000003 ;
      RECT  108500.0 186800.0 107700.0 187600.00000000003 ;
      RECT  90500.0 177600.00000000003 89700.0 178399.99999999997 ;
      RECT  90500.0 177600.00000000003 89700.0 178399.99999999997 ;
      RECT  108500.0 177600.00000000003 107700.0 178399.99999999997 ;
      RECT  108500.0 177600.00000000003 107700.0 178399.99999999997 ;
      RECT  90500.0 186800.0 89700.0 187600.00000000003 ;
      RECT  90500.0 186800.0 89700.0 187600.00000000003 ;
      RECT  108500.0 186800.0 107700.0 187600.00000000003 ;
      RECT  108500.0 186800.0 107700.0 187600.00000000003 ;
      RECT  90500.0 196000.0 89700.0 196800.0 ;
      RECT  90500.0 196000.0 89700.0 196800.0 ;
      RECT  108500.0 196000.0 107700.0 196800.0 ;
      RECT  108500.0 196000.0 107700.0 196800.0 ;
      RECT  81200.0 160800.0 81800.0 196399.99999999997 ;
      RECT  82600.0 160800.0 83200.0 196399.99999999997 ;
      RECT  128600.0 127300.00000000001 129199.99999999999 127900.0 ;
      RECT  130199.99999999999 127300.00000000001 130800.00000000001 127900.0 ;
      RECT  128600.0 127600.00000000001 129199.99999999999 129900.0 ;
      RECT  128900.0 127300.00000000001 130500.0 127900.0 ;
      RECT  130199.99999999999 124900.0 130800.00000000001 127600.00000000001 ;
      RECT  128500.0 129900.0 129300.00000000001 130699.99999999999 ;
      RECT  130100.0 124100.00000000001 130900.0 124900.0 ;
      RECT  130900.0 127200.0 130100.0 128000.0 ;
      RECT  128600.0 136700.0 129199.99999999999 136100.00000000003 ;
      RECT  130199.99999999999 136700.0 130800.00000000001 136100.00000000003 ;
      RECT  128600.0 136400.0 129199.99999999999 134100.00000000003 ;
      RECT  128900.0 136700.0 130500.0 136100.00000000003 ;
      RECT  130199.99999999999 139100.00000000003 130800.00000000001 136400.0 ;
      RECT  128500.0 134100.00000000003 129300.00000000001 133300.0 ;
      RECT  130100.0 139900.0 130900.0 139100.00000000003 ;
      RECT  130900.0 136800.0 130100.0 136000.0 ;
      RECT  128600.0 145700.0 129199.99999999999 146300.0 ;
      RECT  130199.99999999999 145700.0 130800.00000000001 146300.0 ;
      RECT  128600.0 146000.0 129199.99999999999 148300.0 ;
      RECT  128900.0 145700.0 130500.0 146300.0 ;
      RECT  130199.99999999999 143300.0 130800.00000000001 146000.0 ;
      RECT  128500.0 148300.0 129300.00000000001 149100.00000000003 ;
      RECT  130100.0 142500.0 130900.0 143300.0 ;
      RECT  130900.0 145600.00000000003 130100.0 146400.0 ;
      RECT  128600.0 155100.00000000003 129199.99999999999 154500.0 ;
      RECT  130199.99999999999 155100.00000000003 130800.00000000001 154500.0 ;
      RECT  128600.0 154800.0 129199.99999999999 152500.0 ;
      RECT  128900.0 155100.00000000003 130500.0 154500.0 ;
      RECT  130199.99999999999 157500.0 130800.00000000001 154800.0 ;
      RECT  128500.0 152500.0 129300.00000000001 151700.0 ;
      RECT  130100.0 158300.0 130900.0 157500.0 ;
      RECT  130900.0 155200.0 130100.0 154399.99999999997 ;
      RECT  128600.0 164100.00000000003 129199.99999999999 164700.0 ;
      RECT  130199.99999999999 164100.00000000003 130800.00000000001 164700.0 ;
      RECT  128600.0 164399.99999999997 129199.99999999999 166700.0 ;
      RECT  128900.0 164100.00000000003 130500.0 164700.0 ;
      RECT  130199.99999999999 161700.0 130800.00000000001 164399.99999999997 ;
      RECT  128500.0 166700.0 129300.00000000001 167500.0 ;
      RECT  130100.0 160899.99999999997 130900.0 161700.0 ;
      RECT  130900.0 164000.0 130100.0 164800.0 ;
      RECT  128600.0 173500.0 129199.99999999999 172899.99999999997 ;
      RECT  130199.99999999999 173500.0 130800.00000000001 172899.99999999997 ;
      RECT  128600.0 173200.0 129199.99999999999 170899.99999999997 ;
      RECT  128900.0 173500.0 130500.0 172899.99999999997 ;
      RECT  130199.99999999999 175899.99999999997 130800.00000000001 173200.0 ;
      RECT  128500.0 170899.99999999997 129300.00000000001 170100.00000000003 ;
      RECT  130100.0 176700.0 130900.0 175899.99999999997 ;
      RECT  130900.0 173600.00000000003 130100.0 172800.0 ;
      RECT  128600.0 182500.0 129199.99999999999 183100.00000000003 ;
      RECT  130199.99999999999 182500.0 130800.00000000001 183100.00000000003 ;
      RECT  128600.0 182800.0 129199.99999999999 185100.00000000003 ;
      RECT  128900.0 182500.0 130500.0 183100.00000000003 ;
      RECT  130199.99999999999 180100.00000000003 130800.00000000001 182800.0 ;
      RECT  128500.0 185100.00000000003 129300.00000000001 185899.99999999997 ;
      RECT  130100.0 179300.0 130900.0 180100.00000000003 ;
      RECT  130900.0 182399.99999999997 130100.0 183200.0 ;
      RECT  128600.0 191900.00000000003 129199.99999999999 191300.0 ;
      RECT  130199.99999999999 191900.00000000003 130800.00000000001 191300.0 ;
      RECT  128600.0 191600.00000000003 129199.99999999999 189300.0 ;
      RECT  128900.0 191900.00000000003 130500.0 191300.0 ;
      RECT  130199.99999999999 194300.0 130800.00000000001 191600.00000000003 ;
      RECT  128500.0 189300.0 129300.00000000001 188500.0 ;
      RECT  130100.0 195100.00000000003 130900.0 194300.0 ;
      RECT  130900.0 192000.0 130100.0 191200.0 ;
      RECT  128600.0 200900.00000000003 129199.99999999999 201500.0 ;
      RECT  130199.99999999999 200900.00000000003 130800.00000000001 201500.0 ;
      RECT  128600.0 201200.0 129199.99999999999 203500.0 ;
      RECT  128900.0 200900.00000000003 130500.0 201500.0 ;
      RECT  130199.99999999999 198500.0 130800.00000000001 201200.0 ;
      RECT  128500.0 203500.0 129300.00000000001 204300.0 ;
      RECT  130100.0 197700.0 130900.0 198500.0 ;
      RECT  130900.0 200800.0 130100.0 201600.00000000003 ;
      RECT  128600.0 210300.0 129199.99999999999 209700.0 ;
      RECT  130199.99999999999 210300.0 130800.00000000001 209700.0 ;
      RECT  128600.0 210000.0 129199.99999999999 207700.0 ;
      RECT  128900.0 210300.0 130500.0 209700.0 ;
      RECT  130199.99999999999 212700.0 130800.00000000001 210000.0 ;
      RECT  128500.0 207700.0 129300.00000000001 206899.99999999997 ;
      RECT  130100.0 213500.0 130900.0 212700.0 ;
      RECT  130900.0 210399.99999999997 130100.0 209600.00000000003 ;
      RECT  128600.0 219300.0 129199.99999999999 219899.99999999997 ;
      RECT  130199.99999999999 219300.0 130800.00000000001 219899.99999999997 ;
      RECT  128600.0 219600.00000000003 129199.99999999999 221899.99999999997 ;
      RECT  128900.0 219300.0 130500.0 219899.99999999997 ;
      RECT  130199.99999999999 216899.99999999997 130800.00000000001 219600.00000000003 ;
      RECT  128500.0 221899.99999999997 129300.00000000001 222700.0 ;
      RECT  130100.0 216100.00000000003 130900.0 216899.99999999997 ;
      RECT  130900.0 219200.0 130100.0 220000.0 ;
      RECT  128600.0 228700.0 129199.99999999999 228100.00000000003 ;
      RECT  130199.99999999999 228700.0 130800.00000000001 228100.00000000003 ;
      RECT  128600.0 228400.00000000003 129199.99999999999 226100.00000000003 ;
      RECT  128900.0 228700.0 130500.0 228100.00000000003 ;
      RECT  130199.99999999999 231100.00000000003 130800.00000000001 228400.00000000003 ;
      RECT  128500.0 226100.00000000003 129300.00000000001 225300.0 ;
      RECT  130100.0 231900.00000000003 130900.0 231100.00000000003 ;
      RECT  130900.0 228800.0 130100.0 228000.0 ;
      RECT  128600.0 237700.0 129199.99999999999 238300.0 ;
      RECT  130199.99999999999 237700.0 130800.00000000001 238300.0 ;
      RECT  128600.0 238000.0 129199.99999999999 240300.0 ;
      RECT  128900.0 237700.0 130500.0 238300.0 ;
      RECT  130199.99999999999 235300.0 130800.00000000001 238000.0 ;
      RECT  128500.0 240300.0 129300.00000000001 241100.00000000003 ;
      RECT  130100.0 234500.0 130900.0 235300.0 ;
      RECT  130900.0 237600.00000000003 130100.0 238400.00000000003 ;
      RECT  128600.0 247100.00000000003 129199.99999999999 246500.0 ;
      RECT  130199.99999999999 247100.00000000003 130800.00000000001 246500.0 ;
      RECT  128600.0 246800.0 129199.99999999999 244500.0 ;
      RECT  128900.0 247100.00000000003 130500.0 246500.0 ;
      RECT  130199.99999999999 249500.0 130800.00000000001 246800.0 ;
      RECT  128500.0 244500.0 129300.00000000001 243700.0 ;
      RECT  130100.0 250300.0 130900.0 249500.0 ;
      RECT  130900.0 247200.0 130100.0 246400.00000000003 ;
      RECT  128600.0 256100.00000000003 129199.99999999999 256700.0 ;
      RECT  130199.99999999999 256100.00000000003 130800.00000000001 256700.0 ;
      RECT  128600.0 256400.00000000003 129199.99999999999 258700.0 ;
      RECT  128900.0 256100.00000000003 130500.0 256700.0 ;
      RECT  130199.99999999999 253700.0 130800.00000000001 256400.00000000003 ;
      RECT  128500.0 258700.0 129300.00000000001 259500.0 ;
      RECT  130100.0 252900.00000000003 130900.0 253700.0 ;
      RECT  130900.0 256000.0 130100.0 256800.0 ;
      RECT  128600.0 265500.0 129199.99999999999 264900.00000000006 ;
      RECT  130199.99999999999 265500.0 130800.00000000001 264900.00000000006 ;
      RECT  128600.0 265200.0 129199.99999999999 262900.00000000006 ;
      RECT  128900.0 265500.0 130500.0 264900.00000000006 ;
      RECT  130199.99999999999 267900.00000000006 130800.00000000001 265200.0 ;
      RECT  128500.0 262900.00000000006 129300.00000000001 262100.00000000003 ;
      RECT  130100.0 268700.0 130900.0 267900.00000000006 ;
      RECT  130900.0 265600.0 130100.0 264800.0 ;
      RECT  81900.0 132800.0 81100.0 133600.00000000003 ;
      RECT  74600.0 132800.0 73800.0 133600.00000000003 ;
      RECT  83300.0 142000.0 82500.0 142800.0 ;
      RECT  76000.0 142000.0 75200.0 142800.0 ;
      RECT  81900.0 169600.00000000003 81100.0 170399.99999999997 ;
      RECT  77400.0 169600.00000000003 76600.0 170399.99999999997 ;
      RECT  83300.0 178800.0 82500.0 179600.00000000003 ;
      RECT  78800.0 178800.0 78000.0 179600.00000000003 ;
      RECT  112100.0 126800.00000000001 111300.00000000001 127600.00000000001 ;
      RECT  112100.0 131400.0 111300.00000000001 132200.0 ;
      RECT  115500.0 131400.0 114700.0 132200.0 ;
      RECT  112100.0 136400.0 111300.00000000001 137200.0 ;
      RECT  112100.0 141000.0 111300.00000000001 141800.0 ;
      RECT  116900.0 141000.0 116100.0 141800.0 ;
      RECT  112100.0 145200.0 111300.00000000001 146000.0 ;
      RECT  112100.0 149800.0 111300.00000000001 150600.00000000003 ;
      RECT  118300.0 149800.0 117500.0 150600.00000000003 ;
      RECT  112100.0 154800.0 111300.00000000001 155600.00000000003 ;
      RECT  112100.0 159399.99999999997 111300.00000000001 160200.0 ;
      RECT  119700.0 159399.99999999997 118900.0 160200.0 ;
      RECT  112100.0 163600.00000000003 111300.00000000001 164399.99999999997 ;
      RECT  112100.0 168200.0 111300.00000000001 169000.0 ;
      RECT  121100.0 168200.0 120300.00000000001 169000.0 ;
      RECT  112100.0 173200.0 111300.00000000001 174000.0 ;
      RECT  112100.0 177800.0 111300.00000000001 178600.00000000003 ;
      RECT  122500.0 177800.0 121700.0 178600.00000000003 ;
      RECT  112100.0 182000.0 111300.00000000001 182800.0 ;
      RECT  112100.0 186600.00000000003 111300.00000000001 187399.99999999997 ;
      RECT  123900.0 186600.00000000003 123100.0 187399.99999999997 ;
      RECT  112100.0 191600.00000000003 111300.00000000001 192399.99999999997 ;
      RECT  112100.0 196200.0 111300.00000000001 197000.0 ;
      RECT  125300.0 196200.0 124500.0 197000.0 ;
      RECT  115500.0 127200.0 114700.0 128000.0 ;
      RECT  121100.0 125800.00000000001 120300.00000000001 126600.00000000001 ;
      RECT  115500.0 136000.0 114700.0 136800.0 ;
      RECT  122500.0 137400.0 121700.0 138200.0 ;
      RECT  115500.0 145600.00000000003 114700.0 146400.0 ;
      RECT  123900.0 144200.0 123100.0 145000.0 ;
      RECT  115500.0 154399.99999999997 114700.0 155200.0 ;
      RECT  125300.0 155800.0 124500.0 156600.00000000003 ;
      RECT  116900.0 164000.0 116100.0 164800.0 ;
      RECT  121100.0 162600.00000000003 120300.00000000001 163399.99999999997 ;
      RECT  116900.0 172800.0 116100.0 173600.00000000003 ;
      RECT  122500.0 174200.0 121700.0 175000.0 ;
      RECT  116900.0 182399.99999999997 116100.0 183200.0 ;
      RECT  123900.0 181000.0 123100.0 181800.0 ;
      RECT  116900.0 191200.0 116100.0 192000.0 ;
      RECT  125300.0 192600.00000000003 124500.0 193399.99999999997 ;
      RECT  118300.0 200800.0 117500.0 201600.00000000003 ;
      RECT  121100.0 199400.00000000003 120300.00000000001 200200.0 ;
      RECT  118300.0 209600.00000000003 117500.0 210400.00000000003 ;
      RECT  122500.0 211000.0 121700.0 211800.0 ;
      RECT  118300.0 219200.0 117500.0 220000.0 ;
      RECT  123900.0 217800.0 123100.0 218600.00000000003 ;
      RECT  118300.0 228000.0 117500.0 228800.0 ;
      RECT  125300.0 229400.00000000003 124500.0 230200.0 ;
      RECT  119700.0 237600.00000000003 118900.0 238400.00000000003 ;
      RECT  121100.0 236200.0 120300.00000000001 237000.0 ;
      RECT  119700.0 246400.00000000003 118900.0 247200.0 ;
      RECT  122500.0 247800.0 121700.0 248600.00000000003 ;
      RECT  119700.0 256000.0 118900.0 256800.0 ;
      RECT  123900.0 254600.00000000003 123100.0 255400.00000000003 ;
      RECT  119700.0 264800.0 118900.0 265600.0 ;
      RECT  125300.0 266200.0 124500.0 267000.0 ;
      RECT  130900.0 131600.00000000003 130100.00000000003 132400.0 ;
      RECT  130900.0 131600.00000000003 130100.00000000003 132400.0 ;
      RECT  130900.0 122400.0 130100.00000000003 123200.0 ;
      RECT  130900.0 122400.0 130100.00000000003 123200.0 ;
      RECT  130900.0 131600.00000000003 130100.00000000003 132400.0 ;
      RECT  130900.0 131600.00000000003 130100.00000000003 132400.0 ;
      RECT  130900.0 140800.0 130100.00000000003 141600.00000000003 ;
      RECT  130900.0 140800.0 130100.00000000003 141600.00000000003 ;
      RECT  130900.0 150000.0 130100.00000000003 150800.0 ;
      RECT  130900.0 150000.0 130100.00000000003 150800.0 ;
      RECT  130900.0 140800.0 130100.00000000003 141600.00000000003 ;
      RECT  130900.0 140800.0 130100.00000000003 141600.00000000003 ;
      RECT  130900.0 150000.0 130100.00000000003 150800.0 ;
      RECT  130900.0 150000.0 130100.00000000003 150800.0 ;
      RECT  130900.0 159200.0 130100.00000000003 160000.0 ;
      RECT  130900.0 159200.0 130100.00000000003 160000.0 ;
      RECT  130900.0 168399.99999999997 130100.00000000003 169200.0 ;
      RECT  130900.0 168399.99999999997 130100.00000000003 169200.0 ;
      RECT  130900.0 159200.0 130100.00000000003 160000.0 ;
      RECT  130900.0 159200.0 130100.00000000003 160000.0 ;
      RECT  130900.0 168399.99999999997 130100.00000000003 169200.0 ;
      RECT  130900.0 168399.99999999997 130100.00000000003 169200.0 ;
      RECT  130900.0 177600.00000000003 130100.00000000003 178399.99999999997 ;
      RECT  130900.0 177600.00000000003 130100.00000000003 178399.99999999997 ;
      RECT  130900.0 186800.0 130100.00000000003 187600.00000000003 ;
      RECT  130900.0 186800.0 130100.00000000003 187600.00000000003 ;
      RECT  130900.0 177600.00000000003 130100.00000000003 178399.99999999997 ;
      RECT  130900.0 177600.00000000003 130100.00000000003 178399.99999999997 ;
      RECT  130900.0 186800.0 130100.00000000003 187600.00000000003 ;
      RECT  130900.0 186800.0 130100.00000000003 187600.00000000003 ;
      RECT  130900.0 196000.0 130100.00000000003 196800.0 ;
      RECT  130900.0 196000.0 130100.00000000003 196800.0 ;
      RECT  130900.0 205200.0 130100.00000000003 206000.0 ;
      RECT  130900.0 205200.0 130100.00000000003 206000.0 ;
      RECT  130900.0 196000.0 130100.00000000003 196800.0 ;
      RECT  130900.0 196000.0 130100.00000000003 196800.0 ;
      RECT  130900.0 205200.0 130100.00000000003 206000.0 ;
      RECT  130900.0 205200.0 130100.00000000003 206000.0 ;
      RECT  130900.0 214400.00000000003 130100.00000000003 215200.0 ;
      RECT  130900.0 214400.00000000003 130100.00000000003 215200.0 ;
      RECT  130900.0 223600.00000000003 130100.00000000003 224400.00000000003 ;
      RECT  130900.0 223600.00000000003 130100.00000000003 224400.00000000003 ;
      RECT  130900.0 214400.00000000003 130100.00000000003 215200.0 ;
      RECT  130900.0 214400.00000000003 130100.00000000003 215200.0 ;
      RECT  130900.0 223600.00000000003 130100.00000000003 224400.00000000003 ;
      RECT  130900.0 223600.00000000003 130100.00000000003 224400.00000000003 ;
      RECT  130900.0 232800.0 130100.00000000003 233600.00000000003 ;
      RECT  130900.0 232800.0 130100.00000000003 233600.00000000003 ;
      RECT  130900.0 242000.0 130100.00000000003 242800.0 ;
      RECT  130900.0 242000.0 130100.00000000003 242800.0 ;
      RECT  130900.0 232800.0 130100.00000000003 233600.00000000003 ;
      RECT  130900.0 232800.0 130100.00000000003 233600.00000000003 ;
      RECT  130900.0 242000.0 130100.00000000003 242800.0 ;
      RECT  130900.0 242000.0 130100.00000000003 242800.0 ;
      RECT  130900.0 251200.0 130100.00000000003 252000.0 ;
      RECT  130900.0 251200.0 130100.00000000003 252000.0 ;
      RECT  130900.0 260399.99999999997 130100.00000000003 261200.0 ;
      RECT  130900.0 260399.99999999997 130100.00000000003 261200.0 ;
      RECT  130900.0 251200.0 130100.00000000003 252000.0 ;
      RECT  130900.0 251200.0 130100.00000000003 252000.0 ;
      RECT  130900.0 260399.99999999997 130100.00000000003 261200.0 ;
      RECT  130900.0 260399.99999999997 130100.00000000003 261200.0 ;
      RECT  130900.0 269600.0 130100.00000000003 270400.00000000006 ;
      RECT  130900.0 269600.0 130100.00000000003 270400.00000000006 ;
      RECT  73900.0 122800.00000000001 74500.0 196400.00000000003 ;
      RECT  75300.0 122800.00000000001 75900.0 196400.00000000003 ;
      RECT  76699.99999999999 122800.00000000001 77300.0 196400.00000000003 ;
      RECT  78100.0 122800.00000000001 78699.99999999999 196400.00000000003 ;
      RECT  147200.0 125900.0 147800.0 126500.0 ;
      RECT  147200.0 125600.00000000001 147800.0 126200.0 ;
      RECT  147500.0 125900.0 158300.0 126500.0 ;
      RECT  147200.0 137500.0 147800.0 138100.00000000003 ;
      RECT  147200.0 137800.0 147800.0 138400.0 ;
      RECT  147500.0 137500.0 158300.0 138100.00000000003 ;
      RECT  147200.0 144300.0 147800.0 144900.0 ;
      RECT  147200.0 144000.0 147800.0 144600.00000000003 ;
      RECT  147500.0 144300.0 158300.0 144900.0 ;
      RECT  147200.0 155899.99999999997 147800.0 156500.0 ;
      RECT  147200.0 156200.0 147800.0 156800.0 ;
      RECT  147500.0 155899.99999999997 158300.0 156500.0 ;
      RECT  147200.0 162700.0 147800.0 163300.0 ;
      RECT  147200.0 162399.99999999997 147800.0 163000.0 ;
      RECT  147500.0 162700.0 158300.0 163300.0 ;
      RECT  147200.0 174300.0 147800.0 174899.99999999997 ;
      RECT  147200.0 174600.00000000003 147800.0 175200.0 ;
      RECT  147500.0 174300.0 158300.0 174899.99999999997 ;
      RECT  147200.0 181100.00000000003 147800.0 181700.0 ;
      RECT  147200.0 180800.0 147800.0 181399.99999999997 ;
      RECT  147500.0 181100.00000000003 158300.0 181700.0 ;
      RECT  147200.0 192700.0 147800.0 193300.0 ;
      RECT  147200.0 193000.0 147800.0 193600.00000000003 ;
      RECT  147500.0 192700.0 158300.0 193300.0 ;
      RECT  147200.0 199500.0 147800.0 200100.00000000003 ;
      RECT  147200.0 199200.0 147800.0 199800.0 ;
      RECT  147500.0 199500.0 158300.0 200100.00000000003 ;
      RECT  147200.0 211100.00000000003 147800.0 211700.0 ;
      RECT  147200.0 211400.00000000003 147800.0 212000.0 ;
      RECT  147500.0 211100.00000000003 158300.0 211700.0 ;
      RECT  147200.0 217900.00000000003 147800.0 218500.0 ;
      RECT  147200.0 217600.00000000003 147800.0 218200.0 ;
      RECT  147500.0 217900.00000000003 158300.0 218500.0 ;
      RECT  147200.0 229500.0 147800.0 230100.00000000003 ;
      RECT  147200.0 229800.0 147800.0 230399.99999999997 ;
      RECT  147500.0 229500.0 158300.0 230100.00000000003 ;
      RECT  147200.0 236300.0 147800.0 236899.99999999997 ;
      RECT  147200.0 236000.0 147800.0 236600.00000000003 ;
      RECT  147500.0 236300.0 158300.0 236899.99999999997 ;
      RECT  147200.0 247900.00000000003 147800.0 248500.0 ;
      RECT  147200.0 248200.0 147800.0 248800.0 ;
      RECT  147500.0 247900.00000000003 158300.0 248500.0 ;
      RECT  147200.0 254700.0 147800.0 255300.0 ;
      RECT  147200.0 254399.99999999997 147800.0 255000.0 ;
      RECT  147500.0 254700.0 158300.0 255300.0 ;
      RECT  147200.0 266300.0 147800.0 266900.0 ;
      RECT  147200.0 266600.0 147800.0 267200.0 ;
      RECT  147500.0 266300.0 158300.0 266900.0 ;
      RECT  157600.0 127300.00000000001 158200.0 127900.0 ;
      RECT  159200.0 127300.00000000001 159800.0 127900.0 ;
      RECT  157600.0 127600.00000000001 158200.0 129900.0 ;
      RECT  157899.99999999997 127300.00000000001 159500.0 127900.0 ;
      RECT  159200.0 124900.0 159800.0 127600.00000000001 ;
      RECT  157500.0 129900.0 158300.0 130699.99999999999 ;
      RECT  159100.0 124100.00000000001 159899.99999999997 124900.0 ;
      RECT  159899.99999999997 127200.0 159100.0 128000.0 ;
      RECT  157600.0 136700.0 158200.0 136100.00000000003 ;
      RECT  159200.0 136700.0 159800.0 136100.00000000003 ;
      RECT  157600.0 136400.0 158200.0 134100.00000000003 ;
      RECT  157899.99999999997 136700.0 159500.0 136100.00000000003 ;
      RECT  159200.0 139100.00000000003 159800.0 136400.0 ;
      RECT  157500.0 134100.00000000003 158300.0 133300.0 ;
      RECT  159100.0 139900.0 159899.99999999997 139100.00000000003 ;
      RECT  159899.99999999997 136800.0 159100.0 136000.0 ;
      RECT  157600.0 145700.0 158200.0 146300.0 ;
      RECT  159200.0 145700.0 159800.0 146300.0 ;
      RECT  157600.0 146000.0 158200.0 148300.0 ;
      RECT  157899.99999999997 145700.0 159500.0 146300.0 ;
      RECT  159200.0 143300.0 159800.0 146000.0 ;
      RECT  157500.0 148300.0 158300.0 149100.00000000003 ;
      RECT  159100.0 142500.0 159899.99999999997 143300.0 ;
      RECT  159899.99999999997 145600.00000000003 159100.0 146400.0 ;
      RECT  157600.0 155100.00000000003 158200.0 154500.0 ;
      RECT  159200.0 155100.00000000003 159800.0 154500.0 ;
      RECT  157600.0 154800.0 158200.0 152500.0 ;
      RECT  157899.99999999997 155100.00000000003 159500.0 154500.0 ;
      RECT  159200.0 157500.0 159800.0 154800.0 ;
      RECT  157500.0 152500.0 158300.0 151700.0 ;
      RECT  159100.0 158300.0 159899.99999999997 157500.0 ;
      RECT  159899.99999999997 155200.0 159100.0 154399.99999999997 ;
      RECT  157600.0 164100.00000000003 158200.0 164700.0 ;
      RECT  159200.0 164100.00000000003 159800.0 164700.0 ;
      RECT  157600.0 164399.99999999997 158200.0 166700.0 ;
      RECT  157899.99999999997 164100.00000000003 159500.0 164700.0 ;
      RECT  159200.0 161700.0 159800.0 164399.99999999997 ;
      RECT  157500.0 166700.0 158300.0 167500.0 ;
      RECT  159100.0 160899.99999999997 159899.99999999997 161700.0 ;
      RECT  159899.99999999997 164000.0 159100.0 164800.0 ;
      RECT  157600.0 173500.0 158200.0 172899.99999999997 ;
      RECT  159200.0 173500.0 159800.0 172899.99999999997 ;
      RECT  157600.0 173200.0 158200.0 170899.99999999997 ;
      RECT  157899.99999999997 173500.0 159500.0 172899.99999999997 ;
      RECT  159200.0 175899.99999999997 159800.0 173200.0 ;
      RECT  157500.0 170899.99999999997 158300.0 170100.00000000003 ;
      RECT  159100.0 176700.0 159899.99999999997 175899.99999999997 ;
      RECT  159899.99999999997 173600.00000000003 159100.0 172800.0 ;
      RECT  157600.0 182500.0 158200.0 183100.00000000003 ;
      RECT  159200.0 182500.0 159800.0 183100.00000000003 ;
      RECT  157600.0 182800.0 158200.0 185100.00000000003 ;
      RECT  157899.99999999997 182500.0 159500.0 183100.00000000003 ;
      RECT  159200.0 180100.00000000003 159800.0 182800.0 ;
      RECT  157500.0 185100.00000000003 158300.0 185899.99999999997 ;
      RECT  159100.0 179300.0 159899.99999999997 180100.00000000003 ;
      RECT  159899.99999999997 182399.99999999997 159100.0 183200.0 ;
      RECT  157600.0 191900.00000000003 158200.0 191300.0 ;
      RECT  159200.0 191900.00000000003 159800.0 191300.0 ;
      RECT  157600.0 191600.00000000003 158200.0 189300.0 ;
      RECT  157899.99999999997 191900.00000000003 159500.0 191300.0 ;
      RECT  159200.0 194300.0 159800.0 191600.00000000003 ;
      RECT  157500.0 189300.0 158300.0 188500.0 ;
      RECT  159100.0 195100.00000000003 159899.99999999997 194300.0 ;
      RECT  159899.99999999997 192000.0 159100.0 191200.0 ;
      RECT  157600.0 200900.00000000003 158200.0 201500.0 ;
      RECT  159200.0 200900.00000000003 159800.0 201500.0 ;
      RECT  157600.0 201200.0 158200.0 203500.0 ;
      RECT  157899.99999999997 200900.00000000003 159500.0 201500.0 ;
      RECT  159200.0 198500.0 159800.0 201200.0 ;
      RECT  157500.0 203500.0 158300.0 204300.0 ;
      RECT  159100.0 197700.0 159899.99999999997 198500.0 ;
      RECT  159899.99999999997 200800.0 159100.0 201600.00000000003 ;
      RECT  157600.0 210300.0 158200.0 209700.0 ;
      RECT  159200.0 210300.0 159800.0 209700.0 ;
      RECT  157600.0 210000.0 158200.0 207700.0 ;
      RECT  157899.99999999997 210300.0 159500.0 209700.0 ;
      RECT  159200.0 212700.0 159800.0 210000.0 ;
      RECT  157500.0 207700.0 158300.0 206899.99999999997 ;
      RECT  159100.0 213500.0 159899.99999999997 212700.0 ;
      RECT  159899.99999999997 210399.99999999997 159100.0 209600.00000000003 ;
      RECT  157600.0 219300.0 158200.0 219899.99999999997 ;
      RECT  159200.0 219300.0 159800.0 219899.99999999997 ;
      RECT  157600.0 219600.00000000003 158200.0 221899.99999999997 ;
      RECT  157899.99999999997 219300.0 159500.0 219899.99999999997 ;
      RECT  159200.0 216899.99999999997 159800.0 219600.00000000003 ;
      RECT  157500.0 221899.99999999997 158300.0 222700.0 ;
      RECT  159100.0 216100.00000000003 159899.99999999997 216899.99999999997 ;
      RECT  159899.99999999997 219200.0 159100.0 220000.0 ;
      RECT  157600.0 228700.0 158200.0 228100.00000000003 ;
      RECT  159200.0 228700.0 159800.0 228100.00000000003 ;
      RECT  157600.0 228400.00000000003 158200.0 226100.00000000003 ;
      RECT  157899.99999999997 228700.0 159500.0 228100.00000000003 ;
      RECT  159200.0 231100.00000000003 159800.0 228400.00000000003 ;
      RECT  157500.0 226100.00000000003 158300.0 225300.0 ;
      RECT  159100.0 231900.00000000003 159899.99999999997 231100.00000000003 ;
      RECT  159899.99999999997 228800.0 159100.0 228000.0 ;
      RECT  157600.0 237700.0 158200.0 238300.0 ;
      RECT  159200.0 237700.0 159800.0 238300.0 ;
      RECT  157600.0 238000.0 158200.0 240300.0 ;
      RECT  157899.99999999997 237700.0 159500.0 238300.0 ;
      RECT  159200.0 235300.0 159800.0 238000.0 ;
      RECT  157500.0 240300.0 158300.0 241100.00000000003 ;
      RECT  159100.0 234500.0 159899.99999999997 235300.0 ;
      RECT  159899.99999999997 237600.00000000003 159100.0 238400.00000000003 ;
      RECT  157600.0 247100.00000000003 158200.0 246500.0 ;
      RECT  159200.0 247100.00000000003 159800.0 246500.0 ;
      RECT  157600.0 246800.0 158200.0 244500.0 ;
      RECT  157899.99999999997 247100.00000000003 159500.0 246500.0 ;
      RECT  159200.0 249500.0 159800.0 246800.0 ;
      RECT  157500.0 244500.0 158300.0 243700.0 ;
      RECT  159100.0 250300.0 159899.99999999997 249500.0 ;
      RECT  159899.99999999997 247200.0 159100.0 246400.00000000003 ;
      RECT  157600.0 256100.00000000003 158200.0 256700.0 ;
      RECT  159200.0 256100.00000000003 159800.0 256700.0 ;
      RECT  157600.0 256400.00000000003 158200.0 258700.0 ;
      RECT  157899.99999999997 256100.00000000003 159500.0 256700.0 ;
      RECT  159200.0 253700.0 159800.0 256400.00000000003 ;
      RECT  157500.0 258700.0 158300.0 259500.0 ;
      RECT  159100.0 252900.00000000003 159899.99999999997 253700.0 ;
      RECT  159899.99999999997 256000.0 159100.0 256800.0 ;
      RECT  157600.0 265500.0 158200.0 264900.00000000006 ;
      RECT  159200.0 265500.0 159800.0 264900.00000000006 ;
      RECT  157600.0 265200.0 158200.0 262900.00000000006 ;
      RECT  157899.99999999997 265500.0 159500.0 264900.00000000006 ;
      RECT  159200.0 267900.00000000006 159800.0 265200.0 ;
      RECT  157500.0 262900.00000000006 158300.0 262100.00000000003 ;
      RECT  159100.0 268700.0 159899.99999999997 267900.00000000006 ;
      RECT  159899.99999999997 265600.0 159100.0 264800.0 ;
      RECT  145800.0 126800.00000000001 146600.0 127600.00000000001 ;
      RECT  147100.0 125200.0 147899.99999999997 126000.0 ;
      RECT  158300.0 125800.00000000001 157500.0 126600.00000000001 ;
      RECT  145800.0 136400.0 146600.0 137200.0 ;
      RECT  147100.0 138000.0 147899.99999999997 138800.0 ;
      RECT  158300.0 137400.0 157500.0 138200.0 ;
      RECT  145800.0 145200.0 146600.0 146000.0 ;
      RECT  147100.0 143600.00000000003 147899.99999999997 144400.0 ;
      RECT  158300.0 144200.0 157500.0 145000.0 ;
      RECT  145800.0 154800.0 146600.0 155600.00000000003 ;
      RECT  147100.0 156399.99999999997 147899.99999999997 157200.0 ;
      RECT  158300.0 155800.0 157500.0 156600.00000000003 ;
      RECT  145800.0 163600.00000000003 146600.0 164399.99999999997 ;
      RECT  147100.0 162000.0 147899.99999999997 162800.0 ;
      RECT  158300.0 162600.00000000003 157500.0 163399.99999999997 ;
      RECT  145800.0 173200.0 146600.0 174000.0 ;
      RECT  147100.0 174800.0 147899.99999999997 175600.00000000003 ;
      RECT  158300.0 174200.0 157500.0 175000.0 ;
      RECT  145800.0 182000.0 146600.0 182800.0 ;
      RECT  147100.0 180399.99999999997 147899.99999999997 181200.0 ;
      RECT  158300.0 181000.0 157500.0 181800.0 ;
      RECT  145800.0 191600.00000000003 146600.0 192399.99999999997 ;
      RECT  147100.0 193200.0 147899.99999999997 194000.0 ;
      RECT  158300.0 192600.00000000003 157500.0 193399.99999999997 ;
      RECT  145800.0 200400.00000000003 146600.0 201200.0 ;
      RECT  147100.0 198800.0 147899.99999999997 199600.00000000003 ;
      RECT  158300.0 199400.00000000003 157500.0 200200.0 ;
      RECT  145800.0 210000.0 146600.0 210800.0 ;
      RECT  147100.0 211600.00000000003 147899.99999999997 212400.00000000003 ;
      RECT  158300.0 211000.0 157500.0 211800.0 ;
      RECT  145800.0 218800.0 146600.0 219600.00000000003 ;
      RECT  147100.0 217200.0 147899.99999999997 218000.0 ;
      RECT  158300.0 217800.0 157500.0 218600.00000000003 ;
      RECT  145800.0 228400.00000000003 146600.0 229200.0 ;
      RECT  147100.0 230000.0 147899.99999999997 230800.0 ;
      RECT  158300.0 229400.00000000003 157500.0 230200.0 ;
      RECT  145800.0 237200.0 146600.0 238000.0 ;
      RECT  147100.0 235600.00000000003 147899.99999999997 236400.00000000003 ;
      RECT  158300.0 236200.0 157500.0 237000.0 ;
      RECT  145800.0 246800.0 146600.0 247600.00000000003 ;
      RECT  147100.0 248400.00000000003 147899.99999999997 249200.0 ;
      RECT  158300.0 247800.0 157500.0 248600.00000000003 ;
      RECT  145800.0 255600.00000000003 146600.0 256400.00000000003 ;
      RECT  147100.0 254000.0 147899.99999999997 254800.0 ;
      RECT  158300.0 254600.00000000003 157500.0 255400.00000000003 ;
      RECT  145800.0 265200.0 146600.0 266000.0 ;
      RECT  147100.0 266800.0 147899.99999999997 267600.0 ;
      RECT  158300.0 266200.0 157500.0 267000.0 ;
      RECT  155100.0 131600.00000000003 154300.0 132400.0 ;
      RECT  155100.0 131600.00000000003 154300.0 132400.0 ;
      RECT  164700.0 131600.00000000003 163899.99999999997 132400.0 ;
      RECT  164700.0 131600.00000000003 163899.99999999997 132400.0 ;
      RECT  155100.0 122400.0 154300.0 123200.0 ;
      RECT  155100.0 122400.0 154300.0 123200.0 ;
      RECT  164700.0 122400.0 163899.99999999997 123200.0 ;
      RECT  164700.0 122400.0 163899.99999999997 123200.0 ;
      RECT  155100.0 131600.00000000003 154300.0 132400.0 ;
      RECT  155100.0 131600.00000000003 154300.0 132400.0 ;
      RECT  164700.0 131600.00000000003 163899.99999999997 132400.0 ;
      RECT  164700.0 131600.00000000003 163899.99999999997 132400.0 ;
      RECT  155100.0 140800.0 154300.0 141600.00000000003 ;
      RECT  155100.0 140800.0 154300.0 141600.00000000003 ;
      RECT  164700.0 140800.0 163899.99999999997 141600.00000000003 ;
      RECT  164700.0 140800.0 163899.99999999997 141600.00000000003 ;
      RECT  155100.0 150000.0 154300.0 150800.0 ;
      RECT  155100.0 150000.0 154300.0 150800.0 ;
      RECT  164700.0 150000.0 163899.99999999997 150800.0 ;
      RECT  164700.0 150000.0 163899.99999999997 150800.0 ;
      RECT  155100.0 140800.0 154300.0 141600.00000000003 ;
      RECT  155100.0 140800.0 154300.0 141600.00000000003 ;
      RECT  164700.0 140800.0 163899.99999999997 141600.00000000003 ;
      RECT  164700.0 140800.0 163899.99999999997 141600.00000000003 ;
      RECT  155100.0 150000.0 154300.0 150800.0 ;
      RECT  155100.0 150000.0 154300.0 150800.0 ;
      RECT  164700.0 150000.0 163899.99999999997 150800.0 ;
      RECT  164700.0 150000.0 163899.99999999997 150800.0 ;
      RECT  155100.0 159200.0 154300.0 160000.0 ;
      RECT  155100.0 159200.0 154300.0 160000.0 ;
      RECT  164700.0 159200.0 163899.99999999997 160000.0 ;
      RECT  164700.0 159200.0 163899.99999999997 160000.0 ;
      RECT  155100.0 168399.99999999997 154300.0 169200.0 ;
      RECT  155100.0 168399.99999999997 154300.0 169200.0 ;
      RECT  164700.0 168399.99999999997 163899.99999999997 169200.0 ;
      RECT  164700.0 168399.99999999997 163899.99999999997 169200.0 ;
      RECT  155100.0 159200.0 154300.0 160000.0 ;
      RECT  155100.0 159200.0 154300.0 160000.0 ;
      RECT  164700.0 159200.0 163899.99999999997 160000.0 ;
      RECT  164700.0 159200.0 163899.99999999997 160000.0 ;
      RECT  155100.0 168399.99999999997 154300.0 169200.0 ;
      RECT  155100.0 168399.99999999997 154300.0 169200.0 ;
      RECT  164700.0 168399.99999999997 163899.99999999997 169200.0 ;
      RECT  164700.0 168399.99999999997 163899.99999999997 169200.0 ;
      RECT  155100.0 177600.00000000003 154300.0 178399.99999999997 ;
      RECT  155100.0 177600.00000000003 154300.0 178399.99999999997 ;
      RECT  164700.0 177600.00000000003 163899.99999999997 178399.99999999997 ;
      RECT  164700.0 177600.00000000003 163899.99999999997 178399.99999999997 ;
      RECT  155100.0 186800.0 154300.0 187600.00000000003 ;
      RECT  155100.0 186800.0 154300.0 187600.00000000003 ;
      RECT  164700.0 186800.0 163899.99999999997 187600.00000000003 ;
      RECT  164700.0 186800.0 163899.99999999997 187600.00000000003 ;
      RECT  155100.0 177600.00000000003 154300.0 178399.99999999997 ;
      RECT  155100.0 177600.00000000003 154300.0 178399.99999999997 ;
      RECT  164700.0 177600.00000000003 163899.99999999997 178399.99999999997 ;
      RECT  164700.0 177600.00000000003 163899.99999999997 178399.99999999997 ;
      RECT  155100.0 186800.0 154300.0 187600.00000000003 ;
      RECT  155100.0 186800.0 154300.0 187600.00000000003 ;
      RECT  164700.0 186800.0 163899.99999999997 187600.00000000003 ;
      RECT  164700.0 186800.0 163899.99999999997 187600.00000000003 ;
      RECT  155100.0 196000.0 154300.0 196800.0 ;
      RECT  155100.0 196000.0 154300.0 196800.0 ;
      RECT  164700.0 196000.0 163899.99999999997 196800.0 ;
      RECT  164700.0 196000.0 163899.99999999997 196800.0 ;
      RECT  155100.0 205200.0 154300.0 206000.0 ;
      RECT  155100.0 205200.0 154300.0 206000.0 ;
      RECT  164700.0 205200.0 163899.99999999997 206000.0 ;
      RECT  164700.0 205200.0 163899.99999999997 206000.0 ;
      RECT  155100.0 196000.0 154300.0 196800.0 ;
      RECT  155100.0 196000.0 154300.0 196800.0 ;
      RECT  164700.0 196000.0 163899.99999999997 196800.0 ;
      RECT  164700.0 196000.0 163899.99999999997 196800.0 ;
      RECT  155100.0 205200.0 154300.0 206000.0 ;
      RECT  155100.0 205200.0 154300.0 206000.0 ;
      RECT  164700.0 205200.0 163899.99999999997 206000.0 ;
      RECT  164700.0 205200.0 163899.99999999997 206000.0 ;
      RECT  155100.0 214400.00000000003 154300.0 215200.0 ;
      RECT  155100.0 214400.00000000003 154300.0 215200.0 ;
      RECT  164700.0 214400.00000000003 163899.99999999997 215200.0 ;
      RECT  164700.0 214400.00000000003 163899.99999999997 215200.0 ;
      RECT  155100.0 223600.00000000003 154300.0 224400.00000000003 ;
      RECT  155100.0 223600.00000000003 154300.0 224400.00000000003 ;
      RECT  164700.0 223600.00000000003 163899.99999999997 224400.00000000003 ;
      RECT  164700.0 223600.00000000003 163899.99999999997 224400.00000000003 ;
      RECT  155100.0 214400.00000000003 154300.0 215200.0 ;
      RECT  155100.0 214400.00000000003 154300.0 215200.0 ;
      RECT  164700.0 214400.00000000003 163899.99999999997 215200.0 ;
      RECT  164700.0 214400.00000000003 163899.99999999997 215200.0 ;
      RECT  155100.0 223600.00000000003 154300.0 224400.00000000003 ;
      RECT  155100.0 223600.00000000003 154300.0 224400.00000000003 ;
      RECT  164700.0 223600.00000000003 163899.99999999997 224400.00000000003 ;
      RECT  164700.0 223600.00000000003 163899.99999999997 224400.00000000003 ;
      RECT  155100.0 232800.0 154300.0 233600.00000000003 ;
      RECT  155100.0 232800.0 154300.0 233600.00000000003 ;
      RECT  164700.0 232800.0 163899.99999999997 233600.00000000003 ;
      RECT  164700.0 232800.0 163899.99999999997 233600.00000000003 ;
      RECT  155100.0 242000.0 154300.0 242800.0 ;
      RECT  155100.0 242000.0 154300.0 242800.0 ;
      RECT  164700.0 242000.0 163899.99999999997 242800.0 ;
      RECT  164700.0 242000.0 163899.99999999997 242800.0 ;
      RECT  155100.0 232800.0 154300.0 233600.00000000003 ;
      RECT  155100.0 232800.0 154300.0 233600.00000000003 ;
      RECT  164700.0 232800.0 163899.99999999997 233600.00000000003 ;
      RECT  164700.0 232800.0 163899.99999999997 233600.00000000003 ;
      RECT  155100.0 242000.0 154300.0 242800.0 ;
      RECT  155100.0 242000.0 154300.0 242800.0 ;
      RECT  164700.0 242000.0 163899.99999999997 242800.0 ;
      RECT  164700.0 242000.0 163899.99999999997 242800.0 ;
      RECT  155100.0 251200.0 154300.0 252000.0 ;
      RECT  155100.0 251200.0 154300.0 252000.0 ;
      RECT  164700.0 251200.0 163899.99999999997 252000.0 ;
      RECT  164700.0 251200.0 163899.99999999997 252000.0 ;
      RECT  155100.0 260399.99999999997 154300.0 261200.0 ;
      RECT  155100.0 260399.99999999997 154300.0 261200.0 ;
      RECT  164700.0 260399.99999999997 163899.99999999997 261200.0 ;
      RECT  164700.0 260399.99999999997 163899.99999999997 261200.0 ;
      RECT  155100.0 251200.0 154300.0 252000.0 ;
      RECT  155100.0 251200.0 154300.0 252000.0 ;
      RECT  164700.0 251200.0 163899.99999999997 252000.0 ;
      RECT  164700.0 251200.0 163899.99999999997 252000.0 ;
      RECT  155100.0 260399.99999999997 154300.0 261200.0 ;
      RECT  155100.0 260399.99999999997 154300.0 261200.0 ;
      RECT  164700.0 260399.99999999997 163899.99999999997 261200.0 ;
      RECT  164700.0 260399.99999999997 163899.99999999997 261200.0 ;
      RECT  155100.0 269600.0 154300.0 270400.00000000006 ;
      RECT  155100.0 269600.0 154300.0 270400.00000000006 ;
      RECT  164700.0 269600.0 163899.99999999997 270400.00000000006 ;
      RECT  164700.0 269600.0 163899.99999999997 270400.00000000006 ;
      RECT  145899.99999999997 122800.00000000001 146500.0 270000.0 ;
      RECT  174500.0 108700.0 173700.00000000003 109500.0 ;
      RECT  175900.0 28900.000000000007 175100.00000000003 29700.000000000007 ;
      RECT  177300.0 98500.0 176500.0 99300.0 ;
      RECT  146600.00000000003 271000.0 145800.0 271800.0 ;
      RECT  173100.00000000003 271000.0 172300.0 271800.0 ;
      RECT  179200.0 68800.00000000001 180000.0 71800.00000000001 ;
      RECT  186000.0 68800.00000000001 186800.0 71800.00000000001 ;
      RECT  181600.00000000003 24200.000000000004 182400.0 26200.000000000004 ;
      RECT  188400.0 24200.000000000004 189200.0 26200.000000000004 ;
      RECT  73900.0 122800.00000000001 74500.0 196399.99999999997 ;
      RECT  75300.0 122800.00000000001 75900.0 196399.99999999997 ;
      RECT  76700.0 122800.00000000001 77300.0 196399.99999999997 ;
      RECT  78100.00000000001 122800.00000000001 78700.0 196399.99999999997 ;
      RECT  176600.00000000003 24200.000000000004 177200.0 273200.0 ;
      RECT  175200.0 24200.000000000004 175800.0 273200.0 ;
      RECT  173800.0 24200.000000000004 174400.0 273200.0 ;
      RECT  172400.0 24200.000000000004 173000.0 273200.0 ;
      RECT  28200.000000000004 19600.0 28800.000000000004 98200.00000000001 ;
      RECT  29600.0 19600.0 30200.000000000004 98200.00000000001 ;
      RECT  31000.0 19600.0 31600.0 98200.00000000001 ;
      RECT  32400.0 19600.0 33000.0 98200.00000000001 ;
      RECT  32400.0 29200.000000000004 33000.0 58900.00000000001 ;
      RECT  31000.0 50000.0 31600.0 58900.00000000001 ;
      RECT  2800.0000000000005 59600.0 3400.0000000000005 62400.0 ;
      RECT  29600.0 58900.00000000001 30200.000000000004 65300.000000000015 ;
      RECT  32400.0 58900.00000000001 33000.0 64000.0 ;
      RECT  31000.0 58900.00000000001 31600.0 62700.0 ;
      RECT  29600.0 58900.00000000001 30200.000000000004 94800.00000000001 ;
      RECT  32400.0 58900.00000000001 33000.0 96200.00000000001 ;
      RECT  1600.0 89800.00000000001 2200.0 129100.0 ;
      RECT  8900.0 108800.00000000001 9500.0 124500.0 ;
      RECT  28200.000000000004 50400.00000000001 28800.000000000004 58900.0 ;
      RECT  29600.0 28800.000000000004 30200.000000000004 58900.00000000001 ;
      RECT  0.0 19600.0 21800.0 39600.0 ;
      RECT  18800.0 29000.0 19600.0 29800.000000000004 ;
      RECT  23400.000000000004 28800.000000000004 24200.000000000004 29600.0 ;
      RECT  23400.000000000004 28800.000000000004 24200.000000000004 29600.0 ;
      RECT  25000.0 28800.000000000004 25800.0 29600.0 ;
      RECT  7600.000000000001 28200.000000000004 8400.0 29000.0 ;
      RECT  18900.000000000004 29100.0 19500.0 29700.000000000004 ;
      RECT  25100.0 28900.000000000004 25700.000000000004 29500.0 ;
      RECT  2800.0000000000005 26200.000000000004 3600.0 27000.0 ;
      RECT  0.0 59600.0 21800.0 39600.0 ;
      RECT  18800.0 50200.0 19600.0 49400.0 ;
      RECT  23400.000000000004 50400.0 24200.000000000004 49600.0 ;
      RECT  23400.000000000004 50400.0 24200.000000000004 49600.0 ;
      RECT  25000.0 50400.0 25800.0 49600.0 ;
      RECT  7600.000000000001 51000.0 8400.0 50200.0 ;
      RECT  18900.000000000004 50100.0 19500.0 49500.0 ;
      RECT  25100.0 50300.0 25700.000000000004 49700.0 ;
      RECT  2800.0000000000005 53000.0 3600.0 52200.0 ;
      RECT  400.0 39200.0 -400.0 40000.0 ;
      RECT  400.0 39200.0 -400.0 40000.0 ;
      RECT  400.0 19200.000000000004 -400.0 20000.0 ;
      RECT  400.0 19200.000000000004 -400.0 20000.0 ;
      RECT  400.0 39200.0 -400.0 40000.0 ;
      RECT  400.0 39200.0 -400.0 40000.0 ;
      RECT  400.0 59200.0 -400.0 60000.0 ;
      RECT  400.0 59200.0 -400.0 60000.0 ;
      RECT  7600.000000000001 28200.000000000004 8400.0 29000.0 ;
      RECT  7600.000000000001 50200.0 8400.0 51000.0 ;
      RECT  18900.000000000004 29100.0 19500.0 29700.000000000004 ;
      RECT  25100.0 28900.000000000004 25700.000000000004 29500.0 ;
      RECT  18900.000000000004 49500.0 19500.0 50100.0 ;
      RECT  25100.0 49700.0 25700.000000000004 50300.00000000001 ;
      RECT  2800.0000000000005 19600.0 3400.0000000000005 59600.0 ;
      RECT  38500.0 29400.000000000004 39100.0 50400.00000000001 ;
      RECT  39200.0 50000.0 38400.00000000001 50800.00000000001 ;
      RECT  38400.00000000001 29000.0 39200.0 29800.000000000004 ;
      RECT  51200.0 50000.0 52000.0 50800.00000000001 ;
      RECT  51200.0 28400.000000000004 52000.0 29200.000000000004 ;
      RECT  36800.00000000001 29000.0 37600.0 29800.000000000004 ;
      RECT  36900.00000000001 29100.0 37500.0 29700.000000000004 ;
      RECT  51300.00000000001 28500.0 51900.00000000001 29100.0 ;
      RECT  51300.00000000001 50100.0 51900.00000000001 50700.0 ;
      RECT  41300.00000000001 61700.0 41900.00000000001 77500.0 ;
      RECT  38100.0 65000.0 38700.0 65600.0 ;
      RECT  41300.00000000001 65000.0 41900.00000000001 65600.0 ;
      RECT  38100.0 65300.000000000015 38700.0 77500.0 ;
      RECT  38400.00000000001 65000.0 41600.0 65600.0 ;
      RECT  41300.00000000001 61700.0 41900.00000000001 65300.000000000015 ;
      RECT  38000.0 77500.0 38800.00000000001 78300.00000000001 ;
      RECT  41200.0 77500.0 42000.0 78300.00000000001 ;
      RECT  41200.0 60900.0 42000.0 61700.0 ;
      RECT  41200.0 64900.00000000001 42000.0 65700.0 ;
      RECT  38100.0 95100.0 38700.0 94500.0 ;
      RECT  39700.0 95100.0 40300.00000000001 94500.0 ;
      RECT  38100.0 94800.00000000001 38700.0 81699.99999999999 ;
      RECT  38400.00000000001 95100.0 40000.0 94500.0 ;
      RECT  39700.0 97500.0 40300.00000000001 94800.00000000001 ;
      RECT  38000.0 81699.99999999999 38800.00000000001 80900.0 ;
      RECT  39600.0 98300.00000000001 40400.00000000001 97500.0 ;
      RECT  40400.00000000001 95199.99999999999 39600.0 94400.0 ;
      RECT  22700.000000000004 131400.0 23300.000000000004 132000.0 ;
      RECT  22700.000000000004 131700.00000000003 23300.000000000004 133700.00000000003 ;
      RECT  16800.0 131400.0 23000.0 132000.0 ;
      RECT  15700.000000000002 122400.0 16300.0 123000.0 ;
      RECT  29700.000000000004 122400.0 30300.000000000004 123000.0 ;
      RECT  15700.000000000002 122700.00000000001 16300.0 129500.0 ;
      RECT  16000.0 122400.0 30000.0 123000.0 ;
      RECT  29700.000000000004 122700.00000000001 30300.000000000004 124100.00000000003 ;
      RECT  3300.0000000000005 142600.00000000003 3900.0000000000005 143200.00000000003 ;
      RECT  1700.0000000000002 142600.00000000003 2300.0000000000005 143200.00000000003 ;
      RECT  3300.0000000000005 138100.00000000003 3900.0000000000005 142900.0 ;
      RECT  2000.0 142600.00000000003 3600.0 143200.00000000003 ;
      RECT  1700.0000000000002 142900.0 2300.0000000000005 147700.00000000003 ;
      RECT  3300.0000000000005 151800.0 3900.0000000000005 152400.0 ;
      RECT  1700.0000000000002 151800.0 2300.0000000000005 152400.0 ;
      RECT  3300.0000000000005 147700.00000000003 3900.0000000000005 152100.0 ;
      RECT  2000.0 151800.0 3600.0 152400.0 ;
      RECT  1700.0000000000002 152100.0 2300.0000000000005 156500.00000000003 ;
      RECT  3300.0000000000005 161000.0 3900.0000000000005 161600.0 ;
      RECT  1700.0000000000002 161000.0 2300.0000000000005 161600.0 ;
      RECT  3300.0000000000005 156500.0 3900.0000000000005 161300.0 ;
      RECT  2000.0 161000.0 3600.0 161600.0 ;
      RECT  1700.0000000000002 161300.0 2300.0000000000005 166100.0 ;
      RECT  22700.000000000004 165800.0 23300.000000000004 166400.0 ;
      RECT  21200.000000000004 165800.0 23000.000000000004 166400.0 ;
      RECT  22700.000000000004 133700.00000000003 23300.000000000004 166100.0 ;
      RECT  8000.0 137700.00000000003 8800.0 138500.0 ;
      RECT  8000.0 137700.00000000003 8800.0 138500.0 ;
      RECT  14400.0 137700.00000000003 15200.000000000002 138500.0 ;
      RECT  14400.0 137700.00000000003 15200.000000000002 138500.0 ;
      RECT  20800.0 137700.00000000003 21600.0 138500.0 ;
      RECT  20800.0 137700.00000000003 21600.0 138500.0 ;
      RECT  1600.0 137700.00000000003 2400.0000000000005 138500.0 ;
      RECT  3200.0 137700.00000000003 4000.0 138500.0 ;
      RECT  3200.0 137700.00000000003 4000.0 138500.0 ;
      RECT  8000.0 147300.0 8800.0 148100.0 ;
      RECT  8000.0 147300.0 8800.0 148100.0 ;
      RECT  14400.0 147300.0 15200.000000000002 148100.0 ;
      RECT  14400.0 147300.0 15200.000000000002 148100.0 ;
      RECT  20800.0 147300.0 21600.0 148100.0 ;
      RECT  20800.0 147300.0 21600.0 148100.0 ;
      RECT  1600.0 147300.0 2400.0000000000005 148100.0 ;
      RECT  3200.0 147300.0 4000.0 148100.0 ;
      RECT  3200.0 147300.0 4000.0 148100.0 ;
      RECT  8000.0 156100.0 8800.0 156900.0 ;
      RECT  8000.0 156100.0 8800.0 156900.0 ;
      RECT  14400.0 156100.0 15200.000000000002 156900.0 ;
      RECT  14400.0 156100.0 15200.000000000002 156900.0 ;
      RECT  20800.0 156100.0 21600.0 156900.0 ;
      RECT  20800.0 156100.0 21600.0 156900.0 ;
      RECT  1600.0 156100.0 2400.0000000000005 156900.0 ;
      RECT  3200.0 156100.0 4000.0 156900.0 ;
      RECT  3200.0 156100.0 4000.0 156900.0 ;
      RECT  8000.0 165700.00000000003 8800.0 166500.0 ;
      RECT  8000.0 165700.00000000003 8800.0 166500.0 ;
      RECT  14400.0 165700.00000000003 15200.000000000002 166500.0 ;
      RECT  14400.0 165700.00000000003 15200.000000000002 166500.0 ;
      RECT  20800.0 165700.00000000003 21600.0 166500.0 ;
      RECT  20800.0 165700.00000000003 21600.0 166500.0 ;
      RECT  1600.0 165700.00000000003 2400.0000000000005 166500.0 ;
      RECT  3200.0 165700.00000000003 4000.0 166500.0 ;
      RECT  3200.0 165700.00000000003 4000.0 166500.0 ;
      RECT  13200.000000000002 142500.0 12400.0 143300.0 ;
      RECT  13200.000000000002 142500.0 12400.0 143300.0 ;
      RECT  13200.000000000002 133300.0 12400.0 134100.00000000003 ;
      RECT  13200.000000000002 133300.0 12400.0 134100.00000000003 ;
      RECT  19600.0 142500.0 18800.0 143300.0 ;
      RECT  19600.0 142500.0 18800.0 143300.0 ;
      RECT  19600.0 133300.0 18800.0 134100.00000000003 ;
      RECT  19600.0 133300.0 18800.0 134100.00000000003 ;
      RECT  13200.000000000002 160900.0 12400.0 161700.00000000003 ;
      RECT  13200.000000000002 160900.0 12400.0 161700.00000000003 ;
      RECT  13200.000000000002 151700.00000000003 12400.0 152500.0 ;
      RECT  13200.000000000002 151700.00000000003 12400.0 152500.0 ;
      RECT  19600.0 160900.0 18800.0 161700.00000000003 ;
      RECT  19600.0 160900.0 18800.0 161700.00000000003 ;
      RECT  19600.0 151700.00000000003 18800.0 152500.0 ;
      RECT  19600.0 151700.00000000003 18800.0 152500.0 ;
      RECT  13200.000000000002 170100.0 12400.0 170900.0 ;
      RECT  13200.000000000002 170100.0 12400.0 170900.0 ;
      RECT  19600.0 170100.0 18800.0 170900.0 ;
      RECT  19600.0 170100.0 18800.0 170900.0 ;
      RECT  1600.0 137700.00000000003 2400.0000000000005 138500.0 ;
      RECT  20800.0 165700.00000000003 21600.0 166500.0 ;
      RECT  1600.0 133700.00000000003 2200.0 138100.00000000003 ;
      RECT  22700.000000000004 133700.00000000003 23300.0 166100.0 ;
      RECT  28400.000000000004 133700.00000000003 35200.0 124500.0 ;
      RECT  28400.000000000004 133700.00000000003 35200.0 142900.0 ;
      RECT  28400.000000000004 152100.0 35200.0 142900.0 ;
      RECT  28400.000000000004 152100.0 35200.0 161300.0 ;
      RECT  28400.000000000004 170500.00000000003 35200.0 161300.0 ;
      RECT  28400.000000000004 170500.00000000003 35200.0 179700.00000000003 ;
      RECT  28400.000000000004 188900.0 35200.0 179700.00000000003 ;
      RECT  28400.000000000004 188900.0 35200.0 198100.0 ;
      RECT  28400.000000000004 207300.0 35200.0 198100.0 ;
      RECT  31400.000000000004 142500.0 32200.000000000004 143300.0 ;
      RECT  31400.000000000004 142500.0 32200.000000000004 143300.0 ;
      RECT  31400.000000000004 160900.0 32200.000000000004 161700.00000000003 ;
      RECT  31400.000000000004 160900.0 32200.000000000004 161700.00000000003 ;
      RECT  31400.000000000004 179300.0 32200.000000000004 180100.0 ;
      RECT  31400.000000000004 179300.0 32200.000000000004 180100.0 ;
      RECT  31400.000000000004 197700.00000000003 32200.000000000004 198500.0 ;
      RECT  31400.000000000004 197700.00000000003 32200.000000000004 198500.0 ;
      RECT  28000.000000000004 137900.0 28800.0 138700.00000000003 ;
      RECT  34800.00000000001 137900.0 35600.0 138700.00000000003 ;
      RECT  28000.000000000004 147100.00000000003 28800.0 147900.0 ;
      RECT  34800.00000000001 147100.00000000003 35600.0 147900.0 ;
      RECT  28000.000000000004 156300.0 28800.0 157100.0 ;
      RECT  34800.00000000001 156300.0 35600.0 157100.0 ;
      RECT  28000.000000000004 165500.0 28800.0 166300.0 ;
      RECT  34800.00000000001 165500.0 35600.0 166300.0 ;
      RECT  28000.000000000004 174700.00000000003 28800.0 175500.0 ;
      RECT  34800.00000000001 174700.00000000003 35600.0 175500.0 ;
      RECT  28000.000000000004 183900.0 28800.0 184700.00000000003 ;
      RECT  34800.00000000001 183900.0 35600.0 184700.00000000003 ;
      RECT  28000.000000000004 193100.0 28800.0 193900.0 ;
      RECT  34800.00000000001 193100.0 35600.0 193900.0 ;
      RECT  28000.000000000004 202300.0 28800.0 203100.0 ;
      RECT  34800.00000000001 202300.0 35600.0 203100.0 ;
      RECT  29600.0 133300.0 30400.000000000004 208700.00000000003 ;
      RECT  33200.0 134100.00000000003 34000.0 209500.0 ;
      RECT  6800.000000000001 124100.00000000003 6000.000000000001 124900.0 ;
      RECT  6800.000000000001 124100.00000000003 6000.000000000001 124900.0 ;
      RECT  31400.000000000004 122700.00000000001 32200.000000000004 123500.0 ;
      RECT  31400.000000000004 122700.00000000001 32200.000000000004 123500.0 ;
      RECT  28800.0 128700.00000000001 28000.0 129500.0 ;
      RECT  28800.0 128700.00000000001 28000.0 129500.0 ;
      RECT  35600.0 128700.00000000001 34800.00000000001 129500.0 ;
      RECT  35600.0 128700.00000000001 34800.00000000001 129500.0 ;
      RECT  37200.0 134700.00000000003 36400.00000000001 135500.0 ;
      RECT  37200.0 134700.00000000003 36400.00000000001 135500.0 ;
      RECT  37200.0 150300.0 36400.00000000001 151100.0 ;
      RECT  37200.0 150300.0 36400.00000000001 151100.0 ;
      RECT  37200.0 153100.0 36400.00000000001 153900.0 ;
      RECT  37200.0 153100.0 36400.00000000001 153900.0 ;
      RECT  37200.0 168700.00000000003 36400.00000000001 169500.0 ;
      RECT  37200.0 168700.00000000003 36400.00000000001 169500.0 ;
      RECT  37200.0 171500.0 36400.00000000001 172300.0 ;
      RECT  37200.0 171500.0 36400.00000000001 172300.0 ;
      RECT  37200.0 187100.0 36400.00000000001 187900.0 ;
      RECT  37200.0 187100.0 36400.00000000001 187900.0 ;
      RECT  37200.0 189900.0 36400.00000000001 190700.00000000003 ;
      RECT  37200.0 189900.0 36400.00000000001 190700.00000000003 ;
      RECT  37200.0 205500.0 36400.00000000001 206299.99999999997 ;
      RECT  37200.0 205500.0 36400.00000000001 206299.99999999997 ;
      RECT  16400.000000000004 131300.0 17200.000000000004 132100.00000000003 ;
      RECT  17200.000000000004 129100.00000000003 18000.000000000004 129900.0 ;
      RECT  17200.000000000004 129100.00000000003 18000.000000000004 129900.0 ;
      RECT  15600.000000000002 129100.00000000003 16400.000000000004 129900.0 ;
      RECT  8800.0 128900.0 9600.000000000002 129700.00000000001 ;
      RECT  1600.0000000000014 124500.0 2199.999999999999 133700.00000000003 ;
      RECT  8900.000000000002 124500.0 9500.0 129300.00000000001 ;
      RECT  33100.0 28800.000000000004 32300.000000000004 29600.0 ;
      RECT  25000.0 28800.000000000004 25800.0 29600.0 ;
      RECT  31700.000000000004 49600.0 30900.000000000004 50400.00000000001 ;
      RECT  25000.0 49600.0 25800.0 50400.00000000001 ;
      RECT  3500.0 62000.00000000001 2700.0 62800.00000000001 ;
      RECT  28900.000000000004 62000.00000000001 28100.0 62800.00000000001 ;
      RECT  30300.0 64900.00000000001 29500.0 65700.0 ;
      RECT  33100.0 63600.0 32300.000000000004 64400.00000000001 ;
      RECT  31700.000000000004 62300.00000000001 30900.000000000004 63100.0 ;
      RECT  30300.0 94400.0 29500.0 95199.99999999999 ;
      RECT  33100.0 95800.00000000001 32300.000000000004 96600.0 ;
      RECT  2300.0000000000005 89400.0 1500.0000000000002 90199.99999999999 ;
      RECT  48800.00000000001 89400.0 48000.00000000001 90199.99999999999 ;
      RECT  48800.00000000001 89400.0 48000.00000000001 90199.99999999999 ;
      RECT  9600.000000000002 108400.0 8800.0 109200.00000000001 ;
      RECT  28900.000000000004 50000.0 28100.0 50800.00000000001 ;
      RECT  51200.0 50000.0 52000.0 50800.00000000001 ;
      RECT  30300.0 28400.000000000004 29500.0 29200.000000000004 ;
      RECT  51200.0 28400.000000000004 52000.0 29200.000000000004 ;
      RECT  70000.0 39200.0 69200.0 40000.0 ;
      RECT  70000.0 39200.0 69200.0 40000.0 ;
      RECT  70000.0 59200.0 69200.0 60000.0 ;
      RECT  70000.0 59200.0 69200.0 60000.0 ;
      RECT  70000.0 19200.000000000004 69200.0 20000.0 ;
      RECT  70000.0 19200.000000000004 69200.0 20000.0 ;
      RECT  70000.0 79200.0 69200.0 80000.0 ;
      RECT  70000.0 79200.0 69200.0 80000.0 ;
      RECT  70000.0 59200.0 69200.0 60000.0 ;
      RECT  70000.0 59200.0 69200.0 60000.0 ;
      RECT  70000.0 79200.0 69200.0 80000.0 ;
      RECT  70000.0 79200.0 69200.0 80000.0 ;
      RECT  70000.0 99200.00000000001 69200.0 100000.0 ;
      RECT  70000.0 99200.00000000001 69200.0 100000.0 ;
      RECT  70000.0 119200.00000000001 69200.0 120000.0 ;
      RECT  70000.0 119200.00000000001 69200.0 120000.0 ;
      RECT  70000.0 99200.00000000001 69200.0 100000.0 ;
      RECT  70000.0 99200.00000000001 69200.0 100000.0 ;
      RECT  7600.000000000001 28200.000000000004 8400.0 29000.0 ;
      RECT  7600.000000000001 50200.0 8400.0 51000.0 ;
      RECT  36900.0 19600.0 37500.0 29100.0 ;
      RECT  51999.99999999999 211900.00000000003 52599.99999999999 291900.00000000006 ;
      RECT  49199.99999999999 211900.00000000003 71000.0 231900.00000000003 ;
      RECT  49199.99999999999 251900.00000000003 71000.0 231900.00000000003 ;
      RECT  49199.99999999999 251900.00000000003 71000.0 271900.00000000006 ;
      RECT  49199.99999999999 291900.00000000006 71000.0 271900.00000000006 ;
      RECT  60500.0 231500.00000000003 59699.99999999999 232300.00000000003 ;
      RECT  60500.0 231500.00000000003 59699.99999999999 232300.00000000003 ;
      RECT  60500.0 211500.00000000003 59699.99999999999 212300.00000000003 ;
      RECT  60500.0 211500.00000000003 59699.99999999999 212300.00000000003 ;
      RECT  60500.0 231500.00000000003 59699.99999999999 232300.00000000003 ;
      RECT  60500.0 231500.00000000003 59699.99999999999 232300.00000000003 ;
      RECT  60500.0 251500.00000000003 59699.99999999999 252300.00000000003 ;
      RECT  60500.0 251500.00000000003 59699.99999999999 252300.00000000003 ;
      RECT  60500.0 271500.00000000006 59699.99999999999 272300.0 ;
      RECT  60500.0 271500.00000000006 59699.99999999999 272300.0 ;
      RECT  60500.0 251500.00000000003 59699.99999999999 252300.00000000003 ;
      RECT  60500.0 251500.00000000003 59699.99999999999 252300.00000000003 ;
      RECT  60500.0 271500.00000000006 59699.99999999999 272300.0 ;
      RECT  60500.0 271500.00000000006 59699.99999999999 272300.0 ;
      RECT  60500.0 291500.00000000006 59699.99999999999 292300.00000000006 ;
      RECT  60500.0 291500.00000000006 59699.99999999999 292300.00000000006 ;
      RECT  51999.99999999999 214900.00000000003 52800.0 215700.00000000006 ;
      RECT  56800.0 220500.00000000003 57599.99999999999 221300.00000000003 ;
      RECT  56800.0 242500.00000000003 57599.99999999999 243300.00000000003 ;
      RECT  56800.0 260500.00000000006 57599.99999999999 261300.00000000006 ;
      RECT  56800.0 282500.00000000006 57599.99999999999 283300.00000000006 ;
      RECT  68000.0 221300.00000000003 68800.0 222100.00000000003 ;
      RECT  68000.0 241700.00000000006 68800.0 242500.00000000003 ;
      RECT  68000.0 261300.00000000006 68800.0 262100.00000000003 ;
      RECT  68000.0 281700.00000000006 68800.0 282500.00000000006 ;
      RECT  181400.00000000003 0.0 182000.00000000003 20000.0 ;
      RECT  203200.00000000003 0.0 203800.0 20000.0 ;
      RECT  178600.00000000003 0.0 200400.00000000003 20000.0 ;
      RECT  200400.00000000003 0.0 222200.00000000003 20000.0 ;
      RECT  189900.00000000003 19600.0 189100.00000000003 20400.000000000004 ;
      RECT  189900.00000000003 19600.0 189100.00000000003 20400.000000000004 ;
      RECT  189900.00000000003 -400.0 189100.00000000003 400.0 ;
      RECT  189900.00000000003 -400.0 189100.00000000003 400.0 ;
      RECT  211700.00000000003 19600.0 210900.00000000003 20400.000000000004 ;
      RECT  211700.00000000003 19600.0 210900.00000000003 20400.000000000004 ;
      RECT  211700.00000000003 -400.0 210900.00000000003 400.0 ;
      RECT  211700.00000000003 -400.0 210900.00000000003 400.0 ;
      RECT  181400.00000000003 3000.0 182200.00000000003 3800.0 ;
      RECT  203200.00000000003 3000.0 204000.00000000003 3800.0 ;
      RECT  186200.00000000003 8600.0 187000.00000000003 9400.0 ;
      RECT  208000.00000000003 8600.0 208800.0 9400.0 ;
      RECT  197400.00000000003 9400.0 198200.00000000003 10200.000000000002 ;
      RECT  219200.00000000003 9400.0 220000.00000000003 10200.000000000002 ;
      RECT  173100.00000000003 3000.0 172300.0 3800.0 ;
      RECT  72800.0 214900.00000000003 72000.0 215700.00000000006 ;
      RECT  72800.0 50000.0 72000.0 50800.0 ;
      RECT  177300.0 108400.0 176500.0 109200.0 ;
      RECT  71399.99999999999 108400.0 70600.0 109200.0 ;
      RECT  71399.99999999999 108400.0 70600.0 109200.0 ;
      RECT  175900.0 68400.0 175100.0 69200.0 ;
      RECT  71399.99999999999 68400.0 70600.0 69200.0 ;
      RECT  71399.99999999999 68400.0 70600.0 69200.0 ;
      RECT  174500.0 28400.000000000004 173700.0 29200.000000000004 ;
      RECT  71399.99999999999 28400.000000000004 70600.0 29200.000000000004 ;
      RECT  71399.99999999999 28400.000000000004 70600.0 29200.000000000004 ;
      RECT  173100.00000000003 50000.0 172300.0 50800.0 ;
      RECT  71399.99999999999 50000.0 70600.0 50800.0 ;
      RECT  71399.99999999999 50000.0 70600.0 50800.0 ;
      RECT  74600.0 221300.0 73800.0 222100.00000000003 ;
      RECT  68800.0 221300.0 68000.0 222100.00000000003 ;
      RECT  76000.0 241700.0 75200.0 242500.0 ;
      RECT  68800.0 241700.0 68000.0 242500.0 ;
      RECT  77399.99999999999 261300.0 76600.0 262100.00000000003 ;
      RECT  68800.0 261300.0 68000.0 262100.00000000003 ;
      RECT  78800.0 281700.0 78000.0 282500.0 ;
      RECT  68800.0 281700.0 68000.0 282500.0 ;
      RECT  182400.0 22400.000000000004 181600.0 23200.000000000004 ;
      RECT  198200.0 22400.000000000004 197399.99999999997 23200.000000000004 ;
      RECT  189200.0 23800.000000000004 188399.99999999997 24600.000000000004 ;
      RECT  220000.0 23800.000000000004 219200.0 24600.000000000004 ;
   LAYER  metal3 ;
      RECT  172700.0 3100.0000000000014 200399.99999999997 3700.0000000000014 ;
      RECT  71000.0 215000.0 72400.0 215600.0 ;
      RECT  71000.0 50100.00000000001 72400.0 50700.00000000001 ;
      RECT  71000.0 108500.00000000001 176900.0 109100.00000000001 ;
      RECT  71000.0 68500.0 175500.0 69100.0 ;
      RECT  71000.0 28500.000000000004 174100.00000000003 29100.000000000004 ;
      RECT  71000.0 50100.00000000001 172700.0 50700.00000000001 ;
      RECT  68399.99999999999 221400.00000000003 74199.99999999999 222000.00000000003 ;
      RECT  68399.99999999999 241800.0 75600.0 242400.0 ;
      RECT  68399.99999999999 261400.00000000003 76999.99999999999 262000.00000000006 ;
      RECT  68399.99999999999 281800.0 78399.99999999999 282400.00000000006 ;
      RECT  87900.0 131100.0 92100.00000000001 132900.0 ;
      RECT  87900.0 147900.0 92100.00000000001 152100.0 ;
      RECT  18300.0 159900.0 20100.0 164100.0 ;
      RECT  15900.0 128700.00000000001 20100.0 130500.00000000003 ;
      RECT  87900.0 167100.00000000003 92100.00000000001 171300.0 ;
      RECT  59100.0 229500.0 60900.0 233700.0 ;
      RECT  128700.00000000001 167100.00000000003 132900.0 171300.0 ;
      RECT  68700.0 37500.0 70500.0 41700.0 ;
      RECT  30300.0 121500.0 34500.0 125700.0 ;
      RECT  128700.00000000001 186300.0 132900.0 188100.00000000003 ;
      RECT  11100.000000000002 140700.00000000003 15300.0 144900.0 ;
      RECT  179100.00000000003 111900.0 183300.0 113700.0 ;
      RECT  68700.0 119100.00000000001 70500.0 120900.0 ;
      RECT  128700.00000000001 131100.0 132900.0 132900.0 ;
      RECT  107100.00000000001 186300.0 108900.0 188100.00000000003 ;
      RECT  128700.00000000001 241500.0 132900.0 243300.0 ;
      RECT  210300.0 18300.0 212100.00000000003 22500.0 ;
      RECT  -900.0 37500.0 900.0 41700.0 ;
      RECT  128700.00000000001 222300.0 132900.0 226500.0 ;
      RECT  186300.0 111900.0 190500.0 113700.0 ;
      RECT  107100.00000000001 167100.00000000003 108900.0 171300.0 ;
      RECT  18300.0 140700.00000000003 20100.0 144900.0 ;
      RECT  128700.00000000001 203100.00000000003 132900.0 207300.0 ;
      RECT  87900.0 186300.0 92100.00000000001 188100.00000000003 ;
      RECT  59100.0 270300.0 60900.0 274500.0 ;
      RECT  107100.00000000001 131100.0 108900.0 132900.0 ;
      RECT  128700.00000000001 147900.0 132900.0 152100.0 ;
      RECT  188700.00000000003 18300.0 190500.00000000003 22500.0 ;
      RECT  11100.000000000002 159900.0 15300.0 164100.0 ;
      RECT  68700.0 78300.00000000001 70500.0 80100.00000000001 ;
      RECT  3900.0000000000005 123900.0 8100.000000000002 125700.0 ;
      RECT  128700.00000000001 258300.0 132900.0 262500.0 ;
      RECT  107100.00000000001 147900.0 108900.0 152100.0 ;
      RECT  162300.0 241500.0 166500.0 243300.0 ;
      RECT  186300.0 186300.0 190500.0 188100.00000000003 ;
      RECT  183900.0 80700.0 185700.00000000003 82500.0 ;
      RECT  30300.0 179100.00000000003 34500.0 180900.00000000003 ;
      RECT  181500.0 203100.00000000003 183300.0 207300.0 ;
      RECT  186300.0 131100.0 190500.0 132900.0 ;
      RECT  152700.00000000003 203100.00000000003 156900.0 207300.0 ;
      RECT  152700.00000000003 258300.0 156900.0 262500.0 ;
      RECT  152700.00000000003 167100.00000000003 156900.0 171300.0 ;
      RECT  181500.0 222300.0 183300.0 224100.00000000003 ;
      RECT  181500.0 147900.0 183300.0 152100.0 ;
      RECT  162300.0 203100.00000000003 166500.0 207300.0 ;
      RECT  30300.0 140700.00000000003 34500.0 144900.0 ;
      RECT  162300.0 186300.0 166500.0 188100.00000000003 ;
      RECT  181500.0 30300.0 183300.0 32100.0 ;
      RECT  186300.0 47100.0 190500.0 48900.0 ;
      RECT  162300.0 147900.0 166500.0 152100.0 ;
      RECT  162300.0 167100.00000000003 166500.0 171300.0 ;
      RECT  188700.00000000003 30300.0 190500.00000000003 32100.0 ;
      RECT  186300.0 167100.00000000003 190500.0 168900.00000000003 ;
      RECT  152700.00000000003 131100.0 156900.0 132900.0 ;
      RECT  30300.0 195900.0 34500.0 200100.0 ;
      RECT  181500.0 47100.0 183300.0 48900.0 ;
      RECT  152700.00000000003 241500.0 156900.0 243300.0 ;
      RECT  30300.0 159900.0 34500.0 164100.0 ;
      RECT  181500.0 131100.0 183300.0 132900.0 ;
      RECT  162300.0 131100.0 166500.0 132900.0 ;
      RECT  162300.0 222300.0 166500.0 226500.0 ;
      RECT  186300.0 147900.0 190500.0 152100.0 ;
      RECT  188700.00000000003 80700.0 192900.0 82500.0 ;
      RECT  186300.0 241500.0 190500.0 243300.0 ;
      RECT  186300.0 203100.00000000003 190500.0 207300.0 ;
      RECT  181500.0 258300.0 183300.0 262500.0 ;
      RECT  186300.0 258300.0 190500.0 262500.0 ;
      RECT  181500.0 241500.0 183300.0 243300.0 ;
      RECT  152700.00000000003 186300.0 156900.0 188100.00000000003 ;
      RECT  152700.00000000003 222300.0 156900.0 226500.0 ;
      RECT  181500.0 167100.00000000003 183300.0 168900.00000000003 ;
      RECT  186300.0 222300.0 190500.0 224100.00000000003 ;
      RECT  181500.0 186300.0 183300.0 188100.00000000003 ;
      RECT  162300.0 258300.0 166500.0 262500.0 ;
      RECT  152700.00000000003 147900.0 156900.0 152100.0 ;
      RECT  87900.0 140700.00000000003 92100.00000000001 142500.00000000003 ;
      RECT  59100.0 251100.00000000003 60900.0 252900.00000000003 ;
      RECT  107100.00000000001 140700.00000000003 108900.0 142500.00000000003 ;
      RECT  87900.0 195900.0 92100.00000000001 197700.00000000003 ;
      RECT  27900.000000000004 128700.00000000001 29700.000000000004 130500.00000000003 ;
      RECT  188700.00000000003 -900.0 190500.00000000003 900.0 ;
      RECT  59100.0 210300.0 60900.0 212100.00000000003 ;
      RECT  87900.0 176700.00000000003 92100.00000000001 178500.00000000003 ;
      RECT  128700.00000000001 195900.0 132900.0 197700.00000000003 ;
      RECT  107100.00000000001 176700.00000000003 108900.0 178500.00000000003 ;
      RECT  59100.0 289500.0 60900.0 293700.0 ;
      RECT  128700.00000000001 157500.0 132900.0 161700.0 ;
      RECT  68700.0 18300.0 70500.0 20100.0 ;
      RECT  18300.0 150300.0 20100.0 154500.0 ;
      RECT  128700.00000000001 212700.00000000003 132900.0 216900.0 ;
      RECT  11100.000000000002 131100.0 15300.0 135299.99999999997 ;
      RECT  32700.000000000004 128700.00000000001 36900.00000000001 130500.00000000003 ;
      RECT  128700.00000000001 121500.0 132900.0 123300.0 ;
      RECT  11100.000000000002 169500.0 15300.0 171300.0 ;
      RECT  87900.0 157500.0 92100.00000000001 161700.0 ;
      RECT  18300.0 131100.0 20100.0 135299.99999999997 ;
      RECT  18300.0 169500.0 20100.0 171300.0 ;
      RECT  11100.000000000002 150300.0 15300.0 154500.0 ;
      RECT  210300.0 -900.0 212100.00000000003 900.0 ;
      RECT  107100.00000000001 157500.0 108900.0 161700.0 ;
      RECT  68700.0 97500.0 70500.0 101700.0 ;
      RECT  -900.0 18300.0 900.0 20100.0 ;
      RECT  68700.0 59100.0 70500.0 60900.0 ;
      RECT  107100.00000000001 195900.0 108900.0 197700.00000000003 ;
      RECT  128700.00000000001 176700.00000000003 132900.0 178500.00000000003 ;
      RECT  87900.0 121500.0 92100.00000000001 123300.0 ;
      RECT  128700.00000000001 267900.00000000006 132900.0 272100.0 ;
      RECT  128700.00000000001 140700.00000000003 132900.0 142500.00000000003 ;
      RECT  107100.00000000001 121500.0 108900.0 123300.0 ;
      RECT  -900.0 59100.0 900.0 60900.0 ;
      RECT  128700.00000000001 251100.00000000003 132900.0 252900.00000000003 ;
      RECT  128700.00000000001 231900.0 132900.0 233700.00000000003 ;
      RECT  191100.00000000003 198300.0 192900.00000000003 202500.0 ;
      RECT  183900.0 236700.00000000003 188100.0 238500.00000000003 ;
      RECT  191100.00000000003 253500.0 192900.00000000003 257700.0 ;
      RECT  183900.0 207900.0 188100.0 212100.0 ;
      RECT  176700.00000000003 171900.0 180900.0 173700.00000000003 ;
      RECT  191100.00000000003 236700.00000000003 192900.00000000003 238500.00000000003 ;
      RECT  162300.0 231900.0 166500.0 233700.00000000003 ;
      RECT  183900.0 198300.0 188100.0 202500.0 ;
      RECT  191100.00000000003 263100.0 192900.00000000003 267300.0 ;
      RECT  176700.00000000003 152700.00000000003 180900.0 156900.0 ;
      RECT  183900.0 263100.0 188100.0 267300.0 ;
      RECT  183900.0 143100.0 188100.0 147299.99999999997 ;
      RECT  176700.00000000003 243900.0 180900.0 248100.0 ;
      RECT  183900.0 227100.00000000003 188100.0 228900.00000000003 ;
      RECT  176700.00000000003 227100.00000000003 180900.0 228900.00000000003 ;
      RECT  183900.0 133500.0 188100.0 137700.0 ;
      RECT  162300.0 195900.0 166500.0 197700.00000000003 ;
      RECT  191100.00000000003 227100.00000000003 192900.00000000003 228900.00000000003 ;
      RECT  183900.0 243900.0 188100.0 248100.0 ;
      RECT  188700.00000000003 54300.00000000001 192900.0 56100.0 ;
      RECT  191100.00000000003 188700.00000000003 192900.00000000003 192900.0 ;
      RECT  191100.00000000003 143100.0 192900.00000000003 147299.99999999997 ;
      RECT  152700.00000000003 140700.00000000003 156900.0 142500.00000000003 ;
      RECT  27900.000000000004 155100.00000000003 29700.000000000004 159300.0 ;
      RECT  191100.00000000003 162300.0 192900.00000000003 166500.0 ;
      RECT  176700.00000000003 236700.00000000003 180900.0 238500.00000000003 ;
      RECT  176700.00000000003 253500.0 180900.0 257700.0 ;
      RECT  162300.0 157500.0 166500.0 161700.0 ;
      RECT  162300.0 251100.00000000003 166500.0 252900.00000000003 ;
      RECT  152700.00000000003 267900.00000000006 156900.0 272100.0 ;
      RECT  176700.00000000003 207900.0 180900.0 212100.0 ;
      RECT  191100.00000000003 92700.0 192900.00000000003 96900.0 ;
      RECT  152700.00000000003 176700.00000000003 156900.0 178500.00000000003 ;
      RECT  176700.00000000003 126300.00000000001 180900.0 128100.00000000003 ;
      RECT  176700.00000000003 162300.0 180900.0 166500.0 ;
      RECT  176700.00000000003 217500.0 180900.0 221700.0 ;
      RECT  191100.00000000003 181500.0 192900.00000000003 183300.0 ;
      RECT  183900.0 217500.0 188100.0 221700.0 ;
      RECT  27900.000000000004 145500.0 29700.000000000004 149700.0 ;
      RECT  191100.00000000003 126300.00000000001 192900.00000000003 128100.00000000003 ;
      RECT  152700.00000000003 251100.00000000003 156900.0 252900.00000000003 ;
      RECT  191100.00000000003 133500.0 192900.00000000003 137700.0 ;
      RECT  176700.00000000003 133500.0 180900.0 137700.0 ;
      RECT  176700.00000000003 181500.0 180900.0 183300.0 ;
      RECT  162300.0 176700.00000000003 166500.0 178500.00000000003 ;
      RECT  191100.00000000003 207900.0 192900.00000000003 212100.0 ;
      RECT  162300.0 212700.00000000003 166500.0 216900.0 ;
      RECT  183900.0 253500.0 188100.0 257700.0 ;
      RECT  162300.0 121500.0 166500.0 123300.0 ;
      RECT  176700.00000000003 188700.00000000003 180900.0 192900.0 ;
      RECT  183900.0 126300.00000000001 188100.0 128100.00000000003 ;
      RECT  183900.0 181500.0 188100.0 183300.0 ;
      RECT  152700.00000000003 121500.0 156900.0 123300.0 ;
      RECT  176700.00000000003 263100.0 180900.0 267300.0 ;
      RECT  152700.00000000003 231900.0 156900.0 233700.00000000003 ;
      RECT  27900.000000000004 164700.00000000003 29700.000000000004 166500.00000000003 ;
      RECT  162300.0 140700.00000000003 166500.0 142500.00000000003 ;
      RECT  191100.00000000003 243900.0 192900.00000000003 248100.0 ;
      RECT  191100.00000000003 152700.00000000003 192900.00000000003 156900.0 ;
      RECT  27900.000000000004 200700.00000000003 29700.000000000004 204900.0 ;
      RECT  176700.00000000003 198300.0 180900.0 202500.0 ;
      RECT  191100.00000000003 171900.0 192900.00000000003 173700.00000000003 ;
      RECT  27900.000000000004 135900.0 29700.000000000004 140100.0 ;
      RECT  152700.00000000003 157500.0 156900.0 161700.0 ;
      RECT  152700.00000000003 212700.00000000003 156900.0 216900.0 ;
      RECT  183900.0 152700.00000000003 188100.0 156900.0 ;
      RECT  27900.000000000004 174300.0 29700.000000000004 176100.00000000003 ;
      RECT  183900.0 162300.0 188100.0 166500.0 ;
      RECT  176700.00000000003 143100.0 180900.0 147299.99999999997 ;
      RECT  183900.0 188700.00000000003 188100.0 192900.0 ;
      RECT  27900.000000000004 181500.0 29700.000000000004 185700.0 ;
      RECT  191100.00000000003 217500.0 192900.00000000003 221700.0 ;
      RECT  27900.000000000004 191100.00000000003 29700.000000000004 195300.0 ;
      RECT  181500.0 54300.00000000001 185700.0 56100.0 ;
      RECT  162300.0 267900.00000000006 166500.0 272100.0 ;
      RECT  183900.0 171900.0 188100.0 173700.00000000003 ;
      RECT  183900.0 92700.0 188100.0 96900.0 ;
      RECT  152700.00000000003 195900.0 156900.0 197700.00000000003 ;
      RECT  35100.0 205500.0 39300.00000000001 207300.0 ;
      RECT  35100.0 200700.00000000003 36900.0 207300.0 ;
      RECT  32700.000000000004 200700.00000000003 36900.00000000001 204900.0 ;
      RECT  35100.0 133500.0 36900.0 140100.0 ;
      RECT  35100.0 133500.0 39300.00000000001 137700.0 ;
      RECT  32700.000000000004 135900.0 36900.00000000001 140100.0 ;
      RECT  32700.000000000004 135900.0 39300.00000000001 137700.00000000003 ;
      RECT  188700.00000000003 35100.0 190500.00000000003 44100.0 ;
      RECT  188700.00000000003 39900.00000000001 192900.0 44100.00000000001 ;
      RECT  181500.0 35100.0 183300.0 44100.0 ;
      RECT  181500.0 39900.00000000001 185700.0 44100.00000000001 ;
      RECT  32700.000000000004 174300.0 36900.00000000001 176100.00000000003 ;
      RECT  32700.000000000004 164700.00000000003 36900.00000000001 166500.00000000003 ;
      RECT  35100.0 167100.00000000003 39300.00000000001 173700.00000000003 ;
      RECT  35100.0 164700.00000000003 36900.0 176100.00000000003 ;
      RECT  35100.0 186300.0 39300.00000000001 192900.0 ;
      RECT  32700.000000000004 191100.00000000003 36900.00000000001 195300.0 ;
      RECT  32700.000000000004 191100.00000000003 39300.00000000001 192900.00000000003 ;
      RECT  35100.0 181500.0 36900.0 195300.0 ;
      RECT  32700.000000000004 181500.0 36900.00000000001 185700.0 ;
      RECT  35100.0 145500.0 36900.0 159300.0 ;
      RECT  32700.000000000004 155100.00000000003 36900.00000000001 159300.0 ;
      RECT  32700.000000000004 145500.0 36900.00000000001 149700.0 ;
      RECT  35100.0 147900.0 39300.00000000001 154500.0 ;
      RECT  32700.000000000004 147900.0 39300.00000000001 149700.00000000003 ;
      RECT  15900.0 159900.0 17700.0 161700.00000000003 ;
      RECT  16800.0 159900.0 19200.000000000004 161700.00000000003 ;
      RECT  18300.0 159900.0 20100.0 161700.00000000003 ;
      RECT  15900.0 128700.00000000001 17700.0 130500.00000000003 ;
      RECT  59100.0 227100.00000000003 60900.0 228900.00000000003 ;
      RECT  59100.0 228000.0 60900.0 230400.0 ;
      RECT  59100.0 229500.0 60900.0 231300.0 ;
      RECT  59100.0 227100.00000000003 60900.0 228900.00000000003 ;
      RECT  68700.0 35100.0 70500.0 36900.0 ;
      RECT  68700.0 36000.0 70500.0 38400.0 ;
      RECT  68700.0 37500.0 70500.0 39300.0 ;
      RECT  68700.0 35100.0 70500.0 36900.0 ;
      RECT  13500.0 140700.00000000003 15300.0 142500.00000000003 ;
      RECT  104700.0 186300.0 106500.0 188100.00000000003 ;
      RECT  105600.00000000001 186300.0 108000.00000000001 188100.00000000003 ;
      RECT  107100.00000000001 186300.0 108900.0 188100.00000000003 ;
      RECT  104700.0 186300.0 106500.0 188100.00000000003 ;
      RECT  131100.0 243900.0 132900.0 245700.00000000003 ;
      RECT  131100.0 242400.0 132900.0 244800.0 ;
      RECT  131100.0 241500.0 132900.0 243300.0 ;
      RECT  131100.0 243900.0 132900.0 245700.00000000003 ;
      RECT  210300.0 23100.0 212100.00000000003 24900.000000000004 ;
      RECT  210300.0 21600.0 212100.00000000003 24000.0 ;
      RECT  210300.0 20700.000000000004 212100.00000000003 22500.000000000004 ;
      RECT  210300.0 23100.0 212100.00000000003 24900.000000000004 ;
      RECT  -900.0 42300.00000000001 900.0 44100.0 ;
      RECT  -900.0 40800.00000000001 900.0 43200.0 ;
      RECT  -900.0 39900.00000000001 900.0 41700.0 ;
      RECT  -900.0 42300.00000000001 900.0 44100.0 ;
      RECT  104700.0 167100.00000000003 106500.0 168900.00000000003 ;
      RECT  105600.00000000001 167100.00000000003 108000.00000000001 168900.00000000003 ;
      RECT  107100.00000000001 167100.00000000003 108900.0 168900.00000000003 ;
      RECT  104700.0 167100.00000000003 106500.0 168900.00000000003 ;
      RECT  15900.0 140700.00000000003 17700.0 142500.00000000003 ;
      RECT  16800.0 140700.00000000003 19200.000000000004 142500.00000000003 ;
      RECT  18300.0 140700.00000000003 20100.0 142500.00000000003 ;
      RECT  104700.0 131100.0 106500.0 132900.0 ;
      RECT  105600.00000000001 131100.0 108000.00000000001 132900.0 ;
      RECT  107100.00000000001 131100.0 108900.0 132900.0 ;
      RECT  104700.0 131100.0 106500.0 132900.0 ;
      RECT  188700.00000000003 15900.0 190500.00000000003 17700.0 ;
      RECT  188700.00000000003 16800.0 190500.00000000003 19200.000000000004 ;
      RECT  188700.00000000003 18300.0 190500.00000000003 20100.0 ;
      RECT  188700.00000000003 15900.0 190500.00000000003 17700.0 ;
      RECT  13500.0 159900.0 15300.0 161700.00000000003 ;
      RECT  68700.0 80700.0 70500.0 82500.0 ;
      RECT  68700.0 79200.0 70500.0 81600.00000000001 ;
      RECT  68700.0 78300.00000000001 70500.0 80100.00000000001 ;
      RECT  68700.0 80700.0 70500.0 82500.0 ;
      RECT  3900.0000000000005 121500.0 5700.0 123300.0 ;
      RECT  3900.0000000000005 122400.0 5700.0 124800.00000000001 ;
      RECT  3900.0000000000005 123900.0 5700.0 125700.0 ;
      RECT  3900.0000000000005 121500.0 5700.0 123300.0 ;
      RECT  131100.0 255900.0 132900.0 257700.0 ;
      RECT  131100.0 256800.0 132900.0 259200.0 ;
      RECT  131100.0 258300.0 132900.0 260100.00000000003 ;
      RECT  131100.0 255900.0 132900.0 257700.0 ;
      RECT  104700.0 147900.0 106500.0 149700.00000000003 ;
      RECT  105600.00000000001 147900.0 108000.00000000001 149700.00000000003 ;
      RECT  107100.00000000001 147900.0 108900.0 149700.00000000003 ;
      RECT  104700.0 147900.0 106500.0 149700.00000000003 ;
      RECT  164700.00000000003 243900.0 166500.00000000003 245700.00000000003 ;
      RECT  164700.00000000003 242400.0 166500.00000000003 244800.0 ;
      RECT  164700.00000000003 241500.0 166500.00000000003 243300.0 ;
      RECT  164700.00000000003 243900.0 166500.00000000003 245700.00000000003 ;
      RECT  188700.00000000003 186300.0 190500.00000000003 188100.00000000003 ;
      RECT  179100.00000000003 205500.0 180900.00000000003 207300.0 ;
      RECT  180000.0 205500.0 182400.0 207300.0 ;
      RECT  181500.0 205500.0 183300.0 207300.0 ;
      RECT  155100.00000000003 263100.0 156900.00000000003 264900.00000000006 ;
      RECT  155100.00000000003 261600.00000000003 156900.00000000003 264000.0 ;
      RECT  155100.00000000003 260700.0 156900.00000000003 262500.0 ;
      RECT  155100.00000000003 263100.0 156900.00000000003 264900.00000000006 ;
      RECT  179100.00000000003 222300.0 180900.00000000003 224100.00000000003 ;
      RECT  180000.0 222300.0 182400.0 224100.00000000003 ;
      RECT  181500.0 222300.0 183300.0 224100.00000000003 ;
      RECT  32700.000000000004 140700.00000000003 34500.0 142500.00000000003 ;
      RECT  179100.00000000003 30300.0 180900.00000000003 32100.0 ;
      RECT  180000.0 30300.0 182400.0 32100.0 ;
      RECT  181500.0 30300.0 183300.0 32100.0 ;
      RECT  188700.00000000003 47100.0 190500.00000000003 48900.0 ;
      RECT  188700.00000000003 30300.0 190500.00000000003 32100.0 ;
      RECT  179100.00000000003 47100.0 180900.00000000003 48900.0 ;
      RECT  180000.0 47100.0 182400.0 48900.0 ;
      RECT  181500.0 47100.0 183300.0 48900.0 ;
      RECT  155100.00000000003 243900.0 156900.00000000003 245700.00000000003 ;
      RECT  155100.00000000003 242400.0 156900.00000000003 244800.0 ;
      RECT  155100.00000000003 241500.0 156900.00000000003 243300.0 ;
      RECT  155100.00000000003 243900.0 156900.00000000003 245700.00000000003 ;
      RECT  32700.000000000004 159900.0 34500.0 161700.00000000003 ;
      RECT  188700.00000000003 241500.0 190500.00000000003 243300.0 ;
      RECT  188700.00000000003 205500.0 190500.00000000003 207300.0 ;
      RECT  179100.00000000003 260700.0 180900.00000000003 262500.0 ;
      RECT  180000.0 260700.0 182400.0 262500.0 ;
      RECT  181500.0 260700.0 183300.0 262500.0 ;
      RECT  188700.00000000003 260700.0 190500.00000000003 262500.0 ;
      RECT  179100.00000000003 241500.0 180900.00000000003 243300.0 ;
      RECT  180000.0 241500.0 182400.0 243300.0 ;
      RECT  181500.0 241500.0 183300.0 243300.0 ;
      RECT  188700.00000000003 222300.0 190500.00000000003 224100.00000000003 ;
      RECT  179100.00000000003 186300.0 180900.00000000003 188100.00000000003 ;
      RECT  180000.0 186300.0 182400.0 188100.00000000003 ;
      RECT  181500.0 186300.0 183300.0 188100.00000000003 ;
      RECT  164700.00000000003 263100.0 166500.00000000003 264900.00000000006 ;
      RECT  164700.00000000003 261600.00000000003 166500.00000000003 264000.0 ;
      RECT  164700.00000000003 260700.0 166500.00000000003 262500.0 ;
      RECT  164700.00000000003 263100.0 166500.00000000003 264900.00000000006 ;
      RECT  87900.0 143100.0 89700.0 144900.0 ;
      RECT  87900.0 141600.0 89700.0 144000.0 ;
      RECT  87900.0 140700.00000000003 89700.0 142500.00000000003 ;
      RECT  87900.0 143100.0 89700.0 144900.0 ;
      RECT  107100.00000000001 143100.0 108900.0 144900.0 ;
      RECT  107100.00000000001 141600.0 108900.0 144000.0 ;
      RECT  107100.00000000001 140700.00000000003 108900.0 142500.00000000003 ;
      RECT  107100.00000000001 143100.0 108900.0 144900.0 ;
      RECT  87900.0 193500.0 89700.0 195300.0 ;
      RECT  87900.0 194400.0 89700.0 196800.0 ;
      RECT  87900.0 195900.0 89700.0 197700.00000000003 ;
      RECT  87900.0 193500.0 89700.0 195300.0 ;
      RECT  27900.000000000004 128700.00000000001 29700.000000000004 130500.00000000003 ;
      RECT  191100.00000000003 -900.0 192900.00000000003 900.0 ;
      RECT  189600.00000000003 -900.0 192000.00000000003 900.0 ;
      RECT  188700.00000000003 -900.0 190500.00000000003 900.0 ;
      RECT  59100.0 210300.0 60900.0 212100.00000000003 ;
      RECT  87900.0 174300.0 89700.0 176100.00000000003 ;
      RECT  87900.0 175200.00000000003 89700.0 177600.00000000003 ;
      RECT  87900.0 176700.00000000003 89700.0 178500.00000000003 ;
      RECT  87900.0 174300.0 89700.0 176100.00000000003 ;
      RECT  128700.00000000001 193500.0 130500.00000000003 195300.0 ;
      RECT  128700.00000000001 194400.0 130500.00000000003 196800.0 ;
      RECT  128700.00000000001 195900.0 130500.00000000003 197700.00000000003 ;
      RECT  128700.00000000001 193500.0 130500.00000000003 195300.0 ;
      RECT  107100.00000000001 174300.0 108900.0 176100.00000000003 ;
      RECT  107100.00000000001 175200.00000000003 108900.0 177600.00000000003 ;
      RECT  107100.00000000001 176700.00000000003 108900.0 178500.00000000003 ;
      RECT  107100.00000000001 174300.0 108900.0 176100.00000000003 ;
      RECT  128700.00000000001 155100.00000000003 130500.00000000003 156900.00000000003 ;
      RECT  128700.00000000001 156000.0 130500.00000000003 158400.0 ;
      RECT  128700.00000000001 157500.0 130500.00000000003 159300.0 ;
      RECT  128700.00000000001 155100.00000000003 130500.00000000003 156900.00000000003 ;
      RECT  18300.0 152700.00000000003 20100.0 154500.00000000003 ;
      RECT  11100.000000000002 133500.0 12900.000000000002 135300.0 ;
      RECT  37500.0 128700.00000000001 39300.0 130500.00000000003 ;
      RECT  36000.0 128700.00000000001 38400.0 130500.00000000003 ;
      RECT  37500.0 126300.00000000001 39300.0 128100.00000000003 ;
      RECT  37500.0 127200.0 39300.0 129600.0 ;
      RECT  35100.0 128700.00000000001 36900.0 130500.00000000003 ;
      RECT  37500.0 126300.00000000001 39300.0 128100.00000000003 ;
      RECT  128700.00000000001 123900.0 130500.00000000003 125700.0 ;
      RECT  128700.00000000001 122400.0 130500.00000000003 124800.00000000001 ;
      RECT  128700.00000000001 121500.0 130500.00000000003 123300.0 ;
      RECT  128700.00000000001 123900.0 130500.00000000003 125700.0 ;
      RECT  11100.000000000002 171900.0 12900.000000000002 173700.00000000003 ;
      RECT  11100.000000000002 170400.0 12900.000000000002 172800.0 ;
      RECT  11100.000000000002 169500.0 12900.000000000002 171300.0 ;
      RECT  11100.000000000002 171900.0 12900.000000000002 173700.00000000003 ;
      RECT  87900.0 162300.0 89700.0 164100.00000000003 ;
      RECT  87900.0 160800.0 89700.0 163200.00000000003 ;
      RECT  87900.0 159900.0 89700.0 161700.00000000003 ;
      RECT  87900.0 162300.0 89700.0 164100.00000000003 ;
      RECT  18300.0 133500.0 20100.0 135300.0 ;
      RECT  18300.0 171900.0 20100.0 173700.00000000003 ;
      RECT  18300.0 170400.0 20100.0 172800.0 ;
      RECT  18300.0 169500.0 20100.0 171300.0 ;
      RECT  18300.0 171900.0 20100.0 173700.00000000003 ;
      RECT  11100.000000000002 150300.0 12900.000000000002 152100.00000000003 ;
      RECT  210300.0 -900.0 212100.00000000003 900.0 ;
      RECT  107100.00000000001 155100.00000000003 108900.0 156900.00000000003 ;
      RECT  107100.00000000001 156000.0 108900.0 158400.0 ;
      RECT  107100.00000000001 157500.0 108900.0 159300.0 ;
      RECT  107100.00000000001 155100.00000000003 108900.0 156900.00000000003 ;
      RECT  107100.00000000001 193500.0 108900.0 195300.0 ;
      RECT  107100.00000000001 194400.0 108900.0 196800.0 ;
      RECT  107100.00000000001 195900.0 108900.0 197700.00000000003 ;
      RECT  107100.00000000001 193500.0 108900.0 195300.0 ;
      RECT  128700.00000000001 174300.0 130500.00000000003 176100.00000000003 ;
      RECT  128700.00000000001 175200.00000000003 130500.00000000003 177600.00000000003 ;
      RECT  128700.00000000001 176700.00000000003 130500.00000000003 178500.00000000003 ;
      RECT  128700.00000000001 174300.0 130500.00000000003 176100.00000000003 ;
      RECT  87900.0 123900.0 89700.0 125700.0 ;
      RECT  87900.0 122400.0 89700.0 124800.00000000001 ;
      RECT  87900.0 121500.0 89700.0 123300.0 ;
      RECT  87900.0 123900.0 89700.0 125700.0 ;
      RECT  128700.00000000001 143100.0 130500.00000000003 144900.0 ;
      RECT  128700.00000000001 141600.0 130500.00000000003 144000.0 ;
      RECT  128700.00000000001 140700.00000000003 130500.00000000003 142500.00000000003 ;
      RECT  128700.00000000001 143100.0 130500.00000000003 144900.0 ;
      RECT  107100.00000000001 123900.0 108900.0 125700.0 ;
      RECT  107100.00000000001 122400.0 108900.0 124800.00000000001 ;
      RECT  107100.00000000001 121500.0 108900.0 123300.0 ;
      RECT  107100.00000000001 123900.0 108900.0 125700.0 ;
      RECT  191100.00000000003 198300.0 192900.00000000003 200100.00000000003 ;
      RECT  183900.0 236700.00000000003 185700.00000000003 238500.00000000003 ;
      RECT  191100.00000000003 255900.0 192900.00000000003 257700.0 ;
      RECT  191100.00000000003 236700.00000000003 192900.00000000003 238500.00000000003 ;
      RECT  183900.0 200700.00000000003 185700.00000000003 202500.00000000003 ;
      RECT  191100.00000000003 267900.00000000006 192900.00000000003 269700.00000000006 ;
      RECT  191100.00000000003 266400.00000000006 192900.00000000003 268800.0 ;
      RECT  191100.00000000003 265500.0 192900.00000000003 267300.0 ;
      RECT  191100.00000000003 267900.00000000006 192900.00000000003 269700.00000000006 ;
      RECT  183900.0 263100.0 185700.00000000003 264900.00000000006 ;
      RECT  176700.00000000003 248700.00000000003 178500.00000000003 250500.00000000003 ;
      RECT  176700.00000000003 247200.00000000003 178500.00000000003 249600.00000000003 ;
      RECT  176700.00000000003 246300.0 178500.00000000003 248100.00000000003 ;
      RECT  176700.00000000003 248700.00000000003 178500.00000000003 250500.00000000003 ;
      RECT  183900.0 229500.0 185700.00000000003 231300.0 ;
      RECT  183900.0 228000.0 185700.00000000003 230400.0 ;
      RECT  183900.0 227100.00000000003 185700.00000000003 228900.00000000003 ;
      RECT  183900.0 229500.0 185700.00000000003 231300.0 ;
      RECT  176700.00000000003 229500.0 178500.00000000003 231300.0 ;
      RECT  176700.00000000003 228000.0 178500.00000000003 230400.0 ;
      RECT  176700.00000000003 227100.00000000003 178500.00000000003 228900.00000000003 ;
      RECT  176700.00000000003 229500.0 178500.00000000003 231300.0 ;
      RECT  162300.0 193500.0 164100.00000000003 195300.0 ;
      RECT  162300.0 194400.0 164100.00000000003 196800.0 ;
      RECT  162300.0 195900.0 164100.00000000003 197700.00000000003 ;
      RECT  162300.0 193500.0 164100.00000000003 195300.0 ;
      RECT  191100.00000000003 229500.0 192900.00000000003 231300.0 ;
      RECT  191100.00000000003 228000.0 192900.00000000003 230400.0 ;
      RECT  191100.00000000003 227100.00000000003 192900.00000000003 228900.00000000003 ;
      RECT  191100.00000000003 229500.0 192900.00000000003 231300.0 ;
      RECT  183900.0 248700.00000000003 185700.00000000003 250500.00000000003 ;
      RECT  183900.0 247200.00000000003 185700.00000000003 249600.00000000003 ;
      RECT  183900.0 246300.0 185700.00000000003 248100.00000000003 ;
      RECT  183900.0 248700.00000000003 185700.00000000003 250500.00000000003 ;
      RECT  191100.00000000003 56700.0 192900.00000000003 58500.0 ;
      RECT  191100.00000000003 55200.0 192900.00000000003 57600.0 ;
      RECT  191100.00000000003 54300.00000000001 192900.00000000003 56100.0 ;
      RECT  191100.00000000003 56700.0 192900.00000000003 58500.0 ;
      RECT  152700.00000000003 143100.0 154500.00000000003 144900.0 ;
      RECT  152700.00000000003 141600.0 154500.00000000003 144000.0 ;
      RECT  152700.00000000003 140700.00000000003 154500.00000000003 142500.00000000003 ;
      RECT  152700.00000000003 143100.0 154500.00000000003 144900.0 ;
      RECT  181500.0 236700.00000000003 183300.0 238500.00000000003 ;
      RECT  180000.0 236700.00000000003 182400.0 238500.00000000003 ;
      RECT  179100.00000000003 236700.00000000003 180900.00000000003 238500.00000000003 ;
      RECT  179100.00000000003 251100.00000000003 180900.00000000003 252900.00000000003 ;
      RECT  179100.00000000003 252000.0 180900.00000000003 254400.0 ;
      RECT  179100.00000000003 253500.0 180900.00000000003 255300.0 ;
      RECT  179100.00000000003 251100.00000000003 180900.00000000003 252900.00000000003 ;
      RECT  162300.0 155100.00000000003 164100.00000000003 156900.00000000003 ;
      RECT  162300.0 156000.0 164100.00000000003 158400.0 ;
      RECT  162300.0 157500.0 164100.00000000003 159300.0 ;
      RECT  162300.0 155100.00000000003 164100.00000000003 156900.00000000003 ;
      RECT  152700.00000000003 174300.0 154500.00000000003 176100.00000000003 ;
      RECT  152700.00000000003 175200.00000000003 154500.00000000003 177600.00000000003 ;
      RECT  152700.00000000003 176700.00000000003 154500.00000000003 178500.00000000003 ;
      RECT  152700.00000000003 174300.0 154500.00000000003 176100.00000000003 ;
      RECT  174300.0 219900.0 176100.00000000003 221700.00000000003 ;
      RECT  175200.00000000003 219900.0 177600.00000000003 221700.00000000003 ;
      RECT  176700.00000000003 219900.0 178500.00000000003 221700.00000000003 ;
      RECT  183900.0 219900.0 185700.00000000003 221700.00000000003 ;
      RECT  27900.000000000004 147900.0 29700.000000000004 149700.00000000003 ;
      RECT  162300.0 174300.0 164100.00000000003 176100.00000000003 ;
      RECT  162300.0 175200.00000000003 164100.00000000003 177600.00000000003 ;
      RECT  162300.0 176700.00000000003 164100.00000000003 178500.00000000003 ;
      RECT  162300.0 174300.0 164100.00000000003 176100.00000000003 ;
      RECT  183900.0 255900.0 185700.00000000003 257700.0 ;
      RECT  162300.0 123900.0 164100.00000000003 125700.0 ;
      RECT  162300.0 122400.0 164100.00000000003 124800.00000000001 ;
      RECT  162300.0 121500.0 164100.00000000003 123300.0 ;
      RECT  162300.0 123900.0 164100.00000000003 125700.0 ;
      RECT  152700.00000000003 123900.0 154500.00000000003 125700.0 ;
      RECT  152700.00000000003 122400.0 154500.00000000003 124800.00000000001 ;
      RECT  152700.00000000003 121500.0 154500.00000000003 123300.0 ;
      RECT  152700.00000000003 123900.0 154500.00000000003 125700.0 ;
      RECT  179100.00000000003 267900.00000000006 180900.00000000003 269700.00000000006 ;
      RECT  179100.00000000003 266400.00000000006 180900.00000000003 268800.0 ;
      RECT  179100.00000000003 265500.0 180900.00000000003 267300.0 ;
      RECT  179100.00000000003 267900.00000000006 180900.00000000003 269700.00000000006 ;
      RECT  27900.000000000004 164700.00000000003 29700.000000000004 166500.00000000003 ;
      RECT  162300.0 143100.0 164100.00000000003 144900.0 ;
      RECT  162300.0 141600.0 164100.00000000003 144000.0 ;
      RECT  162300.0 140700.00000000003 164100.00000000003 142500.00000000003 ;
      RECT  162300.0 143100.0 164100.00000000003 144900.0 ;
      RECT  191100.00000000003 248700.00000000003 192900.00000000003 250500.00000000003 ;
      RECT  191100.00000000003 247200.00000000003 192900.00000000003 249600.00000000003 ;
      RECT  191100.00000000003 246300.0 192900.00000000003 248100.00000000003 ;
      RECT  191100.00000000003 248700.00000000003 192900.00000000003 250500.00000000003 ;
      RECT  181500.0 198300.0 183300.0 200100.00000000003 ;
      RECT  180000.0 198300.0 182400.0 200100.00000000003 ;
      RECT  179100.00000000003 198300.0 180900.00000000003 200100.00000000003 ;
      RECT  152700.00000000003 155100.00000000003 154500.00000000003 156900.00000000003 ;
      RECT  152700.00000000003 156000.0 154500.00000000003 158400.0 ;
      RECT  152700.00000000003 157500.0 154500.00000000003 159300.0 ;
      RECT  152700.00000000003 155100.00000000003 154500.00000000003 156900.00000000003 ;
      RECT  191100.00000000003 217500.0 192900.00000000003 219300.0 ;
      RECT  181500.0 56700.0 183300.0 58500.0 ;
      RECT  181500.0 55200.0 183300.0 57600.0 ;
      RECT  181500.0 54300.00000000001 183300.0 56100.0 ;
      RECT  181500.0 56700.0 183300.0 58500.0 ;
      RECT  152700.00000000003 193500.0 154500.00000000003 195300.0 ;
      RECT  152700.00000000003 194400.0 154500.00000000003 196800.0 ;
      RECT  152700.00000000003 195900.0 154500.00000000003 197700.00000000003 ;
      RECT  152700.00000000003 193500.0 154500.00000000003 195300.0 ;
      RECT  181600.00000000003 131200.0 182400.0 132000.0 ;
      RECT  188400.0 131200.0 189200.0 132000.0 ;
      RECT  181600.00000000003 131200.0 182400.0 132000.0 ;
      RECT  188400.0 131200.0 189200.0 132000.0 ;
      RECT  181600.00000000003 149600.00000000003 182400.0 150400.0 ;
      RECT  188400.0 149600.00000000003 189200.0 150400.0 ;
      RECT  181600.00000000003 149600.00000000003 182400.0 150400.0 ;
      RECT  188400.0 149600.00000000003 189200.0 150400.0 ;
      RECT  181600.00000000003 168000.0 182400.0 168800.0 ;
      RECT  188400.0 168000.0 189200.0 168800.0 ;
      RECT  181600.00000000003 168000.0 182400.0 168800.0 ;
      RECT  188400.0 168000.0 189200.0 168800.0 ;
      RECT  181600.00000000003 186399.99999999997 182400.0 187200.0 ;
      RECT  188400.0 186399.99999999997 189200.0 187200.0 ;
      RECT  181600.00000000003 186399.99999999997 182400.0 187200.0 ;
      RECT  188400.0 186399.99999999997 189200.0 187200.0 ;
      RECT  181600.00000000003 204800.0 182400.0 205600.00000000003 ;
      RECT  188400.0 204800.0 189200.0 205600.00000000003 ;
      RECT  181600.00000000003 204800.0 182400.0 205600.00000000003 ;
      RECT  188400.0 204800.0 189200.0 205600.00000000003 ;
      RECT  181600.00000000003 223200.0 182400.0 224000.0 ;
      RECT  188400.0 223200.0 189200.0 224000.0 ;
      RECT  181600.00000000003 223200.0 182400.0 224000.0 ;
      RECT  188400.0 223200.0 189200.0 224000.0 ;
      RECT  181600.00000000003 241600.00000000003 182400.0 242399.99999999997 ;
      RECT  188400.0 241600.00000000003 189200.0 242399.99999999997 ;
      RECT  181600.00000000003 241600.00000000003 182400.0 242399.99999999997 ;
      RECT  188400.0 241600.00000000003 189200.0 242399.99999999997 ;
      RECT  181600.00000000003 260000.0 182400.0 260800.0 ;
      RECT  188400.0 260000.0 189200.0 260800.0 ;
      RECT  181600.00000000003 260000.0 182400.0 260800.0 ;
      RECT  188400.0 260000.0 189200.0 260800.0 ;
      RECT  178200.0 126600.00000000001 179000.0 127400.0 ;
      RECT  185000.0 126600.00000000001 185800.0 127400.0 ;
      RECT  185000.0 126600.00000000001 185800.0 127400.0 ;
      RECT  191800.0 126600.00000000001 192600.00000000003 127400.0 ;
      RECT  178200.0 135800.0 179000.0 136600.00000000003 ;
      RECT  185000.0 135800.0 185800.0 136600.00000000003 ;
      RECT  185000.0 135800.0 185800.0 136600.00000000003 ;
      RECT  191800.0 135800.0 192600.00000000003 136600.00000000003 ;
      RECT  178200.0 145000.0 179000.0 145800.0 ;
      RECT  185000.0 145000.0 185800.0 145800.0 ;
      RECT  185000.0 145000.0 185800.0 145800.0 ;
      RECT  191800.0 145000.0 192600.00000000003 145800.0 ;
      RECT  178200.0 154200.0 179000.0 155000.0 ;
      RECT  185000.0 154200.0 185800.0 155000.0 ;
      RECT  185000.0 154200.0 185800.0 155000.0 ;
      RECT  191800.0 154200.0 192600.00000000003 155000.0 ;
      RECT  178200.0 163399.99999999997 179000.0 164200.0 ;
      RECT  185000.0 163399.99999999997 185800.0 164200.0 ;
      RECT  185000.0 163399.99999999997 185800.0 164200.0 ;
      RECT  191800.0 163399.99999999997 192600.00000000003 164200.0 ;
      RECT  178200.0 172600.00000000003 179000.0 173399.99999999997 ;
      RECT  185000.0 172600.00000000003 185800.0 173399.99999999997 ;
      RECT  185000.0 172600.00000000003 185800.0 173399.99999999997 ;
      RECT  191800.0 172600.00000000003 192600.00000000003 173399.99999999997 ;
      RECT  178200.0 181800.0 179000.0 182600.00000000003 ;
      RECT  185000.0 181800.0 185800.0 182600.00000000003 ;
      RECT  185000.0 181800.0 185800.0 182600.00000000003 ;
      RECT  191800.0 181800.0 192600.00000000003 182600.00000000003 ;
      RECT  178200.0 191000.0 179000.0 191800.0 ;
      RECT  185000.0 191000.0 185800.0 191800.0 ;
      RECT  185000.0 191000.0 185800.0 191800.0 ;
      RECT  191800.0 191000.0 192600.00000000003 191800.0 ;
      RECT  178200.0 200200.0 179000.0 201000.0 ;
      RECT  185000.0 200200.0 185800.0 201000.0 ;
      RECT  185000.0 200200.0 185800.0 201000.0 ;
      RECT  191800.0 200200.0 192600.00000000003 201000.0 ;
      RECT  178200.0 209399.99999999997 179000.0 210200.0 ;
      RECT  185000.0 209399.99999999997 185800.0 210200.0 ;
      RECT  185000.0 209399.99999999997 185800.0 210200.0 ;
      RECT  191800.0 209399.99999999997 192600.00000000003 210200.0 ;
      RECT  178200.0 218600.00000000003 179000.0 219399.99999999997 ;
      RECT  185000.0 218600.00000000003 185800.0 219399.99999999997 ;
      RECT  185000.0 218600.00000000003 185800.0 219399.99999999997 ;
      RECT  191800.0 218600.00000000003 192600.00000000003 219399.99999999997 ;
      RECT  178200.0 227800.0 179000.0 228600.00000000003 ;
      RECT  185000.0 227800.0 185800.0 228600.00000000003 ;
      RECT  185000.0 227800.0 185800.0 228600.00000000003 ;
      RECT  191800.0 227800.0 192600.00000000003 228600.00000000003 ;
      RECT  178200.0 237000.0 179000.0 237800.0 ;
      RECT  185000.0 237000.0 185800.0 237800.0 ;
      RECT  185000.0 237000.0 185800.0 237800.0 ;
      RECT  191800.0 237000.0 192600.00000000003 237800.0 ;
      RECT  178200.0 246200.0 179000.0 247000.0 ;
      RECT  185000.0 246200.0 185800.0 247000.0 ;
      RECT  185000.0 246200.0 185800.0 247000.0 ;
      RECT  191800.0 246200.0 192600.00000000003 247000.0 ;
      RECT  178200.0 255399.99999999997 179000.0 256200.0 ;
      RECT  185000.0 255399.99999999997 185800.0 256200.0 ;
      RECT  185000.0 255399.99999999997 185800.0 256200.0 ;
      RECT  191800.0 255399.99999999997 192600.00000000003 256200.0 ;
      RECT  178200.0 264600.0 179000.0 265400.00000000006 ;
      RECT  185000.0 264600.0 185800.0 265400.00000000006 ;
      RECT  185000.0 264600.0 185800.0 265400.00000000006 ;
      RECT  191800.0 264600.0 192600.00000000003 265400.00000000006 ;
      RECT  181700.0 131300.0 182300.0 131900.0 ;
      RECT  188500.0 131300.0 189100.00000000003 131900.0 ;
      RECT  181700.0 149700.0 182300.0 150300.0 ;
      RECT  188500.0 149700.0 189100.00000000003 150300.0 ;
      RECT  181700.0 168100.00000000003 182300.0 168700.0 ;
      RECT  188500.0 168100.00000000003 189100.00000000003 168700.0 ;
      RECT  181700.0 186500.0 182300.0 187100.00000000003 ;
      RECT  188500.0 186500.0 189100.00000000003 187100.00000000003 ;
      RECT  181700.0 204899.99999999997 182300.0 205500.0 ;
      RECT  188500.0 204899.99999999997 189100.00000000003 205500.0 ;
      RECT  181700.0 223300.0 182300.0 223899.99999999997 ;
      RECT  188500.0 223300.0 189100.00000000003 223899.99999999997 ;
      RECT  181700.0 241700.0 182300.0 242300.0 ;
      RECT  188500.0 241700.0 189100.00000000003 242300.0 ;
      RECT  181700.0 260100.00000000003 182300.0 260700.0 ;
      RECT  188500.0 260100.00000000003 189100.00000000003 260700.0 ;
      RECT  178300.0 126700.0 178900.0 127300.00000000001 ;
      RECT  185100.00000000003 126700.0 185700.0 127300.00000000001 ;
      RECT  191900.0 126700.0 192500.0 127300.00000000001 ;
      RECT  178300.0 135900.0 178900.0 136500.0 ;
      RECT  185100.00000000003 135900.0 185700.0 136500.0 ;
      RECT  191900.0 135900.0 192500.0 136500.0 ;
      RECT  178300.0 145100.00000000003 178900.0 145700.0 ;
      RECT  185100.00000000003 145100.00000000003 185700.0 145700.0 ;
      RECT  191900.0 145100.00000000003 192500.0 145700.0 ;
      RECT  178300.0 154300.0 178900.0 154899.99999999997 ;
      RECT  185100.00000000003 154300.0 185700.0 154899.99999999997 ;
      RECT  191900.0 154300.0 192500.0 154899.99999999997 ;
      RECT  178300.0 163500.0 178900.0 164100.00000000003 ;
      RECT  185100.00000000003 163500.0 185700.0 164100.00000000003 ;
      RECT  191900.0 163500.0 192500.0 164100.00000000003 ;
      RECT  178300.0 172700.0 178900.0 173300.0 ;
      RECT  185100.00000000003 172700.0 185700.0 173300.0 ;
      RECT  191900.0 172700.0 192500.0 173300.0 ;
      RECT  178300.0 181899.99999999997 178900.0 182500.0 ;
      RECT  185100.00000000003 181899.99999999997 185700.0 182500.0 ;
      RECT  191900.0 181899.99999999997 192500.0 182500.0 ;
      RECT  178300.0 191100.00000000003 178900.0 191700.0 ;
      RECT  185100.00000000003 191100.00000000003 185700.0 191700.0 ;
      RECT  191900.0 191100.00000000003 192500.0 191700.0 ;
      RECT  178300.0 200300.0 178900.0 200899.99999999997 ;
      RECT  185100.00000000003 200300.0 185700.0 200899.99999999997 ;
      RECT  191900.0 200300.0 192500.0 200899.99999999997 ;
      RECT  178300.0 209500.0 178900.0 210100.00000000003 ;
      RECT  185100.00000000003 209500.0 185700.0 210100.00000000003 ;
      RECT  191900.0 209500.0 192500.0 210100.00000000003 ;
      RECT  178300.0 218700.0 178900.0 219300.0 ;
      RECT  185100.00000000003 218700.0 185700.0 219300.0 ;
      RECT  191900.0 218700.0 192500.0 219300.0 ;
      RECT  178300.0 227899.99999999997 178900.0 228500.0 ;
      RECT  185100.00000000003 227899.99999999997 185700.0 228500.0 ;
      RECT  191900.0 227899.99999999997 192500.0 228500.0 ;
      RECT  178300.0 237100.00000000003 178900.0 237700.0 ;
      RECT  185100.00000000003 237100.00000000003 185700.0 237700.0 ;
      RECT  191900.0 237100.00000000003 192500.0 237700.0 ;
      RECT  178300.0 246300.0 178900.0 246899.99999999997 ;
      RECT  185100.00000000003 246300.0 185700.0 246899.99999999997 ;
      RECT  191900.0 246300.0 192500.0 246899.99999999997 ;
      RECT  178300.0 255500.0 178900.0 256100.00000000003 ;
      RECT  185100.00000000003 255500.0 185700.0 256100.00000000003 ;
      RECT  191900.0 255500.0 192500.0 256100.00000000003 ;
      RECT  178300.0 264700.0 178900.0 265300.0 ;
      RECT  185100.00000000003 264700.0 185700.0 265300.0 ;
      RECT  191900.0 264700.0 192500.0 265300.0 ;
      RECT  181400.0 112000.00000000001 182200.0 112800.00000000001 ;
      RECT  181400.0 112000.00000000001 182200.0 112800.00000000001 ;
      RECT  188200.0 112000.00000000001 189000.0 112800.00000000001 ;
      RECT  188200.0 112000.00000000001 189000.0 112800.00000000001 ;
      RECT  181400.0 112000.00000000001 182200.0 112800.00000000001 ;
      RECT  188200.0 112000.00000000001 189000.0 112800.00000000001 ;
      RECT  185000.0 95000.00000000001 185800.0 95800.00000000001 ;
      RECT  184000.0 81600.00000000001 184800.0 82400.0 ;
      RECT  191800.0 95000.00000000001 192600.00000000003 95800.00000000001 ;
      RECT  190800.0 81600.00000000001 191600.00000000003 82400.0 ;
      RECT  184100.00000000003 81700.0 184700.0 82300.00000000001 ;
      RECT  190900.0 81700.0 191500.0 82300.00000000001 ;
      RECT  185100.00000000003 95100.00000000001 185700.0 95700.0 ;
      RECT  191900.0 95100.00000000001 192500.0 95700.0 ;
      RECT  182400.0 30400.000000000004 183200.0 31200.000000000004 ;
      RECT  181800.0 47800.00000000001 182600.00000000003 48600.00000000001 ;
      RECT  182400.0 37000.0 183200.0 37800.00000000001 ;
      RECT  183800.0 41400.00000000001 184600.00000000003 42200.0 ;
      RECT  183200.0 54800.00000000001 184000.0 55600.00000000001 ;
      RECT  189200.0 30400.000000000004 190000.0 31200.000000000004 ;
      RECT  188600.00000000003 47800.00000000001 189400.0 48600.00000000001 ;
      RECT  189200.0 37000.0 190000.0 37800.00000000001 ;
      RECT  190600.00000000003 41400.00000000001 191400.0 42200.0 ;
      RECT  190000.0 54800.00000000001 190800.0 55600.00000000001 ;
      RECT  182500.0 30500.000000000004 183100.00000000003 31100.0 ;
      RECT  181900.0 47900.00000000001 182500.0 48500.0 ;
      RECT  189300.0 30500.000000000004 189900.0 31100.0 ;
      RECT  188700.0 47900.00000000001 189300.0 48500.0 ;
      RECT  182500.0 37100.0 183100.00000000003 37700.0 ;
      RECT  183900.0 41500.0 184500.0 42100.00000000001 ;
      RECT  183300.0 54900.00000000001 183900.0 55500.0 ;
      RECT  189300.0 37100.0 189900.0 37700.0 ;
      RECT  190700.0 41500.0 191300.0 42100.00000000001 ;
      RECT  190100.00000000003 54900.00000000001 190700.0 55500.0 ;
      RECT  74199.99999999999 132900.0 81500.0 133500.0 ;
      RECT  75600.0 142100.00000000003 82899.99999999999 142700.0 ;
      RECT  77000.0 169700.0 81500.0 170300.0 ;
      RECT  78400.0 178899.99999999997 82900.0 179500.0 ;
      RECT  111700.0 131500.0 115100.0 132100.00000000003 ;
      RECT  111700.0 141100.00000000003 116500.0 141700.0 ;
      RECT  111700.0 149900.0 117900.0 150500.0 ;
      RECT  111700.0 159500.0 119300.00000000001 160100.00000000003 ;
      RECT  111700.0 168300.0 120700.0 168899.99999999997 ;
      RECT  111700.0 177899.99999999997 122100.0 178500.0 ;
      RECT  111700.0 186700.0 123500.0 187300.0 ;
      RECT  111700.0 196300.0 124900.0 196899.99999999997 ;
      RECT  90500.0 131600.00000000003 89700.0 132400.0 ;
      RECT  108500.0 131600.00000000003 107700.0 132400.0 ;
      RECT  90500.0 122400.0 89700.0 123200.0 ;
      RECT  108500.0 122400.0 107700.0 123200.0 ;
      RECT  90500.0 131600.00000000003 89700.0 132400.0 ;
      RECT  108500.0 131600.00000000003 107700.0 132400.0 ;
      RECT  90500.0 140800.0 89700.0 141600.00000000003 ;
      RECT  108500.0 140800.0 107700.0 141600.00000000003 ;
      RECT  90500.0 150000.0 89700.0 150800.0 ;
      RECT  108500.0 150000.0 107700.0 150800.0 ;
      RECT  90500.0 140800.0 89700.0 141600.00000000003 ;
      RECT  108500.0 140800.0 107700.0 141600.00000000003 ;
      RECT  90500.0 150000.0 89700.0 150800.0 ;
      RECT  108500.0 150000.0 107700.0 150800.0 ;
      RECT  90500.0 159200.0 89700.0 160000.0 ;
      RECT  108500.0 159200.0 107700.0 160000.0 ;
      RECT  89700.0 131600.00000000003 90500.0 132400.0 ;
      RECT  107700.0 131600.00000000003 108500.0 132400.0 ;
      RECT  89700.0 150000.0 90500.0 150800.0 ;
      RECT  107700.0 150000.0 108500.0 150800.0 ;
      RECT  89700.0 122400.0 90500.0 123200.0 ;
      RECT  107700.0 122400.0 108500.0 123200.0 ;
      RECT  89700.0 140800.0 90500.0 141600.00000000003 ;
      RECT  107700.0 140800.0 108500.0 141600.00000000003 ;
      RECT  89700.0 159200.0 90500.0 160000.0 ;
      RECT  107700.0 159200.0 108500.0 160000.0 ;
      RECT  90500.0 168399.99999999997 89700.0 169200.0 ;
      RECT  108500.0 168399.99999999997 107700.0 169200.0 ;
      RECT  90500.0 159200.0 89700.0 160000.0 ;
      RECT  108500.0 159200.0 107700.0 160000.0 ;
      RECT  90500.0 168399.99999999997 89700.0 169200.0 ;
      RECT  108500.0 168399.99999999997 107700.0 169200.0 ;
      RECT  90500.0 177600.00000000003 89700.0 178399.99999999997 ;
      RECT  108500.0 177600.00000000003 107700.0 178399.99999999997 ;
      RECT  90500.0 186800.0 89700.0 187600.00000000003 ;
      RECT  108500.0 186800.0 107700.0 187600.00000000003 ;
      RECT  90500.0 177600.00000000003 89700.0 178399.99999999997 ;
      RECT  108500.0 177600.00000000003 107700.0 178399.99999999997 ;
      RECT  90500.0 186800.0 89700.0 187600.00000000003 ;
      RECT  108500.0 186800.0 107700.0 187600.00000000003 ;
      RECT  90500.0 196000.0 89700.0 196800.0 ;
      RECT  108500.0 196000.0 107700.0 196800.0 ;
      RECT  89700.0 168399.99999999997 90500.0 169200.0 ;
      RECT  107700.0 168399.99999999997 108500.0 169200.0 ;
      RECT  89700.0 186800.0 90500.0 187600.00000000003 ;
      RECT  107700.0 186800.0 108500.0 187600.00000000003 ;
      RECT  89700.0 159200.0 90500.0 160000.0 ;
      RECT  107700.0 159200.0 108500.0 160000.0 ;
      RECT  89700.0 177600.00000000003 90500.0 178399.99999999997 ;
      RECT  107700.0 177600.00000000003 108500.0 178399.99999999997 ;
      RECT  89700.0 196000.0 90500.0 196800.0 ;
      RECT  107700.0 196000.0 108500.0 196800.0 ;
      RECT  81900.0 132800.0 81100.0 133600.00000000003 ;
      RECT  74600.0 132800.0 73800.0 133600.00000000003 ;
      RECT  83300.0 142000.0 82500.0 142800.0 ;
      RECT  76000.0 142000.0 75200.0 142800.0 ;
      RECT  81900.0 169600.00000000003 81100.0 170399.99999999997 ;
      RECT  77400.0 169600.00000000003 76600.0 170399.99999999997 ;
      RECT  83300.0 178800.0 82500.0 179600.00000000003 ;
      RECT  78800.0 178800.0 78000.0 179600.00000000003 ;
      RECT  112100.0 131400.0 111300.00000000001 132200.0 ;
      RECT  115500.0 131400.0 114700.0 132200.0 ;
      RECT  112100.0 141000.0 111300.00000000001 141800.0 ;
      RECT  116900.0 141000.0 116100.0 141800.0 ;
      RECT  112100.0 149800.0 111300.00000000001 150600.00000000003 ;
      RECT  118300.0 149800.0 117500.0 150600.00000000003 ;
      RECT  112100.0 159399.99999999997 111300.00000000001 160200.0 ;
      RECT  119700.0 159399.99999999997 118900.0 160200.0 ;
      RECT  112100.0 168200.0 111300.00000000001 169000.0 ;
      RECT  121100.0 168200.0 120300.00000000001 169000.0 ;
      RECT  112100.0 177800.0 111300.00000000001 178600.00000000003 ;
      RECT  122500.0 177800.0 121700.0 178600.00000000003 ;
      RECT  112100.0 186600.00000000003 111300.00000000001 187399.99999999997 ;
      RECT  123900.0 186600.00000000003 123100.0 187399.99999999997 ;
      RECT  112100.0 196200.0 111300.00000000001 197000.0 ;
      RECT  125300.0 196200.0 124500.0 197000.0 ;
      RECT  130900.0 131600.00000000003 130100.00000000003 132400.0 ;
      RECT  130900.0 122400.0 130100.00000000003 123200.0 ;
      RECT  130900.0 131600.00000000003 130100.00000000003 132400.0 ;
      RECT  130900.0 140800.0 130100.00000000003 141600.00000000003 ;
      RECT  130900.0 150000.0 130100.00000000003 150800.0 ;
      RECT  130900.0 140800.0 130100.00000000003 141600.00000000003 ;
      RECT  130900.0 150000.0 130100.00000000003 150800.0 ;
      RECT  130900.0 159200.0 130100.00000000003 160000.0 ;
      RECT  130900.0 168399.99999999997 130100.00000000003 169200.0 ;
      RECT  130900.0 159200.0 130100.00000000003 160000.0 ;
      RECT  130900.0 168399.99999999997 130100.00000000003 169200.0 ;
      RECT  130900.0 177600.00000000003 130100.00000000003 178399.99999999997 ;
      RECT  130900.0 186800.0 130100.00000000003 187600.00000000003 ;
      RECT  130900.0 177600.00000000003 130100.00000000003 178399.99999999997 ;
      RECT  130900.0 186800.0 130100.00000000003 187600.00000000003 ;
      RECT  130900.0 196000.0 130100.00000000003 196800.0 ;
      RECT  130900.0 205200.0 130100.00000000003 206000.0 ;
      RECT  130900.0 196000.0 130100.00000000003 196800.0 ;
      RECT  130900.0 205200.0 130100.00000000003 206000.0 ;
      RECT  130900.0 214400.00000000003 130100.00000000003 215200.0 ;
      RECT  130900.0 223600.00000000003 130100.00000000003 224400.00000000003 ;
      RECT  130900.0 214400.00000000003 130100.00000000003 215200.0 ;
      RECT  130900.0 223600.00000000003 130100.00000000003 224400.00000000003 ;
      RECT  130900.0 232800.0 130100.00000000003 233600.00000000003 ;
      RECT  130900.0 242000.0 130100.00000000003 242800.0 ;
      RECT  130900.0 232800.0 130100.00000000003 233600.00000000003 ;
      RECT  130900.0 242000.0 130100.00000000003 242800.0 ;
      RECT  130900.0 251200.0 130100.00000000003 252000.0 ;
      RECT  130900.0 260399.99999999997 130100.00000000003 261200.0 ;
      RECT  130900.0 251200.0 130100.00000000003 252000.0 ;
      RECT  130900.0 260399.99999999997 130100.00000000003 261200.0 ;
      RECT  130900.0 269600.0 130100.00000000003 270400.00000000006 ;
      RECT  130100.0 131600.00000000003 130900.0 132400.0 ;
      RECT  130100.0 150000.0 130900.0 150800.0 ;
      RECT  130100.0 168399.99999999997 130900.0 169200.0 ;
      RECT  130100.0 186800.0 130900.0 187600.00000000003 ;
      RECT  130100.0 205200.0 130900.0 206000.0 ;
      RECT  130100.0 223600.00000000003 130900.0 224400.00000000003 ;
      RECT  130100.0 242000.0 130900.0 242800.0 ;
      RECT  130100.0 260399.99999999997 130900.0 261200.0 ;
      RECT  89700.0 131600.00000000003 90500.0 132400.0 ;
      RECT  107700.0 131600.00000000003 108500.0 132400.0 ;
      RECT  89700.0 150000.0 90500.0 150800.0 ;
      RECT  107700.0 150000.0 108500.0 150800.0 ;
      RECT  89700.0 168399.99999999997 90500.0 169200.0 ;
      RECT  107700.0 168399.99999999997 108500.0 169200.0 ;
      RECT  89700.0 186800.0 90500.0 187600.00000000003 ;
      RECT  107700.0 186800.0 108500.0 187600.00000000003 ;
      RECT  130100.0 122400.0 130900.0 123200.0 ;
      RECT  130100.0 140800.0 130900.0 141600.00000000003 ;
      RECT  130100.0 159200.0 130900.0 160000.0 ;
      RECT  130100.0 177600.00000000003 130900.0 178399.99999999997 ;
      RECT  130100.0 196000.0 130900.0 196800.0 ;
      RECT  130100.0 214400.00000000003 130900.0 215200.0 ;
      RECT  130100.0 232800.0 130900.0 233600.00000000003 ;
      RECT  130100.0 251200.0 130900.0 252000.0 ;
      RECT  130100.0 269600.0 130900.0 270400.0 ;
      RECT  89700.0 122400.0 90500.0 123200.0 ;
      RECT  107700.0 122400.0 108500.0 123200.0 ;
      RECT  89700.0 140800.0 90500.0 141600.00000000003 ;
      RECT  107700.0 140800.0 108500.0 141600.00000000003 ;
      RECT  89700.0 159200.0 90500.0 160000.0 ;
      RECT  107700.0 159200.0 108500.0 160000.0 ;
      RECT  89700.0 177600.00000000003 90500.0 178399.99999999997 ;
      RECT  107700.0 177600.00000000003 108500.0 178399.99999999997 ;
      RECT  89700.0 196000.0 90500.0 196800.0 ;
      RECT  107700.0 196000.0 108500.0 196800.0 ;
      RECT  155100.0 131600.00000000003 154300.0 132400.0 ;
      RECT  164700.0 131600.00000000003 163899.99999999997 132400.0 ;
      RECT  155100.0 122400.0 154300.0 123200.0 ;
      RECT  164700.0 122400.0 163899.99999999997 123200.0 ;
      RECT  155100.0 131600.00000000003 154300.0 132400.0 ;
      RECT  164700.0 131600.00000000003 163899.99999999997 132400.0 ;
      RECT  155100.0 140800.0 154300.0 141600.00000000003 ;
      RECT  164700.0 140800.0 163899.99999999997 141600.00000000003 ;
      RECT  155100.0 150000.0 154300.0 150800.0 ;
      RECT  164700.0 150000.0 163899.99999999997 150800.0 ;
      RECT  155100.0 140800.0 154300.0 141600.00000000003 ;
      RECT  164700.0 140800.0 163899.99999999997 141600.00000000003 ;
      RECT  155100.0 150000.0 154300.0 150800.0 ;
      RECT  164700.0 150000.0 163899.99999999997 150800.0 ;
      RECT  155100.0 159200.0 154300.0 160000.0 ;
      RECT  164700.0 159200.0 163899.99999999997 160000.0 ;
      RECT  155100.0 168399.99999999997 154300.0 169200.0 ;
      RECT  164700.0 168399.99999999997 163899.99999999997 169200.0 ;
      RECT  155100.0 159200.0 154300.0 160000.0 ;
      RECT  164700.0 159200.0 163899.99999999997 160000.0 ;
      RECT  155100.0 168399.99999999997 154300.0 169200.0 ;
      RECT  164700.0 168399.99999999997 163899.99999999997 169200.0 ;
      RECT  155100.0 177600.00000000003 154300.0 178399.99999999997 ;
      RECT  164700.0 177600.00000000003 163899.99999999997 178399.99999999997 ;
      RECT  155100.0 186800.0 154300.0 187600.00000000003 ;
      RECT  164700.0 186800.0 163899.99999999997 187600.00000000003 ;
      RECT  155100.0 177600.00000000003 154300.0 178399.99999999997 ;
      RECT  164700.0 177600.00000000003 163899.99999999997 178399.99999999997 ;
      RECT  155100.0 186800.0 154300.0 187600.00000000003 ;
      RECT  164700.0 186800.0 163899.99999999997 187600.00000000003 ;
      RECT  155100.0 196000.0 154300.0 196800.0 ;
      RECT  164700.0 196000.0 163899.99999999997 196800.0 ;
      RECT  155100.0 205200.0 154300.0 206000.0 ;
      RECT  164700.0 205200.0 163899.99999999997 206000.0 ;
      RECT  155100.0 196000.0 154300.0 196800.0 ;
      RECT  164700.0 196000.0 163899.99999999997 196800.0 ;
      RECT  155100.0 205200.0 154300.0 206000.0 ;
      RECT  164700.0 205200.0 163899.99999999997 206000.0 ;
      RECT  155100.0 214400.00000000003 154300.0 215200.0 ;
      RECT  164700.0 214400.00000000003 163899.99999999997 215200.0 ;
      RECT  155100.0 223600.00000000003 154300.0 224400.00000000003 ;
      RECT  164700.0 223600.00000000003 163899.99999999997 224400.00000000003 ;
      RECT  155100.0 214400.00000000003 154300.0 215200.0 ;
      RECT  164700.0 214400.00000000003 163899.99999999997 215200.0 ;
      RECT  155100.0 223600.00000000003 154300.0 224400.00000000003 ;
      RECT  164700.0 223600.00000000003 163899.99999999997 224400.00000000003 ;
      RECT  155100.0 232800.0 154300.0 233600.00000000003 ;
      RECT  164700.0 232800.0 163899.99999999997 233600.00000000003 ;
      RECT  155100.0 242000.0 154300.0 242800.0 ;
      RECT  164700.0 242000.0 163899.99999999997 242800.0 ;
      RECT  155100.0 232800.0 154300.0 233600.00000000003 ;
      RECT  164700.0 232800.0 163899.99999999997 233600.00000000003 ;
      RECT  155100.0 242000.0 154300.0 242800.0 ;
      RECT  164700.0 242000.0 163899.99999999997 242800.0 ;
      RECT  155100.0 251200.0 154300.0 252000.0 ;
      RECT  164700.0 251200.0 163899.99999999997 252000.0 ;
      RECT  155100.0 260399.99999999997 154300.0 261200.0 ;
      RECT  164700.0 260399.99999999997 163899.99999999997 261200.0 ;
      RECT  155100.0 251200.0 154300.0 252000.0 ;
      RECT  164700.0 251200.0 163899.99999999997 252000.0 ;
      RECT  155100.0 260399.99999999997 154300.0 261200.0 ;
      RECT  164700.0 260399.99999999997 163899.99999999997 261200.0 ;
      RECT  155100.0 269600.0 154300.0 270400.00000000006 ;
      RECT  164700.0 269600.0 163899.99999999997 270400.00000000006 ;
      RECT  154399.99999999997 131700.0 155000.0 132300.0 ;
      RECT  164000.0 131700.0 164600.0 132300.0 ;
      RECT  154399.99999999997 150100.00000000003 155000.0 150700.0 ;
      RECT  164000.0 150100.00000000003 164600.0 150700.0 ;
      RECT  154399.99999999997 168500.0 155000.0 169100.00000000003 ;
      RECT  164000.0 168500.0 164600.0 169100.00000000003 ;
      RECT  154399.99999999997 186900.00000000003 155000.0 187500.0 ;
      RECT  164000.0 186900.00000000003 164600.0 187500.0 ;
      RECT  154399.99999999997 205300.0 155000.0 205900.00000000003 ;
      RECT  164000.0 205300.0 164600.0 205900.00000000003 ;
      RECT  154399.99999999997 223700.0 155000.0 224300.0 ;
      RECT  164000.0 223700.0 164600.0 224300.0 ;
      RECT  154399.99999999997 242100.00000000003 155000.0 242700.0 ;
      RECT  164000.0 242100.00000000003 164600.0 242700.0 ;
      RECT  154399.99999999997 260500.0 155000.0 261100.00000000003 ;
      RECT  164000.0 260500.0 164600.0 261100.00000000003 ;
      RECT  154399.99999999997 122500.0 155000.0 123100.00000000001 ;
      RECT  164000.0 122500.0 164600.0 123100.00000000001 ;
      RECT  154399.99999999997 140900.0 155000.0 141500.0 ;
      RECT  164000.0 140900.0 164600.0 141500.0 ;
      RECT  154399.99999999997 159300.0 155000.0 159899.99999999997 ;
      RECT  164000.0 159300.0 164600.0 159899.99999999997 ;
      RECT  154399.99999999997 177700.0 155000.0 178300.0 ;
      RECT  164000.0 177700.0 164600.0 178300.0 ;
      RECT  154399.99999999997 196100.00000000003 155000.0 196700.0 ;
      RECT  164000.0 196100.00000000003 164600.0 196700.0 ;
      RECT  154399.99999999997 214500.0 155000.0 215100.00000000003 ;
      RECT  164000.0 214500.0 164600.0 215100.00000000003 ;
      RECT  154399.99999999997 232900.00000000003 155000.0 233500.0 ;
      RECT  164000.0 232900.00000000003 164600.0 233500.0 ;
      RECT  154399.99999999997 251300.0 155000.0 251899.99999999997 ;
      RECT  164000.0 251300.0 164600.0 251899.99999999997 ;
      RECT  154399.99999999997 269700.0 155000.0 270300.0 ;
      RECT  164000.0 269700.0 164600.0 270300.0 ;
      RECT  181700.0 131300.0 182300.0 131900.0 ;
      RECT  188500.0 131300.0 189100.00000000003 131900.0 ;
      RECT  181700.0 149700.0 182300.0 150300.0 ;
      RECT  188500.0 149700.0 189100.00000000003 150300.0 ;
      RECT  181700.0 168100.00000000003 182300.0 168700.0 ;
      RECT  188500.0 168100.00000000003 189100.00000000003 168700.0 ;
      RECT  181700.0 186500.0 182300.0 187100.00000000003 ;
      RECT  188500.0 186500.0 189100.00000000003 187100.00000000003 ;
      RECT  181700.0 204899.99999999997 182300.0 205500.0 ;
      RECT  188500.0 204899.99999999997 189100.00000000003 205500.0 ;
      RECT  181700.0 223300.0 182300.0 223899.99999999997 ;
      RECT  188500.0 223300.0 189100.00000000003 223899.99999999997 ;
      RECT  181700.0 241700.0 182300.0 242300.0 ;
      RECT  188500.0 241700.0 189100.00000000003 242300.0 ;
      RECT  181700.0 260100.00000000003 182300.0 260700.0 ;
      RECT  188500.0 260100.00000000003 189100.00000000003 260700.0 ;
      RECT  181400.0 112000.0 182200.0 112800.0 ;
      RECT  188200.0 112000.0 189000.0 112800.0 ;
      RECT  184100.00000000003 81700.0 184700.0 82300.00000000001 ;
      RECT  190900.0 81700.0 191500.0 82300.00000000001 ;
      RECT  182500.0 30500.0 183100.00000000003 31099.999999999993 ;
      RECT  181900.0 47900.00000000001 182500.0 48500.0 ;
      RECT  189300.0 30500.0 189900.0 31099.999999999993 ;
      RECT  188700.0 47900.00000000001 189300.0 48500.0 ;
      RECT  130100.00000000003 131600.00000000003 130900.0 132400.0 ;
      RECT  130100.00000000003 150000.0 130900.0 150800.0 ;
      RECT  130100.00000000003 168399.99999999997 130900.0 169200.0 ;
      RECT  130100.00000000003 186800.0 130900.0 187600.00000000003 ;
      RECT  130100.00000000003 205200.0 130900.0 206000.0 ;
      RECT  130100.00000000003 223600.00000000003 130900.0 224399.99999999997 ;
      RECT  130100.00000000003 242000.0 130900.0 242800.0 ;
      RECT  130100.00000000003 260399.99999999997 130900.0 261200.0 ;
      RECT  89700.0 131600.00000000003 90500.0 132400.0 ;
      RECT  107700.0 131600.00000000003 108500.0 132400.0 ;
      RECT  89700.0 150000.0 90500.0 150800.0 ;
      RECT  107700.0 150000.0 108500.0 150800.0 ;
      RECT  89700.0 168399.99999999997 90500.0 169200.0 ;
      RECT  107700.0 168399.99999999997 108500.0 169200.0 ;
      RECT  89700.0 186800.0 90500.0 187600.00000000003 ;
      RECT  107700.0 186800.0 108500.0 187600.00000000003 ;
      RECT  154400.0 131700.0 155000.0 132300.0 ;
      RECT  164000.0 131700.0 164600.00000000003 132300.0 ;
      RECT  154400.0 150100.00000000003 155000.0 150700.0 ;
      RECT  164000.0 150100.00000000003 164600.00000000003 150700.0 ;
      RECT  154400.0 168500.0 155000.0 169100.00000000003 ;
      RECT  164000.0 168500.0 164600.00000000003 169100.00000000003 ;
      RECT  154400.0 186899.99999999997 155000.0 187500.0 ;
      RECT  164000.0 186899.99999999997 164600.00000000003 187500.0 ;
      RECT  154400.0 205300.0 155000.0 205899.99999999997 ;
      RECT  164000.0 205300.0 164600.00000000003 205899.99999999997 ;
      RECT  154400.0 223700.0 155000.0 224300.0 ;
      RECT  164000.0 223700.0 164600.00000000003 224300.0 ;
      RECT  154400.0 242100.00000000003 155000.0 242700.0 ;
      RECT  164000.0 242100.00000000003 164600.00000000003 242700.0 ;
      RECT  154400.0 260500.0 155000.0 261100.00000000003 ;
      RECT  164000.0 260500.0 164600.00000000003 261100.00000000003 ;
      RECT  178300.0 126700.0 178900.0 127300.00000000001 ;
      RECT  185100.00000000003 126700.0 185700.0 127300.00000000001 ;
      RECT  191900.0 126700.0 192500.0 127300.00000000001 ;
      RECT  178300.0 135900.0 178900.0 136500.0 ;
      RECT  185100.00000000003 135900.0 185700.0 136500.0 ;
      RECT  191900.0 135900.0 192500.0 136500.0 ;
      RECT  178300.0 145100.00000000003 178900.0 145700.0 ;
      RECT  185100.00000000003 145100.00000000003 185700.0 145700.0 ;
      RECT  191900.0 145100.00000000003 192500.0 145700.0 ;
      RECT  178300.0 154300.0 178900.0 154899.99999999997 ;
      RECT  185100.00000000003 154300.0 185700.0 154899.99999999997 ;
      RECT  191900.0 154300.0 192500.0 154899.99999999997 ;
      RECT  178300.0 163500.0 178900.0 164100.00000000003 ;
      RECT  185100.00000000003 163500.0 185700.0 164100.00000000003 ;
      RECT  191900.0 163500.0 192500.0 164100.00000000003 ;
      RECT  178300.0 172700.0 178900.0 173300.0 ;
      RECT  185100.00000000003 172700.0 185700.0 173300.0 ;
      RECT  191900.0 172700.0 192500.0 173300.0 ;
      RECT  178300.0 181899.99999999997 178900.0 182500.0 ;
      RECT  185100.00000000003 181899.99999999997 185700.0 182500.0 ;
      RECT  191900.0 181899.99999999997 192500.0 182500.0 ;
      RECT  178300.0 191100.00000000003 178900.0 191700.0 ;
      RECT  185100.00000000003 191100.00000000003 185700.0 191700.0 ;
      RECT  191900.0 191100.00000000003 192500.0 191700.0 ;
      RECT  178300.0 200300.0 178900.0 200899.99999999997 ;
      RECT  185100.00000000003 200300.0 185700.0 200899.99999999997 ;
      RECT  191900.0 200300.0 192500.0 200899.99999999997 ;
      RECT  178300.0 209500.0 178900.0 210100.00000000003 ;
      RECT  185100.00000000003 209500.0 185700.0 210100.00000000003 ;
      RECT  191900.0 209500.0 192500.0 210100.00000000003 ;
      RECT  178300.0 218700.0 178900.0 219300.0 ;
      RECT  185100.00000000003 218700.0 185700.0 219300.0 ;
      RECT  191900.0 218700.0 192500.0 219300.0 ;
      RECT  178300.0 227899.99999999997 178900.0 228500.0 ;
      RECT  185100.00000000003 227899.99999999997 185700.0 228500.0 ;
      RECT  191900.0 227899.99999999997 192500.0 228500.0 ;
      RECT  178300.0 237100.00000000003 178900.0 237700.0 ;
      RECT  185100.00000000003 237100.00000000003 185700.0 237700.0 ;
      RECT  191900.0 237100.00000000003 192500.0 237700.0 ;
      RECT  178300.0 246300.0 178900.0 246899.99999999997 ;
      RECT  185100.00000000003 246300.0 185700.0 246899.99999999997 ;
      RECT  191900.0 246300.0 192500.0 246899.99999999997 ;
      RECT  178300.0 255500.0 178900.0 256100.00000000003 ;
      RECT  185100.00000000003 255500.0 185700.0 256100.00000000003 ;
      RECT  191900.0 255500.0 192500.0 256100.00000000003 ;
      RECT  178300.0 264700.0 178900.0 265300.0 ;
      RECT  185100.00000000003 264700.0 185700.0 265300.0 ;
      RECT  191900.0 264700.0 192500.0 265300.0 ;
      RECT  185100.00000000003 95100.00000000001 185700.0 95700.0 ;
      RECT  191900.0 95100.00000000001 192500.0 95700.0 ;
      RECT  182500.0 37099.99999999999 183100.00000000003 37700.0 ;
      RECT  183900.0 41500.0 184500.0 42099.99999999999 ;
      RECT  183300.0 54900.00000000001 183900.0 55500.0 ;
      RECT  189300.0 37099.99999999999 189900.0 37700.0 ;
      RECT  190700.0 41500.0 191300.0 42099.99999999999 ;
      RECT  190100.00000000003 54900.00000000001 190700.0 55500.0 ;
      RECT  130100.00000000003 122400.0 130900.0 123200.0 ;
      RECT  130100.00000000003 140800.0 130900.0 141600.00000000003 ;
      RECT  130100.00000000003 159200.0 130900.0 160000.0 ;
      RECT  130100.00000000003 177600.00000000003 130900.0 178399.99999999997 ;
      RECT  130100.00000000003 196000.0 130900.0 196800.0 ;
      RECT  130100.00000000003 214399.99999999997 130900.0 215200.0 ;
      RECT  130100.00000000003 232800.0 130900.0 233600.00000000003 ;
      RECT  130100.00000000003 251200.0 130900.0 252000.0 ;
      RECT  130100.00000000003 269600.0 130900.0 270400.0 ;
      RECT  89700.0 122400.0 90500.0 123200.0 ;
      RECT  107700.0 122400.0 108500.0 123200.0 ;
      RECT  89700.0 140800.0 90500.0 141600.00000000003 ;
      RECT  107700.0 140800.0 108500.0 141600.00000000003 ;
      RECT  89700.0 159200.0 90500.0 160000.0 ;
      RECT  107700.0 159200.0 108500.0 160000.0 ;
      RECT  89700.0 177600.00000000003 90500.0 178399.99999999997 ;
      RECT  107700.0 177600.00000000003 108500.0 178399.99999999997 ;
      RECT  89700.0 196000.0 90500.0 196800.0 ;
      RECT  107700.0 196000.0 108500.0 196800.0 ;
      RECT  154400.0 122500.0 155000.0 123100.00000000001 ;
      RECT  164000.0 122500.0 164600.00000000003 123100.00000000001 ;
      RECT  154400.0 140900.0 155000.0 141500.0 ;
      RECT  164000.0 140900.0 164600.00000000003 141500.0 ;
      RECT  154400.0 159300.0 155000.0 159899.99999999997 ;
      RECT  164000.0 159300.0 164600.00000000003 159899.99999999997 ;
      RECT  154400.0 177700.0 155000.0 178300.0 ;
      RECT  164000.0 177700.0 164600.00000000003 178300.0 ;
      RECT  154400.0 196100.00000000003 155000.0 196700.0 ;
      RECT  164000.0 196100.00000000003 164600.00000000003 196700.0 ;
      RECT  154400.0 214500.0 155000.0 215100.00000000003 ;
      RECT  164000.0 214500.0 164600.00000000003 215100.00000000003 ;
      RECT  154400.0 232899.99999999997 155000.0 233500.0 ;
      RECT  164000.0 232899.99999999997 164600.00000000003 233500.0 ;
      RECT  154400.0 251300.0 155000.0 251899.99999999997 ;
      RECT  164000.0 251300.0 164600.00000000003 251899.99999999997 ;
      RECT  154400.0 269700.0 155000.0 270300.0 ;
      RECT  164000.0 269700.0 164600.00000000003 270300.0 ;
      RECT  1900.0000000000002 89500.0 48400.0 90100.0 ;
      RECT  28500.0 50100.0 51600.0 50700.0 ;
      RECT  29900.000000000004 28500.0 51600.00000000001 29100.0 ;
      RECT  21200.000000000004 29100.0 21800.000000000004 29700.000000000004 ;
      RECT  21200.000000000004 28900.000000000004 21800.000000000004 29500.0 ;
      RECT  19200.000000000004 29100.0 21500.000000000004 29700.000000000004 ;
      RECT  21200.000000000004 29200.000000000004 21800.000000000004 29400.000000000004 ;
      RECT  21500.0 28900.000000000004 23800.0 29500.0 ;
      RECT  18800.0 29000.0 19600.0 29800.000000000004 ;
      RECT  23400.000000000004 28800.000000000004 24200.000000000004 29600.0 ;
      RECT  21200.000000000004 50100.0 21800.000000000004 49500.0 ;
      RECT  21200.000000000004 50300.0 21800.000000000004 49700.0 ;
      RECT  19200.000000000004 50100.0 21500.000000000004 49500.0 ;
      RECT  21200.000000000004 50000.0 21800.000000000004 49800.0 ;
      RECT  21500.0 50300.0 23800.0 49700.0 ;
      RECT  18800.0 50200.0 19600.0 49400.0 ;
      RECT  23400.000000000004 50400.0 24200.000000000004 49600.0 ;
      RECT  400.0 39200.0 -400.0 40000.0 ;
      RECT  400.0 19200.000000000004 -400.0 20000.0 ;
      RECT  400.0 39200.0 -400.0 40000.0 ;
      RECT  400.0 59200.0 -400.0 60000.0 ;
      RECT  -400.0 39200.0 400.0 40000.0 ;
      RECT  -400.0 19200.000000000004 400.0 20000.0 ;
      RECT  -400.0 59200.0 400.0 60000.00000000001 ;
      RECT  3600.0 137800.0 21200.000000000004 138400.0 ;
      RECT  3600.0 147400.0 21200.000000000004 148000.0 ;
      RECT  3600.0 156200.00000000003 21200.000000000004 156800.0 ;
      RECT  3600.0 165800.0 21200.000000000004 166400.0 ;
      RECT  8000.0 137700.00000000003 8800.0 138500.0 ;
      RECT  14400.0 137700.00000000003 15200.000000000002 138500.0 ;
      RECT  20800.0 137700.00000000003 21600.0 138500.0 ;
      RECT  3200.0 137700.00000000003 4000.0 138500.0 ;
      RECT  8000.0 147300.0 8800.0 148100.0 ;
      RECT  14400.0 147300.0 15200.000000000002 148100.0 ;
      RECT  20800.0 147300.0 21600.0 148100.0 ;
      RECT  3200.0 147300.0 4000.0 148100.0 ;
      RECT  8000.0 156100.0 8800.0 156900.0 ;
      RECT  14400.0 156100.0 15200.000000000002 156900.0 ;
      RECT  20800.0 156100.0 21600.0 156900.0 ;
      RECT  3200.0 156100.0 4000.0 156900.0 ;
      RECT  8000.0 165700.00000000003 8800.0 166500.0 ;
      RECT  14400.0 165700.00000000003 15200.000000000002 166500.0 ;
      RECT  20800.0 165700.00000000003 21600.0 166500.0 ;
      RECT  3200.0 165700.00000000003 4000.0 166500.0 ;
      RECT  13200.000000000002 142500.0 12400.0 143300.0 ;
      RECT  13200.000000000002 133300.0 12400.0 134100.00000000003 ;
      RECT  19600.0 142500.0 18800.0 143300.0 ;
      RECT  19600.0 133300.0 18800.0 134100.00000000003 ;
      RECT  13200.000000000002 160900.0 12400.0 161700.00000000003 ;
      RECT  13200.000000000002 151700.00000000003 12400.0 152500.0 ;
      RECT  19600.0 160900.0 18800.0 161700.00000000003 ;
      RECT  19600.0 151700.00000000003 18800.0 152500.0 ;
      RECT  13200.000000000002 170100.0 12400.0 170900.0 ;
      RECT  19600.0 170100.0 18800.0 170900.0 ;
      RECT  12400.0 142500.0 13200.000000000002 143300.0 ;
      RECT  18800.0 142500.0 19600.0 143300.0 ;
      RECT  12400.0 160900.0 13200.000000000002 161700.00000000003 ;
      RECT  18800.0 160900.0 19600.0 161700.00000000003 ;
      RECT  12400.0 133300.0 13200.000000000002 134100.00000000003 ;
      RECT  18800.0 133300.0 19600.0 134100.00000000003 ;
      RECT  12400.0 151700.00000000003 13200.000000000002 152500.0 ;
      RECT  18800.0 151700.00000000003 19600.0 152500.0 ;
      RECT  12400.0 170100.0 13200.000000000002 170900.0 ;
      RECT  18800.0 170100.0 19600.0 170900.0 ;
      RECT  31400.000000000004 142500.0 32200.000000000004 143300.0 ;
      RECT  31400.000000000004 142500.0 32200.000000000004 143300.0 ;
      RECT  31400.000000000004 160900.0 32200.000000000004 161700.00000000003 ;
      RECT  31400.000000000004 160900.0 32200.000000000004 161700.00000000003 ;
      RECT  31400.000000000004 179300.0 32200.000000000004 180100.0 ;
      RECT  31400.000000000004 179300.0 32200.000000000004 180100.0 ;
      RECT  31400.000000000004 197700.00000000003 32200.000000000004 198500.0 ;
      RECT  31400.000000000004 197700.00000000003 32200.000000000004 198500.0 ;
      RECT  28000.000000000004 137900.0 28800.0 138700.00000000003 ;
      RECT  34800.00000000001 137900.0 35600.0 138700.00000000003 ;
      RECT  28000.000000000004 147100.00000000003 28800.0 147900.0 ;
      RECT  34800.00000000001 147100.00000000003 35600.0 147900.0 ;
      RECT  28000.000000000004 156300.0 28800.0 157100.0 ;
      RECT  34800.00000000001 156300.0 35600.0 157100.0 ;
      RECT  28000.000000000004 165500.0 28800.0 166300.0 ;
      RECT  34800.00000000001 165500.0 35600.0 166300.0 ;
      RECT  28000.000000000004 174700.00000000003 28800.0 175500.0 ;
      RECT  34800.00000000001 174700.00000000003 35600.0 175500.0 ;
      RECT  28000.000000000004 183900.0 28800.0 184700.00000000003 ;
      RECT  34800.00000000001 183900.0 35600.0 184700.00000000003 ;
      RECT  28000.000000000004 193100.0 28800.0 193900.0 ;
      RECT  34800.00000000001 193100.0 35600.0 193900.0 ;
      RECT  28000.000000000004 202300.0 28800.0 203100.0 ;
      RECT  34800.00000000001 202300.0 35600.0 203100.0 ;
      RECT  31500.000000000004 142600.00000000003 32100.0 143200.00000000003 ;
      RECT  31500.000000000004 161000.0 32100.0 161600.0 ;
      RECT  31500.000000000004 179400.0 32100.0 180000.00000000003 ;
      RECT  31500.000000000004 197800.0 32100.0 198400.0 ;
      RECT  28100.0 138000.0 28700.000000000004 138600.00000000003 ;
      RECT  34900.00000000001 138000.0 35500.0 138600.00000000003 ;
      RECT  28100.0 147200.00000000003 28700.000000000004 147800.0 ;
      RECT  34900.00000000001 147200.00000000003 35500.0 147800.0 ;
      RECT  28100.0 156400.0 28700.000000000004 157000.0 ;
      RECT  34900.00000000001 156400.0 35500.0 157000.0 ;
      RECT  28100.0 165600.0 28700.000000000004 166200.00000000003 ;
      RECT  34900.00000000001 165600.0 35500.0 166200.00000000003 ;
      RECT  28100.0 174800.0 28700.000000000004 175400.0 ;
      RECT  34900.00000000001 174800.0 35500.0 175400.0 ;
      RECT  28100.0 184000.00000000003 28700.000000000004 184600.0 ;
      RECT  34900.00000000001 184000.00000000003 35500.0 184600.0 ;
      RECT  28100.0 193200.00000000003 28700.000000000004 193800.0 ;
      RECT  34900.00000000001 193200.00000000003 35500.0 193800.0 ;
      RECT  28100.0 202400.0 28700.000000000004 203000.0 ;
      RECT  34900.00000000001 202400.0 35500.0 203000.0 ;
      RECT  6800.000000000001 124100.00000000003 6000.000000000001 124900.0 ;
      RECT  31400.000000000004 122700.00000000001 32200.000000000004 123500.0 ;
      RECT  28800.0 128700.00000000001 28000.0 129500.0 ;
      RECT  35600.0 128700.00000000001 34800.00000000001 129500.0 ;
      RECT  37200.0 134700.00000000003 36400.00000000001 135500.0 ;
      RECT  37200.0 150300.0 36400.00000000001 151100.0 ;
      RECT  37200.0 153100.0 36400.00000000001 153900.0 ;
      RECT  37200.0 168700.00000000003 36400.00000000001 169500.0 ;
      RECT  37200.0 171500.0 36400.00000000001 172300.0 ;
      RECT  37200.0 187100.0 36400.00000000001 187900.0 ;
      RECT  37200.0 189900.0 36400.00000000001 190700.00000000003 ;
      RECT  37200.0 205500.0 36400.00000000001 206299.99999999997 ;
      RECT  17200.000000000004 129100.00000000003 18000.000000000004 129900.0 ;
      RECT  31500.000000000004 142600.00000000003 32100.0 143200.00000000003 ;
      RECT  31500.000000000004 161000.0 32100.0 161600.0 ;
      RECT  31500.000000000004 179400.0 32100.0 180000.0 ;
      RECT  31500.000000000004 197799.99999999997 32100.0 198400.0 ;
      RECT  12400.000000000002 142500.0 13200.000000000002 143300.0 ;
      RECT  18800.0 142500.0 19600.0 143300.0 ;
      RECT  12400.000000000002 160900.0 13200.000000000002 161700.00000000003 ;
      RECT  18800.0 160900.0 19600.0 161700.00000000003 ;
      RECT  6000.0 124100.00000000003 6800.000000000001 124900.0 ;
      RECT  31400.000000000004 122700.00000000001 32200.000000000004 123500.0 ;
      RECT  17200.000000000004 129100.00000000003 18000.0 129900.0 ;
      RECT  28100.0 138000.0 28700.000000000004 138600.00000000003 ;
      RECT  34900.00000000001 138000.0 35500.0 138600.00000000003 ;
      RECT  28100.0 147200.00000000003 28700.000000000004 147800.0 ;
      RECT  34900.00000000001 147200.00000000003 35500.0 147800.0 ;
      RECT  28100.0 156400.0 28700.000000000004 157000.0 ;
      RECT  34900.00000000001 156400.0 35500.0 157000.0 ;
      RECT  28100.0 165600.0 28700.000000000004 166200.00000000003 ;
      RECT  34900.00000000001 165600.0 35500.0 166200.00000000003 ;
      RECT  28100.0 174800.0 28700.000000000004 175400.0 ;
      RECT  34900.00000000001 174800.0 35500.0 175400.0 ;
      RECT  28100.0 184000.0 28700.000000000004 184600.0 ;
      RECT  34900.00000000001 184000.0 35500.0 184600.0 ;
      RECT  28100.0 193200.00000000003 28700.000000000004 193799.99999999997 ;
      RECT  34900.00000000001 193200.00000000003 35500.0 193799.99999999997 ;
      RECT  28100.0 202400.0 28700.000000000004 203000.0 ;
      RECT  34900.00000000001 202400.0 35500.0 203000.0 ;
      RECT  12400.000000000002 133300.0 13200.000000000002 134100.00000000003 ;
      RECT  18800.0 133300.0 19600.0 134100.00000000003 ;
      RECT  12400.000000000002 151700.00000000003 13200.000000000002 152500.0 ;
      RECT  18800.0 151700.00000000003 19600.0 152500.0 ;
      RECT  12400.000000000002 170100.0 13200.000000000002 170900.0 ;
      RECT  18800.0 170100.0 19600.0 170900.0 ;
      RECT  28000.000000000004 128700.00000000001 28800.0 129500.0 ;
      RECT  34800.00000000001 128700.00000000001 35600.0 129500.0 ;
      RECT  36400.00000000001 134700.00000000003 37200.0 135500.0 ;
      RECT  36400.00000000001 150300.0 37200.0 151100.0 ;
      RECT  36400.00000000001 153100.0 37200.0 153900.0 ;
      RECT  36400.00000000001 168700.00000000003 37200.0 169500.0 ;
      RECT  36400.00000000001 171500.0 37200.0 172300.0 ;
      RECT  36400.00000000001 187100.0 37200.0 187900.0 ;
      RECT  36400.00000000001 189900.0 37200.0 190700.00000000003 ;
      RECT  36400.00000000001 205500.0 37200.0 206300.0 ;
      RECT  2300.0000000000005 89400.0 1500.0000000000002 90199.99999999999 ;
      RECT  48800.00000000001 89400.0 48000.00000000001 90199.99999999999 ;
      RECT  28900.000000000004 50000.0 28100.0 50800.00000000001 ;
      RECT  51200.0 50000.0 52000.0 50800.00000000001 ;
      RECT  30300.0 28400.000000000004 29500.0 29200.000000000004 ;
      RECT  51200.0 28400.000000000004 52000.0 29200.000000000004 ;
      RECT  70000.0 39200.0 69200.0 40000.0 ;
      RECT  70000.0 59200.0 69200.0 60000.0 ;
      RECT  70000.0 19200.000000000004 69200.0 20000.0 ;
      RECT  70000.0 79200.0 69200.0 80000.0 ;
      RECT  70000.0 59200.0 69200.0 60000.0 ;
      RECT  70000.0 79200.0 69200.0 80000.0 ;
      RECT  70000.0 99200.00000000001 69200.0 100000.0 ;
      RECT  70000.0 119200.00000000001 69200.0 120000.0 ;
      RECT  70000.0 99200.00000000001 69200.0 100000.0 ;
      RECT  69200.0 39200.0 70000.0 40000.0 ;
      RECT  69200.0 79200.0 70000.0 80000.0 ;
      RECT  69200.0 119200.00000000001 70000.0 120000.0 ;
      RECT  31500.0 142600.0 32100.0 143200.00000000003 ;
      RECT  31500.0 161000.0 32100.0 161600.0 ;
      RECT  31500.0 179400.0 32100.0 180000.0 ;
      RECT  31500.0 197800.0 32100.0 198400.0 ;
      RECT  12400.0 142500.0 13200.000000000002 143300.0 ;
      RECT  18800.0 142500.0 19600.0 143300.0 ;
      RECT  12400.0 160900.0 13200.000000000002 161700.0 ;
      RECT  18800.0 160900.0 19600.0 161700.0 ;
      RECT  6000.0 124100.0 6800.000000000001 124900.0 ;
      RECT  31400.000000000004 122700.00000000001 32200.000000000004 123500.0 ;
      RECT  17200.0 129100.0 18000.0 129900.0 ;
      RECT  -400.0 39200.0 400.0 40000.0 ;
      RECT  69200.0 59200.0 70000.0 60000.00000000001 ;
      RECT  69200.0 19200.000000000004 70000.0 20000.0 ;
      RECT  69200.0 99200.00000000001 70000.0 100000.0 ;
      RECT  28100.0 138000.0 28700.000000000004 138600.0 ;
      RECT  34900.0 138000.0 35500.0 138600.0 ;
      RECT  28100.0 147200.00000000003 28700.000000000004 147800.0 ;
      RECT  34900.0 147200.00000000003 35500.0 147800.0 ;
      RECT  28100.0 156400.0 28700.000000000004 157000.0 ;
      RECT  34900.0 156400.0 35500.0 157000.0 ;
      RECT  28100.0 165600.0 28700.000000000004 166200.0 ;
      RECT  34900.0 165600.0 35500.0 166200.0 ;
      RECT  28100.0 174800.0 28700.000000000004 175400.0 ;
      RECT  34900.0 174800.0 35500.0 175400.0 ;
      RECT  28100.0 184000.0 28700.000000000004 184600.0 ;
      RECT  34900.0 184000.0 35500.0 184600.0 ;
      RECT  28100.0 193200.00000000003 28700.000000000004 193800.0 ;
      RECT  34900.0 193200.00000000003 35500.0 193800.0 ;
      RECT  28100.0 202400.0 28700.000000000004 203000.0 ;
      RECT  34900.0 202400.0 35500.0 203000.0 ;
      RECT  12400.0 133300.0 13200.000000000002 134100.0 ;
      RECT  18800.0 133300.0 19600.0 134100.0 ;
      RECT  12400.0 151700.0 13200.000000000002 152500.0 ;
      RECT  18800.0 151700.0 19600.0 152500.0 ;
      RECT  12400.0 170100.0 13200.000000000002 170900.0 ;
      RECT  18800.0 170100.0 19600.0 170900.0 ;
      RECT  28000.0 128700.00000000001 28800.0 129500.0 ;
      RECT  34800.00000000001 128700.00000000001 35600.0 129500.0 ;
      RECT  36400.0 134700.00000000003 37200.0 135500.0 ;
      RECT  36400.0 150300.0 37200.0 151100.0 ;
      RECT  36400.0 153100.0 37200.0 153900.0 ;
      RECT  36400.0 168700.0 37200.0 169500.0 ;
      RECT  36400.0 171500.0 37200.0 172300.0 ;
      RECT  36400.0 187100.0 37200.0 187900.0 ;
      RECT  36400.0 189900.0 37200.0 190700.00000000003 ;
      RECT  36400.0 205500.0 37200.0 206300.0 ;
      RECT  -400.0 19200.000000000004 400.0 20000.0 ;
      RECT  -400.0 59200.0 400.0 60000.00000000001 ;
      RECT  60500.0 231500.00000000003 59699.99999999999 232300.00000000003 ;
      RECT  60500.0 211500.00000000003 59699.99999999999 212300.00000000003 ;
      RECT  60500.0 231500.00000000003 59699.99999999999 232300.00000000003 ;
      RECT  60500.0 251500.00000000003 59699.99999999999 252300.00000000003 ;
      RECT  60500.0 271500.00000000006 59699.99999999999 272300.0 ;
      RECT  60500.0 251500.00000000003 59699.99999999999 252300.00000000003 ;
      RECT  60500.0 271500.00000000006 59699.99999999999 272300.0 ;
      RECT  60500.0 291500.00000000006 59699.99999999999 292300.00000000006 ;
      RECT  51999.99999999999 214900.00000000003 52800.0 215700.00000000006 ;
      RECT  49199.99999999999 215000.00000000003 71000.0 215600.00000000003 ;
      RECT  59699.99999999999 231500.00000000003 60500.0 232300.00000000003 ;
      RECT  59699.99999999999 271500.00000000006 60500.0 272300.00000000006 ;
      RECT  59699.99999999999 211500.00000000003 60500.0 212300.00000000003 ;
      RECT  59699.99999999999 251500.00000000003 60500.0 252300.00000000003 ;
      RECT  59699.99999999999 291500.00000000006 60500.0 292300.00000000006 ;
      RECT  189900.00000000003 19600.0 189100.00000000003 20400.000000000004 ;
      RECT  189900.00000000003 -400.0 189100.00000000003 400.0 ;
      RECT  211700.00000000003 19600.0 210900.00000000003 20400.000000000004 ;
      RECT  211700.00000000003 -400.0 210900.00000000003 400.0 ;
      RECT  181400.00000000003 3000.0 182200.00000000003 3800.0 ;
      RECT  203200.00000000003 3000.0 204000.00000000003 3800.0 ;
      RECT  178600.00000000003 3100.0 222200.00000000003 3700.0 ;
      RECT  189100.00000000003 19600.0 189900.00000000003 20400.000000000004 ;
      RECT  210900.00000000003 19600.0 211700.00000000003 20400.000000000004 ;
      RECT  189100.00000000003 -400.0 189900.00000000003 400.0 ;
      RECT  210900.00000000003 -400.0 211700.00000000003 400.0 ;
      RECT  173100.00000000003 3000.0 172300.0 3800.0 ;
      RECT  72800.0 214900.00000000003 72000.0 215700.00000000006 ;
      RECT  72800.0 50000.0 72000.0 50800.0 ;
      RECT  177300.0 108400.0 176500.0 109200.0 ;
      RECT  71399.99999999999 108400.0 70600.0 109200.0 ;
      RECT  175900.0 68400.0 175100.0 69200.0 ;
      RECT  71399.99999999999 68400.0 70600.0 69200.0 ;
      RECT  174500.0 28400.000000000004 173700.0 29200.000000000004 ;
      RECT  71399.99999999999 28400.000000000004 70600.0 29200.000000000004 ;
      RECT  173100.00000000003 50000.0 172300.0 50800.0 ;
      RECT  71399.99999999999 50000.0 70600.0 50800.0 ;
      RECT  74600.0 221300.0 73800.0 222100.00000000003 ;
      RECT  68800.0 221300.0 68000.0 222100.00000000003 ;
      RECT  76000.0 241700.0 75200.0 242500.0 ;
      RECT  68800.0 241700.0 68000.0 242500.0 ;
      RECT  77399.99999999999 261300.0 76600.0 262100.00000000003 ;
      RECT  68800.0 261300.0 68000.0 262100.00000000003 ;
      RECT  78800.0 281700.0 78000.0 282500.0 ;
      RECT  68800.0 281700.0 68000.0 282500.0 ;
      RECT  1500.0 1500.0 3300.0 3300.0 ;
      RECT  9900.0 1500.0 11700.000000000002 3300.0 ;
      RECT  19500.0 1500.0 21300.0 3300.0 ;
      RECT  29100.0 1500.0 30900.000000000004 3300.0 ;
      RECT  38700.0 1500.0 40500.0 3300.0 ;
      RECT  48300.00000000001 1500.0 50100.0 3300.0 ;
      RECT  57900.00000000001 1500.0 59700.0 3300.0 ;
      RECT  67500.0 1500.0 69300.0 3300.0 ;
      RECT  77100.00000000001 1500.0 78900.0 3300.0 ;
      RECT  86700.0 1500.0 88500.0 3300.0 ;
      RECT  96300.00000000001 1500.0 98100.00000000001 3300.0 ;
      RECT  105900.0 1500.0 107700.0 3300.0 ;
      RECT  115500.00000000001 1500.0 117300.00000000001 3300.0 ;
      RECT  125100.00000000001 1500.0 126900.0 3300.0 ;
      RECT  134700.0 1500.0 136500.0 3300.0 ;
      RECT  144299.99999999997 1500.0 146100.0 3300.0 ;
      RECT  153900.0 1500.0 155700.00000000003 3300.0 ;
      RECT  163500.0 1500.0 165300.0 3300.0 ;
      RECT  1500.0 9900.0 3300.0 11700.000000000002 ;
      RECT  9900.0 9900.0 11700.000000000002 11700.000000000002 ;
      RECT  19500.0 9900.0 21300.0 11700.000000000002 ;
      RECT  29100.0 9900.0 30900.000000000004 11700.000000000002 ;
      RECT  38700.0 9900.0 40500.0 11700.000000000002 ;
      RECT  48300.00000000001 9900.0 50100.0 11700.000000000002 ;
      RECT  57900.00000000001 9900.0 59700.0 11700.000000000002 ;
      RECT  67500.0 9900.0 69300.0 11700.000000000002 ;
      RECT  77100.00000000001 9900.0 78900.0 11700.000000000002 ;
      RECT  86700.0 9900.0 88500.0 11700.000000000002 ;
      RECT  96300.00000000001 9900.0 98100.00000000001 11700.000000000002 ;
      RECT  105900.0 9900.0 107700.0 11700.000000000002 ;
      RECT  115500.00000000001 9900.0 117300.00000000001 11700.000000000002 ;
      RECT  125100.00000000001 9900.0 126900.0 11700.000000000002 ;
      RECT  134700.0 9900.0 136500.0 11700.000000000002 ;
      RECT  144299.99999999997 9900.0 146100.0 11700.000000000002 ;
      RECT  153900.0 9900.0 155700.00000000003 11700.000000000002 ;
      RECT  163500.0 9900.0 165300.0 11700.000000000002 ;
      RECT  173100.0 9900.0 174900.0 11700.000000000002 ;
      RECT  182700.0 9900.0 184500.0 11700.000000000002 ;
      RECT  192300.0 9900.0 194100.00000000003 11700.000000000002 ;
      RECT  201900.0 9900.0 203700.00000000003 11700.000000000002 ;
      RECT  211500.0 9900.0 213300.0 11700.000000000002 ;
      RECT  221100.0 9900.0 222900.0 11700.000000000002 ;
      RECT  229500.0 9900.0 231300.0 11700.000000000002 ;
      RECT  1500.0 19500.0 3300.0 21300.0 ;
      RECT  9900.0 19500.0 11700.000000000002 21300.0 ;
      RECT  19500.0 19500.0 21300.0 21300.0 ;
      RECT  29100.0 19500.0 30900.000000000004 21300.0 ;
      RECT  38700.0 19500.0 40500.0 21300.0 ;
      RECT  48300.00000000001 19500.0 50100.0 21300.0 ;
      RECT  57900.00000000001 19500.0 59700.0 21300.0 ;
      RECT  67500.0 19500.0 69300.0 21300.0 ;
      RECT  77100.00000000001 19500.0 78900.0 21300.0 ;
      RECT  86700.0 19500.0 88500.0 21300.0 ;
      RECT  96300.00000000001 19500.0 98100.00000000001 21300.0 ;
      RECT  105900.0 19500.0 107700.0 21300.0 ;
      RECT  115500.00000000001 19500.0 117300.00000000001 21300.0 ;
      RECT  125100.00000000001 19500.0 126900.0 21300.0 ;
      RECT  134700.0 19500.0 136500.0 21300.0 ;
      RECT  144299.99999999997 19500.0 146100.0 21300.0 ;
      RECT  153900.0 19500.0 155700.00000000003 21300.0 ;
      RECT  163500.0 19500.0 165300.0 21300.0 ;
      RECT  173100.0 19500.0 174900.0 21300.0 ;
      RECT  181500.0 19500.0 183300.0 21300.0 ;
      RECT  221100.0 19500.0 222900.0 21300.0 ;
      RECT  229500.0 19500.0 231300.0 21300.0 ;
      RECT  201900.0 29100.0 203700.00000000003 30900.000000000004 ;
      RECT  211500.0 29100.0 213300.0 30900.000000000004 ;
      RECT  221100.0 29100.0 222900.0 30900.000000000004 ;
      RECT  229500.0 29100.0 231300.0 30900.000000000004 ;
      RECT  9900.0 38700.0 11700.000000000002 40500.0 ;
      RECT  19500.0 38700.0 21300.0 40500.0 ;
      RECT  29100.0 38700.0 30900.000000000004 40500.0 ;
      RECT  38700.0 38700.0 40500.0 40500.0 ;
      RECT  48300.00000000001 38700.0 50100.0 40500.0 ;
      RECT  57900.00000000001 38700.0 59700.0 40500.0 ;
      RECT  77100.00000000001 38700.0 78900.0 40500.0 ;
      RECT  86700.0 38700.0 88500.0 40500.0 ;
      RECT  96300.00000000001 38700.0 98100.00000000001 40500.0 ;
      RECT  105900.0 38700.0 107700.0 40500.0 ;
      RECT  115500.00000000001 38700.0 117300.00000000001 40500.0 ;
      RECT  125100.00000000001 38700.0 126900.0 40500.0 ;
      RECT  134700.0 38700.0 136500.0 40500.0 ;
      RECT  144299.99999999997 38700.0 146100.0 40500.0 ;
      RECT  153900.0 38700.0 155700.00000000003 40500.0 ;
      RECT  163500.0 38700.0 165300.0 40500.0 ;
      RECT  173100.0 38700.0 174900.0 40500.0 ;
      RECT  182700.0 38700.0 184500.0 40500.0 ;
      RECT  192300.0 38700.0 194100.00000000003 40500.0 ;
      RECT  201900.0 38700.0 203700.00000000003 40500.0 ;
      RECT  211500.0 38700.0 213300.0 40500.0 ;
      RECT  221100.0 38700.0 222900.0 40500.0 ;
      RECT  229500.0 38700.0 231300.0 40500.0 ;
      RECT  201900.0 48300.00000000001 203700.00000000003 50100.0 ;
      RECT  211500.0 48300.00000000001 213300.0 50100.0 ;
      RECT  221100.0 48300.00000000001 222900.0 50100.0 ;
      RECT  229500.0 48300.00000000001 231300.0 50100.0 ;
      RECT  1500.0 57900.00000000001 3300.0 59700.0 ;
      RECT  9900.0 57900.00000000001 11700.000000000002 59700.0 ;
      RECT  19500.0 57900.00000000001 21300.0 59700.0 ;
      RECT  29100.0 57900.00000000001 30900.000000000004 59700.0 ;
      RECT  38700.0 57900.00000000001 40500.0 59700.0 ;
      RECT  48300.00000000001 57900.00000000001 50100.0 59700.0 ;
      RECT  57900.00000000001 57900.00000000001 59700.0 59700.0 ;
      RECT  67500.0 57900.00000000001 69300.0 59700.0 ;
      RECT  77100.00000000001 57900.00000000001 78900.0 59700.0 ;
      RECT  86700.0 57900.00000000001 88500.0 59700.0 ;
      RECT  96300.00000000001 57900.00000000001 98100.00000000001 59700.0 ;
      RECT  105900.0 57900.00000000001 107700.0 59700.0 ;
      RECT  115500.00000000001 57900.00000000001 117300.00000000001 59700.0 ;
      RECT  125100.00000000001 57900.00000000001 126900.0 59700.0 ;
      RECT  134700.0 57900.00000000001 136500.0 59700.0 ;
      RECT  144299.99999999997 57900.00000000001 146100.0 59700.0 ;
      RECT  153900.0 57900.00000000001 155700.00000000003 59700.0 ;
      RECT  163500.0 57900.00000000001 165300.0 59700.0 ;
      RECT  173100.0 57900.00000000001 174900.0 59700.0 ;
      RECT  182700.0 57900.00000000001 184500.0 59700.0 ;
      RECT  192300.0 57900.00000000001 194100.00000000003 59700.0 ;
      RECT  201900.0 57900.00000000001 203700.00000000003 59700.0 ;
      RECT  211500.0 57900.00000000001 213300.0 59700.0 ;
      RECT  221100.0 57900.00000000001 222900.0 59700.0 ;
      RECT  229500.0 57900.00000000001 231300.0 59700.0 ;
      RECT  1500.0 67500.0 3300.0 69300.0 ;
      RECT  9900.0 67500.0 11700.000000000002 69300.0 ;
      RECT  19500.0 67500.0 21300.0 69300.0 ;
      RECT  29100.0 67500.0 30900.000000000004 69300.0 ;
      RECT  38700.0 67500.0 40500.0 69300.0 ;
      RECT  48300.00000000001 67500.0 50100.0 69300.0 ;
      RECT  57900.00000000001 67500.0 59700.0 69300.0 ;
      RECT  182700.0 67500.0 184500.0 69300.0 ;
      RECT  192300.0 67500.0 194100.00000000003 69300.0 ;
      RECT  201900.0 67500.0 203700.00000000003 69300.0 ;
      RECT  211500.0 67500.0 213300.0 69300.0 ;
      RECT  221100.0 67500.0 222900.0 69300.0 ;
      RECT  229500.0 67500.0 231300.0 69300.0 ;
      RECT  1500.0 77100.00000000001 3300.0 78900.0 ;
      RECT  9900.0 77100.00000000001 11700.000000000002 78900.0 ;
      RECT  19500.0 77100.00000000001 21300.0 78900.0 ;
      RECT  29100.0 77100.00000000001 30900.000000000004 78900.0 ;
      RECT  38700.0 77100.00000000001 40500.0 78900.0 ;
      RECT  48300.00000000001 77100.00000000001 50100.0 78900.0 ;
      RECT  57900.00000000001 77100.00000000001 59700.0 78900.0 ;
      RECT  77100.00000000001 77100.00000000001 78900.0 78900.0 ;
      RECT  86700.0 77100.00000000001 88500.0 78900.0 ;
      RECT  96300.00000000001 77100.00000000001 98100.00000000001 78900.0 ;
      RECT  105900.0 77100.00000000001 107700.0 78900.0 ;
      RECT  115500.00000000001 77100.00000000001 117300.00000000001 78900.0 ;
      RECT  125100.00000000001 77100.00000000001 126900.0 78900.0 ;
      RECT  134700.0 77100.00000000001 136500.0 78900.0 ;
      RECT  144299.99999999997 77100.00000000001 146100.0 78900.0 ;
      RECT  153900.0 77100.00000000001 155700.00000000003 78900.0 ;
      RECT  163500.0 77100.00000000001 165300.0 78900.0 ;
      RECT  173100.0 77100.00000000001 174900.0 78900.0 ;
      RECT  182700.0 77100.00000000001 184500.0 78900.0 ;
      RECT  192300.0 77100.00000000001 194100.00000000003 78900.0 ;
      RECT  201900.0 77100.00000000001 203700.00000000003 78900.0 ;
      RECT  211500.0 77100.00000000001 213300.0 78900.0 ;
      RECT  221100.0 77100.00000000001 222900.0 78900.0 ;
      RECT  229500.0 77100.00000000001 231300.0 78900.0 ;
      RECT  57900.00000000001 86700.0 59700.0 88500.0 ;
      RECT  67500.0 86700.0 69300.0 88500.0 ;
      RECT  77100.00000000001 86700.0 78900.0 88500.0 ;
      RECT  86700.0 86700.0 88500.0 88500.0 ;
      RECT  96300.00000000001 86700.0 98100.00000000001 88500.0 ;
      RECT  105900.0 86700.0 107700.0 88500.0 ;
      RECT  115500.00000000001 86700.0 117300.00000000001 88500.0 ;
      RECT  125100.00000000001 86700.0 126900.0 88500.0 ;
      RECT  134700.0 86700.0 136500.0 88500.0 ;
      RECT  144299.99999999997 86700.0 146100.0 88500.0 ;
      RECT  153900.0 86700.0 155700.00000000003 88500.0 ;
      RECT  163500.0 86700.0 165300.0 88500.0 ;
      RECT  173100.0 86700.0 174900.0 88500.0 ;
      RECT  182700.0 86700.0 184500.0 88500.0 ;
      RECT  192300.0 86700.0 194100.00000000003 88500.0 ;
      RECT  201900.0 86700.0 203700.00000000003 88500.0 ;
      RECT  211500.0 86700.0 213300.0 88500.0 ;
      RECT  221100.0 86700.0 222900.0 88500.0 ;
      RECT  229500.0 86700.0 231300.0 88500.0 ;
      RECT  1500.0 96300.00000000001 3300.0 98100.00000000001 ;
      RECT  9900.0 96300.00000000001 11700.000000000002 98100.00000000001 ;
      RECT  19500.0 96300.00000000001 21300.0 98100.00000000001 ;
      RECT  29100.0 96300.00000000001 30900.000000000004 98100.00000000001 ;
      RECT  38700.0 96300.00000000001 40500.0 98100.00000000001 ;
      RECT  48300.00000000001 96300.00000000001 50100.0 98100.00000000001 ;
      RECT  57900.00000000001 96300.00000000001 59700.0 98100.00000000001 ;
      RECT  67500.0 96300.00000000001 69300.0 98100.00000000001 ;
      RECT  77100.00000000001 96300.00000000001 78900.0 98100.00000000001 ;
      RECT  86700.0 96300.00000000001 88500.0 98100.00000000001 ;
      RECT  96300.00000000001 96300.00000000001 98100.00000000001 98100.00000000001 ;
      RECT  105900.0 96300.00000000001 107700.0 98100.00000000001 ;
      RECT  115500.00000000001 96300.00000000001 117300.00000000001 98100.00000000001 ;
      RECT  125100.00000000001 96300.00000000001 126900.0 98100.00000000001 ;
      RECT  134700.0 96300.00000000001 136500.0 98100.00000000001 ;
      RECT  144299.99999999997 96300.00000000001 146100.0 98100.00000000001 ;
      RECT  153900.0 96300.00000000001 155700.00000000003 98100.00000000001 ;
      RECT  163500.0 96300.00000000001 165300.0 98100.00000000001 ;
      RECT  173100.0 96300.00000000001 174900.0 98100.00000000001 ;
      RECT  182700.0 96300.00000000001 184500.0 98100.00000000001 ;
      RECT  192300.0 96300.00000000001 194100.00000000003 98100.00000000001 ;
      RECT  201900.0 96300.00000000001 203700.00000000003 98100.00000000001 ;
      RECT  211500.0 96300.00000000001 213300.0 98100.00000000001 ;
      RECT  221100.0 96300.00000000001 222900.0 98100.00000000001 ;
      RECT  229500.0 96300.00000000001 231300.0 98100.00000000001 ;
      RECT  1500.0 105900.0 3300.0 107700.0 ;
      RECT  9900.0 105900.0 11700.000000000002 107700.0 ;
      RECT  19500.0 105900.0 21300.0 107700.0 ;
      RECT  29100.0 105900.0 30900.000000000004 107700.0 ;
      RECT  38700.0 105900.0 40500.0 107700.0 ;
      RECT  48300.00000000001 105900.0 50100.0 107700.0 ;
      RECT  57900.00000000001 105900.0 59700.0 107700.0 ;
      RECT  183900.0 105900.0 185700.00000000003 107700.0 ;
      RECT  192300.0 105900.0 194100.00000000003 107700.0 ;
      RECT  201900.0 105900.0 203700.00000000003 107700.0 ;
      RECT  211500.0 105900.0 213300.0 107700.0 ;
      RECT  221100.0 105900.0 222900.0 107700.0 ;
      RECT  229500.0 105900.0 231300.0 107700.0 ;
      RECT  1500.0 115500.00000000001 3300.0 117300.00000000001 ;
      RECT  9900.0 115500.00000000001 11700.000000000002 117300.00000000001 ;
      RECT  19500.0 115500.00000000001 21300.0 117300.00000000001 ;
      RECT  29100.0 115500.00000000001 30900.000000000004 117300.00000000001 ;
      RECT  38700.0 115500.00000000001 40500.0 117300.00000000001 ;
      RECT  48300.00000000001 115500.00000000001 50100.0 117300.00000000001 ;
      RECT  57900.00000000001 115500.00000000001 59700.0 117300.00000000001 ;
      RECT  67500.0 115500.00000000001 69300.0 117300.00000000001 ;
      RECT  77100.00000000001 115500.00000000001 78900.0 117300.00000000001 ;
      RECT  86700.0 115500.00000000001 88500.0 117300.00000000001 ;
      RECT  96300.00000000001 115500.00000000001 98100.00000000001 117300.00000000001 ;
      RECT  105900.0 115500.00000000001 107700.0 117300.00000000001 ;
      RECT  115500.00000000001 115500.00000000001 117300.00000000001 117300.00000000001 ;
      RECT  125100.00000000001 115500.00000000001 126900.0 117300.00000000001 ;
      RECT  134700.0 115500.00000000001 136500.0 117300.00000000001 ;
      RECT  144299.99999999997 115500.00000000001 146100.0 117300.00000000001 ;
      RECT  153900.0 115500.00000000001 155700.00000000003 117300.00000000001 ;
      RECT  163500.0 115500.00000000001 165300.0 117300.00000000001 ;
      RECT  173100.0 115500.00000000001 174900.0 117300.00000000001 ;
      RECT  182700.0 115500.00000000001 184500.0 117300.00000000001 ;
      RECT  192300.0 115500.00000000001 194100.00000000003 117300.00000000001 ;
      RECT  201900.0 115500.00000000001 203700.00000000003 117300.00000000001 ;
      RECT  211500.0 115500.00000000001 213300.0 117300.00000000001 ;
      RECT  221100.0 115500.00000000001 222900.0 117300.00000000001 ;
      RECT  229500.0 115500.00000000001 231300.0 117300.00000000001 ;
      RECT  39900.00000000001 125100.00000000001 41700.0 126900.0 ;
      RECT  48300.00000000001 125100.00000000001 50100.0 126900.0 ;
      RECT  57900.00000000001 125100.00000000001 59700.0 126900.0 ;
      RECT  67500.0 125100.00000000001 69300.0 126900.0 ;
      RECT  77100.00000000001 125100.00000000001 78900.0 126900.0 ;
      RECT  86700.0 125100.00000000001 88500.0 126900.0 ;
      RECT  96300.00000000001 125100.00000000001 98100.00000000001 126900.0 ;
      RECT  105900.0 125100.00000000001 107700.0 126900.0 ;
      RECT  115500.00000000001 125100.00000000001 117300.00000000001 126900.0 ;
      RECT  125100.00000000001 125100.00000000001 126900.0 126900.0 ;
      RECT  134700.0 125100.00000000001 136500.0 126900.0 ;
      RECT  144299.99999999997 125100.00000000001 146100.0 126900.0 ;
      RECT  153900.0 125100.00000000001 155700.00000000003 126900.0 ;
      RECT  163500.0 125100.00000000001 165300.0 126900.0 ;
      RECT  173100.0 125100.00000000001 174900.0 126900.0 ;
      RECT  182700.0 125100.00000000001 184500.0 126900.0 ;
      RECT  192300.0 125100.00000000001 194100.00000000003 126900.0 ;
      RECT  201900.0 125100.00000000001 203700.00000000003 126900.0 ;
      RECT  211500.0 125100.00000000001 213300.0 126900.0 ;
      RECT  221100.0 125100.00000000001 222900.0 126900.0 ;
      RECT  229500.0 125100.00000000001 231300.0 126900.0 ;
      RECT  29100.0 134700.0 30900.000000000004 136500.0 ;
      RECT  38700.0 134700.0 40500.0 136500.0 ;
      RECT  48300.00000000001 134700.0 50100.0 136500.0 ;
      RECT  57900.00000000001 134700.0 59700.0 136500.0 ;
      RECT  66300.00000000001 134700.0 68100.00000000001 136500.0 ;
      RECT  87900.0 134700.0 89700.0 136500.0 ;
      RECT  96300.00000000001 134700.0 98100.00000000001 136500.0 ;
      RECT  105900.0 134700.0 107700.0 136500.0 ;
      RECT  115500.00000000001 134700.0 117300.00000000001 136500.0 ;
      RECT  125100.00000000001 134700.0 126900.0 136500.0 ;
      RECT  134700.0 134700.0 136500.0 136500.0 ;
      RECT  144299.99999999997 134700.0 146100.0 136500.0 ;
      RECT  153900.0 134700.0 155700.00000000003 136500.0 ;
      RECT  163500.0 134700.0 165300.0 136500.0 ;
      RECT  173100.0 134700.0 174900.0 136500.0 ;
      RECT  182700.0 134700.0 184500.0 136500.0 ;
      RECT  192300.0 134700.0 194100.00000000003 136500.0 ;
      RECT  201900.0 134700.0 203700.00000000003 136500.0 ;
      RECT  211500.0 134700.0 213300.0 136500.0 ;
      RECT  221100.0 134700.0 222900.0 136500.0 ;
      RECT  229500.0 134700.0 231300.0 136500.0 ;
      RECT  39900.00000000001 144299.99999999997 41700.0 146100.0 ;
      RECT  48300.00000000001 144299.99999999997 50100.0 146100.0 ;
      RECT  57900.00000000001 144299.99999999997 59700.0 146100.0 ;
      RECT  66300.00000000001 144299.99999999997 68100.00000000001 146100.0 ;
      RECT  96300.00000000001 144299.99999999997 98100.00000000001 146100.0 ;
      RECT  105900.0 144299.99999999997 107700.0 146100.0 ;
      RECT  115500.00000000001 144299.99999999997 117300.00000000001 146100.0 ;
      RECT  125100.00000000001 144299.99999999997 126900.0 146100.0 ;
      RECT  134700.0 144299.99999999997 136500.0 146100.0 ;
      RECT  144299.99999999997 144299.99999999997 146100.0 146100.0 ;
      RECT  153900.0 144299.99999999997 155700.00000000003 146100.0 ;
      RECT  163500.0 144299.99999999997 165300.0 146100.0 ;
      RECT  173100.0 144299.99999999997 174900.0 146100.0 ;
      RECT  182700.0 144299.99999999997 184500.0 146100.0 ;
      RECT  192300.0 144299.99999999997 194100.00000000003 146100.0 ;
      RECT  201900.0 144299.99999999997 203700.00000000003 146100.0 ;
      RECT  211500.0 144299.99999999997 213300.0 146100.0 ;
      RECT  221100.0 144299.99999999997 222900.0 146100.0 ;
      RECT  229500.0 144299.99999999997 231300.0 146100.0 ;
      RECT  29100.0 153900.0 30900.000000000004 155700.00000000003 ;
      RECT  38700.0 153900.0 40500.0 155700.00000000003 ;
      RECT  48300.00000000001 153900.0 50100.0 155700.00000000003 ;
      RECT  57900.00000000001 153900.0 59700.0 155700.00000000003 ;
      RECT  67500.0 153900.0 69300.0 155700.00000000003 ;
      RECT  77100.00000000001 153900.0 78900.0 155700.00000000003 ;
      RECT  86700.0 153900.0 88500.0 155700.00000000003 ;
      RECT  96300.00000000001 153900.0 98100.00000000001 155700.00000000003 ;
      RECT  105900.0 153900.0 107700.0 155700.00000000003 ;
      RECT  115500.00000000001 153900.0 117300.00000000001 155700.00000000003 ;
      RECT  125100.00000000001 153900.0 126900.0 155700.00000000003 ;
      RECT  134700.0 153900.0 136500.0 155700.00000000003 ;
      RECT  144299.99999999997 153900.0 146100.0 155700.00000000003 ;
      RECT  153900.0 153900.0 155700.00000000003 155700.00000000003 ;
      RECT  163500.0 153900.0 165300.0 155700.00000000003 ;
      RECT  173100.0 153900.0 174900.0 155700.00000000003 ;
      RECT  182700.0 153900.0 184500.0 155700.00000000003 ;
      RECT  192300.0 153900.0 194100.00000000003 155700.00000000003 ;
      RECT  201900.0 153900.0 203700.00000000003 155700.00000000003 ;
      RECT  211500.0 153900.0 213300.0 155700.00000000003 ;
      RECT  221100.0 153900.0 222900.0 155700.00000000003 ;
      RECT  229500.0 153900.0 231300.0 155700.00000000003 ;
      RECT  39900.00000000001 163500.0 41700.0 165300.0 ;
      RECT  48300.00000000001 163500.0 50100.0 165300.0 ;
      RECT  57900.00000000001 163500.0 59700.0 165300.0 ;
      RECT  67500.0 163500.0 69300.0 165300.0 ;
      RECT  77100.00000000001 163500.0 78900.0 165300.0 ;
      RECT  86700.0 163500.0 88500.0 165300.0 ;
      RECT  96300.00000000001 163500.0 98100.00000000001 165300.0 ;
      RECT  105900.0 163500.0 107700.0 165300.0 ;
      RECT  115500.00000000001 163500.0 117300.00000000001 165300.0 ;
      RECT  125100.00000000001 163500.0 126900.0 165300.0 ;
      RECT  134700.0 163500.0 136500.0 165300.0 ;
      RECT  144299.99999999997 163500.0 146100.0 165300.0 ;
      RECT  153900.0 163500.0 155700.00000000003 165300.0 ;
      RECT  163500.0 163500.0 165300.0 165300.0 ;
      RECT  173100.0 163500.0 174900.0 165300.0 ;
      RECT  182700.0 163500.0 184500.0 165300.0 ;
      RECT  192300.0 163500.0 194100.00000000003 165300.0 ;
      RECT  201900.0 163500.0 203700.00000000003 165300.0 ;
      RECT  211500.0 163500.0 213300.0 165300.0 ;
      RECT  221100.0 163500.0 222900.0 165300.0 ;
      RECT  229500.0 163500.0 231300.0 165300.0 ;
      RECT  1500.0 173100.0 3300.0 174900.0 ;
      RECT  9900.0 173100.0 11700.000000000002 174900.0 ;
      RECT  19500.0 173100.0 21300.0 174900.0 ;
      RECT  29100.0 173100.0 30900.000000000004 174900.0 ;
      RECT  38700.0 173100.0 40500.0 174900.0 ;
      RECT  48300.00000000001 173100.0 50100.0 174900.0 ;
      RECT  57900.00000000001 173100.0 59700.0 174900.0 ;
      RECT  67500.0 173100.0 69300.0 174900.0 ;
      RECT  77100.00000000001 173100.0 78900.0 174900.0 ;
      RECT  86700.0 173100.0 88500.0 174900.0 ;
      RECT  96300.00000000001 173100.0 98100.00000000001 174900.0 ;
      RECT  105900.0 173100.0 107700.0 174900.0 ;
      RECT  115500.00000000001 173100.0 117300.00000000001 174900.0 ;
      RECT  125100.00000000001 173100.0 126900.0 174900.0 ;
      RECT  134700.0 173100.0 136500.0 174900.0 ;
      RECT  144299.99999999997 173100.0 146100.0 174900.0 ;
      RECT  153900.0 173100.0 155700.00000000003 174900.0 ;
      RECT  163500.0 173100.0 165300.0 174900.0 ;
      RECT  173100.0 173100.0 174900.0 174900.0 ;
      RECT  182700.0 173100.0 184500.0 174900.0 ;
      RECT  192300.0 173100.0 194100.00000000003 174900.0 ;
      RECT  201900.0 173100.0 203700.00000000003 174900.0 ;
      RECT  211500.0 173100.0 213300.0 174900.0 ;
      RECT  221100.0 173100.0 222900.0 174900.0 ;
      RECT  229500.0 173100.0 231300.0 174900.0 ;
      RECT  1500.0 182700.0 3300.0 184500.0 ;
      RECT  9900.0 182700.0 11700.000000000002 184500.0 ;
      RECT  19500.0 182700.0 21300.0 184500.0 ;
      RECT  29100.0 182700.0 30900.000000000004 184500.0 ;
      RECT  38700.0 182700.0 40500.0 184500.0 ;
      RECT  48300.00000000001 182700.0 50100.0 184500.0 ;
      RECT  57900.00000000001 182700.0 59700.0 184500.0 ;
      RECT  67500.0 182700.0 69300.0 184500.0 ;
      RECT  77100.00000000001 182700.0 78900.0 184500.0 ;
      RECT  86700.0 182700.0 88500.0 184500.0 ;
      RECT  96300.00000000001 182700.0 98100.00000000001 184500.0 ;
      RECT  105900.0 182700.0 107700.0 184500.0 ;
      RECT  115500.00000000001 182700.0 117300.00000000001 184500.0 ;
      RECT  125100.00000000001 182700.0 126900.0 184500.0 ;
      RECT  134700.0 182700.0 136500.0 184500.0 ;
      RECT  144299.99999999997 182700.0 146100.0 184500.0 ;
      RECT  153900.0 182700.0 155700.00000000003 184500.0 ;
      RECT  163500.0 182700.0 165300.0 184500.0 ;
      RECT  173100.0 182700.0 174900.0 184500.0 ;
      RECT  182700.0 182700.0 184500.0 184500.0 ;
      RECT  192300.0 182700.0 194100.00000000003 184500.0 ;
      RECT  201900.0 182700.0 203700.00000000003 184500.0 ;
      RECT  211500.0 182700.0 213300.0 184500.0 ;
      RECT  221100.0 182700.0 222900.0 184500.0 ;
      RECT  229500.0 182700.0 231300.0 184500.0 ;
      RECT  1500.0 192300.0 3300.0 194100.00000000003 ;
      RECT  9900.0 192300.0 11700.000000000002 194100.00000000003 ;
      RECT  19500.0 192300.0 21300.0 194100.00000000003 ;
      RECT  29100.0 192300.0 30900.000000000004 194100.00000000003 ;
      RECT  38700.0 192300.0 40500.0 194100.00000000003 ;
      RECT  48300.00000000001 192300.0 50100.0 194100.00000000003 ;
      RECT  57900.00000000001 192300.0 59700.0 194100.00000000003 ;
      RECT  67500.0 192300.0 69300.0 194100.00000000003 ;
      RECT  77100.00000000001 192300.0 78900.0 194100.00000000003 ;
      RECT  86700.0 192300.0 88500.0 194100.00000000003 ;
      RECT  96300.00000000001 192300.0 98100.00000000001 194100.00000000003 ;
      RECT  105900.0 192300.0 107700.0 194100.00000000003 ;
      RECT  115500.00000000001 192300.0 117300.00000000001 194100.00000000003 ;
      RECT  125100.00000000001 192300.0 126900.0 194100.00000000003 ;
      RECT  134700.0 192300.0 136500.0 194100.00000000003 ;
      RECT  144299.99999999997 192300.0 146100.0 194100.00000000003 ;
      RECT  153900.0 192300.0 155700.00000000003 194100.00000000003 ;
      RECT  163500.0 192300.0 165300.0 194100.00000000003 ;
      RECT  173100.0 192300.0 174900.0 194100.00000000003 ;
      RECT  182700.0 192300.0 184500.0 194100.00000000003 ;
      RECT  192300.0 192300.0 194100.00000000003 194100.00000000003 ;
      RECT  201900.0 192300.0 203700.00000000003 194100.00000000003 ;
      RECT  211500.0 192300.0 213300.0 194100.00000000003 ;
      RECT  221100.0 192300.0 222900.0 194100.00000000003 ;
      RECT  229500.0 192300.0 231300.0 194100.00000000003 ;
      RECT  1500.0 201900.0 3300.0 203700.00000000003 ;
      RECT  9900.0 201900.0 11700.000000000002 203700.00000000003 ;
      RECT  19500.0 201900.0 21300.0 203700.00000000003 ;
      RECT  29100.0 201900.0 30900.000000000004 203700.00000000003 ;
      RECT  38700.0 201900.0 40500.0 203700.00000000003 ;
      RECT  48300.00000000001 201900.0 50100.0 203700.00000000003 ;
      RECT  57900.00000000001 201900.0 59700.0 203700.00000000003 ;
      RECT  67500.0 201900.0 69300.0 203700.00000000003 ;
      RECT  77100.00000000001 201900.0 78900.0 203700.00000000003 ;
      RECT  86700.0 201900.0 88500.0 203700.00000000003 ;
      RECT  96300.00000000001 201900.0 98100.00000000001 203700.00000000003 ;
      RECT  105900.0 201900.0 107700.0 203700.00000000003 ;
      RECT  115500.00000000001 201900.0 117300.00000000001 203700.00000000003 ;
      RECT  201900.0 201900.0 203700.00000000003 203700.00000000003 ;
      RECT  211500.0 201900.0 213300.0 203700.00000000003 ;
      RECT  221100.0 201900.0 222900.0 203700.00000000003 ;
      RECT  229500.0 201900.0 231300.0 203700.00000000003 ;
      RECT  1500.0 211500.0 3300.0 213300.0 ;
      RECT  9900.0 211500.0 11700.000000000002 213300.0 ;
      RECT  19500.0 211500.0 21300.0 213300.0 ;
      RECT  29100.0 211500.0 30900.000000000004 213300.0 ;
      RECT  38700.0 211500.0 40500.0 213300.0 ;
      RECT  78300.00000000001 211500.0 80100.00000000001 213300.0 ;
      RECT  86700.0 211500.0 88500.0 213300.0 ;
      RECT  96300.00000000001 211500.0 98100.00000000001 213300.0 ;
      RECT  105900.0 211500.0 107700.0 213300.0 ;
      RECT  115500.00000000001 211500.0 117300.00000000001 213300.0 ;
      RECT  125100.00000000001 211500.0 126900.0 213300.0 ;
      RECT  134700.0 211500.0 136500.0 213300.0 ;
      RECT  144299.99999999997 211500.0 146100.0 213300.0 ;
      RECT  153900.0 211500.0 155700.00000000003 213300.0 ;
      RECT  163500.0 211500.0 165300.0 213300.0 ;
      RECT  173100.0 211500.0 174900.0 213300.0 ;
      RECT  182700.0 211500.0 184500.0 213300.0 ;
      RECT  192300.0 211500.0 194100.00000000003 213300.0 ;
      RECT  201900.0 211500.0 203700.00000000003 213300.0 ;
      RECT  211500.0 211500.0 213300.0 213300.0 ;
      RECT  221100.0 211500.0 222900.0 213300.0 ;
      RECT  229500.0 211500.0 231300.0 213300.0 ;
      RECT  1500.0 221100.0 3300.0 222900.0 ;
      RECT  9900.0 221100.0 11700.000000000002 222900.0 ;
      RECT  19500.0 221100.0 21300.0 222900.0 ;
      RECT  29100.0 221100.0 30900.000000000004 222900.0 ;
      RECT  38700.0 221100.0 40500.0 222900.0 ;
      RECT  48300.00000000001 221100.0 50100.0 222900.0 ;
      RECT  57900.00000000001 221100.0 59700.0 222900.0 ;
      RECT  86700.0 221100.0 88500.0 222900.0 ;
      RECT  96300.00000000001 221100.0 98100.00000000001 222900.0 ;
      RECT  105900.0 221100.0 107700.0 222900.0 ;
      RECT  115500.00000000001 221100.0 117300.00000000001 222900.0 ;
      RECT  201900.0 221100.0 203700.00000000003 222900.0 ;
      RECT  211500.0 221100.0 213300.0 222900.0 ;
      RECT  221100.0 221100.0 222900.0 222900.0 ;
      RECT  229500.0 221100.0 231300.0 222900.0 ;
      RECT  1500.0 230700.0 3300.0 232500.0 ;
      RECT  9900.0 230700.0 11700.000000000002 232500.0 ;
      RECT  19500.0 230700.0 21300.0 232500.0 ;
      RECT  29100.0 230700.0 30900.000000000004 232500.0 ;
      RECT  38700.0 230700.0 40500.0 232500.0 ;
      RECT  48300.00000000001 230700.0 50100.0 232500.0 ;
      RECT  67500.0 230700.0 69300.0 232500.0 ;
      RECT  77100.00000000001 230700.0 78900.0 232500.0 ;
      RECT  86700.0 230700.0 88500.0 232500.0 ;
      RECT  96300.00000000001 230700.0 98100.00000000001 232500.0 ;
      RECT  105900.0 230700.0 107700.0 232500.0 ;
      RECT  115500.00000000001 230700.0 117300.00000000001 232500.0 ;
      RECT  125100.00000000001 230700.0 126900.0 232500.0 ;
      RECT  134700.0 230700.0 136500.0 232500.0 ;
      RECT  144299.99999999997 230700.0 146100.0 232500.0 ;
      RECT  153900.0 230700.0 155700.00000000003 232500.0 ;
      RECT  163500.0 230700.0 165300.0 232500.0 ;
      RECT  173100.0 230700.0 174900.0 232500.0 ;
      RECT  182700.0 230700.0 184500.0 232500.0 ;
      RECT  192300.0 230700.0 194100.00000000003 232500.0 ;
      RECT  201900.0 230700.0 203700.00000000003 232500.0 ;
      RECT  211500.0 230700.0 213300.0 232500.0 ;
      RECT  221100.0 230700.0 222900.0 232500.0 ;
      RECT  229500.0 230700.0 231300.0 232500.0 ;
      RECT  1500.0 240300.0 3300.0 242100.00000000003 ;
      RECT  9900.0 240300.0 11700.000000000002 242100.00000000003 ;
      RECT  19500.0 240300.0 21300.0 242100.00000000003 ;
      RECT  29100.0 240300.0 30900.000000000004 242100.00000000003 ;
      RECT  38700.0 240300.0 40500.0 242100.00000000003 ;
      RECT  48300.00000000001 240300.0 50100.0 242100.00000000003 ;
      RECT  57900.00000000001 240300.0 59700.0 242100.00000000003 ;
      RECT  86700.0 240300.0 88500.0 242100.00000000003 ;
      RECT  96300.00000000001 240300.0 98100.00000000001 242100.00000000003 ;
      RECT  105900.0 240300.0 107700.0 242100.00000000003 ;
      RECT  115500.00000000001 240300.0 117300.00000000001 242100.00000000003 ;
      RECT  201900.0 240300.0 203700.00000000003 242100.00000000003 ;
      RECT  211500.0 240300.0 213300.0 242100.00000000003 ;
      RECT  221100.0 240300.0 222900.0 242100.00000000003 ;
      RECT  229500.0 240300.0 231300.0 242100.00000000003 ;
      RECT  1500.0 249900.0 3300.0 251700.00000000003 ;
      RECT  9900.0 249900.0 11700.000000000002 251700.00000000003 ;
      RECT  19500.0 249900.0 21300.0 251700.00000000003 ;
      RECT  29100.0 249900.0 30900.000000000004 251700.00000000003 ;
      RECT  38700.0 249900.0 40500.0 251700.00000000003 ;
      RECT  48300.00000000001 249900.0 50100.0 251700.00000000003 ;
      RECT  57900.00000000001 249900.0 59700.0 251700.00000000003 ;
      RECT  67500.0 249900.0 69300.0 251700.00000000003 ;
      RECT  77100.00000000001 249900.0 78900.0 251700.00000000003 ;
      RECT  86700.0 249900.0 88500.0 251700.00000000003 ;
      RECT  96300.00000000001 249900.0 98100.00000000001 251700.00000000003 ;
      RECT  105900.0 249900.0 107700.0 251700.00000000003 ;
      RECT  115500.00000000001 249900.0 117300.00000000001 251700.00000000003 ;
      RECT  125100.00000000001 249900.0 126900.0 251700.00000000003 ;
      RECT  134700.0 249900.0 136500.0 251700.00000000003 ;
      RECT  144299.99999999997 249900.0 146100.0 251700.00000000003 ;
      RECT  153900.0 249900.0 155700.00000000003 251700.00000000003 ;
      RECT  163500.0 249900.0 165300.0 251700.00000000003 ;
      RECT  173100.0 249900.0 174900.0 251700.00000000003 ;
      RECT  182700.0 249900.0 184500.0 251700.00000000003 ;
      RECT  192300.0 249900.0 194100.00000000003 251700.00000000003 ;
      RECT  201900.0 249900.0 203700.00000000003 251700.00000000003 ;
      RECT  211500.0 249900.0 213300.0 251700.00000000003 ;
      RECT  221100.0 249900.0 222900.0 251700.00000000003 ;
      RECT  229500.0 249900.0 231300.0 251700.00000000003 ;
      RECT  1500.0 259500.0 3300.0 261300.0 ;
      RECT  9900.0 259500.0 11700.000000000002 261300.0 ;
      RECT  19500.0 259500.0 21300.0 261300.0 ;
      RECT  29100.0 259500.0 30900.000000000004 261300.0 ;
      RECT  38700.0 259500.0 40500.0 261300.0 ;
      RECT  48300.00000000001 259500.0 50100.0 261300.0 ;
      RECT  57900.00000000001 259500.0 59700.0 261300.0 ;
      RECT  86700.0 259500.0 88500.0 261300.0 ;
      RECT  96300.00000000001 259500.0 98100.00000000001 261300.0 ;
      RECT  105900.0 259500.0 107700.0 261300.0 ;
      RECT  115500.00000000001 259500.0 117300.00000000001 261300.0 ;
      RECT  201900.0 259500.0 203700.00000000003 261300.0 ;
      RECT  211500.0 259500.0 213300.0 261300.0 ;
      RECT  221100.0 259500.0 222900.0 261300.0 ;
      RECT  229500.0 259500.0 231300.0 261300.0 ;
      RECT  1500.0 269100.0 3300.0 270900.00000000006 ;
      RECT  9900.0 269100.0 11700.000000000002 270900.00000000006 ;
      RECT  19500.0 269100.0 21300.0 270900.00000000006 ;
      RECT  29100.0 269100.0 30900.000000000004 270900.00000000006 ;
      RECT  38700.0 269100.0 40500.0 270900.00000000006 ;
      RECT  48300.00000000001 269100.0 50100.0 270900.00000000006 ;
      RECT  67500.0 269100.0 69300.0 270900.00000000006 ;
      RECT  77100.00000000001 269100.0 78900.0 270900.00000000006 ;
      RECT  86700.0 269100.0 88500.0 270900.00000000006 ;
      RECT  96300.00000000001 269100.0 98100.00000000001 270900.00000000006 ;
      RECT  105900.0 269100.0 107700.0 270900.00000000006 ;
      RECT  115500.00000000001 269100.0 117300.00000000001 270900.00000000006 ;
      RECT  125100.00000000001 269100.0 126900.0 270900.00000000006 ;
      RECT  134700.0 269100.0 136500.0 270900.00000000006 ;
      RECT  144299.99999999997 269100.0 146100.0 270900.00000000006 ;
      RECT  153900.0 269100.0 155700.00000000003 270900.00000000006 ;
      RECT  163500.0 269100.0 165300.0 270900.00000000006 ;
      RECT  173100.0 269100.0 174900.0 270900.00000000006 ;
      RECT  182700.0 269100.0 184500.0 270900.00000000006 ;
      RECT  192300.0 269100.0 194100.00000000003 270900.00000000006 ;
      RECT  201900.0 269100.0 203700.00000000003 270900.00000000006 ;
      RECT  211500.0 269100.0 213300.0 270900.00000000006 ;
      RECT  221100.0 269100.0 222900.0 270900.00000000006 ;
      RECT  229500.0 269100.0 231300.0 270900.00000000006 ;
      RECT  1500.0 278700.0 3300.0 280500.0 ;
      RECT  9900.0 278700.0 11700.000000000002 280500.0 ;
      RECT  19500.0 278700.0 21300.0 280500.0 ;
      RECT  29100.0 278700.0 30900.000000000004 280500.0 ;
      RECT  38700.0 278700.0 40500.0 280500.0 ;
      RECT  48300.00000000001 278700.0 50100.0 280500.0 ;
      RECT  57900.00000000001 278700.0 59700.0 280500.0 ;
      RECT  86700.0 278700.0 88500.0 280500.0 ;
      RECT  96300.00000000001 278700.0 98100.00000000001 280500.0 ;
      RECT  105900.0 278700.0 107700.0 280500.0 ;
      RECT  115500.00000000001 278700.0 117300.00000000001 280500.0 ;
      RECT  125100.00000000001 278700.0 126900.0 280500.0 ;
      RECT  134700.0 278700.0 136500.0 280500.0 ;
      RECT  144299.99999999997 278700.0 146100.0 280500.0 ;
      RECT  153900.0 278700.0 155700.00000000003 280500.0 ;
      RECT  163500.0 278700.0 165300.0 280500.0 ;
      RECT  173100.0 278700.0 174900.0 280500.0 ;
      RECT  182700.0 278700.0 184500.0 280500.0 ;
      RECT  192300.0 278700.0 194100.00000000003 280500.0 ;
      RECT  201900.0 278700.0 203700.00000000003 280500.0 ;
      RECT  211500.0 278700.0 213300.0 280500.0 ;
      RECT  221100.0 278700.0 222900.0 280500.0 ;
      RECT  229500.0 278700.0 231300.0 280500.0 ;
      RECT  1500.0 288300.0 3300.0 290100.0 ;
      RECT  9900.0 288300.0 11700.000000000002 290100.0 ;
      RECT  19500.0 288300.0 21300.0 290100.0 ;
      RECT  29100.0 288300.0 30900.000000000004 290100.0 ;
      RECT  38700.0 288300.0 40500.0 290100.0 ;
      RECT  48300.00000000001 288300.0 50100.0 290100.0 ;
      RECT  57900.00000000001 288300.0 59700.0 290100.0 ;
      RECT  67500.0 288300.0 69300.0 290100.0 ;
      RECT  77100.00000000001 288300.0 78900.0 290100.0 ;
      RECT  86700.0 288300.0 88500.0 290100.0 ;
      RECT  96300.00000000001 288300.0 98100.00000000001 290100.0 ;
      RECT  105900.0 288300.0 107700.0 290100.0 ;
      RECT  115500.00000000001 288300.0 117300.00000000001 290100.0 ;
      RECT  125100.00000000001 288300.0 126900.0 290100.0 ;
      RECT  134700.0 288300.0 136500.0 290100.0 ;
      RECT  144299.99999999997 288300.0 146100.0 290100.0 ;
      RECT  153900.0 288300.0 155700.00000000003 290100.0 ;
      RECT  163500.0 288300.0 165300.0 290100.0 ;
      RECT  173100.0 288300.0 174900.0 290100.0 ;
      RECT  182700.0 288300.0 184500.0 290100.0 ;
      RECT  192300.0 288300.0 194100.00000000003 290100.0 ;
      RECT  201900.0 288300.0 203700.00000000003 290100.0 ;
      RECT  211500.0 288300.0 213300.0 290100.0 ;
      RECT  221100.0 288300.0 222900.0 290100.0 ;
      RECT  229500.0 288300.0 231300.0 290100.0 ;
      RECT  1500.0 297900.0 3300.0 299700.0 ;
      RECT  9900.0 297900.0 11700.000000000002 299700.0 ;
      RECT  19500.0 297900.0 21300.0 299700.0 ;
      RECT  29100.0 297900.0 30900.000000000004 299700.0 ;
      RECT  38700.0 297900.0 40500.0 299700.0 ;
      RECT  48300.00000000001 297900.0 50100.0 299700.0 ;
      RECT  57900.00000000001 297900.0 59700.0 299700.0 ;
      RECT  67500.0 297900.0 69300.0 299700.0 ;
      RECT  77100.00000000001 297900.0 78900.0 299700.0 ;
      RECT  86700.0 297900.0 88500.0 299700.0 ;
      RECT  96300.00000000001 297900.0 98100.00000000001 299700.0 ;
      RECT  105900.0 297900.0 107700.0 299700.0 ;
      RECT  115500.00000000001 297900.0 117300.00000000001 299700.0 ;
      RECT  125100.00000000001 297900.0 126900.0 299700.0 ;
      RECT  134700.0 297900.0 136500.0 299700.0 ;
      RECT  144299.99999999997 297900.0 146100.0 299700.0 ;
      RECT  153900.0 297900.0 155700.00000000003 299700.0 ;
      RECT  163500.0 297900.0 165300.0 299700.0 ;
      RECT  173100.0 297900.0 174900.0 299700.0 ;
      RECT  182700.0 297900.0 184500.0 299700.0 ;
      RECT  192300.0 297900.0 194100.00000000003 299700.0 ;
      RECT  201900.0 297900.0 203700.00000000003 299700.0 ;
      RECT  211500.0 297900.0 213300.0 299700.0 ;
      RECT  221100.0 297900.0 222900.0 299700.0 ;
      RECT  229500.0 297900.0 231300.0 299700.0 ;
      RECT  5100.000000000001 5100.000000000001 6900.0 6900.0 ;
      RECT  14700.0 5100.000000000001 16500.0 6900.0 ;
      RECT  24300.0 5100.000000000001 26100.0 6900.0 ;
      RECT  33900.00000000001 5100.000000000001 35700.0 6900.0 ;
      RECT  43500.00000000001 5100.000000000001 45300.00000000001 6900.0 ;
      RECT  53100.00000000001 5100.000000000001 54900.00000000001 6900.0 ;
      RECT  62700.0 5100.000000000001 64500.0 6900.0 ;
      RECT  72300.00000000001 5100.000000000001 74100.00000000001 6900.0 ;
      RECT  81900.0 5100.000000000001 83700.0 6900.0 ;
      RECT  91500.00000000001 5100.000000000001 93300.00000000001 6900.0 ;
      RECT  101100.00000000001 5100.000000000001 102900.0 6900.0 ;
      RECT  110700.0 5100.000000000001 112500.0 6900.0 ;
      RECT  120300.00000000001 5100.000000000001 122100.00000000001 6900.0 ;
      RECT  129900.0 5100.000000000001 131700.00000000003 6900.0 ;
      RECT  139500.0 5100.000000000001 141300.0 6900.0 ;
      RECT  149100.0 5100.000000000001 150900.0 6900.0 ;
      RECT  158700.0 5100.000000000001 160500.0 6900.0 ;
      RECT  5100.000000000001 14700.0 6900.0 16500.0 ;
      RECT  14700.0 14700.0 16500.0 16500.0 ;
      RECT  24300.0 14700.0 26100.0 16500.0 ;
      RECT  33900.00000000001 14700.0 35700.0 16500.0 ;
      RECT  43500.00000000001 14700.0 45300.00000000001 16500.0 ;
      RECT  53100.00000000001 14700.0 54900.00000000001 16500.0 ;
      RECT  62700.0 14700.0 64500.0 16500.0 ;
      RECT  72300.00000000001 14700.0 74100.00000000001 16500.0 ;
      RECT  81900.0 14700.0 83700.0 16500.0 ;
      RECT  91500.00000000001 14700.0 93300.00000000001 16500.0 ;
      RECT  101100.00000000001 14700.0 102900.0 16500.0 ;
      RECT  110700.0 14700.0 112500.0 16500.0 ;
      RECT  120300.00000000001 14700.0 122100.00000000001 16500.0 ;
      RECT  129900.0 14700.0 131700.00000000003 16500.0 ;
      RECT  139500.0 14700.0 141300.0 16500.0 ;
      RECT  149100.0 14700.0 150900.0 16500.0 ;
      RECT  158700.0 14700.0 160500.0 16500.0 ;
      RECT  168300.0 14700.0 170100.00000000003 16500.0 ;
      RECT  177900.0 14700.0 179700.00000000003 16500.0 ;
      RECT  187500.0 14700.0 189300.0 16500.0 ;
      RECT  197100.0 14700.0 198900.0 16500.0 ;
      RECT  206700.0 14700.0 208500.0 16500.0 ;
      RECT  216300.0 14700.0 218100.00000000003 16500.0 ;
      RECT  225900.0 14700.0 227700.00000000003 16500.0 ;
      RECT  5100.000000000001 24300.0 6900.0 26100.0 ;
      RECT  14700.0 24300.0 16500.0 26100.0 ;
      RECT  24300.0 24300.0 26100.0 26100.0 ;
      RECT  33900.00000000001 24300.0 35700.0 26100.0 ;
      RECT  43500.00000000001 24300.0 45300.00000000001 26100.0 ;
      RECT  53100.00000000001 24300.0 54900.00000000001 26100.0 ;
      RECT  62700.0 24300.0 64500.0 26100.0 ;
      RECT  72300.00000000001 24300.0 74100.00000000001 26100.0 ;
      RECT  81900.0 24300.0 83700.0 26100.0 ;
      RECT  91500.00000000001 24300.0 93300.00000000001 26100.0 ;
      RECT  101100.00000000001 24300.0 102900.0 26100.0 ;
      RECT  110700.0 24300.0 112500.0 26100.0 ;
      RECT  120300.00000000001 24300.0 122100.00000000001 26100.0 ;
      RECT  129900.0 24300.0 131700.00000000003 26100.0 ;
      RECT  139500.0 24300.0 141300.0 26100.0 ;
      RECT  149100.0 24300.0 150900.0 26100.0 ;
      RECT  158700.0 24300.0 160500.0 26100.0 ;
      RECT  168300.0 24300.0 170100.00000000003 26100.0 ;
      RECT  177900.0 24300.0 179700.00000000003 26100.0 ;
      RECT  187500.0 24300.0 189300.0 26100.0 ;
      RECT  197100.0 24300.0 198900.0 26100.0 ;
      RECT  206700.0 24300.0 208500.0 26100.0 ;
      RECT  216300.0 24300.0 218100.00000000003 26100.0 ;
      RECT  225900.0 24300.0 227700.00000000003 26100.0 ;
      RECT  5100.000000000001 33900.00000000001 6900.0 35700.0 ;
      RECT  14700.0 33900.00000000001 16500.0 35700.0 ;
      RECT  24300.0 33900.00000000001 26100.0 35700.0 ;
      RECT  33900.00000000001 33900.00000000001 35700.0 35700.0 ;
      RECT  43500.00000000001 33900.00000000001 45300.00000000001 35700.0 ;
      RECT  53100.00000000001 33900.00000000001 54900.00000000001 35700.0 ;
      RECT  62700.0 33900.00000000001 64500.0 35700.0 ;
      RECT  72300.00000000001 33900.00000000001 74100.00000000001 35700.0 ;
      RECT  81900.0 33900.00000000001 83700.0 35700.0 ;
      RECT  91500.00000000001 33900.00000000001 93300.00000000001 35700.0 ;
      RECT  101100.00000000001 33900.00000000001 102900.0 35700.0 ;
      RECT  110700.0 33900.00000000001 112500.0 35700.0 ;
      RECT  120300.00000000001 33900.00000000001 122100.00000000001 35700.0 ;
      RECT  129900.0 33900.00000000001 131700.00000000003 35700.0 ;
      RECT  139500.0 33900.00000000001 141300.0 35700.0 ;
      RECT  149100.0 33900.00000000001 150900.0 35700.0 ;
      RECT  158700.0 33900.00000000001 160500.0 35700.0 ;
      RECT  168300.0 33900.00000000001 170100.00000000003 35700.0 ;
      RECT  197100.0 33900.00000000001 198900.0 35700.0 ;
      RECT  206700.0 33900.00000000001 208500.0 35700.0 ;
      RECT  216300.0 33900.00000000001 218100.00000000003 35700.0 ;
      RECT  225900.0 33900.00000000001 227700.00000000003 35700.0 ;
      RECT  5100.000000000001 43500.00000000001 6900.0 45300.00000000001 ;
      RECT  14700.0 43500.00000000001 16500.0 45300.00000000001 ;
      RECT  24300.0 43500.00000000001 26100.0 45300.00000000001 ;
      RECT  33900.00000000001 43500.00000000001 35700.0 45300.00000000001 ;
      RECT  43500.00000000001 43500.00000000001 45300.00000000001 45300.00000000001 ;
      RECT  53100.00000000001 43500.00000000001 54900.00000000001 45300.00000000001 ;
      RECT  62700.0 43500.00000000001 64500.0 45300.00000000001 ;
      RECT  72300.00000000001 43500.00000000001 74100.00000000001 45300.00000000001 ;
      RECT  81900.0 43500.00000000001 83700.0 45300.00000000001 ;
      RECT  91500.00000000001 43500.00000000001 93300.00000000001 45300.00000000001 ;
      RECT  101100.00000000001 43500.00000000001 102900.0 45300.00000000001 ;
      RECT  110700.0 43500.00000000001 112500.0 45300.00000000001 ;
      RECT  120300.00000000001 43500.00000000001 122100.00000000001 45300.00000000001 ;
      RECT  129900.0 43500.00000000001 131700.00000000003 45300.00000000001 ;
      RECT  139500.0 43500.00000000001 141300.0 45300.00000000001 ;
      RECT  149100.0 43500.00000000001 150900.0 45300.00000000001 ;
      RECT  158700.0 43500.00000000001 160500.0 45300.00000000001 ;
      RECT  168300.0 43500.00000000001 170100.00000000003 45300.00000000001 ;
      RECT  198300.0 43500.00000000001 200100.00000000003 45300.00000000001 ;
      RECT  206700.0 43500.00000000001 208500.0 45300.00000000001 ;
      RECT  216300.0 43500.00000000001 218100.00000000003 45300.00000000001 ;
      RECT  225900.0 43500.00000000001 227700.00000000003 45300.00000000001 ;
      RECT  5100.000000000001 53100.00000000001 6900.0 54900.00000000001 ;
      RECT  14700.0 53100.00000000001 16500.0 54900.00000000001 ;
      RECT  24300.0 53100.00000000001 26100.0 54900.00000000001 ;
      RECT  33900.00000000001 53100.00000000001 35700.0 54900.00000000001 ;
      RECT  43500.00000000001 53100.00000000001 45300.00000000001 54900.00000000001 ;
      RECT  53100.00000000001 53100.00000000001 54900.00000000001 54900.00000000001 ;
      RECT  62700.0 53100.00000000001 64500.0 54900.00000000001 ;
      RECT  72300.00000000001 53100.00000000001 74100.00000000001 54900.00000000001 ;
      RECT  81900.0 53100.00000000001 83700.0 54900.00000000001 ;
      RECT  91500.00000000001 53100.00000000001 93300.00000000001 54900.00000000001 ;
      RECT  101100.00000000001 53100.00000000001 102900.0 54900.00000000001 ;
      RECT  110700.0 53100.00000000001 112500.0 54900.00000000001 ;
      RECT  120300.00000000001 53100.00000000001 122100.00000000001 54900.00000000001 ;
      RECT  129900.0 53100.00000000001 131700.00000000003 54900.00000000001 ;
      RECT  139500.0 53100.00000000001 141300.0 54900.00000000001 ;
      RECT  149100.0 53100.00000000001 150900.0 54900.00000000001 ;
      RECT  158700.0 53100.00000000001 160500.0 54900.00000000001 ;
      RECT  168300.0 53100.00000000001 170100.00000000003 54900.00000000001 ;
      RECT  198300.0 53100.00000000001 200100.00000000003 54900.00000000001 ;
      RECT  206700.0 53100.00000000001 208500.0 54900.00000000001 ;
      RECT  216300.0 53100.00000000001 218100.00000000003 54900.00000000001 ;
      RECT  225900.0 53100.00000000001 227700.00000000003 54900.00000000001 ;
      RECT  5100.000000000001 62700.0 6900.0 64500.0 ;
      RECT  14700.0 62700.0 16500.0 64500.0 ;
      RECT  24300.0 62700.0 26100.0 64500.0 ;
      RECT  33900.00000000001 62700.0 35700.0 64500.0 ;
      RECT  43500.00000000001 62700.0 45300.00000000001 64500.0 ;
      RECT  53100.00000000001 62700.0 54900.00000000001 64500.0 ;
      RECT  62700.0 62700.0 64500.0 64500.0 ;
      RECT  72300.00000000001 62700.0 74100.00000000001 64500.0 ;
      RECT  81900.0 62700.0 83700.0 64500.0 ;
      RECT  91500.00000000001 62700.0 93300.00000000001 64500.0 ;
      RECT  101100.00000000001 62700.0 102900.0 64500.0 ;
      RECT  110700.0 62700.0 112500.0 64500.0 ;
      RECT  120300.00000000001 62700.0 122100.00000000001 64500.0 ;
      RECT  129900.0 62700.0 131700.00000000003 64500.0 ;
      RECT  139500.0 62700.0 141300.0 64500.0 ;
      RECT  149100.0 62700.0 150900.0 64500.0 ;
      RECT  158700.0 62700.0 160500.0 64500.0 ;
      RECT  168300.0 62700.0 170100.00000000003 64500.0 ;
      RECT  177900.0 62700.0 179700.00000000003 64500.0 ;
      RECT  187500.0 62700.0 189300.0 64500.0 ;
      RECT  197100.0 62700.0 198900.0 64500.0 ;
      RECT  206700.0 62700.0 208500.0 64500.0 ;
      RECT  216300.0 62700.0 218100.00000000003 64500.0 ;
      RECT  225900.0 62700.0 227700.00000000003 64500.0 ;
      RECT  5100.000000000001 72300.00000000001 6900.0 74100.00000000001 ;
      RECT  14700.0 72300.00000000001 16500.0 74100.00000000001 ;
      RECT  24300.0 72300.00000000001 26100.0 74100.00000000001 ;
      RECT  33900.00000000001 72300.00000000001 35700.0 74100.00000000001 ;
      RECT  43500.00000000001 72300.00000000001 45300.00000000001 74100.00000000001 ;
      RECT  53100.00000000001 72300.00000000001 54900.00000000001 74100.00000000001 ;
      RECT  62700.0 72300.00000000001 64500.0 74100.00000000001 ;
      RECT  72300.00000000001 72300.00000000001 74100.00000000001 74100.00000000001 ;
      RECT  81900.0 72300.00000000001 83700.0 74100.00000000001 ;
      RECT  91500.00000000001 72300.00000000001 93300.00000000001 74100.00000000001 ;
      RECT  101100.00000000001 72300.00000000001 102900.0 74100.00000000001 ;
      RECT  110700.0 72300.00000000001 112500.0 74100.00000000001 ;
      RECT  120300.00000000001 72300.00000000001 122100.00000000001 74100.00000000001 ;
      RECT  129900.0 72300.00000000001 131700.00000000003 74100.00000000001 ;
      RECT  139500.0 72300.00000000001 141300.0 74100.00000000001 ;
      RECT  149100.0 72300.00000000001 150900.0 74100.00000000001 ;
      RECT  158700.0 72300.00000000001 160500.0 74100.00000000001 ;
      RECT  168300.0 72300.00000000001 170100.00000000003 74100.00000000001 ;
      RECT  177900.0 72300.00000000001 179700.00000000003 74100.00000000001 ;
      RECT  187500.0 72300.00000000001 189300.0 74100.00000000001 ;
      RECT  197100.0 72300.00000000001 198900.0 74100.00000000001 ;
      RECT  206700.0 72300.00000000001 208500.0 74100.00000000001 ;
      RECT  216300.0 72300.00000000001 218100.00000000003 74100.00000000001 ;
      RECT  225900.0 72300.00000000001 227700.00000000003 74100.00000000001 ;
      RECT  5100.000000000001 81900.0 6900.0 83700.0 ;
      RECT  14700.0 81900.0 16500.0 83700.0 ;
      RECT  24300.0 81900.0 26100.0 83700.0 ;
      RECT  33900.00000000001 81900.0 35700.0 83700.0 ;
      RECT  43500.00000000001 81900.0 45300.00000000001 83700.0 ;
      RECT  53100.00000000001 81900.0 54900.00000000001 83700.0 ;
      RECT  62700.0 81900.0 64500.0 83700.0 ;
      RECT  72300.00000000001 81900.0 74100.00000000001 83700.0 ;
      RECT  81900.0 81900.0 83700.0 83700.0 ;
      RECT  91500.00000000001 81900.0 93300.00000000001 83700.0 ;
      RECT  101100.00000000001 81900.0 102900.0 83700.0 ;
      RECT  110700.0 81900.0 112500.0 83700.0 ;
      RECT  120300.00000000001 81900.0 122100.00000000001 83700.0 ;
      RECT  129900.0 81900.0 131700.00000000003 83700.0 ;
      RECT  139500.0 81900.0 141300.0 83700.0 ;
      RECT  149100.0 81900.0 150900.0 83700.0 ;
      RECT  158700.0 81900.0 160500.0 83700.0 ;
      RECT  168300.0 81900.0 170100.00000000003 83700.0 ;
      RECT  177900.0 81900.0 179700.00000000003 83700.0 ;
      RECT  187500.0 81900.0 189300.0 83700.0 ;
      RECT  197100.0 81900.0 198900.0 83700.0 ;
      RECT  206700.0 81900.0 208500.0 83700.0 ;
      RECT  216300.0 81900.0 218100.00000000003 83700.0 ;
      RECT  225900.0 81900.0 227700.00000000003 83700.0 ;
      RECT  54300.00000000001 91500.00000000001 56100.0 93300.00000000001 ;
      RECT  62700.0 91500.00000000001 64500.0 93300.00000000001 ;
      RECT  72300.00000000001 91500.00000000001 74100.00000000001 93300.00000000001 ;
      RECT  81900.0 91500.00000000001 83700.0 93300.00000000001 ;
      RECT  91500.00000000001 91500.00000000001 93300.00000000001 93300.00000000001 ;
      RECT  101100.00000000001 91500.00000000001 102900.0 93300.00000000001 ;
      RECT  110700.0 91500.00000000001 112500.0 93300.00000000001 ;
      RECT  120300.00000000001 91500.00000000001 122100.00000000001 93300.00000000001 ;
      RECT  129900.0 91500.00000000001 131700.00000000003 93300.00000000001 ;
      RECT  139500.0 91500.00000000001 141300.0 93300.00000000001 ;
      RECT  149100.0 91500.00000000001 150900.0 93300.00000000001 ;
      RECT  158700.0 91500.00000000001 160500.0 93300.00000000001 ;
      RECT  168300.0 91500.00000000001 170100.00000000003 93300.00000000001 ;
      RECT  176700.0 91500.00000000001 178500.0 93300.00000000001 ;
      RECT  198300.0 91500.00000000001 200100.00000000003 93300.00000000001 ;
      RECT  206700.0 91500.00000000001 208500.0 93300.00000000001 ;
      RECT  216300.0 91500.00000000001 218100.00000000003 93300.00000000001 ;
      RECT  225900.0 91500.00000000001 227700.00000000003 93300.00000000001 ;
      RECT  5100.000000000001 101100.00000000001 6900.0 102900.0 ;
      RECT  14700.0 101100.00000000001 16500.0 102900.0 ;
      RECT  24300.0 101100.00000000001 26100.0 102900.0 ;
      RECT  33900.00000000001 101100.00000000001 35700.0 102900.0 ;
      RECT  43500.00000000001 101100.00000000001 45300.00000000001 102900.0 ;
      RECT  53100.00000000001 101100.00000000001 54900.00000000001 102900.0 ;
      RECT  61500.00000000001 101100.00000000001 63300.00000000001 102900.0 ;
      RECT  81900.0 101100.00000000001 83700.0 102900.0 ;
      RECT  91500.00000000001 101100.00000000001 93300.00000000001 102900.0 ;
      RECT  101100.00000000001 101100.00000000001 102900.0 102900.0 ;
      RECT  110700.0 101100.00000000001 112500.0 102900.0 ;
      RECT  120300.00000000001 101100.00000000001 122100.00000000001 102900.0 ;
      RECT  129900.0 101100.00000000001 131700.00000000003 102900.0 ;
      RECT  139500.0 101100.00000000001 141300.0 102900.0 ;
      RECT  149100.0 101100.00000000001 150900.0 102900.0 ;
      RECT  158700.0 101100.00000000001 160500.0 102900.0 ;
      RECT  168300.0 101100.00000000001 170100.00000000003 102900.0 ;
      RECT  177900.0 101100.00000000001 179700.00000000003 102900.0 ;
      RECT  187500.0 101100.00000000001 189300.0 102900.0 ;
      RECT  197100.0 101100.00000000001 198900.0 102900.0 ;
      RECT  206700.0 101100.00000000001 208500.0 102900.0 ;
      RECT  216300.0 101100.00000000001 218100.00000000003 102900.0 ;
      RECT  225900.0 101100.00000000001 227700.00000000003 102900.0 ;
      RECT  5100.000000000001 110700.0 6900.0 112500.0 ;
      RECT  14700.0 110700.0 16500.0 112500.0 ;
      RECT  24300.0 110700.0 26100.0 112500.0 ;
      RECT  33900.00000000001 110700.0 35700.0 112500.0 ;
      RECT  43500.00000000001 110700.0 45300.00000000001 112500.0 ;
      RECT  53100.00000000001 110700.0 54900.00000000001 112500.0 ;
      RECT  61500.00000000001 110700.0 63300.00000000001 112500.0 ;
      RECT  187500.0 110700.0 189300.0 112500.0 ;
      RECT  197100.0 110700.0 198900.0 112500.0 ;
      RECT  206700.0 110700.0 208500.0 112500.0 ;
      RECT  216300.0 110700.0 218100.00000000003 112500.0 ;
      RECT  225900.0 110700.0 227700.00000000003 112500.0 ;
      RECT  5100.000000000001 120300.00000000001 6900.0 122100.00000000001 ;
      RECT  14700.0 120300.00000000001 16500.0 122100.00000000001 ;
      RECT  24300.0 120300.00000000001 26100.0 122100.00000000001 ;
      RECT  33900.00000000001 120300.00000000001 35700.0 122100.00000000001 ;
      RECT  43500.00000000001 120300.00000000001 45300.00000000001 122100.00000000001 ;
      RECT  53100.00000000001 120300.00000000001 54900.00000000001 122100.00000000001 ;
      RECT  62700.0 120300.00000000001 64500.0 122100.00000000001 ;
      RECT  72300.00000000001 120300.00000000001 74100.00000000001 122100.00000000001 ;
      RECT  80700.0 120300.00000000001 82500.0 122100.00000000001 ;
      RECT  177900.0 120300.00000000001 179700.00000000003 122100.00000000001 ;
      RECT  187500.0 120300.00000000001 189300.0 122100.00000000001 ;
      RECT  197100.0 120300.00000000001 198900.0 122100.00000000001 ;
      RECT  206700.0 120300.00000000001 208500.0 122100.00000000001 ;
      RECT  216300.0 120300.00000000001 218100.00000000003 122100.00000000001 ;
      RECT  225900.0 120300.00000000001 227700.00000000003 122100.00000000001 ;
      RECT  43500.00000000001 129900.0 45300.00000000001 131700.00000000003 ;
      RECT  53100.00000000001 129900.0 54900.00000000001 131700.00000000003 ;
      RECT  62700.0 129900.0 64500.0 131700.00000000003 ;
      RECT  91500.00000000001 129900.0 93300.00000000001 131700.00000000003 ;
      RECT  101100.00000000001 129900.0 102900.0 131700.00000000003 ;
      RECT  121500.00000000001 129900.0 123300.00000000001 131700.00000000003 ;
      RECT  129900.0 129900.0 131700.00000000003 131700.00000000003 ;
      RECT  139500.0 129900.0 141300.0 131700.00000000003 ;
      RECT  149100.0 129900.0 150900.0 131700.00000000003 ;
      RECT  158700.0 129900.0 160500.0 131700.00000000003 ;
      RECT  168300.0 129900.0 170100.00000000003 131700.00000000003 ;
      RECT  177900.0 129900.0 179700.00000000003 131700.00000000003 ;
      RECT  187500.0 129900.0 189300.0 131700.00000000003 ;
      RECT  197100.0 129900.0 198900.0 131700.00000000003 ;
      RECT  206700.0 129900.0 208500.0 131700.00000000003 ;
      RECT  216300.0 129900.0 218100.00000000003 131700.00000000003 ;
      RECT  225900.0 129900.0 227700.00000000003 131700.00000000003 ;
      RECT  43500.00000000001 139500.0 45300.00000000001 141300.0 ;
      RECT  53100.00000000001 139500.0 54900.00000000001 141300.0 ;
      RECT  62700.0 139500.0 64500.0 141300.0 ;
      RECT  177900.0 139500.0 179700.00000000003 141300.0 ;
      RECT  187500.0 139500.0 189300.0 141300.0 ;
      RECT  197100.0 139500.0 198900.0 141300.0 ;
      RECT  206700.0 139500.0 208500.0 141300.0 ;
      RECT  216300.0 139500.0 218100.00000000003 141300.0 ;
      RECT  225900.0 139500.0 227700.00000000003 141300.0 ;
      RECT  44700.0 149100.0 46500.0 150900.0 ;
      RECT  53100.00000000001 149100.0 54900.00000000001 150900.0 ;
      RECT  62700.0 149100.0 64500.0 150900.0 ;
      RECT  72300.00000000001 149100.0 74100.00000000001 150900.0 ;
      RECT  81900.0 149100.0 83700.0 150900.0 ;
      RECT  91500.00000000001 149100.0 93300.00000000001 150900.0 ;
      RECT  101100.00000000001 149100.0 102900.0 150900.0 ;
      RECT  129900.0 149100.0 131700.00000000003 150900.0 ;
      RECT  139500.0 149100.0 141300.0 150900.0 ;
      RECT  149100.0 149100.0 150900.0 150900.0 ;
      RECT  158700.0 149100.0 160500.0 150900.0 ;
      RECT  168300.0 149100.0 170100.00000000003 150900.0 ;
      RECT  177900.0 149100.0 179700.00000000003 150900.0 ;
      RECT  187500.0 149100.0 189300.0 150900.0 ;
      RECT  197100.0 149100.0 198900.0 150900.0 ;
      RECT  206700.0 149100.0 208500.0 150900.0 ;
      RECT  216300.0 149100.0 218100.00000000003 150900.0 ;
      RECT  225900.0 149100.0 227700.00000000003 150900.0 ;
      RECT  43500.00000000001 158700.0 45300.00000000001 160500.0 ;
      RECT  53100.00000000001 158700.0 54900.00000000001 160500.0 ;
      RECT  62700.0 158700.0 64500.0 160500.0 ;
      RECT  72300.00000000001 158700.0 74100.00000000001 160500.0 ;
      RECT  80700.0 158700.0 82500.0 160500.0 ;
      RECT  177900.0 158700.0 179700.00000000003 160500.0 ;
      RECT  187500.0 158700.0 189300.0 160500.0 ;
      RECT  197100.0 158700.0 198900.0 160500.0 ;
      RECT  206700.0 158700.0 208500.0 160500.0 ;
      RECT  216300.0 158700.0 218100.00000000003 160500.0 ;
      RECT  225900.0 158700.0 227700.00000000003 160500.0 ;
      RECT  44700.0 168300.0 46500.0 170100.00000000003 ;
      RECT  53100.00000000001 168300.0 54900.00000000001 170100.00000000003 ;
      RECT  62700.0 168300.0 64500.0 170100.00000000003 ;
      RECT  91500.00000000001 168300.0 93300.00000000001 170100.00000000003 ;
      RECT  101100.00000000001 168300.0 102900.0 170100.00000000003 ;
      RECT  129900.0 168300.0 131700.00000000003 170100.00000000003 ;
      RECT  139500.0 168300.0 141300.0 170100.00000000003 ;
      RECT  149100.0 168300.0 150900.0 170100.00000000003 ;
      RECT  158700.0 168300.0 160500.0 170100.00000000003 ;
      RECT  168300.0 168300.0 170100.00000000003 170100.00000000003 ;
      RECT  177900.0 168300.0 179700.00000000003 170100.00000000003 ;
      RECT  187500.0 168300.0 189300.0 170100.00000000003 ;
      RECT  197100.0 168300.0 198900.0 170100.00000000003 ;
      RECT  206700.0 168300.0 208500.0 170100.00000000003 ;
      RECT  216300.0 168300.0 218100.00000000003 170100.00000000003 ;
      RECT  225900.0 168300.0 227700.00000000003 170100.00000000003 ;
      RECT  5100.000000000001 177900.0 6900.0 179700.00000000003 ;
      RECT  14700.0 177900.0 16500.0 179700.00000000003 ;
      RECT  24300.0 177900.0 26100.0 179700.00000000003 ;
      RECT  33900.00000000001 177900.0 35700.0 179700.00000000003 ;
      RECT  43500.00000000001 177900.0 45300.00000000001 179700.00000000003 ;
      RECT  53100.00000000001 177900.0 54900.00000000001 179700.00000000003 ;
      RECT  62700.0 177900.0 64500.0 179700.00000000003 ;
      RECT  177900.0 177900.0 179700.00000000003 179700.00000000003 ;
      RECT  187500.0 177900.0 189300.0 179700.00000000003 ;
      RECT  197100.0 177900.0 198900.0 179700.00000000003 ;
      RECT  206700.0 177900.0 208500.0 179700.00000000003 ;
      RECT  216300.0 177900.0 218100.00000000003 179700.00000000003 ;
      RECT  225900.0 177900.0 227700.00000000003 179700.00000000003 ;
      RECT  5100.000000000001 187500.0 6900.0 189300.0 ;
      RECT  14700.0 187500.0 16500.0 189300.0 ;
      RECT  24300.0 187500.0 26100.0 189300.0 ;
      RECT  44700.0 187500.0 46500.0 189300.0 ;
      RECT  53100.00000000001 187500.0 54900.00000000001 189300.0 ;
      RECT  62700.0 187500.0 64500.0 189300.0 ;
      RECT  72300.00000000001 187500.0 74100.00000000001 189300.0 ;
      RECT  81900.0 187500.0 83700.0 189300.0 ;
      RECT  91500.00000000001 187500.0 93300.00000000001 189300.0 ;
      RECT  101100.00000000001 187500.0 102900.0 189300.0 ;
      RECT  131100.0 187500.0 132900.0 189300.0 ;
      RECT  139500.0 187500.0 141300.0 189300.0 ;
      RECT  149100.0 187500.0 150900.0 189300.0 ;
      RECT  158700.0 187500.0 160500.0 189300.0 ;
      RECT  168300.0 187500.0 170100.00000000003 189300.0 ;
      RECT  198300.0 187500.0 200100.00000000003 189300.0 ;
      RECT  206700.0 187500.0 208500.0 189300.0 ;
      RECT  216300.0 187500.0 218100.00000000003 189300.0 ;
      RECT  225900.0 187500.0 227700.00000000003 189300.0 ;
      RECT  5100.000000000001 197100.0 6900.0 198900.0 ;
      RECT  14700.0 197100.0 16500.0 198900.0 ;
      RECT  24300.0 197100.0 26100.0 198900.0 ;
      RECT  33900.00000000001 197100.0 35700.0 198900.0 ;
      RECT  43500.00000000001 197100.0 45300.00000000001 198900.0 ;
      RECT  53100.00000000001 197100.0 54900.00000000001 198900.0 ;
      RECT  62700.0 197100.0 64500.0 198900.0 ;
      RECT  72300.00000000001 197100.0 74100.00000000001 198900.0 ;
      RECT  80700.0 197100.0 82500.0 198900.0 ;
      RECT  198300.0 197100.0 200100.00000000003 198900.0 ;
      RECT  206700.0 197100.0 208500.0 198900.0 ;
      RECT  216300.0 197100.0 218100.00000000003 198900.0 ;
      RECT  225900.0 197100.0 227700.00000000003 198900.0 ;
      RECT  5100.000000000001 206700.0 6900.0 208500.0 ;
      RECT  14700.0 206700.0 16500.0 208500.0 ;
      RECT  24300.0 206700.0 26100.0 208500.0 ;
      RECT  44700.0 206700.0 46500.0 208500.0 ;
      RECT  53100.00000000001 206700.0 54900.00000000001 208500.0 ;
      RECT  62700.0 206700.0 64500.0 208500.0 ;
      RECT  72300.00000000001 206700.0 74100.00000000001 208500.0 ;
      RECT  81900.0 206700.0 83700.0 208500.0 ;
      RECT  91500.00000000001 206700.0 93300.00000000001 208500.0 ;
      RECT  101100.00000000001 206700.0 102900.0 208500.0 ;
      RECT  110700.0 206700.0 112500.0 208500.0 ;
      RECT  120300.00000000001 206700.0 122100.00000000001 208500.0 ;
      RECT  129900.0 206700.0 131700.00000000003 208500.0 ;
      RECT  139500.0 206700.0 141300.0 208500.0 ;
      RECT  149100.0 206700.0 150900.0 208500.0 ;
      RECT  158700.0 206700.0 160500.0 208500.0 ;
      RECT  168300.0 206700.0 170100.00000000003 208500.0 ;
      RECT  198300.0 206700.0 200100.00000000003 208500.0 ;
      RECT  206700.0 206700.0 208500.0 208500.0 ;
      RECT  216300.0 206700.0 218100.00000000003 208500.0 ;
      RECT  225900.0 206700.0 227700.00000000003 208500.0 ;
      RECT  5100.000000000001 216300.0 6900.0 218100.00000000003 ;
      RECT  14700.0 216300.0 16500.0 218100.00000000003 ;
      RECT  24300.0 216300.0 26100.0 218100.00000000003 ;
      RECT  33900.00000000001 216300.0 35700.0 218100.00000000003 ;
      RECT  81900.0 216300.0 83700.0 218100.00000000003 ;
      RECT  91500.00000000001 216300.0 93300.00000000001 218100.00000000003 ;
      RECT  101100.00000000001 216300.0 102900.0 218100.00000000003 ;
      RECT  110700.0 216300.0 112500.0 218100.00000000003 ;
      RECT  120300.00000000001 216300.0 122100.00000000001 218100.00000000003 ;
      RECT  198300.0 216300.0 200100.00000000003 218100.00000000003 ;
      RECT  206700.0 216300.0 208500.0 218100.00000000003 ;
      RECT  216300.0 216300.0 218100.00000000003 218100.00000000003 ;
      RECT  225900.0 216300.0 227700.00000000003 218100.00000000003 ;
      RECT  5100.000000000001 225900.0 6900.0 227700.00000000003 ;
      RECT  14700.0 225900.0 16500.0 227700.00000000003 ;
      RECT  24300.0 225900.0 26100.0 227700.00000000003 ;
      RECT  33900.00000000001 225900.0 35700.0 227700.00000000003 ;
      RECT  43500.00000000001 225900.0 45300.00000000001 227700.00000000003 ;
      RECT  53100.00000000001 225900.0 54900.00000000001 227700.00000000003 ;
      RECT  62700.0 225900.0 64500.0 227700.00000000003 ;
      RECT  72300.00000000001 225900.0 74100.00000000001 227700.00000000003 ;
      RECT  81900.0 225900.0 83700.0 227700.00000000003 ;
      RECT  91500.00000000001 225900.0 93300.00000000001 227700.00000000003 ;
      RECT  101100.00000000001 225900.0 102900.0 227700.00000000003 ;
      RECT  110700.0 225900.0 112500.0 227700.00000000003 ;
      RECT  120300.00000000001 225900.0 122100.00000000001 227700.00000000003 ;
      RECT  129900.0 225900.0 131700.00000000003 227700.00000000003 ;
      RECT  139500.0 225900.0 141300.0 227700.00000000003 ;
      RECT  149100.0 225900.0 150900.0 227700.00000000003 ;
      RECT  158700.0 225900.0 160500.0 227700.00000000003 ;
      RECT  168300.0 225900.0 170100.00000000003 227700.00000000003 ;
      RECT  198300.0 225900.0 200100.00000000003 227700.00000000003 ;
      RECT  206700.0 225900.0 208500.0 227700.00000000003 ;
      RECT  216300.0 225900.0 218100.00000000003 227700.00000000003 ;
      RECT  225900.0 225900.0 227700.00000000003 227700.00000000003 ;
      RECT  5100.000000000001 235500.0 6900.0 237300.0 ;
      RECT  14700.0 235500.0 16500.0 237300.0 ;
      RECT  24300.0 235500.0 26100.0 237300.0 ;
      RECT  33900.00000000001 235500.0 35700.0 237300.0 ;
      RECT  43500.00000000001 235500.0 45300.00000000001 237300.0 ;
      RECT  53100.00000000001 235500.0 54900.00000000001 237300.0 ;
      RECT  62700.0 235500.0 64500.0 237300.0 ;
      RECT  72300.00000000001 235500.0 74100.00000000001 237300.0 ;
      RECT  81900.0 235500.0 83700.0 237300.0 ;
      RECT  91500.00000000001 235500.0 93300.00000000001 237300.0 ;
      RECT  101100.00000000001 235500.0 102900.0 237300.0 ;
      RECT  110700.0 235500.0 112500.0 237300.0 ;
      RECT  120300.00000000001 235500.0 122100.00000000001 237300.0 ;
      RECT  129900.0 235500.0 131700.00000000003 237300.0 ;
      RECT  139500.0 235500.0 141300.0 237300.0 ;
      RECT  149100.0 235500.0 150900.0 237300.0 ;
      RECT  158700.0 235500.0 160500.0 237300.0 ;
      RECT  168300.0 235500.0 170100.00000000003 237300.0 ;
      RECT  198300.0 235500.0 200100.00000000003 237300.0 ;
      RECT  206700.0 235500.0 208500.0 237300.0 ;
      RECT  216300.0 235500.0 218100.00000000003 237300.0 ;
      RECT  225900.0 235500.0 227700.00000000003 237300.0 ;
      RECT  5100.000000000001 245100.0 6900.0 246900.0 ;
      RECT  14700.0 245100.0 16500.0 246900.0 ;
      RECT  24300.0 245100.0 26100.0 246900.0 ;
      RECT  33900.00000000001 245100.0 35700.0 246900.0 ;
      RECT  43500.00000000001 245100.0 45300.00000000001 246900.0 ;
      RECT  53100.00000000001 245100.0 54900.00000000001 246900.0 ;
      RECT  62700.0 245100.0 64500.0 246900.0 ;
      RECT  72300.00000000001 245100.0 74100.00000000001 246900.0 ;
      RECT  81900.0 245100.0 83700.0 246900.0 ;
      RECT  91500.00000000001 245100.0 93300.00000000001 246900.0 ;
      RECT  101100.00000000001 245100.0 102900.0 246900.0 ;
      RECT  110700.0 245100.0 112500.0 246900.0 ;
      RECT  120300.00000000001 245100.0 122100.00000000001 246900.0 ;
      RECT  129900.0 245100.0 131700.00000000003 246900.0 ;
      RECT  139500.0 245100.0 141300.0 246900.0 ;
      RECT  149100.0 245100.0 150900.0 246900.0 ;
      RECT  158700.0 245100.0 160500.0 246900.0 ;
      RECT  168300.0 245100.0 170100.00000000003 246900.0 ;
      RECT  198300.0 245100.0 200100.00000000003 246900.0 ;
      RECT  206700.0 245100.0 208500.0 246900.0 ;
      RECT  216300.0 245100.0 218100.00000000003 246900.0 ;
      RECT  225900.0 245100.0 227700.00000000003 246900.0 ;
      RECT  5100.000000000001 254700.0 6900.0 256500.0 ;
      RECT  14700.0 254700.0 16500.0 256500.0 ;
      RECT  24300.0 254700.0 26100.0 256500.0 ;
      RECT  33900.00000000001 254700.0 35700.0 256500.0 ;
      RECT  43500.00000000001 254700.0 45300.00000000001 256500.0 ;
      RECT  53100.00000000001 254700.0 54900.00000000001 256500.0 ;
      RECT  62700.0 254700.0 64500.0 256500.0 ;
      RECT  72300.00000000001 254700.0 74100.00000000001 256500.0 ;
      RECT  81900.0 254700.0 83700.0 256500.0 ;
      RECT  91500.00000000001 254700.0 93300.00000000001 256500.0 ;
      RECT  101100.00000000001 254700.0 102900.0 256500.0 ;
      RECT  110700.0 254700.0 112500.0 256500.0 ;
      RECT  120300.00000000001 254700.0 122100.00000000001 256500.0 ;
      RECT  129900.0 254700.0 131700.00000000003 256500.0 ;
      RECT  139500.0 254700.0 141300.0 256500.0 ;
      RECT  149100.0 254700.0 150900.0 256500.0 ;
      RECT  158700.0 254700.0 160500.0 256500.0 ;
      RECT  168300.0 254700.0 170100.00000000003 256500.0 ;
      RECT  198300.0 254700.0 200100.00000000003 256500.0 ;
      RECT  206700.0 254700.0 208500.0 256500.0 ;
      RECT  216300.0 254700.0 218100.00000000003 256500.0 ;
      RECT  225900.0 254700.0 227700.00000000003 256500.0 ;
      RECT  5100.000000000001 264300.0 6900.0 266100.0 ;
      RECT  14700.0 264300.0 16500.0 266100.0 ;
      RECT  24300.0 264300.0 26100.0 266100.0 ;
      RECT  33900.00000000001 264300.0 35700.0 266100.0 ;
      RECT  43500.00000000001 264300.0 45300.00000000001 266100.0 ;
      RECT  53100.00000000001 264300.0 54900.00000000001 266100.0 ;
      RECT  62700.0 264300.0 64500.0 266100.0 ;
      RECT  72300.00000000001 264300.0 74100.00000000001 266100.0 ;
      RECT  81900.0 264300.0 83700.0 266100.0 ;
      RECT  91500.00000000001 264300.0 93300.00000000001 266100.0 ;
      RECT  101100.00000000001 264300.0 102900.0 266100.0 ;
      RECT  110700.0 264300.0 112500.0 266100.0 ;
      RECT  120300.00000000001 264300.0 122100.00000000001 266100.0 ;
      RECT  129900.0 264300.0 131700.00000000003 266100.0 ;
      RECT  139500.0 264300.0 141300.0 266100.0 ;
      RECT  149100.0 264300.0 150900.0 266100.0 ;
      RECT  158700.0 264300.0 160500.0 266100.0 ;
      RECT  168300.0 264300.0 170100.00000000003 266100.0 ;
      RECT  198300.0 264300.0 200100.00000000003 266100.0 ;
      RECT  206700.0 264300.0 208500.0 266100.0 ;
      RECT  216300.0 264300.0 218100.00000000003 266100.0 ;
      RECT  225900.0 264300.0 227700.00000000003 266100.0 ;
      RECT  5100.000000000001 273900.0 6900.0 275700.0 ;
      RECT  14700.0 273900.0 16500.0 275700.0 ;
      RECT  24300.0 273900.0 26100.0 275700.0 ;
      RECT  33900.00000000001 273900.0 35700.0 275700.0 ;
      RECT  43500.00000000001 273900.0 45300.00000000001 275700.0 ;
      RECT  53100.00000000001 273900.0 54900.00000000001 275700.0 ;
      RECT  62700.0 273900.0 64500.0 275700.0 ;
      RECT  72300.00000000001 273900.0 74100.00000000001 275700.0 ;
      RECT  81900.0 273900.0 83700.0 275700.0 ;
      RECT  91500.00000000001 273900.0 93300.00000000001 275700.0 ;
      RECT  101100.00000000001 273900.0 102900.0 275700.0 ;
      RECT  110700.0 273900.0 112500.0 275700.0 ;
      RECT  120300.00000000001 273900.0 122100.00000000001 275700.0 ;
      RECT  129900.0 273900.0 131700.00000000003 275700.0 ;
      RECT  139500.0 273900.0 141300.0 275700.0 ;
      RECT  149100.0 273900.0 150900.0 275700.0 ;
      RECT  158700.0 273900.0 160500.0 275700.0 ;
      RECT  168300.0 273900.0 170100.00000000003 275700.0 ;
      RECT  177900.0 273900.0 179700.00000000003 275700.0 ;
      RECT  187500.0 273900.0 189300.0 275700.0 ;
      RECT  197100.0 273900.0 198900.0 275700.0 ;
      RECT  206700.0 273900.0 208500.0 275700.0 ;
      RECT  216300.0 273900.0 218100.00000000003 275700.0 ;
      RECT  225900.0 273900.0 227700.00000000003 275700.0 ;
      RECT  5100.000000000001 283500.0 6900.0 285300.0 ;
      RECT  14700.0 283500.0 16500.0 285300.0 ;
      RECT  24300.0 283500.0 26100.0 285300.0 ;
      RECT  33900.00000000001 283500.0 35700.0 285300.0 ;
      RECT  43500.00000000001 283500.0 45300.00000000001 285300.0 ;
      RECT  53100.00000000001 283500.0 54900.00000000001 285300.0 ;
      RECT  91500.00000000001 283500.0 93300.00000000001 285300.0 ;
      RECT  101100.00000000001 283500.0 102900.0 285300.0 ;
      RECT  110700.0 283500.0 112500.0 285300.0 ;
      RECT  120300.00000000001 283500.0 122100.00000000001 285300.0 ;
      RECT  129900.0 283500.0 131700.00000000003 285300.0 ;
      RECT  139500.0 283500.0 141300.0 285300.0 ;
      RECT  149100.0 283500.0 150900.0 285300.0 ;
      RECT  158700.0 283500.0 160500.0 285300.0 ;
      RECT  168300.0 283500.0 170100.00000000003 285300.0 ;
      RECT  177900.0 283500.0 179700.00000000003 285300.0 ;
      RECT  187500.0 283500.0 189300.0 285300.0 ;
      RECT  197100.0 283500.0 198900.0 285300.0 ;
      RECT  206700.0 283500.0 208500.0 285300.0 ;
      RECT  216300.0 283500.0 218100.00000000003 285300.0 ;
      RECT  225900.0 283500.0 227700.00000000003 285300.0 ;
      RECT  5100.000000000001 293100.0 6900.0 294900.00000000006 ;
      RECT  14700.0 293100.0 16500.0 294900.00000000006 ;
      RECT  24300.0 293100.0 26100.0 294900.00000000006 ;
      RECT  33900.00000000001 293100.0 35700.0 294900.00000000006 ;
      RECT  43500.00000000001 293100.0 45300.00000000001 294900.00000000006 ;
      RECT  51900.00000000001 293100.0 53700.0 294900.00000000006 ;
      RECT  72300.00000000001 293100.0 74100.00000000001 294900.00000000006 ;
      RECT  81900.0 293100.0 83700.0 294900.00000000006 ;
      RECT  91500.00000000001 293100.0 93300.00000000001 294900.00000000006 ;
      RECT  101100.00000000001 293100.0 102900.0 294900.00000000006 ;
      RECT  110700.0 293100.0 112500.0 294900.00000000006 ;
      RECT  120300.00000000001 293100.0 122100.00000000001 294900.00000000006 ;
      RECT  129900.0 293100.0 131700.00000000003 294900.00000000006 ;
      RECT  139500.0 293100.0 141300.0 294900.00000000006 ;
      RECT  149100.0 293100.0 150900.0 294900.00000000006 ;
      RECT  158700.0 293100.0 160500.0 294900.00000000006 ;
      RECT  168300.0 293100.0 170100.00000000003 294900.00000000006 ;
      RECT  177900.0 293100.0 179700.00000000003 294900.00000000006 ;
      RECT  187500.0 293100.0 189300.0 294900.00000000006 ;
      RECT  197100.0 293100.0 198900.0 294900.00000000006 ;
      RECT  206700.0 293100.0 208500.0 294900.00000000006 ;
      RECT  216300.0 293100.0 218100.00000000003 294900.00000000006 ;
      RECT  225900.0 293100.0 227700.00000000003 294900.00000000006 ;
      RECT  17200.000000000004 160400.0 16400.000000000004 161200.00000000003 ;
      RECT  17200.000000000004 129199.99999999999 16400.000000000004 130000.0 ;
      RECT  14800.0 141200.0 14000.0 142000.0 ;
      RECT  17200.000000000004 141200.0 16400.000000000004 142000.0 ;
      RECT  14800.0 160400.0 14000.0 161200.00000000003 ;
      RECT  190000.00000000003 186800.0 189200.00000000003 187600.00000000003 ;
      RECT  180400.00000000003 206000.0 179600.00000000003 206800.0 ;
      RECT  180400.00000000003 222800.0 179600.00000000003 223600.00000000003 ;
      RECT  34000.0 141200.0 33200.0 142000.0 ;
      RECT  180400.00000000003 30800.0 179600.00000000003 31600.0 ;
      RECT  190000.00000000003 47600.00000000001 189200.00000000003 48400.00000000001 ;
      RECT  190000.00000000003 30800.0 189200.00000000003 31600.0 ;
      RECT  180400.00000000003 47600.00000000001 179600.00000000003 48400.00000000001 ;
      RECT  34000.0 160400.0 33200.0 161200.00000000003 ;
      RECT  190000.00000000003 242000.0 189200.00000000003 242800.0 ;
      RECT  190000.00000000003 206000.0 189200.00000000003 206800.0 ;
      RECT  180400.00000000003 261200.0 179600.00000000003 262000.0 ;
      RECT  190000.00000000003 261200.0 189200.00000000003 262000.0 ;
      RECT  180400.00000000003 242000.0 179600.00000000003 242800.0 ;
      RECT  190000.00000000003 222800.0 189200.00000000003 223600.00000000003 ;
      RECT  180400.00000000003 186800.0 179600.00000000003 187600.00000000003 ;
      RECT  29200.000000000004 129199.99999999999 28400.000000000004 130000.0 ;
      RECT  192400.00000000003 -400.00000000000006 191600.00000000003 399.9999999999999 ;
      RECT  60400.0 210800.0 59600.0 211600.00000000003 ;
      RECT  19600.0 153200.0 18800.0 154000.0 ;
      RECT  12400.000000000002 134000.0 11600.000000000002 134800.0 ;
      RECT  19600.0 134000.0 18800.0 134800.0 ;
      RECT  12400.000000000002 150799.99999999997 11600.000000000002 151600.0 ;
      RECT  211600.00000000003 -400.00000000000006 210800.0 399.9999999999999 ;
      RECT  192400.00000000003 198800.0 191600.00000000003 199600.00000000003 ;
      RECT  185200.00000000003 237200.0 184400.0 238000.0 ;
      RECT  192400.00000000003 256399.99999999997 191600.00000000003 257200.0 ;
      RECT  192400.00000000003 237200.0 191600.00000000003 238000.0 ;
      RECT  185200.00000000003 201200.0 184400.0 202000.0 ;
      RECT  185200.00000000003 263600.0 184400.0 264400.00000000006 ;
      RECT  182800.0 237200.0 182000.0 238000.0 ;
      RECT  175600.00000000003 220400.0 174800.0 221200.00000000003 ;
      RECT  185200.00000000003 220400.0 184400.0 221200.00000000003 ;
      RECT  29200.000000000004 148400.0 28400.000000000004 149200.00000000003 ;
      RECT  185200.00000000003 256399.99999999997 184400.0 257200.0 ;
      RECT  29200.000000000004 165200.0 28400.000000000004 166000.0 ;
      RECT  182800.0 198800.0 182000.0 199600.00000000003 ;
      RECT  192400.00000000003 218000.0 191600.00000000003 218800.0 ;
   END
   END    sram_2_16_scn4m_subm
END    LIBRARY
