magic
tech gf180mcuD
magscale 1 10
timestamp 1694471735
<< nwell >>
rect 0 674 620 1392
<< nmos >>
rect 220 210 280 380
rect 330 210 390 380
<< pmos >>
rect 190 764 250 1104
rect 360 764 420 1104
<< ndiff >>
rect 120 318 220 380
rect 120 272 142 318
rect 188 272 220 318
rect 120 210 220 272
rect 280 210 330 380
rect 390 318 490 380
rect 390 272 422 318
rect 468 272 490 318
rect 390 210 490 272
<< pdiff >>
rect 90 1051 190 1104
rect 90 817 112 1051
rect 158 817 190 1051
rect 90 764 190 817
rect 250 1051 360 1104
rect 250 817 282 1051
rect 328 817 360 1051
rect 250 764 360 817
rect 420 1051 520 1104
rect 420 817 452 1051
rect 498 817 520 1051
rect 420 764 520 817
<< ndiffc >>
rect 142 272 188 318
rect 422 272 468 318
<< pdiffc >>
rect 112 817 158 1051
rect 282 817 328 1051
rect 452 817 498 1051
<< psubdiff >>
rect 540 159 620 180
rect 540 113 557 159
rect 603 113 620 159
rect 540 73 620 113
<< nsubdiff >>
rect 436 1233 543 1250
rect 436 1187 473 1233
rect 519 1187 543 1233
rect 436 1170 543 1187
<< psubdiffcont >>
rect 557 113 603 159
<< nsubdiffcont >>
rect 473 1187 519 1233
<< polysilicon >>
rect 190 1104 250 1154
rect 360 1104 420 1154
rect 190 470 250 764
rect 360 470 420 764
rect 190 430 280 470
rect 220 380 280 430
rect 330 430 420 470
rect 330 380 390 430
rect 220 170 280 210
rect 180 149 280 170
rect 180 103 207 149
rect 253 103 280 149
rect 180 87 280 103
rect 330 170 390 210
rect 330 149 430 170
rect 330 103 346 149
rect 392 103 430 149
rect 330 87 430 103
<< polycontact >>
rect 207 103 253 149
rect 346 103 392 149
<< metal1 >>
rect 470 1236 522 1248
rect 112 1164 330 1210
rect 112 1051 158 1062
rect 280 1051 330 1164
rect 470 1137 522 1184
rect 158 966 164 978
rect 158 902 164 914
rect 112 806 158 817
rect 280 817 282 1051
rect 328 817 330 1051
rect 452 1051 498 1062
rect 446 966 452 978
rect 446 902 452 914
rect 280 450 330 817
rect 452 806 498 817
rect 140 400 330 450
rect 140 318 190 400
rect 140 272 142 318
rect 188 272 190 318
rect 140 210 190 272
rect 422 324 480 347
rect 474 272 480 324
rect 422 240 480 272
rect 544 162 614 178
rect 155 149 267 152
rect 155 103 207 149
rect 253 103 267 149
rect 155 100 267 103
rect 332 149 451 152
rect 332 103 346 149
rect 392 103 451 149
rect 332 100 451 103
rect 544 110 554 162
rect 606 110 614 162
rect 544 79 614 110
<< via1 >>
rect 470 1233 522 1236
rect 470 1187 473 1233
rect 473 1187 519 1233
rect 519 1187 522 1233
rect 470 1184 522 1187
rect 112 914 158 966
rect 158 914 164 966
rect 446 914 452 966
rect 452 914 498 966
rect 422 318 474 324
rect 422 272 468 318
rect 468 272 474 318
rect 554 159 606 162
rect 554 113 557 159
rect 557 113 603 159
rect 603 113 606 159
rect 554 110 606 113
<< metal2 >>
rect 468 1236 524 1248
rect 468 1184 470 1236
rect 522 1184 524 1236
rect 468 968 524 1184
rect 60 966 572 968
rect 60 914 112 966
rect 164 914 446 966
rect 498 914 572 966
rect 60 912 572 914
rect 60 324 608 326
rect 60 272 422 324
rect 474 272 608 324
rect 60 270 608 272
rect 552 162 608 270
rect 552 110 554 162
rect 606 110 608 162
rect 552 88 608 110
<< labels >>
rlabel metal1 s 230 126 230 126 4 B
rlabel metal1 s 369 126 369 126 4 A
rlabel metal1 s 135 1187 135 1187 4 Y
rlabel metal2 s 547 940 547 940 4 VDD
rlabel metal2 s 524 298 524 298 4 GND
<< properties >>
string FIXED_BBOX 0 0 620 1392
<< end >>
