magic
tech sky130A
magscale 1 2
timestamp 1595931502
<< checkpaint >>
rect -1260 -1286 2166 1652
<< scnmos >>
rect 60 0 90 336
rect 168 0 198 336
rect 276 0 306 336
rect 384 0 414 336
rect 492 0 522 336
rect 600 0 630 336
rect 708 0 738 336
rect 816 0 846 336
<< ndiff >>
rect 0 0 60 336
rect 90 0 168 336
rect 198 0 276 336
rect 306 0 384 336
rect 414 0 492 336
rect 522 0 600 336
rect 630 0 708 336
rect 738 0 816 336
rect 846 0 906 336
<< poly >>
rect 60 362 846 392
rect 60 336 90 362
rect 168 336 198 362
rect 276 336 306 362
rect 384 336 414 362
rect 492 336 522 362
rect 600 336 630 362
rect 708 336 738 362
rect 816 336 846 362
rect 60 -26 90 0
rect 168 -26 198 0
rect 276 -26 306 0
rect 384 -26 414 0
rect 492 -26 522 0
rect 600 -26 630 0
rect 708 -26 738 0
rect 816 -26 846 0
<< locali >>
rect 112 235 794 269
rect 8 135 42 201
rect 112 168 146 235
rect 220 135 254 201
rect 328 168 362 235
rect 436 135 470 201
rect 544 168 578 235
rect 652 135 686 201
rect 760 168 794 235
rect 864 135 898 201
use contact_17  contact_17_8
timestamp 1595931502
transform 1 0 0 0 1 135
box 0 0 50 66
use contact_17  contact_17_7
timestamp 1595931502
transform 1 0 104 0 1 135
box 0 0 50 66
use contact_17  contact_17_6
timestamp 1595931502
transform 1 0 212 0 1 135
box 0 0 50 66
use contact_17  contact_17_5
timestamp 1595931502
transform 1 0 320 0 1 135
box 0 0 50 66
use contact_17  contact_17_4
timestamp 1595931502
transform 1 0 428 0 1 135
box 0 0 50 66
use contact_17  contact_17_3
timestamp 1595931502
transform 1 0 536 0 1 135
box 0 0 50 66
use contact_17  contact_17_2
timestamp 1595931502
transform 1 0 644 0 1 135
box 0 0 50 66
use contact_17  contact_17_1
timestamp 1595931502
transform 1 0 752 0 1 135
box 0 0 50 66
use contact_17  contact_17_0
timestamp 1595931502
transform 1 0 856 0 1 135
box 0 0 50 66
<< labels >>
rlabel poly s 453 377 453 377 4 G
rlabel corelocali s 669 168 669 168 4 S
rlabel corelocali s 881 168 881 168 4 S
rlabel corelocali s 453 168 453 168 4 S
rlabel corelocali s 237 168 237 168 4 S
rlabel corelocali s 25 168 25 168 4 S
rlabel corelocali s 453 252 453 252 4 D
<< properties >>
string FIXED_BBOX -25 -26 931 362
<< end >>
