VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_2_16_1_scn4m_subm
   CLASS BLOCK ;
   SIZE 213.0 BY 424.8 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  108.8 11.4 109.6 12.2 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  130.6 11.4 131.4 12.2 ;
      END
   END din0[1]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  65.2 353.4 66.0 354.2 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  65.2 375.4 66.0 376.2 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  65.2 393.4 66.0 394.2 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  65.2 415.4 66.0 416.2 ;
      END
   END addr0[3]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  10.0 11.4 10.8 12.2 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  10.0 33.4 10.8 34.2 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal2 ;
         RECT  54.1 12.3 54.7 12.9 ;
      END
   END clk0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal2 ;
         RECT  189.3 112.6 190.1 115.6 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal2 ;
         RECT  196.1 112.6 196.9 115.6 ;
      END
   END dout0[1]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  81.6 81.6 188.4 82.8 ;
         LAYER metal3 ;
         RECT  152.0 196.4 152.8 197.2 ;
         LAYER metal4 ;
         RECT  136.8 2.4 138.0 423.6 ;
         LAYER metal3 ;
         RECT  60.0 124.8 210.0 126.0 ;
         LAYER metal3 ;
         RECT  0.0 216.0 121.2 217.2 ;
         LAYER metal3 ;
         RECT  0.0 369.6 210.0 370.8 ;
         LAYER metal3 ;
         RECT  0.0 14.4 27.6 15.6 ;
         LAYER metal3 ;
         RECT  177.6 355.2 205.2 356.4 ;
         LAYER metal3 ;
         RECT  198.7 91.4 199.5 92.2 ;
         LAYER metal3 ;
         RECT  133.5 22.4 134.3 23.2 ;
         LAYER metal3 ;
         RECT  170.4 153.6 210.0 154.8 ;
         LAYER metal3 ;
         RECT  0.0 220.8 116.4 222.0 ;
         LAYER metal3 ;
         RECT  200.9 125.4 201.7 126.2 ;
         LAYER metal3 ;
         RECT  0.0 278.4 121.2 279.6 ;
         LAYER metal3 ;
         RECT  23.2 224.0 24.0 224.8 ;
         LAYER metal3 ;
         RECT  33.6 254.4 116.4 255.6 ;
         LAYER metal4 ;
         RECT  50.4 2.4 51.6 423.6 ;
         LAYER metal3 ;
         RECT  136.8 259.2 210.0 260.4 ;
         LAYER metal3 ;
         RECT  23.2 341.6 24.0 342.4 ;
         LAYER metal4 ;
         RECT  31.2 2.4 32.4 423.6 ;
         LAYER metal3 ;
         RECT  205.3 342.0 206.1 342.8 ;
         LAYER metal4 ;
         RECT  12.0 2.4 13.2 423.6 ;
         LAYER metal3 ;
         RECT  148.8 4.8 210.0 6.0 ;
         LAYER metal3 ;
         RECT  0.0 384.0 63.6 385.2 ;
         LAYER metal4 ;
         RECT  79.2 2.4 80.4 423.6 ;
         LAYER metal3 ;
         RECT  112.8 288.0 147.6 289.2 ;
         LAYER metal3 ;
         RECT  0.0 144.0 210.0 145.2 ;
         LAYER metal3 ;
         RECT  0.0 158.4 210.0 159.6 ;
         LAYER metal3 ;
         RECT  0.0 225.6 87.6 226.8 ;
         LAYER metal4 ;
         RECT  160.8 2.4 162.0 423.6 ;
         LAYER metal3 ;
         RECT  134.4 216.0 210.0 217.2 ;
         LAYER metal3 ;
         RECT  52.8 14.4 210.0 15.6 ;
         LAYER metal3 ;
         RECT  172.8 331.2 210.0 332.4 ;
         LAYER metal3 ;
         RECT  0.0 268.8 90.0 270.0 ;
         LAYER metal3 ;
         RECT  26.4 163.2 73.2 164.4 ;
         LAYER metal3 ;
         RECT  26.4 321.6 210.0 322.8 ;
         LAYER metal3 ;
         RECT  68.1 364.4 68.9 365.2 ;
         LAYER metal3 ;
         RECT  26.4 283.2 116.4 284.4 ;
         LAYER metal3 ;
         RECT  0.0 302.4 210.0 303.6 ;
         LAYER metal3 ;
         RECT  77.6 102.4 78.4 103.2 ;
         LAYER metal3 ;
         RECT  129.6 201.6 169.2 202.8 ;
         LAYER metal3 ;
         RECT  167.2 238.0 168.0 238.8 ;
         LAYER metal3 ;
         RECT  33.6 235.2 210.0 236.4 ;
         LAYER metal3 ;
         RECT  4.8 43.2 73.2 44.4 ;
         LAYER metal3 ;
         RECT  192.2 159.6 193.0 160.4 ;
         LAYER metal4 ;
         RECT  165.6 2.4 166.8 423.6 ;
         LAYER metal3 ;
         RECT  177.6 168.0 205.2 169.2 ;
         LAYER metal3 ;
         RECT  10.0 263.2 10.8 264.0 ;
         LAYER metal3 ;
         RECT  0.0 72.0 75.6 73.2 ;
         LAYER metal3 ;
         RECT  205.3 321.2 206.1 322.0 ;
         LAYER metal3 ;
         RECT  0.0 240.0 210.0 241.2 ;
         LAYER metal3 ;
         RECT  0.0 148.8 27.6 150.0 ;
         LAYER metal3 ;
         RECT  192.5 74.0 193.3 74.8 ;
         LAYER metal3 ;
         RECT  178.1 279.6 178.9 280.4 ;
         LAYER metal3 ;
         RECT  172.8 249.6 210.0 250.8 ;
         LAYER metal4 ;
         RECT  60.0 2.4 61.2 423.6 ;
         LAYER metal3 ;
         RECT  178.1 196.4 178.9 197.2 ;
         LAYER metal3 ;
         RECT  0.0 177.6 210.0 178.8 ;
         LAYER metal3 ;
         RECT  152.0 238.0 152.8 238.8 ;
         LAYER metal4 ;
         RECT  117.6 2.4 118.8 423.6 ;
         LAYER metal3 ;
         RECT  0.0 264.0 116.4 265.2 ;
         LAYER metal3 ;
         RECT  81.6 43.2 210.0 44.4 ;
         LAYER metal4 ;
         RECT  55.2 2.4 56.4 423.6 ;
         LAYER metal4 ;
         RECT  208.8 2.4 210.0 423.6 ;
         LAYER metal3 ;
         RECT  0.0 4.8 44.4 6.0 ;
         LAYER metal3 ;
         RECT  178.1 258.8 178.9 259.6 ;
         LAYER metal3 ;
         RECT  0.0 187.2 87.6 188.4 ;
         LAYER metal3 ;
         RECT  108.1 196.4 108.9 197.2 ;
         LAYER metal3 ;
         RECT  178.1 175.6 178.9 176.4 ;
         LAYER metal3 ;
         RECT  88.8 374.4 210.0 375.6 ;
         LAYER metal3 ;
         RECT  167.2 279.6 168.0 280.4 ;
         LAYER metal3 ;
         RECT  0.0 28.8 27.6 30.0 ;
         LAYER metal3 ;
         RECT  33.6 172.8 210.0 174.0 ;
         LAYER metal3 ;
         RECT  0.0 364.8 210.0 366.0 ;
         LAYER metal3 ;
         RECT  0.0 249.6 87.6 250.8 ;
         LAYER metal3 ;
         RECT  0.0 196.8 121.2 198.0 ;
         LAYER metal3 ;
         RECT  0.0 201.6 116.4 202.8 ;
         LAYER metal4 ;
         RECT  16.8 2.4 18.0 423.6 ;
         LAYER metal3 ;
         RECT  0.0 120.0 73.2 121.2 ;
         LAYER metal4 ;
         RECT  26.4 2.4 27.6 423.6 ;
         LAYER metal3 ;
         RECT  77.6 62.4 78.4 63.2 ;
         LAYER metal3 ;
         RECT  0.0 96.0 210.0 97.2 ;
         LAYER metal3 ;
         RECT  0.0 211.2 116.4 212.4 ;
         LAYER metal4 ;
         RECT  40.8 2.4 42.0 423.6 ;
         LAYER metal3 ;
         RECT  93.1 217.2 93.9 218.0 ;
         LAYER metal3 ;
         RECT  111.7 22.4 112.5 23.2 ;
         LAYER metal3 ;
         RECT  0.0 259.2 121.2 260.4 ;
         LAYER metal3 ;
         RECT  86.4 355.2 166.8 356.4 ;
         LAYER metal4 ;
         RECT  132.0 2.4 133.2 423.6 ;
         LAYER metal3 ;
         RECT  172.8 206.4 210.0 207.6 ;
         LAYER metal3 ;
         RECT  0.0 182.4 169.2 183.6 ;
         LAYER metal4 ;
         RECT  84.0 2.4 85.2 423.6 ;
         LAYER metal3 ;
         RECT  129.6 220.8 169.2 222.0 ;
         LAYER metal3 ;
         RECT  0.0 81.6 73.2 82.8 ;
         LAYER metal3 ;
         RECT  26.4 244.8 169.2 246.0 ;
         LAYER metal3 ;
         RECT  72.0 345.6 169.2 346.8 ;
         LAYER metal3 ;
         RECT  0.0 62.4 210.0 63.6 ;
         LAYER metal3 ;
         RECT  178.1 342.0 178.9 342.8 ;
         LAYER metal3 ;
         RECT  0.0 412.8 70.8 414.0 ;
         LAYER metal3 ;
         RECT  167.2 196.4 168.0 197.2 ;
         LAYER metal3 ;
         RECT  205.3 362.8 206.1 363.6 ;
         LAYER metal3 ;
         RECT  167.2 321.2 168.0 322.0 ;
         LAYER metal3 ;
         RECT  172.8 288.0 210.0 289.2 ;
         LAYER metal3 ;
         RECT  0.0 403.2 210.0 404.4 ;
         LAYER metal4 ;
         RECT  180.0 2.4 181.2 423.6 ;
         LAYER metal3 ;
         RECT  0.0 76.8 210.0 78.0 ;
         LAYER metal3 ;
         RECT  0.0 355.2 70.8 356.4 ;
         LAYER metal3 ;
         RECT  178.1 321.2 178.9 322.0 ;
         LAYER metal3 ;
         RECT  23.2 302.4 24.0 303.2 ;
         LAYER metal3 ;
         RECT  0.0 297.6 210.0 298.8 ;
         LAYER metal3 ;
         RECT  0.0 115.2 210.0 116.4 ;
         LAYER metal3 ;
         RECT  152.0 300.4 152.8 301.2 ;
         LAYER metal4 ;
         RECT  122.4 2.4 123.6 423.6 ;
         LAYER metal3 ;
         RECT  172.8 312.0 210.0 313.2 ;
         LAYER metal3 ;
         RECT  0.0 52.8 39.6 54.0 ;
         LAYER metal3 ;
         RECT  112.8 225.6 147.6 226.8 ;
         LAYER metal3 ;
         RECT  0.0 33.6 210.0 34.8 ;
         LAYER metal3 ;
         RECT  0.0 153.6 75.6 154.8 ;
         LAYER metal3 ;
         RECT  167.2 300.4 168.0 301.2 ;
         LAYER metal3 ;
         RECT  0.0 288.0 87.6 289.2 ;
         LAYER metal3 ;
         RECT  69.6 384.0 210.0 385.2 ;
         LAYER metal4 ;
         RECT  36.0 2.4 37.2 423.6 ;
         LAYER metal3 ;
         RECT  129.6 254.4 169.2 255.6 ;
         LAYER metal4 ;
         RECT  69.6 2.4 70.8 423.6 ;
         LAYER metal3 ;
         RECT  77.6 142.4 78.4 143.2 ;
         LAYER metal4 ;
         RECT  204.0 2.4 205.2 423.6 ;
         LAYER metal3 ;
         RECT  205.3 300.4 206.1 301.2 ;
         LAYER metal3 ;
         RECT  185.4 159.6 186.2 160.4 ;
         LAYER metal3 ;
         RECT  129.6 211.2 169.2 212.4 ;
         LAYER metal3 ;
         RECT  172.8 350.4 210.0 351.6 ;
         LAYER metal3 ;
         RECT  152.0 321.2 152.8 322.0 ;
         LAYER metal3 ;
         RECT  172.8 268.8 210.0 270.0 ;
         LAYER metal4 ;
         RECT  112.8 2.4 114.0 423.6 ;
         LAYER metal4 ;
         RECT  189.6 2.4 190.8 423.6 ;
         LAYER metal3 ;
         RECT  0.0 9.6 210.0 10.8 ;
         LAYER metal3 ;
         RECT  167.2 217.2 168.0 218.0 ;
         LAYER metal3 ;
         RECT  91.2 412.8 210.0 414.0 ;
         LAYER metal3 ;
         RECT  205.3 279.6 206.1 280.4 ;
         LAYER metal3 ;
         RECT  205.3 258.8 206.1 259.6 ;
         LAYER metal3 ;
         RECT  93.1 258.8 93.9 259.6 ;
         LAYER metal3 ;
         RECT  77.6 22.4 78.4 23.2 ;
         LAYER metal3 ;
         RECT  0.0 316.8 169.2 318.0 ;
         LAYER metal4 ;
         RECT  7.2 2.4 8.4 423.6 ;
         LAYER metal3 ;
         RECT  0.0 345.6 63.6 346.8 ;
         LAYER metal3 ;
         RECT  184.9 175.6 185.7 176.4 ;
         LAYER metal3 ;
         RECT  0.0 100.8 186.0 102.0 ;
         LAYER metal3 ;
         RECT  178.1 362.8 178.9 363.6 ;
         LAYER metal3 ;
         RECT  0.0 134.4 210.0 135.6 ;
         LAYER metal3 ;
         RECT  0.0 379.2 210.0 380.4 ;
         LAYER metal3 ;
         RECT  155.2 175.6 156.0 176.4 ;
         LAYER metal3 ;
         RECT  129.6 283.2 169.2 284.4 ;
         LAYER metal3 ;
         RECT  129.6 264.0 169.2 265.2 ;
         LAYER metal3 ;
         RECT  0.0 192.0 116.4 193.2 ;
         LAYER metal3 ;
         RECT  199.3 74.0 200.1 74.8 ;
         LAYER metal3 ;
         RECT  0.0 230.4 210.0 231.6 ;
         LAYER metal3 ;
         RECT  141.6 278.4 210.0 279.6 ;
         LAYER metal3 ;
         RECT  0.0 408.0 210.0 409.2 ;
         LAYER metal3 ;
         RECT  33.6 331.2 147.6 332.4 ;
         LAYER metal3 ;
         RECT  198.5 175.6 199.3 176.4 ;
         LAYER metal3 ;
         RECT  152.0 279.6 152.8 280.4 ;
         LAYER metal3 ;
         RECT  172.8 72.0 210.0 73.2 ;
         LAYER metal3 ;
         RECT  172.8 187.2 210.0 188.4 ;
         LAYER metal3 ;
         RECT  0.0 398.4 210.0 399.6 ;
         LAYER metal4 ;
         RECT  74.4 2.4 75.6 423.6 ;
         LAYER metal3 ;
         RECT  132.0 196.8 210.0 198.0 ;
         LAYER metal3 ;
         RECT  167.2 342.0 168.0 342.8 ;
         LAYER metal3 ;
         RECT  0.0 86.4 188.4 87.6 ;
         LAYER metal3 ;
         RECT  184.9 362.8 185.7 363.6 ;
         LAYER metal3 ;
         RECT  178.1 217.2 178.9 218.0 ;
         LAYER metal3 ;
         RECT  48.0 28.8 210.0 30.0 ;
         LAYER metal3 ;
         RECT  205.3 196.4 206.1 197.2 ;
         LAYER metal3 ;
         RECT  0.0 139.2 190.8 140.4 ;
         LAYER metal3 ;
         RECT  74.4 24.0 210.0 25.2 ;
         LAYER metal3 ;
         RECT  191.9 91.4 192.7 92.2 ;
         LAYER metal3 ;
         RECT  170.4 91.2 210.0 92.4 ;
         LAYER metal3 ;
         RECT  10.0 302.4 10.8 303.2 ;
         LAYER metal3 ;
         RECT  81.6 120.0 210.0 121.2 ;
         LAYER metal3 ;
         RECT  0.0 129.6 210.0 130.8 ;
         LAYER metal3 ;
         RECT  152.0 217.2 152.8 218.0 ;
         LAYER metal3 ;
         RECT  0.0 307.2 169.2 308.4 ;
         LAYER metal3 ;
         RECT  205.3 175.6 206.1 176.4 ;
         LAYER metal3 ;
         RECT  198.5 362.8 199.3 363.6 ;
         LAYER metal3 ;
         RECT  0.0 360.0 210.0 361.2 ;
         LAYER metal3 ;
         RECT  0.0 91.2 75.6 92.4 ;
         LAYER metal4 ;
         RECT  127.2 2.4 128.4 423.6 ;
         LAYER metal3 ;
         RECT  93.1 279.6 93.9 280.4 ;
         LAYER metal3 ;
         RECT  0.0 350.4 147.6 351.6 ;
         LAYER metal3 ;
         RECT  10.0 224.0 10.8 224.8 ;
         LAYER metal3 ;
         RECT  0.0 110.4 210.0 111.6 ;
         LAYER metal3 ;
         RECT  23.2 184.8 24.0 185.6 ;
         LAYER metal3 ;
         RECT  0.0 326.4 169.2 327.6 ;
         LAYER metal3 ;
         RECT  0.0 67.2 210.0 68.4 ;
         LAYER metal3 ;
         RECT  194.1 125.4 194.9 126.2 ;
         LAYER metal3 ;
         RECT  33.6 292.8 210.0 294.0 ;
         LAYER metal3 ;
         RECT  205.3 238.0 206.1 238.8 ;
         LAYER metal3 ;
         RECT  152.0 258.8 152.8 259.6 ;
         LAYER metal4 ;
         RECT  199.2 2.4 200.4 423.6 ;
         LAYER metal3 ;
         RECT  0.0 340.8 210.0 342.0 ;
         LAYER metal3 ;
         RECT  108.1 279.6 108.9 280.4 ;
         LAYER metal3 ;
         RECT  0.0 336.0 169.2 337.2 ;
         LAYER metal3 ;
         RECT  0.0 168.0 166.8 169.2 ;
         LAYER metal3 ;
         RECT  152.0 342.0 152.8 342.8 ;
         LAYER metal3 ;
         RECT  0.0 19.2 210.0 20.4 ;
         LAYER metal3 ;
         RECT  167.2 258.8 168.0 259.6 ;
         LAYER metal3 ;
         RECT  129.6 273.6 169.2 274.8 ;
         LAYER metal3 ;
         RECT  0.0 388.8 210.0 390.0 ;
         LAYER metal3 ;
         RECT  0.0 422.4 63.6 423.6 ;
         LAYER metal4 ;
         RECT  151.2 2.4 152.4 423.6 ;
         LAYER metal4 ;
         RECT  146.4 2.4 147.6 423.6 ;
         LAYER metal3 ;
         RECT  108.1 217.2 108.9 218.0 ;
         LAYER metal3 ;
         RECT  33.6 273.6 116.4 274.8 ;
         LAYER metal3 ;
         RECT  93.1 196.4 93.9 197.2 ;
         LAYER metal4 ;
         RECT  141.6 2.4 142.8 423.6 ;
         LAYER metal3 ;
         RECT  0.0 24.0 37.2 25.2 ;
         LAYER metal3 ;
         RECT  108.1 258.8 108.9 259.6 ;
         LAYER metal3 ;
         RECT  0.0 48.0 210.0 49.2 ;
         LAYER metal3 ;
         RECT  10.0 184.8 10.8 185.6 ;
         LAYER metal3 ;
         RECT  10.0 341.6 10.8 342.4 ;
         LAYER metal4 ;
         RECT  88.8 2.4 90.0 423.6 ;
         LAYER metal3 ;
         RECT  0.0 417.6 210.0 418.8 ;
         LAYER metal3 ;
         RECT  68.1 404.4 68.9 405.2 ;
         LAYER metal3 ;
         RECT  2.0 22.4 2.8 23.2 ;
         LAYER metal3 ;
         RECT  172.8 225.6 210.0 226.8 ;
         LAYER metal4 ;
         RECT  2.4 2.4 3.6 423.6 ;
         LAYER metal3 ;
         RECT  67.2 52.8 210.0 54.0 ;
         LAYER metal4 ;
         RECT  194.4 2.4 195.6 423.6 ;
         LAYER metal4 ;
         RECT  103.2 2.4 104.4 423.6 ;
         LAYER metal4 ;
         RECT  45.6 2.4 46.8 423.6 ;
         LAYER metal4 ;
         RECT  156.0 2.4 157.2 423.6 ;
         LAYER metal3 ;
         RECT  33.6 312.0 147.6 313.2 ;
         LAYER metal4 ;
         RECT  93.6 2.4 94.8 423.6 ;
         LAYER metal3 ;
         RECT  205.3 217.2 206.1 218.0 ;
         LAYER metal3 ;
         RECT  0.0 57.6 210.0 58.8 ;
         LAYER metal4 ;
         RECT  98.4 2.4 99.6 423.6 ;
         LAYER metal3 ;
         RECT  91.2 393.6 210.0 394.8 ;
         LAYER metal3 ;
         RECT  191.7 175.6 192.5 176.4 ;
         LAYER metal3 ;
         RECT  72.0 422.4 210.0 423.6 ;
         LAYER metal3 ;
         RECT  0.0 105.6 210.0 106.8 ;
         LAYER metal4 ;
         RECT  175.2 2.4 176.4 423.6 ;
         LAYER metal3 ;
         RECT  23.2 263.2 24.0 264.0 ;
         LAYER metal3 ;
         RECT  129.6 192.0 169.2 193.2 ;
         LAYER metal4 ;
         RECT  64.8 2.4 66.0 423.6 ;
         LAYER metal4 ;
         RECT  170.4 2.4 171.6 423.6 ;
         LAYER metal3 ;
         RECT  81.6 163.2 210.0 164.4 ;
         LAYER metal4 ;
         RECT  108.0 2.4 109.2 423.6 ;
         LAYER metal3 ;
         RECT  178.1 300.4 178.9 301.2 ;
         LAYER metal3 ;
         RECT  0.0 38.4 210.0 39.6 ;
         LAYER metal3 ;
         RECT  26.4 206.4 90.0 207.6 ;
         LAYER metal4 ;
         RECT  21.6 2.4 22.8 423.6 ;
         LAYER metal3 ;
         RECT  0.0 124.8 34.8 126.0 ;
         LAYER metal3 ;
         RECT  199.0 159.6 199.8 160.4 ;
         LAYER metal3 ;
         RECT  191.7 362.8 192.5 363.6 ;
         LAYER metal3 ;
         RECT  0.0 393.6 70.8 394.8 ;
         LAYER metal3 ;
         RECT  0.0 374.4 70.8 375.6 ;
         LAYER metal4 ;
         RECT  184.8 2.4 186.0 423.6 ;
         LAYER metal3 ;
         RECT  178.1 238.0 178.9 238.8 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal3 ;
         RECT  0.0 98.4 210.0 99.6 ;
         LAYER metal3 ;
         RECT  181.5 243.0 182.3 243.8 ;
         LAYER metal3 ;
         RECT  72.0 362.4 174.0 363.6 ;
         LAYER metal3 ;
         RECT  201.9 253.8 202.7 254.6 ;
         LAYER metal3 ;
         RECT  68.1 344.4 68.9 345.2 ;
         LAYER metal3 ;
         RECT  10.0 165.2 10.8 166.0 ;
         LAYER metal3 ;
         RECT  23.2 322.0 24.0 322.8 ;
         LAYER metal3 ;
         RECT  0.0 237.6 147.6 238.8 ;
         LAYER metal3 ;
         RECT  0.0 295.2 210.0 296.4 ;
         LAYER metal4 ;
         RECT  52.8 2.4 54.0 423.6 ;
         LAYER metal3 ;
         RECT  181.5 253.8 182.3 254.6 ;
         LAYER metal3 ;
         RECT  129.6 189.6 210.0 190.8 ;
         LAYER metal3 ;
         RECT  0.0 367.2 210.0 368.4 ;
         LAYER metal3 ;
         RECT  174.7 170.6 175.5 171.4 ;
         LAYER metal3 ;
         RECT  172.6 167.8 173.4 168.6 ;
         LAYER metal3 ;
         RECT  0.0 136.8 210.0 138.0 ;
         LAYER metal3 ;
         RECT  2.0 42.4 2.8 43.2 ;
         LAYER metal3 ;
         RECT  0.0 333.6 210.0 334.8 ;
         LAYER metal3 ;
         RECT  208.7 263.8 209.5 264.6 ;
         LAYER metal3 ;
         RECT  167.2 310.8 168.0 311.6 ;
         LAYER metal3 ;
         RECT  208.7 180.6 209.5 181.4 ;
         LAYER metal3 ;
         RECT  81.6 103.2 210.0 104.4 ;
         LAYER metal3 ;
         RECT  26.4 184.8 121.2 186.0 ;
         LAYER metal3 ;
         RECT  174.7 326.2 175.5 327.0 ;
         LAYER metal4 ;
         RECT  196.8 2.4 198.0 423.6 ;
         LAYER metal3 ;
         RECT  0.0 338.4 210.0 339.6 ;
         LAYER metal3 ;
         RECT  210.8 355.0 211.6 355.8 ;
         LAYER metal3 ;
         RECT  208.7 337.0 209.5 337.8 ;
         LAYER metal3 ;
         RECT  77.6 162.4 78.4 163.2 ;
         LAYER metal3 ;
         RECT  0.0 160.8 181.2 162.0 ;
         LAYER metal3 ;
         RECT  0.0 199.2 121.2 200.4 ;
         LAYER metal3 ;
         RECT  0.0 266.4 210.0 267.6 ;
         LAYER metal4 ;
         RECT  62.4 2.4 63.6 423.6 ;
         LAYER metal4 ;
         RECT  115.2 2.4 116.4 423.6 ;
         LAYER metal3 ;
         RECT  108.1 206.8 108.9 207.6 ;
         LAYER metal4 ;
         RECT  105.6 2.4 106.8 423.6 ;
         LAYER metal4 ;
         RECT  33.6 2.4 34.8 423.6 ;
         LAYER metal3 ;
         RECT  181.5 263.8 182.3 264.6 ;
         LAYER metal3 ;
         RECT  152.0 331.6 152.8 332.4 ;
         LAYER metal4 ;
         RECT  120.0 2.4 121.2 423.6 ;
         LAYER metal4 ;
         RECT  158.4 2.4 159.6 423.6 ;
         LAYER metal3 ;
         RECT  77.6 42.4 78.4 43.2 ;
         LAYER metal4 ;
         RECT  153.6 2.4 154.8 423.6 ;
         LAYER metal3 ;
         RECT  0.0 228.0 210.0 229.2 ;
         LAYER metal3 ;
         RECT  0.0 328.8 210.0 330.0 ;
         LAYER metal3 ;
         RECT  0.0 180.0 210.0 181.2 ;
         LAYER metal3 ;
         RECT  4.8 21.6 73.2 22.8 ;
         LAYER metal4 ;
         RECT  100.8 2.4 102.0 423.6 ;
         LAYER metal3 ;
         RECT  172.8 112.8 210.0 114.0 ;
         LAYER metal3 ;
         RECT  0.0 117.6 210.0 118.8 ;
         LAYER metal3 ;
         RECT  0.0 247.2 121.2 248.4 ;
         LAYER metal3 ;
         RECT  167.2 227.6 168.0 228.4 ;
         LAYER metal3 ;
         RECT  181.5 337.0 182.3 337.8 ;
         LAYER metal3 ;
         RECT  0.0 60.0 73.2 61.2 ;
         LAYER metal3 ;
         RECT  188.3 357.8 189.1 358.6 ;
         LAYER metal3 ;
         RECT  33.6 271.2 121.2 272.4 ;
         LAYER metal3 ;
         RECT  174.7 233.0 175.5 233.8 ;
         LAYER metal3 ;
         RECT  0.0 386.4 210.0 387.6 ;
         LAYER metal4 ;
         RECT  43.2 2.4 44.4 423.6 ;
         LAYER metal4 ;
         RECT  72.0 2.4 73.2 423.6 ;
         LAYER metal4 ;
         RECT  206.4 2.4 207.6 423.6 ;
         LAYER metal3 ;
         RECT  193.9 85.0 194.7 85.8 ;
         LAYER metal3 ;
         RECT  0.0 31.2 27.6 32.4 ;
         LAYER metal3 ;
         RECT  129.6 285.6 210.0 286.8 ;
         LAYER metal3 ;
         RECT  93.1 227.6 93.9 228.4 ;
         LAYER metal3 ;
         RECT  136.8 247.2 210.0 248.4 ;
         LAYER metal3 ;
         RECT  167.2 352.4 168.0 353.2 ;
         LAYER metal3 ;
         RECT  201.9 233.0 202.7 233.8 ;
         LAYER metal3 ;
         RECT  23.2 204.4 24.0 205.2 ;
         LAYER metal4 ;
         RECT  163.2 2.4 164.4 423.6 ;
         LAYER metal3 ;
         RECT  167.2 206.8 168.0 207.6 ;
         LAYER metal3 ;
         RECT  132.0 184.8 210.0 186.0 ;
         LAYER metal3 ;
         RECT  201.9 138.8 202.7 139.6 ;
         LAYER metal3 ;
         RECT  201.9 316.2 202.7 317.0 ;
         LAYER metal3 ;
         RECT  0.0 16.8 210.0 18.0 ;
         LAYER metal3 ;
         RECT  0.0 45.6 210.0 46.8 ;
         LAYER metal3 ;
         RECT  60.0 122.4 210.0 123.6 ;
         LAYER metal3 ;
         RECT  0.0 218.4 87.6 219.6 ;
         LAYER metal3 ;
         RECT  0.0 108.0 210.0 109.2 ;
         LAYER metal3 ;
         RECT  208.7 253.8 209.5 254.6 ;
         LAYER metal3 ;
         RECT  0.0 141.6 73.2 142.8 ;
         LAYER metal3 ;
         RECT  201.9 222.2 202.7 223.0 ;
         LAYER metal3 ;
         RECT  0.0 381.6 210.0 382.8 ;
         LAYER metal4 ;
         RECT  129.6 2.4 130.8 423.6 ;
         LAYER metal3 ;
         RECT  208.7 274.6 209.5 275.4 ;
         LAYER metal3 ;
         RECT  174.7 305.4 175.5 306.2 ;
         LAYER metal3 ;
         RECT  10.0 243.6 10.8 244.4 ;
         LAYER metal3 ;
         RECT  0.0 103.2 73.2 104.4 ;
         LAYER metal3 ;
         RECT  195.1 138.8 195.9 139.6 ;
         LAYER metal3 ;
         RECT  2.0 2.4 2.8 3.2 ;
         LAYER metal3 ;
         RECT  86.4 348.0 210.0 349.2 ;
         LAYER metal4 ;
         RECT  28.8 2.4 30.0 423.6 ;
         LAYER metal3 ;
         RECT  26.4 223.2 116.4 224.4 ;
         LAYER metal3 ;
         RECT  208.7 222.2 209.5 223.0 ;
         LAYER metal3 ;
         RECT  201.9 170.6 202.7 171.4 ;
         LAYER metal3 ;
         RECT  0.0 324.0 210.0 325.2 ;
         LAYER metal4 ;
         RECT  19.2 2.4 20.4 423.6 ;
         LAYER metal4 ;
         RECT  182.4 2.4 183.6 423.6 ;
         LAYER metal4 ;
         RECT  81.6 2.4 82.8 423.6 ;
         LAYER metal3 ;
         RECT  93.1 248.4 93.9 249.2 ;
         LAYER metal3 ;
         RECT  208.7 295.4 209.5 296.2 ;
         LAYER metal3 ;
         RECT  0.0 55.2 210.0 56.4 ;
         LAYER metal3 ;
         RECT  33.6 252.0 116.4 253.2 ;
         LAYER metal3 ;
         RECT  0.0 319.2 147.6 320.4 ;
         LAYER metal3 ;
         RECT  0.0 396.0 210.0 397.2 ;
         LAYER metal3 ;
         RECT  10.0 322.0 10.8 322.8 ;
         LAYER metal3 ;
         RECT  0.0 348.0 54.0 349.2 ;
         LAYER metal3 ;
         RECT  167.2 186.0 168.0 186.8 ;
         LAYER metal3 ;
         RECT  181.5 180.6 182.3 181.4 ;
         LAYER metal3 ;
         RECT  208.7 212.2 209.5 213.0 ;
         LAYER metal3 ;
         RECT  174.7 347.0 175.5 347.8 ;
         LAYER metal3 ;
         RECT  181.5 274.6 182.3 275.4 ;
         LAYER metal3 ;
         RECT  152.0 269.2 152.8 270.0 ;
         LAYER metal3 ;
         RECT  152.0 290.0 152.8 290.8 ;
         LAYER metal3 ;
         RECT  0.0 309.6 210.0 310.8 ;
         LAYER metal4 ;
         RECT  177.6 2.4 178.8 423.6 ;
         LAYER metal3 ;
         RECT  208.7 201.4 209.5 202.2 ;
         LAYER metal4 ;
         RECT  96.0 2.4 97.2 423.6 ;
         LAYER metal3 ;
         RECT  23.2 282.8 24.0 283.6 ;
         LAYER metal3 ;
         RECT  81.6 141.6 210.0 142.8 ;
         LAYER metal3 ;
         RECT  181.5 347.0 182.3 347.8 ;
         LAYER metal3 ;
         RECT  208.7 191.4 209.5 192.2 ;
         LAYER metal3 ;
         RECT  26.4 261.6 121.2 262.8 ;
         LAYER metal3 ;
         RECT  76.8 2.4 210.0 3.6 ;
         LAYER metal3 ;
         RECT  0.0 314.4 210.0 315.6 ;
         LAYER metal3 ;
         RECT  0.0 405.6 63.6 406.8 ;
         LAYER metal4 ;
         RECT  48.0 2.4 49.2 423.6 ;
         LAYER metal4 ;
         RECT  168.0 2.4 169.2 423.6 ;
         LAYER metal4 ;
         RECT  187.2 2.4 188.4 423.6 ;
         LAYER metal3 ;
         RECT  152.0 352.4 152.8 353.2 ;
         LAYER metal3 ;
         RECT  111.7 2.4 112.5 3.2 ;
         LAYER metal3 ;
         RECT  129.6 208.8 210.0 210.0 ;
         LAYER metal3 ;
         RECT  0.0 2.4 44.4 3.6 ;
         LAYER metal3 ;
         RECT  0.0 357.6 210.0 358.8 ;
         LAYER metal3 ;
         RECT  174.7 337.0 175.5 337.8 ;
         LAYER metal3 ;
         RECT  0.0 26.4 37.2 27.6 ;
         LAYER metal4 ;
         RECT  134.4 2.4 135.6 423.6 ;
         LAYER metal4 ;
         RECT  192.0 2.4 193.2 423.6 ;
         LAYER metal4 ;
         RECT  139.2 2.4 140.4 423.6 ;
         LAYER metal3 ;
         RECT  188.3 170.6 189.1 171.4 ;
         LAYER metal3 ;
         RECT  0.0 242.4 210.0 243.6 ;
         LAYER metal3 ;
         RECT  93.1 269.2 93.9 270.0 ;
         LAYER metal3 ;
         RECT  0.0 420.0 210.0 421.2 ;
         LAYER metal3 ;
         RECT  201.9 347.0 202.7 347.8 ;
         LAYER metal3 ;
         RECT  0.0 132.0 210.0 133.2 ;
         LAYER metal3 ;
         RECT  181.5 357.8 182.3 358.6 ;
         LAYER metal3 ;
         RECT  199.3 80.6 200.1 81.4 ;
         LAYER metal3 ;
         RECT  0.0 146.4 27.6 147.6 ;
         LAYER metal3 ;
         RECT  0.0 12.0 210.0 13.2 ;
         LAYER metal3 ;
         RECT  208.7 233.0 209.5 233.8 ;
         LAYER metal3 ;
         RECT  81.6 60.0 210.0 61.2 ;
         LAYER metal3 ;
         RECT  0.0 112.8 75.6 114.0 ;
         LAYER metal3 ;
         RECT  201.9 284.6 202.7 285.4 ;
         LAYER metal3 ;
         RECT  0.0 204.0 210.0 205.2 ;
         LAYER metal3 ;
         RECT  174.7 274.6 175.5 275.4 ;
         LAYER metal3 ;
         RECT  174.7 253.8 175.5 254.6 ;
         LAYER metal3 ;
         RECT  181.5 212.2 182.3 213.0 ;
         LAYER metal3 ;
         RECT  201.9 212.2 202.7 213.0 ;
         LAYER metal3 ;
         RECT  170.4 151.2 210.0 152.4 ;
         LAYER metal3 ;
         RECT  0.0 156.0 210.0 157.2 ;
         LAYER metal3 ;
         RECT  0.0 93.6 210.0 94.8 ;
         LAYER metal3 ;
         RECT  201.9 243.0 202.7 243.8 ;
         LAYER metal3 ;
         RECT  0.0 285.6 116.4 286.8 ;
         LAYER metal3 ;
         RECT  33.6 232.8 210.0 234.0 ;
         LAYER metal3 ;
         RECT  0.0 372.0 210.0 373.2 ;
         LAYER metal3 ;
         RECT  0.0 415.2 70.8 416.4 ;
         LAYER metal3 ;
         RECT  0.0 304.8 210.0 306.0 ;
         LAYER metal3 ;
         RECT  174.7 191.4 175.5 192.2 ;
         LAYER metal3 ;
         RECT  191.1 99.6 191.9 100.4 ;
         LAYER metal3 ;
         RECT  133.5 2.4 134.3 3.2 ;
         LAYER metal4 ;
         RECT  4.8 2.4 6.0 423.6 ;
         LAYER metal3 ;
         RECT  208.7 347.0 209.5 347.8 ;
         LAYER metal3 ;
         RECT  108.1 186.0 108.9 186.8 ;
         LAYER metal3 ;
         RECT  93.1 206.8 93.9 207.6 ;
         LAYER metal3 ;
         RECT  93.1 186.0 93.9 186.8 ;
         LAYER metal3 ;
         RECT  174.7 243.0 175.5 243.8 ;
         LAYER metal3 ;
         RECT  68.1 424.4 68.9 425.2 ;
         LAYER metal3 ;
         RECT  174.7 201.4 175.5 202.2 ;
         LAYER metal3 ;
         RECT  0.0 36.0 34.8 37.2 ;
         LAYER metal3 ;
         RECT  0.0 64.8 210.0 66.0 ;
         LAYER metal3 ;
         RECT  208.7 170.6 209.5 171.4 ;
         LAYER metal3 ;
         RECT  192.5 80.6 193.3 81.4 ;
         LAYER metal3 ;
         RECT  10.0 282.8 10.8 283.6 ;
         LAYER metal3 ;
         RECT  208.7 243.0 209.5 243.8 ;
         LAYER metal4 ;
         RECT  9.6 2.4 10.8 423.6 ;
         LAYER metal3 ;
         RECT  195.1 357.8 195.9 358.6 ;
         LAYER metal3 ;
         RECT  208.7 305.4 209.5 306.2 ;
         LAYER metal3 ;
         RECT  208.7 284.6 209.5 285.4 ;
         LAYER metal3 ;
         RECT  0.0 391.2 210.0 392.4 ;
         LAYER metal3 ;
         RECT  0.0 170.4 210.0 171.6 ;
         LAYER metal3 ;
         RECT  0.0 127.2 188.4 128.4 ;
         LAYER metal3 ;
         RECT  0.0 276.0 210.0 277.2 ;
         LAYER metal3 ;
         RECT  129.6 223.2 210.0 224.4 ;
         LAYER metal3 ;
         RECT  201.9 180.6 202.7 181.4 ;
         LAYER metal4 ;
         RECT  148.8 2.4 150.0 423.6 ;
         LAYER metal3 ;
         RECT  181.5 233.0 182.3 233.8 ;
         LAYER metal3 ;
         RECT  0.0 122.4 34.8 123.6 ;
         LAYER metal3 ;
         RECT  33.6 194.4 87.6 195.6 ;
         LAYER metal3 ;
         RECT  108.1 227.6 108.9 228.4 ;
         LAYER metal3 ;
         RECT  174.7 357.8 175.5 358.6 ;
         LAYER metal3 ;
         RECT  148.8 7.2 210.0 8.4 ;
         LAYER metal3 ;
         RECT  167.2 331.6 168.0 332.4 ;
         LAYER metal3 ;
         RECT  181.5 170.6 182.3 171.4 ;
         LAYER metal3 ;
         RECT  181.5 305.4 182.3 306.2 ;
         LAYER metal3 ;
         RECT  201.9 305.4 202.7 306.2 ;
         LAYER metal3 ;
         RECT  174.7 284.6 175.5 285.4 ;
         LAYER metal3 ;
         RECT  201.9 201.4 202.7 202.2 ;
         LAYER metal3 ;
         RECT  0.0 151.2 75.6 152.4 ;
         LAYER metal3 ;
         RECT  23.2 165.2 24.0 166.0 ;
         LAYER metal3 ;
         RECT  74.4 26.4 210.0 27.6 ;
         LAYER metal4 ;
         RECT  67.2 2.4 68.4 423.6 ;
         LAYER metal3 ;
         RECT  210.8 167.8 211.6 168.6 ;
         LAYER metal3 ;
         RECT  26.4 300.0 147.6 301.2 ;
         LAYER metal3 ;
         RECT  48.0 31.2 210.0 32.4 ;
         LAYER metal3 ;
         RECT  0.0 400.8 210.0 402.0 ;
         LAYER metal3 ;
         RECT  208.7 357.8 209.5 358.6 ;
         LAYER metal3 ;
         RECT  174.7 222.2 175.5 223.0 ;
         LAYER metal4 ;
         RECT  124.8 2.4 126.0 423.6 ;
         LAYER metal3 ;
         RECT  139.2 21.6 210.0 22.8 ;
         LAYER metal4 ;
         RECT  144.0 2.4 145.2 423.6 ;
         LAYER metal3 ;
         RECT  129.6 199.2 210.0 200.4 ;
         LAYER metal3 ;
         RECT  152.0 248.4 152.8 249.2 ;
         LAYER metal3 ;
         RECT  0.0 165.6 210.0 166.8 ;
         LAYER metal3 ;
         RECT  181.5 222.2 182.3 223.0 ;
         LAYER metal3 ;
         RECT  129.6 271.2 210.0 272.4 ;
         LAYER metal4 ;
         RECT  172.8 2.4 174.0 423.6 ;
         LAYER metal3 ;
         RECT  72.0 405.6 210.0 406.8 ;
         LAYER metal3 ;
         RECT  152.0 186.0 152.8 186.8 ;
         LAYER metal3 ;
         RECT  67.2 36.0 210.0 37.2 ;
         LAYER metal3 ;
         RECT  200.7 85.0 201.5 85.8 ;
         LAYER metal3 ;
         RECT  108.1 290.0 108.9 290.8 ;
         LAYER metal3 ;
         RECT  181.5 295.4 182.3 296.2 ;
         LAYER metal3 ;
         RECT  10.0 204.4 10.8 205.2 ;
         LAYER metal3 ;
         RECT  0.0 352.8 70.8 354.0 ;
         LAYER metal3 ;
         RECT  152.0 206.8 152.8 207.6 ;
         LAYER metal3 ;
         RECT  67.2 50.4 210.0 51.6 ;
         LAYER metal3 ;
         RECT  0.0 189.6 116.4 190.8 ;
         LAYER metal4 ;
         RECT  76.8 2.4 78.0 423.6 ;
         LAYER metal4 ;
         RECT  110.4 2.4 111.6 423.6 ;
         LAYER metal3 ;
         RECT  181.5 284.6 182.3 285.4 ;
         LAYER metal3 ;
         RECT  23.2 243.6 24.0 244.4 ;
         LAYER metal3 ;
         RECT  152.0 227.6 152.8 228.4 ;
         LAYER metal4 ;
         RECT  201.6 2.4 202.8 423.6 ;
         LAYER metal3 ;
         RECT  167.2 269.2 168.0 270.0 ;
         LAYER metal3 ;
         RECT  201.9 337.0 202.7 337.8 ;
         LAYER metal4 ;
         RECT  0.0 2.4 1.2 423.6 ;
         LAYER metal3 ;
         RECT  174.7 212.2 175.5 213.0 ;
         LAYER metal3 ;
         RECT  201.9 263.8 202.7 264.6 ;
         LAYER metal3 ;
         RECT  181.5 326.2 182.3 327.0 ;
         LAYER metal3 ;
         RECT  174.7 295.4 175.5 296.2 ;
         LAYER metal3 ;
         RECT  33.6 175.2 150.0 176.4 ;
         LAYER metal3 ;
         RECT  0.0 88.8 210.0 90.0 ;
         LAYER metal3 ;
         RECT  181.5 201.4 182.3 202.2 ;
         LAYER metal3 ;
         RECT  0.0 84.0 210.0 85.2 ;
         LAYER metal3 ;
         RECT  129.6 252.0 210.0 253.2 ;
         LAYER metal3 ;
         RECT  0.0 7.2 75.6 8.4 ;
         LAYER metal3 ;
         RECT  0.0 79.2 210.0 80.4 ;
         LAYER metal3 ;
         RECT  77.6 82.4 78.4 83.2 ;
         LAYER metal4 ;
         RECT  86.4 2.4 87.6 423.6 ;
         LAYER metal3 ;
         RECT  201.9 326.2 202.7 327.0 ;
         LAYER metal3 ;
         RECT  195.1 170.6 195.9 171.4 ;
         LAYER metal3 ;
         RECT  0.0 40.8 210.0 42.0 ;
         LAYER metal3 ;
         RECT  86.4 352.8 210.0 354.0 ;
         LAYER metal3 ;
         RECT  26.4 343.2 147.6 344.4 ;
         LAYER metal4 ;
         RECT  91.2 2.4 92.4 423.6 ;
         LAYER metal3 ;
         RECT  174.7 263.8 175.5 264.6 ;
         LAYER metal3 ;
         RECT  152.0 310.8 152.8 311.6 ;
         LAYER metal3 ;
         RECT  0.0 74.4 75.6 75.6 ;
         LAYER metal3 ;
         RECT  0.0 280.8 87.6 282.0 ;
         LAYER metal3 ;
         RECT  208.7 326.2 209.5 327.0 ;
         LAYER metal3 ;
         RECT  68.1 384.4 68.9 385.2 ;
         LAYER metal3 ;
         RECT  33.6 290.4 210.0 291.6 ;
         LAYER metal3 ;
         RECT  201.9 191.4 202.7 192.2 ;
         LAYER metal3 ;
         RECT  129.6 261.6 210.0 262.8 ;
         LAYER metal3 ;
         RECT  197.9 99.6 198.7 100.4 ;
         LAYER metal3 ;
         RECT  181.5 191.4 182.3 192.2 ;
         LAYER metal3 ;
         RECT  208.7 316.2 209.5 317.0 ;
         LAYER metal3 ;
         RECT  108.1 248.4 108.9 249.2 ;
         LAYER metal3 ;
         RECT  33.6 213.6 210.0 214.8 ;
         LAYER metal3 ;
         RECT  0.0 208.8 121.2 210.0 ;
         LAYER metal3 ;
         RECT  108.1 269.2 108.9 270.0 ;
         LAYER metal3 ;
         RECT  91.2 415.2 210.0 416.4 ;
         LAYER metal4 ;
         RECT  24.0 2.4 25.2 423.6 ;
         LAYER metal3 ;
         RECT  0.0 410.4 210.0 411.6 ;
         LAYER metal3 ;
         RECT  77.6 2.4 78.4 3.2 ;
         LAYER metal3 ;
         RECT  0.0 256.8 87.6 258.0 ;
         LAYER metal4 ;
         RECT  38.4 2.4 39.6 423.6 ;
         LAYER metal4 ;
         RECT  14.4 2.4 15.6 423.6 ;
         LAYER metal3 ;
         RECT  201.9 295.4 202.7 296.2 ;
         LAYER metal3 ;
         RECT  0.0 362.4 63.6 363.6 ;
         LAYER metal4 ;
         RECT  57.6 2.4 58.8 423.6 ;
         LAYER metal3 ;
         RECT  77.6 122.4 78.4 123.2 ;
         LAYER metal3 ;
         RECT  0.0 50.4 39.6 51.6 ;
         LAYER metal3 ;
         RECT  172.6 355.0 173.4 355.8 ;
         LAYER metal3 ;
         RECT  0.0 376.8 210.0 378.0 ;
         LAYER metal3 ;
         RECT  181.5 316.2 182.3 317.0 ;
         LAYER metal3 ;
         RECT  174.7 180.6 175.5 181.4 ;
         LAYER metal3 ;
         RECT  201.9 357.8 202.7 358.6 ;
         LAYER metal3 ;
         RECT  0.0 69.6 210.0 70.8 ;
         LAYER metal3 ;
         RECT  201.9 274.6 202.7 275.4 ;
         LAYER metal3 ;
         RECT  167.2 248.4 168.0 249.2 ;
         LAYER metal3 ;
         RECT  174.7 316.2 175.5 317.0 ;
         LAYER metal3 ;
         RECT  167.2 290.0 168.0 290.8 ;
         LAYER metal3 ;
         RECT  93.1 290.0 93.9 290.8 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  188.3 196.4 195.9 197.2 ;
      RECT  190.9 193.4 192.5 194.2 ;
      RECT  193.3 192.4 194.1 194.8 ;
      RECT  195.1 190.0 195.9 194.2 ;
      RECT  188.3 188.6 195.9 189.4 ;
      RECT  192.1 189.4 192.9 189.6 ;
      RECT  190.9 194.2 191.7 194.8 ;
      RECT  193.1 194.8 194.1 195.6 ;
      RECT  190.7 190.4 191.7 191.2 ;
      RECT  195.1 194.8 195.9 196.4 ;
      RECT  188.3 194.8 189.1 196.4 ;
      RECT  192.9 191.6 194.1 192.4 ;
      RECT  193.3 191.2 194.1 191.6 ;
      RECT  193.3 190.4 194.3 191.2 ;
      RECT  189.9 187.2 191.5 188.0 ;
      RECT  192.7 187.2 194.3 188.0 ;
      RECT  190.9 194.8 191.9 195.6 ;
      RECT  188.3 190.0 189.1 194.2 ;
      RECT  190.9 191.2 191.7 193.4 ;
      RECT  188.3 197.2 195.9 196.4 ;
      RECT  190.9 200.2 192.5 199.4 ;
      RECT  193.3 201.2 194.1 198.8 ;
      RECT  195.1 203.6 195.9 199.4 ;
      RECT  188.3 205.0 195.9 204.2 ;
      RECT  192.1 204.2 192.9 204.0 ;
      RECT  190.9 199.4 191.7 198.8 ;
      RECT  193.1 198.8 194.1 198.0 ;
      RECT  190.7 203.2 191.7 202.4 ;
      RECT  195.1 198.8 195.9 197.2 ;
      RECT  188.3 198.8 189.1 197.2 ;
      RECT  192.9 202.0 194.1 201.2 ;
      RECT  193.3 202.4 194.1 202.0 ;
      RECT  193.3 203.2 194.3 202.4 ;
      RECT  189.9 206.4 191.5 205.6 ;
      RECT  192.7 206.4 194.3 205.6 ;
      RECT  190.9 198.8 191.9 198.0 ;
      RECT  188.3 203.6 189.1 199.4 ;
      RECT  190.9 202.4 191.7 200.2 ;
      RECT  188.3 217.2 195.9 218.0 ;
      RECT  190.9 214.2 192.5 215.0 ;
      RECT  193.3 213.2 194.1 215.6 ;
      RECT  195.1 210.8 195.9 215.0 ;
      RECT  188.3 209.4 195.9 210.2 ;
      RECT  192.1 210.2 192.9 210.4 ;
      RECT  190.9 215.0 191.7 215.6 ;
      RECT  193.1 215.6 194.1 216.4 ;
      RECT  190.7 211.2 191.7 212.0 ;
      RECT  195.1 215.6 195.9 217.2 ;
      RECT  188.3 215.6 189.1 217.2 ;
      RECT  192.9 212.4 194.1 213.2 ;
      RECT  193.3 212.0 194.1 212.4 ;
      RECT  193.3 211.2 194.3 212.0 ;
      RECT  189.9 208.0 191.5 208.8 ;
      RECT  192.7 208.0 194.3 208.8 ;
      RECT  190.9 215.6 191.9 216.4 ;
      RECT  188.3 210.8 189.1 215.0 ;
      RECT  190.9 212.0 191.7 214.2 ;
      RECT  188.3 218.0 195.9 217.2 ;
      RECT  190.9 221.0 192.5 220.2 ;
      RECT  193.3 222.0 194.1 219.6 ;
      RECT  195.1 224.4 195.9 220.2 ;
      RECT  188.3 225.8 195.9 225.0 ;
      RECT  192.1 225.0 192.9 224.8 ;
      RECT  190.9 220.2 191.7 219.6 ;
      RECT  193.1 219.6 194.1 218.8 ;
      RECT  190.7 224.0 191.7 223.2 ;
      RECT  195.1 219.6 195.9 218.0 ;
      RECT  188.3 219.6 189.1 218.0 ;
      RECT  192.9 222.8 194.1 222.0 ;
      RECT  193.3 223.2 194.1 222.8 ;
      RECT  193.3 224.0 194.3 223.2 ;
      RECT  189.9 227.2 191.5 226.4 ;
      RECT  192.7 227.2 194.3 226.4 ;
      RECT  190.9 219.6 191.9 218.8 ;
      RECT  188.3 224.4 189.1 220.2 ;
      RECT  190.9 223.2 191.7 221.0 ;
      RECT  188.3 238.0 195.9 238.8 ;
      RECT  190.9 235.0 192.5 235.8 ;
      RECT  193.3 234.0 194.1 236.4 ;
      RECT  195.1 231.6 195.9 235.8 ;
      RECT  188.3 230.2 195.9 231.0 ;
      RECT  192.1 231.0 192.9 231.2 ;
      RECT  190.9 235.8 191.7 236.4 ;
      RECT  193.1 236.4 194.1 237.2 ;
      RECT  190.7 232.0 191.7 232.8 ;
      RECT  195.1 236.4 195.9 238.0 ;
      RECT  188.3 236.4 189.1 238.0 ;
      RECT  192.9 233.2 194.1 234.0 ;
      RECT  193.3 232.8 194.1 233.2 ;
      RECT  193.3 232.0 194.3 232.8 ;
      RECT  189.9 228.8 191.5 229.6 ;
      RECT  192.7 228.8 194.3 229.6 ;
      RECT  190.9 236.4 191.9 237.2 ;
      RECT  188.3 231.6 189.1 235.8 ;
      RECT  190.9 232.8 191.7 235.0 ;
      RECT  188.3 238.8 195.9 238.0 ;
      RECT  190.9 241.8 192.5 241.0 ;
      RECT  193.3 242.8 194.1 240.4 ;
      RECT  195.1 245.2 195.9 241.0 ;
      RECT  188.3 246.6 195.9 245.8 ;
      RECT  192.1 245.8 192.9 245.6 ;
      RECT  190.9 241.0 191.7 240.4 ;
      RECT  193.1 240.4 194.1 239.6 ;
      RECT  190.7 244.8 191.7 244.0 ;
      RECT  195.1 240.4 195.9 238.8 ;
      RECT  188.3 240.4 189.1 238.8 ;
      RECT  192.9 243.6 194.1 242.8 ;
      RECT  193.3 244.0 194.1 243.6 ;
      RECT  193.3 244.8 194.3 244.0 ;
      RECT  189.9 248.0 191.5 247.2 ;
      RECT  192.7 248.0 194.3 247.2 ;
      RECT  190.9 240.4 191.9 239.6 ;
      RECT  188.3 245.2 189.1 241.0 ;
      RECT  190.9 244.0 191.7 241.8 ;
      RECT  188.3 258.8 195.9 259.6 ;
      RECT  190.9 255.8 192.5 256.6 ;
      RECT  193.3 254.8 194.1 257.2 ;
      RECT  195.1 252.4 195.9 256.6 ;
      RECT  188.3 251.0 195.9 251.8 ;
      RECT  192.1 251.8 192.9 252.0 ;
      RECT  190.9 256.6 191.7 257.2 ;
      RECT  193.1 257.2 194.1 258.0 ;
      RECT  190.7 252.8 191.7 253.6 ;
      RECT  195.1 257.2 195.9 258.8 ;
      RECT  188.3 257.2 189.1 258.8 ;
      RECT  192.9 254.0 194.1 254.8 ;
      RECT  193.3 253.6 194.1 254.0 ;
      RECT  193.3 252.8 194.3 253.6 ;
      RECT  189.9 249.6 191.5 250.4 ;
      RECT  192.7 249.6 194.3 250.4 ;
      RECT  190.9 257.2 191.9 258.0 ;
      RECT  188.3 252.4 189.1 256.6 ;
      RECT  190.9 253.6 191.7 255.8 ;
      RECT  188.3 259.6 195.9 258.8 ;
      RECT  190.9 262.6 192.5 261.8 ;
      RECT  193.3 263.6 194.1 261.2 ;
      RECT  195.1 266.0 195.9 261.8 ;
      RECT  188.3 267.4 195.9 266.6 ;
      RECT  192.1 266.6 192.9 266.4 ;
      RECT  190.9 261.8 191.7 261.2 ;
      RECT  193.1 261.2 194.1 260.4 ;
      RECT  190.7 265.6 191.7 264.8 ;
      RECT  195.1 261.2 195.9 259.6 ;
      RECT  188.3 261.2 189.1 259.6 ;
      RECT  192.9 264.4 194.1 263.6 ;
      RECT  193.3 264.8 194.1 264.4 ;
      RECT  193.3 265.6 194.3 264.8 ;
      RECT  189.9 268.8 191.5 268.0 ;
      RECT  192.7 268.8 194.3 268.0 ;
      RECT  190.9 261.2 191.9 260.4 ;
      RECT  188.3 266.0 189.1 261.8 ;
      RECT  190.9 264.8 191.7 262.6 ;
      RECT  188.3 279.6 195.9 280.4 ;
      RECT  190.9 276.6 192.5 277.4 ;
      RECT  193.3 275.6 194.1 278.0 ;
      RECT  195.1 273.2 195.9 277.4 ;
      RECT  188.3 271.8 195.9 272.6 ;
      RECT  192.1 272.6 192.9 272.8 ;
      RECT  190.9 277.4 191.7 278.0 ;
      RECT  193.1 278.0 194.1 278.8 ;
      RECT  190.7 273.6 191.7 274.4 ;
      RECT  195.1 278.0 195.9 279.6 ;
      RECT  188.3 278.0 189.1 279.6 ;
      RECT  192.9 274.8 194.1 275.6 ;
      RECT  193.3 274.4 194.1 274.8 ;
      RECT  193.3 273.6 194.3 274.4 ;
      RECT  189.9 270.4 191.5 271.2 ;
      RECT  192.7 270.4 194.3 271.2 ;
      RECT  190.9 278.0 191.9 278.8 ;
      RECT  188.3 273.2 189.1 277.4 ;
      RECT  190.9 274.4 191.7 276.6 ;
      RECT  188.3 280.4 195.9 279.6 ;
      RECT  190.9 283.4 192.5 282.6 ;
      RECT  193.3 284.4 194.1 282.0 ;
      RECT  195.1 286.8 195.9 282.6 ;
      RECT  188.3 288.2 195.9 287.4 ;
      RECT  192.1 287.4 192.9 287.2 ;
      RECT  190.9 282.6 191.7 282.0 ;
      RECT  193.1 282.0 194.1 281.2 ;
      RECT  190.7 286.4 191.7 285.6 ;
      RECT  195.1 282.0 195.9 280.4 ;
      RECT  188.3 282.0 189.1 280.4 ;
      RECT  192.9 285.2 194.1 284.4 ;
      RECT  193.3 285.6 194.1 285.2 ;
      RECT  193.3 286.4 194.3 285.6 ;
      RECT  189.9 289.6 191.5 288.8 ;
      RECT  192.7 289.6 194.3 288.8 ;
      RECT  190.9 282.0 191.9 281.2 ;
      RECT  188.3 286.8 189.1 282.6 ;
      RECT  190.9 285.6 191.7 283.4 ;
      RECT  188.3 300.4 195.9 301.2 ;
      RECT  190.9 297.4 192.5 298.2 ;
      RECT  193.3 296.4 194.1 298.8 ;
      RECT  195.1 294.0 195.9 298.2 ;
      RECT  188.3 292.6 195.9 293.4 ;
      RECT  192.1 293.4 192.9 293.6 ;
      RECT  190.9 298.2 191.7 298.8 ;
      RECT  193.1 298.8 194.1 299.6 ;
      RECT  190.7 294.4 191.7 295.2 ;
      RECT  195.1 298.8 195.9 300.4 ;
      RECT  188.3 298.8 189.1 300.4 ;
      RECT  192.9 295.6 194.1 296.4 ;
      RECT  193.3 295.2 194.1 295.6 ;
      RECT  193.3 294.4 194.3 295.2 ;
      RECT  189.9 291.2 191.5 292.0 ;
      RECT  192.7 291.2 194.3 292.0 ;
      RECT  190.9 298.8 191.9 299.6 ;
      RECT  188.3 294.0 189.1 298.2 ;
      RECT  190.9 295.2 191.7 297.4 ;
      RECT  188.3 301.2 195.9 300.4 ;
      RECT  190.9 304.2 192.5 303.4 ;
      RECT  193.3 305.2 194.1 302.8 ;
      RECT  195.1 307.6 195.9 303.4 ;
      RECT  188.3 309.0 195.9 308.2 ;
      RECT  192.1 308.2 192.9 308.0 ;
      RECT  190.9 303.4 191.7 302.8 ;
      RECT  193.1 302.8 194.1 302.0 ;
      RECT  190.7 307.2 191.7 306.4 ;
      RECT  195.1 302.8 195.9 301.2 ;
      RECT  188.3 302.8 189.1 301.2 ;
      RECT  192.9 306.0 194.1 305.2 ;
      RECT  193.3 306.4 194.1 306.0 ;
      RECT  193.3 307.2 194.3 306.4 ;
      RECT  189.9 310.4 191.5 309.6 ;
      RECT  192.7 310.4 194.3 309.6 ;
      RECT  190.9 302.8 191.9 302.0 ;
      RECT  188.3 307.6 189.1 303.4 ;
      RECT  190.9 306.4 191.7 304.2 ;
      RECT  188.3 321.2 195.9 322.0 ;
      RECT  190.9 318.2 192.5 319.0 ;
      RECT  193.3 317.2 194.1 319.6 ;
      RECT  195.1 314.8 195.9 319.0 ;
      RECT  188.3 313.4 195.9 314.2 ;
      RECT  192.1 314.2 192.9 314.4 ;
      RECT  190.9 319.0 191.7 319.6 ;
      RECT  193.1 319.6 194.1 320.4 ;
      RECT  190.7 315.2 191.7 316.0 ;
      RECT  195.1 319.6 195.9 321.2 ;
      RECT  188.3 319.6 189.1 321.2 ;
      RECT  192.9 316.4 194.1 317.2 ;
      RECT  193.3 316.0 194.1 316.4 ;
      RECT  193.3 315.2 194.3 316.0 ;
      RECT  189.9 312.0 191.5 312.8 ;
      RECT  192.7 312.0 194.3 312.8 ;
      RECT  190.9 319.6 191.9 320.4 ;
      RECT  188.3 314.8 189.1 319.0 ;
      RECT  190.9 316.0 191.7 318.2 ;
      RECT  188.3 322.0 195.9 321.2 ;
      RECT  190.9 325.0 192.5 324.2 ;
      RECT  193.3 326.0 194.1 323.6 ;
      RECT  195.1 328.4 195.9 324.2 ;
      RECT  188.3 329.8 195.9 329.0 ;
      RECT  192.1 329.0 192.9 328.8 ;
      RECT  190.9 324.2 191.7 323.6 ;
      RECT  193.1 323.6 194.1 322.8 ;
      RECT  190.7 328.0 191.7 327.2 ;
      RECT  195.1 323.6 195.9 322.0 ;
      RECT  188.3 323.6 189.1 322.0 ;
      RECT  192.9 326.8 194.1 326.0 ;
      RECT  193.3 327.2 194.1 326.8 ;
      RECT  193.3 328.0 194.3 327.2 ;
      RECT  189.9 331.2 191.5 330.4 ;
      RECT  192.7 331.2 194.3 330.4 ;
      RECT  190.9 323.6 191.9 322.8 ;
      RECT  188.3 328.4 189.1 324.2 ;
      RECT  190.9 327.2 191.7 325.0 ;
      RECT  188.3 342.0 195.9 342.8 ;
      RECT  190.9 339.0 192.5 339.8 ;
      RECT  193.3 338.0 194.1 340.4 ;
      RECT  195.1 335.6 195.9 339.8 ;
      RECT  188.3 334.2 195.9 335.0 ;
      RECT  192.1 335.0 192.9 335.2 ;
      RECT  190.9 339.8 191.7 340.4 ;
      RECT  193.1 340.4 194.1 341.2 ;
      RECT  190.7 336.0 191.7 336.8 ;
      RECT  195.1 340.4 195.9 342.0 ;
      RECT  188.3 340.4 189.1 342.0 ;
      RECT  192.9 337.2 194.1 338.0 ;
      RECT  193.3 336.8 194.1 337.2 ;
      RECT  193.3 336.0 194.3 336.8 ;
      RECT  189.9 332.8 191.5 333.6 ;
      RECT  192.7 332.8 194.3 333.6 ;
      RECT  190.9 340.4 191.9 341.2 ;
      RECT  188.3 335.6 189.1 339.8 ;
      RECT  190.9 336.8 191.7 339.0 ;
      RECT  188.3 342.8 195.9 342.0 ;
      RECT  190.9 345.8 192.5 345.0 ;
      RECT  193.3 346.8 194.1 344.4 ;
      RECT  195.1 349.2 195.9 345.0 ;
      RECT  188.3 350.6 195.9 349.8 ;
      RECT  192.1 349.8 192.9 349.6 ;
      RECT  190.9 345.0 191.7 344.4 ;
      RECT  193.1 344.4 194.1 343.6 ;
      RECT  190.7 348.8 191.7 348.0 ;
      RECT  195.1 344.4 195.9 342.8 ;
      RECT  188.3 344.4 189.1 342.8 ;
      RECT  192.9 347.6 194.1 346.8 ;
      RECT  193.3 348.0 194.1 347.6 ;
      RECT  193.3 348.8 194.3 348.0 ;
      RECT  189.9 352.0 191.5 351.2 ;
      RECT  192.7 352.0 194.3 351.2 ;
      RECT  190.9 344.4 191.9 343.6 ;
      RECT  188.3 349.2 189.1 345.0 ;
      RECT  190.9 348.0 191.7 345.8 ;
      RECT  195.1 196.4 202.7 197.2 ;
      RECT  197.7 193.4 199.3 194.2 ;
      RECT  200.1 192.4 200.9 194.8 ;
      RECT  201.9 190.0 202.7 194.2 ;
      RECT  195.1 188.6 202.7 189.4 ;
      RECT  198.9 189.4 199.7 189.6 ;
      RECT  197.7 194.2 198.5 194.8 ;
      RECT  199.9 194.8 200.9 195.6 ;
      RECT  197.5 190.4 198.5 191.2 ;
      RECT  201.9 194.8 202.7 196.4 ;
      RECT  195.1 194.8 195.9 196.4 ;
      RECT  199.7 191.6 200.9 192.4 ;
      RECT  200.1 191.2 200.9 191.6 ;
      RECT  200.1 190.4 201.1 191.2 ;
      RECT  196.7 187.2 198.3 188.0 ;
      RECT  199.5 187.2 201.1 188.0 ;
      RECT  197.7 194.8 198.7 195.6 ;
      RECT  195.1 190.0 195.9 194.2 ;
      RECT  197.7 191.2 198.5 193.4 ;
      RECT  195.1 197.2 202.7 196.4 ;
      RECT  197.7 200.2 199.3 199.4 ;
      RECT  200.1 201.2 200.9 198.8 ;
      RECT  201.9 203.6 202.7 199.4 ;
      RECT  195.1 205.0 202.7 204.2 ;
      RECT  198.9 204.2 199.7 204.0 ;
      RECT  197.7 199.4 198.5 198.8 ;
      RECT  199.9 198.8 200.9 198.0 ;
      RECT  197.5 203.2 198.5 202.4 ;
      RECT  201.9 198.8 202.7 197.2 ;
      RECT  195.1 198.8 195.9 197.2 ;
      RECT  199.7 202.0 200.9 201.2 ;
      RECT  200.1 202.4 200.9 202.0 ;
      RECT  200.1 203.2 201.1 202.4 ;
      RECT  196.7 206.4 198.3 205.6 ;
      RECT  199.5 206.4 201.1 205.6 ;
      RECT  197.7 198.8 198.7 198.0 ;
      RECT  195.1 203.6 195.9 199.4 ;
      RECT  197.7 202.4 198.5 200.2 ;
      RECT  195.1 217.2 202.7 218.0 ;
      RECT  197.7 214.2 199.3 215.0 ;
      RECT  200.1 213.2 200.9 215.6 ;
      RECT  201.9 210.8 202.7 215.0 ;
      RECT  195.1 209.4 202.7 210.2 ;
      RECT  198.9 210.2 199.7 210.4 ;
      RECT  197.7 215.0 198.5 215.6 ;
      RECT  199.9 215.6 200.9 216.4 ;
      RECT  197.5 211.2 198.5 212.0 ;
      RECT  201.9 215.6 202.7 217.2 ;
      RECT  195.1 215.6 195.9 217.2 ;
      RECT  199.7 212.4 200.9 213.2 ;
      RECT  200.1 212.0 200.9 212.4 ;
      RECT  200.1 211.2 201.1 212.0 ;
      RECT  196.7 208.0 198.3 208.8 ;
      RECT  199.5 208.0 201.1 208.8 ;
      RECT  197.7 215.6 198.7 216.4 ;
      RECT  195.1 210.8 195.9 215.0 ;
      RECT  197.7 212.0 198.5 214.2 ;
      RECT  195.1 218.0 202.7 217.2 ;
      RECT  197.7 221.0 199.3 220.2 ;
      RECT  200.1 222.0 200.9 219.6 ;
      RECT  201.9 224.4 202.7 220.2 ;
      RECT  195.1 225.8 202.7 225.0 ;
      RECT  198.9 225.0 199.7 224.8 ;
      RECT  197.7 220.2 198.5 219.6 ;
      RECT  199.9 219.6 200.9 218.8 ;
      RECT  197.5 224.0 198.5 223.2 ;
      RECT  201.9 219.6 202.7 218.0 ;
      RECT  195.1 219.6 195.9 218.0 ;
      RECT  199.7 222.8 200.9 222.0 ;
      RECT  200.1 223.2 200.9 222.8 ;
      RECT  200.1 224.0 201.1 223.2 ;
      RECT  196.7 227.2 198.3 226.4 ;
      RECT  199.5 227.2 201.1 226.4 ;
      RECT  197.7 219.6 198.7 218.8 ;
      RECT  195.1 224.4 195.9 220.2 ;
      RECT  197.7 223.2 198.5 221.0 ;
      RECT  195.1 238.0 202.7 238.8 ;
      RECT  197.7 235.0 199.3 235.8 ;
      RECT  200.1 234.0 200.9 236.4 ;
      RECT  201.9 231.6 202.7 235.8 ;
      RECT  195.1 230.2 202.7 231.0 ;
      RECT  198.9 231.0 199.7 231.2 ;
      RECT  197.7 235.8 198.5 236.4 ;
      RECT  199.9 236.4 200.9 237.2 ;
      RECT  197.5 232.0 198.5 232.8 ;
      RECT  201.9 236.4 202.7 238.0 ;
      RECT  195.1 236.4 195.9 238.0 ;
      RECT  199.7 233.2 200.9 234.0 ;
      RECT  200.1 232.8 200.9 233.2 ;
      RECT  200.1 232.0 201.1 232.8 ;
      RECT  196.7 228.8 198.3 229.6 ;
      RECT  199.5 228.8 201.1 229.6 ;
      RECT  197.7 236.4 198.7 237.2 ;
      RECT  195.1 231.6 195.9 235.8 ;
      RECT  197.7 232.8 198.5 235.0 ;
      RECT  195.1 238.8 202.7 238.0 ;
      RECT  197.7 241.8 199.3 241.0 ;
      RECT  200.1 242.8 200.9 240.4 ;
      RECT  201.9 245.2 202.7 241.0 ;
      RECT  195.1 246.6 202.7 245.8 ;
      RECT  198.9 245.8 199.7 245.6 ;
      RECT  197.7 241.0 198.5 240.4 ;
      RECT  199.9 240.4 200.9 239.6 ;
      RECT  197.5 244.8 198.5 244.0 ;
      RECT  201.9 240.4 202.7 238.8 ;
      RECT  195.1 240.4 195.9 238.8 ;
      RECT  199.7 243.6 200.9 242.8 ;
      RECT  200.1 244.0 200.9 243.6 ;
      RECT  200.1 244.8 201.1 244.0 ;
      RECT  196.7 248.0 198.3 247.2 ;
      RECT  199.5 248.0 201.1 247.2 ;
      RECT  197.7 240.4 198.7 239.6 ;
      RECT  195.1 245.2 195.9 241.0 ;
      RECT  197.7 244.0 198.5 241.8 ;
      RECT  195.1 258.8 202.7 259.6 ;
      RECT  197.7 255.8 199.3 256.6 ;
      RECT  200.1 254.8 200.9 257.2 ;
      RECT  201.9 252.4 202.7 256.6 ;
      RECT  195.1 251.0 202.7 251.8 ;
      RECT  198.9 251.8 199.7 252.0 ;
      RECT  197.7 256.6 198.5 257.2 ;
      RECT  199.9 257.2 200.9 258.0 ;
      RECT  197.5 252.8 198.5 253.6 ;
      RECT  201.9 257.2 202.7 258.8 ;
      RECT  195.1 257.2 195.9 258.8 ;
      RECT  199.7 254.0 200.9 254.8 ;
      RECT  200.1 253.6 200.9 254.0 ;
      RECT  200.1 252.8 201.1 253.6 ;
      RECT  196.7 249.6 198.3 250.4 ;
      RECT  199.5 249.6 201.1 250.4 ;
      RECT  197.7 257.2 198.7 258.0 ;
      RECT  195.1 252.4 195.9 256.6 ;
      RECT  197.7 253.6 198.5 255.8 ;
      RECT  195.1 259.6 202.7 258.8 ;
      RECT  197.7 262.6 199.3 261.8 ;
      RECT  200.1 263.6 200.9 261.2 ;
      RECT  201.9 266.0 202.7 261.8 ;
      RECT  195.1 267.4 202.7 266.6 ;
      RECT  198.9 266.6 199.7 266.4 ;
      RECT  197.7 261.8 198.5 261.2 ;
      RECT  199.9 261.2 200.9 260.4 ;
      RECT  197.5 265.6 198.5 264.8 ;
      RECT  201.9 261.2 202.7 259.6 ;
      RECT  195.1 261.2 195.9 259.6 ;
      RECT  199.7 264.4 200.9 263.6 ;
      RECT  200.1 264.8 200.9 264.4 ;
      RECT  200.1 265.6 201.1 264.8 ;
      RECT  196.7 268.8 198.3 268.0 ;
      RECT  199.5 268.8 201.1 268.0 ;
      RECT  197.7 261.2 198.7 260.4 ;
      RECT  195.1 266.0 195.9 261.8 ;
      RECT  197.7 264.8 198.5 262.6 ;
      RECT  195.1 279.6 202.7 280.4 ;
      RECT  197.7 276.6 199.3 277.4 ;
      RECT  200.1 275.6 200.9 278.0 ;
      RECT  201.9 273.2 202.7 277.4 ;
      RECT  195.1 271.8 202.7 272.6 ;
      RECT  198.9 272.6 199.7 272.8 ;
      RECT  197.7 277.4 198.5 278.0 ;
      RECT  199.9 278.0 200.9 278.8 ;
      RECT  197.5 273.6 198.5 274.4 ;
      RECT  201.9 278.0 202.7 279.6 ;
      RECT  195.1 278.0 195.9 279.6 ;
      RECT  199.7 274.8 200.9 275.6 ;
      RECT  200.1 274.4 200.9 274.8 ;
      RECT  200.1 273.6 201.1 274.4 ;
      RECT  196.7 270.4 198.3 271.2 ;
      RECT  199.5 270.4 201.1 271.2 ;
      RECT  197.7 278.0 198.7 278.8 ;
      RECT  195.1 273.2 195.9 277.4 ;
      RECT  197.7 274.4 198.5 276.6 ;
      RECT  195.1 280.4 202.7 279.6 ;
      RECT  197.7 283.4 199.3 282.6 ;
      RECT  200.1 284.4 200.9 282.0 ;
      RECT  201.9 286.8 202.7 282.6 ;
      RECT  195.1 288.2 202.7 287.4 ;
      RECT  198.9 287.4 199.7 287.2 ;
      RECT  197.7 282.6 198.5 282.0 ;
      RECT  199.9 282.0 200.9 281.2 ;
      RECT  197.5 286.4 198.5 285.6 ;
      RECT  201.9 282.0 202.7 280.4 ;
      RECT  195.1 282.0 195.9 280.4 ;
      RECT  199.7 285.2 200.9 284.4 ;
      RECT  200.1 285.6 200.9 285.2 ;
      RECT  200.1 286.4 201.1 285.6 ;
      RECT  196.7 289.6 198.3 288.8 ;
      RECT  199.5 289.6 201.1 288.8 ;
      RECT  197.7 282.0 198.7 281.2 ;
      RECT  195.1 286.8 195.9 282.6 ;
      RECT  197.7 285.6 198.5 283.4 ;
      RECT  195.1 300.4 202.7 301.2 ;
      RECT  197.7 297.4 199.3 298.2 ;
      RECT  200.1 296.4 200.9 298.8 ;
      RECT  201.9 294.0 202.7 298.2 ;
      RECT  195.1 292.6 202.7 293.4 ;
      RECT  198.9 293.4 199.7 293.6 ;
      RECT  197.7 298.2 198.5 298.8 ;
      RECT  199.9 298.8 200.9 299.6 ;
      RECT  197.5 294.4 198.5 295.2 ;
      RECT  201.9 298.8 202.7 300.4 ;
      RECT  195.1 298.8 195.9 300.4 ;
      RECT  199.7 295.6 200.9 296.4 ;
      RECT  200.1 295.2 200.9 295.6 ;
      RECT  200.1 294.4 201.1 295.2 ;
      RECT  196.7 291.2 198.3 292.0 ;
      RECT  199.5 291.2 201.1 292.0 ;
      RECT  197.7 298.8 198.7 299.6 ;
      RECT  195.1 294.0 195.9 298.2 ;
      RECT  197.7 295.2 198.5 297.4 ;
      RECT  195.1 301.2 202.7 300.4 ;
      RECT  197.7 304.2 199.3 303.4 ;
      RECT  200.1 305.2 200.9 302.8 ;
      RECT  201.9 307.6 202.7 303.4 ;
      RECT  195.1 309.0 202.7 308.2 ;
      RECT  198.9 308.2 199.7 308.0 ;
      RECT  197.7 303.4 198.5 302.8 ;
      RECT  199.9 302.8 200.9 302.0 ;
      RECT  197.5 307.2 198.5 306.4 ;
      RECT  201.9 302.8 202.7 301.2 ;
      RECT  195.1 302.8 195.9 301.2 ;
      RECT  199.7 306.0 200.9 305.2 ;
      RECT  200.1 306.4 200.9 306.0 ;
      RECT  200.1 307.2 201.1 306.4 ;
      RECT  196.7 310.4 198.3 309.6 ;
      RECT  199.5 310.4 201.1 309.6 ;
      RECT  197.7 302.8 198.7 302.0 ;
      RECT  195.1 307.6 195.9 303.4 ;
      RECT  197.7 306.4 198.5 304.2 ;
      RECT  195.1 321.2 202.7 322.0 ;
      RECT  197.7 318.2 199.3 319.0 ;
      RECT  200.1 317.2 200.9 319.6 ;
      RECT  201.9 314.8 202.7 319.0 ;
      RECT  195.1 313.4 202.7 314.2 ;
      RECT  198.9 314.2 199.7 314.4 ;
      RECT  197.7 319.0 198.5 319.6 ;
      RECT  199.9 319.6 200.9 320.4 ;
      RECT  197.5 315.2 198.5 316.0 ;
      RECT  201.9 319.6 202.7 321.2 ;
      RECT  195.1 319.6 195.9 321.2 ;
      RECT  199.7 316.4 200.9 317.2 ;
      RECT  200.1 316.0 200.9 316.4 ;
      RECT  200.1 315.2 201.1 316.0 ;
      RECT  196.7 312.0 198.3 312.8 ;
      RECT  199.5 312.0 201.1 312.8 ;
      RECT  197.7 319.6 198.7 320.4 ;
      RECT  195.1 314.8 195.9 319.0 ;
      RECT  197.7 316.0 198.5 318.2 ;
      RECT  195.1 322.0 202.7 321.2 ;
      RECT  197.7 325.0 199.3 324.2 ;
      RECT  200.1 326.0 200.9 323.6 ;
      RECT  201.9 328.4 202.7 324.2 ;
      RECT  195.1 329.8 202.7 329.0 ;
      RECT  198.9 329.0 199.7 328.8 ;
      RECT  197.7 324.2 198.5 323.6 ;
      RECT  199.9 323.6 200.9 322.8 ;
      RECT  197.5 328.0 198.5 327.2 ;
      RECT  201.9 323.6 202.7 322.0 ;
      RECT  195.1 323.6 195.9 322.0 ;
      RECT  199.7 326.8 200.9 326.0 ;
      RECT  200.1 327.2 200.9 326.8 ;
      RECT  200.1 328.0 201.1 327.2 ;
      RECT  196.7 331.2 198.3 330.4 ;
      RECT  199.5 331.2 201.1 330.4 ;
      RECT  197.7 323.6 198.7 322.8 ;
      RECT  195.1 328.4 195.9 324.2 ;
      RECT  197.7 327.2 198.5 325.0 ;
      RECT  195.1 342.0 202.7 342.8 ;
      RECT  197.7 339.0 199.3 339.8 ;
      RECT  200.1 338.0 200.9 340.4 ;
      RECT  201.9 335.6 202.7 339.8 ;
      RECT  195.1 334.2 202.7 335.0 ;
      RECT  198.9 335.0 199.7 335.2 ;
      RECT  197.7 339.8 198.5 340.4 ;
      RECT  199.9 340.4 200.9 341.2 ;
      RECT  197.5 336.0 198.5 336.8 ;
      RECT  201.9 340.4 202.7 342.0 ;
      RECT  195.1 340.4 195.9 342.0 ;
      RECT  199.7 337.2 200.9 338.0 ;
      RECT  200.1 336.8 200.9 337.2 ;
      RECT  200.1 336.0 201.1 336.8 ;
      RECT  196.7 332.8 198.3 333.6 ;
      RECT  199.5 332.8 201.1 333.6 ;
      RECT  197.7 340.4 198.7 341.2 ;
      RECT  195.1 335.6 195.9 339.8 ;
      RECT  197.7 336.8 198.5 339.0 ;
      RECT  195.1 342.8 202.7 342.0 ;
      RECT  197.7 345.8 199.3 345.0 ;
      RECT  200.1 346.8 200.9 344.4 ;
      RECT  201.9 349.2 202.7 345.0 ;
      RECT  195.1 350.6 202.7 349.8 ;
      RECT  198.9 349.8 199.7 349.6 ;
      RECT  197.7 345.0 198.5 344.4 ;
      RECT  199.9 344.4 200.9 343.6 ;
      RECT  197.5 348.8 198.5 348.0 ;
      RECT  201.9 344.4 202.7 342.8 ;
      RECT  195.1 344.4 195.9 342.8 ;
      RECT  199.7 347.6 200.9 346.8 ;
      RECT  200.1 348.0 200.9 347.6 ;
      RECT  200.1 348.8 201.1 348.0 ;
      RECT  196.7 352.0 198.3 351.2 ;
      RECT  199.5 352.0 201.1 351.2 ;
      RECT  197.7 344.4 198.7 343.6 ;
      RECT  195.1 349.2 195.9 345.0 ;
      RECT  197.7 348.0 198.5 345.8 ;
      RECT  188.7 188.6 202.3 189.4 ;
      RECT  188.7 204.2 202.3 205.0 ;
      RECT  188.7 209.4 202.3 210.2 ;
      RECT  188.7 225.0 202.3 225.8 ;
      RECT  188.7 230.2 202.3 231.0 ;
      RECT  188.7 245.8 202.3 246.6 ;
      RECT  188.7 251.0 202.3 251.8 ;
      RECT  188.7 266.6 202.3 267.4 ;
      RECT  188.7 271.8 202.3 272.6 ;
      RECT  188.7 287.4 202.3 288.2 ;
      RECT  188.7 292.6 202.3 293.4 ;
      RECT  188.7 308.2 202.3 309.0 ;
      RECT  188.7 313.4 202.3 314.2 ;
      RECT  188.7 329.0 202.3 329.8 ;
      RECT  188.7 334.2 202.3 335.0 ;
      RECT  188.7 349.8 202.3 350.6 ;
      RECT  181.5 175.6 189.1 176.4 ;
      RECT  184.1 172.6 185.7 173.4 ;
      RECT  186.5 171.6 187.3 174.0 ;
      RECT  188.3 169.2 189.1 173.4 ;
      RECT  181.5 167.8 189.1 168.6 ;
      RECT  185.3 168.6 186.1 168.8 ;
      RECT  184.1 173.4 184.9 174.0 ;
      RECT  186.3 174.0 187.3 174.8 ;
      RECT  183.9 169.6 184.9 170.4 ;
      RECT  188.3 174.0 189.1 175.6 ;
      RECT  181.5 174.0 182.3 175.6 ;
      RECT  186.1 170.8 187.3 171.6 ;
      RECT  186.5 170.4 187.3 170.8 ;
      RECT  186.5 169.6 187.5 170.4 ;
      RECT  183.9 166.4 184.7 167.2 ;
      RECT  186.7 166.4 187.5 167.2 ;
      RECT  184.1 174.0 185.1 174.8 ;
      RECT  181.5 169.2 182.3 173.4 ;
      RECT  184.1 170.4 184.9 172.6 ;
      RECT  181.5 176.4 189.1 175.6 ;
      RECT  184.1 179.4 185.7 178.6 ;
      RECT  186.5 180.4 187.3 178.0 ;
      RECT  188.3 182.8 189.1 178.6 ;
      RECT  181.5 184.2 189.1 183.4 ;
      RECT  185.3 183.4 186.1 183.2 ;
      RECT  184.1 178.6 184.9 178.0 ;
      RECT  186.3 178.0 187.3 177.2 ;
      RECT  183.9 182.4 184.9 181.6 ;
      RECT  186.3 177.2 187.1 176.4 ;
      RECT  181.5 178.0 182.3 176.4 ;
      RECT  188.3 178.0 189.1 176.4 ;
      RECT  186.1 181.2 187.3 180.4 ;
      RECT  186.5 181.6 187.3 181.2 ;
      RECT  186.5 182.4 187.5 181.6 ;
      RECT  183.1 185.6 184.7 184.8 ;
      RECT  185.9 185.6 187.5 184.8 ;
      RECT  184.1 178.0 185.1 177.2 ;
      RECT  181.5 182.8 182.3 178.6 ;
      RECT  184.1 181.6 184.9 179.4 ;
      RECT  181.5 196.4 189.1 197.2 ;
      RECT  184.1 193.4 185.7 194.2 ;
      RECT  186.5 192.4 187.3 194.8 ;
      RECT  188.3 190.0 189.1 194.2 ;
      RECT  181.5 188.6 189.1 189.4 ;
      RECT  185.3 189.4 186.1 189.6 ;
      RECT  184.1 194.2 184.9 194.8 ;
      RECT  186.3 194.8 187.3 195.6 ;
      RECT  183.9 190.4 184.9 191.2 ;
      RECT  186.3 195.6 187.1 196.4 ;
      RECT  181.5 194.8 182.3 196.4 ;
      RECT  188.3 194.8 189.1 196.4 ;
      RECT  186.1 191.6 187.3 192.4 ;
      RECT  186.5 191.2 187.3 191.6 ;
      RECT  186.5 190.4 187.5 191.2 ;
      RECT  183.1 187.2 184.7 188.0 ;
      RECT  185.9 187.2 187.5 188.0 ;
      RECT  184.1 194.8 185.1 195.6 ;
      RECT  181.5 190.0 182.3 194.2 ;
      RECT  184.1 191.2 184.9 193.4 ;
      RECT  181.5 197.2 189.1 196.4 ;
      RECT  184.1 200.2 185.7 199.4 ;
      RECT  186.5 201.2 187.3 198.8 ;
      RECT  188.3 203.6 189.1 199.4 ;
      RECT  181.5 205.0 189.1 204.2 ;
      RECT  185.3 204.2 186.1 204.0 ;
      RECT  184.1 199.4 184.9 198.8 ;
      RECT  186.3 198.8 187.3 198.0 ;
      RECT  183.9 203.2 184.9 202.4 ;
      RECT  186.3 198.0 187.1 197.2 ;
      RECT  181.5 198.8 182.3 197.2 ;
      RECT  188.3 198.8 189.1 197.2 ;
      RECT  186.1 202.0 187.3 201.2 ;
      RECT  186.5 202.4 187.3 202.0 ;
      RECT  186.5 203.2 187.5 202.4 ;
      RECT  183.1 206.4 184.7 205.6 ;
      RECT  185.9 206.4 187.5 205.6 ;
      RECT  184.1 198.8 185.1 198.0 ;
      RECT  181.5 203.6 182.3 199.4 ;
      RECT  184.1 202.4 184.9 200.2 ;
      RECT  181.5 217.2 189.1 218.0 ;
      RECT  184.1 214.2 185.7 215.0 ;
      RECT  186.5 213.2 187.3 215.6 ;
      RECT  188.3 210.8 189.1 215.0 ;
      RECT  181.5 209.4 189.1 210.2 ;
      RECT  185.3 210.2 186.1 210.4 ;
      RECT  184.1 215.0 184.9 215.6 ;
      RECT  186.3 215.6 187.3 216.4 ;
      RECT  183.9 211.2 184.9 212.0 ;
      RECT  186.3 216.4 187.1 217.2 ;
      RECT  181.5 215.6 182.3 217.2 ;
      RECT  188.3 215.6 189.1 217.2 ;
      RECT  186.1 212.4 187.3 213.2 ;
      RECT  186.5 212.0 187.3 212.4 ;
      RECT  186.5 211.2 187.5 212.0 ;
      RECT  183.1 208.0 184.7 208.8 ;
      RECT  185.9 208.0 187.5 208.8 ;
      RECT  184.1 215.6 185.1 216.4 ;
      RECT  181.5 210.8 182.3 215.0 ;
      RECT  184.1 212.0 184.9 214.2 ;
      RECT  181.5 218.0 189.1 217.2 ;
      RECT  184.1 221.0 185.7 220.2 ;
      RECT  186.5 222.0 187.3 219.6 ;
      RECT  188.3 224.4 189.1 220.2 ;
      RECT  181.5 225.8 189.1 225.0 ;
      RECT  185.3 225.0 186.1 224.8 ;
      RECT  184.1 220.2 184.9 219.6 ;
      RECT  186.3 219.6 187.3 218.8 ;
      RECT  183.9 224.0 184.9 223.2 ;
      RECT  186.3 218.8 187.1 218.0 ;
      RECT  181.5 219.6 182.3 218.0 ;
      RECT  188.3 219.6 189.1 218.0 ;
      RECT  186.1 222.8 187.3 222.0 ;
      RECT  186.5 223.2 187.3 222.8 ;
      RECT  186.5 224.0 187.5 223.2 ;
      RECT  183.1 227.2 184.7 226.4 ;
      RECT  185.9 227.2 187.5 226.4 ;
      RECT  184.1 219.6 185.1 218.8 ;
      RECT  181.5 224.4 182.3 220.2 ;
      RECT  184.1 223.2 184.9 221.0 ;
      RECT  181.5 238.0 189.1 238.8 ;
      RECT  184.1 235.0 185.7 235.8 ;
      RECT  186.5 234.0 187.3 236.4 ;
      RECT  188.3 231.6 189.1 235.8 ;
      RECT  181.5 230.2 189.1 231.0 ;
      RECT  185.3 231.0 186.1 231.2 ;
      RECT  184.1 235.8 184.9 236.4 ;
      RECT  186.3 236.4 187.3 237.2 ;
      RECT  183.9 232.0 184.9 232.8 ;
      RECT  186.3 237.2 187.1 238.0 ;
      RECT  181.5 236.4 182.3 238.0 ;
      RECT  188.3 236.4 189.1 238.0 ;
      RECT  186.1 233.2 187.3 234.0 ;
      RECT  186.5 232.8 187.3 233.2 ;
      RECT  186.5 232.0 187.5 232.8 ;
      RECT  183.1 228.8 184.7 229.6 ;
      RECT  185.9 228.8 187.5 229.6 ;
      RECT  184.1 236.4 185.1 237.2 ;
      RECT  181.5 231.6 182.3 235.8 ;
      RECT  184.1 232.8 184.9 235.0 ;
      RECT  181.5 238.8 189.1 238.0 ;
      RECT  184.1 241.8 185.7 241.0 ;
      RECT  186.5 242.8 187.3 240.4 ;
      RECT  188.3 245.2 189.1 241.0 ;
      RECT  181.5 246.6 189.1 245.8 ;
      RECT  185.3 245.8 186.1 245.6 ;
      RECT  184.1 241.0 184.9 240.4 ;
      RECT  186.3 240.4 187.3 239.6 ;
      RECT  183.9 244.8 184.9 244.0 ;
      RECT  186.3 239.6 187.1 238.8 ;
      RECT  181.5 240.4 182.3 238.8 ;
      RECT  188.3 240.4 189.1 238.8 ;
      RECT  186.1 243.6 187.3 242.8 ;
      RECT  186.5 244.0 187.3 243.6 ;
      RECT  186.5 244.8 187.5 244.0 ;
      RECT  183.1 248.0 184.7 247.2 ;
      RECT  185.9 248.0 187.5 247.2 ;
      RECT  184.1 240.4 185.1 239.6 ;
      RECT  181.5 245.2 182.3 241.0 ;
      RECT  184.1 244.0 184.9 241.8 ;
      RECT  181.5 258.8 189.1 259.6 ;
      RECT  184.1 255.8 185.7 256.6 ;
      RECT  186.5 254.8 187.3 257.2 ;
      RECT  188.3 252.4 189.1 256.6 ;
      RECT  181.5 251.0 189.1 251.8 ;
      RECT  185.3 251.8 186.1 252.0 ;
      RECT  184.1 256.6 184.9 257.2 ;
      RECT  186.3 257.2 187.3 258.0 ;
      RECT  183.9 252.8 184.9 253.6 ;
      RECT  186.3 258.0 187.1 258.8 ;
      RECT  181.5 257.2 182.3 258.8 ;
      RECT  188.3 257.2 189.1 258.8 ;
      RECT  186.1 254.0 187.3 254.8 ;
      RECT  186.5 253.6 187.3 254.0 ;
      RECT  186.5 252.8 187.5 253.6 ;
      RECT  183.1 249.6 184.7 250.4 ;
      RECT  185.9 249.6 187.5 250.4 ;
      RECT  184.1 257.2 185.1 258.0 ;
      RECT  181.5 252.4 182.3 256.6 ;
      RECT  184.1 253.6 184.9 255.8 ;
      RECT  181.5 259.6 189.1 258.8 ;
      RECT  184.1 262.6 185.7 261.8 ;
      RECT  186.5 263.6 187.3 261.2 ;
      RECT  188.3 266.0 189.1 261.8 ;
      RECT  181.5 267.4 189.1 266.6 ;
      RECT  185.3 266.6 186.1 266.4 ;
      RECT  184.1 261.8 184.9 261.2 ;
      RECT  186.3 261.2 187.3 260.4 ;
      RECT  183.9 265.6 184.9 264.8 ;
      RECT  186.3 260.4 187.1 259.6 ;
      RECT  181.5 261.2 182.3 259.6 ;
      RECT  188.3 261.2 189.1 259.6 ;
      RECT  186.1 264.4 187.3 263.6 ;
      RECT  186.5 264.8 187.3 264.4 ;
      RECT  186.5 265.6 187.5 264.8 ;
      RECT  183.1 268.8 184.7 268.0 ;
      RECT  185.9 268.8 187.5 268.0 ;
      RECT  184.1 261.2 185.1 260.4 ;
      RECT  181.5 266.0 182.3 261.8 ;
      RECT  184.1 264.8 184.9 262.6 ;
      RECT  181.5 279.6 189.1 280.4 ;
      RECT  184.1 276.6 185.7 277.4 ;
      RECT  186.5 275.6 187.3 278.0 ;
      RECT  188.3 273.2 189.1 277.4 ;
      RECT  181.5 271.8 189.1 272.6 ;
      RECT  185.3 272.6 186.1 272.8 ;
      RECT  184.1 277.4 184.9 278.0 ;
      RECT  186.3 278.0 187.3 278.8 ;
      RECT  183.9 273.6 184.9 274.4 ;
      RECT  186.3 278.8 187.1 279.6 ;
      RECT  181.5 278.0 182.3 279.6 ;
      RECT  188.3 278.0 189.1 279.6 ;
      RECT  186.1 274.8 187.3 275.6 ;
      RECT  186.5 274.4 187.3 274.8 ;
      RECT  186.5 273.6 187.5 274.4 ;
      RECT  183.1 270.4 184.7 271.2 ;
      RECT  185.9 270.4 187.5 271.2 ;
      RECT  184.1 278.0 185.1 278.8 ;
      RECT  181.5 273.2 182.3 277.4 ;
      RECT  184.1 274.4 184.9 276.6 ;
      RECT  181.5 280.4 189.1 279.6 ;
      RECT  184.1 283.4 185.7 282.6 ;
      RECT  186.5 284.4 187.3 282.0 ;
      RECT  188.3 286.8 189.1 282.6 ;
      RECT  181.5 288.2 189.1 287.4 ;
      RECT  185.3 287.4 186.1 287.2 ;
      RECT  184.1 282.6 184.9 282.0 ;
      RECT  186.3 282.0 187.3 281.2 ;
      RECT  183.9 286.4 184.9 285.6 ;
      RECT  186.3 281.2 187.1 280.4 ;
      RECT  181.5 282.0 182.3 280.4 ;
      RECT  188.3 282.0 189.1 280.4 ;
      RECT  186.1 285.2 187.3 284.4 ;
      RECT  186.5 285.6 187.3 285.2 ;
      RECT  186.5 286.4 187.5 285.6 ;
      RECT  183.1 289.6 184.7 288.8 ;
      RECT  185.9 289.6 187.5 288.8 ;
      RECT  184.1 282.0 185.1 281.2 ;
      RECT  181.5 286.8 182.3 282.6 ;
      RECT  184.1 285.6 184.9 283.4 ;
      RECT  181.5 300.4 189.1 301.2 ;
      RECT  184.1 297.4 185.7 298.2 ;
      RECT  186.5 296.4 187.3 298.8 ;
      RECT  188.3 294.0 189.1 298.2 ;
      RECT  181.5 292.6 189.1 293.4 ;
      RECT  185.3 293.4 186.1 293.6 ;
      RECT  184.1 298.2 184.9 298.8 ;
      RECT  186.3 298.8 187.3 299.6 ;
      RECT  183.9 294.4 184.9 295.2 ;
      RECT  186.3 299.6 187.1 300.4 ;
      RECT  181.5 298.8 182.3 300.4 ;
      RECT  188.3 298.8 189.1 300.4 ;
      RECT  186.1 295.6 187.3 296.4 ;
      RECT  186.5 295.2 187.3 295.6 ;
      RECT  186.5 294.4 187.5 295.2 ;
      RECT  183.1 291.2 184.7 292.0 ;
      RECT  185.9 291.2 187.5 292.0 ;
      RECT  184.1 298.8 185.1 299.6 ;
      RECT  181.5 294.0 182.3 298.2 ;
      RECT  184.1 295.2 184.9 297.4 ;
      RECT  181.5 301.2 189.1 300.4 ;
      RECT  184.1 304.2 185.7 303.4 ;
      RECT  186.5 305.2 187.3 302.8 ;
      RECT  188.3 307.6 189.1 303.4 ;
      RECT  181.5 309.0 189.1 308.2 ;
      RECT  185.3 308.2 186.1 308.0 ;
      RECT  184.1 303.4 184.9 302.8 ;
      RECT  186.3 302.8 187.3 302.0 ;
      RECT  183.9 307.2 184.9 306.4 ;
      RECT  186.3 302.0 187.1 301.2 ;
      RECT  181.5 302.8 182.3 301.2 ;
      RECT  188.3 302.8 189.1 301.2 ;
      RECT  186.1 306.0 187.3 305.2 ;
      RECT  186.5 306.4 187.3 306.0 ;
      RECT  186.5 307.2 187.5 306.4 ;
      RECT  183.1 310.4 184.7 309.6 ;
      RECT  185.9 310.4 187.5 309.6 ;
      RECT  184.1 302.8 185.1 302.0 ;
      RECT  181.5 307.6 182.3 303.4 ;
      RECT  184.1 306.4 184.9 304.2 ;
      RECT  181.5 321.2 189.1 322.0 ;
      RECT  184.1 318.2 185.7 319.0 ;
      RECT  186.5 317.2 187.3 319.6 ;
      RECT  188.3 314.8 189.1 319.0 ;
      RECT  181.5 313.4 189.1 314.2 ;
      RECT  185.3 314.2 186.1 314.4 ;
      RECT  184.1 319.0 184.9 319.6 ;
      RECT  186.3 319.6 187.3 320.4 ;
      RECT  183.9 315.2 184.9 316.0 ;
      RECT  186.3 320.4 187.1 321.2 ;
      RECT  181.5 319.6 182.3 321.2 ;
      RECT  188.3 319.6 189.1 321.2 ;
      RECT  186.1 316.4 187.3 317.2 ;
      RECT  186.5 316.0 187.3 316.4 ;
      RECT  186.5 315.2 187.5 316.0 ;
      RECT  183.1 312.0 184.7 312.8 ;
      RECT  185.9 312.0 187.5 312.8 ;
      RECT  184.1 319.6 185.1 320.4 ;
      RECT  181.5 314.8 182.3 319.0 ;
      RECT  184.1 316.0 184.9 318.2 ;
      RECT  181.5 322.0 189.1 321.2 ;
      RECT  184.1 325.0 185.7 324.2 ;
      RECT  186.5 326.0 187.3 323.6 ;
      RECT  188.3 328.4 189.1 324.2 ;
      RECT  181.5 329.8 189.1 329.0 ;
      RECT  185.3 329.0 186.1 328.8 ;
      RECT  184.1 324.2 184.9 323.6 ;
      RECT  186.3 323.6 187.3 322.8 ;
      RECT  183.9 328.0 184.9 327.2 ;
      RECT  186.3 322.8 187.1 322.0 ;
      RECT  181.5 323.6 182.3 322.0 ;
      RECT  188.3 323.6 189.1 322.0 ;
      RECT  186.1 326.8 187.3 326.0 ;
      RECT  186.5 327.2 187.3 326.8 ;
      RECT  186.5 328.0 187.5 327.2 ;
      RECT  183.1 331.2 184.7 330.4 ;
      RECT  185.9 331.2 187.5 330.4 ;
      RECT  184.1 323.6 185.1 322.8 ;
      RECT  181.5 328.4 182.3 324.2 ;
      RECT  184.1 327.2 184.9 325.0 ;
      RECT  181.5 342.0 189.1 342.8 ;
      RECT  184.1 339.0 185.7 339.8 ;
      RECT  186.5 338.0 187.3 340.4 ;
      RECT  188.3 335.6 189.1 339.8 ;
      RECT  181.5 334.2 189.1 335.0 ;
      RECT  185.3 335.0 186.1 335.2 ;
      RECT  184.1 339.8 184.9 340.4 ;
      RECT  186.3 340.4 187.3 341.2 ;
      RECT  183.9 336.0 184.9 336.8 ;
      RECT  186.3 341.2 187.1 342.0 ;
      RECT  181.5 340.4 182.3 342.0 ;
      RECT  188.3 340.4 189.1 342.0 ;
      RECT  186.1 337.2 187.3 338.0 ;
      RECT  186.5 336.8 187.3 337.2 ;
      RECT  186.5 336.0 187.5 336.8 ;
      RECT  183.1 332.8 184.7 333.6 ;
      RECT  185.9 332.8 187.5 333.6 ;
      RECT  184.1 340.4 185.1 341.2 ;
      RECT  181.5 335.6 182.3 339.8 ;
      RECT  184.1 336.8 184.9 339.0 ;
      RECT  181.5 342.8 189.1 342.0 ;
      RECT  184.1 345.8 185.7 345.0 ;
      RECT  186.5 346.8 187.3 344.4 ;
      RECT  188.3 349.2 189.1 345.0 ;
      RECT  181.5 350.6 189.1 349.8 ;
      RECT  185.3 349.8 186.1 349.6 ;
      RECT  184.1 345.0 184.9 344.4 ;
      RECT  186.3 344.4 187.3 343.6 ;
      RECT  183.9 348.8 184.9 348.0 ;
      RECT  186.3 343.6 187.1 342.8 ;
      RECT  181.5 344.4 182.3 342.8 ;
      RECT  188.3 344.4 189.1 342.8 ;
      RECT  186.1 347.6 187.3 346.8 ;
      RECT  186.5 348.0 187.3 347.6 ;
      RECT  186.5 348.8 187.5 348.0 ;
      RECT  183.1 352.0 184.7 351.2 ;
      RECT  185.9 352.0 187.5 351.2 ;
      RECT  184.1 344.4 185.1 343.6 ;
      RECT  181.5 349.2 182.3 345.0 ;
      RECT  184.1 348.0 184.9 345.8 ;
      RECT  181.5 362.8 189.1 363.6 ;
      RECT  184.1 359.8 185.7 360.6 ;
      RECT  186.5 358.8 187.3 361.2 ;
      RECT  188.3 356.4 189.1 360.6 ;
      RECT  181.5 355.0 189.1 355.8 ;
      RECT  185.3 355.8 186.1 356.0 ;
      RECT  184.1 360.6 184.9 361.2 ;
      RECT  186.3 361.2 187.3 362.0 ;
      RECT  183.9 356.8 184.9 357.6 ;
      RECT  188.3 361.2 189.1 362.8 ;
      RECT  181.5 361.2 182.3 362.8 ;
      RECT  186.1 358.0 187.3 358.8 ;
      RECT  186.5 357.6 187.3 358.0 ;
      RECT  186.5 356.8 187.5 357.6 ;
      RECT  183.9 353.6 184.7 354.4 ;
      RECT  186.7 353.6 187.5 354.4 ;
      RECT  184.1 361.2 185.1 362.0 ;
      RECT  181.5 356.4 182.3 360.6 ;
      RECT  184.1 357.6 184.9 359.8 ;
      RECT  181.9 167.8 188.7 168.6 ;
      RECT  181.9 183.4 188.7 184.2 ;
      RECT  181.9 188.6 188.7 189.4 ;
      RECT  181.9 204.2 188.7 205.0 ;
      RECT  181.9 209.4 188.7 210.2 ;
      RECT  181.9 225.0 188.7 225.8 ;
      RECT  181.9 230.2 188.7 231.0 ;
      RECT  181.9 245.8 188.7 246.6 ;
      RECT  181.9 251.0 188.7 251.8 ;
      RECT  181.9 266.6 188.7 267.4 ;
      RECT  181.9 271.8 188.7 272.6 ;
      RECT  181.9 287.4 188.7 288.2 ;
      RECT  181.9 292.6 188.7 293.4 ;
      RECT  181.9 308.2 188.7 309.0 ;
      RECT  181.9 313.4 188.7 314.2 ;
      RECT  181.9 329.0 188.7 329.8 ;
      RECT  181.9 334.2 188.7 335.0 ;
      RECT  181.9 349.8 188.7 350.6 ;
      RECT  181.9 355.0 188.7 355.8 ;
      RECT  188.3 176.4 195.9 175.6 ;
      RECT  190.9 179.4 192.5 178.6 ;
      RECT  193.3 180.4 194.1 178.0 ;
      RECT  195.1 182.8 195.9 178.6 ;
      RECT  188.3 184.2 195.9 183.4 ;
      RECT  192.1 183.4 192.9 183.2 ;
      RECT  190.9 178.6 191.7 178.0 ;
      RECT  193.1 178.0 194.1 177.2 ;
      RECT  190.7 182.4 191.7 181.6 ;
      RECT  195.1 178.0 195.9 176.4 ;
      RECT  188.3 178.0 189.1 176.4 ;
      RECT  192.9 181.2 194.1 180.4 ;
      RECT  193.3 181.6 194.1 181.2 ;
      RECT  193.3 182.4 194.3 181.6 ;
      RECT  190.7 185.6 191.5 184.8 ;
      RECT  193.5 185.6 194.3 184.8 ;
      RECT  190.9 178.0 191.9 177.2 ;
      RECT  188.3 182.8 189.1 178.6 ;
      RECT  190.9 181.6 191.7 179.4 ;
      RECT  195.1 176.4 202.7 175.6 ;
      RECT  197.7 179.4 199.3 178.6 ;
      RECT  200.1 180.4 200.9 178.0 ;
      RECT  201.9 182.8 202.7 178.6 ;
      RECT  195.1 184.2 202.7 183.4 ;
      RECT  198.9 183.4 199.7 183.2 ;
      RECT  197.7 178.6 198.5 178.0 ;
      RECT  199.9 178.0 200.9 177.2 ;
      RECT  197.5 182.4 198.5 181.6 ;
      RECT  201.9 178.0 202.7 176.4 ;
      RECT  195.1 178.0 195.9 176.4 ;
      RECT  199.7 181.2 200.9 180.4 ;
      RECT  200.1 181.6 200.9 181.2 ;
      RECT  200.1 182.4 201.1 181.6 ;
      RECT  197.5 185.6 198.3 184.8 ;
      RECT  200.3 185.6 201.1 184.8 ;
      RECT  197.7 178.0 198.7 177.2 ;
      RECT  195.1 182.8 195.9 178.6 ;
      RECT  197.7 181.6 198.5 179.4 ;
      RECT  188.7 184.2 202.3 183.4 ;
      RECT  188.3 175.6 195.9 176.4 ;
      RECT  190.9 172.6 192.5 173.4 ;
      RECT  193.3 171.6 194.1 174.0 ;
      RECT  195.1 169.2 195.9 173.4 ;
      RECT  188.3 167.8 195.9 168.6 ;
      RECT  192.1 168.6 192.9 168.8 ;
      RECT  190.9 173.4 191.7 174.0 ;
      RECT  193.1 174.0 194.1 174.8 ;
      RECT  190.7 169.6 191.7 170.4 ;
      RECT  195.1 174.0 195.9 175.6 ;
      RECT  188.3 174.0 189.1 175.6 ;
      RECT  192.9 170.8 194.1 171.6 ;
      RECT  193.3 170.4 194.1 170.8 ;
      RECT  193.3 169.6 194.3 170.4 ;
      RECT  190.7 166.4 191.5 167.2 ;
      RECT  193.5 166.4 194.3 167.2 ;
      RECT  190.9 174.0 191.9 174.8 ;
      RECT  188.3 169.2 189.1 173.4 ;
      RECT  190.9 170.4 191.7 172.6 ;
      RECT  195.1 175.6 202.7 176.4 ;
      RECT  197.7 172.6 199.3 173.4 ;
      RECT  200.1 171.6 200.9 174.0 ;
      RECT  201.9 169.2 202.7 173.4 ;
      RECT  195.1 167.8 202.7 168.6 ;
      RECT  198.9 168.6 199.7 168.8 ;
      RECT  197.7 173.4 198.5 174.0 ;
      RECT  199.9 174.0 200.9 174.8 ;
      RECT  197.5 169.6 198.5 170.4 ;
      RECT  201.9 174.0 202.7 175.6 ;
      RECT  195.1 174.0 195.9 175.6 ;
      RECT  199.7 170.8 200.9 171.6 ;
      RECT  200.1 170.4 200.9 170.8 ;
      RECT  200.1 169.6 201.1 170.4 ;
      RECT  197.5 166.4 198.3 167.2 ;
      RECT  200.3 166.4 201.1 167.2 ;
      RECT  197.7 174.0 198.7 174.8 ;
      RECT  195.1 169.2 195.9 173.4 ;
      RECT  197.7 170.4 198.5 172.6 ;
      RECT  188.7 167.8 202.3 168.6 ;
      RECT  188.3 362.8 195.9 363.6 ;
      RECT  190.9 359.8 192.5 360.6 ;
      RECT  193.3 358.8 194.1 361.2 ;
      RECT  195.1 356.4 195.9 360.6 ;
      RECT  188.3 355.0 195.9 355.8 ;
      RECT  192.1 355.8 192.9 356.0 ;
      RECT  190.9 360.6 191.7 361.2 ;
      RECT  193.1 361.2 194.1 362.0 ;
      RECT  190.7 356.8 191.7 357.6 ;
      RECT  195.1 361.2 195.9 362.8 ;
      RECT  188.3 361.2 189.1 362.8 ;
      RECT  192.9 358.0 194.1 358.8 ;
      RECT  193.3 357.6 194.1 358.0 ;
      RECT  193.3 356.8 194.3 357.6 ;
      RECT  190.7 353.6 191.5 354.4 ;
      RECT  193.5 353.6 194.3 354.4 ;
      RECT  190.9 361.2 191.9 362.0 ;
      RECT  188.3 356.4 189.1 360.6 ;
      RECT  190.9 357.6 191.7 359.8 ;
      RECT  195.1 362.8 202.7 363.6 ;
      RECT  197.7 359.8 199.3 360.6 ;
      RECT  200.1 358.8 200.9 361.2 ;
      RECT  201.9 356.4 202.7 360.6 ;
      RECT  195.1 355.0 202.7 355.8 ;
      RECT  198.9 355.8 199.7 356.0 ;
      RECT  197.7 360.6 198.5 361.2 ;
      RECT  199.9 361.2 200.9 362.0 ;
      RECT  197.5 356.8 198.5 357.6 ;
      RECT  201.9 361.2 202.7 362.8 ;
      RECT  195.1 361.2 195.9 362.8 ;
      RECT  199.7 358.0 200.9 358.8 ;
      RECT  200.1 357.6 200.9 358.0 ;
      RECT  200.1 356.8 201.1 357.6 ;
      RECT  197.5 353.6 198.3 354.4 ;
      RECT  200.3 353.6 201.1 354.4 ;
      RECT  197.7 361.2 198.7 362.0 ;
      RECT  195.1 356.4 195.9 360.6 ;
      RECT  197.7 357.6 198.5 359.8 ;
      RECT  188.7 355.0 202.3 355.8 ;
      RECT  174.7 175.6 182.3 176.4 ;
      RECT  177.3 172.6 178.9 173.4 ;
      RECT  179.7 171.6 180.5 174.0 ;
      RECT  181.5 169.2 182.3 173.4 ;
      RECT  174.7 167.8 182.3 168.6 ;
      RECT  178.5 168.6 179.3 168.8 ;
      RECT  177.3 173.4 178.1 174.0 ;
      RECT  179.5 174.0 180.5 174.8 ;
      RECT  177.1 169.6 178.1 170.4 ;
      RECT  181.5 174.0 182.3 175.6 ;
      RECT  174.7 174.0 175.5 175.6 ;
      RECT  179.3 170.8 180.5 171.6 ;
      RECT  179.7 170.4 180.5 170.8 ;
      RECT  179.7 169.6 180.7 170.4 ;
      RECT  177.1 166.4 177.9 167.2 ;
      RECT  179.9 166.4 180.7 167.2 ;
      RECT  177.3 174.0 178.3 174.8 ;
      RECT  174.7 169.2 175.5 173.4 ;
      RECT  177.3 170.4 178.1 172.6 ;
      RECT  174.7 176.4 182.3 175.6 ;
      RECT  177.3 179.4 178.9 178.6 ;
      RECT  179.7 180.4 180.5 178.0 ;
      RECT  181.5 182.8 182.3 178.6 ;
      RECT  174.7 184.2 182.3 183.4 ;
      RECT  178.5 183.4 179.3 183.2 ;
      RECT  177.3 178.6 178.1 178.0 ;
      RECT  179.5 178.0 180.5 177.2 ;
      RECT  177.1 182.4 178.1 181.6 ;
      RECT  181.5 178.0 182.3 176.4 ;
      RECT  174.7 178.0 175.5 176.4 ;
      RECT  179.3 181.2 180.5 180.4 ;
      RECT  179.7 181.6 180.5 181.2 ;
      RECT  179.7 182.4 180.7 181.6 ;
      RECT  177.1 185.6 177.9 184.8 ;
      RECT  179.9 185.6 180.7 184.8 ;
      RECT  177.3 178.0 178.3 177.2 ;
      RECT  174.7 182.8 175.5 178.6 ;
      RECT  177.3 181.6 178.1 179.4 ;
      RECT  174.7 196.4 182.3 197.2 ;
      RECT  177.3 193.4 178.9 194.2 ;
      RECT  179.7 192.4 180.5 194.8 ;
      RECT  181.5 190.0 182.3 194.2 ;
      RECT  174.7 188.6 182.3 189.4 ;
      RECT  178.5 189.4 179.3 189.6 ;
      RECT  177.3 194.2 178.1 194.8 ;
      RECT  179.5 194.8 180.5 195.6 ;
      RECT  177.1 190.4 178.1 191.2 ;
      RECT  181.5 194.8 182.3 196.4 ;
      RECT  174.7 194.8 175.5 196.4 ;
      RECT  179.3 191.6 180.5 192.4 ;
      RECT  179.7 191.2 180.5 191.6 ;
      RECT  179.7 190.4 180.7 191.2 ;
      RECT  177.1 187.2 177.9 188.0 ;
      RECT  179.9 187.2 180.7 188.0 ;
      RECT  177.3 194.8 178.3 195.6 ;
      RECT  174.7 190.0 175.5 194.2 ;
      RECT  177.3 191.2 178.1 193.4 ;
      RECT  174.7 197.2 182.3 196.4 ;
      RECT  177.3 200.2 178.9 199.4 ;
      RECT  179.7 201.2 180.5 198.8 ;
      RECT  181.5 203.6 182.3 199.4 ;
      RECT  174.7 205.0 182.3 204.2 ;
      RECT  178.5 204.2 179.3 204.0 ;
      RECT  177.3 199.4 178.1 198.8 ;
      RECT  179.5 198.8 180.5 198.0 ;
      RECT  177.1 203.2 178.1 202.4 ;
      RECT  181.5 198.8 182.3 197.2 ;
      RECT  174.7 198.8 175.5 197.2 ;
      RECT  179.3 202.0 180.5 201.2 ;
      RECT  179.7 202.4 180.5 202.0 ;
      RECT  179.7 203.2 180.7 202.4 ;
      RECT  177.1 206.4 177.9 205.6 ;
      RECT  179.9 206.4 180.7 205.6 ;
      RECT  177.3 198.8 178.3 198.0 ;
      RECT  174.7 203.6 175.5 199.4 ;
      RECT  177.3 202.4 178.1 200.2 ;
      RECT  174.7 217.2 182.3 218.0 ;
      RECT  177.3 214.2 178.9 215.0 ;
      RECT  179.7 213.2 180.5 215.6 ;
      RECT  181.5 210.8 182.3 215.0 ;
      RECT  174.7 209.4 182.3 210.2 ;
      RECT  178.5 210.2 179.3 210.4 ;
      RECT  177.3 215.0 178.1 215.6 ;
      RECT  179.5 215.6 180.5 216.4 ;
      RECT  177.1 211.2 178.1 212.0 ;
      RECT  181.5 215.6 182.3 217.2 ;
      RECT  174.7 215.6 175.5 217.2 ;
      RECT  179.3 212.4 180.5 213.2 ;
      RECT  179.7 212.0 180.5 212.4 ;
      RECT  179.7 211.2 180.7 212.0 ;
      RECT  177.1 208.0 177.9 208.8 ;
      RECT  179.9 208.0 180.7 208.8 ;
      RECT  177.3 215.6 178.3 216.4 ;
      RECT  174.7 210.8 175.5 215.0 ;
      RECT  177.3 212.0 178.1 214.2 ;
      RECT  174.7 218.0 182.3 217.2 ;
      RECT  177.3 221.0 178.9 220.2 ;
      RECT  179.7 222.0 180.5 219.6 ;
      RECT  181.5 224.4 182.3 220.2 ;
      RECT  174.7 225.8 182.3 225.0 ;
      RECT  178.5 225.0 179.3 224.8 ;
      RECT  177.3 220.2 178.1 219.6 ;
      RECT  179.5 219.6 180.5 218.8 ;
      RECT  177.1 224.0 178.1 223.2 ;
      RECT  181.5 219.6 182.3 218.0 ;
      RECT  174.7 219.6 175.5 218.0 ;
      RECT  179.3 222.8 180.5 222.0 ;
      RECT  179.7 223.2 180.5 222.8 ;
      RECT  179.7 224.0 180.7 223.2 ;
      RECT  177.1 227.2 177.9 226.4 ;
      RECT  179.9 227.2 180.7 226.4 ;
      RECT  177.3 219.6 178.3 218.8 ;
      RECT  174.7 224.4 175.5 220.2 ;
      RECT  177.3 223.2 178.1 221.0 ;
      RECT  174.7 238.0 182.3 238.8 ;
      RECT  177.3 235.0 178.9 235.8 ;
      RECT  179.7 234.0 180.5 236.4 ;
      RECT  181.5 231.6 182.3 235.8 ;
      RECT  174.7 230.2 182.3 231.0 ;
      RECT  178.5 231.0 179.3 231.2 ;
      RECT  177.3 235.8 178.1 236.4 ;
      RECT  179.5 236.4 180.5 237.2 ;
      RECT  177.1 232.0 178.1 232.8 ;
      RECT  181.5 236.4 182.3 238.0 ;
      RECT  174.7 236.4 175.5 238.0 ;
      RECT  179.3 233.2 180.5 234.0 ;
      RECT  179.7 232.8 180.5 233.2 ;
      RECT  179.7 232.0 180.7 232.8 ;
      RECT  177.1 228.8 177.9 229.6 ;
      RECT  179.9 228.8 180.7 229.6 ;
      RECT  177.3 236.4 178.3 237.2 ;
      RECT  174.7 231.6 175.5 235.8 ;
      RECT  177.3 232.8 178.1 235.0 ;
      RECT  174.7 238.8 182.3 238.0 ;
      RECT  177.3 241.8 178.9 241.0 ;
      RECT  179.7 242.8 180.5 240.4 ;
      RECT  181.5 245.2 182.3 241.0 ;
      RECT  174.7 246.6 182.3 245.8 ;
      RECT  178.5 245.8 179.3 245.6 ;
      RECT  177.3 241.0 178.1 240.4 ;
      RECT  179.5 240.4 180.5 239.6 ;
      RECT  177.1 244.8 178.1 244.0 ;
      RECT  181.5 240.4 182.3 238.8 ;
      RECT  174.7 240.4 175.5 238.8 ;
      RECT  179.3 243.6 180.5 242.8 ;
      RECT  179.7 244.0 180.5 243.6 ;
      RECT  179.7 244.8 180.7 244.0 ;
      RECT  177.1 248.0 177.9 247.2 ;
      RECT  179.9 248.0 180.7 247.2 ;
      RECT  177.3 240.4 178.3 239.6 ;
      RECT  174.7 245.2 175.5 241.0 ;
      RECT  177.3 244.0 178.1 241.8 ;
      RECT  174.7 258.8 182.3 259.6 ;
      RECT  177.3 255.8 178.9 256.6 ;
      RECT  179.7 254.8 180.5 257.2 ;
      RECT  181.5 252.4 182.3 256.6 ;
      RECT  174.7 251.0 182.3 251.8 ;
      RECT  178.5 251.8 179.3 252.0 ;
      RECT  177.3 256.6 178.1 257.2 ;
      RECT  179.5 257.2 180.5 258.0 ;
      RECT  177.1 252.8 178.1 253.6 ;
      RECT  181.5 257.2 182.3 258.8 ;
      RECT  174.7 257.2 175.5 258.8 ;
      RECT  179.3 254.0 180.5 254.8 ;
      RECT  179.7 253.6 180.5 254.0 ;
      RECT  179.7 252.8 180.7 253.6 ;
      RECT  177.1 249.6 177.9 250.4 ;
      RECT  179.9 249.6 180.7 250.4 ;
      RECT  177.3 257.2 178.3 258.0 ;
      RECT  174.7 252.4 175.5 256.6 ;
      RECT  177.3 253.6 178.1 255.8 ;
      RECT  174.7 259.6 182.3 258.8 ;
      RECT  177.3 262.6 178.9 261.8 ;
      RECT  179.7 263.6 180.5 261.2 ;
      RECT  181.5 266.0 182.3 261.8 ;
      RECT  174.7 267.4 182.3 266.6 ;
      RECT  178.5 266.6 179.3 266.4 ;
      RECT  177.3 261.8 178.1 261.2 ;
      RECT  179.5 261.2 180.5 260.4 ;
      RECT  177.1 265.6 178.1 264.8 ;
      RECT  181.5 261.2 182.3 259.6 ;
      RECT  174.7 261.2 175.5 259.6 ;
      RECT  179.3 264.4 180.5 263.6 ;
      RECT  179.7 264.8 180.5 264.4 ;
      RECT  179.7 265.6 180.7 264.8 ;
      RECT  177.1 268.8 177.9 268.0 ;
      RECT  179.9 268.8 180.7 268.0 ;
      RECT  177.3 261.2 178.3 260.4 ;
      RECT  174.7 266.0 175.5 261.8 ;
      RECT  177.3 264.8 178.1 262.6 ;
      RECT  174.7 279.6 182.3 280.4 ;
      RECT  177.3 276.6 178.9 277.4 ;
      RECT  179.7 275.6 180.5 278.0 ;
      RECT  181.5 273.2 182.3 277.4 ;
      RECT  174.7 271.8 182.3 272.6 ;
      RECT  178.5 272.6 179.3 272.8 ;
      RECT  177.3 277.4 178.1 278.0 ;
      RECT  179.5 278.0 180.5 278.8 ;
      RECT  177.1 273.6 178.1 274.4 ;
      RECT  181.5 278.0 182.3 279.6 ;
      RECT  174.7 278.0 175.5 279.6 ;
      RECT  179.3 274.8 180.5 275.6 ;
      RECT  179.7 274.4 180.5 274.8 ;
      RECT  179.7 273.6 180.7 274.4 ;
      RECT  177.1 270.4 177.9 271.2 ;
      RECT  179.9 270.4 180.7 271.2 ;
      RECT  177.3 278.0 178.3 278.8 ;
      RECT  174.7 273.2 175.5 277.4 ;
      RECT  177.3 274.4 178.1 276.6 ;
      RECT  174.7 280.4 182.3 279.6 ;
      RECT  177.3 283.4 178.9 282.6 ;
      RECT  179.7 284.4 180.5 282.0 ;
      RECT  181.5 286.8 182.3 282.6 ;
      RECT  174.7 288.2 182.3 287.4 ;
      RECT  178.5 287.4 179.3 287.2 ;
      RECT  177.3 282.6 178.1 282.0 ;
      RECT  179.5 282.0 180.5 281.2 ;
      RECT  177.1 286.4 178.1 285.6 ;
      RECT  181.5 282.0 182.3 280.4 ;
      RECT  174.7 282.0 175.5 280.4 ;
      RECT  179.3 285.2 180.5 284.4 ;
      RECT  179.7 285.6 180.5 285.2 ;
      RECT  179.7 286.4 180.7 285.6 ;
      RECT  177.1 289.6 177.9 288.8 ;
      RECT  179.9 289.6 180.7 288.8 ;
      RECT  177.3 282.0 178.3 281.2 ;
      RECT  174.7 286.8 175.5 282.6 ;
      RECT  177.3 285.6 178.1 283.4 ;
      RECT  174.7 300.4 182.3 301.2 ;
      RECT  177.3 297.4 178.9 298.2 ;
      RECT  179.7 296.4 180.5 298.8 ;
      RECT  181.5 294.0 182.3 298.2 ;
      RECT  174.7 292.6 182.3 293.4 ;
      RECT  178.5 293.4 179.3 293.6 ;
      RECT  177.3 298.2 178.1 298.8 ;
      RECT  179.5 298.8 180.5 299.6 ;
      RECT  177.1 294.4 178.1 295.2 ;
      RECT  181.5 298.8 182.3 300.4 ;
      RECT  174.7 298.8 175.5 300.4 ;
      RECT  179.3 295.6 180.5 296.4 ;
      RECT  179.7 295.2 180.5 295.6 ;
      RECT  179.7 294.4 180.7 295.2 ;
      RECT  177.1 291.2 177.9 292.0 ;
      RECT  179.9 291.2 180.7 292.0 ;
      RECT  177.3 298.8 178.3 299.6 ;
      RECT  174.7 294.0 175.5 298.2 ;
      RECT  177.3 295.2 178.1 297.4 ;
      RECT  174.7 301.2 182.3 300.4 ;
      RECT  177.3 304.2 178.9 303.4 ;
      RECT  179.7 305.2 180.5 302.8 ;
      RECT  181.5 307.6 182.3 303.4 ;
      RECT  174.7 309.0 182.3 308.2 ;
      RECT  178.5 308.2 179.3 308.0 ;
      RECT  177.3 303.4 178.1 302.8 ;
      RECT  179.5 302.8 180.5 302.0 ;
      RECT  177.1 307.2 178.1 306.4 ;
      RECT  181.5 302.8 182.3 301.2 ;
      RECT  174.7 302.8 175.5 301.2 ;
      RECT  179.3 306.0 180.5 305.2 ;
      RECT  179.7 306.4 180.5 306.0 ;
      RECT  179.7 307.2 180.7 306.4 ;
      RECT  177.1 310.4 177.9 309.6 ;
      RECT  179.9 310.4 180.7 309.6 ;
      RECT  177.3 302.8 178.3 302.0 ;
      RECT  174.7 307.6 175.5 303.4 ;
      RECT  177.3 306.4 178.1 304.2 ;
      RECT  174.7 321.2 182.3 322.0 ;
      RECT  177.3 318.2 178.9 319.0 ;
      RECT  179.7 317.2 180.5 319.6 ;
      RECT  181.5 314.8 182.3 319.0 ;
      RECT  174.7 313.4 182.3 314.2 ;
      RECT  178.5 314.2 179.3 314.4 ;
      RECT  177.3 319.0 178.1 319.6 ;
      RECT  179.5 319.6 180.5 320.4 ;
      RECT  177.1 315.2 178.1 316.0 ;
      RECT  181.5 319.6 182.3 321.2 ;
      RECT  174.7 319.6 175.5 321.2 ;
      RECT  179.3 316.4 180.5 317.2 ;
      RECT  179.7 316.0 180.5 316.4 ;
      RECT  179.7 315.2 180.7 316.0 ;
      RECT  177.1 312.0 177.9 312.8 ;
      RECT  179.9 312.0 180.7 312.8 ;
      RECT  177.3 319.6 178.3 320.4 ;
      RECT  174.7 314.8 175.5 319.0 ;
      RECT  177.3 316.0 178.1 318.2 ;
      RECT  174.7 322.0 182.3 321.2 ;
      RECT  177.3 325.0 178.9 324.2 ;
      RECT  179.7 326.0 180.5 323.6 ;
      RECT  181.5 328.4 182.3 324.2 ;
      RECT  174.7 329.8 182.3 329.0 ;
      RECT  178.5 329.0 179.3 328.8 ;
      RECT  177.3 324.2 178.1 323.6 ;
      RECT  179.5 323.6 180.5 322.8 ;
      RECT  177.1 328.0 178.1 327.2 ;
      RECT  181.5 323.6 182.3 322.0 ;
      RECT  174.7 323.6 175.5 322.0 ;
      RECT  179.3 326.8 180.5 326.0 ;
      RECT  179.7 327.2 180.5 326.8 ;
      RECT  179.7 328.0 180.7 327.2 ;
      RECT  177.1 331.2 177.9 330.4 ;
      RECT  179.9 331.2 180.7 330.4 ;
      RECT  177.3 323.6 178.3 322.8 ;
      RECT  174.7 328.4 175.5 324.2 ;
      RECT  177.3 327.2 178.1 325.0 ;
      RECT  174.7 342.0 182.3 342.8 ;
      RECT  177.3 339.0 178.9 339.8 ;
      RECT  179.7 338.0 180.5 340.4 ;
      RECT  181.5 335.6 182.3 339.8 ;
      RECT  174.7 334.2 182.3 335.0 ;
      RECT  178.5 335.0 179.3 335.2 ;
      RECT  177.3 339.8 178.1 340.4 ;
      RECT  179.5 340.4 180.5 341.2 ;
      RECT  177.1 336.0 178.1 336.8 ;
      RECT  181.5 340.4 182.3 342.0 ;
      RECT  174.7 340.4 175.5 342.0 ;
      RECT  179.3 337.2 180.5 338.0 ;
      RECT  179.7 336.8 180.5 337.2 ;
      RECT  179.7 336.0 180.7 336.8 ;
      RECT  177.1 332.8 177.9 333.6 ;
      RECT  179.9 332.8 180.7 333.6 ;
      RECT  177.3 340.4 178.3 341.2 ;
      RECT  174.7 335.6 175.5 339.8 ;
      RECT  177.3 336.8 178.1 339.0 ;
      RECT  174.7 342.8 182.3 342.0 ;
      RECT  177.3 345.8 178.9 345.0 ;
      RECT  179.7 346.8 180.5 344.4 ;
      RECT  181.5 349.2 182.3 345.0 ;
      RECT  174.7 350.6 182.3 349.8 ;
      RECT  178.5 349.8 179.3 349.6 ;
      RECT  177.3 345.0 178.1 344.4 ;
      RECT  179.5 344.4 180.5 343.6 ;
      RECT  177.1 348.8 178.1 348.0 ;
      RECT  181.5 344.4 182.3 342.8 ;
      RECT  174.7 344.4 175.5 342.8 ;
      RECT  179.3 347.6 180.5 346.8 ;
      RECT  179.7 348.0 180.5 347.6 ;
      RECT  179.7 348.8 180.7 348.0 ;
      RECT  177.1 352.0 177.9 351.2 ;
      RECT  179.9 352.0 180.7 351.2 ;
      RECT  177.3 344.4 178.3 343.6 ;
      RECT  174.7 349.2 175.5 345.0 ;
      RECT  177.3 348.0 178.1 345.8 ;
      RECT  174.7 362.8 182.3 363.6 ;
      RECT  177.3 359.8 178.9 360.6 ;
      RECT  179.7 358.8 180.5 361.2 ;
      RECT  181.5 356.4 182.3 360.6 ;
      RECT  174.7 355.0 182.3 355.8 ;
      RECT  178.5 355.8 179.3 356.0 ;
      RECT  177.3 360.6 178.1 361.2 ;
      RECT  179.5 361.2 180.5 362.0 ;
      RECT  177.1 356.8 178.1 357.6 ;
      RECT  181.5 361.2 182.3 362.8 ;
      RECT  174.7 361.2 175.5 362.8 ;
      RECT  179.3 358.0 180.5 358.8 ;
      RECT  179.7 357.6 180.5 358.0 ;
      RECT  179.7 356.8 180.7 357.6 ;
      RECT  177.1 353.6 177.9 354.4 ;
      RECT  179.9 353.6 180.7 354.4 ;
      RECT  177.3 361.2 178.3 362.0 ;
      RECT  174.7 356.4 175.5 360.6 ;
      RECT  177.3 357.6 178.1 359.8 ;
      RECT  175.1 167.8 181.9 168.6 ;
      RECT  175.1 183.4 181.9 184.2 ;
      RECT  175.1 188.6 181.9 189.4 ;
      RECT  175.1 204.2 181.9 205.0 ;
      RECT  175.1 209.4 181.9 210.2 ;
      RECT  175.1 225.0 181.9 225.8 ;
      RECT  175.1 230.2 181.9 231.0 ;
      RECT  175.1 245.8 181.9 246.6 ;
      RECT  175.1 251.0 181.9 251.8 ;
      RECT  175.1 266.6 181.9 267.4 ;
      RECT  175.1 271.8 181.9 272.6 ;
      RECT  175.1 287.4 181.9 288.2 ;
      RECT  175.1 292.6 181.9 293.4 ;
      RECT  175.1 308.2 181.9 309.0 ;
      RECT  175.1 313.4 181.9 314.2 ;
      RECT  175.1 329.0 181.9 329.8 ;
      RECT  175.1 334.2 181.9 335.0 ;
      RECT  175.1 349.8 181.9 350.6 ;
      RECT  175.1 355.0 181.9 355.8 ;
      RECT  201.9 175.6 209.5 176.4 ;
      RECT  204.5 172.6 206.1 173.4 ;
      RECT  206.9 171.6 207.7 174.0 ;
      RECT  208.7 169.2 209.5 173.4 ;
      RECT  201.9 167.8 209.5 168.6 ;
      RECT  205.7 168.6 206.5 168.8 ;
      RECT  204.5 173.4 205.3 174.0 ;
      RECT  206.7 174.0 207.7 174.8 ;
      RECT  204.3 169.6 205.3 170.4 ;
      RECT  208.7 174.0 209.5 175.6 ;
      RECT  201.9 174.0 202.7 175.6 ;
      RECT  206.5 170.8 207.7 171.6 ;
      RECT  206.9 170.4 207.7 170.8 ;
      RECT  206.9 169.6 207.9 170.4 ;
      RECT  204.3 166.4 205.1 167.2 ;
      RECT  207.1 166.4 207.9 167.2 ;
      RECT  204.5 174.0 205.5 174.8 ;
      RECT  201.9 169.2 202.7 173.4 ;
      RECT  204.5 170.4 205.3 172.6 ;
      RECT  201.9 176.4 209.5 175.6 ;
      RECT  204.5 179.4 206.1 178.6 ;
      RECT  206.9 180.4 207.7 178.0 ;
      RECT  208.7 182.8 209.5 178.6 ;
      RECT  201.9 184.2 209.5 183.4 ;
      RECT  205.7 183.4 206.5 183.2 ;
      RECT  204.5 178.6 205.3 178.0 ;
      RECT  206.7 178.0 207.7 177.2 ;
      RECT  204.3 182.4 205.3 181.6 ;
      RECT  208.7 178.0 209.5 176.4 ;
      RECT  201.9 178.0 202.7 176.4 ;
      RECT  206.5 181.2 207.7 180.4 ;
      RECT  206.9 181.6 207.7 181.2 ;
      RECT  206.9 182.4 207.9 181.6 ;
      RECT  204.3 185.6 205.1 184.8 ;
      RECT  207.1 185.6 207.9 184.8 ;
      RECT  204.5 178.0 205.5 177.2 ;
      RECT  201.9 182.8 202.7 178.6 ;
      RECT  204.5 181.6 205.3 179.4 ;
      RECT  201.9 196.4 209.5 197.2 ;
      RECT  204.5 193.4 206.1 194.2 ;
      RECT  206.9 192.4 207.7 194.8 ;
      RECT  208.7 190.0 209.5 194.2 ;
      RECT  201.9 188.6 209.5 189.4 ;
      RECT  205.7 189.4 206.5 189.6 ;
      RECT  204.5 194.2 205.3 194.8 ;
      RECT  206.7 194.8 207.7 195.6 ;
      RECT  204.3 190.4 205.3 191.2 ;
      RECT  208.7 194.8 209.5 196.4 ;
      RECT  201.9 194.8 202.7 196.4 ;
      RECT  206.5 191.6 207.7 192.4 ;
      RECT  206.9 191.2 207.7 191.6 ;
      RECT  206.9 190.4 207.9 191.2 ;
      RECT  204.3 187.2 205.1 188.0 ;
      RECT  207.1 187.2 207.9 188.0 ;
      RECT  204.5 194.8 205.5 195.6 ;
      RECT  201.9 190.0 202.7 194.2 ;
      RECT  204.5 191.2 205.3 193.4 ;
      RECT  201.9 197.2 209.5 196.4 ;
      RECT  204.5 200.2 206.1 199.4 ;
      RECT  206.9 201.2 207.7 198.8 ;
      RECT  208.7 203.6 209.5 199.4 ;
      RECT  201.9 205.0 209.5 204.2 ;
      RECT  205.7 204.2 206.5 204.0 ;
      RECT  204.5 199.4 205.3 198.8 ;
      RECT  206.7 198.8 207.7 198.0 ;
      RECT  204.3 203.2 205.3 202.4 ;
      RECT  208.7 198.8 209.5 197.2 ;
      RECT  201.9 198.8 202.7 197.2 ;
      RECT  206.5 202.0 207.7 201.2 ;
      RECT  206.9 202.4 207.7 202.0 ;
      RECT  206.9 203.2 207.9 202.4 ;
      RECT  204.3 206.4 205.1 205.6 ;
      RECT  207.1 206.4 207.9 205.6 ;
      RECT  204.5 198.8 205.5 198.0 ;
      RECT  201.9 203.6 202.7 199.4 ;
      RECT  204.5 202.4 205.3 200.2 ;
      RECT  201.9 217.2 209.5 218.0 ;
      RECT  204.5 214.2 206.1 215.0 ;
      RECT  206.9 213.2 207.7 215.6 ;
      RECT  208.7 210.8 209.5 215.0 ;
      RECT  201.9 209.4 209.5 210.2 ;
      RECT  205.7 210.2 206.5 210.4 ;
      RECT  204.5 215.0 205.3 215.6 ;
      RECT  206.7 215.6 207.7 216.4 ;
      RECT  204.3 211.2 205.3 212.0 ;
      RECT  208.7 215.6 209.5 217.2 ;
      RECT  201.9 215.6 202.7 217.2 ;
      RECT  206.5 212.4 207.7 213.2 ;
      RECT  206.9 212.0 207.7 212.4 ;
      RECT  206.9 211.2 207.9 212.0 ;
      RECT  204.3 208.0 205.1 208.8 ;
      RECT  207.1 208.0 207.9 208.8 ;
      RECT  204.5 215.6 205.5 216.4 ;
      RECT  201.9 210.8 202.7 215.0 ;
      RECT  204.5 212.0 205.3 214.2 ;
      RECT  201.9 218.0 209.5 217.2 ;
      RECT  204.5 221.0 206.1 220.2 ;
      RECT  206.9 222.0 207.7 219.6 ;
      RECT  208.7 224.4 209.5 220.2 ;
      RECT  201.9 225.8 209.5 225.0 ;
      RECT  205.7 225.0 206.5 224.8 ;
      RECT  204.5 220.2 205.3 219.6 ;
      RECT  206.7 219.6 207.7 218.8 ;
      RECT  204.3 224.0 205.3 223.2 ;
      RECT  208.7 219.6 209.5 218.0 ;
      RECT  201.9 219.6 202.7 218.0 ;
      RECT  206.5 222.8 207.7 222.0 ;
      RECT  206.9 223.2 207.7 222.8 ;
      RECT  206.9 224.0 207.9 223.2 ;
      RECT  204.3 227.2 205.1 226.4 ;
      RECT  207.1 227.2 207.9 226.4 ;
      RECT  204.5 219.6 205.5 218.8 ;
      RECT  201.9 224.4 202.7 220.2 ;
      RECT  204.5 223.2 205.3 221.0 ;
      RECT  201.9 238.0 209.5 238.8 ;
      RECT  204.5 235.0 206.1 235.8 ;
      RECT  206.9 234.0 207.7 236.4 ;
      RECT  208.7 231.6 209.5 235.8 ;
      RECT  201.9 230.2 209.5 231.0 ;
      RECT  205.7 231.0 206.5 231.2 ;
      RECT  204.5 235.8 205.3 236.4 ;
      RECT  206.7 236.4 207.7 237.2 ;
      RECT  204.3 232.0 205.3 232.8 ;
      RECT  208.7 236.4 209.5 238.0 ;
      RECT  201.9 236.4 202.7 238.0 ;
      RECT  206.5 233.2 207.7 234.0 ;
      RECT  206.9 232.8 207.7 233.2 ;
      RECT  206.9 232.0 207.9 232.8 ;
      RECT  204.3 228.8 205.1 229.6 ;
      RECT  207.1 228.8 207.9 229.6 ;
      RECT  204.5 236.4 205.5 237.2 ;
      RECT  201.9 231.6 202.7 235.8 ;
      RECT  204.5 232.8 205.3 235.0 ;
      RECT  201.9 238.8 209.5 238.0 ;
      RECT  204.5 241.8 206.1 241.0 ;
      RECT  206.9 242.8 207.7 240.4 ;
      RECT  208.7 245.2 209.5 241.0 ;
      RECT  201.9 246.6 209.5 245.8 ;
      RECT  205.7 245.8 206.5 245.6 ;
      RECT  204.5 241.0 205.3 240.4 ;
      RECT  206.7 240.4 207.7 239.6 ;
      RECT  204.3 244.8 205.3 244.0 ;
      RECT  208.7 240.4 209.5 238.8 ;
      RECT  201.9 240.4 202.7 238.8 ;
      RECT  206.5 243.6 207.7 242.8 ;
      RECT  206.9 244.0 207.7 243.6 ;
      RECT  206.9 244.8 207.9 244.0 ;
      RECT  204.3 248.0 205.1 247.2 ;
      RECT  207.1 248.0 207.9 247.2 ;
      RECT  204.5 240.4 205.5 239.6 ;
      RECT  201.9 245.2 202.7 241.0 ;
      RECT  204.5 244.0 205.3 241.8 ;
      RECT  201.9 258.8 209.5 259.6 ;
      RECT  204.5 255.8 206.1 256.6 ;
      RECT  206.9 254.8 207.7 257.2 ;
      RECT  208.7 252.4 209.5 256.6 ;
      RECT  201.9 251.0 209.5 251.8 ;
      RECT  205.7 251.8 206.5 252.0 ;
      RECT  204.5 256.6 205.3 257.2 ;
      RECT  206.7 257.2 207.7 258.0 ;
      RECT  204.3 252.8 205.3 253.6 ;
      RECT  208.7 257.2 209.5 258.8 ;
      RECT  201.9 257.2 202.7 258.8 ;
      RECT  206.5 254.0 207.7 254.8 ;
      RECT  206.9 253.6 207.7 254.0 ;
      RECT  206.9 252.8 207.9 253.6 ;
      RECT  204.3 249.6 205.1 250.4 ;
      RECT  207.1 249.6 207.9 250.4 ;
      RECT  204.5 257.2 205.5 258.0 ;
      RECT  201.9 252.4 202.7 256.6 ;
      RECT  204.5 253.6 205.3 255.8 ;
      RECT  201.9 259.6 209.5 258.8 ;
      RECT  204.5 262.6 206.1 261.8 ;
      RECT  206.9 263.6 207.7 261.2 ;
      RECT  208.7 266.0 209.5 261.8 ;
      RECT  201.9 267.4 209.5 266.6 ;
      RECT  205.7 266.6 206.5 266.4 ;
      RECT  204.5 261.8 205.3 261.2 ;
      RECT  206.7 261.2 207.7 260.4 ;
      RECT  204.3 265.6 205.3 264.8 ;
      RECT  208.7 261.2 209.5 259.6 ;
      RECT  201.9 261.2 202.7 259.6 ;
      RECT  206.5 264.4 207.7 263.6 ;
      RECT  206.9 264.8 207.7 264.4 ;
      RECT  206.9 265.6 207.9 264.8 ;
      RECT  204.3 268.8 205.1 268.0 ;
      RECT  207.1 268.8 207.9 268.0 ;
      RECT  204.5 261.2 205.5 260.4 ;
      RECT  201.9 266.0 202.7 261.8 ;
      RECT  204.5 264.8 205.3 262.6 ;
      RECT  201.9 279.6 209.5 280.4 ;
      RECT  204.5 276.6 206.1 277.4 ;
      RECT  206.9 275.6 207.7 278.0 ;
      RECT  208.7 273.2 209.5 277.4 ;
      RECT  201.9 271.8 209.5 272.6 ;
      RECT  205.7 272.6 206.5 272.8 ;
      RECT  204.5 277.4 205.3 278.0 ;
      RECT  206.7 278.0 207.7 278.8 ;
      RECT  204.3 273.6 205.3 274.4 ;
      RECT  208.7 278.0 209.5 279.6 ;
      RECT  201.9 278.0 202.7 279.6 ;
      RECT  206.5 274.8 207.7 275.6 ;
      RECT  206.9 274.4 207.7 274.8 ;
      RECT  206.9 273.6 207.9 274.4 ;
      RECT  204.3 270.4 205.1 271.2 ;
      RECT  207.1 270.4 207.9 271.2 ;
      RECT  204.5 278.0 205.5 278.8 ;
      RECT  201.9 273.2 202.7 277.4 ;
      RECT  204.5 274.4 205.3 276.6 ;
      RECT  201.9 280.4 209.5 279.6 ;
      RECT  204.5 283.4 206.1 282.6 ;
      RECT  206.9 284.4 207.7 282.0 ;
      RECT  208.7 286.8 209.5 282.6 ;
      RECT  201.9 288.2 209.5 287.4 ;
      RECT  205.7 287.4 206.5 287.2 ;
      RECT  204.5 282.6 205.3 282.0 ;
      RECT  206.7 282.0 207.7 281.2 ;
      RECT  204.3 286.4 205.3 285.6 ;
      RECT  208.7 282.0 209.5 280.4 ;
      RECT  201.9 282.0 202.7 280.4 ;
      RECT  206.5 285.2 207.7 284.4 ;
      RECT  206.9 285.6 207.7 285.2 ;
      RECT  206.9 286.4 207.9 285.6 ;
      RECT  204.3 289.6 205.1 288.8 ;
      RECT  207.1 289.6 207.9 288.8 ;
      RECT  204.5 282.0 205.5 281.2 ;
      RECT  201.9 286.8 202.7 282.6 ;
      RECT  204.5 285.6 205.3 283.4 ;
      RECT  201.9 300.4 209.5 301.2 ;
      RECT  204.5 297.4 206.1 298.2 ;
      RECT  206.9 296.4 207.7 298.8 ;
      RECT  208.7 294.0 209.5 298.2 ;
      RECT  201.9 292.6 209.5 293.4 ;
      RECT  205.7 293.4 206.5 293.6 ;
      RECT  204.5 298.2 205.3 298.8 ;
      RECT  206.7 298.8 207.7 299.6 ;
      RECT  204.3 294.4 205.3 295.2 ;
      RECT  208.7 298.8 209.5 300.4 ;
      RECT  201.9 298.8 202.7 300.4 ;
      RECT  206.5 295.6 207.7 296.4 ;
      RECT  206.9 295.2 207.7 295.6 ;
      RECT  206.9 294.4 207.9 295.2 ;
      RECT  204.3 291.2 205.1 292.0 ;
      RECT  207.1 291.2 207.9 292.0 ;
      RECT  204.5 298.8 205.5 299.6 ;
      RECT  201.9 294.0 202.7 298.2 ;
      RECT  204.5 295.2 205.3 297.4 ;
      RECT  201.9 301.2 209.5 300.4 ;
      RECT  204.5 304.2 206.1 303.4 ;
      RECT  206.9 305.2 207.7 302.8 ;
      RECT  208.7 307.6 209.5 303.4 ;
      RECT  201.9 309.0 209.5 308.2 ;
      RECT  205.7 308.2 206.5 308.0 ;
      RECT  204.5 303.4 205.3 302.8 ;
      RECT  206.7 302.8 207.7 302.0 ;
      RECT  204.3 307.2 205.3 306.4 ;
      RECT  208.7 302.8 209.5 301.2 ;
      RECT  201.9 302.8 202.7 301.2 ;
      RECT  206.5 306.0 207.7 305.2 ;
      RECT  206.9 306.4 207.7 306.0 ;
      RECT  206.9 307.2 207.9 306.4 ;
      RECT  204.3 310.4 205.1 309.6 ;
      RECT  207.1 310.4 207.9 309.6 ;
      RECT  204.5 302.8 205.5 302.0 ;
      RECT  201.9 307.6 202.7 303.4 ;
      RECT  204.5 306.4 205.3 304.2 ;
      RECT  201.9 321.2 209.5 322.0 ;
      RECT  204.5 318.2 206.1 319.0 ;
      RECT  206.9 317.2 207.7 319.6 ;
      RECT  208.7 314.8 209.5 319.0 ;
      RECT  201.9 313.4 209.5 314.2 ;
      RECT  205.7 314.2 206.5 314.4 ;
      RECT  204.5 319.0 205.3 319.6 ;
      RECT  206.7 319.6 207.7 320.4 ;
      RECT  204.3 315.2 205.3 316.0 ;
      RECT  208.7 319.6 209.5 321.2 ;
      RECT  201.9 319.6 202.7 321.2 ;
      RECT  206.5 316.4 207.7 317.2 ;
      RECT  206.9 316.0 207.7 316.4 ;
      RECT  206.9 315.2 207.9 316.0 ;
      RECT  204.3 312.0 205.1 312.8 ;
      RECT  207.1 312.0 207.9 312.8 ;
      RECT  204.5 319.6 205.5 320.4 ;
      RECT  201.9 314.8 202.7 319.0 ;
      RECT  204.5 316.0 205.3 318.2 ;
      RECT  201.9 322.0 209.5 321.2 ;
      RECT  204.5 325.0 206.1 324.2 ;
      RECT  206.9 326.0 207.7 323.6 ;
      RECT  208.7 328.4 209.5 324.2 ;
      RECT  201.9 329.8 209.5 329.0 ;
      RECT  205.7 329.0 206.5 328.8 ;
      RECT  204.5 324.2 205.3 323.6 ;
      RECT  206.7 323.6 207.7 322.8 ;
      RECT  204.3 328.0 205.3 327.2 ;
      RECT  208.7 323.6 209.5 322.0 ;
      RECT  201.9 323.6 202.7 322.0 ;
      RECT  206.5 326.8 207.7 326.0 ;
      RECT  206.9 327.2 207.7 326.8 ;
      RECT  206.9 328.0 207.9 327.2 ;
      RECT  204.3 331.2 205.1 330.4 ;
      RECT  207.1 331.2 207.9 330.4 ;
      RECT  204.5 323.6 205.5 322.8 ;
      RECT  201.9 328.4 202.7 324.2 ;
      RECT  204.5 327.2 205.3 325.0 ;
      RECT  201.9 342.0 209.5 342.8 ;
      RECT  204.5 339.0 206.1 339.8 ;
      RECT  206.9 338.0 207.7 340.4 ;
      RECT  208.7 335.6 209.5 339.8 ;
      RECT  201.9 334.2 209.5 335.0 ;
      RECT  205.7 335.0 206.5 335.2 ;
      RECT  204.5 339.8 205.3 340.4 ;
      RECT  206.7 340.4 207.7 341.2 ;
      RECT  204.3 336.0 205.3 336.8 ;
      RECT  208.7 340.4 209.5 342.0 ;
      RECT  201.9 340.4 202.7 342.0 ;
      RECT  206.5 337.2 207.7 338.0 ;
      RECT  206.9 336.8 207.7 337.2 ;
      RECT  206.9 336.0 207.9 336.8 ;
      RECT  204.3 332.8 205.1 333.6 ;
      RECT  207.1 332.8 207.9 333.6 ;
      RECT  204.5 340.4 205.5 341.2 ;
      RECT  201.9 335.6 202.7 339.8 ;
      RECT  204.5 336.8 205.3 339.0 ;
      RECT  201.9 342.8 209.5 342.0 ;
      RECT  204.5 345.8 206.1 345.0 ;
      RECT  206.9 346.8 207.7 344.4 ;
      RECT  208.7 349.2 209.5 345.0 ;
      RECT  201.9 350.6 209.5 349.8 ;
      RECT  205.7 349.8 206.5 349.6 ;
      RECT  204.5 345.0 205.3 344.4 ;
      RECT  206.7 344.4 207.7 343.6 ;
      RECT  204.3 348.8 205.3 348.0 ;
      RECT  208.7 344.4 209.5 342.8 ;
      RECT  201.9 344.4 202.7 342.8 ;
      RECT  206.5 347.6 207.7 346.8 ;
      RECT  206.9 348.0 207.7 347.6 ;
      RECT  206.9 348.8 207.9 348.0 ;
      RECT  204.3 352.0 205.1 351.2 ;
      RECT  207.1 352.0 207.9 351.2 ;
      RECT  204.5 344.4 205.5 343.6 ;
      RECT  201.9 349.2 202.7 345.0 ;
      RECT  204.5 348.0 205.3 345.8 ;
      RECT  201.9 362.8 209.5 363.6 ;
      RECT  204.5 359.8 206.1 360.6 ;
      RECT  206.9 358.8 207.7 361.2 ;
      RECT  208.7 356.4 209.5 360.6 ;
      RECT  201.9 355.0 209.5 355.8 ;
      RECT  205.7 355.8 206.5 356.0 ;
      RECT  204.5 360.6 205.3 361.2 ;
      RECT  206.7 361.2 207.7 362.0 ;
      RECT  204.3 356.8 205.3 357.6 ;
      RECT  208.7 361.2 209.5 362.8 ;
      RECT  201.9 361.2 202.7 362.8 ;
      RECT  206.5 358.0 207.7 358.8 ;
      RECT  206.9 357.6 207.7 358.0 ;
      RECT  206.9 356.8 207.9 357.6 ;
      RECT  204.3 353.6 205.1 354.4 ;
      RECT  207.1 353.6 207.9 354.4 ;
      RECT  204.5 361.2 205.5 362.0 ;
      RECT  201.9 356.4 202.7 360.6 ;
      RECT  204.5 357.6 205.3 359.8 ;
      RECT  202.3 167.8 209.1 168.6 ;
      RECT  202.3 183.4 209.1 184.2 ;
      RECT  202.3 188.6 209.1 189.4 ;
      RECT  202.3 204.2 209.1 205.0 ;
      RECT  202.3 209.4 209.1 210.2 ;
      RECT  202.3 225.0 209.1 225.8 ;
      RECT  202.3 230.2 209.1 231.0 ;
      RECT  202.3 245.8 209.1 246.6 ;
      RECT  202.3 251.0 209.1 251.8 ;
      RECT  202.3 266.6 209.1 267.4 ;
      RECT  202.3 271.8 209.1 272.6 ;
      RECT  202.3 287.4 209.1 288.2 ;
      RECT  202.3 292.6 209.1 293.4 ;
      RECT  202.3 308.2 209.1 309.0 ;
      RECT  202.3 313.4 209.1 314.2 ;
      RECT  202.3 329.0 209.1 329.8 ;
      RECT  202.3 334.2 209.1 335.0 ;
      RECT  202.3 349.8 209.1 350.6 ;
      RECT  202.3 355.0 209.1 355.8 ;
      RECT  173.0 183.4 211.2 184.2 ;
      RECT  173.0 188.6 211.2 189.4 ;
      RECT  173.0 204.2 211.2 205.0 ;
      RECT  173.0 209.4 211.2 210.2 ;
      RECT  173.0 225.0 211.2 225.8 ;
      RECT  173.0 230.2 211.2 231.0 ;
      RECT  173.0 245.8 211.2 246.6 ;
      RECT  173.0 251.0 211.2 251.8 ;
      RECT  173.0 266.6 211.2 267.4 ;
      RECT  173.0 271.8 211.2 272.6 ;
      RECT  173.0 287.4 211.2 288.2 ;
      RECT  173.0 292.6 211.2 293.4 ;
      RECT  173.0 308.2 211.2 309.0 ;
      RECT  173.0 313.4 211.2 314.2 ;
      RECT  173.0 329.0 211.2 329.8 ;
      RECT  173.0 334.2 211.2 335.0 ;
      RECT  173.0 349.8 211.2 350.6 ;
      RECT  185.4 152.4 186.2 153.2 ;
      RECT  183.4 152.4 184.2 153.2 ;
      RECT  185.4 156.8 186.2 157.6 ;
      RECT  183.4 156.8 184.2 157.6 ;
      RECT  187.4 156.8 188.2 157.6 ;
      RECT  185.4 156.8 186.2 157.6 ;
      RECT  181.9 150.3 188.7 150.9 ;
      RECT  192.2 152.4 193.0 153.2 ;
      RECT  190.2 152.4 191.0 153.2 ;
      RECT  192.2 156.8 193.0 157.6 ;
      RECT  190.2 156.8 191.0 157.6 ;
      RECT  194.2 156.8 195.0 157.6 ;
      RECT  192.2 156.8 193.0 157.6 ;
      RECT  188.7 150.3 195.5 150.9 ;
      RECT  199.0 152.4 199.8 153.2 ;
      RECT  197.0 152.4 197.8 153.2 ;
      RECT  199.0 156.8 199.8 157.6 ;
      RECT  197.0 156.8 197.8 157.6 ;
      RECT  201.0 156.8 201.8 157.6 ;
      RECT  199.0 156.8 199.8 157.6 ;
      RECT  195.5 150.3 202.3 150.9 ;
      RECT  173.0 150.3 202.3 150.9 ;
      RECT  193.3 133.6 194.1 136.0 ;
      RECT  189.9 122.8 191.3 123.4 ;
      RECT  191.7 134.2 192.5 136.0 ;
      RECT  194.1 125.8 194.9 127.0 ;
      RECT  189.9 121.4 190.5 122.8 ;
      RECT  189.3 116.6 190.7 117.2 ;
      RECT  194.9 121.4 195.5 122.8 ;
      RECT  191.9 138.6 192.7 140.4 ;
      RECT  188.3 142.4 195.9 143.2 ;
      RECT  190.5 123.4 191.3 123.6 ;
      RECT  189.9 117.2 190.7 121.4 ;
      RECT  190.1 125.6 191.3 126.4 ;
      RECT  193.1 116.6 193.9 122.2 ;
      RECT  191.7 127.0 194.9 127.6 ;
      RECT  191.3 121.4 192.1 122.2 ;
      RECT  193.3 132.8 194.7 133.6 ;
      RECT  195.1 140.0 195.9 140.8 ;
      RECT  193.5 139.2 195.9 140.0 ;
      RECT  191.9 136.0 192.5 138.6 ;
      RECT  191.5 116.6 192.3 121.4 ;
      RECT  194.7 116.6 195.5 121.4 ;
      RECT  194.5 122.8 195.5 123.6 ;
      RECT  193.3 128.2 194.1 132.8 ;
      RECT  189.3 114.8 190.1 116.6 ;
      RECT  193.5 140.0 194.3 140.4 ;
      RECT  190.1 126.4 190.9 136.0 ;
      RECT  191.7 127.6 192.3 128.2 ;
      RECT  193.5 138.6 194.3 139.2 ;
      RECT  191.7 128.2 192.5 131.8 ;
      RECT  200.1 133.6 200.9 136.0 ;
      RECT  196.7 122.8 198.1 123.4 ;
      RECT  198.5 134.2 199.3 136.0 ;
      RECT  200.9 125.8 201.7 127.0 ;
      RECT  196.7 121.4 197.3 122.8 ;
      RECT  196.1 116.6 197.5 117.2 ;
      RECT  201.7 121.4 202.3 122.8 ;
      RECT  198.7 138.6 199.5 140.4 ;
      RECT  195.1 142.4 202.7 143.2 ;
      RECT  197.3 123.4 198.1 123.6 ;
      RECT  196.7 117.2 197.5 121.4 ;
      RECT  196.9 125.6 198.1 126.4 ;
      RECT  199.9 116.6 200.7 122.2 ;
      RECT  198.5 127.0 201.7 127.6 ;
      RECT  198.1 121.4 198.9 122.2 ;
      RECT  200.1 132.8 201.5 133.6 ;
      RECT  201.9 140.0 202.7 140.8 ;
      RECT  200.3 139.2 202.7 140.0 ;
      RECT  198.7 136.0 199.3 138.6 ;
      RECT  198.3 116.6 199.1 121.4 ;
      RECT  201.5 116.6 202.3 121.4 ;
      RECT  201.3 122.8 202.3 123.6 ;
      RECT  200.1 128.2 200.9 132.8 ;
      RECT  196.1 114.8 196.9 116.6 ;
      RECT  200.3 140.0 201.1 140.4 ;
      RECT  196.9 126.4 197.7 136.0 ;
      RECT  198.5 127.6 199.1 128.2 ;
      RECT  200.3 138.6 201.1 139.2 ;
      RECT  198.5 128.2 199.3 131.8 ;
      RECT  173.0 142.5 202.3 143.1 ;
      RECT  192.5 79.2 193.3 81.4 ;
      RECT  191.1 91.4 192.7 92.2 ;
      RECT  192.9 87.0 194.1 87.8 ;
      RECT  189.7 84.2 190.5 88.0 ;
      RECT  191.1 92.2 191.9 94.2 ;
      RECT  192.9 84.2 194.7 85.6 ;
      RECT  193.3 82.8 194.9 83.6 ;
      RECT  189.7 88.0 193.7 88.6 ;
      RECT  192.9 87.8 193.7 88.0 ;
      RECT  190.9 79.2 191.7 80.6 ;
      RECT  189.5 103.4 190.3 105.8 ;
      RECT  189.7 88.6 190.5 90.6 ;
      RECT  192.9 88.6 193.7 90.6 ;
      RECT  190.9 75.4 191.7 77.4 ;
      RECT  191.3 84.2 192.1 85.6 ;
      RECT  189.3 78.0 190.1 80.6 ;
      RECT  192.7 96.2 193.5 97.4 ;
      RECT  189.3 82.0 190.1 82.8 ;
      RECT  189.3 74.0 193.3 74.8 ;
      RECT  191.7 69.0 192.5 70.6 ;
      RECT  192.7 92.8 193.5 95.4 ;
      RECT  192.7 103.4 193.5 106.6 ;
      RECT  189.3 74.8 190.1 76.8 ;
      RECT  192.5 74.8 193.3 76.8 ;
      RECT  192.7 95.4 195.3 96.2 ;
      RECT  194.3 104.2 195.3 105.0 ;
      RECT  189.5 92.8 190.3 101.4 ;
      RECT  189.3 77.4 191.7 78.0 ;
      RECT  191.1 96.6 191.9 105.8 ;
      RECT  193.7 85.6 194.7 85.8 ;
      RECT  189.3 72.6 194.9 73.4 ;
      RECT  194.7 96.2 195.3 104.2 ;
      RECT  191.3 89.2 192.1 91.4 ;
      RECT  194.1 75.4 194.9 82.8 ;
      RECT  189.7 105.8 190.3 106.4 ;
      RECT  189.5 80.6 190.1 82.0 ;
      RECT  189.7 106.4 191.5 107.2 ;
      RECT  199.3 79.2 200.1 81.4 ;
      RECT  197.9 91.4 199.5 92.2 ;
      RECT  199.7 87.0 200.9 87.8 ;
      RECT  196.5 84.2 197.3 88.0 ;
      RECT  197.9 92.2 198.7 94.2 ;
      RECT  199.7 84.2 201.5 85.6 ;
      RECT  200.1 82.8 201.7 83.6 ;
      RECT  196.5 88.0 200.5 88.6 ;
      RECT  199.7 87.8 200.5 88.0 ;
      RECT  197.7 79.2 198.5 80.6 ;
      RECT  196.3 103.4 197.1 105.8 ;
      RECT  196.5 88.6 197.3 90.6 ;
      RECT  199.7 88.6 200.5 90.6 ;
      RECT  197.7 75.4 198.5 77.4 ;
      RECT  198.1 84.2 198.9 85.6 ;
      RECT  196.1 78.0 196.9 80.6 ;
      RECT  199.5 96.2 200.3 97.4 ;
      RECT  196.1 82.0 196.9 82.8 ;
      RECT  196.1 74.0 200.1 74.8 ;
      RECT  198.5 69.0 199.3 70.6 ;
      RECT  199.5 92.8 200.3 95.4 ;
      RECT  199.5 103.4 200.3 106.6 ;
      RECT  196.1 74.8 196.9 76.8 ;
      RECT  199.3 74.8 200.1 76.8 ;
      RECT  199.5 95.4 202.1 96.2 ;
      RECT  201.1 104.2 202.1 105.0 ;
      RECT  196.3 92.8 197.1 101.4 ;
      RECT  196.1 77.4 198.5 78.0 ;
      RECT  197.9 96.6 198.7 105.8 ;
      RECT  200.5 85.6 201.5 85.8 ;
      RECT  196.1 72.6 201.7 73.4 ;
      RECT  201.5 96.2 202.1 104.2 ;
      RECT  198.1 89.2 198.9 91.4 ;
      RECT  200.9 75.4 201.7 82.8 ;
      RECT  196.5 105.8 197.1 106.4 ;
      RECT  196.3 80.6 196.9 82.0 ;
      RECT  196.5 106.4 198.3 107.2 ;
      RECT  173.0 72.6 202.3 73.2 ;
      RECT  173.0 143.1 202.3 142.5 ;
      RECT  173.0 150.9 202.3 150.3 ;
      RECT  173.0 73.2 202.3 72.6 ;
      RECT  97.3 194.7 98.1 195.5 ;
      RECT  95.3 194.7 96.1 195.5 ;
      RECT  97.3 187.3 98.1 188.1 ;
      RECT  95.3 187.3 96.1 188.1 ;
      RECT  95.7 191.0 96.5 191.8 ;
      RECT  97.7 191.1 98.3 191.7 ;
      RECT  94.1 196.5 100.7 197.1 ;
      RECT  94.1 186.1 100.7 186.7 ;
      RECT  97.3 198.9 98.1 198.1 ;
      RECT  95.3 198.9 96.1 198.1 ;
      RECT  97.3 206.3 98.1 205.5 ;
      RECT  95.3 206.3 96.1 205.5 ;
      RECT  95.7 202.6 96.5 201.8 ;
      RECT  97.7 202.5 98.3 201.9 ;
      RECT  94.1 197.1 100.7 196.5 ;
      RECT  94.1 207.5 100.7 206.9 ;
      RECT  112.3 194.7 113.1 195.5 ;
      RECT  110.3 194.7 111.1 195.5 ;
      RECT  114.3 194.7 115.1 195.5 ;
      RECT  112.3 194.7 113.1 195.5 ;
      RECT  110.3 187.7 111.1 188.5 ;
      RECT  114.3 187.7 115.1 188.5 ;
      RECT  111.3 189.2 112.1 190.0 ;
      RECT  113.3 192.0 114.1 192.8 ;
      RECT  115.8 193.4 116.4 194.0 ;
      RECT  109.1 196.5 117.7 197.1 ;
      RECT  109.1 186.1 117.7 186.7 ;
      RECT  120.9 194.7 121.7 195.5 ;
      RECT  118.9 194.7 119.7 195.5 ;
      RECT  120.9 187.3 121.7 188.1 ;
      RECT  118.9 187.3 119.7 188.1 ;
      RECT  119.3 191.0 120.1 191.8 ;
      RECT  121.3 191.1 121.9 191.7 ;
      RECT  117.7 196.5 124.3 197.1 ;
      RECT  117.7 186.1 124.3 186.7 ;
      RECT  111.3 189.2 112.1 190.0 ;
      RECT  113.3 192.0 114.1 192.8 ;
      RECT  121.3 191.1 121.9 191.7 ;
      RECT  109.1 196.5 124.3 197.1 ;
      RECT  109.1 186.1 124.3 186.7 ;
      RECT  112.3 198.9 113.1 198.1 ;
      RECT  110.3 198.9 111.1 198.1 ;
      RECT  114.3 198.9 115.1 198.1 ;
      RECT  112.3 198.9 113.1 198.1 ;
      RECT  110.3 205.9 111.1 205.1 ;
      RECT  114.3 205.9 115.1 205.1 ;
      RECT  111.3 204.4 112.1 203.6 ;
      RECT  113.3 201.6 114.1 200.8 ;
      RECT  115.8 200.2 116.4 199.6 ;
      RECT  109.1 197.1 117.7 196.5 ;
      RECT  109.1 207.5 117.7 206.9 ;
      RECT  120.9 198.9 121.7 198.1 ;
      RECT  118.9 198.9 119.7 198.1 ;
      RECT  120.9 206.3 121.7 205.5 ;
      RECT  118.9 206.3 119.7 205.5 ;
      RECT  119.3 202.6 120.1 201.8 ;
      RECT  121.3 202.5 121.9 201.9 ;
      RECT  117.7 197.1 124.3 196.5 ;
      RECT  117.7 207.5 124.3 206.9 ;
      RECT  111.3 204.4 112.1 203.6 ;
      RECT  113.3 201.6 114.1 200.8 ;
      RECT  121.3 202.5 121.9 201.9 ;
      RECT  109.1 197.1 124.3 196.5 ;
      RECT  109.1 207.5 124.3 206.9 ;
      RECT  112.3 215.5 113.1 216.3 ;
      RECT  110.3 215.5 111.1 216.3 ;
      RECT  114.3 215.5 115.1 216.3 ;
      RECT  112.3 215.5 113.1 216.3 ;
      RECT  110.3 208.5 111.1 209.3 ;
      RECT  114.3 208.5 115.1 209.3 ;
      RECT  111.3 210.0 112.1 210.8 ;
      RECT  113.3 212.8 114.1 213.6 ;
      RECT  115.8 214.2 116.4 214.8 ;
      RECT  109.1 217.3 117.7 217.9 ;
      RECT  109.1 206.9 117.7 207.5 ;
      RECT  120.9 215.5 121.7 216.3 ;
      RECT  118.9 215.5 119.7 216.3 ;
      RECT  120.9 208.1 121.7 208.9 ;
      RECT  118.9 208.1 119.7 208.9 ;
      RECT  119.3 211.8 120.1 212.6 ;
      RECT  121.3 211.9 121.9 212.5 ;
      RECT  117.7 217.3 124.3 217.9 ;
      RECT  117.7 206.9 124.3 207.5 ;
      RECT  111.3 210.0 112.1 210.8 ;
      RECT  113.3 212.8 114.1 213.6 ;
      RECT  121.3 211.9 121.9 212.5 ;
      RECT  109.1 217.3 124.3 217.9 ;
      RECT  109.1 206.9 124.3 207.5 ;
      RECT  112.3 219.7 113.1 218.9 ;
      RECT  110.3 219.7 111.1 218.9 ;
      RECT  114.3 219.7 115.1 218.9 ;
      RECT  112.3 219.7 113.1 218.9 ;
      RECT  110.3 226.7 111.1 225.9 ;
      RECT  114.3 226.7 115.1 225.9 ;
      RECT  111.3 225.2 112.1 224.4 ;
      RECT  113.3 222.4 114.1 221.6 ;
      RECT  115.8 221.0 116.4 220.4 ;
      RECT  109.1 217.9 117.7 217.3 ;
      RECT  109.1 228.3 117.7 227.7 ;
      RECT  120.9 219.7 121.7 218.9 ;
      RECT  118.9 219.7 119.7 218.9 ;
      RECT  120.9 227.1 121.7 226.3 ;
      RECT  118.9 227.1 119.7 226.3 ;
      RECT  119.3 223.4 120.1 222.6 ;
      RECT  121.3 223.3 121.9 222.7 ;
      RECT  117.7 217.9 124.3 217.3 ;
      RECT  117.7 228.3 124.3 227.7 ;
      RECT  111.3 225.2 112.1 224.4 ;
      RECT  113.3 222.4 114.1 221.6 ;
      RECT  121.3 223.3 121.9 222.7 ;
      RECT  109.1 217.9 124.3 217.3 ;
      RECT  109.1 228.3 124.3 227.7 ;
      RECT  121.3 191.1 121.9 191.7 ;
      RECT  121.3 201.9 121.9 202.5 ;
      RECT  121.3 211.9 121.9 212.5 ;
      RECT  121.3 222.7 121.9 223.3 ;
      RECT  97.3 257.1 98.1 257.9 ;
      RECT  95.3 257.1 96.1 257.9 ;
      RECT  97.3 249.7 98.1 250.5 ;
      RECT  95.3 249.7 96.1 250.5 ;
      RECT  95.7 253.4 96.5 254.2 ;
      RECT  97.7 253.5 98.3 254.1 ;
      RECT  94.1 258.9 100.7 259.5 ;
      RECT  94.1 248.5 100.7 249.1 ;
      RECT  97.3 261.3 98.1 260.5 ;
      RECT  95.3 261.3 96.1 260.5 ;
      RECT  97.3 268.7 98.1 267.9 ;
      RECT  95.3 268.7 96.1 267.9 ;
      RECT  95.7 265.0 96.5 264.2 ;
      RECT  97.7 264.9 98.3 264.3 ;
      RECT  94.1 259.5 100.7 258.9 ;
      RECT  94.1 269.9 100.7 269.3 ;
      RECT  112.3 257.1 113.1 257.9 ;
      RECT  110.3 257.1 111.1 257.9 ;
      RECT  114.3 257.1 115.1 257.9 ;
      RECT  112.3 257.1 113.1 257.9 ;
      RECT  110.3 250.1 111.1 250.9 ;
      RECT  114.3 250.1 115.1 250.9 ;
      RECT  111.3 251.6 112.1 252.4 ;
      RECT  113.3 254.4 114.1 255.2 ;
      RECT  115.8 255.8 116.4 256.4 ;
      RECT  109.1 258.9 117.7 259.5 ;
      RECT  109.1 248.5 117.7 249.1 ;
      RECT  120.9 257.1 121.7 257.9 ;
      RECT  118.9 257.1 119.7 257.9 ;
      RECT  120.9 249.7 121.7 250.5 ;
      RECT  118.9 249.7 119.7 250.5 ;
      RECT  119.3 253.4 120.1 254.2 ;
      RECT  121.3 253.5 121.9 254.1 ;
      RECT  117.7 258.9 124.3 259.5 ;
      RECT  117.7 248.5 124.3 249.1 ;
      RECT  111.3 251.6 112.1 252.4 ;
      RECT  113.3 254.4 114.1 255.2 ;
      RECT  121.3 253.5 121.9 254.1 ;
      RECT  109.1 258.9 124.3 259.5 ;
      RECT  109.1 248.5 124.3 249.1 ;
      RECT  112.3 261.3 113.1 260.5 ;
      RECT  110.3 261.3 111.1 260.5 ;
      RECT  114.3 261.3 115.1 260.5 ;
      RECT  112.3 261.3 113.1 260.5 ;
      RECT  110.3 268.3 111.1 267.5 ;
      RECT  114.3 268.3 115.1 267.5 ;
      RECT  111.3 266.8 112.1 266.0 ;
      RECT  113.3 264.0 114.1 263.2 ;
      RECT  115.8 262.6 116.4 262.0 ;
      RECT  109.1 259.5 117.7 258.9 ;
      RECT  109.1 269.9 117.7 269.3 ;
      RECT  120.9 261.3 121.7 260.5 ;
      RECT  118.9 261.3 119.7 260.5 ;
      RECT  120.9 268.7 121.7 267.9 ;
      RECT  118.9 268.7 119.7 267.9 ;
      RECT  119.3 265.0 120.1 264.2 ;
      RECT  121.3 264.9 121.9 264.3 ;
      RECT  117.7 259.5 124.3 258.9 ;
      RECT  117.7 269.9 124.3 269.3 ;
      RECT  111.3 266.8 112.1 266.0 ;
      RECT  113.3 264.0 114.1 263.2 ;
      RECT  121.3 264.9 121.9 264.3 ;
      RECT  109.1 259.5 124.3 258.9 ;
      RECT  109.1 269.9 124.3 269.3 ;
      RECT  112.3 277.9 113.1 278.7 ;
      RECT  110.3 277.9 111.1 278.7 ;
      RECT  114.3 277.9 115.1 278.7 ;
      RECT  112.3 277.9 113.1 278.7 ;
      RECT  110.3 270.9 111.1 271.7 ;
      RECT  114.3 270.9 115.1 271.7 ;
      RECT  111.3 272.4 112.1 273.2 ;
      RECT  113.3 275.2 114.1 276.0 ;
      RECT  115.8 276.6 116.4 277.2 ;
      RECT  109.1 279.7 117.7 280.3 ;
      RECT  109.1 269.3 117.7 269.9 ;
      RECT  120.9 277.9 121.7 278.7 ;
      RECT  118.9 277.9 119.7 278.7 ;
      RECT  120.9 270.5 121.7 271.3 ;
      RECT  118.9 270.5 119.7 271.3 ;
      RECT  119.3 274.2 120.1 275.0 ;
      RECT  121.3 274.3 121.9 274.9 ;
      RECT  117.7 279.7 124.3 280.3 ;
      RECT  117.7 269.3 124.3 269.9 ;
      RECT  111.3 272.4 112.1 273.2 ;
      RECT  113.3 275.2 114.1 276.0 ;
      RECT  121.3 274.3 121.9 274.9 ;
      RECT  109.1 279.7 124.3 280.3 ;
      RECT  109.1 269.3 124.3 269.9 ;
      RECT  112.3 282.1 113.1 281.3 ;
      RECT  110.3 282.1 111.1 281.3 ;
      RECT  114.3 282.1 115.1 281.3 ;
      RECT  112.3 282.1 113.1 281.3 ;
      RECT  110.3 289.1 111.1 288.3 ;
      RECT  114.3 289.1 115.1 288.3 ;
      RECT  111.3 287.6 112.1 286.8 ;
      RECT  113.3 284.8 114.1 284.0 ;
      RECT  115.8 283.4 116.4 282.8 ;
      RECT  109.1 280.3 117.7 279.7 ;
      RECT  109.1 290.7 117.7 290.1 ;
      RECT  120.9 282.1 121.7 281.3 ;
      RECT  118.9 282.1 119.7 281.3 ;
      RECT  120.9 289.5 121.7 288.7 ;
      RECT  118.9 289.5 119.7 288.7 ;
      RECT  119.3 285.8 120.1 285.0 ;
      RECT  121.3 285.7 121.9 285.1 ;
      RECT  117.7 280.3 124.3 279.7 ;
      RECT  117.7 290.7 124.3 290.1 ;
      RECT  111.3 287.6 112.1 286.8 ;
      RECT  113.3 284.8 114.1 284.0 ;
      RECT  121.3 285.7 121.9 285.1 ;
      RECT  109.1 280.3 124.3 279.7 ;
      RECT  109.1 290.7 124.3 290.1 ;
      RECT  121.3 253.5 121.9 254.1 ;
      RECT  121.3 264.3 121.9 264.9 ;
      RECT  121.3 274.3 121.9 274.9 ;
      RECT  121.3 285.1 121.9 285.7 ;
      RECT  140.1 194.7 140.9 195.5 ;
      RECT  138.1 194.7 138.9 195.5 ;
      RECT  142.1 194.7 142.9 195.5 ;
      RECT  140.1 194.7 140.9 195.5 ;
      RECT  138.1 187.7 138.9 188.5 ;
      RECT  142.1 187.7 142.9 188.5 ;
      RECT  139.1 189.2 139.9 190.0 ;
      RECT  141.1 192.0 141.9 192.8 ;
      RECT  143.6 193.4 144.2 194.0 ;
      RECT  136.9 196.5 145.5 197.1 ;
      RECT  136.9 186.1 145.5 186.7 ;
      RECT  148.7 194.7 149.5 195.5 ;
      RECT  146.7 194.7 147.5 195.5 ;
      RECT  148.7 187.3 149.5 188.1 ;
      RECT  146.7 187.3 147.5 188.1 ;
      RECT  147.1 191.0 147.9 191.8 ;
      RECT  149.1 191.1 149.7 191.7 ;
      RECT  145.5 196.5 152.1 197.1 ;
      RECT  145.5 186.1 152.1 186.7 ;
      RECT  139.1 189.2 139.9 190.0 ;
      RECT  141.1 192.0 141.9 192.8 ;
      RECT  149.1 191.1 149.7 191.7 ;
      RECT  136.9 196.5 152.1 197.1 ;
      RECT  136.9 186.1 152.1 186.7 ;
      RECT  140.1 198.9 140.9 198.1 ;
      RECT  138.1 198.9 138.9 198.1 ;
      RECT  142.1 198.9 142.9 198.1 ;
      RECT  140.1 198.9 140.9 198.1 ;
      RECT  138.1 205.9 138.9 205.1 ;
      RECT  142.1 205.9 142.9 205.1 ;
      RECT  139.1 204.4 139.9 203.6 ;
      RECT  141.1 201.6 141.9 200.8 ;
      RECT  143.6 200.2 144.2 199.6 ;
      RECT  136.9 197.1 145.5 196.5 ;
      RECT  136.9 207.5 145.5 206.9 ;
      RECT  148.7 198.9 149.5 198.1 ;
      RECT  146.7 198.9 147.5 198.1 ;
      RECT  148.7 206.3 149.5 205.5 ;
      RECT  146.7 206.3 147.5 205.5 ;
      RECT  147.1 202.6 147.9 201.8 ;
      RECT  149.1 202.5 149.7 201.9 ;
      RECT  145.5 197.1 152.1 196.5 ;
      RECT  145.5 207.5 152.1 206.9 ;
      RECT  139.1 204.4 139.9 203.6 ;
      RECT  141.1 201.6 141.9 200.8 ;
      RECT  149.1 202.5 149.7 201.9 ;
      RECT  136.9 197.1 152.1 196.5 ;
      RECT  136.9 207.5 152.1 206.9 ;
      RECT  140.1 215.5 140.9 216.3 ;
      RECT  138.1 215.5 138.9 216.3 ;
      RECT  142.1 215.5 142.9 216.3 ;
      RECT  140.1 215.5 140.9 216.3 ;
      RECT  138.1 208.5 138.9 209.3 ;
      RECT  142.1 208.5 142.9 209.3 ;
      RECT  139.1 210.0 139.9 210.8 ;
      RECT  141.1 212.8 141.9 213.6 ;
      RECT  143.6 214.2 144.2 214.8 ;
      RECT  136.9 217.3 145.5 217.9 ;
      RECT  136.9 206.9 145.5 207.5 ;
      RECT  148.7 215.5 149.5 216.3 ;
      RECT  146.7 215.5 147.5 216.3 ;
      RECT  148.7 208.1 149.5 208.9 ;
      RECT  146.7 208.1 147.5 208.9 ;
      RECT  147.1 211.8 147.9 212.6 ;
      RECT  149.1 211.9 149.7 212.5 ;
      RECT  145.5 217.3 152.1 217.9 ;
      RECT  145.5 206.9 152.1 207.5 ;
      RECT  139.1 210.0 139.9 210.8 ;
      RECT  141.1 212.8 141.9 213.6 ;
      RECT  149.1 211.9 149.7 212.5 ;
      RECT  136.9 217.3 152.1 217.9 ;
      RECT  136.9 206.9 152.1 207.5 ;
      RECT  140.1 219.7 140.9 218.9 ;
      RECT  138.1 219.7 138.9 218.9 ;
      RECT  142.1 219.7 142.9 218.9 ;
      RECT  140.1 219.7 140.9 218.9 ;
      RECT  138.1 226.7 138.9 225.9 ;
      RECT  142.1 226.7 142.9 225.9 ;
      RECT  139.1 225.2 139.9 224.4 ;
      RECT  141.1 222.4 141.9 221.6 ;
      RECT  143.6 221.0 144.2 220.4 ;
      RECT  136.9 217.9 145.5 217.3 ;
      RECT  136.9 228.3 145.5 227.7 ;
      RECT  148.7 219.7 149.5 218.9 ;
      RECT  146.7 219.7 147.5 218.9 ;
      RECT  148.7 227.1 149.5 226.3 ;
      RECT  146.7 227.1 147.5 226.3 ;
      RECT  147.1 223.4 147.9 222.6 ;
      RECT  149.1 223.3 149.7 222.7 ;
      RECT  145.5 217.9 152.1 217.3 ;
      RECT  145.5 228.3 152.1 227.7 ;
      RECT  139.1 225.2 139.9 224.4 ;
      RECT  141.1 222.4 141.9 221.6 ;
      RECT  149.1 223.3 149.7 222.7 ;
      RECT  136.9 217.9 152.1 217.3 ;
      RECT  136.9 228.3 152.1 227.7 ;
      RECT  140.1 236.3 140.9 237.1 ;
      RECT  138.1 236.3 138.9 237.1 ;
      RECT  142.1 236.3 142.9 237.1 ;
      RECT  140.1 236.3 140.9 237.1 ;
      RECT  138.1 229.3 138.9 230.1 ;
      RECT  142.1 229.3 142.9 230.1 ;
      RECT  139.1 230.8 139.9 231.6 ;
      RECT  141.1 233.6 141.9 234.4 ;
      RECT  143.6 235.0 144.2 235.6 ;
      RECT  136.9 238.1 145.5 238.7 ;
      RECT  136.9 227.7 145.5 228.3 ;
      RECT  148.7 236.3 149.5 237.1 ;
      RECT  146.7 236.3 147.5 237.1 ;
      RECT  148.7 228.9 149.5 229.7 ;
      RECT  146.7 228.9 147.5 229.7 ;
      RECT  147.1 232.6 147.9 233.4 ;
      RECT  149.1 232.7 149.7 233.3 ;
      RECT  145.5 238.1 152.1 238.7 ;
      RECT  145.5 227.7 152.1 228.3 ;
      RECT  139.1 230.8 139.9 231.6 ;
      RECT  141.1 233.6 141.9 234.4 ;
      RECT  149.1 232.7 149.7 233.3 ;
      RECT  136.9 238.1 152.1 238.7 ;
      RECT  136.9 227.7 152.1 228.3 ;
      RECT  140.1 240.5 140.9 239.7 ;
      RECT  138.1 240.5 138.9 239.7 ;
      RECT  142.1 240.5 142.9 239.7 ;
      RECT  140.1 240.5 140.9 239.7 ;
      RECT  138.1 247.5 138.9 246.7 ;
      RECT  142.1 247.5 142.9 246.7 ;
      RECT  139.1 246.0 139.9 245.2 ;
      RECT  141.1 243.2 141.9 242.4 ;
      RECT  143.6 241.8 144.2 241.2 ;
      RECT  136.9 238.7 145.5 238.1 ;
      RECT  136.9 249.1 145.5 248.5 ;
      RECT  148.7 240.5 149.5 239.7 ;
      RECT  146.7 240.5 147.5 239.7 ;
      RECT  148.7 247.9 149.5 247.1 ;
      RECT  146.7 247.9 147.5 247.1 ;
      RECT  147.1 244.2 147.9 243.4 ;
      RECT  149.1 244.1 149.7 243.5 ;
      RECT  145.5 238.7 152.1 238.1 ;
      RECT  145.5 249.1 152.1 248.5 ;
      RECT  139.1 246.0 139.9 245.2 ;
      RECT  141.1 243.2 141.9 242.4 ;
      RECT  149.1 244.1 149.7 243.5 ;
      RECT  136.9 238.7 152.1 238.1 ;
      RECT  136.9 249.1 152.1 248.5 ;
      RECT  140.1 257.1 140.9 257.9 ;
      RECT  138.1 257.1 138.9 257.9 ;
      RECT  142.1 257.1 142.9 257.9 ;
      RECT  140.1 257.1 140.9 257.9 ;
      RECT  138.1 250.1 138.9 250.9 ;
      RECT  142.1 250.1 142.9 250.9 ;
      RECT  139.1 251.6 139.9 252.4 ;
      RECT  141.1 254.4 141.9 255.2 ;
      RECT  143.6 255.8 144.2 256.4 ;
      RECT  136.9 258.9 145.5 259.5 ;
      RECT  136.9 248.5 145.5 249.1 ;
      RECT  148.7 257.1 149.5 257.9 ;
      RECT  146.7 257.1 147.5 257.9 ;
      RECT  148.7 249.7 149.5 250.5 ;
      RECT  146.7 249.7 147.5 250.5 ;
      RECT  147.1 253.4 147.9 254.2 ;
      RECT  149.1 253.5 149.7 254.1 ;
      RECT  145.5 258.9 152.1 259.5 ;
      RECT  145.5 248.5 152.1 249.1 ;
      RECT  139.1 251.6 139.9 252.4 ;
      RECT  141.1 254.4 141.9 255.2 ;
      RECT  149.1 253.5 149.7 254.1 ;
      RECT  136.9 258.9 152.1 259.5 ;
      RECT  136.9 248.5 152.1 249.1 ;
      RECT  140.1 261.3 140.9 260.5 ;
      RECT  138.1 261.3 138.9 260.5 ;
      RECT  142.1 261.3 142.9 260.5 ;
      RECT  140.1 261.3 140.9 260.5 ;
      RECT  138.1 268.3 138.9 267.5 ;
      RECT  142.1 268.3 142.9 267.5 ;
      RECT  139.1 266.8 139.9 266.0 ;
      RECT  141.1 264.0 141.9 263.2 ;
      RECT  143.6 262.6 144.2 262.0 ;
      RECT  136.9 259.5 145.5 258.9 ;
      RECT  136.9 269.9 145.5 269.3 ;
      RECT  148.7 261.3 149.5 260.5 ;
      RECT  146.7 261.3 147.5 260.5 ;
      RECT  148.7 268.7 149.5 267.9 ;
      RECT  146.7 268.7 147.5 267.9 ;
      RECT  147.1 265.0 147.9 264.2 ;
      RECT  149.1 264.9 149.7 264.3 ;
      RECT  145.5 259.5 152.1 258.9 ;
      RECT  145.5 269.9 152.1 269.3 ;
      RECT  139.1 266.8 139.9 266.0 ;
      RECT  141.1 264.0 141.9 263.2 ;
      RECT  149.1 264.9 149.7 264.3 ;
      RECT  136.9 259.5 152.1 258.9 ;
      RECT  136.9 269.9 152.1 269.3 ;
      RECT  140.1 277.9 140.9 278.7 ;
      RECT  138.1 277.9 138.9 278.7 ;
      RECT  142.1 277.9 142.9 278.7 ;
      RECT  140.1 277.9 140.9 278.7 ;
      RECT  138.1 270.9 138.9 271.7 ;
      RECT  142.1 270.9 142.9 271.7 ;
      RECT  139.1 272.4 139.9 273.2 ;
      RECT  141.1 275.2 141.9 276.0 ;
      RECT  143.6 276.6 144.2 277.2 ;
      RECT  136.9 279.7 145.5 280.3 ;
      RECT  136.9 269.3 145.5 269.9 ;
      RECT  148.7 277.9 149.5 278.7 ;
      RECT  146.7 277.9 147.5 278.7 ;
      RECT  148.7 270.5 149.5 271.3 ;
      RECT  146.7 270.5 147.5 271.3 ;
      RECT  147.1 274.2 147.9 275.0 ;
      RECT  149.1 274.3 149.7 274.9 ;
      RECT  145.5 279.7 152.1 280.3 ;
      RECT  145.5 269.3 152.1 269.9 ;
      RECT  139.1 272.4 139.9 273.2 ;
      RECT  141.1 275.2 141.9 276.0 ;
      RECT  149.1 274.3 149.7 274.9 ;
      RECT  136.9 279.7 152.1 280.3 ;
      RECT  136.9 269.3 152.1 269.9 ;
      RECT  140.1 282.1 140.9 281.3 ;
      RECT  138.1 282.1 138.9 281.3 ;
      RECT  142.1 282.1 142.9 281.3 ;
      RECT  140.1 282.1 140.9 281.3 ;
      RECT  138.1 289.1 138.9 288.3 ;
      RECT  142.1 289.1 142.9 288.3 ;
      RECT  139.1 287.6 139.9 286.8 ;
      RECT  141.1 284.8 141.9 284.0 ;
      RECT  143.6 283.4 144.2 282.8 ;
      RECT  136.9 280.3 145.5 279.7 ;
      RECT  136.9 290.7 145.5 290.1 ;
      RECT  148.7 282.1 149.5 281.3 ;
      RECT  146.7 282.1 147.5 281.3 ;
      RECT  148.7 289.5 149.5 288.7 ;
      RECT  146.7 289.5 147.5 288.7 ;
      RECT  147.1 285.8 147.9 285.0 ;
      RECT  149.1 285.7 149.7 285.1 ;
      RECT  145.5 280.3 152.1 279.7 ;
      RECT  145.5 290.7 152.1 290.1 ;
      RECT  139.1 287.6 139.9 286.8 ;
      RECT  141.1 284.8 141.9 284.0 ;
      RECT  149.1 285.7 149.7 285.1 ;
      RECT  136.9 280.3 152.1 279.7 ;
      RECT  136.9 290.7 152.1 290.1 ;
      RECT  140.1 298.7 140.9 299.5 ;
      RECT  138.1 298.7 138.9 299.5 ;
      RECT  142.1 298.7 142.9 299.5 ;
      RECT  140.1 298.7 140.9 299.5 ;
      RECT  138.1 291.7 138.9 292.5 ;
      RECT  142.1 291.7 142.9 292.5 ;
      RECT  139.1 293.2 139.9 294.0 ;
      RECT  141.1 296.0 141.9 296.8 ;
      RECT  143.6 297.4 144.2 298.0 ;
      RECT  136.9 300.5 145.5 301.1 ;
      RECT  136.9 290.1 145.5 290.7 ;
      RECT  148.7 298.7 149.5 299.5 ;
      RECT  146.7 298.7 147.5 299.5 ;
      RECT  148.7 291.3 149.5 292.1 ;
      RECT  146.7 291.3 147.5 292.1 ;
      RECT  147.1 295.0 147.9 295.8 ;
      RECT  149.1 295.1 149.7 295.7 ;
      RECT  145.5 300.5 152.1 301.1 ;
      RECT  145.5 290.1 152.1 290.7 ;
      RECT  139.1 293.2 139.9 294.0 ;
      RECT  141.1 296.0 141.9 296.8 ;
      RECT  149.1 295.1 149.7 295.7 ;
      RECT  136.9 300.5 152.1 301.1 ;
      RECT  136.9 290.1 152.1 290.7 ;
      RECT  140.1 302.9 140.9 302.1 ;
      RECT  138.1 302.9 138.9 302.1 ;
      RECT  142.1 302.9 142.9 302.1 ;
      RECT  140.1 302.9 140.9 302.1 ;
      RECT  138.1 309.9 138.9 309.1 ;
      RECT  142.1 309.9 142.9 309.1 ;
      RECT  139.1 308.4 139.9 307.6 ;
      RECT  141.1 305.6 141.9 304.8 ;
      RECT  143.6 304.2 144.2 303.6 ;
      RECT  136.9 301.1 145.5 300.5 ;
      RECT  136.9 311.5 145.5 310.9 ;
      RECT  148.7 302.9 149.5 302.1 ;
      RECT  146.7 302.9 147.5 302.1 ;
      RECT  148.7 310.3 149.5 309.5 ;
      RECT  146.7 310.3 147.5 309.5 ;
      RECT  147.1 306.6 147.9 305.8 ;
      RECT  149.1 306.5 149.7 305.9 ;
      RECT  145.5 301.1 152.1 300.5 ;
      RECT  145.5 311.5 152.1 310.9 ;
      RECT  139.1 308.4 139.9 307.6 ;
      RECT  141.1 305.6 141.9 304.8 ;
      RECT  149.1 306.5 149.7 305.9 ;
      RECT  136.9 301.1 152.1 300.5 ;
      RECT  136.9 311.5 152.1 310.9 ;
      RECT  140.1 319.5 140.9 320.3 ;
      RECT  138.1 319.5 138.9 320.3 ;
      RECT  142.1 319.5 142.9 320.3 ;
      RECT  140.1 319.5 140.9 320.3 ;
      RECT  138.1 312.5 138.9 313.3 ;
      RECT  142.1 312.5 142.9 313.3 ;
      RECT  139.1 314.0 139.9 314.8 ;
      RECT  141.1 316.8 141.9 317.6 ;
      RECT  143.6 318.2 144.2 318.8 ;
      RECT  136.9 321.3 145.5 321.9 ;
      RECT  136.9 310.9 145.5 311.5 ;
      RECT  148.7 319.5 149.5 320.3 ;
      RECT  146.7 319.5 147.5 320.3 ;
      RECT  148.7 312.1 149.5 312.9 ;
      RECT  146.7 312.1 147.5 312.9 ;
      RECT  147.1 315.8 147.9 316.6 ;
      RECT  149.1 315.9 149.7 316.5 ;
      RECT  145.5 321.3 152.1 321.9 ;
      RECT  145.5 310.9 152.1 311.5 ;
      RECT  139.1 314.0 139.9 314.8 ;
      RECT  141.1 316.8 141.9 317.6 ;
      RECT  149.1 315.9 149.7 316.5 ;
      RECT  136.9 321.3 152.1 321.9 ;
      RECT  136.9 310.9 152.1 311.5 ;
      RECT  140.1 323.7 140.9 322.9 ;
      RECT  138.1 323.7 138.9 322.9 ;
      RECT  142.1 323.7 142.9 322.9 ;
      RECT  140.1 323.7 140.9 322.9 ;
      RECT  138.1 330.7 138.9 329.9 ;
      RECT  142.1 330.7 142.9 329.9 ;
      RECT  139.1 329.2 139.9 328.4 ;
      RECT  141.1 326.4 141.9 325.6 ;
      RECT  143.6 325.0 144.2 324.4 ;
      RECT  136.9 321.9 145.5 321.3 ;
      RECT  136.9 332.3 145.5 331.7 ;
      RECT  148.7 323.7 149.5 322.9 ;
      RECT  146.7 323.7 147.5 322.9 ;
      RECT  148.7 331.1 149.5 330.3 ;
      RECT  146.7 331.1 147.5 330.3 ;
      RECT  147.1 327.4 147.9 326.6 ;
      RECT  149.1 327.3 149.7 326.7 ;
      RECT  145.5 321.9 152.1 321.3 ;
      RECT  145.5 332.3 152.1 331.7 ;
      RECT  139.1 329.2 139.9 328.4 ;
      RECT  141.1 326.4 141.9 325.6 ;
      RECT  149.1 327.3 149.7 326.7 ;
      RECT  136.9 321.9 152.1 321.3 ;
      RECT  136.9 332.3 152.1 331.7 ;
      RECT  140.1 340.3 140.9 341.1 ;
      RECT  138.1 340.3 138.9 341.1 ;
      RECT  142.1 340.3 142.9 341.1 ;
      RECT  140.1 340.3 140.9 341.1 ;
      RECT  138.1 333.3 138.9 334.1 ;
      RECT  142.1 333.3 142.9 334.1 ;
      RECT  139.1 334.8 139.9 335.6 ;
      RECT  141.1 337.6 141.9 338.4 ;
      RECT  143.6 339.0 144.2 339.6 ;
      RECT  136.9 342.1 145.5 342.7 ;
      RECT  136.9 331.7 145.5 332.3 ;
      RECT  148.7 340.3 149.5 341.1 ;
      RECT  146.7 340.3 147.5 341.1 ;
      RECT  148.7 332.9 149.5 333.7 ;
      RECT  146.7 332.9 147.5 333.7 ;
      RECT  147.1 336.6 147.9 337.4 ;
      RECT  149.1 336.7 149.7 337.3 ;
      RECT  145.5 342.1 152.1 342.7 ;
      RECT  145.5 331.7 152.1 332.3 ;
      RECT  139.1 334.8 139.9 335.6 ;
      RECT  141.1 337.6 141.9 338.4 ;
      RECT  149.1 336.7 149.7 337.3 ;
      RECT  136.9 342.1 152.1 342.7 ;
      RECT  136.9 331.7 152.1 332.3 ;
      RECT  140.1 344.5 140.9 343.7 ;
      RECT  138.1 344.5 138.9 343.7 ;
      RECT  142.1 344.5 142.9 343.7 ;
      RECT  140.1 344.5 140.9 343.7 ;
      RECT  138.1 351.5 138.9 350.7 ;
      RECT  142.1 351.5 142.9 350.7 ;
      RECT  139.1 350.0 139.9 349.2 ;
      RECT  141.1 347.2 141.9 346.4 ;
      RECT  143.6 345.8 144.2 345.2 ;
      RECT  136.9 342.7 145.5 342.1 ;
      RECT  136.9 353.1 145.5 352.5 ;
      RECT  148.7 344.5 149.5 343.7 ;
      RECT  146.7 344.5 147.5 343.7 ;
      RECT  148.7 351.9 149.5 351.1 ;
      RECT  146.7 351.9 147.5 351.1 ;
      RECT  147.1 348.2 147.9 347.4 ;
      RECT  149.1 348.1 149.7 347.5 ;
      RECT  145.5 342.7 152.1 342.1 ;
      RECT  145.5 353.1 152.1 352.5 ;
      RECT  139.1 350.0 139.9 349.2 ;
      RECT  141.1 347.2 141.9 346.4 ;
      RECT  149.1 348.1 149.7 347.5 ;
      RECT  136.9 342.7 152.1 342.1 ;
      RECT  136.9 353.1 152.1 352.5 ;
      RECT  149.1 191.1 149.7 191.7 ;
      RECT  149.1 201.9 149.7 202.5 ;
      RECT  149.1 211.9 149.7 212.5 ;
      RECT  149.1 222.7 149.7 223.3 ;
      RECT  149.1 232.7 149.7 233.3 ;
      RECT  149.1 243.5 149.7 244.1 ;
      RECT  149.1 253.5 149.7 254.1 ;
      RECT  149.1 264.3 149.7 264.9 ;
      RECT  149.1 274.3 149.7 274.9 ;
      RECT  149.1 285.1 149.7 285.7 ;
      RECT  149.1 295.1 149.7 295.7 ;
      RECT  149.1 305.9 149.7 306.5 ;
      RECT  149.1 315.9 149.7 316.5 ;
      RECT  149.1 326.7 149.7 327.3 ;
      RECT  149.1 336.7 149.7 337.3 ;
      RECT  149.1 347.5 149.7 348.1 ;
      RECT  155.6 194.7 156.4 195.5 ;
      RECT  153.6 194.7 154.4 195.5 ;
      RECT  157.6 194.7 158.4 195.5 ;
      RECT  155.6 194.7 156.4 195.5 ;
      RECT  153.6 187.7 154.4 188.5 ;
      RECT  157.6 187.7 158.4 188.5 ;
      RECT  154.6 189.2 155.4 190.0 ;
      RECT  156.6 192.0 157.4 192.8 ;
      RECT  159.1 193.4 159.7 194.0 ;
      RECT  152.4 196.5 161.0 197.1 ;
      RECT  152.4 186.1 161.0 186.7 ;
      RECT  164.2 194.7 165.0 195.5 ;
      RECT  162.2 194.7 163.0 195.5 ;
      RECT  164.2 187.3 165.0 188.1 ;
      RECT  162.2 187.3 163.0 188.1 ;
      RECT  162.6 191.0 163.4 191.8 ;
      RECT  164.6 191.1 165.2 191.7 ;
      RECT  161.0 196.5 167.6 197.1 ;
      RECT  161.0 186.1 167.6 186.7 ;
      RECT  154.6 189.2 155.4 190.0 ;
      RECT  156.6 192.0 157.4 192.8 ;
      RECT  164.6 191.1 165.2 191.7 ;
      RECT  152.4 196.5 167.6 197.1 ;
      RECT  152.4 186.1 167.6 186.7 ;
      RECT  155.6 198.9 156.4 198.1 ;
      RECT  153.6 198.9 154.4 198.1 ;
      RECT  157.6 198.9 158.4 198.1 ;
      RECT  155.6 198.9 156.4 198.1 ;
      RECT  153.6 205.9 154.4 205.1 ;
      RECT  157.6 205.9 158.4 205.1 ;
      RECT  154.6 204.4 155.4 203.6 ;
      RECT  156.6 201.6 157.4 200.8 ;
      RECT  159.1 200.2 159.7 199.6 ;
      RECT  152.4 197.1 161.0 196.5 ;
      RECT  152.4 207.5 161.0 206.9 ;
      RECT  164.2 198.9 165.0 198.1 ;
      RECT  162.2 198.9 163.0 198.1 ;
      RECT  164.2 206.3 165.0 205.5 ;
      RECT  162.2 206.3 163.0 205.5 ;
      RECT  162.6 202.6 163.4 201.8 ;
      RECT  164.6 202.5 165.2 201.9 ;
      RECT  161.0 197.1 167.6 196.5 ;
      RECT  161.0 207.5 167.6 206.9 ;
      RECT  154.6 204.4 155.4 203.6 ;
      RECT  156.6 201.6 157.4 200.8 ;
      RECT  164.6 202.5 165.2 201.9 ;
      RECT  152.4 197.1 167.6 196.5 ;
      RECT  152.4 207.5 167.6 206.9 ;
      RECT  155.6 215.5 156.4 216.3 ;
      RECT  153.6 215.5 154.4 216.3 ;
      RECT  157.6 215.5 158.4 216.3 ;
      RECT  155.6 215.5 156.4 216.3 ;
      RECT  153.6 208.5 154.4 209.3 ;
      RECT  157.6 208.5 158.4 209.3 ;
      RECT  154.6 210.0 155.4 210.8 ;
      RECT  156.6 212.8 157.4 213.6 ;
      RECT  159.1 214.2 159.7 214.8 ;
      RECT  152.4 217.3 161.0 217.9 ;
      RECT  152.4 206.9 161.0 207.5 ;
      RECT  164.2 215.5 165.0 216.3 ;
      RECT  162.2 215.5 163.0 216.3 ;
      RECT  164.2 208.1 165.0 208.9 ;
      RECT  162.2 208.1 163.0 208.9 ;
      RECT  162.6 211.8 163.4 212.6 ;
      RECT  164.6 211.9 165.2 212.5 ;
      RECT  161.0 217.3 167.6 217.9 ;
      RECT  161.0 206.9 167.6 207.5 ;
      RECT  154.6 210.0 155.4 210.8 ;
      RECT  156.6 212.8 157.4 213.6 ;
      RECT  164.6 211.9 165.2 212.5 ;
      RECT  152.4 217.3 167.6 217.9 ;
      RECT  152.4 206.9 167.6 207.5 ;
      RECT  155.6 219.7 156.4 218.9 ;
      RECT  153.6 219.7 154.4 218.9 ;
      RECT  157.6 219.7 158.4 218.9 ;
      RECT  155.6 219.7 156.4 218.9 ;
      RECT  153.6 226.7 154.4 225.9 ;
      RECT  157.6 226.7 158.4 225.9 ;
      RECT  154.6 225.2 155.4 224.4 ;
      RECT  156.6 222.4 157.4 221.6 ;
      RECT  159.1 221.0 159.7 220.4 ;
      RECT  152.4 217.9 161.0 217.3 ;
      RECT  152.4 228.3 161.0 227.7 ;
      RECT  164.2 219.7 165.0 218.9 ;
      RECT  162.2 219.7 163.0 218.9 ;
      RECT  164.2 227.1 165.0 226.3 ;
      RECT  162.2 227.1 163.0 226.3 ;
      RECT  162.6 223.4 163.4 222.6 ;
      RECT  164.6 223.3 165.2 222.7 ;
      RECT  161.0 217.9 167.6 217.3 ;
      RECT  161.0 228.3 167.6 227.7 ;
      RECT  154.6 225.2 155.4 224.4 ;
      RECT  156.6 222.4 157.4 221.6 ;
      RECT  164.6 223.3 165.2 222.7 ;
      RECT  152.4 217.9 167.6 217.3 ;
      RECT  152.4 228.3 167.6 227.7 ;
      RECT  155.6 236.3 156.4 237.1 ;
      RECT  153.6 236.3 154.4 237.1 ;
      RECT  157.6 236.3 158.4 237.1 ;
      RECT  155.6 236.3 156.4 237.1 ;
      RECT  153.6 229.3 154.4 230.1 ;
      RECT  157.6 229.3 158.4 230.1 ;
      RECT  154.6 230.8 155.4 231.6 ;
      RECT  156.6 233.6 157.4 234.4 ;
      RECT  159.1 235.0 159.7 235.6 ;
      RECT  152.4 238.1 161.0 238.7 ;
      RECT  152.4 227.7 161.0 228.3 ;
      RECT  164.2 236.3 165.0 237.1 ;
      RECT  162.2 236.3 163.0 237.1 ;
      RECT  164.2 228.9 165.0 229.7 ;
      RECT  162.2 228.9 163.0 229.7 ;
      RECT  162.6 232.6 163.4 233.4 ;
      RECT  164.6 232.7 165.2 233.3 ;
      RECT  161.0 238.1 167.6 238.7 ;
      RECT  161.0 227.7 167.6 228.3 ;
      RECT  154.6 230.8 155.4 231.6 ;
      RECT  156.6 233.6 157.4 234.4 ;
      RECT  164.6 232.7 165.2 233.3 ;
      RECT  152.4 238.1 167.6 238.7 ;
      RECT  152.4 227.7 167.6 228.3 ;
      RECT  155.6 240.5 156.4 239.7 ;
      RECT  153.6 240.5 154.4 239.7 ;
      RECT  157.6 240.5 158.4 239.7 ;
      RECT  155.6 240.5 156.4 239.7 ;
      RECT  153.6 247.5 154.4 246.7 ;
      RECT  157.6 247.5 158.4 246.7 ;
      RECT  154.6 246.0 155.4 245.2 ;
      RECT  156.6 243.2 157.4 242.4 ;
      RECT  159.1 241.8 159.7 241.2 ;
      RECT  152.4 238.7 161.0 238.1 ;
      RECT  152.4 249.1 161.0 248.5 ;
      RECT  164.2 240.5 165.0 239.7 ;
      RECT  162.2 240.5 163.0 239.7 ;
      RECT  164.2 247.9 165.0 247.1 ;
      RECT  162.2 247.9 163.0 247.1 ;
      RECT  162.6 244.2 163.4 243.4 ;
      RECT  164.6 244.1 165.2 243.5 ;
      RECT  161.0 238.7 167.6 238.1 ;
      RECT  161.0 249.1 167.6 248.5 ;
      RECT  154.6 246.0 155.4 245.2 ;
      RECT  156.6 243.2 157.4 242.4 ;
      RECT  164.6 244.1 165.2 243.5 ;
      RECT  152.4 238.7 167.6 238.1 ;
      RECT  152.4 249.1 167.6 248.5 ;
      RECT  155.6 257.1 156.4 257.9 ;
      RECT  153.6 257.1 154.4 257.9 ;
      RECT  157.6 257.1 158.4 257.9 ;
      RECT  155.6 257.1 156.4 257.9 ;
      RECT  153.6 250.1 154.4 250.9 ;
      RECT  157.6 250.1 158.4 250.9 ;
      RECT  154.6 251.6 155.4 252.4 ;
      RECT  156.6 254.4 157.4 255.2 ;
      RECT  159.1 255.8 159.7 256.4 ;
      RECT  152.4 258.9 161.0 259.5 ;
      RECT  152.4 248.5 161.0 249.1 ;
      RECT  164.2 257.1 165.0 257.9 ;
      RECT  162.2 257.1 163.0 257.9 ;
      RECT  164.2 249.7 165.0 250.5 ;
      RECT  162.2 249.7 163.0 250.5 ;
      RECT  162.6 253.4 163.4 254.2 ;
      RECT  164.6 253.5 165.2 254.1 ;
      RECT  161.0 258.9 167.6 259.5 ;
      RECT  161.0 248.5 167.6 249.1 ;
      RECT  154.6 251.6 155.4 252.4 ;
      RECT  156.6 254.4 157.4 255.2 ;
      RECT  164.6 253.5 165.2 254.1 ;
      RECT  152.4 258.9 167.6 259.5 ;
      RECT  152.4 248.5 167.6 249.1 ;
      RECT  155.6 261.3 156.4 260.5 ;
      RECT  153.6 261.3 154.4 260.5 ;
      RECT  157.6 261.3 158.4 260.5 ;
      RECT  155.6 261.3 156.4 260.5 ;
      RECT  153.6 268.3 154.4 267.5 ;
      RECT  157.6 268.3 158.4 267.5 ;
      RECT  154.6 266.8 155.4 266.0 ;
      RECT  156.6 264.0 157.4 263.2 ;
      RECT  159.1 262.6 159.7 262.0 ;
      RECT  152.4 259.5 161.0 258.9 ;
      RECT  152.4 269.9 161.0 269.3 ;
      RECT  164.2 261.3 165.0 260.5 ;
      RECT  162.2 261.3 163.0 260.5 ;
      RECT  164.2 268.7 165.0 267.9 ;
      RECT  162.2 268.7 163.0 267.9 ;
      RECT  162.6 265.0 163.4 264.2 ;
      RECT  164.6 264.9 165.2 264.3 ;
      RECT  161.0 259.5 167.6 258.9 ;
      RECT  161.0 269.9 167.6 269.3 ;
      RECT  154.6 266.8 155.4 266.0 ;
      RECT  156.6 264.0 157.4 263.2 ;
      RECT  164.6 264.9 165.2 264.3 ;
      RECT  152.4 259.5 167.6 258.9 ;
      RECT  152.4 269.9 167.6 269.3 ;
      RECT  155.6 277.9 156.4 278.7 ;
      RECT  153.6 277.9 154.4 278.7 ;
      RECT  157.6 277.9 158.4 278.7 ;
      RECT  155.6 277.9 156.4 278.7 ;
      RECT  153.6 270.9 154.4 271.7 ;
      RECT  157.6 270.9 158.4 271.7 ;
      RECT  154.6 272.4 155.4 273.2 ;
      RECT  156.6 275.2 157.4 276.0 ;
      RECT  159.1 276.6 159.7 277.2 ;
      RECT  152.4 279.7 161.0 280.3 ;
      RECT  152.4 269.3 161.0 269.9 ;
      RECT  164.2 277.9 165.0 278.7 ;
      RECT  162.2 277.9 163.0 278.7 ;
      RECT  164.2 270.5 165.0 271.3 ;
      RECT  162.2 270.5 163.0 271.3 ;
      RECT  162.6 274.2 163.4 275.0 ;
      RECT  164.6 274.3 165.2 274.9 ;
      RECT  161.0 279.7 167.6 280.3 ;
      RECT  161.0 269.3 167.6 269.9 ;
      RECT  154.6 272.4 155.4 273.2 ;
      RECT  156.6 275.2 157.4 276.0 ;
      RECT  164.6 274.3 165.2 274.9 ;
      RECT  152.4 279.7 167.6 280.3 ;
      RECT  152.4 269.3 167.6 269.9 ;
      RECT  155.6 282.1 156.4 281.3 ;
      RECT  153.6 282.1 154.4 281.3 ;
      RECT  157.6 282.1 158.4 281.3 ;
      RECT  155.6 282.1 156.4 281.3 ;
      RECT  153.6 289.1 154.4 288.3 ;
      RECT  157.6 289.1 158.4 288.3 ;
      RECT  154.6 287.6 155.4 286.8 ;
      RECT  156.6 284.8 157.4 284.0 ;
      RECT  159.1 283.4 159.7 282.8 ;
      RECT  152.4 280.3 161.0 279.7 ;
      RECT  152.4 290.7 161.0 290.1 ;
      RECT  164.2 282.1 165.0 281.3 ;
      RECT  162.2 282.1 163.0 281.3 ;
      RECT  164.2 289.5 165.0 288.7 ;
      RECT  162.2 289.5 163.0 288.7 ;
      RECT  162.6 285.8 163.4 285.0 ;
      RECT  164.6 285.7 165.2 285.1 ;
      RECT  161.0 280.3 167.6 279.7 ;
      RECT  161.0 290.7 167.6 290.1 ;
      RECT  154.6 287.6 155.4 286.8 ;
      RECT  156.6 284.8 157.4 284.0 ;
      RECT  164.6 285.7 165.2 285.1 ;
      RECT  152.4 280.3 167.6 279.7 ;
      RECT  152.4 290.7 167.6 290.1 ;
      RECT  155.6 298.7 156.4 299.5 ;
      RECT  153.6 298.7 154.4 299.5 ;
      RECT  157.6 298.7 158.4 299.5 ;
      RECT  155.6 298.7 156.4 299.5 ;
      RECT  153.6 291.7 154.4 292.5 ;
      RECT  157.6 291.7 158.4 292.5 ;
      RECT  154.6 293.2 155.4 294.0 ;
      RECT  156.6 296.0 157.4 296.8 ;
      RECT  159.1 297.4 159.7 298.0 ;
      RECT  152.4 300.5 161.0 301.1 ;
      RECT  152.4 290.1 161.0 290.7 ;
      RECT  164.2 298.7 165.0 299.5 ;
      RECT  162.2 298.7 163.0 299.5 ;
      RECT  164.2 291.3 165.0 292.1 ;
      RECT  162.2 291.3 163.0 292.1 ;
      RECT  162.6 295.0 163.4 295.8 ;
      RECT  164.6 295.1 165.2 295.7 ;
      RECT  161.0 300.5 167.6 301.1 ;
      RECT  161.0 290.1 167.6 290.7 ;
      RECT  154.6 293.2 155.4 294.0 ;
      RECT  156.6 296.0 157.4 296.8 ;
      RECT  164.6 295.1 165.2 295.7 ;
      RECT  152.4 300.5 167.6 301.1 ;
      RECT  152.4 290.1 167.6 290.7 ;
      RECT  155.6 302.9 156.4 302.1 ;
      RECT  153.6 302.9 154.4 302.1 ;
      RECT  157.6 302.9 158.4 302.1 ;
      RECT  155.6 302.9 156.4 302.1 ;
      RECT  153.6 309.9 154.4 309.1 ;
      RECT  157.6 309.9 158.4 309.1 ;
      RECT  154.6 308.4 155.4 307.6 ;
      RECT  156.6 305.6 157.4 304.8 ;
      RECT  159.1 304.2 159.7 303.6 ;
      RECT  152.4 301.1 161.0 300.5 ;
      RECT  152.4 311.5 161.0 310.9 ;
      RECT  164.2 302.9 165.0 302.1 ;
      RECT  162.2 302.9 163.0 302.1 ;
      RECT  164.2 310.3 165.0 309.5 ;
      RECT  162.2 310.3 163.0 309.5 ;
      RECT  162.6 306.6 163.4 305.8 ;
      RECT  164.6 306.5 165.2 305.9 ;
      RECT  161.0 301.1 167.6 300.5 ;
      RECT  161.0 311.5 167.6 310.9 ;
      RECT  154.6 308.4 155.4 307.6 ;
      RECT  156.6 305.6 157.4 304.8 ;
      RECT  164.6 306.5 165.2 305.9 ;
      RECT  152.4 301.1 167.6 300.5 ;
      RECT  152.4 311.5 167.6 310.9 ;
      RECT  155.6 319.5 156.4 320.3 ;
      RECT  153.6 319.5 154.4 320.3 ;
      RECT  157.6 319.5 158.4 320.3 ;
      RECT  155.6 319.5 156.4 320.3 ;
      RECT  153.6 312.5 154.4 313.3 ;
      RECT  157.6 312.5 158.4 313.3 ;
      RECT  154.6 314.0 155.4 314.8 ;
      RECT  156.6 316.8 157.4 317.6 ;
      RECT  159.1 318.2 159.7 318.8 ;
      RECT  152.4 321.3 161.0 321.9 ;
      RECT  152.4 310.9 161.0 311.5 ;
      RECT  164.2 319.5 165.0 320.3 ;
      RECT  162.2 319.5 163.0 320.3 ;
      RECT  164.2 312.1 165.0 312.9 ;
      RECT  162.2 312.1 163.0 312.9 ;
      RECT  162.6 315.8 163.4 316.6 ;
      RECT  164.6 315.9 165.2 316.5 ;
      RECT  161.0 321.3 167.6 321.9 ;
      RECT  161.0 310.9 167.6 311.5 ;
      RECT  154.6 314.0 155.4 314.8 ;
      RECT  156.6 316.8 157.4 317.6 ;
      RECT  164.6 315.9 165.2 316.5 ;
      RECT  152.4 321.3 167.6 321.9 ;
      RECT  152.4 310.9 167.6 311.5 ;
      RECT  155.6 323.7 156.4 322.9 ;
      RECT  153.6 323.7 154.4 322.9 ;
      RECT  157.6 323.7 158.4 322.9 ;
      RECT  155.6 323.7 156.4 322.9 ;
      RECT  153.6 330.7 154.4 329.9 ;
      RECT  157.6 330.7 158.4 329.9 ;
      RECT  154.6 329.2 155.4 328.4 ;
      RECT  156.6 326.4 157.4 325.6 ;
      RECT  159.1 325.0 159.7 324.4 ;
      RECT  152.4 321.9 161.0 321.3 ;
      RECT  152.4 332.3 161.0 331.7 ;
      RECT  164.2 323.7 165.0 322.9 ;
      RECT  162.2 323.7 163.0 322.9 ;
      RECT  164.2 331.1 165.0 330.3 ;
      RECT  162.2 331.1 163.0 330.3 ;
      RECT  162.6 327.4 163.4 326.6 ;
      RECT  164.6 327.3 165.2 326.7 ;
      RECT  161.0 321.9 167.6 321.3 ;
      RECT  161.0 332.3 167.6 331.7 ;
      RECT  154.6 329.2 155.4 328.4 ;
      RECT  156.6 326.4 157.4 325.6 ;
      RECT  164.6 327.3 165.2 326.7 ;
      RECT  152.4 321.9 167.6 321.3 ;
      RECT  152.4 332.3 167.6 331.7 ;
      RECT  155.6 340.3 156.4 341.1 ;
      RECT  153.6 340.3 154.4 341.1 ;
      RECT  157.6 340.3 158.4 341.1 ;
      RECT  155.6 340.3 156.4 341.1 ;
      RECT  153.6 333.3 154.4 334.1 ;
      RECT  157.6 333.3 158.4 334.1 ;
      RECT  154.6 334.8 155.4 335.6 ;
      RECT  156.6 337.6 157.4 338.4 ;
      RECT  159.1 339.0 159.7 339.6 ;
      RECT  152.4 342.1 161.0 342.7 ;
      RECT  152.4 331.7 161.0 332.3 ;
      RECT  164.2 340.3 165.0 341.1 ;
      RECT  162.2 340.3 163.0 341.1 ;
      RECT  164.2 332.9 165.0 333.7 ;
      RECT  162.2 332.9 163.0 333.7 ;
      RECT  162.6 336.6 163.4 337.4 ;
      RECT  164.6 336.7 165.2 337.3 ;
      RECT  161.0 342.1 167.6 342.7 ;
      RECT  161.0 331.7 167.6 332.3 ;
      RECT  154.6 334.8 155.4 335.6 ;
      RECT  156.6 337.6 157.4 338.4 ;
      RECT  164.6 336.7 165.2 337.3 ;
      RECT  152.4 342.1 167.6 342.7 ;
      RECT  152.4 331.7 167.6 332.3 ;
      RECT  155.6 344.5 156.4 343.7 ;
      RECT  153.6 344.5 154.4 343.7 ;
      RECT  157.6 344.5 158.4 343.7 ;
      RECT  155.6 344.5 156.4 343.7 ;
      RECT  153.6 351.5 154.4 350.7 ;
      RECT  157.6 351.5 158.4 350.7 ;
      RECT  154.6 350.0 155.4 349.2 ;
      RECT  156.6 347.2 157.4 346.4 ;
      RECT  159.1 345.8 159.7 345.2 ;
      RECT  152.4 342.7 161.0 342.1 ;
      RECT  152.4 353.1 161.0 352.5 ;
      RECT  164.2 344.5 165.0 343.7 ;
      RECT  162.2 344.5 163.0 343.7 ;
      RECT  164.2 351.9 165.0 351.1 ;
      RECT  162.2 351.9 163.0 351.1 ;
      RECT  162.6 348.2 163.4 347.4 ;
      RECT  164.6 348.1 165.2 347.5 ;
      RECT  161.0 342.7 167.6 342.1 ;
      RECT  161.0 353.1 167.6 352.5 ;
      RECT  154.6 350.0 155.4 349.2 ;
      RECT  156.6 347.2 157.4 346.4 ;
      RECT  164.6 348.1 165.2 347.5 ;
      RECT  152.4 342.7 167.6 342.1 ;
      RECT  152.4 353.1 167.6 352.5 ;
      RECT  154.6 189.2 155.4 190.0 ;
      RECT  154.6 203.6 155.4 204.4 ;
      RECT  154.6 210.0 155.4 210.8 ;
      RECT  154.6 224.4 155.4 225.2 ;
      RECT  154.6 230.8 155.4 231.6 ;
      RECT  154.6 245.2 155.4 246.0 ;
      RECT  154.6 251.6 155.4 252.4 ;
      RECT  154.6 266.0 155.4 266.8 ;
      RECT  154.6 272.4 155.4 273.2 ;
      RECT  154.6 286.8 155.4 287.6 ;
      RECT  154.6 293.2 155.4 294.0 ;
      RECT  154.6 307.6 155.4 308.4 ;
      RECT  154.6 314.0 155.4 314.8 ;
      RECT  154.6 328.4 155.4 329.2 ;
      RECT  154.6 334.8 155.4 335.6 ;
      RECT  154.6 349.2 155.4 350.0 ;
      RECT  164.6 191.1 165.2 191.7 ;
      RECT  164.6 201.9 165.2 202.5 ;
      RECT  164.6 211.9 165.2 212.5 ;
      RECT  164.6 222.7 165.2 223.3 ;
      RECT  164.6 232.7 165.2 233.3 ;
      RECT  164.6 243.5 165.2 244.1 ;
      RECT  164.6 253.5 165.2 254.1 ;
      RECT  164.6 264.3 165.2 264.9 ;
      RECT  164.6 274.3 165.2 274.9 ;
      RECT  164.6 285.1 165.2 285.7 ;
      RECT  164.6 295.1 165.2 295.7 ;
      RECT  164.6 305.9 165.2 306.5 ;
      RECT  164.6 315.9 165.2 316.5 ;
      RECT  164.6 326.7 165.2 327.3 ;
      RECT  164.6 336.7 165.2 337.3 ;
      RECT  164.6 347.5 165.2 348.1 ;
      RECT  158.8 178.1 159.6 177.3 ;
      RECT  156.8 178.1 157.6 177.3 ;
      RECT  158.8 185.5 159.6 184.7 ;
      RECT  156.8 185.5 157.6 184.7 ;
      RECT  157.2 181.8 158.0 181.0 ;
      RECT  159.2 181.7 159.8 181.1 ;
      RECT  155.6 176.3 162.2 175.7 ;
      RECT  155.6 186.7 162.2 186.1 ;
      RECT  165.4 178.1 166.2 177.3 ;
      RECT  163.4 178.1 164.2 177.3 ;
      RECT  165.4 185.5 166.2 184.7 ;
      RECT  163.4 185.5 164.2 184.7 ;
      RECT  163.8 181.8 164.6 181.0 ;
      RECT  165.8 181.7 166.4 181.1 ;
      RECT  162.2 176.3 167.4 175.7 ;
      RECT  162.2 186.7 167.4 186.1 ;
      RECT  157.2 181.8 158.0 181.0 ;
      RECT  165.8 181.7 166.4 181.1 ;
      RECT  155.6 176.3 167.4 175.7 ;
      RECT  155.6 186.7 167.4 186.1 ;
      RECT  164.6 191.1 165.2 191.7 ;
      RECT  164.6 201.9 165.2 202.5 ;
      RECT  164.6 211.9 165.2 212.5 ;
      RECT  164.6 222.7 165.2 223.3 ;
      RECT  164.6 232.7 165.2 233.3 ;
      RECT  164.6 243.5 165.2 244.1 ;
      RECT  164.6 253.5 165.2 254.1 ;
      RECT  164.6 264.3 165.2 264.9 ;
      RECT  164.6 274.3 165.2 274.9 ;
      RECT  164.6 285.1 165.2 285.7 ;
      RECT  164.6 295.1 165.2 295.7 ;
      RECT  164.6 305.9 165.2 306.5 ;
      RECT  164.6 315.9 165.2 316.5 ;
      RECT  164.6 326.7 165.2 327.3 ;
      RECT  164.6 336.7 165.2 337.3 ;
      RECT  164.6 347.5 165.2 348.1 ;
      RECT  165.8 181.1 166.4 181.7 ;
      RECT  3.6 13.0 13.4 13.2 ;
      RECT  17.8 12.4 22.0 13.0 ;
      RECT  21.2 4.0 22.0 8.4 ;
      RECT  10.2 16.4 13.8 17.0 ;
      RECT  21.2 9.0 22.0 12.4 ;
      RECT  10.2 7.2 11.0 7.4 ;
      RECT  12.8 14.8 15.0 15.4 ;
      RECT  3.6 4.0 4.4 8.8 ;
      RECT  14.2 9.4 15.0 9.6 ;
      RECT  10.2 16.2 11.0 16.4 ;
      RECT  14.2 14.6 15.0 14.8 ;
      RECT  6.8 14.8 7.6 15.0 ;
      RECT  14.8 13.4 17.2 14.0 ;
      RECT  7.4 10.2 8.2 10.4 ;
      RECT  21.2 13.0 22.0 21.6 ;
      RECT  18.2 8.2 19.0 8.4 ;
      RECT  16.4 11.0 20.2 11.6 ;
      RECT  8.6 7.4 9.2 9.6 ;
      RECT  10.6 3.4 11.6 6.0 ;
      RECT  19.6 3.4 20.4 7.8 ;
      RECT  11.4 14.8 12.2 15.0 ;
      RECT  19.4 11.6 20.2 11.8 ;
      RECT  12.4 17.6 13.2 21.6 ;
      RECT  6.8 16.8 7.6 17.6 ;
      RECT  16.4 16.8 17.2 17.6 ;
      RECT  8.6 13.2 13.4 13.6 ;
      RECT  3.6 12.8 9.4 13.0 ;
      RECT  5.8 11.4 10.8 12.0 ;
      RECT  13.0 16.2 13.8 16.4 ;
      RECT  6.8 17.6 8.8 18.2 ;
      RECT  5.2 3.4 6.0 8.0 ;
      RECT  10.2 6.6 13.0 7.2 ;
      RECT  22.8 3.4 23.6 4.8 ;
      RECT  3.6 13.2 4.4 21.6 ;
      RECT  5.2 13.8 6.0 22.2 ;
      RECT  16.6 14.0 17.2 15.0 ;
      RECT  16.4 5.4 17.8 6.0 ;
      RECT  10.8 17.6 11.6 22.2 ;
      RECT  14.0 17.6 14.8 22.2 ;
      RECT  16.6 15.0 18.0 15.8 ;
      RECT  14.8 10.2 15.4 13.4 ;
      RECT  4.4 9.4 6.0 9.6 ;
      RECT  6.8 5.4 8.8 6.0 ;
      RECT  8.0 4.0 8.8 5.4 ;
      RECT  16.6 17.6 17.8 21.6 ;
      RECT  8.4 6.6 9.2 7.4 ;
      RECT  12.8 13.6 13.4 14.8 ;
      RECT  10.0 12.0 10.8 12.2 ;
      RECT  16.4 10.8 17.2 11.0 ;
      RECT  12.4 17.0 13.0 17.6 ;
      RECT  6.8 14.2 12.2 14.8 ;
      RECT  12.4 4.0 13.2 6.0 ;
      RECT  2.4 22.2 24.2 23.4 ;
      RECT  8.0 18.2 8.8 21.6 ;
      RECT  19.6 13.6 20.4 22.2 ;
      RECT  3.6 12.6 9.2 12.8 ;
      RECT  5.8 11.2 6.6 11.4 ;
      RECT  14.0 3.4 14.8 6.0 ;
      RECT  16.6 4.0 17.8 5.4 ;
      RECT  2.4 2.2 24.2 3.4 ;
      RECT  22.8 20.6 23.6 22.2 ;
      RECT  4.4 9.6 15.4 10.2 ;
      RECT  18.2 8.4 22.0 9.0 ;
      RECT  6.8 6.0 7.6 6.8 ;
      RECT  12.4 6.0 13.0 6.6 ;
      RECT  16.4 6.0 17.2 6.8 ;
      RECT  17.8 12.2 18.6 12.4 ;
      RECT  29.8 19.9 30.6 20.7 ;
      RECT  27.8 19.9 28.6 20.7 ;
      RECT  29.8 4.1 30.6 4.9 ;
      RECT  27.8 4.1 28.6 4.9 ;
      RECT  28.2 12.0 29.0 12.8 ;
      RECT  30.2 12.1 30.8 12.7 ;
      RECT  26.6 22.5 33.2 23.1 ;
      RECT  26.6 2.5 33.2 3.1 ;
      RECT  36.4 18.3 37.2 19.1 ;
      RECT  34.4 18.3 35.2 19.1 ;
      RECT  36.4 4.9 37.2 5.7 ;
      RECT  34.4 4.9 35.2 5.7 ;
      RECT  34.8 11.6 35.6 12.4 ;
      RECT  36.8 11.7 37.4 12.3 ;
      RECT  33.2 22.5 39.8 23.1 ;
      RECT  33.2 2.5 39.8 3.1 ;
      RECT  2.4 22.2 39.8 23.4 ;
      RECT  2.4 2.2 39.8 3.4 ;
      RECT  3.6 32.6 13.4 32.4 ;
      RECT  17.8 33.2 22.0 32.6 ;
      RECT  21.2 41.6 22.0 37.2 ;
      RECT  10.2 29.2 13.8 28.6 ;
      RECT  21.2 36.6 22.0 33.2 ;
      RECT  10.2 38.4 11.0 38.2 ;
      RECT  12.8 30.8 15.0 30.2 ;
      RECT  3.6 41.6 4.4 36.8 ;
      RECT  14.2 36.2 15.0 36.0 ;
      RECT  10.2 29.4 11.0 29.2 ;
      RECT  14.2 31.0 15.0 30.8 ;
      RECT  6.8 30.8 7.6 30.6 ;
      RECT  14.8 32.2 17.2 31.6 ;
      RECT  7.4 35.4 8.2 35.2 ;
      RECT  21.2 32.6 22.0 24.0 ;
      RECT  18.2 37.4 19.0 37.2 ;
      RECT  16.4 34.6 20.2 34.0 ;
      RECT  8.6 38.2 9.2 36.0 ;
      RECT  10.6 42.2 11.6 39.6 ;
      RECT  19.6 42.2 20.4 37.8 ;
      RECT  11.4 30.8 12.2 30.6 ;
      RECT  19.4 34.0 20.2 33.8 ;
      RECT  12.4 28.0 13.2 24.0 ;
      RECT  6.8 28.8 7.6 28.0 ;
      RECT  16.4 28.8 17.2 28.0 ;
      RECT  8.6 32.4 13.4 32.0 ;
      RECT  3.6 32.8 9.4 32.6 ;
      RECT  5.8 34.2 10.8 33.6 ;
      RECT  13.0 29.4 13.8 29.2 ;
      RECT  6.8 28.0 8.8 27.4 ;
      RECT  5.2 42.2 6.0 37.6 ;
      RECT  10.2 39.0 13.0 38.4 ;
      RECT  22.8 42.2 23.6 40.8 ;
      RECT  3.6 32.4 4.4 24.0 ;
      RECT  5.2 31.8 6.0 23.4 ;
      RECT  16.6 31.6 17.2 30.6 ;
      RECT  16.4 40.2 17.8 39.6 ;
      RECT  10.8 28.0 11.6 23.4 ;
      RECT  14.0 28.0 14.8 23.4 ;
      RECT  16.6 30.6 18.0 29.8 ;
      RECT  14.8 35.4 15.4 32.2 ;
      RECT  4.4 36.2 6.0 36.0 ;
      RECT  6.8 40.2 8.8 39.6 ;
      RECT  8.0 41.6 8.8 40.2 ;
      RECT  16.6 28.0 17.8 24.0 ;
      RECT  8.4 39.0 9.2 38.2 ;
      RECT  12.8 32.0 13.4 30.8 ;
      RECT  10.0 33.6 10.8 33.4 ;
      RECT  16.4 34.8 17.2 34.6 ;
      RECT  12.4 28.6 13.0 28.0 ;
      RECT  6.8 31.4 12.2 30.8 ;
      RECT  12.4 41.6 13.2 39.6 ;
      RECT  2.4 23.4 24.2 22.2 ;
      RECT  8.0 27.4 8.8 24.0 ;
      RECT  19.6 32.0 20.4 23.4 ;
      RECT  3.6 33.0 9.2 32.8 ;
      RECT  5.8 34.4 6.6 34.2 ;
      RECT  14.0 42.2 14.8 39.6 ;
      RECT  16.6 41.6 17.8 40.2 ;
      RECT  2.4 43.4 24.2 42.2 ;
      RECT  22.8 25.0 23.6 23.4 ;
      RECT  4.4 36.0 15.4 35.4 ;
      RECT  18.2 37.2 22.0 36.6 ;
      RECT  6.8 39.6 7.6 38.8 ;
      RECT  12.4 39.6 13.0 39.0 ;
      RECT  16.4 39.6 17.2 38.8 ;
      RECT  17.8 33.4 18.6 33.2 ;
      RECT  29.8 25.7 30.6 24.9 ;
      RECT  27.8 25.7 28.6 24.9 ;
      RECT  29.8 41.5 30.6 40.7 ;
      RECT  27.8 41.5 28.6 40.7 ;
      RECT  28.2 33.6 29.0 32.8 ;
      RECT  30.2 33.5 30.8 32.9 ;
      RECT  26.6 23.1 33.2 22.5 ;
      RECT  26.6 43.1 33.2 42.5 ;
      RECT  36.4 27.3 37.2 26.5 ;
      RECT  34.4 27.3 35.2 26.5 ;
      RECT  36.4 40.7 37.2 39.9 ;
      RECT  34.4 40.7 35.2 39.9 ;
      RECT  34.8 34.0 35.6 33.2 ;
      RECT  36.8 33.9 37.4 33.3 ;
      RECT  33.2 23.1 39.8 22.5 ;
      RECT  33.2 43.1 39.8 42.5 ;
      RECT  2.4 23.4 39.8 22.2 ;
      RECT  2.4 43.4 39.8 42.2 ;
      RECT  55.6 20.7 56.4 21.5 ;
      RECT  53.6 20.7 54.4 21.5 ;
      RECT  55.6 3.7 56.4 4.5 ;
      RECT  53.6 3.7 54.4 4.5 ;
      RECT  54.0 12.2 54.8 13.0 ;
      RECT  56.0 12.3 56.6 12.9 ;
      RECT  52.4 22.5 59.0 23.1 ;
      RECT  52.4 2.5 59.0 3.1 ;
      RECT  62.2 19.9 63.0 20.7 ;
      RECT  60.2 19.9 61.0 20.7 ;
      RECT  62.2 4.1 63.0 4.9 ;
      RECT  60.2 4.1 61.0 4.9 ;
      RECT  60.6 12.0 61.4 12.8 ;
      RECT  62.6 12.1 63.2 12.7 ;
      RECT  59.0 22.5 64.2 23.1 ;
      RECT  59.0 2.5 64.2 3.1 ;
      RECT  67.4 17.5 68.2 18.3 ;
      RECT  65.4 17.5 66.2 18.3 ;
      RECT  67.4 5.3 68.2 6.1 ;
      RECT  65.4 5.3 66.2 6.1 ;
      RECT  65.8 11.4 66.6 12.2 ;
      RECT  67.8 11.5 68.4 12.1 ;
      RECT  64.2 22.5 69.4 23.1 ;
      RECT  64.2 2.5 69.4 3.1 ;
      RECT  72.5 16.3 76.5 16.9 ;
      RECT  74.0 17.5 74.8 18.3 ;
      RECT  70.6 17.5 71.4 18.3 ;
      RECT  72.5 6.7 76.5 7.3 ;
      RECT  70.6 5.3 71.4 6.1 ;
      RECT  74.0 5.3 74.8 6.1 ;
      RECT  71.0 11.4 71.8 12.2 ;
      RECT  74.5 11.5 75.1 12.1 ;
      RECT  69.4 22.5 78.0 23.1 ;
      RECT  69.4 2.5 78.0 3.1 ;
      RECT  54.0 12.2 54.8 13.0 ;
      RECT  74.5 11.5 75.1 12.1 ;
      RECT  52.4 22.5 78.0 23.1 ;
      RECT  52.4 2.5 78.0 3.1 ;
      RECT  55.6 24.9 56.4 24.1 ;
      RECT  53.6 24.9 54.4 24.1 ;
      RECT  55.6 41.9 56.4 41.1 ;
      RECT  53.6 41.9 54.4 41.1 ;
      RECT  54.0 33.4 54.8 32.6 ;
      RECT  56.0 33.3 56.6 32.7 ;
      RECT  52.4 23.1 59.0 22.5 ;
      RECT  52.4 43.1 59.0 42.5 ;
      RECT  62.2 24.9 63.0 24.1 ;
      RECT  60.2 24.9 61.0 24.1 ;
      RECT  64.2 24.9 65.0 24.1 ;
      RECT  62.2 24.9 63.0 24.1 ;
      RECT  60.2 41.5 61.0 40.7 ;
      RECT  64.2 41.5 65.0 40.7 ;
      RECT  61.2 40.0 62.0 39.2 ;
      RECT  63.2 37.2 64.0 36.4 ;
      RECT  65.7 26.2 66.3 25.6 ;
      RECT  59.0 23.1 66.6 22.5 ;
      RECT  59.0 43.1 66.6 42.5 ;
      RECT  69.7 28.5 73.7 27.9 ;
      RECT  67.8 27.3 68.6 26.5 ;
      RECT  71.2 27.3 72.0 26.5 ;
      RECT  69.7 39.3 73.7 38.7 ;
      RECT  67.8 40.7 68.6 39.9 ;
      RECT  71.2 40.7 72.0 39.9 ;
      RECT  68.2 34.0 69.0 33.2 ;
      RECT  71.7 33.9 72.3 33.3 ;
      RECT  66.6 23.1 76.4 22.5 ;
      RECT  66.6 43.1 76.4 42.5 ;
      RECT  68.2 34.0 69.0 33.2 ;
      RECT  71.7 33.9 72.3 33.3 ;
      RECT  66.6 23.1 76.4 22.5 ;
      RECT  66.6 43.1 76.4 42.5 ;
      RECT  61.2 40.0 62.0 39.2 ;
      RECT  63.2 37.2 64.0 36.4 ;
      RECT  71.7 33.9 72.3 33.3 ;
      RECT  59.0 23.1 76.4 22.5 ;
      RECT  59.0 43.1 76.4 42.5 ;
      RECT  55.6 60.7 56.4 61.5 ;
      RECT  53.6 60.7 54.4 61.5 ;
      RECT  57.6 60.7 58.4 61.5 ;
      RECT  55.6 60.7 56.4 61.5 ;
      RECT  53.6 44.1 54.4 44.9 ;
      RECT  57.6 44.1 58.4 44.9 ;
      RECT  54.6 45.6 55.4 46.4 ;
      RECT  56.6 48.4 57.4 49.2 ;
      RECT  59.1 59.4 59.7 60.0 ;
      RECT  52.4 62.5 60.0 63.1 ;
      RECT  52.4 42.5 60.0 43.1 ;
      RECT  63.1 57.1 67.1 57.7 ;
      RECT  61.2 58.3 62.0 59.1 ;
      RECT  64.6 58.3 65.4 59.1 ;
      RECT  63.1 46.3 67.1 46.9 ;
      RECT  61.2 44.9 62.0 45.7 ;
      RECT  64.6 44.9 65.4 45.7 ;
      RECT  61.6 51.6 62.4 52.4 ;
      RECT  65.1 51.7 65.7 52.3 ;
      RECT  60.0 62.5 69.8 63.1 ;
      RECT  60.0 42.5 69.8 43.1 ;
      RECT  61.6 51.6 62.4 52.4 ;
      RECT  65.1 51.7 65.7 52.3 ;
      RECT  60.0 62.5 69.8 63.1 ;
      RECT  60.0 42.5 69.8 43.1 ;
      RECT  54.6 45.6 55.4 46.4 ;
      RECT  56.6 48.4 57.4 49.2 ;
      RECT  65.1 51.7 65.7 52.3 ;
      RECT  52.4 62.5 69.8 63.1 ;
      RECT  52.4 42.5 69.8 43.1 ;
      RECT  55.6 64.9 56.4 64.1 ;
      RECT  53.6 64.9 54.4 64.1 ;
      RECT  55.6 81.9 56.4 81.1 ;
      RECT  53.6 81.9 54.4 81.1 ;
      RECT  54.0 73.4 54.8 72.6 ;
      RECT  56.0 73.3 56.6 72.7 ;
      RECT  52.4 63.1 59.0 62.5 ;
      RECT  52.4 83.1 59.0 82.5 ;
      RECT  62.2 64.9 63.0 64.1 ;
      RECT  60.2 64.9 61.0 64.1 ;
      RECT  62.2 81.9 63.0 81.1 ;
      RECT  60.2 81.9 61.0 81.1 ;
      RECT  60.6 73.4 61.4 72.6 ;
      RECT  62.6 73.3 63.2 72.7 ;
      RECT  59.0 63.1 64.2 62.5 ;
      RECT  59.0 83.1 64.2 82.5 ;
      RECT  67.4 65.7 68.2 64.9 ;
      RECT  65.4 65.7 66.2 64.9 ;
      RECT  67.4 81.5 68.2 80.7 ;
      RECT  65.4 81.5 66.2 80.7 ;
      RECT  65.8 73.6 66.6 72.8 ;
      RECT  67.8 73.5 68.4 72.9 ;
      RECT  64.2 63.1 69.4 62.5 ;
      RECT  64.2 83.1 69.4 82.5 ;
      RECT  72.6 68.1 73.4 67.3 ;
      RECT  70.6 68.1 71.4 67.3 ;
      RECT  72.6 80.3 73.4 79.5 ;
      RECT  70.6 80.3 71.4 79.5 ;
      RECT  71.0 74.2 71.8 73.4 ;
      RECT  73.0 74.1 73.6 73.5 ;
      RECT  69.4 63.1 74.6 62.5 ;
      RECT  69.4 83.1 74.6 82.5 ;
      RECT  54.0 73.4 54.8 72.6 ;
      RECT  73.0 74.1 73.6 73.5 ;
      RECT  52.4 63.1 74.6 62.5 ;
      RECT  52.4 83.1 74.6 82.5 ;
      RECT  55.6 140.7 56.4 141.5 ;
      RECT  53.6 140.7 54.4 141.5 ;
      RECT  55.6 123.7 56.4 124.5 ;
      RECT  53.6 123.7 54.4 124.5 ;
      RECT  54.0 132.2 54.8 133.0 ;
      RECT  56.0 132.3 56.6 132.9 ;
      RECT  52.4 142.5 59.0 143.1 ;
      RECT  52.4 122.5 59.0 123.1 ;
      RECT  55.6 100.7 56.4 101.5 ;
      RECT  53.6 100.7 54.4 101.5 ;
      RECT  57.6 100.7 58.4 101.5 ;
      RECT  55.6 100.7 56.4 101.5 ;
      RECT  59.6 100.7 60.4 101.5 ;
      RECT  57.6 100.7 58.4 101.5 ;
      RECT  53.6 84.1 54.4 84.9 ;
      RECT  59.6 84.1 60.4 84.9 ;
      RECT  54.2 85.6 55.0 86.4 ;
      RECT  56.6 87.0 57.4 87.8 ;
      RECT  59.0 88.4 59.8 89.2 ;
      RECT  61.1 99.5 61.7 100.1 ;
      RECT  52.4 102.5 62.0 103.1 ;
      RECT  52.4 82.5 62.0 83.1 ;
      RECT  65.0 97.5 65.8 98.3 ;
      RECT  66.8 97.5 67.6 98.3 ;
      RECT  63.2 97.5 64.0 98.3 ;
      RECT  65.0 85.3 65.8 86.1 ;
      RECT  63.2 85.3 64.0 86.1 ;
      RECT  66.8 85.3 67.6 86.1 ;
      RECT  63.6 91.4 64.4 92.2 ;
      RECT  65.4 91.5 66.0 92.1 ;
      RECT  62.0 102.5 70.2 103.1 ;
      RECT  62.0 82.5 70.2 83.1 ;
      RECT  63.6 91.4 64.4 92.2 ;
      RECT  65.4 91.5 66.0 92.1 ;
      RECT  62.0 102.5 70.2 103.1 ;
      RECT  62.0 82.5 70.2 83.1 ;
      RECT  54.2 85.6 55.0 86.4 ;
      RECT  56.6 87.0 57.4 87.8 ;
      RECT  59.0 88.4 59.8 89.2 ;
      RECT  65.4 91.5 66.0 92.1 ;
      RECT  52.4 102.5 70.2 103.1 ;
      RECT  52.4 82.5 70.2 83.1 ;
      RECT  55.6 144.9 56.4 144.1 ;
      RECT  53.6 144.9 54.4 144.1 ;
      RECT  57.6 144.9 58.4 144.1 ;
      RECT  55.6 144.9 56.4 144.1 ;
      RECT  59.6 144.9 60.4 144.1 ;
      RECT  57.6 144.9 58.4 144.1 ;
      RECT  53.6 161.5 54.4 160.7 ;
      RECT  59.6 161.5 60.4 160.7 ;
      RECT  54.2 160.0 55.0 159.2 ;
      RECT  56.6 158.6 57.4 157.8 ;
      RECT  59.0 157.2 59.8 156.4 ;
      RECT  61.1 146.1 61.7 145.5 ;
      RECT  52.4 143.1 62.0 142.5 ;
      RECT  52.4 163.1 62.0 162.5 ;
      RECT  65.2 145.7 66.0 144.9 ;
      RECT  63.2 145.7 64.0 144.9 ;
      RECT  65.2 161.5 66.0 160.7 ;
      RECT  63.2 161.5 64.0 160.7 ;
      RECT  63.6 153.6 64.4 152.8 ;
      RECT  65.6 153.5 66.2 152.9 ;
      RECT  62.0 143.1 68.6 142.5 ;
      RECT  62.0 163.1 68.6 162.5 ;
      RECT  63.6 153.6 64.4 152.8 ;
      RECT  65.6 153.5 66.2 152.9 ;
      RECT  62.0 143.1 68.6 142.5 ;
      RECT  62.0 163.1 68.6 162.5 ;
      RECT  54.2 160.0 55.0 159.2 ;
      RECT  56.6 158.6 57.4 157.8 ;
      RECT  59.0 157.2 59.8 156.4 ;
      RECT  65.6 153.5 66.2 152.9 ;
      RECT  52.4 143.1 68.6 142.5 ;
      RECT  52.4 163.1 68.6 162.5 ;
      RECT  32.2 183.1 31.4 183.9 ;
      RECT  34.2 183.1 33.4 183.9 ;
      RECT  32.2 166.5 31.4 167.3 ;
      RECT  34.2 166.5 33.4 167.3 ;
      RECT  33.8 174.8 33.0 175.6 ;
      RECT  31.8 174.9 31.2 175.5 ;
      RECT  35.4 184.9 28.8 185.5 ;
      RECT  35.4 165.3 28.8 165.9 ;
      RECT  25.6 183.1 24.8 183.9 ;
      RECT  27.6 183.1 26.8 183.9 ;
      RECT  25.6 166.5 24.8 167.3 ;
      RECT  27.6 166.5 26.8 167.3 ;
      RECT  27.2 174.8 26.4 175.6 ;
      RECT  25.2 174.9 24.6 175.5 ;
      RECT  28.8 184.9 22.2 185.5 ;
      RECT  28.8 165.3 22.2 165.9 ;
      RECT  19.0 183.1 18.2 183.9 ;
      RECT  21.0 183.1 20.2 183.9 ;
      RECT  19.0 166.5 18.2 167.3 ;
      RECT  21.0 166.5 20.2 167.3 ;
      RECT  20.6 174.8 19.8 175.6 ;
      RECT  18.6 174.9 18.0 175.5 ;
      RECT  22.2 184.9 15.6 185.5 ;
      RECT  22.2 165.3 15.6 165.9 ;
      RECT  12.4 183.1 11.6 183.9 ;
      RECT  14.4 183.1 13.6 183.9 ;
      RECT  12.4 166.5 11.6 167.3 ;
      RECT  14.4 166.5 13.6 167.3 ;
      RECT  14.0 174.8 13.2 175.6 ;
      RECT  12.0 174.9 11.4 175.5 ;
      RECT  15.6 184.9 9.0 185.5 ;
      RECT  15.6 165.3 9.0 165.9 ;
      RECT  5.8 183.1 5.0 183.9 ;
      RECT  7.8 183.1 7.0 183.9 ;
      RECT  5.8 166.5 5.0 167.3 ;
      RECT  7.8 166.5 7.0 167.3 ;
      RECT  7.4 174.8 6.6 175.6 ;
      RECT  5.4 174.9 4.8 175.5 ;
      RECT  9.0 184.9 2.4 185.5 ;
      RECT  9.0 165.3 2.4 165.9 ;
      RECT  32.2 187.3 31.4 186.5 ;
      RECT  34.2 187.3 33.4 186.5 ;
      RECT  32.2 203.9 31.4 203.1 ;
      RECT  34.2 203.9 33.4 203.1 ;
      RECT  33.8 195.6 33.0 194.8 ;
      RECT  31.8 195.5 31.2 194.9 ;
      RECT  35.4 185.5 28.8 184.9 ;
      RECT  35.4 205.1 28.8 204.5 ;
      RECT  25.6 187.3 24.8 186.5 ;
      RECT  27.6 187.3 26.8 186.5 ;
      RECT  25.6 203.9 24.8 203.1 ;
      RECT  27.6 203.9 26.8 203.1 ;
      RECT  27.2 195.6 26.4 194.8 ;
      RECT  25.2 195.5 24.6 194.9 ;
      RECT  28.8 185.5 22.2 184.9 ;
      RECT  28.8 205.1 22.2 204.5 ;
      RECT  19.0 187.3 18.2 186.5 ;
      RECT  21.0 187.3 20.2 186.5 ;
      RECT  19.0 203.9 18.2 203.1 ;
      RECT  21.0 203.9 20.2 203.1 ;
      RECT  20.6 195.6 19.8 194.8 ;
      RECT  18.6 195.5 18.0 194.9 ;
      RECT  22.2 185.5 15.6 184.9 ;
      RECT  22.2 205.1 15.6 204.5 ;
      RECT  12.4 187.3 11.6 186.5 ;
      RECT  14.4 187.3 13.6 186.5 ;
      RECT  12.4 203.9 11.6 203.1 ;
      RECT  14.4 203.9 13.6 203.1 ;
      RECT  14.0 195.6 13.2 194.8 ;
      RECT  12.0 195.5 11.4 194.9 ;
      RECT  15.6 185.5 9.0 184.9 ;
      RECT  15.6 205.1 9.0 204.5 ;
      RECT  5.8 187.3 5.0 186.5 ;
      RECT  7.8 187.3 7.0 186.5 ;
      RECT  5.8 203.9 5.0 203.1 ;
      RECT  7.8 203.9 7.0 203.1 ;
      RECT  7.4 195.6 6.6 194.8 ;
      RECT  5.4 195.5 4.8 194.9 ;
      RECT  9.0 185.5 2.4 184.9 ;
      RECT  9.0 205.1 2.4 204.5 ;
      RECT  32.2 222.3 31.4 223.1 ;
      RECT  34.2 222.3 33.4 223.1 ;
      RECT  32.2 205.7 31.4 206.5 ;
      RECT  34.2 205.7 33.4 206.5 ;
      RECT  33.8 214.0 33.0 214.8 ;
      RECT  31.8 214.1 31.2 214.7 ;
      RECT  35.4 224.1 28.8 224.7 ;
      RECT  35.4 204.5 28.8 205.1 ;
      RECT  25.6 222.3 24.8 223.1 ;
      RECT  27.6 222.3 26.8 223.1 ;
      RECT  25.6 205.7 24.8 206.5 ;
      RECT  27.6 205.7 26.8 206.5 ;
      RECT  27.2 214.0 26.4 214.8 ;
      RECT  25.2 214.1 24.6 214.7 ;
      RECT  28.8 224.1 22.2 224.7 ;
      RECT  28.8 204.5 22.2 205.1 ;
      RECT  19.0 222.3 18.2 223.1 ;
      RECT  21.0 222.3 20.2 223.1 ;
      RECT  19.0 205.7 18.2 206.5 ;
      RECT  21.0 205.7 20.2 206.5 ;
      RECT  20.6 214.0 19.8 214.8 ;
      RECT  18.6 214.1 18.0 214.7 ;
      RECT  22.2 224.1 15.6 224.7 ;
      RECT  22.2 204.5 15.6 205.1 ;
      RECT  12.4 222.3 11.6 223.1 ;
      RECT  14.4 222.3 13.6 223.1 ;
      RECT  12.4 205.7 11.6 206.5 ;
      RECT  14.4 205.7 13.6 206.5 ;
      RECT  14.0 214.0 13.2 214.8 ;
      RECT  12.0 214.1 11.4 214.7 ;
      RECT  15.6 224.1 9.0 224.7 ;
      RECT  15.6 204.5 9.0 205.1 ;
      RECT  5.8 222.3 5.0 223.1 ;
      RECT  7.8 222.3 7.0 223.1 ;
      RECT  5.8 205.7 5.0 206.5 ;
      RECT  7.8 205.7 7.0 206.5 ;
      RECT  7.4 214.0 6.6 214.8 ;
      RECT  5.4 214.1 4.8 214.7 ;
      RECT  9.0 224.1 2.4 224.7 ;
      RECT  9.0 204.5 2.4 205.1 ;
      RECT  32.2 226.5 31.4 225.7 ;
      RECT  34.2 226.5 33.4 225.7 ;
      RECT  32.2 243.1 31.4 242.3 ;
      RECT  34.2 243.1 33.4 242.3 ;
      RECT  33.8 234.8 33.0 234.0 ;
      RECT  31.8 234.7 31.2 234.1 ;
      RECT  35.4 224.7 28.8 224.1 ;
      RECT  35.4 244.3 28.8 243.7 ;
      RECT  25.6 226.5 24.8 225.7 ;
      RECT  27.6 226.5 26.8 225.7 ;
      RECT  25.6 243.1 24.8 242.3 ;
      RECT  27.6 243.1 26.8 242.3 ;
      RECT  27.2 234.8 26.4 234.0 ;
      RECT  25.2 234.7 24.6 234.1 ;
      RECT  28.8 224.7 22.2 224.1 ;
      RECT  28.8 244.3 22.2 243.7 ;
      RECT  19.0 226.5 18.2 225.7 ;
      RECT  21.0 226.5 20.2 225.7 ;
      RECT  19.0 243.1 18.2 242.3 ;
      RECT  21.0 243.1 20.2 242.3 ;
      RECT  20.6 234.8 19.8 234.0 ;
      RECT  18.6 234.7 18.0 234.1 ;
      RECT  22.2 224.7 15.6 224.1 ;
      RECT  22.2 244.3 15.6 243.7 ;
      RECT  12.4 226.5 11.6 225.7 ;
      RECT  14.4 226.5 13.6 225.7 ;
      RECT  12.4 243.1 11.6 242.3 ;
      RECT  14.4 243.1 13.6 242.3 ;
      RECT  14.0 234.8 13.2 234.0 ;
      RECT  12.0 234.7 11.4 234.1 ;
      RECT  15.6 224.7 9.0 224.1 ;
      RECT  15.6 244.3 9.0 243.7 ;
      RECT  5.8 226.5 5.0 225.7 ;
      RECT  7.8 226.5 7.0 225.7 ;
      RECT  5.8 243.1 5.0 242.3 ;
      RECT  7.8 243.1 7.0 242.3 ;
      RECT  7.4 234.8 6.6 234.0 ;
      RECT  5.4 234.7 4.8 234.1 ;
      RECT  9.0 224.7 2.4 224.1 ;
      RECT  9.0 244.3 2.4 243.7 ;
      RECT  32.2 261.5 31.4 262.3 ;
      RECT  34.2 261.5 33.4 262.3 ;
      RECT  32.2 244.9 31.4 245.7 ;
      RECT  34.2 244.9 33.4 245.7 ;
      RECT  33.8 253.2 33.0 254.0 ;
      RECT  31.8 253.3 31.2 253.9 ;
      RECT  35.4 263.3 28.8 263.9 ;
      RECT  35.4 243.7 28.8 244.3 ;
      RECT  25.6 261.5 24.8 262.3 ;
      RECT  27.6 261.5 26.8 262.3 ;
      RECT  25.6 244.9 24.8 245.7 ;
      RECT  27.6 244.9 26.8 245.7 ;
      RECT  27.2 253.2 26.4 254.0 ;
      RECT  25.2 253.3 24.6 253.9 ;
      RECT  28.8 263.3 22.2 263.9 ;
      RECT  28.8 243.7 22.2 244.3 ;
      RECT  19.0 261.5 18.2 262.3 ;
      RECT  21.0 261.5 20.2 262.3 ;
      RECT  19.0 244.9 18.2 245.7 ;
      RECT  21.0 244.9 20.2 245.7 ;
      RECT  20.6 253.2 19.8 254.0 ;
      RECT  18.6 253.3 18.0 253.9 ;
      RECT  22.2 263.3 15.6 263.9 ;
      RECT  22.2 243.7 15.6 244.3 ;
      RECT  12.4 261.5 11.6 262.3 ;
      RECT  14.4 261.5 13.6 262.3 ;
      RECT  12.4 244.9 11.6 245.7 ;
      RECT  14.4 244.9 13.6 245.7 ;
      RECT  14.0 253.2 13.2 254.0 ;
      RECT  12.0 253.3 11.4 253.9 ;
      RECT  15.6 263.3 9.0 263.9 ;
      RECT  15.6 243.7 9.0 244.3 ;
      RECT  5.8 261.5 5.0 262.3 ;
      RECT  7.8 261.5 7.0 262.3 ;
      RECT  5.8 244.9 5.0 245.7 ;
      RECT  7.8 244.9 7.0 245.7 ;
      RECT  7.4 253.2 6.6 254.0 ;
      RECT  5.4 253.3 4.8 253.9 ;
      RECT  9.0 263.3 2.4 263.9 ;
      RECT  9.0 243.7 2.4 244.3 ;
      RECT  32.2 265.7 31.4 264.9 ;
      RECT  34.2 265.7 33.4 264.9 ;
      RECT  32.2 282.3 31.4 281.5 ;
      RECT  34.2 282.3 33.4 281.5 ;
      RECT  33.8 274.0 33.0 273.2 ;
      RECT  31.8 273.9 31.2 273.3 ;
      RECT  35.4 263.9 28.8 263.3 ;
      RECT  35.4 283.5 28.8 282.9 ;
      RECT  25.6 265.7 24.8 264.9 ;
      RECT  27.6 265.7 26.8 264.9 ;
      RECT  25.6 282.3 24.8 281.5 ;
      RECT  27.6 282.3 26.8 281.5 ;
      RECT  27.2 274.0 26.4 273.2 ;
      RECT  25.2 273.9 24.6 273.3 ;
      RECT  28.8 263.9 22.2 263.3 ;
      RECT  28.8 283.5 22.2 282.9 ;
      RECT  19.0 265.7 18.2 264.9 ;
      RECT  21.0 265.7 20.2 264.9 ;
      RECT  19.0 282.3 18.2 281.5 ;
      RECT  21.0 282.3 20.2 281.5 ;
      RECT  20.6 274.0 19.8 273.2 ;
      RECT  18.6 273.9 18.0 273.3 ;
      RECT  22.2 263.9 15.6 263.3 ;
      RECT  22.2 283.5 15.6 282.9 ;
      RECT  12.4 265.7 11.6 264.9 ;
      RECT  14.4 265.7 13.6 264.9 ;
      RECT  12.4 282.3 11.6 281.5 ;
      RECT  14.4 282.3 13.6 281.5 ;
      RECT  14.0 274.0 13.2 273.2 ;
      RECT  12.0 273.9 11.4 273.3 ;
      RECT  15.6 263.9 9.0 263.3 ;
      RECT  15.6 283.5 9.0 282.9 ;
      RECT  5.8 265.7 5.0 264.9 ;
      RECT  7.8 265.7 7.0 264.9 ;
      RECT  5.8 282.3 5.0 281.5 ;
      RECT  7.8 282.3 7.0 281.5 ;
      RECT  7.4 274.0 6.6 273.2 ;
      RECT  5.4 273.9 4.8 273.3 ;
      RECT  9.0 263.9 2.4 263.3 ;
      RECT  9.0 283.5 2.4 282.9 ;
      RECT  32.2 300.7 31.4 301.5 ;
      RECT  34.2 300.7 33.4 301.5 ;
      RECT  32.2 284.1 31.4 284.9 ;
      RECT  34.2 284.1 33.4 284.9 ;
      RECT  33.8 292.4 33.0 293.2 ;
      RECT  31.8 292.5 31.2 293.1 ;
      RECT  35.4 302.5 28.8 303.1 ;
      RECT  35.4 282.9 28.8 283.5 ;
      RECT  25.6 300.7 24.8 301.5 ;
      RECT  27.6 300.7 26.8 301.5 ;
      RECT  25.6 284.1 24.8 284.9 ;
      RECT  27.6 284.1 26.8 284.9 ;
      RECT  27.2 292.4 26.4 293.2 ;
      RECT  25.2 292.5 24.6 293.1 ;
      RECT  28.8 302.5 22.2 303.1 ;
      RECT  28.8 282.9 22.2 283.5 ;
      RECT  19.0 300.7 18.2 301.5 ;
      RECT  21.0 300.7 20.2 301.5 ;
      RECT  19.0 284.1 18.2 284.9 ;
      RECT  21.0 284.1 20.2 284.9 ;
      RECT  20.6 292.4 19.8 293.2 ;
      RECT  18.6 292.5 18.0 293.1 ;
      RECT  22.2 302.5 15.6 303.1 ;
      RECT  22.2 282.9 15.6 283.5 ;
      RECT  12.4 300.7 11.6 301.5 ;
      RECT  14.4 300.7 13.6 301.5 ;
      RECT  12.4 284.1 11.6 284.9 ;
      RECT  14.4 284.1 13.6 284.9 ;
      RECT  14.0 292.4 13.2 293.2 ;
      RECT  12.0 292.5 11.4 293.1 ;
      RECT  15.6 302.5 9.0 303.1 ;
      RECT  15.6 282.9 9.0 283.5 ;
      RECT  5.8 300.7 5.0 301.5 ;
      RECT  7.8 300.7 7.0 301.5 ;
      RECT  5.8 284.1 5.0 284.9 ;
      RECT  7.8 284.1 7.0 284.9 ;
      RECT  7.4 292.4 6.6 293.2 ;
      RECT  5.4 292.5 4.8 293.1 ;
      RECT  9.0 302.5 2.4 303.1 ;
      RECT  9.0 282.9 2.4 283.5 ;
      RECT  32.2 304.9 31.4 304.1 ;
      RECT  34.2 304.9 33.4 304.1 ;
      RECT  32.2 321.5 31.4 320.7 ;
      RECT  34.2 321.5 33.4 320.7 ;
      RECT  33.8 313.2 33.0 312.4 ;
      RECT  31.8 313.1 31.2 312.5 ;
      RECT  35.4 303.1 28.8 302.5 ;
      RECT  35.4 322.7 28.8 322.1 ;
      RECT  25.6 304.9 24.8 304.1 ;
      RECT  27.6 304.9 26.8 304.1 ;
      RECT  25.6 321.5 24.8 320.7 ;
      RECT  27.6 321.5 26.8 320.7 ;
      RECT  27.2 313.2 26.4 312.4 ;
      RECT  25.2 313.1 24.6 312.5 ;
      RECT  28.8 303.1 22.2 302.5 ;
      RECT  28.8 322.7 22.2 322.1 ;
      RECT  19.0 304.9 18.2 304.1 ;
      RECT  21.0 304.9 20.2 304.1 ;
      RECT  19.0 321.5 18.2 320.7 ;
      RECT  21.0 321.5 20.2 320.7 ;
      RECT  20.6 313.2 19.8 312.4 ;
      RECT  18.6 313.1 18.0 312.5 ;
      RECT  22.2 303.1 15.6 302.5 ;
      RECT  22.2 322.7 15.6 322.1 ;
      RECT  12.4 304.9 11.6 304.1 ;
      RECT  14.4 304.9 13.6 304.1 ;
      RECT  12.4 321.5 11.6 320.7 ;
      RECT  14.4 321.5 13.6 320.7 ;
      RECT  14.0 313.2 13.2 312.4 ;
      RECT  12.0 313.1 11.4 312.5 ;
      RECT  15.6 303.1 9.0 302.5 ;
      RECT  15.6 322.7 9.0 322.1 ;
      RECT  5.8 304.9 5.0 304.1 ;
      RECT  7.8 304.9 7.0 304.1 ;
      RECT  5.8 321.5 5.0 320.7 ;
      RECT  7.8 321.5 7.0 320.7 ;
      RECT  7.4 313.2 6.6 312.4 ;
      RECT  5.4 313.1 4.8 312.5 ;
      RECT  9.0 303.1 2.4 302.5 ;
      RECT  9.0 322.7 2.4 322.1 ;
      RECT  32.2 339.9 31.4 340.7 ;
      RECT  34.2 339.9 33.4 340.7 ;
      RECT  32.2 323.3 31.4 324.1 ;
      RECT  34.2 323.3 33.4 324.1 ;
      RECT  33.8 331.6 33.0 332.4 ;
      RECT  31.8 331.7 31.2 332.3 ;
      RECT  35.4 341.7 28.8 342.3 ;
      RECT  35.4 322.1 28.8 322.7 ;
      RECT  25.6 339.9 24.8 340.7 ;
      RECT  27.6 339.9 26.8 340.7 ;
      RECT  25.6 323.3 24.8 324.1 ;
      RECT  27.6 323.3 26.8 324.1 ;
      RECT  27.2 331.6 26.4 332.4 ;
      RECT  25.2 331.7 24.6 332.3 ;
      RECT  28.8 341.7 22.2 342.3 ;
      RECT  28.8 322.1 22.2 322.7 ;
      RECT  19.0 339.9 18.2 340.7 ;
      RECT  21.0 339.9 20.2 340.7 ;
      RECT  19.0 323.3 18.2 324.1 ;
      RECT  21.0 323.3 20.2 324.1 ;
      RECT  20.6 331.6 19.8 332.4 ;
      RECT  18.6 331.7 18.0 332.3 ;
      RECT  22.2 341.7 15.6 342.3 ;
      RECT  22.2 322.1 15.6 322.7 ;
      RECT  12.4 339.9 11.6 340.7 ;
      RECT  14.4 339.9 13.6 340.7 ;
      RECT  12.4 323.3 11.6 324.1 ;
      RECT  14.4 323.3 13.6 324.1 ;
      RECT  14.0 331.6 13.2 332.4 ;
      RECT  12.0 331.7 11.4 332.3 ;
      RECT  15.6 341.7 9.0 342.3 ;
      RECT  15.6 322.1 9.0 322.7 ;
      RECT  5.8 339.9 5.0 340.7 ;
      RECT  7.8 339.9 7.0 340.7 ;
      RECT  5.8 323.3 5.0 324.1 ;
      RECT  7.8 323.3 7.0 324.1 ;
      RECT  7.4 331.6 6.6 332.4 ;
      RECT  5.4 331.7 4.8 332.3 ;
      RECT  9.0 341.7 2.4 342.3 ;
      RECT  9.0 322.1 2.4 322.7 ;
      RECT  55.6 104.9 56.4 104.1 ;
      RECT  53.6 104.9 54.4 104.1 ;
      RECT  57.6 104.9 58.4 104.1 ;
      RECT  55.6 104.9 56.4 104.1 ;
      RECT  53.6 121.5 54.4 120.7 ;
      RECT  57.6 121.5 58.4 120.7 ;
      RECT  54.6 120.0 55.4 119.2 ;
      RECT  56.6 117.2 57.4 116.4 ;
      RECT  59.1 106.2 59.7 105.6 ;
      RECT  52.4 103.1 61.0 102.5 ;
      RECT  52.4 123.1 61.0 122.5 ;
      RECT  64.2 104.9 65.0 104.1 ;
      RECT  62.2 104.9 63.0 104.1 ;
      RECT  64.2 121.9 65.0 121.1 ;
      RECT  62.2 121.9 63.0 121.1 ;
      RECT  62.6 113.4 63.4 112.6 ;
      RECT  64.6 113.3 65.2 112.7 ;
      RECT  61.0 103.1 67.6 102.5 ;
      RECT  61.0 123.1 67.6 122.5 ;
      RECT  70.8 104.9 71.6 104.1 ;
      RECT  68.8 104.9 69.6 104.1 ;
      RECT  70.8 121.9 71.6 121.1 ;
      RECT  68.8 121.9 69.6 121.1 ;
      RECT  69.2 113.4 70.0 112.6 ;
      RECT  71.2 113.3 71.8 112.7 ;
      RECT  67.6 103.1 72.8 102.5 ;
      RECT  67.6 123.1 72.8 122.5 ;
      RECT  62.6 113.4 63.4 112.6 ;
      RECT  71.2 113.3 71.8 112.7 ;
      RECT  61.0 103.1 72.8 102.5 ;
      RECT  61.0 123.1 72.8 122.5 ;
      RECT  58.8 355.0 68.6 355.2 ;
      RECT  73.0 354.4 77.2 355.0 ;
      RECT  76.4 346.0 77.2 350.4 ;
      RECT  65.4 358.4 69.0 359.0 ;
      RECT  76.4 351.0 77.2 354.4 ;
      RECT  65.4 349.2 66.2 349.4 ;
      RECT  68.0 356.8 70.2 357.4 ;
      RECT  58.8 346.0 59.6 350.8 ;
      RECT  69.4 351.4 70.2 351.6 ;
      RECT  65.4 358.2 66.2 358.4 ;
      RECT  69.4 356.6 70.2 356.8 ;
      RECT  62.0 356.8 62.8 357.0 ;
      RECT  70.0 355.4 72.4 356.0 ;
      RECT  62.6 352.2 63.4 352.4 ;
      RECT  76.4 355.0 77.2 363.6 ;
      RECT  73.4 350.2 74.2 350.4 ;
      RECT  71.6 353.0 75.4 353.6 ;
      RECT  63.8 349.4 64.4 351.6 ;
      RECT  65.8 345.4 66.8 348.0 ;
      RECT  74.8 345.4 75.6 349.8 ;
      RECT  66.6 356.8 67.4 357.0 ;
      RECT  74.6 353.6 75.4 353.8 ;
      RECT  67.6 359.6 68.4 363.6 ;
      RECT  62.0 358.8 62.8 359.6 ;
      RECT  71.6 358.8 72.4 359.6 ;
      RECT  63.8 355.2 68.6 355.6 ;
      RECT  58.8 354.8 64.6 355.0 ;
      RECT  61.0 353.4 66.0 354.0 ;
      RECT  68.2 358.2 69.0 358.4 ;
      RECT  62.0 359.6 64.0 360.2 ;
      RECT  60.4 345.4 61.2 350.0 ;
      RECT  65.4 348.6 68.2 349.2 ;
      RECT  78.0 345.4 78.8 346.8 ;
      RECT  58.8 355.2 59.6 363.6 ;
      RECT  60.4 355.8 61.2 364.2 ;
      RECT  71.8 356.0 72.4 357.0 ;
      RECT  71.6 347.4 73.0 348.0 ;
      RECT  66.0 359.6 66.8 364.2 ;
      RECT  69.2 359.6 70.0 364.2 ;
      RECT  71.8 357.0 73.2 357.8 ;
      RECT  70.0 352.2 70.6 355.4 ;
      RECT  59.6 351.4 61.2 351.6 ;
      RECT  62.0 347.4 64.0 348.0 ;
      RECT  63.2 346.0 64.0 347.4 ;
      RECT  71.8 359.6 73.0 363.6 ;
      RECT  63.6 348.6 64.4 349.4 ;
      RECT  68.0 355.6 68.6 356.8 ;
      RECT  65.2 354.0 66.0 354.2 ;
      RECT  71.6 352.8 72.4 353.0 ;
      RECT  67.6 359.0 68.2 359.6 ;
      RECT  62.0 356.2 67.4 356.8 ;
      RECT  67.6 346.0 68.4 348.0 ;
      RECT  57.6 364.2 79.4 365.4 ;
      RECT  63.2 360.2 64.0 363.6 ;
      RECT  74.8 355.6 75.6 364.2 ;
      RECT  58.8 354.6 64.4 354.8 ;
      RECT  61.0 353.2 61.8 353.4 ;
      RECT  69.2 345.4 70.0 348.0 ;
      RECT  71.8 346.0 73.0 347.4 ;
      RECT  57.6 344.2 79.4 345.4 ;
      RECT  78.0 362.6 78.8 364.2 ;
      RECT  59.6 351.6 70.6 352.2 ;
      RECT  73.4 350.4 77.2 351.0 ;
      RECT  62.0 348.0 62.8 348.8 ;
      RECT  67.6 348.0 68.2 348.6 ;
      RECT  71.6 348.0 72.4 348.8 ;
      RECT  73.0 354.2 73.8 354.4 ;
      RECT  58.8 374.6 68.6 374.4 ;
      RECT  73.0 375.2 77.2 374.6 ;
      RECT  76.4 383.6 77.2 379.2 ;
      RECT  65.4 371.2 69.0 370.6 ;
      RECT  76.4 378.6 77.2 375.2 ;
      RECT  65.4 380.4 66.2 380.2 ;
      RECT  68.0 372.8 70.2 372.2 ;
      RECT  58.8 383.6 59.6 378.8 ;
      RECT  69.4 378.2 70.2 378.0 ;
      RECT  65.4 371.4 66.2 371.2 ;
      RECT  69.4 373.0 70.2 372.8 ;
      RECT  62.0 372.8 62.8 372.6 ;
      RECT  70.0 374.2 72.4 373.6 ;
      RECT  62.6 377.4 63.4 377.2 ;
      RECT  76.4 374.6 77.2 366.0 ;
      RECT  73.4 379.4 74.2 379.2 ;
      RECT  71.6 376.6 75.4 376.0 ;
      RECT  63.8 380.2 64.4 378.0 ;
      RECT  65.8 384.2 66.8 381.6 ;
      RECT  74.8 384.2 75.6 379.8 ;
      RECT  66.6 372.8 67.4 372.6 ;
      RECT  74.6 376.0 75.4 375.8 ;
      RECT  67.6 370.0 68.4 366.0 ;
      RECT  62.0 370.8 62.8 370.0 ;
      RECT  71.6 370.8 72.4 370.0 ;
      RECT  63.8 374.4 68.6 374.0 ;
      RECT  58.8 374.8 64.6 374.6 ;
      RECT  61.0 376.2 66.0 375.6 ;
      RECT  68.2 371.4 69.0 371.2 ;
      RECT  62.0 370.0 64.0 369.4 ;
      RECT  60.4 384.2 61.2 379.6 ;
      RECT  65.4 381.0 68.2 380.4 ;
      RECT  78.0 384.2 78.8 382.8 ;
      RECT  58.8 374.4 59.6 366.0 ;
      RECT  60.4 373.8 61.2 365.4 ;
      RECT  71.8 373.6 72.4 372.6 ;
      RECT  71.6 382.2 73.0 381.6 ;
      RECT  66.0 370.0 66.8 365.4 ;
      RECT  69.2 370.0 70.0 365.4 ;
      RECT  71.8 372.6 73.2 371.8 ;
      RECT  70.0 377.4 70.6 374.2 ;
      RECT  59.6 378.2 61.2 378.0 ;
      RECT  62.0 382.2 64.0 381.6 ;
      RECT  63.2 383.6 64.0 382.2 ;
      RECT  71.8 370.0 73.0 366.0 ;
      RECT  63.6 381.0 64.4 380.2 ;
      RECT  68.0 374.0 68.6 372.8 ;
      RECT  65.2 375.6 66.0 375.4 ;
      RECT  71.6 376.8 72.4 376.6 ;
      RECT  67.6 370.6 68.2 370.0 ;
      RECT  62.0 373.4 67.4 372.8 ;
      RECT  67.6 383.6 68.4 381.6 ;
      RECT  57.6 365.4 79.4 364.2 ;
      RECT  63.2 369.4 64.0 366.0 ;
      RECT  74.8 374.0 75.6 365.4 ;
      RECT  58.8 375.0 64.4 374.8 ;
      RECT  61.0 376.4 61.8 376.2 ;
      RECT  69.2 384.2 70.0 381.6 ;
      RECT  71.8 383.6 73.0 382.2 ;
      RECT  57.6 385.4 79.4 384.2 ;
      RECT  78.0 367.0 78.8 365.4 ;
      RECT  59.6 378.0 70.6 377.4 ;
      RECT  73.4 379.2 77.2 378.6 ;
      RECT  62.0 381.6 62.8 380.8 ;
      RECT  67.6 381.6 68.2 381.0 ;
      RECT  71.6 381.6 72.4 380.8 ;
      RECT  73.0 375.4 73.8 375.2 ;
      RECT  58.8 395.0 68.6 395.2 ;
      RECT  73.0 394.4 77.2 395.0 ;
      RECT  76.4 386.0 77.2 390.4 ;
      RECT  65.4 398.4 69.0 399.0 ;
      RECT  76.4 391.0 77.2 394.4 ;
      RECT  65.4 389.2 66.2 389.4 ;
      RECT  68.0 396.8 70.2 397.4 ;
      RECT  58.8 386.0 59.6 390.8 ;
      RECT  69.4 391.4 70.2 391.6 ;
      RECT  65.4 398.2 66.2 398.4 ;
      RECT  69.4 396.6 70.2 396.8 ;
      RECT  62.0 396.8 62.8 397.0 ;
      RECT  70.0 395.4 72.4 396.0 ;
      RECT  62.6 392.2 63.4 392.4 ;
      RECT  76.4 395.0 77.2 403.6 ;
      RECT  73.4 390.2 74.2 390.4 ;
      RECT  71.6 393.0 75.4 393.6 ;
      RECT  63.8 389.4 64.4 391.6 ;
      RECT  65.8 385.4 66.8 388.0 ;
      RECT  74.8 385.4 75.6 389.8 ;
      RECT  66.6 396.8 67.4 397.0 ;
      RECT  74.6 393.6 75.4 393.8 ;
      RECT  67.6 399.6 68.4 403.6 ;
      RECT  62.0 398.8 62.8 399.6 ;
      RECT  71.6 398.8 72.4 399.6 ;
      RECT  63.8 395.2 68.6 395.6 ;
      RECT  58.8 394.8 64.6 395.0 ;
      RECT  61.0 393.4 66.0 394.0 ;
      RECT  68.2 398.2 69.0 398.4 ;
      RECT  62.0 399.6 64.0 400.2 ;
      RECT  60.4 385.4 61.2 390.0 ;
      RECT  65.4 388.6 68.2 389.2 ;
      RECT  78.0 385.4 78.8 386.8 ;
      RECT  58.8 395.2 59.6 403.6 ;
      RECT  60.4 395.8 61.2 404.2 ;
      RECT  71.8 396.0 72.4 397.0 ;
      RECT  71.6 387.4 73.0 388.0 ;
      RECT  66.0 399.6 66.8 404.2 ;
      RECT  69.2 399.6 70.0 404.2 ;
      RECT  71.8 397.0 73.2 397.8 ;
      RECT  70.0 392.2 70.6 395.4 ;
      RECT  59.6 391.4 61.2 391.6 ;
      RECT  62.0 387.4 64.0 388.0 ;
      RECT  63.2 386.0 64.0 387.4 ;
      RECT  71.8 399.6 73.0 403.6 ;
      RECT  63.6 388.6 64.4 389.4 ;
      RECT  68.0 395.6 68.6 396.8 ;
      RECT  65.2 394.0 66.0 394.2 ;
      RECT  71.6 392.8 72.4 393.0 ;
      RECT  67.6 399.0 68.2 399.6 ;
      RECT  62.0 396.2 67.4 396.8 ;
      RECT  67.6 386.0 68.4 388.0 ;
      RECT  57.6 404.2 79.4 405.4 ;
      RECT  63.2 400.2 64.0 403.6 ;
      RECT  74.8 395.6 75.6 404.2 ;
      RECT  58.8 394.6 64.4 394.8 ;
      RECT  61.0 393.2 61.8 393.4 ;
      RECT  69.2 385.4 70.0 388.0 ;
      RECT  71.8 386.0 73.0 387.4 ;
      RECT  57.6 384.2 79.4 385.4 ;
      RECT  78.0 402.6 78.8 404.2 ;
      RECT  59.6 391.6 70.6 392.2 ;
      RECT  73.4 390.4 77.2 391.0 ;
      RECT  62.0 388.0 62.8 388.8 ;
      RECT  67.6 388.0 68.2 388.6 ;
      RECT  71.6 388.0 72.4 388.8 ;
      RECT  73.0 394.2 73.8 394.4 ;
      RECT  58.8 414.6 68.6 414.4 ;
      RECT  73.0 415.2 77.2 414.6 ;
      RECT  76.4 423.6 77.2 419.2 ;
      RECT  65.4 411.2 69.0 410.6 ;
      RECT  76.4 418.6 77.2 415.2 ;
      RECT  65.4 420.4 66.2 420.2 ;
      RECT  68.0 412.8 70.2 412.2 ;
      RECT  58.8 423.6 59.6 418.8 ;
      RECT  69.4 418.2 70.2 418.0 ;
      RECT  65.4 411.4 66.2 411.2 ;
      RECT  69.4 413.0 70.2 412.8 ;
      RECT  62.0 412.8 62.8 412.6 ;
      RECT  70.0 414.2 72.4 413.6 ;
      RECT  62.6 417.4 63.4 417.2 ;
      RECT  76.4 414.6 77.2 406.0 ;
      RECT  73.4 419.4 74.2 419.2 ;
      RECT  71.6 416.6 75.4 416.0 ;
      RECT  63.8 420.2 64.4 418.0 ;
      RECT  65.8 424.2 66.8 421.6 ;
      RECT  74.8 424.2 75.6 419.8 ;
      RECT  66.6 412.8 67.4 412.6 ;
      RECT  74.6 416.0 75.4 415.8 ;
      RECT  67.6 410.0 68.4 406.0 ;
      RECT  62.0 410.8 62.8 410.0 ;
      RECT  71.6 410.8 72.4 410.0 ;
      RECT  63.8 414.4 68.6 414.0 ;
      RECT  58.8 414.8 64.6 414.6 ;
      RECT  61.0 416.2 66.0 415.6 ;
      RECT  68.2 411.4 69.0 411.2 ;
      RECT  62.0 410.0 64.0 409.4 ;
      RECT  60.4 424.2 61.2 419.6 ;
      RECT  65.4 421.0 68.2 420.4 ;
      RECT  78.0 424.2 78.8 422.8 ;
      RECT  58.8 414.4 59.6 406.0 ;
      RECT  60.4 413.8 61.2 405.4 ;
      RECT  71.8 413.6 72.4 412.6 ;
      RECT  71.6 422.2 73.0 421.6 ;
      RECT  66.0 410.0 66.8 405.4 ;
      RECT  69.2 410.0 70.0 405.4 ;
      RECT  71.8 412.6 73.2 411.8 ;
      RECT  70.0 417.4 70.6 414.2 ;
      RECT  59.6 418.2 61.2 418.0 ;
      RECT  62.0 422.2 64.0 421.6 ;
      RECT  63.2 423.6 64.0 422.2 ;
      RECT  71.8 410.0 73.0 406.0 ;
      RECT  63.6 421.0 64.4 420.2 ;
      RECT  68.0 414.0 68.6 412.8 ;
      RECT  65.2 415.6 66.0 415.4 ;
      RECT  71.6 416.8 72.4 416.6 ;
      RECT  67.6 410.6 68.2 410.0 ;
      RECT  62.0 413.4 67.4 412.8 ;
      RECT  67.6 423.6 68.4 421.6 ;
      RECT  57.6 405.4 79.4 404.2 ;
      RECT  63.2 409.4 64.0 406.0 ;
      RECT  74.8 414.0 75.6 405.4 ;
      RECT  58.8 415.0 64.4 414.8 ;
      RECT  61.0 416.4 61.8 416.2 ;
      RECT  69.2 424.2 70.0 421.6 ;
      RECT  71.8 423.6 73.0 422.2 ;
      RECT  57.6 425.4 79.4 424.2 ;
      RECT  78.0 407.0 78.8 405.4 ;
      RECT  59.6 418.0 70.6 417.4 ;
      RECT  73.4 419.2 77.2 418.6 ;
      RECT  62.0 421.6 62.8 420.8 ;
      RECT  67.6 421.6 68.2 421.0 ;
      RECT  71.6 421.6 72.4 420.8 ;
      RECT  73.0 415.4 73.8 415.2 ;
      RECT  102.4 13.0 112.2 13.2 ;
      RECT  116.6 12.4 120.8 13.0 ;
      RECT  120.0 4.0 120.8 8.4 ;
      RECT  109.0 16.4 112.6 17.0 ;
      RECT  120.0 9.0 120.8 12.4 ;
      RECT  109.0 7.2 109.8 7.4 ;
      RECT  111.6 14.8 113.8 15.4 ;
      RECT  102.4 4.0 103.2 8.8 ;
      RECT  113.0 9.4 113.8 9.6 ;
      RECT  109.0 16.2 109.8 16.4 ;
      RECT  113.0 14.6 113.8 14.8 ;
      RECT  105.6 14.8 106.4 15.0 ;
      RECT  113.6 13.4 116.0 14.0 ;
      RECT  106.2 10.2 107.0 10.4 ;
      RECT  120.0 13.0 120.8 21.6 ;
      RECT  117.0 8.2 117.8 8.4 ;
      RECT  115.2 11.0 119.0 11.6 ;
      RECT  107.4 7.4 108.0 9.6 ;
      RECT  109.4 3.4 110.4 6.0 ;
      RECT  118.4 3.4 119.2 7.8 ;
      RECT  110.2 14.8 111.0 15.0 ;
      RECT  118.2 11.6 119.0 11.8 ;
      RECT  111.2 17.6 112.0 21.6 ;
      RECT  105.6 16.8 106.4 17.6 ;
      RECT  115.2 16.8 116.0 17.6 ;
      RECT  107.4 13.2 112.2 13.6 ;
      RECT  102.4 12.8 108.2 13.0 ;
      RECT  104.6 11.4 109.6 12.0 ;
      RECT  111.8 16.2 112.6 16.4 ;
      RECT  105.6 17.6 107.6 18.2 ;
      RECT  104.0 3.4 104.8 8.0 ;
      RECT  109.0 6.6 111.8 7.2 ;
      RECT  121.6 3.4 122.4 4.8 ;
      RECT  102.4 13.2 103.2 21.6 ;
      RECT  104.0 13.8 104.8 22.2 ;
      RECT  115.4 14.0 116.0 15.0 ;
      RECT  115.2 5.4 116.6 6.0 ;
      RECT  109.6 17.6 110.4 22.2 ;
      RECT  112.8 17.6 113.6 22.2 ;
      RECT  115.4 15.0 116.8 15.8 ;
      RECT  113.6 10.2 114.2 13.4 ;
      RECT  103.2 9.4 104.8 9.6 ;
      RECT  105.6 5.4 107.6 6.0 ;
      RECT  106.8 4.0 107.6 5.4 ;
      RECT  115.4 17.6 116.6 21.6 ;
      RECT  107.2 6.6 108.0 7.4 ;
      RECT  111.6 13.6 112.2 14.8 ;
      RECT  108.8 12.0 109.6 12.2 ;
      RECT  115.2 10.8 116.0 11.0 ;
      RECT  111.2 17.0 111.8 17.6 ;
      RECT  105.6 14.2 111.0 14.8 ;
      RECT  111.2 4.0 112.0 6.0 ;
      RECT  101.2 22.2 123.0 23.4 ;
      RECT  106.8 18.2 107.6 21.6 ;
      RECT  118.4 13.6 119.2 22.2 ;
      RECT  102.4 12.6 108.0 12.8 ;
      RECT  104.6 11.2 105.4 11.4 ;
      RECT  112.8 3.4 113.6 6.0 ;
      RECT  115.4 4.0 116.6 5.4 ;
      RECT  101.2 2.2 123.0 3.4 ;
      RECT  121.6 20.6 122.4 22.2 ;
      RECT  103.2 9.6 114.2 10.2 ;
      RECT  117.0 8.4 120.8 9.0 ;
      RECT  105.6 6.0 106.4 6.8 ;
      RECT  111.2 6.0 111.8 6.6 ;
      RECT  115.2 6.0 116.0 6.8 ;
      RECT  116.6 12.2 117.4 12.4 ;
      RECT  124.2 13.0 134.0 13.2 ;
      RECT  138.4 12.4 142.6 13.0 ;
      RECT  141.8 4.0 142.6 8.4 ;
      RECT  130.8 16.4 134.4 17.0 ;
      RECT  141.8 9.0 142.6 12.4 ;
      RECT  130.8 7.2 131.6 7.4 ;
      RECT  133.4 14.8 135.6 15.4 ;
      RECT  124.2 4.0 125.0 8.8 ;
      RECT  134.8 9.4 135.6 9.6 ;
      RECT  130.8 16.2 131.6 16.4 ;
      RECT  134.8 14.6 135.6 14.8 ;
      RECT  127.4 14.8 128.2 15.0 ;
      RECT  135.4 13.4 137.8 14.0 ;
      RECT  128.0 10.2 128.8 10.4 ;
      RECT  141.8 13.0 142.6 21.6 ;
      RECT  138.8 8.2 139.6 8.4 ;
      RECT  137.0 11.0 140.8 11.6 ;
      RECT  129.2 7.4 129.8 9.6 ;
      RECT  131.2 3.4 132.2 6.0 ;
      RECT  140.2 3.4 141.0 7.8 ;
      RECT  132.0 14.8 132.8 15.0 ;
      RECT  140.0 11.6 140.8 11.8 ;
      RECT  133.0 17.6 133.8 21.6 ;
      RECT  127.4 16.8 128.2 17.6 ;
      RECT  137.0 16.8 137.8 17.6 ;
      RECT  129.2 13.2 134.0 13.6 ;
      RECT  124.2 12.8 130.0 13.0 ;
      RECT  126.4 11.4 131.4 12.0 ;
      RECT  133.6 16.2 134.4 16.4 ;
      RECT  127.4 17.6 129.4 18.2 ;
      RECT  125.8 3.4 126.6 8.0 ;
      RECT  130.8 6.6 133.6 7.2 ;
      RECT  143.4 3.4 144.2 4.8 ;
      RECT  124.2 13.2 125.0 21.6 ;
      RECT  125.8 13.8 126.6 22.2 ;
      RECT  137.2 14.0 137.8 15.0 ;
      RECT  137.0 5.4 138.4 6.0 ;
      RECT  131.4 17.6 132.2 22.2 ;
      RECT  134.6 17.6 135.4 22.2 ;
      RECT  137.2 15.0 138.6 15.8 ;
      RECT  135.4 10.2 136.0 13.4 ;
      RECT  125.0 9.4 126.6 9.6 ;
      RECT  127.4 5.4 129.4 6.0 ;
      RECT  128.6 4.0 129.4 5.4 ;
      RECT  137.2 17.6 138.4 21.6 ;
      RECT  129.0 6.6 129.8 7.4 ;
      RECT  133.4 13.6 134.0 14.8 ;
      RECT  130.6 12.0 131.4 12.2 ;
      RECT  137.0 10.8 137.8 11.0 ;
      RECT  133.0 17.0 133.6 17.6 ;
      RECT  127.4 14.2 132.8 14.8 ;
      RECT  133.0 4.0 133.8 6.0 ;
      RECT  123.0 22.2 144.8 23.4 ;
      RECT  128.6 18.2 129.4 21.6 ;
      RECT  140.2 13.6 141.0 22.2 ;
      RECT  124.2 12.6 129.8 12.8 ;
      RECT  126.4 11.2 127.2 11.4 ;
      RECT  134.6 3.4 135.4 6.0 ;
      RECT  137.2 4.0 138.4 5.4 ;
      RECT  123.0 2.2 144.8 3.4 ;
      RECT  143.4 20.6 144.2 22.2 ;
      RECT  125.0 9.6 136.0 10.2 ;
      RECT  138.8 8.4 142.6 9.0 ;
      RECT  127.4 6.0 128.2 6.8 ;
      RECT  133.0 6.0 133.6 6.6 ;
      RECT  137.0 6.0 137.8 6.8 ;
      RECT  138.4 12.2 139.2 12.4 ;
   LAYER  metal2 ;
      RECT  188.3 186.4 189.1 197.2 ;
      RECT  191.7 196.4 192.5 197.2 ;
      RECT  193.5 188.0 194.3 197.2 ;
      RECT  189.9 186.4 190.7 197.2 ;
      RECT  195.1 186.4 195.9 197.2 ;
      RECT  192.7 187.2 194.3 188.0 ;
      RECT  193.5 186.4 194.3 187.2 ;
      RECT  188.3 207.2 189.1 196.4 ;
      RECT  191.7 197.2 192.5 196.4 ;
      RECT  193.5 205.6 194.3 196.4 ;
      RECT  189.9 207.2 190.7 196.4 ;
      RECT  195.1 207.2 195.9 196.4 ;
      RECT  192.7 206.4 194.3 205.6 ;
      RECT  193.5 207.2 194.3 206.4 ;
      RECT  188.3 207.2 189.1 218.0 ;
      RECT  191.7 217.2 192.5 218.0 ;
      RECT  193.5 208.8 194.3 218.0 ;
      RECT  189.9 207.2 190.7 218.0 ;
      RECT  195.1 207.2 195.9 218.0 ;
      RECT  192.7 208.0 194.3 208.8 ;
      RECT  193.5 207.2 194.3 208.0 ;
      RECT  188.3 228.0 189.1 217.2 ;
      RECT  191.7 218.0 192.5 217.2 ;
      RECT  193.5 226.4 194.3 217.2 ;
      RECT  189.9 228.0 190.7 217.2 ;
      RECT  195.1 228.0 195.9 217.2 ;
      RECT  192.7 227.2 194.3 226.4 ;
      RECT  193.5 228.0 194.3 227.2 ;
      RECT  188.3 228.0 189.1 238.8 ;
      RECT  191.7 238.0 192.5 238.8 ;
      RECT  193.5 229.6 194.3 238.8 ;
      RECT  189.9 228.0 190.7 238.8 ;
      RECT  195.1 228.0 195.9 238.8 ;
      RECT  192.7 228.8 194.3 229.6 ;
      RECT  193.5 228.0 194.3 228.8 ;
      RECT  188.3 248.8 189.1 238.0 ;
      RECT  191.7 238.8 192.5 238.0 ;
      RECT  193.5 247.2 194.3 238.0 ;
      RECT  189.9 248.8 190.7 238.0 ;
      RECT  195.1 248.8 195.9 238.0 ;
      RECT  192.7 248.0 194.3 247.2 ;
      RECT  193.5 248.8 194.3 248.0 ;
      RECT  188.3 248.8 189.1 259.6 ;
      RECT  191.7 258.8 192.5 259.6 ;
      RECT  193.5 250.4 194.3 259.6 ;
      RECT  189.9 248.8 190.7 259.6 ;
      RECT  195.1 248.8 195.9 259.6 ;
      RECT  192.7 249.6 194.3 250.4 ;
      RECT  193.5 248.8 194.3 249.6 ;
      RECT  188.3 269.6 189.1 258.8 ;
      RECT  191.7 259.6 192.5 258.8 ;
      RECT  193.5 268.0 194.3 258.8 ;
      RECT  189.9 269.6 190.7 258.8 ;
      RECT  195.1 269.6 195.9 258.8 ;
      RECT  192.7 268.8 194.3 268.0 ;
      RECT  193.5 269.6 194.3 268.8 ;
      RECT  188.3 269.6 189.1 280.4 ;
      RECT  191.7 279.6 192.5 280.4 ;
      RECT  193.5 271.2 194.3 280.4 ;
      RECT  189.9 269.6 190.7 280.4 ;
      RECT  195.1 269.6 195.9 280.4 ;
      RECT  192.7 270.4 194.3 271.2 ;
      RECT  193.5 269.6 194.3 270.4 ;
      RECT  188.3 290.4 189.1 279.6 ;
      RECT  191.7 280.4 192.5 279.6 ;
      RECT  193.5 288.8 194.3 279.6 ;
      RECT  189.9 290.4 190.7 279.6 ;
      RECT  195.1 290.4 195.9 279.6 ;
      RECT  192.7 289.6 194.3 288.8 ;
      RECT  193.5 290.4 194.3 289.6 ;
      RECT  188.3 290.4 189.1 301.2 ;
      RECT  191.7 300.4 192.5 301.2 ;
      RECT  193.5 292.0 194.3 301.2 ;
      RECT  189.9 290.4 190.7 301.2 ;
      RECT  195.1 290.4 195.9 301.2 ;
      RECT  192.7 291.2 194.3 292.0 ;
      RECT  193.5 290.4 194.3 291.2 ;
      RECT  188.3 311.2 189.1 300.4 ;
      RECT  191.7 301.2 192.5 300.4 ;
      RECT  193.5 309.6 194.3 300.4 ;
      RECT  189.9 311.2 190.7 300.4 ;
      RECT  195.1 311.2 195.9 300.4 ;
      RECT  192.7 310.4 194.3 309.6 ;
      RECT  193.5 311.2 194.3 310.4 ;
      RECT  188.3 311.2 189.1 322.0 ;
      RECT  191.7 321.2 192.5 322.0 ;
      RECT  193.5 312.8 194.3 322.0 ;
      RECT  189.9 311.2 190.7 322.0 ;
      RECT  195.1 311.2 195.9 322.0 ;
      RECT  192.7 312.0 194.3 312.8 ;
      RECT  193.5 311.2 194.3 312.0 ;
      RECT  188.3 332.0 189.1 321.2 ;
      RECT  191.7 322.0 192.5 321.2 ;
      RECT  193.5 330.4 194.3 321.2 ;
      RECT  189.9 332.0 190.7 321.2 ;
      RECT  195.1 332.0 195.9 321.2 ;
      RECT  192.7 331.2 194.3 330.4 ;
      RECT  193.5 332.0 194.3 331.2 ;
      RECT  188.3 332.0 189.1 342.8 ;
      RECT  191.7 342.0 192.5 342.8 ;
      RECT  193.5 333.6 194.3 342.8 ;
      RECT  189.9 332.0 190.7 342.8 ;
      RECT  195.1 332.0 195.9 342.8 ;
      RECT  192.7 332.8 194.3 333.6 ;
      RECT  193.5 332.0 194.3 332.8 ;
      RECT  188.3 352.8 189.1 342.0 ;
      RECT  191.7 342.8 192.5 342.0 ;
      RECT  193.5 351.2 194.3 342.0 ;
      RECT  189.9 352.8 190.7 342.0 ;
      RECT  195.1 352.8 195.9 342.0 ;
      RECT  192.7 352.0 194.3 351.2 ;
      RECT  193.5 352.8 194.3 352.0 ;
      RECT  195.1 186.4 195.9 197.2 ;
      RECT  198.5 196.4 199.3 197.2 ;
      RECT  200.3 188.0 201.1 197.2 ;
      RECT  196.7 186.4 197.5 197.2 ;
      RECT  201.9 186.4 202.7 197.2 ;
      RECT  199.5 187.2 201.1 188.0 ;
      RECT  200.3 186.4 201.1 187.2 ;
      RECT  195.1 207.2 195.9 196.4 ;
      RECT  198.5 197.2 199.3 196.4 ;
      RECT  200.3 205.6 201.1 196.4 ;
      RECT  196.7 207.2 197.5 196.4 ;
      RECT  201.9 207.2 202.7 196.4 ;
      RECT  199.5 206.4 201.1 205.6 ;
      RECT  200.3 207.2 201.1 206.4 ;
      RECT  195.1 207.2 195.9 218.0 ;
      RECT  198.5 217.2 199.3 218.0 ;
      RECT  200.3 208.8 201.1 218.0 ;
      RECT  196.7 207.2 197.5 218.0 ;
      RECT  201.9 207.2 202.7 218.0 ;
      RECT  199.5 208.0 201.1 208.8 ;
      RECT  200.3 207.2 201.1 208.0 ;
      RECT  195.1 228.0 195.9 217.2 ;
      RECT  198.5 218.0 199.3 217.2 ;
      RECT  200.3 226.4 201.1 217.2 ;
      RECT  196.7 228.0 197.5 217.2 ;
      RECT  201.9 228.0 202.7 217.2 ;
      RECT  199.5 227.2 201.1 226.4 ;
      RECT  200.3 228.0 201.1 227.2 ;
      RECT  195.1 228.0 195.9 238.8 ;
      RECT  198.5 238.0 199.3 238.8 ;
      RECT  200.3 229.6 201.1 238.8 ;
      RECT  196.7 228.0 197.5 238.8 ;
      RECT  201.9 228.0 202.7 238.8 ;
      RECT  199.5 228.8 201.1 229.6 ;
      RECT  200.3 228.0 201.1 228.8 ;
      RECT  195.1 248.8 195.9 238.0 ;
      RECT  198.5 238.8 199.3 238.0 ;
      RECT  200.3 247.2 201.1 238.0 ;
      RECT  196.7 248.8 197.5 238.0 ;
      RECT  201.9 248.8 202.7 238.0 ;
      RECT  199.5 248.0 201.1 247.2 ;
      RECT  200.3 248.8 201.1 248.0 ;
      RECT  195.1 248.8 195.9 259.6 ;
      RECT  198.5 258.8 199.3 259.6 ;
      RECT  200.3 250.4 201.1 259.6 ;
      RECT  196.7 248.8 197.5 259.6 ;
      RECT  201.9 248.8 202.7 259.6 ;
      RECT  199.5 249.6 201.1 250.4 ;
      RECT  200.3 248.8 201.1 249.6 ;
      RECT  195.1 269.6 195.9 258.8 ;
      RECT  198.5 259.6 199.3 258.8 ;
      RECT  200.3 268.0 201.1 258.8 ;
      RECT  196.7 269.6 197.5 258.8 ;
      RECT  201.9 269.6 202.7 258.8 ;
      RECT  199.5 268.8 201.1 268.0 ;
      RECT  200.3 269.6 201.1 268.8 ;
      RECT  195.1 269.6 195.9 280.4 ;
      RECT  198.5 279.6 199.3 280.4 ;
      RECT  200.3 271.2 201.1 280.4 ;
      RECT  196.7 269.6 197.5 280.4 ;
      RECT  201.9 269.6 202.7 280.4 ;
      RECT  199.5 270.4 201.1 271.2 ;
      RECT  200.3 269.6 201.1 270.4 ;
      RECT  195.1 290.4 195.9 279.6 ;
      RECT  198.5 280.4 199.3 279.6 ;
      RECT  200.3 288.8 201.1 279.6 ;
      RECT  196.7 290.4 197.5 279.6 ;
      RECT  201.9 290.4 202.7 279.6 ;
      RECT  199.5 289.6 201.1 288.8 ;
      RECT  200.3 290.4 201.1 289.6 ;
      RECT  195.1 290.4 195.9 301.2 ;
      RECT  198.5 300.4 199.3 301.2 ;
      RECT  200.3 292.0 201.1 301.2 ;
      RECT  196.7 290.4 197.5 301.2 ;
      RECT  201.9 290.4 202.7 301.2 ;
      RECT  199.5 291.2 201.1 292.0 ;
      RECT  200.3 290.4 201.1 291.2 ;
      RECT  195.1 311.2 195.9 300.4 ;
      RECT  198.5 301.2 199.3 300.4 ;
      RECT  200.3 309.6 201.1 300.4 ;
      RECT  196.7 311.2 197.5 300.4 ;
      RECT  201.9 311.2 202.7 300.4 ;
      RECT  199.5 310.4 201.1 309.6 ;
      RECT  200.3 311.2 201.1 310.4 ;
      RECT  195.1 311.2 195.9 322.0 ;
      RECT  198.5 321.2 199.3 322.0 ;
      RECT  200.3 312.8 201.1 322.0 ;
      RECT  196.7 311.2 197.5 322.0 ;
      RECT  201.9 311.2 202.7 322.0 ;
      RECT  199.5 312.0 201.1 312.8 ;
      RECT  200.3 311.2 201.1 312.0 ;
      RECT  195.1 332.0 195.9 321.2 ;
      RECT  198.5 322.0 199.3 321.2 ;
      RECT  200.3 330.4 201.1 321.2 ;
      RECT  196.7 332.0 197.5 321.2 ;
      RECT  201.9 332.0 202.7 321.2 ;
      RECT  199.5 331.2 201.1 330.4 ;
      RECT  200.3 332.0 201.1 331.2 ;
      RECT  195.1 332.0 195.9 342.8 ;
      RECT  198.5 342.0 199.3 342.8 ;
      RECT  200.3 333.6 201.1 342.8 ;
      RECT  196.7 332.0 197.5 342.8 ;
      RECT  201.9 332.0 202.7 342.8 ;
      RECT  199.5 332.8 201.1 333.6 ;
      RECT  200.3 332.0 201.1 332.8 ;
      RECT  195.1 352.8 195.9 342.0 ;
      RECT  198.5 342.8 199.3 342.0 ;
      RECT  200.3 351.2 201.1 342.0 ;
      RECT  196.7 352.8 197.5 342.0 ;
      RECT  201.9 352.8 202.7 342.0 ;
      RECT  199.5 352.0 201.1 351.2 ;
      RECT  200.3 352.8 201.1 352.0 ;
      RECT  189.9 186.4 190.7 352.8 ;
      RECT  193.5 186.4 194.3 352.8 ;
      RECT  196.7 186.4 197.5 352.8 ;
      RECT  200.3 186.4 201.1 352.8 ;
      RECT  198.5 196.4 199.3 197.2 ;
      RECT  191.7 217.2 192.5 218.0 ;
      RECT  191.7 279.6 192.5 280.4 ;
      RECT  191.7 321.2 192.5 322.0 ;
      RECT  191.7 321.2 192.5 322.0 ;
      RECT  191.7 342.0 192.5 342.8 ;
      RECT  198.5 300.4 199.3 301.2 ;
      RECT  198.5 300.4 199.3 301.2 ;
      RECT  191.7 300.4 192.5 301.2 ;
      RECT  191.7 300.4 192.5 301.2 ;
      RECT  191.7 238.0 192.5 238.8 ;
      RECT  191.7 238.0 192.5 238.8 ;
      RECT  198.5 279.6 199.3 280.4 ;
      RECT  198.5 258.8 199.3 259.6 ;
      RECT  198.5 321.2 199.3 322.0 ;
      RECT  198.5 321.2 199.3 322.0 ;
      RECT  191.7 258.8 192.5 259.6 ;
      RECT  198.5 342.0 199.3 342.8 ;
      RECT  198.5 238.0 199.3 238.8 ;
      RECT  198.5 238.0 199.3 238.8 ;
      RECT  198.5 217.2 199.3 218.0 ;
      RECT  191.7 196.4 192.5 197.2 ;
      RECT  188.3 300.4 189.1 311.2 ;
      RECT  201.9 217.2 202.7 228.0 ;
      RECT  195.1 217.2 195.9 228.0 ;
      RECT  195.1 217.2 195.9 228.0 ;
      RECT  201.9 186.4 202.7 197.2 ;
      RECT  188.3 248.8 189.1 259.6 ;
      RECT  195.1 300.4 195.9 311.2 ;
      RECT  195.1 300.4 195.9 311.2 ;
      RECT  195.1 342.0 195.9 352.8 ;
      RECT  195.1 342.0 195.9 352.8 ;
      RECT  201.9 279.6 202.7 290.4 ;
      RECT  195.1 290.4 195.9 301.2 ;
      RECT  195.1 290.4 195.9 301.2 ;
      RECT  195.1 196.4 195.9 207.2 ;
      RECT  195.1 196.4 195.9 207.2 ;
      RECT  195.1 238.0 195.9 248.8 ;
      RECT  201.9 228.0 202.7 238.8 ;
      RECT  195.1 238.0 195.9 248.8 ;
      RECT  195.1 269.6 195.9 280.4 ;
      RECT  195.1 269.6 195.9 280.4 ;
      RECT  195.1 279.6 195.9 290.4 ;
      RECT  195.1 279.6 195.9 290.4 ;
      RECT  188.3 321.2 189.1 332.0 ;
      RECT  188.3 332.0 189.1 342.8 ;
      RECT  201.9 196.4 202.7 207.2 ;
      RECT  188.3 228.0 189.1 238.8 ;
      RECT  188.3 196.4 189.1 207.2 ;
      RECT  195.1 248.8 195.9 259.6 ;
      RECT  201.9 238.0 202.7 248.8 ;
      RECT  195.1 248.8 195.9 259.6 ;
      RECT  188.3 311.2 189.1 322.0 ;
      RECT  195.1 311.2 195.9 322.0 ;
      RECT  195.1 311.2 195.9 322.0 ;
      RECT  201.9 332.0 202.7 342.8 ;
      RECT  201.9 342.0 202.7 352.8 ;
      RECT  188.3 217.2 189.1 228.0 ;
      RECT  195.1 258.8 195.9 269.6 ;
      RECT  188.3 207.2 189.1 218.0 ;
      RECT  201.9 248.8 202.7 259.6 ;
      RECT  195.1 258.8 195.9 269.6 ;
      RECT  188.3 238.0 189.1 248.8 ;
      RECT  201.9 311.2 202.7 322.0 ;
      RECT  188.3 258.8 189.1 269.6 ;
      RECT  195.1 186.4 195.9 197.2 ;
      RECT  195.1 186.4 195.9 197.2 ;
      RECT  188.3 269.6 189.1 280.4 ;
      RECT  201.9 207.2 202.7 218.0 ;
      RECT  188.3 342.0 189.1 352.8 ;
      RECT  201.9 258.8 202.7 269.6 ;
      RECT  195.1 332.0 195.9 342.8 ;
      RECT  195.1 321.2 195.9 332.0 ;
      RECT  195.1 228.0 195.9 238.8 ;
      RECT  195.1 228.0 195.9 238.8 ;
      RECT  188.3 279.6 189.1 290.4 ;
      RECT  188.3 290.4 189.1 301.2 ;
      RECT  195.1 321.2 195.9 332.0 ;
      RECT  195.1 207.2 195.9 218.0 ;
      RECT  195.1 207.2 195.9 218.0 ;
      RECT  201.9 321.2 202.7 332.0 ;
      RECT  201.9 290.4 202.7 301.2 ;
      RECT  201.9 300.4 202.7 311.2 ;
      RECT  195.1 332.0 195.9 342.8 ;
      RECT  201.9 269.6 202.7 280.4 ;
      RECT  188.3 186.4 189.1 197.2 ;
      RECT  188.3 165.6 189.1 176.4 ;
      RECT  181.5 165.6 182.3 176.4 ;
      RECT  184.9 175.6 185.7 176.4 ;
      RECT  186.7 165.6 187.5 176.4 ;
      RECT  183.1 165.6 183.9 176.4 ;
      RECT  181.5 186.4 182.3 175.6 ;
      RECT  184.9 176.4 185.7 175.6 ;
      RECT  186.7 184.8 187.5 175.6 ;
      RECT  183.1 186.4 183.9 175.6 ;
      RECT  188.3 186.4 189.1 175.6 ;
      RECT  185.9 185.6 187.5 184.8 ;
      RECT  186.7 186.4 187.5 185.6 ;
      RECT  181.5 186.4 182.3 197.2 ;
      RECT  184.9 196.4 185.7 197.2 ;
      RECT  186.7 188.0 187.5 197.2 ;
      RECT  183.1 186.4 183.9 197.2 ;
      RECT  188.3 186.4 189.1 197.2 ;
      RECT  185.9 187.2 187.5 188.0 ;
      RECT  186.7 186.4 187.5 187.2 ;
      RECT  181.5 207.2 182.3 196.4 ;
      RECT  184.9 197.2 185.7 196.4 ;
      RECT  186.7 205.6 187.5 196.4 ;
      RECT  183.1 207.2 183.9 196.4 ;
      RECT  188.3 207.2 189.1 196.4 ;
      RECT  185.9 206.4 187.5 205.6 ;
      RECT  186.7 207.2 187.5 206.4 ;
      RECT  181.5 207.2 182.3 218.0 ;
      RECT  184.9 217.2 185.7 218.0 ;
      RECT  186.7 208.8 187.5 218.0 ;
      RECT  183.1 207.2 183.9 218.0 ;
      RECT  188.3 207.2 189.1 218.0 ;
      RECT  185.9 208.0 187.5 208.8 ;
      RECT  186.7 207.2 187.5 208.0 ;
      RECT  181.5 228.0 182.3 217.2 ;
      RECT  184.9 218.0 185.7 217.2 ;
      RECT  186.7 226.4 187.5 217.2 ;
      RECT  183.1 228.0 183.9 217.2 ;
      RECT  188.3 228.0 189.1 217.2 ;
      RECT  185.9 227.2 187.5 226.4 ;
      RECT  186.7 228.0 187.5 227.2 ;
      RECT  181.5 228.0 182.3 238.8 ;
      RECT  184.9 238.0 185.7 238.8 ;
      RECT  186.7 229.6 187.5 238.8 ;
      RECT  183.1 228.0 183.9 238.8 ;
      RECT  188.3 228.0 189.1 238.8 ;
      RECT  185.9 228.8 187.5 229.6 ;
      RECT  186.7 228.0 187.5 228.8 ;
      RECT  181.5 248.8 182.3 238.0 ;
      RECT  184.9 238.8 185.7 238.0 ;
      RECT  186.7 247.2 187.5 238.0 ;
      RECT  183.1 248.8 183.9 238.0 ;
      RECT  188.3 248.8 189.1 238.0 ;
      RECT  185.9 248.0 187.5 247.2 ;
      RECT  186.7 248.8 187.5 248.0 ;
      RECT  181.5 248.8 182.3 259.6 ;
      RECT  184.9 258.8 185.7 259.6 ;
      RECT  186.7 250.4 187.5 259.6 ;
      RECT  183.1 248.8 183.9 259.6 ;
      RECT  188.3 248.8 189.1 259.6 ;
      RECT  185.9 249.6 187.5 250.4 ;
      RECT  186.7 248.8 187.5 249.6 ;
      RECT  181.5 269.6 182.3 258.8 ;
      RECT  184.9 259.6 185.7 258.8 ;
      RECT  186.7 268.0 187.5 258.8 ;
      RECT  183.1 269.6 183.9 258.8 ;
      RECT  188.3 269.6 189.1 258.8 ;
      RECT  185.9 268.8 187.5 268.0 ;
      RECT  186.7 269.6 187.5 268.8 ;
      RECT  181.5 269.6 182.3 280.4 ;
      RECT  184.9 279.6 185.7 280.4 ;
      RECT  186.7 271.2 187.5 280.4 ;
      RECT  183.1 269.6 183.9 280.4 ;
      RECT  188.3 269.6 189.1 280.4 ;
      RECT  185.9 270.4 187.5 271.2 ;
      RECT  186.7 269.6 187.5 270.4 ;
      RECT  181.5 290.4 182.3 279.6 ;
      RECT  184.9 280.4 185.7 279.6 ;
      RECT  186.7 288.8 187.5 279.6 ;
      RECT  183.1 290.4 183.9 279.6 ;
      RECT  188.3 290.4 189.1 279.6 ;
      RECT  185.9 289.6 187.5 288.8 ;
      RECT  186.7 290.4 187.5 289.6 ;
      RECT  181.5 290.4 182.3 301.2 ;
      RECT  184.9 300.4 185.7 301.2 ;
      RECT  186.7 292.0 187.5 301.2 ;
      RECT  183.1 290.4 183.9 301.2 ;
      RECT  188.3 290.4 189.1 301.2 ;
      RECT  185.9 291.2 187.5 292.0 ;
      RECT  186.7 290.4 187.5 291.2 ;
      RECT  181.5 311.2 182.3 300.4 ;
      RECT  184.9 301.2 185.7 300.4 ;
      RECT  186.7 309.6 187.5 300.4 ;
      RECT  183.1 311.2 183.9 300.4 ;
      RECT  188.3 311.2 189.1 300.4 ;
      RECT  185.9 310.4 187.5 309.6 ;
      RECT  186.7 311.2 187.5 310.4 ;
      RECT  181.5 311.2 182.3 322.0 ;
      RECT  184.9 321.2 185.7 322.0 ;
      RECT  186.7 312.8 187.5 322.0 ;
      RECT  183.1 311.2 183.9 322.0 ;
      RECT  188.3 311.2 189.1 322.0 ;
      RECT  185.9 312.0 187.5 312.8 ;
      RECT  186.7 311.2 187.5 312.0 ;
      RECT  181.5 332.0 182.3 321.2 ;
      RECT  184.9 322.0 185.7 321.2 ;
      RECT  186.7 330.4 187.5 321.2 ;
      RECT  183.1 332.0 183.9 321.2 ;
      RECT  188.3 332.0 189.1 321.2 ;
      RECT  185.9 331.2 187.5 330.4 ;
      RECT  186.7 332.0 187.5 331.2 ;
      RECT  181.5 332.0 182.3 342.8 ;
      RECT  184.9 342.0 185.7 342.8 ;
      RECT  186.7 333.6 187.5 342.8 ;
      RECT  183.1 332.0 183.9 342.8 ;
      RECT  188.3 332.0 189.1 342.8 ;
      RECT  185.9 332.8 187.5 333.6 ;
      RECT  186.7 332.0 187.5 332.8 ;
      RECT  181.5 352.8 182.3 342.0 ;
      RECT  184.9 342.8 185.7 342.0 ;
      RECT  186.7 351.2 187.5 342.0 ;
      RECT  183.1 352.8 183.9 342.0 ;
      RECT  188.3 352.8 189.1 342.0 ;
      RECT  185.9 352.0 187.5 351.2 ;
      RECT  186.7 352.8 187.5 352.0 ;
      RECT  188.3 352.8 189.1 363.6 ;
      RECT  181.5 352.8 182.3 363.6 ;
      RECT  184.9 362.8 185.7 363.6 ;
      RECT  186.7 352.8 187.5 363.6 ;
      RECT  183.1 352.8 183.9 363.6 ;
      RECT  183.1 165.6 183.9 363.2 ;
      RECT  186.7 165.6 187.5 363.2 ;
      RECT  184.9 279.6 185.7 280.4 ;
      RECT  184.9 279.6 185.7 280.4 ;
      RECT  184.9 217.2 185.7 218.0 ;
      RECT  184.9 217.2 185.7 218.0 ;
      RECT  184.9 342.0 185.7 342.8 ;
      RECT  184.9 300.4 185.7 301.2 ;
      RECT  184.9 300.4 185.7 301.2 ;
      RECT  184.9 175.6 185.7 176.4 ;
      RECT  184.9 196.4 185.7 197.2 ;
      RECT  184.9 321.2 185.7 322.0 ;
      RECT  184.9 238.0 185.7 238.8 ;
      RECT  184.9 258.8 185.7 259.6 ;
      RECT  181.5 279.6 182.3 290.4 ;
      RECT  181.5 332.0 182.3 342.8 ;
      RECT  188.3 196.4 189.1 207.2 ;
      RECT  181.5 228.0 182.3 238.8 ;
      RECT  188.3 279.6 189.1 290.4 ;
      RECT  188.3 321.2 189.1 332.0 ;
      RECT  188.3 269.6 189.1 280.4 ;
      RECT  188.3 175.6 189.1 186.4 ;
      RECT  188.3 217.2 189.1 228.0 ;
      RECT  188.3 248.8 189.1 259.6 ;
      RECT  181.5 300.4 182.3 311.2 ;
      RECT  188.3 258.8 189.1 269.6 ;
      RECT  181.5 311.2 182.3 322.0 ;
      RECT  181.5 207.2 182.3 218.0 ;
      RECT  181.5 175.6 182.3 186.4 ;
      RECT  188.3 228.0 189.1 238.8 ;
      RECT  181.5 342.0 182.3 352.8 ;
      RECT  181.5 290.4 182.3 301.2 ;
      RECT  188.3 290.4 189.1 301.2 ;
      RECT  188.3 342.0 189.1 352.8 ;
      RECT  181.5 196.4 182.3 207.2 ;
      RECT  188.3 238.0 189.1 248.8 ;
      RECT  181.5 186.4 182.3 197.2 ;
      RECT  188.3 332.0 189.1 342.8 ;
      RECT  181.5 217.2 182.3 228.0 ;
      RECT  181.5 238.0 182.3 248.8 ;
      RECT  181.5 248.8 182.3 259.6 ;
      RECT  181.5 321.2 182.3 332.0 ;
      RECT  188.3 300.4 189.1 311.2 ;
      RECT  188.3 207.2 189.1 218.0 ;
      RECT  181.5 258.8 182.3 269.6 ;
      RECT  181.5 269.6 182.3 280.4 ;
      RECT  188.3 186.4 189.1 197.2 ;
      RECT  188.3 311.2 189.1 322.0 ;
      RECT  195.1 186.4 195.9 175.6 ;
      RECT  188.3 186.4 189.1 175.6 ;
      RECT  191.7 176.4 192.5 175.6 ;
      RECT  193.5 186.4 194.3 175.6 ;
      RECT  189.9 186.4 190.7 175.6 ;
      RECT  201.9 186.4 202.7 175.6 ;
      RECT  195.1 186.4 195.9 175.6 ;
      RECT  198.5 176.4 199.3 175.6 ;
      RECT  200.3 186.4 201.1 175.6 ;
      RECT  196.7 186.4 197.5 175.6 ;
      RECT  191.7 176.4 192.5 175.6 ;
      RECT  198.5 176.4 199.3 175.6 ;
      RECT  195.1 186.4 195.9 175.6 ;
      RECT  201.9 186.4 202.7 175.6 ;
      RECT  195.1 186.4 195.9 175.6 ;
      RECT  188.3 186.4 189.1 175.6 ;
      RECT  195.1 165.6 195.9 176.4 ;
      RECT  188.3 165.6 189.1 176.4 ;
      RECT  191.7 175.6 192.5 176.4 ;
      RECT  193.5 165.6 194.3 176.4 ;
      RECT  189.9 165.6 190.7 176.4 ;
      RECT  201.9 165.6 202.7 176.4 ;
      RECT  195.1 165.6 195.9 176.4 ;
      RECT  198.5 175.6 199.3 176.4 ;
      RECT  200.3 165.6 201.1 176.4 ;
      RECT  196.7 165.6 197.5 176.4 ;
      RECT  191.7 175.6 192.5 176.4 ;
      RECT  198.5 175.6 199.3 176.4 ;
      RECT  195.1 165.6 195.9 176.4 ;
      RECT  201.9 165.6 202.7 176.4 ;
      RECT  195.1 165.6 195.9 176.4 ;
      RECT  188.3 165.6 189.1 176.4 ;
      RECT  195.1 352.8 195.9 363.6 ;
      RECT  188.3 352.8 189.1 363.6 ;
      RECT  191.7 362.8 192.5 363.6 ;
      RECT  193.5 352.8 194.3 363.6 ;
      RECT  189.9 352.8 190.7 363.6 ;
      RECT  201.9 352.8 202.7 363.6 ;
      RECT  195.1 352.8 195.9 363.6 ;
      RECT  198.5 362.8 199.3 363.6 ;
      RECT  200.3 352.8 201.1 363.6 ;
      RECT  196.7 352.8 197.5 363.6 ;
      RECT  191.7 362.8 192.5 363.6 ;
      RECT  198.5 362.8 199.3 363.6 ;
      RECT  195.1 352.8 195.9 363.6 ;
      RECT  201.9 352.8 202.7 363.6 ;
      RECT  195.1 352.8 195.9 363.6 ;
      RECT  188.3 352.8 189.1 363.6 ;
      RECT  181.5 165.6 182.3 176.4 ;
      RECT  174.7 165.6 175.5 176.4 ;
      RECT  178.1 175.6 178.9 176.4 ;
      RECT  179.9 165.6 180.7 176.4 ;
      RECT  176.3 165.6 177.1 176.4 ;
      RECT  181.5 186.4 182.3 175.6 ;
      RECT  174.7 186.4 175.5 175.6 ;
      RECT  178.1 176.4 178.9 175.6 ;
      RECT  179.9 186.4 180.7 175.6 ;
      RECT  176.3 186.4 177.1 175.6 ;
      RECT  181.5 186.4 182.3 197.2 ;
      RECT  174.7 186.4 175.5 197.2 ;
      RECT  178.1 196.4 178.9 197.2 ;
      RECT  179.9 186.4 180.7 197.2 ;
      RECT  176.3 186.4 177.1 197.2 ;
      RECT  181.5 207.2 182.3 196.4 ;
      RECT  174.7 207.2 175.5 196.4 ;
      RECT  178.1 197.2 178.9 196.4 ;
      RECT  179.9 207.2 180.7 196.4 ;
      RECT  176.3 207.2 177.1 196.4 ;
      RECT  181.5 207.2 182.3 218.0 ;
      RECT  174.7 207.2 175.5 218.0 ;
      RECT  178.1 217.2 178.9 218.0 ;
      RECT  179.9 207.2 180.7 218.0 ;
      RECT  176.3 207.2 177.1 218.0 ;
      RECT  181.5 228.0 182.3 217.2 ;
      RECT  174.7 228.0 175.5 217.2 ;
      RECT  178.1 218.0 178.9 217.2 ;
      RECT  179.9 228.0 180.7 217.2 ;
      RECT  176.3 228.0 177.1 217.2 ;
      RECT  181.5 228.0 182.3 238.8 ;
      RECT  174.7 228.0 175.5 238.8 ;
      RECT  178.1 238.0 178.9 238.8 ;
      RECT  179.9 228.0 180.7 238.8 ;
      RECT  176.3 228.0 177.1 238.8 ;
      RECT  181.5 248.8 182.3 238.0 ;
      RECT  174.7 248.8 175.5 238.0 ;
      RECT  178.1 238.8 178.9 238.0 ;
      RECT  179.9 248.8 180.7 238.0 ;
      RECT  176.3 248.8 177.1 238.0 ;
      RECT  181.5 248.8 182.3 259.6 ;
      RECT  174.7 248.8 175.5 259.6 ;
      RECT  178.1 258.8 178.9 259.6 ;
      RECT  179.9 248.8 180.7 259.6 ;
      RECT  176.3 248.8 177.1 259.6 ;
      RECT  181.5 269.6 182.3 258.8 ;
      RECT  174.7 269.6 175.5 258.8 ;
      RECT  178.1 259.6 178.9 258.8 ;
      RECT  179.9 269.6 180.7 258.8 ;
      RECT  176.3 269.6 177.1 258.8 ;
      RECT  181.5 269.6 182.3 280.4 ;
      RECT  174.7 269.6 175.5 280.4 ;
      RECT  178.1 279.6 178.9 280.4 ;
      RECT  179.9 269.6 180.7 280.4 ;
      RECT  176.3 269.6 177.1 280.4 ;
      RECT  181.5 290.4 182.3 279.6 ;
      RECT  174.7 290.4 175.5 279.6 ;
      RECT  178.1 280.4 178.9 279.6 ;
      RECT  179.9 290.4 180.7 279.6 ;
      RECT  176.3 290.4 177.1 279.6 ;
      RECT  181.5 290.4 182.3 301.2 ;
      RECT  174.7 290.4 175.5 301.2 ;
      RECT  178.1 300.4 178.9 301.2 ;
      RECT  179.9 290.4 180.7 301.2 ;
      RECT  176.3 290.4 177.1 301.2 ;
      RECT  181.5 311.2 182.3 300.4 ;
      RECT  174.7 311.2 175.5 300.4 ;
      RECT  178.1 301.2 178.9 300.4 ;
      RECT  179.9 311.2 180.7 300.4 ;
      RECT  176.3 311.2 177.1 300.4 ;
      RECT  181.5 311.2 182.3 322.0 ;
      RECT  174.7 311.2 175.5 322.0 ;
      RECT  178.1 321.2 178.9 322.0 ;
      RECT  179.9 311.2 180.7 322.0 ;
      RECT  176.3 311.2 177.1 322.0 ;
      RECT  181.5 332.0 182.3 321.2 ;
      RECT  174.7 332.0 175.5 321.2 ;
      RECT  178.1 322.0 178.9 321.2 ;
      RECT  179.9 332.0 180.7 321.2 ;
      RECT  176.3 332.0 177.1 321.2 ;
      RECT  181.5 332.0 182.3 342.8 ;
      RECT  174.7 332.0 175.5 342.8 ;
      RECT  178.1 342.0 178.9 342.8 ;
      RECT  179.9 332.0 180.7 342.8 ;
      RECT  176.3 332.0 177.1 342.8 ;
      RECT  181.5 352.8 182.3 342.0 ;
      RECT  174.7 352.8 175.5 342.0 ;
      RECT  178.1 342.8 178.9 342.0 ;
      RECT  179.9 352.8 180.7 342.0 ;
      RECT  176.3 352.8 177.1 342.0 ;
      RECT  181.5 352.8 182.3 363.6 ;
      RECT  174.7 352.8 175.5 363.6 ;
      RECT  178.1 362.8 178.9 363.6 ;
      RECT  179.9 352.8 180.7 363.6 ;
      RECT  176.3 352.8 177.1 363.6 ;
      RECT  178.1 279.6 178.9 280.4 ;
      RECT  178.1 279.6 178.9 280.4 ;
      RECT  178.1 217.2 178.9 218.0 ;
      RECT  178.1 217.2 178.9 218.0 ;
      RECT  178.1 342.0 178.9 342.8 ;
      RECT  178.1 300.4 178.9 301.2 ;
      RECT  178.1 300.4 178.9 301.2 ;
      RECT  178.1 362.8 178.9 363.6 ;
      RECT  178.1 175.6 178.9 176.4 ;
      RECT  178.1 196.4 178.9 197.2 ;
      RECT  178.1 321.2 178.9 322.0 ;
      RECT  178.1 238.0 178.9 238.8 ;
      RECT  178.1 258.8 178.9 259.6 ;
      RECT  174.7 279.6 175.5 290.4 ;
      RECT  174.7 332.0 175.5 342.8 ;
      RECT  181.5 196.4 182.3 207.2 ;
      RECT  174.7 228.0 175.5 238.8 ;
      RECT  181.5 279.6 182.3 290.4 ;
      RECT  181.5 321.2 182.3 332.0 ;
      RECT  181.5 269.6 182.3 280.4 ;
      RECT  181.5 175.6 182.3 186.4 ;
      RECT  181.5 217.2 182.3 228.0 ;
      RECT  181.5 248.8 182.3 259.6 ;
      RECT  174.7 300.4 175.5 311.2 ;
      RECT  181.5 258.8 182.3 269.6 ;
      RECT  174.7 311.2 175.5 322.0 ;
      RECT  174.7 207.2 175.5 218.0 ;
      RECT  174.7 175.6 175.5 186.4 ;
      RECT  181.5 228.0 182.3 238.8 ;
      RECT  174.7 342.0 175.5 352.8 ;
      RECT  174.7 352.8 175.5 363.6 ;
      RECT  174.7 290.4 175.5 301.2 ;
      RECT  181.5 290.4 182.3 301.2 ;
      RECT  181.5 342.0 182.3 352.8 ;
      RECT  174.7 196.4 175.5 207.2 ;
      RECT  181.5 238.0 182.3 248.8 ;
      RECT  174.7 186.4 175.5 197.2 ;
      RECT  181.5 332.0 182.3 342.8 ;
      RECT  181.5 352.8 182.3 363.6 ;
      RECT  174.7 217.2 175.5 228.0 ;
      RECT  174.7 238.0 175.5 248.8 ;
      RECT  181.5 165.6 182.3 176.4 ;
      RECT  174.7 248.8 175.5 259.6 ;
      RECT  174.7 321.2 175.5 332.0 ;
      RECT  181.5 300.4 182.3 311.2 ;
      RECT  181.5 207.2 182.3 218.0 ;
      RECT  174.7 258.8 175.5 269.6 ;
      RECT  174.7 269.6 175.5 280.4 ;
      RECT  181.5 186.4 182.3 197.2 ;
      RECT  181.5 311.2 182.3 322.0 ;
      RECT  174.7 165.6 175.5 176.4 ;
      RECT  208.7 165.6 209.5 176.4 ;
      RECT  201.9 165.6 202.7 176.4 ;
      RECT  205.3 175.6 206.1 176.4 ;
      RECT  207.1 165.6 207.9 176.4 ;
      RECT  203.5 165.6 204.3 176.4 ;
      RECT  208.7 186.4 209.5 175.6 ;
      RECT  201.9 186.4 202.7 175.6 ;
      RECT  205.3 176.4 206.1 175.6 ;
      RECT  207.1 186.4 207.9 175.6 ;
      RECT  203.5 186.4 204.3 175.6 ;
      RECT  208.7 186.4 209.5 197.2 ;
      RECT  201.9 186.4 202.7 197.2 ;
      RECT  205.3 196.4 206.1 197.2 ;
      RECT  207.1 186.4 207.9 197.2 ;
      RECT  203.5 186.4 204.3 197.2 ;
      RECT  208.7 207.2 209.5 196.4 ;
      RECT  201.9 207.2 202.7 196.4 ;
      RECT  205.3 197.2 206.1 196.4 ;
      RECT  207.1 207.2 207.9 196.4 ;
      RECT  203.5 207.2 204.3 196.4 ;
      RECT  208.7 207.2 209.5 218.0 ;
      RECT  201.9 207.2 202.7 218.0 ;
      RECT  205.3 217.2 206.1 218.0 ;
      RECT  207.1 207.2 207.9 218.0 ;
      RECT  203.5 207.2 204.3 218.0 ;
      RECT  208.7 228.0 209.5 217.2 ;
      RECT  201.9 228.0 202.7 217.2 ;
      RECT  205.3 218.0 206.1 217.2 ;
      RECT  207.1 228.0 207.9 217.2 ;
      RECT  203.5 228.0 204.3 217.2 ;
      RECT  208.7 228.0 209.5 238.8 ;
      RECT  201.9 228.0 202.7 238.8 ;
      RECT  205.3 238.0 206.1 238.8 ;
      RECT  207.1 228.0 207.9 238.8 ;
      RECT  203.5 228.0 204.3 238.8 ;
      RECT  208.7 248.8 209.5 238.0 ;
      RECT  201.9 248.8 202.7 238.0 ;
      RECT  205.3 238.8 206.1 238.0 ;
      RECT  207.1 248.8 207.9 238.0 ;
      RECT  203.5 248.8 204.3 238.0 ;
      RECT  208.7 248.8 209.5 259.6 ;
      RECT  201.9 248.8 202.7 259.6 ;
      RECT  205.3 258.8 206.1 259.6 ;
      RECT  207.1 248.8 207.9 259.6 ;
      RECT  203.5 248.8 204.3 259.6 ;
      RECT  208.7 269.6 209.5 258.8 ;
      RECT  201.9 269.6 202.7 258.8 ;
      RECT  205.3 259.6 206.1 258.8 ;
      RECT  207.1 269.6 207.9 258.8 ;
      RECT  203.5 269.6 204.3 258.8 ;
      RECT  208.7 269.6 209.5 280.4 ;
      RECT  201.9 269.6 202.7 280.4 ;
      RECT  205.3 279.6 206.1 280.4 ;
      RECT  207.1 269.6 207.9 280.4 ;
      RECT  203.5 269.6 204.3 280.4 ;
      RECT  208.7 290.4 209.5 279.6 ;
      RECT  201.9 290.4 202.7 279.6 ;
      RECT  205.3 280.4 206.1 279.6 ;
      RECT  207.1 290.4 207.9 279.6 ;
      RECT  203.5 290.4 204.3 279.6 ;
      RECT  208.7 290.4 209.5 301.2 ;
      RECT  201.9 290.4 202.7 301.2 ;
      RECT  205.3 300.4 206.1 301.2 ;
      RECT  207.1 290.4 207.9 301.2 ;
      RECT  203.5 290.4 204.3 301.2 ;
      RECT  208.7 311.2 209.5 300.4 ;
      RECT  201.9 311.2 202.7 300.4 ;
      RECT  205.3 301.2 206.1 300.4 ;
      RECT  207.1 311.2 207.9 300.4 ;
      RECT  203.5 311.2 204.3 300.4 ;
      RECT  208.7 311.2 209.5 322.0 ;
      RECT  201.9 311.2 202.7 322.0 ;
      RECT  205.3 321.2 206.1 322.0 ;
      RECT  207.1 311.2 207.9 322.0 ;
      RECT  203.5 311.2 204.3 322.0 ;
      RECT  208.7 332.0 209.5 321.2 ;
      RECT  201.9 332.0 202.7 321.2 ;
      RECT  205.3 322.0 206.1 321.2 ;
      RECT  207.1 332.0 207.9 321.2 ;
      RECT  203.5 332.0 204.3 321.2 ;
      RECT  208.7 332.0 209.5 342.8 ;
      RECT  201.9 332.0 202.7 342.8 ;
      RECT  205.3 342.0 206.1 342.8 ;
      RECT  207.1 332.0 207.9 342.8 ;
      RECT  203.5 332.0 204.3 342.8 ;
      RECT  208.7 352.8 209.5 342.0 ;
      RECT  201.9 352.8 202.7 342.0 ;
      RECT  205.3 342.8 206.1 342.0 ;
      RECT  207.1 352.8 207.9 342.0 ;
      RECT  203.5 352.8 204.3 342.0 ;
      RECT  208.7 352.8 209.5 363.6 ;
      RECT  201.9 352.8 202.7 363.6 ;
      RECT  205.3 362.8 206.1 363.6 ;
      RECT  207.1 352.8 207.9 363.6 ;
      RECT  203.5 352.8 204.3 363.6 ;
      RECT  205.3 279.6 206.1 280.4 ;
      RECT  205.3 279.6 206.1 280.4 ;
      RECT  205.3 217.2 206.1 218.0 ;
      RECT  205.3 217.2 206.1 218.0 ;
      RECT  205.3 342.0 206.1 342.8 ;
      RECT  205.3 300.4 206.1 301.2 ;
      RECT  205.3 300.4 206.1 301.2 ;
      RECT  205.3 362.8 206.1 363.6 ;
      RECT  205.3 175.6 206.1 176.4 ;
      RECT  205.3 196.4 206.1 197.2 ;
      RECT  205.3 321.2 206.1 322.0 ;
      RECT  205.3 238.0 206.1 238.8 ;
      RECT  205.3 258.8 206.1 259.6 ;
      RECT  201.9 279.6 202.7 290.4 ;
      RECT  201.9 332.0 202.7 342.8 ;
      RECT  208.7 196.4 209.5 207.2 ;
      RECT  201.9 228.0 202.7 238.8 ;
      RECT  208.7 279.6 209.5 290.4 ;
      RECT  208.7 321.2 209.5 332.0 ;
      RECT  208.7 269.6 209.5 280.4 ;
      RECT  208.7 175.6 209.5 186.4 ;
      RECT  208.7 217.2 209.5 228.0 ;
      RECT  208.7 248.8 209.5 259.6 ;
      RECT  201.9 300.4 202.7 311.2 ;
      RECT  208.7 258.8 209.5 269.6 ;
      RECT  201.9 311.2 202.7 322.0 ;
      RECT  201.9 207.2 202.7 218.0 ;
      RECT  201.9 175.6 202.7 186.4 ;
      RECT  208.7 228.0 209.5 238.8 ;
      RECT  201.9 342.0 202.7 352.8 ;
      RECT  201.9 352.8 202.7 363.6 ;
      RECT  201.9 290.4 202.7 301.2 ;
      RECT  208.7 290.4 209.5 301.2 ;
      RECT  208.7 342.0 209.5 352.8 ;
      RECT  201.9 196.4 202.7 207.2 ;
      RECT  208.7 238.0 209.5 248.8 ;
      RECT  201.9 186.4 202.7 197.2 ;
      RECT  208.7 332.0 209.5 342.8 ;
      RECT  208.7 352.8 209.5 363.6 ;
      RECT  201.9 217.2 202.7 228.0 ;
      RECT  201.9 238.0 202.7 248.8 ;
      RECT  208.7 165.6 209.5 176.4 ;
      RECT  201.9 248.8 202.7 259.6 ;
      RECT  201.9 321.2 202.7 332.0 ;
      RECT  208.7 300.4 209.5 311.2 ;
      RECT  208.7 207.2 209.5 218.0 ;
      RECT  201.9 258.8 202.7 269.6 ;
      RECT  201.9 269.6 202.7 280.4 ;
      RECT  208.7 186.4 209.5 197.2 ;
      RECT  208.7 311.2 209.5 322.0 ;
      RECT  201.9 165.6 202.7 176.4 ;
      RECT  183.1 165.6 183.9 363.2 ;
      RECT  186.7 165.6 187.5 363.2 ;
      RECT  189.9 165.6 190.7 363.2 ;
      RECT  193.5 165.6 194.3 363.2 ;
      RECT  196.7 165.6 197.5 363.2 ;
      RECT  200.3 165.6 201.1 363.2 ;
      RECT  184.9 321.2 185.7 322.0 ;
      RECT  184.9 279.6 185.7 280.4 ;
      RECT  184.9 196.4 185.7 197.2 ;
      RECT  184.9 300.4 185.7 301.2 ;
      RECT  184.9 258.8 185.7 259.6 ;
      RECT  184.9 238.0 185.7 238.8 ;
      RECT  184.9 342.0 185.7 342.8 ;
      RECT  184.9 175.6 185.7 176.4 ;
      RECT  184.9 217.2 185.7 218.0 ;
      RECT  188.3 311.2 189.1 322.0 ;
      RECT  181.5 207.2 182.3 218.0 ;
      RECT  181.5 342.0 182.3 352.8 ;
      RECT  188.3 238.0 189.1 248.8 ;
      RECT  181.5 238.0 182.3 248.8 ;
      RECT  188.3 228.0 189.1 238.8 ;
      RECT  188.3 175.6 189.1 186.4 ;
      RECT  188.3 207.2 189.1 218.0 ;
      RECT  188.3 186.4 189.1 197.2 ;
      RECT  188.3 258.8 189.1 269.6 ;
      RECT  181.5 269.6 182.3 280.4 ;
      RECT  188.3 300.4 189.1 311.2 ;
      RECT  188.3 279.6 189.1 290.4 ;
      RECT  188.3 269.6 189.1 280.4 ;
      RECT  181.5 258.8 182.3 269.6 ;
      RECT  188.3 196.4 189.1 207.2 ;
      RECT  188.3 248.8 189.1 259.6 ;
      RECT  181.5 186.4 182.3 197.2 ;
      RECT  188.3 290.4 189.1 301.2 ;
      RECT  181.5 279.6 182.3 290.4 ;
      RECT  181.5 228.0 182.3 238.8 ;
      RECT  188.3 321.2 189.1 332.0 ;
      RECT  181.5 321.2 182.3 332.0 ;
      RECT  181.5 290.4 182.3 301.2 ;
      RECT  181.5 311.2 182.3 322.0 ;
      RECT  181.5 175.6 182.3 186.4 ;
      RECT  188.3 332.0 189.1 342.8 ;
      RECT  181.5 332.0 182.3 342.8 ;
      RECT  181.5 300.4 182.3 311.2 ;
      RECT  181.5 196.4 182.3 207.2 ;
      RECT  188.3 342.0 189.1 352.8 ;
      RECT  188.3 217.2 189.1 228.0 ;
      RECT  181.5 217.2 182.3 228.0 ;
      RECT  181.5 248.8 182.3 259.6 ;
      RECT  183.0 149.4 183.6 161.4 ;
      RECT  187.0 149.4 187.6 161.4 ;
      RECT  189.8 149.4 190.4 161.4 ;
      RECT  193.8 149.4 194.4 161.4 ;
      RECT  196.6 149.4 197.2 161.4 ;
      RECT  200.6 149.4 201.2 161.4 ;
      RECT  183.0 149.4 183.6 161.4 ;
      RECT  187.0 149.4 187.6 161.4 ;
      RECT  189.8 149.4 190.4 161.4 ;
      RECT  193.8 149.4 194.4 161.4 ;
      RECT  196.6 149.4 197.2 161.4 ;
      RECT  200.6 149.4 201.2 161.4 ;
      RECT  194.1 125.0 194.9 126.6 ;
      RECT  192.7 121.4 193.9 122.2 ;
      RECT  190.7 121.4 192.1 122.2 ;
      RECT  190.7 122.2 191.5 145.2 ;
      RECT  192.7 122.2 193.5 145.2 ;
      RECT  195.1 138.4 195.9 140.0 ;
      RECT  190.7 112.6 191.5 121.4 ;
      RECT  192.7 112.6 193.5 121.4 ;
      RECT  189.3 112.6 190.1 115.6 ;
      RECT  200.9 125.0 201.7 126.6 ;
      RECT  199.5 121.4 200.7 122.2 ;
      RECT  197.5 121.4 198.9 122.2 ;
      RECT  197.5 122.2 198.3 145.2 ;
      RECT  199.5 122.2 200.3 145.2 ;
      RECT  201.9 138.4 202.7 140.0 ;
      RECT  197.5 112.6 198.3 121.4 ;
      RECT  199.5 112.6 200.3 121.4 ;
      RECT  196.1 112.6 196.9 115.6 ;
      RECT  189.3 112.6 190.1 115.6 ;
      RECT  190.7 122.2 191.5 145.2 ;
      RECT  192.7 122.2 193.5 145.2 ;
      RECT  196.1 112.6 196.9 115.6 ;
      RECT  197.5 122.2 198.3 145.2 ;
      RECT  199.5 122.2 200.3 145.2 ;
      RECT  190.7 106.4 191.5 108.4 ;
      RECT  192.5 80.6 193.3 81.4 ;
      RECT  192.5 74.0 193.3 74.8 ;
      RECT  191.1 99.6 191.9 100.4 ;
      RECT  193.9 85.0 194.7 85.8 ;
      RECT  191.9 91.4 192.7 92.2 ;
      RECT  191.7 67.8 192.5 69.8 ;
      RECT  192.7 103.4 193.5 108.4 ;
      RECT  197.5 106.4 198.3 108.4 ;
      RECT  199.3 80.6 200.1 81.4 ;
      RECT  199.3 74.0 200.1 74.8 ;
      RECT  197.9 99.6 198.7 100.4 ;
      RECT  200.7 85.0 201.5 85.8 ;
      RECT  198.7 91.4 199.5 92.2 ;
      RECT  198.5 67.8 199.3 69.8 ;
      RECT  199.5 103.4 200.3 108.4 ;
      RECT  191.7 67.8 192.5 69.8 ;
      RECT  198.5 67.8 199.3 69.8 ;
      RECT  190.7 106.4 191.5 108.4 ;
      RECT  192.7 103.4 193.5 108.4 ;
      RECT  197.5 106.4 198.3 108.4 ;
      RECT  199.5 103.4 200.3 108.4 ;
      RECT  183.0 161.4 183.6 149.4 ;
      RECT  187.0 161.4 187.6 149.4 ;
      RECT  189.8 161.4 190.4 149.4 ;
      RECT  193.8 161.4 194.4 149.4 ;
      RECT  196.6 161.4 197.2 149.4 ;
      RECT  200.6 161.4 201.2 149.4 ;
      RECT  189.3 115.6 190.1 112.6 ;
      RECT  196.1 115.6 196.9 112.6 ;
      RECT  191.7 69.8 192.5 67.8 ;
      RECT  198.5 69.8 199.3 67.8 ;
      RECT  89.8 191.0 90.6 191.8 ;
      RECT  91.2 201.8 92.0 202.6 ;
      RECT  89.8 253.4 90.6 254.2 ;
      RECT  91.2 264.2 92.0 265.0 ;
      RECT  82.3 186.4 82.9 290.4 ;
      RECT  83.7 186.4 84.3 290.4 ;
      RECT  85.1 186.4 85.7 290.4 ;
      RECT  86.5 186.4 87.1 290.4 ;
      RECT  156.6 186.4 157.2 352.8 ;
      RECT  82.3 186.4 82.9 290.4 ;
      RECT  83.7 186.4 84.3 290.4 ;
      RECT  85.1 186.4 85.7 290.4 ;
      RECT  86.5 186.4 87.1 290.4 ;
      RECT  157.3 181.1 157.9 181.7 ;
      RECT  189.3 112.6 190.1 115.6 ;
      RECT  196.1 112.6 196.9 115.6 ;
      RECT  191.7 67.8 192.5 69.8 ;
      RECT  198.5 67.8 199.3 69.8 ;
      RECT  82.3 186.4 82.9 290.4 ;
      RECT  83.7 186.4 84.3 290.4 ;
      RECT  85.1 186.4 85.7 290.4 ;
      RECT  86.5 186.4 87.1 290.4 ;
      RECT  164.6 67.8 165.2 165.6 ;
      RECT  167.4 67.8 168.0 165.6 ;
      RECT  166.0 67.8 166.6 165.6 ;
      RECT  168.8 67.8 169.4 165.6 ;
      RECT  6.8 6.0 7.6 17.6 ;
      RECT  16.4 6.0 17.2 17.6 ;
      RECT  5.2 9.4 6.0 10.2 ;
      RECT  10.0 11.4 10.8 12.2 ;
      RECT  3.6 8.0 4.4 13.6 ;
      RECT  21.2 12.2 22.0 13.0 ;
      RECT  10.0 11.4 10.8 12.2 ;
      RECT  38.2 8.9 38.8 9.5 ;
      RECT  32.6 14.9 33.2 15.5 ;
      RECT  5.2 9.4 6.0 10.2 ;
      RECT  6.8 39.6 7.6 28.0 ;
      RECT  16.4 39.6 17.2 28.0 ;
      RECT  5.2 36.2 6.0 35.4 ;
      RECT  10.0 34.2 10.8 33.4 ;
      RECT  3.6 37.6 4.4 32.0 ;
      RECT  21.2 33.4 22.0 32.6 ;
      RECT  10.0 34.2 10.8 33.4 ;
      RECT  38.2 36.7 38.8 36.1 ;
      RECT  32.6 30.7 33.2 30.1 ;
      RECT  5.2 36.2 6.0 35.4 ;
      RECT  10.0 11.4 10.8 12.2 ;
      RECT  10.0 33.4 10.8 34.2 ;
      RECT  38.2 8.9 38.8 9.5 ;
      RECT  32.6 14.9 33.2 15.5 ;
      RECT  38.2 36.1 38.8 36.7 ;
      RECT  32.6 30.1 33.2 30.7 ;
      RECT  5.2 2.8 5.8 42.8 ;
      RECT  33.8 165.6 33.2 175.2 ;
      RECT  5.5 165.6 4.9 332.0 ;
      RECT  10.0 11.4 10.8 12.2 ;
      RECT  10.0 33.4 10.8 34.2 ;
      RECT  54.1 12.3 54.7 12.9 ;
      RECT  33.2 165.6 33.8 175.2 ;
      RECT  65.9 152.9 79.4 153.5 ;
      RECT  65.7 91.5 79.4 92.1 ;
      RECT  71.5 112.7 79.4 113.3 ;
      RECT  73.3 73.5 79.4 74.1 ;
      RECT  74.8 11.5 79.4 12.1 ;
      RECT  62.0 348.0 62.8 359.6 ;
      RECT  71.6 348.0 72.4 359.6 ;
      RECT  60.4 351.4 61.2 352.2 ;
      RECT  65.2 353.4 66.0 354.2 ;
      RECT  58.8 350.0 59.6 355.6 ;
      RECT  76.4 354.2 77.2 355.0 ;
      RECT  62.0 381.6 62.8 370.0 ;
      RECT  71.6 381.6 72.4 370.0 ;
      RECT  60.4 378.2 61.2 377.4 ;
      RECT  65.2 376.2 66.0 375.4 ;
      RECT  58.8 379.6 59.6 374.0 ;
      RECT  76.4 375.4 77.2 374.6 ;
      RECT  62.0 388.0 62.8 399.6 ;
      RECT  71.6 388.0 72.4 399.6 ;
      RECT  60.4 391.4 61.2 392.2 ;
      RECT  65.2 393.4 66.0 394.2 ;
      RECT  58.8 390.0 59.6 395.6 ;
      RECT  76.4 394.2 77.2 395.0 ;
      RECT  62.0 421.6 62.8 410.0 ;
      RECT  71.6 421.6 72.4 410.0 ;
      RECT  60.4 418.2 61.2 417.4 ;
      RECT  65.2 416.2 66.0 415.4 ;
      RECT  58.8 419.6 59.6 414.0 ;
      RECT  76.4 415.4 77.2 414.6 ;
      RECT  65.2 353.4 66.0 354.2 ;
      RECT  65.2 375.4 66.0 376.2 ;
      RECT  65.2 393.4 66.0 394.2 ;
      RECT  65.2 415.4 66.0 416.2 ;
      RECT  76.4 354.2 77.2 355.0 ;
      RECT  76.4 374.6 77.2 375.4 ;
      RECT  76.4 394.2 77.2 395.0 ;
      RECT  76.4 414.6 77.2 415.4 ;
      RECT  105.6 6.0 106.4 17.6 ;
      RECT  115.2 6.0 116.0 17.6 ;
      RECT  104.0 9.4 104.8 10.2 ;
      RECT  108.8 11.4 109.6 12.2 ;
      RECT  102.4 8.0 103.2 13.6 ;
      RECT  120.0 12.2 120.8 13.0 ;
      RECT  127.4 6.0 128.2 17.6 ;
      RECT  137.0 6.0 137.8 17.6 ;
      RECT  125.8 9.4 126.6 10.2 ;
      RECT  130.6 11.4 131.4 12.2 ;
      RECT  124.2 8.0 125.0 13.6 ;
      RECT  141.8 12.2 142.6 13.0 ;
      RECT  108.8 11.4 109.6 12.2 ;
      RECT  130.6 11.4 131.4 12.2 ;
      RECT  120.0 12.2 120.8 13.0 ;
      RECT  141.8 12.2 142.6 13.0 ;
   LAYER  metal3 ;
      RECT  184.9 175.6 185.7 176.4 ;
      RECT  184.9 362.8 185.7 363.6 ;
      RECT  188.3 357.8 189.1 358.6 ;
      RECT  181.5 170.6 182.3 171.4 ;
      RECT  188.3 170.6 189.1 171.4 ;
      RECT  181.5 357.8 182.3 358.6 ;
      RECT  205.3 196.4 206.1 197.2 ;
      RECT  184.9 362.8 185.7 363.6 ;
      RECT  178.1 279.6 178.9 280.4 ;
      RECT  205.3 238.0 206.1 238.8 ;
      RECT  178.1 238.0 178.9 238.8 ;
      RECT  198.5 175.6 199.3 176.4 ;
      RECT  178.1 175.6 178.9 176.4 ;
      RECT  205.3 258.8 206.1 259.6 ;
      RECT  178.1 300.4 178.9 301.2 ;
      RECT  191.7 362.8 192.5 363.6 ;
      RECT  205.3 175.6 206.1 176.4 ;
      RECT  178.1 342.0 178.9 342.8 ;
      RECT  205.3 362.8 206.1 363.6 ;
      RECT  178.1 321.2 178.9 322.0 ;
      RECT  191.7 175.6 192.5 176.4 ;
      RECT  178.1 362.8 178.9 363.6 ;
      RECT  205.3 342.0 206.1 342.8 ;
      RECT  178.1 258.8 178.9 259.6 ;
      RECT  178.1 217.2 178.9 218.0 ;
      RECT  205.3 217.2 206.1 218.0 ;
      RECT  205.3 321.2 206.1 322.0 ;
      RECT  205.3 300.4 206.1 301.2 ;
      RECT  198.5 362.8 199.3 363.6 ;
      RECT  184.9 175.6 185.7 176.4 ;
      RECT  205.3 279.6 206.1 280.4 ;
      RECT  178.1 196.4 178.9 197.2 ;
      RECT  181.5 263.8 182.3 264.6 ;
      RECT  208.7 284.6 209.5 285.4 ;
      RECT  201.9 170.6 202.7 171.4 ;
      RECT  201.9 347.0 202.7 347.8 ;
      RECT  201.9 170.6 202.7 171.4 ;
      RECT  201.9 253.8 202.7 254.6 ;
      RECT  181.5 253.8 182.3 254.6 ;
      RECT  201.9 263.8 202.7 264.6 ;
      RECT  201.9 222.2 202.7 223.0 ;
      RECT  181.5 295.4 182.3 296.2 ;
      RECT  174.7 243.0 175.5 243.8 ;
      RECT  174.7 337.0 175.5 337.8 ;
      RECT  181.5 316.2 182.3 317.0 ;
      RECT  181.5 243.0 182.3 243.8 ;
      RECT  174.7 347.0 175.5 347.8 ;
      RECT  201.9 212.2 202.7 213.0 ;
      RECT  181.5 347.0 182.3 347.8 ;
      RECT  208.7 347.0 209.5 347.8 ;
      RECT  172.6 167.8 173.4 168.6 ;
      RECT  181.5 170.6 182.3 171.4 ;
      RECT  181.5 170.6 182.3 171.4 ;
      RECT  208.7 274.6 209.5 275.4 ;
      RECT  201.9 337.0 202.7 337.8 ;
      RECT  174.7 263.8 175.5 264.6 ;
      RECT  181.5 357.8 182.3 358.6 ;
      RECT  181.5 357.8 182.3 358.6 ;
      RECT  208.7 222.2 209.5 223.0 ;
      RECT  174.7 357.8 175.5 358.6 ;
      RECT  201.9 357.8 202.7 358.6 ;
      RECT  201.9 357.8 202.7 358.6 ;
      RECT  208.7 243.0 209.5 243.8 ;
      RECT  174.7 316.2 175.5 317.0 ;
      RECT  174.7 326.2 175.5 327.0 ;
      RECT  181.5 337.0 182.3 337.8 ;
      RECT  201.9 243.0 202.7 243.8 ;
      RECT  195.1 170.6 195.9 171.4 ;
      RECT  195.1 357.8 195.9 358.6 ;
      RECT  210.8 167.8 211.6 168.6 ;
      RECT  201.9 233.0 202.7 233.8 ;
      RECT  201.9 316.2 202.7 317.0 ;
      RECT  208.7 191.4 209.5 192.2 ;
      RECT  181.5 284.6 182.3 285.4 ;
      RECT  208.7 180.6 209.5 181.4 ;
      RECT  208.7 305.4 209.5 306.2 ;
      RECT  208.7 201.4 209.5 202.2 ;
      RECT  174.7 233.0 175.5 233.8 ;
      RECT  208.7 253.8 209.5 254.6 ;
      RECT  174.7 305.4 175.5 306.2 ;
      RECT  181.5 233.0 182.3 233.8 ;
      RECT  201.9 274.6 202.7 275.4 ;
      RECT  208.7 233.0 209.5 233.8 ;
      RECT  208.7 212.2 209.5 213.0 ;
      RECT  208.7 337.0 209.5 337.8 ;
      RECT  181.5 305.4 182.3 306.2 ;
      RECT  174.7 284.6 175.5 285.4 ;
      RECT  208.7 326.2 209.5 327.0 ;
      RECT  201.9 191.4 202.7 192.2 ;
      RECT  201.9 284.6 202.7 285.4 ;
      RECT  201.9 295.4 202.7 296.2 ;
      RECT  174.7 170.6 175.5 171.4 ;
      RECT  208.7 316.2 209.5 317.0 ;
      RECT  174.7 274.6 175.5 275.4 ;
      RECT  208.7 170.6 209.5 171.4 ;
      RECT  174.7 191.4 175.5 192.2 ;
      RECT  174.7 201.4 175.5 202.2 ;
      RECT  181.5 191.4 182.3 192.2 ;
      RECT  188.3 170.6 189.1 171.4 ;
      RECT  188.3 170.6 189.1 171.4 ;
      RECT  174.7 222.2 175.5 223.0 ;
      RECT  201.9 305.4 202.7 306.2 ;
      RECT  174.7 212.2 175.5 213.0 ;
      RECT  181.5 212.2 182.3 213.0 ;
      RECT  174.7 180.6 175.5 181.4 ;
      RECT  201.9 201.4 202.7 202.2 ;
      RECT  208.7 295.4 209.5 296.2 ;
      RECT  181.5 326.2 182.3 327.0 ;
      RECT  201.9 326.2 202.7 327.0 ;
      RECT  188.3 357.8 189.1 358.6 ;
      RECT  188.3 357.8 189.1 358.6 ;
      RECT  181.5 180.6 182.3 181.4 ;
      RECT  181.5 201.4 182.3 202.2 ;
      RECT  208.7 357.8 209.5 358.6 ;
      RECT  181.5 274.6 182.3 275.4 ;
      RECT  181.5 222.2 182.3 223.0 ;
      RECT  210.8 355.0 211.6 355.8 ;
      RECT  172.6 355.0 173.4 355.8 ;
      RECT  174.7 295.4 175.5 296.2 ;
      RECT  201.9 180.6 202.7 181.4 ;
      RECT  174.7 253.8 175.5 254.6 ;
      RECT  208.7 263.8 209.5 264.6 ;
      RECT  185.4 159.6 186.2 160.4 ;
      RECT  192.2 159.6 193.0 160.4 ;
      RECT  199.0 159.6 199.8 160.4 ;
      RECT  192.2 159.6 193.0 160.4 ;
      RECT  199.0 159.6 199.8 160.4 ;
      RECT  185.4 159.6 186.2 160.4 ;
      RECT  200.9 125.4 201.7 126.2 ;
      RECT  194.1 125.4 194.9 126.2 ;
      RECT  201.9 138.8 202.7 139.6 ;
      RECT  195.1 138.8 195.9 139.6 ;
      RECT  198.7 91.4 199.5 92.2 ;
      RECT  191.9 91.4 192.7 92.2 ;
      RECT  192.5 74.0 193.3 74.8 ;
      RECT  199.3 74.0 200.1 74.8 ;
      RECT  200.7 85.0 201.5 85.8 ;
      RECT  191.1 99.6 191.9 100.4 ;
      RECT  197.9 99.6 198.7 100.4 ;
      RECT  193.9 85.0 194.7 85.8 ;
      RECT  192.5 80.6 193.3 81.4 ;
      RECT  199.3 80.6 200.1 81.4 ;
      RECT  198.7 92.2 199.5 91.4 ;
      RECT  199.3 74.8 200.1 74.0 ;
      RECT  192.2 160.4 193.0 159.6 ;
      RECT  192.5 74.8 193.3 74.0 ;
      RECT  200.9 126.2 201.7 125.4 ;
      RECT  191.9 92.2 192.7 91.4 ;
      RECT  199.0 160.4 199.8 159.6 ;
      RECT  185.4 160.4 186.2 159.6 ;
      RECT  194.1 126.2 194.9 125.4 ;
      RECT  192.5 81.4 193.3 80.6 ;
      RECT  197.9 100.4 198.7 99.6 ;
      RECT  201.9 139.6 202.7 138.8 ;
      RECT  195.1 139.6 195.9 138.8 ;
      RECT  200.7 85.8 201.5 85.0 ;
      RECT  191.1 100.4 191.9 99.6 ;
      RECT  199.3 81.4 200.1 80.6 ;
      RECT  193.9 85.8 194.7 85.0 ;
      RECT  108.1 196.4 108.9 197.2 ;
      RECT  108.1 196.4 108.9 197.2 ;
      RECT  93.1 217.2 93.9 218.0 ;
      RECT  93.1 217.2 93.9 218.0 ;
      RECT  93.1 196.4 93.9 197.2 ;
      RECT  93.1 196.4 93.9 197.2 ;
      RECT  108.1 217.2 108.9 218.0 ;
      RECT  108.1 217.2 108.9 218.0 ;
      RECT  108.1 227.6 108.9 228.4 ;
      RECT  93.1 227.6 93.9 228.4 ;
      RECT  93.1 186.0 93.9 186.8 ;
      RECT  108.1 206.8 108.9 207.6 ;
      RECT  108.1 186.0 108.9 186.8 ;
      RECT  93.1 206.8 93.9 207.6 ;
      RECT  108.1 258.8 108.9 259.6 ;
      RECT  108.1 258.8 108.9 259.6 ;
      RECT  93.1 279.6 93.9 280.4 ;
      RECT  93.1 279.6 93.9 280.4 ;
      RECT  93.1 258.8 93.9 259.6 ;
      RECT  93.1 258.8 93.9 259.6 ;
      RECT  108.1 279.6 108.9 280.4 ;
      RECT  108.1 279.6 108.9 280.4 ;
      RECT  108.1 290.0 108.9 290.8 ;
      RECT  93.1 290.0 93.9 290.8 ;
      RECT  93.1 248.4 93.9 249.2 ;
      RECT  108.1 269.2 108.9 270.0 ;
      RECT  108.1 248.4 108.9 249.2 ;
      RECT  93.1 269.2 93.9 270.0 ;
      RECT  108.1 217.2 108.9 218.0 ;
      RECT  152.0 258.8 152.8 259.6 ;
      RECT  152.0 258.8 152.8 259.6 ;
      RECT  108.1 196.4 108.9 197.2 ;
      RECT  152.0 321.2 152.8 322.0 ;
      RECT  152.0 196.4 152.8 197.2 ;
      RECT  152.0 196.4 152.8 197.2 ;
      RECT  93.1 258.8 93.9 259.6 ;
      RECT  108.1 279.6 108.9 280.4 ;
      RECT  152.0 279.6 152.8 280.4 ;
      RECT  93.1 196.4 93.9 197.2 ;
      RECT  93.1 279.6 93.9 280.4 ;
      RECT  152.0 217.2 152.8 218.0 ;
      RECT  152.0 217.2 152.8 218.0 ;
      RECT  152.0 279.6 152.8 280.4 ;
      RECT  152.0 300.4 152.8 301.2 ;
      RECT  108.1 258.8 108.9 259.6 ;
      RECT  152.0 342.0 152.8 342.8 ;
      RECT  152.0 238.0 152.8 238.8 ;
      RECT  93.1 217.2 93.9 218.0 ;
      RECT  152.0 206.8 152.8 207.6 ;
      RECT  108.1 290.0 108.9 290.8 ;
      RECT  93.1 206.8 93.9 207.6 ;
      RECT  108.1 206.8 108.9 207.6 ;
      RECT  108.1 186.0 108.9 186.8 ;
      RECT  152.0 269.2 152.8 270.0 ;
      RECT  93.1 248.4 93.9 249.2 ;
      RECT  93.1 269.2 93.9 270.0 ;
      RECT  93.1 227.6 93.9 228.4 ;
      RECT  108.1 248.4 108.9 249.2 ;
      RECT  93.1 186.0 93.9 186.8 ;
      RECT  152.0 331.6 152.8 332.4 ;
      RECT  108.1 269.2 108.9 270.0 ;
      RECT  93.1 290.0 93.9 290.8 ;
      RECT  108.1 227.6 108.9 228.4 ;
      RECT  152.0 310.8 152.8 311.6 ;
      RECT  152.0 186.0 152.8 186.8 ;
      RECT  152.0 290.0 152.8 290.8 ;
      RECT  152.0 352.4 152.8 353.2 ;
      RECT  152.0 248.4 152.8 249.2 ;
      RECT  152.0 227.6 152.8 228.4 ;
      RECT  167.2 258.8 168.0 259.6 ;
      RECT  167.2 279.6 168.0 280.4 ;
      RECT  167.2 279.6 168.0 280.4 ;
      RECT  167.2 300.4 168.0 301.2 ;
      RECT  167.2 238.0 168.0 238.8 ;
      RECT  167.2 342.0 168.0 342.8 ;
      RECT  167.2 217.2 168.0 218.0 ;
      RECT  167.2 196.4 168.0 197.2 ;
      RECT  167.2 217.2 168.0 218.0 ;
      RECT  167.2 196.4 168.0 197.2 ;
      RECT  167.2 321.2 168.0 322.0 ;
      RECT  167.2 258.8 168.0 259.6 ;
      RECT  167.2 269.2 168.0 270.0 ;
      RECT  167.2 331.6 168.0 332.4 ;
      RECT  167.2 310.8 168.0 311.6 ;
      RECT  167.2 227.6 168.0 228.4 ;
      RECT  167.2 248.4 168.0 249.2 ;
      RECT  167.2 206.8 168.0 207.6 ;
      RECT  167.2 352.4 168.0 353.2 ;
      RECT  167.2 186.0 168.0 186.8 ;
      RECT  167.2 290.0 168.0 290.8 ;
      RECT  155.2 175.6 156.0 176.4 ;
      RECT  152.0 258.8 152.8 259.6 ;
      RECT  152.0 279.6 152.8 280.4 ;
      RECT  167.2 196.4 168.0 197.2 ;
      RECT  152.0 300.4 152.8 301.2 ;
      RECT  152.0 321.2 152.8 322.0 ;
      RECT  93.1 258.8 93.9 259.6 ;
      RECT  167.2 342.0 168.0 342.8 ;
      RECT  167.2 238.0 168.0 238.8 ;
      RECT  152.0 238.0 152.8 238.8 ;
      RECT  93.1 196.4 93.9 197.2 ;
      RECT  108.1 258.8 108.9 259.6 ;
      RECT  167.2 321.2 168.0 322.0 ;
      RECT  152.0 217.2 152.8 218.0 ;
      RECT  93.1 217.2 93.9 218.0 ;
      RECT  167.2 279.6 168.0 280.4 ;
      RECT  93.1 279.6 93.9 280.4 ;
      RECT  167.2 258.8 168.0 259.6 ;
      RECT  152.0 196.4 152.8 197.2 ;
      RECT  108.1 196.4 108.9 197.2 ;
      RECT  167.2 300.4 168.0 301.2 ;
      RECT  167.2 217.2 168.0 218.0 ;
      RECT  152.0 342.0 152.8 342.8 ;
      RECT  108.1 279.6 108.9 280.4 ;
      RECT  108.1 217.2 108.9 218.0 ;
      RECT  152.0 227.6 152.8 228.4 ;
      RECT  108.1 248.4 108.9 249.2 ;
      RECT  93.1 186.0 93.9 186.8 ;
      RECT  152.0 331.6 152.8 332.4 ;
      RECT  152.0 290.0 152.8 290.8 ;
      RECT  167.2 227.6 168.0 228.4 ;
      RECT  167.2 206.8 168.0 207.6 ;
      RECT  167.2 352.4 168.0 353.2 ;
      RECT  108.1 227.6 108.9 228.4 ;
      RECT  152.0 352.4 152.8 353.2 ;
      RECT  93.1 269.2 93.9 270.0 ;
      RECT  167.2 269.2 168.0 270.0 ;
      RECT  152.0 310.8 152.8 311.6 ;
      RECT  152.0 206.8 152.8 207.6 ;
      RECT  167.2 290.0 168.0 290.8 ;
      RECT  108.1 290.0 108.9 290.8 ;
      RECT  167.2 331.6 168.0 332.4 ;
      RECT  167.2 310.8 168.0 311.6 ;
      RECT  152.0 248.4 152.8 249.2 ;
      RECT  152.0 269.2 152.8 270.0 ;
      RECT  108.1 186.0 108.9 186.8 ;
      RECT  167.2 186.0 168.0 186.8 ;
      RECT  93.1 290.0 93.9 290.8 ;
      RECT  108.1 269.2 108.9 270.0 ;
      RECT  167.2 248.4 168.0 249.2 ;
      RECT  93.1 227.6 93.9 228.4 ;
      RECT  108.1 206.8 108.9 207.6 ;
      RECT  93.1 206.8 93.9 207.6 ;
      RECT  93.1 248.4 93.9 249.2 ;
      RECT  152.0 186.0 152.8 186.8 ;
      RECT  82.2 147.7 183.3 148.3 ;
      RECT  199.0 159.6 199.8 160.4 ;
      RECT  191.9 91.4 192.7 92.2 ;
      RECT  205.3 196.4 206.1 197.2 ;
      RECT  194.1 125.4 194.9 126.2 ;
      RECT  184.9 362.8 185.7 363.6 ;
      RECT  178.1 279.6 178.9 280.4 ;
      RECT  152.0 321.2 152.8 322.0 ;
      RECT  205.3 238.0 206.1 238.8 ;
      RECT  178.1 238.0 178.9 238.8 ;
      RECT  198.5 175.6 199.3 176.4 ;
      RECT  192.5 74.0 193.3 74.8 ;
      RECT  178.1 175.6 178.9 176.4 ;
      RECT  205.3 258.8 206.1 259.6 ;
      RECT  200.9 125.4 201.7 126.2 ;
      RECT  167.2 279.6 168.0 280.4 ;
      RECT  152.0 196.4 152.8 197.2 ;
      RECT  167.2 300.4 168.0 301.2 ;
      RECT  178.1 300.4 178.9 301.2 ;
      RECT  108.1 279.6 108.9 280.4 ;
      RECT  192.2 159.6 193.0 160.4 ;
      RECT  167.2 217.2 168.0 218.0 ;
      RECT  93.1 196.4 93.9 197.2 ;
      RECT  93.1 279.6 93.9 280.4 ;
      RECT  152.0 217.2 152.8 218.0 ;
      RECT  191.7 362.8 192.5 363.6 ;
      RECT  167.2 258.8 168.0 259.6 ;
      RECT  199.3 74.0 200.1 74.8 ;
      RECT  93.1 217.2 93.9 218.0 ;
      RECT  205.3 175.6 206.1 176.4 ;
      RECT  152.0 300.4 152.8 301.2 ;
      RECT  178.1 342.0 178.9 342.8 ;
      RECT  205.3 362.8 206.1 363.6 ;
      RECT  178.1 321.2 178.9 322.0 ;
      RECT  191.7 175.6 192.5 176.4 ;
      RECT  108.1 258.8 108.9 259.6 ;
      RECT  93.1 258.8 93.9 259.6 ;
      RECT  178.1 362.8 178.9 363.6 ;
      RECT  205.3 342.0 206.1 342.8 ;
      RECT  198.7 91.4 199.5 92.2 ;
      RECT  178.1 258.8 178.9 259.6 ;
      RECT  185.4 159.6 186.2 160.4 ;
      RECT  178.1 217.2 178.9 218.0 ;
      RECT  155.2 175.6 156.0 176.4 ;
      RECT  152.0 279.6 152.8 280.4 ;
      RECT  167.2 196.4 168.0 197.2 ;
      RECT  205.3 217.2 206.1 218.0 ;
      RECT  108.1 217.2 108.9 218.0 ;
      RECT  167.2 342.0 168.0 342.8 ;
      RECT  152.0 258.8 152.8 259.6 ;
      RECT  205.3 321.2 206.1 322.0 ;
      RECT  205.3 300.4 206.1 301.2 ;
      RECT  167.2 238.0 168.0 238.8 ;
      RECT  152.0 238.0 152.8 238.8 ;
      RECT  198.5 362.8 199.3 363.6 ;
      RECT  184.9 175.6 185.7 176.4 ;
      RECT  167.2 321.2 168.0 322.0 ;
      RECT  152.0 342.0 152.8 342.8 ;
      RECT  108.1 196.4 108.9 197.2 ;
      RECT  205.3 279.6 206.1 280.4 ;
      RECT  178.1 196.4 178.9 197.2 ;
      RECT  181.5 263.8 182.3 264.6 ;
      RECT  208.7 284.6 209.5 285.4 ;
      RECT  201.9 170.6 202.7 171.4 ;
      RECT  201.9 347.0 202.7 347.8 ;
      RECT  201.9 253.8 202.7 254.6 ;
      RECT  181.5 253.8 182.3 254.6 ;
      RECT  201.9 263.8 202.7 264.6 ;
      RECT  201.9 222.2 202.7 223.0 ;
      RECT  181.5 295.4 182.3 296.2 ;
      RECT  174.7 243.0 175.5 243.8 ;
      RECT  174.7 337.0 175.5 337.8 ;
      RECT  181.5 316.2 182.3 317.0 ;
      RECT  193.9 85.0 194.7 85.8 ;
      RECT  152.0 290.0 152.8 290.8 ;
      RECT  108.1 269.2 108.9 270.0 ;
      RECT  181.5 243.0 182.3 243.8 ;
      RECT  174.7 347.0 175.5 347.8 ;
      RECT  201.9 212.2 202.7 213.0 ;
      RECT  181.5 347.0 182.3 347.8 ;
      RECT  152.0 227.6 152.8 228.4 ;
      RECT  208.7 347.0 209.5 347.8 ;
      RECT  172.6 167.8 173.4 168.6 ;
      RECT  181.5 170.6 182.3 171.4 ;
      RECT  195.1 138.8 195.9 139.6 ;
      RECT  208.7 274.6 209.5 275.4 ;
      RECT  201.9 138.8 202.7 139.6 ;
      RECT  201.9 337.0 202.7 337.8 ;
      RECT  174.7 263.8 175.5 264.6 ;
      RECT  181.5 357.8 182.3 358.6 ;
      RECT  208.7 222.2 209.5 223.0 ;
      RECT  93.1 248.4 93.9 249.2 ;
      RECT  174.7 357.8 175.5 358.6 ;
      RECT  201.9 357.8 202.7 358.6 ;
      RECT  208.7 243.0 209.5 243.8 ;
      RECT  174.7 316.2 175.5 317.0 ;
      RECT  174.7 326.2 175.5 327.0 ;
      RECT  181.5 337.0 182.3 337.8 ;
      RECT  201.9 243.0 202.7 243.8 ;
      RECT  195.1 170.6 195.9 171.4 ;
      RECT  195.1 357.8 195.9 358.6 ;
      RECT  210.8 167.8 211.6 168.6 ;
      RECT  201.9 233.0 202.7 233.8 ;
      RECT  201.9 316.2 202.7 317.0 ;
      RECT  208.7 191.4 209.5 192.2 ;
      RECT  181.5 284.6 182.3 285.4 ;
      RECT  191.1 99.6 191.9 100.4 ;
      RECT  167.2 186.0 168.0 186.8 ;
      RECT  208.7 180.6 209.5 181.4 ;
      RECT  93.1 186.0 93.9 186.8 ;
      RECT  208.7 305.4 209.5 306.2 ;
      RECT  208.7 201.4 209.5 202.2 ;
      RECT  174.7 233.0 175.5 233.8 ;
      RECT  208.7 253.8 209.5 254.6 ;
      RECT  174.7 305.4 175.5 306.2 ;
      RECT  181.5 233.0 182.3 233.8 ;
      RECT  152.0 310.8 152.8 311.6 ;
      RECT  152.0 206.8 152.8 207.6 ;
      RECT  201.9 274.6 202.7 275.4 ;
      RECT  208.7 233.0 209.5 233.8 ;
      RECT  208.7 212.2 209.5 213.0 ;
      RECT  208.7 337.0 209.5 337.8 ;
      RECT  181.5 305.4 182.3 306.2 ;
      RECT  174.7 284.6 175.5 285.4 ;
      RECT  167.2 290.0 168.0 290.8 ;
      RECT  208.7 326.2 209.5 327.0 ;
      RECT  201.9 191.4 202.7 192.2 ;
      RECT  200.7 85.0 201.5 85.8 ;
      RECT  201.9 284.6 202.7 285.4 ;
      RECT  201.9 295.4 202.7 296.2 ;
      RECT  108.1 206.8 108.9 207.6 ;
      RECT  174.7 170.6 175.5 171.4 ;
      RECT  208.7 316.2 209.5 317.0 ;
      RECT  174.7 274.6 175.5 275.4 ;
      RECT  208.7 170.6 209.5 171.4 ;
      RECT  167.2 227.6 168.0 228.4 ;
      RECT  174.7 191.4 175.5 192.2 ;
      RECT  108.1 186.0 108.9 186.8 ;
      RECT  174.7 201.4 175.5 202.2 ;
      RECT  181.5 191.4 182.3 192.2 ;
      RECT  197.9 99.6 198.7 100.4 ;
      RECT  93.1 269.2 93.9 270.0 ;
      RECT  188.3 170.6 189.1 171.4 ;
      RECT  167.2 269.2 168.0 270.0 ;
      RECT  93.1 206.8 93.9 207.6 ;
      RECT  174.7 222.2 175.5 223.0 ;
      RECT  201.9 305.4 202.7 306.2 ;
      RECT  174.7 212.2 175.5 213.0 ;
      RECT  167.2 310.8 168.0 311.6 ;
      RECT  108.1 290.0 108.9 290.8 ;
      RECT  108.1 248.4 108.9 249.2 ;
      RECT  199.3 80.6 200.1 81.4 ;
      RECT  181.5 212.2 182.3 213.0 ;
      RECT  152.0 352.4 152.8 353.2 ;
      RECT  174.7 180.6 175.5 181.4 ;
      RECT  201.9 201.4 202.7 202.2 ;
      RECT  152.0 186.0 152.8 186.8 ;
      RECT  192.5 80.6 193.3 81.4 ;
      RECT  93.1 290.0 93.9 290.8 ;
      RECT  208.7 295.4 209.5 296.2 ;
      RECT  181.5 326.2 182.3 327.0 ;
      RECT  152.0 269.2 152.8 270.0 ;
      RECT  201.9 326.2 202.7 327.0 ;
      RECT  188.3 357.8 189.1 358.6 ;
      RECT  152.0 248.4 152.8 249.2 ;
      RECT  181.5 180.6 182.3 181.4 ;
      RECT  108.1 227.6 108.9 228.4 ;
      RECT  152.0 331.6 152.8 332.4 ;
      RECT  181.5 201.4 182.3 202.2 ;
      RECT  167.2 206.8 168.0 207.6 ;
      RECT  208.7 357.8 209.5 358.6 ;
      RECT  181.5 274.6 182.3 275.4 ;
      RECT  167.2 331.6 168.0 332.4 ;
      RECT  167.2 352.4 168.0 353.2 ;
      RECT  181.5 222.2 182.3 223.0 ;
      RECT  210.8 355.0 211.6 355.8 ;
      RECT  167.2 248.4 168.0 249.2 ;
      RECT  93.1 227.6 93.9 228.4 ;
      RECT  172.6 355.0 173.4 355.8 ;
      RECT  174.7 295.4 175.5 296.2 ;
      RECT  201.9 180.6 202.7 181.4 ;
      RECT  174.7 253.8 175.5 254.6 ;
      RECT  208.7 263.8 209.5 264.6 ;
      RECT  2.0 22.4 2.8 23.2 ;
      RECT  2.0 42.4 2.8 43.2 ;
      RECT  2.0 2.4 2.8 3.2 ;
      RECT  24.0 224.0 23.2 224.8 ;
      RECT  24.0 302.4 23.2 303.2 ;
      RECT  10.8 263.2 10.0 264.0 ;
      RECT  24.0 184.8 23.2 185.6 ;
      RECT  10.8 184.8 10.0 185.6 ;
      RECT  10.8 341.6 10.0 342.4 ;
      RECT  24.0 263.2 23.2 264.0 ;
      RECT  10.8 224.0 10.0 224.8 ;
      RECT  24.0 341.6 23.2 342.4 ;
      RECT  10.8 302.4 10.0 303.2 ;
      RECT  10.8 322.0 10.0 322.8 ;
      RECT  10.8 165.2 10.0 166.0 ;
      RECT  10.8 243.6 10.0 244.4 ;
      RECT  24.0 204.4 23.2 205.2 ;
      RECT  10.8 282.8 10.0 283.6 ;
      RECT  24.0 322.0 23.2 322.8 ;
      RECT  24.0 243.6 23.2 244.4 ;
      RECT  10.8 204.4 10.0 205.2 ;
      RECT  24.0 282.8 23.2 283.6 ;
      RECT  24.0 165.2 23.2 166.0 ;
      RECT  23.2 341.6 24.0 342.4 ;
      RECT  77.6 62.4 78.4 63.2 ;
      RECT  77.6 102.4 78.4 103.2 ;
      RECT  23.2 302.4 24.0 303.2 ;
      RECT  77.6 142.4 78.4 143.2 ;
      RECT  10.0 224.0 10.8 224.8 ;
      RECT  10.0 302.4 10.8 303.2 ;
      RECT  10.0 263.2 10.8 264.0 ;
      RECT  23.2 184.8 24.0 185.6 ;
      RECT  77.6 22.4 78.4 23.2 ;
      RECT  10.0 341.6 10.8 342.4 ;
      RECT  2.0 22.4 2.8 23.2 ;
      RECT  10.0 184.8 10.8 185.6 ;
      RECT  23.2 263.2 24.0 264.0 ;
      RECT  23.2 224.0 24.0 224.8 ;
      RECT  23.2 322.0 24.0 322.8 ;
      RECT  10.0 243.6 10.8 244.4 ;
      RECT  2.0 2.4 2.8 3.2 ;
      RECT  10.0 282.8 10.8 283.6 ;
      RECT  23.2 243.6 24.0 244.4 ;
      RECT  10.0 204.4 10.8 205.2 ;
      RECT  23.2 165.2 24.0 166.0 ;
      RECT  77.6 162.4 78.4 163.2 ;
      RECT  77.6 2.4 78.4 3.2 ;
      RECT  77.6 42.4 78.4 43.2 ;
      RECT  77.6 122.4 78.4 123.2 ;
      RECT  10.0 322.0 10.8 322.8 ;
      RECT  10.0 165.2 10.8 166.0 ;
      RECT  23.2 282.8 24.0 283.6 ;
      RECT  23.2 204.4 24.0 205.2 ;
      RECT  2.0 42.4 2.8 43.2 ;
      RECT  77.6 82.4 78.4 83.2 ;
      RECT  57.6 347.9 79.4 348.5 ;
      RECT  68.1 404.4 68.9 405.2 ;
      RECT  68.1 364.4 68.9 365.2 ;
      RECT  68.1 424.4 68.9 425.2 ;
      RECT  68.1 344.4 68.9 345.2 ;
      RECT  68.1 384.4 68.9 385.2 ;
      RECT  101.2 5.9 144.8 6.5 ;
      RECT  133.5 22.4 134.3 23.2 ;
      RECT  111.7 22.4 112.5 23.2 ;
      RECT  111.7 2.4 112.5 3.2 ;
      RECT  133.5 2.4 134.3 3.2 ;
   LAYER  metal4 ;
   END
   END    sram_2_16_1_scn4m_subm
END    LIBRARY
