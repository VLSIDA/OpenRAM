magic
tech sky130A
magscale 1 2
timestamp 1595931502
<< checkpaint >>
rect -1260 -1286 2274 1716
<< scnmos >>
rect 60 0 90 400
rect 168 0 198 400
rect 276 0 306 400
rect 384 0 414 400
rect 492 0 522 400
rect 600 0 630 400
rect 708 0 738 400
rect 816 0 846 400
rect 924 0 954 400
<< ndiff >>
rect 0 0 60 400
rect 90 0 168 400
rect 198 0 276 400
rect 306 0 384 400
rect 414 0 492 400
rect 522 0 600 400
rect 630 0 708 400
rect 738 0 816 400
rect 846 0 924 400
rect 954 0 1014 400
<< poly >>
rect 60 426 954 456
rect 60 400 90 426
rect 168 400 198 426
rect 276 400 306 426
rect 384 400 414 426
rect 492 400 522 426
rect 600 400 630 426
rect 708 400 738 426
rect 816 400 846 426
rect 924 400 954 426
rect 60 -26 90 0
rect 168 -26 198 0
rect 276 -26 306 0
rect 384 -26 414 0
rect 492 -26 522 0
rect 600 -26 630 0
rect 708 -26 738 0
rect 816 -26 846 0
rect 924 -26 954 0
<< locali >>
rect 112 267 1006 301
rect 8 167 42 233
rect 112 200 146 267
rect 220 167 254 233
rect 328 200 362 267
rect 436 167 470 233
rect 544 200 578 267
rect 652 167 686 233
rect 760 200 794 267
rect 868 167 902 233
rect 972 200 1006 267
use contact_17  contact_17_0
timestamp 1595931502
transform 1 0 964 0 1 167
box 0 0 50 66
use contact_17  contact_17_1
timestamp 1595931502
transform 1 0 860 0 1 167
box 0 0 50 66
use contact_17  contact_17_2
timestamp 1595931502
transform 1 0 752 0 1 167
box 0 0 50 66
use contact_17  contact_17_3
timestamp 1595931502
transform 1 0 644 0 1 167
box 0 0 50 66
use contact_17  contact_17_4
timestamp 1595931502
transform 1 0 536 0 1 167
box 0 0 50 66
use contact_17  contact_17_5
timestamp 1595931502
transform 1 0 428 0 1 167
box 0 0 50 66
use contact_17  contact_17_6
timestamp 1595931502
transform 1 0 320 0 1 167
box 0 0 50 66
use contact_17  contact_17_7
timestamp 1595931502
transform 1 0 212 0 1 167
box 0 0 50 66
use contact_17  contact_17_8
timestamp 1595931502
transform 1 0 104 0 1 167
box 0 0 50 66
use contact_17  contact_17_9
timestamp 1595931502
transform 1 0 0 0 1 167
box 0 0 50 66
<< labels >>
rlabel poly s 507 441 507 441 4 G
rlabel corelocali s 669 200 669 200 4 S
rlabel corelocali s 453 200 453 200 4 S
rlabel corelocali s 25 200 25 200 4 S
rlabel corelocali s 885 200 885 200 4 S
rlabel corelocali s 237 200 237 200 4 S
rlabel corelocali s 559 284 559 284 4 D
<< properties >>
string FIXED_BBOX -25 -26 1039 426
<< end >>
