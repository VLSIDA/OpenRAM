magic
tech sky130A
magscale 1 2
timestamp 1595931502
<< checkpaint >>
rect -1260 -1286 1626 1716
<< scnmos >>
rect 60 0 90 400
rect 168 0 198 400
rect 276 0 306 400
<< ndiff >>
rect 0 0 60 400
rect 90 0 168 400
rect 198 0 276 400
rect 306 0 366 400
<< poly >>
rect 60 426 306 456
rect 60 400 90 426
rect 168 400 198 426
rect 276 400 306 426
rect 60 -26 90 0
rect 168 -26 198 0
rect 276 -26 306 0
<< locali >>
rect 112 267 358 301
rect 8 167 42 233
rect 112 200 146 267
rect 220 167 254 233
rect 324 200 358 267
use contact_17  contact_17_3
timestamp 1595931502
transform 1 0 0 0 1 167
box 0 0 50 66
use contact_17  contact_17_2
timestamp 1595931502
transform 1 0 104 0 1 167
box 0 0 50 66
use contact_17  contact_17_1
timestamp 1595931502
transform 1 0 212 0 1 167
box 0 0 50 66
use contact_17  contact_17_0
timestamp 1595931502
transform 1 0 316 0 1 167
box 0 0 50 66
<< labels >>
rlabel poly s 183 441 183 441 4 G
rlabel corelocali s 25 200 25 200 4 S
rlabel corelocali s 237 200 237 200 4 S
rlabel corelocali s 235 284 235 284 4 D
<< properties >>
string FIXED_BBOX -25 -26 391 426
<< end >>
