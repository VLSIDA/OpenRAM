magic
tech sky130A
magscale 1 2
timestamp 1595931502
<< checkpaint >>
rect -1296 -1277 3638 2731
<< nwell >>
rect -36 679 2378 1471
<< locali >>
rect 0 1397 2342 1431
rect 64 636 98 702
rect 179 664 449 698
rect 551 690 815 724
rect 1040 690 1295 724
rect 1827 690 1861 724
rect 551 681 585 690
rect 0 -17 2342 17
use pinv_4  pinv_4_0
timestamp 1595931502
transform 1 0 0 0 1 0
box -36 -17 404 1471
use pinv_3  pinv_3_0
timestamp 1595931502
transform 1 0 368 0 1 0
box -36 -17 402 1471
use pinv_6  pinv_6_0
timestamp 1595931502
transform 1 0 1214 0 1 0
box -36 -17 1164 1471
use pinv_5  pinv_5_0
timestamp 1595931502
transform 1 0 734 0 1 0
box -36 -17 516 1471
<< labels >>
rlabel corelocali s 1171 0 1171 0 4 gnd
rlabel corelocali s 1844 707 1844 707 4 Z
rlabel corelocali s 1171 1414 1171 1414 4 vdd
rlabel corelocali s 81 669 81 669 4 A
<< properties >>
string FIXED_BBOX 0 0 2342 1414
<< end >>
