**************************************************
* OpenRAM generated memory.
* Words: 2048
* Data bits: 32
* Banks: 1
* Column mux: 4:1
**************************************************

* ptx M{0} {1} nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.0225p ad=0.0225p

* ptx M{0} {1} pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p

.SUBCKT pnand2_1 A B Z vdd gnd
Mpnand2_pmos1 vdd A Z vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpnand2_pmos2 Z B vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpnand2_nmos1 Z B net1 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.0225p ad=0.0225p
Mpnand2_nmos2 net1 A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.0225p ad=0.0225p
.ENDS pnand2_1

.SUBCKT pnand3_1 A B C Z vdd gnd
Mpnand3_pmos1 vdd A Z vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpnand3_pmos2 Z B vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpnand3_pmos3 Z C vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpnand3_nmos1 Z C net1 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.0225p ad=0.0225p
Mpnand3_nmos2 net1 B net2 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.0225p ad=0.0225p
Mpnand3_nmos3 net2 A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.0225p ad=0.0225p
.ENDS pnand3_1

* ptx M{0} {1} nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01125p ad=0.01125p

* ptx M{0} {1} pmos_vtg m=1 w=0.405u l=0.05u pd=0.91u ps=0.91u as=0.050625p ad=0.050625p

.SUBCKT pnor2_1 A B Z vdd gnd
Mpnor2_pmos1 vdd A net1 vdd pmos_vtg m=1 w=0.405u l=0.05u pd=0.91u ps=0.91u as=0.050625p ad=0.050625p
Mpnor2_pmos2 net1 B Z vdd pmos_vtg m=1 w=0.405u l=0.05u pd=0.91u ps=0.91u as=0.050625p ad=0.050625p
Mpnor2_nmos1 Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01125p ad=0.01125p
Mpnor2_nmos2 Z B gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01125p ad=0.01125p
.ENDS pnor2_1

.SUBCKT pinv_1 A Z vdd gnd
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01125p ad=0.01125p
.ENDS pinv_1

* ptx M{0} {1} nmos_vtg m=2 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01125p ad=0.01125p

* ptx M{0} {1} pmos_vtg m=2 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p

.SUBCKT pinv_2 A Z vdd gnd
Mpinv_pmos Z A vdd vdd pmos_vtg m=2 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpinv_nmos Z A gnd gnd nmos_vtg m=2 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01125p ad=0.01125p
.ENDS pinv_2

* ptx M{0} {1} nmos_vtg m=3 w=0.12u l=0.05u pd=0.34u ps=0.34u as=0.015p ad=0.015p

* ptx M{0} {1} pmos_vtg m=3 w=0.36u l=0.05u pd=0.82u ps=0.82u as=0.045p ad=0.045p

.SUBCKT pinv_3 A Z vdd gnd
Mpinv_pmos Z A vdd vdd pmos_vtg m=3 w=0.36u l=0.05u pd=0.82u ps=0.82u as=0.045p ad=0.045p
Mpinv_nmos Z A gnd gnd nmos_vtg m=3 w=0.12u l=0.05u pd=0.34u ps=0.34u as=0.015p ad=0.015p
.ENDS pinv_3

* ptx M{0} {1} nmos_vtg m=6 w=0.12u l=0.05u pd=0.34u ps=0.34u as=0.015p ad=0.015p

* ptx M{0} {1} pmos_vtg m=6 w=0.36u l=0.05u pd=0.82u ps=0.82u as=0.045p ad=0.045p

.SUBCKT pinv_4 A Z vdd gnd
Mpinv_pmos Z A vdd vdd pmos_vtg m=6 w=0.36u l=0.05u pd=0.82u ps=0.82u as=0.045p ad=0.045p
Mpinv_nmos Z A gnd gnd nmos_vtg m=6 w=0.12u l=0.05u pd=0.34u ps=0.34u as=0.015p ad=0.015p
.ENDS pinv_4

* ptx M{0} {1} nmos_vtg m=12 w=0.12u l=0.05u pd=0.34u ps=0.34u as=0.015p ad=0.015p

* ptx M{0} {1} pmos_vtg m=12 w=0.36u l=0.05u pd=0.82u ps=0.82u as=0.045p ad=0.045p

.SUBCKT pinv_5 A Z vdd gnd
Mpinv_pmos Z A vdd vdd pmos_vtg m=12 w=0.36u l=0.05u pd=0.82u ps=0.82u as=0.045p ad=0.045p
Mpinv_nmos Z A gnd gnd nmos_vtg m=12 w=0.12u l=0.05u pd=0.34u ps=0.34u as=0.015p ad=0.015p
.ENDS pinv_5
*master-slave flip-flop with both output and inverted ouput

.SUBCKT ms_flop din dout dout_bar clk vdd gnd
xmaster din mout mout_bar clk clk_bar vdd gnd dlatch
xslave mout_bar dout_bar dout clk_bar clk_nn vdd gnd dlatch
.ENDS flop

.SUBCKT dlatch din dout dout_bar clk clk_bar vdd gnd
*clk inverter
mPff1 clk_bar clk vdd vdd PMOS_VTG W=180.0n L=50n m=1
mNff1 clk_bar clk gnd gnd NMOS_VTG W=90n L=50n m=1

*transmission gate 1
mtmP1 din clk int1 vdd PMOS_VTG W=180.0n L=50n m=1
mtmN1 din clk_bar int1 gnd NMOS_VTG W=90n L=50n m=1

*foward inverter
mPff3 dout_bar int1 vdd vdd PMOS_VTG W=180.0n L=50n m=1
mNff3 dout_bar int1 gnd gnd NMOS_VTG W=90n L=50n m=1

*backward inverter
mPff4 dout dout_bar vdd vdd PMOS_VTG W=180.0n L=50n m=1
mNf4 dout dout_bar gnd gnd NMOS_VTG W=90n L=50n m=1

*transmission gate 2
mtmP2 int1 clk_bar dout vdd PMOS_VTG W=180.0n L=50n m=1
mtmN2 int1 clk dout gnd NMOS_VTG W=90n L=50n m=1
.ENDS dlatch


.SUBCKT msf_control din[0] din[1] din[2] dout[0] dout_bar[0] dout[1] dout_bar[1] dout[2] dout_bar[2] clk vdd gnd
XXdff0 din[0] dout[0] dout_bar[0] clk vdd gnd ms_flop
XXdff1 din[1] dout[1] dout_bar[1] clk vdd gnd ms_flop
XXdff2 din[2] dout[2] dout_bar[2] clk vdd gnd ms_flop
.ENDS msf_control

.SUBCKT replica_cell_6t bl br wl vdd gnd
MM3 bl wl gnd gnd NMOS_VTG W=135.00n L=50n
MM2 br wl net4 gnd NMOS_VTG W=135.00n L=50n
MM1 gnd net4 gnd gnd NMOS_VTG W=205.00n L=50n
MM0 net4 gnd gnd gnd NMOS_VTG W=205.00n L=50n
MM5 gnd net4 vdd vdd PMOS_VTG W=90n L=50n
MM4 net4 gnd vdd vdd PMOS_VTG W=90n L=50n
.ENDS replica_cell_6t


.SUBCKT cell_6t bl br wl vdd gnd
MM3 bl wl net10 gnd NMOS_VTG W=135.00n L=50n
MM2 br wl net4 gnd NMOS_VTG W=135.00n L=50n
MM1 net10 net4 gnd gnd NMOS_VTG W=205.00n L=50n
MM0 net4 net10 gnd gnd NMOS_VTG W=205.00n L=50n
MM5 net10 net4 vdd vdd PMOS_VTG W=90n L=50n
MM4 net4 net10 vdd vdd PMOS_VTG W=90n L=50n
.ENDS cell_6t


.SUBCKT bitline_load bl[0] br[0] wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] vdd gnd
Xbit_r0_c0 bl[0] br[0] wl[0] vdd gnd cell_6t
Xbit_r1_c0 bl[0] br[0] wl[1] vdd gnd cell_6t
Xbit_r2_c0 bl[0] br[0] wl[2] vdd gnd cell_6t
Xbit_r3_c0 bl[0] br[0] wl[3] vdd gnd cell_6t
Xbit_r4_c0 bl[0] br[0] wl[4] vdd gnd cell_6t
Xbit_r5_c0 bl[0] br[0] wl[5] vdd gnd cell_6t
Xbit_r6_c0 bl[0] br[0] wl[6] vdd gnd cell_6t
Xbit_r7_c0 bl[0] br[0] wl[7] vdd gnd cell_6t
Xbit_r8_c0 bl[0] br[0] wl[8] vdd gnd cell_6t
Xbit_r9_c0 bl[0] br[0] wl[9] vdd gnd cell_6t
Xbit_r10_c0 bl[0] br[0] wl[10] vdd gnd cell_6t
Xbit_r11_c0 bl[0] br[0] wl[11] vdd gnd cell_6t
Xbit_r12_c0 bl[0] br[0] wl[12] vdd gnd cell_6t
Xbit_r13_c0 bl[0] br[0] wl[13] vdd gnd cell_6t
Xbit_r14_c0 bl[0] br[0] wl[14] vdd gnd cell_6t
Xbit_r15_c0 bl[0] br[0] wl[15] vdd gnd cell_6t
Xbit_r16_c0 bl[0] br[0] wl[16] vdd gnd cell_6t
Xbit_r17_c0 bl[0] br[0] wl[17] vdd gnd cell_6t
Xbit_r18_c0 bl[0] br[0] wl[18] vdd gnd cell_6t
Xbit_r19_c0 bl[0] br[0] wl[19] vdd gnd cell_6t
Xbit_r20_c0 bl[0] br[0] wl[20] vdd gnd cell_6t
Xbit_r21_c0 bl[0] br[0] wl[21] vdd gnd cell_6t
Xbit_r22_c0 bl[0] br[0] wl[22] vdd gnd cell_6t
Xbit_r23_c0 bl[0] br[0] wl[23] vdd gnd cell_6t
Xbit_r24_c0 bl[0] br[0] wl[24] vdd gnd cell_6t
Xbit_r25_c0 bl[0] br[0] wl[25] vdd gnd cell_6t
Xbit_r26_c0 bl[0] br[0] wl[26] vdd gnd cell_6t
Xbit_r27_c0 bl[0] br[0] wl[27] vdd gnd cell_6t
Xbit_r28_c0 bl[0] br[0] wl[28] vdd gnd cell_6t
Xbit_r29_c0 bl[0] br[0] wl[29] vdd gnd cell_6t
Xbit_r30_c0 bl[0] br[0] wl[30] vdd gnd cell_6t
Xbit_r31_c0 bl[0] br[0] wl[31] vdd gnd cell_6t
Xbit_r32_c0 bl[0] br[0] wl[32] vdd gnd cell_6t
Xbit_r33_c0 bl[0] br[0] wl[33] vdd gnd cell_6t
Xbit_r34_c0 bl[0] br[0] wl[34] vdd gnd cell_6t
Xbit_r35_c0 bl[0] br[0] wl[35] vdd gnd cell_6t
Xbit_r36_c0 bl[0] br[0] wl[36] vdd gnd cell_6t
Xbit_r37_c0 bl[0] br[0] wl[37] vdd gnd cell_6t
Xbit_r38_c0 bl[0] br[0] wl[38] vdd gnd cell_6t
Xbit_r39_c0 bl[0] br[0] wl[39] vdd gnd cell_6t
Xbit_r40_c0 bl[0] br[0] wl[40] vdd gnd cell_6t
Xbit_r41_c0 bl[0] br[0] wl[41] vdd gnd cell_6t
Xbit_r42_c0 bl[0] br[0] wl[42] vdd gnd cell_6t
Xbit_r43_c0 bl[0] br[0] wl[43] vdd gnd cell_6t
Xbit_r44_c0 bl[0] br[0] wl[44] vdd gnd cell_6t
Xbit_r45_c0 bl[0] br[0] wl[45] vdd gnd cell_6t
Xbit_r46_c0 bl[0] br[0] wl[46] vdd gnd cell_6t
Xbit_r47_c0 bl[0] br[0] wl[47] vdd gnd cell_6t
Xbit_r48_c0 bl[0] br[0] wl[48] vdd gnd cell_6t
Xbit_r49_c0 bl[0] br[0] wl[49] vdd gnd cell_6t
Xbit_r50_c0 bl[0] br[0] wl[50] vdd gnd cell_6t
Xbit_r51_c0 bl[0] br[0] wl[51] vdd gnd cell_6t
Xbit_r52_c0 bl[0] br[0] wl[52] vdd gnd cell_6t
Xbit_r53_c0 bl[0] br[0] wl[53] vdd gnd cell_6t
Xbit_r54_c0 bl[0] br[0] wl[54] vdd gnd cell_6t
Xbit_r55_c0 bl[0] br[0] wl[55] vdd gnd cell_6t
Xbit_r56_c0 bl[0] br[0] wl[56] vdd gnd cell_6t
Xbit_r57_c0 bl[0] br[0] wl[57] vdd gnd cell_6t
Xbit_r58_c0 bl[0] br[0] wl[58] vdd gnd cell_6t
Xbit_r59_c0 bl[0] br[0] wl[59] vdd gnd cell_6t
Xbit_r60_c0 bl[0] br[0] wl[60] vdd gnd cell_6t
Xbit_r61_c0 bl[0] br[0] wl[61] vdd gnd cell_6t
Xbit_r62_c0 bl[0] br[0] wl[62] vdd gnd cell_6t
Xbit_r63_c0 bl[0] br[0] wl[63] vdd gnd cell_6t
Xbit_r64_c0 bl[0] br[0] wl[64] vdd gnd cell_6t
Xbit_r65_c0 bl[0] br[0] wl[65] vdd gnd cell_6t
Xbit_r66_c0 bl[0] br[0] wl[66] vdd gnd cell_6t
Xbit_r67_c0 bl[0] br[0] wl[67] vdd gnd cell_6t
Xbit_r68_c0 bl[0] br[0] wl[68] vdd gnd cell_6t
Xbit_r69_c0 bl[0] br[0] wl[69] vdd gnd cell_6t
Xbit_r70_c0 bl[0] br[0] wl[70] vdd gnd cell_6t
Xbit_r71_c0 bl[0] br[0] wl[71] vdd gnd cell_6t
Xbit_r72_c0 bl[0] br[0] wl[72] vdd gnd cell_6t
Xbit_r73_c0 bl[0] br[0] wl[73] vdd gnd cell_6t
Xbit_r74_c0 bl[0] br[0] wl[74] vdd gnd cell_6t
Xbit_r75_c0 bl[0] br[0] wl[75] vdd gnd cell_6t
Xbit_r76_c0 bl[0] br[0] wl[76] vdd gnd cell_6t
Xbit_r77_c0 bl[0] br[0] wl[77] vdd gnd cell_6t
Xbit_r78_c0 bl[0] br[0] wl[78] vdd gnd cell_6t
Xbit_r79_c0 bl[0] br[0] wl[79] vdd gnd cell_6t
Xbit_r80_c0 bl[0] br[0] wl[80] vdd gnd cell_6t
Xbit_r81_c0 bl[0] br[0] wl[81] vdd gnd cell_6t
Xbit_r82_c0 bl[0] br[0] wl[82] vdd gnd cell_6t
Xbit_r83_c0 bl[0] br[0] wl[83] vdd gnd cell_6t
Xbit_r84_c0 bl[0] br[0] wl[84] vdd gnd cell_6t
Xbit_r85_c0 bl[0] br[0] wl[85] vdd gnd cell_6t
Xbit_r86_c0 bl[0] br[0] wl[86] vdd gnd cell_6t
Xbit_r87_c0 bl[0] br[0] wl[87] vdd gnd cell_6t
Xbit_r88_c0 bl[0] br[0] wl[88] vdd gnd cell_6t
Xbit_r89_c0 bl[0] br[0] wl[89] vdd gnd cell_6t
Xbit_r90_c0 bl[0] br[0] wl[90] vdd gnd cell_6t
Xbit_r91_c0 bl[0] br[0] wl[91] vdd gnd cell_6t
Xbit_r92_c0 bl[0] br[0] wl[92] vdd gnd cell_6t
Xbit_r93_c0 bl[0] br[0] wl[93] vdd gnd cell_6t
Xbit_r94_c0 bl[0] br[0] wl[94] vdd gnd cell_6t
Xbit_r95_c0 bl[0] br[0] wl[95] vdd gnd cell_6t
Xbit_r96_c0 bl[0] br[0] wl[96] vdd gnd cell_6t
Xbit_r97_c0 bl[0] br[0] wl[97] vdd gnd cell_6t
Xbit_r98_c0 bl[0] br[0] wl[98] vdd gnd cell_6t
Xbit_r99_c0 bl[0] br[0] wl[99] vdd gnd cell_6t
Xbit_r100_c0 bl[0] br[0] wl[100] vdd gnd cell_6t
Xbit_r101_c0 bl[0] br[0] wl[101] vdd gnd cell_6t
Xbit_r102_c0 bl[0] br[0] wl[102] vdd gnd cell_6t
.ENDS bitline_load

.SUBCKT pinv_6 A Z vdd gnd
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01125p ad=0.01125p
.ENDS pinv_6

.SUBCKT delay_chain in out vdd gnd
Xdinv0 in s1 vdd gnd pinv_6
Xdinv1 s1 s2n1 vdd gnd pinv_6
Xdinv2 s1 s2n2 vdd gnd pinv_6
Xdinv3 s1 s2 vdd gnd pinv_6
Xdinv4 s2 s3n1 vdd gnd pinv_6
Xdinv5 s2 s3n2 vdd gnd pinv_6
Xdinv6 s2 s3 vdd gnd pinv_6
Xdinv7 s3 s4n1 vdd gnd pinv_6
Xdinv8 s3 s4n2 vdd gnd pinv_6
Xdinv9 s3 s4 vdd gnd pinv_6
Xdinv10 s4 s5n1 vdd gnd pinv_6
Xdinv11 s4 s5n2 vdd gnd pinv_6
Xdinv12 s4 out vdd gnd pinv_6
.ENDS delay_chain

.SUBCKT pinv_7 A Z vdd gnd
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01125p ad=0.01125p
.ENDS pinv_7

* ptx M{0} {1} pmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01125p ad=0.01125p

.SUBCKT replica_bitline en out vdd gnd
Xrbl_inv bl[0] out vdd gnd pinv_7
Mrbl_access_tx vdd delayed_en bl[0] vdd pmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01125p ad=0.01125p
Xdelay_chain en delayed_en vdd gnd delay_chain
Xbitcell bl[0] br[0] delayed_en vdd gnd replica_cell_6t
Xload bl[0] br[0] gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd gnd vdd gnd bitline_load
.ENDS replica_bitline

.SUBCKT control_logic csb web oeb clk s_en w_en tri_en tri_en_bar clk_bar clk_buf vdd gnd
Xmsf_control oeb csb web oe_bar oe cs_bar cs we_bar we clk_buf vdd gnd msf_control
Xinv_clk1_bar clk clk1_bar vdd gnd pinv_2
Xinv_clk2 clk1_bar clk2 vdd gnd pinv_3
Xinv_clk_bar clk2 clk_bar vdd gnd pinv_4
Xinv_clk_buf clk_bar clk_buf vdd gnd pinv_5
Xnand3_rblk_bar clk_bar oe cs rblk_bar vdd gnd pnand3_1
Xinv_rblk rblk_bar rblk vdd gnd pinv_1
Xnor2_tri_en clk_buf oe_bar tri_en vdd gnd pnor2_1
Xnand2_tri_en clk_bar oe tri_en_bar vdd gnd pnand2_1
Xinv_s_en pre_s_en_bar s_en vdd gnd pinv_1
Xinv_pre_s_en_bar pre_s_en pre_s_en_bar vdd gnd pinv_1
Xnand3_w_en_bar clk_bar cs we w_en_bar vdd gnd pnand3_1
Xinv_pre_w_en w_en_bar pre_w_en vdd gnd pinv_1
Xinv_pre_w_en_bar pre_w_en pre_w_en_bar vdd gnd pinv_1
Xinv_w_en2 pre_w_en_bar w_en vdd gnd pinv_1
Xreplica_bitline rblk pre_s_en vdd gnd replica_bitline
.ENDS control_logic

.SUBCKT bitcell_array bl[0] br[0] bl[1] br[1] bl[2] br[2] bl[3] br[3] bl[4] br[4] bl[5] br[5] bl[6] br[6] bl[7] br[7] bl[8] br[8] bl[9] br[9] bl[10] br[10] bl[11] br[11] bl[12] br[12] bl[13] br[13] bl[14] br[14] bl[15] br[15] bl[16] br[16] bl[17] br[17] bl[18] br[18] bl[19] br[19] bl[20] br[20] bl[21] br[21] bl[22] br[22] bl[23] br[23] bl[24] br[24] bl[25] br[25] bl[26] br[26] bl[27] br[27] bl[28] br[28] bl[29] br[29] bl[30] br[30] bl[31] br[31] bl[32] br[32] bl[33] br[33] bl[34] br[34] bl[35] br[35] bl[36] br[36] bl[37] br[37] bl[38] br[38] bl[39] br[39] bl[40] br[40] bl[41] br[41] bl[42] br[42] bl[43] br[43] bl[44] br[44] bl[45] br[45] bl[46] br[46] bl[47] br[47] bl[48] br[48] bl[49] br[49] bl[50] br[50] bl[51] br[51] bl[52] br[52] bl[53] br[53] bl[54] br[54] bl[55] br[55] bl[56] br[56] bl[57] br[57] bl[58] br[58] bl[59] br[59] bl[60] br[60] bl[61] br[61] bl[62] br[62] bl[63] br[63] bl[64] br[64] bl[65] br[65] bl[66] br[66] bl[67] br[67] bl[68] br[68] bl[69] br[69] bl[70] br[70] bl[71] br[71] bl[72] br[72] bl[73] br[73] bl[74] br[74] bl[75] br[75] bl[76] br[76] bl[77] br[77] bl[78] br[78] bl[79] br[79] bl[80] br[80] bl[81] br[81] bl[82] br[82] bl[83] br[83] bl[84] br[84] bl[85] br[85] bl[86] br[86] bl[87] br[87] bl[88] br[88] bl[89] br[89] bl[90] br[90] bl[91] br[91] bl[92] br[92] bl[93] br[93] bl[94] br[94] bl[95] br[95] bl[96] br[96] bl[97] br[97] bl[98] br[98] bl[99] br[99] bl[100] br[100] bl[101] br[101] bl[102] br[102] bl[103] br[103] bl[104] br[104] bl[105] br[105] bl[106] br[106] bl[107] br[107] bl[108] br[108] bl[109] br[109] bl[110] br[110] bl[111] br[111] bl[112] br[112] bl[113] br[113] bl[114] br[114] bl[115] br[115] bl[116] br[116] bl[117] br[117] bl[118] br[118] bl[119] br[119] bl[120] br[120] bl[121] br[121] bl[122] br[122] bl[123] br[123] bl[124] br[124] bl[125] br[125] bl[126] br[126] bl[127] br[127] wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] wl[128] wl[129] wl[130] wl[131] wl[132] wl[133] wl[134] wl[135] wl[136] wl[137] wl[138] wl[139] wl[140] wl[141] wl[142] wl[143] wl[144] wl[145] wl[146] wl[147] wl[148] wl[149] wl[150] wl[151] wl[152] wl[153] wl[154] wl[155] wl[156] wl[157] wl[158] wl[159] wl[160] wl[161] wl[162] wl[163] wl[164] wl[165] wl[166] wl[167] wl[168] wl[169] wl[170] wl[171] wl[172] wl[173] wl[174] wl[175] wl[176] wl[177] wl[178] wl[179] wl[180] wl[181] wl[182] wl[183] wl[184] wl[185] wl[186] wl[187] wl[188] wl[189] wl[190] wl[191] wl[192] wl[193] wl[194] wl[195] wl[196] wl[197] wl[198] wl[199] wl[200] wl[201] wl[202] wl[203] wl[204] wl[205] wl[206] wl[207] wl[208] wl[209] wl[210] wl[211] wl[212] wl[213] wl[214] wl[215] wl[216] wl[217] wl[218] wl[219] wl[220] wl[221] wl[222] wl[223] wl[224] wl[225] wl[226] wl[227] wl[228] wl[229] wl[230] wl[231] wl[232] wl[233] wl[234] wl[235] wl[236] wl[237] wl[238] wl[239] wl[240] wl[241] wl[242] wl[243] wl[244] wl[245] wl[246] wl[247] wl[248] wl[249] wl[250] wl[251] wl[252] wl[253] wl[254] wl[255] wl[256] wl[257] wl[258] wl[259] wl[260] wl[261] wl[262] wl[263] wl[264] wl[265] wl[266] wl[267] wl[268] wl[269] wl[270] wl[271] wl[272] wl[273] wl[274] wl[275] wl[276] wl[277] wl[278] wl[279] wl[280] wl[281] wl[282] wl[283] wl[284] wl[285] wl[286] wl[287] wl[288] wl[289] wl[290] wl[291] wl[292] wl[293] wl[294] wl[295] wl[296] wl[297] wl[298] wl[299] wl[300] wl[301] wl[302] wl[303] wl[304] wl[305] wl[306] wl[307] wl[308] wl[309] wl[310] wl[311] wl[312] wl[313] wl[314] wl[315] wl[316] wl[317] wl[318] wl[319] wl[320] wl[321] wl[322] wl[323] wl[324] wl[325] wl[326] wl[327] wl[328] wl[329] wl[330] wl[331] wl[332] wl[333] wl[334] wl[335] wl[336] wl[337] wl[338] wl[339] wl[340] wl[341] wl[342] wl[343] wl[344] wl[345] wl[346] wl[347] wl[348] wl[349] wl[350] wl[351] wl[352] wl[353] wl[354] wl[355] wl[356] wl[357] wl[358] wl[359] wl[360] wl[361] wl[362] wl[363] wl[364] wl[365] wl[366] wl[367] wl[368] wl[369] wl[370] wl[371] wl[372] wl[373] wl[374] wl[375] wl[376] wl[377] wl[378] wl[379] wl[380] wl[381] wl[382] wl[383] wl[384] wl[385] wl[386] wl[387] wl[388] wl[389] wl[390] wl[391] wl[392] wl[393] wl[394] wl[395] wl[396] wl[397] wl[398] wl[399] wl[400] wl[401] wl[402] wl[403] wl[404] wl[405] wl[406] wl[407] wl[408] wl[409] wl[410] wl[411] wl[412] wl[413] wl[414] wl[415] wl[416] wl[417] wl[418] wl[419] wl[420] wl[421] wl[422] wl[423] wl[424] wl[425] wl[426] wl[427] wl[428] wl[429] wl[430] wl[431] wl[432] wl[433] wl[434] wl[435] wl[436] wl[437] wl[438] wl[439] wl[440] wl[441] wl[442] wl[443] wl[444] wl[445] wl[446] wl[447] wl[448] wl[449] wl[450] wl[451] wl[452] wl[453] wl[454] wl[455] wl[456] wl[457] wl[458] wl[459] wl[460] wl[461] wl[462] wl[463] wl[464] wl[465] wl[466] wl[467] wl[468] wl[469] wl[470] wl[471] wl[472] wl[473] wl[474] wl[475] wl[476] wl[477] wl[478] wl[479] wl[480] wl[481] wl[482] wl[483] wl[484] wl[485] wl[486] wl[487] wl[488] wl[489] wl[490] wl[491] wl[492] wl[493] wl[494] wl[495] wl[496] wl[497] wl[498] wl[499] wl[500] wl[501] wl[502] wl[503] wl[504] wl[505] wl[506] wl[507] wl[508] wl[509] wl[510] wl[511] vdd gnd
Xbit_r0_c0 bl[0] br[0] wl[0] vdd gnd cell_6t
Xbit_r1_c0 bl[0] br[0] wl[1] vdd gnd cell_6t
Xbit_r2_c0 bl[0] br[0] wl[2] vdd gnd cell_6t
Xbit_r3_c0 bl[0] br[0] wl[3] vdd gnd cell_6t
Xbit_r4_c0 bl[0] br[0] wl[4] vdd gnd cell_6t
Xbit_r5_c0 bl[0] br[0] wl[5] vdd gnd cell_6t
Xbit_r6_c0 bl[0] br[0] wl[6] vdd gnd cell_6t
Xbit_r7_c0 bl[0] br[0] wl[7] vdd gnd cell_6t
Xbit_r8_c0 bl[0] br[0] wl[8] vdd gnd cell_6t
Xbit_r9_c0 bl[0] br[0] wl[9] vdd gnd cell_6t
Xbit_r10_c0 bl[0] br[0] wl[10] vdd gnd cell_6t
Xbit_r11_c0 bl[0] br[0] wl[11] vdd gnd cell_6t
Xbit_r12_c0 bl[0] br[0] wl[12] vdd gnd cell_6t
Xbit_r13_c0 bl[0] br[0] wl[13] vdd gnd cell_6t
Xbit_r14_c0 bl[0] br[0] wl[14] vdd gnd cell_6t
Xbit_r15_c0 bl[0] br[0] wl[15] vdd gnd cell_6t
Xbit_r16_c0 bl[0] br[0] wl[16] vdd gnd cell_6t
Xbit_r17_c0 bl[0] br[0] wl[17] vdd gnd cell_6t
Xbit_r18_c0 bl[0] br[0] wl[18] vdd gnd cell_6t
Xbit_r19_c0 bl[0] br[0] wl[19] vdd gnd cell_6t
Xbit_r20_c0 bl[0] br[0] wl[20] vdd gnd cell_6t
Xbit_r21_c0 bl[0] br[0] wl[21] vdd gnd cell_6t
Xbit_r22_c0 bl[0] br[0] wl[22] vdd gnd cell_6t
Xbit_r23_c0 bl[0] br[0] wl[23] vdd gnd cell_6t
Xbit_r24_c0 bl[0] br[0] wl[24] vdd gnd cell_6t
Xbit_r25_c0 bl[0] br[0] wl[25] vdd gnd cell_6t
Xbit_r26_c0 bl[0] br[0] wl[26] vdd gnd cell_6t
Xbit_r27_c0 bl[0] br[0] wl[27] vdd gnd cell_6t
Xbit_r28_c0 bl[0] br[0] wl[28] vdd gnd cell_6t
Xbit_r29_c0 bl[0] br[0] wl[29] vdd gnd cell_6t
Xbit_r30_c0 bl[0] br[0] wl[30] vdd gnd cell_6t
Xbit_r31_c0 bl[0] br[0] wl[31] vdd gnd cell_6t
Xbit_r32_c0 bl[0] br[0] wl[32] vdd gnd cell_6t
Xbit_r33_c0 bl[0] br[0] wl[33] vdd gnd cell_6t
Xbit_r34_c0 bl[0] br[0] wl[34] vdd gnd cell_6t
Xbit_r35_c0 bl[0] br[0] wl[35] vdd gnd cell_6t
Xbit_r36_c0 bl[0] br[0] wl[36] vdd gnd cell_6t
Xbit_r37_c0 bl[0] br[0] wl[37] vdd gnd cell_6t
Xbit_r38_c0 bl[0] br[0] wl[38] vdd gnd cell_6t
Xbit_r39_c0 bl[0] br[0] wl[39] vdd gnd cell_6t
Xbit_r40_c0 bl[0] br[0] wl[40] vdd gnd cell_6t
Xbit_r41_c0 bl[0] br[0] wl[41] vdd gnd cell_6t
Xbit_r42_c0 bl[0] br[0] wl[42] vdd gnd cell_6t
Xbit_r43_c0 bl[0] br[0] wl[43] vdd gnd cell_6t
Xbit_r44_c0 bl[0] br[0] wl[44] vdd gnd cell_6t
Xbit_r45_c0 bl[0] br[0] wl[45] vdd gnd cell_6t
Xbit_r46_c0 bl[0] br[0] wl[46] vdd gnd cell_6t
Xbit_r47_c0 bl[0] br[0] wl[47] vdd gnd cell_6t
Xbit_r48_c0 bl[0] br[0] wl[48] vdd gnd cell_6t
Xbit_r49_c0 bl[0] br[0] wl[49] vdd gnd cell_6t
Xbit_r50_c0 bl[0] br[0] wl[50] vdd gnd cell_6t
Xbit_r51_c0 bl[0] br[0] wl[51] vdd gnd cell_6t
Xbit_r52_c0 bl[0] br[0] wl[52] vdd gnd cell_6t
Xbit_r53_c0 bl[0] br[0] wl[53] vdd gnd cell_6t
Xbit_r54_c0 bl[0] br[0] wl[54] vdd gnd cell_6t
Xbit_r55_c0 bl[0] br[0] wl[55] vdd gnd cell_6t
Xbit_r56_c0 bl[0] br[0] wl[56] vdd gnd cell_6t
Xbit_r57_c0 bl[0] br[0] wl[57] vdd gnd cell_6t
Xbit_r58_c0 bl[0] br[0] wl[58] vdd gnd cell_6t
Xbit_r59_c0 bl[0] br[0] wl[59] vdd gnd cell_6t
Xbit_r60_c0 bl[0] br[0] wl[60] vdd gnd cell_6t
Xbit_r61_c0 bl[0] br[0] wl[61] vdd gnd cell_6t
Xbit_r62_c0 bl[0] br[0] wl[62] vdd gnd cell_6t
Xbit_r63_c0 bl[0] br[0] wl[63] vdd gnd cell_6t
Xbit_r64_c0 bl[0] br[0] wl[64] vdd gnd cell_6t
Xbit_r65_c0 bl[0] br[0] wl[65] vdd gnd cell_6t
Xbit_r66_c0 bl[0] br[0] wl[66] vdd gnd cell_6t
Xbit_r67_c0 bl[0] br[0] wl[67] vdd gnd cell_6t
Xbit_r68_c0 bl[0] br[0] wl[68] vdd gnd cell_6t
Xbit_r69_c0 bl[0] br[0] wl[69] vdd gnd cell_6t
Xbit_r70_c0 bl[0] br[0] wl[70] vdd gnd cell_6t
Xbit_r71_c0 bl[0] br[0] wl[71] vdd gnd cell_6t
Xbit_r72_c0 bl[0] br[0] wl[72] vdd gnd cell_6t
Xbit_r73_c0 bl[0] br[0] wl[73] vdd gnd cell_6t
Xbit_r74_c0 bl[0] br[0] wl[74] vdd gnd cell_6t
Xbit_r75_c0 bl[0] br[0] wl[75] vdd gnd cell_6t
Xbit_r76_c0 bl[0] br[0] wl[76] vdd gnd cell_6t
Xbit_r77_c0 bl[0] br[0] wl[77] vdd gnd cell_6t
Xbit_r78_c0 bl[0] br[0] wl[78] vdd gnd cell_6t
Xbit_r79_c0 bl[0] br[0] wl[79] vdd gnd cell_6t
Xbit_r80_c0 bl[0] br[0] wl[80] vdd gnd cell_6t
Xbit_r81_c0 bl[0] br[0] wl[81] vdd gnd cell_6t
Xbit_r82_c0 bl[0] br[0] wl[82] vdd gnd cell_6t
Xbit_r83_c0 bl[0] br[0] wl[83] vdd gnd cell_6t
Xbit_r84_c0 bl[0] br[0] wl[84] vdd gnd cell_6t
Xbit_r85_c0 bl[0] br[0] wl[85] vdd gnd cell_6t
Xbit_r86_c0 bl[0] br[0] wl[86] vdd gnd cell_6t
Xbit_r87_c0 bl[0] br[0] wl[87] vdd gnd cell_6t
Xbit_r88_c0 bl[0] br[0] wl[88] vdd gnd cell_6t
Xbit_r89_c0 bl[0] br[0] wl[89] vdd gnd cell_6t
Xbit_r90_c0 bl[0] br[0] wl[90] vdd gnd cell_6t
Xbit_r91_c0 bl[0] br[0] wl[91] vdd gnd cell_6t
Xbit_r92_c0 bl[0] br[0] wl[92] vdd gnd cell_6t
Xbit_r93_c0 bl[0] br[0] wl[93] vdd gnd cell_6t
Xbit_r94_c0 bl[0] br[0] wl[94] vdd gnd cell_6t
Xbit_r95_c0 bl[0] br[0] wl[95] vdd gnd cell_6t
Xbit_r96_c0 bl[0] br[0] wl[96] vdd gnd cell_6t
Xbit_r97_c0 bl[0] br[0] wl[97] vdd gnd cell_6t
Xbit_r98_c0 bl[0] br[0] wl[98] vdd gnd cell_6t
Xbit_r99_c0 bl[0] br[0] wl[99] vdd gnd cell_6t
Xbit_r100_c0 bl[0] br[0] wl[100] vdd gnd cell_6t
Xbit_r101_c0 bl[0] br[0] wl[101] vdd gnd cell_6t
Xbit_r102_c0 bl[0] br[0] wl[102] vdd gnd cell_6t
Xbit_r103_c0 bl[0] br[0] wl[103] vdd gnd cell_6t
Xbit_r104_c0 bl[0] br[0] wl[104] vdd gnd cell_6t
Xbit_r105_c0 bl[0] br[0] wl[105] vdd gnd cell_6t
Xbit_r106_c0 bl[0] br[0] wl[106] vdd gnd cell_6t
Xbit_r107_c0 bl[0] br[0] wl[107] vdd gnd cell_6t
Xbit_r108_c0 bl[0] br[0] wl[108] vdd gnd cell_6t
Xbit_r109_c0 bl[0] br[0] wl[109] vdd gnd cell_6t
Xbit_r110_c0 bl[0] br[0] wl[110] vdd gnd cell_6t
Xbit_r111_c0 bl[0] br[0] wl[111] vdd gnd cell_6t
Xbit_r112_c0 bl[0] br[0] wl[112] vdd gnd cell_6t
Xbit_r113_c0 bl[0] br[0] wl[113] vdd gnd cell_6t
Xbit_r114_c0 bl[0] br[0] wl[114] vdd gnd cell_6t
Xbit_r115_c0 bl[0] br[0] wl[115] vdd gnd cell_6t
Xbit_r116_c0 bl[0] br[0] wl[116] vdd gnd cell_6t
Xbit_r117_c0 bl[0] br[0] wl[117] vdd gnd cell_6t
Xbit_r118_c0 bl[0] br[0] wl[118] vdd gnd cell_6t
Xbit_r119_c0 bl[0] br[0] wl[119] vdd gnd cell_6t
Xbit_r120_c0 bl[0] br[0] wl[120] vdd gnd cell_6t
Xbit_r121_c0 bl[0] br[0] wl[121] vdd gnd cell_6t
Xbit_r122_c0 bl[0] br[0] wl[122] vdd gnd cell_6t
Xbit_r123_c0 bl[0] br[0] wl[123] vdd gnd cell_6t
Xbit_r124_c0 bl[0] br[0] wl[124] vdd gnd cell_6t
Xbit_r125_c0 bl[0] br[0] wl[125] vdd gnd cell_6t
Xbit_r126_c0 bl[0] br[0] wl[126] vdd gnd cell_6t
Xbit_r127_c0 bl[0] br[0] wl[127] vdd gnd cell_6t
Xbit_r128_c0 bl[0] br[0] wl[128] vdd gnd cell_6t
Xbit_r129_c0 bl[0] br[0] wl[129] vdd gnd cell_6t
Xbit_r130_c0 bl[0] br[0] wl[130] vdd gnd cell_6t
Xbit_r131_c0 bl[0] br[0] wl[131] vdd gnd cell_6t
Xbit_r132_c0 bl[0] br[0] wl[132] vdd gnd cell_6t
Xbit_r133_c0 bl[0] br[0] wl[133] vdd gnd cell_6t
Xbit_r134_c0 bl[0] br[0] wl[134] vdd gnd cell_6t
Xbit_r135_c0 bl[0] br[0] wl[135] vdd gnd cell_6t
Xbit_r136_c0 bl[0] br[0] wl[136] vdd gnd cell_6t
Xbit_r137_c0 bl[0] br[0] wl[137] vdd gnd cell_6t
Xbit_r138_c0 bl[0] br[0] wl[138] vdd gnd cell_6t
Xbit_r139_c0 bl[0] br[0] wl[139] vdd gnd cell_6t
Xbit_r140_c0 bl[0] br[0] wl[140] vdd gnd cell_6t
Xbit_r141_c0 bl[0] br[0] wl[141] vdd gnd cell_6t
Xbit_r142_c0 bl[0] br[0] wl[142] vdd gnd cell_6t
Xbit_r143_c0 bl[0] br[0] wl[143] vdd gnd cell_6t
Xbit_r144_c0 bl[0] br[0] wl[144] vdd gnd cell_6t
Xbit_r145_c0 bl[0] br[0] wl[145] vdd gnd cell_6t
Xbit_r146_c0 bl[0] br[0] wl[146] vdd gnd cell_6t
Xbit_r147_c0 bl[0] br[0] wl[147] vdd gnd cell_6t
Xbit_r148_c0 bl[0] br[0] wl[148] vdd gnd cell_6t
Xbit_r149_c0 bl[0] br[0] wl[149] vdd gnd cell_6t
Xbit_r150_c0 bl[0] br[0] wl[150] vdd gnd cell_6t
Xbit_r151_c0 bl[0] br[0] wl[151] vdd gnd cell_6t
Xbit_r152_c0 bl[0] br[0] wl[152] vdd gnd cell_6t
Xbit_r153_c0 bl[0] br[0] wl[153] vdd gnd cell_6t
Xbit_r154_c0 bl[0] br[0] wl[154] vdd gnd cell_6t
Xbit_r155_c0 bl[0] br[0] wl[155] vdd gnd cell_6t
Xbit_r156_c0 bl[0] br[0] wl[156] vdd gnd cell_6t
Xbit_r157_c0 bl[0] br[0] wl[157] vdd gnd cell_6t
Xbit_r158_c0 bl[0] br[0] wl[158] vdd gnd cell_6t
Xbit_r159_c0 bl[0] br[0] wl[159] vdd gnd cell_6t
Xbit_r160_c0 bl[0] br[0] wl[160] vdd gnd cell_6t
Xbit_r161_c0 bl[0] br[0] wl[161] vdd gnd cell_6t
Xbit_r162_c0 bl[0] br[0] wl[162] vdd gnd cell_6t
Xbit_r163_c0 bl[0] br[0] wl[163] vdd gnd cell_6t
Xbit_r164_c0 bl[0] br[0] wl[164] vdd gnd cell_6t
Xbit_r165_c0 bl[0] br[0] wl[165] vdd gnd cell_6t
Xbit_r166_c0 bl[0] br[0] wl[166] vdd gnd cell_6t
Xbit_r167_c0 bl[0] br[0] wl[167] vdd gnd cell_6t
Xbit_r168_c0 bl[0] br[0] wl[168] vdd gnd cell_6t
Xbit_r169_c0 bl[0] br[0] wl[169] vdd gnd cell_6t
Xbit_r170_c0 bl[0] br[0] wl[170] vdd gnd cell_6t
Xbit_r171_c0 bl[0] br[0] wl[171] vdd gnd cell_6t
Xbit_r172_c0 bl[0] br[0] wl[172] vdd gnd cell_6t
Xbit_r173_c0 bl[0] br[0] wl[173] vdd gnd cell_6t
Xbit_r174_c0 bl[0] br[0] wl[174] vdd gnd cell_6t
Xbit_r175_c0 bl[0] br[0] wl[175] vdd gnd cell_6t
Xbit_r176_c0 bl[0] br[0] wl[176] vdd gnd cell_6t
Xbit_r177_c0 bl[0] br[0] wl[177] vdd gnd cell_6t
Xbit_r178_c0 bl[0] br[0] wl[178] vdd gnd cell_6t
Xbit_r179_c0 bl[0] br[0] wl[179] vdd gnd cell_6t
Xbit_r180_c0 bl[0] br[0] wl[180] vdd gnd cell_6t
Xbit_r181_c0 bl[0] br[0] wl[181] vdd gnd cell_6t
Xbit_r182_c0 bl[0] br[0] wl[182] vdd gnd cell_6t
Xbit_r183_c0 bl[0] br[0] wl[183] vdd gnd cell_6t
Xbit_r184_c0 bl[0] br[0] wl[184] vdd gnd cell_6t
Xbit_r185_c0 bl[0] br[0] wl[185] vdd gnd cell_6t
Xbit_r186_c0 bl[0] br[0] wl[186] vdd gnd cell_6t
Xbit_r187_c0 bl[0] br[0] wl[187] vdd gnd cell_6t
Xbit_r188_c0 bl[0] br[0] wl[188] vdd gnd cell_6t
Xbit_r189_c0 bl[0] br[0] wl[189] vdd gnd cell_6t
Xbit_r190_c0 bl[0] br[0] wl[190] vdd gnd cell_6t
Xbit_r191_c0 bl[0] br[0] wl[191] vdd gnd cell_6t
Xbit_r192_c0 bl[0] br[0] wl[192] vdd gnd cell_6t
Xbit_r193_c0 bl[0] br[0] wl[193] vdd gnd cell_6t
Xbit_r194_c0 bl[0] br[0] wl[194] vdd gnd cell_6t
Xbit_r195_c0 bl[0] br[0] wl[195] vdd gnd cell_6t
Xbit_r196_c0 bl[0] br[0] wl[196] vdd gnd cell_6t
Xbit_r197_c0 bl[0] br[0] wl[197] vdd gnd cell_6t
Xbit_r198_c0 bl[0] br[0] wl[198] vdd gnd cell_6t
Xbit_r199_c0 bl[0] br[0] wl[199] vdd gnd cell_6t
Xbit_r200_c0 bl[0] br[0] wl[200] vdd gnd cell_6t
Xbit_r201_c0 bl[0] br[0] wl[201] vdd gnd cell_6t
Xbit_r202_c0 bl[0] br[0] wl[202] vdd gnd cell_6t
Xbit_r203_c0 bl[0] br[0] wl[203] vdd gnd cell_6t
Xbit_r204_c0 bl[0] br[0] wl[204] vdd gnd cell_6t
Xbit_r205_c0 bl[0] br[0] wl[205] vdd gnd cell_6t
Xbit_r206_c0 bl[0] br[0] wl[206] vdd gnd cell_6t
Xbit_r207_c0 bl[0] br[0] wl[207] vdd gnd cell_6t
Xbit_r208_c0 bl[0] br[0] wl[208] vdd gnd cell_6t
Xbit_r209_c0 bl[0] br[0] wl[209] vdd gnd cell_6t
Xbit_r210_c0 bl[0] br[0] wl[210] vdd gnd cell_6t
Xbit_r211_c0 bl[0] br[0] wl[211] vdd gnd cell_6t
Xbit_r212_c0 bl[0] br[0] wl[212] vdd gnd cell_6t
Xbit_r213_c0 bl[0] br[0] wl[213] vdd gnd cell_6t
Xbit_r214_c0 bl[0] br[0] wl[214] vdd gnd cell_6t
Xbit_r215_c0 bl[0] br[0] wl[215] vdd gnd cell_6t
Xbit_r216_c0 bl[0] br[0] wl[216] vdd gnd cell_6t
Xbit_r217_c0 bl[0] br[0] wl[217] vdd gnd cell_6t
Xbit_r218_c0 bl[0] br[0] wl[218] vdd gnd cell_6t
Xbit_r219_c0 bl[0] br[0] wl[219] vdd gnd cell_6t
Xbit_r220_c0 bl[0] br[0] wl[220] vdd gnd cell_6t
Xbit_r221_c0 bl[0] br[0] wl[221] vdd gnd cell_6t
Xbit_r222_c0 bl[0] br[0] wl[222] vdd gnd cell_6t
Xbit_r223_c0 bl[0] br[0] wl[223] vdd gnd cell_6t
Xbit_r224_c0 bl[0] br[0] wl[224] vdd gnd cell_6t
Xbit_r225_c0 bl[0] br[0] wl[225] vdd gnd cell_6t
Xbit_r226_c0 bl[0] br[0] wl[226] vdd gnd cell_6t
Xbit_r227_c0 bl[0] br[0] wl[227] vdd gnd cell_6t
Xbit_r228_c0 bl[0] br[0] wl[228] vdd gnd cell_6t
Xbit_r229_c0 bl[0] br[0] wl[229] vdd gnd cell_6t
Xbit_r230_c0 bl[0] br[0] wl[230] vdd gnd cell_6t
Xbit_r231_c0 bl[0] br[0] wl[231] vdd gnd cell_6t
Xbit_r232_c0 bl[0] br[0] wl[232] vdd gnd cell_6t
Xbit_r233_c0 bl[0] br[0] wl[233] vdd gnd cell_6t
Xbit_r234_c0 bl[0] br[0] wl[234] vdd gnd cell_6t
Xbit_r235_c0 bl[0] br[0] wl[235] vdd gnd cell_6t
Xbit_r236_c0 bl[0] br[0] wl[236] vdd gnd cell_6t
Xbit_r237_c0 bl[0] br[0] wl[237] vdd gnd cell_6t
Xbit_r238_c0 bl[0] br[0] wl[238] vdd gnd cell_6t
Xbit_r239_c0 bl[0] br[0] wl[239] vdd gnd cell_6t
Xbit_r240_c0 bl[0] br[0] wl[240] vdd gnd cell_6t
Xbit_r241_c0 bl[0] br[0] wl[241] vdd gnd cell_6t
Xbit_r242_c0 bl[0] br[0] wl[242] vdd gnd cell_6t
Xbit_r243_c0 bl[0] br[0] wl[243] vdd gnd cell_6t
Xbit_r244_c0 bl[0] br[0] wl[244] vdd gnd cell_6t
Xbit_r245_c0 bl[0] br[0] wl[245] vdd gnd cell_6t
Xbit_r246_c0 bl[0] br[0] wl[246] vdd gnd cell_6t
Xbit_r247_c0 bl[0] br[0] wl[247] vdd gnd cell_6t
Xbit_r248_c0 bl[0] br[0] wl[248] vdd gnd cell_6t
Xbit_r249_c0 bl[0] br[0] wl[249] vdd gnd cell_6t
Xbit_r250_c0 bl[0] br[0] wl[250] vdd gnd cell_6t
Xbit_r251_c0 bl[0] br[0] wl[251] vdd gnd cell_6t
Xbit_r252_c0 bl[0] br[0] wl[252] vdd gnd cell_6t
Xbit_r253_c0 bl[0] br[0] wl[253] vdd gnd cell_6t
Xbit_r254_c0 bl[0] br[0] wl[254] vdd gnd cell_6t
Xbit_r255_c0 bl[0] br[0] wl[255] vdd gnd cell_6t
Xbit_r256_c0 bl[0] br[0] wl[256] vdd gnd cell_6t
Xbit_r257_c0 bl[0] br[0] wl[257] vdd gnd cell_6t
Xbit_r258_c0 bl[0] br[0] wl[258] vdd gnd cell_6t
Xbit_r259_c0 bl[0] br[0] wl[259] vdd gnd cell_6t
Xbit_r260_c0 bl[0] br[0] wl[260] vdd gnd cell_6t
Xbit_r261_c0 bl[0] br[0] wl[261] vdd gnd cell_6t
Xbit_r262_c0 bl[0] br[0] wl[262] vdd gnd cell_6t
Xbit_r263_c0 bl[0] br[0] wl[263] vdd gnd cell_6t
Xbit_r264_c0 bl[0] br[0] wl[264] vdd gnd cell_6t
Xbit_r265_c0 bl[0] br[0] wl[265] vdd gnd cell_6t
Xbit_r266_c0 bl[0] br[0] wl[266] vdd gnd cell_6t
Xbit_r267_c0 bl[0] br[0] wl[267] vdd gnd cell_6t
Xbit_r268_c0 bl[0] br[0] wl[268] vdd gnd cell_6t
Xbit_r269_c0 bl[0] br[0] wl[269] vdd gnd cell_6t
Xbit_r270_c0 bl[0] br[0] wl[270] vdd gnd cell_6t
Xbit_r271_c0 bl[0] br[0] wl[271] vdd gnd cell_6t
Xbit_r272_c0 bl[0] br[0] wl[272] vdd gnd cell_6t
Xbit_r273_c0 bl[0] br[0] wl[273] vdd gnd cell_6t
Xbit_r274_c0 bl[0] br[0] wl[274] vdd gnd cell_6t
Xbit_r275_c0 bl[0] br[0] wl[275] vdd gnd cell_6t
Xbit_r276_c0 bl[0] br[0] wl[276] vdd gnd cell_6t
Xbit_r277_c0 bl[0] br[0] wl[277] vdd gnd cell_6t
Xbit_r278_c0 bl[0] br[0] wl[278] vdd gnd cell_6t
Xbit_r279_c0 bl[0] br[0] wl[279] vdd gnd cell_6t
Xbit_r280_c0 bl[0] br[0] wl[280] vdd gnd cell_6t
Xbit_r281_c0 bl[0] br[0] wl[281] vdd gnd cell_6t
Xbit_r282_c0 bl[0] br[0] wl[282] vdd gnd cell_6t
Xbit_r283_c0 bl[0] br[0] wl[283] vdd gnd cell_6t
Xbit_r284_c0 bl[0] br[0] wl[284] vdd gnd cell_6t
Xbit_r285_c0 bl[0] br[0] wl[285] vdd gnd cell_6t
Xbit_r286_c0 bl[0] br[0] wl[286] vdd gnd cell_6t
Xbit_r287_c0 bl[0] br[0] wl[287] vdd gnd cell_6t
Xbit_r288_c0 bl[0] br[0] wl[288] vdd gnd cell_6t
Xbit_r289_c0 bl[0] br[0] wl[289] vdd gnd cell_6t
Xbit_r290_c0 bl[0] br[0] wl[290] vdd gnd cell_6t
Xbit_r291_c0 bl[0] br[0] wl[291] vdd gnd cell_6t
Xbit_r292_c0 bl[0] br[0] wl[292] vdd gnd cell_6t
Xbit_r293_c0 bl[0] br[0] wl[293] vdd gnd cell_6t
Xbit_r294_c0 bl[0] br[0] wl[294] vdd gnd cell_6t
Xbit_r295_c0 bl[0] br[0] wl[295] vdd gnd cell_6t
Xbit_r296_c0 bl[0] br[0] wl[296] vdd gnd cell_6t
Xbit_r297_c0 bl[0] br[0] wl[297] vdd gnd cell_6t
Xbit_r298_c0 bl[0] br[0] wl[298] vdd gnd cell_6t
Xbit_r299_c0 bl[0] br[0] wl[299] vdd gnd cell_6t
Xbit_r300_c0 bl[0] br[0] wl[300] vdd gnd cell_6t
Xbit_r301_c0 bl[0] br[0] wl[301] vdd gnd cell_6t
Xbit_r302_c0 bl[0] br[0] wl[302] vdd gnd cell_6t
Xbit_r303_c0 bl[0] br[0] wl[303] vdd gnd cell_6t
Xbit_r304_c0 bl[0] br[0] wl[304] vdd gnd cell_6t
Xbit_r305_c0 bl[0] br[0] wl[305] vdd gnd cell_6t
Xbit_r306_c0 bl[0] br[0] wl[306] vdd gnd cell_6t
Xbit_r307_c0 bl[0] br[0] wl[307] vdd gnd cell_6t
Xbit_r308_c0 bl[0] br[0] wl[308] vdd gnd cell_6t
Xbit_r309_c0 bl[0] br[0] wl[309] vdd gnd cell_6t
Xbit_r310_c0 bl[0] br[0] wl[310] vdd gnd cell_6t
Xbit_r311_c0 bl[0] br[0] wl[311] vdd gnd cell_6t
Xbit_r312_c0 bl[0] br[0] wl[312] vdd gnd cell_6t
Xbit_r313_c0 bl[0] br[0] wl[313] vdd gnd cell_6t
Xbit_r314_c0 bl[0] br[0] wl[314] vdd gnd cell_6t
Xbit_r315_c0 bl[0] br[0] wl[315] vdd gnd cell_6t
Xbit_r316_c0 bl[0] br[0] wl[316] vdd gnd cell_6t
Xbit_r317_c0 bl[0] br[0] wl[317] vdd gnd cell_6t
Xbit_r318_c0 bl[0] br[0] wl[318] vdd gnd cell_6t
Xbit_r319_c0 bl[0] br[0] wl[319] vdd gnd cell_6t
Xbit_r320_c0 bl[0] br[0] wl[320] vdd gnd cell_6t
Xbit_r321_c0 bl[0] br[0] wl[321] vdd gnd cell_6t
Xbit_r322_c0 bl[0] br[0] wl[322] vdd gnd cell_6t
Xbit_r323_c0 bl[0] br[0] wl[323] vdd gnd cell_6t
Xbit_r324_c0 bl[0] br[0] wl[324] vdd gnd cell_6t
Xbit_r325_c0 bl[0] br[0] wl[325] vdd gnd cell_6t
Xbit_r326_c0 bl[0] br[0] wl[326] vdd gnd cell_6t
Xbit_r327_c0 bl[0] br[0] wl[327] vdd gnd cell_6t
Xbit_r328_c0 bl[0] br[0] wl[328] vdd gnd cell_6t
Xbit_r329_c0 bl[0] br[0] wl[329] vdd gnd cell_6t
Xbit_r330_c0 bl[0] br[0] wl[330] vdd gnd cell_6t
Xbit_r331_c0 bl[0] br[0] wl[331] vdd gnd cell_6t
Xbit_r332_c0 bl[0] br[0] wl[332] vdd gnd cell_6t
Xbit_r333_c0 bl[0] br[0] wl[333] vdd gnd cell_6t
Xbit_r334_c0 bl[0] br[0] wl[334] vdd gnd cell_6t
Xbit_r335_c0 bl[0] br[0] wl[335] vdd gnd cell_6t
Xbit_r336_c0 bl[0] br[0] wl[336] vdd gnd cell_6t
Xbit_r337_c0 bl[0] br[0] wl[337] vdd gnd cell_6t
Xbit_r338_c0 bl[0] br[0] wl[338] vdd gnd cell_6t
Xbit_r339_c0 bl[0] br[0] wl[339] vdd gnd cell_6t
Xbit_r340_c0 bl[0] br[0] wl[340] vdd gnd cell_6t
Xbit_r341_c0 bl[0] br[0] wl[341] vdd gnd cell_6t
Xbit_r342_c0 bl[0] br[0] wl[342] vdd gnd cell_6t
Xbit_r343_c0 bl[0] br[0] wl[343] vdd gnd cell_6t
Xbit_r344_c0 bl[0] br[0] wl[344] vdd gnd cell_6t
Xbit_r345_c0 bl[0] br[0] wl[345] vdd gnd cell_6t
Xbit_r346_c0 bl[0] br[0] wl[346] vdd gnd cell_6t
Xbit_r347_c0 bl[0] br[0] wl[347] vdd gnd cell_6t
Xbit_r348_c0 bl[0] br[0] wl[348] vdd gnd cell_6t
Xbit_r349_c0 bl[0] br[0] wl[349] vdd gnd cell_6t
Xbit_r350_c0 bl[0] br[0] wl[350] vdd gnd cell_6t
Xbit_r351_c0 bl[0] br[0] wl[351] vdd gnd cell_6t
Xbit_r352_c0 bl[0] br[0] wl[352] vdd gnd cell_6t
Xbit_r353_c0 bl[0] br[0] wl[353] vdd gnd cell_6t
Xbit_r354_c0 bl[0] br[0] wl[354] vdd gnd cell_6t
Xbit_r355_c0 bl[0] br[0] wl[355] vdd gnd cell_6t
Xbit_r356_c0 bl[0] br[0] wl[356] vdd gnd cell_6t
Xbit_r357_c0 bl[0] br[0] wl[357] vdd gnd cell_6t
Xbit_r358_c0 bl[0] br[0] wl[358] vdd gnd cell_6t
Xbit_r359_c0 bl[0] br[0] wl[359] vdd gnd cell_6t
Xbit_r360_c0 bl[0] br[0] wl[360] vdd gnd cell_6t
Xbit_r361_c0 bl[0] br[0] wl[361] vdd gnd cell_6t
Xbit_r362_c0 bl[0] br[0] wl[362] vdd gnd cell_6t
Xbit_r363_c0 bl[0] br[0] wl[363] vdd gnd cell_6t
Xbit_r364_c0 bl[0] br[0] wl[364] vdd gnd cell_6t
Xbit_r365_c0 bl[0] br[0] wl[365] vdd gnd cell_6t
Xbit_r366_c0 bl[0] br[0] wl[366] vdd gnd cell_6t
Xbit_r367_c0 bl[0] br[0] wl[367] vdd gnd cell_6t
Xbit_r368_c0 bl[0] br[0] wl[368] vdd gnd cell_6t
Xbit_r369_c0 bl[0] br[0] wl[369] vdd gnd cell_6t
Xbit_r370_c0 bl[0] br[0] wl[370] vdd gnd cell_6t
Xbit_r371_c0 bl[0] br[0] wl[371] vdd gnd cell_6t
Xbit_r372_c0 bl[0] br[0] wl[372] vdd gnd cell_6t
Xbit_r373_c0 bl[0] br[0] wl[373] vdd gnd cell_6t
Xbit_r374_c0 bl[0] br[0] wl[374] vdd gnd cell_6t
Xbit_r375_c0 bl[0] br[0] wl[375] vdd gnd cell_6t
Xbit_r376_c0 bl[0] br[0] wl[376] vdd gnd cell_6t
Xbit_r377_c0 bl[0] br[0] wl[377] vdd gnd cell_6t
Xbit_r378_c0 bl[0] br[0] wl[378] vdd gnd cell_6t
Xbit_r379_c0 bl[0] br[0] wl[379] vdd gnd cell_6t
Xbit_r380_c0 bl[0] br[0] wl[380] vdd gnd cell_6t
Xbit_r381_c0 bl[0] br[0] wl[381] vdd gnd cell_6t
Xbit_r382_c0 bl[0] br[0] wl[382] vdd gnd cell_6t
Xbit_r383_c0 bl[0] br[0] wl[383] vdd gnd cell_6t
Xbit_r384_c0 bl[0] br[0] wl[384] vdd gnd cell_6t
Xbit_r385_c0 bl[0] br[0] wl[385] vdd gnd cell_6t
Xbit_r386_c0 bl[0] br[0] wl[386] vdd gnd cell_6t
Xbit_r387_c0 bl[0] br[0] wl[387] vdd gnd cell_6t
Xbit_r388_c0 bl[0] br[0] wl[388] vdd gnd cell_6t
Xbit_r389_c0 bl[0] br[0] wl[389] vdd gnd cell_6t
Xbit_r390_c0 bl[0] br[0] wl[390] vdd gnd cell_6t
Xbit_r391_c0 bl[0] br[0] wl[391] vdd gnd cell_6t
Xbit_r392_c0 bl[0] br[0] wl[392] vdd gnd cell_6t
Xbit_r393_c0 bl[0] br[0] wl[393] vdd gnd cell_6t
Xbit_r394_c0 bl[0] br[0] wl[394] vdd gnd cell_6t
Xbit_r395_c0 bl[0] br[0] wl[395] vdd gnd cell_6t
Xbit_r396_c0 bl[0] br[0] wl[396] vdd gnd cell_6t
Xbit_r397_c0 bl[0] br[0] wl[397] vdd gnd cell_6t
Xbit_r398_c0 bl[0] br[0] wl[398] vdd gnd cell_6t
Xbit_r399_c0 bl[0] br[0] wl[399] vdd gnd cell_6t
Xbit_r400_c0 bl[0] br[0] wl[400] vdd gnd cell_6t
Xbit_r401_c0 bl[0] br[0] wl[401] vdd gnd cell_6t
Xbit_r402_c0 bl[0] br[0] wl[402] vdd gnd cell_6t
Xbit_r403_c0 bl[0] br[0] wl[403] vdd gnd cell_6t
Xbit_r404_c0 bl[0] br[0] wl[404] vdd gnd cell_6t
Xbit_r405_c0 bl[0] br[0] wl[405] vdd gnd cell_6t
Xbit_r406_c0 bl[0] br[0] wl[406] vdd gnd cell_6t
Xbit_r407_c0 bl[0] br[0] wl[407] vdd gnd cell_6t
Xbit_r408_c0 bl[0] br[0] wl[408] vdd gnd cell_6t
Xbit_r409_c0 bl[0] br[0] wl[409] vdd gnd cell_6t
Xbit_r410_c0 bl[0] br[0] wl[410] vdd gnd cell_6t
Xbit_r411_c0 bl[0] br[0] wl[411] vdd gnd cell_6t
Xbit_r412_c0 bl[0] br[0] wl[412] vdd gnd cell_6t
Xbit_r413_c0 bl[0] br[0] wl[413] vdd gnd cell_6t
Xbit_r414_c0 bl[0] br[0] wl[414] vdd gnd cell_6t
Xbit_r415_c0 bl[0] br[0] wl[415] vdd gnd cell_6t
Xbit_r416_c0 bl[0] br[0] wl[416] vdd gnd cell_6t
Xbit_r417_c0 bl[0] br[0] wl[417] vdd gnd cell_6t
Xbit_r418_c0 bl[0] br[0] wl[418] vdd gnd cell_6t
Xbit_r419_c0 bl[0] br[0] wl[419] vdd gnd cell_6t
Xbit_r420_c0 bl[0] br[0] wl[420] vdd gnd cell_6t
Xbit_r421_c0 bl[0] br[0] wl[421] vdd gnd cell_6t
Xbit_r422_c0 bl[0] br[0] wl[422] vdd gnd cell_6t
Xbit_r423_c0 bl[0] br[0] wl[423] vdd gnd cell_6t
Xbit_r424_c0 bl[0] br[0] wl[424] vdd gnd cell_6t
Xbit_r425_c0 bl[0] br[0] wl[425] vdd gnd cell_6t
Xbit_r426_c0 bl[0] br[0] wl[426] vdd gnd cell_6t
Xbit_r427_c0 bl[0] br[0] wl[427] vdd gnd cell_6t
Xbit_r428_c0 bl[0] br[0] wl[428] vdd gnd cell_6t
Xbit_r429_c0 bl[0] br[0] wl[429] vdd gnd cell_6t
Xbit_r430_c0 bl[0] br[0] wl[430] vdd gnd cell_6t
Xbit_r431_c0 bl[0] br[0] wl[431] vdd gnd cell_6t
Xbit_r432_c0 bl[0] br[0] wl[432] vdd gnd cell_6t
Xbit_r433_c0 bl[0] br[0] wl[433] vdd gnd cell_6t
Xbit_r434_c0 bl[0] br[0] wl[434] vdd gnd cell_6t
Xbit_r435_c0 bl[0] br[0] wl[435] vdd gnd cell_6t
Xbit_r436_c0 bl[0] br[0] wl[436] vdd gnd cell_6t
Xbit_r437_c0 bl[0] br[0] wl[437] vdd gnd cell_6t
Xbit_r438_c0 bl[0] br[0] wl[438] vdd gnd cell_6t
Xbit_r439_c0 bl[0] br[0] wl[439] vdd gnd cell_6t
Xbit_r440_c0 bl[0] br[0] wl[440] vdd gnd cell_6t
Xbit_r441_c0 bl[0] br[0] wl[441] vdd gnd cell_6t
Xbit_r442_c0 bl[0] br[0] wl[442] vdd gnd cell_6t
Xbit_r443_c0 bl[0] br[0] wl[443] vdd gnd cell_6t
Xbit_r444_c0 bl[0] br[0] wl[444] vdd gnd cell_6t
Xbit_r445_c0 bl[0] br[0] wl[445] vdd gnd cell_6t
Xbit_r446_c0 bl[0] br[0] wl[446] vdd gnd cell_6t
Xbit_r447_c0 bl[0] br[0] wl[447] vdd gnd cell_6t
Xbit_r448_c0 bl[0] br[0] wl[448] vdd gnd cell_6t
Xbit_r449_c0 bl[0] br[0] wl[449] vdd gnd cell_6t
Xbit_r450_c0 bl[0] br[0] wl[450] vdd gnd cell_6t
Xbit_r451_c0 bl[0] br[0] wl[451] vdd gnd cell_6t
Xbit_r452_c0 bl[0] br[0] wl[452] vdd gnd cell_6t
Xbit_r453_c0 bl[0] br[0] wl[453] vdd gnd cell_6t
Xbit_r454_c0 bl[0] br[0] wl[454] vdd gnd cell_6t
Xbit_r455_c0 bl[0] br[0] wl[455] vdd gnd cell_6t
Xbit_r456_c0 bl[0] br[0] wl[456] vdd gnd cell_6t
Xbit_r457_c0 bl[0] br[0] wl[457] vdd gnd cell_6t
Xbit_r458_c0 bl[0] br[0] wl[458] vdd gnd cell_6t
Xbit_r459_c0 bl[0] br[0] wl[459] vdd gnd cell_6t
Xbit_r460_c0 bl[0] br[0] wl[460] vdd gnd cell_6t
Xbit_r461_c0 bl[0] br[0] wl[461] vdd gnd cell_6t
Xbit_r462_c0 bl[0] br[0] wl[462] vdd gnd cell_6t
Xbit_r463_c0 bl[0] br[0] wl[463] vdd gnd cell_6t
Xbit_r464_c0 bl[0] br[0] wl[464] vdd gnd cell_6t
Xbit_r465_c0 bl[0] br[0] wl[465] vdd gnd cell_6t
Xbit_r466_c0 bl[0] br[0] wl[466] vdd gnd cell_6t
Xbit_r467_c0 bl[0] br[0] wl[467] vdd gnd cell_6t
Xbit_r468_c0 bl[0] br[0] wl[468] vdd gnd cell_6t
Xbit_r469_c0 bl[0] br[0] wl[469] vdd gnd cell_6t
Xbit_r470_c0 bl[0] br[0] wl[470] vdd gnd cell_6t
Xbit_r471_c0 bl[0] br[0] wl[471] vdd gnd cell_6t
Xbit_r472_c0 bl[0] br[0] wl[472] vdd gnd cell_6t
Xbit_r473_c0 bl[0] br[0] wl[473] vdd gnd cell_6t
Xbit_r474_c0 bl[0] br[0] wl[474] vdd gnd cell_6t
Xbit_r475_c0 bl[0] br[0] wl[475] vdd gnd cell_6t
Xbit_r476_c0 bl[0] br[0] wl[476] vdd gnd cell_6t
Xbit_r477_c0 bl[0] br[0] wl[477] vdd gnd cell_6t
Xbit_r478_c0 bl[0] br[0] wl[478] vdd gnd cell_6t
Xbit_r479_c0 bl[0] br[0] wl[479] vdd gnd cell_6t
Xbit_r480_c0 bl[0] br[0] wl[480] vdd gnd cell_6t
Xbit_r481_c0 bl[0] br[0] wl[481] vdd gnd cell_6t
Xbit_r482_c0 bl[0] br[0] wl[482] vdd gnd cell_6t
Xbit_r483_c0 bl[0] br[0] wl[483] vdd gnd cell_6t
Xbit_r484_c0 bl[0] br[0] wl[484] vdd gnd cell_6t
Xbit_r485_c0 bl[0] br[0] wl[485] vdd gnd cell_6t
Xbit_r486_c0 bl[0] br[0] wl[486] vdd gnd cell_6t
Xbit_r487_c0 bl[0] br[0] wl[487] vdd gnd cell_6t
Xbit_r488_c0 bl[0] br[0] wl[488] vdd gnd cell_6t
Xbit_r489_c0 bl[0] br[0] wl[489] vdd gnd cell_6t
Xbit_r490_c0 bl[0] br[0] wl[490] vdd gnd cell_6t
Xbit_r491_c0 bl[0] br[0] wl[491] vdd gnd cell_6t
Xbit_r492_c0 bl[0] br[0] wl[492] vdd gnd cell_6t
Xbit_r493_c0 bl[0] br[0] wl[493] vdd gnd cell_6t
Xbit_r494_c0 bl[0] br[0] wl[494] vdd gnd cell_6t
Xbit_r495_c0 bl[0] br[0] wl[495] vdd gnd cell_6t
Xbit_r496_c0 bl[0] br[0] wl[496] vdd gnd cell_6t
Xbit_r497_c0 bl[0] br[0] wl[497] vdd gnd cell_6t
Xbit_r498_c0 bl[0] br[0] wl[498] vdd gnd cell_6t
Xbit_r499_c0 bl[0] br[0] wl[499] vdd gnd cell_6t
Xbit_r500_c0 bl[0] br[0] wl[500] vdd gnd cell_6t
Xbit_r501_c0 bl[0] br[0] wl[501] vdd gnd cell_6t
Xbit_r502_c0 bl[0] br[0] wl[502] vdd gnd cell_6t
Xbit_r503_c0 bl[0] br[0] wl[503] vdd gnd cell_6t
Xbit_r504_c0 bl[0] br[0] wl[504] vdd gnd cell_6t
Xbit_r505_c0 bl[0] br[0] wl[505] vdd gnd cell_6t
Xbit_r506_c0 bl[0] br[0] wl[506] vdd gnd cell_6t
Xbit_r507_c0 bl[0] br[0] wl[507] vdd gnd cell_6t
Xbit_r508_c0 bl[0] br[0] wl[508] vdd gnd cell_6t
Xbit_r509_c0 bl[0] br[0] wl[509] vdd gnd cell_6t
Xbit_r510_c0 bl[0] br[0] wl[510] vdd gnd cell_6t
Xbit_r511_c0 bl[0] br[0] wl[511] vdd gnd cell_6t
Xbit_r0_c1 bl[1] br[1] wl[0] vdd gnd cell_6t
Xbit_r1_c1 bl[1] br[1] wl[1] vdd gnd cell_6t
Xbit_r2_c1 bl[1] br[1] wl[2] vdd gnd cell_6t
Xbit_r3_c1 bl[1] br[1] wl[3] vdd gnd cell_6t
Xbit_r4_c1 bl[1] br[1] wl[4] vdd gnd cell_6t
Xbit_r5_c1 bl[1] br[1] wl[5] vdd gnd cell_6t
Xbit_r6_c1 bl[1] br[1] wl[6] vdd gnd cell_6t
Xbit_r7_c1 bl[1] br[1] wl[7] vdd gnd cell_6t
Xbit_r8_c1 bl[1] br[1] wl[8] vdd gnd cell_6t
Xbit_r9_c1 bl[1] br[1] wl[9] vdd gnd cell_6t
Xbit_r10_c1 bl[1] br[1] wl[10] vdd gnd cell_6t
Xbit_r11_c1 bl[1] br[1] wl[11] vdd gnd cell_6t
Xbit_r12_c1 bl[1] br[1] wl[12] vdd gnd cell_6t
Xbit_r13_c1 bl[1] br[1] wl[13] vdd gnd cell_6t
Xbit_r14_c1 bl[1] br[1] wl[14] vdd gnd cell_6t
Xbit_r15_c1 bl[1] br[1] wl[15] vdd gnd cell_6t
Xbit_r16_c1 bl[1] br[1] wl[16] vdd gnd cell_6t
Xbit_r17_c1 bl[1] br[1] wl[17] vdd gnd cell_6t
Xbit_r18_c1 bl[1] br[1] wl[18] vdd gnd cell_6t
Xbit_r19_c1 bl[1] br[1] wl[19] vdd gnd cell_6t
Xbit_r20_c1 bl[1] br[1] wl[20] vdd gnd cell_6t
Xbit_r21_c1 bl[1] br[1] wl[21] vdd gnd cell_6t
Xbit_r22_c1 bl[1] br[1] wl[22] vdd gnd cell_6t
Xbit_r23_c1 bl[1] br[1] wl[23] vdd gnd cell_6t
Xbit_r24_c1 bl[1] br[1] wl[24] vdd gnd cell_6t
Xbit_r25_c1 bl[1] br[1] wl[25] vdd gnd cell_6t
Xbit_r26_c1 bl[1] br[1] wl[26] vdd gnd cell_6t
Xbit_r27_c1 bl[1] br[1] wl[27] vdd gnd cell_6t
Xbit_r28_c1 bl[1] br[1] wl[28] vdd gnd cell_6t
Xbit_r29_c1 bl[1] br[1] wl[29] vdd gnd cell_6t
Xbit_r30_c1 bl[1] br[1] wl[30] vdd gnd cell_6t
Xbit_r31_c1 bl[1] br[1] wl[31] vdd gnd cell_6t
Xbit_r32_c1 bl[1] br[1] wl[32] vdd gnd cell_6t
Xbit_r33_c1 bl[1] br[1] wl[33] vdd gnd cell_6t
Xbit_r34_c1 bl[1] br[1] wl[34] vdd gnd cell_6t
Xbit_r35_c1 bl[1] br[1] wl[35] vdd gnd cell_6t
Xbit_r36_c1 bl[1] br[1] wl[36] vdd gnd cell_6t
Xbit_r37_c1 bl[1] br[1] wl[37] vdd gnd cell_6t
Xbit_r38_c1 bl[1] br[1] wl[38] vdd gnd cell_6t
Xbit_r39_c1 bl[1] br[1] wl[39] vdd gnd cell_6t
Xbit_r40_c1 bl[1] br[1] wl[40] vdd gnd cell_6t
Xbit_r41_c1 bl[1] br[1] wl[41] vdd gnd cell_6t
Xbit_r42_c1 bl[1] br[1] wl[42] vdd gnd cell_6t
Xbit_r43_c1 bl[1] br[1] wl[43] vdd gnd cell_6t
Xbit_r44_c1 bl[1] br[1] wl[44] vdd gnd cell_6t
Xbit_r45_c1 bl[1] br[1] wl[45] vdd gnd cell_6t
Xbit_r46_c1 bl[1] br[1] wl[46] vdd gnd cell_6t
Xbit_r47_c1 bl[1] br[1] wl[47] vdd gnd cell_6t
Xbit_r48_c1 bl[1] br[1] wl[48] vdd gnd cell_6t
Xbit_r49_c1 bl[1] br[1] wl[49] vdd gnd cell_6t
Xbit_r50_c1 bl[1] br[1] wl[50] vdd gnd cell_6t
Xbit_r51_c1 bl[1] br[1] wl[51] vdd gnd cell_6t
Xbit_r52_c1 bl[1] br[1] wl[52] vdd gnd cell_6t
Xbit_r53_c1 bl[1] br[1] wl[53] vdd gnd cell_6t
Xbit_r54_c1 bl[1] br[1] wl[54] vdd gnd cell_6t
Xbit_r55_c1 bl[1] br[1] wl[55] vdd gnd cell_6t
Xbit_r56_c1 bl[1] br[1] wl[56] vdd gnd cell_6t
Xbit_r57_c1 bl[1] br[1] wl[57] vdd gnd cell_6t
Xbit_r58_c1 bl[1] br[1] wl[58] vdd gnd cell_6t
Xbit_r59_c1 bl[1] br[1] wl[59] vdd gnd cell_6t
Xbit_r60_c1 bl[1] br[1] wl[60] vdd gnd cell_6t
Xbit_r61_c1 bl[1] br[1] wl[61] vdd gnd cell_6t
Xbit_r62_c1 bl[1] br[1] wl[62] vdd gnd cell_6t
Xbit_r63_c1 bl[1] br[1] wl[63] vdd gnd cell_6t
Xbit_r64_c1 bl[1] br[1] wl[64] vdd gnd cell_6t
Xbit_r65_c1 bl[1] br[1] wl[65] vdd gnd cell_6t
Xbit_r66_c1 bl[1] br[1] wl[66] vdd gnd cell_6t
Xbit_r67_c1 bl[1] br[1] wl[67] vdd gnd cell_6t
Xbit_r68_c1 bl[1] br[1] wl[68] vdd gnd cell_6t
Xbit_r69_c1 bl[1] br[1] wl[69] vdd gnd cell_6t
Xbit_r70_c1 bl[1] br[1] wl[70] vdd gnd cell_6t
Xbit_r71_c1 bl[1] br[1] wl[71] vdd gnd cell_6t
Xbit_r72_c1 bl[1] br[1] wl[72] vdd gnd cell_6t
Xbit_r73_c1 bl[1] br[1] wl[73] vdd gnd cell_6t
Xbit_r74_c1 bl[1] br[1] wl[74] vdd gnd cell_6t
Xbit_r75_c1 bl[1] br[1] wl[75] vdd gnd cell_6t
Xbit_r76_c1 bl[1] br[1] wl[76] vdd gnd cell_6t
Xbit_r77_c1 bl[1] br[1] wl[77] vdd gnd cell_6t
Xbit_r78_c1 bl[1] br[1] wl[78] vdd gnd cell_6t
Xbit_r79_c1 bl[1] br[1] wl[79] vdd gnd cell_6t
Xbit_r80_c1 bl[1] br[1] wl[80] vdd gnd cell_6t
Xbit_r81_c1 bl[1] br[1] wl[81] vdd gnd cell_6t
Xbit_r82_c1 bl[1] br[1] wl[82] vdd gnd cell_6t
Xbit_r83_c1 bl[1] br[1] wl[83] vdd gnd cell_6t
Xbit_r84_c1 bl[1] br[1] wl[84] vdd gnd cell_6t
Xbit_r85_c1 bl[1] br[1] wl[85] vdd gnd cell_6t
Xbit_r86_c1 bl[1] br[1] wl[86] vdd gnd cell_6t
Xbit_r87_c1 bl[1] br[1] wl[87] vdd gnd cell_6t
Xbit_r88_c1 bl[1] br[1] wl[88] vdd gnd cell_6t
Xbit_r89_c1 bl[1] br[1] wl[89] vdd gnd cell_6t
Xbit_r90_c1 bl[1] br[1] wl[90] vdd gnd cell_6t
Xbit_r91_c1 bl[1] br[1] wl[91] vdd gnd cell_6t
Xbit_r92_c1 bl[1] br[1] wl[92] vdd gnd cell_6t
Xbit_r93_c1 bl[1] br[1] wl[93] vdd gnd cell_6t
Xbit_r94_c1 bl[1] br[1] wl[94] vdd gnd cell_6t
Xbit_r95_c1 bl[1] br[1] wl[95] vdd gnd cell_6t
Xbit_r96_c1 bl[1] br[1] wl[96] vdd gnd cell_6t
Xbit_r97_c1 bl[1] br[1] wl[97] vdd gnd cell_6t
Xbit_r98_c1 bl[1] br[1] wl[98] vdd gnd cell_6t
Xbit_r99_c1 bl[1] br[1] wl[99] vdd gnd cell_6t
Xbit_r100_c1 bl[1] br[1] wl[100] vdd gnd cell_6t
Xbit_r101_c1 bl[1] br[1] wl[101] vdd gnd cell_6t
Xbit_r102_c1 bl[1] br[1] wl[102] vdd gnd cell_6t
Xbit_r103_c1 bl[1] br[1] wl[103] vdd gnd cell_6t
Xbit_r104_c1 bl[1] br[1] wl[104] vdd gnd cell_6t
Xbit_r105_c1 bl[1] br[1] wl[105] vdd gnd cell_6t
Xbit_r106_c1 bl[1] br[1] wl[106] vdd gnd cell_6t
Xbit_r107_c1 bl[1] br[1] wl[107] vdd gnd cell_6t
Xbit_r108_c1 bl[1] br[1] wl[108] vdd gnd cell_6t
Xbit_r109_c1 bl[1] br[1] wl[109] vdd gnd cell_6t
Xbit_r110_c1 bl[1] br[1] wl[110] vdd gnd cell_6t
Xbit_r111_c1 bl[1] br[1] wl[111] vdd gnd cell_6t
Xbit_r112_c1 bl[1] br[1] wl[112] vdd gnd cell_6t
Xbit_r113_c1 bl[1] br[1] wl[113] vdd gnd cell_6t
Xbit_r114_c1 bl[1] br[1] wl[114] vdd gnd cell_6t
Xbit_r115_c1 bl[1] br[1] wl[115] vdd gnd cell_6t
Xbit_r116_c1 bl[1] br[1] wl[116] vdd gnd cell_6t
Xbit_r117_c1 bl[1] br[1] wl[117] vdd gnd cell_6t
Xbit_r118_c1 bl[1] br[1] wl[118] vdd gnd cell_6t
Xbit_r119_c1 bl[1] br[1] wl[119] vdd gnd cell_6t
Xbit_r120_c1 bl[1] br[1] wl[120] vdd gnd cell_6t
Xbit_r121_c1 bl[1] br[1] wl[121] vdd gnd cell_6t
Xbit_r122_c1 bl[1] br[1] wl[122] vdd gnd cell_6t
Xbit_r123_c1 bl[1] br[1] wl[123] vdd gnd cell_6t
Xbit_r124_c1 bl[1] br[1] wl[124] vdd gnd cell_6t
Xbit_r125_c1 bl[1] br[1] wl[125] vdd gnd cell_6t
Xbit_r126_c1 bl[1] br[1] wl[126] vdd gnd cell_6t
Xbit_r127_c1 bl[1] br[1] wl[127] vdd gnd cell_6t
Xbit_r128_c1 bl[1] br[1] wl[128] vdd gnd cell_6t
Xbit_r129_c1 bl[1] br[1] wl[129] vdd gnd cell_6t
Xbit_r130_c1 bl[1] br[1] wl[130] vdd gnd cell_6t
Xbit_r131_c1 bl[1] br[1] wl[131] vdd gnd cell_6t
Xbit_r132_c1 bl[1] br[1] wl[132] vdd gnd cell_6t
Xbit_r133_c1 bl[1] br[1] wl[133] vdd gnd cell_6t
Xbit_r134_c1 bl[1] br[1] wl[134] vdd gnd cell_6t
Xbit_r135_c1 bl[1] br[1] wl[135] vdd gnd cell_6t
Xbit_r136_c1 bl[1] br[1] wl[136] vdd gnd cell_6t
Xbit_r137_c1 bl[1] br[1] wl[137] vdd gnd cell_6t
Xbit_r138_c1 bl[1] br[1] wl[138] vdd gnd cell_6t
Xbit_r139_c1 bl[1] br[1] wl[139] vdd gnd cell_6t
Xbit_r140_c1 bl[1] br[1] wl[140] vdd gnd cell_6t
Xbit_r141_c1 bl[1] br[1] wl[141] vdd gnd cell_6t
Xbit_r142_c1 bl[1] br[1] wl[142] vdd gnd cell_6t
Xbit_r143_c1 bl[1] br[1] wl[143] vdd gnd cell_6t
Xbit_r144_c1 bl[1] br[1] wl[144] vdd gnd cell_6t
Xbit_r145_c1 bl[1] br[1] wl[145] vdd gnd cell_6t
Xbit_r146_c1 bl[1] br[1] wl[146] vdd gnd cell_6t
Xbit_r147_c1 bl[1] br[1] wl[147] vdd gnd cell_6t
Xbit_r148_c1 bl[1] br[1] wl[148] vdd gnd cell_6t
Xbit_r149_c1 bl[1] br[1] wl[149] vdd gnd cell_6t
Xbit_r150_c1 bl[1] br[1] wl[150] vdd gnd cell_6t
Xbit_r151_c1 bl[1] br[1] wl[151] vdd gnd cell_6t
Xbit_r152_c1 bl[1] br[1] wl[152] vdd gnd cell_6t
Xbit_r153_c1 bl[1] br[1] wl[153] vdd gnd cell_6t
Xbit_r154_c1 bl[1] br[1] wl[154] vdd gnd cell_6t
Xbit_r155_c1 bl[1] br[1] wl[155] vdd gnd cell_6t
Xbit_r156_c1 bl[1] br[1] wl[156] vdd gnd cell_6t
Xbit_r157_c1 bl[1] br[1] wl[157] vdd gnd cell_6t
Xbit_r158_c1 bl[1] br[1] wl[158] vdd gnd cell_6t
Xbit_r159_c1 bl[1] br[1] wl[159] vdd gnd cell_6t
Xbit_r160_c1 bl[1] br[1] wl[160] vdd gnd cell_6t
Xbit_r161_c1 bl[1] br[1] wl[161] vdd gnd cell_6t
Xbit_r162_c1 bl[1] br[1] wl[162] vdd gnd cell_6t
Xbit_r163_c1 bl[1] br[1] wl[163] vdd gnd cell_6t
Xbit_r164_c1 bl[1] br[1] wl[164] vdd gnd cell_6t
Xbit_r165_c1 bl[1] br[1] wl[165] vdd gnd cell_6t
Xbit_r166_c1 bl[1] br[1] wl[166] vdd gnd cell_6t
Xbit_r167_c1 bl[1] br[1] wl[167] vdd gnd cell_6t
Xbit_r168_c1 bl[1] br[1] wl[168] vdd gnd cell_6t
Xbit_r169_c1 bl[1] br[1] wl[169] vdd gnd cell_6t
Xbit_r170_c1 bl[1] br[1] wl[170] vdd gnd cell_6t
Xbit_r171_c1 bl[1] br[1] wl[171] vdd gnd cell_6t
Xbit_r172_c1 bl[1] br[1] wl[172] vdd gnd cell_6t
Xbit_r173_c1 bl[1] br[1] wl[173] vdd gnd cell_6t
Xbit_r174_c1 bl[1] br[1] wl[174] vdd gnd cell_6t
Xbit_r175_c1 bl[1] br[1] wl[175] vdd gnd cell_6t
Xbit_r176_c1 bl[1] br[1] wl[176] vdd gnd cell_6t
Xbit_r177_c1 bl[1] br[1] wl[177] vdd gnd cell_6t
Xbit_r178_c1 bl[1] br[1] wl[178] vdd gnd cell_6t
Xbit_r179_c1 bl[1] br[1] wl[179] vdd gnd cell_6t
Xbit_r180_c1 bl[1] br[1] wl[180] vdd gnd cell_6t
Xbit_r181_c1 bl[1] br[1] wl[181] vdd gnd cell_6t
Xbit_r182_c1 bl[1] br[1] wl[182] vdd gnd cell_6t
Xbit_r183_c1 bl[1] br[1] wl[183] vdd gnd cell_6t
Xbit_r184_c1 bl[1] br[1] wl[184] vdd gnd cell_6t
Xbit_r185_c1 bl[1] br[1] wl[185] vdd gnd cell_6t
Xbit_r186_c1 bl[1] br[1] wl[186] vdd gnd cell_6t
Xbit_r187_c1 bl[1] br[1] wl[187] vdd gnd cell_6t
Xbit_r188_c1 bl[1] br[1] wl[188] vdd gnd cell_6t
Xbit_r189_c1 bl[1] br[1] wl[189] vdd gnd cell_6t
Xbit_r190_c1 bl[1] br[1] wl[190] vdd gnd cell_6t
Xbit_r191_c1 bl[1] br[1] wl[191] vdd gnd cell_6t
Xbit_r192_c1 bl[1] br[1] wl[192] vdd gnd cell_6t
Xbit_r193_c1 bl[1] br[1] wl[193] vdd gnd cell_6t
Xbit_r194_c1 bl[1] br[1] wl[194] vdd gnd cell_6t
Xbit_r195_c1 bl[1] br[1] wl[195] vdd gnd cell_6t
Xbit_r196_c1 bl[1] br[1] wl[196] vdd gnd cell_6t
Xbit_r197_c1 bl[1] br[1] wl[197] vdd gnd cell_6t
Xbit_r198_c1 bl[1] br[1] wl[198] vdd gnd cell_6t
Xbit_r199_c1 bl[1] br[1] wl[199] vdd gnd cell_6t
Xbit_r200_c1 bl[1] br[1] wl[200] vdd gnd cell_6t
Xbit_r201_c1 bl[1] br[1] wl[201] vdd gnd cell_6t
Xbit_r202_c1 bl[1] br[1] wl[202] vdd gnd cell_6t
Xbit_r203_c1 bl[1] br[1] wl[203] vdd gnd cell_6t
Xbit_r204_c1 bl[1] br[1] wl[204] vdd gnd cell_6t
Xbit_r205_c1 bl[1] br[1] wl[205] vdd gnd cell_6t
Xbit_r206_c1 bl[1] br[1] wl[206] vdd gnd cell_6t
Xbit_r207_c1 bl[1] br[1] wl[207] vdd gnd cell_6t
Xbit_r208_c1 bl[1] br[1] wl[208] vdd gnd cell_6t
Xbit_r209_c1 bl[1] br[1] wl[209] vdd gnd cell_6t
Xbit_r210_c1 bl[1] br[1] wl[210] vdd gnd cell_6t
Xbit_r211_c1 bl[1] br[1] wl[211] vdd gnd cell_6t
Xbit_r212_c1 bl[1] br[1] wl[212] vdd gnd cell_6t
Xbit_r213_c1 bl[1] br[1] wl[213] vdd gnd cell_6t
Xbit_r214_c1 bl[1] br[1] wl[214] vdd gnd cell_6t
Xbit_r215_c1 bl[1] br[1] wl[215] vdd gnd cell_6t
Xbit_r216_c1 bl[1] br[1] wl[216] vdd gnd cell_6t
Xbit_r217_c1 bl[1] br[1] wl[217] vdd gnd cell_6t
Xbit_r218_c1 bl[1] br[1] wl[218] vdd gnd cell_6t
Xbit_r219_c1 bl[1] br[1] wl[219] vdd gnd cell_6t
Xbit_r220_c1 bl[1] br[1] wl[220] vdd gnd cell_6t
Xbit_r221_c1 bl[1] br[1] wl[221] vdd gnd cell_6t
Xbit_r222_c1 bl[1] br[1] wl[222] vdd gnd cell_6t
Xbit_r223_c1 bl[1] br[1] wl[223] vdd gnd cell_6t
Xbit_r224_c1 bl[1] br[1] wl[224] vdd gnd cell_6t
Xbit_r225_c1 bl[1] br[1] wl[225] vdd gnd cell_6t
Xbit_r226_c1 bl[1] br[1] wl[226] vdd gnd cell_6t
Xbit_r227_c1 bl[1] br[1] wl[227] vdd gnd cell_6t
Xbit_r228_c1 bl[1] br[1] wl[228] vdd gnd cell_6t
Xbit_r229_c1 bl[1] br[1] wl[229] vdd gnd cell_6t
Xbit_r230_c1 bl[1] br[1] wl[230] vdd gnd cell_6t
Xbit_r231_c1 bl[1] br[1] wl[231] vdd gnd cell_6t
Xbit_r232_c1 bl[1] br[1] wl[232] vdd gnd cell_6t
Xbit_r233_c1 bl[1] br[1] wl[233] vdd gnd cell_6t
Xbit_r234_c1 bl[1] br[1] wl[234] vdd gnd cell_6t
Xbit_r235_c1 bl[1] br[1] wl[235] vdd gnd cell_6t
Xbit_r236_c1 bl[1] br[1] wl[236] vdd gnd cell_6t
Xbit_r237_c1 bl[1] br[1] wl[237] vdd gnd cell_6t
Xbit_r238_c1 bl[1] br[1] wl[238] vdd gnd cell_6t
Xbit_r239_c1 bl[1] br[1] wl[239] vdd gnd cell_6t
Xbit_r240_c1 bl[1] br[1] wl[240] vdd gnd cell_6t
Xbit_r241_c1 bl[1] br[1] wl[241] vdd gnd cell_6t
Xbit_r242_c1 bl[1] br[1] wl[242] vdd gnd cell_6t
Xbit_r243_c1 bl[1] br[1] wl[243] vdd gnd cell_6t
Xbit_r244_c1 bl[1] br[1] wl[244] vdd gnd cell_6t
Xbit_r245_c1 bl[1] br[1] wl[245] vdd gnd cell_6t
Xbit_r246_c1 bl[1] br[1] wl[246] vdd gnd cell_6t
Xbit_r247_c1 bl[1] br[1] wl[247] vdd gnd cell_6t
Xbit_r248_c1 bl[1] br[1] wl[248] vdd gnd cell_6t
Xbit_r249_c1 bl[1] br[1] wl[249] vdd gnd cell_6t
Xbit_r250_c1 bl[1] br[1] wl[250] vdd gnd cell_6t
Xbit_r251_c1 bl[1] br[1] wl[251] vdd gnd cell_6t
Xbit_r252_c1 bl[1] br[1] wl[252] vdd gnd cell_6t
Xbit_r253_c1 bl[1] br[1] wl[253] vdd gnd cell_6t
Xbit_r254_c1 bl[1] br[1] wl[254] vdd gnd cell_6t
Xbit_r255_c1 bl[1] br[1] wl[255] vdd gnd cell_6t
Xbit_r256_c1 bl[1] br[1] wl[256] vdd gnd cell_6t
Xbit_r257_c1 bl[1] br[1] wl[257] vdd gnd cell_6t
Xbit_r258_c1 bl[1] br[1] wl[258] vdd gnd cell_6t
Xbit_r259_c1 bl[1] br[1] wl[259] vdd gnd cell_6t
Xbit_r260_c1 bl[1] br[1] wl[260] vdd gnd cell_6t
Xbit_r261_c1 bl[1] br[1] wl[261] vdd gnd cell_6t
Xbit_r262_c1 bl[1] br[1] wl[262] vdd gnd cell_6t
Xbit_r263_c1 bl[1] br[1] wl[263] vdd gnd cell_6t
Xbit_r264_c1 bl[1] br[1] wl[264] vdd gnd cell_6t
Xbit_r265_c1 bl[1] br[1] wl[265] vdd gnd cell_6t
Xbit_r266_c1 bl[1] br[1] wl[266] vdd gnd cell_6t
Xbit_r267_c1 bl[1] br[1] wl[267] vdd gnd cell_6t
Xbit_r268_c1 bl[1] br[1] wl[268] vdd gnd cell_6t
Xbit_r269_c1 bl[1] br[1] wl[269] vdd gnd cell_6t
Xbit_r270_c1 bl[1] br[1] wl[270] vdd gnd cell_6t
Xbit_r271_c1 bl[1] br[1] wl[271] vdd gnd cell_6t
Xbit_r272_c1 bl[1] br[1] wl[272] vdd gnd cell_6t
Xbit_r273_c1 bl[1] br[1] wl[273] vdd gnd cell_6t
Xbit_r274_c1 bl[1] br[1] wl[274] vdd gnd cell_6t
Xbit_r275_c1 bl[1] br[1] wl[275] vdd gnd cell_6t
Xbit_r276_c1 bl[1] br[1] wl[276] vdd gnd cell_6t
Xbit_r277_c1 bl[1] br[1] wl[277] vdd gnd cell_6t
Xbit_r278_c1 bl[1] br[1] wl[278] vdd gnd cell_6t
Xbit_r279_c1 bl[1] br[1] wl[279] vdd gnd cell_6t
Xbit_r280_c1 bl[1] br[1] wl[280] vdd gnd cell_6t
Xbit_r281_c1 bl[1] br[1] wl[281] vdd gnd cell_6t
Xbit_r282_c1 bl[1] br[1] wl[282] vdd gnd cell_6t
Xbit_r283_c1 bl[1] br[1] wl[283] vdd gnd cell_6t
Xbit_r284_c1 bl[1] br[1] wl[284] vdd gnd cell_6t
Xbit_r285_c1 bl[1] br[1] wl[285] vdd gnd cell_6t
Xbit_r286_c1 bl[1] br[1] wl[286] vdd gnd cell_6t
Xbit_r287_c1 bl[1] br[1] wl[287] vdd gnd cell_6t
Xbit_r288_c1 bl[1] br[1] wl[288] vdd gnd cell_6t
Xbit_r289_c1 bl[1] br[1] wl[289] vdd gnd cell_6t
Xbit_r290_c1 bl[1] br[1] wl[290] vdd gnd cell_6t
Xbit_r291_c1 bl[1] br[1] wl[291] vdd gnd cell_6t
Xbit_r292_c1 bl[1] br[1] wl[292] vdd gnd cell_6t
Xbit_r293_c1 bl[1] br[1] wl[293] vdd gnd cell_6t
Xbit_r294_c1 bl[1] br[1] wl[294] vdd gnd cell_6t
Xbit_r295_c1 bl[1] br[1] wl[295] vdd gnd cell_6t
Xbit_r296_c1 bl[1] br[1] wl[296] vdd gnd cell_6t
Xbit_r297_c1 bl[1] br[1] wl[297] vdd gnd cell_6t
Xbit_r298_c1 bl[1] br[1] wl[298] vdd gnd cell_6t
Xbit_r299_c1 bl[1] br[1] wl[299] vdd gnd cell_6t
Xbit_r300_c1 bl[1] br[1] wl[300] vdd gnd cell_6t
Xbit_r301_c1 bl[1] br[1] wl[301] vdd gnd cell_6t
Xbit_r302_c1 bl[1] br[1] wl[302] vdd gnd cell_6t
Xbit_r303_c1 bl[1] br[1] wl[303] vdd gnd cell_6t
Xbit_r304_c1 bl[1] br[1] wl[304] vdd gnd cell_6t
Xbit_r305_c1 bl[1] br[1] wl[305] vdd gnd cell_6t
Xbit_r306_c1 bl[1] br[1] wl[306] vdd gnd cell_6t
Xbit_r307_c1 bl[1] br[1] wl[307] vdd gnd cell_6t
Xbit_r308_c1 bl[1] br[1] wl[308] vdd gnd cell_6t
Xbit_r309_c1 bl[1] br[1] wl[309] vdd gnd cell_6t
Xbit_r310_c1 bl[1] br[1] wl[310] vdd gnd cell_6t
Xbit_r311_c1 bl[1] br[1] wl[311] vdd gnd cell_6t
Xbit_r312_c1 bl[1] br[1] wl[312] vdd gnd cell_6t
Xbit_r313_c1 bl[1] br[1] wl[313] vdd gnd cell_6t
Xbit_r314_c1 bl[1] br[1] wl[314] vdd gnd cell_6t
Xbit_r315_c1 bl[1] br[1] wl[315] vdd gnd cell_6t
Xbit_r316_c1 bl[1] br[1] wl[316] vdd gnd cell_6t
Xbit_r317_c1 bl[1] br[1] wl[317] vdd gnd cell_6t
Xbit_r318_c1 bl[1] br[1] wl[318] vdd gnd cell_6t
Xbit_r319_c1 bl[1] br[1] wl[319] vdd gnd cell_6t
Xbit_r320_c1 bl[1] br[1] wl[320] vdd gnd cell_6t
Xbit_r321_c1 bl[1] br[1] wl[321] vdd gnd cell_6t
Xbit_r322_c1 bl[1] br[1] wl[322] vdd gnd cell_6t
Xbit_r323_c1 bl[1] br[1] wl[323] vdd gnd cell_6t
Xbit_r324_c1 bl[1] br[1] wl[324] vdd gnd cell_6t
Xbit_r325_c1 bl[1] br[1] wl[325] vdd gnd cell_6t
Xbit_r326_c1 bl[1] br[1] wl[326] vdd gnd cell_6t
Xbit_r327_c1 bl[1] br[1] wl[327] vdd gnd cell_6t
Xbit_r328_c1 bl[1] br[1] wl[328] vdd gnd cell_6t
Xbit_r329_c1 bl[1] br[1] wl[329] vdd gnd cell_6t
Xbit_r330_c1 bl[1] br[1] wl[330] vdd gnd cell_6t
Xbit_r331_c1 bl[1] br[1] wl[331] vdd gnd cell_6t
Xbit_r332_c1 bl[1] br[1] wl[332] vdd gnd cell_6t
Xbit_r333_c1 bl[1] br[1] wl[333] vdd gnd cell_6t
Xbit_r334_c1 bl[1] br[1] wl[334] vdd gnd cell_6t
Xbit_r335_c1 bl[1] br[1] wl[335] vdd gnd cell_6t
Xbit_r336_c1 bl[1] br[1] wl[336] vdd gnd cell_6t
Xbit_r337_c1 bl[1] br[1] wl[337] vdd gnd cell_6t
Xbit_r338_c1 bl[1] br[1] wl[338] vdd gnd cell_6t
Xbit_r339_c1 bl[1] br[1] wl[339] vdd gnd cell_6t
Xbit_r340_c1 bl[1] br[1] wl[340] vdd gnd cell_6t
Xbit_r341_c1 bl[1] br[1] wl[341] vdd gnd cell_6t
Xbit_r342_c1 bl[1] br[1] wl[342] vdd gnd cell_6t
Xbit_r343_c1 bl[1] br[1] wl[343] vdd gnd cell_6t
Xbit_r344_c1 bl[1] br[1] wl[344] vdd gnd cell_6t
Xbit_r345_c1 bl[1] br[1] wl[345] vdd gnd cell_6t
Xbit_r346_c1 bl[1] br[1] wl[346] vdd gnd cell_6t
Xbit_r347_c1 bl[1] br[1] wl[347] vdd gnd cell_6t
Xbit_r348_c1 bl[1] br[1] wl[348] vdd gnd cell_6t
Xbit_r349_c1 bl[1] br[1] wl[349] vdd gnd cell_6t
Xbit_r350_c1 bl[1] br[1] wl[350] vdd gnd cell_6t
Xbit_r351_c1 bl[1] br[1] wl[351] vdd gnd cell_6t
Xbit_r352_c1 bl[1] br[1] wl[352] vdd gnd cell_6t
Xbit_r353_c1 bl[1] br[1] wl[353] vdd gnd cell_6t
Xbit_r354_c1 bl[1] br[1] wl[354] vdd gnd cell_6t
Xbit_r355_c1 bl[1] br[1] wl[355] vdd gnd cell_6t
Xbit_r356_c1 bl[1] br[1] wl[356] vdd gnd cell_6t
Xbit_r357_c1 bl[1] br[1] wl[357] vdd gnd cell_6t
Xbit_r358_c1 bl[1] br[1] wl[358] vdd gnd cell_6t
Xbit_r359_c1 bl[1] br[1] wl[359] vdd gnd cell_6t
Xbit_r360_c1 bl[1] br[1] wl[360] vdd gnd cell_6t
Xbit_r361_c1 bl[1] br[1] wl[361] vdd gnd cell_6t
Xbit_r362_c1 bl[1] br[1] wl[362] vdd gnd cell_6t
Xbit_r363_c1 bl[1] br[1] wl[363] vdd gnd cell_6t
Xbit_r364_c1 bl[1] br[1] wl[364] vdd gnd cell_6t
Xbit_r365_c1 bl[1] br[1] wl[365] vdd gnd cell_6t
Xbit_r366_c1 bl[1] br[1] wl[366] vdd gnd cell_6t
Xbit_r367_c1 bl[1] br[1] wl[367] vdd gnd cell_6t
Xbit_r368_c1 bl[1] br[1] wl[368] vdd gnd cell_6t
Xbit_r369_c1 bl[1] br[1] wl[369] vdd gnd cell_6t
Xbit_r370_c1 bl[1] br[1] wl[370] vdd gnd cell_6t
Xbit_r371_c1 bl[1] br[1] wl[371] vdd gnd cell_6t
Xbit_r372_c1 bl[1] br[1] wl[372] vdd gnd cell_6t
Xbit_r373_c1 bl[1] br[1] wl[373] vdd gnd cell_6t
Xbit_r374_c1 bl[1] br[1] wl[374] vdd gnd cell_6t
Xbit_r375_c1 bl[1] br[1] wl[375] vdd gnd cell_6t
Xbit_r376_c1 bl[1] br[1] wl[376] vdd gnd cell_6t
Xbit_r377_c1 bl[1] br[1] wl[377] vdd gnd cell_6t
Xbit_r378_c1 bl[1] br[1] wl[378] vdd gnd cell_6t
Xbit_r379_c1 bl[1] br[1] wl[379] vdd gnd cell_6t
Xbit_r380_c1 bl[1] br[1] wl[380] vdd gnd cell_6t
Xbit_r381_c1 bl[1] br[1] wl[381] vdd gnd cell_6t
Xbit_r382_c1 bl[1] br[1] wl[382] vdd gnd cell_6t
Xbit_r383_c1 bl[1] br[1] wl[383] vdd gnd cell_6t
Xbit_r384_c1 bl[1] br[1] wl[384] vdd gnd cell_6t
Xbit_r385_c1 bl[1] br[1] wl[385] vdd gnd cell_6t
Xbit_r386_c1 bl[1] br[1] wl[386] vdd gnd cell_6t
Xbit_r387_c1 bl[1] br[1] wl[387] vdd gnd cell_6t
Xbit_r388_c1 bl[1] br[1] wl[388] vdd gnd cell_6t
Xbit_r389_c1 bl[1] br[1] wl[389] vdd gnd cell_6t
Xbit_r390_c1 bl[1] br[1] wl[390] vdd gnd cell_6t
Xbit_r391_c1 bl[1] br[1] wl[391] vdd gnd cell_6t
Xbit_r392_c1 bl[1] br[1] wl[392] vdd gnd cell_6t
Xbit_r393_c1 bl[1] br[1] wl[393] vdd gnd cell_6t
Xbit_r394_c1 bl[1] br[1] wl[394] vdd gnd cell_6t
Xbit_r395_c1 bl[1] br[1] wl[395] vdd gnd cell_6t
Xbit_r396_c1 bl[1] br[1] wl[396] vdd gnd cell_6t
Xbit_r397_c1 bl[1] br[1] wl[397] vdd gnd cell_6t
Xbit_r398_c1 bl[1] br[1] wl[398] vdd gnd cell_6t
Xbit_r399_c1 bl[1] br[1] wl[399] vdd gnd cell_6t
Xbit_r400_c1 bl[1] br[1] wl[400] vdd gnd cell_6t
Xbit_r401_c1 bl[1] br[1] wl[401] vdd gnd cell_6t
Xbit_r402_c1 bl[1] br[1] wl[402] vdd gnd cell_6t
Xbit_r403_c1 bl[1] br[1] wl[403] vdd gnd cell_6t
Xbit_r404_c1 bl[1] br[1] wl[404] vdd gnd cell_6t
Xbit_r405_c1 bl[1] br[1] wl[405] vdd gnd cell_6t
Xbit_r406_c1 bl[1] br[1] wl[406] vdd gnd cell_6t
Xbit_r407_c1 bl[1] br[1] wl[407] vdd gnd cell_6t
Xbit_r408_c1 bl[1] br[1] wl[408] vdd gnd cell_6t
Xbit_r409_c1 bl[1] br[1] wl[409] vdd gnd cell_6t
Xbit_r410_c1 bl[1] br[1] wl[410] vdd gnd cell_6t
Xbit_r411_c1 bl[1] br[1] wl[411] vdd gnd cell_6t
Xbit_r412_c1 bl[1] br[1] wl[412] vdd gnd cell_6t
Xbit_r413_c1 bl[1] br[1] wl[413] vdd gnd cell_6t
Xbit_r414_c1 bl[1] br[1] wl[414] vdd gnd cell_6t
Xbit_r415_c1 bl[1] br[1] wl[415] vdd gnd cell_6t
Xbit_r416_c1 bl[1] br[1] wl[416] vdd gnd cell_6t
Xbit_r417_c1 bl[1] br[1] wl[417] vdd gnd cell_6t
Xbit_r418_c1 bl[1] br[1] wl[418] vdd gnd cell_6t
Xbit_r419_c1 bl[1] br[1] wl[419] vdd gnd cell_6t
Xbit_r420_c1 bl[1] br[1] wl[420] vdd gnd cell_6t
Xbit_r421_c1 bl[1] br[1] wl[421] vdd gnd cell_6t
Xbit_r422_c1 bl[1] br[1] wl[422] vdd gnd cell_6t
Xbit_r423_c1 bl[1] br[1] wl[423] vdd gnd cell_6t
Xbit_r424_c1 bl[1] br[1] wl[424] vdd gnd cell_6t
Xbit_r425_c1 bl[1] br[1] wl[425] vdd gnd cell_6t
Xbit_r426_c1 bl[1] br[1] wl[426] vdd gnd cell_6t
Xbit_r427_c1 bl[1] br[1] wl[427] vdd gnd cell_6t
Xbit_r428_c1 bl[1] br[1] wl[428] vdd gnd cell_6t
Xbit_r429_c1 bl[1] br[1] wl[429] vdd gnd cell_6t
Xbit_r430_c1 bl[1] br[1] wl[430] vdd gnd cell_6t
Xbit_r431_c1 bl[1] br[1] wl[431] vdd gnd cell_6t
Xbit_r432_c1 bl[1] br[1] wl[432] vdd gnd cell_6t
Xbit_r433_c1 bl[1] br[1] wl[433] vdd gnd cell_6t
Xbit_r434_c1 bl[1] br[1] wl[434] vdd gnd cell_6t
Xbit_r435_c1 bl[1] br[1] wl[435] vdd gnd cell_6t
Xbit_r436_c1 bl[1] br[1] wl[436] vdd gnd cell_6t
Xbit_r437_c1 bl[1] br[1] wl[437] vdd gnd cell_6t
Xbit_r438_c1 bl[1] br[1] wl[438] vdd gnd cell_6t
Xbit_r439_c1 bl[1] br[1] wl[439] vdd gnd cell_6t
Xbit_r440_c1 bl[1] br[1] wl[440] vdd gnd cell_6t
Xbit_r441_c1 bl[1] br[1] wl[441] vdd gnd cell_6t
Xbit_r442_c1 bl[1] br[1] wl[442] vdd gnd cell_6t
Xbit_r443_c1 bl[1] br[1] wl[443] vdd gnd cell_6t
Xbit_r444_c1 bl[1] br[1] wl[444] vdd gnd cell_6t
Xbit_r445_c1 bl[1] br[1] wl[445] vdd gnd cell_6t
Xbit_r446_c1 bl[1] br[1] wl[446] vdd gnd cell_6t
Xbit_r447_c1 bl[1] br[1] wl[447] vdd gnd cell_6t
Xbit_r448_c1 bl[1] br[1] wl[448] vdd gnd cell_6t
Xbit_r449_c1 bl[1] br[1] wl[449] vdd gnd cell_6t
Xbit_r450_c1 bl[1] br[1] wl[450] vdd gnd cell_6t
Xbit_r451_c1 bl[1] br[1] wl[451] vdd gnd cell_6t
Xbit_r452_c1 bl[1] br[1] wl[452] vdd gnd cell_6t
Xbit_r453_c1 bl[1] br[1] wl[453] vdd gnd cell_6t
Xbit_r454_c1 bl[1] br[1] wl[454] vdd gnd cell_6t
Xbit_r455_c1 bl[1] br[1] wl[455] vdd gnd cell_6t
Xbit_r456_c1 bl[1] br[1] wl[456] vdd gnd cell_6t
Xbit_r457_c1 bl[1] br[1] wl[457] vdd gnd cell_6t
Xbit_r458_c1 bl[1] br[1] wl[458] vdd gnd cell_6t
Xbit_r459_c1 bl[1] br[1] wl[459] vdd gnd cell_6t
Xbit_r460_c1 bl[1] br[1] wl[460] vdd gnd cell_6t
Xbit_r461_c1 bl[1] br[1] wl[461] vdd gnd cell_6t
Xbit_r462_c1 bl[1] br[1] wl[462] vdd gnd cell_6t
Xbit_r463_c1 bl[1] br[1] wl[463] vdd gnd cell_6t
Xbit_r464_c1 bl[1] br[1] wl[464] vdd gnd cell_6t
Xbit_r465_c1 bl[1] br[1] wl[465] vdd gnd cell_6t
Xbit_r466_c1 bl[1] br[1] wl[466] vdd gnd cell_6t
Xbit_r467_c1 bl[1] br[1] wl[467] vdd gnd cell_6t
Xbit_r468_c1 bl[1] br[1] wl[468] vdd gnd cell_6t
Xbit_r469_c1 bl[1] br[1] wl[469] vdd gnd cell_6t
Xbit_r470_c1 bl[1] br[1] wl[470] vdd gnd cell_6t
Xbit_r471_c1 bl[1] br[1] wl[471] vdd gnd cell_6t
Xbit_r472_c1 bl[1] br[1] wl[472] vdd gnd cell_6t
Xbit_r473_c1 bl[1] br[1] wl[473] vdd gnd cell_6t
Xbit_r474_c1 bl[1] br[1] wl[474] vdd gnd cell_6t
Xbit_r475_c1 bl[1] br[1] wl[475] vdd gnd cell_6t
Xbit_r476_c1 bl[1] br[1] wl[476] vdd gnd cell_6t
Xbit_r477_c1 bl[1] br[1] wl[477] vdd gnd cell_6t
Xbit_r478_c1 bl[1] br[1] wl[478] vdd gnd cell_6t
Xbit_r479_c1 bl[1] br[1] wl[479] vdd gnd cell_6t
Xbit_r480_c1 bl[1] br[1] wl[480] vdd gnd cell_6t
Xbit_r481_c1 bl[1] br[1] wl[481] vdd gnd cell_6t
Xbit_r482_c1 bl[1] br[1] wl[482] vdd gnd cell_6t
Xbit_r483_c1 bl[1] br[1] wl[483] vdd gnd cell_6t
Xbit_r484_c1 bl[1] br[1] wl[484] vdd gnd cell_6t
Xbit_r485_c1 bl[1] br[1] wl[485] vdd gnd cell_6t
Xbit_r486_c1 bl[1] br[1] wl[486] vdd gnd cell_6t
Xbit_r487_c1 bl[1] br[1] wl[487] vdd gnd cell_6t
Xbit_r488_c1 bl[1] br[1] wl[488] vdd gnd cell_6t
Xbit_r489_c1 bl[1] br[1] wl[489] vdd gnd cell_6t
Xbit_r490_c1 bl[1] br[1] wl[490] vdd gnd cell_6t
Xbit_r491_c1 bl[1] br[1] wl[491] vdd gnd cell_6t
Xbit_r492_c1 bl[1] br[1] wl[492] vdd gnd cell_6t
Xbit_r493_c1 bl[1] br[1] wl[493] vdd gnd cell_6t
Xbit_r494_c1 bl[1] br[1] wl[494] vdd gnd cell_6t
Xbit_r495_c1 bl[1] br[1] wl[495] vdd gnd cell_6t
Xbit_r496_c1 bl[1] br[1] wl[496] vdd gnd cell_6t
Xbit_r497_c1 bl[1] br[1] wl[497] vdd gnd cell_6t
Xbit_r498_c1 bl[1] br[1] wl[498] vdd gnd cell_6t
Xbit_r499_c1 bl[1] br[1] wl[499] vdd gnd cell_6t
Xbit_r500_c1 bl[1] br[1] wl[500] vdd gnd cell_6t
Xbit_r501_c1 bl[1] br[1] wl[501] vdd gnd cell_6t
Xbit_r502_c1 bl[1] br[1] wl[502] vdd gnd cell_6t
Xbit_r503_c1 bl[1] br[1] wl[503] vdd gnd cell_6t
Xbit_r504_c1 bl[1] br[1] wl[504] vdd gnd cell_6t
Xbit_r505_c1 bl[1] br[1] wl[505] vdd gnd cell_6t
Xbit_r506_c1 bl[1] br[1] wl[506] vdd gnd cell_6t
Xbit_r507_c1 bl[1] br[1] wl[507] vdd gnd cell_6t
Xbit_r508_c1 bl[1] br[1] wl[508] vdd gnd cell_6t
Xbit_r509_c1 bl[1] br[1] wl[509] vdd gnd cell_6t
Xbit_r510_c1 bl[1] br[1] wl[510] vdd gnd cell_6t
Xbit_r511_c1 bl[1] br[1] wl[511] vdd gnd cell_6t
Xbit_r0_c2 bl[2] br[2] wl[0] vdd gnd cell_6t
Xbit_r1_c2 bl[2] br[2] wl[1] vdd gnd cell_6t
Xbit_r2_c2 bl[2] br[2] wl[2] vdd gnd cell_6t
Xbit_r3_c2 bl[2] br[2] wl[3] vdd gnd cell_6t
Xbit_r4_c2 bl[2] br[2] wl[4] vdd gnd cell_6t
Xbit_r5_c2 bl[2] br[2] wl[5] vdd gnd cell_6t
Xbit_r6_c2 bl[2] br[2] wl[6] vdd gnd cell_6t
Xbit_r7_c2 bl[2] br[2] wl[7] vdd gnd cell_6t
Xbit_r8_c2 bl[2] br[2] wl[8] vdd gnd cell_6t
Xbit_r9_c2 bl[2] br[2] wl[9] vdd gnd cell_6t
Xbit_r10_c2 bl[2] br[2] wl[10] vdd gnd cell_6t
Xbit_r11_c2 bl[2] br[2] wl[11] vdd gnd cell_6t
Xbit_r12_c2 bl[2] br[2] wl[12] vdd gnd cell_6t
Xbit_r13_c2 bl[2] br[2] wl[13] vdd gnd cell_6t
Xbit_r14_c2 bl[2] br[2] wl[14] vdd gnd cell_6t
Xbit_r15_c2 bl[2] br[2] wl[15] vdd gnd cell_6t
Xbit_r16_c2 bl[2] br[2] wl[16] vdd gnd cell_6t
Xbit_r17_c2 bl[2] br[2] wl[17] vdd gnd cell_6t
Xbit_r18_c2 bl[2] br[2] wl[18] vdd gnd cell_6t
Xbit_r19_c2 bl[2] br[2] wl[19] vdd gnd cell_6t
Xbit_r20_c2 bl[2] br[2] wl[20] vdd gnd cell_6t
Xbit_r21_c2 bl[2] br[2] wl[21] vdd gnd cell_6t
Xbit_r22_c2 bl[2] br[2] wl[22] vdd gnd cell_6t
Xbit_r23_c2 bl[2] br[2] wl[23] vdd gnd cell_6t
Xbit_r24_c2 bl[2] br[2] wl[24] vdd gnd cell_6t
Xbit_r25_c2 bl[2] br[2] wl[25] vdd gnd cell_6t
Xbit_r26_c2 bl[2] br[2] wl[26] vdd gnd cell_6t
Xbit_r27_c2 bl[2] br[2] wl[27] vdd gnd cell_6t
Xbit_r28_c2 bl[2] br[2] wl[28] vdd gnd cell_6t
Xbit_r29_c2 bl[2] br[2] wl[29] vdd gnd cell_6t
Xbit_r30_c2 bl[2] br[2] wl[30] vdd gnd cell_6t
Xbit_r31_c2 bl[2] br[2] wl[31] vdd gnd cell_6t
Xbit_r32_c2 bl[2] br[2] wl[32] vdd gnd cell_6t
Xbit_r33_c2 bl[2] br[2] wl[33] vdd gnd cell_6t
Xbit_r34_c2 bl[2] br[2] wl[34] vdd gnd cell_6t
Xbit_r35_c2 bl[2] br[2] wl[35] vdd gnd cell_6t
Xbit_r36_c2 bl[2] br[2] wl[36] vdd gnd cell_6t
Xbit_r37_c2 bl[2] br[2] wl[37] vdd gnd cell_6t
Xbit_r38_c2 bl[2] br[2] wl[38] vdd gnd cell_6t
Xbit_r39_c2 bl[2] br[2] wl[39] vdd gnd cell_6t
Xbit_r40_c2 bl[2] br[2] wl[40] vdd gnd cell_6t
Xbit_r41_c2 bl[2] br[2] wl[41] vdd gnd cell_6t
Xbit_r42_c2 bl[2] br[2] wl[42] vdd gnd cell_6t
Xbit_r43_c2 bl[2] br[2] wl[43] vdd gnd cell_6t
Xbit_r44_c2 bl[2] br[2] wl[44] vdd gnd cell_6t
Xbit_r45_c2 bl[2] br[2] wl[45] vdd gnd cell_6t
Xbit_r46_c2 bl[2] br[2] wl[46] vdd gnd cell_6t
Xbit_r47_c2 bl[2] br[2] wl[47] vdd gnd cell_6t
Xbit_r48_c2 bl[2] br[2] wl[48] vdd gnd cell_6t
Xbit_r49_c2 bl[2] br[2] wl[49] vdd gnd cell_6t
Xbit_r50_c2 bl[2] br[2] wl[50] vdd gnd cell_6t
Xbit_r51_c2 bl[2] br[2] wl[51] vdd gnd cell_6t
Xbit_r52_c2 bl[2] br[2] wl[52] vdd gnd cell_6t
Xbit_r53_c2 bl[2] br[2] wl[53] vdd gnd cell_6t
Xbit_r54_c2 bl[2] br[2] wl[54] vdd gnd cell_6t
Xbit_r55_c2 bl[2] br[2] wl[55] vdd gnd cell_6t
Xbit_r56_c2 bl[2] br[2] wl[56] vdd gnd cell_6t
Xbit_r57_c2 bl[2] br[2] wl[57] vdd gnd cell_6t
Xbit_r58_c2 bl[2] br[2] wl[58] vdd gnd cell_6t
Xbit_r59_c2 bl[2] br[2] wl[59] vdd gnd cell_6t
Xbit_r60_c2 bl[2] br[2] wl[60] vdd gnd cell_6t
Xbit_r61_c2 bl[2] br[2] wl[61] vdd gnd cell_6t
Xbit_r62_c2 bl[2] br[2] wl[62] vdd gnd cell_6t
Xbit_r63_c2 bl[2] br[2] wl[63] vdd gnd cell_6t
Xbit_r64_c2 bl[2] br[2] wl[64] vdd gnd cell_6t
Xbit_r65_c2 bl[2] br[2] wl[65] vdd gnd cell_6t
Xbit_r66_c2 bl[2] br[2] wl[66] vdd gnd cell_6t
Xbit_r67_c2 bl[2] br[2] wl[67] vdd gnd cell_6t
Xbit_r68_c2 bl[2] br[2] wl[68] vdd gnd cell_6t
Xbit_r69_c2 bl[2] br[2] wl[69] vdd gnd cell_6t
Xbit_r70_c2 bl[2] br[2] wl[70] vdd gnd cell_6t
Xbit_r71_c2 bl[2] br[2] wl[71] vdd gnd cell_6t
Xbit_r72_c2 bl[2] br[2] wl[72] vdd gnd cell_6t
Xbit_r73_c2 bl[2] br[2] wl[73] vdd gnd cell_6t
Xbit_r74_c2 bl[2] br[2] wl[74] vdd gnd cell_6t
Xbit_r75_c2 bl[2] br[2] wl[75] vdd gnd cell_6t
Xbit_r76_c2 bl[2] br[2] wl[76] vdd gnd cell_6t
Xbit_r77_c2 bl[2] br[2] wl[77] vdd gnd cell_6t
Xbit_r78_c2 bl[2] br[2] wl[78] vdd gnd cell_6t
Xbit_r79_c2 bl[2] br[2] wl[79] vdd gnd cell_6t
Xbit_r80_c2 bl[2] br[2] wl[80] vdd gnd cell_6t
Xbit_r81_c2 bl[2] br[2] wl[81] vdd gnd cell_6t
Xbit_r82_c2 bl[2] br[2] wl[82] vdd gnd cell_6t
Xbit_r83_c2 bl[2] br[2] wl[83] vdd gnd cell_6t
Xbit_r84_c2 bl[2] br[2] wl[84] vdd gnd cell_6t
Xbit_r85_c2 bl[2] br[2] wl[85] vdd gnd cell_6t
Xbit_r86_c2 bl[2] br[2] wl[86] vdd gnd cell_6t
Xbit_r87_c2 bl[2] br[2] wl[87] vdd gnd cell_6t
Xbit_r88_c2 bl[2] br[2] wl[88] vdd gnd cell_6t
Xbit_r89_c2 bl[2] br[2] wl[89] vdd gnd cell_6t
Xbit_r90_c2 bl[2] br[2] wl[90] vdd gnd cell_6t
Xbit_r91_c2 bl[2] br[2] wl[91] vdd gnd cell_6t
Xbit_r92_c2 bl[2] br[2] wl[92] vdd gnd cell_6t
Xbit_r93_c2 bl[2] br[2] wl[93] vdd gnd cell_6t
Xbit_r94_c2 bl[2] br[2] wl[94] vdd gnd cell_6t
Xbit_r95_c2 bl[2] br[2] wl[95] vdd gnd cell_6t
Xbit_r96_c2 bl[2] br[2] wl[96] vdd gnd cell_6t
Xbit_r97_c2 bl[2] br[2] wl[97] vdd gnd cell_6t
Xbit_r98_c2 bl[2] br[2] wl[98] vdd gnd cell_6t
Xbit_r99_c2 bl[2] br[2] wl[99] vdd gnd cell_6t
Xbit_r100_c2 bl[2] br[2] wl[100] vdd gnd cell_6t
Xbit_r101_c2 bl[2] br[2] wl[101] vdd gnd cell_6t
Xbit_r102_c2 bl[2] br[2] wl[102] vdd gnd cell_6t
Xbit_r103_c2 bl[2] br[2] wl[103] vdd gnd cell_6t
Xbit_r104_c2 bl[2] br[2] wl[104] vdd gnd cell_6t
Xbit_r105_c2 bl[2] br[2] wl[105] vdd gnd cell_6t
Xbit_r106_c2 bl[2] br[2] wl[106] vdd gnd cell_6t
Xbit_r107_c2 bl[2] br[2] wl[107] vdd gnd cell_6t
Xbit_r108_c2 bl[2] br[2] wl[108] vdd gnd cell_6t
Xbit_r109_c2 bl[2] br[2] wl[109] vdd gnd cell_6t
Xbit_r110_c2 bl[2] br[2] wl[110] vdd gnd cell_6t
Xbit_r111_c2 bl[2] br[2] wl[111] vdd gnd cell_6t
Xbit_r112_c2 bl[2] br[2] wl[112] vdd gnd cell_6t
Xbit_r113_c2 bl[2] br[2] wl[113] vdd gnd cell_6t
Xbit_r114_c2 bl[2] br[2] wl[114] vdd gnd cell_6t
Xbit_r115_c2 bl[2] br[2] wl[115] vdd gnd cell_6t
Xbit_r116_c2 bl[2] br[2] wl[116] vdd gnd cell_6t
Xbit_r117_c2 bl[2] br[2] wl[117] vdd gnd cell_6t
Xbit_r118_c2 bl[2] br[2] wl[118] vdd gnd cell_6t
Xbit_r119_c2 bl[2] br[2] wl[119] vdd gnd cell_6t
Xbit_r120_c2 bl[2] br[2] wl[120] vdd gnd cell_6t
Xbit_r121_c2 bl[2] br[2] wl[121] vdd gnd cell_6t
Xbit_r122_c2 bl[2] br[2] wl[122] vdd gnd cell_6t
Xbit_r123_c2 bl[2] br[2] wl[123] vdd gnd cell_6t
Xbit_r124_c2 bl[2] br[2] wl[124] vdd gnd cell_6t
Xbit_r125_c2 bl[2] br[2] wl[125] vdd gnd cell_6t
Xbit_r126_c2 bl[2] br[2] wl[126] vdd gnd cell_6t
Xbit_r127_c2 bl[2] br[2] wl[127] vdd gnd cell_6t
Xbit_r128_c2 bl[2] br[2] wl[128] vdd gnd cell_6t
Xbit_r129_c2 bl[2] br[2] wl[129] vdd gnd cell_6t
Xbit_r130_c2 bl[2] br[2] wl[130] vdd gnd cell_6t
Xbit_r131_c2 bl[2] br[2] wl[131] vdd gnd cell_6t
Xbit_r132_c2 bl[2] br[2] wl[132] vdd gnd cell_6t
Xbit_r133_c2 bl[2] br[2] wl[133] vdd gnd cell_6t
Xbit_r134_c2 bl[2] br[2] wl[134] vdd gnd cell_6t
Xbit_r135_c2 bl[2] br[2] wl[135] vdd gnd cell_6t
Xbit_r136_c2 bl[2] br[2] wl[136] vdd gnd cell_6t
Xbit_r137_c2 bl[2] br[2] wl[137] vdd gnd cell_6t
Xbit_r138_c2 bl[2] br[2] wl[138] vdd gnd cell_6t
Xbit_r139_c2 bl[2] br[2] wl[139] vdd gnd cell_6t
Xbit_r140_c2 bl[2] br[2] wl[140] vdd gnd cell_6t
Xbit_r141_c2 bl[2] br[2] wl[141] vdd gnd cell_6t
Xbit_r142_c2 bl[2] br[2] wl[142] vdd gnd cell_6t
Xbit_r143_c2 bl[2] br[2] wl[143] vdd gnd cell_6t
Xbit_r144_c2 bl[2] br[2] wl[144] vdd gnd cell_6t
Xbit_r145_c2 bl[2] br[2] wl[145] vdd gnd cell_6t
Xbit_r146_c2 bl[2] br[2] wl[146] vdd gnd cell_6t
Xbit_r147_c2 bl[2] br[2] wl[147] vdd gnd cell_6t
Xbit_r148_c2 bl[2] br[2] wl[148] vdd gnd cell_6t
Xbit_r149_c2 bl[2] br[2] wl[149] vdd gnd cell_6t
Xbit_r150_c2 bl[2] br[2] wl[150] vdd gnd cell_6t
Xbit_r151_c2 bl[2] br[2] wl[151] vdd gnd cell_6t
Xbit_r152_c2 bl[2] br[2] wl[152] vdd gnd cell_6t
Xbit_r153_c2 bl[2] br[2] wl[153] vdd gnd cell_6t
Xbit_r154_c2 bl[2] br[2] wl[154] vdd gnd cell_6t
Xbit_r155_c2 bl[2] br[2] wl[155] vdd gnd cell_6t
Xbit_r156_c2 bl[2] br[2] wl[156] vdd gnd cell_6t
Xbit_r157_c2 bl[2] br[2] wl[157] vdd gnd cell_6t
Xbit_r158_c2 bl[2] br[2] wl[158] vdd gnd cell_6t
Xbit_r159_c2 bl[2] br[2] wl[159] vdd gnd cell_6t
Xbit_r160_c2 bl[2] br[2] wl[160] vdd gnd cell_6t
Xbit_r161_c2 bl[2] br[2] wl[161] vdd gnd cell_6t
Xbit_r162_c2 bl[2] br[2] wl[162] vdd gnd cell_6t
Xbit_r163_c2 bl[2] br[2] wl[163] vdd gnd cell_6t
Xbit_r164_c2 bl[2] br[2] wl[164] vdd gnd cell_6t
Xbit_r165_c2 bl[2] br[2] wl[165] vdd gnd cell_6t
Xbit_r166_c2 bl[2] br[2] wl[166] vdd gnd cell_6t
Xbit_r167_c2 bl[2] br[2] wl[167] vdd gnd cell_6t
Xbit_r168_c2 bl[2] br[2] wl[168] vdd gnd cell_6t
Xbit_r169_c2 bl[2] br[2] wl[169] vdd gnd cell_6t
Xbit_r170_c2 bl[2] br[2] wl[170] vdd gnd cell_6t
Xbit_r171_c2 bl[2] br[2] wl[171] vdd gnd cell_6t
Xbit_r172_c2 bl[2] br[2] wl[172] vdd gnd cell_6t
Xbit_r173_c2 bl[2] br[2] wl[173] vdd gnd cell_6t
Xbit_r174_c2 bl[2] br[2] wl[174] vdd gnd cell_6t
Xbit_r175_c2 bl[2] br[2] wl[175] vdd gnd cell_6t
Xbit_r176_c2 bl[2] br[2] wl[176] vdd gnd cell_6t
Xbit_r177_c2 bl[2] br[2] wl[177] vdd gnd cell_6t
Xbit_r178_c2 bl[2] br[2] wl[178] vdd gnd cell_6t
Xbit_r179_c2 bl[2] br[2] wl[179] vdd gnd cell_6t
Xbit_r180_c2 bl[2] br[2] wl[180] vdd gnd cell_6t
Xbit_r181_c2 bl[2] br[2] wl[181] vdd gnd cell_6t
Xbit_r182_c2 bl[2] br[2] wl[182] vdd gnd cell_6t
Xbit_r183_c2 bl[2] br[2] wl[183] vdd gnd cell_6t
Xbit_r184_c2 bl[2] br[2] wl[184] vdd gnd cell_6t
Xbit_r185_c2 bl[2] br[2] wl[185] vdd gnd cell_6t
Xbit_r186_c2 bl[2] br[2] wl[186] vdd gnd cell_6t
Xbit_r187_c2 bl[2] br[2] wl[187] vdd gnd cell_6t
Xbit_r188_c2 bl[2] br[2] wl[188] vdd gnd cell_6t
Xbit_r189_c2 bl[2] br[2] wl[189] vdd gnd cell_6t
Xbit_r190_c2 bl[2] br[2] wl[190] vdd gnd cell_6t
Xbit_r191_c2 bl[2] br[2] wl[191] vdd gnd cell_6t
Xbit_r192_c2 bl[2] br[2] wl[192] vdd gnd cell_6t
Xbit_r193_c2 bl[2] br[2] wl[193] vdd gnd cell_6t
Xbit_r194_c2 bl[2] br[2] wl[194] vdd gnd cell_6t
Xbit_r195_c2 bl[2] br[2] wl[195] vdd gnd cell_6t
Xbit_r196_c2 bl[2] br[2] wl[196] vdd gnd cell_6t
Xbit_r197_c2 bl[2] br[2] wl[197] vdd gnd cell_6t
Xbit_r198_c2 bl[2] br[2] wl[198] vdd gnd cell_6t
Xbit_r199_c2 bl[2] br[2] wl[199] vdd gnd cell_6t
Xbit_r200_c2 bl[2] br[2] wl[200] vdd gnd cell_6t
Xbit_r201_c2 bl[2] br[2] wl[201] vdd gnd cell_6t
Xbit_r202_c2 bl[2] br[2] wl[202] vdd gnd cell_6t
Xbit_r203_c2 bl[2] br[2] wl[203] vdd gnd cell_6t
Xbit_r204_c2 bl[2] br[2] wl[204] vdd gnd cell_6t
Xbit_r205_c2 bl[2] br[2] wl[205] vdd gnd cell_6t
Xbit_r206_c2 bl[2] br[2] wl[206] vdd gnd cell_6t
Xbit_r207_c2 bl[2] br[2] wl[207] vdd gnd cell_6t
Xbit_r208_c2 bl[2] br[2] wl[208] vdd gnd cell_6t
Xbit_r209_c2 bl[2] br[2] wl[209] vdd gnd cell_6t
Xbit_r210_c2 bl[2] br[2] wl[210] vdd gnd cell_6t
Xbit_r211_c2 bl[2] br[2] wl[211] vdd gnd cell_6t
Xbit_r212_c2 bl[2] br[2] wl[212] vdd gnd cell_6t
Xbit_r213_c2 bl[2] br[2] wl[213] vdd gnd cell_6t
Xbit_r214_c2 bl[2] br[2] wl[214] vdd gnd cell_6t
Xbit_r215_c2 bl[2] br[2] wl[215] vdd gnd cell_6t
Xbit_r216_c2 bl[2] br[2] wl[216] vdd gnd cell_6t
Xbit_r217_c2 bl[2] br[2] wl[217] vdd gnd cell_6t
Xbit_r218_c2 bl[2] br[2] wl[218] vdd gnd cell_6t
Xbit_r219_c2 bl[2] br[2] wl[219] vdd gnd cell_6t
Xbit_r220_c2 bl[2] br[2] wl[220] vdd gnd cell_6t
Xbit_r221_c2 bl[2] br[2] wl[221] vdd gnd cell_6t
Xbit_r222_c2 bl[2] br[2] wl[222] vdd gnd cell_6t
Xbit_r223_c2 bl[2] br[2] wl[223] vdd gnd cell_6t
Xbit_r224_c2 bl[2] br[2] wl[224] vdd gnd cell_6t
Xbit_r225_c2 bl[2] br[2] wl[225] vdd gnd cell_6t
Xbit_r226_c2 bl[2] br[2] wl[226] vdd gnd cell_6t
Xbit_r227_c2 bl[2] br[2] wl[227] vdd gnd cell_6t
Xbit_r228_c2 bl[2] br[2] wl[228] vdd gnd cell_6t
Xbit_r229_c2 bl[2] br[2] wl[229] vdd gnd cell_6t
Xbit_r230_c2 bl[2] br[2] wl[230] vdd gnd cell_6t
Xbit_r231_c2 bl[2] br[2] wl[231] vdd gnd cell_6t
Xbit_r232_c2 bl[2] br[2] wl[232] vdd gnd cell_6t
Xbit_r233_c2 bl[2] br[2] wl[233] vdd gnd cell_6t
Xbit_r234_c2 bl[2] br[2] wl[234] vdd gnd cell_6t
Xbit_r235_c2 bl[2] br[2] wl[235] vdd gnd cell_6t
Xbit_r236_c2 bl[2] br[2] wl[236] vdd gnd cell_6t
Xbit_r237_c2 bl[2] br[2] wl[237] vdd gnd cell_6t
Xbit_r238_c2 bl[2] br[2] wl[238] vdd gnd cell_6t
Xbit_r239_c2 bl[2] br[2] wl[239] vdd gnd cell_6t
Xbit_r240_c2 bl[2] br[2] wl[240] vdd gnd cell_6t
Xbit_r241_c2 bl[2] br[2] wl[241] vdd gnd cell_6t
Xbit_r242_c2 bl[2] br[2] wl[242] vdd gnd cell_6t
Xbit_r243_c2 bl[2] br[2] wl[243] vdd gnd cell_6t
Xbit_r244_c2 bl[2] br[2] wl[244] vdd gnd cell_6t
Xbit_r245_c2 bl[2] br[2] wl[245] vdd gnd cell_6t
Xbit_r246_c2 bl[2] br[2] wl[246] vdd gnd cell_6t
Xbit_r247_c2 bl[2] br[2] wl[247] vdd gnd cell_6t
Xbit_r248_c2 bl[2] br[2] wl[248] vdd gnd cell_6t
Xbit_r249_c2 bl[2] br[2] wl[249] vdd gnd cell_6t
Xbit_r250_c2 bl[2] br[2] wl[250] vdd gnd cell_6t
Xbit_r251_c2 bl[2] br[2] wl[251] vdd gnd cell_6t
Xbit_r252_c2 bl[2] br[2] wl[252] vdd gnd cell_6t
Xbit_r253_c2 bl[2] br[2] wl[253] vdd gnd cell_6t
Xbit_r254_c2 bl[2] br[2] wl[254] vdd gnd cell_6t
Xbit_r255_c2 bl[2] br[2] wl[255] vdd gnd cell_6t
Xbit_r256_c2 bl[2] br[2] wl[256] vdd gnd cell_6t
Xbit_r257_c2 bl[2] br[2] wl[257] vdd gnd cell_6t
Xbit_r258_c2 bl[2] br[2] wl[258] vdd gnd cell_6t
Xbit_r259_c2 bl[2] br[2] wl[259] vdd gnd cell_6t
Xbit_r260_c2 bl[2] br[2] wl[260] vdd gnd cell_6t
Xbit_r261_c2 bl[2] br[2] wl[261] vdd gnd cell_6t
Xbit_r262_c2 bl[2] br[2] wl[262] vdd gnd cell_6t
Xbit_r263_c2 bl[2] br[2] wl[263] vdd gnd cell_6t
Xbit_r264_c2 bl[2] br[2] wl[264] vdd gnd cell_6t
Xbit_r265_c2 bl[2] br[2] wl[265] vdd gnd cell_6t
Xbit_r266_c2 bl[2] br[2] wl[266] vdd gnd cell_6t
Xbit_r267_c2 bl[2] br[2] wl[267] vdd gnd cell_6t
Xbit_r268_c2 bl[2] br[2] wl[268] vdd gnd cell_6t
Xbit_r269_c2 bl[2] br[2] wl[269] vdd gnd cell_6t
Xbit_r270_c2 bl[2] br[2] wl[270] vdd gnd cell_6t
Xbit_r271_c2 bl[2] br[2] wl[271] vdd gnd cell_6t
Xbit_r272_c2 bl[2] br[2] wl[272] vdd gnd cell_6t
Xbit_r273_c2 bl[2] br[2] wl[273] vdd gnd cell_6t
Xbit_r274_c2 bl[2] br[2] wl[274] vdd gnd cell_6t
Xbit_r275_c2 bl[2] br[2] wl[275] vdd gnd cell_6t
Xbit_r276_c2 bl[2] br[2] wl[276] vdd gnd cell_6t
Xbit_r277_c2 bl[2] br[2] wl[277] vdd gnd cell_6t
Xbit_r278_c2 bl[2] br[2] wl[278] vdd gnd cell_6t
Xbit_r279_c2 bl[2] br[2] wl[279] vdd gnd cell_6t
Xbit_r280_c2 bl[2] br[2] wl[280] vdd gnd cell_6t
Xbit_r281_c2 bl[2] br[2] wl[281] vdd gnd cell_6t
Xbit_r282_c2 bl[2] br[2] wl[282] vdd gnd cell_6t
Xbit_r283_c2 bl[2] br[2] wl[283] vdd gnd cell_6t
Xbit_r284_c2 bl[2] br[2] wl[284] vdd gnd cell_6t
Xbit_r285_c2 bl[2] br[2] wl[285] vdd gnd cell_6t
Xbit_r286_c2 bl[2] br[2] wl[286] vdd gnd cell_6t
Xbit_r287_c2 bl[2] br[2] wl[287] vdd gnd cell_6t
Xbit_r288_c2 bl[2] br[2] wl[288] vdd gnd cell_6t
Xbit_r289_c2 bl[2] br[2] wl[289] vdd gnd cell_6t
Xbit_r290_c2 bl[2] br[2] wl[290] vdd gnd cell_6t
Xbit_r291_c2 bl[2] br[2] wl[291] vdd gnd cell_6t
Xbit_r292_c2 bl[2] br[2] wl[292] vdd gnd cell_6t
Xbit_r293_c2 bl[2] br[2] wl[293] vdd gnd cell_6t
Xbit_r294_c2 bl[2] br[2] wl[294] vdd gnd cell_6t
Xbit_r295_c2 bl[2] br[2] wl[295] vdd gnd cell_6t
Xbit_r296_c2 bl[2] br[2] wl[296] vdd gnd cell_6t
Xbit_r297_c2 bl[2] br[2] wl[297] vdd gnd cell_6t
Xbit_r298_c2 bl[2] br[2] wl[298] vdd gnd cell_6t
Xbit_r299_c2 bl[2] br[2] wl[299] vdd gnd cell_6t
Xbit_r300_c2 bl[2] br[2] wl[300] vdd gnd cell_6t
Xbit_r301_c2 bl[2] br[2] wl[301] vdd gnd cell_6t
Xbit_r302_c2 bl[2] br[2] wl[302] vdd gnd cell_6t
Xbit_r303_c2 bl[2] br[2] wl[303] vdd gnd cell_6t
Xbit_r304_c2 bl[2] br[2] wl[304] vdd gnd cell_6t
Xbit_r305_c2 bl[2] br[2] wl[305] vdd gnd cell_6t
Xbit_r306_c2 bl[2] br[2] wl[306] vdd gnd cell_6t
Xbit_r307_c2 bl[2] br[2] wl[307] vdd gnd cell_6t
Xbit_r308_c2 bl[2] br[2] wl[308] vdd gnd cell_6t
Xbit_r309_c2 bl[2] br[2] wl[309] vdd gnd cell_6t
Xbit_r310_c2 bl[2] br[2] wl[310] vdd gnd cell_6t
Xbit_r311_c2 bl[2] br[2] wl[311] vdd gnd cell_6t
Xbit_r312_c2 bl[2] br[2] wl[312] vdd gnd cell_6t
Xbit_r313_c2 bl[2] br[2] wl[313] vdd gnd cell_6t
Xbit_r314_c2 bl[2] br[2] wl[314] vdd gnd cell_6t
Xbit_r315_c2 bl[2] br[2] wl[315] vdd gnd cell_6t
Xbit_r316_c2 bl[2] br[2] wl[316] vdd gnd cell_6t
Xbit_r317_c2 bl[2] br[2] wl[317] vdd gnd cell_6t
Xbit_r318_c2 bl[2] br[2] wl[318] vdd gnd cell_6t
Xbit_r319_c2 bl[2] br[2] wl[319] vdd gnd cell_6t
Xbit_r320_c2 bl[2] br[2] wl[320] vdd gnd cell_6t
Xbit_r321_c2 bl[2] br[2] wl[321] vdd gnd cell_6t
Xbit_r322_c2 bl[2] br[2] wl[322] vdd gnd cell_6t
Xbit_r323_c2 bl[2] br[2] wl[323] vdd gnd cell_6t
Xbit_r324_c2 bl[2] br[2] wl[324] vdd gnd cell_6t
Xbit_r325_c2 bl[2] br[2] wl[325] vdd gnd cell_6t
Xbit_r326_c2 bl[2] br[2] wl[326] vdd gnd cell_6t
Xbit_r327_c2 bl[2] br[2] wl[327] vdd gnd cell_6t
Xbit_r328_c2 bl[2] br[2] wl[328] vdd gnd cell_6t
Xbit_r329_c2 bl[2] br[2] wl[329] vdd gnd cell_6t
Xbit_r330_c2 bl[2] br[2] wl[330] vdd gnd cell_6t
Xbit_r331_c2 bl[2] br[2] wl[331] vdd gnd cell_6t
Xbit_r332_c2 bl[2] br[2] wl[332] vdd gnd cell_6t
Xbit_r333_c2 bl[2] br[2] wl[333] vdd gnd cell_6t
Xbit_r334_c2 bl[2] br[2] wl[334] vdd gnd cell_6t
Xbit_r335_c2 bl[2] br[2] wl[335] vdd gnd cell_6t
Xbit_r336_c2 bl[2] br[2] wl[336] vdd gnd cell_6t
Xbit_r337_c2 bl[2] br[2] wl[337] vdd gnd cell_6t
Xbit_r338_c2 bl[2] br[2] wl[338] vdd gnd cell_6t
Xbit_r339_c2 bl[2] br[2] wl[339] vdd gnd cell_6t
Xbit_r340_c2 bl[2] br[2] wl[340] vdd gnd cell_6t
Xbit_r341_c2 bl[2] br[2] wl[341] vdd gnd cell_6t
Xbit_r342_c2 bl[2] br[2] wl[342] vdd gnd cell_6t
Xbit_r343_c2 bl[2] br[2] wl[343] vdd gnd cell_6t
Xbit_r344_c2 bl[2] br[2] wl[344] vdd gnd cell_6t
Xbit_r345_c2 bl[2] br[2] wl[345] vdd gnd cell_6t
Xbit_r346_c2 bl[2] br[2] wl[346] vdd gnd cell_6t
Xbit_r347_c2 bl[2] br[2] wl[347] vdd gnd cell_6t
Xbit_r348_c2 bl[2] br[2] wl[348] vdd gnd cell_6t
Xbit_r349_c2 bl[2] br[2] wl[349] vdd gnd cell_6t
Xbit_r350_c2 bl[2] br[2] wl[350] vdd gnd cell_6t
Xbit_r351_c2 bl[2] br[2] wl[351] vdd gnd cell_6t
Xbit_r352_c2 bl[2] br[2] wl[352] vdd gnd cell_6t
Xbit_r353_c2 bl[2] br[2] wl[353] vdd gnd cell_6t
Xbit_r354_c2 bl[2] br[2] wl[354] vdd gnd cell_6t
Xbit_r355_c2 bl[2] br[2] wl[355] vdd gnd cell_6t
Xbit_r356_c2 bl[2] br[2] wl[356] vdd gnd cell_6t
Xbit_r357_c2 bl[2] br[2] wl[357] vdd gnd cell_6t
Xbit_r358_c2 bl[2] br[2] wl[358] vdd gnd cell_6t
Xbit_r359_c2 bl[2] br[2] wl[359] vdd gnd cell_6t
Xbit_r360_c2 bl[2] br[2] wl[360] vdd gnd cell_6t
Xbit_r361_c2 bl[2] br[2] wl[361] vdd gnd cell_6t
Xbit_r362_c2 bl[2] br[2] wl[362] vdd gnd cell_6t
Xbit_r363_c2 bl[2] br[2] wl[363] vdd gnd cell_6t
Xbit_r364_c2 bl[2] br[2] wl[364] vdd gnd cell_6t
Xbit_r365_c2 bl[2] br[2] wl[365] vdd gnd cell_6t
Xbit_r366_c2 bl[2] br[2] wl[366] vdd gnd cell_6t
Xbit_r367_c2 bl[2] br[2] wl[367] vdd gnd cell_6t
Xbit_r368_c2 bl[2] br[2] wl[368] vdd gnd cell_6t
Xbit_r369_c2 bl[2] br[2] wl[369] vdd gnd cell_6t
Xbit_r370_c2 bl[2] br[2] wl[370] vdd gnd cell_6t
Xbit_r371_c2 bl[2] br[2] wl[371] vdd gnd cell_6t
Xbit_r372_c2 bl[2] br[2] wl[372] vdd gnd cell_6t
Xbit_r373_c2 bl[2] br[2] wl[373] vdd gnd cell_6t
Xbit_r374_c2 bl[2] br[2] wl[374] vdd gnd cell_6t
Xbit_r375_c2 bl[2] br[2] wl[375] vdd gnd cell_6t
Xbit_r376_c2 bl[2] br[2] wl[376] vdd gnd cell_6t
Xbit_r377_c2 bl[2] br[2] wl[377] vdd gnd cell_6t
Xbit_r378_c2 bl[2] br[2] wl[378] vdd gnd cell_6t
Xbit_r379_c2 bl[2] br[2] wl[379] vdd gnd cell_6t
Xbit_r380_c2 bl[2] br[2] wl[380] vdd gnd cell_6t
Xbit_r381_c2 bl[2] br[2] wl[381] vdd gnd cell_6t
Xbit_r382_c2 bl[2] br[2] wl[382] vdd gnd cell_6t
Xbit_r383_c2 bl[2] br[2] wl[383] vdd gnd cell_6t
Xbit_r384_c2 bl[2] br[2] wl[384] vdd gnd cell_6t
Xbit_r385_c2 bl[2] br[2] wl[385] vdd gnd cell_6t
Xbit_r386_c2 bl[2] br[2] wl[386] vdd gnd cell_6t
Xbit_r387_c2 bl[2] br[2] wl[387] vdd gnd cell_6t
Xbit_r388_c2 bl[2] br[2] wl[388] vdd gnd cell_6t
Xbit_r389_c2 bl[2] br[2] wl[389] vdd gnd cell_6t
Xbit_r390_c2 bl[2] br[2] wl[390] vdd gnd cell_6t
Xbit_r391_c2 bl[2] br[2] wl[391] vdd gnd cell_6t
Xbit_r392_c2 bl[2] br[2] wl[392] vdd gnd cell_6t
Xbit_r393_c2 bl[2] br[2] wl[393] vdd gnd cell_6t
Xbit_r394_c2 bl[2] br[2] wl[394] vdd gnd cell_6t
Xbit_r395_c2 bl[2] br[2] wl[395] vdd gnd cell_6t
Xbit_r396_c2 bl[2] br[2] wl[396] vdd gnd cell_6t
Xbit_r397_c2 bl[2] br[2] wl[397] vdd gnd cell_6t
Xbit_r398_c2 bl[2] br[2] wl[398] vdd gnd cell_6t
Xbit_r399_c2 bl[2] br[2] wl[399] vdd gnd cell_6t
Xbit_r400_c2 bl[2] br[2] wl[400] vdd gnd cell_6t
Xbit_r401_c2 bl[2] br[2] wl[401] vdd gnd cell_6t
Xbit_r402_c2 bl[2] br[2] wl[402] vdd gnd cell_6t
Xbit_r403_c2 bl[2] br[2] wl[403] vdd gnd cell_6t
Xbit_r404_c2 bl[2] br[2] wl[404] vdd gnd cell_6t
Xbit_r405_c2 bl[2] br[2] wl[405] vdd gnd cell_6t
Xbit_r406_c2 bl[2] br[2] wl[406] vdd gnd cell_6t
Xbit_r407_c2 bl[2] br[2] wl[407] vdd gnd cell_6t
Xbit_r408_c2 bl[2] br[2] wl[408] vdd gnd cell_6t
Xbit_r409_c2 bl[2] br[2] wl[409] vdd gnd cell_6t
Xbit_r410_c2 bl[2] br[2] wl[410] vdd gnd cell_6t
Xbit_r411_c2 bl[2] br[2] wl[411] vdd gnd cell_6t
Xbit_r412_c2 bl[2] br[2] wl[412] vdd gnd cell_6t
Xbit_r413_c2 bl[2] br[2] wl[413] vdd gnd cell_6t
Xbit_r414_c2 bl[2] br[2] wl[414] vdd gnd cell_6t
Xbit_r415_c2 bl[2] br[2] wl[415] vdd gnd cell_6t
Xbit_r416_c2 bl[2] br[2] wl[416] vdd gnd cell_6t
Xbit_r417_c2 bl[2] br[2] wl[417] vdd gnd cell_6t
Xbit_r418_c2 bl[2] br[2] wl[418] vdd gnd cell_6t
Xbit_r419_c2 bl[2] br[2] wl[419] vdd gnd cell_6t
Xbit_r420_c2 bl[2] br[2] wl[420] vdd gnd cell_6t
Xbit_r421_c2 bl[2] br[2] wl[421] vdd gnd cell_6t
Xbit_r422_c2 bl[2] br[2] wl[422] vdd gnd cell_6t
Xbit_r423_c2 bl[2] br[2] wl[423] vdd gnd cell_6t
Xbit_r424_c2 bl[2] br[2] wl[424] vdd gnd cell_6t
Xbit_r425_c2 bl[2] br[2] wl[425] vdd gnd cell_6t
Xbit_r426_c2 bl[2] br[2] wl[426] vdd gnd cell_6t
Xbit_r427_c2 bl[2] br[2] wl[427] vdd gnd cell_6t
Xbit_r428_c2 bl[2] br[2] wl[428] vdd gnd cell_6t
Xbit_r429_c2 bl[2] br[2] wl[429] vdd gnd cell_6t
Xbit_r430_c2 bl[2] br[2] wl[430] vdd gnd cell_6t
Xbit_r431_c2 bl[2] br[2] wl[431] vdd gnd cell_6t
Xbit_r432_c2 bl[2] br[2] wl[432] vdd gnd cell_6t
Xbit_r433_c2 bl[2] br[2] wl[433] vdd gnd cell_6t
Xbit_r434_c2 bl[2] br[2] wl[434] vdd gnd cell_6t
Xbit_r435_c2 bl[2] br[2] wl[435] vdd gnd cell_6t
Xbit_r436_c2 bl[2] br[2] wl[436] vdd gnd cell_6t
Xbit_r437_c2 bl[2] br[2] wl[437] vdd gnd cell_6t
Xbit_r438_c2 bl[2] br[2] wl[438] vdd gnd cell_6t
Xbit_r439_c2 bl[2] br[2] wl[439] vdd gnd cell_6t
Xbit_r440_c2 bl[2] br[2] wl[440] vdd gnd cell_6t
Xbit_r441_c2 bl[2] br[2] wl[441] vdd gnd cell_6t
Xbit_r442_c2 bl[2] br[2] wl[442] vdd gnd cell_6t
Xbit_r443_c2 bl[2] br[2] wl[443] vdd gnd cell_6t
Xbit_r444_c2 bl[2] br[2] wl[444] vdd gnd cell_6t
Xbit_r445_c2 bl[2] br[2] wl[445] vdd gnd cell_6t
Xbit_r446_c2 bl[2] br[2] wl[446] vdd gnd cell_6t
Xbit_r447_c2 bl[2] br[2] wl[447] vdd gnd cell_6t
Xbit_r448_c2 bl[2] br[2] wl[448] vdd gnd cell_6t
Xbit_r449_c2 bl[2] br[2] wl[449] vdd gnd cell_6t
Xbit_r450_c2 bl[2] br[2] wl[450] vdd gnd cell_6t
Xbit_r451_c2 bl[2] br[2] wl[451] vdd gnd cell_6t
Xbit_r452_c2 bl[2] br[2] wl[452] vdd gnd cell_6t
Xbit_r453_c2 bl[2] br[2] wl[453] vdd gnd cell_6t
Xbit_r454_c2 bl[2] br[2] wl[454] vdd gnd cell_6t
Xbit_r455_c2 bl[2] br[2] wl[455] vdd gnd cell_6t
Xbit_r456_c2 bl[2] br[2] wl[456] vdd gnd cell_6t
Xbit_r457_c2 bl[2] br[2] wl[457] vdd gnd cell_6t
Xbit_r458_c2 bl[2] br[2] wl[458] vdd gnd cell_6t
Xbit_r459_c2 bl[2] br[2] wl[459] vdd gnd cell_6t
Xbit_r460_c2 bl[2] br[2] wl[460] vdd gnd cell_6t
Xbit_r461_c2 bl[2] br[2] wl[461] vdd gnd cell_6t
Xbit_r462_c2 bl[2] br[2] wl[462] vdd gnd cell_6t
Xbit_r463_c2 bl[2] br[2] wl[463] vdd gnd cell_6t
Xbit_r464_c2 bl[2] br[2] wl[464] vdd gnd cell_6t
Xbit_r465_c2 bl[2] br[2] wl[465] vdd gnd cell_6t
Xbit_r466_c2 bl[2] br[2] wl[466] vdd gnd cell_6t
Xbit_r467_c2 bl[2] br[2] wl[467] vdd gnd cell_6t
Xbit_r468_c2 bl[2] br[2] wl[468] vdd gnd cell_6t
Xbit_r469_c2 bl[2] br[2] wl[469] vdd gnd cell_6t
Xbit_r470_c2 bl[2] br[2] wl[470] vdd gnd cell_6t
Xbit_r471_c2 bl[2] br[2] wl[471] vdd gnd cell_6t
Xbit_r472_c2 bl[2] br[2] wl[472] vdd gnd cell_6t
Xbit_r473_c2 bl[2] br[2] wl[473] vdd gnd cell_6t
Xbit_r474_c2 bl[2] br[2] wl[474] vdd gnd cell_6t
Xbit_r475_c2 bl[2] br[2] wl[475] vdd gnd cell_6t
Xbit_r476_c2 bl[2] br[2] wl[476] vdd gnd cell_6t
Xbit_r477_c2 bl[2] br[2] wl[477] vdd gnd cell_6t
Xbit_r478_c2 bl[2] br[2] wl[478] vdd gnd cell_6t
Xbit_r479_c2 bl[2] br[2] wl[479] vdd gnd cell_6t
Xbit_r480_c2 bl[2] br[2] wl[480] vdd gnd cell_6t
Xbit_r481_c2 bl[2] br[2] wl[481] vdd gnd cell_6t
Xbit_r482_c2 bl[2] br[2] wl[482] vdd gnd cell_6t
Xbit_r483_c2 bl[2] br[2] wl[483] vdd gnd cell_6t
Xbit_r484_c2 bl[2] br[2] wl[484] vdd gnd cell_6t
Xbit_r485_c2 bl[2] br[2] wl[485] vdd gnd cell_6t
Xbit_r486_c2 bl[2] br[2] wl[486] vdd gnd cell_6t
Xbit_r487_c2 bl[2] br[2] wl[487] vdd gnd cell_6t
Xbit_r488_c2 bl[2] br[2] wl[488] vdd gnd cell_6t
Xbit_r489_c2 bl[2] br[2] wl[489] vdd gnd cell_6t
Xbit_r490_c2 bl[2] br[2] wl[490] vdd gnd cell_6t
Xbit_r491_c2 bl[2] br[2] wl[491] vdd gnd cell_6t
Xbit_r492_c2 bl[2] br[2] wl[492] vdd gnd cell_6t
Xbit_r493_c2 bl[2] br[2] wl[493] vdd gnd cell_6t
Xbit_r494_c2 bl[2] br[2] wl[494] vdd gnd cell_6t
Xbit_r495_c2 bl[2] br[2] wl[495] vdd gnd cell_6t
Xbit_r496_c2 bl[2] br[2] wl[496] vdd gnd cell_6t
Xbit_r497_c2 bl[2] br[2] wl[497] vdd gnd cell_6t
Xbit_r498_c2 bl[2] br[2] wl[498] vdd gnd cell_6t
Xbit_r499_c2 bl[2] br[2] wl[499] vdd gnd cell_6t
Xbit_r500_c2 bl[2] br[2] wl[500] vdd gnd cell_6t
Xbit_r501_c2 bl[2] br[2] wl[501] vdd gnd cell_6t
Xbit_r502_c2 bl[2] br[2] wl[502] vdd gnd cell_6t
Xbit_r503_c2 bl[2] br[2] wl[503] vdd gnd cell_6t
Xbit_r504_c2 bl[2] br[2] wl[504] vdd gnd cell_6t
Xbit_r505_c2 bl[2] br[2] wl[505] vdd gnd cell_6t
Xbit_r506_c2 bl[2] br[2] wl[506] vdd gnd cell_6t
Xbit_r507_c2 bl[2] br[2] wl[507] vdd gnd cell_6t
Xbit_r508_c2 bl[2] br[2] wl[508] vdd gnd cell_6t
Xbit_r509_c2 bl[2] br[2] wl[509] vdd gnd cell_6t
Xbit_r510_c2 bl[2] br[2] wl[510] vdd gnd cell_6t
Xbit_r511_c2 bl[2] br[2] wl[511] vdd gnd cell_6t
Xbit_r0_c3 bl[3] br[3] wl[0] vdd gnd cell_6t
Xbit_r1_c3 bl[3] br[3] wl[1] vdd gnd cell_6t
Xbit_r2_c3 bl[3] br[3] wl[2] vdd gnd cell_6t
Xbit_r3_c3 bl[3] br[3] wl[3] vdd gnd cell_6t
Xbit_r4_c3 bl[3] br[3] wl[4] vdd gnd cell_6t
Xbit_r5_c3 bl[3] br[3] wl[5] vdd gnd cell_6t
Xbit_r6_c3 bl[3] br[3] wl[6] vdd gnd cell_6t
Xbit_r7_c3 bl[3] br[3] wl[7] vdd gnd cell_6t
Xbit_r8_c3 bl[3] br[3] wl[8] vdd gnd cell_6t
Xbit_r9_c3 bl[3] br[3] wl[9] vdd gnd cell_6t
Xbit_r10_c3 bl[3] br[3] wl[10] vdd gnd cell_6t
Xbit_r11_c3 bl[3] br[3] wl[11] vdd gnd cell_6t
Xbit_r12_c3 bl[3] br[3] wl[12] vdd gnd cell_6t
Xbit_r13_c3 bl[3] br[3] wl[13] vdd gnd cell_6t
Xbit_r14_c3 bl[3] br[3] wl[14] vdd gnd cell_6t
Xbit_r15_c3 bl[3] br[3] wl[15] vdd gnd cell_6t
Xbit_r16_c3 bl[3] br[3] wl[16] vdd gnd cell_6t
Xbit_r17_c3 bl[3] br[3] wl[17] vdd gnd cell_6t
Xbit_r18_c3 bl[3] br[3] wl[18] vdd gnd cell_6t
Xbit_r19_c3 bl[3] br[3] wl[19] vdd gnd cell_6t
Xbit_r20_c3 bl[3] br[3] wl[20] vdd gnd cell_6t
Xbit_r21_c3 bl[3] br[3] wl[21] vdd gnd cell_6t
Xbit_r22_c3 bl[3] br[3] wl[22] vdd gnd cell_6t
Xbit_r23_c3 bl[3] br[3] wl[23] vdd gnd cell_6t
Xbit_r24_c3 bl[3] br[3] wl[24] vdd gnd cell_6t
Xbit_r25_c3 bl[3] br[3] wl[25] vdd gnd cell_6t
Xbit_r26_c3 bl[3] br[3] wl[26] vdd gnd cell_6t
Xbit_r27_c3 bl[3] br[3] wl[27] vdd gnd cell_6t
Xbit_r28_c3 bl[3] br[3] wl[28] vdd gnd cell_6t
Xbit_r29_c3 bl[3] br[3] wl[29] vdd gnd cell_6t
Xbit_r30_c3 bl[3] br[3] wl[30] vdd gnd cell_6t
Xbit_r31_c3 bl[3] br[3] wl[31] vdd gnd cell_6t
Xbit_r32_c3 bl[3] br[3] wl[32] vdd gnd cell_6t
Xbit_r33_c3 bl[3] br[3] wl[33] vdd gnd cell_6t
Xbit_r34_c3 bl[3] br[3] wl[34] vdd gnd cell_6t
Xbit_r35_c3 bl[3] br[3] wl[35] vdd gnd cell_6t
Xbit_r36_c3 bl[3] br[3] wl[36] vdd gnd cell_6t
Xbit_r37_c3 bl[3] br[3] wl[37] vdd gnd cell_6t
Xbit_r38_c3 bl[3] br[3] wl[38] vdd gnd cell_6t
Xbit_r39_c3 bl[3] br[3] wl[39] vdd gnd cell_6t
Xbit_r40_c3 bl[3] br[3] wl[40] vdd gnd cell_6t
Xbit_r41_c3 bl[3] br[3] wl[41] vdd gnd cell_6t
Xbit_r42_c3 bl[3] br[3] wl[42] vdd gnd cell_6t
Xbit_r43_c3 bl[3] br[3] wl[43] vdd gnd cell_6t
Xbit_r44_c3 bl[3] br[3] wl[44] vdd gnd cell_6t
Xbit_r45_c3 bl[3] br[3] wl[45] vdd gnd cell_6t
Xbit_r46_c3 bl[3] br[3] wl[46] vdd gnd cell_6t
Xbit_r47_c3 bl[3] br[3] wl[47] vdd gnd cell_6t
Xbit_r48_c3 bl[3] br[3] wl[48] vdd gnd cell_6t
Xbit_r49_c3 bl[3] br[3] wl[49] vdd gnd cell_6t
Xbit_r50_c3 bl[3] br[3] wl[50] vdd gnd cell_6t
Xbit_r51_c3 bl[3] br[3] wl[51] vdd gnd cell_6t
Xbit_r52_c3 bl[3] br[3] wl[52] vdd gnd cell_6t
Xbit_r53_c3 bl[3] br[3] wl[53] vdd gnd cell_6t
Xbit_r54_c3 bl[3] br[3] wl[54] vdd gnd cell_6t
Xbit_r55_c3 bl[3] br[3] wl[55] vdd gnd cell_6t
Xbit_r56_c3 bl[3] br[3] wl[56] vdd gnd cell_6t
Xbit_r57_c3 bl[3] br[3] wl[57] vdd gnd cell_6t
Xbit_r58_c3 bl[3] br[3] wl[58] vdd gnd cell_6t
Xbit_r59_c3 bl[3] br[3] wl[59] vdd gnd cell_6t
Xbit_r60_c3 bl[3] br[3] wl[60] vdd gnd cell_6t
Xbit_r61_c3 bl[3] br[3] wl[61] vdd gnd cell_6t
Xbit_r62_c3 bl[3] br[3] wl[62] vdd gnd cell_6t
Xbit_r63_c3 bl[3] br[3] wl[63] vdd gnd cell_6t
Xbit_r64_c3 bl[3] br[3] wl[64] vdd gnd cell_6t
Xbit_r65_c3 bl[3] br[3] wl[65] vdd gnd cell_6t
Xbit_r66_c3 bl[3] br[3] wl[66] vdd gnd cell_6t
Xbit_r67_c3 bl[3] br[3] wl[67] vdd gnd cell_6t
Xbit_r68_c3 bl[3] br[3] wl[68] vdd gnd cell_6t
Xbit_r69_c3 bl[3] br[3] wl[69] vdd gnd cell_6t
Xbit_r70_c3 bl[3] br[3] wl[70] vdd gnd cell_6t
Xbit_r71_c3 bl[3] br[3] wl[71] vdd gnd cell_6t
Xbit_r72_c3 bl[3] br[3] wl[72] vdd gnd cell_6t
Xbit_r73_c3 bl[3] br[3] wl[73] vdd gnd cell_6t
Xbit_r74_c3 bl[3] br[3] wl[74] vdd gnd cell_6t
Xbit_r75_c3 bl[3] br[3] wl[75] vdd gnd cell_6t
Xbit_r76_c3 bl[3] br[3] wl[76] vdd gnd cell_6t
Xbit_r77_c3 bl[3] br[3] wl[77] vdd gnd cell_6t
Xbit_r78_c3 bl[3] br[3] wl[78] vdd gnd cell_6t
Xbit_r79_c3 bl[3] br[3] wl[79] vdd gnd cell_6t
Xbit_r80_c3 bl[3] br[3] wl[80] vdd gnd cell_6t
Xbit_r81_c3 bl[3] br[3] wl[81] vdd gnd cell_6t
Xbit_r82_c3 bl[3] br[3] wl[82] vdd gnd cell_6t
Xbit_r83_c3 bl[3] br[3] wl[83] vdd gnd cell_6t
Xbit_r84_c3 bl[3] br[3] wl[84] vdd gnd cell_6t
Xbit_r85_c3 bl[3] br[3] wl[85] vdd gnd cell_6t
Xbit_r86_c3 bl[3] br[3] wl[86] vdd gnd cell_6t
Xbit_r87_c3 bl[3] br[3] wl[87] vdd gnd cell_6t
Xbit_r88_c3 bl[3] br[3] wl[88] vdd gnd cell_6t
Xbit_r89_c3 bl[3] br[3] wl[89] vdd gnd cell_6t
Xbit_r90_c3 bl[3] br[3] wl[90] vdd gnd cell_6t
Xbit_r91_c3 bl[3] br[3] wl[91] vdd gnd cell_6t
Xbit_r92_c3 bl[3] br[3] wl[92] vdd gnd cell_6t
Xbit_r93_c3 bl[3] br[3] wl[93] vdd gnd cell_6t
Xbit_r94_c3 bl[3] br[3] wl[94] vdd gnd cell_6t
Xbit_r95_c3 bl[3] br[3] wl[95] vdd gnd cell_6t
Xbit_r96_c3 bl[3] br[3] wl[96] vdd gnd cell_6t
Xbit_r97_c3 bl[3] br[3] wl[97] vdd gnd cell_6t
Xbit_r98_c3 bl[3] br[3] wl[98] vdd gnd cell_6t
Xbit_r99_c3 bl[3] br[3] wl[99] vdd gnd cell_6t
Xbit_r100_c3 bl[3] br[3] wl[100] vdd gnd cell_6t
Xbit_r101_c3 bl[3] br[3] wl[101] vdd gnd cell_6t
Xbit_r102_c3 bl[3] br[3] wl[102] vdd gnd cell_6t
Xbit_r103_c3 bl[3] br[3] wl[103] vdd gnd cell_6t
Xbit_r104_c3 bl[3] br[3] wl[104] vdd gnd cell_6t
Xbit_r105_c3 bl[3] br[3] wl[105] vdd gnd cell_6t
Xbit_r106_c3 bl[3] br[3] wl[106] vdd gnd cell_6t
Xbit_r107_c3 bl[3] br[3] wl[107] vdd gnd cell_6t
Xbit_r108_c3 bl[3] br[3] wl[108] vdd gnd cell_6t
Xbit_r109_c3 bl[3] br[3] wl[109] vdd gnd cell_6t
Xbit_r110_c3 bl[3] br[3] wl[110] vdd gnd cell_6t
Xbit_r111_c3 bl[3] br[3] wl[111] vdd gnd cell_6t
Xbit_r112_c3 bl[3] br[3] wl[112] vdd gnd cell_6t
Xbit_r113_c3 bl[3] br[3] wl[113] vdd gnd cell_6t
Xbit_r114_c3 bl[3] br[3] wl[114] vdd gnd cell_6t
Xbit_r115_c3 bl[3] br[3] wl[115] vdd gnd cell_6t
Xbit_r116_c3 bl[3] br[3] wl[116] vdd gnd cell_6t
Xbit_r117_c3 bl[3] br[3] wl[117] vdd gnd cell_6t
Xbit_r118_c3 bl[3] br[3] wl[118] vdd gnd cell_6t
Xbit_r119_c3 bl[3] br[3] wl[119] vdd gnd cell_6t
Xbit_r120_c3 bl[3] br[3] wl[120] vdd gnd cell_6t
Xbit_r121_c3 bl[3] br[3] wl[121] vdd gnd cell_6t
Xbit_r122_c3 bl[3] br[3] wl[122] vdd gnd cell_6t
Xbit_r123_c3 bl[3] br[3] wl[123] vdd gnd cell_6t
Xbit_r124_c3 bl[3] br[3] wl[124] vdd gnd cell_6t
Xbit_r125_c3 bl[3] br[3] wl[125] vdd gnd cell_6t
Xbit_r126_c3 bl[3] br[3] wl[126] vdd gnd cell_6t
Xbit_r127_c3 bl[3] br[3] wl[127] vdd gnd cell_6t
Xbit_r128_c3 bl[3] br[3] wl[128] vdd gnd cell_6t
Xbit_r129_c3 bl[3] br[3] wl[129] vdd gnd cell_6t
Xbit_r130_c3 bl[3] br[3] wl[130] vdd gnd cell_6t
Xbit_r131_c3 bl[3] br[3] wl[131] vdd gnd cell_6t
Xbit_r132_c3 bl[3] br[3] wl[132] vdd gnd cell_6t
Xbit_r133_c3 bl[3] br[3] wl[133] vdd gnd cell_6t
Xbit_r134_c3 bl[3] br[3] wl[134] vdd gnd cell_6t
Xbit_r135_c3 bl[3] br[3] wl[135] vdd gnd cell_6t
Xbit_r136_c3 bl[3] br[3] wl[136] vdd gnd cell_6t
Xbit_r137_c3 bl[3] br[3] wl[137] vdd gnd cell_6t
Xbit_r138_c3 bl[3] br[3] wl[138] vdd gnd cell_6t
Xbit_r139_c3 bl[3] br[3] wl[139] vdd gnd cell_6t
Xbit_r140_c3 bl[3] br[3] wl[140] vdd gnd cell_6t
Xbit_r141_c3 bl[3] br[3] wl[141] vdd gnd cell_6t
Xbit_r142_c3 bl[3] br[3] wl[142] vdd gnd cell_6t
Xbit_r143_c3 bl[3] br[3] wl[143] vdd gnd cell_6t
Xbit_r144_c3 bl[3] br[3] wl[144] vdd gnd cell_6t
Xbit_r145_c3 bl[3] br[3] wl[145] vdd gnd cell_6t
Xbit_r146_c3 bl[3] br[3] wl[146] vdd gnd cell_6t
Xbit_r147_c3 bl[3] br[3] wl[147] vdd gnd cell_6t
Xbit_r148_c3 bl[3] br[3] wl[148] vdd gnd cell_6t
Xbit_r149_c3 bl[3] br[3] wl[149] vdd gnd cell_6t
Xbit_r150_c3 bl[3] br[3] wl[150] vdd gnd cell_6t
Xbit_r151_c3 bl[3] br[3] wl[151] vdd gnd cell_6t
Xbit_r152_c3 bl[3] br[3] wl[152] vdd gnd cell_6t
Xbit_r153_c3 bl[3] br[3] wl[153] vdd gnd cell_6t
Xbit_r154_c3 bl[3] br[3] wl[154] vdd gnd cell_6t
Xbit_r155_c3 bl[3] br[3] wl[155] vdd gnd cell_6t
Xbit_r156_c3 bl[3] br[3] wl[156] vdd gnd cell_6t
Xbit_r157_c3 bl[3] br[3] wl[157] vdd gnd cell_6t
Xbit_r158_c3 bl[3] br[3] wl[158] vdd gnd cell_6t
Xbit_r159_c3 bl[3] br[3] wl[159] vdd gnd cell_6t
Xbit_r160_c3 bl[3] br[3] wl[160] vdd gnd cell_6t
Xbit_r161_c3 bl[3] br[3] wl[161] vdd gnd cell_6t
Xbit_r162_c3 bl[3] br[3] wl[162] vdd gnd cell_6t
Xbit_r163_c3 bl[3] br[3] wl[163] vdd gnd cell_6t
Xbit_r164_c3 bl[3] br[3] wl[164] vdd gnd cell_6t
Xbit_r165_c3 bl[3] br[3] wl[165] vdd gnd cell_6t
Xbit_r166_c3 bl[3] br[3] wl[166] vdd gnd cell_6t
Xbit_r167_c3 bl[3] br[3] wl[167] vdd gnd cell_6t
Xbit_r168_c3 bl[3] br[3] wl[168] vdd gnd cell_6t
Xbit_r169_c3 bl[3] br[3] wl[169] vdd gnd cell_6t
Xbit_r170_c3 bl[3] br[3] wl[170] vdd gnd cell_6t
Xbit_r171_c3 bl[3] br[3] wl[171] vdd gnd cell_6t
Xbit_r172_c3 bl[3] br[3] wl[172] vdd gnd cell_6t
Xbit_r173_c3 bl[3] br[3] wl[173] vdd gnd cell_6t
Xbit_r174_c3 bl[3] br[3] wl[174] vdd gnd cell_6t
Xbit_r175_c3 bl[3] br[3] wl[175] vdd gnd cell_6t
Xbit_r176_c3 bl[3] br[3] wl[176] vdd gnd cell_6t
Xbit_r177_c3 bl[3] br[3] wl[177] vdd gnd cell_6t
Xbit_r178_c3 bl[3] br[3] wl[178] vdd gnd cell_6t
Xbit_r179_c3 bl[3] br[3] wl[179] vdd gnd cell_6t
Xbit_r180_c3 bl[3] br[3] wl[180] vdd gnd cell_6t
Xbit_r181_c3 bl[3] br[3] wl[181] vdd gnd cell_6t
Xbit_r182_c3 bl[3] br[3] wl[182] vdd gnd cell_6t
Xbit_r183_c3 bl[3] br[3] wl[183] vdd gnd cell_6t
Xbit_r184_c3 bl[3] br[3] wl[184] vdd gnd cell_6t
Xbit_r185_c3 bl[3] br[3] wl[185] vdd gnd cell_6t
Xbit_r186_c3 bl[3] br[3] wl[186] vdd gnd cell_6t
Xbit_r187_c3 bl[3] br[3] wl[187] vdd gnd cell_6t
Xbit_r188_c3 bl[3] br[3] wl[188] vdd gnd cell_6t
Xbit_r189_c3 bl[3] br[3] wl[189] vdd gnd cell_6t
Xbit_r190_c3 bl[3] br[3] wl[190] vdd gnd cell_6t
Xbit_r191_c3 bl[3] br[3] wl[191] vdd gnd cell_6t
Xbit_r192_c3 bl[3] br[3] wl[192] vdd gnd cell_6t
Xbit_r193_c3 bl[3] br[3] wl[193] vdd gnd cell_6t
Xbit_r194_c3 bl[3] br[3] wl[194] vdd gnd cell_6t
Xbit_r195_c3 bl[3] br[3] wl[195] vdd gnd cell_6t
Xbit_r196_c3 bl[3] br[3] wl[196] vdd gnd cell_6t
Xbit_r197_c3 bl[3] br[3] wl[197] vdd gnd cell_6t
Xbit_r198_c3 bl[3] br[3] wl[198] vdd gnd cell_6t
Xbit_r199_c3 bl[3] br[3] wl[199] vdd gnd cell_6t
Xbit_r200_c3 bl[3] br[3] wl[200] vdd gnd cell_6t
Xbit_r201_c3 bl[3] br[3] wl[201] vdd gnd cell_6t
Xbit_r202_c3 bl[3] br[3] wl[202] vdd gnd cell_6t
Xbit_r203_c3 bl[3] br[3] wl[203] vdd gnd cell_6t
Xbit_r204_c3 bl[3] br[3] wl[204] vdd gnd cell_6t
Xbit_r205_c3 bl[3] br[3] wl[205] vdd gnd cell_6t
Xbit_r206_c3 bl[3] br[3] wl[206] vdd gnd cell_6t
Xbit_r207_c3 bl[3] br[3] wl[207] vdd gnd cell_6t
Xbit_r208_c3 bl[3] br[3] wl[208] vdd gnd cell_6t
Xbit_r209_c3 bl[3] br[3] wl[209] vdd gnd cell_6t
Xbit_r210_c3 bl[3] br[3] wl[210] vdd gnd cell_6t
Xbit_r211_c3 bl[3] br[3] wl[211] vdd gnd cell_6t
Xbit_r212_c3 bl[3] br[3] wl[212] vdd gnd cell_6t
Xbit_r213_c3 bl[3] br[3] wl[213] vdd gnd cell_6t
Xbit_r214_c3 bl[3] br[3] wl[214] vdd gnd cell_6t
Xbit_r215_c3 bl[3] br[3] wl[215] vdd gnd cell_6t
Xbit_r216_c3 bl[3] br[3] wl[216] vdd gnd cell_6t
Xbit_r217_c3 bl[3] br[3] wl[217] vdd gnd cell_6t
Xbit_r218_c3 bl[3] br[3] wl[218] vdd gnd cell_6t
Xbit_r219_c3 bl[3] br[3] wl[219] vdd gnd cell_6t
Xbit_r220_c3 bl[3] br[3] wl[220] vdd gnd cell_6t
Xbit_r221_c3 bl[3] br[3] wl[221] vdd gnd cell_6t
Xbit_r222_c3 bl[3] br[3] wl[222] vdd gnd cell_6t
Xbit_r223_c3 bl[3] br[3] wl[223] vdd gnd cell_6t
Xbit_r224_c3 bl[3] br[3] wl[224] vdd gnd cell_6t
Xbit_r225_c3 bl[3] br[3] wl[225] vdd gnd cell_6t
Xbit_r226_c3 bl[3] br[3] wl[226] vdd gnd cell_6t
Xbit_r227_c3 bl[3] br[3] wl[227] vdd gnd cell_6t
Xbit_r228_c3 bl[3] br[3] wl[228] vdd gnd cell_6t
Xbit_r229_c3 bl[3] br[3] wl[229] vdd gnd cell_6t
Xbit_r230_c3 bl[3] br[3] wl[230] vdd gnd cell_6t
Xbit_r231_c3 bl[3] br[3] wl[231] vdd gnd cell_6t
Xbit_r232_c3 bl[3] br[3] wl[232] vdd gnd cell_6t
Xbit_r233_c3 bl[3] br[3] wl[233] vdd gnd cell_6t
Xbit_r234_c3 bl[3] br[3] wl[234] vdd gnd cell_6t
Xbit_r235_c3 bl[3] br[3] wl[235] vdd gnd cell_6t
Xbit_r236_c3 bl[3] br[3] wl[236] vdd gnd cell_6t
Xbit_r237_c3 bl[3] br[3] wl[237] vdd gnd cell_6t
Xbit_r238_c3 bl[3] br[3] wl[238] vdd gnd cell_6t
Xbit_r239_c3 bl[3] br[3] wl[239] vdd gnd cell_6t
Xbit_r240_c3 bl[3] br[3] wl[240] vdd gnd cell_6t
Xbit_r241_c3 bl[3] br[3] wl[241] vdd gnd cell_6t
Xbit_r242_c3 bl[3] br[3] wl[242] vdd gnd cell_6t
Xbit_r243_c3 bl[3] br[3] wl[243] vdd gnd cell_6t
Xbit_r244_c3 bl[3] br[3] wl[244] vdd gnd cell_6t
Xbit_r245_c3 bl[3] br[3] wl[245] vdd gnd cell_6t
Xbit_r246_c3 bl[3] br[3] wl[246] vdd gnd cell_6t
Xbit_r247_c3 bl[3] br[3] wl[247] vdd gnd cell_6t
Xbit_r248_c3 bl[3] br[3] wl[248] vdd gnd cell_6t
Xbit_r249_c3 bl[3] br[3] wl[249] vdd gnd cell_6t
Xbit_r250_c3 bl[3] br[3] wl[250] vdd gnd cell_6t
Xbit_r251_c3 bl[3] br[3] wl[251] vdd gnd cell_6t
Xbit_r252_c3 bl[3] br[3] wl[252] vdd gnd cell_6t
Xbit_r253_c3 bl[3] br[3] wl[253] vdd gnd cell_6t
Xbit_r254_c3 bl[3] br[3] wl[254] vdd gnd cell_6t
Xbit_r255_c3 bl[3] br[3] wl[255] vdd gnd cell_6t
Xbit_r256_c3 bl[3] br[3] wl[256] vdd gnd cell_6t
Xbit_r257_c3 bl[3] br[3] wl[257] vdd gnd cell_6t
Xbit_r258_c3 bl[3] br[3] wl[258] vdd gnd cell_6t
Xbit_r259_c3 bl[3] br[3] wl[259] vdd gnd cell_6t
Xbit_r260_c3 bl[3] br[3] wl[260] vdd gnd cell_6t
Xbit_r261_c3 bl[3] br[3] wl[261] vdd gnd cell_6t
Xbit_r262_c3 bl[3] br[3] wl[262] vdd gnd cell_6t
Xbit_r263_c3 bl[3] br[3] wl[263] vdd gnd cell_6t
Xbit_r264_c3 bl[3] br[3] wl[264] vdd gnd cell_6t
Xbit_r265_c3 bl[3] br[3] wl[265] vdd gnd cell_6t
Xbit_r266_c3 bl[3] br[3] wl[266] vdd gnd cell_6t
Xbit_r267_c3 bl[3] br[3] wl[267] vdd gnd cell_6t
Xbit_r268_c3 bl[3] br[3] wl[268] vdd gnd cell_6t
Xbit_r269_c3 bl[3] br[3] wl[269] vdd gnd cell_6t
Xbit_r270_c3 bl[3] br[3] wl[270] vdd gnd cell_6t
Xbit_r271_c3 bl[3] br[3] wl[271] vdd gnd cell_6t
Xbit_r272_c3 bl[3] br[3] wl[272] vdd gnd cell_6t
Xbit_r273_c3 bl[3] br[3] wl[273] vdd gnd cell_6t
Xbit_r274_c3 bl[3] br[3] wl[274] vdd gnd cell_6t
Xbit_r275_c3 bl[3] br[3] wl[275] vdd gnd cell_6t
Xbit_r276_c3 bl[3] br[3] wl[276] vdd gnd cell_6t
Xbit_r277_c3 bl[3] br[3] wl[277] vdd gnd cell_6t
Xbit_r278_c3 bl[3] br[3] wl[278] vdd gnd cell_6t
Xbit_r279_c3 bl[3] br[3] wl[279] vdd gnd cell_6t
Xbit_r280_c3 bl[3] br[3] wl[280] vdd gnd cell_6t
Xbit_r281_c3 bl[3] br[3] wl[281] vdd gnd cell_6t
Xbit_r282_c3 bl[3] br[3] wl[282] vdd gnd cell_6t
Xbit_r283_c3 bl[3] br[3] wl[283] vdd gnd cell_6t
Xbit_r284_c3 bl[3] br[3] wl[284] vdd gnd cell_6t
Xbit_r285_c3 bl[3] br[3] wl[285] vdd gnd cell_6t
Xbit_r286_c3 bl[3] br[3] wl[286] vdd gnd cell_6t
Xbit_r287_c3 bl[3] br[3] wl[287] vdd gnd cell_6t
Xbit_r288_c3 bl[3] br[3] wl[288] vdd gnd cell_6t
Xbit_r289_c3 bl[3] br[3] wl[289] vdd gnd cell_6t
Xbit_r290_c3 bl[3] br[3] wl[290] vdd gnd cell_6t
Xbit_r291_c3 bl[3] br[3] wl[291] vdd gnd cell_6t
Xbit_r292_c3 bl[3] br[3] wl[292] vdd gnd cell_6t
Xbit_r293_c3 bl[3] br[3] wl[293] vdd gnd cell_6t
Xbit_r294_c3 bl[3] br[3] wl[294] vdd gnd cell_6t
Xbit_r295_c3 bl[3] br[3] wl[295] vdd gnd cell_6t
Xbit_r296_c3 bl[3] br[3] wl[296] vdd gnd cell_6t
Xbit_r297_c3 bl[3] br[3] wl[297] vdd gnd cell_6t
Xbit_r298_c3 bl[3] br[3] wl[298] vdd gnd cell_6t
Xbit_r299_c3 bl[3] br[3] wl[299] vdd gnd cell_6t
Xbit_r300_c3 bl[3] br[3] wl[300] vdd gnd cell_6t
Xbit_r301_c3 bl[3] br[3] wl[301] vdd gnd cell_6t
Xbit_r302_c3 bl[3] br[3] wl[302] vdd gnd cell_6t
Xbit_r303_c3 bl[3] br[3] wl[303] vdd gnd cell_6t
Xbit_r304_c3 bl[3] br[3] wl[304] vdd gnd cell_6t
Xbit_r305_c3 bl[3] br[3] wl[305] vdd gnd cell_6t
Xbit_r306_c3 bl[3] br[3] wl[306] vdd gnd cell_6t
Xbit_r307_c3 bl[3] br[3] wl[307] vdd gnd cell_6t
Xbit_r308_c3 bl[3] br[3] wl[308] vdd gnd cell_6t
Xbit_r309_c3 bl[3] br[3] wl[309] vdd gnd cell_6t
Xbit_r310_c3 bl[3] br[3] wl[310] vdd gnd cell_6t
Xbit_r311_c3 bl[3] br[3] wl[311] vdd gnd cell_6t
Xbit_r312_c3 bl[3] br[3] wl[312] vdd gnd cell_6t
Xbit_r313_c3 bl[3] br[3] wl[313] vdd gnd cell_6t
Xbit_r314_c3 bl[3] br[3] wl[314] vdd gnd cell_6t
Xbit_r315_c3 bl[3] br[3] wl[315] vdd gnd cell_6t
Xbit_r316_c3 bl[3] br[3] wl[316] vdd gnd cell_6t
Xbit_r317_c3 bl[3] br[3] wl[317] vdd gnd cell_6t
Xbit_r318_c3 bl[3] br[3] wl[318] vdd gnd cell_6t
Xbit_r319_c3 bl[3] br[3] wl[319] vdd gnd cell_6t
Xbit_r320_c3 bl[3] br[3] wl[320] vdd gnd cell_6t
Xbit_r321_c3 bl[3] br[3] wl[321] vdd gnd cell_6t
Xbit_r322_c3 bl[3] br[3] wl[322] vdd gnd cell_6t
Xbit_r323_c3 bl[3] br[3] wl[323] vdd gnd cell_6t
Xbit_r324_c3 bl[3] br[3] wl[324] vdd gnd cell_6t
Xbit_r325_c3 bl[3] br[3] wl[325] vdd gnd cell_6t
Xbit_r326_c3 bl[3] br[3] wl[326] vdd gnd cell_6t
Xbit_r327_c3 bl[3] br[3] wl[327] vdd gnd cell_6t
Xbit_r328_c3 bl[3] br[3] wl[328] vdd gnd cell_6t
Xbit_r329_c3 bl[3] br[3] wl[329] vdd gnd cell_6t
Xbit_r330_c3 bl[3] br[3] wl[330] vdd gnd cell_6t
Xbit_r331_c3 bl[3] br[3] wl[331] vdd gnd cell_6t
Xbit_r332_c3 bl[3] br[3] wl[332] vdd gnd cell_6t
Xbit_r333_c3 bl[3] br[3] wl[333] vdd gnd cell_6t
Xbit_r334_c3 bl[3] br[3] wl[334] vdd gnd cell_6t
Xbit_r335_c3 bl[3] br[3] wl[335] vdd gnd cell_6t
Xbit_r336_c3 bl[3] br[3] wl[336] vdd gnd cell_6t
Xbit_r337_c3 bl[3] br[3] wl[337] vdd gnd cell_6t
Xbit_r338_c3 bl[3] br[3] wl[338] vdd gnd cell_6t
Xbit_r339_c3 bl[3] br[3] wl[339] vdd gnd cell_6t
Xbit_r340_c3 bl[3] br[3] wl[340] vdd gnd cell_6t
Xbit_r341_c3 bl[3] br[3] wl[341] vdd gnd cell_6t
Xbit_r342_c3 bl[3] br[3] wl[342] vdd gnd cell_6t
Xbit_r343_c3 bl[3] br[3] wl[343] vdd gnd cell_6t
Xbit_r344_c3 bl[3] br[3] wl[344] vdd gnd cell_6t
Xbit_r345_c3 bl[3] br[3] wl[345] vdd gnd cell_6t
Xbit_r346_c3 bl[3] br[3] wl[346] vdd gnd cell_6t
Xbit_r347_c3 bl[3] br[3] wl[347] vdd gnd cell_6t
Xbit_r348_c3 bl[3] br[3] wl[348] vdd gnd cell_6t
Xbit_r349_c3 bl[3] br[3] wl[349] vdd gnd cell_6t
Xbit_r350_c3 bl[3] br[3] wl[350] vdd gnd cell_6t
Xbit_r351_c3 bl[3] br[3] wl[351] vdd gnd cell_6t
Xbit_r352_c3 bl[3] br[3] wl[352] vdd gnd cell_6t
Xbit_r353_c3 bl[3] br[3] wl[353] vdd gnd cell_6t
Xbit_r354_c3 bl[3] br[3] wl[354] vdd gnd cell_6t
Xbit_r355_c3 bl[3] br[3] wl[355] vdd gnd cell_6t
Xbit_r356_c3 bl[3] br[3] wl[356] vdd gnd cell_6t
Xbit_r357_c3 bl[3] br[3] wl[357] vdd gnd cell_6t
Xbit_r358_c3 bl[3] br[3] wl[358] vdd gnd cell_6t
Xbit_r359_c3 bl[3] br[3] wl[359] vdd gnd cell_6t
Xbit_r360_c3 bl[3] br[3] wl[360] vdd gnd cell_6t
Xbit_r361_c3 bl[3] br[3] wl[361] vdd gnd cell_6t
Xbit_r362_c3 bl[3] br[3] wl[362] vdd gnd cell_6t
Xbit_r363_c3 bl[3] br[3] wl[363] vdd gnd cell_6t
Xbit_r364_c3 bl[3] br[3] wl[364] vdd gnd cell_6t
Xbit_r365_c3 bl[3] br[3] wl[365] vdd gnd cell_6t
Xbit_r366_c3 bl[3] br[3] wl[366] vdd gnd cell_6t
Xbit_r367_c3 bl[3] br[3] wl[367] vdd gnd cell_6t
Xbit_r368_c3 bl[3] br[3] wl[368] vdd gnd cell_6t
Xbit_r369_c3 bl[3] br[3] wl[369] vdd gnd cell_6t
Xbit_r370_c3 bl[3] br[3] wl[370] vdd gnd cell_6t
Xbit_r371_c3 bl[3] br[3] wl[371] vdd gnd cell_6t
Xbit_r372_c3 bl[3] br[3] wl[372] vdd gnd cell_6t
Xbit_r373_c3 bl[3] br[3] wl[373] vdd gnd cell_6t
Xbit_r374_c3 bl[3] br[3] wl[374] vdd gnd cell_6t
Xbit_r375_c3 bl[3] br[3] wl[375] vdd gnd cell_6t
Xbit_r376_c3 bl[3] br[3] wl[376] vdd gnd cell_6t
Xbit_r377_c3 bl[3] br[3] wl[377] vdd gnd cell_6t
Xbit_r378_c3 bl[3] br[3] wl[378] vdd gnd cell_6t
Xbit_r379_c3 bl[3] br[3] wl[379] vdd gnd cell_6t
Xbit_r380_c3 bl[3] br[3] wl[380] vdd gnd cell_6t
Xbit_r381_c3 bl[3] br[3] wl[381] vdd gnd cell_6t
Xbit_r382_c3 bl[3] br[3] wl[382] vdd gnd cell_6t
Xbit_r383_c3 bl[3] br[3] wl[383] vdd gnd cell_6t
Xbit_r384_c3 bl[3] br[3] wl[384] vdd gnd cell_6t
Xbit_r385_c3 bl[3] br[3] wl[385] vdd gnd cell_6t
Xbit_r386_c3 bl[3] br[3] wl[386] vdd gnd cell_6t
Xbit_r387_c3 bl[3] br[3] wl[387] vdd gnd cell_6t
Xbit_r388_c3 bl[3] br[3] wl[388] vdd gnd cell_6t
Xbit_r389_c3 bl[3] br[3] wl[389] vdd gnd cell_6t
Xbit_r390_c3 bl[3] br[3] wl[390] vdd gnd cell_6t
Xbit_r391_c3 bl[3] br[3] wl[391] vdd gnd cell_6t
Xbit_r392_c3 bl[3] br[3] wl[392] vdd gnd cell_6t
Xbit_r393_c3 bl[3] br[3] wl[393] vdd gnd cell_6t
Xbit_r394_c3 bl[3] br[3] wl[394] vdd gnd cell_6t
Xbit_r395_c3 bl[3] br[3] wl[395] vdd gnd cell_6t
Xbit_r396_c3 bl[3] br[3] wl[396] vdd gnd cell_6t
Xbit_r397_c3 bl[3] br[3] wl[397] vdd gnd cell_6t
Xbit_r398_c3 bl[3] br[3] wl[398] vdd gnd cell_6t
Xbit_r399_c3 bl[3] br[3] wl[399] vdd gnd cell_6t
Xbit_r400_c3 bl[3] br[3] wl[400] vdd gnd cell_6t
Xbit_r401_c3 bl[3] br[3] wl[401] vdd gnd cell_6t
Xbit_r402_c3 bl[3] br[3] wl[402] vdd gnd cell_6t
Xbit_r403_c3 bl[3] br[3] wl[403] vdd gnd cell_6t
Xbit_r404_c3 bl[3] br[3] wl[404] vdd gnd cell_6t
Xbit_r405_c3 bl[3] br[3] wl[405] vdd gnd cell_6t
Xbit_r406_c3 bl[3] br[3] wl[406] vdd gnd cell_6t
Xbit_r407_c3 bl[3] br[3] wl[407] vdd gnd cell_6t
Xbit_r408_c3 bl[3] br[3] wl[408] vdd gnd cell_6t
Xbit_r409_c3 bl[3] br[3] wl[409] vdd gnd cell_6t
Xbit_r410_c3 bl[3] br[3] wl[410] vdd gnd cell_6t
Xbit_r411_c3 bl[3] br[3] wl[411] vdd gnd cell_6t
Xbit_r412_c3 bl[3] br[3] wl[412] vdd gnd cell_6t
Xbit_r413_c3 bl[3] br[3] wl[413] vdd gnd cell_6t
Xbit_r414_c3 bl[3] br[3] wl[414] vdd gnd cell_6t
Xbit_r415_c3 bl[3] br[3] wl[415] vdd gnd cell_6t
Xbit_r416_c3 bl[3] br[3] wl[416] vdd gnd cell_6t
Xbit_r417_c3 bl[3] br[3] wl[417] vdd gnd cell_6t
Xbit_r418_c3 bl[3] br[3] wl[418] vdd gnd cell_6t
Xbit_r419_c3 bl[3] br[3] wl[419] vdd gnd cell_6t
Xbit_r420_c3 bl[3] br[3] wl[420] vdd gnd cell_6t
Xbit_r421_c3 bl[3] br[3] wl[421] vdd gnd cell_6t
Xbit_r422_c3 bl[3] br[3] wl[422] vdd gnd cell_6t
Xbit_r423_c3 bl[3] br[3] wl[423] vdd gnd cell_6t
Xbit_r424_c3 bl[3] br[3] wl[424] vdd gnd cell_6t
Xbit_r425_c3 bl[3] br[3] wl[425] vdd gnd cell_6t
Xbit_r426_c3 bl[3] br[3] wl[426] vdd gnd cell_6t
Xbit_r427_c3 bl[3] br[3] wl[427] vdd gnd cell_6t
Xbit_r428_c3 bl[3] br[3] wl[428] vdd gnd cell_6t
Xbit_r429_c3 bl[3] br[3] wl[429] vdd gnd cell_6t
Xbit_r430_c3 bl[3] br[3] wl[430] vdd gnd cell_6t
Xbit_r431_c3 bl[3] br[3] wl[431] vdd gnd cell_6t
Xbit_r432_c3 bl[3] br[3] wl[432] vdd gnd cell_6t
Xbit_r433_c3 bl[3] br[3] wl[433] vdd gnd cell_6t
Xbit_r434_c3 bl[3] br[3] wl[434] vdd gnd cell_6t
Xbit_r435_c3 bl[3] br[3] wl[435] vdd gnd cell_6t
Xbit_r436_c3 bl[3] br[3] wl[436] vdd gnd cell_6t
Xbit_r437_c3 bl[3] br[3] wl[437] vdd gnd cell_6t
Xbit_r438_c3 bl[3] br[3] wl[438] vdd gnd cell_6t
Xbit_r439_c3 bl[3] br[3] wl[439] vdd gnd cell_6t
Xbit_r440_c3 bl[3] br[3] wl[440] vdd gnd cell_6t
Xbit_r441_c3 bl[3] br[3] wl[441] vdd gnd cell_6t
Xbit_r442_c3 bl[3] br[3] wl[442] vdd gnd cell_6t
Xbit_r443_c3 bl[3] br[3] wl[443] vdd gnd cell_6t
Xbit_r444_c3 bl[3] br[3] wl[444] vdd gnd cell_6t
Xbit_r445_c3 bl[3] br[3] wl[445] vdd gnd cell_6t
Xbit_r446_c3 bl[3] br[3] wl[446] vdd gnd cell_6t
Xbit_r447_c3 bl[3] br[3] wl[447] vdd gnd cell_6t
Xbit_r448_c3 bl[3] br[3] wl[448] vdd gnd cell_6t
Xbit_r449_c3 bl[3] br[3] wl[449] vdd gnd cell_6t
Xbit_r450_c3 bl[3] br[3] wl[450] vdd gnd cell_6t
Xbit_r451_c3 bl[3] br[3] wl[451] vdd gnd cell_6t
Xbit_r452_c3 bl[3] br[3] wl[452] vdd gnd cell_6t
Xbit_r453_c3 bl[3] br[3] wl[453] vdd gnd cell_6t
Xbit_r454_c3 bl[3] br[3] wl[454] vdd gnd cell_6t
Xbit_r455_c3 bl[3] br[3] wl[455] vdd gnd cell_6t
Xbit_r456_c3 bl[3] br[3] wl[456] vdd gnd cell_6t
Xbit_r457_c3 bl[3] br[3] wl[457] vdd gnd cell_6t
Xbit_r458_c3 bl[3] br[3] wl[458] vdd gnd cell_6t
Xbit_r459_c3 bl[3] br[3] wl[459] vdd gnd cell_6t
Xbit_r460_c3 bl[3] br[3] wl[460] vdd gnd cell_6t
Xbit_r461_c3 bl[3] br[3] wl[461] vdd gnd cell_6t
Xbit_r462_c3 bl[3] br[3] wl[462] vdd gnd cell_6t
Xbit_r463_c3 bl[3] br[3] wl[463] vdd gnd cell_6t
Xbit_r464_c3 bl[3] br[3] wl[464] vdd gnd cell_6t
Xbit_r465_c3 bl[3] br[3] wl[465] vdd gnd cell_6t
Xbit_r466_c3 bl[3] br[3] wl[466] vdd gnd cell_6t
Xbit_r467_c3 bl[3] br[3] wl[467] vdd gnd cell_6t
Xbit_r468_c3 bl[3] br[3] wl[468] vdd gnd cell_6t
Xbit_r469_c3 bl[3] br[3] wl[469] vdd gnd cell_6t
Xbit_r470_c3 bl[3] br[3] wl[470] vdd gnd cell_6t
Xbit_r471_c3 bl[3] br[3] wl[471] vdd gnd cell_6t
Xbit_r472_c3 bl[3] br[3] wl[472] vdd gnd cell_6t
Xbit_r473_c3 bl[3] br[3] wl[473] vdd gnd cell_6t
Xbit_r474_c3 bl[3] br[3] wl[474] vdd gnd cell_6t
Xbit_r475_c3 bl[3] br[3] wl[475] vdd gnd cell_6t
Xbit_r476_c3 bl[3] br[3] wl[476] vdd gnd cell_6t
Xbit_r477_c3 bl[3] br[3] wl[477] vdd gnd cell_6t
Xbit_r478_c3 bl[3] br[3] wl[478] vdd gnd cell_6t
Xbit_r479_c3 bl[3] br[3] wl[479] vdd gnd cell_6t
Xbit_r480_c3 bl[3] br[3] wl[480] vdd gnd cell_6t
Xbit_r481_c3 bl[3] br[3] wl[481] vdd gnd cell_6t
Xbit_r482_c3 bl[3] br[3] wl[482] vdd gnd cell_6t
Xbit_r483_c3 bl[3] br[3] wl[483] vdd gnd cell_6t
Xbit_r484_c3 bl[3] br[3] wl[484] vdd gnd cell_6t
Xbit_r485_c3 bl[3] br[3] wl[485] vdd gnd cell_6t
Xbit_r486_c3 bl[3] br[3] wl[486] vdd gnd cell_6t
Xbit_r487_c3 bl[3] br[3] wl[487] vdd gnd cell_6t
Xbit_r488_c3 bl[3] br[3] wl[488] vdd gnd cell_6t
Xbit_r489_c3 bl[3] br[3] wl[489] vdd gnd cell_6t
Xbit_r490_c3 bl[3] br[3] wl[490] vdd gnd cell_6t
Xbit_r491_c3 bl[3] br[3] wl[491] vdd gnd cell_6t
Xbit_r492_c3 bl[3] br[3] wl[492] vdd gnd cell_6t
Xbit_r493_c3 bl[3] br[3] wl[493] vdd gnd cell_6t
Xbit_r494_c3 bl[3] br[3] wl[494] vdd gnd cell_6t
Xbit_r495_c3 bl[3] br[3] wl[495] vdd gnd cell_6t
Xbit_r496_c3 bl[3] br[3] wl[496] vdd gnd cell_6t
Xbit_r497_c3 bl[3] br[3] wl[497] vdd gnd cell_6t
Xbit_r498_c3 bl[3] br[3] wl[498] vdd gnd cell_6t
Xbit_r499_c3 bl[3] br[3] wl[499] vdd gnd cell_6t
Xbit_r500_c3 bl[3] br[3] wl[500] vdd gnd cell_6t
Xbit_r501_c3 bl[3] br[3] wl[501] vdd gnd cell_6t
Xbit_r502_c3 bl[3] br[3] wl[502] vdd gnd cell_6t
Xbit_r503_c3 bl[3] br[3] wl[503] vdd gnd cell_6t
Xbit_r504_c3 bl[3] br[3] wl[504] vdd gnd cell_6t
Xbit_r505_c3 bl[3] br[3] wl[505] vdd gnd cell_6t
Xbit_r506_c3 bl[3] br[3] wl[506] vdd gnd cell_6t
Xbit_r507_c3 bl[3] br[3] wl[507] vdd gnd cell_6t
Xbit_r508_c3 bl[3] br[3] wl[508] vdd gnd cell_6t
Xbit_r509_c3 bl[3] br[3] wl[509] vdd gnd cell_6t
Xbit_r510_c3 bl[3] br[3] wl[510] vdd gnd cell_6t
Xbit_r511_c3 bl[3] br[3] wl[511] vdd gnd cell_6t
Xbit_r0_c4 bl[4] br[4] wl[0] vdd gnd cell_6t
Xbit_r1_c4 bl[4] br[4] wl[1] vdd gnd cell_6t
Xbit_r2_c4 bl[4] br[4] wl[2] vdd gnd cell_6t
Xbit_r3_c4 bl[4] br[4] wl[3] vdd gnd cell_6t
Xbit_r4_c4 bl[4] br[4] wl[4] vdd gnd cell_6t
Xbit_r5_c4 bl[4] br[4] wl[5] vdd gnd cell_6t
Xbit_r6_c4 bl[4] br[4] wl[6] vdd gnd cell_6t
Xbit_r7_c4 bl[4] br[4] wl[7] vdd gnd cell_6t
Xbit_r8_c4 bl[4] br[4] wl[8] vdd gnd cell_6t
Xbit_r9_c4 bl[4] br[4] wl[9] vdd gnd cell_6t
Xbit_r10_c4 bl[4] br[4] wl[10] vdd gnd cell_6t
Xbit_r11_c4 bl[4] br[4] wl[11] vdd gnd cell_6t
Xbit_r12_c4 bl[4] br[4] wl[12] vdd gnd cell_6t
Xbit_r13_c4 bl[4] br[4] wl[13] vdd gnd cell_6t
Xbit_r14_c4 bl[4] br[4] wl[14] vdd gnd cell_6t
Xbit_r15_c4 bl[4] br[4] wl[15] vdd gnd cell_6t
Xbit_r16_c4 bl[4] br[4] wl[16] vdd gnd cell_6t
Xbit_r17_c4 bl[4] br[4] wl[17] vdd gnd cell_6t
Xbit_r18_c4 bl[4] br[4] wl[18] vdd gnd cell_6t
Xbit_r19_c4 bl[4] br[4] wl[19] vdd gnd cell_6t
Xbit_r20_c4 bl[4] br[4] wl[20] vdd gnd cell_6t
Xbit_r21_c4 bl[4] br[4] wl[21] vdd gnd cell_6t
Xbit_r22_c4 bl[4] br[4] wl[22] vdd gnd cell_6t
Xbit_r23_c4 bl[4] br[4] wl[23] vdd gnd cell_6t
Xbit_r24_c4 bl[4] br[4] wl[24] vdd gnd cell_6t
Xbit_r25_c4 bl[4] br[4] wl[25] vdd gnd cell_6t
Xbit_r26_c4 bl[4] br[4] wl[26] vdd gnd cell_6t
Xbit_r27_c4 bl[4] br[4] wl[27] vdd gnd cell_6t
Xbit_r28_c4 bl[4] br[4] wl[28] vdd gnd cell_6t
Xbit_r29_c4 bl[4] br[4] wl[29] vdd gnd cell_6t
Xbit_r30_c4 bl[4] br[4] wl[30] vdd gnd cell_6t
Xbit_r31_c4 bl[4] br[4] wl[31] vdd gnd cell_6t
Xbit_r32_c4 bl[4] br[4] wl[32] vdd gnd cell_6t
Xbit_r33_c4 bl[4] br[4] wl[33] vdd gnd cell_6t
Xbit_r34_c4 bl[4] br[4] wl[34] vdd gnd cell_6t
Xbit_r35_c4 bl[4] br[4] wl[35] vdd gnd cell_6t
Xbit_r36_c4 bl[4] br[4] wl[36] vdd gnd cell_6t
Xbit_r37_c4 bl[4] br[4] wl[37] vdd gnd cell_6t
Xbit_r38_c4 bl[4] br[4] wl[38] vdd gnd cell_6t
Xbit_r39_c4 bl[4] br[4] wl[39] vdd gnd cell_6t
Xbit_r40_c4 bl[4] br[4] wl[40] vdd gnd cell_6t
Xbit_r41_c4 bl[4] br[4] wl[41] vdd gnd cell_6t
Xbit_r42_c4 bl[4] br[4] wl[42] vdd gnd cell_6t
Xbit_r43_c4 bl[4] br[4] wl[43] vdd gnd cell_6t
Xbit_r44_c4 bl[4] br[4] wl[44] vdd gnd cell_6t
Xbit_r45_c4 bl[4] br[4] wl[45] vdd gnd cell_6t
Xbit_r46_c4 bl[4] br[4] wl[46] vdd gnd cell_6t
Xbit_r47_c4 bl[4] br[4] wl[47] vdd gnd cell_6t
Xbit_r48_c4 bl[4] br[4] wl[48] vdd gnd cell_6t
Xbit_r49_c4 bl[4] br[4] wl[49] vdd gnd cell_6t
Xbit_r50_c4 bl[4] br[4] wl[50] vdd gnd cell_6t
Xbit_r51_c4 bl[4] br[4] wl[51] vdd gnd cell_6t
Xbit_r52_c4 bl[4] br[4] wl[52] vdd gnd cell_6t
Xbit_r53_c4 bl[4] br[4] wl[53] vdd gnd cell_6t
Xbit_r54_c4 bl[4] br[4] wl[54] vdd gnd cell_6t
Xbit_r55_c4 bl[4] br[4] wl[55] vdd gnd cell_6t
Xbit_r56_c4 bl[4] br[4] wl[56] vdd gnd cell_6t
Xbit_r57_c4 bl[4] br[4] wl[57] vdd gnd cell_6t
Xbit_r58_c4 bl[4] br[4] wl[58] vdd gnd cell_6t
Xbit_r59_c4 bl[4] br[4] wl[59] vdd gnd cell_6t
Xbit_r60_c4 bl[4] br[4] wl[60] vdd gnd cell_6t
Xbit_r61_c4 bl[4] br[4] wl[61] vdd gnd cell_6t
Xbit_r62_c4 bl[4] br[4] wl[62] vdd gnd cell_6t
Xbit_r63_c4 bl[4] br[4] wl[63] vdd gnd cell_6t
Xbit_r64_c4 bl[4] br[4] wl[64] vdd gnd cell_6t
Xbit_r65_c4 bl[4] br[4] wl[65] vdd gnd cell_6t
Xbit_r66_c4 bl[4] br[4] wl[66] vdd gnd cell_6t
Xbit_r67_c4 bl[4] br[4] wl[67] vdd gnd cell_6t
Xbit_r68_c4 bl[4] br[4] wl[68] vdd gnd cell_6t
Xbit_r69_c4 bl[4] br[4] wl[69] vdd gnd cell_6t
Xbit_r70_c4 bl[4] br[4] wl[70] vdd gnd cell_6t
Xbit_r71_c4 bl[4] br[4] wl[71] vdd gnd cell_6t
Xbit_r72_c4 bl[4] br[4] wl[72] vdd gnd cell_6t
Xbit_r73_c4 bl[4] br[4] wl[73] vdd gnd cell_6t
Xbit_r74_c4 bl[4] br[4] wl[74] vdd gnd cell_6t
Xbit_r75_c4 bl[4] br[4] wl[75] vdd gnd cell_6t
Xbit_r76_c4 bl[4] br[4] wl[76] vdd gnd cell_6t
Xbit_r77_c4 bl[4] br[4] wl[77] vdd gnd cell_6t
Xbit_r78_c4 bl[4] br[4] wl[78] vdd gnd cell_6t
Xbit_r79_c4 bl[4] br[4] wl[79] vdd gnd cell_6t
Xbit_r80_c4 bl[4] br[4] wl[80] vdd gnd cell_6t
Xbit_r81_c4 bl[4] br[4] wl[81] vdd gnd cell_6t
Xbit_r82_c4 bl[4] br[4] wl[82] vdd gnd cell_6t
Xbit_r83_c4 bl[4] br[4] wl[83] vdd gnd cell_6t
Xbit_r84_c4 bl[4] br[4] wl[84] vdd gnd cell_6t
Xbit_r85_c4 bl[4] br[4] wl[85] vdd gnd cell_6t
Xbit_r86_c4 bl[4] br[4] wl[86] vdd gnd cell_6t
Xbit_r87_c4 bl[4] br[4] wl[87] vdd gnd cell_6t
Xbit_r88_c4 bl[4] br[4] wl[88] vdd gnd cell_6t
Xbit_r89_c4 bl[4] br[4] wl[89] vdd gnd cell_6t
Xbit_r90_c4 bl[4] br[4] wl[90] vdd gnd cell_6t
Xbit_r91_c4 bl[4] br[4] wl[91] vdd gnd cell_6t
Xbit_r92_c4 bl[4] br[4] wl[92] vdd gnd cell_6t
Xbit_r93_c4 bl[4] br[4] wl[93] vdd gnd cell_6t
Xbit_r94_c4 bl[4] br[4] wl[94] vdd gnd cell_6t
Xbit_r95_c4 bl[4] br[4] wl[95] vdd gnd cell_6t
Xbit_r96_c4 bl[4] br[4] wl[96] vdd gnd cell_6t
Xbit_r97_c4 bl[4] br[4] wl[97] vdd gnd cell_6t
Xbit_r98_c4 bl[4] br[4] wl[98] vdd gnd cell_6t
Xbit_r99_c4 bl[4] br[4] wl[99] vdd gnd cell_6t
Xbit_r100_c4 bl[4] br[4] wl[100] vdd gnd cell_6t
Xbit_r101_c4 bl[4] br[4] wl[101] vdd gnd cell_6t
Xbit_r102_c4 bl[4] br[4] wl[102] vdd gnd cell_6t
Xbit_r103_c4 bl[4] br[4] wl[103] vdd gnd cell_6t
Xbit_r104_c4 bl[4] br[4] wl[104] vdd gnd cell_6t
Xbit_r105_c4 bl[4] br[4] wl[105] vdd gnd cell_6t
Xbit_r106_c4 bl[4] br[4] wl[106] vdd gnd cell_6t
Xbit_r107_c4 bl[4] br[4] wl[107] vdd gnd cell_6t
Xbit_r108_c4 bl[4] br[4] wl[108] vdd gnd cell_6t
Xbit_r109_c4 bl[4] br[4] wl[109] vdd gnd cell_6t
Xbit_r110_c4 bl[4] br[4] wl[110] vdd gnd cell_6t
Xbit_r111_c4 bl[4] br[4] wl[111] vdd gnd cell_6t
Xbit_r112_c4 bl[4] br[4] wl[112] vdd gnd cell_6t
Xbit_r113_c4 bl[4] br[4] wl[113] vdd gnd cell_6t
Xbit_r114_c4 bl[4] br[4] wl[114] vdd gnd cell_6t
Xbit_r115_c4 bl[4] br[4] wl[115] vdd gnd cell_6t
Xbit_r116_c4 bl[4] br[4] wl[116] vdd gnd cell_6t
Xbit_r117_c4 bl[4] br[4] wl[117] vdd gnd cell_6t
Xbit_r118_c4 bl[4] br[4] wl[118] vdd gnd cell_6t
Xbit_r119_c4 bl[4] br[4] wl[119] vdd gnd cell_6t
Xbit_r120_c4 bl[4] br[4] wl[120] vdd gnd cell_6t
Xbit_r121_c4 bl[4] br[4] wl[121] vdd gnd cell_6t
Xbit_r122_c4 bl[4] br[4] wl[122] vdd gnd cell_6t
Xbit_r123_c4 bl[4] br[4] wl[123] vdd gnd cell_6t
Xbit_r124_c4 bl[4] br[4] wl[124] vdd gnd cell_6t
Xbit_r125_c4 bl[4] br[4] wl[125] vdd gnd cell_6t
Xbit_r126_c4 bl[4] br[4] wl[126] vdd gnd cell_6t
Xbit_r127_c4 bl[4] br[4] wl[127] vdd gnd cell_6t
Xbit_r128_c4 bl[4] br[4] wl[128] vdd gnd cell_6t
Xbit_r129_c4 bl[4] br[4] wl[129] vdd gnd cell_6t
Xbit_r130_c4 bl[4] br[4] wl[130] vdd gnd cell_6t
Xbit_r131_c4 bl[4] br[4] wl[131] vdd gnd cell_6t
Xbit_r132_c4 bl[4] br[4] wl[132] vdd gnd cell_6t
Xbit_r133_c4 bl[4] br[4] wl[133] vdd gnd cell_6t
Xbit_r134_c4 bl[4] br[4] wl[134] vdd gnd cell_6t
Xbit_r135_c4 bl[4] br[4] wl[135] vdd gnd cell_6t
Xbit_r136_c4 bl[4] br[4] wl[136] vdd gnd cell_6t
Xbit_r137_c4 bl[4] br[4] wl[137] vdd gnd cell_6t
Xbit_r138_c4 bl[4] br[4] wl[138] vdd gnd cell_6t
Xbit_r139_c4 bl[4] br[4] wl[139] vdd gnd cell_6t
Xbit_r140_c4 bl[4] br[4] wl[140] vdd gnd cell_6t
Xbit_r141_c4 bl[4] br[4] wl[141] vdd gnd cell_6t
Xbit_r142_c4 bl[4] br[4] wl[142] vdd gnd cell_6t
Xbit_r143_c4 bl[4] br[4] wl[143] vdd gnd cell_6t
Xbit_r144_c4 bl[4] br[4] wl[144] vdd gnd cell_6t
Xbit_r145_c4 bl[4] br[4] wl[145] vdd gnd cell_6t
Xbit_r146_c4 bl[4] br[4] wl[146] vdd gnd cell_6t
Xbit_r147_c4 bl[4] br[4] wl[147] vdd gnd cell_6t
Xbit_r148_c4 bl[4] br[4] wl[148] vdd gnd cell_6t
Xbit_r149_c4 bl[4] br[4] wl[149] vdd gnd cell_6t
Xbit_r150_c4 bl[4] br[4] wl[150] vdd gnd cell_6t
Xbit_r151_c4 bl[4] br[4] wl[151] vdd gnd cell_6t
Xbit_r152_c4 bl[4] br[4] wl[152] vdd gnd cell_6t
Xbit_r153_c4 bl[4] br[4] wl[153] vdd gnd cell_6t
Xbit_r154_c4 bl[4] br[4] wl[154] vdd gnd cell_6t
Xbit_r155_c4 bl[4] br[4] wl[155] vdd gnd cell_6t
Xbit_r156_c4 bl[4] br[4] wl[156] vdd gnd cell_6t
Xbit_r157_c4 bl[4] br[4] wl[157] vdd gnd cell_6t
Xbit_r158_c4 bl[4] br[4] wl[158] vdd gnd cell_6t
Xbit_r159_c4 bl[4] br[4] wl[159] vdd gnd cell_6t
Xbit_r160_c4 bl[4] br[4] wl[160] vdd gnd cell_6t
Xbit_r161_c4 bl[4] br[4] wl[161] vdd gnd cell_6t
Xbit_r162_c4 bl[4] br[4] wl[162] vdd gnd cell_6t
Xbit_r163_c4 bl[4] br[4] wl[163] vdd gnd cell_6t
Xbit_r164_c4 bl[4] br[4] wl[164] vdd gnd cell_6t
Xbit_r165_c4 bl[4] br[4] wl[165] vdd gnd cell_6t
Xbit_r166_c4 bl[4] br[4] wl[166] vdd gnd cell_6t
Xbit_r167_c4 bl[4] br[4] wl[167] vdd gnd cell_6t
Xbit_r168_c4 bl[4] br[4] wl[168] vdd gnd cell_6t
Xbit_r169_c4 bl[4] br[4] wl[169] vdd gnd cell_6t
Xbit_r170_c4 bl[4] br[4] wl[170] vdd gnd cell_6t
Xbit_r171_c4 bl[4] br[4] wl[171] vdd gnd cell_6t
Xbit_r172_c4 bl[4] br[4] wl[172] vdd gnd cell_6t
Xbit_r173_c4 bl[4] br[4] wl[173] vdd gnd cell_6t
Xbit_r174_c4 bl[4] br[4] wl[174] vdd gnd cell_6t
Xbit_r175_c4 bl[4] br[4] wl[175] vdd gnd cell_6t
Xbit_r176_c4 bl[4] br[4] wl[176] vdd gnd cell_6t
Xbit_r177_c4 bl[4] br[4] wl[177] vdd gnd cell_6t
Xbit_r178_c4 bl[4] br[4] wl[178] vdd gnd cell_6t
Xbit_r179_c4 bl[4] br[4] wl[179] vdd gnd cell_6t
Xbit_r180_c4 bl[4] br[4] wl[180] vdd gnd cell_6t
Xbit_r181_c4 bl[4] br[4] wl[181] vdd gnd cell_6t
Xbit_r182_c4 bl[4] br[4] wl[182] vdd gnd cell_6t
Xbit_r183_c4 bl[4] br[4] wl[183] vdd gnd cell_6t
Xbit_r184_c4 bl[4] br[4] wl[184] vdd gnd cell_6t
Xbit_r185_c4 bl[4] br[4] wl[185] vdd gnd cell_6t
Xbit_r186_c4 bl[4] br[4] wl[186] vdd gnd cell_6t
Xbit_r187_c4 bl[4] br[4] wl[187] vdd gnd cell_6t
Xbit_r188_c4 bl[4] br[4] wl[188] vdd gnd cell_6t
Xbit_r189_c4 bl[4] br[4] wl[189] vdd gnd cell_6t
Xbit_r190_c4 bl[4] br[4] wl[190] vdd gnd cell_6t
Xbit_r191_c4 bl[4] br[4] wl[191] vdd gnd cell_6t
Xbit_r192_c4 bl[4] br[4] wl[192] vdd gnd cell_6t
Xbit_r193_c4 bl[4] br[4] wl[193] vdd gnd cell_6t
Xbit_r194_c4 bl[4] br[4] wl[194] vdd gnd cell_6t
Xbit_r195_c4 bl[4] br[4] wl[195] vdd gnd cell_6t
Xbit_r196_c4 bl[4] br[4] wl[196] vdd gnd cell_6t
Xbit_r197_c4 bl[4] br[4] wl[197] vdd gnd cell_6t
Xbit_r198_c4 bl[4] br[4] wl[198] vdd gnd cell_6t
Xbit_r199_c4 bl[4] br[4] wl[199] vdd gnd cell_6t
Xbit_r200_c4 bl[4] br[4] wl[200] vdd gnd cell_6t
Xbit_r201_c4 bl[4] br[4] wl[201] vdd gnd cell_6t
Xbit_r202_c4 bl[4] br[4] wl[202] vdd gnd cell_6t
Xbit_r203_c4 bl[4] br[4] wl[203] vdd gnd cell_6t
Xbit_r204_c4 bl[4] br[4] wl[204] vdd gnd cell_6t
Xbit_r205_c4 bl[4] br[4] wl[205] vdd gnd cell_6t
Xbit_r206_c4 bl[4] br[4] wl[206] vdd gnd cell_6t
Xbit_r207_c4 bl[4] br[4] wl[207] vdd gnd cell_6t
Xbit_r208_c4 bl[4] br[4] wl[208] vdd gnd cell_6t
Xbit_r209_c4 bl[4] br[4] wl[209] vdd gnd cell_6t
Xbit_r210_c4 bl[4] br[4] wl[210] vdd gnd cell_6t
Xbit_r211_c4 bl[4] br[4] wl[211] vdd gnd cell_6t
Xbit_r212_c4 bl[4] br[4] wl[212] vdd gnd cell_6t
Xbit_r213_c4 bl[4] br[4] wl[213] vdd gnd cell_6t
Xbit_r214_c4 bl[4] br[4] wl[214] vdd gnd cell_6t
Xbit_r215_c4 bl[4] br[4] wl[215] vdd gnd cell_6t
Xbit_r216_c4 bl[4] br[4] wl[216] vdd gnd cell_6t
Xbit_r217_c4 bl[4] br[4] wl[217] vdd gnd cell_6t
Xbit_r218_c4 bl[4] br[4] wl[218] vdd gnd cell_6t
Xbit_r219_c4 bl[4] br[4] wl[219] vdd gnd cell_6t
Xbit_r220_c4 bl[4] br[4] wl[220] vdd gnd cell_6t
Xbit_r221_c4 bl[4] br[4] wl[221] vdd gnd cell_6t
Xbit_r222_c4 bl[4] br[4] wl[222] vdd gnd cell_6t
Xbit_r223_c4 bl[4] br[4] wl[223] vdd gnd cell_6t
Xbit_r224_c4 bl[4] br[4] wl[224] vdd gnd cell_6t
Xbit_r225_c4 bl[4] br[4] wl[225] vdd gnd cell_6t
Xbit_r226_c4 bl[4] br[4] wl[226] vdd gnd cell_6t
Xbit_r227_c4 bl[4] br[4] wl[227] vdd gnd cell_6t
Xbit_r228_c4 bl[4] br[4] wl[228] vdd gnd cell_6t
Xbit_r229_c4 bl[4] br[4] wl[229] vdd gnd cell_6t
Xbit_r230_c4 bl[4] br[4] wl[230] vdd gnd cell_6t
Xbit_r231_c4 bl[4] br[4] wl[231] vdd gnd cell_6t
Xbit_r232_c4 bl[4] br[4] wl[232] vdd gnd cell_6t
Xbit_r233_c4 bl[4] br[4] wl[233] vdd gnd cell_6t
Xbit_r234_c4 bl[4] br[4] wl[234] vdd gnd cell_6t
Xbit_r235_c4 bl[4] br[4] wl[235] vdd gnd cell_6t
Xbit_r236_c4 bl[4] br[4] wl[236] vdd gnd cell_6t
Xbit_r237_c4 bl[4] br[4] wl[237] vdd gnd cell_6t
Xbit_r238_c4 bl[4] br[4] wl[238] vdd gnd cell_6t
Xbit_r239_c4 bl[4] br[4] wl[239] vdd gnd cell_6t
Xbit_r240_c4 bl[4] br[4] wl[240] vdd gnd cell_6t
Xbit_r241_c4 bl[4] br[4] wl[241] vdd gnd cell_6t
Xbit_r242_c4 bl[4] br[4] wl[242] vdd gnd cell_6t
Xbit_r243_c4 bl[4] br[4] wl[243] vdd gnd cell_6t
Xbit_r244_c4 bl[4] br[4] wl[244] vdd gnd cell_6t
Xbit_r245_c4 bl[4] br[4] wl[245] vdd gnd cell_6t
Xbit_r246_c4 bl[4] br[4] wl[246] vdd gnd cell_6t
Xbit_r247_c4 bl[4] br[4] wl[247] vdd gnd cell_6t
Xbit_r248_c4 bl[4] br[4] wl[248] vdd gnd cell_6t
Xbit_r249_c4 bl[4] br[4] wl[249] vdd gnd cell_6t
Xbit_r250_c4 bl[4] br[4] wl[250] vdd gnd cell_6t
Xbit_r251_c4 bl[4] br[4] wl[251] vdd gnd cell_6t
Xbit_r252_c4 bl[4] br[4] wl[252] vdd gnd cell_6t
Xbit_r253_c4 bl[4] br[4] wl[253] vdd gnd cell_6t
Xbit_r254_c4 bl[4] br[4] wl[254] vdd gnd cell_6t
Xbit_r255_c4 bl[4] br[4] wl[255] vdd gnd cell_6t
Xbit_r256_c4 bl[4] br[4] wl[256] vdd gnd cell_6t
Xbit_r257_c4 bl[4] br[4] wl[257] vdd gnd cell_6t
Xbit_r258_c4 bl[4] br[4] wl[258] vdd gnd cell_6t
Xbit_r259_c4 bl[4] br[4] wl[259] vdd gnd cell_6t
Xbit_r260_c4 bl[4] br[4] wl[260] vdd gnd cell_6t
Xbit_r261_c4 bl[4] br[4] wl[261] vdd gnd cell_6t
Xbit_r262_c4 bl[4] br[4] wl[262] vdd gnd cell_6t
Xbit_r263_c4 bl[4] br[4] wl[263] vdd gnd cell_6t
Xbit_r264_c4 bl[4] br[4] wl[264] vdd gnd cell_6t
Xbit_r265_c4 bl[4] br[4] wl[265] vdd gnd cell_6t
Xbit_r266_c4 bl[4] br[4] wl[266] vdd gnd cell_6t
Xbit_r267_c4 bl[4] br[4] wl[267] vdd gnd cell_6t
Xbit_r268_c4 bl[4] br[4] wl[268] vdd gnd cell_6t
Xbit_r269_c4 bl[4] br[4] wl[269] vdd gnd cell_6t
Xbit_r270_c4 bl[4] br[4] wl[270] vdd gnd cell_6t
Xbit_r271_c4 bl[4] br[4] wl[271] vdd gnd cell_6t
Xbit_r272_c4 bl[4] br[4] wl[272] vdd gnd cell_6t
Xbit_r273_c4 bl[4] br[4] wl[273] vdd gnd cell_6t
Xbit_r274_c4 bl[4] br[4] wl[274] vdd gnd cell_6t
Xbit_r275_c4 bl[4] br[4] wl[275] vdd gnd cell_6t
Xbit_r276_c4 bl[4] br[4] wl[276] vdd gnd cell_6t
Xbit_r277_c4 bl[4] br[4] wl[277] vdd gnd cell_6t
Xbit_r278_c4 bl[4] br[4] wl[278] vdd gnd cell_6t
Xbit_r279_c4 bl[4] br[4] wl[279] vdd gnd cell_6t
Xbit_r280_c4 bl[4] br[4] wl[280] vdd gnd cell_6t
Xbit_r281_c4 bl[4] br[4] wl[281] vdd gnd cell_6t
Xbit_r282_c4 bl[4] br[4] wl[282] vdd gnd cell_6t
Xbit_r283_c4 bl[4] br[4] wl[283] vdd gnd cell_6t
Xbit_r284_c4 bl[4] br[4] wl[284] vdd gnd cell_6t
Xbit_r285_c4 bl[4] br[4] wl[285] vdd gnd cell_6t
Xbit_r286_c4 bl[4] br[4] wl[286] vdd gnd cell_6t
Xbit_r287_c4 bl[4] br[4] wl[287] vdd gnd cell_6t
Xbit_r288_c4 bl[4] br[4] wl[288] vdd gnd cell_6t
Xbit_r289_c4 bl[4] br[4] wl[289] vdd gnd cell_6t
Xbit_r290_c4 bl[4] br[4] wl[290] vdd gnd cell_6t
Xbit_r291_c4 bl[4] br[4] wl[291] vdd gnd cell_6t
Xbit_r292_c4 bl[4] br[4] wl[292] vdd gnd cell_6t
Xbit_r293_c4 bl[4] br[4] wl[293] vdd gnd cell_6t
Xbit_r294_c4 bl[4] br[4] wl[294] vdd gnd cell_6t
Xbit_r295_c4 bl[4] br[4] wl[295] vdd gnd cell_6t
Xbit_r296_c4 bl[4] br[4] wl[296] vdd gnd cell_6t
Xbit_r297_c4 bl[4] br[4] wl[297] vdd gnd cell_6t
Xbit_r298_c4 bl[4] br[4] wl[298] vdd gnd cell_6t
Xbit_r299_c4 bl[4] br[4] wl[299] vdd gnd cell_6t
Xbit_r300_c4 bl[4] br[4] wl[300] vdd gnd cell_6t
Xbit_r301_c4 bl[4] br[4] wl[301] vdd gnd cell_6t
Xbit_r302_c4 bl[4] br[4] wl[302] vdd gnd cell_6t
Xbit_r303_c4 bl[4] br[4] wl[303] vdd gnd cell_6t
Xbit_r304_c4 bl[4] br[4] wl[304] vdd gnd cell_6t
Xbit_r305_c4 bl[4] br[4] wl[305] vdd gnd cell_6t
Xbit_r306_c4 bl[4] br[4] wl[306] vdd gnd cell_6t
Xbit_r307_c4 bl[4] br[4] wl[307] vdd gnd cell_6t
Xbit_r308_c4 bl[4] br[4] wl[308] vdd gnd cell_6t
Xbit_r309_c4 bl[4] br[4] wl[309] vdd gnd cell_6t
Xbit_r310_c4 bl[4] br[4] wl[310] vdd gnd cell_6t
Xbit_r311_c4 bl[4] br[4] wl[311] vdd gnd cell_6t
Xbit_r312_c4 bl[4] br[4] wl[312] vdd gnd cell_6t
Xbit_r313_c4 bl[4] br[4] wl[313] vdd gnd cell_6t
Xbit_r314_c4 bl[4] br[4] wl[314] vdd gnd cell_6t
Xbit_r315_c4 bl[4] br[4] wl[315] vdd gnd cell_6t
Xbit_r316_c4 bl[4] br[4] wl[316] vdd gnd cell_6t
Xbit_r317_c4 bl[4] br[4] wl[317] vdd gnd cell_6t
Xbit_r318_c4 bl[4] br[4] wl[318] vdd gnd cell_6t
Xbit_r319_c4 bl[4] br[4] wl[319] vdd gnd cell_6t
Xbit_r320_c4 bl[4] br[4] wl[320] vdd gnd cell_6t
Xbit_r321_c4 bl[4] br[4] wl[321] vdd gnd cell_6t
Xbit_r322_c4 bl[4] br[4] wl[322] vdd gnd cell_6t
Xbit_r323_c4 bl[4] br[4] wl[323] vdd gnd cell_6t
Xbit_r324_c4 bl[4] br[4] wl[324] vdd gnd cell_6t
Xbit_r325_c4 bl[4] br[4] wl[325] vdd gnd cell_6t
Xbit_r326_c4 bl[4] br[4] wl[326] vdd gnd cell_6t
Xbit_r327_c4 bl[4] br[4] wl[327] vdd gnd cell_6t
Xbit_r328_c4 bl[4] br[4] wl[328] vdd gnd cell_6t
Xbit_r329_c4 bl[4] br[4] wl[329] vdd gnd cell_6t
Xbit_r330_c4 bl[4] br[4] wl[330] vdd gnd cell_6t
Xbit_r331_c4 bl[4] br[4] wl[331] vdd gnd cell_6t
Xbit_r332_c4 bl[4] br[4] wl[332] vdd gnd cell_6t
Xbit_r333_c4 bl[4] br[4] wl[333] vdd gnd cell_6t
Xbit_r334_c4 bl[4] br[4] wl[334] vdd gnd cell_6t
Xbit_r335_c4 bl[4] br[4] wl[335] vdd gnd cell_6t
Xbit_r336_c4 bl[4] br[4] wl[336] vdd gnd cell_6t
Xbit_r337_c4 bl[4] br[4] wl[337] vdd gnd cell_6t
Xbit_r338_c4 bl[4] br[4] wl[338] vdd gnd cell_6t
Xbit_r339_c4 bl[4] br[4] wl[339] vdd gnd cell_6t
Xbit_r340_c4 bl[4] br[4] wl[340] vdd gnd cell_6t
Xbit_r341_c4 bl[4] br[4] wl[341] vdd gnd cell_6t
Xbit_r342_c4 bl[4] br[4] wl[342] vdd gnd cell_6t
Xbit_r343_c4 bl[4] br[4] wl[343] vdd gnd cell_6t
Xbit_r344_c4 bl[4] br[4] wl[344] vdd gnd cell_6t
Xbit_r345_c4 bl[4] br[4] wl[345] vdd gnd cell_6t
Xbit_r346_c4 bl[4] br[4] wl[346] vdd gnd cell_6t
Xbit_r347_c4 bl[4] br[4] wl[347] vdd gnd cell_6t
Xbit_r348_c4 bl[4] br[4] wl[348] vdd gnd cell_6t
Xbit_r349_c4 bl[4] br[4] wl[349] vdd gnd cell_6t
Xbit_r350_c4 bl[4] br[4] wl[350] vdd gnd cell_6t
Xbit_r351_c4 bl[4] br[4] wl[351] vdd gnd cell_6t
Xbit_r352_c4 bl[4] br[4] wl[352] vdd gnd cell_6t
Xbit_r353_c4 bl[4] br[4] wl[353] vdd gnd cell_6t
Xbit_r354_c4 bl[4] br[4] wl[354] vdd gnd cell_6t
Xbit_r355_c4 bl[4] br[4] wl[355] vdd gnd cell_6t
Xbit_r356_c4 bl[4] br[4] wl[356] vdd gnd cell_6t
Xbit_r357_c4 bl[4] br[4] wl[357] vdd gnd cell_6t
Xbit_r358_c4 bl[4] br[4] wl[358] vdd gnd cell_6t
Xbit_r359_c4 bl[4] br[4] wl[359] vdd gnd cell_6t
Xbit_r360_c4 bl[4] br[4] wl[360] vdd gnd cell_6t
Xbit_r361_c4 bl[4] br[4] wl[361] vdd gnd cell_6t
Xbit_r362_c4 bl[4] br[4] wl[362] vdd gnd cell_6t
Xbit_r363_c4 bl[4] br[4] wl[363] vdd gnd cell_6t
Xbit_r364_c4 bl[4] br[4] wl[364] vdd gnd cell_6t
Xbit_r365_c4 bl[4] br[4] wl[365] vdd gnd cell_6t
Xbit_r366_c4 bl[4] br[4] wl[366] vdd gnd cell_6t
Xbit_r367_c4 bl[4] br[4] wl[367] vdd gnd cell_6t
Xbit_r368_c4 bl[4] br[4] wl[368] vdd gnd cell_6t
Xbit_r369_c4 bl[4] br[4] wl[369] vdd gnd cell_6t
Xbit_r370_c4 bl[4] br[4] wl[370] vdd gnd cell_6t
Xbit_r371_c4 bl[4] br[4] wl[371] vdd gnd cell_6t
Xbit_r372_c4 bl[4] br[4] wl[372] vdd gnd cell_6t
Xbit_r373_c4 bl[4] br[4] wl[373] vdd gnd cell_6t
Xbit_r374_c4 bl[4] br[4] wl[374] vdd gnd cell_6t
Xbit_r375_c4 bl[4] br[4] wl[375] vdd gnd cell_6t
Xbit_r376_c4 bl[4] br[4] wl[376] vdd gnd cell_6t
Xbit_r377_c4 bl[4] br[4] wl[377] vdd gnd cell_6t
Xbit_r378_c4 bl[4] br[4] wl[378] vdd gnd cell_6t
Xbit_r379_c4 bl[4] br[4] wl[379] vdd gnd cell_6t
Xbit_r380_c4 bl[4] br[4] wl[380] vdd gnd cell_6t
Xbit_r381_c4 bl[4] br[4] wl[381] vdd gnd cell_6t
Xbit_r382_c4 bl[4] br[4] wl[382] vdd gnd cell_6t
Xbit_r383_c4 bl[4] br[4] wl[383] vdd gnd cell_6t
Xbit_r384_c4 bl[4] br[4] wl[384] vdd gnd cell_6t
Xbit_r385_c4 bl[4] br[4] wl[385] vdd gnd cell_6t
Xbit_r386_c4 bl[4] br[4] wl[386] vdd gnd cell_6t
Xbit_r387_c4 bl[4] br[4] wl[387] vdd gnd cell_6t
Xbit_r388_c4 bl[4] br[4] wl[388] vdd gnd cell_6t
Xbit_r389_c4 bl[4] br[4] wl[389] vdd gnd cell_6t
Xbit_r390_c4 bl[4] br[4] wl[390] vdd gnd cell_6t
Xbit_r391_c4 bl[4] br[4] wl[391] vdd gnd cell_6t
Xbit_r392_c4 bl[4] br[4] wl[392] vdd gnd cell_6t
Xbit_r393_c4 bl[4] br[4] wl[393] vdd gnd cell_6t
Xbit_r394_c4 bl[4] br[4] wl[394] vdd gnd cell_6t
Xbit_r395_c4 bl[4] br[4] wl[395] vdd gnd cell_6t
Xbit_r396_c4 bl[4] br[4] wl[396] vdd gnd cell_6t
Xbit_r397_c4 bl[4] br[4] wl[397] vdd gnd cell_6t
Xbit_r398_c4 bl[4] br[4] wl[398] vdd gnd cell_6t
Xbit_r399_c4 bl[4] br[4] wl[399] vdd gnd cell_6t
Xbit_r400_c4 bl[4] br[4] wl[400] vdd gnd cell_6t
Xbit_r401_c4 bl[4] br[4] wl[401] vdd gnd cell_6t
Xbit_r402_c4 bl[4] br[4] wl[402] vdd gnd cell_6t
Xbit_r403_c4 bl[4] br[4] wl[403] vdd gnd cell_6t
Xbit_r404_c4 bl[4] br[4] wl[404] vdd gnd cell_6t
Xbit_r405_c4 bl[4] br[4] wl[405] vdd gnd cell_6t
Xbit_r406_c4 bl[4] br[4] wl[406] vdd gnd cell_6t
Xbit_r407_c4 bl[4] br[4] wl[407] vdd gnd cell_6t
Xbit_r408_c4 bl[4] br[4] wl[408] vdd gnd cell_6t
Xbit_r409_c4 bl[4] br[4] wl[409] vdd gnd cell_6t
Xbit_r410_c4 bl[4] br[4] wl[410] vdd gnd cell_6t
Xbit_r411_c4 bl[4] br[4] wl[411] vdd gnd cell_6t
Xbit_r412_c4 bl[4] br[4] wl[412] vdd gnd cell_6t
Xbit_r413_c4 bl[4] br[4] wl[413] vdd gnd cell_6t
Xbit_r414_c4 bl[4] br[4] wl[414] vdd gnd cell_6t
Xbit_r415_c4 bl[4] br[4] wl[415] vdd gnd cell_6t
Xbit_r416_c4 bl[4] br[4] wl[416] vdd gnd cell_6t
Xbit_r417_c4 bl[4] br[4] wl[417] vdd gnd cell_6t
Xbit_r418_c4 bl[4] br[4] wl[418] vdd gnd cell_6t
Xbit_r419_c4 bl[4] br[4] wl[419] vdd gnd cell_6t
Xbit_r420_c4 bl[4] br[4] wl[420] vdd gnd cell_6t
Xbit_r421_c4 bl[4] br[4] wl[421] vdd gnd cell_6t
Xbit_r422_c4 bl[4] br[4] wl[422] vdd gnd cell_6t
Xbit_r423_c4 bl[4] br[4] wl[423] vdd gnd cell_6t
Xbit_r424_c4 bl[4] br[4] wl[424] vdd gnd cell_6t
Xbit_r425_c4 bl[4] br[4] wl[425] vdd gnd cell_6t
Xbit_r426_c4 bl[4] br[4] wl[426] vdd gnd cell_6t
Xbit_r427_c4 bl[4] br[4] wl[427] vdd gnd cell_6t
Xbit_r428_c4 bl[4] br[4] wl[428] vdd gnd cell_6t
Xbit_r429_c4 bl[4] br[4] wl[429] vdd gnd cell_6t
Xbit_r430_c4 bl[4] br[4] wl[430] vdd gnd cell_6t
Xbit_r431_c4 bl[4] br[4] wl[431] vdd gnd cell_6t
Xbit_r432_c4 bl[4] br[4] wl[432] vdd gnd cell_6t
Xbit_r433_c4 bl[4] br[4] wl[433] vdd gnd cell_6t
Xbit_r434_c4 bl[4] br[4] wl[434] vdd gnd cell_6t
Xbit_r435_c4 bl[4] br[4] wl[435] vdd gnd cell_6t
Xbit_r436_c4 bl[4] br[4] wl[436] vdd gnd cell_6t
Xbit_r437_c4 bl[4] br[4] wl[437] vdd gnd cell_6t
Xbit_r438_c4 bl[4] br[4] wl[438] vdd gnd cell_6t
Xbit_r439_c4 bl[4] br[4] wl[439] vdd gnd cell_6t
Xbit_r440_c4 bl[4] br[4] wl[440] vdd gnd cell_6t
Xbit_r441_c4 bl[4] br[4] wl[441] vdd gnd cell_6t
Xbit_r442_c4 bl[4] br[4] wl[442] vdd gnd cell_6t
Xbit_r443_c4 bl[4] br[4] wl[443] vdd gnd cell_6t
Xbit_r444_c4 bl[4] br[4] wl[444] vdd gnd cell_6t
Xbit_r445_c4 bl[4] br[4] wl[445] vdd gnd cell_6t
Xbit_r446_c4 bl[4] br[4] wl[446] vdd gnd cell_6t
Xbit_r447_c4 bl[4] br[4] wl[447] vdd gnd cell_6t
Xbit_r448_c4 bl[4] br[4] wl[448] vdd gnd cell_6t
Xbit_r449_c4 bl[4] br[4] wl[449] vdd gnd cell_6t
Xbit_r450_c4 bl[4] br[4] wl[450] vdd gnd cell_6t
Xbit_r451_c4 bl[4] br[4] wl[451] vdd gnd cell_6t
Xbit_r452_c4 bl[4] br[4] wl[452] vdd gnd cell_6t
Xbit_r453_c4 bl[4] br[4] wl[453] vdd gnd cell_6t
Xbit_r454_c4 bl[4] br[4] wl[454] vdd gnd cell_6t
Xbit_r455_c4 bl[4] br[4] wl[455] vdd gnd cell_6t
Xbit_r456_c4 bl[4] br[4] wl[456] vdd gnd cell_6t
Xbit_r457_c4 bl[4] br[4] wl[457] vdd gnd cell_6t
Xbit_r458_c4 bl[4] br[4] wl[458] vdd gnd cell_6t
Xbit_r459_c4 bl[4] br[4] wl[459] vdd gnd cell_6t
Xbit_r460_c4 bl[4] br[4] wl[460] vdd gnd cell_6t
Xbit_r461_c4 bl[4] br[4] wl[461] vdd gnd cell_6t
Xbit_r462_c4 bl[4] br[4] wl[462] vdd gnd cell_6t
Xbit_r463_c4 bl[4] br[4] wl[463] vdd gnd cell_6t
Xbit_r464_c4 bl[4] br[4] wl[464] vdd gnd cell_6t
Xbit_r465_c4 bl[4] br[4] wl[465] vdd gnd cell_6t
Xbit_r466_c4 bl[4] br[4] wl[466] vdd gnd cell_6t
Xbit_r467_c4 bl[4] br[4] wl[467] vdd gnd cell_6t
Xbit_r468_c4 bl[4] br[4] wl[468] vdd gnd cell_6t
Xbit_r469_c4 bl[4] br[4] wl[469] vdd gnd cell_6t
Xbit_r470_c4 bl[4] br[4] wl[470] vdd gnd cell_6t
Xbit_r471_c4 bl[4] br[4] wl[471] vdd gnd cell_6t
Xbit_r472_c4 bl[4] br[4] wl[472] vdd gnd cell_6t
Xbit_r473_c4 bl[4] br[4] wl[473] vdd gnd cell_6t
Xbit_r474_c4 bl[4] br[4] wl[474] vdd gnd cell_6t
Xbit_r475_c4 bl[4] br[4] wl[475] vdd gnd cell_6t
Xbit_r476_c4 bl[4] br[4] wl[476] vdd gnd cell_6t
Xbit_r477_c4 bl[4] br[4] wl[477] vdd gnd cell_6t
Xbit_r478_c4 bl[4] br[4] wl[478] vdd gnd cell_6t
Xbit_r479_c4 bl[4] br[4] wl[479] vdd gnd cell_6t
Xbit_r480_c4 bl[4] br[4] wl[480] vdd gnd cell_6t
Xbit_r481_c4 bl[4] br[4] wl[481] vdd gnd cell_6t
Xbit_r482_c4 bl[4] br[4] wl[482] vdd gnd cell_6t
Xbit_r483_c4 bl[4] br[4] wl[483] vdd gnd cell_6t
Xbit_r484_c4 bl[4] br[4] wl[484] vdd gnd cell_6t
Xbit_r485_c4 bl[4] br[4] wl[485] vdd gnd cell_6t
Xbit_r486_c4 bl[4] br[4] wl[486] vdd gnd cell_6t
Xbit_r487_c4 bl[4] br[4] wl[487] vdd gnd cell_6t
Xbit_r488_c4 bl[4] br[4] wl[488] vdd gnd cell_6t
Xbit_r489_c4 bl[4] br[4] wl[489] vdd gnd cell_6t
Xbit_r490_c4 bl[4] br[4] wl[490] vdd gnd cell_6t
Xbit_r491_c4 bl[4] br[4] wl[491] vdd gnd cell_6t
Xbit_r492_c4 bl[4] br[4] wl[492] vdd gnd cell_6t
Xbit_r493_c4 bl[4] br[4] wl[493] vdd gnd cell_6t
Xbit_r494_c4 bl[4] br[4] wl[494] vdd gnd cell_6t
Xbit_r495_c4 bl[4] br[4] wl[495] vdd gnd cell_6t
Xbit_r496_c4 bl[4] br[4] wl[496] vdd gnd cell_6t
Xbit_r497_c4 bl[4] br[4] wl[497] vdd gnd cell_6t
Xbit_r498_c4 bl[4] br[4] wl[498] vdd gnd cell_6t
Xbit_r499_c4 bl[4] br[4] wl[499] vdd gnd cell_6t
Xbit_r500_c4 bl[4] br[4] wl[500] vdd gnd cell_6t
Xbit_r501_c4 bl[4] br[4] wl[501] vdd gnd cell_6t
Xbit_r502_c4 bl[4] br[4] wl[502] vdd gnd cell_6t
Xbit_r503_c4 bl[4] br[4] wl[503] vdd gnd cell_6t
Xbit_r504_c4 bl[4] br[4] wl[504] vdd gnd cell_6t
Xbit_r505_c4 bl[4] br[4] wl[505] vdd gnd cell_6t
Xbit_r506_c4 bl[4] br[4] wl[506] vdd gnd cell_6t
Xbit_r507_c4 bl[4] br[4] wl[507] vdd gnd cell_6t
Xbit_r508_c4 bl[4] br[4] wl[508] vdd gnd cell_6t
Xbit_r509_c4 bl[4] br[4] wl[509] vdd gnd cell_6t
Xbit_r510_c4 bl[4] br[4] wl[510] vdd gnd cell_6t
Xbit_r511_c4 bl[4] br[4] wl[511] vdd gnd cell_6t
Xbit_r0_c5 bl[5] br[5] wl[0] vdd gnd cell_6t
Xbit_r1_c5 bl[5] br[5] wl[1] vdd gnd cell_6t
Xbit_r2_c5 bl[5] br[5] wl[2] vdd gnd cell_6t
Xbit_r3_c5 bl[5] br[5] wl[3] vdd gnd cell_6t
Xbit_r4_c5 bl[5] br[5] wl[4] vdd gnd cell_6t
Xbit_r5_c5 bl[5] br[5] wl[5] vdd gnd cell_6t
Xbit_r6_c5 bl[5] br[5] wl[6] vdd gnd cell_6t
Xbit_r7_c5 bl[5] br[5] wl[7] vdd gnd cell_6t
Xbit_r8_c5 bl[5] br[5] wl[8] vdd gnd cell_6t
Xbit_r9_c5 bl[5] br[5] wl[9] vdd gnd cell_6t
Xbit_r10_c5 bl[5] br[5] wl[10] vdd gnd cell_6t
Xbit_r11_c5 bl[5] br[5] wl[11] vdd gnd cell_6t
Xbit_r12_c5 bl[5] br[5] wl[12] vdd gnd cell_6t
Xbit_r13_c5 bl[5] br[5] wl[13] vdd gnd cell_6t
Xbit_r14_c5 bl[5] br[5] wl[14] vdd gnd cell_6t
Xbit_r15_c5 bl[5] br[5] wl[15] vdd gnd cell_6t
Xbit_r16_c5 bl[5] br[5] wl[16] vdd gnd cell_6t
Xbit_r17_c5 bl[5] br[5] wl[17] vdd gnd cell_6t
Xbit_r18_c5 bl[5] br[5] wl[18] vdd gnd cell_6t
Xbit_r19_c5 bl[5] br[5] wl[19] vdd gnd cell_6t
Xbit_r20_c5 bl[5] br[5] wl[20] vdd gnd cell_6t
Xbit_r21_c5 bl[5] br[5] wl[21] vdd gnd cell_6t
Xbit_r22_c5 bl[5] br[5] wl[22] vdd gnd cell_6t
Xbit_r23_c5 bl[5] br[5] wl[23] vdd gnd cell_6t
Xbit_r24_c5 bl[5] br[5] wl[24] vdd gnd cell_6t
Xbit_r25_c5 bl[5] br[5] wl[25] vdd gnd cell_6t
Xbit_r26_c5 bl[5] br[5] wl[26] vdd gnd cell_6t
Xbit_r27_c5 bl[5] br[5] wl[27] vdd gnd cell_6t
Xbit_r28_c5 bl[5] br[5] wl[28] vdd gnd cell_6t
Xbit_r29_c5 bl[5] br[5] wl[29] vdd gnd cell_6t
Xbit_r30_c5 bl[5] br[5] wl[30] vdd gnd cell_6t
Xbit_r31_c5 bl[5] br[5] wl[31] vdd gnd cell_6t
Xbit_r32_c5 bl[5] br[5] wl[32] vdd gnd cell_6t
Xbit_r33_c5 bl[5] br[5] wl[33] vdd gnd cell_6t
Xbit_r34_c5 bl[5] br[5] wl[34] vdd gnd cell_6t
Xbit_r35_c5 bl[5] br[5] wl[35] vdd gnd cell_6t
Xbit_r36_c5 bl[5] br[5] wl[36] vdd gnd cell_6t
Xbit_r37_c5 bl[5] br[5] wl[37] vdd gnd cell_6t
Xbit_r38_c5 bl[5] br[5] wl[38] vdd gnd cell_6t
Xbit_r39_c5 bl[5] br[5] wl[39] vdd gnd cell_6t
Xbit_r40_c5 bl[5] br[5] wl[40] vdd gnd cell_6t
Xbit_r41_c5 bl[5] br[5] wl[41] vdd gnd cell_6t
Xbit_r42_c5 bl[5] br[5] wl[42] vdd gnd cell_6t
Xbit_r43_c5 bl[5] br[5] wl[43] vdd gnd cell_6t
Xbit_r44_c5 bl[5] br[5] wl[44] vdd gnd cell_6t
Xbit_r45_c5 bl[5] br[5] wl[45] vdd gnd cell_6t
Xbit_r46_c5 bl[5] br[5] wl[46] vdd gnd cell_6t
Xbit_r47_c5 bl[5] br[5] wl[47] vdd gnd cell_6t
Xbit_r48_c5 bl[5] br[5] wl[48] vdd gnd cell_6t
Xbit_r49_c5 bl[5] br[5] wl[49] vdd gnd cell_6t
Xbit_r50_c5 bl[5] br[5] wl[50] vdd gnd cell_6t
Xbit_r51_c5 bl[5] br[5] wl[51] vdd gnd cell_6t
Xbit_r52_c5 bl[5] br[5] wl[52] vdd gnd cell_6t
Xbit_r53_c5 bl[5] br[5] wl[53] vdd gnd cell_6t
Xbit_r54_c5 bl[5] br[5] wl[54] vdd gnd cell_6t
Xbit_r55_c5 bl[5] br[5] wl[55] vdd gnd cell_6t
Xbit_r56_c5 bl[5] br[5] wl[56] vdd gnd cell_6t
Xbit_r57_c5 bl[5] br[5] wl[57] vdd gnd cell_6t
Xbit_r58_c5 bl[5] br[5] wl[58] vdd gnd cell_6t
Xbit_r59_c5 bl[5] br[5] wl[59] vdd gnd cell_6t
Xbit_r60_c5 bl[5] br[5] wl[60] vdd gnd cell_6t
Xbit_r61_c5 bl[5] br[5] wl[61] vdd gnd cell_6t
Xbit_r62_c5 bl[5] br[5] wl[62] vdd gnd cell_6t
Xbit_r63_c5 bl[5] br[5] wl[63] vdd gnd cell_6t
Xbit_r64_c5 bl[5] br[5] wl[64] vdd gnd cell_6t
Xbit_r65_c5 bl[5] br[5] wl[65] vdd gnd cell_6t
Xbit_r66_c5 bl[5] br[5] wl[66] vdd gnd cell_6t
Xbit_r67_c5 bl[5] br[5] wl[67] vdd gnd cell_6t
Xbit_r68_c5 bl[5] br[5] wl[68] vdd gnd cell_6t
Xbit_r69_c5 bl[5] br[5] wl[69] vdd gnd cell_6t
Xbit_r70_c5 bl[5] br[5] wl[70] vdd gnd cell_6t
Xbit_r71_c5 bl[5] br[5] wl[71] vdd gnd cell_6t
Xbit_r72_c5 bl[5] br[5] wl[72] vdd gnd cell_6t
Xbit_r73_c5 bl[5] br[5] wl[73] vdd gnd cell_6t
Xbit_r74_c5 bl[5] br[5] wl[74] vdd gnd cell_6t
Xbit_r75_c5 bl[5] br[5] wl[75] vdd gnd cell_6t
Xbit_r76_c5 bl[5] br[5] wl[76] vdd gnd cell_6t
Xbit_r77_c5 bl[5] br[5] wl[77] vdd gnd cell_6t
Xbit_r78_c5 bl[5] br[5] wl[78] vdd gnd cell_6t
Xbit_r79_c5 bl[5] br[5] wl[79] vdd gnd cell_6t
Xbit_r80_c5 bl[5] br[5] wl[80] vdd gnd cell_6t
Xbit_r81_c5 bl[5] br[5] wl[81] vdd gnd cell_6t
Xbit_r82_c5 bl[5] br[5] wl[82] vdd gnd cell_6t
Xbit_r83_c5 bl[5] br[5] wl[83] vdd gnd cell_6t
Xbit_r84_c5 bl[5] br[5] wl[84] vdd gnd cell_6t
Xbit_r85_c5 bl[5] br[5] wl[85] vdd gnd cell_6t
Xbit_r86_c5 bl[5] br[5] wl[86] vdd gnd cell_6t
Xbit_r87_c5 bl[5] br[5] wl[87] vdd gnd cell_6t
Xbit_r88_c5 bl[5] br[5] wl[88] vdd gnd cell_6t
Xbit_r89_c5 bl[5] br[5] wl[89] vdd gnd cell_6t
Xbit_r90_c5 bl[5] br[5] wl[90] vdd gnd cell_6t
Xbit_r91_c5 bl[5] br[5] wl[91] vdd gnd cell_6t
Xbit_r92_c5 bl[5] br[5] wl[92] vdd gnd cell_6t
Xbit_r93_c5 bl[5] br[5] wl[93] vdd gnd cell_6t
Xbit_r94_c5 bl[5] br[5] wl[94] vdd gnd cell_6t
Xbit_r95_c5 bl[5] br[5] wl[95] vdd gnd cell_6t
Xbit_r96_c5 bl[5] br[5] wl[96] vdd gnd cell_6t
Xbit_r97_c5 bl[5] br[5] wl[97] vdd gnd cell_6t
Xbit_r98_c5 bl[5] br[5] wl[98] vdd gnd cell_6t
Xbit_r99_c5 bl[5] br[5] wl[99] vdd gnd cell_6t
Xbit_r100_c5 bl[5] br[5] wl[100] vdd gnd cell_6t
Xbit_r101_c5 bl[5] br[5] wl[101] vdd gnd cell_6t
Xbit_r102_c5 bl[5] br[5] wl[102] vdd gnd cell_6t
Xbit_r103_c5 bl[5] br[5] wl[103] vdd gnd cell_6t
Xbit_r104_c5 bl[5] br[5] wl[104] vdd gnd cell_6t
Xbit_r105_c5 bl[5] br[5] wl[105] vdd gnd cell_6t
Xbit_r106_c5 bl[5] br[5] wl[106] vdd gnd cell_6t
Xbit_r107_c5 bl[5] br[5] wl[107] vdd gnd cell_6t
Xbit_r108_c5 bl[5] br[5] wl[108] vdd gnd cell_6t
Xbit_r109_c5 bl[5] br[5] wl[109] vdd gnd cell_6t
Xbit_r110_c5 bl[5] br[5] wl[110] vdd gnd cell_6t
Xbit_r111_c5 bl[5] br[5] wl[111] vdd gnd cell_6t
Xbit_r112_c5 bl[5] br[5] wl[112] vdd gnd cell_6t
Xbit_r113_c5 bl[5] br[5] wl[113] vdd gnd cell_6t
Xbit_r114_c5 bl[5] br[5] wl[114] vdd gnd cell_6t
Xbit_r115_c5 bl[5] br[5] wl[115] vdd gnd cell_6t
Xbit_r116_c5 bl[5] br[5] wl[116] vdd gnd cell_6t
Xbit_r117_c5 bl[5] br[5] wl[117] vdd gnd cell_6t
Xbit_r118_c5 bl[5] br[5] wl[118] vdd gnd cell_6t
Xbit_r119_c5 bl[5] br[5] wl[119] vdd gnd cell_6t
Xbit_r120_c5 bl[5] br[5] wl[120] vdd gnd cell_6t
Xbit_r121_c5 bl[5] br[5] wl[121] vdd gnd cell_6t
Xbit_r122_c5 bl[5] br[5] wl[122] vdd gnd cell_6t
Xbit_r123_c5 bl[5] br[5] wl[123] vdd gnd cell_6t
Xbit_r124_c5 bl[5] br[5] wl[124] vdd gnd cell_6t
Xbit_r125_c5 bl[5] br[5] wl[125] vdd gnd cell_6t
Xbit_r126_c5 bl[5] br[5] wl[126] vdd gnd cell_6t
Xbit_r127_c5 bl[5] br[5] wl[127] vdd gnd cell_6t
Xbit_r128_c5 bl[5] br[5] wl[128] vdd gnd cell_6t
Xbit_r129_c5 bl[5] br[5] wl[129] vdd gnd cell_6t
Xbit_r130_c5 bl[5] br[5] wl[130] vdd gnd cell_6t
Xbit_r131_c5 bl[5] br[5] wl[131] vdd gnd cell_6t
Xbit_r132_c5 bl[5] br[5] wl[132] vdd gnd cell_6t
Xbit_r133_c5 bl[5] br[5] wl[133] vdd gnd cell_6t
Xbit_r134_c5 bl[5] br[5] wl[134] vdd gnd cell_6t
Xbit_r135_c5 bl[5] br[5] wl[135] vdd gnd cell_6t
Xbit_r136_c5 bl[5] br[5] wl[136] vdd gnd cell_6t
Xbit_r137_c5 bl[5] br[5] wl[137] vdd gnd cell_6t
Xbit_r138_c5 bl[5] br[5] wl[138] vdd gnd cell_6t
Xbit_r139_c5 bl[5] br[5] wl[139] vdd gnd cell_6t
Xbit_r140_c5 bl[5] br[5] wl[140] vdd gnd cell_6t
Xbit_r141_c5 bl[5] br[5] wl[141] vdd gnd cell_6t
Xbit_r142_c5 bl[5] br[5] wl[142] vdd gnd cell_6t
Xbit_r143_c5 bl[5] br[5] wl[143] vdd gnd cell_6t
Xbit_r144_c5 bl[5] br[5] wl[144] vdd gnd cell_6t
Xbit_r145_c5 bl[5] br[5] wl[145] vdd gnd cell_6t
Xbit_r146_c5 bl[5] br[5] wl[146] vdd gnd cell_6t
Xbit_r147_c5 bl[5] br[5] wl[147] vdd gnd cell_6t
Xbit_r148_c5 bl[5] br[5] wl[148] vdd gnd cell_6t
Xbit_r149_c5 bl[5] br[5] wl[149] vdd gnd cell_6t
Xbit_r150_c5 bl[5] br[5] wl[150] vdd gnd cell_6t
Xbit_r151_c5 bl[5] br[5] wl[151] vdd gnd cell_6t
Xbit_r152_c5 bl[5] br[5] wl[152] vdd gnd cell_6t
Xbit_r153_c5 bl[5] br[5] wl[153] vdd gnd cell_6t
Xbit_r154_c5 bl[5] br[5] wl[154] vdd gnd cell_6t
Xbit_r155_c5 bl[5] br[5] wl[155] vdd gnd cell_6t
Xbit_r156_c5 bl[5] br[5] wl[156] vdd gnd cell_6t
Xbit_r157_c5 bl[5] br[5] wl[157] vdd gnd cell_6t
Xbit_r158_c5 bl[5] br[5] wl[158] vdd gnd cell_6t
Xbit_r159_c5 bl[5] br[5] wl[159] vdd gnd cell_6t
Xbit_r160_c5 bl[5] br[5] wl[160] vdd gnd cell_6t
Xbit_r161_c5 bl[5] br[5] wl[161] vdd gnd cell_6t
Xbit_r162_c5 bl[5] br[5] wl[162] vdd gnd cell_6t
Xbit_r163_c5 bl[5] br[5] wl[163] vdd gnd cell_6t
Xbit_r164_c5 bl[5] br[5] wl[164] vdd gnd cell_6t
Xbit_r165_c5 bl[5] br[5] wl[165] vdd gnd cell_6t
Xbit_r166_c5 bl[5] br[5] wl[166] vdd gnd cell_6t
Xbit_r167_c5 bl[5] br[5] wl[167] vdd gnd cell_6t
Xbit_r168_c5 bl[5] br[5] wl[168] vdd gnd cell_6t
Xbit_r169_c5 bl[5] br[5] wl[169] vdd gnd cell_6t
Xbit_r170_c5 bl[5] br[5] wl[170] vdd gnd cell_6t
Xbit_r171_c5 bl[5] br[5] wl[171] vdd gnd cell_6t
Xbit_r172_c5 bl[5] br[5] wl[172] vdd gnd cell_6t
Xbit_r173_c5 bl[5] br[5] wl[173] vdd gnd cell_6t
Xbit_r174_c5 bl[5] br[5] wl[174] vdd gnd cell_6t
Xbit_r175_c5 bl[5] br[5] wl[175] vdd gnd cell_6t
Xbit_r176_c5 bl[5] br[5] wl[176] vdd gnd cell_6t
Xbit_r177_c5 bl[5] br[5] wl[177] vdd gnd cell_6t
Xbit_r178_c5 bl[5] br[5] wl[178] vdd gnd cell_6t
Xbit_r179_c5 bl[5] br[5] wl[179] vdd gnd cell_6t
Xbit_r180_c5 bl[5] br[5] wl[180] vdd gnd cell_6t
Xbit_r181_c5 bl[5] br[5] wl[181] vdd gnd cell_6t
Xbit_r182_c5 bl[5] br[5] wl[182] vdd gnd cell_6t
Xbit_r183_c5 bl[5] br[5] wl[183] vdd gnd cell_6t
Xbit_r184_c5 bl[5] br[5] wl[184] vdd gnd cell_6t
Xbit_r185_c5 bl[5] br[5] wl[185] vdd gnd cell_6t
Xbit_r186_c5 bl[5] br[5] wl[186] vdd gnd cell_6t
Xbit_r187_c5 bl[5] br[5] wl[187] vdd gnd cell_6t
Xbit_r188_c5 bl[5] br[5] wl[188] vdd gnd cell_6t
Xbit_r189_c5 bl[5] br[5] wl[189] vdd gnd cell_6t
Xbit_r190_c5 bl[5] br[5] wl[190] vdd gnd cell_6t
Xbit_r191_c5 bl[5] br[5] wl[191] vdd gnd cell_6t
Xbit_r192_c5 bl[5] br[5] wl[192] vdd gnd cell_6t
Xbit_r193_c5 bl[5] br[5] wl[193] vdd gnd cell_6t
Xbit_r194_c5 bl[5] br[5] wl[194] vdd gnd cell_6t
Xbit_r195_c5 bl[5] br[5] wl[195] vdd gnd cell_6t
Xbit_r196_c5 bl[5] br[5] wl[196] vdd gnd cell_6t
Xbit_r197_c5 bl[5] br[5] wl[197] vdd gnd cell_6t
Xbit_r198_c5 bl[5] br[5] wl[198] vdd gnd cell_6t
Xbit_r199_c5 bl[5] br[5] wl[199] vdd gnd cell_6t
Xbit_r200_c5 bl[5] br[5] wl[200] vdd gnd cell_6t
Xbit_r201_c5 bl[5] br[5] wl[201] vdd gnd cell_6t
Xbit_r202_c5 bl[5] br[5] wl[202] vdd gnd cell_6t
Xbit_r203_c5 bl[5] br[5] wl[203] vdd gnd cell_6t
Xbit_r204_c5 bl[5] br[5] wl[204] vdd gnd cell_6t
Xbit_r205_c5 bl[5] br[5] wl[205] vdd gnd cell_6t
Xbit_r206_c5 bl[5] br[5] wl[206] vdd gnd cell_6t
Xbit_r207_c5 bl[5] br[5] wl[207] vdd gnd cell_6t
Xbit_r208_c5 bl[5] br[5] wl[208] vdd gnd cell_6t
Xbit_r209_c5 bl[5] br[5] wl[209] vdd gnd cell_6t
Xbit_r210_c5 bl[5] br[5] wl[210] vdd gnd cell_6t
Xbit_r211_c5 bl[5] br[5] wl[211] vdd gnd cell_6t
Xbit_r212_c5 bl[5] br[5] wl[212] vdd gnd cell_6t
Xbit_r213_c5 bl[5] br[5] wl[213] vdd gnd cell_6t
Xbit_r214_c5 bl[5] br[5] wl[214] vdd gnd cell_6t
Xbit_r215_c5 bl[5] br[5] wl[215] vdd gnd cell_6t
Xbit_r216_c5 bl[5] br[5] wl[216] vdd gnd cell_6t
Xbit_r217_c5 bl[5] br[5] wl[217] vdd gnd cell_6t
Xbit_r218_c5 bl[5] br[5] wl[218] vdd gnd cell_6t
Xbit_r219_c5 bl[5] br[5] wl[219] vdd gnd cell_6t
Xbit_r220_c5 bl[5] br[5] wl[220] vdd gnd cell_6t
Xbit_r221_c5 bl[5] br[5] wl[221] vdd gnd cell_6t
Xbit_r222_c5 bl[5] br[5] wl[222] vdd gnd cell_6t
Xbit_r223_c5 bl[5] br[5] wl[223] vdd gnd cell_6t
Xbit_r224_c5 bl[5] br[5] wl[224] vdd gnd cell_6t
Xbit_r225_c5 bl[5] br[5] wl[225] vdd gnd cell_6t
Xbit_r226_c5 bl[5] br[5] wl[226] vdd gnd cell_6t
Xbit_r227_c5 bl[5] br[5] wl[227] vdd gnd cell_6t
Xbit_r228_c5 bl[5] br[5] wl[228] vdd gnd cell_6t
Xbit_r229_c5 bl[5] br[5] wl[229] vdd gnd cell_6t
Xbit_r230_c5 bl[5] br[5] wl[230] vdd gnd cell_6t
Xbit_r231_c5 bl[5] br[5] wl[231] vdd gnd cell_6t
Xbit_r232_c5 bl[5] br[5] wl[232] vdd gnd cell_6t
Xbit_r233_c5 bl[5] br[5] wl[233] vdd gnd cell_6t
Xbit_r234_c5 bl[5] br[5] wl[234] vdd gnd cell_6t
Xbit_r235_c5 bl[5] br[5] wl[235] vdd gnd cell_6t
Xbit_r236_c5 bl[5] br[5] wl[236] vdd gnd cell_6t
Xbit_r237_c5 bl[5] br[5] wl[237] vdd gnd cell_6t
Xbit_r238_c5 bl[5] br[5] wl[238] vdd gnd cell_6t
Xbit_r239_c5 bl[5] br[5] wl[239] vdd gnd cell_6t
Xbit_r240_c5 bl[5] br[5] wl[240] vdd gnd cell_6t
Xbit_r241_c5 bl[5] br[5] wl[241] vdd gnd cell_6t
Xbit_r242_c5 bl[5] br[5] wl[242] vdd gnd cell_6t
Xbit_r243_c5 bl[5] br[5] wl[243] vdd gnd cell_6t
Xbit_r244_c5 bl[5] br[5] wl[244] vdd gnd cell_6t
Xbit_r245_c5 bl[5] br[5] wl[245] vdd gnd cell_6t
Xbit_r246_c5 bl[5] br[5] wl[246] vdd gnd cell_6t
Xbit_r247_c5 bl[5] br[5] wl[247] vdd gnd cell_6t
Xbit_r248_c5 bl[5] br[5] wl[248] vdd gnd cell_6t
Xbit_r249_c5 bl[5] br[5] wl[249] vdd gnd cell_6t
Xbit_r250_c5 bl[5] br[5] wl[250] vdd gnd cell_6t
Xbit_r251_c5 bl[5] br[5] wl[251] vdd gnd cell_6t
Xbit_r252_c5 bl[5] br[5] wl[252] vdd gnd cell_6t
Xbit_r253_c5 bl[5] br[5] wl[253] vdd gnd cell_6t
Xbit_r254_c5 bl[5] br[5] wl[254] vdd gnd cell_6t
Xbit_r255_c5 bl[5] br[5] wl[255] vdd gnd cell_6t
Xbit_r256_c5 bl[5] br[5] wl[256] vdd gnd cell_6t
Xbit_r257_c5 bl[5] br[5] wl[257] vdd gnd cell_6t
Xbit_r258_c5 bl[5] br[5] wl[258] vdd gnd cell_6t
Xbit_r259_c5 bl[5] br[5] wl[259] vdd gnd cell_6t
Xbit_r260_c5 bl[5] br[5] wl[260] vdd gnd cell_6t
Xbit_r261_c5 bl[5] br[5] wl[261] vdd gnd cell_6t
Xbit_r262_c5 bl[5] br[5] wl[262] vdd gnd cell_6t
Xbit_r263_c5 bl[5] br[5] wl[263] vdd gnd cell_6t
Xbit_r264_c5 bl[5] br[5] wl[264] vdd gnd cell_6t
Xbit_r265_c5 bl[5] br[5] wl[265] vdd gnd cell_6t
Xbit_r266_c5 bl[5] br[5] wl[266] vdd gnd cell_6t
Xbit_r267_c5 bl[5] br[5] wl[267] vdd gnd cell_6t
Xbit_r268_c5 bl[5] br[5] wl[268] vdd gnd cell_6t
Xbit_r269_c5 bl[5] br[5] wl[269] vdd gnd cell_6t
Xbit_r270_c5 bl[5] br[5] wl[270] vdd gnd cell_6t
Xbit_r271_c5 bl[5] br[5] wl[271] vdd gnd cell_6t
Xbit_r272_c5 bl[5] br[5] wl[272] vdd gnd cell_6t
Xbit_r273_c5 bl[5] br[5] wl[273] vdd gnd cell_6t
Xbit_r274_c5 bl[5] br[5] wl[274] vdd gnd cell_6t
Xbit_r275_c5 bl[5] br[5] wl[275] vdd gnd cell_6t
Xbit_r276_c5 bl[5] br[5] wl[276] vdd gnd cell_6t
Xbit_r277_c5 bl[5] br[5] wl[277] vdd gnd cell_6t
Xbit_r278_c5 bl[5] br[5] wl[278] vdd gnd cell_6t
Xbit_r279_c5 bl[5] br[5] wl[279] vdd gnd cell_6t
Xbit_r280_c5 bl[5] br[5] wl[280] vdd gnd cell_6t
Xbit_r281_c5 bl[5] br[5] wl[281] vdd gnd cell_6t
Xbit_r282_c5 bl[5] br[5] wl[282] vdd gnd cell_6t
Xbit_r283_c5 bl[5] br[5] wl[283] vdd gnd cell_6t
Xbit_r284_c5 bl[5] br[5] wl[284] vdd gnd cell_6t
Xbit_r285_c5 bl[5] br[5] wl[285] vdd gnd cell_6t
Xbit_r286_c5 bl[5] br[5] wl[286] vdd gnd cell_6t
Xbit_r287_c5 bl[5] br[5] wl[287] vdd gnd cell_6t
Xbit_r288_c5 bl[5] br[5] wl[288] vdd gnd cell_6t
Xbit_r289_c5 bl[5] br[5] wl[289] vdd gnd cell_6t
Xbit_r290_c5 bl[5] br[5] wl[290] vdd gnd cell_6t
Xbit_r291_c5 bl[5] br[5] wl[291] vdd gnd cell_6t
Xbit_r292_c5 bl[5] br[5] wl[292] vdd gnd cell_6t
Xbit_r293_c5 bl[5] br[5] wl[293] vdd gnd cell_6t
Xbit_r294_c5 bl[5] br[5] wl[294] vdd gnd cell_6t
Xbit_r295_c5 bl[5] br[5] wl[295] vdd gnd cell_6t
Xbit_r296_c5 bl[5] br[5] wl[296] vdd gnd cell_6t
Xbit_r297_c5 bl[5] br[5] wl[297] vdd gnd cell_6t
Xbit_r298_c5 bl[5] br[5] wl[298] vdd gnd cell_6t
Xbit_r299_c5 bl[5] br[5] wl[299] vdd gnd cell_6t
Xbit_r300_c5 bl[5] br[5] wl[300] vdd gnd cell_6t
Xbit_r301_c5 bl[5] br[5] wl[301] vdd gnd cell_6t
Xbit_r302_c5 bl[5] br[5] wl[302] vdd gnd cell_6t
Xbit_r303_c5 bl[5] br[5] wl[303] vdd gnd cell_6t
Xbit_r304_c5 bl[5] br[5] wl[304] vdd gnd cell_6t
Xbit_r305_c5 bl[5] br[5] wl[305] vdd gnd cell_6t
Xbit_r306_c5 bl[5] br[5] wl[306] vdd gnd cell_6t
Xbit_r307_c5 bl[5] br[5] wl[307] vdd gnd cell_6t
Xbit_r308_c5 bl[5] br[5] wl[308] vdd gnd cell_6t
Xbit_r309_c5 bl[5] br[5] wl[309] vdd gnd cell_6t
Xbit_r310_c5 bl[5] br[5] wl[310] vdd gnd cell_6t
Xbit_r311_c5 bl[5] br[5] wl[311] vdd gnd cell_6t
Xbit_r312_c5 bl[5] br[5] wl[312] vdd gnd cell_6t
Xbit_r313_c5 bl[5] br[5] wl[313] vdd gnd cell_6t
Xbit_r314_c5 bl[5] br[5] wl[314] vdd gnd cell_6t
Xbit_r315_c5 bl[5] br[5] wl[315] vdd gnd cell_6t
Xbit_r316_c5 bl[5] br[5] wl[316] vdd gnd cell_6t
Xbit_r317_c5 bl[5] br[5] wl[317] vdd gnd cell_6t
Xbit_r318_c5 bl[5] br[5] wl[318] vdd gnd cell_6t
Xbit_r319_c5 bl[5] br[5] wl[319] vdd gnd cell_6t
Xbit_r320_c5 bl[5] br[5] wl[320] vdd gnd cell_6t
Xbit_r321_c5 bl[5] br[5] wl[321] vdd gnd cell_6t
Xbit_r322_c5 bl[5] br[5] wl[322] vdd gnd cell_6t
Xbit_r323_c5 bl[5] br[5] wl[323] vdd gnd cell_6t
Xbit_r324_c5 bl[5] br[5] wl[324] vdd gnd cell_6t
Xbit_r325_c5 bl[5] br[5] wl[325] vdd gnd cell_6t
Xbit_r326_c5 bl[5] br[5] wl[326] vdd gnd cell_6t
Xbit_r327_c5 bl[5] br[5] wl[327] vdd gnd cell_6t
Xbit_r328_c5 bl[5] br[5] wl[328] vdd gnd cell_6t
Xbit_r329_c5 bl[5] br[5] wl[329] vdd gnd cell_6t
Xbit_r330_c5 bl[5] br[5] wl[330] vdd gnd cell_6t
Xbit_r331_c5 bl[5] br[5] wl[331] vdd gnd cell_6t
Xbit_r332_c5 bl[5] br[5] wl[332] vdd gnd cell_6t
Xbit_r333_c5 bl[5] br[5] wl[333] vdd gnd cell_6t
Xbit_r334_c5 bl[5] br[5] wl[334] vdd gnd cell_6t
Xbit_r335_c5 bl[5] br[5] wl[335] vdd gnd cell_6t
Xbit_r336_c5 bl[5] br[5] wl[336] vdd gnd cell_6t
Xbit_r337_c5 bl[5] br[5] wl[337] vdd gnd cell_6t
Xbit_r338_c5 bl[5] br[5] wl[338] vdd gnd cell_6t
Xbit_r339_c5 bl[5] br[5] wl[339] vdd gnd cell_6t
Xbit_r340_c5 bl[5] br[5] wl[340] vdd gnd cell_6t
Xbit_r341_c5 bl[5] br[5] wl[341] vdd gnd cell_6t
Xbit_r342_c5 bl[5] br[5] wl[342] vdd gnd cell_6t
Xbit_r343_c5 bl[5] br[5] wl[343] vdd gnd cell_6t
Xbit_r344_c5 bl[5] br[5] wl[344] vdd gnd cell_6t
Xbit_r345_c5 bl[5] br[5] wl[345] vdd gnd cell_6t
Xbit_r346_c5 bl[5] br[5] wl[346] vdd gnd cell_6t
Xbit_r347_c5 bl[5] br[5] wl[347] vdd gnd cell_6t
Xbit_r348_c5 bl[5] br[5] wl[348] vdd gnd cell_6t
Xbit_r349_c5 bl[5] br[5] wl[349] vdd gnd cell_6t
Xbit_r350_c5 bl[5] br[5] wl[350] vdd gnd cell_6t
Xbit_r351_c5 bl[5] br[5] wl[351] vdd gnd cell_6t
Xbit_r352_c5 bl[5] br[5] wl[352] vdd gnd cell_6t
Xbit_r353_c5 bl[5] br[5] wl[353] vdd gnd cell_6t
Xbit_r354_c5 bl[5] br[5] wl[354] vdd gnd cell_6t
Xbit_r355_c5 bl[5] br[5] wl[355] vdd gnd cell_6t
Xbit_r356_c5 bl[5] br[5] wl[356] vdd gnd cell_6t
Xbit_r357_c5 bl[5] br[5] wl[357] vdd gnd cell_6t
Xbit_r358_c5 bl[5] br[5] wl[358] vdd gnd cell_6t
Xbit_r359_c5 bl[5] br[5] wl[359] vdd gnd cell_6t
Xbit_r360_c5 bl[5] br[5] wl[360] vdd gnd cell_6t
Xbit_r361_c5 bl[5] br[5] wl[361] vdd gnd cell_6t
Xbit_r362_c5 bl[5] br[5] wl[362] vdd gnd cell_6t
Xbit_r363_c5 bl[5] br[5] wl[363] vdd gnd cell_6t
Xbit_r364_c5 bl[5] br[5] wl[364] vdd gnd cell_6t
Xbit_r365_c5 bl[5] br[5] wl[365] vdd gnd cell_6t
Xbit_r366_c5 bl[5] br[5] wl[366] vdd gnd cell_6t
Xbit_r367_c5 bl[5] br[5] wl[367] vdd gnd cell_6t
Xbit_r368_c5 bl[5] br[5] wl[368] vdd gnd cell_6t
Xbit_r369_c5 bl[5] br[5] wl[369] vdd gnd cell_6t
Xbit_r370_c5 bl[5] br[5] wl[370] vdd gnd cell_6t
Xbit_r371_c5 bl[5] br[5] wl[371] vdd gnd cell_6t
Xbit_r372_c5 bl[5] br[5] wl[372] vdd gnd cell_6t
Xbit_r373_c5 bl[5] br[5] wl[373] vdd gnd cell_6t
Xbit_r374_c5 bl[5] br[5] wl[374] vdd gnd cell_6t
Xbit_r375_c5 bl[5] br[5] wl[375] vdd gnd cell_6t
Xbit_r376_c5 bl[5] br[5] wl[376] vdd gnd cell_6t
Xbit_r377_c5 bl[5] br[5] wl[377] vdd gnd cell_6t
Xbit_r378_c5 bl[5] br[5] wl[378] vdd gnd cell_6t
Xbit_r379_c5 bl[5] br[5] wl[379] vdd gnd cell_6t
Xbit_r380_c5 bl[5] br[5] wl[380] vdd gnd cell_6t
Xbit_r381_c5 bl[5] br[5] wl[381] vdd gnd cell_6t
Xbit_r382_c5 bl[5] br[5] wl[382] vdd gnd cell_6t
Xbit_r383_c5 bl[5] br[5] wl[383] vdd gnd cell_6t
Xbit_r384_c5 bl[5] br[5] wl[384] vdd gnd cell_6t
Xbit_r385_c5 bl[5] br[5] wl[385] vdd gnd cell_6t
Xbit_r386_c5 bl[5] br[5] wl[386] vdd gnd cell_6t
Xbit_r387_c5 bl[5] br[5] wl[387] vdd gnd cell_6t
Xbit_r388_c5 bl[5] br[5] wl[388] vdd gnd cell_6t
Xbit_r389_c5 bl[5] br[5] wl[389] vdd gnd cell_6t
Xbit_r390_c5 bl[5] br[5] wl[390] vdd gnd cell_6t
Xbit_r391_c5 bl[5] br[5] wl[391] vdd gnd cell_6t
Xbit_r392_c5 bl[5] br[5] wl[392] vdd gnd cell_6t
Xbit_r393_c5 bl[5] br[5] wl[393] vdd gnd cell_6t
Xbit_r394_c5 bl[5] br[5] wl[394] vdd gnd cell_6t
Xbit_r395_c5 bl[5] br[5] wl[395] vdd gnd cell_6t
Xbit_r396_c5 bl[5] br[5] wl[396] vdd gnd cell_6t
Xbit_r397_c5 bl[5] br[5] wl[397] vdd gnd cell_6t
Xbit_r398_c5 bl[5] br[5] wl[398] vdd gnd cell_6t
Xbit_r399_c5 bl[5] br[5] wl[399] vdd gnd cell_6t
Xbit_r400_c5 bl[5] br[5] wl[400] vdd gnd cell_6t
Xbit_r401_c5 bl[5] br[5] wl[401] vdd gnd cell_6t
Xbit_r402_c5 bl[5] br[5] wl[402] vdd gnd cell_6t
Xbit_r403_c5 bl[5] br[5] wl[403] vdd gnd cell_6t
Xbit_r404_c5 bl[5] br[5] wl[404] vdd gnd cell_6t
Xbit_r405_c5 bl[5] br[5] wl[405] vdd gnd cell_6t
Xbit_r406_c5 bl[5] br[5] wl[406] vdd gnd cell_6t
Xbit_r407_c5 bl[5] br[5] wl[407] vdd gnd cell_6t
Xbit_r408_c5 bl[5] br[5] wl[408] vdd gnd cell_6t
Xbit_r409_c5 bl[5] br[5] wl[409] vdd gnd cell_6t
Xbit_r410_c5 bl[5] br[5] wl[410] vdd gnd cell_6t
Xbit_r411_c5 bl[5] br[5] wl[411] vdd gnd cell_6t
Xbit_r412_c5 bl[5] br[5] wl[412] vdd gnd cell_6t
Xbit_r413_c5 bl[5] br[5] wl[413] vdd gnd cell_6t
Xbit_r414_c5 bl[5] br[5] wl[414] vdd gnd cell_6t
Xbit_r415_c5 bl[5] br[5] wl[415] vdd gnd cell_6t
Xbit_r416_c5 bl[5] br[5] wl[416] vdd gnd cell_6t
Xbit_r417_c5 bl[5] br[5] wl[417] vdd gnd cell_6t
Xbit_r418_c5 bl[5] br[5] wl[418] vdd gnd cell_6t
Xbit_r419_c5 bl[5] br[5] wl[419] vdd gnd cell_6t
Xbit_r420_c5 bl[5] br[5] wl[420] vdd gnd cell_6t
Xbit_r421_c5 bl[5] br[5] wl[421] vdd gnd cell_6t
Xbit_r422_c5 bl[5] br[5] wl[422] vdd gnd cell_6t
Xbit_r423_c5 bl[5] br[5] wl[423] vdd gnd cell_6t
Xbit_r424_c5 bl[5] br[5] wl[424] vdd gnd cell_6t
Xbit_r425_c5 bl[5] br[5] wl[425] vdd gnd cell_6t
Xbit_r426_c5 bl[5] br[5] wl[426] vdd gnd cell_6t
Xbit_r427_c5 bl[5] br[5] wl[427] vdd gnd cell_6t
Xbit_r428_c5 bl[5] br[5] wl[428] vdd gnd cell_6t
Xbit_r429_c5 bl[5] br[5] wl[429] vdd gnd cell_6t
Xbit_r430_c5 bl[5] br[5] wl[430] vdd gnd cell_6t
Xbit_r431_c5 bl[5] br[5] wl[431] vdd gnd cell_6t
Xbit_r432_c5 bl[5] br[5] wl[432] vdd gnd cell_6t
Xbit_r433_c5 bl[5] br[5] wl[433] vdd gnd cell_6t
Xbit_r434_c5 bl[5] br[5] wl[434] vdd gnd cell_6t
Xbit_r435_c5 bl[5] br[5] wl[435] vdd gnd cell_6t
Xbit_r436_c5 bl[5] br[5] wl[436] vdd gnd cell_6t
Xbit_r437_c5 bl[5] br[5] wl[437] vdd gnd cell_6t
Xbit_r438_c5 bl[5] br[5] wl[438] vdd gnd cell_6t
Xbit_r439_c5 bl[5] br[5] wl[439] vdd gnd cell_6t
Xbit_r440_c5 bl[5] br[5] wl[440] vdd gnd cell_6t
Xbit_r441_c5 bl[5] br[5] wl[441] vdd gnd cell_6t
Xbit_r442_c5 bl[5] br[5] wl[442] vdd gnd cell_6t
Xbit_r443_c5 bl[5] br[5] wl[443] vdd gnd cell_6t
Xbit_r444_c5 bl[5] br[5] wl[444] vdd gnd cell_6t
Xbit_r445_c5 bl[5] br[5] wl[445] vdd gnd cell_6t
Xbit_r446_c5 bl[5] br[5] wl[446] vdd gnd cell_6t
Xbit_r447_c5 bl[5] br[5] wl[447] vdd gnd cell_6t
Xbit_r448_c5 bl[5] br[5] wl[448] vdd gnd cell_6t
Xbit_r449_c5 bl[5] br[5] wl[449] vdd gnd cell_6t
Xbit_r450_c5 bl[5] br[5] wl[450] vdd gnd cell_6t
Xbit_r451_c5 bl[5] br[5] wl[451] vdd gnd cell_6t
Xbit_r452_c5 bl[5] br[5] wl[452] vdd gnd cell_6t
Xbit_r453_c5 bl[5] br[5] wl[453] vdd gnd cell_6t
Xbit_r454_c5 bl[5] br[5] wl[454] vdd gnd cell_6t
Xbit_r455_c5 bl[5] br[5] wl[455] vdd gnd cell_6t
Xbit_r456_c5 bl[5] br[5] wl[456] vdd gnd cell_6t
Xbit_r457_c5 bl[5] br[5] wl[457] vdd gnd cell_6t
Xbit_r458_c5 bl[5] br[5] wl[458] vdd gnd cell_6t
Xbit_r459_c5 bl[5] br[5] wl[459] vdd gnd cell_6t
Xbit_r460_c5 bl[5] br[5] wl[460] vdd gnd cell_6t
Xbit_r461_c5 bl[5] br[5] wl[461] vdd gnd cell_6t
Xbit_r462_c5 bl[5] br[5] wl[462] vdd gnd cell_6t
Xbit_r463_c5 bl[5] br[5] wl[463] vdd gnd cell_6t
Xbit_r464_c5 bl[5] br[5] wl[464] vdd gnd cell_6t
Xbit_r465_c5 bl[5] br[5] wl[465] vdd gnd cell_6t
Xbit_r466_c5 bl[5] br[5] wl[466] vdd gnd cell_6t
Xbit_r467_c5 bl[5] br[5] wl[467] vdd gnd cell_6t
Xbit_r468_c5 bl[5] br[5] wl[468] vdd gnd cell_6t
Xbit_r469_c5 bl[5] br[5] wl[469] vdd gnd cell_6t
Xbit_r470_c5 bl[5] br[5] wl[470] vdd gnd cell_6t
Xbit_r471_c5 bl[5] br[5] wl[471] vdd gnd cell_6t
Xbit_r472_c5 bl[5] br[5] wl[472] vdd gnd cell_6t
Xbit_r473_c5 bl[5] br[5] wl[473] vdd gnd cell_6t
Xbit_r474_c5 bl[5] br[5] wl[474] vdd gnd cell_6t
Xbit_r475_c5 bl[5] br[5] wl[475] vdd gnd cell_6t
Xbit_r476_c5 bl[5] br[5] wl[476] vdd gnd cell_6t
Xbit_r477_c5 bl[5] br[5] wl[477] vdd gnd cell_6t
Xbit_r478_c5 bl[5] br[5] wl[478] vdd gnd cell_6t
Xbit_r479_c5 bl[5] br[5] wl[479] vdd gnd cell_6t
Xbit_r480_c5 bl[5] br[5] wl[480] vdd gnd cell_6t
Xbit_r481_c5 bl[5] br[5] wl[481] vdd gnd cell_6t
Xbit_r482_c5 bl[5] br[5] wl[482] vdd gnd cell_6t
Xbit_r483_c5 bl[5] br[5] wl[483] vdd gnd cell_6t
Xbit_r484_c5 bl[5] br[5] wl[484] vdd gnd cell_6t
Xbit_r485_c5 bl[5] br[5] wl[485] vdd gnd cell_6t
Xbit_r486_c5 bl[5] br[5] wl[486] vdd gnd cell_6t
Xbit_r487_c5 bl[5] br[5] wl[487] vdd gnd cell_6t
Xbit_r488_c5 bl[5] br[5] wl[488] vdd gnd cell_6t
Xbit_r489_c5 bl[5] br[5] wl[489] vdd gnd cell_6t
Xbit_r490_c5 bl[5] br[5] wl[490] vdd gnd cell_6t
Xbit_r491_c5 bl[5] br[5] wl[491] vdd gnd cell_6t
Xbit_r492_c5 bl[5] br[5] wl[492] vdd gnd cell_6t
Xbit_r493_c5 bl[5] br[5] wl[493] vdd gnd cell_6t
Xbit_r494_c5 bl[5] br[5] wl[494] vdd gnd cell_6t
Xbit_r495_c5 bl[5] br[5] wl[495] vdd gnd cell_6t
Xbit_r496_c5 bl[5] br[5] wl[496] vdd gnd cell_6t
Xbit_r497_c5 bl[5] br[5] wl[497] vdd gnd cell_6t
Xbit_r498_c5 bl[5] br[5] wl[498] vdd gnd cell_6t
Xbit_r499_c5 bl[5] br[5] wl[499] vdd gnd cell_6t
Xbit_r500_c5 bl[5] br[5] wl[500] vdd gnd cell_6t
Xbit_r501_c5 bl[5] br[5] wl[501] vdd gnd cell_6t
Xbit_r502_c5 bl[5] br[5] wl[502] vdd gnd cell_6t
Xbit_r503_c5 bl[5] br[5] wl[503] vdd gnd cell_6t
Xbit_r504_c5 bl[5] br[5] wl[504] vdd gnd cell_6t
Xbit_r505_c5 bl[5] br[5] wl[505] vdd gnd cell_6t
Xbit_r506_c5 bl[5] br[5] wl[506] vdd gnd cell_6t
Xbit_r507_c5 bl[5] br[5] wl[507] vdd gnd cell_6t
Xbit_r508_c5 bl[5] br[5] wl[508] vdd gnd cell_6t
Xbit_r509_c5 bl[5] br[5] wl[509] vdd gnd cell_6t
Xbit_r510_c5 bl[5] br[5] wl[510] vdd gnd cell_6t
Xbit_r511_c5 bl[5] br[5] wl[511] vdd gnd cell_6t
Xbit_r0_c6 bl[6] br[6] wl[0] vdd gnd cell_6t
Xbit_r1_c6 bl[6] br[6] wl[1] vdd gnd cell_6t
Xbit_r2_c6 bl[6] br[6] wl[2] vdd gnd cell_6t
Xbit_r3_c6 bl[6] br[6] wl[3] vdd gnd cell_6t
Xbit_r4_c6 bl[6] br[6] wl[4] vdd gnd cell_6t
Xbit_r5_c6 bl[6] br[6] wl[5] vdd gnd cell_6t
Xbit_r6_c6 bl[6] br[6] wl[6] vdd gnd cell_6t
Xbit_r7_c6 bl[6] br[6] wl[7] vdd gnd cell_6t
Xbit_r8_c6 bl[6] br[6] wl[8] vdd gnd cell_6t
Xbit_r9_c6 bl[6] br[6] wl[9] vdd gnd cell_6t
Xbit_r10_c6 bl[6] br[6] wl[10] vdd gnd cell_6t
Xbit_r11_c6 bl[6] br[6] wl[11] vdd gnd cell_6t
Xbit_r12_c6 bl[6] br[6] wl[12] vdd gnd cell_6t
Xbit_r13_c6 bl[6] br[6] wl[13] vdd gnd cell_6t
Xbit_r14_c6 bl[6] br[6] wl[14] vdd gnd cell_6t
Xbit_r15_c6 bl[6] br[6] wl[15] vdd gnd cell_6t
Xbit_r16_c6 bl[6] br[6] wl[16] vdd gnd cell_6t
Xbit_r17_c6 bl[6] br[6] wl[17] vdd gnd cell_6t
Xbit_r18_c6 bl[6] br[6] wl[18] vdd gnd cell_6t
Xbit_r19_c6 bl[6] br[6] wl[19] vdd gnd cell_6t
Xbit_r20_c6 bl[6] br[6] wl[20] vdd gnd cell_6t
Xbit_r21_c6 bl[6] br[6] wl[21] vdd gnd cell_6t
Xbit_r22_c6 bl[6] br[6] wl[22] vdd gnd cell_6t
Xbit_r23_c6 bl[6] br[6] wl[23] vdd gnd cell_6t
Xbit_r24_c6 bl[6] br[6] wl[24] vdd gnd cell_6t
Xbit_r25_c6 bl[6] br[6] wl[25] vdd gnd cell_6t
Xbit_r26_c6 bl[6] br[6] wl[26] vdd gnd cell_6t
Xbit_r27_c6 bl[6] br[6] wl[27] vdd gnd cell_6t
Xbit_r28_c6 bl[6] br[6] wl[28] vdd gnd cell_6t
Xbit_r29_c6 bl[6] br[6] wl[29] vdd gnd cell_6t
Xbit_r30_c6 bl[6] br[6] wl[30] vdd gnd cell_6t
Xbit_r31_c6 bl[6] br[6] wl[31] vdd gnd cell_6t
Xbit_r32_c6 bl[6] br[6] wl[32] vdd gnd cell_6t
Xbit_r33_c6 bl[6] br[6] wl[33] vdd gnd cell_6t
Xbit_r34_c6 bl[6] br[6] wl[34] vdd gnd cell_6t
Xbit_r35_c6 bl[6] br[6] wl[35] vdd gnd cell_6t
Xbit_r36_c6 bl[6] br[6] wl[36] vdd gnd cell_6t
Xbit_r37_c6 bl[6] br[6] wl[37] vdd gnd cell_6t
Xbit_r38_c6 bl[6] br[6] wl[38] vdd gnd cell_6t
Xbit_r39_c6 bl[6] br[6] wl[39] vdd gnd cell_6t
Xbit_r40_c6 bl[6] br[6] wl[40] vdd gnd cell_6t
Xbit_r41_c6 bl[6] br[6] wl[41] vdd gnd cell_6t
Xbit_r42_c6 bl[6] br[6] wl[42] vdd gnd cell_6t
Xbit_r43_c6 bl[6] br[6] wl[43] vdd gnd cell_6t
Xbit_r44_c6 bl[6] br[6] wl[44] vdd gnd cell_6t
Xbit_r45_c6 bl[6] br[6] wl[45] vdd gnd cell_6t
Xbit_r46_c6 bl[6] br[6] wl[46] vdd gnd cell_6t
Xbit_r47_c6 bl[6] br[6] wl[47] vdd gnd cell_6t
Xbit_r48_c6 bl[6] br[6] wl[48] vdd gnd cell_6t
Xbit_r49_c6 bl[6] br[6] wl[49] vdd gnd cell_6t
Xbit_r50_c6 bl[6] br[6] wl[50] vdd gnd cell_6t
Xbit_r51_c6 bl[6] br[6] wl[51] vdd gnd cell_6t
Xbit_r52_c6 bl[6] br[6] wl[52] vdd gnd cell_6t
Xbit_r53_c6 bl[6] br[6] wl[53] vdd gnd cell_6t
Xbit_r54_c6 bl[6] br[6] wl[54] vdd gnd cell_6t
Xbit_r55_c6 bl[6] br[6] wl[55] vdd gnd cell_6t
Xbit_r56_c6 bl[6] br[6] wl[56] vdd gnd cell_6t
Xbit_r57_c6 bl[6] br[6] wl[57] vdd gnd cell_6t
Xbit_r58_c6 bl[6] br[6] wl[58] vdd gnd cell_6t
Xbit_r59_c6 bl[6] br[6] wl[59] vdd gnd cell_6t
Xbit_r60_c6 bl[6] br[6] wl[60] vdd gnd cell_6t
Xbit_r61_c6 bl[6] br[6] wl[61] vdd gnd cell_6t
Xbit_r62_c6 bl[6] br[6] wl[62] vdd gnd cell_6t
Xbit_r63_c6 bl[6] br[6] wl[63] vdd gnd cell_6t
Xbit_r64_c6 bl[6] br[6] wl[64] vdd gnd cell_6t
Xbit_r65_c6 bl[6] br[6] wl[65] vdd gnd cell_6t
Xbit_r66_c6 bl[6] br[6] wl[66] vdd gnd cell_6t
Xbit_r67_c6 bl[6] br[6] wl[67] vdd gnd cell_6t
Xbit_r68_c6 bl[6] br[6] wl[68] vdd gnd cell_6t
Xbit_r69_c6 bl[6] br[6] wl[69] vdd gnd cell_6t
Xbit_r70_c6 bl[6] br[6] wl[70] vdd gnd cell_6t
Xbit_r71_c6 bl[6] br[6] wl[71] vdd gnd cell_6t
Xbit_r72_c6 bl[6] br[6] wl[72] vdd gnd cell_6t
Xbit_r73_c6 bl[6] br[6] wl[73] vdd gnd cell_6t
Xbit_r74_c6 bl[6] br[6] wl[74] vdd gnd cell_6t
Xbit_r75_c6 bl[6] br[6] wl[75] vdd gnd cell_6t
Xbit_r76_c6 bl[6] br[6] wl[76] vdd gnd cell_6t
Xbit_r77_c6 bl[6] br[6] wl[77] vdd gnd cell_6t
Xbit_r78_c6 bl[6] br[6] wl[78] vdd gnd cell_6t
Xbit_r79_c6 bl[6] br[6] wl[79] vdd gnd cell_6t
Xbit_r80_c6 bl[6] br[6] wl[80] vdd gnd cell_6t
Xbit_r81_c6 bl[6] br[6] wl[81] vdd gnd cell_6t
Xbit_r82_c6 bl[6] br[6] wl[82] vdd gnd cell_6t
Xbit_r83_c6 bl[6] br[6] wl[83] vdd gnd cell_6t
Xbit_r84_c6 bl[6] br[6] wl[84] vdd gnd cell_6t
Xbit_r85_c6 bl[6] br[6] wl[85] vdd gnd cell_6t
Xbit_r86_c6 bl[6] br[6] wl[86] vdd gnd cell_6t
Xbit_r87_c6 bl[6] br[6] wl[87] vdd gnd cell_6t
Xbit_r88_c6 bl[6] br[6] wl[88] vdd gnd cell_6t
Xbit_r89_c6 bl[6] br[6] wl[89] vdd gnd cell_6t
Xbit_r90_c6 bl[6] br[6] wl[90] vdd gnd cell_6t
Xbit_r91_c6 bl[6] br[6] wl[91] vdd gnd cell_6t
Xbit_r92_c6 bl[6] br[6] wl[92] vdd gnd cell_6t
Xbit_r93_c6 bl[6] br[6] wl[93] vdd gnd cell_6t
Xbit_r94_c6 bl[6] br[6] wl[94] vdd gnd cell_6t
Xbit_r95_c6 bl[6] br[6] wl[95] vdd gnd cell_6t
Xbit_r96_c6 bl[6] br[6] wl[96] vdd gnd cell_6t
Xbit_r97_c6 bl[6] br[6] wl[97] vdd gnd cell_6t
Xbit_r98_c6 bl[6] br[6] wl[98] vdd gnd cell_6t
Xbit_r99_c6 bl[6] br[6] wl[99] vdd gnd cell_6t
Xbit_r100_c6 bl[6] br[6] wl[100] vdd gnd cell_6t
Xbit_r101_c6 bl[6] br[6] wl[101] vdd gnd cell_6t
Xbit_r102_c6 bl[6] br[6] wl[102] vdd gnd cell_6t
Xbit_r103_c6 bl[6] br[6] wl[103] vdd gnd cell_6t
Xbit_r104_c6 bl[6] br[6] wl[104] vdd gnd cell_6t
Xbit_r105_c6 bl[6] br[6] wl[105] vdd gnd cell_6t
Xbit_r106_c6 bl[6] br[6] wl[106] vdd gnd cell_6t
Xbit_r107_c6 bl[6] br[6] wl[107] vdd gnd cell_6t
Xbit_r108_c6 bl[6] br[6] wl[108] vdd gnd cell_6t
Xbit_r109_c6 bl[6] br[6] wl[109] vdd gnd cell_6t
Xbit_r110_c6 bl[6] br[6] wl[110] vdd gnd cell_6t
Xbit_r111_c6 bl[6] br[6] wl[111] vdd gnd cell_6t
Xbit_r112_c6 bl[6] br[6] wl[112] vdd gnd cell_6t
Xbit_r113_c6 bl[6] br[6] wl[113] vdd gnd cell_6t
Xbit_r114_c6 bl[6] br[6] wl[114] vdd gnd cell_6t
Xbit_r115_c6 bl[6] br[6] wl[115] vdd gnd cell_6t
Xbit_r116_c6 bl[6] br[6] wl[116] vdd gnd cell_6t
Xbit_r117_c6 bl[6] br[6] wl[117] vdd gnd cell_6t
Xbit_r118_c6 bl[6] br[6] wl[118] vdd gnd cell_6t
Xbit_r119_c6 bl[6] br[6] wl[119] vdd gnd cell_6t
Xbit_r120_c6 bl[6] br[6] wl[120] vdd gnd cell_6t
Xbit_r121_c6 bl[6] br[6] wl[121] vdd gnd cell_6t
Xbit_r122_c6 bl[6] br[6] wl[122] vdd gnd cell_6t
Xbit_r123_c6 bl[6] br[6] wl[123] vdd gnd cell_6t
Xbit_r124_c6 bl[6] br[6] wl[124] vdd gnd cell_6t
Xbit_r125_c6 bl[6] br[6] wl[125] vdd gnd cell_6t
Xbit_r126_c6 bl[6] br[6] wl[126] vdd gnd cell_6t
Xbit_r127_c6 bl[6] br[6] wl[127] vdd gnd cell_6t
Xbit_r128_c6 bl[6] br[6] wl[128] vdd gnd cell_6t
Xbit_r129_c6 bl[6] br[6] wl[129] vdd gnd cell_6t
Xbit_r130_c6 bl[6] br[6] wl[130] vdd gnd cell_6t
Xbit_r131_c6 bl[6] br[6] wl[131] vdd gnd cell_6t
Xbit_r132_c6 bl[6] br[6] wl[132] vdd gnd cell_6t
Xbit_r133_c6 bl[6] br[6] wl[133] vdd gnd cell_6t
Xbit_r134_c6 bl[6] br[6] wl[134] vdd gnd cell_6t
Xbit_r135_c6 bl[6] br[6] wl[135] vdd gnd cell_6t
Xbit_r136_c6 bl[6] br[6] wl[136] vdd gnd cell_6t
Xbit_r137_c6 bl[6] br[6] wl[137] vdd gnd cell_6t
Xbit_r138_c6 bl[6] br[6] wl[138] vdd gnd cell_6t
Xbit_r139_c6 bl[6] br[6] wl[139] vdd gnd cell_6t
Xbit_r140_c6 bl[6] br[6] wl[140] vdd gnd cell_6t
Xbit_r141_c6 bl[6] br[6] wl[141] vdd gnd cell_6t
Xbit_r142_c6 bl[6] br[6] wl[142] vdd gnd cell_6t
Xbit_r143_c6 bl[6] br[6] wl[143] vdd gnd cell_6t
Xbit_r144_c6 bl[6] br[6] wl[144] vdd gnd cell_6t
Xbit_r145_c6 bl[6] br[6] wl[145] vdd gnd cell_6t
Xbit_r146_c6 bl[6] br[6] wl[146] vdd gnd cell_6t
Xbit_r147_c6 bl[6] br[6] wl[147] vdd gnd cell_6t
Xbit_r148_c6 bl[6] br[6] wl[148] vdd gnd cell_6t
Xbit_r149_c6 bl[6] br[6] wl[149] vdd gnd cell_6t
Xbit_r150_c6 bl[6] br[6] wl[150] vdd gnd cell_6t
Xbit_r151_c6 bl[6] br[6] wl[151] vdd gnd cell_6t
Xbit_r152_c6 bl[6] br[6] wl[152] vdd gnd cell_6t
Xbit_r153_c6 bl[6] br[6] wl[153] vdd gnd cell_6t
Xbit_r154_c6 bl[6] br[6] wl[154] vdd gnd cell_6t
Xbit_r155_c6 bl[6] br[6] wl[155] vdd gnd cell_6t
Xbit_r156_c6 bl[6] br[6] wl[156] vdd gnd cell_6t
Xbit_r157_c6 bl[6] br[6] wl[157] vdd gnd cell_6t
Xbit_r158_c6 bl[6] br[6] wl[158] vdd gnd cell_6t
Xbit_r159_c6 bl[6] br[6] wl[159] vdd gnd cell_6t
Xbit_r160_c6 bl[6] br[6] wl[160] vdd gnd cell_6t
Xbit_r161_c6 bl[6] br[6] wl[161] vdd gnd cell_6t
Xbit_r162_c6 bl[6] br[6] wl[162] vdd gnd cell_6t
Xbit_r163_c6 bl[6] br[6] wl[163] vdd gnd cell_6t
Xbit_r164_c6 bl[6] br[6] wl[164] vdd gnd cell_6t
Xbit_r165_c6 bl[6] br[6] wl[165] vdd gnd cell_6t
Xbit_r166_c6 bl[6] br[6] wl[166] vdd gnd cell_6t
Xbit_r167_c6 bl[6] br[6] wl[167] vdd gnd cell_6t
Xbit_r168_c6 bl[6] br[6] wl[168] vdd gnd cell_6t
Xbit_r169_c6 bl[6] br[6] wl[169] vdd gnd cell_6t
Xbit_r170_c6 bl[6] br[6] wl[170] vdd gnd cell_6t
Xbit_r171_c6 bl[6] br[6] wl[171] vdd gnd cell_6t
Xbit_r172_c6 bl[6] br[6] wl[172] vdd gnd cell_6t
Xbit_r173_c6 bl[6] br[6] wl[173] vdd gnd cell_6t
Xbit_r174_c6 bl[6] br[6] wl[174] vdd gnd cell_6t
Xbit_r175_c6 bl[6] br[6] wl[175] vdd gnd cell_6t
Xbit_r176_c6 bl[6] br[6] wl[176] vdd gnd cell_6t
Xbit_r177_c6 bl[6] br[6] wl[177] vdd gnd cell_6t
Xbit_r178_c6 bl[6] br[6] wl[178] vdd gnd cell_6t
Xbit_r179_c6 bl[6] br[6] wl[179] vdd gnd cell_6t
Xbit_r180_c6 bl[6] br[6] wl[180] vdd gnd cell_6t
Xbit_r181_c6 bl[6] br[6] wl[181] vdd gnd cell_6t
Xbit_r182_c6 bl[6] br[6] wl[182] vdd gnd cell_6t
Xbit_r183_c6 bl[6] br[6] wl[183] vdd gnd cell_6t
Xbit_r184_c6 bl[6] br[6] wl[184] vdd gnd cell_6t
Xbit_r185_c6 bl[6] br[6] wl[185] vdd gnd cell_6t
Xbit_r186_c6 bl[6] br[6] wl[186] vdd gnd cell_6t
Xbit_r187_c6 bl[6] br[6] wl[187] vdd gnd cell_6t
Xbit_r188_c6 bl[6] br[6] wl[188] vdd gnd cell_6t
Xbit_r189_c6 bl[6] br[6] wl[189] vdd gnd cell_6t
Xbit_r190_c6 bl[6] br[6] wl[190] vdd gnd cell_6t
Xbit_r191_c6 bl[6] br[6] wl[191] vdd gnd cell_6t
Xbit_r192_c6 bl[6] br[6] wl[192] vdd gnd cell_6t
Xbit_r193_c6 bl[6] br[6] wl[193] vdd gnd cell_6t
Xbit_r194_c6 bl[6] br[6] wl[194] vdd gnd cell_6t
Xbit_r195_c6 bl[6] br[6] wl[195] vdd gnd cell_6t
Xbit_r196_c6 bl[6] br[6] wl[196] vdd gnd cell_6t
Xbit_r197_c6 bl[6] br[6] wl[197] vdd gnd cell_6t
Xbit_r198_c6 bl[6] br[6] wl[198] vdd gnd cell_6t
Xbit_r199_c6 bl[6] br[6] wl[199] vdd gnd cell_6t
Xbit_r200_c6 bl[6] br[6] wl[200] vdd gnd cell_6t
Xbit_r201_c6 bl[6] br[6] wl[201] vdd gnd cell_6t
Xbit_r202_c6 bl[6] br[6] wl[202] vdd gnd cell_6t
Xbit_r203_c6 bl[6] br[6] wl[203] vdd gnd cell_6t
Xbit_r204_c6 bl[6] br[6] wl[204] vdd gnd cell_6t
Xbit_r205_c6 bl[6] br[6] wl[205] vdd gnd cell_6t
Xbit_r206_c6 bl[6] br[6] wl[206] vdd gnd cell_6t
Xbit_r207_c6 bl[6] br[6] wl[207] vdd gnd cell_6t
Xbit_r208_c6 bl[6] br[6] wl[208] vdd gnd cell_6t
Xbit_r209_c6 bl[6] br[6] wl[209] vdd gnd cell_6t
Xbit_r210_c6 bl[6] br[6] wl[210] vdd gnd cell_6t
Xbit_r211_c6 bl[6] br[6] wl[211] vdd gnd cell_6t
Xbit_r212_c6 bl[6] br[6] wl[212] vdd gnd cell_6t
Xbit_r213_c6 bl[6] br[6] wl[213] vdd gnd cell_6t
Xbit_r214_c6 bl[6] br[6] wl[214] vdd gnd cell_6t
Xbit_r215_c6 bl[6] br[6] wl[215] vdd gnd cell_6t
Xbit_r216_c6 bl[6] br[6] wl[216] vdd gnd cell_6t
Xbit_r217_c6 bl[6] br[6] wl[217] vdd gnd cell_6t
Xbit_r218_c6 bl[6] br[6] wl[218] vdd gnd cell_6t
Xbit_r219_c6 bl[6] br[6] wl[219] vdd gnd cell_6t
Xbit_r220_c6 bl[6] br[6] wl[220] vdd gnd cell_6t
Xbit_r221_c6 bl[6] br[6] wl[221] vdd gnd cell_6t
Xbit_r222_c6 bl[6] br[6] wl[222] vdd gnd cell_6t
Xbit_r223_c6 bl[6] br[6] wl[223] vdd gnd cell_6t
Xbit_r224_c6 bl[6] br[6] wl[224] vdd gnd cell_6t
Xbit_r225_c6 bl[6] br[6] wl[225] vdd gnd cell_6t
Xbit_r226_c6 bl[6] br[6] wl[226] vdd gnd cell_6t
Xbit_r227_c6 bl[6] br[6] wl[227] vdd gnd cell_6t
Xbit_r228_c6 bl[6] br[6] wl[228] vdd gnd cell_6t
Xbit_r229_c6 bl[6] br[6] wl[229] vdd gnd cell_6t
Xbit_r230_c6 bl[6] br[6] wl[230] vdd gnd cell_6t
Xbit_r231_c6 bl[6] br[6] wl[231] vdd gnd cell_6t
Xbit_r232_c6 bl[6] br[6] wl[232] vdd gnd cell_6t
Xbit_r233_c6 bl[6] br[6] wl[233] vdd gnd cell_6t
Xbit_r234_c6 bl[6] br[6] wl[234] vdd gnd cell_6t
Xbit_r235_c6 bl[6] br[6] wl[235] vdd gnd cell_6t
Xbit_r236_c6 bl[6] br[6] wl[236] vdd gnd cell_6t
Xbit_r237_c6 bl[6] br[6] wl[237] vdd gnd cell_6t
Xbit_r238_c6 bl[6] br[6] wl[238] vdd gnd cell_6t
Xbit_r239_c6 bl[6] br[6] wl[239] vdd gnd cell_6t
Xbit_r240_c6 bl[6] br[6] wl[240] vdd gnd cell_6t
Xbit_r241_c6 bl[6] br[6] wl[241] vdd gnd cell_6t
Xbit_r242_c6 bl[6] br[6] wl[242] vdd gnd cell_6t
Xbit_r243_c6 bl[6] br[6] wl[243] vdd gnd cell_6t
Xbit_r244_c6 bl[6] br[6] wl[244] vdd gnd cell_6t
Xbit_r245_c6 bl[6] br[6] wl[245] vdd gnd cell_6t
Xbit_r246_c6 bl[6] br[6] wl[246] vdd gnd cell_6t
Xbit_r247_c6 bl[6] br[6] wl[247] vdd gnd cell_6t
Xbit_r248_c6 bl[6] br[6] wl[248] vdd gnd cell_6t
Xbit_r249_c6 bl[6] br[6] wl[249] vdd gnd cell_6t
Xbit_r250_c6 bl[6] br[6] wl[250] vdd gnd cell_6t
Xbit_r251_c6 bl[6] br[6] wl[251] vdd gnd cell_6t
Xbit_r252_c6 bl[6] br[6] wl[252] vdd gnd cell_6t
Xbit_r253_c6 bl[6] br[6] wl[253] vdd gnd cell_6t
Xbit_r254_c6 bl[6] br[6] wl[254] vdd gnd cell_6t
Xbit_r255_c6 bl[6] br[6] wl[255] vdd gnd cell_6t
Xbit_r256_c6 bl[6] br[6] wl[256] vdd gnd cell_6t
Xbit_r257_c6 bl[6] br[6] wl[257] vdd gnd cell_6t
Xbit_r258_c6 bl[6] br[6] wl[258] vdd gnd cell_6t
Xbit_r259_c6 bl[6] br[6] wl[259] vdd gnd cell_6t
Xbit_r260_c6 bl[6] br[6] wl[260] vdd gnd cell_6t
Xbit_r261_c6 bl[6] br[6] wl[261] vdd gnd cell_6t
Xbit_r262_c6 bl[6] br[6] wl[262] vdd gnd cell_6t
Xbit_r263_c6 bl[6] br[6] wl[263] vdd gnd cell_6t
Xbit_r264_c6 bl[6] br[6] wl[264] vdd gnd cell_6t
Xbit_r265_c6 bl[6] br[6] wl[265] vdd gnd cell_6t
Xbit_r266_c6 bl[6] br[6] wl[266] vdd gnd cell_6t
Xbit_r267_c6 bl[6] br[6] wl[267] vdd gnd cell_6t
Xbit_r268_c6 bl[6] br[6] wl[268] vdd gnd cell_6t
Xbit_r269_c6 bl[6] br[6] wl[269] vdd gnd cell_6t
Xbit_r270_c6 bl[6] br[6] wl[270] vdd gnd cell_6t
Xbit_r271_c6 bl[6] br[6] wl[271] vdd gnd cell_6t
Xbit_r272_c6 bl[6] br[6] wl[272] vdd gnd cell_6t
Xbit_r273_c6 bl[6] br[6] wl[273] vdd gnd cell_6t
Xbit_r274_c6 bl[6] br[6] wl[274] vdd gnd cell_6t
Xbit_r275_c6 bl[6] br[6] wl[275] vdd gnd cell_6t
Xbit_r276_c6 bl[6] br[6] wl[276] vdd gnd cell_6t
Xbit_r277_c6 bl[6] br[6] wl[277] vdd gnd cell_6t
Xbit_r278_c6 bl[6] br[6] wl[278] vdd gnd cell_6t
Xbit_r279_c6 bl[6] br[6] wl[279] vdd gnd cell_6t
Xbit_r280_c6 bl[6] br[6] wl[280] vdd gnd cell_6t
Xbit_r281_c6 bl[6] br[6] wl[281] vdd gnd cell_6t
Xbit_r282_c6 bl[6] br[6] wl[282] vdd gnd cell_6t
Xbit_r283_c6 bl[6] br[6] wl[283] vdd gnd cell_6t
Xbit_r284_c6 bl[6] br[6] wl[284] vdd gnd cell_6t
Xbit_r285_c6 bl[6] br[6] wl[285] vdd gnd cell_6t
Xbit_r286_c6 bl[6] br[6] wl[286] vdd gnd cell_6t
Xbit_r287_c6 bl[6] br[6] wl[287] vdd gnd cell_6t
Xbit_r288_c6 bl[6] br[6] wl[288] vdd gnd cell_6t
Xbit_r289_c6 bl[6] br[6] wl[289] vdd gnd cell_6t
Xbit_r290_c6 bl[6] br[6] wl[290] vdd gnd cell_6t
Xbit_r291_c6 bl[6] br[6] wl[291] vdd gnd cell_6t
Xbit_r292_c6 bl[6] br[6] wl[292] vdd gnd cell_6t
Xbit_r293_c6 bl[6] br[6] wl[293] vdd gnd cell_6t
Xbit_r294_c6 bl[6] br[6] wl[294] vdd gnd cell_6t
Xbit_r295_c6 bl[6] br[6] wl[295] vdd gnd cell_6t
Xbit_r296_c6 bl[6] br[6] wl[296] vdd gnd cell_6t
Xbit_r297_c6 bl[6] br[6] wl[297] vdd gnd cell_6t
Xbit_r298_c6 bl[6] br[6] wl[298] vdd gnd cell_6t
Xbit_r299_c6 bl[6] br[6] wl[299] vdd gnd cell_6t
Xbit_r300_c6 bl[6] br[6] wl[300] vdd gnd cell_6t
Xbit_r301_c6 bl[6] br[6] wl[301] vdd gnd cell_6t
Xbit_r302_c6 bl[6] br[6] wl[302] vdd gnd cell_6t
Xbit_r303_c6 bl[6] br[6] wl[303] vdd gnd cell_6t
Xbit_r304_c6 bl[6] br[6] wl[304] vdd gnd cell_6t
Xbit_r305_c6 bl[6] br[6] wl[305] vdd gnd cell_6t
Xbit_r306_c6 bl[6] br[6] wl[306] vdd gnd cell_6t
Xbit_r307_c6 bl[6] br[6] wl[307] vdd gnd cell_6t
Xbit_r308_c6 bl[6] br[6] wl[308] vdd gnd cell_6t
Xbit_r309_c6 bl[6] br[6] wl[309] vdd gnd cell_6t
Xbit_r310_c6 bl[6] br[6] wl[310] vdd gnd cell_6t
Xbit_r311_c6 bl[6] br[6] wl[311] vdd gnd cell_6t
Xbit_r312_c6 bl[6] br[6] wl[312] vdd gnd cell_6t
Xbit_r313_c6 bl[6] br[6] wl[313] vdd gnd cell_6t
Xbit_r314_c6 bl[6] br[6] wl[314] vdd gnd cell_6t
Xbit_r315_c6 bl[6] br[6] wl[315] vdd gnd cell_6t
Xbit_r316_c6 bl[6] br[6] wl[316] vdd gnd cell_6t
Xbit_r317_c6 bl[6] br[6] wl[317] vdd gnd cell_6t
Xbit_r318_c6 bl[6] br[6] wl[318] vdd gnd cell_6t
Xbit_r319_c6 bl[6] br[6] wl[319] vdd gnd cell_6t
Xbit_r320_c6 bl[6] br[6] wl[320] vdd gnd cell_6t
Xbit_r321_c6 bl[6] br[6] wl[321] vdd gnd cell_6t
Xbit_r322_c6 bl[6] br[6] wl[322] vdd gnd cell_6t
Xbit_r323_c6 bl[6] br[6] wl[323] vdd gnd cell_6t
Xbit_r324_c6 bl[6] br[6] wl[324] vdd gnd cell_6t
Xbit_r325_c6 bl[6] br[6] wl[325] vdd gnd cell_6t
Xbit_r326_c6 bl[6] br[6] wl[326] vdd gnd cell_6t
Xbit_r327_c6 bl[6] br[6] wl[327] vdd gnd cell_6t
Xbit_r328_c6 bl[6] br[6] wl[328] vdd gnd cell_6t
Xbit_r329_c6 bl[6] br[6] wl[329] vdd gnd cell_6t
Xbit_r330_c6 bl[6] br[6] wl[330] vdd gnd cell_6t
Xbit_r331_c6 bl[6] br[6] wl[331] vdd gnd cell_6t
Xbit_r332_c6 bl[6] br[6] wl[332] vdd gnd cell_6t
Xbit_r333_c6 bl[6] br[6] wl[333] vdd gnd cell_6t
Xbit_r334_c6 bl[6] br[6] wl[334] vdd gnd cell_6t
Xbit_r335_c6 bl[6] br[6] wl[335] vdd gnd cell_6t
Xbit_r336_c6 bl[6] br[6] wl[336] vdd gnd cell_6t
Xbit_r337_c6 bl[6] br[6] wl[337] vdd gnd cell_6t
Xbit_r338_c6 bl[6] br[6] wl[338] vdd gnd cell_6t
Xbit_r339_c6 bl[6] br[6] wl[339] vdd gnd cell_6t
Xbit_r340_c6 bl[6] br[6] wl[340] vdd gnd cell_6t
Xbit_r341_c6 bl[6] br[6] wl[341] vdd gnd cell_6t
Xbit_r342_c6 bl[6] br[6] wl[342] vdd gnd cell_6t
Xbit_r343_c6 bl[6] br[6] wl[343] vdd gnd cell_6t
Xbit_r344_c6 bl[6] br[6] wl[344] vdd gnd cell_6t
Xbit_r345_c6 bl[6] br[6] wl[345] vdd gnd cell_6t
Xbit_r346_c6 bl[6] br[6] wl[346] vdd gnd cell_6t
Xbit_r347_c6 bl[6] br[6] wl[347] vdd gnd cell_6t
Xbit_r348_c6 bl[6] br[6] wl[348] vdd gnd cell_6t
Xbit_r349_c6 bl[6] br[6] wl[349] vdd gnd cell_6t
Xbit_r350_c6 bl[6] br[6] wl[350] vdd gnd cell_6t
Xbit_r351_c6 bl[6] br[6] wl[351] vdd gnd cell_6t
Xbit_r352_c6 bl[6] br[6] wl[352] vdd gnd cell_6t
Xbit_r353_c6 bl[6] br[6] wl[353] vdd gnd cell_6t
Xbit_r354_c6 bl[6] br[6] wl[354] vdd gnd cell_6t
Xbit_r355_c6 bl[6] br[6] wl[355] vdd gnd cell_6t
Xbit_r356_c6 bl[6] br[6] wl[356] vdd gnd cell_6t
Xbit_r357_c6 bl[6] br[6] wl[357] vdd gnd cell_6t
Xbit_r358_c6 bl[6] br[6] wl[358] vdd gnd cell_6t
Xbit_r359_c6 bl[6] br[6] wl[359] vdd gnd cell_6t
Xbit_r360_c6 bl[6] br[6] wl[360] vdd gnd cell_6t
Xbit_r361_c6 bl[6] br[6] wl[361] vdd gnd cell_6t
Xbit_r362_c6 bl[6] br[6] wl[362] vdd gnd cell_6t
Xbit_r363_c6 bl[6] br[6] wl[363] vdd gnd cell_6t
Xbit_r364_c6 bl[6] br[6] wl[364] vdd gnd cell_6t
Xbit_r365_c6 bl[6] br[6] wl[365] vdd gnd cell_6t
Xbit_r366_c6 bl[6] br[6] wl[366] vdd gnd cell_6t
Xbit_r367_c6 bl[6] br[6] wl[367] vdd gnd cell_6t
Xbit_r368_c6 bl[6] br[6] wl[368] vdd gnd cell_6t
Xbit_r369_c6 bl[6] br[6] wl[369] vdd gnd cell_6t
Xbit_r370_c6 bl[6] br[6] wl[370] vdd gnd cell_6t
Xbit_r371_c6 bl[6] br[6] wl[371] vdd gnd cell_6t
Xbit_r372_c6 bl[6] br[6] wl[372] vdd gnd cell_6t
Xbit_r373_c6 bl[6] br[6] wl[373] vdd gnd cell_6t
Xbit_r374_c6 bl[6] br[6] wl[374] vdd gnd cell_6t
Xbit_r375_c6 bl[6] br[6] wl[375] vdd gnd cell_6t
Xbit_r376_c6 bl[6] br[6] wl[376] vdd gnd cell_6t
Xbit_r377_c6 bl[6] br[6] wl[377] vdd gnd cell_6t
Xbit_r378_c6 bl[6] br[6] wl[378] vdd gnd cell_6t
Xbit_r379_c6 bl[6] br[6] wl[379] vdd gnd cell_6t
Xbit_r380_c6 bl[6] br[6] wl[380] vdd gnd cell_6t
Xbit_r381_c6 bl[6] br[6] wl[381] vdd gnd cell_6t
Xbit_r382_c6 bl[6] br[6] wl[382] vdd gnd cell_6t
Xbit_r383_c6 bl[6] br[6] wl[383] vdd gnd cell_6t
Xbit_r384_c6 bl[6] br[6] wl[384] vdd gnd cell_6t
Xbit_r385_c6 bl[6] br[6] wl[385] vdd gnd cell_6t
Xbit_r386_c6 bl[6] br[6] wl[386] vdd gnd cell_6t
Xbit_r387_c6 bl[6] br[6] wl[387] vdd gnd cell_6t
Xbit_r388_c6 bl[6] br[6] wl[388] vdd gnd cell_6t
Xbit_r389_c6 bl[6] br[6] wl[389] vdd gnd cell_6t
Xbit_r390_c6 bl[6] br[6] wl[390] vdd gnd cell_6t
Xbit_r391_c6 bl[6] br[6] wl[391] vdd gnd cell_6t
Xbit_r392_c6 bl[6] br[6] wl[392] vdd gnd cell_6t
Xbit_r393_c6 bl[6] br[6] wl[393] vdd gnd cell_6t
Xbit_r394_c6 bl[6] br[6] wl[394] vdd gnd cell_6t
Xbit_r395_c6 bl[6] br[6] wl[395] vdd gnd cell_6t
Xbit_r396_c6 bl[6] br[6] wl[396] vdd gnd cell_6t
Xbit_r397_c6 bl[6] br[6] wl[397] vdd gnd cell_6t
Xbit_r398_c6 bl[6] br[6] wl[398] vdd gnd cell_6t
Xbit_r399_c6 bl[6] br[6] wl[399] vdd gnd cell_6t
Xbit_r400_c6 bl[6] br[6] wl[400] vdd gnd cell_6t
Xbit_r401_c6 bl[6] br[6] wl[401] vdd gnd cell_6t
Xbit_r402_c6 bl[6] br[6] wl[402] vdd gnd cell_6t
Xbit_r403_c6 bl[6] br[6] wl[403] vdd gnd cell_6t
Xbit_r404_c6 bl[6] br[6] wl[404] vdd gnd cell_6t
Xbit_r405_c6 bl[6] br[6] wl[405] vdd gnd cell_6t
Xbit_r406_c6 bl[6] br[6] wl[406] vdd gnd cell_6t
Xbit_r407_c6 bl[6] br[6] wl[407] vdd gnd cell_6t
Xbit_r408_c6 bl[6] br[6] wl[408] vdd gnd cell_6t
Xbit_r409_c6 bl[6] br[6] wl[409] vdd gnd cell_6t
Xbit_r410_c6 bl[6] br[6] wl[410] vdd gnd cell_6t
Xbit_r411_c6 bl[6] br[6] wl[411] vdd gnd cell_6t
Xbit_r412_c6 bl[6] br[6] wl[412] vdd gnd cell_6t
Xbit_r413_c6 bl[6] br[6] wl[413] vdd gnd cell_6t
Xbit_r414_c6 bl[6] br[6] wl[414] vdd gnd cell_6t
Xbit_r415_c6 bl[6] br[6] wl[415] vdd gnd cell_6t
Xbit_r416_c6 bl[6] br[6] wl[416] vdd gnd cell_6t
Xbit_r417_c6 bl[6] br[6] wl[417] vdd gnd cell_6t
Xbit_r418_c6 bl[6] br[6] wl[418] vdd gnd cell_6t
Xbit_r419_c6 bl[6] br[6] wl[419] vdd gnd cell_6t
Xbit_r420_c6 bl[6] br[6] wl[420] vdd gnd cell_6t
Xbit_r421_c6 bl[6] br[6] wl[421] vdd gnd cell_6t
Xbit_r422_c6 bl[6] br[6] wl[422] vdd gnd cell_6t
Xbit_r423_c6 bl[6] br[6] wl[423] vdd gnd cell_6t
Xbit_r424_c6 bl[6] br[6] wl[424] vdd gnd cell_6t
Xbit_r425_c6 bl[6] br[6] wl[425] vdd gnd cell_6t
Xbit_r426_c6 bl[6] br[6] wl[426] vdd gnd cell_6t
Xbit_r427_c6 bl[6] br[6] wl[427] vdd gnd cell_6t
Xbit_r428_c6 bl[6] br[6] wl[428] vdd gnd cell_6t
Xbit_r429_c6 bl[6] br[6] wl[429] vdd gnd cell_6t
Xbit_r430_c6 bl[6] br[6] wl[430] vdd gnd cell_6t
Xbit_r431_c6 bl[6] br[6] wl[431] vdd gnd cell_6t
Xbit_r432_c6 bl[6] br[6] wl[432] vdd gnd cell_6t
Xbit_r433_c6 bl[6] br[6] wl[433] vdd gnd cell_6t
Xbit_r434_c6 bl[6] br[6] wl[434] vdd gnd cell_6t
Xbit_r435_c6 bl[6] br[6] wl[435] vdd gnd cell_6t
Xbit_r436_c6 bl[6] br[6] wl[436] vdd gnd cell_6t
Xbit_r437_c6 bl[6] br[6] wl[437] vdd gnd cell_6t
Xbit_r438_c6 bl[6] br[6] wl[438] vdd gnd cell_6t
Xbit_r439_c6 bl[6] br[6] wl[439] vdd gnd cell_6t
Xbit_r440_c6 bl[6] br[6] wl[440] vdd gnd cell_6t
Xbit_r441_c6 bl[6] br[6] wl[441] vdd gnd cell_6t
Xbit_r442_c6 bl[6] br[6] wl[442] vdd gnd cell_6t
Xbit_r443_c6 bl[6] br[6] wl[443] vdd gnd cell_6t
Xbit_r444_c6 bl[6] br[6] wl[444] vdd gnd cell_6t
Xbit_r445_c6 bl[6] br[6] wl[445] vdd gnd cell_6t
Xbit_r446_c6 bl[6] br[6] wl[446] vdd gnd cell_6t
Xbit_r447_c6 bl[6] br[6] wl[447] vdd gnd cell_6t
Xbit_r448_c6 bl[6] br[6] wl[448] vdd gnd cell_6t
Xbit_r449_c6 bl[6] br[6] wl[449] vdd gnd cell_6t
Xbit_r450_c6 bl[6] br[6] wl[450] vdd gnd cell_6t
Xbit_r451_c6 bl[6] br[6] wl[451] vdd gnd cell_6t
Xbit_r452_c6 bl[6] br[6] wl[452] vdd gnd cell_6t
Xbit_r453_c6 bl[6] br[6] wl[453] vdd gnd cell_6t
Xbit_r454_c6 bl[6] br[6] wl[454] vdd gnd cell_6t
Xbit_r455_c6 bl[6] br[6] wl[455] vdd gnd cell_6t
Xbit_r456_c6 bl[6] br[6] wl[456] vdd gnd cell_6t
Xbit_r457_c6 bl[6] br[6] wl[457] vdd gnd cell_6t
Xbit_r458_c6 bl[6] br[6] wl[458] vdd gnd cell_6t
Xbit_r459_c6 bl[6] br[6] wl[459] vdd gnd cell_6t
Xbit_r460_c6 bl[6] br[6] wl[460] vdd gnd cell_6t
Xbit_r461_c6 bl[6] br[6] wl[461] vdd gnd cell_6t
Xbit_r462_c6 bl[6] br[6] wl[462] vdd gnd cell_6t
Xbit_r463_c6 bl[6] br[6] wl[463] vdd gnd cell_6t
Xbit_r464_c6 bl[6] br[6] wl[464] vdd gnd cell_6t
Xbit_r465_c6 bl[6] br[6] wl[465] vdd gnd cell_6t
Xbit_r466_c6 bl[6] br[6] wl[466] vdd gnd cell_6t
Xbit_r467_c6 bl[6] br[6] wl[467] vdd gnd cell_6t
Xbit_r468_c6 bl[6] br[6] wl[468] vdd gnd cell_6t
Xbit_r469_c6 bl[6] br[6] wl[469] vdd gnd cell_6t
Xbit_r470_c6 bl[6] br[6] wl[470] vdd gnd cell_6t
Xbit_r471_c6 bl[6] br[6] wl[471] vdd gnd cell_6t
Xbit_r472_c6 bl[6] br[6] wl[472] vdd gnd cell_6t
Xbit_r473_c6 bl[6] br[6] wl[473] vdd gnd cell_6t
Xbit_r474_c6 bl[6] br[6] wl[474] vdd gnd cell_6t
Xbit_r475_c6 bl[6] br[6] wl[475] vdd gnd cell_6t
Xbit_r476_c6 bl[6] br[6] wl[476] vdd gnd cell_6t
Xbit_r477_c6 bl[6] br[6] wl[477] vdd gnd cell_6t
Xbit_r478_c6 bl[6] br[6] wl[478] vdd gnd cell_6t
Xbit_r479_c6 bl[6] br[6] wl[479] vdd gnd cell_6t
Xbit_r480_c6 bl[6] br[6] wl[480] vdd gnd cell_6t
Xbit_r481_c6 bl[6] br[6] wl[481] vdd gnd cell_6t
Xbit_r482_c6 bl[6] br[6] wl[482] vdd gnd cell_6t
Xbit_r483_c6 bl[6] br[6] wl[483] vdd gnd cell_6t
Xbit_r484_c6 bl[6] br[6] wl[484] vdd gnd cell_6t
Xbit_r485_c6 bl[6] br[6] wl[485] vdd gnd cell_6t
Xbit_r486_c6 bl[6] br[6] wl[486] vdd gnd cell_6t
Xbit_r487_c6 bl[6] br[6] wl[487] vdd gnd cell_6t
Xbit_r488_c6 bl[6] br[6] wl[488] vdd gnd cell_6t
Xbit_r489_c6 bl[6] br[6] wl[489] vdd gnd cell_6t
Xbit_r490_c6 bl[6] br[6] wl[490] vdd gnd cell_6t
Xbit_r491_c6 bl[6] br[6] wl[491] vdd gnd cell_6t
Xbit_r492_c6 bl[6] br[6] wl[492] vdd gnd cell_6t
Xbit_r493_c6 bl[6] br[6] wl[493] vdd gnd cell_6t
Xbit_r494_c6 bl[6] br[6] wl[494] vdd gnd cell_6t
Xbit_r495_c6 bl[6] br[6] wl[495] vdd gnd cell_6t
Xbit_r496_c6 bl[6] br[6] wl[496] vdd gnd cell_6t
Xbit_r497_c6 bl[6] br[6] wl[497] vdd gnd cell_6t
Xbit_r498_c6 bl[6] br[6] wl[498] vdd gnd cell_6t
Xbit_r499_c6 bl[6] br[6] wl[499] vdd gnd cell_6t
Xbit_r500_c6 bl[6] br[6] wl[500] vdd gnd cell_6t
Xbit_r501_c6 bl[6] br[6] wl[501] vdd gnd cell_6t
Xbit_r502_c6 bl[6] br[6] wl[502] vdd gnd cell_6t
Xbit_r503_c6 bl[6] br[6] wl[503] vdd gnd cell_6t
Xbit_r504_c6 bl[6] br[6] wl[504] vdd gnd cell_6t
Xbit_r505_c6 bl[6] br[6] wl[505] vdd gnd cell_6t
Xbit_r506_c6 bl[6] br[6] wl[506] vdd gnd cell_6t
Xbit_r507_c6 bl[6] br[6] wl[507] vdd gnd cell_6t
Xbit_r508_c6 bl[6] br[6] wl[508] vdd gnd cell_6t
Xbit_r509_c6 bl[6] br[6] wl[509] vdd gnd cell_6t
Xbit_r510_c6 bl[6] br[6] wl[510] vdd gnd cell_6t
Xbit_r511_c6 bl[6] br[6] wl[511] vdd gnd cell_6t
Xbit_r0_c7 bl[7] br[7] wl[0] vdd gnd cell_6t
Xbit_r1_c7 bl[7] br[7] wl[1] vdd gnd cell_6t
Xbit_r2_c7 bl[7] br[7] wl[2] vdd gnd cell_6t
Xbit_r3_c7 bl[7] br[7] wl[3] vdd gnd cell_6t
Xbit_r4_c7 bl[7] br[7] wl[4] vdd gnd cell_6t
Xbit_r5_c7 bl[7] br[7] wl[5] vdd gnd cell_6t
Xbit_r6_c7 bl[7] br[7] wl[6] vdd gnd cell_6t
Xbit_r7_c7 bl[7] br[7] wl[7] vdd gnd cell_6t
Xbit_r8_c7 bl[7] br[7] wl[8] vdd gnd cell_6t
Xbit_r9_c7 bl[7] br[7] wl[9] vdd gnd cell_6t
Xbit_r10_c7 bl[7] br[7] wl[10] vdd gnd cell_6t
Xbit_r11_c7 bl[7] br[7] wl[11] vdd gnd cell_6t
Xbit_r12_c7 bl[7] br[7] wl[12] vdd gnd cell_6t
Xbit_r13_c7 bl[7] br[7] wl[13] vdd gnd cell_6t
Xbit_r14_c7 bl[7] br[7] wl[14] vdd gnd cell_6t
Xbit_r15_c7 bl[7] br[7] wl[15] vdd gnd cell_6t
Xbit_r16_c7 bl[7] br[7] wl[16] vdd gnd cell_6t
Xbit_r17_c7 bl[7] br[7] wl[17] vdd gnd cell_6t
Xbit_r18_c7 bl[7] br[7] wl[18] vdd gnd cell_6t
Xbit_r19_c7 bl[7] br[7] wl[19] vdd gnd cell_6t
Xbit_r20_c7 bl[7] br[7] wl[20] vdd gnd cell_6t
Xbit_r21_c7 bl[7] br[7] wl[21] vdd gnd cell_6t
Xbit_r22_c7 bl[7] br[7] wl[22] vdd gnd cell_6t
Xbit_r23_c7 bl[7] br[7] wl[23] vdd gnd cell_6t
Xbit_r24_c7 bl[7] br[7] wl[24] vdd gnd cell_6t
Xbit_r25_c7 bl[7] br[7] wl[25] vdd gnd cell_6t
Xbit_r26_c7 bl[7] br[7] wl[26] vdd gnd cell_6t
Xbit_r27_c7 bl[7] br[7] wl[27] vdd gnd cell_6t
Xbit_r28_c7 bl[7] br[7] wl[28] vdd gnd cell_6t
Xbit_r29_c7 bl[7] br[7] wl[29] vdd gnd cell_6t
Xbit_r30_c7 bl[7] br[7] wl[30] vdd gnd cell_6t
Xbit_r31_c7 bl[7] br[7] wl[31] vdd gnd cell_6t
Xbit_r32_c7 bl[7] br[7] wl[32] vdd gnd cell_6t
Xbit_r33_c7 bl[7] br[7] wl[33] vdd gnd cell_6t
Xbit_r34_c7 bl[7] br[7] wl[34] vdd gnd cell_6t
Xbit_r35_c7 bl[7] br[7] wl[35] vdd gnd cell_6t
Xbit_r36_c7 bl[7] br[7] wl[36] vdd gnd cell_6t
Xbit_r37_c7 bl[7] br[7] wl[37] vdd gnd cell_6t
Xbit_r38_c7 bl[7] br[7] wl[38] vdd gnd cell_6t
Xbit_r39_c7 bl[7] br[7] wl[39] vdd gnd cell_6t
Xbit_r40_c7 bl[7] br[7] wl[40] vdd gnd cell_6t
Xbit_r41_c7 bl[7] br[7] wl[41] vdd gnd cell_6t
Xbit_r42_c7 bl[7] br[7] wl[42] vdd gnd cell_6t
Xbit_r43_c7 bl[7] br[7] wl[43] vdd gnd cell_6t
Xbit_r44_c7 bl[7] br[7] wl[44] vdd gnd cell_6t
Xbit_r45_c7 bl[7] br[7] wl[45] vdd gnd cell_6t
Xbit_r46_c7 bl[7] br[7] wl[46] vdd gnd cell_6t
Xbit_r47_c7 bl[7] br[7] wl[47] vdd gnd cell_6t
Xbit_r48_c7 bl[7] br[7] wl[48] vdd gnd cell_6t
Xbit_r49_c7 bl[7] br[7] wl[49] vdd gnd cell_6t
Xbit_r50_c7 bl[7] br[7] wl[50] vdd gnd cell_6t
Xbit_r51_c7 bl[7] br[7] wl[51] vdd gnd cell_6t
Xbit_r52_c7 bl[7] br[7] wl[52] vdd gnd cell_6t
Xbit_r53_c7 bl[7] br[7] wl[53] vdd gnd cell_6t
Xbit_r54_c7 bl[7] br[7] wl[54] vdd gnd cell_6t
Xbit_r55_c7 bl[7] br[7] wl[55] vdd gnd cell_6t
Xbit_r56_c7 bl[7] br[7] wl[56] vdd gnd cell_6t
Xbit_r57_c7 bl[7] br[7] wl[57] vdd gnd cell_6t
Xbit_r58_c7 bl[7] br[7] wl[58] vdd gnd cell_6t
Xbit_r59_c7 bl[7] br[7] wl[59] vdd gnd cell_6t
Xbit_r60_c7 bl[7] br[7] wl[60] vdd gnd cell_6t
Xbit_r61_c7 bl[7] br[7] wl[61] vdd gnd cell_6t
Xbit_r62_c7 bl[7] br[7] wl[62] vdd gnd cell_6t
Xbit_r63_c7 bl[7] br[7] wl[63] vdd gnd cell_6t
Xbit_r64_c7 bl[7] br[7] wl[64] vdd gnd cell_6t
Xbit_r65_c7 bl[7] br[7] wl[65] vdd gnd cell_6t
Xbit_r66_c7 bl[7] br[7] wl[66] vdd gnd cell_6t
Xbit_r67_c7 bl[7] br[7] wl[67] vdd gnd cell_6t
Xbit_r68_c7 bl[7] br[7] wl[68] vdd gnd cell_6t
Xbit_r69_c7 bl[7] br[7] wl[69] vdd gnd cell_6t
Xbit_r70_c7 bl[7] br[7] wl[70] vdd gnd cell_6t
Xbit_r71_c7 bl[7] br[7] wl[71] vdd gnd cell_6t
Xbit_r72_c7 bl[7] br[7] wl[72] vdd gnd cell_6t
Xbit_r73_c7 bl[7] br[7] wl[73] vdd gnd cell_6t
Xbit_r74_c7 bl[7] br[7] wl[74] vdd gnd cell_6t
Xbit_r75_c7 bl[7] br[7] wl[75] vdd gnd cell_6t
Xbit_r76_c7 bl[7] br[7] wl[76] vdd gnd cell_6t
Xbit_r77_c7 bl[7] br[7] wl[77] vdd gnd cell_6t
Xbit_r78_c7 bl[7] br[7] wl[78] vdd gnd cell_6t
Xbit_r79_c7 bl[7] br[7] wl[79] vdd gnd cell_6t
Xbit_r80_c7 bl[7] br[7] wl[80] vdd gnd cell_6t
Xbit_r81_c7 bl[7] br[7] wl[81] vdd gnd cell_6t
Xbit_r82_c7 bl[7] br[7] wl[82] vdd gnd cell_6t
Xbit_r83_c7 bl[7] br[7] wl[83] vdd gnd cell_6t
Xbit_r84_c7 bl[7] br[7] wl[84] vdd gnd cell_6t
Xbit_r85_c7 bl[7] br[7] wl[85] vdd gnd cell_6t
Xbit_r86_c7 bl[7] br[7] wl[86] vdd gnd cell_6t
Xbit_r87_c7 bl[7] br[7] wl[87] vdd gnd cell_6t
Xbit_r88_c7 bl[7] br[7] wl[88] vdd gnd cell_6t
Xbit_r89_c7 bl[7] br[7] wl[89] vdd gnd cell_6t
Xbit_r90_c7 bl[7] br[7] wl[90] vdd gnd cell_6t
Xbit_r91_c7 bl[7] br[7] wl[91] vdd gnd cell_6t
Xbit_r92_c7 bl[7] br[7] wl[92] vdd gnd cell_6t
Xbit_r93_c7 bl[7] br[7] wl[93] vdd gnd cell_6t
Xbit_r94_c7 bl[7] br[7] wl[94] vdd gnd cell_6t
Xbit_r95_c7 bl[7] br[7] wl[95] vdd gnd cell_6t
Xbit_r96_c7 bl[7] br[7] wl[96] vdd gnd cell_6t
Xbit_r97_c7 bl[7] br[7] wl[97] vdd gnd cell_6t
Xbit_r98_c7 bl[7] br[7] wl[98] vdd gnd cell_6t
Xbit_r99_c7 bl[7] br[7] wl[99] vdd gnd cell_6t
Xbit_r100_c7 bl[7] br[7] wl[100] vdd gnd cell_6t
Xbit_r101_c7 bl[7] br[7] wl[101] vdd gnd cell_6t
Xbit_r102_c7 bl[7] br[7] wl[102] vdd gnd cell_6t
Xbit_r103_c7 bl[7] br[7] wl[103] vdd gnd cell_6t
Xbit_r104_c7 bl[7] br[7] wl[104] vdd gnd cell_6t
Xbit_r105_c7 bl[7] br[7] wl[105] vdd gnd cell_6t
Xbit_r106_c7 bl[7] br[7] wl[106] vdd gnd cell_6t
Xbit_r107_c7 bl[7] br[7] wl[107] vdd gnd cell_6t
Xbit_r108_c7 bl[7] br[7] wl[108] vdd gnd cell_6t
Xbit_r109_c7 bl[7] br[7] wl[109] vdd gnd cell_6t
Xbit_r110_c7 bl[7] br[7] wl[110] vdd gnd cell_6t
Xbit_r111_c7 bl[7] br[7] wl[111] vdd gnd cell_6t
Xbit_r112_c7 bl[7] br[7] wl[112] vdd gnd cell_6t
Xbit_r113_c7 bl[7] br[7] wl[113] vdd gnd cell_6t
Xbit_r114_c7 bl[7] br[7] wl[114] vdd gnd cell_6t
Xbit_r115_c7 bl[7] br[7] wl[115] vdd gnd cell_6t
Xbit_r116_c7 bl[7] br[7] wl[116] vdd gnd cell_6t
Xbit_r117_c7 bl[7] br[7] wl[117] vdd gnd cell_6t
Xbit_r118_c7 bl[7] br[7] wl[118] vdd gnd cell_6t
Xbit_r119_c7 bl[7] br[7] wl[119] vdd gnd cell_6t
Xbit_r120_c7 bl[7] br[7] wl[120] vdd gnd cell_6t
Xbit_r121_c7 bl[7] br[7] wl[121] vdd gnd cell_6t
Xbit_r122_c7 bl[7] br[7] wl[122] vdd gnd cell_6t
Xbit_r123_c7 bl[7] br[7] wl[123] vdd gnd cell_6t
Xbit_r124_c7 bl[7] br[7] wl[124] vdd gnd cell_6t
Xbit_r125_c7 bl[7] br[7] wl[125] vdd gnd cell_6t
Xbit_r126_c7 bl[7] br[7] wl[126] vdd gnd cell_6t
Xbit_r127_c7 bl[7] br[7] wl[127] vdd gnd cell_6t
Xbit_r128_c7 bl[7] br[7] wl[128] vdd gnd cell_6t
Xbit_r129_c7 bl[7] br[7] wl[129] vdd gnd cell_6t
Xbit_r130_c7 bl[7] br[7] wl[130] vdd gnd cell_6t
Xbit_r131_c7 bl[7] br[7] wl[131] vdd gnd cell_6t
Xbit_r132_c7 bl[7] br[7] wl[132] vdd gnd cell_6t
Xbit_r133_c7 bl[7] br[7] wl[133] vdd gnd cell_6t
Xbit_r134_c7 bl[7] br[7] wl[134] vdd gnd cell_6t
Xbit_r135_c7 bl[7] br[7] wl[135] vdd gnd cell_6t
Xbit_r136_c7 bl[7] br[7] wl[136] vdd gnd cell_6t
Xbit_r137_c7 bl[7] br[7] wl[137] vdd gnd cell_6t
Xbit_r138_c7 bl[7] br[7] wl[138] vdd gnd cell_6t
Xbit_r139_c7 bl[7] br[7] wl[139] vdd gnd cell_6t
Xbit_r140_c7 bl[7] br[7] wl[140] vdd gnd cell_6t
Xbit_r141_c7 bl[7] br[7] wl[141] vdd gnd cell_6t
Xbit_r142_c7 bl[7] br[7] wl[142] vdd gnd cell_6t
Xbit_r143_c7 bl[7] br[7] wl[143] vdd gnd cell_6t
Xbit_r144_c7 bl[7] br[7] wl[144] vdd gnd cell_6t
Xbit_r145_c7 bl[7] br[7] wl[145] vdd gnd cell_6t
Xbit_r146_c7 bl[7] br[7] wl[146] vdd gnd cell_6t
Xbit_r147_c7 bl[7] br[7] wl[147] vdd gnd cell_6t
Xbit_r148_c7 bl[7] br[7] wl[148] vdd gnd cell_6t
Xbit_r149_c7 bl[7] br[7] wl[149] vdd gnd cell_6t
Xbit_r150_c7 bl[7] br[7] wl[150] vdd gnd cell_6t
Xbit_r151_c7 bl[7] br[7] wl[151] vdd gnd cell_6t
Xbit_r152_c7 bl[7] br[7] wl[152] vdd gnd cell_6t
Xbit_r153_c7 bl[7] br[7] wl[153] vdd gnd cell_6t
Xbit_r154_c7 bl[7] br[7] wl[154] vdd gnd cell_6t
Xbit_r155_c7 bl[7] br[7] wl[155] vdd gnd cell_6t
Xbit_r156_c7 bl[7] br[7] wl[156] vdd gnd cell_6t
Xbit_r157_c7 bl[7] br[7] wl[157] vdd gnd cell_6t
Xbit_r158_c7 bl[7] br[7] wl[158] vdd gnd cell_6t
Xbit_r159_c7 bl[7] br[7] wl[159] vdd gnd cell_6t
Xbit_r160_c7 bl[7] br[7] wl[160] vdd gnd cell_6t
Xbit_r161_c7 bl[7] br[7] wl[161] vdd gnd cell_6t
Xbit_r162_c7 bl[7] br[7] wl[162] vdd gnd cell_6t
Xbit_r163_c7 bl[7] br[7] wl[163] vdd gnd cell_6t
Xbit_r164_c7 bl[7] br[7] wl[164] vdd gnd cell_6t
Xbit_r165_c7 bl[7] br[7] wl[165] vdd gnd cell_6t
Xbit_r166_c7 bl[7] br[7] wl[166] vdd gnd cell_6t
Xbit_r167_c7 bl[7] br[7] wl[167] vdd gnd cell_6t
Xbit_r168_c7 bl[7] br[7] wl[168] vdd gnd cell_6t
Xbit_r169_c7 bl[7] br[7] wl[169] vdd gnd cell_6t
Xbit_r170_c7 bl[7] br[7] wl[170] vdd gnd cell_6t
Xbit_r171_c7 bl[7] br[7] wl[171] vdd gnd cell_6t
Xbit_r172_c7 bl[7] br[7] wl[172] vdd gnd cell_6t
Xbit_r173_c7 bl[7] br[7] wl[173] vdd gnd cell_6t
Xbit_r174_c7 bl[7] br[7] wl[174] vdd gnd cell_6t
Xbit_r175_c7 bl[7] br[7] wl[175] vdd gnd cell_6t
Xbit_r176_c7 bl[7] br[7] wl[176] vdd gnd cell_6t
Xbit_r177_c7 bl[7] br[7] wl[177] vdd gnd cell_6t
Xbit_r178_c7 bl[7] br[7] wl[178] vdd gnd cell_6t
Xbit_r179_c7 bl[7] br[7] wl[179] vdd gnd cell_6t
Xbit_r180_c7 bl[7] br[7] wl[180] vdd gnd cell_6t
Xbit_r181_c7 bl[7] br[7] wl[181] vdd gnd cell_6t
Xbit_r182_c7 bl[7] br[7] wl[182] vdd gnd cell_6t
Xbit_r183_c7 bl[7] br[7] wl[183] vdd gnd cell_6t
Xbit_r184_c7 bl[7] br[7] wl[184] vdd gnd cell_6t
Xbit_r185_c7 bl[7] br[7] wl[185] vdd gnd cell_6t
Xbit_r186_c7 bl[7] br[7] wl[186] vdd gnd cell_6t
Xbit_r187_c7 bl[7] br[7] wl[187] vdd gnd cell_6t
Xbit_r188_c7 bl[7] br[7] wl[188] vdd gnd cell_6t
Xbit_r189_c7 bl[7] br[7] wl[189] vdd gnd cell_6t
Xbit_r190_c7 bl[7] br[7] wl[190] vdd gnd cell_6t
Xbit_r191_c7 bl[7] br[7] wl[191] vdd gnd cell_6t
Xbit_r192_c7 bl[7] br[7] wl[192] vdd gnd cell_6t
Xbit_r193_c7 bl[7] br[7] wl[193] vdd gnd cell_6t
Xbit_r194_c7 bl[7] br[7] wl[194] vdd gnd cell_6t
Xbit_r195_c7 bl[7] br[7] wl[195] vdd gnd cell_6t
Xbit_r196_c7 bl[7] br[7] wl[196] vdd gnd cell_6t
Xbit_r197_c7 bl[7] br[7] wl[197] vdd gnd cell_6t
Xbit_r198_c7 bl[7] br[7] wl[198] vdd gnd cell_6t
Xbit_r199_c7 bl[7] br[7] wl[199] vdd gnd cell_6t
Xbit_r200_c7 bl[7] br[7] wl[200] vdd gnd cell_6t
Xbit_r201_c7 bl[7] br[7] wl[201] vdd gnd cell_6t
Xbit_r202_c7 bl[7] br[7] wl[202] vdd gnd cell_6t
Xbit_r203_c7 bl[7] br[7] wl[203] vdd gnd cell_6t
Xbit_r204_c7 bl[7] br[7] wl[204] vdd gnd cell_6t
Xbit_r205_c7 bl[7] br[7] wl[205] vdd gnd cell_6t
Xbit_r206_c7 bl[7] br[7] wl[206] vdd gnd cell_6t
Xbit_r207_c7 bl[7] br[7] wl[207] vdd gnd cell_6t
Xbit_r208_c7 bl[7] br[7] wl[208] vdd gnd cell_6t
Xbit_r209_c7 bl[7] br[7] wl[209] vdd gnd cell_6t
Xbit_r210_c7 bl[7] br[7] wl[210] vdd gnd cell_6t
Xbit_r211_c7 bl[7] br[7] wl[211] vdd gnd cell_6t
Xbit_r212_c7 bl[7] br[7] wl[212] vdd gnd cell_6t
Xbit_r213_c7 bl[7] br[7] wl[213] vdd gnd cell_6t
Xbit_r214_c7 bl[7] br[7] wl[214] vdd gnd cell_6t
Xbit_r215_c7 bl[7] br[7] wl[215] vdd gnd cell_6t
Xbit_r216_c7 bl[7] br[7] wl[216] vdd gnd cell_6t
Xbit_r217_c7 bl[7] br[7] wl[217] vdd gnd cell_6t
Xbit_r218_c7 bl[7] br[7] wl[218] vdd gnd cell_6t
Xbit_r219_c7 bl[7] br[7] wl[219] vdd gnd cell_6t
Xbit_r220_c7 bl[7] br[7] wl[220] vdd gnd cell_6t
Xbit_r221_c7 bl[7] br[7] wl[221] vdd gnd cell_6t
Xbit_r222_c7 bl[7] br[7] wl[222] vdd gnd cell_6t
Xbit_r223_c7 bl[7] br[7] wl[223] vdd gnd cell_6t
Xbit_r224_c7 bl[7] br[7] wl[224] vdd gnd cell_6t
Xbit_r225_c7 bl[7] br[7] wl[225] vdd gnd cell_6t
Xbit_r226_c7 bl[7] br[7] wl[226] vdd gnd cell_6t
Xbit_r227_c7 bl[7] br[7] wl[227] vdd gnd cell_6t
Xbit_r228_c7 bl[7] br[7] wl[228] vdd gnd cell_6t
Xbit_r229_c7 bl[7] br[7] wl[229] vdd gnd cell_6t
Xbit_r230_c7 bl[7] br[7] wl[230] vdd gnd cell_6t
Xbit_r231_c7 bl[7] br[7] wl[231] vdd gnd cell_6t
Xbit_r232_c7 bl[7] br[7] wl[232] vdd gnd cell_6t
Xbit_r233_c7 bl[7] br[7] wl[233] vdd gnd cell_6t
Xbit_r234_c7 bl[7] br[7] wl[234] vdd gnd cell_6t
Xbit_r235_c7 bl[7] br[7] wl[235] vdd gnd cell_6t
Xbit_r236_c7 bl[7] br[7] wl[236] vdd gnd cell_6t
Xbit_r237_c7 bl[7] br[7] wl[237] vdd gnd cell_6t
Xbit_r238_c7 bl[7] br[7] wl[238] vdd gnd cell_6t
Xbit_r239_c7 bl[7] br[7] wl[239] vdd gnd cell_6t
Xbit_r240_c7 bl[7] br[7] wl[240] vdd gnd cell_6t
Xbit_r241_c7 bl[7] br[7] wl[241] vdd gnd cell_6t
Xbit_r242_c7 bl[7] br[7] wl[242] vdd gnd cell_6t
Xbit_r243_c7 bl[7] br[7] wl[243] vdd gnd cell_6t
Xbit_r244_c7 bl[7] br[7] wl[244] vdd gnd cell_6t
Xbit_r245_c7 bl[7] br[7] wl[245] vdd gnd cell_6t
Xbit_r246_c7 bl[7] br[7] wl[246] vdd gnd cell_6t
Xbit_r247_c7 bl[7] br[7] wl[247] vdd gnd cell_6t
Xbit_r248_c7 bl[7] br[7] wl[248] vdd gnd cell_6t
Xbit_r249_c7 bl[7] br[7] wl[249] vdd gnd cell_6t
Xbit_r250_c7 bl[7] br[7] wl[250] vdd gnd cell_6t
Xbit_r251_c7 bl[7] br[7] wl[251] vdd gnd cell_6t
Xbit_r252_c7 bl[7] br[7] wl[252] vdd gnd cell_6t
Xbit_r253_c7 bl[7] br[7] wl[253] vdd gnd cell_6t
Xbit_r254_c7 bl[7] br[7] wl[254] vdd gnd cell_6t
Xbit_r255_c7 bl[7] br[7] wl[255] vdd gnd cell_6t
Xbit_r256_c7 bl[7] br[7] wl[256] vdd gnd cell_6t
Xbit_r257_c7 bl[7] br[7] wl[257] vdd gnd cell_6t
Xbit_r258_c7 bl[7] br[7] wl[258] vdd gnd cell_6t
Xbit_r259_c7 bl[7] br[7] wl[259] vdd gnd cell_6t
Xbit_r260_c7 bl[7] br[7] wl[260] vdd gnd cell_6t
Xbit_r261_c7 bl[7] br[7] wl[261] vdd gnd cell_6t
Xbit_r262_c7 bl[7] br[7] wl[262] vdd gnd cell_6t
Xbit_r263_c7 bl[7] br[7] wl[263] vdd gnd cell_6t
Xbit_r264_c7 bl[7] br[7] wl[264] vdd gnd cell_6t
Xbit_r265_c7 bl[7] br[7] wl[265] vdd gnd cell_6t
Xbit_r266_c7 bl[7] br[7] wl[266] vdd gnd cell_6t
Xbit_r267_c7 bl[7] br[7] wl[267] vdd gnd cell_6t
Xbit_r268_c7 bl[7] br[7] wl[268] vdd gnd cell_6t
Xbit_r269_c7 bl[7] br[7] wl[269] vdd gnd cell_6t
Xbit_r270_c7 bl[7] br[7] wl[270] vdd gnd cell_6t
Xbit_r271_c7 bl[7] br[7] wl[271] vdd gnd cell_6t
Xbit_r272_c7 bl[7] br[7] wl[272] vdd gnd cell_6t
Xbit_r273_c7 bl[7] br[7] wl[273] vdd gnd cell_6t
Xbit_r274_c7 bl[7] br[7] wl[274] vdd gnd cell_6t
Xbit_r275_c7 bl[7] br[7] wl[275] vdd gnd cell_6t
Xbit_r276_c7 bl[7] br[7] wl[276] vdd gnd cell_6t
Xbit_r277_c7 bl[7] br[7] wl[277] vdd gnd cell_6t
Xbit_r278_c7 bl[7] br[7] wl[278] vdd gnd cell_6t
Xbit_r279_c7 bl[7] br[7] wl[279] vdd gnd cell_6t
Xbit_r280_c7 bl[7] br[7] wl[280] vdd gnd cell_6t
Xbit_r281_c7 bl[7] br[7] wl[281] vdd gnd cell_6t
Xbit_r282_c7 bl[7] br[7] wl[282] vdd gnd cell_6t
Xbit_r283_c7 bl[7] br[7] wl[283] vdd gnd cell_6t
Xbit_r284_c7 bl[7] br[7] wl[284] vdd gnd cell_6t
Xbit_r285_c7 bl[7] br[7] wl[285] vdd gnd cell_6t
Xbit_r286_c7 bl[7] br[7] wl[286] vdd gnd cell_6t
Xbit_r287_c7 bl[7] br[7] wl[287] vdd gnd cell_6t
Xbit_r288_c7 bl[7] br[7] wl[288] vdd gnd cell_6t
Xbit_r289_c7 bl[7] br[7] wl[289] vdd gnd cell_6t
Xbit_r290_c7 bl[7] br[7] wl[290] vdd gnd cell_6t
Xbit_r291_c7 bl[7] br[7] wl[291] vdd gnd cell_6t
Xbit_r292_c7 bl[7] br[7] wl[292] vdd gnd cell_6t
Xbit_r293_c7 bl[7] br[7] wl[293] vdd gnd cell_6t
Xbit_r294_c7 bl[7] br[7] wl[294] vdd gnd cell_6t
Xbit_r295_c7 bl[7] br[7] wl[295] vdd gnd cell_6t
Xbit_r296_c7 bl[7] br[7] wl[296] vdd gnd cell_6t
Xbit_r297_c7 bl[7] br[7] wl[297] vdd gnd cell_6t
Xbit_r298_c7 bl[7] br[7] wl[298] vdd gnd cell_6t
Xbit_r299_c7 bl[7] br[7] wl[299] vdd gnd cell_6t
Xbit_r300_c7 bl[7] br[7] wl[300] vdd gnd cell_6t
Xbit_r301_c7 bl[7] br[7] wl[301] vdd gnd cell_6t
Xbit_r302_c7 bl[7] br[7] wl[302] vdd gnd cell_6t
Xbit_r303_c7 bl[7] br[7] wl[303] vdd gnd cell_6t
Xbit_r304_c7 bl[7] br[7] wl[304] vdd gnd cell_6t
Xbit_r305_c7 bl[7] br[7] wl[305] vdd gnd cell_6t
Xbit_r306_c7 bl[7] br[7] wl[306] vdd gnd cell_6t
Xbit_r307_c7 bl[7] br[7] wl[307] vdd gnd cell_6t
Xbit_r308_c7 bl[7] br[7] wl[308] vdd gnd cell_6t
Xbit_r309_c7 bl[7] br[7] wl[309] vdd gnd cell_6t
Xbit_r310_c7 bl[7] br[7] wl[310] vdd gnd cell_6t
Xbit_r311_c7 bl[7] br[7] wl[311] vdd gnd cell_6t
Xbit_r312_c7 bl[7] br[7] wl[312] vdd gnd cell_6t
Xbit_r313_c7 bl[7] br[7] wl[313] vdd gnd cell_6t
Xbit_r314_c7 bl[7] br[7] wl[314] vdd gnd cell_6t
Xbit_r315_c7 bl[7] br[7] wl[315] vdd gnd cell_6t
Xbit_r316_c7 bl[7] br[7] wl[316] vdd gnd cell_6t
Xbit_r317_c7 bl[7] br[7] wl[317] vdd gnd cell_6t
Xbit_r318_c7 bl[7] br[7] wl[318] vdd gnd cell_6t
Xbit_r319_c7 bl[7] br[7] wl[319] vdd gnd cell_6t
Xbit_r320_c7 bl[7] br[7] wl[320] vdd gnd cell_6t
Xbit_r321_c7 bl[7] br[7] wl[321] vdd gnd cell_6t
Xbit_r322_c7 bl[7] br[7] wl[322] vdd gnd cell_6t
Xbit_r323_c7 bl[7] br[7] wl[323] vdd gnd cell_6t
Xbit_r324_c7 bl[7] br[7] wl[324] vdd gnd cell_6t
Xbit_r325_c7 bl[7] br[7] wl[325] vdd gnd cell_6t
Xbit_r326_c7 bl[7] br[7] wl[326] vdd gnd cell_6t
Xbit_r327_c7 bl[7] br[7] wl[327] vdd gnd cell_6t
Xbit_r328_c7 bl[7] br[7] wl[328] vdd gnd cell_6t
Xbit_r329_c7 bl[7] br[7] wl[329] vdd gnd cell_6t
Xbit_r330_c7 bl[7] br[7] wl[330] vdd gnd cell_6t
Xbit_r331_c7 bl[7] br[7] wl[331] vdd gnd cell_6t
Xbit_r332_c7 bl[7] br[7] wl[332] vdd gnd cell_6t
Xbit_r333_c7 bl[7] br[7] wl[333] vdd gnd cell_6t
Xbit_r334_c7 bl[7] br[7] wl[334] vdd gnd cell_6t
Xbit_r335_c7 bl[7] br[7] wl[335] vdd gnd cell_6t
Xbit_r336_c7 bl[7] br[7] wl[336] vdd gnd cell_6t
Xbit_r337_c7 bl[7] br[7] wl[337] vdd gnd cell_6t
Xbit_r338_c7 bl[7] br[7] wl[338] vdd gnd cell_6t
Xbit_r339_c7 bl[7] br[7] wl[339] vdd gnd cell_6t
Xbit_r340_c7 bl[7] br[7] wl[340] vdd gnd cell_6t
Xbit_r341_c7 bl[7] br[7] wl[341] vdd gnd cell_6t
Xbit_r342_c7 bl[7] br[7] wl[342] vdd gnd cell_6t
Xbit_r343_c7 bl[7] br[7] wl[343] vdd gnd cell_6t
Xbit_r344_c7 bl[7] br[7] wl[344] vdd gnd cell_6t
Xbit_r345_c7 bl[7] br[7] wl[345] vdd gnd cell_6t
Xbit_r346_c7 bl[7] br[7] wl[346] vdd gnd cell_6t
Xbit_r347_c7 bl[7] br[7] wl[347] vdd gnd cell_6t
Xbit_r348_c7 bl[7] br[7] wl[348] vdd gnd cell_6t
Xbit_r349_c7 bl[7] br[7] wl[349] vdd gnd cell_6t
Xbit_r350_c7 bl[7] br[7] wl[350] vdd gnd cell_6t
Xbit_r351_c7 bl[7] br[7] wl[351] vdd gnd cell_6t
Xbit_r352_c7 bl[7] br[7] wl[352] vdd gnd cell_6t
Xbit_r353_c7 bl[7] br[7] wl[353] vdd gnd cell_6t
Xbit_r354_c7 bl[7] br[7] wl[354] vdd gnd cell_6t
Xbit_r355_c7 bl[7] br[7] wl[355] vdd gnd cell_6t
Xbit_r356_c7 bl[7] br[7] wl[356] vdd gnd cell_6t
Xbit_r357_c7 bl[7] br[7] wl[357] vdd gnd cell_6t
Xbit_r358_c7 bl[7] br[7] wl[358] vdd gnd cell_6t
Xbit_r359_c7 bl[7] br[7] wl[359] vdd gnd cell_6t
Xbit_r360_c7 bl[7] br[7] wl[360] vdd gnd cell_6t
Xbit_r361_c7 bl[7] br[7] wl[361] vdd gnd cell_6t
Xbit_r362_c7 bl[7] br[7] wl[362] vdd gnd cell_6t
Xbit_r363_c7 bl[7] br[7] wl[363] vdd gnd cell_6t
Xbit_r364_c7 bl[7] br[7] wl[364] vdd gnd cell_6t
Xbit_r365_c7 bl[7] br[7] wl[365] vdd gnd cell_6t
Xbit_r366_c7 bl[7] br[7] wl[366] vdd gnd cell_6t
Xbit_r367_c7 bl[7] br[7] wl[367] vdd gnd cell_6t
Xbit_r368_c7 bl[7] br[7] wl[368] vdd gnd cell_6t
Xbit_r369_c7 bl[7] br[7] wl[369] vdd gnd cell_6t
Xbit_r370_c7 bl[7] br[7] wl[370] vdd gnd cell_6t
Xbit_r371_c7 bl[7] br[7] wl[371] vdd gnd cell_6t
Xbit_r372_c7 bl[7] br[7] wl[372] vdd gnd cell_6t
Xbit_r373_c7 bl[7] br[7] wl[373] vdd gnd cell_6t
Xbit_r374_c7 bl[7] br[7] wl[374] vdd gnd cell_6t
Xbit_r375_c7 bl[7] br[7] wl[375] vdd gnd cell_6t
Xbit_r376_c7 bl[7] br[7] wl[376] vdd gnd cell_6t
Xbit_r377_c7 bl[7] br[7] wl[377] vdd gnd cell_6t
Xbit_r378_c7 bl[7] br[7] wl[378] vdd gnd cell_6t
Xbit_r379_c7 bl[7] br[7] wl[379] vdd gnd cell_6t
Xbit_r380_c7 bl[7] br[7] wl[380] vdd gnd cell_6t
Xbit_r381_c7 bl[7] br[7] wl[381] vdd gnd cell_6t
Xbit_r382_c7 bl[7] br[7] wl[382] vdd gnd cell_6t
Xbit_r383_c7 bl[7] br[7] wl[383] vdd gnd cell_6t
Xbit_r384_c7 bl[7] br[7] wl[384] vdd gnd cell_6t
Xbit_r385_c7 bl[7] br[7] wl[385] vdd gnd cell_6t
Xbit_r386_c7 bl[7] br[7] wl[386] vdd gnd cell_6t
Xbit_r387_c7 bl[7] br[7] wl[387] vdd gnd cell_6t
Xbit_r388_c7 bl[7] br[7] wl[388] vdd gnd cell_6t
Xbit_r389_c7 bl[7] br[7] wl[389] vdd gnd cell_6t
Xbit_r390_c7 bl[7] br[7] wl[390] vdd gnd cell_6t
Xbit_r391_c7 bl[7] br[7] wl[391] vdd gnd cell_6t
Xbit_r392_c7 bl[7] br[7] wl[392] vdd gnd cell_6t
Xbit_r393_c7 bl[7] br[7] wl[393] vdd gnd cell_6t
Xbit_r394_c7 bl[7] br[7] wl[394] vdd gnd cell_6t
Xbit_r395_c7 bl[7] br[7] wl[395] vdd gnd cell_6t
Xbit_r396_c7 bl[7] br[7] wl[396] vdd gnd cell_6t
Xbit_r397_c7 bl[7] br[7] wl[397] vdd gnd cell_6t
Xbit_r398_c7 bl[7] br[7] wl[398] vdd gnd cell_6t
Xbit_r399_c7 bl[7] br[7] wl[399] vdd gnd cell_6t
Xbit_r400_c7 bl[7] br[7] wl[400] vdd gnd cell_6t
Xbit_r401_c7 bl[7] br[7] wl[401] vdd gnd cell_6t
Xbit_r402_c7 bl[7] br[7] wl[402] vdd gnd cell_6t
Xbit_r403_c7 bl[7] br[7] wl[403] vdd gnd cell_6t
Xbit_r404_c7 bl[7] br[7] wl[404] vdd gnd cell_6t
Xbit_r405_c7 bl[7] br[7] wl[405] vdd gnd cell_6t
Xbit_r406_c7 bl[7] br[7] wl[406] vdd gnd cell_6t
Xbit_r407_c7 bl[7] br[7] wl[407] vdd gnd cell_6t
Xbit_r408_c7 bl[7] br[7] wl[408] vdd gnd cell_6t
Xbit_r409_c7 bl[7] br[7] wl[409] vdd gnd cell_6t
Xbit_r410_c7 bl[7] br[7] wl[410] vdd gnd cell_6t
Xbit_r411_c7 bl[7] br[7] wl[411] vdd gnd cell_6t
Xbit_r412_c7 bl[7] br[7] wl[412] vdd gnd cell_6t
Xbit_r413_c7 bl[7] br[7] wl[413] vdd gnd cell_6t
Xbit_r414_c7 bl[7] br[7] wl[414] vdd gnd cell_6t
Xbit_r415_c7 bl[7] br[7] wl[415] vdd gnd cell_6t
Xbit_r416_c7 bl[7] br[7] wl[416] vdd gnd cell_6t
Xbit_r417_c7 bl[7] br[7] wl[417] vdd gnd cell_6t
Xbit_r418_c7 bl[7] br[7] wl[418] vdd gnd cell_6t
Xbit_r419_c7 bl[7] br[7] wl[419] vdd gnd cell_6t
Xbit_r420_c7 bl[7] br[7] wl[420] vdd gnd cell_6t
Xbit_r421_c7 bl[7] br[7] wl[421] vdd gnd cell_6t
Xbit_r422_c7 bl[7] br[7] wl[422] vdd gnd cell_6t
Xbit_r423_c7 bl[7] br[7] wl[423] vdd gnd cell_6t
Xbit_r424_c7 bl[7] br[7] wl[424] vdd gnd cell_6t
Xbit_r425_c7 bl[7] br[7] wl[425] vdd gnd cell_6t
Xbit_r426_c7 bl[7] br[7] wl[426] vdd gnd cell_6t
Xbit_r427_c7 bl[7] br[7] wl[427] vdd gnd cell_6t
Xbit_r428_c7 bl[7] br[7] wl[428] vdd gnd cell_6t
Xbit_r429_c7 bl[7] br[7] wl[429] vdd gnd cell_6t
Xbit_r430_c7 bl[7] br[7] wl[430] vdd gnd cell_6t
Xbit_r431_c7 bl[7] br[7] wl[431] vdd gnd cell_6t
Xbit_r432_c7 bl[7] br[7] wl[432] vdd gnd cell_6t
Xbit_r433_c7 bl[7] br[7] wl[433] vdd gnd cell_6t
Xbit_r434_c7 bl[7] br[7] wl[434] vdd gnd cell_6t
Xbit_r435_c7 bl[7] br[7] wl[435] vdd gnd cell_6t
Xbit_r436_c7 bl[7] br[7] wl[436] vdd gnd cell_6t
Xbit_r437_c7 bl[7] br[7] wl[437] vdd gnd cell_6t
Xbit_r438_c7 bl[7] br[7] wl[438] vdd gnd cell_6t
Xbit_r439_c7 bl[7] br[7] wl[439] vdd gnd cell_6t
Xbit_r440_c7 bl[7] br[7] wl[440] vdd gnd cell_6t
Xbit_r441_c7 bl[7] br[7] wl[441] vdd gnd cell_6t
Xbit_r442_c7 bl[7] br[7] wl[442] vdd gnd cell_6t
Xbit_r443_c7 bl[7] br[7] wl[443] vdd gnd cell_6t
Xbit_r444_c7 bl[7] br[7] wl[444] vdd gnd cell_6t
Xbit_r445_c7 bl[7] br[7] wl[445] vdd gnd cell_6t
Xbit_r446_c7 bl[7] br[7] wl[446] vdd gnd cell_6t
Xbit_r447_c7 bl[7] br[7] wl[447] vdd gnd cell_6t
Xbit_r448_c7 bl[7] br[7] wl[448] vdd gnd cell_6t
Xbit_r449_c7 bl[7] br[7] wl[449] vdd gnd cell_6t
Xbit_r450_c7 bl[7] br[7] wl[450] vdd gnd cell_6t
Xbit_r451_c7 bl[7] br[7] wl[451] vdd gnd cell_6t
Xbit_r452_c7 bl[7] br[7] wl[452] vdd gnd cell_6t
Xbit_r453_c7 bl[7] br[7] wl[453] vdd gnd cell_6t
Xbit_r454_c7 bl[7] br[7] wl[454] vdd gnd cell_6t
Xbit_r455_c7 bl[7] br[7] wl[455] vdd gnd cell_6t
Xbit_r456_c7 bl[7] br[7] wl[456] vdd gnd cell_6t
Xbit_r457_c7 bl[7] br[7] wl[457] vdd gnd cell_6t
Xbit_r458_c7 bl[7] br[7] wl[458] vdd gnd cell_6t
Xbit_r459_c7 bl[7] br[7] wl[459] vdd gnd cell_6t
Xbit_r460_c7 bl[7] br[7] wl[460] vdd gnd cell_6t
Xbit_r461_c7 bl[7] br[7] wl[461] vdd gnd cell_6t
Xbit_r462_c7 bl[7] br[7] wl[462] vdd gnd cell_6t
Xbit_r463_c7 bl[7] br[7] wl[463] vdd gnd cell_6t
Xbit_r464_c7 bl[7] br[7] wl[464] vdd gnd cell_6t
Xbit_r465_c7 bl[7] br[7] wl[465] vdd gnd cell_6t
Xbit_r466_c7 bl[7] br[7] wl[466] vdd gnd cell_6t
Xbit_r467_c7 bl[7] br[7] wl[467] vdd gnd cell_6t
Xbit_r468_c7 bl[7] br[7] wl[468] vdd gnd cell_6t
Xbit_r469_c7 bl[7] br[7] wl[469] vdd gnd cell_6t
Xbit_r470_c7 bl[7] br[7] wl[470] vdd gnd cell_6t
Xbit_r471_c7 bl[7] br[7] wl[471] vdd gnd cell_6t
Xbit_r472_c7 bl[7] br[7] wl[472] vdd gnd cell_6t
Xbit_r473_c7 bl[7] br[7] wl[473] vdd gnd cell_6t
Xbit_r474_c7 bl[7] br[7] wl[474] vdd gnd cell_6t
Xbit_r475_c7 bl[7] br[7] wl[475] vdd gnd cell_6t
Xbit_r476_c7 bl[7] br[7] wl[476] vdd gnd cell_6t
Xbit_r477_c7 bl[7] br[7] wl[477] vdd gnd cell_6t
Xbit_r478_c7 bl[7] br[7] wl[478] vdd gnd cell_6t
Xbit_r479_c7 bl[7] br[7] wl[479] vdd gnd cell_6t
Xbit_r480_c7 bl[7] br[7] wl[480] vdd gnd cell_6t
Xbit_r481_c7 bl[7] br[7] wl[481] vdd gnd cell_6t
Xbit_r482_c7 bl[7] br[7] wl[482] vdd gnd cell_6t
Xbit_r483_c7 bl[7] br[7] wl[483] vdd gnd cell_6t
Xbit_r484_c7 bl[7] br[7] wl[484] vdd gnd cell_6t
Xbit_r485_c7 bl[7] br[7] wl[485] vdd gnd cell_6t
Xbit_r486_c7 bl[7] br[7] wl[486] vdd gnd cell_6t
Xbit_r487_c7 bl[7] br[7] wl[487] vdd gnd cell_6t
Xbit_r488_c7 bl[7] br[7] wl[488] vdd gnd cell_6t
Xbit_r489_c7 bl[7] br[7] wl[489] vdd gnd cell_6t
Xbit_r490_c7 bl[7] br[7] wl[490] vdd gnd cell_6t
Xbit_r491_c7 bl[7] br[7] wl[491] vdd gnd cell_6t
Xbit_r492_c7 bl[7] br[7] wl[492] vdd gnd cell_6t
Xbit_r493_c7 bl[7] br[7] wl[493] vdd gnd cell_6t
Xbit_r494_c7 bl[7] br[7] wl[494] vdd gnd cell_6t
Xbit_r495_c7 bl[7] br[7] wl[495] vdd gnd cell_6t
Xbit_r496_c7 bl[7] br[7] wl[496] vdd gnd cell_6t
Xbit_r497_c7 bl[7] br[7] wl[497] vdd gnd cell_6t
Xbit_r498_c7 bl[7] br[7] wl[498] vdd gnd cell_6t
Xbit_r499_c7 bl[7] br[7] wl[499] vdd gnd cell_6t
Xbit_r500_c7 bl[7] br[7] wl[500] vdd gnd cell_6t
Xbit_r501_c7 bl[7] br[7] wl[501] vdd gnd cell_6t
Xbit_r502_c7 bl[7] br[7] wl[502] vdd gnd cell_6t
Xbit_r503_c7 bl[7] br[7] wl[503] vdd gnd cell_6t
Xbit_r504_c7 bl[7] br[7] wl[504] vdd gnd cell_6t
Xbit_r505_c7 bl[7] br[7] wl[505] vdd gnd cell_6t
Xbit_r506_c7 bl[7] br[7] wl[506] vdd gnd cell_6t
Xbit_r507_c7 bl[7] br[7] wl[507] vdd gnd cell_6t
Xbit_r508_c7 bl[7] br[7] wl[508] vdd gnd cell_6t
Xbit_r509_c7 bl[7] br[7] wl[509] vdd gnd cell_6t
Xbit_r510_c7 bl[7] br[7] wl[510] vdd gnd cell_6t
Xbit_r511_c7 bl[7] br[7] wl[511] vdd gnd cell_6t
Xbit_r0_c8 bl[8] br[8] wl[0] vdd gnd cell_6t
Xbit_r1_c8 bl[8] br[8] wl[1] vdd gnd cell_6t
Xbit_r2_c8 bl[8] br[8] wl[2] vdd gnd cell_6t
Xbit_r3_c8 bl[8] br[8] wl[3] vdd gnd cell_6t
Xbit_r4_c8 bl[8] br[8] wl[4] vdd gnd cell_6t
Xbit_r5_c8 bl[8] br[8] wl[5] vdd gnd cell_6t
Xbit_r6_c8 bl[8] br[8] wl[6] vdd gnd cell_6t
Xbit_r7_c8 bl[8] br[8] wl[7] vdd gnd cell_6t
Xbit_r8_c8 bl[8] br[8] wl[8] vdd gnd cell_6t
Xbit_r9_c8 bl[8] br[8] wl[9] vdd gnd cell_6t
Xbit_r10_c8 bl[8] br[8] wl[10] vdd gnd cell_6t
Xbit_r11_c8 bl[8] br[8] wl[11] vdd gnd cell_6t
Xbit_r12_c8 bl[8] br[8] wl[12] vdd gnd cell_6t
Xbit_r13_c8 bl[8] br[8] wl[13] vdd gnd cell_6t
Xbit_r14_c8 bl[8] br[8] wl[14] vdd gnd cell_6t
Xbit_r15_c8 bl[8] br[8] wl[15] vdd gnd cell_6t
Xbit_r16_c8 bl[8] br[8] wl[16] vdd gnd cell_6t
Xbit_r17_c8 bl[8] br[8] wl[17] vdd gnd cell_6t
Xbit_r18_c8 bl[8] br[8] wl[18] vdd gnd cell_6t
Xbit_r19_c8 bl[8] br[8] wl[19] vdd gnd cell_6t
Xbit_r20_c8 bl[8] br[8] wl[20] vdd gnd cell_6t
Xbit_r21_c8 bl[8] br[8] wl[21] vdd gnd cell_6t
Xbit_r22_c8 bl[8] br[8] wl[22] vdd gnd cell_6t
Xbit_r23_c8 bl[8] br[8] wl[23] vdd gnd cell_6t
Xbit_r24_c8 bl[8] br[8] wl[24] vdd gnd cell_6t
Xbit_r25_c8 bl[8] br[8] wl[25] vdd gnd cell_6t
Xbit_r26_c8 bl[8] br[8] wl[26] vdd gnd cell_6t
Xbit_r27_c8 bl[8] br[8] wl[27] vdd gnd cell_6t
Xbit_r28_c8 bl[8] br[8] wl[28] vdd gnd cell_6t
Xbit_r29_c8 bl[8] br[8] wl[29] vdd gnd cell_6t
Xbit_r30_c8 bl[8] br[8] wl[30] vdd gnd cell_6t
Xbit_r31_c8 bl[8] br[8] wl[31] vdd gnd cell_6t
Xbit_r32_c8 bl[8] br[8] wl[32] vdd gnd cell_6t
Xbit_r33_c8 bl[8] br[8] wl[33] vdd gnd cell_6t
Xbit_r34_c8 bl[8] br[8] wl[34] vdd gnd cell_6t
Xbit_r35_c8 bl[8] br[8] wl[35] vdd gnd cell_6t
Xbit_r36_c8 bl[8] br[8] wl[36] vdd gnd cell_6t
Xbit_r37_c8 bl[8] br[8] wl[37] vdd gnd cell_6t
Xbit_r38_c8 bl[8] br[8] wl[38] vdd gnd cell_6t
Xbit_r39_c8 bl[8] br[8] wl[39] vdd gnd cell_6t
Xbit_r40_c8 bl[8] br[8] wl[40] vdd gnd cell_6t
Xbit_r41_c8 bl[8] br[8] wl[41] vdd gnd cell_6t
Xbit_r42_c8 bl[8] br[8] wl[42] vdd gnd cell_6t
Xbit_r43_c8 bl[8] br[8] wl[43] vdd gnd cell_6t
Xbit_r44_c8 bl[8] br[8] wl[44] vdd gnd cell_6t
Xbit_r45_c8 bl[8] br[8] wl[45] vdd gnd cell_6t
Xbit_r46_c8 bl[8] br[8] wl[46] vdd gnd cell_6t
Xbit_r47_c8 bl[8] br[8] wl[47] vdd gnd cell_6t
Xbit_r48_c8 bl[8] br[8] wl[48] vdd gnd cell_6t
Xbit_r49_c8 bl[8] br[8] wl[49] vdd gnd cell_6t
Xbit_r50_c8 bl[8] br[8] wl[50] vdd gnd cell_6t
Xbit_r51_c8 bl[8] br[8] wl[51] vdd gnd cell_6t
Xbit_r52_c8 bl[8] br[8] wl[52] vdd gnd cell_6t
Xbit_r53_c8 bl[8] br[8] wl[53] vdd gnd cell_6t
Xbit_r54_c8 bl[8] br[8] wl[54] vdd gnd cell_6t
Xbit_r55_c8 bl[8] br[8] wl[55] vdd gnd cell_6t
Xbit_r56_c8 bl[8] br[8] wl[56] vdd gnd cell_6t
Xbit_r57_c8 bl[8] br[8] wl[57] vdd gnd cell_6t
Xbit_r58_c8 bl[8] br[8] wl[58] vdd gnd cell_6t
Xbit_r59_c8 bl[8] br[8] wl[59] vdd gnd cell_6t
Xbit_r60_c8 bl[8] br[8] wl[60] vdd gnd cell_6t
Xbit_r61_c8 bl[8] br[8] wl[61] vdd gnd cell_6t
Xbit_r62_c8 bl[8] br[8] wl[62] vdd gnd cell_6t
Xbit_r63_c8 bl[8] br[8] wl[63] vdd gnd cell_6t
Xbit_r64_c8 bl[8] br[8] wl[64] vdd gnd cell_6t
Xbit_r65_c8 bl[8] br[8] wl[65] vdd gnd cell_6t
Xbit_r66_c8 bl[8] br[8] wl[66] vdd gnd cell_6t
Xbit_r67_c8 bl[8] br[8] wl[67] vdd gnd cell_6t
Xbit_r68_c8 bl[8] br[8] wl[68] vdd gnd cell_6t
Xbit_r69_c8 bl[8] br[8] wl[69] vdd gnd cell_6t
Xbit_r70_c8 bl[8] br[8] wl[70] vdd gnd cell_6t
Xbit_r71_c8 bl[8] br[8] wl[71] vdd gnd cell_6t
Xbit_r72_c8 bl[8] br[8] wl[72] vdd gnd cell_6t
Xbit_r73_c8 bl[8] br[8] wl[73] vdd gnd cell_6t
Xbit_r74_c8 bl[8] br[8] wl[74] vdd gnd cell_6t
Xbit_r75_c8 bl[8] br[8] wl[75] vdd gnd cell_6t
Xbit_r76_c8 bl[8] br[8] wl[76] vdd gnd cell_6t
Xbit_r77_c8 bl[8] br[8] wl[77] vdd gnd cell_6t
Xbit_r78_c8 bl[8] br[8] wl[78] vdd gnd cell_6t
Xbit_r79_c8 bl[8] br[8] wl[79] vdd gnd cell_6t
Xbit_r80_c8 bl[8] br[8] wl[80] vdd gnd cell_6t
Xbit_r81_c8 bl[8] br[8] wl[81] vdd gnd cell_6t
Xbit_r82_c8 bl[8] br[8] wl[82] vdd gnd cell_6t
Xbit_r83_c8 bl[8] br[8] wl[83] vdd gnd cell_6t
Xbit_r84_c8 bl[8] br[8] wl[84] vdd gnd cell_6t
Xbit_r85_c8 bl[8] br[8] wl[85] vdd gnd cell_6t
Xbit_r86_c8 bl[8] br[8] wl[86] vdd gnd cell_6t
Xbit_r87_c8 bl[8] br[8] wl[87] vdd gnd cell_6t
Xbit_r88_c8 bl[8] br[8] wl[88] vdd gnd cell_6t
Xbit_r89_c8 bl[8] br[8] wl[89] vdd gnd cell_6t
Xbit_r90_c8 bl[8] br[8] wl[90] vdd gnd cell_6t
Xbit_r91_c8 bl[8] br[8] wl[91] vdd gnd cell_6t
Xbit_r92_c8 bl[8] br[8] wl[92] vdd gnd cell_6t
Xbit_r93_c8 bl[8] br[8] wl[93] vdd gnd cell_6t
Xbit_r94_c8 bl[8] br[8] wl[94] vdd gnd cell_6t
Xbit_r95_c8 bl[8] br[8] wl[95] vdd gnd cell_6t
Xbit_r96_c8 bl[8] br[8] wl[96] vdd gnd cell_6t
Xbit_r97_c8 bl[8] br[8] wl[97] vdd gnd cell_6t
Xbit_r98_c8 bl[8] br[8] wl[98] vdd gnd cell_6t
Xbit_r99_c8 bl[8] br[8] wl[99] vdd gnd cell_6t
Xbit_r100_c8 bl[8] br[8] wl[100] vdd gnd cell_6t
Xbit_r101_c8 bl[8] br[8] wl[101] vdd gnd cell_6t
Xbit_r102_c8 bl[8] br[8] wl[102] vdd gnd cell_6t
Xbit_r103_c8 bl[8] br[8] wl[103] vdd gnd cell_6t
Xbit_r104_c8 bl[8] br[8] wl[104] vdd gnd cell_6t
Xbit_r105_c8 bl[8] br[8] wl[105] vdd gnd cell_6t
Xbit_r106_c8 bl[8] br[8] wl[106] vdd gnd cell_6t
Xbit_r107_c8 bl[8] br[8] wl[107] vdd gnd cell_6t
Xbit_r108_c8 bl[8] br[8] wl[108] vdd gnd cell_6t
Xbit_r109_c8 bl[8] br[8] wl[109] vdd gnd cell_6t
Xbit_r110_c8 bl[8] br[8] wl[110] vdd gnd cell_6t
Xbit_r111_c8 bl[8] br[8] wl[111] vdd gnd cell_6t
Xbit_r112_c8 bl[8] br[8] wl[112] vdd gnd cell_6t
Xbit_r113_c8 bl[8] br[8] wl[113] vdd gnd cell_6t
Xbit_r114_c8 bl[8] br[8] wl[114] vdd gnd cell_6t
Xbit_r115_c8 bl[8] br[8] wl[115] vdd gnd cell_6t
Xbit_r116_c8 bl[8] br[8] wl[116] vdd gnd cell_6t
Xbit_r117_c8 bl[8] br[8] wl[117] vdd gnd cell_6t
Xbit_r118_c8 bl[8] br[8] wl[118] vdd gnd cell_6t
Xbit_r119_c8 bl[8] br[8] wl[119] vdd gnd cell_6t
Xbit_r120_c8 bl[8] br[8] wl[120] vdd gnd cell_6t
Xbit_r121_c8 bl[8] br[8] wl[121] vdd gnd cell_6t
Xbit_r122_c8 bl[8] br[8] wl[122] vdd gnd cell_6t
Xbit_r123_c8 bl[8] br[8] wl[123] vdd gnd cell_6t
Xbit_r124_c8 bl[8] br[8] wl[124] vdd gnd cell_6t
Xbit_r125_c8 bl[8] br[8] wl[125] vdd gnd cell_6t
Xbit_r126_c8 bl[8] br[8] wl[126] vdd gnd cell_6t
Xbit_r127_c8 bl[8] br[8] wl[127] vdd gnd cell_6t
Xbit_r128_c8 bl[8] br[8] wl[128] vdd gnd cell_6t
Xbit_r129_c8 bl[8] br[8] wl[129] vdd gnd cell_6t
Xbit_r130_c8 bl[8] br[8] wl[130] vdd gnd cell_6t
Xbit_r131_c8 bl[8] br[8] wl[131] vdd gnd cell_6t
Xbit_r132_c8 bl[8] br[8] wl[132] vdd gnd cell_6t
Xbit_r133_c8 bl[8] br[8] wl[133] vdd gnd cell_6t
Xbit_r134_c8 bl[8] br[8] wl[134] vdd gnd cell_6t
Xbit_r135_c8 bl[8] br[8] wl[135] vdd gnd cell_6t
Xbit_r136_c8 bl[8] br[8] wl[136] vdd gnd cell_6t
Xbit_r137_c8 bl[8] br[8] wl[137] vdd gnd cell_6t
Xbit_r138_c8 bl[8] br[8] wl[138] vdd gnd cell_6t
Xbit_r139_c8 bl[8] br[8] wl[139] vdd gnd cell_6t
Xbit_r140_c8 bl[8] br[8] wl[140] vdd gnd cell_6t
Xbit_r141_c8 bl[8] br[8] wl[141] vdd gnd cell_6t
Xbit_r142_c8 bl[8] br[8] wl[142] vdd gnd cell_6t
Xbit_r143_c8 bl[8] br[8] wl[143] vdd gnd cell_6t
Xbit_r144_c8 bl[8] br[8] wl[144] vdd gnd cell_6t
Xbit_r145_c8 bl[8] br[8] wl[145] vdd gnd cell_6t
Xbit_r146_c8 bl[8] br[8] wl[146] vdd gnd cell_6t
Xbit_r147_c8 bl[8] br[8] wl[147] vdd gnd cell_6t
Xbit_r148_c8 bl[8] br[8] wl[148] vdd gnd cell_6t
Xbit_r149_c8 bl[8] br[8] wl[149] vdd gnd cell_6t
Xbit_r150_c8 bl[8] br[8] wl[150] vdd gnd cell_6t
Xbit_r151_c8 bl[8] br[8] wl[151] vdd gnd cell_6t
Xbit_r152_c8 bl[8] br[8] wl[152] vdd gnd cell_6t
Xbit_r153_c8 bl[8] br[8] wl[153] vdd gnd cell_6t
Xbit_r154_c8 bl[8] br[8] wl[154] vdd gnd cell_6t
Xbit_r155_c8 bl[8] br[8] wl[155] vdd gnd cell_6t
Xbit_r156_c8 bl[8] br[8] wl[156] vdd gnd cell_6t
Xbit_r157_c8 bl[8] br[8] wl[157] vdd gnd cell_6t
Xbit_r158_c8 bl[8] br[8] wl[158] vdd gnd cell_6t
Xbit_r159_c8 bl[8] br[8] wl[159] vdd gnd cell_6t
Xbit_r160_c8 bl[8] br[8] wl[160] vdd gnd cell_6t
Xbit_r161_c8 bl[8] br[8] wl[161] vdd gnd cell_6t
Xbit_r162_c8 bl[8] br[8] wl[162] vdd gnd cell_6t
Xbit_r163_c8 bl[8] br[8] wl[163] vdd gnd cell_6t
Xbit_r164_c8 bl[8] br[8] wl[164] vdd gnd cell_6t
Xbit_r165_c8 bl[8] br[8] wl[165] vdd gnd cell_6t
Xbit_r166_c8 bl[8] br[8] wl[166] vdd gnd cell_6t
Xbit_r167_c8 bl[8] br[8] wl[167] vdd gnd cell_6t
Xbit_r168_c8 bl[8] br[8] wl[168] vdd gnd cell_6t
Xbit_r169_c8 bl[8] br[8] wl[169] vdd gnd cell_6t
Xbit_r170_c8 bl[8] br[8] wl[170] vdd gnd cell_6t
Xbit_r171_c8 bl[8] br[8] wl[171] vdd gnd cell_6t
Xbit_r172_c8 bl[8] br[8] wl[172] vdd gnd cell_6t
Xbit_r173_c8 bl[8] br[8] wl[173] vdd gnd cell_6t
Xbit_r174_c8 bl[8] br[8] wl[174] vdd gnd cell_6t
Xbit_r175_c8 bl[8] br[8] wl[175] vdd gnd cell_6t
Xbit_r176_c8 bl[8] br[8] wl[176] vdd gnd cell_6t
Xbit_r177_c8 bl[8] br[8] wl[177] vdd gnd cell_6t
Xbit_r178_c8 bl[8] br[8] wl[178] vdd gnd cell_6t
Xbit_r179_c8 bl[8] br[8] wl[179] vdd gnd cell_6t
Xbit_r180_c8 bl[8] br[8] wl[180] vdd gnd cell_6t
Xbit_r181_c8 bl[8] br[8] wl[181] vdd gnd cell_6t
Xbit_r182_c8 bl[8] br[8] wl[182] vdd gnd cell_6t
Xbit_r183_c8 bl[8] br[8] wl[183] vdd gnd cell_6t
Xbit_r184_c8 bl[8] br[8] wl[184] vdd gnd cell_6t
Xbit_r185_c8 bl[8] br[8] wl[185] vdd gnd cell_6t
Xbit_r186_c8 bl[8] br[8] wl[186] vdd gnd cell_6t
Xbit_r187_c8 bl[8] br[8] wl[187] vdd gnd cell_6t
Xbit_r188_c8 bl[8] br[8] wl[188] vdd gnd cell_6t
Xbit_r189_c8 bl[8] br[8] wl[189] vdd gnd cell_6t
Xbit_r190_c8 bl[8] br[8] wl[190] vdd gnd cell_6t
Xbit_r191_c8 bl[8] br[8] wl[191] vdd gnd cell_6t
Xbit_r192_c8 bl[8] br[8] wl[192] vdd gnd cell_6t
Xbit_r193_c8 bl[8] br[8] wl[193] vdd gnd cell_6t
Xbit_r194_c8 bl[8] br[8] wl[194] vdd gnd cell_6t
Xbit_r195_c8 bl[8] br[8] wl[195] vdd gnd cell_6t
Xbit_r196_c8 bl[8] br[8] wl[196] vdd gnd cell_6t
Xbit_r197_c8 bl[8] br[8] wl[197] vdd gnd cell_6t
Xbit_r198_c8 bl[8] br[8] wl[198] vdd gnd cell_6t
Xbit_r199_c8 bl[8] br[8] wl[199] vdd gnd cell_6t
Xbit_r200_c8 bl[8] br[8] wl[200] vdd gnd cell_6t
Xbit_r201_c8 bl[8] br[8] wl[201] vdd gnd cell_6t
Xbit_r202_c8 bl[8] br[8] wl[202] vdd gnd cell_6t
Xbit_r203_c8 bl[8] br[8] wl[203] vdd gnd cell_6t
Xbit_r204_c8 bl[8] br[8] wl[204] vdd gnd cell_6t
Xbit_r205_c8 bl[8] br[8] wl[205] vdd gnd cell_6t
Xbit_r206_c8 bl[8] br[8] wl[206] vdd gnd cell_6t
Xbit_r207_c8 bl[8] br[8] wl[207] vdd gnd cell_6t
Xbit_r208_c8 bl[8] br[8] wl[208] vdd gnd cell_6t
Xbit_r209_c8 bl[8] br[8] wl[209] vdd gnd cell_6t
Xbit_r210_c8 bl[8] br[8] wl[210] vdd gnd cell_6t
Xbit_r211_c8 bl[8] br[8] wl[211] vdd gnd cell_6t
Xbit_r212_c8 bl[8] br[8] wl[212] vdd gnd cell_6t
Xbit_r213_c8 bl[8] br[8] wl[213] vdd gnd cell_6t
Xbit_r214_c8 bl[8] br[8] wl[214] vdd gnd cell_6t
Xbit_r215_c8 bl[8] br[8] wl[215] vdd gnd cell_6t
Xbit_r216_c8 bl[8] br[8] wl[216] vdd gnd cell_6t
Xbit_r217_c8 bl[8] br[8] wl[217] vdd gnd cell_6t
Xbit_r218_c8 bl[8] br[8] wl[218] vdd gnd cell_6t
Xbit_r219_c8 bl[8] br[8] wl[219] vdd gnd cell_6t
Xbit_r220_c8 bl[8] br[8] wl[220] vdd gnd cell_6t
Xbit_r221_c8 bl[8] br[8] wl[221] vdd gnd cell_6t
Xbit_r222_c8 bl[8] br[8] wl[222] vdd gnd cell_6t
Xbit_r223_c8 bl[8] br[8] wl[223] vdd gnd cell_6t
Xbit_r224_c8 bl[8] br[8] wl[224] vdd gnd cell_6t
Xbit_r225_c8 bl[8] br[8] wl[225] vdd gnd cell_6t
Xbit_r226_c8 bl[8] br[8] wl[226] vdd gnd cell_6t
Xbit_r227_c8 bl[8] br[8] wl[227] vdd gnd cell_6t
Xbit_r228_c8 bl[8] br[8] wl[228] vdd gnd cell_6t
Xbit_r229_c8 bl[8] br[8] wl[229] vdd gnd cell_6t
Xbit_r230_c8 bl[8] br[8] wl[230] vdd gnd cell_6t
Xbit_r231_c8 bl[8] br[8] wl[231] vdd gnd cell_6t
Xbit_r232_c8 bl[8] br[8] wl[232] vdd gnd cell_6t
Xbit_r233_c8 bl[8] br[8] wl[233] vdd gnd cell_6t
Xbit_r234_c8 bl[8] br[8] wl[234] vdd gnd cell_6t
Xbit_r235_c8 bl[8] br[8] wl[235] vdd gnd cell_6t
Xbit_r236_c8 bl[8] br[8] wl[236] vdd gnd cell_6t
Xbit_r237_c8 bl[8] br[8] wl[237] vdd gnd cell_6t
Xbit_r238_c8 bl[8] br[8] wl[238] vdd gnd cell_6t
Xbit_r239_c8 bl[8] br[8] wl[239] vdd gnd cell_6t
Xbit_r240_c8 bl[8] br[8] wl[240] vdd gnd cell_6t
Xbit_r241_c8 bl[8] br[8] wl[241] vdd gnd cell_6t
Xbit_r242_c8 bl[8] br[8] wl[242] vdd gnd cell_6t
Xbit_r243_c8 bl[8] br[8] wl[243] vdd gnd cell_6t
Xbit_r244_c8 bl[8] br[8] wl[244] vdd gnd cell_6t
Xbit_r245_c8 bl[8] br[8] wl[245] vdd gnd cell_6t
Xbit_r246_c8 bl[8] br[8] wl[246] vdd gnd cell_6t
Xbit_r247_c8 bl[8] br[8] wl[247] vdd gnd cell_6t
Xbit_r248_c8 bl[8] br[8] wl[248] vdd gnd cell_6t
Xbit_r249_c8 bl[8] br[8] wl[249] vdd gnd cell_6t
Xbit_r250_c8 bl[8] br[8] wl[250] vdd gnd cell_6t
Xbit_r251_c8 bl[8] br[8] wl[251] vdd gnd cell_6t
Xbit_r252_c8 bl[8] br[8] wl[252] vdd gnd cell_6t
Xbit_r253_c8 bl[8] br[8] wl[253] vdd gnd cell_6t
Xbit_r254_c8 bl[8] br[8] wl[254] vdd gnd cell_6t
Xbit_r255_c8 bl[8] br[8] wl[255] vdd gnd cell_6t
Xbit_r256_c8 bl[8] br[8] wl[256] vdd gnd cell_6t
Xbit_r257_c8 bl[8] br[8] wl[257] vdd gnd cell_6t
Xbit_r258_c8 bl[8] br[8] wl[258] vdd gnd cell_6t
Xbit_r259_c8 bl[8] br[8] wl[259] vdd gnd cell_6t
Xbit_r260_c8 bl[8] br[8] wl[260] vdd gnd cell_6t
Xbit_r261_c8 bl[8] br[8] wl[261] vdd gnd cell_6t
Xbit_r262_c8 bl[8] br[8] wl[262] vdd gnd cell_6t
Xbit_r263_c8 bl[8] br[8] wl[263] vdd gnd cell_6t
Xbit_r264_c8 bl[8] br[8] wl[264] vdd gnd cell_6t
Xbit_r265_c8 bl[8] br[8] wl[265] vdd gnd cell_6t
Xbit_r266_c8 bl[8] br[8] wl[266] vdd gnd cell_6t
Xbit_r267_c8 bl[8] br[8] wl[267] vdd gnd cell_6t
Xbit_r268_c8 bl[8] br[8] wl[268] vdd gnd cell_6t
Xbit_r269_c8 bl[8] br[8] wl[269] vdd gnd cell_6t
Xbit_r270_c8 bl[8] br[8] wl[270] vdd gnd cell_6t
Xbit_r271_c8 bl[8] br[8] wl[271] vdd gnd cell_6t
Xbit_r272_c8 bl[8] br[8] wl[272] vdd gnd cell_6t
Xbit_r273_c8 bl[8] br[8] wl[273] vdd gnd cell_6t
Xbit_r274_c8 bl[8] br[8] wl[274] vdd gnd cell_6t
Xbit_r275_c8 bl[8] br[8] wl[275] vdd gnd cell_6t
Xbit_r276_c8 bl[8] br[8] wl[276] vdd gnd cell_6t
Xbit_r277_c8 bl[8] br[8] wl[277] vdd gnd cell_6t
Xbit_r278_c8 bl[8] br[8] wl[278] vdd gnd cell_6t
Xbit_r279_c8 bl[8] br[8] wl[279] vdd gnd cell_6t
Xbit_r280_c8 bl[8] br[8] wl[280] vdd gnd cell_6t
Xbit_r281_c8 bl[8] br[8] wl[281] vdd gnd cell_6t
Xbit_r282_c8 bl[8] br[8] wl[282] vdd gnd cell_6t
Xbit_r283_c8 bl[8] br[8] wl[283] vdd gnd cell_6t
Xbit_r284_c8 bl[8] br[8] wl[284] vdd gnd cell_6t
Xbit_r285_c8 bl[8] br[8] wl[285] vdd gnd cell_6t
Xbit_r286_c8 bl[8] br[8] wl[286] vdd gnd cell_6t
Xbit_r287_c8 bl[8] br[8] wl[287] vdd gnd cell_6t
Xbit_r288_c8 bl[8] br[8] wl[288] vdd gnd cell_6t
Xbit_r289_c8 bl[8] br[8] wl[289] vdd gnd cell_6t
Xbit_r290_c8 bl[8] br[8] wl[290] vdd gnd cell_6t
Xbit_r291_c8 bl[8] br[8] wl[291] vdd gnd cell_6t
Xbit_r292_c8 bl[8] br[8] wl[292] vdd gnd cell_6t
Xbit_r293_c8 bl[8] br[8] wl[293] vdd gnd cell_6t
Xbit_r294_c8 bl[8] br[8] wl[294] vdd gnd cell_6t
Xbit_r295_c8 bl[8] br[8] wl[295] vdd gnd cell_6t
Xbit_r296_c8 bl[8] br[8] wl[296] vdd gnd cell_6t
Xbit_r297_c8 bl[8] br[8] wl[297] vdd gnd cell_6t
Xbit_r298_c8 bl[8] br[8] wl[298] vdd gnd cell_6t
Xbit_r299_c8 bl[8] br[8] wl[299] vdd gnd cell_6t
Xbit_r300_c8 bl[8] br[8] wl[300] vdd gnd cell_6t
Xbit_r301_c8 bl[8] br[8] wl[301] vdd gnd cell_6t
Xbit_r302_c8 bl[8] br[8] wl[302] vdd gnd cell_6t
Xbit_r303_c8 bl[8] br[8] wl[303] vdd gnd cell_6t
Xbit_r304_c8 bl[8] br[8] wl[304] vdd gnd cell_6t
Xbit_r305_c8 bl[8] br[8] wl[305] vdd gnd cell_6t
Xbit_r306_c8 bl[8] br[8] wl[306] vdd gnd cell_6t
Xbit_r307_c8 bl[8] br[8] wl[307] vdd gnd cell_6t
Xbit_r308_c8 bl[8] br[8] wl[308] vdd gnd cell_6t
Xbit_r309_c8 bl[8] br[8] wl[309] vdd gnd cell_6t
Xbit_r310_c8 bl[8] br[8] wl[310] vdd gnd cell_6t
Xbit_r311_c8 bl[8] br[8] wl[311] vdd gnd cell_6t
Xbit_r312_c8 bl[8] br[8] wl[312] vdd gnd cell_6t
Xbit_r313_c8 bl[8] br[8] wl[313] vdd gnd cell_6t
Xbit_r314_c8 bl[8] br[8] wl[314] vdd gnd cell_6t
Xbit_r315_c8 bl[8] br[8] wl[315] vdd gnd cell_6t
Xbit_r316_c8 bl[8] br[8] wl[316] vdd gnd cell_6t
Xbit_r317_c8 bl[8] br[8] wl[317] vdd gnd cell_6t
Xbit_r318_c8 bl[8] br[8] wl[318] vdd gnd cell_6t
Xbit_r319_c8 bl[8] br[8] wl[319] vdd gnd cell_6t
Xbit_r320_c8 bl[8] br[8] wl[320] vdd gnd cell_6t
Xbit_r321_c8 bl[8] br[8] wl[321] vdd gnd cell_6t
Xbit_r322_c8 bl[8] br[8] wl[322] vdd gnd cell_6t
Xbit_r323_c8 bl[8] br[8] wl[323] vdd gnd cell_6t
Xbit_r324_c8 bl[8] br[8] wl[324] vdd gnd cell_6t
Xbit_r325_c8 bl[8] br[8] wl[325] vdd gnd cell_6t
Xbit_r326_c8 bl[8] br[8] wl[326] vdd gnd cell_6t
Xbit_r327_c8 bl[8] br[8] wl[327] vdd gnd cell_6t
Xbit_r328_c8 bl[8] br[8] wl[328] vdd gnd cell_6t
Xbit_r329_c8 bl[8] br[8] wl[329] vdd gnd cell_6t
Xbit_r330_c8 bl[8] br[8] wl[330] vdd gnd cell_6t
Xbit_r331_c8 bl[8] br[8] wl[331] vdd gnd cell_6t
Xbit_r332_c8 bl[8] br[8] wl[332] vdd gnd cell_6t
Xbit_r333_c8 bl[8] br[8] wl[333] vdd gnd cell_6t
Xbit_r334_c8 bl[8] br[8] wl[334] vdd gnd cell_6t
Xbit_r335_c8 bl[8] br[8] wl[335] vdd gnd cell_6t
Xbit_r336_c8 bl[8] br[8] wl[336] vdd gnd cell_6t
Xbit_r337_c8 bl[8] br[8] wl[337] vdd gnd cell_6t
Xbit_r338_c8 bl[8] br[8] wl[338] vdd gnd cell_6t
Xbit_r339_c8 bl[8] br[8] wl[339] vdd gnd cell_6t
Xbit_r340_c8 bl[8] br[8] wl[340] vdd gnd cell_6t
Xbit_r341_c8 bl[8] br[8] wl[341] vdd gnd cell_6t
Xbit_r342_c8 bl[8] br[8] wl[342] vdd gnd cell_6t
Xbit_r343_c8 bl[8] br[8] wl[343] vdd gnd cell_6t
Xbit_r344_c8 bl[8] br[8] wl[344] vdd gnd cell_6t
Xbit_r345_c8 bl[8] br[8] wl[345] vdd gnd cell_6t
Xbit_r346_c8 bl[8] br[8] wl[346] vdd gnd cell_6t
Xbit_r347_c8 bl[8] br[8] wl[347] vdd gnd cell_6t
Xbit_r348_c8 bl[8] br[8] wl[348] vdd gnd cell_6t
Xbit_r349_c8 bl[8] br[8] wl[349] vdd gnd cell_6t
Xbit_r350_c8 bl[8] br[8] wl[350] vdd gnd cell_6t
Xbit_r351_c8 bl[8] br[8] wl[351] vdd gnd cell_6t
Xbit_r352_c8 bl[8] br[8] wl[352] vdd gnd cell_6t
Xbit_r353_c8 bl[8] br[8] wl[353] vdd gnd cell_6t
Xbit_r354_c8 bl[8] br[8] wl[354] vdd gnd cell_6t
Xbit_r355_c8 bl[8] br[8] wl[355] vdd gnd cell_6t
Xbit_r356_c8 bl[8] br[8] wl[356] vdd gnd cell_6t
Xbit_r357_c8 bl[8] br[8] wl[357] vdd gnd cell_6t
Xbit_r358_c8 bl[8] br[8] wl[358] vdd gnd cell_6t
Xbit_r359_c8 bl[8] br[8] wl[359] vdd gnd cell_6t
Xbit_r360_c8 bl[8] br[8] wl[360] vdd gnd cell_6t
Xbit_r361_c8 bl[8] br[8] wl[361] vdd gnd cell_6t
Xbit_r362_c8 bl[8] br[8] wl[362] vdd gnd cell_6t
Xbit_r363_c8 bl[8] br[8] wl[363] vdd gnd cell_6t
Xbit_r364_c8 bl[8] br[8] wl[364] vdd gnd cell_6t
Xbit_r365_c8 bl[8] br[8] wl[365] vdd gnd cell_6t
Xbit_r366_c8 bl[8] br[8] wl[366] vdd gnd cell_6t
Xbit_r367_c8 bl[8] br[8] wl[367] vdd gnd cell_6t
Xbit_r368_c8 bl[8] br[8] wl[368] vdd gnd cell_6t
Xbit_r369_c8 bl[8] br[8] wl[369] vdd gnd cell_6t
Xbit_r370_c8 bl[8] br[8] wl[370] vdd gnd cell_6t
Xbit_r371_c8 bl[8] br[8] wl[371] vdd gnd cell_6t
Xbit_r372_c8 bl[8] br[8] wl[372] vdd gnd cell_6t
Xbit_r373_c8 bl[8] br[8] wl[373] vdd gnd cell_6t
Xbit_r374_c8 bl[8] br[8] wl[374] vdd gnd cell_6t
Xbit_r375_c8 bl[8] br[8] wl[375] vdd gnd cell_6t
Xbit_r376_c8 bl[8] br[8] wl[376] vdd gnd cell_6t
Xbit_r377_c8 bl[8] br[8] wl[377] vdd gnd cell_6t
Xbit_r378_c8 bl[8] br[8] wl[378] vdd gnd cell_6t
Xbit_r379_c8 bl[8] br[8] wl[379] vdd gnd cell_6t
Xbit_r380_c8 bl[8] br[8] wl[380] vdd gnd cell_6t
Xbit_r381_c8 bl[8] br[8] wl[381] vdd gnd cell_6t
Xbit_r382_c8 bl[8] br[8] wl[382] vdd gnd cell_6t
Xbit_r383_c8 bl[8] br[8] wl[383] vdd gnd cell_6t
Xbit_r384_c8 bl[8] br[8] wl[384] vdd gnd cell_6t
Xbit_r385_c8 bl[8] br[8] wl[385] vdd gnd cell_6t
Xbit_r386_c8 bl[8] br[8] wl[386] vdd gnd cell_6t
Xbit_r387_c8 bl[8] br[8] wl[387] vdd gnd cell_6t
Xbit_r388_c8 bl[8] br[8] wl[388] vdd gnd cell_6t
Xbit_r389_c8 bl[8] br[8] wl[389] vdd gnd cell_6t
Xbit_r390_c8 bl[8] br[8] wl[390] vdd gnd cell_6t
Xbit_r391_c8 bl[8] br[8] wl[391] vdd gnd cell_6t
Xbit_r392_c8 bl[8] br[8] wl[392] vdd gnd cell_6t
Xbit_r393_c8 bl[8] br[8] wl[393] vdd gnd cell_6t
Xbit_r394_c8 bl[8] br[8] wl[394] vdd gnd cell_6t
Xbit_r395_c8 bl[8] br[8] wl[395] vdd gnd cell_6t
Xbit_r396_c8 bl[8] br[8] wl[396] vdd gnd cell_6t
Xbit_r397_c8 bl[8] br[8] wl[397] vdd gnd cell_6t
Xbit_r398_c8 bl[8] br[8] wl[398] vdd gnd cell_6t
Xbit_r399_c8 bl[8] br[8] wl[399] vdd gnd cell_6t
Xbit_r400_c8 bl[8] br[8] wl[400] vdd gnd cell_6t
Xbit_r401_c8 bl[8] br[8] wl[401] vdd gnd cell_6t
Xbit_r402_c8 bl[8] br[8] wl[402] vdd gnd cell_6t
Xbit_r403_c8 bl[8] br[8] wl[403] vdd gnd cell_6t
Xbit_r404_c8 bl[8] br[8] wl[404] vdd gnd cell_6t
Xbit_r405_c8 bl[8] br[8] wl[405] vdd gnd cell_6t
Xbit_r406_c8 bl[8] br[8] wl[406] vdd gnd cell_6t
Xbit_r407_c8 bl[8] br[8] wl[407] vdd gnd cell_6t
Xbit_r408_c8 bl[8] br[8] wl[408] vdd gnd cell_6t
Xbit_r409_c8 bl[8] br[8] wl[409] vdd gnd cell_6t
Xbit_r410_c8 bl[8] br[8] wl[410] vdd gnd cell_6t
Xbit_r411_c8 bl[8] br[8] wl[411] vdd gnd cell_6t
Xbit_r412_c8 bl[8] br[8] wl[412] vdd gnd cell_6t
Xbit_r413_c8 bl[8] br[8] wl[413] vdd gnd cell_6t
Xbit_r414_c8 bl[8] br[8] wl[414] vdd gnd cell_6t
Xbit_r415_c8 bl[8] br[8] wl[415] vdd gnd cell_6t
Xbit_r416_c8 bl[8] br[8] wl[416] vdd gnd cell_6t
Xbit_r417_c8 bl[8] br[8] wl[417] vdd gnd cell_6t
Xbit_r418_c8 bl[8] br[8] wl[418] vdd gnd cell_6t
Xbit_r419_c8 bl[8] br[8] wl[419] vdd gnd cell_6t
Xbit_r420_c8 bl[8] br[8] wl[420] vdd gnd cell_6t
Xbit_r421_c8 bl[8] br[8] wl[421] vdd gnd cell_6t
Xbit_r422_c8 bl[8] br[8] wl[422] vdd gnd cell_6t
Xbit_r423_c8 bl[8] br[8] wl[423] vdd gnd cell_6t
Xbit_r424_c8 bl[8] br[8] wl[424] vdd gnd cell_6t
Xbit_r425_c8 bl[8] br[8] wl[425] vdd gnd cell_6t
Xbit_r426_c8 bl[8] br[8] wl[426] vdd gnd cell_6t
Xbit_r427_c8 bl[8] br[8] wl[427] vdd gnd cell_6t
Xbit_r428_c8 bl[8] br[8] wl[428] vdd gnd cell_6t
Xbit_r429_c8 bl[8] br[8] wl[429] vdd gnd cell_6t
Xbit_r430_c8 bl[8] br[8] wl[430] vdd gnd cell_6t
Xbit_r431_c8 bl[8] br[8] wl[431] vdd gnd cell_6t
Xbit_r432_c8 bl[8] br[8] wl[432] vdd gnd cell_6t
Xbit_r433_c8 bl[8] br[8] wl[433] vdd gnd cell_6t
Xbit_r434_c8 bl[8] br[8] wl[434] vdd gnd cell_6t
Xbit_r435_c8 bl[8] br[8] wl[435] vdd gnd cell_6t
Xbit_r436_c8 bl[8] br[8] wl[436] vdd gnd cell_6t
Xbit_r437_c8 bl[8] br[8] wl[437] vdd gnd cell_6t
Xbit_r438_c8 bl[8] br[8] wl[438] vdd gnd cell_6t
Xbit_r439_c8 bl[8] br[8] wl[439] vdd gnd cell_6t
Xbit_r440_c8 bl[8] br[8] wl[440] vdd gnd cell_6t
Xbit_r441_c8 bl[8] br[8] wl[441] vdd gnd cell_6t
Xbit_r442_c8 bl[8] br[8] wl[442] vdd gnd cell_6t
Xbit_r443_c8 bl[8] br[8] wl[443] vdd gnd cell_6t
Xbit_r444_c8 bl[8] br[8] wl[444] vdd gnd cell_6t
Xbit_r445_c8 bl[8] br[8] wl[445] vdd gnd cell_6t
Xbit_r446_c8 bl[8] br[8] wl[446] vdd gnd cell_6t
Xbit_r447_c8 bl[8] br[8] wl[447] vdd gnd cell_6t
Xbit_r448_c8 bl[8] br[8] wl[448] vdd gnd cell_6t
Xbit_r449_c8 bl[8] br[8] wl[449] vdd gnd cell_6t
Xbit_r450_c8 bl[8] br[8] wl[450] vdd gnd cell_6t
Xbit_r451_c8 bl[8] br[8] wl[451] vdd gnd cell_6t
Xbit_r452_c8 bl[8] br[8] wl[452] vdd gnd cell_6t
Xbit_r453_c8 bl[8] br[8] wl[453] vdd gnd cell_6t
Xbit_r454_c8 bl[8] br[8] wl[454] vdd gnd cell_6t
Xbit_r455_c8 bl[8] br[8] wl[455] vdd gnd cell_6t
Xbit_r456_c8 bl[8] br[8] wl[456] vdd gnd cell_6t
Xbit_r457_c8 bl[8] br[8] wl[457] vdd gnd cell_6t
Xbit_r458_c8 bl[8] br[8] wl[458] vdd gnd cell_6t
Xbit_r459_c8 bl[8] br[8] wl[459] vdd gnd cell_6t
Xbit_r460_c8 bl[8] br[8] wl[460] vdd gnd cell_6t
Xbit_r461_c8 bl[8] br[8] wl[461] vdd gnd cell_6t
Xbit_r462_c8 bl[8] br[8] wl[462] vdd gnd cell_6t
Xbit_r463_c8 bl[8] br[8] wl[463] vdd gnd cell_6t
Xbit_r464_c8 bl[8] br[8] wl[464] vdd gnd cell_6t
Xbit_r465_c8 bl[8] br[8] wl[465] vdd gnd cell_6t
Xbit_r466_c8 bl[8] br[8] wl[466] vdd gnd cell_6t
Xbit_r467_c8 bl[8] br[8] wl[467] vdd gnd cell_6t
Xbit_r468_c8 bl[8] br[8] wl[468] vdd gnd cell_6t
Xbit_r469_c8 bl[8] br[8] wl[469] vdd gnd cell_6t
Xbit_r470_c8 bl[8] br[8] wl[470] vdd gnd cell_6t
Xbit_r471_c8 bl[8] br[8] wl[471] vdd gnd cell_6t
Xbit_r472_c8 bl[8] br[8] wl[472] vdd gnd cell_6t
Xbit_r473_c8 bl[8] br[8] wl[473] vdd gnd cell_6t
Xbit_r474_c8 bl[8] br[8] wl[474] vdd gnd cell_6t
Xbit_r475_c8 bl[8] br[8] wl[475] vdd gnd cell_6t
Xbit_r476_c8 bl[8] br[8] wl[476] vdd gnd cell_6t
Xbit_r477_c8 bl[8] br[8] wl[477] vdd gnd cell_6t
Xbit_r478_c8 bl[8] br[8] wl[478] vdd gnd cell_6t
Xbit_r479_c8 bl[8] br[8] wl[479] vdd gnd cell_6t
Xbit_r480_c8 bl[8] br[8] wl[480] vdd gnd cell_6t
Xbit_r481_c8 bl[8] br[8] wl[481] vdd gnd cell_6t
Xbit_r482_c8 bl[8] br[8] wl[482] vdd gnd cell_6t
Xbit_r483_c8 bl[8] br[8] wl[483] vdd gnd cell_6t
Xbit_r484_c8 bl[8] br[8] wl[484] vdd gnd cell_6t
Xbit_r485_c8 bl[8] br[8] wl[485] vdd gnd cell_6t
Xbit_r486_c8 bl[8] br[8] wl[486] vdd gnd cell_6t
Xbit_r487_c8 bl[8] br[8] wl[487] vdd gnd cell_6t
Xbit_r488_c8 bl[8] br[8] wl[488] vdd gnd cell_6t
Xbit_r489_c8 bl[8] br[8] wl[489] vdd gnd cell_6t
Xbit_r490_c8 bl[8] br[8] wl[490] vdd gnd cell_6t
Xbit_r491_c8 bl[8] br[8] wl[491] vdd gnd cell_6t
Xbit_r492_c8 bl[8] br[8] wl[492] vdd gnd cell_6t
Xbit_r493_c8 bl[8] br[8] wl[493] vdd gnd cell_6t
Xbit_r494_c8 bl[8] br[8] wl[494] vdd gnd cell_6t
Xbit_r495_c8 bl[8] br[8] wl[495] vdd gnd cell_6t
Xbit_r496_c8 bl[8] br[8] wl[496] vdd gnd cell_6t
Xbit_r497_c8 bl[8] br[8] wl[497] vdd gnd cell_6t
Xbit_r498_c8 bl[8] br[8] wl[498] vdd gnd cell_6t
Xbit_r499_c8 bl[8] br[8] wl[499] vdd gnd cell_6t
Xbit_r500_c8 bl[8] br[8] wl[500] vdd gnd cell_6t
Xbit_r501_c8 bl[8] br[8] wl[501] vdd gnd cell_6t
Xbit_r502_c8 bl[8] br[8] wl[502] vdd gnd cell_6t
Xbit_r503_c8 bl[8] br[8] wl[503] vdd gnd cell_6t
Xbit_r504_c8 bl[8] br[8] wl[504] vdd gnd cell_6t
Xbit_r505_c8 bl[8] br[8] wl[505] vdd gnd cell_6t
Xbit_r506_c8 bl[8] br[8] wl[506] vdd gnd cell_6t
Xbit_r507_c8 bl[8] br[8] wl[507] vdd gnd cell_6t
Xbit_r508_c8 bl[8] br[8] wl[508] vdd gnd cell_6t
Xbit_r509_c8 bl[8] br[8] wl[509] vdd gnd cell_6t
Xbit_r510_c8 bl[8] br[8] wl[510] vdd gnd cell_6t
Xbit_r511_c8 bl[8] br[8] wl[511] vdd gnd cell_6t
Xbit_r0_c9 bl[9] br[9] wl[0] vdd gnd cell_6t
Xbit_r1_c9 bl[9] br[9] wl[1] vdd gnd cell_6t
Xbit_r2_c9 bl[9] br[9] wl[2] vdd gnd cell_6t
Xbit_r3_c9 bl[9] br[9] wl[3] vdd gnd cell_6t
Xbit_r4_c9 bl[9] br[9] wl[4] vdd gnd cell_6t
Xbit_r5_c9 bl[9] br[9] wl[5] vdd gnd cell_6t
Xbit_r6_c9 bl[9] br[9] wl[6] vdd gnd cell_6t
Xbit_r7_c9 bl[9] br[9] wl[7] vdd gnd cell_6t
Xbit_r8_c9 bl[9] br[9] wl[8] vdd gnd cell_6t
Xbit_r9_c9 bl[9] br[9] wl[9] vdd gnd cell_6t
Xbit_r10_c9 bl[9] br[9] wl[10] vdd gnd cell_6t
Xbit_r11_c9 bl[9] br[9] wl[11] vdd gnd cell_6t
Xbit_r12_c9 bl[9] br[9] wl[12] vdd gnd cell_6t
Xbit_r13_c9 bl[9] br[9] wl[13] vdd gnd cell_6t
Xbit_r14_c9 bl[9] br[9] wl[14] vdd gnd cell_6t
Xbit_r15_c9 bl[9] br[9] wl[15] vdd gnd cell_6t
Xbit_r16_c9 bl[9] br[9] wl[16] vdd gnd cell_6t
Xbit_r17_c9 bl[9] br[9] wl[17] vdd gnd cell_6t
Xbit_r18_c9 bl[9] br[9] wl[18] vdd gnd cell_6t
Xbit_r19_c9 bl[9] br[9] wl[19] vdd gnd cell_6t
Xbit_r20_c9 bl[9] br[9] wl[20] vdd gnd cell_6t
Xbit_r21_c9 bl[9] br[9] wl[21] vdd gnd cell_6t
Xbit_r22_c9 bl[9] br[9] wl[22] vdd gnd cell_6t
Xbit_r23_c9 bl[9] br[9] wl[23] vdd gnd cell_6t
Xbit_r24_c9 bl[9] br[9] wl[24] vdd gnd cell_6t
Xbit_r25_c9 bl[9] br[9] wl[25] vdd gnd cell_6t
Xbit_r26_c9 bl[9] br[9] wl[26] vdd gnd cell_6t
Xbit_r27_c9 bl[9] br[9] wl[27] vdd gnd cell_6t
Xbit_r28_c9 bl[9] br[9] wl[28] vdd gnd cell_6t
Xbit_r29_c9 bl[9] br[9] wl[29] vdd gnd cell_6t
Xbit_r30_c9 bl[9] br[9] wl[30] vdd gnd cell_6t
Xbit_r31_c9 bl[9] br[9] wl[31] vdd gnd cell_6t
Xbit_r32_c9 bl[9] br[9] wl[32] vdd gnd cell_6t
Xbit_r33_c9 bl[9] br[9] wl[33] vdd gnd cell_6t
Xbit_r34_c9 bl[9] br[9] wl[34] vdd gnd cell_6t
Xbit_r35_c9 bl[9] br[9] wl[35] vdd gnd cell_6t
Xbit_r36_c9 bl[9] br[9] wl[36] vdd gnd cell_6t
Xbit_r37_c9 bl[9] br[9] wl[37] vdd gnd cell_6t
Xbit_r38_c9 bl[9] br[9] wl[38] vdd gnd cell_6t
Xbit_r39_c9 bl[9] br[9] wl[39] vdd gnd cell_6t
Xbit_r40_c9 bl[9] br[9] wl[40] vdd gnd cell_6t
Xbit_r41_c9 bl[9] br[9] wl[41] vdd gnd cell_6t
Xbit_r42_c9 bl[9] br[9] wl[42] vdd gnd cell_6t
Xbit_r43_c9 bl[9] br[9] wl[43] vdd gnd cell_6t
Xbit_r44_c9 bl[9] br[9] wl[44] vdd gnd cell_6t
Xbit_r45_c9 bl[9] br[9] wl[45] vdd gnd cell_6t
Xbit_r46_c9 bl[9] br[9] wl[46] vdd gnd cell_6t
Xbit_r47_c9 bl[9] br[9] wl[47] vdd gnd cell_6t
Xbit_r48_c9 bl[9] br[9] wl[48] vdd gnd cell_6t
Xbit_r49_c9 bl[9] br[9] wl[49] vdd gnd cell_6t
Xbit_r50_c9 bl[9] br[9] wl[50] vdd gnd cell_6t
Xbit_r51_c9 bl[9] br[9] wl[51] vdd gnd cell_6t
Xbit_r52_c9 bl[9] br[9] wl[52] vdd gnd cell_6t
Xbit_r53_c9 bl[9] br[9] wl[53] vdd gnd cell_6t
Xbit_r54_c9 bl[9] br[9] wl[54] vdd gnd cell_6t
Xbit_r55_c9 bl[9] br[9] wl[55] vdd gnd cell_6t
Xbit_r56_c9 bl[9] br[9] wl[56] vdd gnd cell_6t
Xbit_r57_c9 bl[9] br[9] wl[57] vdd gnd cell_6t
Xbit_r58_c9 bl[9] br[9] wl[58] vdd gnd cell_6t
Xbit_r59_c9 bl[9] br[9] wl[59] vdd gnd cell_6t
Xbit_r60_c9 bl[9] br[9] wl[60] vdd gnd cell_6t
Xbit_r61_c9 bl[9] br[9] wl[61] vdd gnd cell_6t
Xbit_r62_c9 bl[9] br[9] wl[62] vdd gnd cell_6t
Xbit_r63_c9 bl[9] br[9] wl[63] vdd gnd cell_6t
Xbit_r64_c9 bl[9] br[9] wl[64] vdd gnd cell_6t
Xbit_r65_c9 bl[9] br[9] wl[65] vdd gnd cell_6t
Xbit_r66_c9 bl[9] br[9] wl[66] vdd gnd cell_6t
Xbit_r67_c9 bl[9] br[9] wl[67] vdd gnd cell_6t
Xbit_r68_c9 bl[9] br[9] wl[68] vdd gnd cell_6t
Xbit_r69_c9 bl[9] br[9] wl[69] vdd gnd cell_6t
Xbit_r70_c9 bl[9] br[9] wl[70] vdd gnd cell_6t
Xbit_r71_c9 bl[9] br[9] wl[71] vdd gnd cell_6t
Xbit_r72_c9 bl[9] br[9] wl[72] vdd gnd cell_6t
Xbit_r73_c9 bl[9] br[9] wl[73] vdd gnd cell_6t
Xbit_r74_c9 bl[9] br[9] wl[74] vdd gnd cell_6t
Xbit_r75_c9 bl[9] br[9] wl[75] vdd gnd cell_6t
Xbit_r76_c9 bl[9] br[9] wl[76] vdd gnd cell_6t
Xbit_r77_c9 bl[9] br[9] wl[77] vdd gnd cell_6t
Xbit_r78_c9 bl[9] br[9] wl[78] vdd gnd cell_6t
Xbit_r79_c9 bl[9] br[9] wl[79] vdd gnd cell_6t
Xbit_r80_c9 bl[9] br[9] wl[80] vdd gnd cell_6t
Xbit_r81_c9 bl[9] br[9] wl[81] vdd gnd cell_6t
Xbit_r82_c9 bl[9] br[9] wl[82] vdd gnd cell_6t
Xbit_r83_c9 bl[9] br[9] wl[83] vdd gnd cell_6t
Xbit_r84_c9 bl[9] br[9] wl[84] vdd gnd cell_6t
Xbit_r85_c9 bl[9] br[9] wl[85] vdd gnd cell_6t
Xbit_r86_c9 bl[9] br[9] wl[86] vdd gnd cell_6t
Xbit_r87_c9 bl[9] br[9] wl[87] vdd gnd cell_6t
Xbit_r88_c9 bl[9] br[9] wl[88] vdd gnd cell_6t
Xbit_r89_c9 bl[9] br[9] wl[89] vdd gnd cell_6t
Xbit_r90_c9 bl[9] br[9] wl[90] vdd gnd cell_6t
Xbit_r91_c9 bl[9] br[9] wl[91] vdd gnd cell_6t
Xbit_r92_c9 bl[9] br[9] wl[92] vdd gnd cell_6t
Xbit_r93_c9 bl[9] br[9] wl[93] vdd gnd cell_6t
Xbit_r94_c9 bl[9] br[9] wl[94] vdd gnd cell_6t
Xbit_r95_c9 bl[9] br[9] wl[95] vdd gnd cell_6t
Xbit_r96_c9 bl[9] br[9] wl[96] vdd gnd cell_6t
Xbit_r97_c9 bl[9] br[9] wl[97] vdd gnd cell_6t
Xbit_r98_c9 bl[9] br[9] wl[98] vdd gnd cell_6t
Xbit_r99_c9 bl[9] br[9] wl[99] vdd gnd cell_6t
Xbit_r100_c9 bl[9] br[9] wl[100] vdd gnd cell_6t
Xbit_r101_c9 bl[9] br[9] wl[101] vdd gnd cell_6t
Xbit_r102_c9 bl[9] br[9] wl[102] vdd gnd cell_6t
Xbit_r103_c9 bl[9] br[9] wl[103] vdd gnd cell_6t
Xbit_r104_c9 bl[9] br[9] wl[104] vdd gnd cell_6t
Xbit_r105_c9 bl[9] br[9] wl[105] vdd gnd cell_6t
Xbit_r106_c9 bl[9] br[9] wl[106] vdd gnd cell_6t
Xbit_r107_c9 bl[9] br[9] wl[107] vdd gnd cell_6t
Xbit_r108_c9 bl[9] br[9] wl[108] vdd gnd cell_6t
Xbit_r109_c9 bl[9] br[9] wl[109] vdd gnd cell_6t
Xbit_r110_c9 bl[9] br[9] wl[110] vdd gnd cell_6t
Xbit_r111_c9 bl[9] br[9] wl[111] vdd gnd cell_6t
Xbit_r112_c9 bl[9] br[9] wl[112] vdd gnd cell_6t
Xbit_r113_c9 bl[9] br[9] wl[113] vdd gnd cell_6t
Xbit_r114_c9 bl[9] br[9] wl[114] vdd gnd cell_6t
Xbit_r115_c9 bl[9] br[9] wl[115] vdd gnd cell_6t
Xbit_r116_c9 bl[9] br[9] wl[116] vdd gnd cell_6t
Xbit_r117_c9 bl[9] br[9] wl[117] vdd gnd cell_6t
Xbit_r118_c9 bl[9] br[9] wl[118] vdd gnd cell_6t
Xbit_r119_c9 bl[9] br[9] wl[119] vdd gnd cell_6t
Xbit_r120_c9 bl[9] br[9] wl[120] vdd gnd cell_6t
Xbit_r121_c9 bl[9] br[9] wl[121] vdd gnd cell_6t
Xbit_r122_c9 bl[9] br[9] wl[122] vdd gnd cell_6t
Xbit_r123_c9 bl[9] br[9] wl[123] vdd gnd cell_6t
Xbit_r124_c9 bl[9] br[9] wl[124] vdd gnd cell_6t
Xbit_r125_c9 bl[9] br[9] wl[125] vdd gnd cell_6t
Xbit_r126_c9 bl[9] br[9] wl[126] vdd gnd cell_6t
Xbit_r127_c9 bl[9] br[9] wl[127] vdd gnd cell_6t
Xbit_r128_c9 bl[9] br[9] wl[128] vdd gnd cell_6t
Xbit_r129_c9 bl[9] br[9] wl[129] vdd gnd cell_6t
Xbit_r130_c9 bl[9] br[9] wl[130] vdd gnd cell_6t
Xbit_r131_c9 bl[9] br[9] wl[131] vdd gnd cell_6t
Xbit_r132_c9 bl[9] br[9] wl[132] vdd gnd cell_6t
Xbit_r133_c9 bl[9] br[9] wl[133] vdd gnd cell_6t
Xbit_r134_c9 bl[9] br[9] wl[134] vdd gnd cell_6t
Xbit_r135_c9 bl[9] br[9] wl[135] vdd gnd cell_6t
Xbit_r136_c9 bl[9] br[9] wl[136] vdd gnd cell_6t
Xbit_r137_c9 bl[9] br[9] wl[137] vdd gnd cell_6t
Xbit_r138_c9 bl[9] br[9] wl[138] vdd gnd cell_6t
Xbit_r139_c9 bl[9] br[9] wl[139] vdd gnd cell_6t
Xbit_r140_c9 bl[9] br[9] wl[140] vdd gnd cell_6t
Xbit_r141_c9 bl[9] br[9] wl[141] vdd gnd cell_6t
Xbit_r142_c9 bl[9] br[9] wl[142] vdd gnd cell_6t
Xbit_r143_c9 bl[9] br[9] wl[143] vdd gnd cell_6t
Xbit_r144_c9 bl[9] br[9] wl[144] vdd gnd cell_6t
Xbit_r145_c9 bl[9] br[9] wl[145] vdd gnd cell_6t
Xbit_r146_c9 bl[9] br[9] wl[146] vdd gnd cell_6t
Xbit_r147_c9 bl[9] br[9] wl[147] vdd gnd cell_6t
Xbit_r148_c9 bl[9] br[9] wl[148] vdd gnd cell_6t
Xbit_r149_c9 bl[9] br[9] wl[149] vdd gnd cell_6t
Xbit_r150_c9 bl[9] br[9] wl[150] vdd gnd cell_6t
Xbit_r151_c9 bl[9] br[9] wl[151] vdd gnd cell_6t
Xbit_r152_c9 bl[9] br[9] wl[152] vdd gnd cell_6t
Xbit_r153_c9 bl[9] br[9] wl[153] vdd gnd cell_6t
Xbit_r154_c9 bl[9] br[9] wl[154] vdd gnd cell_6t
Xbit_r155_c9 bl[9] br[9] wl[155] vdd gnd cell_6t
Xbit_r156_c9 bl[9] br[9] wl[156] vdd gnd cell_6t
Xbit_r157_c9 bl[9] br[9] wl[157] vdd gnd cell_6t
Xbit_r158_c9 bl[9] br[9] wl[158] vdd gnd cell_6t
Xbit_r159_c9 bl[9] br[9] wl[159] vdd gnd cell_6t
Xbit_r160_c9 bl[9] br[9] wl[160] vdd gnd cell_6t
Xbit_r161_c9 bl[9] br[9] wl[161] vdd gnd cell_6t
Xbit_r162_c9 bl[9] br[9] wl[162] vdd gnd cell_6t
Xbit_r163_c9 bl[9] br[9] wl[163] vdd gnd cell_6t
Xbit_r164_c9 bl[9] br[9] wl[164] vdd gnd cell_6t
Xbit_r165_c9 bl[9] br[9] wl[165] vdd gnd cell_6t
Xbit_r166_c9 bl[9] br[9] wl[166] vdd gnd cell_6t
Xbit_r167_c9 bl[9] br[9] wl[167] vdd gnd cell_6t
Xbit_r168_c9 bl[9] br[9] wl[168] vdd gnd cell_6t
Xbit_r169_c9 bl[9] br[9] wl[169] vdd gnd cell_6t
Xbit_r170_c9 bl[9] br[9] wl[170] vdd gnd cell_6t
Xbit_r171_c9 bl[9] br[9] wl[171] vdd gnd cell_6t
Xbit_r172_c9 bl[9] br[9] wl[172] vdd gnd cell_6t
Xbit_r173_c9 bl[9] br[9] wl[173] vdd gnd cell_6t
Xbit_r174_c9 bl[9] br[9] wl[174] vdd gnd cell_6t
Xbit_r175_c9 bl[9] br[9] wl[175] vdd gnd cell_6t
Xbit_r176_c9 bl[9] br[9] wl[176] vdd gnd cell_6t
Xbit_r177_c9 bl[9] br[9] wl[177] vdd gnd cell_6t
Xbit_r178_c9 bl[9] br[9] wl[178] vdd gnd cell_6t
Xbit_r179_c9 bl[9] br[9] wl[179] vdd gnd cell_6t
Xbit_r180_c9 bl[9] br[9] wl[180] vdd gnd cell_6t
Xbit_r181_c9 bl[9] br[9] wl[181] vdd gnd cell_6t
Xbit_r182_c9 bl[9] br[9] wl[182] vdd gnd cell_6t
Xbit_r183_c9 bl[9] br[9] wl[183] vdd gnd cell_6t
Xbit_r184_c9 bl[9] br[9] wl[184] vdd gnd cell_6t
Xbit_r185_c9 bl[9] br[9] wl[185] vdd gnd cell_6t
Xbit_r186_c9 bl[9] br[9] wl[186] vdd gnd cell_6t
Xbit_r187_c9 bl[9] br[9] wl[187] vdd gnd cell_6t
Xbit_r188_c9 bl[9] br[9] wl[188] vdd gnd cell_6t
Xbit_r189_c9 bl[9] br[9] wl[189] vdd gnd cell_6t
Xbit_r190_c9 bl[9] br[9] wl[190] vdd gnd cell_6t
Xbit_r191_c9 bl[9] br[9] wl[191] vdd gnd cell_6t
Xbit_r192_c9 bl[9] br[9] wl[192] vdd gnd cell_6t
Xbit_r193_c9 bl[9] br[9] wl[193] vdd gnd cell_6t
Xbit_r194_c9 bl[9] br[9] wl[194] vdd gnd cell_6t
Xbit_r195_c9 bl[9] br[9] wl[195] vdd gnd cell_6t
Xbit_r196_c9 bl[9] br[9] wl[196] vdd gnd cell_6t
Xbit_r197_c9 bl[9] br[9] wl[197] vdd gnd cell_6t
Xbit_r198_c9 bl[9] br[9] wl[198] vdd gnd cell_6t
Xbit_r199_c9 bl[9] br[9] wl[199] vdd gnd cell_6t
Xbit_r200_c9 bl[9] br[9] wl[200] vdd gnd cell_6t
Xbit_r201_c9 bl[9] br[9] wl[201] vdd gnd cell_6t
Xbit_r202_c9 bl[9] br[9] wl[202] vdd gnd cell_6t
Xbit_r203_c9 bl[9] br[9] wl[203] vdd gnd cell_6t
Xbit_r204_c9 bl[9] br[9] wl[204] vdd gnd cell_6t
Xbit_r205_c9 bl[9] br[9] wl[205] vdd gnd cell_6t
Xbit_r206_c9 bl[9] br[9] wl[206] vdd gnd cell_6t
Xbit_r207_c9 bl[9] br[9] wl[207] vdd gnd cell_6t
Xbit_r208_c9 bl[9] br[9] wl[208] vdd gnd cell_6t
Xbit_r209_c9 bl[9] br[9] wl[209] vdd gnd cell_6t
Xbit_r210_c9 bl[9] br[9] wl[210] vdd gnd cell_6t
Xbit_r211_c9 bl[9] br[9] wl[211] vdd gnd cell_6t
Xbit_r212_c9 bl[9] br[9] wl[212] vdd gnd cell_6t
Xbit_r213_c9 bl[9] br[9] wl[213] vdd gnd cell_6t
Xbit_r214_c9 bl[9] br[9] wl[214] vdd gnd cell_6t
Xbit_r215_c9 bl[9] br[9] wl[215] vdd gnd cell_6t
Xbit_r216_c9 bl[9] br[9] wl[216] vdd gnd cell_6t
Xbit_r217_c9 bl[9] br[9] wl[217] vdd gnd cell_6t
Xbit_r218_c9 bl[9] br[9] wl[218] vdd gnd cell_6t
Xbit_r219_c9 bl[9] br[9] wl[219] vdd gnd cell_6t
Xbit_r220_c9 bl[9] br[9] wl[220] vdd gnd cell_6t
Xbit_r221_c9 bl[9] br[9] wl[221] vdd gnd cell_6t
Xbit_r222_c9 bl[9] br[9] wl[222] vdd gnd cell_6t
Xbit_r223_c9 bl[9] br[9] wl[223] vdd gnd cell_6t
Xbit_r224_c9 bl[9] br[9] wl[224] vdd gnd cell_6t
Xbit_r225_c9 bl[9] br[9] wl[225] vdd gnd cell_6t
Xbit_r226_c9 bl[9] br[9] wl[226] vdd gnd cell_6t
Xbit_r227_c9 bl[9] br[9] wl[227] vdd gnd cell_6t
Xbit_r228_c9 bl[9] br[9] wl[228] vdd gnd cell_6t
Xbit_r229_c9 bl[9] br[9] wl[229] vdd gnd cell_6t
Xbit_r230_c9 bl[9] br[9] wl[230] vdd gnd cell_6t
Xbit_r231_c9 bl[9] br[9] wl[231] vdd gnd cell_6t
Xbit_r232_c9 bl[9] br[9] wl[232] vdd gnd cell_6t
Xbit_r233_c9 bl[9] br[9] wl[233] vdd gnd cell_6t
Xbit_r234_c9 bl[9] br[9] wl[234] vdd gnd cell_6t
Xbit_r235_c9 bl[9] br[9] wl[235] vdd gnd cell_6t
Xbit_r236_c9 bl[9] br[9] wl[236] vdd gnd cell_6t
Xbit_r237_c9 bl[9] br[9] wl[237] vdd gnd cell_6t
Xbit_r238_c9 bl[9] br[9] wl[238] vdd gnd cell_6t
Xbit_r239_c9 bl[9] br[9] wl[239] vdd gnd cell_6t
Xbit_r240_c9 bl[9] br[9] wl[240] vdd gnd cell_6t
Xbit_r241_c9 bl[9] br[9] wl[241] vdd gnd cell_6t
Xbit_r242_c9 bl[9] br[9] wl[242] vdd gnd cell_6t
Xbit_r243_c9 bl[9] br[9] wl[243] vdd gnd cell_6t
Xbit_r244_c9 bl[9] br[9] wl[244] vdd gnd cell_6t
Xbit_r245_c9 bl[9] br[9] wl[245] vdd gnd cell_6t
Xbit_r246_c9 bl[9] br[9] wl[246] vdd gnd cell_6t
Xbit_r247_c9 bl[9] br[9] wl[247] vdd gnd cell_6t
Xbit_r248_c9 bl[9] br[9] wl[248] vdd gnd cell_6t
Xbit_r249_c9 bl[9] br[9] wl[249] vdd gnd cell_6t
Xbit_r250_c9 bl[9] br[9] wl[250] vdd gnd cell_6t
Xbit_r251_c9 bl[9] br[9] wl[251] vdd gnd cell_6t
Xbit_r252_c9 bl[9] br[9] wl[252] vdd gnd cell_6t
Xbit_r253_c9 bl[9] br[9] wl[253] vdd gnd cell_6t
Xbit_r254_c9 bl[9] br[9] wl[254] vdd gnd cell_6t
Xbit_r255_c9 bl[9] br[9] wl[255] vdd gnd cell_6t
Xbit_r256_c9 bl[9] br[9] wl[256] vdd gnd cell_6t
Xbit_r257_c9 bl[9] br[9] wl[257] vdd gnd cell_6t
Xbit_r258_c9 bl[9] br[9] wl[258] vdd gnd cell_6t
Xbit_r259_c9 bl[9] br[9] wl[259] vdd gnd cell_6t
Xbit_r260_c9 bl[9] br[9] wl[260] vdd gnd cell_6t
Xbit_r261_c9 bl[9] br[9] wl[261] vdd gnd cell_6t
Xbit_r262_c9 bl[9] br[9] wl[262] vdd gnd cell_6t
Xbit_r263_c9 bl[9] br[9] wl[263] vdd gnd cell_6t
Xbit_r264_c9 bl[9] br[9] wl[264] vdd gnd cell_6t
Xbit_r265_c9 bl[9] br[9] wl[265] vdd gnd cell_6t
Xbit_r266_c9 bl[9] br[9] wl[266] vdd gnd cell_6t
Xbit_r267_c9 bl[9] br[9] wl[267] vdd gnd cell_6t
Xbit_r268_c9 bl[9] br[9] wl[268] vdd gnd cell_6t
Xbit_r269_c9 bl[9] br[9] wl[269] vdd gnd cell_6t
Xbit_r270_c9 bl[9] br[9] wl[270] vdd gnd cell_6t
Xbit_r271_c9 bl[9] br[9] wl[271] vdd gnd cell_6t
Xbit_r272_c9 bl[9] br[9] wl[272] vdd gnd cell_6t
Xbit_r273_c9 bl[9] br[9] wl[273] vdd gnd cell_6t
Xbit_r274_c9 bl[9] br[9] wl[274] vdd gnd cell_6t
Xbit_r275_c9 bl[9] br[9] wl[275] vdd gnd cell_6t
Xbit_r276_c9 bl[9] br[9] wl[276] vdd gnd cell_6t
Xbit_r277_c9 bl[9] br[9] wl[277] vdd gnd cell_6t
Xbit_r278_c9 bl[9] br[9] wl[278] vdd gnd cell_6t
Xbit_r279_c9 bl[9] br[9] wl[279] vdd gnd cell_6t
Xbit_r280_c9 bl[9] br[9] wl[280] vdd gnd cell_6t
Xbit_r281_c9 bl[9] br[9] wl[281] vdd gnd cell_6t
Xbit_r282_c9 bl[9] br[9] wl[282] vdd gnd cell_6t
Xbit_r283_c9 bl[9] br[9] wl[283] vdd gnd cell_6t
Xbit_r284_c9 bl[9] br[9] wl[284] vdd gnd cell_6t
Xbit_r285_c9 bl[9] br[9] wl[285] vdd gnd cell_6t
Xbit_r286_c9 bl[9] br[9] wl[286] vdd gnd cell_6t
Xbit_r287_c9 bl[9] br[9] wl[287] vdd gnd cell_6t
Xbit_r288_c9 bl[9] br[9] wl[288] vdd gnd cell_6t
Xbit_r289_c9 bl[9] br[9] wl[289] vdd gnd cell_6t
Xbit_r290_c9 bl[9] br[9] wl[290] vdd gnd cell_6t
Xbit_r291_c9 bl[9] br[9] wl[291] vdd gnd cell_6t
Xbit_r292_c9 bl[9] br[9] wl[292] vdd gnd cell_6t
Xbit_r293_c9 bl[9] br[9] wl[293] vdd gnd cell_6t
Xbit_r294_c9 bl[9] br[9] wl[294] vdd gnd cell_6t
Xbit_r295_c9 bl[9] br[9] wl[295] vdd gnd cell_6t
Xbit_r296_c9 bl[9] br[9] wl[296] vdd gnd cell_6t
Xbit_r297_c9 bl[9] br[9] wl[297] vdd gnd cell_6t
Xbit_r298_c9 bl[9] br[9] wl[298] vdd gnd cell_6t
Xbit_r299_c9 bl[9] br[9] wl[299] vdd gnd cell_6t
Xbit_r300_c9 bl[9] br[9] wl[300] vdd gnd cell_6t
Xbit_r301_c9 bl[9] br[9] wl[301] vdd gnd cell_6t
Xbit_r302_c9 bl[9] br[9] wl[302] vdd gnd cell_6t
Xbit_r303_c9 bl[9] br[9] wl[303] vdd gnd cell_6t
Xbit_r304_c9 bl[9] br[9] wl[304] vdd gnd cell_6t
Xbit_r305_c9 bl[9] br[9] wl[305] vdd gnd cell_6t
Xbit_r306_c9 bl[9] br[9] wl[306] vdd gnd cell_6t
Xbit_r307_c9 bl[9] br[9] wl[307] vdd gnd cell_6t
Xbit_r308_c9 bl[9] br[9] wl[308] vdd gnd cell_6t
Xbit_r309_c9 bl[9] br[9] wl[309] vdd gnd cell_6t
Xbit_r310_c9 bl[9] br[9] wl[310] vdd gnd cell_6t
Xbit_r311_c9 bl[9] br[9] wl[311] vdd gnd cell_6t
Xbit_r312_c9 bl[9] br[9] wl[312] vdd gnd cell_6t
Xbit_r313_c9 bl[9] br[9] wl[313] vdd gnd cell_6t
Xbit_r314_c9 bl[9] br[9] wl[314] vdd gnd cell_6t
Xbit_r315_c9 bl[9] br[9] wl[315] vdd gnd cell_6t
Xbit_r316_c9 bl[9] br[9] wl[316] vdd gnd cell_6t
Xbit_r317_c9 bl[9] br[9] wl[317] vdd gnd cell_6t
Xbit_r318_c9 bl[9] br[9] wl[318] vdd gnd cell_6t
Xbit_r319_c9 bl[9] br[9] wl[319] vdd gnd cell_6t
Xbit_r320_c9 bl[9] br[9] wl[320] vdd gnd cell_6t
Xbit_r321_c9 bl[9] br[9] wl[321] vdd gnd cell_6t
Xbit_r322_c9 bl[9] br[9] wl[322] vdd gnd cell_6t
Xbit_r323_c9 bl[9] br[9] wl[323] vdd gnd cell_6t
Xbit_r324_c9 bl[9] br[9] wl[324] vdd gnd cell_6t
Xbit_r325_c9 bl[9] br[9] wl[325] vdd gnd cell_6t
Xbit_r326_c9 bl[9] br[9] wl[326] vdd gnd cell_6t
Xbit_r327_c9 bl[9] br[9] wl[327] vdd gnd cell_6t
Xbit_r328_c9 bl[9] br[9] wl[328] vdd gnd cell_6t
Xbit_r329_c9 bl[9] br[9] wl[329] vdd gnd cell_6t
Xbit_r330_c9 bl[9] br[9] wl[330] vdd gnd cell_6t
Xbit_r331_c9 bl[9] br[9] wl[331] vdd gnd cell_6t
Xbit_r332_c9 bl[9] br[9] wl[332] vdd gnd cell_6t
Xbit_r333_c9 bl[9] br[9] wl[333] vdd gnd cell_6t
Xbit_r334_c9 bl[9] br[9] wl[334] vdd gnd cell_6t
Xbit_r335_c9 bl[9] br[9] wl[335] vdd gnd cell_6t
Xbit_r336_c9 bl[9] br[9] wl[336] vdd gnd cell_6t
Xbit_r337_c9 bl[9] br[9] wl[337] vdd gnd cell_6t
Xbit_r338_c9 bl[9] br[9] wl[338] vdd gnd cell_6t
Xbit_r339_c9 bl[9] br[9] wl[339] vdd gnd cell_6t
Xbit_r340_c9 bl[9] br[9] wl[340] vdd gnd cell_6t
Xbit_r341_c9 bl[9] br[9] wl[341] vdd gnd cell_6t
Xbit_r342_c9 bl[9] br[9] wl[342] vdd gnd cell_6t
Xbit_r343_c9 bl[9] br[9] wl[343] vdd gnd cell_6t
Xbit_r344_c9 bl[9] br[9] wl[344] vdd gnd cell_6t
Xbit_r345_c9 bl[9] br[9] wl[345] vdd gnd cell_6t
Xbit_r346_c9 bl[9] br[9] wl[346] vdd gnd cell_6t
Xbit_r347_c9 bl[9] br[9] wl[347] vdd gnd cell_6t
Xbit_r348_c9 bl[9] br[9] wl[348] vdd gnd cell_6t
Xbit_r349_c9 bl[9] br[9] wl[349] vdd gnd cell_6t
Xbit_r350_c9 bl[9] br[9] wl[350] vdd gnd cell_6t
Xbit_r351_c9 bl[9] br[9] wl[351] vdd gnd cell_6t
Xbit_r352_c9 bl[9] br[9] wl[352] vdd gnd cell_6t
Xbit_r353_c9 bl[9] br[9] wl[353] vdd gnd cell_6t
Xbit_r354_c9 bl[9] br[9] wl[354] vdd gnd cell_6t
Xbit_r355_c9 bl[9] br[9] wl[355] vdd gnd cell_6t
Xbit_r356_c9 bl[9] br[9] wl[356] vdd gnd cell_6t
Xbit_r357_c9 bl[9] br[9] wl[357] vdd gnd cell_6t
Xbit_r358_c9 bl[9] br[9] wl[358] vdd gnd cell_6t
Xbit_r359_c9 bl[9] br[9] wl[359] vdd gnd cell_6t
Xbit_r360_c9 bl[9] br[9] wl[360] vdd gnd cell_6t
Xbit_r361_c9 bl[9] br[9] wl[361] vdd gnd cell_6t
Xbit_r362_c9 bl[9] br[9] wl[362] vdd gnd cell_6t
Xbit_r363_c9 bl[9] br[9] wl[363] vdd gnd cell_6t
Xbit_r364_c9 bl[9] br[9] wl[364] vdd gnd cell_6t
Xbit_r365_c9 bl[9] br[9] wl[365] vdd gnd cell_6t
Xbit_r366_c9 bl[9] br[9] wl[366] vdd gnd cell_6t
Xbit_r367_c9 bl[9] br[9] wl[367] vdd gnd cell_6t
Xbit_r368_c9 bl[9] br[9] wl[368] vdd gnd cell_6t
Xbit_r369_c9 bl[9] br[9] wl[369] vdd gnd cell_6t
Xbit_r370_c9 bl[9] br[9] wl[370] vdd gnd cell_6t
Xbit_r371_c9 bl[9] br[9] wl[371] vdd gnd cell_6t
Xbit_r372_c9 bl[9] br[9] wl[372] vdd gnd cell_6t
Xbit_r373_c9 bl[9] br[9] wl[373] vdd gnd cell_6t
Xbit_r374_c9 bl[9] br[9] wl[374] vdd gnd cell_6t
Xbit_r375_c9 bl[9] br[9] wl[375] vdd gnd cell_6t
Xbit_r376_c9 bl[9] br[9] wl[376] vdd gnd cell_6t
Xbit_r377_c9 bl[9] br[9] wl[377] vdd gnd cell_6t
Xbit_r378_c9 bl[9] br[9] wl[378] vdd gnd cell_6t
Xbit_r379_c9 bl[9] br[9] wl[379] vdd gnd cell_6t
Xbit_r380_c9 bl[9] br[9] wl[380] vdd gnd cell_6t
Xbit_r381_c9 bl[9] br[9] wl[381] vdd gnd cell_6t
Xbit_r382_c9 bl[9] br[9] wl[382] vdd gnd cell_6t
Xbit_r383_c9 bl[9] br[9] wl[383] vdd gnd cell_6t
Xbit_r384_c9 bl[9] br[9] wl[384] vdd gnd cell_6t
Xbit_r385_c9 bl[9] br[9] wl[385] vdd gnd cell_6t
Xbit_r386_c9 bl[9] br[9] wl[386] vdd gnd cell_6t
Xbit_r387_c9 bl[9] br[9] wl[387] vdd gnd cell_6t
Xbit_r388_c9 bl[9] br[9] wl[388] vdd gnd cell_6t
Xbit_r389_c9 bl[9] br[9] wl[389] vdd gnd cell_6t
Xbit_r390_c9 bl[9] br[9] wl[390] vdd gnd cell_6t
Xbit_r391_c9 bl[9] br[9] wl[391] vdd gnd cell_6t
Xbit_r392_c9 bl[9] br[9] wl[392] vdd gnd cell_6t
Xbit_r393_c9 bl[9] br[9] wl[393] vdd gnd cell_6t
Xbit_r394_c9 bl[9] br[9] wl[394] vdd gnd cell_6t
Xbit_r395_c9 bl[9] br[9] wl[395] vdd gnd cell_6t
Xbit_r396_c9 bl[9] br[9] wl[396] vdd gnd cell_6t
Xbit_r397_c9 bl[9] br[9] wl[397] vdd gnd cell_6t
Xbit_r398_c9 bl[9] br[9] wl[398] vdd gnd cell_6t
Xbit_r399_c9 bl[9] br[9] wl[399] vdd gnd cell_6t
Xbit_r400_c9 bl[9] br[9] wl[400] vdd gnd cell_6t
Xbit_r401_c9 bl[9] br[9] wl[401] vdd gnd cell_6t
Xbit_r402_c9 bl[9] br[9] wl[402] vdd gnd cell_6t
Xbit_r403_c9 bl[9] br[9] wl[403] vdd gnd cell_6t
Xbit_r404_c9 bl[9] br[9] wl[404] vdd gnd cell_6t
Xbit_r405_c9 bl[9] br[9] wl[405] vdd gnd cell_6t
Xbit_r406_c9 bl[9] br[9] wl[406] vdd gnd cell_6t
Xbit_r407_c9 bl[9] br[9] wl[407] vdd gnd cell_6t
Xbit_r408_c9 bl[9] br[9] wl[408] vdd gnd cell_6t
Xbit_r409_c9 bl[9] br[9] wl[409] vdd gnd cell_6t
Xbit_r410_c9 bl[9] br[9] wl[410] vdd gnd cell_6t
Xbit_r411_c9 bl[9] br[9] wl[411] vdd gnd cell_6t
Xbit_r412_c9 bl[9] br[9] wl[412] vdd gnd cell_6t
Xbit_r413_c9 bl[9] br[9] wl[413] vdd gnd cell_6t
Xbit_r414_c9 bl[9] br[9] wl[414] vdd gnd cell_6t
Xbit_r415_c9 bl[9] br[9] wl[415] vdd gnd cell_6t
Xbit_r416_c9 bl[9] br[9] wl[416] vdd gnd cell_6t
Xbit_r417_c9 bl[9] br[9] wl[417] vdd gnd cell_6t
Xbit_r418_c9 bl[9] br[9] wl[418] vdd gnd cell_6t
Xbit_r419_c9 bl[9] br[9] wl[419] vdd gnd cell_6t
Xbit_r420_c9 bl[9] br[9] wl[420] vdd gnd cell_6t
Xbit_r421_c9 bl[9] br[9] wl[421] vdd gnd cell_6t
Xbit_r422_c9 bl[9] br[9] wl[422] vdd gnd cell_6t
Xbit_r423_c9 bl[9] br[9] wl[423] vdd gnd cell_6t
Xbit_r424_c9 bl[9] br[9] wl[424] vdd gnd cell_6t
Xbit_r425_c9 bl[9] br[9] wl[425] vdd gnd cell_6t
Xbit_r426_c9 bl[9] br[9] wl[426] vdd gnd cell_6t
Xbit_r427_c9 bl[9] br[9] wl[427] vdd gnd cell_6t
Xbit_r428_c9 bl[9] br[9] wl[428] vdd gnd cell_6t
Xbit_r429_c9 bl[9] br[9] wl[429] vdd gnd cell_6t
Xbit_r430_c9 bl[9] br[9] wl[430] vdd gnd cell_6t
Xbit_r431_c9 bl[9] br[9] wl[431] vdd gnd cell_6t
Xbit_r432_c9 bl[9] br[9] wl[432] vdd gnd cell_6t
Xbit_r433_c9 bl[9] br[9] wl[433] vdd gnd cell_6t
Xbit_r434_c9 bl[9] br[9] wl[434] vdd gnd cell_6t
Xbit_r435_c9 bl[9] br[9] wl[435] vdd gnd cell_6t
Xbit_r436_c9 bl[9] br[9] wl[436] vdd gnd cell_6t
Xbit_r437_c9 bl[9] br[9] wl[437] vdd gnd cell_6t
Xbit_r438_c9 bl[9] br[9] wl[438] vdd gnd cell_6t
Xbit_r439_c9 bl[9] br[9] wl[439] vdd gnd cell_6t
Xbit_r440_c9 bl[9] br[9] wl[440] vdd gnd cell_6t
Xbit_r441_c9 bl[9] br[9] wl[441] vdd gnd cell_6t
Xbit_r442_c9 bl[9] br[9] wl[442] vdd gnd cell_6t
Xbit_r443_c9 bl[9] br[9] wl[443] vdd gnd cell_6t
Xbit_r444_c9 bl[9] br[9] wl[444] vdd gnd cell_6t
Xbit_r445_c9 bl[9] br[9] wl[445] vdd gnd cell_6t
Xbit_r446_c9 bl[9] br[9] wl[446] vdd gnd cell_6t
Xbit_r447_c9 bl[9] br[9] wl[447] vdd gnd cell_6t
Xbit_r448_c9 bl[9] br[9] wl[448] vdd gnd cell_6t
Xbit_r449_c9 bl[9] br[9] wl[449] vdd gnd cell_6t
Xbit_r450_c9 bl[9] br[9] wl[450] vdd gnd cell_6t
Xbit_r451_c9 bl[9] br[9] wl[451] vdd gnd cell_6t
Xbit_r452_c9 bl[9] br[9] wl[452] vdd gnd cell_6t
Xbit_r453_c9 bl[9] br[9] wl[453] vdd gnd cell_6t
Xbit_r454_c9 bl[9] br[9] wl[454] vdd gnd cell_6t
Xbit_r455_c9 bl[9] br[9] wl[455] vdd gnd cell_6t
Xbit_r456_c9 bl[9] br[9] wl[456] vdd gnd cell_6t
Xbit_r457_c9 bl[9] br[9] wl[457] vdd gnd cell_6t
Xbit_r458_c9 bl[9] br[9] wl[458] vdd gnd cell_6t
Xbit_r459_c9 bl[9] br[9] wl[459] vdd gnd cell_6t
Xbit_r460_c9 bl[9] br[9] wl[460] vdd gnd cell_6t
Xbit_r461_c9 bl[9] br[9] wl[461] vdd gnd cell_6t
Xbit_r462_c9 bl[9] br[9] wl[462] vdd gnd cell_6t
Xbit_r463_c9 bl[9] br[9] wl[463] vdd gnd cell_6t
Xbit_r464_c9 bl[9] br[9] wl[464] vdd gnd cell_6t
Xbit_r465_c9 bl[9] br[9] wl[465] vdd gnd cell_6t
Xbit_r466_c9 bl[9] br[9] wl[466] vdd gnd cell_6t
Xbit_r467_c9 bl[9] br[9] wl[467] vdd gnd cell_6t
Xbit_r468_c9 bl[9] br[9] wl[468] vdd gnd cell_6t
Xbit_r469_c9 bl[9] br[9] wl[469] vdd gnd cell_6t
Xbit_r470_c9 bl[9] br[9] wl[470] vdd gnd cell_6t
Xbit_r471_c9 bl[9] br[9] wl[471] vdd gnd cell_6t
Xbit_r472_c9 bl[9] br[9] wl[472] vdd gnd cell_6t
Xbit_r473_c9 bl[9] br[9] wl[473] vdd gnd cell_6t
Xbit_r474_c9 bl[9] br[9] wl[474] vdd gnd cell_6t
Xbit_r475_c9 bl[9] br[9] wl[475] vdd gnd cell_6t
Xbit_r476_c9 bl[9] br[9] wl[476] vdd gnd cell_6t
Xbit_r477_c9 bl[9] br[9] wl[477] vdd gnd cell_6t
Xbit_r478_c9 bl[9] br[9] wl[478] vdd gnd cell_6t
Xbit_r479_c9 bl[9] br[9] wl[479] vdd gnd cell_6t
Xbit_r480_c9 bl[9] br[9] wl[480] vdd gnd cell_6t
Xbit_r481_c9 bl[9] br[9] wl[481] vdd gnd cell_6t
Xbit_r482_c9 bl[9] br[9] wl[482] vdd gnd cell_6t
Xbit_r483_c9 bl[9] br[9] wl[483] vdd gnd cell_6t
Xbit_r484_c9 bl[9] br[9] wl[484] vdd gnd cell_6t
Xbit_r485_c9 bl[9] br[9] wl[485] vdd gnd cell_6t
Xbit_r486_c9 bl[9] br[9] wl[486] vdd gnd cell_6t
Xbit_r487_c9 bl[9] br[9] wl[487] vdd gnd cell_6t
Xbit_r488_c9 bl[9] br[9] wl[488] vdd gnd cell_6t
Xbit_r489_c9 bl[9] br[9] wl[489] vdd gnd cell_6t
Xbit_r490_c9 bl[9] br[9] wl[490] vdd gnd cell_6t
Xbit_r491_c9 bl[9] br[9] wl[491] vdd gnd cell_6t
Xbit_r492_c9 bl[9] br[9] wl[492] vdd gnd cell_6t
Xbit_r493_c9 bl[9] br[9] wl[493] vdd gnd cell_6t
Xbit_r494_c9 bl[9] br[9] wl[494] vdd gnd cell_6t
Xbit_r495_c9 bl[9] br[9] wl[495] vdd gnd cell_6t
Xbit_r496_c9 bl[9] br[9] wl[496] vdd gnd cell_6t
Xbit_r497_c9 bl[9] br[9] wl[497] vdd gnd cell_6t
Xbit_r498_c9 bl[9] br[9] wl[498] vdd gnd cell_6t
Xbit_r499_c9 bl[9] br[9] wl[499] vdd gnd cell_6t
Xbit_r500_c9 bl[9] br[9] wl[500] vdd gnd cell_6t
Xbit_r501_c9 bl[9] br[9] wl[501] vdd gnd cell_6t
Xbit_r502_c9 bl[9] br[9] wl[502] vdd gnd cell_6t
Xbit_r503_c9 bl[9] br[9] wl[503] vdd gnd cell_6t
Xbit_r504_c9 bl[9] br[9] wl[504] vdd gnd cell_6t
Xbit_r505_c9 bl[9] br[9] wl[505] vdd gnd cell_6t
Xbit_r506_c9 bl[9] br[9] wl[506] vdd gnd cell_6t
Xbit_r507_c9 bl[9] br[9] wl[507] vdd gnd cell_6t
Xbit_r508_c9 bl[9] br[9] wl[508] vdd gnd cell_6t
Xbit_r509_c9 bl[9] br[9] wl[509] vdd gnd cell_6t
Xbit_r510_c9 bl[9] br[9] wl[510] vdd gnd cell_6t
Xbit_r511_c9 bl[9] br[9] wl[511] vdd gnd cell_6t
Xbit_r0_c10 bl[10] br[10] wl[0] vdd gnd cell_6t
Xbit_r1_c10 bl[10] br[10] wl[1] vdd gnd cell_6t
Xbit_r2_c10 bl[10] br[10] wl[2] vdd gnd cell_6t
Xbit_r3_c10 bl[10] br[10] wl[3] vdd gnd cell_6t
Xbit_r4_c10 bl[10] br[10] wl[4] vdd gnd cell_6t
Xbit_r5_c10 bl[10] br[10] wl[5] vdd gnd cell_6t
Xbit_r6_c10 bl[10] br[10] wl[6] vdd gnd cell_6t
Xbit_r7_c10 bl[10] br[10] wl[7] vdd gnd cell_6t
Xbit_r8_c10 bl[10] br[10] wl[8] vdd gnd cell_6t
Xbit_r9_c10 bl[10] br[10] wl[9] vdd gnd cell_6t
Xbit_r10_c10 bl[10] br[10] wl[10] vdd gnd cell_6t
Xbit_r11_c10 bl[10] br[10] wl[11] vdd gnd cell_6t
Xbit_r12_c10 bl[10] br[10] wl[12] vdd gnd cell_6t
Xbit_r13_c10 bl[10] br[10] wl[13] vdd gnd cell_6t
Xbit_r14_c10 bl[10] br[10] wl[14] vdd gnd cell_6t
Xbit_r15_c10 bl[10] br[10] wl[15] vdd gnd cell_6t
Xbit_r16_c10 bl[10] br[10] wl[16] vdd gnd cell_6t
Xbit_r17_c10 bl[10] br[10] wl[17] vdd gnd cell_6t
Xbit_r18_c10 bl[10] br[10] wl[18] vdd gnd cell_6t
Xbit_r19_c10 bl[10] br[10] wl[19] vdd gnd cell_6t
Xbit_r20_c10 bl[10] br[10] wl[20] vdd gnd cell_6t
Xbit_r21_c10 bl[10] br[10] wl[21] vdd gnd cell_6t
Xbit_r22_c10 bl[10] br[10] wl[22] vdd gnd cell_6t
Xbit_r23_c10 bl[10] br[10] wl[23] vdd gnd cell_6t
Xbit_r24_c10 bl[10] br[10] wl[24] vdd gnd cell_6t
Xbit_r25_c10 bl[10] br[10] wl[25] vdd gnd cell_6t
Xbit_r26_c10 bl[10] br[10] wl[26] vdd gnd cell_6t
Xbit_r27_c10 bl[10] br[10] wl[27] vdd gnd cell_6t
Xbit_r28_c10 bl[10] br[10] wl[28] vdd gnd cell_6t
Xbit_r29_c10 bl[10] br[10] wl[29] vdd gnd cell_6t
Xbit_r30_c10 bl[10] br[10] wl[30] vdd gnd cell_6t
Xbit_r31_c10 bl[10] br[10] wl[31] vdd gnd cell_6t
Xbit_r32_c10 bl[10] br[10] wl[32] vdd gnd cell_6t
Xbit_r33_c10 bl[10] br[10] wl[33] vdd gnd cell_6t
Xbit_r34_c10 bl[10] br[10] wl[34] vdd gnd cell_6t
Xbit_r35_c10 bl[10] br[10] wl[35] vdd gnd cell_6t
Xbit_r36_c10 bl[10] br[10] wl[36] vdd gnd cell_6t
Xbit_r37_c10 bl[10] br[10] wl[37] vdd gnd cell_6t
Xbit_r38_c10 bl[10] br[10] wl[38] vdd gnd cell_6t
Xbit_r39_c10 bl[10] br[10] wl[39] vdd gnd cell_6t
Xbit_r40_c10 bl[10] br[10] wl[40] vdd gnd cell_6t
Xbit_r41_c10 bl[10] br[10] wl[41] vdd gnd cell_6t
Xbit_r42_c10 bl[10] br[10] wl[42] vdd gnd cell_6t
Xbit_r43_c10 bl[10] br[10] wl[43] vdd gnd cell_6t
Xbit_r44_c10 bl[10] br[10] wl[44] vdd gnd cell_6t
Xbit_r45_c10 bl[10] br[10] wl[45] vdd gnd cell_6t
Xbit_r46_c10 bl[10] br[10] wl[46] vdd gnd cell_6t
Xbit_r47_c10 bl[10] br[10] wl[47] vdd gnd cell_6t
Xbit_r48_c10 bl[10] br[10] wl[48] vdd gnd cell_6t
Xbit_r49_c10 bl[10] br[10] wl[49] vdd gnd cell_6t
Xbit_r50_c10 bl[10] br[10] wl[50] vdd gnd cell_6t
Xbit_r51_c10 bl[10] br[10] wl[51] vdd gnd cell_6t
Xbit_r52_c10 bl[10] br[10] wl[52] vdd gnd cell_6t
Xbit_r53_c10 bl[10] br[10] wl[53] vdd gnd cell_6t
Xbit_r54_c10 bl[10] br[10] wl[54] vdd gnd cell_6t
Xbit_r55_c10 bl[10] br[10] wl[55] vdd gnd cell_6t
Xbit_r56_c10 bl[10] br[10] wl[56] vdd gnd cell_6t
Xbit_r57_c10 bl[10] br[10] wl[57] vdd gnd cell_6t
Xbit_r58_c10 bl[10] br[10] wl[58] vdd gnd cell_6t
Xbit_r59_c10 bl[10] br[10] wl[59] vdd gnd cell_6t
Xbit_r60_c10 bl[10] br[10] wl[60] vdd gnd cell_6t
Xbit_r61_c10 bl[10] br[10] wl[61] vdd gnd cell_6t
Xbit_r62_c10 bl[10] br[10] wl[62] vdd gnd cell_6t
Xbit_r63_c10 bl[10] br[10] wl[63] vdd gnd cell_6t
Xbit_r64_c10 bl[10] br[10] wl[64] vdd gnd cell_6t
Xbit_r65_c10 bl[10] br[10] wl[65] vdd gnd cell_6t
Xbit_r66_c10 bl[10] br[10] wl[66] vdd gnd cell_6t
Xbit_r67_c10 bl[10] br[10] wl[67] vdd gnd cell_6t
Xbit_r68_c10 bl[10] br[10] wl[68] vdd gnd cell_6t
Xbit_r69_c10 bl[10] br[10] wl[69] vdd gnd cell_6t
Xbit_r70_c10 bl[10] br[10] wl[70] vdd gnd cell_6t
Xbit_r71_c10 bl[10] br[10] wl[71] vdd gnd cell_6t
Xbit_r72_c10 bl[10] br[10] wl[72] vdd gnd cell_6t
Xbit_r73_c10 bl[10] br[10] wl[73] vdd gnd cell_6t
Xbit_r74_c10 bl[10] br[10] wl[74] vdd gnd cell_6t
Xbit_r75_c10 bl[10] br[10] wl[75] vdd gnd cell_6t
Xbit_r76_c10 bl[10] br[10] wl[76] vdd gnd cell_6t
Xbit_r77_c10 bl[10] br[10] wl[77] vdd gnd cell_6t
Xbit_r78_c10 bl[10] br[10] wl[78] vdd gnd cell_6t
Xbit_r79_c10 bl[10] br[10] wl[79] vdd gnd cell_6t
Xbit_r80_c10 bl[10] br[10] wl[80] vdd gnd cell_6t
Xbit_r81_c10 bl[10] br[10] wl[81] vdd gnd cell_6t
Xbit_r82_c10 bl[10] br[10] wl[82] vdd gnd cell_6t
Xbit_r83_c10 bl[10] br[10] wl[83] vdd gnd cell_6t
Xbit_r84_c10 bl[10] br[10] wl[84] vdd gnd cell_6t
Xbit_r85_c10 bl[10] br[10] wl[85] vdd gnd cell_6t
Xbit_r86_c10 bl[10] br[10] wl[86] vdd gnd cell_6t
Xbit_r87_c10 bl[10] br[10] wl[87] vdd gnd cell_6t
Xbit_r88_c10 bl[10] br[10] wl[88] vdd gnd cell_6t
Xbit_r89_c10 bl[10] br[10] wl[89] vdd gnd cell_6t
Xbit_r90_c10 bl[10] br[10] wl[90] vdd gnd cell_6t
Xbit_r91_c10 bl[10] br[10] wl[91] vdd gnd cell_6t
Xbit_r92_c10 bl[10] br[10] wl[92] vdd gnd cell_6t
Xbit_r93_c10 bl[10] br[10] wl[93] vdd gnd cell_6t
Xbit_r94_c10 bl[10] br[10] wl[94] vdd gnd cell_6t
Xbit_r95_c10 bl[10] br[10] wl[95] vdd gnd cell_6t
Xbit_r96_c10 bl[10] br[10] wl[96] vdd gnd cell_6t
Xbit_r97_c10 bl[10] br[10] wl[97] vdd gnd cell_6t
Xbit_r98_c10 bl[10] br[10] wl[98] vdd gnd cell_6t
Xbit_r99_c10 bl[10] br[10] wl[99] vdd gnd cell_6t
Xbit_r100_c10 bl[10] br[10] wl[100] vdd gnd cell_6t
Xbit_r101_c10 bl[10] br[10] wl[101] vdd gnd cell_6t
Xbit_r102_c10 bl[10] br[10] wl[102] vdd gnd cell_6t
Xbit_r103_c10 bl[10] br[10] wl[103] vdd gnd cell_6t
Xbit_r104_c10 bl[10] br[10] wl[104] vdd gnd cell_6t
Xbit_r105_c10 bl[10] br[10] wl[105] vdd gnd cell_6t
Xbit_r106_c10 bl[10] br[10] wl[106] vdd gnd cell_6t
Xbit_r107_c10 bl[10] br[10] wl[107] vdd gnd cell_6t
Xbit_r108_c10 bl[10] br[10] wl[108] vdd gnd cell_6t
Xbit_r109_c10 bl[10] br[10] wl[109] vdd gnd cell_6t
Xbit_r110_c10 bl[10] br[10] wl[110] vdd gnd cell_6t
Xbit_r111_c10 bl[10] br[10] wl[111] vdd gnd cell_6t
Xbit_r112_c10 bl[10] br[10] wl[112] vdd gnd cell_6t
Xbit_r113_c10 bl[10] br[10] wl[113] vdd gnd cell_6t
Xbit_r114_c10 bl[10] br[10] wl[114] vdd gnd cell_6t
Xbit_r115_c10 bl[10] br[10] wl[115] vdd gnd cell_6t
Xbit_r116_c10 bl[10] br[10] wl[116] vdd gnd cell_6t
Xbit_r117_c10 bl[10] br[10] wl[117] vdd gnd cell_6t
Xbit_r118_c10 bl[10] br[10] wl[118] vdd gnd cell_6t
Xbit_r119_c10 bl[10] br[10] wl[119] vdd gnd cell_6t
Xbit_r120_c10 bl[10] br[10] wl[120] vdd gnd cell_6t
Xbit_r121_c10 bl[10] br[10] wl[121] vdd gnd cell_6t
Xbit_r122_c10 bl[10] br[10] wl[122] vdd gnd cell_6t
Xbit_r123_c10 bl[10] br[10] wl[123] vdd gnd cell_6t
Xbit_r124_c10 bl[10] br[10] wl[124] vdd gnd cell_6t
Xbit_r125_c10 bl[10] br[10] wl[125] vdd gnd cell_6t
Xbit_r126_c10 bl[10] br[10] wl[126] vdd gnd cell_6t
Xbit_r127_c10 bl[10] br[10] wl[127] vdd gnd cell_6t
Xbit_r128_c10 bl[10] br[10] wl[128] vdd gnd cell_6t
Xbit_r129_c10 bl[10] br[10] wl[129] vdd gnd cell_6t
Xbit_r130_c10 bl[10] br[10] wl[130] vdd gnd cell_6t
Xbit_r131_c10 bl[10] br[10] wl[131] vdd gnd cell_6t
Xbit_r132_c10 bl[10] br[10] wl[132] vdd gnd cell_6t
Xbit_r133_c10 bl[10] br[10] wl[133] vdd gnd cell_6t
Xbit_r134_c10 bl[10] br[10] wl[134] vdd gnd cell_6t
Xbit_r135_c10 bl[10] br[10] wl[135] vdd gnd cell_6t
Xbit_r136_c10 bl[10] br[10] wl[136] vdd gnd cell_6t
Xbit_r137_c10 bl[10] br[10] wl[137] vdd gnd cell_6t
Xbit_r138_c10 bl[10] br[10] wl[138] vdd gnd cell_6t
Xbit_r139_c10 bl[10] br[10] wl[139] vdd gnd cell_6t
Xbit_r140_c10 bl[10] br[10] wl[140] vdd gnd cell_6t
Xbit_r141_c10 bl[10] br[10] wl[141] vdd gnd cell_6t
Xbit_r142_c10 bl[10] br[10] wl[142] vdd gnd cell_6t
Xbit_r143_c10 bl[10] br[10] wl[143] vdd gnd cell_6t
Xbit_r144_c10 bl[10] br[10] wl[144] vdd gnd cell_6t
Xbit_r145_c10 bl[10] br[10] wl[145] vdd gnd cell_6t
Xbit_r146_c10 bl[10] br[10] wl[146] vdd gnd cell_6t
Xbit_r147_c10 bl[10] br[10] wl[147] vdd gnd cell_6t
Xbit_r148_c10 bl[10] br[10] wl[148] vdd gnd cell_6t
Xbit_r149_c10 bl[10] br[10] wl[149] vdd gnd cell_6t
Xbit_r150_c10 bl[10] br[10] wl[150] vdd gnd cell_6t
Xbit_r151_c10 bl[10] br[10] wl[151] vdd gnd cell_6t
Xbit_r152_c10 bl[10] br[10] wl[152] vdd gnd cell_6t
Xbit_r153_c10 bl[10] br[10] wl[153] vdd gnd cell_6t
Xbit_r154_c10 bl[10] br[10] wl[154] vdd gnd cell_6t
Xbit_r155_c10 bl[10] br[10] wl[155] vdd gnd cell_6t
Xbit_r156_c10 bl[10] br[10] wl[156] vdd gnd cell_6t
Xbit_r157_c10 bl[10] br[10] wl[157] vdd gnd cell_6t
Xbit_r158_c10 bl[10] br[10] wl[158] vdd gnd cell_6t
Xbit_r159_c10 bl[10] br[10] wl[159] vdd gnd cell_6t
Xbit_r160_c10 bl[10] br[10] wl[160] vdd gnd cell_6t
Xbit_r161_c10 bl[10] br[10] wl[161] vdd gnd cell_6t
Xbit_r162_c10 bl[10] br[10] wl[162] vdd gnd cell_6t
Xbit_r163_c10 bl[10] br[10] wl[163] vdd gnd cell_6t
Xbit_r164_c10 bl[10] br[10] wl[164] vdd gnd cell_6t
Xbit_r165_c10 bl[10] br[10] wl[165] vdd gnd cell_6t
Xbit_r166_c10 bl[10] br[10] wl[166] vdd gnd cell_6t
Xbit_r167_c10 bl[10] br[10] wl[167] vdd gnd cell_6t
Xbit_r168_c10 bl[10] br[10] wl[168] vdd gnd cell_6t
Xbit_r169_c10 bl[10] br[10] wl[169] vdd gnd cell_6t
Xbit_r170_c10 bl[10] br[10] wl[170] vdd gnd cell_6t
Xbit_r171_c10 bl[10] br[10] wl[171] vdd gnd cell_6t
Xbit_r172_c10 bl[10] br[10] wl[172] vdd gnd cell_6t
Xbit_r173_c10 bl[10] br[10] wl[173] vdd gnd cell_6t
Xbit_r174_c10 bl[10] br[10] wl[174] vdd gnd cell_6t
Xbit_r175_c10 bl[10] br[10] wl[175] vdd gnd cell_6t
Xbit_r176_c10 bl[10] br[10] wl[176] vdd gnd cell_6t
Xbit_r177_c10 bl[10] br[10] wl[177] vdd gnd cell_6t
Xbit_r178_c10 bl[10] br[10] wl[178] vdd gnd cell_6t
Xbit_r179_c10 bl[10] br[10] wl[179] vdd gnd cell_6t
Xbit_r180_c10 bl[10] br[10] wl[180] vdd gnd cell_6t
Xbit_r181_c10 bl[10] br[10] wl[181] vdd gnd cell_6t
Xbit_r182_c10 bl[10] br[10] wl[182] vdd gnd cell_6t
Xbit_r183_c10 bl[10] br[10] wl[183] vdd gnd cell_6t
Xbit_r184_c10 bl[10] br[10] wl[184] vdd gnd cell_6t
Xbit_r185_c10 bl[10] br[10] wl[185] vdd gnd cell_6t
Xbit_r186_c10 bl[10] br[10] wl[186] vdd gnd cell_6t
Xbit_r187_c10 bl[10] br[10] wl[187] vdd gnd cell_6t
Xbit_r188_c10 bl[10] br[10] wl[188] vdd gnd cell_6t
Xbit_r189_c10 bl[10] br[10] wl[189] vdd gnd cell_6t
Xbit_r190_c10 bl[10] br[10] wl[190] vdd gnd cell_6t
Xbit_r191_c10 bl[10] br[10] wl[191] vdd gnd cell_6t
Xbit_r192_c10 bl[10] br[10] wl[192] vdd gnd cell_6t
Xbit_r193_c10 bl[10] br[10] wl[193] vdd gnd cell_6t
Xbit_r194_c10 bl[10] br[10] wl[194] vdd gnd cell_6t
Xbit_r195_c10 bl[10] br[10] wl[195] vdd gnd cell_6t
Xbit_r196_c10 bl[10] br[10] wl[196] vdd gnd cell_6t
Xbit_r197_c10 bl[10] br[10] wl[197] vdd gnd cell_6t
Xbit_r198_c10 bl[10] br[10] wl[198] vdd gnd cell_6t
Xbit_r199_c10 bl[10] br[10] wl[199] vdd gnd cell_6t
Xbit_r200_c10 bl[10] br[10] wl[200] vdd gnd cell_6t
Xbit_r201_c10 bl[10] br[10] wl[201] vdd gnd cell_6t
Xbit_r202_c10 bl[10] br[10] wl[202] vdd gnd cell_6t
Xbit_r203_c10 bl[10] br[10] wl[203] vdd gnd cell_6t
Xbit_r204_c10 bl[10] br[10] wl[204] vdd gnd cell_6t
Xbit_r205_c10 bl[10] br[10] wl[205] vdd gnd cell_6t
Xbit_r206_c10 bl[10] br[10] wl[206] vdd gnd cell_6t
Xbit_r207_c10 bl[10] br[10] wl[207] vdd gnd cell_6t
Xbit_r208_c10 bl[10] br[10] wl[208] vdd gnd cell_6t
Xbit_r209_c10 bl[10] br[10] wl[209] vdd gnd cell_6t
Xbit_r210_c10 bl[10] br[10] wl[210] vdd gnd cell_6t
Xbit_r211_c10 bl[10] br[10] wl[211] vdd gnd cell_6t
Xbit_r212_c10 bl[10] br[10] wl[212] vdd gnd cell_6t
Xbit_r213_c10 bl[10] br[10] wl[213] vdd gnd cell_6t
Xbit_r214_c10 bl[10] br[10] wl[214] vdd gnd cell_6t
Xbit_r215_c10 bl[10] br[10] wl[215] vdd gnd cell_6t
Xbit_r216_c10 bl[10] br[10] wl[216] vdd gnd cell_6t
Xbit_r217_c10 bl[10] br[10] wl[217] vdd gnd cell_6t
Xbit_r218_c10 bl[10] br[10] wl[218] vdd gnd cell_6t
Xbit_r219_c10 bl[10] br[10] wl[219] vdd gnd cell_6t
Xbit_r220_c10 bl[10] br[10] wl[220] vdd gnd cell_6t
Xbit_r221_c10 bl[10] br[10] wl[221] vdd gnd cell_6t
Xbit_r222_c10 bl[10] br[10] wl[222] vdd gnd cell_6t
Xbit_r223_c10 bl[10] br[10] wl[223] vdd gnd cell_6t
Xbit_r224_c10 bl[10] br[10] wl[224] vdd gnd cell_6t
Xbit_r225_c10 bl[10] br[10] wl[225] vdd gnd cell_6t
Xbit_r226_c10 bl[10] br[10] wl[226] vdd gnd cell_6t
Xbit_r227_c10 bl[10] br[10] wl[227] vdd gnd cell_6t
Xbit_r228_c10 bl[10] br[10] wl[228] vdd gnd cell_6t
Xbit_r229_c10 bl[10] br[10] wl[229] vdd gnd cell_6t
Xbit_r230_c10 bl[10] br[10] wl[230] vdd gnd cell_6t
Xbit_r231_c10 bl[10] br[10] wl[231] vdd gnd cell_6t
Xbit_r232_c10 bl[10] br[10] wl[232] vdd gnd cell_6t
Xbit_r233_c10 bl[10] br[10] wl[233] vdd gnd cell_6t
Xbit_r234_c10 bl[10] br[10] wl[234] vdd gnd cell_6t
Xbit_r235_c10 bl[10] br[10] wl[235] vdd gnd cell_6t
Xbit_r236_c10 bl[10] br[10] wl[236] vdd gnd cell_6t
Xbit_r237_c10 bl[10] br[10] wl[237] vdd gnd cell_6t
Xbit_r238_c10 bl[10] br[10] wl[238] vdd gnd cell_6t
Xbit_r239_c10 bl[10] br[10] wl[239] vdd gnd cell_6t
Xbit_r240_c10 bl[10] br[10] wl[240] vdd gnd cell_6t
Xbit_r241_c10 bl[10] br[10] wl[241] vdd gnd cell_6t
Xbit_r242_c10 bl[10] br[10] wl[242] vdd gnd cell_6t
Xbit_r243_c10 bl[10] br[10] wl[243] vdd gnd cell_6t
Xbit_r244_c10 bl[10] br[10] wl[244] vdd gnd cell_6t
Xbit_r245_c10 bl[10] br[10] wl[245] vdd gnd cell_6t
Xbit_r246_c10 bl[10] br[10] wl[246] vdd gnd cell_6t
Xbit_r247_c10 bl[10] br[10] wl[247] vdd gnd cell_6t
Xbit_r248_c10 bl[10] br[10] wl[248] vdd gnd cell_6t
Xbit_r249_c10 bl[10] br[10] wl[249] vdd gnd cell_6t
Xbit_r250_c10 bl[10] br[10] wl[250] vdd gnd cell_6t
Xbit_r251_c10 bl[10] br[10] wl[251] vdd gnd cell_6t
Xbit_r252_c10 bl[10] br[10] wl[252] vdd gnd cell_6t
Xbit_r253_c10 bl[10] br[10] wl[253] vdd gnd cell_6t
Xbit_r254_c10 bl[10] br[10] wl[254] vdd gnd cell_6t
Xbit_r255_c10 bl[10] br[10] wl[255] vdd gnd cell_6t
Xbit_r256_c10 bl[10] br[10] wl[256] vdd gnd cell_6t
Xbit_r257_c10 bl[10] br[10] wl[257] vdd gnd cell_6t
Xbit_r258_c10 bl[10] br[10] wl[258] vdd gnd cell_6t
Xbit_r259_c10 bl[10] br[10] wl[259] vdd gnd cell_6t
Xbit_r260_c10 bl[10] br[10] wl[260] vdd gnd cell_6t
Xbit_r261_c10 bl[10] br[10] wl[261] vdd gnd cell_6t
Xbit_r262_c10 bl[10] br[10] wl[262] vdd gnd cell_6t
Xbit_r263_c10 bl[10] br[10] wl[263] vdd gnd cell_6t
Xbit_r264_c10 bl[10] br[10] wl[264] vdd gnd cell_6t
Xbit_r265_c10 bl[10] br[10] wl[265] vdd gnd cell_6t
Xbit_r266_c10 bl[10] br[10] wl[266] vdd gnd cell_6t
Xbit_r267_c10 bl[10] br[10] wl[267] vdd gnd cell_6t
Xbit_r268_c10 bl[10] br[10] wl[268] vdd gnd cell_6t
Xbit_r269_c10 bl[10] br[10] wl[269] vdd gnd cell_6t
Xbit_r270_c10 bl[10] br[10] wl[270] vdd gnd cell_6t
Xbit_r271_c10 bl[10] br[10] wl[271] vdd gnd cell_6t
Xbit_r272_c10 bl[10] br[10] wl[272] vdd gnd cell_6t
Xbit_r273_c10 bl[10] br[10] wl[273] vdd gnd cell_6t
Xbit_r274_c10 bl[10] br[10] wl[274] vdd gnd cell_6t
Xbit_r275_c10 bl[10] br[10] wl[275] vdd gnd cell_6t
Xbit_r276_c10 bl[10] br[10] wl[276] vdd gnd cell_6t
Xbit_r277_c10 bl[10] br[10] wl[277] vdd gnd cell_6t
Xbit_r278_c10 bl[10] br[10] wl[278] vdd gnd cell_6t
Xbit_r279_c10 bl[10] br[10] wl[279] vdd gnd cell_6t
Xbit_r280_c10 bl[10] br[10] wl[280] vdd gnd cell_6t
Xbit_r281_c10 bl[10] br[10] wl[281] vdd gnd cell_6t
Xbit_r282_c10 bl[10] br[10] wl[282] vdd gnd cell_6t
Xbit_r283_c10 bl[10] br[10] wl[283] vdd gnd cell_6t
Xbit_r284_c10 bl[10] br[10] wl[284] vdd gnd cell_6t
Xbit_r285_c10 bl[10] br[10] wl[285] vdd gnd cell_6t
Xbit_r286_c10 bl[10] br[10] wl[286] vdd gnd cell_6t
Xbit_r287_c10 bl[10] br[10] wl[287] vdd gnd cell_6t
Xbit_r288_c10 bl[10] br[10] wl[288] vdd gnd cell_6t
Xbit_r289_c10 bl[10] br[10] wl[289] vdd gnd cell_6t
Xbit_r290_c10 bl[10] br[10] wl[290] vdd gnd cell_6t
Xbit_r291_c10 bl[10] br[10] wl[291] vdd gnd cell_6t
Xbit_r292_c10 bl[10] br[10] wl[292] vdd gnd cell_6t
Xbit_r293_c10 bl[10] br[10] wl[293] vdd gnd cell_6t
Xbit_r294_c10 bl[10] br[10] wl[294] vdd gnd cell_6t
Xbit_r295_c10 bl[10] br[10] wl[295] vdd gnd cell_6t
Xbit_r296_c10 bl[10] br[10] wl[296] vdd gnd cell_6t
Xbit_r297_c10 bl[10] br[10] wl[297] vdd gnd cell_6t
Xbit_r298_c10 bl[10] br[10] wl[298] vdd gnd cell_6t
Xbit_r299_c10 bl[10] br[10] wl[299] vdd gnd cell_6t
Xbit_r300_c10 bl[10] br[10] wl[300] vdd gnd cell_6t
Xbit_r301_c10 bl[10] br[10] wl[301] vdd gnd cell_6t
Xbit_r302_c10 bl[10] br[10] wl[302] vdd gnd cell_6t
Xbit_r303_c10 bl[10] br[10] wl[303] vdd gnd cell_6t
Xbit_r304_c10 bl[10] br[10] wl[304] vdd gnd cell_6t
Xbit_r305_c10 bl[10] br[10] wl[305] vdd gnd cell_6t
Xbit_r306_c10 bl[10] br[10] wl[306] vdd gnd cell_6t
Xbit_r307_c10 bl[10] br[10] wl[307] vdd gnd cell_6t
Xbit_r308_c10 bl[10] br[10] wl[308] vdd gnd cell_6t
Xbit_r309_c10 bl[10] br[10] wl[309] vdd gnd cell_6t
Xbit_r310_c10 bl[10] br[10] wl[310] vdd gnd cell_6t
Xbit_r311_c10 bl[10] br[10] wl[311] vdd gnd cell_6t
Xbit_r312_c10 bl[10] br[10] wl[312] vdd gnd cell_6t
Xbit_r313_c10 bl[10] br[10] wl[313] vdd gnd cell_6t
Xbit_r314_c10 bl[10] br[10] wl[314] vdd gnd cell_6t
Xbit_r315_c10 bl[10] br[10] wl[315] vdd gnd cell_6t
Xbit_r316_c10 bl[10] br[10] wl[316] vdd gnd cell_6t
Xbit_r317_c10 bl[10] br[10] wl[317] vdd gnd cell_6t
Xbit_r318_c10 bl[10] br[10] wl[318] vdd gnd cell_6t
Xbit_r319_c10 bl[10] br[10] wl[319] vdd gnd cell_6t
Xbit_r320_c10 bl[10] br[10] wl[320] vdd gnd cell_6t
Xbit_r321_c10 bl[10] br[10] wl[321] vdd gnd cell_6t
Xbit_r322_c10 bl[10] br[10] wl[322] vdd gnd cell_6t
Xbit_r323_c10 bl[10] br[10] wl[323] vdd gnd cell_6t
Xbit_r324_c10 bl[10] br[10] wl[324] vdd gnd cell_6t
Xbit_r325_c10 bl[10] br[10] wl[325] vdd gnd cell_6t
Xbit_r326_c10 bl[10] br[10] wl[326] vdd gnd cell_6t
Xbit_r327_c10 bl[10] br[10] wl[327] vdd gnd cell_6t
Xbit_r328_c10 bl[10] br[10] wl[328] vdd gnd cell_6t
Xbit_r329_c10 bl[10] br[10] wl[329] vdd gnd cell_6t
Xbit_r330_c10 bl[10] br[10] wl[330] vdd gnd cell_6t
Xbit_r331_c10 bl[10] br[10] wl[331] vdd gnd cell_6t
Xbit_r332_c10 bl[10] br[10] wl[332] vdd gnd cell_6t
Xbit_r333_c10 bl[10] br[10] wl[333] vdd gnd cell_6t
Xbit_r334_c10 bl[10] br[10] wl[334] vdd gnd cell_6t
Xbit_r335_c10 bl[10] br[10] wl[335] vdd gnd cell_6t
Xbit_r336_c10 bl[10] br[10] wl[336] vdd gnd cell_6t
Xbit_r337_c10 bl[10] br[10] wl[337] vdd gnd cell_6t
Xbit_r338_c10 bl[10] br[10] wl[338] vdd gnd cell_6t
Xbit_r339_c10 bl[10] br[10] wl[339] vdd gnd cell_6t
Xbit_r340_c10 bl[10] br[10] wl[340] vdd gnd cell_6t
Xbit_r341_c10 bl[10] br[10] wl[341] vdd gnd cell_6t
Xbit_r342_c10 bl[10] br[10] wl[342] vdd gnd cell_6t
Xbit_r343_c10 bl[10] br[10] wl[343] vdd gnd cell_6t
Xbit_r344_c10 bl[10] br[10] wl[344] vdd gnd cell_6t
Xbit_r345_c10 bl[10] br[10] wl[345] vdd gnd cell_6t
Xbit_r346_c10 bl[10] br[10] wl[346] vdd gnd cell_6t
Xbit_r347_c10 bl[10] br[10] wl[347] vdd gnd cell_6t
Xbit_r348_c10 bl[10] br[10] wl[348] vdd gnd cell_6t
Xbit_r349_c10 bl[10] br[10] wl[349] vdd gnd cell_6t
Xbit_r350_c10 bl[10] br[10] wl[350] vdd gnd cell_6t
Xbit_r351_c10 bl[10] br[10] wl[351] vdd gnd cell_6t
Xbit_r352_c10 bl[10] br[10] wl[352] vdd gnd cell_6t
Xbit_r353_c10 bl[10] br[10] wl[353] vdd gnd cell_6t
Xbit_r354_c10 bl[10] br[10] wl[354] vdd gnd cell_6t
Xbit_r355_c10 bl[10] br[10] wl[355] vdd gnd cell_6t
Xbit_r356_c10 bl[10] br[10] wl[356] vdd gnd cell_6t
Xbit_r357_c10 bl[10] br[10] wl[357] vdd gnd cell_6t
Xbit_r358_c10 bl[10] br[10] wl[358] vdd gnd cell_6t
Xbit_r359_c10 bl[10] br[10] wl[359] vdd gnd cell_6t
Xbit_r360_c10 bl[10] br[10] wl[360] vdd gnd cell_6t
Xbit_r361_c10 bl[10] br[10] wl[361] vdd gnd cell_6t
Xbit_r362_c10 bl[10] br[10] wl[362] vdd gnd cell_6t
Xbit_r363_c10 bl[10] br[10] wl[363] vdd gnd cell_6t
Xbit_r364_c10 bl[10] br[10] wl[364] vdd gnd cell_6t
Xbit_r365_c10 bl[10] br[10] wl[365] vdd gnd cell_6t
Xbit_r366_c10 bl[10] br[10] wl[366] vdd gnd cell_6t
Xbit_r367_c10 bl[10] br[10] wl[367] vdd gnd cell_6t
Xbit_r368_c10 bl[10] br[10] wl[368] vdd gnd cell_6t
Xbit_r369_c10 bl[10] br[10] wl[369] vdd gnd cell_6t
Xbit_r370_c10 bl[10] br[10] wl[370] vdd gnd cell_6t
Xbit_r371_c10 bl[10] br[10] wl[371] vdd gnd cell_6t
Xbit_r372_c10 bl[10] br[10] wl[372] vdd gnd cell_6t
Xbit_r373_c10 bl[10] br[10] wl[373] vdd gnd cell_6t
Xbit_r374_c10 bl[10] br[10] wl[374] vdd gnd cell_6t
Xbit_r375_c10 bl[10] br[10] wl[375] vdd gnd cell_6t
Xbit_r376_c10 bl[10] br[10] wl[376] vdd gnd cell_6t
Xbit_r377_c10 bl[10] br[10] wl[377] vdd gnd cell_6t
Xbit_r378_c10 bl[10] br[10] wl[378] vdd gnd cell_6t
Xbit_r379_c10 bl[10] br[10] wl[379] vdd gnd cell_6t
Xbit_r380_c10 bl[10] br[10] wl[380] vdd gnd cell_6t
Xbit_r381_c10 bl[10] br[10] wl[381] vdd gnd cell_6t
Xbit_r382_c10 bl[10] br[10] wl[382] vdd gnd cell_6t
Xbit_r383_c10 bl[10] br[10] wl[383] vdd gnd cell_6t
Xbit_r384_c10 bl[10] br[10] wl[384] vdd gnd cell_6t
Xbit_r385_c10 bl[10] br[10] wl[385] vdd gnd cell_6t
Xbit_r386_c10 bl[10] br[10] wl[386] vdd gnd cell_6t
Xbit_r387_c10 bl[10] br[10] wl[387] vdd gnd cell_6t
Xbit_r388_c10 bl[10] br[10] wl[388] vdd gnd cell_6t
Xbit_r389_c10 bl[10] br[10] wl[389] vdd gnd cell_6t
Xbit_r390_c10 bl[10] br[10] wl[390] vdd gnd cell_6t
Xbit_r391_c10 bl[10] br[10] wl[391] vdd gnd cell_6t
Xbit_r392_c10 bl[10] br[10] wl[392] vdd gnd cell_6t
Xbit_r393_c10 bl[10] br[10] wl[393] vdd gnd cell_6t
Xbit_r394_c10 bl[10] br[10] wl[394] vdd gnd cell_6t
Xbit_r395_c10 bl[10] br[10] wl[395] vdd gnd cell_6t
Xbit_r396_c10 bl[10] br[10] wl[396] vdd gnd cell_6t
Xbit_r397_c10 bl[10] br[10] wl[397] vdd gnd cell_6t
Xbit_r398_c10 bl[10] br[10] wl[398] vdd gnd cell_6t
Xbit_r399_c10 bl[10] br[10] wl[399] vdd gnd cell_6t
Xbit_r400_c10 bl[10] br[10] wl[400] vdd gnd cell_6t
Xbit_r401_c10 bl[10] br[10] wl[401] vdd gnd cell_6t
Xbit_r402_c10 bl[10] br[10] wl[402] vdd gnd cell_6t
Xbit_r403_c10 bl[10] br[10] wl[403] vdd gnd cell_6t
Xbit_r404_c10 bl[10] br[10] wl[404] vdd gnd cell_6t
Xbit_r405_c10 bl[10] br[10] wl[405] vdd gnd cell_6t
Xbit_r406_c10 bl[10] br[10] wl[406] vdd gnd cell_6t
Xbit_r407_c10 bl[10] br[10] wl[407] vdd gnd cell_6t
Xbit_r408_c10 bl[10] br[10] wl[408] vdd gnd cell_6t
Xbit_r409_c10 bl[10] br[10] wl[409] vdd gnd cell_6t
Xbit_r410_c10 bl[10] br[10] wl[410] vdd gnd cell_6t
Xbit_r411_c10 bl[10] br[10] wl[411] vdd gnd cell_6t
Xbit_r412_c10 bl[10] br[10] wl[412] vdd gnd cell_6t
Xbit_r413_c10 bl[10] br[10] wl[413] vdd gnd cell_6t
Xbit_r414_c10 bl[10] br[10] wl[414] vdd gnd cell_6t
Xbit_r415_c10 bl[10] br[10] wl[415] vdd gnd cell_6t
Xbit_r416_c10 bl[10] br[10] wl[416] vdd gnd cell_6t
Xbit_r417_c10 bl[10] br[10] wl[417] vdd gnd cell_6t
Xbit_r418_c10 bl[10] br[10] wl[418] vdd gnd cell_6t
Xbit_r419_c10 bl[10] br[10] wl[419] vdd gnd cell_6t
Xbit_r420_c10 bl[10] br[10] wl[420] vdd gnd cell_6t
Xbit_r421_c10 bl[10] br[10] wl[421] vdd gnd cell_6t
Xbit_r422_c10 bl[10] br[10] wl[422] vdd gnd cell_6t
Xbit_r423_c10 bl[10] br[10] wl[423] vdd gnd cell_6t
Xbit_r424_c10 bl[10] br[10] wl[424] vdd gnd cell_6t
Xbit_r425_c10 bl[10] br[10] wl[425] vdd gnd cell_6t
Xbit_r426_c10 bl[10] br[10] wl[426] vdd gnd cell_6t
Xbit_r427_c10 bl[10] br[10] wl[427] vdd gnd cell_6t
Xbit_r428_c10 bl[10] br[10] wl[428] vdd gnd cell_6t
Xbit_r429_c10 bl[10] br[10] wl[429] vdd gnd cell_6t
Xbit_r430_c10 bl[10] br[10] wl[430] vdd gnd cell_6t
Xbit_r431_c10 bl[10] br[10] wl[431] vdd gnd cell_6t
Xbit_r432_c10 bl[10] br[10] wl[432] vdd gnd cell_6t
Xbit_r433_c10 bl[10] br[10] wl[433] vdd gnd cell_6t
Xbit_r434_c10 bl[10] br[10] wl[434] vdd gnd cell_6t
Xbit_r435_c10 bl[10] br[10] wl[435] vdd gnd cell_6t
Xbit_r436_c10 bl[10] br[10] wl[436] vdd gnd cell_6t
Xbit_r437_c10 bl[10] br[10] wl[437] vdd gnd cell_6t
Xbit_r438_c10 bl[10] br[10] wl[438] vdd gnd cell_6t
Xbit_r439_c10 bl[10] br[10] wl[439] vdd gnd cell_6t
Xbit_r440_c10 bl[10] br[10] wl[440] vdd gnd cell_6t
Xbit_r441_c10 bl[10] br[10] wl[441] vdd gnd cell_6t
Xbit_r442_c10 bl[10] br[10] wl[442] vdd gnd cell_6t
Xbit_r443_c10 bl[10] br[10] wl[443] vdd gnd cell_6t
Xbit_r444_c10 bl[10] br[10] wl[444] vdd gnd cell_6t
Xbit_r445_c10 bl[10] br[10] wl[445] vdd gnd cell_6t
Xbit_r446_c10 bl[10] br[10] wl[446] vdd gnd cell_6t
Xbit_r447_c10 bl[10] br[10] wl[447] vdd gnd cell_6t
Xbit_r448_c10 bl[10] br[10] wl[448] vdd gnd cell_6t
Xbit_r449_c10 bl[10] br[10] wl[449] vdd gnd cell_6t
Xbit_r450_c10 bl[10] br[10] wl[450] vdd gnd cell_6t
Xbit_r451_c10 bl[10] br[10] wl[451] vdd gnd cell_6t
Xbit_r452_c10 bl[10] br[10] wl[452] vdd gnd cell_6t
Xbit_r453_c10 bl[10] br[10] wl[453] vdd gnd cell_6t
Xbit_r454_c10 bl[10] br[10] wl[454] vdd gnd cell_6t
Xbit_r455_c10 bl[10] br[10] wl[455] vdd gnd cell_6t
Xbit_r456_c10 bl[10] br[10] wl[456] vdd gnd cell_6t
Xbit_r457_c10 bl[10] br[10] wl[457] vdd gnd cell_6t
Xbit_r458_c10 bl[10] br[10] wl[458] vdd gnd cell_6t
Xbit_r459_c10 bl[10] br[10] wl[459] vdd gnd cell_6t
Xbit_r460_c10 bl[10] br[10] wl[460] vdd gnd cell_6t
Xbit_r461_c10 bl[10] br[10] wl[461] vdd gnd cell_6t
Xbit_r462_c10 bl[10] br[10] wl[462] vdd gnd cell_6t
Xbit_r463_c10 bl[10] br[10] wl[463] vdd gnd cell_6t
Xbit_r464_c10 bl[10] br[10] wl[464] vdd gnd cell_6t
Xbit_r465_c10 bl[10] br[10] wl[465] vdd gnd cell_6t
Xbit_r466_c10 bl[10] br[10] wl[466] vdd gnd cell_6t
Xbit_r467_c10 bl[10] br[10] wl[467] vdd gnd cell_6t
Xbit_r468_c10 bl[10] br[10] wl[468] vdd gnd cell_6t
Xbit_r469_c10 bl[10] br[10] wl[469] vdd gnd cell_6t
Xbit_r470_c10 bl[10] br[10] wl[470] vdd gnd cell_6t
Xbit_r471_c10 bl[10] br[10] wl[471] vdd gnd cell_6t
Xbit_r472_c10 bl[10] br[10] wl[472] vdd gnd cell_6t
Xbit_r473_c10 bl[10] br[10] wl[473] vdd gnd cell_6t
Xbit_r474_c10 bl[10] br[10] wl[474] vdd gnd cell_6t
Xbit_r475_c10 bl[10] br[10] wl[475] vdd gnd cell_6t
Xbit_r476_c10 bl[10] br[10] wl[476] vdd gnd cell_6t
Xbit_r477_c10 bl[10] br[10] wl[477] vdd gnd cell_6t
Xbit_r478_c10 bl[10] br[10] wl[478] vdd gnd cell_6t
Xbit_r479_c10 bl[10] br[10] wl[479] vdd gnd cell_6t
Xbit_r480_c10 bl[10] br[10] wl[480] vdd gnd cell_6t
Xbit_r481_c10 bl[10] br[10] wl[481] vdd gnd cell_6t
Xbit_r482_c10 bl[10] br[10] wl[482] vdd gnd cell_6t
Xbit_r483_c10 bl[10] br[10] wl[483] vdd gnd cell_6t
Xbit_r484_c10 bl[10] br[10] wl[484] vdd gnd cell_6t
Xbit_r485_c10 bl[10] br[10] wl[485] vdd gnd cell_6t
Xbit_r486_c10 bl[10] br[10] wl[486] vdd gnd cell_6t
Xbit_r487_c10 bl[10] br[10] wl[487] vdd gnd cell_6t
Xbit_r488_c10 bl[10] br[10] wl[488] vdd gnd cell_6t
Xbit_r489_c10 bl[10] br[10] wl[489] vdd gnd cell_6t
Xbit_r490_c10 bl[10] br[10] wl[490] vdd gnd cell_6t
Xbit_r491_c10 bl[10] br[10] wl[491] vdd gnd cell_6t
Xbit_r492_c10 bl[10] br[10] wl[492] vdd gnd cell_6t
Xbit_r493_c10 bl[10] br[10] wl[493] vdd gnd cell_6t
Xbit_r494_c10 bl[10] br[10] wl[494] vdd gnd cell_6t
Xbit_r495_c10 bl[10] br[10] wl[495] vdd gnd cell_6t
Xbit_r496_c10 bl[10] br[10] wl[496] vdd gnd cell_6t
Xbit_r497_c10 bl[10] br[10] wl[497] vdd gnd cell_6t
Xbit_r498_c10 bl[10] br[10] wl[498] vdd gnd cell_6t
Xbit_r499_c10 bl[10] br[10] wl[499] vdd gnd cell_6t
Xbit_r500_c10 bl[10] br[10] wl[500] vdd gnd cell_6t
Xbit_r501_c10 bl[10] br[10] wl[501] vdd gnd cell_6t
Xbit_r502_c10 bl[10] br[10] wl[502] vdd gnd cell_6t
Xbit_r503_c10 bl[10] br[10] wl[503] vdd gnd cell_6t
Xbit_r504_c10 bl[10] br[10] wl[504] vdd gnd cell_6t
Xbit_r505_c10 bl[10] br[10] wl[505] vdd gnd cell_6t
Xbit_r506_c10 bl[10] br[10] wl[506] vdd gnd cell_6t
Xbit_r507_c10 bl[10] br[10] wl[507] vdd gnd cell_6t
Xbit_r508_c10 bl[10] br[10] wl[508] vdd gnd cell_6t
Xbit_r509_c10 bl[10] br[10] wl[509] vdd gnd cell_6t
Xbit_r510_c10 bl[10] br[10] wl[510] vdd gnd cell_6t
Xbit_r511_c10 bl[10] br[10] wl[511] vdd gnd cell_6t
Xbit_r0_c11 bl[11] br[11] wl[0] vdd gnd cell_6t
Xbit_r1_c11 bl[11] br[11] wl[1] vdd gnd cell_6t
Xbit_r2_c11 bl[11] br[11] wl[2] vdd gnd cell_6t
Xbit_r3_c11 bl[11] br[11] wl[3] vdd gnd cell_6t
Xbit_r4_c11 bl[11] br[11] wl[4] vdd gnd cell_6t
Xbit_r5_c11 bl[11] br[11] wl[5] vdd gnd cell_6t
Xbit_r6_c11 bl[11] br[11] wl[6] vdd gnd cell_6t
Xbit_r7_c11 bl[11] br[11] wl[7] vdd gnd cell_6t
Xbit_r8_c11 bl[11] br[11] wl[8] vdd gnd cell_6t
Xbit_r9_c11 bl[11] br[11] wl[9] vdd gnd cell_6t
Xbit_r10_c11 bl[11] br[11] wl[10] vdd gnd cell_6t
Xbit_r11_c11 bl[11] br[11] wl[11] vdd gnd cell_6t
Xbit_r12_c11 bl[11] br[11] wl[12] vdd gnd cell_6t
Xbit_r13_c11 bl[11] br[11] wl[13] vdd gnd cell_6t
Xbit_r14_c11 bl[11] br[11] wl[14] vdd gnd cell_6t
Xbit_r15_c11 bl[11] br[11] wl[15] vdd gnd cell_6t
Xbit_r16_c11 bl[11] br[11] wl[16] vdd gnd cell_6t
Xbit_r17_c11 bl[11] br[11] wl[17] vdd gnd cell_6t
Xbit_r18_c11 bl[11] br[11] wl[18] vdd gnd cell_6t
Xbit_r19_c11 bl[11] br[11] wl[19] vdd gnd cell_6t
Xbit_r20_c11 bl[11] br[11] wl[20] vdd gnd cell_6t
Xbit_r21_c11 bl[11] br[11] wl[21] vdd gnd cell_6t
Xbit_r22_c11 bl[11] br[11] wl[22] vdd gnd cell_6t
Xbit_r23_c11 bl[11] br[11] wl[23] vdd gnd cell_6t
Xbit_r24_c11 bl[11] br[11] wl[24] vdd gnd cell_6t
Xbit_r25_c11 bl[11] br[11] wl[25] vdd gnd cell_6t
Xbit_r26_c11 bl[11] br[11] wl[26] vdd gnd cell_6t
Xbit_r27_c11 bl[11] br[11] wl[27] vdd gnd cell_6t
Xbit_r28_c11 bl[11] br[11] wl[28] vdd gnd cell_6t
Xbit_r29_c11 bl[11] br[11] wl[29] vdd gnd cell_6t
Xbit_r30_c11 bl[11] br[11] wl[30] vdd gnd cell_6t
Xbit_r31_c11 bl[11] br[11] wl[31] vdd gnd cell_6t
Xbit_r32_c11 bl[11] br[11] wl[32] vdd gnd cell_6t
Xbit_r33_c11 bl[11] br[11] wl[33] vdd gnd cell_6t
Xbit_r34_c11 bl[11] br[11] wl[34] vdd gnd cell_6t
Xbit_r35_c11 bl[11] br[11] wl[35] vdd gnd cell_6t
Xbit_r36_c11 bl[11] br[11] wl[36] vdd gnd cell_6t
Xbit_r37_c11 bl[11] br[11] wl[37] vdd gnd cell_6t
Xbit_r38_c11 bl[11] br[11] wl[38] vdd gnd cell_6t
Xbit_r39_c11 bl[11] br[11] wl[39] vdd gnd cell_6t
Xbit_r40_c11 bl[11] br[11] wl[40] vdd gnd cell_6t
Xbit_r41_c11 bl[11] br[11] wl[41] vdd gnd cell_6t
Xbit_r42_c11 bl[11] br[11] wl[42] vdd gnd cell_6t
Xbit_r43_c11 bl[11] br[11] wl[43] vdd gnd cell_6t
Xbit_r44_c11 bl[11] br[11] wl[44] vdd gnd cell_6t
Xbit_r45_c11 bl[11] br[11] wl[45] vdd gnd cell_6t
Xbit_r46_c11 bl[11] br[11] wl[46] vdd gnd cell_6t
Xbit_r47_c11 bl[11] br[11] wl[47] vdd gnd cell_6t
Xbit_r48_c11 bl[11] br[11] wl[48] vdd gnd cell_6t
Xbit_r49_c11 bl[11] br[11] wl[49] vdd gnd cell_6t
Xbit_r50_c11 bl[11] br[11] wl[50] vdd gnd cell_6t
Xbit_r51_c11 bl[11] br[11] wl[51] vdd gnd cell_6t
Xbit_r52_c11 bl[11] br[11] wl[52] vdd gnd cell_6t
Xbit_r53_c11 bl[11] br[11] wl[53] vdd gnd cell_6t
Xbit_r54_c11 bl[11] br[11] wl[54] vdd gnd cell_6t
Xbit_r55_c11 bl[11] br[11] wl[55] vdd gnd cell_6t
Xbit_r56_c11 bl[11] br[11] wl[56] vdd gnd cell_6t
Xbit_r57_c11 bl[11] br[11] wl[57] vdd gnd cell_6t
Xbit_r58_c11 bl[11] br[11] wl[58] vdd gnd cell_6t
Xbit_r59_c11 bl[11] br[11] wl[59] vdd gnd cell_6t
Xbit_r60_c11 bl[11] br[11] wl[60] vdd gnd cell_6t
Xbit_r61_c11 bl[11] br[11] wl[61] vdd gnd cell_6t
Xbit_r62_c11 bl[11] br[11] wl[62] vdd gnd cell_6t
Xbit_r63_c11 bl[11] br[11] wl[63] vdd gnd cell_6t
Xbit_r64_c11 bl[11] br[11] wl[64] vdd gnd cell_6t
Xbit_r65_c11 bl[11] br[11] wl[65] vdd gnd cell_6t
Xbit_r66_c11 bl[11] br[11] wl[66] vdd gnd cell_6t
Xbit_r67_c11 bl[11] br[11] wl[67] vdd gnd cell_6t
Xbit_r68_c11 bl[11] br[11] wl[68] vdd gnd cell_6t
Xbit_r69_c11 bl[11] br[11] wl[69] vdd gnd cell_6t
Xbit_r70_c11 bl[11] br[11] wl[70] vdd gnd cell_6t
Xbit_r71_c11 bl[11] br[11] wl[71] vdd gnd cell_6t
Xbit_r72_c11 bl[11] br[11] wl[72] vdd gnd cell_6t
Xbit_r73_c11 bl[11] br[11] wl[73] vdd gnd cell_6t
Xbit_r74_c11 bl[11] br[11] wl[74] vdd gnd cell_6t
Xbit_r75_c11 bl[11] br[11] wl[75] vdd gnd cell_6t
Xbit_r76_c11 bl[11] br[11] wl[76] vdd gnd cell_6t
Xbit_r77_c11 bl[11] br[11] wl[77] vdd gnd cell_6t
Xbit_r78_c11 bl[11] br[11] wl[78] vdd gnd cell_6t
Xbit_r79_c11 bl[11] br[11] wl[79] vdd gnd cell_6t
Xbit_r80_c11 bl[11] br[11] wl[80] vdd gnd cell_6t
Xbit_r81_c11 bl[11] br[11] wl[81] vdd gnd cell_6t
Xbit_r82_c11 bl[11] br[11] wl[82] vdd gnd cell_6t
Xbit_r83_c11 bl[11] br[11] wl[83] vdd gnd cell_6t
Xbit_r84_c11 bl[11] br[11] wl[84] vdd gnd cell_6t
Xbit_r85_c11 bl[11] br[11] wl[85] vdd gnd cell_6t
Xbit_r86_c11 bl[11] br[11] wl[86] vdd gnd cell_6t
Xbit_r87_c11 bl[11] br[11] wl[87] vdd gnd cell_6t
Xbit_r88_c11 bl[11] br[11] wl[88] vdd gnd cell_6t
Xbit_r89_c11 bl[11] br[11] wl[89] vdd gnd cell_6t
Xbit_r90_c11 bl[11] br[11] wl[90] vdd gnd cell_6t
Xbit_r91_c11 bl[11] br[11] wl[91] vdd gnd cell_6t
Xbit_r92_c11 bl[11] br[11] wl[92] vdd gnd cell_6t
Xbit_r93_c11 bl[11] br[11] wl[93] vdd gnd cell_6t
Xbit_r94_c11 bl[11] br[11] wl[94] vdd gnd cell_6t
Xbit_r95_c11 bl[11] br[11] wl[95] vdd gnd cell_6t
Xbit_r96_c11 bl[11] br[11] wl[96] vdd gnd cell_6t
Xbit_r97_c11 bl[11] br[11] wl[97] vdd gnd cell_6t
Xbit_r98_c11 bl[11] br[11] wl[98] vdd gnd cell_6t
Xbit_r99_c11 bl[11] br[11] wl[99] vdd gnd cell_6t
Xbit_r100_c11 bl[11] br[11] wl[100] vdd gnd cell_6t
Xbit_r101_c11 bl[11] br[11] wl[101] vdd gnd cell_6t
Xbit_r102_c11 bl[11] br[11] wl[102] vdd gnd cell_6t
Xbit_r103_c11 bl[11] br[11] wl[103] vdd gnd cell_6t
Xbit_r104_c11 bl[11] br[11] wl[104] vdd gnd cell_6t
Xbit_r105_c11 bl[11] br[11] wl[105] vdd gnd cell_6t
Xbit_r106_c11 bl[11] br[11] wl[106] vdd gnd cell_6t
Xbit_r107_c11 bl[11] br[11] wl[107] vdd gnd cell_6t
Xbit_r108_c11 bl[11] br[11] wl[108] vdd gnd cell_6t
Xbit_r109_c11 bl[11] br[11] wl[109] vdd gnd cell_6t
Xbit_r110_c11 bl[11] br[11] wl[110] vdd gnd cell_6t
Xbit_r111_c11 bl[11] br[11] wl[111] vdd gnd cell_6t
Xbit_r112_c11 bl[11] br[11] wl[112] vdd gnd cell_6t
Xbit_r113_c11 bl[11] br[11] wl[113] vdd gnd cell_6t
Xbit_r114_c11 bl[11] br[11] wl[114] vdd gnd cell_6t
Xbit_r115_c11 bl[11] br[11] wl[115] vdd gnd cell_6t
Xbit_r116_c11 bl[11] br[11] wl[116] vdd gnd cell_6t
Xbit_r117_c11 bl[11] br[11] wl[117] vdd gnd cell_6t
Xbit_r118_c11 bl[11] br[11] wl[118] vdd gnd cell_6t
Xbit_r119_c11 bl[11] br[11] wl[119] vdd gnd cell_6t
Xbit_r120_c11 bl[11] br[11] wl[120] vdd gnd cell_6t
Xbit_r121_c11 bl[11] br[11] wl[121] vdd gnd cell_6t
Xbit_r122_c11 bl[11] br[11] wl[122] vdd gnd cell_6t
Xbit_r123_c11 bl[11] br[11] wl[123] vdd gnd cell_6t
Xbit_r124_c11 bl[11] br[11] wl[124] vdd gnd cell_6t
Xbit_r125_c11 bl[11] br[11] wl[125] vdd gnd cell_6t
Xbit_r126_c11 bl[11] br[11] wl[126] vdd gnd cell_6t
Xbit_r127_c11 bl[11] br[11] wl[127] vdd gnd cell_6t
Xbit_r128_c11 bl[11] br[11] wl[128] vdd gnd cell_6t
Xbit_r129_c11 bl[11] br[11] wl[129] vdd gnd cell_6t
Xbit_r130_c11 bl[11] br[11] wl[130] vdd gnd cell_6t
Xbit_r131_c11 bl[11] br[11] wl[131] vdd gnd cell_6t
Xbit_r132_c11 bl[11] br[11] wl[132] vdd gnd cell_6t
Xbit_r133_c11 bl[11] br[11] wl[133] vdd gnd cell_6t
Xbit_r134_c11 bl[11] br[11] wl[134] vdd gnd cell_6t
Xbit_r135_c11 bl[11] br[11] wl[135] vdd gnd cell_6t
Xbit_r136_c11 bl[11] br[11] wl[136] vdd gnd cell_6t
Xbit_r137_c11 bl[11] br[11] wl[137] vdd gnd cell_6t
Xbit_r138_c11 bl[11] br[11] wl[138] vdd gnd cell_6t
Xbit_r139_c11 bl[11] br[11] wl[139] vdd gnd cell_6t
Xbit_r140_c11 bl[11] br[11] wl[140] vdd gnd cell_6t
Xbit_r141_c11 bl[11] br[11] wl[141] vdd gnd cell_6t
Xbit_r142_c11 bl[11] br[11] wl[142] vdd gnd cell_6t
Xbit_r143_c11 bl[11] br[11] wl[143] vdd gnd cell_6t
Xbit_r144_c11 bl[11] br[11] wl[144] vdd gnd cell_6t
Xbit_r145_c11 bl[11] br[11] wl[145] vdd gnd cell_6t
Xbit_r146_c11 bl[11] br[11] wl[146] vdd gnd cell_6t
Xbit_r147_c11 bl[11] br[11] wl[147] vdd gnd cell_6t
Xbit_r148_c11 bl[11] br[11] wl[148] vdd gnd cell_6t
Xbit_r149_c11 bl[11] br[11] wl[149] vdd gnd cell_6t
Xbit_r150_c11 bl[11] br[11] wl[150] vdd gnd cell_6t
Xbit_r151_c11 bl[11] br[11] wl[151] vdd gnd cell_6t
Xbit_r152_c11 bl[11] br[11] wl[152] vdd gnd cell_6t
Xbit_r153_c11 bl[11] br[11] wl[153] vdd gnd cell_6t
Xbit_r154_c11 bl[11] br[11] wl[154] vdd gnd cell_6t
Xbit_r155_c11 bl[11] br[11] wl[155] vdd gnd cell_6t
Xbit_r156_c11 bl[11] br[11] wl[156] vdd gnd cell_6t
Xbit_r157_c11 bl[11] br[11] wl[157] vdd gnd cell_6t
Xbit_r158_c11 bl[11] br[11] wl[158] vdd gnd cell_6t
Xbit_r159_c11 bl[11] br[11] wl[159] vdd gnd cell_6t
Xbit_r160_c11 bl[11] br[11] wl[160] vdd gnd cell_6t
Xbit_r161_c11 bl[11] br[11] wl[161] vdd gnd cell_6t
Xbit_r162_c11 bl[11] br[11] wl[162] vdd gnd cell_6t
Xbit_r163_c11 bl[11] br[11] wl[163] vdd gnd cell_6t
Xbit_r164_c11 bl[11] br[11] wl[164] vdd gnd cell_6t
Xbit_r165_c11 bl[11] br[11] wl[165] vdd gnd cell_6t
Xbit_r166_c11 bl[11] br[11] wl[166] vdd gnd cell_6t
Xbit_r167_c11 bl[11] br[11] wl[167] vdd gnd cell_6t
Xbit_r168_c11 bl[11] br[11] wl[168] vdd gnd cell_6t
Xbit_r169_c11 bl[11] br[11] wl[169] vdd gnd cell_6t
Xbit_r170_c11 bl[11] br[11] wl[170] vdd gnd cell_6t
Xbit_r171_c11 bl[11] br[11] wl[171] vdd gnd cell_6t
Xbit_r172_c11 bl[11] br[11] wl[172] vdd gnd cell_6t
Xbit_r173_c11 bl[11] br[11] wl[173] vdd gnd cell_6t
Xbit_r174_c11 bl[11] br[11] wl[174] vdd gnd cell_6t
Xbit_r175_c11 bl[11] br[11] wl[175] vdd gnd cell_6t
Xbit_r176_c11 bl[11] br[11] wl[176] vdd gnd cell_6t
Xbit_r177_c11 bl[11] br[11] wl[177] vdd gnd cell_6t
Xbit_r178_c11 bl[11] br[11] wl[178] vdd gnd cell_6t
Xbit_r179_c11 bl[11] br[11] wl[179] vdd gnd cell_6t
Xbit_r180_c11 bl[11] br[11] wl[180] vdd gnd cell_6t
Xbit_r181_c11 bl[11] br[11] wl[181] vdd gnd cell_6t
Xbit_r182_c11 bl[11] br[11] wl[182] vdd gnd cell_6t
Xbit_r183_c11 bl[11] br[11] wl[183] vdd gnd cell_6t
Xbit_r184_c11 bl[11] br[11] wl[184] vdd gnd cell_6t
Xbit_r185_c11 bl[11] br[11] wl[185] vdd gnd cell_6t
Xbit_r186_c11 bl[11] br[11] wl[186] vdd gnd cell_6t
Xbit_r187_c11 bl[11] br[11] wl[187] vdd gnd cell_6t
Xbit_r188_c11 bl[11] br[11] wl[188] vdd gnd cell_6t
Xbit_r189_c11 bl[11] br[11] wl[189] vdd gnd cell_6t
Xbit_r190_c11 bl[11] br[11] wl[190] vdd gnd cell_6t
Xbit_r191_c11 bl[11] br[11] wl[191] vdd gnd cell_6t
Xbit_r192_c11 bl[11] br[11] wl[192] vdd gnd cell_6t
Xbit_r193_c11 bl[11] br[11] wl[193] vdd gnd cell_6t
Xbit_r194_c11 bl[11] br[11] wl[194] vdd gnd cell_6t
Xbit_r195_c11 bl[11] br[11] wl[195] vdd gnd cell_6t
Xbit_r196_c11 bl[11] br[11] wl[196] vdd gnd cell_6t
Xbit_r197_c11 bl[11] br[11] wl[197] vdd gnd cell_6t
Xbit_r198_c11 bl[11] br[11] wl[198] vdd gnd cell_6t
Xbit_r199_c11 bl[11] br[11] wl[199] vdd gnd cell_6t
Xbit_r200_c11 bl[11] br[11] wl[200] vdd gnd cell_6t
Xbit_r201_c11 bl[11] br[11] wl[201] vdd gnd cell_6t
Xbit_r202_c11 bl[11] br[11] wl[202] vdd gnd cell_6t
Xbit_r203_c11 bl[11] br[11] wl[203] vdd gnd cell_6t
Xbit_r204_c11 bl[11] br[11] wl[204] vdd gnd cell_6t
Xbit_r205_c11 bl[11] br[11] wl[205] vdd gnd cell_6t
Xbit_r206_c11 bl[11] br[11] wl[206] vdd gnd cell_6t
Xbit_r207_c11 bl[11] br[11] wl[207] vdd gnd cell_6t
Xbit_r208_c11 bl[11] br[11] wl[208] vdd gnd cell_6t
Xbit_r209_c11 bl[11] br[11] wl[209] vdd gnd cell_6t
Xbit_r210_c11 bl[11] br[11] wl[210] vdd gnd cell_6t
Xbit_r211_c11 bl[11] br[11] wl[211] vdd gnd cell_6t
Xbit_r212_c11 bl[11] br[11] wl[212] vdd gnd cell_6t
Xbit_r213_c11 bl[11] br[11] wl[213] vdd gnd cell_6t
Xbit_r214_c11 bl[11] br[11] wl[214] vdd gnd cell_6t
Xbit_r215_c11 bl[11] br[11] wl[215] vdd gnd cell_6t
Xbit_r216_c11 bl[11] br[11] wl[216] vdd gnd cell_6t
Xbit_r217_c11 bl[11] br[11] wl[217] vdd gnd cell_6t
Xbit_r218_c11 bl[11] br[11] wl[218] vdd gnd cell_6t
Xbit_r219_c11 bl[11] br[11] wl[219] vdd gnd cell_6t
Xbit_r220_c11 bl[11] br[11] wl[220] vdd gnd cell_6t
Xbit_r221_c11 bl[11] br[11] wl[221] vdd gnd cell_6t
Xbit_r222_c11 bl[11] br[11] wl[222] vdd gnd cell_6t
Xbit_r223_c11 bl[11] br[11] wl[223] vdd gnd cell_6t
Xbit_r224_c11 bl[11] br[11] wl[224] vdd gnd cell_6t
Xbit_r225_c11 bl[11] br[11] wl[225] vdd gnd cell_6t
Xbit_r226_c11 bl[11] br[11] wl[226] vdd gnd cell_6t
Xbit_r227_c11 bl[11] br[11] wl[227] vdd gnd cell_6t
Xbit_r228_c11 bl[11] br[11] wl[228] vdd gnd cell_6t
Xbit_r229_c11 bl[11] br[11] wl[229] vdd gnd cell_6t
Xbit_r230_c11 bl[11] br[11] wl[230] vdd gnd cell_6t
Xbit_r231_c11 bl[11] br[11] wl[231] vdd gnd cell_6t
Xbit_r232_c11 bl[11] br[11] wl[232] vdd gnd cell_6t
Xbit_r233_c11 bl[11] br[11] wl[233] vdd gnd cell_6t
Xbit_r234_c11 bl[11] br[11] wl[234] vdd gnd cell_6t
Xbit_r235_c11 bl[11] br[11] wl[235] vdd gnd cell_6t
Xbit_r236_c11 bl[11] br[11] wl[236] vdd gnd cell_6t
Xbit_r237_c11 bl[11] br[11] wl[237] vdd gnd cell_6t
Xbit_r238_c11 bl[11] br[11] wl[238] vdd gnd cell_6t
Xbit_r239_c11 bl[11] br[11] wl[239] vdd gnd cell_6t
Xbit_r240_c11 bl[11] br[11] wl[240] vdd gnd cell_6t
Xbit_r241_c11 bl[11] br[11] wl[241] vdd gnd cell_6t
Xbit_r242_c11 bl[11] br[11] wl[242] vdd gnd cell_6t
Xbit_r243_c11 bl[11] br[11] wl[243] vdd gnd cell_6t
Xbit_r244_c11 bl[11] br[11] wl[244] vdd gnd cell_6t
Xbit_r245_c11 bl[11] br[11] wl[245] vdd gnd cell_6t
Xbit_r246_c11 bl[11] br[11] wl[246] vdd gnd cell_6t
Xbit_r247_c11 bl[11] br[11] wl[247] vdd gnd cell_6t
Xbit_r248_c11 bl[11] br[11] wl[248] vdd gnd cell_6t
Xbit_r249_c11 bl[11] br[11] wl[249] vdd gnd cell_6t
Xbit_r250_c11 bl[11] br[11] wl[250] vdd gnd cell_6t
Xbit_r251_c11 bl[11] br[11] wl[251] vdd gnd cell_6t
Xbit_r252_c11 bl[11] br[11] wl[252] vdd gnd cell_6t
Xbit_r253_c11 bl[11] br[11] wl[253] vdd gnd cell_6t
Xbit_r254_c11 bl[11] br[11] wl[254] vdd gnd cell_6t
Xbit_r255_c11 bl[11] br[11] wl[255] vdd gnd cell_6t
Xbit_r256_c11 bl[11] br[11] wl[256] vdd gnd cell_6t
Xbit_r257_c11 bl[11] br[11] wl[257] vdd gnd cell_6t
Xbit_r258_c11 bl[11] br[11] wl[258] vdd gnd cell_6t
Xbit_r259_c11 bl[11] br[11] wl[259] vdd gnd cell_6t
Xbit_r260_c11 bl[11] br[11] wl[260] vdd gnd cell_6t
Xbit_r261_c11 bl[11] br[11] wl[261] vdd gnd cell_6t
Xbit_r262_c11 bl[11] br[11] wl[262] vdd gnd cell_6t
Xbit_r263_c11 bl[11] br[11] wl[263] vdd gnd cell_6t
Xbit_r264_c11 bl[11] br[11] wl[264] vdd gnd cell_6t
Xbit_r265_c11 bl[11] br[11] wl[265] vdd gnd cell_6t
Xbit_r266_c11 bl[11] br[11] wl[266] vdd gnd cell_6t
Xbit_r267_c11 bl[11] br[11] wl[267] vdd gnd cell_6t
Xbit_r268_c11 bl[11] br[11] wl[268] vdd gnd cell_6t
Xbit_r269_c11 bl[11] br[11] wl[269] vdd gnd cell_6t
Xbit_r270_c11 bl[11] br[11] wl[270] vdd gnd cell_6t
Xbit_r271_c11 bl[11] br[11] wl[271] vdd gnd cell_6t
Xbit_r272_c11 bl[11] br[11] wl[272] vdd gnd cell_6t
Xbit_r273_c11 bl[11] br[11] wl[273] vdd gnd cell_6t
Xbit_r274_c11 bl[11] br[11] wl[274] vdd gnd cell_6t
Xbit_r275_c11 bl[11] br[11] wl[275] vdd gnd cell_6t
Xbit_r276_c11 bl[11] br[11] wl[276] vdd gnd cell_6t
Xbit_r277_c11 bl[11] br[11] wl[277] vdd gnd cell_6t
Xbit_r278_c11 bl[11] br[11] wl[278] vdd gnd cell_6t
Xbit_r279_c11 bl[11] br[11] wl[279] vdd gnd cell_6t
Xbit_r280_c11 bl[11] br[11] wl[280] vdd gnd cell_6t
Xbit_r281_c11 bl[11] br[11] wl[281] vdd gnd cell_6t
Xbit_r282_c11 bl[11] br[11] wl[282] vdd gnd cell_6t
Xbit_r283_c11 bl[11] br[11] wl[283] vdd gnd cell_6t
Xbit_r284_c11 bl[11] br[11] wl[284] vdd gnd cell_6t
Xbit_r285_c11 bl[11] br[11] wl[285] vdd gnd cell_6t
Xbit_r286_c11 bl[11] br[11] wl[286] vdd gnd cell_6t
Xbit_r287_c11 bl[11] br[11] wl[287] vdd gnd cell_6t
Xbit_r288_c11 bl[11] br[11] wl[288] vdd gnd cell_6t
Xbit_r289_c11 bl[11] br[11] wl[289] vdd gnd cell_6t
Xbit_r290_c11 bl[11] br[11] wl[290] vdd gnd cell_6t
Xbit_r291_c11 bl[11] br[11] wl[291] vdd gnd cell_6t
Xbit_r292_c11 bl[11] br[11] wl[292] vdd gnd cell_6t
Xbit_r293_c11 bl[11] br[11] wl[293] vdd gnd cell_6t
Xbit_r294_c11 bl[11] br[11] wl[294] vdd gnd cell_6t
Xbit_r295_c11 bl[11] br[11] wl[295] vdd gnd cell_6t
Xbit_r296_c11 bl[11] br[11] wl[296] vdd gnd cell_6t
Xbit_r297_c11 bl[11] br[11] wl[297] vdd gnd cell_6t
Xbit_r298_c11 bl[11] br[11] wl[298] vdd gnd cell_6t
Xbit_r299_c11 bl[11] br[11] wl[299] vdd gnd cell_6t
Xbit_r300_c11 bl[11] br[11] wl[300] vdd gnd cell_6t
Xbit_r301_c11 bl[11] br[11] wl[301] vdd gnd cell_6t
Xbit_r302_c11 bl[11] br[11] wl[302] vdd gnd cell_6t
Xbit_r303_c11 bl[11] br[11] wl[303] vdd gnd cell_6t
Xbit_r304_c11 bl[11] br[11] wl[304] vdd gnd cell_6t
Xbit_r305_c11 bl[11] br[11] wl[305] vdd gnd cell_6t
Xbit_r306_c11 bl[11] br[11] wl[306] vdd gnd cell_6t
Xbit_r307_c11 bl[11] br[11] wl[307] vdd gnd cell_6t
Xbit_r308_c11 bl[11] br[11] wl[308] vdd gnd cell_6t
Xbit_r309_c11 bl[11] br[11] wl[309] vdd gnd cell_6t
Xbit_r310_c11 bl[11] br[11] wl[310] vdd gnd cell_6t
Xbit_r311_c11 bl[11] br[11] wl[311] vdd gnd cell_6t
Xbit_r312_c11 bl[11] br[11] wl[312] vdd gnd cell_6t
Xbit_r313_c11 bl[11] br[11] wl[313] vdd gnd cell_6t
Xbit_r314_c11 bl[11] br[11] wl[314] vdd gnd cell_6t
Xbit_r315_c11 bl[11] br[11] wl[315] vdd gnd cell_6t
Xbit_r316_c11 bl[11] br[11] wl[316] vdd gnd cell_6t
Xbit_r317_c11 bl[11] br[11] wl[317] vdd gnd cell_6t
Xbit_r318_c11 bl[11] br[11] wl[318] vdd gnd cell_6t
Xbit_r319_c11 bl[11] br[11] wl[319] vdd gnd cell_6t
Xbit_r320_c11 bl[11] br[11] wl[320] vdd gnd cell_6t
Xbit_r321_c11 bl[11] br[11] wl[321] vdd gnd cell_6t
Xbit_r322_c11 bl[11] br[11] wl[322] vdd gnd cell_6t
Xbit_r323_c11 bl[11] br[11] wl[323] vdd gnd cell_6t
Xbit_r324_c11 bl[11] br[11] wl[324] vdd gnd cell_6t
Xbit_r325_c11 bl[11] br[11] wl[325] vdd gnd cell_6t
Xbit_r326_c11 bl[11] br[11] wl[326] vdd gnd cell_6t
Xbit_r327_c11 bl[11] br[11] wl[327] vdd gnd cell_6t
Xbit_r328_c11 bl[11] br[11] wl[328] vdd gnd cell_6t
Xbit_r329_c11 bl[11] br[11] wl[329] vdd gnd cell_6t
Xbit_r330_c11 bl[11] br[11] wl[330] vdd gnd cell_6t
Xbit_r331_c11 bl[11] br[11] wl[331] vdd gnd cell_6t
Xbit_r332_c11 bl[11] br[11] wl[332] vdd gnd cell_6t
Xbit_r333_c11 bl[11] br[11] wl[333] vdd gnd cell_6t
Xbit_r334_c11 bl[11] br[11] wl[334] vdd gnd cell_6t
Xbit_r335_c11 bl[11] br[11] wl[335] vdd gnd cell_6t
Xbit_r336_c11 bl[11] br[11] wl[336] vdd gnd cell_6t
Xbit_r337_c11 bl[11] br[11] wl[337] vdd gnd cell_6t
Xbit_r338_c11 bl[11] br[11] wl[338] vdd gnd cell_6t
Xbit_r339_c11 bl[11] br[11] wl[339] vdd gnd cell_6t
Xbit_r340_c11 bl[11] br[11] wl[340] vdd gnd cell_6t
Xbit_r341_c11 bl[11] br[11] wl[341] vdd gnd cell_6t
Xbit_r342_c11 bl[11] br[11] wl[342] vdd gnd cell_6t
Xbit_r343_c11 bl[11] br[11] wl[343] vdd gnd cell_6t
Xbit_r344_c11 bl[11] br[11] wl[344] vdd gnd cell_6t
Xbit_r345_c11 bl[11] br[11] wl[345] vdd gnd cell_6t
Xbit_r346_c11 bl[11] br[11] wl[346] vdd gnd cell_6t
Xbit_r347_c11 bl[11] br[11] wl[347] vdd gnd cell_6t
Xbit_r348_c11 bl[11] br[11] wl[348] vdd gnd cell_6t
Xbit_r349_c11 bl[11] br[11] wl[349] vdd gnd cell_6t
Xbit_r350_c11 bl[11] br[11] wl[350] vdd gnd cell_6t
Xbit_r351_c11 bl[11] br[11] wl[351] vdd gnd cell_6t
Xbit_r352_c11 bl[11] br[11] wl[352] vdd gnd cell_6t
Xbit_r353_c11 bl[11] br[11] wl[353] vdd gnd cell_6t
Xbit_r354_c11 bl[11] br[11] wl[354] vdd gnd cell_6t
Xbit_r355_c11 bl[11] br[11] wl[355] vdd gnd cell_6t
Xbit_r356_c11 bl[11] br[11] wl[356] vdd gnd cell_6t
Xbit_r357_c11 bl[11] br[11] wl[357] vdd gnd cell_6t
Xbit_r358_c11 bl[11] br[11] wl[358] vdd gnd cell_6t
Xbit_r359_c11 bl[11] br[11] wl[359] vdd gnd cell_6t
Xbit_r360_c11 bl[11] br[11] wl[360] vdd gnd cell_6t
Xbit_r361_c11 bl[11] br[11] wl[361] vdd gnd cell_6t
Xbit_r362_c11 bl[11] br[11] wl[362] vdd gnd cell_6t
Xbit_r363_c11 bl[11] br[11] wl[363] vdd gnd cell_6t
Xbit_r364_c11 bl[11] br[11] wl[364] vdd gnd cell_6t
Xbit_r365_c11 bl[11] br[11] wl[365] vdd gnd cell_6t
Xbit_r366_c11 bl[11] br[11] wl[366] vdd gnd cell_6t
Xbit_r367_c11 bl[11] br[11] wl[367] vdd gnd cell_6t
Xbit_r368_c11 bl[11] br[11] wl[368] vdd gnd cell_6t
Xbit_r369_c11 bl[11] br[11] wl[369] vdd gnd cell_6t
Xbit_r370_c11 bl[11] br[11] wl[370] vdd gnd cell_6t
Xbit_r371_c11 bl[11] br[11] wl[371] vdd gnd cell_6t
Xbit_r372_c11 bl[11] br[11] wl[372] vdd gnd cell_6t
Xbit_r373_c11 bl[11] br[11] wl[373] vdd gnd cell_6t
Xbit_r374_c11 bl[11] br[11] wl[374] vdd gnd cell_6t
Xbit_r375_c11 bl[11] br[11] wl[375] vdd gnd cell_6t
Xbit_r376_c11 bl[11] br[11] wl[376] vdd gnd cell_6t
Xbit_r377_c11 bl[11] br[11] wl[377] vdd gnd cell_6t
Xbit_r378_c11 bl[11] br[11] wl[378] vdd gnd cell_6t
Xbit_r379_c11 bl[11] br[11] wl[379] vdd gnd cell_6t
Xbit_r380_c11 bl[11] br[11] wl[380] vdd gnd cell_6t
Xbit_r381_c11 bl[11] br[11] wl[381] vdd gnd cell_6t
Xbit_r382_c11 bl[11] br[11] wl[382] vdd gnd cell_6t
Xbit_r383_c11 bl[11] br[11] wl[383] vdd gnd cell_6t
Xbit_r384_c11 bl[11] br[11] wl[384] vdd gnd cell_6t
Xbit_r385_c11 bl[11] br[11] wl[385] vdd gnd cell_6t
Xbit_r386_c11 bl[11] br[11] wl[386] vdd gnd cell_6t
Xbit_r387_c11 bl[11] br[11] wl[387] vdd gnd cell_6t
Xbit_r388_c11 bl[11] br[11] wl[388] vdd gnd cell_6t
Xbit_r389_c11 bl[11] br[11] wl[389] vdd gnd cell_6t
Xbit_r390_c11 bl[11] br[11] wl[390] vdd gnd cell_6t
Xbit_r391_c11 bl[11] br[11] wl[391] vdd gnd cell_6t
Xbit_r392_c11 bl[11] br[11] wl[392] vdd gnd cell_6t
Xbit_r393_c11 bl[11] br[11] wl[393] vdd gnd cell_6t
Xbit_r394_c11 bl[11] br[11] wl[394] vdd gnd cell_6t
Xbit_r395_c11 bl[11] br[11] wl[395] vdd gnd cell_6t
Xbit_r396_c11 bl[11] br[11] wl[396] vdd gnd cell_6t
Xbit_r397_c11 bl[11] br[11] wl[397] vdd gnd cell_6t
Xbit_r398_c11 bl[11] br[11] wl[398] vdd gnd cell_6t
Xbit_r399_c11 bl[11] br[11] wl[399] vdd gnd cell_6t
Xbit_r400_c11 bl[11] br[11] wl[400] vdd gnd cell_6t
Xbit_r401_c11 bl[11] br[11] wl[401] vdd gnd cell_6t
Xbit_r402_c11 bl[11] br[11] wl[402] vdd gnd cell_6t
Xbit_r403_c11 bl[11] br[11] wl[403] vdd gnd cell_6t
Xbit_r404_c11 bl[11] br[11] wl[404] vdd gnd cell_6t
Xbit_r405_c11 bl[11] br[11] wl[405] vdd gnd cell_6t
Xbit_r406_c11 bl[11] br[11] wl[406] vdd gnd cell_6t
Xbit_r407_c11 bl[11] br[11] wl[407] vdd gnd cell_6t
Xbit_r408_c11 bl[11] br[11] wl[408] vdd gnd cell_6t
Xbit_r409_c11 bl[11] br[11] wl[409] vdd gnd cell_6t
Xbit_r410_c11 bl[11] br[11] wl[410] vdd gnd cell_6t
Xbit_r411_c11 bl[11] br[11] wl[411] vdd gnd cell_6t
Xbit_r412_c11 bl[11] br[11] wl[412] vdd gnd cell_6t
Xbit_r413_c11 bl[11] br[11] wl[413] vdd gnd cell_6t
Xbit_r414_c11 bl[11] br[11] wl[414] vdd gnd cell_6t
Xbit_r415_c11 bl[11] br[11] wl[415] vdd gnd cell_6t
Xbit_r416_c11 bl[11] br[11] wl[416] vdd gnd cell_6t
Xbit_r417_c11 bl[11] br[11] wl[417] vdd gnd cell_6t
Xbit_r418_c11 bl[11] br[11] wl[418] vdd gnd cell_6t
Xbit_r419_c11 bl[11] br[11] wl[419] vdd gnd cell_6t
Xbit_r420_c11 bl[11] br[11] wl[420] vdd gnd cell_6t
Xbit_r421_c11 bl[11] br[11] wl[421] vdd gnd cell_6t
Xbit_r422_c11 bl[11] br[11] wl[422] vdd gnd cell_6t
Xbit_r423_c11 bl[11] br[11] wl[423] vdd gnd cell_6t
Xbit_r424_c11 bl[11] br[11] wl[424] vdd gnd cell_6t
Xbit_r425_c11 bl[11] br[11] wl[425] vdd gnd cell_6t
Xbit_r426_c11 bl[11] br[11] wl[426] vdd gnd cell_6t
Xbit_r427_c11 bl[11] br[11] wl[427] vdd gnd cell_6t
Xbit_r428_c11 bl[11] br[11] wl[428] vdd gnd cell_6t
Xbit_r429_c11 bl[11] br[11] wl[429] vdd gnd cell_6t
Xbit_r430_c11 bl[11] br[11] wl[430] vdd gnd cell_6t
Xbit_r431_c11 bl[11] br[11] wl[431] vdd gnd cell_6t
Xbit_r432_c11 bl[11] br[11] wl[432] vdd gnd cell_6t
Xbit_r433_c11 bl[11] br[11] wl[433] vdd gnd cell_6t
Xbit_r434_c11 bl[11] br[11] wl[434] vdd gnd cell_6t
Xbit_r435_c11 bl[11] br[11] wl[435] vdd gnd cell_6t
Xbit_r436_c11 bl[11] br[11] wl[436] vdd gnd cell_6t
Xbit_r437_c11 bl[11] br[11] wl[437] vdd gnd cell_6t
Xbit_r438_c11 bl[11] br[11] wl[438] vdd gnd cell_6t
Xbit_r439_c11 bl[11] br[11] wl[439] vdd gnd cell_6t
Xbit_r440_c11 bl[11] br[11] wl[440] vdd gnd cell_6t
Xbit_r441_c11 bl[11] br[11] wl[441] vdd gnd cell_6t
Xbit_r442_c11 bl[11] br[11] wl[442] vdd gnd cell_6t
Xbit_r443_c11 bl[11] br[11] wl[443] vdd gnd cell_6t
Xbit_r444_c11 bl[11] br[11] wl[444] vdd gnd cell_6t
Xbit_r445_c11 bl[11] br[11] wl[445] vdd gnd cell_6t
Xbit_r446_c11 bl[11] br[11] wl[446] vdd gnd cell_6t
Xbit_r447_c11 bl[11] br[11] wl[447] vdd gnd cell_6t
Xbit_r448_c11 bl[11] br[11] wl[448] vdd gnd cell_6t
Xbit_r449_c11 bl[11] br[11] wl[449] vdd gnd cell_6t
Xbit_r450_c11 bl[11] br[11] wl[450] vdd gnd cell_6t
Xbit_r451_c11 bl[11] br[11] wl[451] vdd gnd cell_6t
Xbit_r452_c11 bl[11] br[11] wl[452] vdd gnd cell_6t
Xbit_r453_c11 bl[11] br[11] wl[453] vdd gnd cell_6t
Xbit_r454_c11 bl[11] br[11] wl[454] vdd gnd cell_6t
Xbit_r455_c11 bl[11] br[11] wl[455] vdd gnd cell_6t
Xbit_r456_c11 bl[11] br[11] wl[456] vdd gnd cell_6t
Xbit_r457_c11 bl[11] br[11] wl[457] vdd gnd cell_6t
Xbit_r458_c11 bl[11] br[11] wl[458] vdd gnd cell_6t
Xbit_r459_c11 bl[11] br[11] wl[459] vdd gnd cell_6t
Xbit_r460_c11 bl[11] br[11] wl[460] vdd gnd cell_6t
Xbit_r461_c11 bl[11] br[11] wl[461] vdd gnd cell_6t
Xbit_r462_c11 bl[11] br[11] wl[462] vdd gnd cell_6t
Xbit_r463_c11 bl[11] br[11] wl[463] vdd gnd cell_6t
Xbit_r464_c11 bl[11] br[11] wl[464] vdd gnd cell_6t
Xbit_r465_c11 bl[11] br[11] wl[465] vdd gnd cell_6t
Xbit_r466_c11 bl[11] br[11] wl[466] vdd gnd cell_6t
Xbit_r467_c11 bl[11] br[11] wl[467] vdd gnd cell_6t
Xbit_r468_c11 bl[11] br[11] wl[468] vdd gnd cell_6t
Xbit_r469_c11 bl[11] br[11] wl[469] vdd gnd cell_6t
Xbit_r470_c11 bl[11] br[11] wl[470] vdd gnd cell_6t
Xbit_r471_c11 bl[11] br[11] wl[471] vdd gnd cell_6t
Xbit_r472_c11 bl[11] br[11] wl[472] vdd gnd cell_6t
Xbit_r473_c11 bl[11] br[11] wl[473] vdd gnd cell_6t
Xbit_r474_c11 bl[11] br[11] wl[474] vdd gnd cell_6t
Xbit_r475_c11 bl[11] br[11] wl[475] vdd gnd cell_6t
Xbit_r476_c11 bl[11] br[11] wl[476] vdd gnd cell_6t
Xbit_r477_c11 bl[11] br[11] wl[477] vdd gnd cell_6t
Xbit_r478_c11 bl[11] br[11] wl[478] vdd gnd cell_6t
Xbit_r479_c11 bl[11] br[11] wl[479] vdd gnd cell_6t
Xbit_r480_c11 bl[11] br[11] wl[480] vdd gnd cell_6t
Xbit_r481_c11 bl[11] br[11] wl[481] vdd gnd cell_6t
Xbit_r482_c11 bl[11] br[11] wl[482] vdd gnd cell_6t
Xbit_r483_c11 bl[11] br[11] wl[483] vdd gnd cell_6t
Xbit_r484_c11 bl[11] br[11] wl[484] vdd gnd cell_6t
Xbit_r485_c11 bl[11] br[11] wl[485] vdd gnd cell_6t
Xbit_r486_c11 bl[11] br[11] wl[486] vdd gnd cell_6t
Xbit_r487_c11 bl[11] br[11] wl[487] vdd gnd cell_6t
Xbit_r488_c11 bl[11] br[11] wl[488] vdd gnd cell_6t
Xbit_r489_c11 bl[11] br[11] wl[489] vdd gnd cell_6t
Xbit_r490_c11 bl[11] br[11] wl[490] vdd gnd cell_6t
Xbit_r491_c11 bl[11] br[11] wl[491] vdd gnd cell_6t
Xbit_r492_c11 bl[11] br[11] wl[492] vdd gnd cell_6t
Xbit_r493_c11 bl[11] br[11] wl[493] vdd gnd cell_6t
Xbit_r494_c11 bl[11] br[11] wl[494] vdd gnd cell_6t
Xbit_r495_c11 bl[11] br[11] wl[495] vdd gnd cell_6t
Xbit_r496_c11 bl[11] br[11] wl[496] vdd gnd cell_6t
Xbit_r497_c11 bl[11] br[11] wl[497] vdd gnd cell_6t
Xbit_r498_c11 bl[11] br[11] wl[498] vdd gnd cell_6t
Xbit_r499_c11 bl[11] br[11] wl[499] vdd gnd cell_6t
Xbit_r500_c11 bl[11] br[11] wl[500] vdd gnd cell_6t
Xbit_r501_c11 bl[11] br[11] wl[501] vdd gnd cell_6t
Xbit_r502_c11 bl[11] br[11] wl[502] vdd gnd cell_6t
Xbit_r503_c11 bl[11] br[11] wl[503] vdd gnd cell_6t
Xbit_r504_c11 bl[11] br[11] wl[504] vdd gnd cell_6t
Xbit_r505_c11 bl[11] br[11] wl[505] vdd gnd cell_6t
Xbit_r506_c11 bl[11] br[11] wl[506] vdd gnd cell_6t
Xbit_r507_c11 bl[11] br[11] wl[507] vdd gnd cell_6t
Xbit_r508_c11 bl[11] br[11] wl[508] vdd gnd cell_6t
Xbit_r509_c11 bl[11] br[11] wl[509] vdd gnd cell_6t
Xbit_r510_c11 bl[11] br[11] wl[510] vdd gnd cell_6t
Xbit_r511_c11 bl[11] br[11] wl[511] vdd gnd cell_6t
Xbit_r0_c12 bl[12] br[12] wl[0] vdd gnd cell_6t
Xbit_r1_c12 bl[12] br[12] wl[1] vdd gnd cell_6t
Xbit_r2_c12 bl[12] br[12] wl[2] vdd gnd cell_6t
Xbit_r3_c12 bl[12] br[12] wl[3] vdd gnd cell_6t
Xbit_r4_c12 bl[12] br[12] wl[4] vdd gnd cell_6t
Xbit_r5_c12 bl[12] br[12] wl[5] vdd gnd cell_6t
Xbit_r6_c12 bl[12] br[12] wl[6] vdd gnd cell_6t
Xbit_r7_c12 bl[12] br[12] wl[7] vdd gnd cell_6t
Xbit_r8_c12 bl[12] br[12] wl[8] vdd gnd cell_6t
Xbit_r9_c12 bl[12] br[12] wl[9] vdd gnd cell_6t
Xbit_r10_c12 bl[12] br[12] wl[10] vdd gnd cell_6t
Xbit_r11_c12 bl[12] br[12] wl[11] vdd gnd cell_6t
Xbit_r12_c12 bl[12] br[12] wl[12] vdd gnd cell_6t
Xbit_r13_c12 bl[12] br[12] wl[13] vdd gnd cell_6t
Xbit_r14_c12 bl[12] br[12] wl[14] vdd gnd cell_6t
Xbit_r15_c12 bl[12] br[12] wl[15] vdd gnd cell_6t
Xbit_r16_c12 bl[12] br[12] wl[16] vdd gnd cell_6t
Xbit_r17_c12 bl[12] br[12] wl[17] vdd gnd cell_6t
Xbit_r18_c12 bl[12] br[12] wl[18] vdd gnd cell_6t
Xbit_r19_c12 bl[12] br[12] wl[19] vdd gnd cell_6t
Xbit_r20_c12 bl[12] br[12] wl[20] vdd gnd cell_6t
Xbit_r21_c12 bl[12] br[12] wl[21] vdd gnd cell_6t
Xbit_r22_c12 bl[12] br[12] wl[22] vdd gnd cell_6t
Xbit_r23_c12 bl[12] br[12] wl[23] vdd gnd cell_6t
Xbit_r24_c12 bl[12] br[12] wl[24] vdd gnd cell_6t
Xbit_r25_c12 bl[12] br[12] wl[25] vdd gnd cell_6t
Xbit_r26_c12 bl[12] br[12] wl[26] vdd gnd cell_6t
Xbit_r27_c12 bl[12] br[12] wl[27] vdd gnd cell_6t
Xbit_r28_c12 bl[12] br[12] wl[28] vdd gnd cell_6t
Xbit_r29_c12 bl[12] br[12] wl[29] vdd gnd cell_6t
Xbit_r30_c12 bl[12] br[12] wl[30] vdd gnd cell_6t
Xbit_r31_c12 bl[12] br[12] wl[31] vdd gnd cell_6t
Xbit_r32_c12 bl[12] br[12] wl[32] vdd gnd cell_6t
Xbit_r33_c12 bl[12] br[12] wl[33] vdd gnd cell_6t
Xbit_r34_c12 bl[12] br[12] wl[34] vdd gnd cell_6t
Xbit_r35_c12 bl[12] br[12] wl[35] vdd gnd cell_6t
Xbit_r36_c12 bl[12] br[12] wl[36] vdd gnd cell_6t
Xbit_r37_c12 bl[12] br[12] wl[37] vdd gnd cell_6t
Xbit_r38_c12 bl[12] br[12] wl[38] vdd gnd cell_6t
Xbit_r39_c12 bl[12] br[12] wl[39] vdd gnd cell_6t
Xbit_r40_c12 bl[12] br[12] wl[40] vdd gnd cell_6t
Xbit_r41_c12 bl[12] br[12] wl[41] vdd gnd cell_6t
Xbit_r42_c12 bl[12] br[12] wl[42] vdd gnd cell_6t
Xbit_r43_c12 bl[12] br[12] wl[43] vdd gnd cell_6t
Xbit_r44_c12 bl[12] br[12] wl[44] vdd gnd cell_6t
Xbit_r45_c12 bl[12] br[12] wl[45] vdd gnd cell_6t
Xbit_r46_c12 bl[12] br[12] wl[46] vdd gnd cell_6t
Xbit_r47_c12 bl[12] br[12] wl[47] vdd gnd cell_6t
Xbit_r48_c12 bl[12] br[12] wl[48] vdd gnd cell_6t
Xbit_r49_c12 bl[12] br[12] wl[49] vdd gnd cell_6t
Xbit_r50_c12 bl[12] br[12] wl[50] vdd gnd cell_6t
Xbit_r51_c12 bl[12] br[12] wl[51] vdd gnd cell_6t
Xbit_r52_c12 bl[12] br[12] wl[52] vdd gnd cell_6t
Xbit_r53_c12 bl[12] br[12] wl[53] vdd gnd cell_6t
Xbit_r54_c12 bl[12] br[12] wl[54] vdd gnd cell_6t
Xbit_r55_c12 bl[12] br[12] wl[55] vdd gnd cell_6t
Xbit_r56_c12 bl[12] br[12] wl[56] vdd gnd cell_6t
Xbit_r57_c12 bl[12] br[12] wl[57] vdd gnd cell_6t
Xbit_r58_c12 bl[12] br[12] wl[58] vdd gnd cell_6t
Xbit_r59_c12 bl[12] br[12] wl[59] vdd gnd cell_6t
Xbit_r60_c12 bl[12] br[12] wl[60] vdd gnd cell_6t
Xbit_r61_c12 bl[12] br[12] wl[61] vdd gnd cell_6t
Xbit_r62_c12 bl[12] br[12] wl[62] vdd gnd cell_6t
Xbit_r63_c12 bl[12] br[12] wl[63] vdd gnd cell_6t
Xbit_r64_c12 bl[12] br[12] wl[64] vdd gnd cell_6t
Xbit_r65_c12 bl[12] br[12] wl[65] vdd gnd cell_6t
Xbit_r66_c12 bl[12] br[12] wl[66] vdd gnd cell_6t
Xbit_r67_c12 bl[12] br[12] wl[67] vdd gnd cell_6t
Xbit_r68_c12 bl[12] br[12] wl[68] vdd gnd cell_6t
Xbit_r69_c12 bl[12] br[12] wl[69] vdd gnd cell_6t
Xbit_r70_c12 bl[12] br[12] wl[70] vdd gnd cell_6t
Xbit_r71_c12 bl[12] br[12] wl[71] vdd gnd cell_6t
Xbit_r72_c12 bl[12] br[12] wl[72] vdd gnd cell_6t
Xbit_r73_c12 bl[12] br[12] wl[73] vdd gnd cell_6t
Xbit_r74_c12 bl[12] br[12] wl[74] vdd gnd cell_6t
Xbit_r75_c12 bl[12] br[12] wl[75] vdd gnd cell_6t
Xbit_r76_c12 bl[12] br[12] wl[76] vdd gnd cell_6t
Xbit_r77_c12 bl[12] br[12] wl[77] vdd gnd cell_6t
Xbit_r78_c12 bl[12] br[12] wl[78] vdd gnd cell_6t
Xbit_r79_c12 bl[12] br[12] wl[79] vdd gnd cell_6t
Xbit_r80_c12 bl[12] br[12] wl[80] vdd gnd cell_6t
Xbit_r81_c12 bl[12] br[12] wl[81] vdd gnd cell_6t
Xbit_r82_c12 bl[12] br[12] wl[82] vdd gnd cell_6t
Xbit_r83_c12 bl[12] br[12] wl[83] vdd gnd cell_6t
Xbit_r84_c12 bl[12] br[12] wl[84] vdd gnd cell_6t
Xbit_r85_c12 bl[12] br[12] wl[85] vdd gnd cell_6t
Xbit_r86_c12 bl[12] br[12] wl[86] vdd gnd cell_6t
Xbit_r87_c12 bl[12] br[12] wl[87] vdd gnd cell_6t
Xbit_r88_c12 bl[12] br[12] wl[88] vdd gnd cell_6t
Xbit_r89_c12 bl[12] br[12] wl[89] vdd gnd cell_6t
Xbit_r90_c12 bl[12] br[12] wl[90] vdd gnd cell_6t
Xbit_r91_c12 bl[12] br[12] wl[91] vdd gnd cell_6t
Xbit_r92_c12 bl[12] br[12] wl[92] vdd gnd cell_6t
Xbit_r93_c12 bl[12] br[12] wl[93] vdd gnd cell_6t
Xbit_r94_c12 bl[12] br[12] wl[94] vdd gnd cell_6t
Xbit_r95_c12 bl[12] br[12] wl[95] vdd gnd cell_6t
Xbit_r96_c12 bl[12] br[12] wl[96] vdd gnd cell_6t
Xbit_r97_c12 bl[12] br[12] wl[97] vdd gnd cell_6t
Xbit_r98_c12 bl[12] br[12] wl[98] vdd gnd cell_6t
Xbit_r99_c12 bl[12] br[12] wl[99] vdd gnd cell_6t
Xbit_r100_c12 bl[12] br[12] wl[100] vdd gnd cell_6t
Xbit_r101_c12 bl[12] br[12] wl[101] vdd gnd cell_6t
Xbit_r102_c12 bl[12] br[12] wl[102] vdd gnd cell_6t
Xbit_r103_c12 bl[12] br[12] wl[103] vdd gnd cell_6t
Xbit_r104_c12 bl[12] br[12] wl[104] vdd gnd cell_6t
Xbit_r105_c12 bl[12] br[12] wl[105] vdd gnd cell_6t
Xbit_r106_c12 bl[12] br[12] wl[106] vdd gnd cell_6t
Xbit_r107_c12 bl[12] br[12] wl[107] vdd gnd cell_6t
Xbit_r108_c12 bl[12] br[12] wl[108] vdd gnd cell_6t
Xbit_r109_c12 bl[12] br[12] wl[109] vdd gnd cell_6t
Xbit_r110_c12 bl[12] br[12] wl[110] vdd gnd cell_6t
Xbit_r111_c12 bl[12] br[12] wl[111] vdd gnd cell_6t
Xbit_r112_c12 bl[12] br[12] wl[112] vdd gnd cell_6t
Xbit_r113_c12 bl[12] br[12] wl[113] vdd gnd cell_6t
Xbit_r114_c12 bl[12] br[12] wl[114] vdd gnd cell_6t
Xbit_r115_c12 bl[12] br[12] wl[115] vdd gnd cell_6t
Xbit_r116_c12 bl[12] br[12] wl[116] vdd gnd cell_6t
Xbit_r117_c12 bl[12] br[12] wl[117] vdd gnd cell_6t
Xbit_r118_c12 bl[12] br[12] wl[118] vdd gnd cell_6t
Xbit_r119_c12 bl[12] br[12] wl[119] vdd gnd cell_6t
Xbit_r120_c12 bl[12] br[12] wl[120] vdd gnd cell_6t
Xbit_r121_c12 bl[12] br[12] wl[121] vdd gnd cell_6t
Xbit_r122_c12 bl[12] br[12] wl[122] vdd gnd cell_6t
Xbit_r123_c12 bl[12] br[12] wl[123] vdd gnd cell_6t
Xbit_r124_c12 bl[12] br[12] wl[124] vdd gnd cell_6t
Xbit_r125_c12 bl[12] br[12] wl[125] vdd gnd cell_6t
Xbit_r126_c12 bl[12] br[12] wl[126] vdd gnd cell_6t
Xbit_r127_c12 bl[12] br[12] wl[127] vdd gnd cell_6t
Xbit_r128_c12 bl[12] br[12] wl[128] vdd gnd cell_6t
Xbit_r129_c12 bl[12] br[12] wl[129] vdd gnd cell_6t
Xbit_r130_c12 bl[12] br[12] wl[130] vdd gnd cell_6t
Xbit_r131_c12 bl[12] br[12] wl[131] vdd gnd cell_6t
Xbit_r132_c12 bl[12] br[12] wl[132] vdd gnd cell_6t
Xbit_r133_c12 bl[12] br[12] wl[133] vdd gnd cell_6t
Xbit_r134_c12 bl[12] br[12] wl[134] vdd gnd cell_6t
Xbit_r135_c12 bl[12] br[12] wl[135] vdd gnd cell_6t
Xbit_r136_c12 bl[12] br[12] wl[136] vdd gnd cell_6t
Xbit_r137_c12 bl[12] br[12] wl[137] vdd gnd cell_6t
Xbit_r138_c12 bl[12] br[12] wl[138] vdd gnd cell_6t
Xbit_r139_c12 bl[12] br[12] wl[139] vdd gnd cell_6t
Xbit_r140_c12 bl[12] br[12] wl[140] vdd gnd cell_6t
Xbit_r141_c12 bl[12] br[12] wl[141] vdd gnd cell_6t
Xbit_r142_c12 bl[12] br[12] wl[142] vdd gnd cell_6t
Xbit_r143_c12 bl[12] br[12] wl[143] vdd gnd cell_6t
Xbit_r144_c12 bl[12] br[12] wl[144] vdd gnd cell_6t
Xbit_r145_c12 bl[12] br[12] wl[145] vdd gnd cell_6t
Xbit_r146_c12 bl[12] br[12] wl[146] vdd gnd cell_6t
Xbit_r147_c12 bl[12] br[12] wl[147] vdd gnd cell_6t
Xbit_r148_c12 bl[12] br[12] wl[148] vdd gnd cell_6t
Xbit_r149_c12 bl[12] br[12] wl[149] vdd gnd cell_6t
Xbit_r150_c12 bl[12] br[12] wl[150] vdd gnd cell_6t
Xbit_r151_c12 bl[12] br[12] wl[151] vdd gnd cell_6t
Xbit_r152_c12 bl[12] br[12] wl[152] vdd gnd cell_6t
Xbit_r153_c12 bl[12] br[12] wl[153] vdd gnd cell_6t
Xbit_r154_c12 bl[12] br[12] wl[154] vdd gnd cell_6t
Xbit_r155_c12 bl[12] br[12] wl[155] vdd gnd cell_6t
Xbit_r156_c12 bl[12] br[12] wl[156] vdd gnd cell_6t
Xbit_r157_c12 bl[12] br[12] wl[157] vdd gnd cell_6t
Xbit_r158_c12 bl[12] br[12] wl[158] vdd gnd cell_6t
Xbit_r159_c12 bl[12] br[12] wl[159] vdd gnd cell_6t
Xbit_r160_c12 bl[12] br[12] wl[160] vdd gnd cell_6t
Xbit_r161_c12 bl[12] br[12] wl[161] vdd gnd cell_6t
Xbit_r162_c12 bl[12] br[12] wl[162] vdd gnd cell_6t
Xbit_r163_c12 bl[12] br[12] wl[163] vdd gnd cell_6t
Xbit_r164_c12 bl[12] br[12] wl[164] vdd gnd cell_6t
Xbit_r165_c12 bl[12] br[12] wl[165] vdd gnd cell_6t
Xbit_r166_c12 bl[12] br[12] wl[166] vdd gnd cell_6t
Xbit_r167_c12 bl[12] br[12] wl[167] vdd gnd cell_6t
Xbit_r168_c12 bl[12] br[12] wl[168] vdd gnd cell_6t
Xbit_r169_c12 bl[12] br[12] wl[169] vdd gnd cell_6t
Xbit_r170_c12 bl[12] br[12] wl[170] vdd gnd cell_6t
Xbit_r171_c12 bl[12] br[12] wl[171] vdd gnd cell_6t
Xbit_r172_c12 bl[12] br[12] wl[172] vdd gnd cell_6t
Xbit_r173_c12 bl[12] br[12] wl[173] vdd gnd cell_6t
Xbit_r174_c12 bl[12] br[12] wl[174] vdd gnd cell_6t
Xbit_r175_c12 bl[12] br[12] wl[175] vdd gnd cell_6t
Xbit_r176_c12 bl[12] br[12] wl[176] vdd gnd cell_6t
Xbit_r177_c12 bl[12] br[12] wl[177] vdd gnd cell_6t
Xbit_r178_c12 bl[12] br[12] wl[178] vdd gnd cell_6t
Xbit_r179_c12 bl[12] br[12] wl[179] vdd gnd cell_6t
Xbit_r180_c12 bl[12] br[12] wl[180] vdd gnd cell_6t
Xbit_r181_c12 bl[12] br[12] wl[181] vdd gnd cell_6t
Xbit_r182_c12 bl[12] br[12] wl[182] vdd gnd cell_6t
Xbit_r183_c12 bl[12] br[12] wl[183] vdd gnd cell_6t
Xbit_r184_c12 bl[12] br[12] wl[184] vdd gnd cell_6t
Xbit_r185_c12 bl[12] br[12] wl[185] vdd gnd cell_6t
Xbit_r186_c12 bl[12] br[12] wl[186] vdd gnd cell_6t
Xbit_r187_c12 bl[12] br[12] wl[187] vdd gnd cell_6t
Xbit_r188_c12 bl[12] br[12] wl[188] vdd gnd cell_6t
Xbit_r189_c12 bl[12] br[12] wl[189] vdd gnd cell_6t
Xbit_r190_c12 bl[12] br[12] wl[190] vdd gnd cell_6t
Xbit_r191_c12 bl[12] br[12] wl[191] vdd gnd cell_6t
Xbit_r192_c12 bl[12] br[12] wl[192] vdd gnd cell_6t
Xbit_r193_c12 bl[12] br[12] wl[193] vdd gnd cell_6t
Xbit_r194_c12 bl[12] br[12] wl[194] vdd gnd cell_6t
Xbit_r195_c12 bl[12] br[12] wl[195] vdd gnd cell_6t
Xbit_r196_c12 bl[12] br[12] wl[196] vdd gnd cell_6t
Xbit_r197_c12 bl[12] br[12] wl[197] vdd gnd cell_6t
Xbit_r198_c12 bl[12] br[12] wl[198] vdd gnd cell_6t
Xbit_r199_c12 bl[12] br[12] wl[199] vdd gnd cell_6t
Xbit_r200_c12 bl[12] br[12] wl[200] vdd gnd cell_6t
Xbit_r201_c12 bl[12] br[12] wl[201] vdd gnd cell_6t
Xbit_r202_c12 bl[12] br[12] wl[202] vdd gnd cell_6t
Xbit_r203_c12 bl[12] br[12] wl[203] vdd gnd cell_6t
Xbit_r204_c12 bl[12] br[12] wl[204] vdd gnd cell_6t
Xbit_r205_c12 bl[12] br[12] wl[205] vdd gnd cell_6t
Xbit_r206_c12 bl[12] br[12] wl[206] vdd gnd cell_6t
Xbit_r207_c12 bl[12] br[12] wl[207] vdd gnd cell_6t
Xbit_r208_c12 bl[12] br[12] wl[208] vdd gnd cell_6t
Xbit_r209_c12 bl[12] br[12] wl[209] vdd gnd cell_6t
Xbit_r210_c12 bl[12] br[12] wl[210] vdd gnd cell_6t
Xbit_r211_c12 bl[12] br[12] wl[211] vdd gnd cell_6t
Xbit_r212_c12 bl[12] br[12] wl[212] vdd gnd cell_6t
Xbit_r213_c12 bl[12] br[12] wl[213] vdd gnd cell_6t
Xbit_r214_c12 bl[12] br[12] wl[214] vdd gnd cell_6t
Xbit_r215_c12 bl[12] br[12] wl[215] vdd gnd cell_6t
Xbit_r216_c12 bl[12] br[12] wl[216] vdd gnd cell_6t
Xbit_r217_c12 bl[12] br[12] wl[217] vdd gnd cell_6t
Xbit_r218_c12 bl[12] br[12] wl[218] vdd gnd cell_6t
Xbit_r219_c12 bl[12] br[12] wl[219] vdd gnd cell_6t
Xbit_r220_c12 bl[12] br[12] wl[220] vdd gnd cell_6t
Xbit_r221_c12 bl[12] br[12] wl[221] vdd gnd cell_6t
Xbit_r222_c12 bl[12] br[12] wl[222] vdd gnd cell_6t
Xbit_r223_c12 bl[12] br[12] wl[223] vdd gnd cell_6t
Xbit_r224_c12 bl[12] br[12] wl[224] vdd gnd cell_6t
Xbit_r225_c12 bl[12] br[12] wl[225] vdd gnd cell_6t
Xbit_r226_c12 bl[12] br[12] wl[226] vdd gnd cell_6t
Xbit_r227_c12 bl[12] br[12] wl[227] vdd gnd cell_6t
Xbit_r228_c12 bl[12] br[12] wl[228] vdd gnd cell_6t
Xbit_r229_c12 bl[12] br[12] wl[229] vdd gnd cell_6t
Xbit_r230_c12 bl[12] br[12] wl[230] vdd gnd cell_6t
Xbit_r231_c12 bl[12] br[12] wl[231] vdd gnd cell_6t
Xbit_r232_c12 bl[12] br[12] wl[232] vdd gnd cell_6t
Xbit_r233_c12 bl[12] br[12] wl[233] vdd gnd cell_6t
Xbit_r234_c12 bl[12] br[12] wl[234] vdd gnd cell_6t
Xbit_r235_c12 bl[12] br[12] wl[235] vdd gnd cell_6t
Xbit_r236_c12 bl[12] br[12] wl[236] vdd gnd cell_6t
Xbit_r237_c12 bl[12] br[12] wl[237] vdd gnd cell_6t
Xbit_r238_c12 bl[12] br[12] wl[238] vdd gnd cell_6t
Xbit_r239_c12 bl[12] br[12] wl[239] vdd gnd cell_6t
Xbit_r240_c12 bl[12] br[12] wl[240] vdd gnd cell_6t
Xbit_r241_c12 bl[12] br[12] wl[241] vdd gnd cell_6t
Xbit_r242_c12 bl[12] br[12] wl[242] vdd gnd cell_6t
Xbit_r243_c12 bl[12] br[12] wl[243] vdd gnd cell_6t
Xbit_r244_c12 bl[12] br[12] wl[244] vdd gnd cell_6t
Xbit_r245_c12 bl[12] br[12] wl[245] vdd gnd cell_6t
Xbit_r246_c12 bl[12] br[12] wl[246] vdd gnd cell_6t
Xbit_r247_c12 bl[12] br[12] wl[247] vdd gnd cell_6t
Xbit_r248_c12 bl[12] br[12] wl[248] vdd gnd cell_6t
Xbit_r249_c12 bl[12] br[12] wl[249] vdd gnd cell_6t
Xbit_r250_c12 bl[12] br[12] wl[250] vdd gnd cell_6t
Xbit_r251_c12 bl[12] br[12] wl[251] vdd gnd cell_6t
Xbit_r252_c12 bl[12] br[12] wl[252] vdd gnd cell_6t
Xbit_r253_c12 bl[12] br[12] wl[253] vdd gnd cell_6t
Xbit_r254_c12 bl[12] br[12] wl[254] vdd gnd cell_6t
Xbit_r255_c12 bl[12] br[12] wl[255] vdd gnd cell_6t
Xbit_r256_c12 bl[12] br[12] wl[256] vdd gnd cell_6t
Xbit_r257_c12 bl[12] br[12] wl[257] vdd gnd cell_6t
Xbit_r258_c12 bl[12] br[12] wl[258] vdd gnd cell_6t
Xbit_r259_c12 bl[12] br[12] wl[259] vdd gnd cell_6t
Xbit_r260_c12 bl[12] br[12] wl[260] vdd gnd cell_6t
Xbit_r261_c12 bl[12] br[12] wl[261] vdd gnd cell_6t
Xbit_r262_c12 bl[12] br[12] wl[262] vdd gnd cell_6t
Xbit_r263_c12 bl[12] br[12] wl[263] vdd gnd cell_6t
Xbit_r264_c12 bl[12] br[12] wl[264] vdd gnd cell_6t
Xbit_r265_c12 bl[12] br[12] wl[265] vdd gnd cell_6t
Xbit_r266_c12 bl[12] br[12] wl[266] vdd gnd cell_6t
Xbit_r267_c12 bl[12] br[12] wl[267] vdd gnd cell_6t
Xbit_r268_c12 bl[12] br[12] wl[268] vdd gnd cell_6t
Xbit_r269_c12 bl[12] br[12] wl[269] vdd gnd cell_6t
Xbit_r270_c12 bl[12] br[12] wl[270] vdd gnd cell_6t
Xbit_r271_c12 bl[12] br[12] wl[271] vdd gnd cell_6t
Xbit_r272_c12 bl[12] br[12] wl[272] vdd gnd cell_6t
Xbit_r273_c12 bl[12] br[12] wl[273] vdd gnd cell_6t
Xbit_r274_c12 bl[12] br[12] wl[274] vdd gnd cell_6t
Xbit_r275_c12 bl[12] br[12] wl[275] vdd gnd cell_6t
Xbit_r276_c12 bl[12] br[12] wl[276] vdd gnd cell_6t
Xbit_r277_c12 bl[12] br[12] wl[277] vdd gnd cell_6t
Xbit_r278_c12 bl[12] br[12] wl[278] vdd gnd cell_6t
Xbit_r279_c12 bl[12] br[12] wl[279] vdd gnd cell_6t
Xbit_r280_c12 bl[12] br[12] wl[280] vdd gnd cell_6t
Xbit_r281_c12 bl[12] br[12] wl[281] vdd gnd cell_6t
Xbit_r282_c12 bl[12] br[12] wl[282] vdd gnd cell_6t
Xbit_r283_c12 bl[12] br[12] wl[283] vdd gnd cell_6t
Xbit_r284_c12 bl[12] br[12] wl[284] vdd gnd cell_6t
Xbit_r285_c12 bl[12] br[12] wl[285] vdd gnd cell_6t
Xbit_r286_c12 bl[12] br[12] wl[286] vdd gnd cell_6t
Xbit_r287_c12 bl[12] br[12] wl[287] vdd gnd cell_6t
Xbit_r288_c12 bl[12] br[12] wl[288] vdd gnd cell_6t
Xbit_r289_c12 bl[12] br[12] wl[289] vdd gnd cell_6t
Xbit_r290_c12 bl[12] br[12] wl[290] vdd gnd cell_6t
Xbit_r291_c12 bl[12] br[12] wl[291] vdd gnd cell_6t
Xbit_r292_c12 bl[12] br[12] wl[292] vdd gnd cell_6t
Xbit_r293_c12 bl[12] br[12] wl[293] vdd gnd cell_6t
Xbit_r294_c12 bl[12] br[12] wl[294] vdd gnd cell_6t
Xbit_r295_c12 bl[12] br[12] wl[295] vdd gnd cell_6t
Xbit_r296_c12 bl[12] br[12] wl[296] vdd gnd cell_6t
Xbit_r297_c12 bl[12] br[12] wl[297] vdd gnd cell_6t
Xbit_r298_c12 bl[12] br[12] wl[298] vdd gnd cell_6t
Xbit_r299_c12 bl[12] br[12] wl[299] vdd gnd cell_6t
Xbit_r300_c12 bl[12] br[12] wl[300] vdd gnd cell_6t
Xbit_r301_c12 bl[12] br[12] wl[301] vdd gnd cell_6t
Xbit_r302_c12 bl[12] br[12] wl[302] vdd gnd cell_6t
Xbit_r303_c12 bl[12] br[12] wl[303] vdd gnd cell_6t
Xbit_r304_c12 bl[12] br[12] wl[304] vdd gnd cell_6t
Xbit_r305_c12 bl[12] br[12] wl[305] vdd gnd cell_6t
Xbit_r306_c12 bl[12] br[12] wl[306] vdd gnd cell_6t
Xbit_r307_c12 bl[12] br[12] wl[307] vdd gnd cell_6t
Xbit_r308_c12 bl[12] br[12] wl[308] vdd gnd cell_6t
Xbit_r309_c12 bl[12] br[12] wl[309] vdd gnd cell_6t
Xbit_r310_c12 bl[12] br[12] wl[310] vdd gnd cell_6t
Xbit_r311_c12 bl[12] br[12] wl[311] vdd gnd cell_6t
Xbit_r312_c12 bl[12] br[12] wl[312] vdd gnd cell_6t
Xbit_r313_c12 bl[12] br[12] wl[313] vdd gnd cell_6t
Xbit_r314_c12 bl[12] br[12] wl[314] vdd gnd cell_6t
Xbit_r315_c12 bl[12] br[12] wl[315] vdd gnd cell_6t
Xbit_r316_c12 bl[12] br[12] wl[316] vdd gnd cell_6t
Xbit_r317_c12 bl[12] br[12] wl[317] vdd gnd cell_6t
Xbit_r318_c12 bl[12] br[12] wl[318] vdd gnd cell_6t
Xbit_r319_c12 bl[12] br[12] wl[319] vdd gnd cell_6t
Xbit_r320_c12 bl[12] br[12] wl[320] vdd gnd cell_6t
Xbit_r321_c12 bl[12] br[12] wl[321] vdd gnd cell_6t
Xbit_r322_c12 bl[12] br[12] wl[322] vdd gnd cell_6t
Xbit_r323_c12 bl[12] br[12] wl[323] vdd gnd cell_6t
Xbit_r324_c12 bl[12] br[12] wl[324] vdd gnd cell_6t
Xbit_r325_c12 bl[12] br[12] wl[325] vdd gnd cell_6t
Xbit_r326_c12 bl[12] br[12] wl[326] vdd gnd cell_6t
Xbit_r327_c12 bl[12] br[12] wl[327] vdd gnd cell_6t
Xbit_r328_c12 bl[12] br[12] wl[328] vdd gnd cell_6t
Xbit_r329_c12 bl[12] br[12] wl[329] vdd gnd cell_6t
Xbit_r330_c12 bl[12] br[12] wl[330] vdd gnd cell_6t
Xbit_r331_c12 bl[12] br[12] wl[331] vdd gnd cell_6t
Xbit_r332_c12 bl[12] br[12] wl[332] vdd gnd cell_6t
Xbit_r333_c12 bl[12] br[12] wl[333] vdd gnd cell_6t
Xbit_r334_c12 bl[12] br[12] wl[334] vdd gnd cell_6t
Xbit_r335_c12 bl[12] br[12] wl[335] vdd gnd cell_6t
Xbit_r336_c12 bl[12] br[12] wl[336] vdd gnd cell_6t
Xbit_r337_c12 bl[12] br[12] wl[337] vdd gnd cell_6t
Xbit_r338_c12 bl[12] br[12] wl[338] vdd gnd cell_6t
Xbit_r339_c12 bl[12] br[12] wl[339] vdd gnd cell_6t
Xbit_r340_c12 bl[12] br[12] wl[340] vdd gnd cell_6t
Xbit_r341_c12 bl[12] br[12] wl[341] vdd gnd cell_6t
Xbit_r342_c12 bl[12] br[12] wl[342] vdd gnd cell_6t
Xbit_r343_c12 bl[12] br[12] wl[343] vdd gnd cell_6t
Xbit_r344_c12 bl[12] br[12] wl[344] vdd gnd cell_6t
Xbit_r345_c12 bl[12] br[12] wl[345] vdd gnd cell_6t
Xbit_r346_c12 bl[12] br[12] wl[346] vdd gnd cell_6t
Xbit_r347_c12 bl[12] br[12] wl[347] vdd gnd cell_6t
Xbit_r348_c12 bl[12] br[12] wl[348] vdd gnd cell_6t
Xbit_r349_c12 bl[12] br[12] wl[349] vdd gnd cell_6t
Xbit_r350_c12 bl[12] br[12] wl[350] vdd gnd cell_6t
Xbit_r351_c12 bl[12] br[12] wl[351] vdd gnd cell_6t
Xbit_r352_c12 bl[12] br[12] wl[352] vdd gnd cell_6t
Xbit_r353_c12 bl[12] br[12] wl[353] vdd gnd cell_6t
Xbit_r354_c12 bl[12] br[12] wl[354] vdd gnd cell_6t
Xbit_r355_c12 bl[12] br[12] wl[355] vdd gnd cell_6t
Xbit_r356_c12 bl[12] br[12] wl[356] vdd gnd cell_6t
Xbit_r357_c12 bl[12] br[12] wl[357] vdd gnd cell_6t
Xbit_r358_c12 bl[12] br[12] wl[358] vdd gnd cell_6t
Xbit_r359_c12 bl[12] br[12] wl[359] vdd gnd cell_6t
Xbit_r360_c12 bl[12] br[12] wl[360] vdd gnd cell_6t
Xbit_r361_c12 bl[12] br[12] wl[361] vdd gnd cell_6t
Xbit_r362_c12 bl[12] br[12] wl[362] vdd gnd cell_6t
Xbit_r363_c12 bl[12] br[12] wl[363] vdd gnd cell_6t
Xbit_r364_c12 bl[12] br[12] wl[364] vdd gnd cell_6t
Xbit_r365_c12 bl[12] br[12] wl[365] vdd gnd cell_6t
Xbit_r366_c12 bl[12] br[12] wl[366] vdd gnd cell_6t
Xbit_r367_c12 bl[12] br[12] wl[367] vdd gnd cell_6t
Xbit_r368_c12 bl[12] br[12] wl[368] vdd gnd cell_6t
Xbit_r369_c12 bl[12] br[12] wl[369] vdd gnd cell_6t
Xbit_r370_c12 bl[12] br[12] wl[370] vdd gnd cell_6t
Xbit_r371_c12 bl[12] br[12] wl[371] vdd gnd cell_6t
Xbit_r372_c12 bl[12] br[12] wl[372] vdd gnd cell_6t
Xbit_r373_c12 bl[12] br[12] wl[373] vdd gnd cell_6t
Xbit_r374_c12 bl[12] br[12] wl[374] vdd gnd cell_6t
Xbit_r375_c12 bl[12] br[12] wl[375] vdd gnd cell_6t
Xbit_r376_c12 bl[12] br[12] wl[376] vdd gnd cell_6t
Xbit_r377_c12 bl[12] br[12] wl[377] vdd gnd cell_6t
Xbit_r378_c12 bl[12] br[12] wl[378] vdd gnd cell_6t
Xbit_r379_c12 bl[12] br[12] wl[379] vdd gnd cell_6t
Xbit_r380_c12 bl[12] br[12] wl[380] vdd gnd cell_6t
Xbit_r381_c12 bl[12] br[12] wl[381] vdd gnd cell_6t
Xbit_r382_c12 bl[12] br[12] wl[382] vdd gnd cell_6t
Xbit_r383_c12 bl[12] br[12] wl[383] vdd gnd cell_6t
Xbit_r384_c12 bl[12] br[12] wl[384] vdd gnd cell_6t
Xbit_r385_c12 bl[12] br[12] wl[385] vdd gnd cell_6t
Xbit_r386_c12 bl[12] br[12] wl[386] vdd gnd cell_6t
Xbit_r387_c12 bl[12] br[12] wl[387] vdd gnd cell_6t
Xbit_r388_c12 bl[12] br[12] wl[388] vdd gnd cell_6t
Xbit_r389_c12 bl[12] br[12] wl[389] vdd gnd cell_6t
Xbit_r390_c12 bl[12] br[12] wl[390] vdd gnd cell_6t
Xbit_r391_c12 bl[12] br[12] wl[391] vdd gnd cell_6t
Xbit_r392_c12 bl[12] br[12] wl[392] vdd gnd cell_6t
Xbit_r393_c12 bl[12] br[12] wl[393] vdd gnd cell_6t
Xbit_r394_c12 bl[12] br[12] wl[394] vdd gnd cell_6t
Xbit_r395_c12 bl[12] br[12] wl[395] vdd gnd cell_6t
Xbit_r396_c12 bl[12] br[12] wl[396] vdd gnd cell_6t
Xbit_r397_c12 bl[12] br[12] wl[397] vdd gnd cell_6t
Xbit_r398_c12 bl[12] br[12] wl[398] vdd gnd cell_6t
Xbit_r399_c12 bl[12] br[12] wl[399] vdd gnd cell_6t
Xbit_r400_c12 bl[12] br[12] wl[400] vdd gnd cell_6t
Xbit_r401_c12 bl[12] br[12] wl[401] vdd gnd cell_6t
Xbit_r402_c12 bl[12] br[12] wl[402] vdd gnd cell_6t
Xbit_r403_c12 bl[12] br[12] wl[403] vdd gnd cell_6t
Xbit_r404_c12 bl[12] br[12] wl[404] vdd gnd cell_6t
Xbit_r405_c12 bl[12] br[12] wl[405] vdd gnd cell_6t
Xbit_r406_c12 bl[12] br[12] wl[406] vdd gnd cell_6t
Xbit_r407_c12 bl[12] br[12] wl[407] vdd gnd cell_6t
Xbit_r408_c12 bl[12] br[12] wl[408] vdd gnd cell_6t
Xbit_r409_c12 bl[12] br[12] wl[409] vdd gnd cell_6t
Xbit_r410_c12 bl[12] br[12] wl[410] vdd gnd cell_6t
Xbit_r411_c12 bl[12] br[12] wl[411] vdd gnd cell_6t
Xbit_r412_c12 bl[12] br[12] wl[412] vdd gnd cell_6t
Xbit_r413_c12 bl[12] br[12] wl[413] vdd gnd cell_6t
Xbit_r414_c12 bl[12] br[12] wl[414] vdd gnd cell_6t
Xbit_r415_c12 bl[12] br[12] wl[415] vdd gnd cell_6t
Xbit_r416_c12 bl[12] br[12] wl[416] vdd gnd cell_6t
Xbit_r417_c12 bl[12] br[12] wl[417] vdd gnd cell_6t
Xbit_r418_c12 bl[12] br[12] wl[418] vdd gnd cell_6t
Xbit_r419_c12 bl[12] br[12] wl[419] vdd gnd cell_6t
Xbit_r420_c12 bl[12] br[12] wl[420] vdd gnd cell_6t
Xbit_r421_c12 bl[12] br[12] wl[421] vdd gnd cell_6t
Xbit_r422_c12 bl[12] br[12] wl[422] vdd gnd cell_6t
Xbit_r423_c12 bl[12] br[12] wl[423] vdd gnd cell_6t
Xbit_r424_c12 bl[12] br[12] wl[424] vdd gnd cell_6t
Xbit_r425_c12 bl[12] br[12] wl[425] vdd gnd cell_6t
Xbit_r426_c12 bl[12] br[12] wl[426] vdd gnd cell_6t
Xbit_r427_c12 bl[12] br[12] wl[427] vdd gnd cell_6t
Xbit_r428_c12 bl[12] br[12] wl[428] vdd gnd cell_6t
Xbit_r429_c12 bl[12] br[12] wl[429] vdd gnd cell_6t
Xbit_r430_c12 bl[12] br[12] wl[430] vdd gnd cell_6t
Xbit_r431_c12 bl[12] br[12] wl[431] vdd gnd cell_6t
Xbit_r432_c12 bl[12] br[12] wl[432] vdd gnd cell_6t
Xbit_r433_c12 bl[12] br[12] wl[433] vdd gnd cell_6t
Xbit_r434_c12 bl[12] br[12] wl[434] vdd gnd cell_6t
Xbit_r435_c12 bl[12] br[12] wl[435] vdd gnd cell_6t
Xbit_r436_c12 bl[12] br[12] wl[436] vdd gnd cell_6t
Xbit_r437_c12 bl[12] br[12] wl[437] vdd gnd cell_6t
Xbit_r438_c12 bl[12] br[12] wl[438] vdd gnd cell_6t
Xbit_r439_c12 bl[12] br[12] wl[439] vdd gnd cell_6t
Xbit_r440_c12 bl[12] br[12] wl[440] vdd gnd cell_6t
Xbit_r441_c12 bl[12] br[12] wl[441] vdd gnd cell_6t
Xbit_r442_c12 bl[12] br[12] wl[442] vdd gnd cell_6t
Xbit_r443_c12 bl[12] br[12] wl[443] vdd gnd cell_6t
Xbit_r444_c12 bl[12] br[12] wl[444] vdd gnd cell_6t
Xbit_r445_c12 bl[12] br[12] wl[445] vdd gnd cell_6t
Xbit_r446_c12 bl[12] br[12] wl[446] vdd gnd cell_6t
Xbit_r447_c12 bl[12] br[12] wl[447] vdd gnd cell_6t
Xbit_r448_c12 bl[12] br[12] wl[448] vdd gnd cell_6t
Xbit_r449_c12 bl[12] br[12] wl[449] vdd gnd cell_6t
Xbit_r450_c12 bl[12] br[12] wl[450] vdd gnd cell_6t
Xbit_r451_c12 bl[12] br[12] wl[451] vdd gnd cell_6t
Xbit_r452_c12 bl[12] br[12] wl[452] vdd gnd cell_6t
Xbit_r453_c12 bl[12] br[12] wl[453] vdd gnd cell_6t
Xbit_r454_c12 bl[12] br[12] wl[454] vdd gnd cell_6t
Xbit_r455_c12 bl[12] br[12] wl[455] vdd gnd cell_6t
Xbit_r456_c12 bl[12] br[12] wl[456] vdd gnd cell_6t
Xbit_r457_c12 bl[12] br[12] wl[457] vdd gnd cell_6t
Xbit_r458_c12 bl[12] br[12] wl[458] vdd gnd cell_6t
Xbit_r459_c12 bl[12] br[12] wl[459] vdd gnd cell_6t
Xbit_r460_c12 bl[12] br[12] wl[460] vdd gnd cell_6t
Xbit_r461_c12 bl[12] br[12] wl[461] vdd gnd cell_6t
Xbit_r462_c12 bl[12] br[12] wl[462] vdd gnd cell_6t
Xbit_r463_c12 bl[12] br[12] wl[463] vdd gnd cell_6t
Xbit_r464_c12 bl[12] br[12] wl[464] vdd gnd cell_6t
Xbit_r465_c12 bl[12] br[12] wl[465] vdd gnd cell_6t
Xbit_r466_c12 bl[12] br[12] wl[466] vdd gnd cell_6t
Xbit_r467_c12 bl[12] br[12] wl[467] vdd gnd cell_6t
Xbit_r468_c12 bl[12] br[12] wl[468] vdd gnd cell_6t
Xbit_r469_c12 bl[12] br[12] wl[469] vdd gnd cell_6t
Xbit_r470_c12 bl[12] br[12] wl[470] vdd gnd cell_6t
Xbit_r471_c12 bl[12] br[12] wl[471] vdd gnd cell_6t
Xbit_r472_c12 bl[12] br[12] wl[472] vdd gnd cell_6t
Xbit_r473_c12 bl[12] br[12] wl[473] vdd gnd cell_6t
Xbit_r474_c12 bl[12] br[12] wl[474] vdd gnd cell_6t
Xbit_r475_c12 bl[12] br[12] wl[475] vdd gnd cell_6t
Xbit_r476_c12 bl[12] br[12] wl[476] vdd gnd cell_6t
Xbit_r477_c12 bl[12] br[12] wl[477] vdd gnd cell_6t
Xbit_r478_c12 bl[12] br[12] wl[478] vdd gnd cell_6t
Xbit_r479_c12 bl[12] br[12] wl[479] vdd gnd cell_6t
Xbit_r480_c12 bl[12] br[12] wl[480] vdd gnd cell_6t
Xbit_r481_c12 bl[12] br[12] wl[481] vdd gnd cell_6t
Xbit_r482_c12 bl[12] br[12] wl[482] vdd gnd cell_6t
Xbit_r483_c12 bl[12] br[12] wl[483] vdd gnd cell_6t
Xbit_r484_c12 bl[12] br[12] wl[484] vdd gnd cell_6t
Xbit_r485_c12 bl[12] br[12] wl[485] vdd gnd cell_6t
Xbit_r486_c12 bl[12] br[12] wl[486] vdd gnd cell_6t
Xbit_r487_c12 bl[12] br[12] wl[487] vdd gnd cell_6t
Xbit_r488_c12 bl[12] br[12] wl[488] vdd gnd cell_6t
Xbit_r489_c12 bl[12] br[12] wl[489] vdd gnd cell_6t
Xbit_r490_c12 bl[12] br[12] wl[490] vdd gnd cell_6t
Xbit_r491_c12 bl[12] br[12] wl[491] vdd gnd cell_6t
Xbit_r492_c12 bl[12] br[12] wl[492] vdd gnd cell_6t
Xbit_r493_c12 bl[12] br[12] wl[493] vdd gnd cell_6t
Xbit_r494_c12 bl[12] br[12] wl[494] vdd gnd cell_6t
Xbit_r495_c12 bl[12] br[12] wl[495] vdd gnd cell_6t
Xbit_r496_c12 bl[12] br[12] wl[496] vdd gnd cell_6t
Xbit_r497_c12 bl[12] br[12] wl[497] vdd gnd cell_6t
Xbit_r498_c12 bl[12] br[12] wl[498] vdd gnd cell_6t
Xbit_r499_c12 bl[12] br[12] wl[499] vdd gnd cell_6t
Xbit_r500_c12 bl[12] br[12] wl[500] vdd gnd cell_6t
Xbit_r501_c12 bl[12] br[12] wl[501] vdd gnd cell_6t
Xbit_r502_c12 bl[12] br[12] wl[502] vdd gnd cell_6t
Xbit_r503_c12 bl[12] br[12] wl[503] vdd gnd cell_6t
Xbit_r504_c12 bl[12] br[12] wl[504] vdd gnd cell_6t
Xbit_r505_c12 bl[12] br[12] wl[505] vdd gnd cell_6t
Xbit_r506_c12 bl[12] br[12] wl[506] vdd gnd cell_6t
Xbit_r507_c12 bl[12] br[12] wl[507] vdd gnd cell_6t
Xbit_r508_c12 bl[12] br[12] wl[508] vdd gnd cell_6t
Xbit_r509_c12 bl[12] br[12] wl[509] vdd gnd cell_6t
Xbit_r510_c12 bl[12] br[12] wl[510] vdd gnd cell_6t
Xbit_r511_c12 bl[12] br[12] wl[511] vdd gnd cell_6t
Xbit_r0_c13 bl[13] br[13] wl[0] vdd gnd cell_6t
Xbit_r1_c13 bl[13] br[13] wl[1] vdd gnd cell_6t
Xbit_r2_c13 bl[13] br[13] wl[2] vdd gnd cell_6t
Xbit_r3_c13 bl[13] br[13] wl[3] vdd gnd cell_6t
Xbit_r4_c13 bl[13] br[13] wl[4] vdd gnd cell_6t
Xbit_r5_c13 bl[13] br[13] wl[5] vdd gnd cell_6t
Xbit_r6_c13 bl[13] br[13] wl[6] vdd gnd cell_6t
Xbit_r7_c13 bl[13] br[13] wl[7] vdd gnd cell_6t
Xbit_r8_c13 bl[13] br[13] wl[8] vdd gnd cell_6t
Xbit_r9_c13 bl[13] br[13] wl[9] vdd gnd cell_6t
Xbit_r10_c13 bl[13] br[13] wl[10] vdd gnd cell_6t
Xbit_r11_c13 bl[13] br[13] wl[11] vdd gnd cell_6t
Xbit_r12_c13 bl[13] br[13] wl[12] vdd gnd cell_6t
Xbit_r13_c13 bl[13] br[13] wl[13] vdd gnd cell_6t
Xbit_r14_c13 bl[13] br[13] wl[14] vdd gnd cell_6t
Xbit_r15_c13 bl[13] br[13] wl[15] vdd gnd cell_6t
Xbit_r16_c13 bl[13] br[13] wl[16] vdd gnd cell_6t
Xbit_r17_c13 bl[13] br[13] wl[17] vdd gnd cell_6t
Xbit_r18_c13 bl[13] br[13] wl[18] vdd gnd cell_6t
Xbit_r19_c13 bl[13] br[13] wl[19] vdd gnd cell_6t
Xbit_r20_c13 bl[13] br[13] wl[20] vdd gnd cell_6t
Xbit_r21_c13 bl[13] br[13] wl[21] vdd gnd cell_6t
Xbit_r22_c13 bl[13] br[13] wl[22] vdd gnd cell_6t
Xbit_r23_c13 bl[13] br[13] wl[23] vdd gnd cell_6t
Xbit_r24_c13 bl[13] br[13] wl[24] vdd gnd cell_6t
Xbit_r25_c13 bl[13] br[13] wl[25] vdd gnd cell_6t
Xbit_r26_c13 bl[13] br[13] wl[26] vdd gnd cell_6t
Xbit_r27_c13 bl[13] br[13] wl[27] vdd gnd cell_6t
Xbit_r28_c13 bl[13] br[13] wl[28] vdd gnd cell_6t
Xbit_r29_c13 bl[13] br[13] wl[29] vdd gnd cell_6t
Xbit_r30_c13 bl[13] br[13] wl[30] vdd gnd cell_6t
Xbit_r31_c13 bl[13] br[13] wl[31] vdd gnd cell_6t
Xbit_r32_c13 bl[13] br[13] wl[32] vdd gnd cell_6t
Xbit_r33_c13 bl[13] br[13] wl[33] vdd gnd cell_6t
Xbit_r34_c13 bl[13] br[13] wl[34] vdd gnd cell_6t
Xbit_r35_c13 bl[13] br[13] wl[35] vdd gnd cell_6t
Xbit_r36_c13 bl[13] br[13] wl[36] vdd gnd cell_6t
Xbit_r37_c13 bl[13] br[13] wl[37] vdd gnd cell_6t
Xbit_r38_c13 bl[13] br[13] wl[38] vdd gnd cell_6t
Xbit_r39_c13 bl[13] br[13] wl[39] vdd gnd cell_6t
Xbit_r40_c13 bl[13] br[13] wl[40] vdd gnd cell_6t
Xbit_r41_c13 bl[13] br[13] wl[41] vdd gnd cell_6t
Xbit_r42_c13 bl[13] br[13] wl[42] vdd gnd cell_6t
Xbit_r43_c13 bl[13] br[13] wl[43] vdd gnd cell_6t
Xbit_r44_c13 bl[13] br[13] wl[44] vdd gnd cell_6t
Xbit_r45_c13 bl[13] br[13] wl[45] vdd gnd cell_6t
Xbit_r46_c13 bl[13] br[13] wl[46] vdd gnd cell_6t
Xbit_r47_c13 bl[13] br[13] wl[47] vdd gnd cell_6t
Xbit_r48_c13 bl[13] br[13] wl[48] vdd gnd cell_6t
Xbit_r49_c13 bl[13] br[13] wl[49] vdd gnd cell_6t
Xbit_r50_c13 bl[13] br[13] wl[50] vdd gnd cell_6t
Xbit_r51_c13 bl[13] br[13] wl[51] vdd gnd cell_6t
Xbit_r52_c13 bl[13] br[13] wl[52] vdd gnd cell_6t
Xbit_r53_c13 bl[13] br[13] wl[53] vdd gnd cell_6t
Xbit_r54_c13 bl[13] br[13] wl[54] vdd gnd cell_6t
Xbit_r55_c13 bl[13] br[13] wl[55] vdd gnd cell_6t
Xbit_r56_c13 bl[13] br[13] wl[56] vdd gnd cell_6t
Xbit_r57_c13 bl[13] br[13] wl[57] vdd gnd cell_6t
Xbit_r58_c13 bl[13] br[13] wl[58] vdd gnd cell_6t
Xbit_r59_c13 bl[13] br[13] wl[59] vdd gnd cell_6t
Xbit_r60_c13 bl[13] br[13] wl[60] vdd gnd cell_6t
Xbit_r61_c13 bl[13] br[13] wl[61] vdd gnd cell_6t
Xbit_r62_c13 bl[13] br[13] wl[62] vdd gnd cell_6t
Xbit_r63_c13 bl[13] br[13] wl[63] vdd gnd cell_6t
Xbit_r64_c13 bl[13] br[13] wl[64] vdd gnd cell_6t
Xbit_r65_c13 bl[13] br[13] wl[65] vdd gnd cell_6t
Xbit_r66_c13 bl[13] br[13] wl[66] vdd gnd cell_6t
Xbit_r67_c13 bl[13] br[13] wl[67] vdd gnd cell_6t
Xbit_r68_c13 bl[13] br[13] wl[68] vdd gnd cell_6t
Xbit_r69_c13 bl[13] br[13] wl[69] vdd gnd cell_6t
Xbit_r70_c13 bl[13] br[13] wl[70] vdd gnd cell_6t
Xbit_r71_c13 bl[13] br[13] wl[71] vdd gnd cell_6t
Xbit_r72_c13 bl[13] br[13] wl[72] vdd gnd cell_6t
Xbit_r73_c13 bl[13] br[13] wl[73] vdd gnd cell_6t
Xbit_r74_c13 bl[13] br[13] wl[74] vdd gnd cell_6t
Xbit_r75_c13 bl[13] br[13] wl[75] vdd gnd cell_6t
Xbit_r76_c13 bl[13] br[13] wl[76] vdd gnd cell_6t
Xbit_r77_c13 bl[13] br[13] wl[77] vdd gnd cell_6t
Xbit_r78_c13 bl[13] br[13] wl[78] vdd gnd cell_6t
Xbit_r79_c13 bl[13] br[13] wl[79] vdd gnd cell_6t
Xbit_r80_c13 bl[13] br[13] wl[80] vdd gnd cell_6t
Xbit_r81_c13 bl[13] br[13] wl[81] vdd gnd cell_6t
Xbit_r82_c13 bl[13] br[13] wl[82] vdd gnd cell_6t
Xbit_r83_c13 bl[13] br[13] wl[83] vdd gnd cell_6t
Xbit_r84_c13 bl[13] br[13] wl[84] vdd gnd cell_6t
Xbit_r85_c13 bl[13] br[13] wl[85] vdd gnd cell_6t
Xbit_r86_c13 bl[13] br[13] wl[86] vdd gnd cell_6t
Xbit_r87_c13 bl[13] br[13] wl[87] vdd gnd cell_6t
Xbit_r88_c13 bl[13] br[13] wl[88] vdd gnd cell_6t
Xbit_r89_c13 bl[13] br[13] wl[89] vdd gnd cell_6t
Xbit_r90_c13 bl[13] br[13] wl[90] vdd gnd cell_6t
Xbit_r91_c13 bl[13] br[13] wl[91] vdd gnd cell_6t
Xbit_r92_c13 bl[13] br[13] wl[92] vdd gnd cell_6t
Xbit_r93_c13 bl[13] br[13] wl[93] vdd gnd cell_6t
Xbit_r94_c13 bl[13] br[13] wl[94] vdd gnd cell_6t
Xbit_r95_c13 bl[13] br[13] wl[95] vdd gnd cell_6t
Xbit_r96_c13 bl[13] br[13] wl[96] vdd gnd cell_6t
Xbit_r97_c13 bl[13] br[13] wl[97] vdd gnd cell_6t
Xbit_r98_c13 bl[13] br[13] wl[98] vdd gnd cell_6t
Xbit_r99_c13 bl[13] br[13] wl[99] vdd gnd cell_6t
Xbit_r100_c13 bl[13] br[13] wl[100] vdd gnd cell_6t
Xbit_r101_c13 bl[13] br[13] wl[101] vdd gnd cell_6t
Xbit_r102_c13 bl[13] br[13] wl[102] vdd gnd cell_6t
Xbit_r103_c13 bl[13] br[13] wl[103] vdd gnd cell_6t
Xbit_r104_c13 bl[13] br[13] wl[104] vdd gnd cell_6t
Xbit_r105_c13 bl[13] br[13] wl[105] vdd gnd cell_6t
Xbit_r106_c13 bl[13] br[13] wl[106] vdd gnd cell_6t
Xbit_r107_c13 bl[13] br[13] wl[107] vdd gnd cell_6t
Xbit_r108_c13 bl[13] br[13] wl[108] vdd gnd cell_6t
Xbit_r109_c13 bl[13] br[13] wl[109] vdd gnd cell_6t
Xbit_r110_c13 bl[13] br[13] wl[110] vdd gnd cell_6t
Xbit_r111_c13 bl[13] br[13] wl[111] vdd gnd cell_6t
Xbit_r112_c13 bl[13] br[13] wl[112] vdd gnd cell_6t
Xbit_r113_c13 bl[13] br[13] wl[113] vdd gnd cell_6t
Xbit_r114_c13 bl[13] br[13] wl[114] vdd gnd cell_6t
Xbit_r115_c13 bl[13] br[13] wl[115] vdd gnd cell_6t
Xbit_r116_c13 bl[13] br[13] wl[116] vdd gnd cell_6t
Xbit_r117_c13 bl[13] br[13] wl[117] vdd gnd cell_6t
Xbit_r118_c13 bl[13] br[13] wl[118] vdd gnd cell_6t
Xbit_r119_c13 bl[13] br[13] wl[119] vdd gnd cell_6t
Xbit_r120_c13 bl[13] br[13] wl[120] vdd gnd cell_6t
Xbit_r121_c13 bl[13] br[13] wl[121] vdd gnd cell_6t
Xbit_r122_c13 bl[13] br[13] wl[122] vdd gnd cell_6t
Xbit_r123_c13 bl[13] br[13] wl[123] vdd gnd cell_6t
Xbit_r124_c13 bl[13] br[13] wl[124] vdd gnd cell_6t
Xbit_r125_c13 bl[13] br[13] wl[125] vdd gnd cell_6t
Xbit_r126_c13 bl[13] br[13] wl[126] vdd gnd cell_6t
Xbit_r127_c13 bl[13] br[13] wl[127] vdd gnd cell_6t
Xbit_r128_c13 bl[13] br[13] wl[128] vdd gnd cell_6t
Xbit_r129_c13 bl[13] br[13] wl[129] vdd gnd cell_6t
Xbit_r130_c13 bl[13] br[13] wl[130] vdd gnd cell_6t
Xbit_r131_c13 bl[13] br[13] wl[131] vdd gnd cell_6t
Xbit_r132_c13 bl[13] br[13] wl[132] vdd gnd cell_6t
Xbit_r133_c13 bl[13] br[13] wl[133] vdd gnd cell_6t
Xbit_r134_c13 bl[13] br[13] wl[134] vdd gnd cell_6t
Xbit_r135_c13 bl[13] br[13] wl[135] vdd gnd cell_6t
Xbit_r136_c13 bl[13] br[13] wl[136] vdd gnd cell_6t
Xbit_r137_c13 bl[13] br[13] wl[137] vdd gnd cell_6t
Xbit_r138_c13 bl[13] br[13] wl[138] vdd gnd cell_6t
Xbit_r139_c13 bl[13] br[13] wl[139] vdd gnd cell_6t
Xbit_r140_c13 bl[13] br[13] wl[140] vdd gnd cell_6t
Xbit_r141_c13 bl[13] br[13] wl[141] vdd gnd cell_6t
Xbit_r142_c13 bl[13] br[13] wl[142] vdd gnd cell_6t
Xbit_r143_c13 bl[13] br[13] wl[143] vdd gnd cell_6t
Xbit_r144_c13 bl[13] br[13] wl[144] vdd gnd cell_6t
Xbit_r145_c13 bl[13] br[13] wl[145] vdd gnd cell_6t
Xbit_r146_c13 bl[13] br[13] wl[146] vdd gnd cell_6t
Xbit_r147_c13 bl[13] br[13] wl[147] vdd gnd cell_6t
Xbit_r148_c13 bl[13] br[13] wl[148] vdd gnd cell_6t
Xbit_r149_c13 bl[13] br[13] wl[149] vdd gnd cell_6t
Xbit_r150_c13 bl[13] br[13] wl[150] vdd gnd cell_6t
Xbit_r151_c13 bl[13] br[13] wl[151] vdd gnd cell_6t
Xbit_r152_c13 bl[13] br[13] wl[152] vdd gnd cell_6t
Xbit_r153_c13 bl[13] br[13] wl[153] vdd gnd cell_6t
Xbit_r154_c13 bl[13] br[13] wl[154] vdd gnd cell_6t
Xbit_r155_c13 bl[13] br[13] wl[155] vdd gnd cell_6t
Xbit_r156_c13 bl[13] br[13] wl[156] vdd gnd cell_6t
Xbit_r157_c13 bl[13] br[13] wl[157] vdd gnd cell_6t
Xbit_r158_c13 bl[13] br[13] wl[158] vdd gnd cell_6t
Xbit_r159_c13 bl[13] br[13] wl[159] vdd gnd cell_6t
Xbit_r160_c13 bl[13] br[13] wl[160] vdd gnd cell_6t
Xbit_r161_c13 bl[13] br[13] wl[161] vdd gnd cell_6t
Xbit_r162_c13 bl[13] br[13] wl[162] vdd gnd cell_6t
Xbit_r163_c13 bl[13] br[13] wl[163] vdd gnd cell_6t
Xbit_r164_c13 bl[13] br[13] wl[164] vdd gnd cell_6t
Xbit_r165_c13 bl[13] br[13] wl[165] vdd gnd cell_6t
Xbit_r166_c13 bl[13] br[13] wl[166] vdd gnd cell_6t
Xbit_r167_c13 bl[13] br[13] wl[167] vdd gnd cell_6t
Xbit_r168_c13 bl[13] br[13] wl[168] vdd gnd cell_6t
Xbit_r169_c13 bl[13] br[13] wl[169] vdd gnd cell_6t
Xbit_r170_c13 bl[13] br[13] wl[170] vdd gnd cell_6t
Xbit_r171_c13 bl[13] br[13] wl[171] vdd gnd cell_6t
Xbit_r172_c13 bl[13] br[13] wl[172] vdd gnd cell_6t
Xbit_r173_c13 bl[13] br[13] wl[173] vdd gnd cell_6t
Xbit_r174_c13 bl[13] br[13] wl[174] vdd gnd cell_6t
Xbit_r175_c13 bl[13] br[13] wl[175] vdd gnd cell_6t
Xbit_r176_c13 bl[13] br[13] wl[176] vdd gnd cell_6t
Xbit_r177_c13 bl[13] br[13] wl[177] vdd gnd cell_6t
Xbit_r178_c13 bl[13] br[13] wl[178] vdd gnd cell_6t
Xbit_r179_c13 bl[13] br[13] wl[179] vdd gnd cell_6t
Xbit_r180_c13 bl[13] br[13] wl[180] vdd gnd cell_6t
Xbit_r181_c13 bl[13] br[13] wl[181] vdd gnd cell_6t
Xbit_r182_c13 bl[13] br[13] wl[182] vdd gnd cell_6t
Xbit_r183_c13 bl[13] br[13] wl[183] vdd gnd cell_6t
Xbit_r184_c13 bl[13] br[13] wl[184] vdd gnd cell_6t
Xbit_r185_c13 bl[13] br[13] wl[185] vdd gnd cell_6t
Xbit_r186_c13 bl[13] br[13] wl[186] vdd gnd cell_6t
Xbit_r187_c13 bl[13] br[13] wl[187] vdd gnd cell_6t
Xbit_r188_c13 bl[13] br[13] wl[188] vdd gnd cell_6t
Xbit_r189_c13 bl[13] br[13] wl[189] vdd gnd cell_6t
Xbit_r190_c13 bl[13] br[13] wl[190] vdd gnd cell_6t
Xbit_r191_c13 bl[13] br[13] wl[191] vdd gnd cell_6t
Xbit_r192_c13 bl[13] br[13] wl[192] vdd gnd cell_6t
Xbit_r193_c13 bl[13] br[13] wl[193] vdd gnd cell_6t
Xbit_r194_c13 bl[13] br[13] wl[194] vdd gnd cell_6t
Xbit_r195_c13 bl[13] br[13] wl[195] vdd gnd cell_6t
Xbit_r196_c13 bl[13] br[13] wl[196] vdd gnd cell_6t
Xbit_r197_c13 bl[13] br[13] wl[197] vdd gnd cell_6t
Xbit_r198_c13 bl[13] br[13] wl[198] vdd gnd cell_6t
Xbit_r199_c13 bl[13] br[13] wl[199] vdd gnd cell_6t
Xbit_r200_c13 bl[13] br[13] wl[200] vdd gnd cell_6t
Xbit_r201_c13 bl[13] br[13] wl[201] vdd gnd cell_6t
Xbit_r202_c13 bl[13] br[13] wl[202] vdd gnd cell_6t
Xbit_r203_c13 bl[13] br[13] wl[203] vdd gnd cell_6t
Xbit_r204_c13 bl[13] br[13] wl[204] vdd gnd cell_6t
Xbit_r205_c13 bl[13] br[13] wl[205] vdd gnd cell_6t
Xbit_r206_c13 bl[13] br[13] wl[206] vdd gnd cell_6t
Xbit_r207_c13 bl[13] br[13] wl[207] vdd gnd cell_6t
Xbit_r208_c13 bl[13] br[13] wl[208] vdd gnd cell_6t
Xbit_r209_c13 bl[13] br[13] wl[209] vdd gnd cell_6t
Xbit_r210_c13 bl[13] br[13] wl[210] vdd gnd cell_6t
Xbit_r211_c13 bl[13] br[13] wl[211] vdd gnd cell_6t
Xbit_r212_c13 bl[13] br[13] wl[212] vdd gnd cell_6t
Xbit_r213_c13 bl[13] br[13] wl[213] vdd gnd cell_6t
Xbit_r214_c13 bl[13] br[13] wl[214] vdd gnd cell_6t
Xbit_r215_c13 bl[13] br[13] wl[215] vdd gnd cell_6t
Xbit_r216_c13 bl[13] br[13] wl[216] vdd gnd cell_6t
Xbit_r217_c13 bl[13] br[13] wl[217] vdd gnd cell_6t
Xbit_r218_c13 bl[13] br[13] wl[218] vdd gnd cell_6t
Xbit_r219_c13 bl[13] br[13] wl[219] vdd gnd cell_6t
Xbit_r220_c13 bl[13] br[13] wl[220] vdd gnd cell_6t
Xbit_r221_c13 bl[13] br[13] wl[221] vdd gnd cell_6t
Xbit_r222_c13 bl[13] br[13] wl[222] vdd gnd cell_6t
Xbit_r223_c13 bl[13] br[13] wl[223] vdd gnd cell_6t
Xbit_r224_c13 bl[13] br[13] wl[224] vdd gnd cell_6t
Xbit_r225_c13 bl[13] br[13] wl[225] vdd gnd cell_6t
Xbit_r226_c13 bl[13] br[13] wl[226] vdd gnd cell_6t
Xbit_r227_c13 bl[13] br[13] wl[227] vdd gnd cell_6t
Xbit_r228_c13 bl[13] br[13] wl[228] vdd gnd cell_6t
Xbit_r229_c13 bl[13] br[13] wl[229] vdd gnd cell_6t
Xbit_r230_c13 bl[13] br[13] wl[230] vdd gnd cell_6t
Xbit_r231_c13 bl[13] br[13] wl[231] vdd gnd cell_6t
Xbit_r232_c13 bl[13] br[13] wl[232] vdd gnd cell_6t
Xbit_r233_c13 bl[13] br[13] wl[233] vdd gnd cell_6t
Xbit_r234_c13 bl[13] br[13] wl[234] vdd gnd cell_6t
Xbit_r235_c13 bl[13] br[13] wl[235] vdd gnd cell_6t
Xbit_r236_c13 bl[13] br[13] wl[236] vdd gnd cell_6t
Xbit_r237_c13 bl[13] br[13] wl[237] vdd gnd cell_6t
Xbit_r238_c13 bl[13] br[13] wl[238] vdd gnd cell_6t
Xbit_r239_c13 bl[13] br[13] wl[239] vdd gnd cell_6t
Xbit_r240_c13 bl[13] br[13] wl[240] vdd gnd cell_6t
Xbit_r241_c13 bl[13] br[13] wl[241] vdd gnd cell_6t
Xbit_r242_c13 bl[13] br[13] wl[242] vdd gnd cell_6t
Xbit_r243_c13 bl[13] br[13] wl[243] vdd gnd cell_6t
Xbit_r244_c13 bl[13] br[13] wl[244] vdd gnd cell_6t
Xbit_r245_c13 bl[13] br[13] wl[245] vdd gnd cell_6t
Xbit_r246_c13 bl[13] br[13] wl[246] vdd gnd cell_6t
Xbit_r247_c13 bl[13] br[13] wl[247] vdd gnd cell_6t
Xbit_r248_c13 bl[13] br[13] wl[248] vdd gnd cell_6t
Xbit_r249_c13 bl[13] br[13] wl[249] vdd gnd cell_6t
Xbit_r250_c13 bl[13] br[13] wl[250] vdd gnd cell_6t
Xbit_r251_c13 bl[13] br[13] wl[251] vdd gnd cell_6t
Xbit_r252_c13 bl[13] br[13] wl[252] vdd gnd cell_6t
Xbit_r253_c13 bl[13] br[13] wl[253] vdd gnd cell_6t
Xbit_r254_c13 bl[13] br[13] wl[254] vdd gnd cell_6t
Xbit_r255_c13 bl[13] br[13] wl[255] vdd gnd cell_6t
Xbit_r256_c13 bl[13] br[13] wl[256] vdd gnd cell_6t
Xbit_r257_c13 bl[13] br[13] wl[257] vdd gnd cell_6t
Xbit_r258_c13 bl[13] br[13] wl[258] vdd gnd cell_6t
Xbit_r259_c13 bl[13] br[13] wl[259] vdd gnd cell_6t
Xbit_r260_c13 bl[13] br[13] wl[260] vdd gnd cell_6t
Xbit_r261_c13 bl[13] br[13] wl[261] vdd gnd cell_6t
Xbit_r262_c13 bl[13] br[13] wl[262] vdd gnd cell_6t
Xbit_r263_c13 bl[13] br[13] wl[263] vdd gnd cell_6t
Xbit_r264_c13 bl[13] br[13] wl[264] vdd gnd cell_6t
Xbit_r265_c13 bl[13] br[13] wl[265] vdd gnd cell_6t
Xbit_r266_c13 bl[13] br[13] wl[266] vdd gnd cell_6t
Xbit_r267_c13 bl[13] br[13] wl[267] vdd gnd cell_6t
Xbit_r268_c13 bl[13] br[13] wl[268] vdd gnd cell_6t
Xbit_r269_c13 bl[13] br[13] wl[269] vdd gnd cell_6t
Xbit_r270_c13 bl[13] br[13] wl[270] vdd gnd cell_6t
Xbit_r271_c13 bl[13] br[13] wl[271] vdd gnd cell_6t
Xbit_r272_c13 bl[13] br[13] wl[272] vdd gnd cell_6t
Xbit_r273_c13 bl[13] br[13] wl[273] vdd gnd cell_6t
Xbit_r274_c13 bl[13] br[13] wl[274] vdd gnd cell_6t
Xbit_r275_c13 bl[13] br[13] wl[275] vdd gnd cell_6t
Xbit_r276_c13 bl[13] br[13] wl[276] vdd gnd cell_6t
Xbit_r277_c13 bl[13] br[13] wl[277] vdd gnd cell_6t
Xbit_r278_c13 bl[13] br[13] wl[278] vdd gnd cell_6t
Xbit_r279_c13 bl[13] br[13] wl[279] vdd gnd cell_6t
Xbit_r280_c13 bl[13] br[13] wl[280] vdd gnd cell_6t
Xbit_r281_c13 bl[13] br[13] wl[281] vdd gnd cell_6t
Xbit_r282_c13 bl[13] br[13] wl[282] vdd gnd cell_6t
Xbit_r283_c13 bl[13] br[13] wl[283] vdd gnd cell_6t
Xbit_r284_c13 bl[13] br[13] wl[284] vdd gnd cell_6t
Xbit_r285_c13 bl[13] br[13] wl[285] vdd gnd cell_6t
Xbit_r286_c13 bl[13] br[13] wl[286] vdd gnd cell_6t
Xbit_r287_c13 bl[13] br[13] wl[287] vdd gnd cell_6t
Xbit_r288_c13 bl[13] br[13] wl[288] vdd gnd cell_6t
Xbit_r289_c13 bl[13] br[13] wl[289] vdd gnd cell_6t
Xbit_r290_c13 bl[13] br[13] wl[290] vdd gnd cell_6t
Xbit_r291_c13 bl[13] br[13] wl[291] vdd gnd cell_6t
Xbit_r292_c13 bl[13] br[13] wl[292] vdd gnd cell_6t
Xbit_r293_c13 bl[13] br[13] wl[293] vdd gnd cell_6t
Xbit_r294_c13 bl[13] br[13] wl[294] vdd gnd cell_6t
Xbit_r295_c13 bl[13] br[13] wl[295] vdd gnd cell_6t
Xbit_r296_c13 bl[13] br[13] wl[296] vdd gnd cell_6t
Xbit_r297_c13 bl[13] br[13] wl[297] vdd gnd cell_6t
Xbit_r298_c13 bl[13] br[13] wl[298] vdd gnd cell_6t
Xbit_r299_c13 bl[13] br[13] wl[299] vdd gnd cell_6t
Xbit_r300_c13 bl[13] br[13] wl[300] vdd gnd cell_6t
Xbit_r301_c13 bl[13] br[13] wl[301] vdd gnd cell_6t
Xbit_r302_c13 bl[13] br[13] wl[302] vdd gnd cell_6t
Xbit_r303_c13 bl[13] br[13] wl[303] vdd gnd cell_6t
Xbit_r304_c13 bl[13] br[13] wl[304] vdd gnd cell_6t
Xbit_r305_c13 bl[13] br[13] wl[305] vdd gnd cell_6t
Xbit_r306_c13 bl[13] br[13] wl[306] vdd gnd cell_6t
Xbit_r307_c13 bl[13] br[13] wl[307] vdd gnd cell_6t
Xbit_r308_c13 bl[13] br[13] wl[308] vdd gnd cell_6t
Xbit_r309_c13 bl[13] br[13] wl[309] vdd gnd cell_6t
Xbit_r310_c13 bl[13] br[13] wl[310] vdd gnd cell_6t
Xbit_r311_c13 bl[13] br[13] wl[311] vdd gnd cell_6t
Xbit_r312_c13 bl[13] br[13] wl[312] vdd gnd cell_6t
Xbit_r313_c13 bl[13] br[13] wl[313] vdd gnd cell_6t
Xbit_r314_c13 bl[13] br[13] wl[314] vdd gnd cell_6t
Xbit_r315_c13 bl[13] br[13] wl[315] vdd gnd cell_6t
Xbit_r316_c13 bl[13] br[13] wl[316] vdd gnd cell_6t
Xbit_r317_c13 bl[13] br[13] wl[317] vdd gnd cell_6t
Xbit_r318_c13 bl[13] br[13] wl[318] vdd gnd cell_6t
Xbit_r319_c13 bl[13] br[13] wl[319] vdd gnd cell_6t
Xbit_r320_c13 bl[13] br[13] wl[320] vdd gnd cell_6t
Xbit_r321_c13 bl[13] br[13] wl[321] vdd gnd cell_6t
Xbit_r322_c13 bl[13] br[13] wl[322] vdd gnd cell_6t
Xbit_r323_c13 bl[13] br[13] wl[323] vdd gnd cell_6t
Xbit_r324_c13 bl[13] br[13] wl[324] vdd gnd cell_6t
Xbit_r325_c13 bl[13] br[13] wl[325] vdd gnd cell_6t
Xbit_r326_c13 bl[13] br[13] wl[326] vdd gnd cell_6t
Xbit_r327_c13 bl[13] br[13] wl[327] vdd gnd cell_6t
Xbit_r328_c13 bl[13] br[13] wl[328] vdd gnd cell_6t
Xbit_r329_c13 bl[13] br[13] wl[329] vdd gnd cell_6t
Xbit_r330_c13 bl[13] br[13] wl[330] vdd gnd cell_6t
Xbit_r331_c13 bl[13] br[13] wl[331] vdd gnd cell_6t
Xbit_r332_c13 bl[13] br[13] wl[332] vdd gnd cell_6t
Xbit_r333_c13 bl[13] br[13] wl[333] vdd gnd cell_6t
Xbit_r334_c13 bl[13] br[13] wl[334] vdd gnd cell_6t
Xbit_r335_c13 bl[13] br[13] wl[335] vdd gnd cell_6t
Xbit_r336_c13 bl[13] br[13] wl[336] vdd gnd cell_6t
Xbit_r337_c13 bl[13] br[13] wl[337] vdd gnd cell_6t
Xbit_r338_c13 bl[13] br[13] wl[338] vdd gnd cell_6t
Xbit_r339_c13 bl[13] br[13] wl[339] vdd gnd cell_6t
Xbit_r340_c13 bl[13] br[13] wl[340] vdd gnd cell_6t
Xbit_r341_c13 bl[13] br[13] wl[341] vdd gnd cell_6t
Xbit_r342_c13 bl[13] br[13] wl[342] vdd gnd cell_6t
Xbit_r343_c13 bl[13] br[13] wl[343] vdd gnd cell_6t
Xbit_r344_c13 bl[13] br[13] wl[344] vdd gnd cell_6t
Xbit_r345_c13 bl[13] br[13] wl[345] vdd gnd cell_6t
Xbit_r346_c13 bl[13] br[13] wl[346] vdd gnd cell_6t
Xbit_r347_c13 bl[13] br[13] wl[347] vdd gnd cell_6t
Xbit_r348_c13 bl[13] br[13] wl[348] vdd gnd cell_6t
Xbit_r349_c13 bl[13] br[13] wl[349] vdd gnd cell_6t
Xbit_r350_c13 bl[13] br[13] wl[350] vdd gnd cell_6t
Xbit_r351_c13 bl[13] br[13] wl[351] vdd gnd cell_6t
Xbit_r352_c13 bl[13] br[13] wl[352] vdd gnd cell_6t
Xbit_r353_c13 bl[13] br[13] wl[353] vdd gnd cell_6t
Xbit_r354_c13 bl[13] br[13] wl[354] vdd gnd cell_6t
Xbit_r355_c13 bl[13] br[13] wl[355] vdd gnd cell_6t
Xbit_r356_c13 bl[13] br[13] wl[356] vdd gnd cell_6t
Xbit_r357_c13 bl[13] br[13] wl[357] vdd gnd cell_6t
Xbit_r358_c13 bl[13] br[13] wl[358] vdd gnd cell_6t
Xbit_r359_c13 bl[13] br[13] wl[359] vdd gnd cell_6t
Xbit_r360_c13 bl[13] br[13] wl[360] vdd gnd cell_6t
Xbit_r361_c13 bl[13] br[13] wl[361] vdd gnd cell_6t
Xbit_r362_c13 bl[13] br[13] wl[362] vdd gnd cell_6t
Xbit_r363_c13 bl[13] br[13] wl[363] vdd gnd cell_6t
Xbit_r364_c13 bl[13] br[13] wl[364] vdd gnd cell_6t
Xbit_r365_c13 bl[13] br[13] wl[365] vdd gnd cell_6t
Xbit_r366_c13 bl[13] br[13] wl[366] vdd gnd cell_6t
Xbit_r367_c13 bl[13] br[13] wl[367] vdd gnd cell_6t
Xbit_r368_c13 bl[13] br[13] wl[368] vdd gnd cell_6t
Xbit_r369_c13 bl[13] br[13] wl[369] vdd gnd cell_6t
Xbit_r370_c13 bl[13] br[13] wl[370] vdd gnd cell_6t
Xbit_r371_c13 bl[13] br[13] wl[371] vdd gnd cell_6t
Xbit_r372_c13 bl[13] br[13] wl[372] vdd gnd cell_6t
Xbit_r373_c13 bl[13] br[13] wl[373] vdd gnd cell_6t
Xbit_r374_c13 bl[13] br[13] wl[374] vdd gnd cell_6t
Xbit_r375_c13 bl[13] br[13] wl[375] vdd gnd cell_6t
Xbit_r376_c13 bl[13] br[13] wl[376] vdd gnd cell_6t
Xbit_r377_c13 bl[13] br[13] wl[377] vdd gnd cell_6t
Xbit_r378_c13 bl[13] br[13] wl[378] vdd gnd cell_6t
Xbit_r379_c13 bl[13] br[13] wl[379] vdd gnd cell_6t
Xbit_r380_c13 bl[13] br[13] wl[380] vdd gnd cell_6t
Xbit_r381_c13 bl[13] br[13] wl[381] vdd gnd cell_6t
Xbit_r382_c13 bl[13] br[13] wl[382] vdd gnd cell_6t
Xbit_r383_c13 bl[13] br[13] wl[383] vdd gnd cell_6t
Xbit_r384_c13 bl[13] br[13] wl[384] vdd gnd cell_6t
Xbit_r385_c13 bl[13] br[13] wl[385] vdd gnd cell_6t
Xbit_r386_c13 bl[13] br[13] wl[386] vdd gnd cell_6t
Xbit_r387_c13 bl[13] br[13] wl[387] vdd gnd cell_6t
Xbit_r388_c13 bl[13] br[13] wl[388] vdd gnd cell_6t
Xbit_r389_c13 bl[13] br[13] wl[389] vdd gnd cell_6t
Xbit_r390_c13 bl[13] br[13] wl[390] vdd gnd cell_6t
Xbit_r391_c13 bl[13] br[13] wl[391] vdd gnd cell_6t
Xbit_r392_c13 bl[13] br[13] wl[392] vdd gnd cell_6t
Xbit_r393_c13 bl[13] br[13] wl[393] vdd gnd cell_6t
Xbit_r394_c13 bl[13] br[13] wl[394] vdd gnd cell_6t
Xbit_r395_c13 bl[13] br[13] wl[395] vdd gnd cell_6t
Xbit_r396_c13 bl[13] br[13] wl[396] vdd gnd cell_6t
Xbit_r397_c13 bl[13] br[13] wl[397] vdd gnd cell_6t
Xbit_r398_c13 bl[13] br[13] wl[398] vdd gnd cell_6t
Xbit_r399_c13 bl[13] br[13] wl[399] vdd gnd cell_6t
Xbit_r400_c13 bl[13] br[13] wl[400] vdd gnd cell_6t
Xbit_r401_c13 bl[13] br[13] wl[401] vdd gnd cell_6t
Xbit_r402_c13 bl[13] br[13] wl[402] vdd gnd cell_6t
Xbit_r403_c13 bl[13] br[13] wl[403] vdd gnd cell_6t
Xbit_r404_c13 bl[13] br[13] wl[404] vdd gnd cell_6t
Xbit_r405_c13 bl[13] br[13] wl[405] vdd gnd cell_6t
Xbit_r406_c13 bl[13] br[13] wl[406] vdd gnd cell_6t
Xbit_r407_c13 bl[13] br[13] wl[407] vdd gnd cell_6t
Xbit_r408_c13 bl[13] br[13] wl[408] vdd gnd cell_6t
Xbit_r409_c13 bl[13] br[13] wl[409] vdd gnd cell_6t
Xbit_r410_c13 bl[13] br[13] wl[410] vdd gnd cell_6t
Xbit_r411_c13 bl[13] br[13] wl[411] vdd gnd cell_6t
Xbit_r412_c13 bl[13] br[13] wl[412] vdd gnd cell_6t
Xbit_r413_c13 bl[13] br[13] wl[413] vdd gnd cell_6t
Xbit_r414_c13 bl[13] br[13] wl[414] vdd gnd cell_6t
Xbit_r415_c13 bl[13] br[13] wl[415] vdd gnd cell_6t
Xbit_r416_c13 bl[13] br[13] wl[416] vdd gnd cell_6t
Xbit_r417_c13 bl[13] br[13] wl[417] vdd gnd cell_6t
Xbit_r418_c13 bl[13] br[13] wl[418] vdd gnd cell_6t
Xbit_r419_c13 bl[13] br[13] wl[419] vdd gnd cell_6t
Xbit_r420_c13 bl[13] br[13] wl[420] vdd gnd cell_6t
Xbit_r421_c13 bl[13] br[13] wl[421] vdd gnd cell_6t
Xbit_r422_c13 bl[13] br[13] wl[422] vdd gnd cell_6t
Xbit_r423_c13 bl[13] br[13] wl[423] vdd gnd cell_6t
Xbit_r424_c13 bl[13] br[13] wl[424] vdd gnd cell_6t
Xbit_r425_c13 bl[13] br[13] wl[425] vdd gnd cell_6t
Xbit_r426_c13 bl[13] br[13] wl[426] vdd gnd cell_6t
Xbit_r427_c13 bl[13] br[13] wl[427] vdd gnd cell_6t
Xbit_r428_c13 bl[13] br[13] wl[428] vdd gnd cell_6t
Xbit_r429_c13 bl[13] br[13] wl[429] vdd gnd cell_6t
Xbit_r430_c13 bl[13] br[13] wl[430] vdd gnd cell_6t
Xbit_r431_c13 bl[13] br[13] wl[431] vdd gnd cell_6t
Xbit_r432_c13 bl[13] br[13] wl[432] vdd gnd cell_6t
Xbit_r433_c13 bl[13] br[13] wl[433] vdd gnd cell_6t
Xbit_r434_c13 bl[13] br[13] wl[434] vdd gnd cell_6t
Xbit_r435_c13 bl[13] br[13] wl[435] vdd gnd cell_6t
Xbit_r436_c13 bl[13] br[13] wl[436] vdd gnd cell_6t
Xbit_r437_c13 bl[13] br[13] wl[437] vdd gnd cell_6t
Xbit_r438_c13 bl[13] br[13] wl[438] vdd gnd cell_6t
Xbit_r439_c13 bl[13] br[13] wl[439] vdd gnd cell_6t
Xbit_r440_c13 bl[13] br[13] wl[440] vdd gnd cell_6t
Xbit_r441_c13 bl[13] br[13] wl[441] vdd gnd cell_6t
Xbit_r442_c13 bl[13] br[13] wl[442] vdd gnd cell_6t
Xbit_r443_c13 bl[13] br[13] wl[443] vdd gnd cell_6t
Xbit_r444_c13 bl[13] br[13] wl[444] vdd gnd cell_6t
Xbit_r445_c13 bl[13] br[13] wl[445] vdd gnd cell_6t
Xbit_r446_c13 bl[13] br[13] wl[446] vdd gnd cell_6t
Xbit_r447_c13 bl[13] br[13] wl[447] vdd gnd cell_6t
Xbit_r448_c13 bl[13] br[13] wl[448] vdd gnd cell_6t
Xbit_r449_c13 bl[13] br[13] wl[449] vdd gnd cell_6t
Xbit_r450_c13 bl[13] br[13] wl[450] vdd gnd cell_6t
Xbit_r451_c13 bl[13] br[13] wl[451] vdd gnd cell_6t
Xbit_r452_c13 bl[13] br[13] wl[452] vdd gnd cell_6t
Xbit_r453_c13 bl[13] br[13] wl[453] vdd gnd cell_6t
Xbit_r454_c13 bl[13] br[13] wl[454] vdd gnd cell_6t
Xbit_r455_c13 bl[13] br[13] wl[455] vdd gnd cell_6t
Xbit_r456_c13 bl[13] br[13] wl[456] vdd gnd cell_6t
Xbit_r457_c13 bl[13] br[13] wl[457] vdd gnd cell_6t
Xbit_r458_c13 bl[13] br[13] wl[458] vdd gnd cell_6t
Xbit_r459_c13 bl[13] br[13] wl[459] vdd gnd cell_6t
Xbit_r460_c13 bl[13] br[13] wl[460] vdd gnd cell_6t
Xbit_r461_c13 bl[13] br[13] wl[461] vdd gnd cell_6t
Xbit_r462_c13 bl[13] br[13] wl[462] vdd gnd cell_6t
Xbit_r463_c13 bl[13] br[13] wl[463] vdd gnd cell_6t
Xbit_r464_c13 bl[13] br[13] wl[464] vdd gnd cell_6t
Xbit_r465_c13 bl[13] br[13] wl[465] vdd gnd cell_6t
Xbit_r466_c13 bl[13] br[13] wl[466] vdd gnd cell_6t
Xbit_r467_c13 bl[13] br[13] wl[467] vdd gnd cell_6t
Xbit_r468_c13 bl[13] br[13] wl[468] vdd gnd cell_6t
Xbit_r469_c13 bl[13] br[13] wl[469] vdd gnd cell_6t
Xbit_r470_c13 bl[13] br[13] wl[470] vdd gnd cell_6t
Xbit_r471_c13 bl[13] br[13] wl[471] vdd gnd cell_6t
Xbit_r472_c13 bl[13] br[13] wl[472] vdd gnd cell_6t
Xbit_r473_c13 bl[13] br[13] wl[473] vdd gnd cell_6t
Xbit_r474_c13 bl[13] br[13] wl[474] vdd gnd cell_6t
Xbit_r475_c13 bl[13] br[13] wl[475] vdd gnd cell_6t
Xbit_r476_c13 bl[13] br[13] wl[476] vdd gnd cell_6t
Xbit_r477_c13 bl[13] br[13] wl[477] vdd gnd cell_6t
Xbit_r478_c13 bl[13] br[13] wl[478] vdd gnd cell_6t
Xbit_r479_c13 bl[13] br[13] wl[479] vdd gnd cell_6t
Xbit_r480_c13 bl[13] br[13] wl[480] vdd gnd cell_6t
Xbit_r481_c13 bl[13] br[13] wl[481] vdd gnd cell_6t
Xbit_r482_c13 bl[13] br[13] wl[482] vdd gnd cell_6t
Xbit_r483_c13 bl[13] br[13] wl[483] vdd gnd cell_6t
Xbit_r484_c13 bl[13] br[13] wl[484] vdd gnd cell_6t
Xbit_r485_c13 bl[13] br[13] wl[485] vdd gnd cell_6t
Xbit_r486_c13 bl[13] br[13] wl[486] vdd gnd cell_6t
Xbit_r487_c13 bl[13] br[13] wl[487] vdd gnd cell_6t
Xbit_r488_c13 bl[13] br[13] wl[488] vdd gnd cell_6t
Xbit_r489_c13 bl[13] br[13] wl[489] vdd gnd cell_6t
Xbit_r490_c13 bl[13] br[13] wl[490] vdd gnd cell_6t
Xbit_r491_c13 bl[13] br[13] wl[491] vdd gnd cell_6t
Xbit_r492_c13 bl[13] br[13] wl[492] vdd gnd cell_6t
Xbit_r493_c13 bl[13] br[13] wl[493] vdd gnd cell_6t
Xbit_r494_c13 bl[13] br[13] wl[494] vdd gnd cell_6t
Xbit_r495_c13 bl[13] br[13] wl[495] vdd gnd cell_6t
Xbit_r496_c13 bl[13] br[13] wl[496] vdd gnd cell_6t
Xbit_r497_c13 bl[13] br[13] wl[497] vdd gnd cell_6t
Xbit_r498_c13 bl[13] br[13] wl[498] vdd gnd cell_6t
Xbit_r499_c13 bl[13] br[13] wl[499] vdd gnd cell_6t
Xbit_r500_c13 bl[13] br[13] wl[500] vdd gnd cell_6t
Xbit_r501_c13 bl[13] br[13] wl[501] vdd gnd cell_6t
Xbit_r502_c13 bl[13] br[13] wl[502] vdd gnd cell_6t
Xbit_r503_c13 bl[13] br[13] wl[503] vdd gnd cell_6t
Xbit_r504_c13 bl[13] br[13] wl[504] vdd gnd cell_6t
Xbit_r505_c13 bl[13] br[13] wl[505] vdd gnd cell_6t
Xbit_r506_c13 bl[13] br[13] wl[506] vdd gnd cell_6t
Xbit_r507_c13 bl[13] br[13] wl[507] vdd gnd cell_6t
Xbit_r508_c13 bl[13] br[13] wl[508] vdd gnd cell_6t
Xbit_r509_c13 bl[13] br[13] wl[509] vdd gnd cell_6t
Xbit_r510_c13 bl[13] br[13] wl[510] vdd gnd cell_6t
Xbit_r511_c13 bl[13] br[13] wl[511] vdd gnd cell_6t
Xbit_r0_c14 bl[14] br[14] wl[0] vdd gnd cell_6t
Xbit_r1_c14 bl[14] br[14] wl[1] vdd gnd cell_6t
Xbit_r2_c14 bl[14] br[14] wl[2] vdd gnd cell_6t
Xbit_r3_c14 bl[14] br[14] wl[3] vdd gnd cell_6t
Xbit_r4_c14 bl[14] br[14] wl[4] vdd gnd cell_6t
Xbit_r5_c14 bl[14] br[14] wl[5] vdd gnd cell_6t
Xbit_r6_c14 bl[14] br[14] wl[6] vdd gnd cell_6t
Xbit_r7_c14 bl[14] br[14] wl[7] vdd gnd cell_6t
Xbit_r8_c14 bl[14] br[14] wl[8] vdd gnd cell_6t
Xbit_r9_c14 bl[14] br[14] wl[9] vdd gnd cell_6t
Xbit_r10_c14 bl[14] br[14] wl[10] vdd gnd cell_6t
Xbit_r11_c14 bl[14] br[14] wl[11] vdd gnd cell_6t
Xbit_r12_c14 bl[14] br[14] wl[12] vdd gnd cell_6t
Xbit_r13_c14 bl[14] br[14] wl[13] vdd gnd cell_6t
Xbit_r14_c14 bl[14] br[14] wl[14] vdd gnd cell_6t
Xbit_r15_c14 bl[14] br[14] wl[15] vdd gnd cell_6t
Xbit_r16_c14 bl[14] br[14] wl[16] vdd gnd cell_6t
Xbit_r17_c14 bl[14] br[14] wl[17] vdd gnd cell_6t
Xbit_r18_c14 bl[14] br[14] wl[18] vdd gnd cell_6t
Xbit_r19_c14 bl[14] br[14] wl[19] vdd gnd cell_6t
Xbit_r20_c14 bl[14] br[14] wl[20] vdd gnd cell_6t
Xbit_r21_c14 bl[14] br[14] wl[21] vdd gnd cell_6t
Xbit_r22_c14 bl[14] br[14] wl[22] vdd gnd cell_6t
Xbit_r23_c14 bl[14] br[14] wl[23] vdd gnd cell_6t
Xbit_r24_c14 bl[14] br[14] wl[24] vdd gnd cell_6t
Xbit_r25_c14 bl[14] br[14] wl[25] vdd gnd cell_6t
Xbit_r26_c14 bl[14] br[14] wl[26] vdd gnd cell_6t
Xbit_r27_c14 bl[14] br[14] wl[27] vdd gnd cell_6t
Xbit_r28_c14 bl[14] br[14] wl[28] vdd gnd cell_6t
Xbit_r29_c14 bl[14] br[14] wl[29] vdd gnd cell_6t
Xbit_r30_c14 bl[14] br[14] wl[30] vdd gnd cell_6t
Xbit_r31_c14 bl[14] br[14] wl[31] vdd gnd cell_6t
Xbit_r32_c14 bl[14] br[14] wl[32] vdd gnd cell_6t
Xbit_r33_c14 bl[14] br[14] wl[33] vdd gnd cell_6t
Xbit_r34_c14 bl[14] br[14] wl[34] vdd gnd cell_6t
Xbit_r35_c14 bl[14] br[14] wl[35] vdd gnd cell_6t
Xbit_r36_c14 bl[14] br[14] wl[36] vdd gnd cell_6t
Xbit_r37_c14 bl[14] br[14] wl[37] vdd gnd cell_6t
Xbit_r38_c14 bl[14] br[14] wl[38] vdd gnd cell_6t
Xbit_r39_c14 bl[14] br[14] wl[39] vdd gnd cell_6t
Xbit_r40_c14 bl[14] br[14] wl[40] vdd gnd cell_6t
Xbit_r41_c14 bl[14] br[14] wl[41] vdd gnd cell_6t
Xbit_r42_c14 bl[14] br[14] wl[42] vdd gnd cell_6t
Xbit_r43_c14 bl[14] br[14] wl[43] vdd gnd cell_6t
Xbit_r44_c14 bl[14] br[14] wl[44] vdd gnd cell_6t
Xbit_r45_c14 bl[14] br[14] wl[45] vdd gnd cell_6t
Xbit_r46_c14 bl[14] br[14] wl[46] vdd gnd cell_6t
Xbit_r47_c14 bl[14] br[14] wl[47] vdd gnd cell_6t
Xbit_r48_c14 bl[14] br[14] wl[48] vdd gnd cell_6t
Xbit_r49_c14 bl[14] br[14] wl[49] vdd gnd cell_6t
Xbit_r50_c14 bl[14] br[14] wl[50] vdd gnd cell_6t
Xbit_r51_c14 bl[14] br[14] wl[51] vdd gnd cell_6t
Xbit_r52_c14 bl[14] br[14] wl[52] vdd gnd cell_6t
Xbit_r53_c14 bl[14] br[14] wl[53] vdd gnd cell_6t
Xbit_r54_c14 bl[14] br[14] wl[54] vdd gnd cell_6t
Xbit_r55_c14 bl[14] br[14] wl[55] vdd gnd cell_6t
Xbit_r56_c14 bl[14] br[14] wl[56] vdd gnd cell_6t
Xbit_r57_c14 bl[14] br[14] wl[57] vdd gnd cell_6t
Xbit_r58_c14 bl[14] br[14] wl[58] vdd gnd cell_6t
Xbit_r59_c14 bl[14] br[14] wl[59] vdd gnd cell_6t
Xbit_r60_c14 bl[14] br[14] wl[60] vdd gnd cell_6t
Xbit_r61_c14 bl[14] br[14] wl[61] vdd gnd cell_6t
Xbit_r62_c14 bl[14] br[14] wl[62] vdd gnd cell_6t
Xbit_r63_c14 bl[14] br[14] wl[63] vdd gnd cell_6t
Xbit_r64_c14 bl[14] br[14] wl[64] vdd gnd cell_6t
Xbit_r65_c14 bl[14] br[14] wl[65] vdd gnd cell_6t
Xbit_r66_c14 bl[14] br[14] wl[66] vdd gnd cell_6t
Xbit_r67_c14 bl[14] br[14] wl[67] vdd gnd cell_6t
Xbit_r68_c14 bl[14] br[14] wl[68] vdd gnd cell_6t
Xbit_r69_c14 bl[14] br[14] wl[69] vdd gnd cell_6t
Xbit_r70_c14 bl[14] br[14] wl[70] vdd gnd cell_6t
Xbit_r71_c14 bl[14] br[14] wl[71] vdd gnd cell_6t
Xbit_r72_c14 bl[14] br[14] wl[72] vdd gnd cell_6t
Xbit_r73_c14 bl[14] br[14] wl[73] vdd gnd cell_6t
Xbit_r74_c14 bl[14] br[14] wl[74] vdd gnd cell_6t
Xbit_r75_c14 bl[14] br[14] wl[75] vdd gnd cell_6t
Xbit_r76_c14 bl[14] br[14] wl[76] vdd gnd cell_6t
Xbit_r77_c14 bl[14] br[14] wl[77] vdd gnd cell_6t
Xbit_r78_c14 bl[14] br[14] wl[78] vdd gnd cell_6t
Xbit_r79_c14 bl[14] br[14] wl[79] vdd gnd cell_6t
Xbit_r80_c14 bl[14] br[14] wl[80] vdd gnd cell_6t
Xbit_r81_c14 bl[14] br[14] wl[81] vdd gnd cell_6t
Xbit_r82_c14 bl[14] br[14] wl[82] vdd gnd cell_6t
Xbit_r83_c14 bl[14] br[14] wl[83] vdd gnd cell_6t
Xbit_r84_c14 bl[14] br[14] wl[84] vdd gnd cell_6t
Xbit_r85_c14 bl[14] br[14] wl[85] vdd gnd cell_6t
Xbit_r86_c14 bl[14] br[14] wl[86] vdd gnd cell_6t
Xbit_r87_c14 bl[14] br[14] wl[87] vdd gnd cell_6t
Xbit_r88_c14 bl[14] br[14] wl[88] vdd gnd cell_6t
Xbit_r89_c14 bl[14] br[14] wl[89] vdd gnd cell_6t
Xbit_r90_c14 bl[14] br[14] wl[90] vdd gnd cell_6t
Xbit_r91_c14 bl[14] br[14] wl[91] vdd gnd cell_6t
Xbit_r92_c14 bl[14] br[14] wl[92] vdd gnd cell_6t
Xbit_r93_c14 bl[14] br[14] wl[93] vdd gnd cell_6t
Xbit_r94_c14 bl[14] br[14] wl[94] vdd gnd cell_6t
Xbit_r95_c14 bl[14] br[14] wl[95] vdd gnd cell_6t
Xbit_r96_c14 bl[14] br[14] wl[96] vdd gnd cell_6t
Xbit_r97_c14 bl[14] br[14] wl[97] vdd gnd cell_6t
Xbit_r98_c14 bl[14] br[14] wl[98] vdd gnd cell_6t
Xbit_r99_c14 bl[14] br[14] wl[99] vdd gnd cell_6t
Xbit_r100_c14 bl[14] br[14] wl[100] vdd gnd cell_6t
Xbit_r101_c14 bl[14] br[14] wl[101] vdd gnd cell_6t
Xbit_r102_c14 bl[14] br[14] wl[102] vdd gnd cell_6t
Xbit_r103_c14 bl[14] br[14] wl[103] vdd gnd cell_6t
Xbit_r104_c14 bl[14] br[14] wl[104] vdd gnd cell_6t
Xbit_r105_c14 bl[14] br[14] wl[105] vdd gnd cell_6t
Xbit_r106_c14 bl[14] br[14] wl[106] vdd gnd cell_6t
Xbit_r107_c14 bl[14] br[14] wl[107] vdd gnd cell_6t
Xbit_r108_c14 bl[14] br[14] wl[108] vdd gnd cell_6t
Xbit_r109_c14 bl[14] br[14] wl[109] vdd gnd cell_6t
Xbit_r110_c14 bl[14] br[14] wl[110] vdd gnd cell_6t
Xbit_r111_c14 bl[14] br[14] wl[111] vdd gnd cell_6t
Xbit_r112_c14 bl[14] br[14] wl[112] vdd gnd cell_6t
Xbit_r113_c14 bl[14] br[14] wl[113] vdd gnd cell_6t
Xbit_r114_c14 bl[14] br[14] wl[114] vdd gnd cell_6t
Xbit_r115_c14 bl[14] br[14] wl[115] vdd gnd cell_6t
Xbit_r116_c14 bl[14] br[14] wl[116] vdd gnd cell_6t
Xbit_r117_c14 bl[14] br[14] wl[117] vdd gnd cell_6t
Xbit_r118_c14 bl[14] br[14] wl[118] vdd gnd cell_6t
Xbit_r119_c14 bl[14] br[14] wl[119] vdd gnd cell_6t
Xbit_r120_c14 bl[14] br[14] wl[120] vdd gnd cell_6t
Xbit_r121_c14 bl[14] br[14] wl[121] vdd gnd cell_6t
Xbit_r122_c14 bl[14] br[14] wl[122] vdd gnd cell_6t
Xbit_r123_c14 bl[14] br[14] wl[123] vdd gnd cell_6t
Xbit_r124_c14 bl[14] br[14] wl[124] vdd gnd cell_6t
Xbit_r125_c14 bl[14] br[14] wl[125] vdd gnd cell_6t
Xbit_r126_c14 bl[14] br[14] wl[126] vdd gnd cell_6t
Xbit_r127_c14 bl[14] br[14] wl[127] vdd gnd cell_6t
Xbit_r128_c14 bl[14] br[14] wl[128] vdd gnd cell_6t
Xbit_r129_c14 bl[14] br[14] wl[129] vdd gnd cell_6t
Xbit_r130_c14 bl[14] br[14] wl[130] vdd gnd cell_6t
Xbit_r131_c14 bl[14] br[14] wl[131] vdd gnd cell_6t
Xbit_r132_c14 bl[14] br[14] wl[132] vdd gnd cell_6t
Xbit_r133_c14 bl[14] br[14] wl[133] vdd gnd cell_6t
Xbit_r134_c14 bl[14] br[14] wl[134] vdd gnd cell_6t
Xbit_r135_c14 bl[14] br[14] wl[135] vdd gnd cell_6t
Xbit_r136_c14 bl[14] br[14] wl[136] vdd gnd cell_6t
Xbit_r137_c14 bl[14] br[14] wl[137] vdd gnd cell_6t
Xbit_r138_c14 bl[14] br[14] wl[138] vdd gnd cell_6t
Xbit_r139_c14 bl[14] br[14] wl[139] vdd gnd cell_6t
Xbit_r140_c14 bl[14] br[14] wl[140] vdd gnd cell_6t
Xbit_r141_c14 bl[14] br[14] wl[141] vdd gnd cell_6t
Xbit_r142_c14 bl[14] br[14] wl[142] vdd gnd cell_6t
Xbit_r143_c14 bl[14] br[14] wl[143] vdd gnd cell_6t
Xbit_r144_c14 bl[14] br[14] wl[144] vdd gnd cell_6t
Xbit_r145_c14 bl[14] br[14] wl[145] vdd gnd cell_6t
Xbit_r146_c14 bl[14] br[14] wl[146] vdd gnd cell_6t
Xbit_r147_c14 bl[14] br[14] wl[147] vdd gnd cell_6t
Xbit_r148_c14 bl[14] br[14] wl[148] vdd gnd cell_6t
Xbit_r149_c14 bl[14] br[14] wl[149] vdd gnd cell_6t
Xbit_r150_c14 bl[14] br[14] wl[150] vdd gnd cell_6t
Xbit_r151_c14 bl[14] br[14] wl[151] vdd gnd cell_6t
Xbit_r152_c14 bl[14] br[14] wl[152] vdd gnd cell_6t
Xbit_r153_c14 bl[14] br[14] wl[153] vdd gnd cell_6t
Xbit_r154_c14 bl[14] br[14] wl[154] vdd gnd cell_6t
Xbit_r155_c14 bl[14] br[14] wl[155] vdd gnd cell_6t
Xbit_r156_c14 bl[14] br[14] wl[156] vdd gnd cell_6t
Xbit_r157_c14 bl[14] br[14] wl[157] vdd gnd cell_6t
Xbit_r158_c14 bl[14] br[14] wl[158] vdd gnd cell_6t
Xbit_r159_c14 bl[14] br[14] wl[159] vdd gnd cell_6t
Xbit_r160_c14 bl[14] br[14] wl[160] vdd gnd cell_6t
Xbit_r161_c14 bl[14] br[14] wl[161] vdd gnd cell_6t
Xbit_r162_c14 bl[14] br[14] wl[162] vdd gnd cell_6t
Xbit_r163_c14 bl[14] br[14] wl[163] vdd gnd cell_6t
Xbit_r164_c14 bl[14] br[14] wl[164] vdd gnd cell_6t
Xbit_r165_c14 bl[14] br[14] wl[165] vdd gnd cell_6t
Xbit_r166_c14 bl[14] br[14] wl[166] vdd gnd cell_6t
Xbit_r167_c14 bl[14] br[14] wl[167] vdd gnd cell_6t
Xbit_r168_c14 bl[14] br[14] wl[168] vdd gnd cell_6t
Xbit_r169_c14 bl[14] br[14] wl[169] vdd gnd cell_6t
Xbit_r170_c14 bl[14] br[14] wl[170] vdd gnd cell_6t
Xbit_r171_c14 bl[14] br[14] wl[171] vdd gnd cell_6t
Xbit_r172_c14 bl[14] br[14] wl[172] vdd gnd cell_6t
Xbit_r173_c14 bl[14] br[14] wl[173] vdd gnd cell_6t
Xbit_r174_c14 bl[14] br[14] wl[174] vdd gnd cell_6t
Xbit_r175_c14 bl[14] br[14] wl[175] vdd gnd cell_6t
Xbit_r176_c14 bl[14] br[14] wl[176] vdd gnd cell_6t
Xbit_r177_c14 bl[14] br[14] wl[177] vdd gnd cell_6t
Xbit_r178_c14 bl[14] br[14] wl[178] vdd gnd cell_6t
Xbit_r179_c14 bl[14] br[14] wl[179] vdd gnd cell_6t
Xbit_r180_c14 bl[14] br[14] wl[180] vdd gnd cell_6t
Xbit_r181_c14 bl[14] br[14] wl[181] vdd gnd cell_6t
Xbit_r182_c14 bl[14] br[14] wl[182] vdd gnd cell_6t
Xbit_r183_c14 bl[14] br[14] wl[183] vdd gnd cell_6t
Xbit_r184_c14 bl[14] br[14] wl[184] vdd gnd cell_6t
Xbit_r185_c14 bl[14] br[14] wl[185] vdd gnd cell_6t
Xbit_r186_c14 bl[14] br[14] wl[186] vdd gnd cell_6t
Xbit_r187_c14 bl[14] br[14] wl[187] vdd gnd cell_6t
Xbit_r188_c14 bl[14] br[14] wl[188] vdd gnd cell_6t
Xbit_r189_c14 bl[14] br[14] wl[189] vdd gnd cell_6t
Xbit_r190_c14 bl[14] br[14] wl[190] vdd gnd cell_6t
Xbit_r191_c14 bl[14] br[14] wl[191] vdd gnd cell_6t
Xbit_r192_c14 bl[14] br[14] wl[192] vdd gnd cell_6t
Xbit_r193_c14 bl[14] br[14] wl[193] vdd gnd cell_6t
Xbit_r194_c14 bl[14] br[14] wl[194] vdd gnd cell_6t
Xbit_r195_c14 bl[14] br[14] wl[195] vdd gnd cell_6t
Xbit_r196_c14 bl[14] br[14] wl[196] vdd gnd cell_6t
Xbit_r197_c14 bl[14] br[14] wl[197] vdd gnd cell_6t
Xbit_r198_c14 bl[14] br[14] wl[198] vdd gnd cell_6t
Xbit_r199_c14 bl[14] br[14] wl[199] vdd gnd cell_6t
Xbit_r200_c14 bl[14] br[14] wl[200] vdd gnd cell_6t
Xbit_r201_c14 bl[14] br[14] wl[201] vdd gnd cell_6t
Xbit_r202_c14 bl[14] br[14] wl[202] vdd gnd cell_6t
Xbit_r203_c14 bl[14] br[14] wl[203] vdd gnd cell_6t
Xbit_r204_c14 bl[14] br[14] wl[204] vdd gnd cell_6t
Xbit_r205_c14 bl[14] br[14] wl[205] vdd gnd cell_6t
Xbit_r206_c14 bl[14] br[14] wl[206] vdd gnd cell_6t
Xbit_r207_c14 bl[14] br[14] wl[207] vdd gnd cell_6t
Xbit_r208_c14 bl[14] br[14] wl[208] vdd gnd cell_6t
Xbit_r209_c14 bl[14] br[14] wl[209] vdd gnd cell_6t
Xbit_r210_c14 bl[14] br[14] wl[210] vdd gnd cell_6t
Xbit_r211_c14 bl[14] br[14] wl[211] vdd gnd cell_6t
Xbit_r212_c14 bl[14] br[14] wl[212] vdd gnd cell_6t
Xbit_r213_c14 bl[14] br[14] wl[213] vdd gnd cell_6t
Xbit_r214_c14 bl[14] br[14] wl[214] vdd gnd cell_6t
Xbit_r215_c14 bl[14] br[14] wl[215] vdd gnd cell_6t
Xbit_r216_c14 bl[14] br[14] wl[216] vdd gnd cell_6t
Xbit_r217_c14 bl[14] br[14] wl[217] vdd gnd cell_6t
Xbit_r218_c14 bl[14] br[14] wl[218] vdd gnd cell_6t
Xbit_r219_c14 bl[14] br[14] wl[219] vdd gnd cell_6t
Xbit_r220_c14 bl[14] br[14] wl[220] vdd gnd cell_6t
Xbit_r221_c14 bl[14] br[14] wl[221] vdd gnd cell_6t
Xbit_r222_c14 bl[14] br[14] wl[222] vdd gnd cell_6t
Xbit_r223_c14 bl[14] br[14] wl[223] vdd gnd cell_6t
Xbit_r224_c14 bl[14] br[14] wl[224] vdd gnd cell_6t
Xbit_r225_c14 bl[14] br[14] wl[225] vdd gnd cell_6t
Xbit_r226_c14 bl[14] br[14] wl[226] vdd gnd cell_6t
Xbit_r227_c14 bl[14] br[14] wl[227] vdd gnd cell_6t
Xbit_r228_c14 bl[14] br[14] wl[228] vdd gnd cell_6t
Xbit_r229_c14 bl[14] br[14] wl[229] vdd gnd cell_6t
Xbit_r230_c14 bl[14] br[14] wl[230] vdd gnd cell_6t
Xbit_r231_c14 bl[14] br[14] wl[231] vdd gnd cell_6t
Xbit_r232_c14 bl[14] br[14] wl[232] vdd gnd cell_6t
Xbit_r233_c14 bl[14] br[14] wl[233] vdd gnd cell_6t
Xbit_r234_c14 bl[14] br[14] wl[234] vdd gnd cell_6t
Xbit_r235_c14 bl[14] br[14] wl[235] vdd gnd cell_6t
Xbit_r236_c14 bl[14] br[14] wl[236] vdd gnd cell_6t
Xbit_r237_c14 bl[14] br[14] wl[237] vdd gnd cell_6t
Xbit_r238_c14 bl[14] br[14] wl[238] vdd gnd cell_6t
Xbit_r239_c14 bl[14] br[14] wl[239] vdd gnd cell_6t
Xbit_r240_c14 bl[14] br[14] wl[240] vdd gnd cell_6t
Xbit_r241_c14 bl[14] br[14] wl[241] vdd gnd cell_6t
Xbit_r242_c14 bl[14] br[14] wl[242] vdd gnd cell_6t
Xbit_r243_c14 bl[14] br[14] wl[243] vdd gnd cell_6t
Xbit_r244_c14 bl[14] br[14] wl[244] vdd gnd cell_6t
Xbit_r245_c14 bl[14] br[14] wl[245] vdd gnd cell_6t
Xbit_r246_c14 bl[14] br[14] wl[246] vdd gnd cell_6t
Xbit_r247_c14 bl[14] br[14] wl[247] vdd gnd cell_6t
Xbit_r248_c14 bl[14] br[14] wl[248] vdd gnd cell_6t
Xbit_r249_c14 bl[14] br[14] wl[249] vdd gnd cell_6t
Xbit_r250_c14 bl[14] br[14] wl[250] vdd gnd cell_6t
Xbit_r251_c14 bl[14] br[14] wl[251] vdd gnd cell_6t
Xbit_r252_c14 bl[14] br[14] wl[252] vdd gnd cell_6t
Xbit_r253_c14 bl[14] br[14] wl[253] vdd gnd cell_6t
Xbit_r254_c14 bl[14] br[14] wl[254] vdd gnd cell_6t
Xbit_r255_c14 bl[14] br[14] wl[255] vdd gnd cell_6t
Xbit_r256_c14 bl[14] br[14] wl[256] vdd gnd cell_6t
Xbit_r257_c14 bl[14] br[14] wl[257] vdd gnd cell_6t
Xbit_r258_c14 bl[14] br[14] wl[258] vdd gnd cell_6t
Xbit_r259_c14 bl[14] br[14] wl[259] vdd gnd cell_6t
Xbit_r260_c14 bl[14] br[14] wl[260] vdd gnd cell_6t
Xbit_r261_c14 bl[14] br[14] wl[261] vdd gnd cell_6t
Xbit_r262_c14 bl[14] br[14] wl[262] vdd gnd cell_6t
Xbit_r263_c14 bl[14] br[14] wl[263] vdd gnd cell_6t
Xbit_r264_c14 bl[14] br[14] wl[264] vdd gnd cell_6t
Xbit_r265_c14 bl[14] br[14] wl[265] vdd gnd cell_6t
Xbit_r266_c14 bl[14] br[14] wl[266] vdd gnd cell_6t
Xbit_r267_c14 bl[14] br[14] wl[267] vdd gnd cell_6t
Xbit_r268_c14 bl[14] br[14] wl[268] vdd gnd cell_6t
Xbit_r269_c14 bl[14] br[14] wl[269] vdd gnd cell_6t
Xbit_r270_c14 bl[14] br[14] wl[270] vdd gnd cell_6t
Xbit_r271_c14 bl[14] br[14] wl[271] vdd gnd cell_6t
Xbit_r272_c14 bl[14] br[14] wl[272] vdd gnd cell_6t
Xbit_r273_c14 bl[14] br[14] wl[273] vdd gnd cell_6t
Xbit_r274_c14 bl[14] br[14] wl[274] vdd gnd cell_6t
Xbit_r275_c14 bl[14] br[14] wl[275] vdd gnd cell_6t
Xbit_r276_c14 bl[14] br[14] wl[276] vdd gnd cell_6t
Xbit_r277_c14 bl[14] br[14] wl[277] vdd gnd cell_6t
Xbit_r278_c14 bl[14] br[14] wl[278] vdd gnd cell_6t
Xbit_r279_c14 bl[14] br[14] wl[279] vdd gnd cell_6t
Xbit_r280_c14 bl[14] br[14] wl[280] vdd gnd cell_6t
Xbit_r281_c14 bl[14] br[14] wl[281] vdd gnd cell_6t
Xbit_r282_c14 bl[14] br[14] wl[282] vdd gnd cell_6t
Xbit_r283_c14 bl[14] br[14] wl[283] vdd gnd cell_6t
Xbit_r284_c14 bl[14] br[14] wl[284] vdd gnd cell_6t
Xbit_r285_c14 bl[14] br[14] wl[285] vdd gnd cell_6t
Xbit_r286_c14 bl[14] br[14] wl[286] vdd gnd cell_6t
Xbit_r287_c14 bl[14] br[14] wl[287] vdd gnd cell_6t
Xbit_r288_c14 bl[14] br[14] wl[288] vdd gnd cell_6t
Xbit_r289_c14 bl[14] br[14] wl[289] vdd gnd cell_6t
Xbit_r290_c14 bl[14] br[14] wl[290] vdd gnd cell_6t
Xbit_r291_c14 bl[14] br[14] wl[291] vdd gnd cell_6t
Xbit_r292_c14 bl[14] br[14] wl[292] vdd gnd cell_6t
Xbit_r293_c14 bl[14] br[14] wl[293] vdd gnd cell_6t
Xbit_r294_c14 bl[14] br[14] wl[294] vdd gnd cell_6t
Xbit_r295_c14 bl[14] br[14] wl[295] vdd gnd cell_6t
Xbit_r296_c14 bl[14] br[14] wl[296] vdd gnd cell_6t
Xbit_r297_c14 bl[14] br[14] wl[297] vdd gnd cell_6t
Xbit_r298_c14 bl[14] br[14] wl[298] vdd gnd cell_6t
Xbit_r299_c14 bl[14] br[14] wl[299] vdd gnd cell_6t
Xbit_r300_c14 bl[14] br[14] wl[300] vdd gnd cell_6t
Xbit_r301_c14 bl[14] br[14] wl[301] vdd gnd cell_6t
Xbit_r302_c14 bl[14] br[14] wl[302] vdd gnd cell_6t
Xbit_r303_c14 bl[14] br[14] wl[303] vdd gnd cell_6t
Xbit_r304_c14 bl[14] br[14] wl[304] vdd gnd cell_6t
Xbit_r305_c14 bl[14] br[14] wl[305] vdd gnd cell_6t
Xbit_r306_c14 bl[14] br[14] wl[306] vdd gnd cell_6t
Xbit_r307_c14 bl[14] br[14] wl[307] vdd gnd cell_6t
Xbit_r308_c14 bl[14] br[14] wl[308] vdd gnd cell_6t
Xbit_r309_c14 bl[14] br[14] wl[309] vdd gnd cell_6t
Xbit_r310_c14 bl[14] br[14] wl[310] vdd gnd cell_6t
Xbit_r311_c14 bl[14] br[14] wl[311] vdd gnd cell_6t
Xbit_r312_c14 bl[14] br[14] wl[312] vdd gnd cell_6t
Xbit_r313_c14 bl[14] br[14] wl[313] vdd gnd cell_6t
Xbit_r314_c14 bl[14] br[14] wl[314] vdd gnd cell_6t
Xbit_r315_c14 bl[14] br[14] wl[315] vdd gnd cell_6t
Xbit_r316_c14 bl[14] br[14] wl[316] vdd gnd cell_6t
Xbit_r317_c14 bl[14] br[14] wl[317] vdd gnd cell_6t
Xbit_r318_c14 bl[14] br[14] wl[318] vdd gnd cell_6t
Xbit_r319_c14 bl[14] br[14] wl[319] vdd gnd cell_6t
Xbit_r320_c14 bl[14] br[14] wl[320] vdd gnd cell_6t
Xbit_r321_c14 bl[14] br[14] wl[321] vdd gnd cell_6t
Xbit_r322_c14 bl[14] br[14] wl[322] vdd gnd cell_6t
Xbit_r323_c14 bl[14] br[14] wl[323] vdd gnd cell_6t
Xbit_r324_c14 bl[14] br[14] wl[324] vdd gnd cell_6t
Xbit_r325_c14 bl[14] br[14] wl[325] vdd gnd cell_6t
Xbit_r326_c14 bl[14] br[14] wl[326] vdd gnd cell_6t
Xbit_r327_c14 bl[14] br[14] wl[327] vdd gnd cell_6t
Xbit_r328_c14 bl[14] br[14] wl[328] vdd gnd cell_6t
Xbit_r329_c14 bl[14] br[14] wl[329] vdd gnd cell_6t
Xbit_r330_c14 bl[14] br[14] wl[330] vdd gnd cell_6t
Xbit_r331_c14 bl[14] br[14] wl[331] vdd gnd cell_6t
Xbit_r332_c14 bl[14] br[14] wl[332] vdd gnd cell_6t
Xbit_r333_c14 bl[14] br[14] wl[333] vdd gnd cell_6t
Xbit_r334_c14 bl[14] br[14] wl[334] vdd gnd cell_6t
Xbit_r335_c14 bl[14] br[14] wl[335] vdd gnd cell_6t
Xbit_r336_c14 bl[14] br[14] wl[336] vdd gnd cell_6t
Xbit_r337_c14 bl[14] br[14] wl[337] vdd gnd cell_6t
Xbit_r338_c14 bl[14] br[14] wl[338] vdd gnd cell_6t
Xbit_r339_c14 bl[14] br[14] wl[339] vdd gnd cell_6t
Xbit_r340_c14 bl[14] br[14] wl[340] vdd gnd cell_6t
Xbit_r341_c14 bl[14] br[14] wl[341] vdd gnd cell_6t
Xbit_r342_c14 bl[14] br[14] wl[342] vdd gnd cell_6t
Xbit_r343_c14 bl[14] br[14] wl[343] vdd gnd cell_6t
Xbit_r344_c14 bl[14] br[14] wl[344] vdd gnd cell_6t
Xbit_r345_c14 bl[14] br[14] wl[345] vdd gnd cell_6t
Xbit_r346_c14 bl[14] br[14] wl[346] vdd gnd cell_6t
Xbit_r347_c14 bl[14] br[14] wl[347] vdd gnd cell_6t
Xbit_r348_c14 bl[14] br[14] wl[348] vdd gnd cell_6t
Xbit_r349_c14 bl[14] br[14] wl[349] vdd gnd cell_6t
Xbit_r350_c14 bl[14] br[14] wl[350] vdd gnd cell_6t
Xbit_r351_c14 bl[14] br[14] wl[351] vdd gnd cell_6t
Xbit_r352_c14 bl[14] br[14] wl[352] vdd gnd cell_6t
Xbit_r353_c14 bl[14] br[14] wl[353] vdd gnd cell_6t
Xbit_r354_c14 bl[14] br[14] wl[354] vdd gnd cell_6t
Xbit_r355_c14 bl[14] br[14] wl[355] vdd gnd cell_6t
Xbit_r356_c14 bl[14] br[14] wl[356] vdd gnd cell_6t
Xbit_r357_c14 bl[14] br[14] wl[357] vdd gnd cell_6t
Xbit_r358_c14 bl[14] br[14] wl[358] vdd gnd cell_6t
Xbit_r359_c14 bl[14] br[14] wl[359] vdd gnd cell_6t
Xbit_r360_c14 bl[14] br[14] wl[360] vdd gnd cell_6t
Xbit_r361_c14 bl[14] br[14] wl[361] vdd gnd cell_6t
Xbit_r362_c14 bl[14] br[14] wl[362] vdd gnd cell_6t
Xbit_r363_c14 bl[14] br[14] wl[363] vdd gnd cell_6t
Xbit_r364_c14 bl[14] br[14] wl[364] vdd gnd cell_6t
Xbit_r365_c14 bl[14] br[14] wl[365] vdd gnd cell_6t
Xbit_r366_c14 bl[14] br[14] wl[366] vdd gnd cell_6t
Xbit_r367_c14 bl[14] br[14] wl[367] vdd gnd cell_6t
Xbit_r368_c14 bl[14] br[14] wl[368] vdd gnd cell_6t
Xbit_r369_c14 bl[14] br[14] wl[369] vdd gnd cell_6t
Xbit_r370_c14 bl[14] br[14] wl[370] vdd gnd cell_6t
Xbit_r371_c14 bl[14] br[14] wl[371] vdd gnd cell_6t
Xbit_r372_c14 bl[14] br[14] wl[372] vdd gnd cell_6t
Xbit_r373_c14 bl[14] br[14] wl[373] vdd gnd cell_6t
Xbit_r374_c14 bl[14] br[14] wl[374] vdd gnd cell_6t
Xbit_r375_c14 bl[14] br[14] wl[375] vdd gnd cell_6t
Xbit_r376_c14 bl[14] br[14] wl[376] vdd gnd cell_6t
Xbit_r377_c14 bl[14] br[14] wl[377] vdd gnd cell_6t
Xbit_r378_c14 bl[14] br[14] wl[378] vdd gnd cell_6t
Xbit_r379_c14 bl[14] br[14] wl[379] vdd gnd cell_6t
Xbit_r380_c14 bl[14] br[14] wl[380] vdd gnd cell_6t
Xbit_r381_c14 bl[14] br[14] wl[381] vdd gnd cell_6t
Xbit_r382_c14 bl[14] br[14] wl[382] vdd gnd cell_6t
Xbit_r383_c14 bl[14] br[14] wl[383] vdd gnd cell_6t
Xbit_r384_c14 bl[14] br[14] wl[384] vdd gnd cell_6t
Xbit_r385_c14 bl[14] br[14] wl[385] vdd gnd cell_6t
Xbit_r386_c14 bl[14] br[14] wl[386] vdd gnd cell_6t
Xbit_r387_c14 bl[14] br[14] wl[387] vdd gnd cell_6t
Xbit_r388_c14 bl[14] br[14] wl[388] vdd gnd cell_6t
Xbit_r389_c14 bl[14] br[14] wl[389] vdd gnd cell_6t
Xbit_r390_c14 bl[14] br[14] wl[390] vdd gnd cell_6t
Xbit_r391_c14 bl[14] br[14] wl[391] vdd gnd cell_6t
Xbit_r392_c14 bl[14] br[14] wl[392] vdd gnd cell_6t
Xbit_r393_c14 bl[14] br[14] wl[393] vdd gnd cell_6t
Xbit_r394_c14 bl[14] br[14] wl[394] vdd gnd cell_6t
Xbit_r395_c14 bl[14] br[14] wl[395] vdd gnd cell_6t
Xbit_r396_c14 bl[14] br[14] wl[396] vdd gnd cell_6t
Xbit_r397_c14 bl[14] br[14] wl[397] vdd gnd cell_6t
Xbit_r398_c14 bl[14] br[14] wl[398] vdd gnd cell_6t
Xbit_r399_c14 bl[14] br[14] wl[399] vdd gnd cell_6t
Xbit_r400_c14 bl[14] br[14] wl[400] vdd gnd cell_6t
Xbit_r401_c14 bl[14] br[14] wl[401] vdd gnd cell_6t
Xbit_r402_c14 bl[14] br[14] wl[402] vdd gnd cell_6t
Xbit_r403_c14 bl[14] br[14] wl[403] vdd gnd cell_6t
Xbit_r404_c14 bl[14] br[14] wl[404] vdd gnd cell_6t
Xbit_r405_c14 bl[14] br[14] wl[405] vdd gnd cell_6t
Xbit_r406_c14 bl[14] br[14] wl[406] vdd gnd cell_6t
Xbit_r407_c14 bl[14] br[14] wl[407] vdd gnd cell_6t
Xbit_r408_c14 bl[14] br[14] wl[408] vdd gnd cell_6t
Xbit_r409_c14 bl[14] br[14] wl[409] vdd gnd cell_6t
Xbit_r410_c14 bl[14] br[14] wl[410] vdd gnd cell_6t
Xbit_r411_c14 bl[14] br[14] wl[411] vdd gnd cell_6t
Xbit_r412_c14 bl[14] br[14] wl[412] vdd gnd cell_6t
Xbit_r413_c14 bl[14] br[14] wl[413] vdd gnd cell_6t
Xbit_r414_c14 bl[14] br[14] wl[414] vdd gnd cell_6t
Xbit_r415_c14 bl[14] br[14] wl[415] vdd gnd cell_6t
Xbit_r416_c14 bl[14] br[14] wl[416] vdd gnd cell_6t
Xbit_r417_c14 bl[14] br[14] wl[417] vdd gnd cell_6t
Xbit_r418_c14 bl[14] br[14] wl[418] vdd gnd cell_6t
Xbit_r419_c14 bl[14] br[14] wl[419] vdd gnd cell_6t
Xbit_r420_c14 bl[14] br[14] wl[420] vdd gnd cell_6t
Xbit_r421_c14 bl[14] br[14] wl[421] vdd gnd cell_6t
Xbit_r422_c14 bl[14] br[14] wl[422] vdd gnd cell_6t
Xbit_r423_c14 bl[14] br[14] wl[423] vdd gnd cell_6t
Xbit_r424_c14 bl[14] br[14] wl[424] vdd gnd cell_6t
Xbit_r425_c14 bl[14] br[14] wl[425] vdd gnd cell_6t
Xbit_r426_c14 bl[14] br[14] wl[426] vdd gnd cell_6t
Xbit_r427_c14 bl[14] br[14] wl[427] vdd gnd cell_6t
Xbit_r428_c14 bl[14] br[14] wl[428] vdd gnd cell_6t
Xbit_r429_c14 bl[14] br[14] wl[429] vdd gnd cell_6t
Xbit_r430_c14 bl[14] br[14] wl[430] vdd gnd cell_6t
Xbit_r431_c14 bl[14] br[14] wl[431] vdd gnd cell_6t
Xbit_r432_c14 bl[14] br[14] wl[432] vdd gnd cell_6t
Xbit_r433_c14 bl[14] br[14] wl[433] vdd gnd cell_6t
Xbit_r434_c14 bl[14] br[14] wl[434] vdd gnd cell_6t
Xbit_r435_c14 bl[14] br[14] wl[435] vdd gnd cell_6t
Xbit_r436_c14 bl[14] br[14] wl[436] vdd gnd cell_6t
Xbit_r437_c14 bl[14] br[14] wl[437] vdd gnd cell_6t
Xbit_r438_c14 bl[14] br[14] wl[438] vdd gnd cell_6t
Xbit_r439_c14 bl[14] br[14] wl[439] vdd gnd cell_6t
Xbit_r440_c14 bl[14] br[14] wl[440] vdd gnd cell_6t
Xbit_r441_c14 bl[14] br[14] wl[441] vdd gnd cell_6t
Xbit_r442_c14 bl[14] br[14] wl[442] vdd gnd cell_6t
Xbit_r443_c14 bl[14] br[14] wl[443] vdd gnd cell_6t
Xbit_r444_c14 bl[14] br[14] wl[444] vdd gnd cell_6t
Xbit_r445_c14 bl[14] br[14] wl[445] vdd gnd cell_6t
Xbit_r446_c14 bl[14] br[14] wl[446] vdd gnd cell_6t
Xbit_r447_c14 bl[14] br[14] wl[447] vdd gnd cell_6t
Xbit_r448_c14 bl[14] br[14] wl[448] vdd gnd cell_6t
Xbit_r449_c14 bl[14] br[14] wl[449] vdd gnd cell_6t
Xbit_r450_c14 bl[14] br[14] wl[450] vdd gnd cell_6t
Xbit_r451_c14 bl[14] br[14] wl[451] vdd gnd cell_6t
Xbit_r452_c14 bl[14] br[14] wl[452] vdd gnd cell_6t
Xbit_r453_c14 bl[14] br[14] wl[453] vdd gnd cell_6t
Xbit_r454_c14 bl[14] br[14] wl[454] vdd gnd cell_6t
Xbit_r455_c14 bl[14] br[14] wl[455] vdd gnd cell_6t
Xbit_r456_c14 bl[14] br[14] wl[456] vdd gnd cell_6t
Xbit_r457_c14 bl[14] br[14] wl[457] vdd gnd cell_6t
Xbit_r458_c14 bl[14] br[14] wl[458] vdd gnd cell_6t
Xbit_r459_c14 bl[14] br[14] wl[459] vdd gnd cell_6t
Xbit_r460_c14 bl[14] br[14] wl[460] vdd gnd cell_6t
Xbit_r461_c14 bl[14] br[14] wl[461] vdd gnd cell_6t
Xbit_r462_c14 bl[14] br[14] wl[462] vdd gnd cell_6t
Xbit_r463_c14 bl[14] br[14] wl[463] vdd gnd cell_6t
Xbit_r464_c14 bl[14] br[14] wl[464] vdd gnd cell_6t
Xbit_r465_c14 bl[14] br[14] wl[465] vdd gnd cell_6t
Xbit_r466_c14 bl[14] br[14] wl[466] vdd gnd cell_6t
Xbit_r467_c14 bl[14] br[14] wl[467] vdd gnd cell_6t
Xbit_r468_c14 bl[14] br[14] wl[468] vdd gnd cell_6t
Xbit_r469_c14 bl[14] br[14] wl[469] vdd gnd cell_6t
Xbit_r470_c14 bl[14] br[14] wl[470] vdd gnd cell_6t
Xbit_r471_c14 bl[14] br[14] wl[471] vdd gnd cell_6t
Xbit_r472_c14 bl[14] br[14] wl[472] vdd gnd cell_6t
Xbit_r473_c14 bl[14] br[14] wl[473] vdd gnd cell_6t
Xbit_r474_c14 bl[14] br[14] wl[474] vdd gnd cell_6t
Xbit_r475_c14 bl[14] br[14] wl[475] vdd gnd cell_6t
Xbit_r476_c14 bl[14] br[14] wl[476] vdd gnd cell_6t
Xbit_r477_c14 bl[14] br[14] wl[477] vdd gnd cell_6t
Xbit_r478_c14 bl[14] br[14] wl[478] vdd gnd cell_6t
Xbit_r479_c14 bl[14] br[14] wl[479] vdd gnd cell_6t
Xbit_r480_c14 bl[14] br[14] wl[480] vdd gnd cell_6t
Xbit_r481_c14 bl[14] br[14] wl[481] vdd gnd cell_6t
Xbit_r482_c14 bl[14] br[14] wl[482] vdd gnd cell_6t
Xbit_r483_c14 bl[14] br[14] wl[483] vdd gnd cell_6t
Xbit_r484_c14 bl[14] br[14] wl[484] vdd gnd cell_6t
Xbit_r485_c14 bl[14] br[14] wl[485] vdd gnd cell_6t
Xbit_r486_c14 bl[14] br[14] wl[486] vdd gnd cell_6t
Xbit_r487_c14 bl[14] br[14] wl[487] vdd gnd cell_6t
Xbit_r488_c14 bl[14] br[14] wl[488] vdd gnd cell_6t
Xbit_r489_c14 bl[14] br[14] wl[489] vdd gnd cell_6t
Xbit_r490_c14 bl[14] br[14] wl[490] vdd gnd cell_6t
Xbit_r491_c14 bl[14] br[14] wl[491] vdd gnd cell_6t
Xbit_r492_c14 bl[14] br[14] wl[492] vdd gnd cell_6t
Xbit_r493_c14 bl[14] br[14] wl[493] vdd gnd cell_6t
Xbit_r494_c14 bl[14] br[14] wl[494] vdd gnd cell_6t
Xbit_r495_c14 bl[14] br[14] wl[495] vdd gnd cell_6t
Xbit_r496_c14 bl[14] br[14] wl[496] vdd gnd cell_6t
Xbit_r497_c14 bl[14] br[14] wl[497] vdd gnd cell_6t
Xbit_r498_c14 bl[14] br[14] wl[498] vdd gnd cell_6t
Xbit_r499_c14 bl[14] br[14] wl[499] vdd gnd cell_6t
Xbit_r500_c14 bl[14] br[14] wl[500] vdd gnd cell_6t
Xbit_r501_c14 bl[14] br[14] wl[501] vdd gnd cell_6t
Xbit_r502_c14 bl[14] br[14] wl[502] vdd gnd cell_6t
Xbit_r503_c14 bl[14] br[14] wl[503] vdd gnd cell_6t
Xbit_r504_c14 bl[14] br[14] wl[504] vdd gnd cell_6t
Xbit_r505_c14 bl[14] br[14] wl[505] vdd gnd cell_6t
Xbit_r506_c14 bl[14] br[14] wl[506] vdd gnd cell_6t
Xbit_r507_c14 bl[14] br[14] wl[507] vdd gnd cell_6t
Xbit_r508_c14 bl[14] br[14] wl[508] vdd gnd cell_6t
Xbit_r509_c14 bl[14] br[14] wl[509] vdd gnd cell_6t
Xbit_r510_c14 bl[14] br[14] wl[510] vdd gnd cell_6t
Xbit_r511_c14 bl[14] br[14] wl[511] vdd gnd cell_6t
Xbit_r0_c15 bl[15] br[15] wl[0] vdd gnd cell_6t
Xbit_r1_c15 bl[15] br[15] wl[1] vdd gnd cell_6t
Xbit_r2_c15 bl[15] br[15] wl[2] vdd gnd cell_6t
Xbit_r3_c15 bl[15] br[15] wl[3] vdd gnd cell_6t
Xbit_r4_c15 bl[15] br[15] wl[4] vdd gnd cell_6t
Xbit_r5_c15 bl[15] br[15] wl[5] vdd gnd cell_6t
Xbit_r6_c15 bl[15] br[15] wl[6] vdd gnd cell_6t
Xbit_r7_c15 bl[15] br[15] wl[7] vdd gnd cell_6t
Xbit_r8_c15 bl[15] br[15] wl[8] vdd gnd cell_6t
Xbit_r9_c15 bl[15] br[15] wl[9] vdd gnd cell_6t
Xbit_r10_c15 bl[15] br[15] wl[10] vdd gnd cell_6t
Xbit_r11_c15 bl[15] br[15] wl[11] vdd gnd cell_6t
Xbit_r12_c15 bl[15] br[15] wl[12] vdd gnd cell_6t
Xbit_r13_c15 bl[15] br[15] wl[13] vdd gnd cell_6t
Xbit_r14_c15 bl[15] br[15] wl[14] vdd gnd cell_6t
Xbit_r15_c15 bl[15] br[15] wl[15] vdd gnd cell_6t
Xbit_r16_c15 bl[15] br[15] wl[16] vdd gnd cell_6t
Xbit_r17_c15 bl[15] br[15] wl[17] vdd gnd cell_6t
Xbit_r18_c15 bl[15] br[15] wl[18] vdd gnd cell_6t
Xbit_r19_c15 bl[15] br[15] wl[19] vdd gnd cell_6t
Xbit_r20_c15 bl[15] br[15] wl[20] vdd gnd cell_6t
Xbit_r21_c15 bl[15] br[15] wl[21] vdd gnd cell_6t
Xbit_r22_c15 bl[15] br[15] wl[22] vdd gnd cell_6t
Xbit_r23_c15 bl[15] br[15] wl[23] vdd gnd cell_6t
Xbit_r24_c15 bl[15] br[15] wl[24] vdd gnd cell_6t
Xbit_r25_c15 bl[15] br[15] wl[25] vdd gnd cell_6t
Xbit_r26_c15 bl[15] br[15] wl[26] vdd gnd cell_6t
Xbit_r27_c15 bl[15] br[15] wl[27] vdd gnd cell_6t
Xbit_r28_c15 bl[15] br[15] wl[28] vdd gnd cell_6t
Xbit_r29_c15 bl[15] br[15] wl[29] vdd gnd cell_6t
Xbit_r30_c15 bl[15] br[15] wl[30] vdd gnd cell_6t
Xbit_r31_c15 bl[15] br[15] wl[31] vdd gnd cell_6t
Xbit_r32_c15 bl[15] br[15] wl[32] vdd gnd cell_6t
Xbit_r33_c15 bl[15] br[15] wl[33] vdd gnd cell_6t
Xbit_r34_c15 bl[15] br[15] wl[34] vdd gnd cell_6t
Xbit_r35_c15 bl[15] br[15] wl[35] vdd gnd cell_6t
Xbit_r36_c15 bl[15] br[15] wl[36] vdd gnd cell_6t
Xbit_r37_c15 bl[15] br[15] wl[37] vdd gnd cell_6t
Xbit_r38_c15 bl[15] br[15] wl[38] vdd gnd cell_6t
Xbit_r39_c15 bl[15] br[15] wl[39] vdd gnd cell_6t
Xbit_r40_c15 bl[15] br[15] wl[40] vdd gnd cell_6t
Xbit_r41_c15 bl[15] br[15] wl[41] vdd gnd cell_6t
Xbit_r42_c15 bl[15] br[15] wl[42] vdd gnd cell_6t
Xbit_r43_c15 bl[15] br[15] wl[43] vdd gnd cell_6t
Xbit_r44_c15 bl[15] br[15] wl[44] vdd gnd cell_6t
Xbit_r45_c15 bl[15] br[15] wl[45] vdd gnd cell_6t
Xbit_r46_c15 bl[15] br[15] wl[46] vdd gnd cell_6t
Xbit_r47_c15 bl[15] br[15] wl[47] vdd gnd cell_6t
Xbit_r48_c15 bl[15] br[15] wl[48] vdd gnd cell_6t
Xbit_r49_c15 bl[15] br[15] wl[49] vdd gnd cell_6t
Xbit_r50_c15 bl[15] br[15] wl[50] vdd gnd cell_6t
Xbit_r51_c15 bl[15] br[15] wl[51] vdd gnd cell_6t
Xbit_r52_c15 bl[15] br[15] wl[52] vdd gnd cell_6t
Xbit_r53_c15 bl[15] br[15] wl[53] vdd gnd cell_6t
Xbit_r54_c15 bl[15] br[15] wl[54] vdd gnd cell_6t
Xbit_r55_c15 bl[15] br[15] wl[55] vdd gnd cell_6t
Xbit_r56_c15 bl[15] br[15] wl[56] vdd gnd cell_6t
Xbit_r57_c15 bl[15] br[15] wl[57] vdd gnd cell_6t
Xbit_r58_c15 bl[15] br[15] wl[58] vdd gnd cell_6t
Xbit_r59_c15 bl[15] br[15] wl[59] vdd gnd cell_6t
Xbit_r60_c15 bl[15] br[15] wl[60] vdd gnd cell_6t
Xbit_r61_c15 bl[15] br[15] wl[61] vdd gnd cell_6t
Xbit_r62_c15 bl[15] br[15] wl[62] vdd gnd cell_6t
Xbit_r63_c15 bl[15] br[15] wl[63] vdd gnd cell_6t
Xbit_r64_c15 bl[15] br[15] wl[64] vdd gnd cell_6t
Xbit_r65_c15 bl[15] br[15] wl[65] vdd gnd cell_6t
Xbit_r66_c15 bl[15] br[15] wl[66] vdd gnd cell_6t
Xbit_r67_c15 bl[15] br[15] wl[67] vdd gnd cell_6t
Xbit_r68_c15 bl[15] br[15] wl[68] vdd gnd cell_6t
Xbit_r69_c15 bl[15] br[15] wl[69] vdd gnd cell_6t
Xbit_r70_c15 bl[15] br[15] wl[70] vdd gnd cell_6t
Xbit_r71_c15 bl[15] br[15] wl[71] vdd gnd cell_6t
Xbit_r72_c15 bl[15] br[15] wl[72] vdd gnd cell_6t
Xbit_r73_c15 bl[15] br[15] wl[73] vdd gnd cell_6t
Xbit_r74_c15 bl[15] br[15] wl[74] vdd gnd cell_6t
Xbit_r75_c15 bl[15] br[15] wl[75] vdd gnd cell_6t
Xbit_r76_c15 bl[15] br[15] wl[76] vdd gnd cell_6t
Xbit_r77_c15 bl[15] br[15] wl[77] vdd gnd cell_6t
Xbit_r78_c15 bl[15] br[15] wl[78] vdd gnd cell_6t
Xbit_r79_c15 bl[15] br[15] wl[79] vdd gnd cell_6t
Xbit_r80_c15 bl[15] br[15] wl[80] vdd gnd cell_6t
Xbit_r81_c15 bl[15] br[15] wl[81] vdd gnd cell_6t
Xbit_r82_c15 bl[15] br[15] wl[82] vdd gnd cell_6t
Xbit_r83_c15 bl[15] br[15] wl[83] vdd gnd cell_6t
Xbit_r84_c15 bl[15] br[15] wl[84] vdd gnd cell_6t
Xbit_r85_c15 bl[15] br[15] wl[85] vdd gnd cell_6t
Xbit_r86_c15 bl[15] br[15] wl[86] vdd gnd cell_6t
Xbit_r87_c15 bl[15] br[15] wl[87] vdd gnd cell_6t
Xbit_r88_c15 bl[15] br[15] wl[88] vdd gnd cell_6t
Xbit_r89_c15 bl[15] br[15] wl[89] vdd gnd cell_6t
Xbit_r90_c15 bl[15] br[15] wl[90] vdd gnd cell_6t
Xbit_r91_c15 bl[15] br[15] wl[91] vdd gnd cell_6t
Xbit_r92_c15 bl[15] br[15] wl[92] vdd gnd cell_6t
Xbit_r93_c15 bl[15] br[15] wl[93] vdd gnd cell_6t
Xbit_r94_c15 bl[15] br[15] wl[94] vdd gnd cell_6t
Xbit_r95_c15 bl[15] br[15] wl[95] vdd gnd cell_6t
Xbit_r96_c15 bl[15] br[15] wl[96] vdd gnd cell_6t
Xbit_r97_c15 bl[15] br[15] wl[97] vdd gnd cell_6t
Xbit_r98_c15 bl[15] br[15] wl[98] vdd gnd cell_6t
Xbit_r99_c15 bl[15] br[15] wl[99] vdd gnd cell_6t
Xbit_r100_c15 bl[15] br[15] wl[100] vdd gnd cell_6t
Xbit_r101_c15 bl[15] br[15] wl[101] vdd gnd cell_6t
Xbit_r102_c15 bl[15] br[15] wl[102] vdd gnd cell_6t
Xbit_r103_c15 bl[15] br[15] wl[103] vdd gnd cell_6t
Xbit_r104_c15 bl[15] br[15] wl[104] vdd gnd cell_6t
Xbit_r105_c15 bl[15] br[15] wl[105] vdd gnd cell_6t
Xbit_r106_c15 bl[15] br[15] wl[106] vdd gnd cell_6t
Xbit_r107_c15 bl[15] br[15] wl[107] vdd gnd cell_6t
Xbit_r108_c15 bl[15] br[15] wl[108] vdd gnd cell_6t
Xbit_r109_c15 bl[15] br[15] wl[109] vdd gnd cell_6t
Xbit_r110_c15 bl[15] br[15] wl[110] vdd gnd cell_6t
Xbit_r111_c15 bl[15] br[15] wl[111] vdd gnd cell_6t
Xbit_r112_c15 bl[15] br[15] wl[112] vdd gnd cell_6t
Xbit_r113_c15 bl[15] br[15] wl[113] vdd gnd cell_6t
Xbit_r114_c15 bl[15] br[15] wl[114] vdd gnd cell_6t
Xbit_r115_c15 bl[15] br[15] wl[115] vdd gnd cell_6t
Xbit_r116_c15 bl[15] br[15] wl[116] vdd gnd cell_6t
Xbit_r117_c15 bl[15] br[15] wl[117] vdd gnd cell_6t
Xbit_r118_c15 bl[15] br[15] wl[118] vdd gnd cell_6t
Xbit_r119_c15 bl[15] br[15] wl[119] vdd gnd cell_6t
Xbit_r120_c15 bl[15] br[15] wl[120] vdd gnd cell_6t
Xbit_r121_c15 bl[15] br[15] wl[121] vdd gnd cell_6t
Xbit_r122_c15 bl[15] br[15] wl[122] vdd gnd cell_6t
Xbit_r123_c15 bl[15] br[15] wl[123] vdd gnd cell_6t
Xbit_r124_c15 bl[15] br[15] wl[124] vdd gnd cell_6t
Xbit_r125_c15 bl[15] br[15] wl[125] vdd gnd cell_6t
Xbit_r126_c15 bl[15] br[15] wl[126] vdd gnd cell_6t
Xbit_r127_c15 bl[15] br[15] wl[127] vdd gnd cell_6t
Xbit_r128_c15 bl[15] br[15] wl[128] vdd gnd cell_6t
Xbit_r129_c15 bl[15] br[15] wl[129] vdd gnd cell_6t
Xbit_r130_c15 bl[15] br[15] wl[130] vdd gnd cell_6t
Xbit_r131_c15 bl[15] br[15] wl[131] vdd gnd cell_6t
Xbit_r132_c15 bl[15] br[15] wl[132] vdd gnd cell_6t
Xbit_r133_c15 bl[15] br[15] wl[133] vdd gnd cell_6t
Xbit_r134_c15 bl[15] br[15] wl[134] vdd gnd cell_6t
Xbit_r135_c15 bl[15] br[15] wl[135] vdd gnd cell_6t
Xbit_r136_c15 bl[15] br[15] wl[136] vdd gnd cell_6t
Xbit_r137_c15 bl[15] br[15] wl[137] vdd gnd cell_6t
Xbit_r138_c15 bl[15] br[15] wl[138] vdd gnd cell_6t
Xbit_r139_c15 bl[15] br[15] wl[139] vdd gnd cell_6t
Xbit_r140_c15 bl[15] br[15] wl[140] vdd gnd cell_6t
Xbit_r141_c15 bl[15] br[15] wl[141] vdd gnd cell_6t
Xbit_r142_c15 bl[15] br[15] wl[142] vdd gnd cell_6t
Xbit_r143_c15 bl[15] br[15] wl[143] vdd gnd cell_6t
Xbit_r144_c15 bl[15] br[15] wl[144] vdd gnd cell_6t
Xbit_r145_c15 bl[15] br[15] wl[145] vdd gnd cell_6t
Xbit_r146_c15 bl[15] br[15] wl[146] vdd gnd cell_6t
Xbit_r147_c15 bl[15] br[15] wl[147] vdd gnd cell_6t
Xbit_r148_c15 bl[15] br[15] wl[148] vdd gnd cell_6t
Xbit_r149_c15 bl[15] br[15] wl[149] vdd gnd cell_6t
Xbit_r150_c15 bl[15] br[15] wl[150] vdd gnd cell_6t
Xbit_r151_c15 bl[15] br[15] wl[151] vdd gnd cell_6t
Xbit_r152_c15 bl[15] br[15] wl[152] vdd gnd cell_6t
Xbit_r153_c15 bl[15] br[15] wl[153] vdd gnd cell_6t
Xbit_r154_c15 bl[15] br[15] wl[154] vdd gnd cell_6t
Xbit_r155_c15 bl[15] br[15] wl[155] vdd gnd cell_6t
Xbit_r156_c15 bl[15] br[15] wl[156] vdd gnd cell_6t
Xbit_r157_c15 bl[15] br[15] wl[157] vdd gnd cell_6t
Xbit_r158_c15 bl[15] br[15] wl[158] vdd gnd cell_6t
Xbit_r159_c15 bl[15] br[15] wl[159] vdd gnd cell_6t
Xbit_r160_c15 bl[15] br[15] wl[160] vdd gnd cell_6t
Xbit_r161_c15 bl[15] br[15] wl[161] vdd gnd cell_6t
Xbit_r162_c15 bl[15] br[15] wl[162] vdd gnd cell_6t
Xbit_r163_c15 bl[15] br[15] wl[163] vdd gnd cell_6t
Xbit_r164_c15 bl[15] br[15] wl[164] vdd gnd cell_6t
Xbit_r165_c15 bl[15] br[15] wl[165] vdd gnd cell_6t
Xbit_r166_c15 bl[15] br[15] wl[166] vdd gnd cell_6t
Xbit_r167_c15 bl[15] br[15] wl[167] vdd gnd cell_6t
Xbit_r168_c15 bl[15] br[15] wl[168] vdd gnd cell_6t
Xbit_r169_c15 bl[15] br[15] wl[169] vdd gnd cell_6t
Xbit_r170_c15 bl[15] br[15] wl[170] vdd gnd cell_6t
Xbit_r171_c15 bl[15] br[15] wl[171] vdd gnd cell_6t
Xbit_r172_c15 bl[15] br[15] wl[172] vdd gnd cell_6t
Xbit_r173_c15 bl[15] br[15] wl[173] vdd gnd cell_6t
Xbit_r174_c15 bl[15] br[15] wl[174] vdd gnd cell_6t
Xbit_r175_c15 bl[15] br[15] wl[175] vdd gnd cell_6t
Xbit_r176_c15 bl[15] br[15] wl[176] vdd gnd cell_6t
Xbit_r177_c15 bl[15] br[15] wl[177] vdd gnd cell_6t
Xbit_r178_c15 bl[15] br[15] wl[178] vdd gnd cell_6t
Xbit_r179_c15 bl[15] br[15] wl[179] vdd gnd cell_6t
Xbit_r180_c15 bl[15] br[15] wl[180] vdd gnd cell_6t
Xbit_r181_c15 bl[15] br[15] wl[181] vdd gnd cell_6t
Xbit_r182_c15 bl[15] br[15] wl[182] vdd gnd cell_6t
Xbit_r183_c15 bl[15] br[15] wl[183] vdd gnd cell_6t
Xbit_r184_c15 bl[15] br[15] wl[184] vdd gnd cell_6t
Xbit_r185_c15 bl[15] br[15] wl[185] vdd gnd cell_6t
Xbit_r186_c15 bl[15] br[15] wl[186] vdd gnd cell_6t
Xbit_r187_c15 bl[15] br[15] wl[187] vdd gnd cell_6t
Xbit_r188_c15 bl[15] br[15] wl[188] vdd gnd cell_6t
Xbit_r189_c15 bl[15] br[15] wl[189] vdd gnd cell_6t
Xbit_r190_c15 bl[15] br[15] wl[190] vdd gnd cell_6t
Xbit_r191_c15 bl[15] br[15] wl[191] vdd gnd cell_6t
Xbit_r192_c15 bl[15] br[15] wl[192] vdd gnd cell_6t
Xbit_r193_c15 bl[15] br[15] wl[193] vdd gnd cell_6t
Xbit_r194_c15 bl[15] br[15] wl[194] vdd gnd cell_6t
Xbit_r195_c15 bl[15] br[15] wl[195] vdd gnd cell_6t
Xbit_r196_c15 bl[15] br[15] wl[196] vdd gnd cell_6t
Xbit_r197_c15 bl[15] br[15] wl[197] vdd gnd cell_6t
Xbit_r198_c15 bl[15] br[15] wl[198] vdd gnd cell_6t
Xbit_r199_c15 bl[15] br[15] wl[199] vdd gnd cell_6t
Xbit_r200_c15 bl[15] br[15] wl[200] vdd gnd cell_6t
Xbit_r201_c15 bl[15] br[15] wl[201] vdd gnd cell_6t
Xbit_r202_c15 bl[15] br[15] wl[202] vdd gnd cell_6t
Xbit_r203_c15 bl[15] br[15] wl[203] vdd gnd cell_6t
Xbit_r204_c15 bl[15] br[15] wl[204] vdd gnd cell_6t
Xbit_r205_c15 bl[15] br[15] wl[205] vdd gnd cell_6t
Xbit_r206_c15 bl[15] br[15] wl[206] vdd gnd cell_6t
Xbit_r207_c15 bl[15] br[15] wl[207] vdd gnd cell_6t
Xbit_r208_c15 bl[15] br[15] wl[208] vdd gnd cell_6t
Xbit_r209_c15 bl[15] br[15] wl[209] vdd gnd cell_6t
Xbit_r210_c15 bl[15] br[15] wl[210] vdd gnd cell_6t
Xbit_r211_c15 bl[15] br[15] wl[211] vdd gnd cell_6t
Xbit_r212_c15 bl[15] br[15] wl[212] vdd gnd cell_6t
Xbit_r213_c15 bl[15] br[15] wl[213] vdd gnd cell_6t
Xbit_r214_c15 bl[15] br[15] wl[214] vdd gnd cell_6t
Xbit_r215_c15 bl[15] br[15] wl[215] vdd gnd cell_6t
Xbit_r216_c15 bl[15] br[15] wl[216] vdd gnd cell_6t
Xbit_r217_c15 bl[15] br[15] wl[217] vdd gnd cell_6t
Xbit_r218_c15 bl[15] br[15] wl[218] vdd gnd cell_6t
Xbit_r219_c15 bl[15] br[15] wl[219] vdd gnd cell_6t
Xbit_r220_c15 bl[15] br[15] wl[220] vdd gnd cell_6t
Xbit_r221_c15 bl[15] br[15] wl[221] vdd gnd cell_6t
Xbit_r222_c15 bl[15] br[15] wl[222] vdd gnd cell_6t
Xbit_r223_c15 bl[15] br[15] wl[223] vdd gnd cell_6t
Xbit_r224_c15 bl[15] br[15] wl[224] vdd gnd cell_6t
Xbit_r225_c15 bl[15] br[15] wl[225] vdd gnd cell_6t
Xbit_r226_c15 bl[15] br[15] wl[226] vdd gnd cell_6t
Xbit_r227_c15 bl[15] br[15] wl[227] vdd gnd cell_6t
Xbit_r228_c15 bl[15] br[15] wl[228] vdd gnd cell_6t
Xbit_r229_c15 bl[15] br[15] wl[229] vdd gnd cell_6t
Xbit_r230_c15 bl[15] br[15] wl[230] vdd gnd cell_6t
Xbit_r231_c15 bl[15] br[15] wl[231] vdd gnd cell_6t
Xbit_r232_c15 bl[15] br[15] wl[232] vdd gnd cell_6t
Xbit_r233_c15 bl[15] br[15] wl[233] vdd gnd cell_6t
Xbit_r234_c15 bl[15] br[15] wl[234] vdd gnd cell_6t
Xbit_r235_c15 bl[15] br[15] wl[235] vdd gnd cell_6t
Xbit_r236_c15 bl[15] br[15] wl[236] vdd gnd cell_6t
Xbit_r237_c15 bl[15] br[15] wl[237] vdd gnd cell_6t
Xbit_r238_c15 bl[15] br[15] wl[238] vdd gnd cell_6t
Xbit_r239_c15 bl[15] br[15] wl[239] vdd gnd cell_6t
Xbit_r240_c15 bl[15] br[15] wl[240] vdd gnd cell_6t
Xbit_r241_c15 bl[15] br[15] wl[241] vdd gnd cell_6t
Xbit_r242_c15 bl[15] br[15] wl[242] vdd gnd cell_6t
Xbit_r243_c15 bl[15] br[15] wl[243] vdd gnd cell_6t
Xbit_r244_c15 bl[15] br[15] wl[244] vdd gnd cell_6t
Xbit_r245_c15 bl[15] br[15] wl[245] vdd gnd cell_6t
Xbit_r246_c15 bl[15] br[15] wl[246] vdd gnd cell_6t
Xbit_r247_c15 bl[15] br[15] wl[247] vdd gnd cell_6t
Xbit_r248_c15 bl[15] br[15] wl[248] vdd gnd cell_6t
Xbit_r249_c15 bl[15] br[15] wl[249] vdd gnd cell_6t
Xbit_r250_c15 bl[15] br[15] wl[250] vdd gnd cell_6t
Xbit_r251_c15 bl[15] br[15] wl[251] vdd gnd cell_6t
Xbit_r252_c15 bl[15] br[15] wl[252] vdd gnd cell_6t
Xbit_r253_c15 bl[15] br[15] wl[253] vdd gnd cell_6t
Xbit_r254_c15 bl[15] br[15] wl[254] vdd gnd cell_6t
Xbit_r255_c15 bl[15] br[15] wl[255] vdd gnd cell_6t
Xbit_r256_c15 bl[15] br[15] wl[256] vdd gnd cell_6t
Xbit_r257_c15 bl[15] br[15] wl[257] vdd gnd cell_6t
Xbit_r258_c15 bl[15] br[15] wl[258] vdd gnd cell_6t
Xbit_r259_c15 bl[15] br[15] wl[259] vdd gnd cell_6t
Xbit_r260_c15 bl[15] br[15] wl[260] vdd gnd cell_6t
Xbit_r261_c15 bl[15] br[15] wl[261] vdd gnd cell_6t
Xbit_r262_c15 bl[15] br[15] wl[262] vdd gnd cell_6t
Xbit_r263_c15 bl[15] br[15] wl[263] vdd gnd cell_6t
Xbit_r264_c15 bl[15] br[15] wl[264] vdd gnd cell_6t
Xbit_r265_c15 bl[15] br[15] wl[265] vdd gnd cell_6t
Xbit_r266_c15 bl[15] br[15] wl[266] vdd gnd cell_6t
Xbit_r267_c15 bl[15] br[15] wl[267] vdd gnd cell_6t
Xbit_r268_c15 bl[15] br[15] wl[268] vdd gnd cell_6t
Xbit_r269_c15 bl[15] br[15] wl[269] vdd gnd cell_6t
Xbit_r270_c15 bl[15] br[15] wl[270] vdd gnd cell_6t
Xbit_r271_c15 bl[15] br[15] wl[271] vdd gnd cell_6t
Xbit_r272_c15 bl[15] br[15] wl[272] vdd gnd cell_6t
Xbit_r273_c15 bl[15] br[15] wl[273] vdd gnd cell_6t
Xbit_r274_c15 bl[15] br[15] wl[274] vdd gnd cell_6t
Xbit_r275_c15 bl[15] br[15] wl[275] vdd gnd cell_6t
Xbit_r276_c15 bl[15] br[15] wl[276] vdd gnd cell_6t
Xbit_r277_c15 bl[15] br[15] wl[277] vdd gnd cell_6t
Xbit_r278_c15 bl[15] br[15] wl[278] vdd gnd cell_6t
Xbit_r279_c15 bl[15] br[15] wl[279] vdd gnd cell_6t
Xbit_r280_c15 bl[15] br[15] wl[280] vdd gnd cell_6t
Xbit_r281_c15 bl[15] br[15] wl[281] vdd gnd cell_6t
Xbit_r282_c15 bl[15] br[15] wl[282] vdd gnd cell_6t
Xbit_r283_c15 bl[15] br[15] wl[283] vdd gnd cell_6t
Xbit_r284_c15 bl[15] br[15] wl[284] vdd gnd cell_6t
Xbit_r285_c15 bl[15] br[15] wl[285] vdd gnd cell_6t
Xbit_r286_c15 bl[15] br[15] wl[286] vdd gnd cell_6t
Xbit_r287_c15 bl[15] br[15] wl[287] vdd gnd cell_6t
Xbit_r288_c15 bl[15] br[15] wl[288] vdd gnd cell_6t
Xbit_r289_c15 bl[15] br[15] wl[289] vdd gnd cell_6t
Xbit_r290_c15 bl[15] br[15] wl[290] vdd gnd cell_6t
Xbit_r291_c15 bl[15] br[15] wl[291] vdd gnd cell_6t
Xbit_r292_c15 bl[15] br[15] wl[292] vdd gnd cell_6t
Xbit_r293_c15 bl[15] br[15] wl[293] vdd gnd cell_6t
Xbit_r294_c15 bl[15] br[15] wl[294] vdd gnd cell_6t
Xbit_r295_c15 bl[15] br[15] wl[295] vdd gnd cell_6t
Xbit_r296_c15 bl[15] br[15] wl[296] vdd gnd cell_6t
Xbit_r297_c15 bl[15] br[15] wl[297] vdd gnd cell_6t
Xbit_r298_c15 bl[15] br[15] wl[298] vdd gnd cell_6t
Xbit_r299_c15 bl[15] br[15] wl[299] vdd gnd cell_6t
Xbit_r300_c15 bl[15] br[15] wl[300] vdd gnd cell_6t
Xbit_r301_c15 bl[15] br[15] wl[301] vdd gnd cell_6t
Xbit_r302_c15 bl[15] br[15] wl[302] vdd gnd cell_6t
Xbit_r303_c15 bl[15] br[15] wl[303] vdd gnd cell_6t
Xbit_r304_c15 bl[15] br[15] wl[304] vdd gnd cell_6t
Xbit_r305_c15 bl[15] br[15] wl[305] vdd gnd cell_6t
Xbit_r306_c15 bl[15] br[15] wl[306] vdd gnd cell_6t
Xbit_r307_c15 bl[15] br[15] wl[307] vdd gnd cell_6t
Xbit_r308_c15 bl[15] br[15] wl[308] vdd gnd cell_6t
Xbit_r309_c15 bl[15] br[15] wl[309] vdd gnd cell_6t
Xbit_r310_c15 bl[15] br[15] wl[310] vdd gnd cell_6t
Xbit_r311_c15 bl[15] br[15] wl[311] vdd gnd cell_6t
Xbit_r312_c15 bl[15] br[15] wl[312] vdd gnd cell_6t
Xbit_r313_c15 bl[15] br[15] wl[313] vdd gnd cell_6t
Xbit_r314_c15 bl[15] br[15] wl[314] vdd gnd cell_6t
Xbit_r315_c15 bl[15] br[15] wl[315] vdd gnd cell_6t
Xbit_r316_c15 bl[15] br[15] wl[316] vdd gnd cell_6t
Xbit_r317_c15 bl[15] br[15] wl[317] vdd gnd cell_6t
Xbit_r318_c15 bl[15] br[15] wl[318] vdd gnd cell_6t
Xbit_r319_c15 bl[15] br[15] wl[319] vdd gnd cell_6t
Xbit_r320_c15 bl[15] br[15] wl[320] vdd gnd cell_6t
Xbit_r321_c15 bl[15] br[15] wl[321] vdd gnd cell_6t
Xbit_r322_c15 bl[15] br[15] wl[322] vdd gnd cell_6t
Xbit_r323_c15 bl[15] br[15] wl[323] vdd gnd cell_6t
Xbit_r324_c15 bl[15] br[15] wl[324] vdd gnd cell_6t
Xbit_r325_c15 bl[15] br[15] wl[325] vdd gnd cell_6t
Xbit_r326_c15 bl[15] br[15] wl[326] vdd gnd cell_6t
Xbit_r327_c15 bl[15] br[15] wl[327] vdd gnd cell_6t
Xbit_r328_c15 bl[15] br[15] wl[328] vdd gnd cell_6t
Xbit_r329_c15 bl[15] br[15] wl[329] vdd gnd cell_6t
Xbit_r330_c15 bl[15] br[15] wl[330] vdd gnd cell_6t
Xbit_r331_c15 bl[15] br[15] wl[331] vdd gnd cell_6t
Xbit_r332_c15 bl[15] br[15] wl[332] vdd gnd cell_6t
Xbit_r333_c15 bl[15] br[15] wl[333] vdd gnd cell_6t
Xbit_r334_c15 bl[15] br[15] wl[334] vdd gnd cell_6t
Xbit_r335_c15 bl[15] br[15] wl[335] vdd gnd cell_6t
Xbit_r336_c15 bl[15] br[15] wl[336] vdd gnd cell_6t
Xbit_r337_c15 bl[15] br[15] wl[337] vdd gnd cell_6t
Xbit_r338_c15 bl[15] br[15] wl[338] vdd gnd cell_6t
Xbit_r339_c15 bl[15] br[15] wl[339] vdd gnd cell_6t
Xbit_r340_c15 bl[15] br[15] wl[340] vdd gnd cell_6t
Xbit_r341_c15 bl[15] br[15] wl[341] vdd gnd cell_6t
Xbit_r342_c15 bl[15] br[15] wl[342] vdd gnd cell_6t
Xbit_r343_c15 bl[15] br[15] wl[343] vdd gnd cell_6t
Xbit_r344_c15 bl[15] br[15] wl[344] vdd gnd cell_6t
Xbit_r345_c15 bl[15] br[15] wl[345] vdd gnd cell_6t
Xbit_r346_c15 bl[15] br[15] wl[346] vdd gnd cell_6t
Xbit_r347_c15 bl[15] br[15] wl[347] vdd gnd cell_6t
Xbit_r348_c15 bl[15] br[15] wl[348] vdd gnd cell_6t
Xbit_r349_c15 bl[15] br[15] wl[349] vdd gnd cell_6t
Xbit_r350_c15 bl[15] br[15] wl[350] vdd gnd cell_6t
Xbit_r351_c15 bl[15] br[15] wl[351] vdd gnd cell_6t
Xbit_r352_c15 bl[15] br[15] wl[352] vdd gnd cell_6t
Xbit_r353_c15 bl[15] br[15] wl[353] vdd gnd cell_6t
Xbit_r354_c15 bl[15] br[15] wl[354] vdd gnd cell_6t
Xbit_r355_c15 bl[15] br[15] wl[355] vdd gnd cell_6t
Xbit_r356_c15 bl[15] br[15] wl[356] vdd gnd cell_6t
Xbit_r357_c15 bl[15] br[15] wl[357] vdd gnd cell_6t
Xbit_r358_c15 bl[15] br[15] wl[358] vdd gnd cell_6t
Xbit_r359_c15 bl[15] br[15] wl[359] vdd gnd cell_6t
Xbit_r360_c15 bl[15] br[15] wl[360] vdd gnd cell_6t
Xbit_r361_c15 bl[15] br[15] wl[361] vdd gnd cell_6t
Xbit_r362_c15 bl[15] br[15] wl[362] vdd gnd cell_6t
Xbit_r363_c15 bl[15] br[15] wl[363] vdd gnd cell_6t
Xbit_r364_c15 bl[15] br[15] wl[364] vdd gnd cell_6t
Xbit_r365_c15 bl[15] br[15] wl[365] vdd gnd cell_6t
Xbit_r366_c15 bl[15] br[15] wl[366] vdd gnd cell_6t
Xbit_r367_c15 bl[15] br[15] wl[367] vdd gnd cell_6t
Xbit_r368_c15 bl[15] br[15] wl[368] vdd gnd cell_6t
Xbit_r369_c15 bl[15] br[15] wl[369] vdd gnd cell_6t
Xbit_r370_c15 bl[15] br[15] wl[370] vdd gnd cell_6t
Xbit_r371_c15 bl[15] br[15] wl[371] vdd gnd cell_6t
Xbit_r372_c15 bl[15] br[15] wl[372] vdd gnd cell_6t
Xbit_r373_c15 bl[15] br[15] wl[373] vdd gnd cell_6t
Xbit_r374_c15 bl[15] br[15] wl[374] vdd gnd cell_6t
Xbit_r375_c15 bl[15] br[15] wl[375] vdd gnd cell_6t
Xbit_r376_c15 bl[15] br[15] wl[376] vdd gnd cell_6t
Xbit_r377_c15 bl[15] br[15] wl[377] vdd gnd cell_6t
Xbit_r378_c15 bl[15] br[15] wl[378] vdd gnd cell_6t
Xbit_r379_c15 bl[15] br[15] wl[379] vdd gnd cell_6t
Xbit_r380_c15 bl[15] br[15] wl[380] vdd gnd cell_6t
Xbit_r381_c15 bl[15] br[15] wl[381] vdd gnd cell_6t
Xbit_r382_c15 bl[15] br[15] wl[382] vdd gnd cell_6t
Xbit_r383_c15 bl[15] br[15] wl[383] vdd gnd cell_6t
Xbit_r384_c15 bl[15] br[15] wl[384] vdd gnd cell_6t
Xbit_r385_c15 bl[15] br[15] wl[385] vdd gnd cell_6t
Xbit_r386_c15 bl[15] br[15] wl[386] vdd gnd cell_6t
Xbit_r387_c15 bl[15] br[15] wl[387] vdd gnd cell_6t
Xbit_r388_c15 bl[15] br[15] wl[388] vdd gnd cell_6t
Xbit_r389_c15 bl[15] br[15] wl[389] vdd gnd cell_6t
Xbit_r390_c15 bl[15] br[15] wl[390] vdd gnd cell_6t
Xbit_r391_c15 bl[15] br[15] wl[391] vdd gnd cell_6t
Xbit_r392_c15 bl[15] br[15] wl[392] vdd gnd cell_6t
Xbit_r393_c15 bl[15] br[15] wl[393] vdd gnd cell_6t
Xbit_r394_c15 bl[15] br[15] wl[394] vdd gnd cell_6t
Xbit_r395_c15 bl[15] br[15] wl[395] vdd gnd cell_6t
Xbit_r396_c15 bl[15] br[15] wl[396] vdd gnd cell_6t
Xbit_r397_c15 bl[15] br[15] wl[397] vdd gnd cell_6t
Xbit_r398_c15 bl[15] br[15] wl[398] vdd gnd cell_6t
Xbit_r399_c15 bl[15] br[15] wl[399] vdd gnd cell_6t
Xbit_r400_c15 bl[15] br[15] wl[400] vdd gnd cell_6t
Xbit_r401_c15 bl[15] br[15] wl[401] vdd gnd cell_6t
Xbit_r402_c15 bl[15] br[15] wl[402] vdd gnd cell_6t
Xbit_r403_c15 bl[15] br[15] wl[403] vdd gnd cell_6t
Xbit_r404_c15 bl[15] br[15] wl[404] vdd gnd cell_6t
Xbit_r405_c15 bl[15] br[15] wl[405] vdd gnd cell_6t
Xbit_r406_c15 bl[15] br[15] wl[406] vdd gnd cell_6t
Xbit_r407_c15 bl[15] br[15] wl[407] vdd gnd cell_6t
Xbit_r408_c15 bl[15] br[15] wl[408] vdd gnd cell_6t
Xbit_r409_c15 bl[15] br[15] wl[409] vdd gnd cell_6t
Xbit_r410_c15 bl[15] br[15] wl[410] vdd gnd cell_6t
Xbit_r411_c15 bl[15] br[15] wl[411] vdd gnd cell_6t
Xbit_r412_c15 bl[15] br[15] wl[412] vdd gnd cell_6t
Xbit_r413_c15 bl[15] br[15] wl[413] vdd gnd cell_6t
Xbit_r414_c15 bl[15] br[15] wl[414] vdd gnd cell_6t
Xbit_r415_c15 bl[15] br[15] wl[415] vdd gnd cell_6t
Xbit_r416_c15 bl[15] br[15] wl[416] vdd gnd cell_6t
Xbit_r417_c15 bl[15] br[15] wl[417] vdd gnd cell_6t
Xbit_r418_c15 bl[15] br[15] wl[418] vdd gnd cell_6t
Xbit_r419_c15 bl[15] br[15] wl[419] vdd gnd cell_6t
Xbit_r420_c15 bl[15] br[15] wl[420] vdd gnd cell_6t
Xbit_r421_c15 bl[15] br[15] wl[421] vdd gnd cell_6t
Xbit_r422_c15 bl[15] br[15] wl[422] vdd gnd cell_6t
Xbit_r423_c15 bl[15] br[15] wl[423] vdd gnd cell_6t
Xbit_r424_c15 bl[15] br[15] wl[424] vdd gnd cell_6t
Xbit_r425_c15 bl[15] br[15] wl[425] vdd gnd cell_6t
Xbit_r426_c15 bl[15] br[15] wl[426] vdd gnd cell_6t
Xbit_r427_c15 bl[15] br[15] wl[427] vdd gnd cell_6t
Xbit_r428_c15 bl[15] br[15] wl[428] vdd gnd cell_6t
Xbit_r429_c15 bl[15] br[15] wl[429] vdd gnd cell_6t
Xbit_r430_c15 bl[15] br[15] wl[430] vdd gnd cell_6t
Xbit_r431_c15 bl[15] br[15] wl[431] vdd gnd cell_6t
Xbit_r432_c15 bl[15] br[15] wl[432] vdd gnd cell_6t
Xbit_r433_c15 bl[15] br[15] wl[433] vdd gnd cell_6t
Xbit_r434_c15 bl[15] br[15] wl[434] vdd gnd cell_6t
Xbit_r435_c15 bl[15] br[15] wl[435] vdd gnd cell_6t
Xbit_r436_c15 bl[15] br[15] wl[436] vdd gnd cell_6t
Xbit_r437_c15 bl[15] br[15] wl[437] vdd gnd cell_6t
Xbit_r438_c15 bl[15] br[15] wl[438] vdd gnd cell_6t
Xbit_r439_c15 bl[15] br[15] wl[439] vdd gnd cell_6t
Xbit_r440_c15 bl[15] br[15] wl[440] vdd gnd cell_6t
Xbit_r441_c15 bl[15] br[15] wl[441] vdd gnd cell_6t
Xbit_r442_c15 bl[15] br[15] wl[442] vdd gnd cell_6t
Xbit_r443_c15 bl[15] br[15] wl[443] vdd gnd cell_6t
Xbit_r444_c15 bl[15] br[15] wl[444] vdd gnd cell_6t
Xbit_r445_c15 bl[15] br[15] wl[445] vdd gnd cell_6t
Xbit_r446_c15 bl[15] br[15] wl[446] vdd gnd cell_6t
Xbit_r447_c15 bl[15] br[15] wl[447] vdd gnd cell_6t
Xbit_r448_c15 bl[15] br[15] wl[448] vdd gnd cell_6t
Xbit_r449_c15 bl[15] br[15] wl[449] vdd gnd cell_6t
Xbit_r450_c15 bl[15] br[15] wl[450] vdd gnd cell_6t
Xbit_r451_c15 bl[15] br[15] wl[451] vdd gnd cell_6t
Xbit_r452_c15 bl[15] br[15] wl[452] vdd gnd cell_6t
Xbit_r453_c15 bl[15] br[15] wl[453] vdd gnd cell_6t
Xbit_r454_c15 bl[15] br[15] wl[454] vdd gnd cell_6t
Xbit_r455_c15 bl[15] br[15] wl[455] vdd gnd cell_6t
Xbit_r456_c15 bl[15] br[15] wl[456] vdd gnd cell_6t
Xbit_r457_c15 bl[15] br[15] wl[457] vdd gnd cell_6t
Xbit_r458_c15 bl[15] br[15] wl[458] vdd gnd cell_6t
Xbit_r459_c15 bl[15] br[15] wl[459] vdd gnd cell_6t
Xbit_r460_c15 bl[15] br[15] wl[460] vdd gnd cell_6t
Xbit_r461_c15 bl[15] br[15] wl[461] vdd gnd cell_6t
Xbit_r462_c15 bl[15] br[15] wl[462] vdd gnd cell_6t
Xbit_r463_c15 bl[15] br[15] wl[463] vdd gnd cell_6t
Xbit_r464_c15 bl[15] br[15] wl[464] vdd gnd cell_6t
Xbit_r465_c15 bl[15] br[15] wl[465] vdd gnd cell_6t
Xbit_r466_c15 bl[15] br[15] wl[466] vdd gnd cell_6t
Xbit_r467_c15 bl[15] br[15] wl[467] vdd gnd cell_6t
Xbit_r468_c15 bl[15] br[15] wl[468] vdd gnd cell_6t
Xbit_r469_c15 bl[15] br[15] wl[469] vdd gnd cell_6t
Xbit_r470_c15 bl[15] br[15] wl[470] vdd gnd cell_6t
Xbit_r471_c15 bl[15] br[15] wl[471] vdd gnd cell_6t
Xbit_r472_c15 bl[15] br[15] wl[472] vdd gnd cell_6t
Xbit_r473_c15 bl[15] br[15] wl[473] vdd gnd cell_6t
Xbit_r474_c15 bl[15] br[15] wl[474] vdd gnd cell_6t
Xbit_r475_c15 bl[15] br[15] wl[475] vdd gnd cell_6t
Xbit_r476_c15 bl[15] br[15] wl[476] vdd gnd cell_6t
Xbit_r477_c15 bl[15] br[15] wl[477] vdd gnd cell_6t
Xbit_r478_c15 bl[15] br[15] wl[478] vdd gnd cell_6t
Xbit_r479_c15 bl[15] br[15] wl[479] vdd gnd cell_6t
Xbit_r480_c15 bl[15] br[15] wl[480] vdd gnd cell_6t
Xbit_r481_c15 bl[15] br[15] wl[481] vdd gnd cell_6t
Xbit_r482_c15 bl[15] br[15] wl[482] vdd gnd cell_6t
Xbit_r483_c15 bl[15] br[15] wl[483] vdd gnd cell_6t
Xbit_r484_c15 bl[15] br[15] wl[484] vdd gnd cell_6t
Xbit_r485_c15 bl[15] br[15] wl[485] vdd gnd cell_6t
Xbit_r486_c15 bl[15] br[15] wl[486] vdd gnd cell_6t
Xbit_r487_c15 bl[15] br[15] wl[487] vdd gnd cell_6t
Xbit_r488_c15 bl[15] br[15] wl[488] vdd gnd cell_6t
Xbit_r489_c15 bl[15] br[15] wl[489] vdd gnd cell_6t
Xbit_r490_c15 bl[15] br[15] wl[490] vdd gnd cell_6t
Xbit_r491_c15 bl[15] br[15] wl[491] vdd gnd cell_6t
Xbit_r492_c15 bl[15] br[15] wl[492] vdd gnd cell_6t
Xbit_r493_c15 bl[15] br[15] wl[493] vdd gnd cell_6t
Xbit_r494_c15 bl[15] br[15] wl[494] vdd gnd cell_6t
Xbit_r495_c15 bl[15] br[15] wl[495] vdd gnd cell_6t
Xbit_r496_c15 bl[15] br[15] wl[496] vdd gnd cell_6t
Xbit_r497_c15 bl[15] br[15] wl[497] vdd gnd cell_6t
Xbit_r498_c15 bl[15] br[15] wl[498] vdd gnd cell_6t
Xbit_r499_c15 bl[15] br[15] wl[499] vdd gnd cell_6t
Xbit_r500_c15 bl[15] br[15] wl[500] vdd gnd cell_6t
Xbit_r501_c15 bl[15] br[15] wl[501] vdd gnd cell_6t
Xbit_r502_c15 bl[15] br[15] wl[502] vdd gnd cell_6t
Xbit_r503_c15 bl[15] br[15] wl[503] vdd gnd cell_6t
Xbit_r504_c15 bl[15] br[15] wl[504] vdd gnd cell_6t
Xbit_r505_c15 bl[15] br[15] wl[505] vdd gnd cell_6t
Xbit_r506_c15 bl[15] br[15] wl[506] vdd gnd cell_6t
Xbit_r507_c15 bl[15] br[15] wl[507] vdd gnd cell_6t
Xbit_r508_c15 bl[15] br[15] wl[508] vdd gnd cell_6t
Xbit_r509_c15 bl[15] br[15] wl[509] vdd gnd cell_6t
Xbit_r510_c15 bl[15] br[15] wl[510] vdd gnd cell_6t
Xbit_r511_c15 bl[15] br[15] wl[511] vdd gnd cell_6t
Xbit_r0_c16 bl[16] br[16] wl[0] vdd gnd cell_6t
Xbit_r1_c16 bl[16] br[16] wl[1] vdd gnd cell_6t
Xbit_r2_c16 bl[16] br[16] wl[2] vdd gnd cell_6t
Xbit_r3_c16 bl[16] br[16] wl[3] vdd gnd cell_6t
Xbit_r4_c16 bl[16] br[16] wl[4] vdd gnd cell_6t
Xbit_r5_c16 bl[16] br[16] wl[5] vdd gnd cell_6t
Xbit_r6_c16 bl[16] br[16] wl[6] vdd gnd cell_6t
Xbit_r7_c16 bl[16] br[16] wl[7] vdd gnd cell_6t
Xbit_r8_c16 bl[16] br[16] wl[8] vdd gnd cell_6t
Xbit_r9_c16 bl[16] br[16] wl[9] vdd gnd cell_6t
Xbit_r10_c16 bl[16] br[16] wl[10] vdd gnd cell_6t
Xbit_r11_c16 bl[16] br[16] wl[11] vdd gnd cell_6t
Xbit_r12_c16 bl[16] br[16] wl[12] vdd gnd cell_6t
Xbit_r13_c16 bl[16] br[16] wl[13] vdd gnd cell_6t
Xbit_r14_c16 bl[16] br[16] wl[14] vdd gnd cell_6t
Xbit_r15_c16 bl[16] br[16] wl[15] vdd gnd cell_6t
Xbit_r16_c16 bl[16] br[16] wl[16] vdd gnd cell_6t
Xbit_r17_c16 bl[16] br[16] wl[17] vdd gnd cell_6t
Xbit_r18_c16 bl[16] br[16] wl[18] vdd gnd cell_6t
Xbit_r19_c16 bl[16] br[16] wl[19] vdd gnd cell_6t
Xbit_r20_c16 bl[16] br[16] wl[20] vdd gnd cell_6t
Xbit_r21_c16 bl[16] br[16] wl[21] vdd gnd cell_6t
Xbit_r22_c16 bl[16] br[16] wl[22] vdd gnd cell_6t
Xbit_r23_c16 bl[16] br[16] wl[23] vdd gnd cell_6t
Xbit_r24_c16 bl[16] br[16] wl[24] vdd gnd cell_6t
Xbit_r25_c16 bl[16] br[16] wl[25] vdd gnd cell_6t
Xbit_r26_c16 bl[16] br[16] wl[26] vdd gnd cell_6t
Xbit_r27_c16 bl[16] br[16] wl[27] vdd gnd cell_6t
Xbit_r28_c16 bl[16] br[16] wl[28] vdd gnd cell_6t
Xbit_r29_c16 bl[16] br[16] wl[29] vdd gnd cell_6t
Xbit_r30_c16 bl[16] br[16] wl[30] vdd gnd cell_6t
Xbit_r31_c16 bl[16] br[16] wl[31] vdd gnd cell_6t
Xbit_r32_c16 bl[16] br[16] wl[32] vdd gnd cell_6t
Xbit_r33_c16 bl[16] br[16] wl[33] vdd gnd cell_6t
Xbit_r34_c16 bl[16] br[16] wl[34] vdd gnd cell_6t
Xbit_r35_c16 bl[16] br[16] wl[35] vdd gnd cell_6t
Xbit_r36_c16 bl[16] br[16] wl[36] vdd gnd cell_6t
Xbit_r37_c16 bl[16] br[16] wl[37] vdd gnd cell_6t
Xbit_r38_c16 bl[16] br[16] wl[38] vdd gnd cell_6t
Xbit_r39_c16 bl[16] br[16] wl[39] vdd gnd cell_6t
Xbit_r40_c16 bl[16] br[16] wl[40] vdd gnd cell_6t
Xbit_r41_c16 bl[16] br[16] wl[41] vdd gnd cell_6t
Xbit_r42_c16 bl[16] br[16] wl[42] vdd gnd cell_6t
Xbit_r43_c16 bl[16] br[16] wl[43] vdd gnd cell_6t
Xbit_r44_c16 bl[16] br[16] wl[44] vdd gnd cell_6t
Xbit_r45_c16 bl[16] br[16] wl[45] vdd gnd cell_6t
Xbit_r46_c16 bl[16] br[16] wl[46] vdd gnd cell_6t
Xbit_r47_c16 bl[16] br[16] wl[47] vdd gnd cell_6t
Xbit_r48_c16 bl[16] br[16] wl[48] vdd gnd cell_6t
Xbit_r49_c16 bl[16] br[16] wl[49] vdd gnd cell_6t
Xbit_r50_c16 bl[16] br[16] wl[50] vdd gnd cell_6t
Xbit_r51_c16 bl[16] br[16] wl[51] vdd gnd cell_6t
Xbit_r52_c16 bl[16] br[16] wl[52] vdd gnd cell_6t
Xbit_r53_c16 bl[16] br[16] wl[53] vdd gnd cell_6t
Xbit_r54_c16 bl[16] br[16] wl[54] vdd gnd cell_6t
Xbit_r55_c16 bl[16] br[16] wl[55] vdd gnd cell_6t
Xbit_r56_c16 bl[16] br[16] wl[56] vdd gnd cell_6t
Xbit_r57_c16 bl[16] br[16] wl[57] vdd gnd cell_6t
Xbit_r58_c16 bl[16] br[16] wl[58] vdd gnd cell_6t
Xbit_r59_c16 bl[16] br[16] wl[59] vdd gnd cell_6t
Xbit_r60_c16 bl[16] br[16] wl[60] vdd gnd cell_6t
Xbit_r61_c16 bl[16] br[16] wl[61] vdd gnd cell_6t
Xbit_r62_c16 bl[16] br[16] wl[62] vdd gnd cell_6t
Xbit_r63_c16 bl[16] br[16] wl[63] vdd gnd cell_6t
Xbit_r64_c16 bl[16] br[16] wl[64] vdd gnd cell_6t
Xbit_r65_c16 bl[16] br[16] wl[65] vdd gnd cell_6t
Xbit_r66_c16 bl[16] br[16] wl[66] vdd gnd cell_6t
Xbit_r67_c16 bl[16] br[16] wl[67] vdd gnd cell_6t
Xbit_r68_c16 bl[16] br[16] wl[68] vdd gnd cell_6t
Xbit_r69_c16 bl[16] br[16] wl[69] vdd gnd cell_6t
Xbit_r70_c16 bl[16] br[16] wl[70] vdd gnd cell_6t
Xbit_r71_c16 bl[16] br[16] wl[71] vdd gnd cell_6t
Xbit_r72_c16 bl[16] br[16] wl[72] vdd gnd cell_6t
Xbit_r73_c16 bl[16] br[16] wl[73] vdd gnd cell_6t
Xbit_r74_c16 bl[16] br[16] wl[74] vdd gnd cell_6t
Xbit_r75_c16 bl[16] br[16] wl[75] vdd gnd cell_6t
Xbit_r76_c16 bl[16] br[16] wl[76] vdd gnd cell_6t
Xbit_r77_c16 bl[16] br[16] wl[77] vdd gnd cell_6t
Xbit_r78_c16 bl[16] br[16] wl[78] vdd gnd cell_6t
Xbit_r79_c16 bl[16] br[16] wl[79] vdd gnd cell_6t
Xbit_r80_c16 bl[16] br[16] wl[80] vdd gnd cell_6t
Xbit_r81_c16 bl[16] br[16] wl[81] vdd gnd cell_6t
Xbit_r82_c16 bl[16] br[16] wl[82] vdd gnd cell_6t
Xbit_r83_c16 bl[16] br[16] wl[83] vdd gnd cell_6t
Xbit_r84_c16 bl[16] br[16] wl[84] vdd gnd cell_6t
Xbit_r85_c16 bl[16] br[16] wl[85] vdd gnd cell_6t
Xbit_r86_c16 bl[16] br[16] wl[86] vdd gnd cell_6t
Xbit_r87_c16 bl[16] br[16] wl[87] vdd gnd cell_6t
Xbit_r88_c16 bl[16] br[16] wl[88] vdd gnd cell_6t
Xbit_r89_c16 bl[16] br[16] wl[89] vdd gnd cell_6t
Xbit_r90_c16 bl[16] br[16] wl[90] vdd gnd cell_6t
Xbit_r91_c16 bl[16] br[16] wl[91] vdd gnd cell_6t
Xbit_r92_c16 bl[16] br[16] wl[92] vdd gnd cell_6t
Xbit_r93_c16 bl[16] br[16] wl[93] vdd gnd cell_6t
Xbit_r94_c16 bl[16] br[16] wl[94] vdd gnd cell_6t
Xbit_r95_c16 bl[16] br[16] wl[95] vdd gnd cell_6t
Xbit_r96_c16 bl[16] br[16] wl[96] vdd gnd cell_6t
Xbit_r97_c16 bl[16] br[16] wl[97] vdd gnd cell_6t
Xbit_r98_c16 bl[16] br[16] wl[98] vdd gnd cell_6t
Xbit_r99_c16 bl[16] br[16] wl[99] vdd gnd cell_6t
Xbit_r100_c16 bl[16] br[16] wl[100] vdd gnd cell_6t
Xbit_r101_c16 bl[16] br[16] wl[101] vdd gnd cell_6t
Xbit_r102_c16 bl[16] br[16] wl[102] vdd gnd cell_6t
Xbit_r103_c16 bl[16] br[16] wl[103] vdd gnd cell_6t
Xbit_r104_c16 bl[16] br[16] wl[104] vdd gnd cell_6t
Xbit_r105_c16 bl[16] br[16] wl[105] vdd gnd cell_6t
Xbit_r106_c16 bl[16] br[16] wl[106] vdd gnd cell_6t
Xbit_r107_c16 bl[16] br[16] wl[107] vdd gnd cell_6t
Xbit_r108_c16 bl[16] br[16] wl[108] vdd gnd cell_6t
Xbit_r109_c16 bl[16] br[16] wl[109] vdd gnd cell_6t
Xbit_r110_c16 bl[16] br[16] wl[110] vdd gnd cell_6t
Xbit_r111_c16 bl[16] br[16] wl[111] vdd gnd cell_6t
Xbit_r112_c16 bl[16] br[16] wl[112] vdd gnd cell_6t
Xbit_r113_c16 bl[16] br[16] wl[113] vdd gnd cell_6t
Xbit_r114_c16 bl[16] br[16] wl[114] vdd gnd cell_6t
Xbit_r115_c16 bl[16] br[16] wl[115] vdd gnd cell_6t
Xbit_r116_c16 bl[16] br[16] wl[116] vdd gnd cell_6t
Xbit_r117_c16 bl[16] br[16] wl[117] vdd gnd cell_6t
Xbit_r118_c16 bl[16] br[16] wl[118] vdd gnd cell_6t
Xbit_r119_c16 bl[16] br[16] wl[119] vdd gnd cell_6t
Xbit_r120_c16 bl[16] br[16] wl[120] vdd gnd cell_6t
Xbit_r121_c16 bl[16] br[16] wl[121] vdd gnd cell_6t
Xbit_r122_c16 bl[16] br[16] wl[122] vdd gnd cell_6t
Xbit_r123_c16 bl[16] br[16] wl[123] vdd gnd cell_6t
Xbit_r124_c16 bl[16] br[16] wl[124] vdd gnd cell_6t
Xbit_r125_c16 bl[16] br[16] wl[125] vdd gnd cell_6t
Xbit_r126_c16 bl[16] br[16] wl[126] vdd gnd cell_6t
Xbit_r127_c16 bl[16] br[16] wl[127] vdd gnd cell_6t
Xbit_r128_c16 bl[16] br[16] wl[128] vdd gnd cell_6t
Xbit_r129_c16 bl[16] br[16] wl[129] vdd gnd cell_6t
Xbit_r130_c16 bl[16] br[16] wl[130] vdd gnd cell_6t
Xbit_r131_c16 bl[16] br[16] wl[131] vdd gnd cell_6t
Xbit_r132_c16 bl[16] br[16] wl[132] vdd gnd cell_6t
Xbit_r133_c16 bl[16] br[16] wl[133] vdd gnd cell_6t
Xbit_r134_c16 bl[16] br[16] wl[134] vdd gnd cell_6t
Xbit_r135_c16 bl[16] br[16] wl[135] vdd gnd cell_6t
Xbit_r136_c16 bl[16] br[16] wl[136] vdd gnd cell_6t
Xbit_r137_c16 bl[16] br[16] wl[137] vdd gnd cell_6t
Xbit_r138_c16 bl[16] br[16] wl[138] vdd gnd cell_6t
Xbit_r139_c16 bl[16] br[16] wl[139] vdd gnd cell_6t
Xbit_r140_c16 bl[16] br[16] wl[140] vdd gnd cell_6t
Xbit_r141_c16 bl[16] br[16] wl[141] vdd gnd cell_6t
Xbit_r142_c16 bl[16] br[16] wl[142] vdd gnd cell_6t
Xbit_r143_c16 bl[16] br[16] wl[143] vdd gnd cell_6t
Xbit_r144_c16 bl[16] br[16] wl[144] vdd gnd cell_6t
Xbit_r145_c16 bl[16] br[16] wl[145] vdd gnd cell_6t
Xbit_r146_c16 bl[16] br[16] wl[146] vdd gnd cell_6t
Xbit_r147_c16 bl[16] br[16] wl[147] vdd gnd cell_6t
Xbit_r148_c16 bl[16] br[16] wl[148] vdd gnd cell_6t
Xbit_r149_c16 bl[16] br[16] wl[149] vdd gnd cell_6t
Xbit_r150_c16 bl[16] br[16] wl[150] vdd gnd cell_6t
Xbit_r151_c16 bl[16] br[16] wl[151] vdd gnd cell_6t
Xbit_r152_c16 bl[16] br[16] wl[152] vdd gnd cell_6t
Xbit_r153_c16 bl[16] br[16] wl[153] vdd gnd cell_6t
Xbit_r154_c16 bl[16] br[16] wl[154] vdd gnd cell_6t
Xbit_r155_c16 bl[16] br[16] wl[155] vdd gnd cell_6t
Xbit_r156_c16 bl[16] br[16] wl[156] vdd gnd cell_6t
Xbit_r157_c16 bl[16] br[16] wl[157] vdd gnd cell_6t
Xbit_r158_c16 bl[16] br[16] wl[158] vdd gnd cell_6t
Xbit_r159_c16 bl[16] br[16] wl[159] vdd gnd cell_6t
Xbit_r160_c16 bl[16] br[16] wl[160] vdd gnd cell_6t
Xbit_r161_c16 bl[16] br[16] wl[161] vdd gnd cell_6t
Xbit_r162_c16 bl[16] br[16] wl[162] vdd gnd cell_6t
Xbit_r163_c16 bl[16] br[16] wl[163] vdd gnd cell_6t
Xbit_r164_c16 bl[16] br[16] wl[164] vdd gnd cell_6t
Xbit_r165_c16 bl[16] br[16] wl[165] vdd gnd cell_6t
Xbit_r166_c16 bl[16] br[16] wl[166] vdd gnd cell_6t
Xbit_r167_c16 bl[16] br[16] wl[167] vdd gnd cell_6t
Xbit_r168_c16 bl[16] br[16] wl[168] vdd gnd cell_6t
Xbit_r169_c16 bl[16] br[16] wl[169] vdd gnd cell_6t
Xbit_r170_c16 bl[16] br[16] wl[170] vdd gnd cell_6t
Xbit_r171_c16 bl[16] br[16] wl[171] vdd gnd cell_6t
Xbit_r172_c16 bl[16] br[16] wl[172] vdd gnd cell_6t
Xbit_r173_c16 bl[16] br[16] wl[173] vdd gnd cell_6t
Xbit_r174_c16 bl[16] br[16] wl[174] vdd gnd cell_6t
Xbit_r175_c16 bl[16] br[16] wl[175] vdd gnd cell_6t
Xbit_r176_c16 bl[16] br[16] wl[176] vdd gnd cell_6t
Xbit_r177_c16 bl[16] br[16] wl[177] vdd gnd cell_6t
Xbit_r178_c16 bl[16] br[16] wl[178] vdd gnd cell_6t
Xbit_r179_c16 bl[16] br[16] wl[179] vdd gnd cell_6t
Xbit_r180_c16 bl[16] br[16] wl[180] vdd gnd cell_6t
Xbit_r181_c16 bl[16] br[16] wl[181] vdd gnd cell_6t
Xbit_r182_c16 bl[16] br[16] wl[182] vdd gnd cell_6t
Xbit_r183_c16 bl[16] br[16] wl[183] vdd gnd cell_6t
Xbit_r184_c16 bl[16] br[16] wl[184] vdd gnd cell_6t
Xbit_r185_c16 bl[16] br[16] wl[185] vdd gnd cell_6t
Xbit_r186_c16 bl[16] br[16] wl[186] vdd gnd cell_6t
Xbit_r187_c16 bl[16] br[16] wl[187] vdd gnd cell_6t
Xbit_r188_c16 bl[16] br[16] wl[188] vdd gnd cell_6t
Xbit_r189_c16 bl[16] br[16] wl[189] vdd gnd cell_6t
Xbit_r190_c16 bl[16] br[16] wl[190] vdd gnd cell_6t
Xbit_r191_c16 bl[16] br[16] wl[191] vdd gnd cell_6t
Xbit_r192_c16 bl[16] br[16] wl[192] vdd gnd cell_6t
Xbit_r193_c16 bl[16] br[16] wl[193] vdd gnd cell_6t
Xbit_r194_c16 bl[16] br[16] wl[194] vdd gnd cell_6t
Xbit_r195_c16 bl[16] br[16] wl[195] vdd gnd cell_6t
Xbit_r196_c16 bl[16] br[16] wl[196] vdd gnd cell_6t
Xbit_r197_c16 bl[16] br[16] wl[197] vdd gnd cell_6t
Xbit_r198_c16 bl[16] br[16] wl[198] vdd gnd cell_6t
Xbit_r199_c16 bl[16] br[16] wl[199] vdd gnd cell_6t
Xbit_r200_c16 bl[16] br[16] wl[200] vdd gnd cell_6t
Xbit_r201_c16 bl[16] br[16] wl[201] vdd gnd cell_6t
Xbit_r202_c16 bl[16] br[16] wl[202] vdd gnd cell_6t
Xbit_r203_c16 bl[16] br[16] wl[203] vdd gnd cell_6t
Xbit_r204_c16 bl[16] br[16] wl[204] vdd gnd cell_6t
Xbit_r205_c16 bl[16] br[16] wl[205] vdd gnd cell_6t
Xbit_r206_c16 bl[16] br[16] wl[206] vdd gnd cell_6t
Xbit_r207_c16 bl[16] br[16] wl[207] vdd gnd cell_6t
Xbit_r208_c16 bl[16] br[16] wl[208] vdd gnd cell_6t
Xbit_r209_c16 bl[16] br[16] wl[209] vdd gnd cell_6t
Xbit_r210_c16 bl[16] br[16] wl[210] vdd gnd cell_6t
Xbit_r211_c16 bl[16] br[16] wl[211] vdd gnd cell_6t
Xbit_r212_c16 bl[16] br[16] wl[212] vdd gnd cell_6t
Xbit_r213_c16 bl[16] br[16] wl[213] vdd gnd cell_6t
Xbit_r214_c16 bl[16] br[16] wl[214] vdd gnd cell_6t
Xbit_r215_c16 bl[16] br[16] wl[215] vdd gnd cell_6t
Xbit_r216_c16 bl[16] br[16] wl[216] vdd gnd cell_6t
Xbit_r217_c16 bl[16] br[16] wl[217] vdd gnd cell_6t
Xbit_r218_c16 bl[16] br[16] wl[218] vdd gnd cell_6t
Xbit_r219_c16 bl[16] br[16] wl[219] vdd gnd cell_6t
Xbit_r220_c16 bl[16] br[16] wl[220] vdd gnd cell_6t
Xbit_r221_c16 bl[16] br[16] wl[221] vdd gnd cell_6t
Xbit_r222_c16 bl[16] br[16] wl[222] vdd gnd cell_6t
Xbit_r223_c16 bl[16] br[16] wl[223] vdd gnd cell_6t
Xbit_r224_c16 bl[16] br[16] wl[224] vdd gnd cell_6t
Xbit_r225_c16 bl[16] br[16] wl[225] vdd gnd cell_6t
Xbit_r226_c16 bl[16] br[16] wl[226] vdd gnd cell_6t
Xbit_r227_c16 bl[16] br[16] wl[227] vdd gnd cell_6t
Xbit_r228_c16 bl[16] br[16] wl[228] vdd gnd cell_6t
Xbit_r229_c16 bl[16] br[16] wl[229] vdd gnd cell_6t
Xbit_r230_c16 bl[16] br[16] wl[230] vdd gnd cell_6t
Xbit_r231_c16 bl[16] br[16] wl[231] vdd gnd cell_6t
Xbit_r232_c16 bl[16] br[16] wl[232] vdd gnd cell_6t
Xbit_r233_c16 bl[16] br[16] wl[233] vdd gnd cell_6t
Xbit_r234_c16 bl[16] br[16] wl[234] vdd gnd cell_6t
Xbit_r235_c16 bl[16] br[16] wl[235] vdd gnd cell_6t
Xbit_r236_c16 bl[16] br[16] wl[236] vdd gnd cell_6t
Xbit_r237_c16 bl[16] br[16] wl[237] vdd gnd cell_6t
Xbit_r238_c16 bl[16] br[16] wl[238] vdd gnd cell_6t
Xbit_r239_c16 bl[16] br[16] wl[239] vdd gnd cell_6t
Xbit_r240_c16 bl[16] br[16] wl[240] vdd gnd cell_6t
Xbit_r241_c16 bl[16] br[16] wl[241] vdd gnd cell_6t
Xbit_r242_c16 bl[16] br[16] wl[242] vdd gnd cell_6t
Xbit_r243_c16 bl[16] br[16] wl[243] vdd gnd cell_6t
Xbit_r244_c16 bl[16] br[16] wl[244] vdd gnd cell_6t
Xbit_r245_c16 bl[16] br[16] wl[245] vdd gnd cell_6t
Xbit_r246_c16 bl[16] br[16] wl[246] vdd gnd cell_6t
Xbit_r247_c16 bl[16] br[16] wl[247] vdd gnd cell_6t
Xbit_r248_c16 bl[16] br[16] wl[248] vdd gnd cell_6t
Xbit_r249_c16 bl[16] br[16] wl[249] vdd gnd cell_6t
Xbit_r250_c16 bl[16] br[16] wl[250] vdd gnd cell_6t
Xbit_r251_c16 bl[16] br[16] wl[251] vdd gnd cell_6t
Xbit_r252_c16 bl[16] br[16] wl[252] vdd gnd cell_6t
Xbit_r253_c16 bl[16] br[16] wl[253] vdd gnd cell_6t
Xbit_r254_c16 bl[16] br[16] wl[254] vdd gnd cell_6t
Xbit_r255_c16 bl[16] br[16] wl[255] vdd gnd cell_6t
Xbit_r256_c16 bl[16] br[16] wl[256] vdd gnd cell_6t
Xbit_r257_c16 bl[16] br[16] wl[257] vdd gnd cell_6t
Xbit_r258_c16 bl[16] br[16] wl[258] vdd gnd cell_6t
Xbit_r259_c16 bl[16] br[16] wl[259] vdd gnd cell_6t
Xbit_r260_c16 bl[16] br[16] wl[260] vdd gnd cell_6t
Xbit_r261_c16 bl[16] br[16] wl[261] vdd gnd cell_6t
Xbit_r262_c16 bl[16] br[16] wl[262] vdd gnd cell_6t
Xbit_r263_c16 bl[16] br[16] wl[263] vdd gnd cell_6t
Xbit_r264_c16 bl[16] br[16] wl[264] vdd gnd cell_6t
Xbit_r265_c16 bl[16] br[16] wl[265] vdd gnd cell_6t
Xbit_r266_c16 bl[16] br[16] wl[266] vdd gnd cell_6t
Xbit_r267_c16 bl[16] br[16] wl[267] vdd gnd cell_6t
Xbit_r268_c16 bl[16] br[16] wl[268] vdd gnd cell_6t
Xbit_r269_c16 bl[16] br[16] wl[269] vdd gnd cell_6t
Xbit_r270_c16 bl[16] br[16] wl[270] vdd gnd cell_6t
Xbit_r271_c16 bl[16] br[16] wl[271] vdd gnd cell_6t
Xbit_r272_c16 bl[16] br[16] wl[272] vdd gnd cell_6t
Xbit_r273_c16 bl[16] br[16] wl[273] vdd gnd cell_6t
Xbit_r274_c16 bl[16] br[16] wl[274] vdd gnd cell_6t
Xbit_r275_c16 bl[16] br[16] wl[275] vdd gnd cell_6t
Xbit_r276_c16 bl[16] br[16] wl[276] vdd gnd cell_6t
Xbit_r277_c16 bl[16] br[16] wl[277] vdd gnd cell_6t
Xbit_r278_c16 bl[16] br[16] wl[278] vdd gnd cell_6t
Xbit_r279_c16 bl[16] br[16] wl[279] vdd gnd cell_6t
Xbit_r280_c16 bl[16] br[16] wl[280] vdd gnd cell_6t
Xbit_r281_c16 bl[16] br[16] wl[281] vdd gnd cell_6t
Xbit_r282_c16 bl[16] br[16] wl[282] vdd gnd cell_6t
Xbit_r283_c16 bl[16] br[16] wl[283] vdd gnd cell_6t
Xbit_r284_c16 bl[16] br[16] wl[284] vdd gnd cell_6t
Xbit_r285_c16 bl[16] br[16] wl[285] vdd gnd cell_6t
Xbit_r286_c16 bl[16] br[16] wl[286] vdd gnd cell_6t
Xbit_r287_c16 bl[16] br[16] wl[287] vdd gnd cell_6t
Xbit_r288_c16 bl[16] br[16] wl[288] vdd gnd cell_6t
Xbit_r289_c16 bl[16] br[16] wl[289] vdd gnd cell_6t
Xbit_r290_c16 bl[16] br[16] wl[290] vdd gnd cell_6t
Xbit_r291_c16 bl[16] br[16] wl[291] vdd gnd cell_6t
Xbit_r292_c16 bl[16] br[16] wl[292] vdd gnd cell_6t
Xbit_r293_c16 bl[16] br[16] wl[293] vdd gnd cell_6t
Xbit_r294_c16 bl[16] br[16] wl[294] vdd gnd cell_6t
Xbit_r295_c16 bl[16] br[16] wl[295] vdd gnd cell_6t
Xbit_r296_c16 bl[16] br[16] wl[296] vdd gnd cell_6t
Xbit_r297_c16 bl[16] br[16] wl[297] vdd gnd cell_6t
Xbit_r298_c16 bl[16] br[16] wl[298] vdd gnd cell_6t
Xbit_r299_c16 bl[16] br[16] wl[299] vdd gnd cell_6t
Xbit_r300_c16 bl[16] br[16] wl[300] vdd gnd cell_6t
Xbit_r301_c16 bl[16] br[16] wl[301] vdd gnd cell_6t
Xbit_r302_c16 bl[16] br[16] wl[302] vdd gnd cell_6t
Xbit_r303_c16 bl[16] br[16] wl[303] vdd gnd cell_6t
Xbit_r304_c16 bl[16] br[16] wl[304] vdd gnd cell_6t
Xbit_r305_c16 bl[16] br[16] wl[305] vdd gnd cell_6t
Xbit_r306_c16 bl[16] br[16] wl[306] vdd gnd cell_6t
Xbit_r307_c16 bl[16] br[16] wl[307] vdd gnd cell_6t
Xbit_r308_c16 bl[16] br[16] wl[308] vdd gnd cell_6t
Xbit_r309_c16 bl[16] br[16] wl[309] vdd gnd cell_6t
Xbit_r310_c16 bl[16] br[16] wl[310] vdd gnd cell_6t
Xbit_r311_c16 bl[16] br[16] wl[311] vdd gnd cell_6t
Xbit_r312_c16 bl[16] br[16] wl[312] vdd gnd cell_6t
Xbit_r313_c16 bl[16] br[16] wl[313] vdd gnd cell_6t
Xbit_r314_c16 bl[16] br[16] wl[314] vdd gnd cell_6t
Xbit_r315_c16 bl[16] br[16] wl[315] vdd gnd cell_6t
Xbit_r316_c16 bl[16] br[16] wl[316] vdd gnd cell_6t
Xbit_r317_c16 bl[16] br[16] wl[317] vdd gnd cell_6t
Xbit_r318_c16 bl[16] br[16] wl[318] vdd gnd cell_6t
Xbit_r319_c16 bl[16] br[16] wl[319] vdd gnd cell_6t
Xbit_r320_c16 bl[16] br[16] wl[320] vdd gnd cell_6t
Xbit_r321_c16 bl[16] br[16] wl[321] vdd gnd cell_6t
Xbit_r322_c16 bl[16] br[16] wl[322] vdd gnd cell_6t
Xbit_r323_c16 bl[16] br[16] wl[323] vdd gnd cell_6t
Xbit_r324_c16 bl[16] br[16] wl[324] vdd gnd cell_6t
Xbit_r325_c16 bl[16] br[16] wl[325] vdd gnd cell_6t
Xbit_r326_c16 bl[16] br[16] wl[326] vdd gnd cell_6t
Xbit_r327_c16 bl[16] br[16] wl[327] vdd gnd cell_6t
Xbit_r328_c16 bl[16] br[16] wl[328] vdd gnd cell_6t
Xbit_r329_c16 bl[16] br[16] wl[329] vdd gnd cell_6t
Xbit_r330_c16 bl[16] br[16] wl[330] vdd gnd cell_6t
Xbit_r331_c16 bl[16] br[16] wl[331] vdd gnd cell_6t
Xbit_r332_c16 bl[16] br[16] wl[332] vdd gnd cell_6t
Xbit_r333_c16 bl[16] br[16] wl[333] vdd gnd cell_6t
Xbit_r334_c16 bl[16] br[16] wl[334] vdd gnd cell_6t
Xbit_r335_c16 bl[16] br[16] wl[335] vdd gnd cell_6t
Xbit_r336_c16 bl[16] br[16] wl[336] vdd gnd cell_6t
Xbit_r337_c16 bl[16] br[16] wl[337] vdd gnd cell_6t
Xbit_r338_c16 bl[16] br[16] wl[338] vdd gnd cell_6t
Xbit_r339_c16 bl[16] br[16] wl[339] vdd gnd cell_6t
Xbit_r340_c16 bl[16] br[16] wl[340] vdd gnd cell_6t
Xbit_r341_c16 bl[16] br[16] wl[341] vdd gnd cell_6t
Xbit_r342_c16 bl[16] br[16] wl[342] vdd gnd cell_6t
Xbit_r343_c16 bl[16] br[16] wl[343] vdd gnd cell_6t
Xbit_r344_c16 bl[16] br[16] wl[344] vdd gnd cell_6t
Xbit_r345_c16 bl[16] br[16] wl[345] vdd gnd cell_6t
Xbit_r346_c16 bl[16] br[16] wl[346] vdd gnd cell_6t
Xbit_r347_c16 bl[16] br[16] wl[347] vdd gnd cell_6t
Xbit_r348_c16 bl[16] br[16] wl[348] vdd gnd cell_6t
Xbit_r349_c16 bl[16] br[16] wl[349] vdd gnd cell_6t
Xbit_r350_c16 bl[16] br[16] wl[350] vdd gnd cell_6t
Xbit_r351_c16 bl[16] br[16] wl[351] vdd gnd cell_6t
Xbit_r352_c16 bl[16] br[16] wl[352] vdd gnd cell_6t
Xbit_r353_c16 bl[16] br[16] wl[353] vdd gnd cell_6t
Xbit_r354_c16 bl[16] br[16] wl[354] vdd gnd cell_6t
Xbit_r355_c16 bl[16] br[16] wl[355] vdd gnd cell_6t
Xbit_r356_c16 bl[16] br[16] wl[356] vdd gnd cell_6t
Xbit_r357_c16 bl[16] br[16] wl[357] vdd gnd cell_6t
Xbit_r358_c16 bl[16] br[16] wl[358] vdd gnd cell_6t
Xbit_r359_c16 bl[16] br[16] wl[359] vdd gnd cell_6t
Xbit_r360_c16 bl[16] br[16] wl[360] vdd gnd cell_6t
Xbit_r361_c16 bl[16] br[16] wl[361] vdd gnd cell_6t
Xbit_r362_c16 bl[16] br[16] wl[362] vdd gnd cell_6t
Xbit_r363_c16 bl[16] br[16] wl[363] vdd gnd cell_6t
Xbit_r364_c16 bl[16] br[16] wl[364] vdd gnd cell_6t
Xbit_r365_c16 bl[16] br[16] wl[365] vdd gnd cell_6t
Xbit_r366_c16 bl[16] br[16] wl[366] vdd gnd cell_6t
Xbit_r367_c16 bl[16] br[16] wl[367] vdd gnd cell_6t
Xbit_r368_c16 bl[16] br[16] wl[368] vdd gnd cell_6t
Xbit_r369_c16 bl[16] br[16] wl[369] vdd gnd cell_6t
Xbit_r370_c16 bl[16] br[16] wl[370] vdd gnd cell_6t
Xbit_r371_c16 bl[16] br[16] wl[371] vdd gnd cell_6t
Xbit_r372_c16 bl[16] br[16] wl[372] vdd gnd cell_6t
Xbit_r373_c16 bl[16] br[16] wl[373] vdd gnd cell_6t
Xbit_r374_c16 bl[16] br[16] wl[374] vdd gnd cell_6t
Xbit_r375_c16 bl[16] br[16] wl[375] vdd gnd cell_6t
Xbit_r376_c16 bl[16] br[16] wl[376] vdd gnd cell_6t
Xbit_r377_c16 bl[16] br[16] wl[377] vdd gnd cell_6t
Xbit_r378_c16 bl[16] br[16] wl[378] vdd gnd cell_6t
Xbit_r379_c16 bl[16] br[16] wl[379] vdd gnd cell_6t
Xbit_r380_c16 bl[16] br[16] wl[380] vdd gnd cell_6t
Xbit_r381_c16 bl[16] br[16] wl[381] vdd gnd cell_6t
Xbit_r382_c16 bl[16] br[16] wl[382] vdd gnd cell_6t
Xbit_r383_c16 bl[16] br[16] wl[383] vdd gnd cell_6t
Xbit_r384_c16 bl[16] br[16] wl[384] vdd gnd cell_6t
Xbit_r385_c16 bl[16] br[16] wl[385] vdd gnd cell_6t
Xbit_r386_c16 bl[16] br[16] wl[386] vdd gnd cell_6t
Xbit_r387_c16 bl[16] br[16] wl[387] vdd gnd cell_6t
Xbit_r388_c16 bl[16] br[16] wl[388] vdd gnd cell_6t
Xbit_r389_c16 bl[16] br[16] wl[389] vdd gnd cell_6t
Xbit_r390_c16 bl[16] br[16] wl[390] vdd gnd cell_6t
Xbit_r391_c16 bl[16] br[16] wl[391] vdd gnd cell_6t
Xbit_r392_c16 bl[16] br[16] wl[392] vdd gnd cell_6t
Xbit_r393_c16 bl[16] br[16] wl[393] vdd gnd cell_6t
Xbit_r394_c16 bl[16] br[16] wl[394] vdd gnd cell_6t
Xbit_r395_c16 bl[16] br[16] wl[395] vdd gnd cell_6t
Xbit_r396_c16 bl[16] br[16] wl[396] vdd gnd cell_6t
Xbit_r397_c16 bl[16] br[16] wl[397] vdd gnd cell_6t
Xbit_r398_c16 bl[16] br[16] wl[398] vdd gnd cell_6t
Xbit_r399_c16 bl[16] br[16] wl[399] vdd gnd cell_6t
Xbit_r400_c16 bl[16] br[16] wl[400] vdd gnd cell_6t
Xbit_r401_c16 bl[16] br[16] wl[401] vdd gnd cell_6t
Xbit_r402_c16 bl[16] br[16] wl[402] vdd gnd cell_6t
Xbit_r403_c16 bl[16] br[16] wl[403] vdd gnd cell_6t
Xbit_r404_c16 bl[16] br[16] wl[404] vdd gnd cell_6t
Xbit_r405_c16 bl[16] br[16] wl[405] vdd gnd cell_6t
Xbit_r406_c16 bl[16] br[16] wl[406] vdd gnd cell_6t
Xbit_r407_c16 bl[16] br[16] wl[407] vdd gnd cell_6t
Xbit_r408_c16 bl[16] br[16] wl[408] vdd gnd cell_6t
Xbit_r409_c16 bl[16] br[16] wl[409] vdd gnd cell_6t
Xbit_r410_c16 bl[16] br[16] wl[410] vdd gnd cell_6t
Xbit_r411_c16 bl[16] br[16] wl[411] vdd gnd cell_6t
Xbit_r412_c16 bl[16] br[16] wl[412] vdd gnd cell_6t
Xbit_r413_c16 bl[16] br[16] wl[413] vdd gnd cell_6t
Xbit_r414_c16 bl[16] br[16] wl[414] vdd gnd cell_6t
Xbit_r415_c16 bl[16] br[16] wl[415] vdd gnd cell_6t
Xbit_r416_c16 bl[16] br[16] wl[416] vdd gnd cell_6t
Xbit_r417_c16 bl[16] br[16] wl[417] vdd gnd cell_6t
Xbit_r418_c16 bl[16] br[16] wl[418] vdd gnd cell_6t
Xbit_r419_c16 bl[16] br[16] wl[419] vdd gnd cell_6t
Xbit_r420_c16 bl[16] br[16] wl[420] vdd gnd cell_6t
Xbit_r421_c16 bl[16] br[16] wl[421] vdd gnd cell_6t
Xbit_r422_c16 bl[16] br[16] wl[422] vdd gnd cell_6t
Xbit_r423_c16 bl[16] br[16] wl[423] vdd gnd cell_6t
Xbit_r424_c16 bl[16] br[16] wl[424] vdd gnd cell_6t
Xbit_r425_c16 bl[16] br[16] wl[425] vdd gnd cell_6t
Xbit_r426_c16 bl[16] br[16] wl[426] vdd gnd cell_6t
Xbit_r427_c16 bl[16] br[16] wl[427] vdd gnd cell_6t
Xbit_r428_c16 bl[16] br[16] wl[428] vdd gnd cell_6t
Xbit_r429_c16 bl[16] br[16] wl[429] vdd gnd cell_6t
Xbit_r430_c16 bl[16] br[16] wl[430] vdd gnd cell_6t
Xbit_r431_c16 bl[16] br[16] wl[431] vdd gnd cell_6t
Xbit_r432_c16 bl[16] br[16] wl[432] vdd gnd cell_6t
Xbit_r433_c16 bl[16] br[16] wl[433] vdd gnd cell_6t
Xbit_r434_c16 bl[16] br[16] wl[434] vdd gnd cell_6t
Xbit_r435_c16 bl[16] br[16] wl[435] vdd gnd cell_6t
Xbit_r436_c16 bl[16] br[16] wl[436] vdd gnd cell_6t
Xbit_r437_c16 bl[16] br[16] wl[437] vdd gnd cell_6t
Xbit_r438_c16 bl[16] br[16] wl[438] vdd gnd cell_6t
Xbit_r439_c16 bl[16] br[16] wl[439] vdd gnd cell_6t
Xbit_r440_c16 bl[16] br[16] wl[440] vdd gnd cell_6t
Xbit_r441_c16 bl[16] br[16] wl[441] vdd gnd cell_6t
Xbit_r442_c16 bl[16] br[16] wl[442] vdd gnd cell_6t
Xbit_r443_c16 bl[16] br[16] wl[443] vdd gnd cell_6t
Xbit_r444_c16 bl[16] br[16] wl[444] vdd gnd cell_6t
Xbit_r445_c16 bl[16] br[16] wl[445] vdd gnd cell_6t
Xbit_r446_c16 bl[16] br[16] wl[446] vdd gnd cell_6t
Xbit_r447_c16 bl[16] br[16] wl[447] vdd gnd cell_6t
Xbit_r448_c16 bl[16] br[16] wl[448] vdd gnd cell_6t
Xbit_r449_c16 bl[16] br[16] wl[449] vdd gnd cell_6t
Xbit_r450_c16 bl[16] br[16] wl[450] vdd gnd cell_6t
Xbit_r451_c16 bl[16] br[16] wl[451] vdd gnd cell_6t
Xbit_r452_c16 bl[16] br[16] wl[452] vdd gnd cell_6t
Xbit_r453_c16 bl[16] br[16] wl[453] vdd gnd cell_6t
Xbit_r454_c16 bl[16] br[16] wl[454] vdd gnd cell_6t
Xbit_r455_c16 bl[16] br[16] wl[455] vdd gnd cell_6t
Xbit_r456_c16 bl[16] br[16] wl[456] vdd gnd cell_6t
Xbit_r457_c16 bl[16] br[16] wl[457] vdd gnd cell_6t
Xbit_r458_c16 bl[16] br[16] wl[458] vdd gnd cell_6t
Xbit_r459_c16 bl[16] br[16] wl[459] vdd gnd cell_6t
Xbit_r460_c16 bl[16] br[16] wl[460] vdd gnd cell_6t
Xbit_r461_c16 bl[16] br[16] wl[461] vdd gnd cell_6t
Xbit_r462_c16 bl[16] br[16] wl[462] vdd gnd cell_6t
Xbit_r463_c16 bl[16] br[16] wl[463] vdd gnd cell_6t
Xbit_r464_c16 bl[16] br[16] wl[464] vdd gnd cell_6t
Xbit_r465_c16 bl[16] br[16] wl[465] vdd gnd cell_6t
Xbit_r466_c16 bl[16] br[16] wl[466] vdd gnd cell_6t
Xbit_r467_c16 bl[16] br[16] wl[467] vdd gnd cell_6t
Xbit_r468_c16 bl[16] br[16] wl[468] vdd gnd cell_6t
Xbit_r469_c16 bl[16] br[16] wl[469] vdd gnd cell_6t
Xbit_r470_c16 bl[16] br[16] wl[470] vdd gnd cell_6t
Xbit_r471_c16 bl[16] br[16] wl[471] vdd gnd cell_6t
Xbit_r472_c16 bl[16] br[16] wl[472] vdd gnd cell_6t
Xbit_r473_c16 bl[16] br[16] wl[473] vdd gnd cell_6t
Xbit_r474_c16 bl[16] br[16] wl[474] vdd gnd cell_6t
Xbit_r475_c16 bl[16] br[16] wl[475] vdd gnd cell_6t
Xbit_r476_c16 bl[16] br[16] wl[476] vdd gnd cell_6t
Xbit_r477_c16 bl[16] br[16] wl[477] vdd gnd cell_6t
Xbit_r478_c16 bl[16] br[16] wl[478] vdd gnd cell_6t
Xbit_r479_c16 bl[16] br[16] wl[479] vdd gnd cell_6t
Xbit_r480_c16 bl[16] br[16] wl[480] vdd gnd cell_6t
Xbit_r481_c16 bl[16] br[16] wl[481] vdd gnd cell_6t
Xbit_r482_c16 bl[16] br[16] wl[482] vdd gnd cell_6t
Xbit_r483_c16 bl[16] br[16] wl[483] vdd gnd cell_6t
Xbit_r484_c16 bl[16] br[16] wl[484] vdd gnd cell_6t
Xbit_r485_c16 bl[16] br[16] wl[485] vdd gnd cell_6t
Xbit_r486_c16 bl[16] br[16] wl[486] vdd gnd cell_6t
Xbit_r487_c16 bl[16] br[16] wl[487] vdd gnd cell_6t
Xbit_r488_c16 bl[16] br[16] wl[488] vdd gnd cell_6t
Xbit_r489_c16 bl[16] br[16] wl[489] vdd gnd cell_6t
Xbit_r490_c16 bl[16] br[16] wl[490] vdd gnd cell_6t
Xbit_r491_c16 bl[16] br[16] wl[491] vdd gnd cell_6t
Xbit_r492_c16 bl[16] br[16] wl[492] vdd gnd cell_6t
Xbit_r493_c16 bl[16] br[16] wl[493] vdd gnd cell_6t
Xbit_r494_c16 bl[16] br[16] wl[494] vdd gnd cell_6t
Xbit_r495_c16 bl[16] br[16] wl[495] vdd gnd cell_6t
Xbit_r496_c16 bl[16] br[16] wl[496] vdd gnd cell_6t
Xbit_r497_c16 bl[16] br[16] wl[497] vdd gnd cell_6t
Xbit_r498_c16 bl[16] br[16] wl[498] vdd gnd cell_6t
Xbit_r499_c16 bl[16] br[16] wl[499] vdd gnd cell_6t
Xbit_r500_c16 bl[16] br[16] wl[500] vdd gnd cell_6t
Xbit_r501_c16 bl[16] br[16] wl[501] vdd gnd cell_6t
Xbit_r502_c16 bl[16] br[16] wl[502] vdd gnd cell_6t
Xbit_r503_c16 bl[16] br[16] wl[503] vdd gnd cell_6t
Xbit_r504_c16 bl[16] br[16] wl[504] vdd gnd cell_6t
Xbit_r505_c16 bl[16] br[16] wl[505] vdd gnd cell_6t
Xbit_r506_c16 bl[16] br[16] wl[506] vdd gnd cell_6t
Xbit_r507_c16 bl[16] br[16] wl[507] vdd gnd cell_6t
Xbit_r508_c16 bl[16] br[16] wl[508] vdd gnd cell_6t
Xbit_r509_c16 bl[16] br[16] wl[509] vdd gnd cell_6t
Xbit_r510_c16 bl[16] br[16] wl[510] vdd gnd cell_6t
Xbit_r511_c16 bl[16] br[16] wl[511] vdd gnd cell_6t
Xbit_r0_c17 bl[17] br[17] wl[0] vdd gnd cell_6t
Xbit_r1_c17 bl[17] br[17] wl[1] vdd gnd cell_6t
Xbit_r2_c17 bl[17] br[17] wl[2] vdd gnd cell_6t
Xbit_r3_c17 bl[17] br[17] wl[3] vdd gnd cell_6t
Xbit_r4_c17 bl[17] br[17] wl[4] vdd gnd cell_6t
Xbit_r5_c17 bl[17] br[17] wl[5] vdd gnd cell_6t
Xbit_r6_c17 bl[17] br[17] wl[6] vdd gnd cell_6t
Xbit_r7_c17 bl[17] br[17] wl[7] vdd gnd cell_6t
Xbit_r8_c17 bl[17] br[17] wl[8] vdd gnd cell_6t
Xbit_r9_c17 bl[17] br[17] wl[9] vdd gnd cell_6t
Xbit_r10_c17 bl[17] br[17] wl[10] vdd gnd cell_6t
Xbit_r11_c17 bl[17] br[17] wl[11] vdd gnd cell_6t
Xbit_r12_c17 bl[17] br[17] wl[12] vdd gnd cell_6t
Xbit_r13_c17 bl[17] br[17] wl[13] vdd gnd cell_6t
Xbit_r14_c17 bl[17] br[17] wl[14] vdd gnd cell_6t
Xbit_r15_c17 bl[17] br[17] wl[15] vdd gnd cell_6t
Xbit_r16_c17 bl[17] br[17] wl[16] vdd gnd cell_6t
Xbit_r17_c17 bl[17] br[17] wl[17] vdd gnd cell_6t
Xbit_r18_c17 bl[17] br[17] wl[18] vdd gnd cell_6t
Xbit_r19_c17 bl[17] br[17] wl[19] vdd gnd cell_6t
Xbit_r20_c17 bl[17] br[17] wl[20] vdd gnd cell_6t
Xbit_r21_c17 bl[17] br[17] wl[21] vdd gnd cell_6t
Xbit_r22_c17 bl[17] br[17] wl[22] vdd gnd cell_6t
Xbit_r23_c17 bl[17] br[17] wl[23] vdd gnd cell_6t
Xbit_r24_c17 bl[17] br[17] wl[24] vdd gnd cell_6t
Xbit_r25_c17 bl[17] br[17] wl[25] vdd gnd cell_6t
Xbit_r26_c17 bl[17] br[17] wl[26] vdd gnd cell_6t
Xbit_r27_c17 bl[17] br[17] wl[27] vdd gnd cell_6t
Xbit_r28_c17 bl[17] br[17] wl[28] vdd gnd cell_6t
Xbit_r29_c17 bl[17] br[17] wl[29] vdd gnd cell_6t
Xbit_r30_c17 bl[17] br[17] wl[30] vdd gnd cell_6t
Xbit_r31_c17 bl[17] br[17] wl[31] vdd gnd cell_6t
Xbit_r32_c17 bl[17] br[17] wl[32] vdd gnd cell_6t
Xbit_r33_c17 bl[17] br[17] wl[33] vdd gnd cell_6t
Xbit_r34_c17 bl[17] br[17] wl[34] vdd gnd cell_6t
Xbit_r35_c17 bl[17] br[17] wl[35] vdd gnd cell_6t
Xbit_r36_c17 bl[17] br[17] wl[36] vdd gnd cell_6t
Xbit_r37_c17 bl[17] br[17] wl[37] vdd gnd cell_6t
Xbit_r38_c17 bl[17] br[17] wl[38] vdd gnd cell_6t
Xbit_r39_c17 bl[17] br[17] wl[39] vdd gnd cell_6t
Xbit_r40_c17 bl[17] br[17] wl[40] vdd gnd cell_6t
Xbit_r41_c17 bl[17] br[17] wl[41] vdd gnd cell_6t
Xbit_r42_c17 bl[17] br[17] wl[42] vdd gnd cell_6t
Xbit_r43_c17 bl[17] br[17] wl[43] vdd gnd cell_6t
Xbit_r44_c17 bl[17] br[17] wl[44] vdd gnd cell_6t
Xbit_r45_c17 bl[17] br[17] wl[45] vdd gnd cell_6t
Xbit_r46_c17 bl[17] br[17] wl[46] vdd gnd cell_6t
Xbit_r47_c17 bl[17] br[17] wl[47] vdd gnd cell_6t
Xbit_r48_c17 bl[17] br[17] wl[48] vdd gnd cell_6t
Xbit_r49_c17 bl[17] br[17] wl[49] vdd gnd cell_6t
Xbit_r50_c17 bl[17] br[17] wl[50] vdd gnd cell_6t
Xbit_r51_c17 bl[17] br[17] wl[51] vdd gnd cell_6t
Xbit_r52_c17 bl[17] br[17] wl[52] vdd gnd cell_6t
Xbit_r53_c17 bl[17] br[17] wl[53] vdd gnd cell_6t
Xbit_r54_c17 bl[17] br[17] wl[54] vdd gnd cell_6t
Xbit_r55_c17 bl[17] br[17] wl[55] vdd gnd cell_6t
Xbit_r56_c17 bl[17] br[17] wl[56] vdd gnd cell_6t
Xbit_r57_c17 bl[17] br[17] wl[57] vdd gnd cell_6t
Xbit_r58_c17 bl[17] br[17] wl[58] vdd gnd cell_6t
Xbit_r59_c17 bl[17] br[17] wl[59] vdd gnd cell_6t
Xbit_r60_c17 bl[17] br[17] wl[60] vdd gnd cell_6t
Xbit_r61_c17 bl[17] br[17] wl[61] vdd gnd cell_6t
Xbit_r62_c17 bl[17] br[17] wl[62] vdd gnd cell_6t
Xbit_r63_c17 bl[17] br[17] wl[63] vdd gnd cell_6t
Xbit_r64_c17 bl[17] br[17] wl[64] vdd gnd cell_6t
Xbit_r65_c17 bl[17] br[17] wl[65] vdd gnd cell_6t
Xbit_r66_c17 bl[17] br[17] wl[66] vdd gnd cell_6t
Xbit_r67_c17 bl[17] br[17] wl[67] vdd gnd cell_6t
Xbit_r68_c17 bl[17] br[17] wl[68] vdd gnd cell_6t
Xbit_r69_c17 bl[17] br[17] wl[69] vdd gnd cell_6t
Xbit_r70_c17 bl[17] br[17] wl[70] vdd gnd cell_6t
Xbit_r71_c17 bl[17] br[17] wl[71] vdd gnd cell_6t
Xbit_r72_c17 bl[17] br[17] wl[72] vdd gnd cell_6t
Xbit_r73_c17 bl[17] br[17] wl[73] vdd gnd cell_6t
Xbit_r74_c17 bl[17] br[17] wl[74] vdd gnd cell_6t
Xbit_r75_c17 bl[17] br[17] wl[75] vdd gnd cell_6t
Xbit_r76_c17 bl[17] br[17] wl[76] vdd gnd cell_6t
Xbit_r77_c17 bl[17] br[17] wl[77] vdd gnd cell_6t
Xbit_r78_c17 bl[17] br[17] wl[78] vdd gnd cell_6t
Xbit_r79_c17 bl[17] br[17] wl[79] vdd gnd cell_6t
Xbit_r80_c17 bl[17] br[17] wl[80] vdd gnd cell_6t
Xbit_r81_c17 bl[17] br[17] wl[81] vdd gnd cell_6t
Xbit_r82_c17 bl[17] br[17] wl[82] vdd gnd cell_6t
Xbit_r83_c17 bl[17] br[17] wl[83] vdd gnd cell_6t
Xbit_r84_c17 bl[17] br[17] wl[84] vdd gnd cell_6t
Xbit_r85_c17 bl[17] br[17] wl[85] vdd gnd cell_6t
Xbit_r86_c17 bl[17] br[17] wl[86] vdd gnd cell_6t
Xbit_r87_c17 bl[17] br[17] wl[87] vdd gnd cell_6t
Xbit_r88_c17 bl[17] br[17] wl[88] vdd gnd cell_6t
Xbit_r89_c17 bl[17] br[17] wl[89] vdd gnd cell_6t
Xbit_r90_c17 bl[17] br[17] wl[90] vdd gnd cell_6t
Xbit_r91_c17 bl[17] br[17] wl[91] vdd gnd cell_6t
Xbit_r92_c17 bl[17] br[17] wl[92] vdd gnd cell_6t
Xbit_r93_c17 bl[17] br[17] wl[93] vdd gnd cell_6t
Xbit_r94_c17 bl[17] br[17] wl[94] vdd gnd cell_6t
Xbit_r95_c17 bl[17] br[17] wl[95] vdd gnd cell_6t
Xbit_r96_c17 bl[17] br[17] wl[96] vdd gnd cell_6t
Xbit_r97_c17 bl[17] br[17] wl[97] vdd gnd cell_6t
Xbit_r98_c17 bl[17] br[17] wl[98] vdd gnd cell_6t
Xbit_r99_c17 bl[17] br[17] wl[99] vdd gnd cell_6t
Xbit_r100_c17 bl[17] br[17] wl[100] vdd gnd cell_6t
Xbit_r101_c17 bl[17] br[17] wl[101] vdd gnd cell_6t
Xbit_r102_c17 bl[17] br[17] wl[102] vdd gnd cell_6t
Xbit_r103_c17 bl[17] br[17] wl[103] vdd gnd cell_6t
Xbit_r104_c17 bl[17] br[17] wl[104] vdd gnd cell_6t
Xbit_r105_c17 bl[17] br[17] wl[105] vdd gnd cell_6t
Xbit_r106_c17 bl[17] br[17] wl[106] vdd gnd cell_6t
Xbit_r107_c17 bl[17] br[17] wl[107] vdd gnd cell_6t
Xbit_r108_c17 bl[17] br[17] wl[108] vdd gnd cell_6t
Xbit_r109_c17 bl[17] br[17] wl[109] vdd gnd cell_6t
Xbit_r110_c17 bl[17] br[17] wl[110] vdd gnd cell_6t
Xbit_r111_c17 bl[17] br[17] wl[111] vdd gnd cell_6t
Xbit_r112_c17 bl[17] br[17] wl[112] vdd gnd cell_6t
Xbit_r113_c17 bl[17] br[17] wl[113] vdd gnd cell_6t
Xbit_r114_c17 bl[17] br[17] wl[114] vdd gnd cell_6t
Xbit_r115_c17 bl[17] br[17] wl[115] vdd gnd cell_6t
Xbit_r116_c17 bl[17] br[17] wl[116] vdd gnd cell_6t
Xbit_r117_c17 bl[17] br[17] wl[117] vdd gnd cell_6t
Xbit_r118_c17 bl[17] br[17] wl[118] vdd gnd cell_6t
Xbit_r119_c17 bl[17] br[17] wl[119] vdd gnd cell_6t
Xbit_r120_c17 bl[17] br[17] wl[120] vdd gnd cell_6t
Xbit_r121_c17 bl[17] br[17] wl[121] vdd gnd cell_6t
Xbit_r122_c17 bl[17] br[17] wl[122] vdd gnd cell_6t
Xbit_r123_c17 bl[17] br[17] wl[123] vdd gnd cell_6t
Xbit_r124_c17 bl[17] br[17] wl[124] vdd gnd cell_6t
Xbit_r125_c17 bl[17] br[17] wl[125] vdd gnd cell_6t
Xbit_r126_c17 bl[17] br[17] wl[126] vdd gnd cell_6t
Xbit_r127_c17 bl[17] br[17] wl[127] vdd gnd cell_6t
Xbit_r128_c17 bl[17] br[17] wl[128] vdd gnd cell_6t
Xbit_r129_c17 bl[17] br[17] wl[129] vdd gnd cell_6t
Xbit_r130_c17 bl[17] br[17] wl[130] vdd gnd cell_6t
Xbit_r131_c17 bl[17] br[17] wl[131] vdd gnd cell_6t
Xbit_r132_c17 bl[17] br[17] wl[132] vdd gnd cell_6t
Xbit_r133_c17 bl[17] br[17] wl[133] vdd gnd cell_6t
Xbit_r134_c17 bl[17] br[17] wl[134] vdd gnd cell_6t
Xbit_r135_c17 bl[17] br[17] wl[135] vdd gnd cell_6t
Xbit_r136_c17 bl[17] br[17] wl[136] vdd gnd cell_6t
Xbit_r137_c17 bl[17] br[17] wl[137] vdd gnd cell_6t
Xbit_r138_c17 bl[17] br[17] wl[138] vdd gnd cell_6t
Xbit_r139_c17 bl[17] br[17] wl[139] vdd gnd cell_6t
Xbit_r140_c17 bl[17] br[17] wl[140] vdd gnd cell_6t
Xbit_r141_c17 bl[17] br[17] wl[141] vdd gnd cell_6t
Xbit_r142_c17 bl[17] br[17] wl[142] vdd gnd cell_6t
Xbit_r143_c17 bl[17] br[17] wl[143] vdd gnd cell_6t
Xbit_r144_c17 bl[17] br[17] wl[144] vdd gnd cell_6t
Xbit_r145_c17 bl[17] br[17] wl[145] vdd gnd cell_6t
Xbit_r146_c17 bl[17] br[17] wl[146] vdd gnd cell_6t
Xbit_r147_c17 bl[17] br[17] wl[147] vdd gnd cell_6t
Xbit_r148_c17 bl[17] br[17] wl[148] vdd gnd cell_6t
Xbit_r149_c17 bl[17] br[17] wl[149] vdd gnd cell_6t
Xbit_r150_c17 bl[17] br[17] wl[150] vdd gnd cell_6t
Xbit_r151_c17 bl[17] br[17] wl[151] vdd gnd cell_6t
Xbit_r152_c17 bl[17] br[17] wl[152] vdd gnd cell_6t
Xbit_r153_c17 bl[17] br[17] wl[153] vdd gnd cell_6t
Xbit_r154_c17 bl[17] br[17] wl[154] vdd gnd cell_6t
Xbit_r155_c17 bl[17] br[17] wl[155] vdd gnd cell_6t
Xbit_r156_c17 bl[17] br[17] wl[156] vdd gnd cell_6t
Xbit_r157_c17 bl[17] br[17] wl[157] vdd gnd cell_6t
Xbit_r158_c17 bl[17] br[17] wl[158] vdd gnd cell_6t
Xbit_r159_c17 bl[17] br[17] wl[159] vdd gnd cell_6t
Xbit_r160_c17 bl[17] br[17] wl[160] vdd gnd cell_6t
Xbit_r161_c17 bl[17] br[17] wl[161] vdd gnd cell_6t
Xbit_r162_c17 bl[17] br[17] wl[162] vdd gnd cell_6t
Xbit_r163_c17 bl[17] br[17] wl[163] vdd gnd cell_6t
Xbit_r164_c17 bl[17] br[17] wl[164] vdd gnd cell_6t
Xbit_r165_c17 bl[17] br[17] wl[165] vdd gnd cell_6t
Xbit_r166_c17 bl[17] br[17] wl[166] vdd gnd cell_6t
Xbit_r167_c17 bl[17] br[17] wl[167] vdd gnd cell_6t
Xbit_r168_c17 bl[17] br[17] wl[168] vdd gnd cell_6t
Xbit_r169_c17 bl[17] br[17] wl[169] vdd gnd cell_6t
Xbit_r170_c17 bl[17] br[17] wl[170] vdd gnd cell_6t
Xbit_r171_c17 bl[17] br[17] wl[171] vdd gnd cell_6t
Xbit_r172_c17 bl[17] br[17] wl[172] vdd gnd cell_6t
Xbit_r173_c17 bl[17] br[17] wl[173] vdd gnd cell_6t
Xbit_r174_c17 bl[17] br[17] wl[174] vdd gnd cell_6t
Xbit_r175_c17 bl[17] br[17] wl[175] vdd gnd cell_6t
Xbit_r176_c17 bl[17] br[17] wl[176] vdd gnd cell_6t
Xbit_r177_c17 bl[17] br[17] wl[177] vdd gnd cell_6t
Xbit_r178_c17 bl[17] br[17] wl[178] vdd gnd cell_6t
Xbit_r179_c17 bl[17] br[17] wl[179] vdd gnd cell_6t
Xbit_r180_c17 bl[17] br[17] wl[180] vdd gnd cell_6t
Xbit_r181_c17 bl[17] br[17] wl[181] vdd gnd cell_6t
Xbit_r182_c17 bl[17] br[17] wl[182] vdd gnd cell_6t
Xbit_r183_c17 bl[17] br[17] wl[183] vdd gnd cell_6t
Xbit_r184_c17 bl[17] br[17] wl[184] vdd gnd cell_6t
Xbit_r185_c17 bl[17] br[17] wl[185] vdd gnd cell_6t
Xbit_r186_c17 bl[17] br[17] wl[186] vdd gnd cell_6t
Xbit_r187_c17 bl[17] br[17] wl[187] vdd gnd cell_6t
Xbit_r188_c17 bl[17] br[17] wl[188] vdd gnd cell_6t
Xbit_r189_c17 bl[17] br[17] wl[189] vdd gnd cell_6t
Xbit_r190_c17 bl[17] br[17] wl[190] vdd gnd cell_6t
Xbit_r191_c17 bl[17] br[17] wl[191] vdd gnd cell_6t
Xbit_r192_c17 bl[17] br[17] wl[192] vdd gnd cell_6t
Xbit_r193_c17 bl[17] br[17] wl[193] vdd gnd cell_6t
Xbit_r194_c17 bl[17] br[17] wl[194] vdd gnd cell_6t
Xbit_r195_c17 bl[17] br[17] wl[195] vdd gnd cell_6t
Xbit_r196_c17 bl[17] br[17] wl[196] vdd gnd cell_6t
Xbit_r197_c17 bl[17] br[17] wl[197] vdd gnd cell_6t
Xbit_r198_c17 bl[17] br[17] wl[198] vdd gnd cell_6t
Xbit_r199_c17 bl[17] br[17] wl[199] vdd gnd cell_6t
Xbit_r200_c17 bl[17] br[17] wl[200] vdd gnd cell_6t
Xbit_r201_c17 bl[17] br[17] wl[201] vdd gnd cell_6t
Xbit_r202_c17 bl[17] br[17] wl[202] vdd gnd cell_6t
Xbit_r203_c17 bl[17] br[17] wl[203] vdd gnd cell_6t
Xbit_r204_c17 bl[17] br[17] wl[204] vdd gnd cell_6t
Xbit_r205_c17 bl[17] br[17] wl[205] vdd gnd cell_6t
Xbit_r206_c17 bl[17] br[17] wl[206] vdd gnd cell_6t
Xbit_r207_c17 bl[17] br[17] wl[207] vdd gnd cell_6t
Xbit_r208_c17 bl[17] br[17] wl[208] vdd gnd cell_6t
Xbit_r209_c17 bl[17] br[17] wl[209] vdd gnd cell_6t
Xbit_r210_c17 bl[17] br[17] wl[210] vdd gnd cell_6t
Xbit_r211_c17 bl[17] br[17] wl[211] vdd gnd cell_6t
Xbit_r212_c17 bl[17] br[17] wl[212] vdd gnd cell_6t
Xbit_r213_c17 bl[17] br[17] wl[213] vdd gnd cell_6t
Xbit_r214_c17 bl[17] br[17] wl[214] vdd gnd cell_6t
Xbit_r215_c17 bl[17] br[17] wl[215] vdd gnd cell_6t
Xbit_r216_c17 bl[17] br[17] wl[216] vdd gnd cell_6t
Xbit_r217_c17 bl[17] br[17] wl[217] vdd gnd cell_6t
Xbit_r218_c17 bl[17] br[17] wl[218] vdd gnd cell_6t
Xbit_r219_c17 bl[17] br[17] wl[219] vdd gnd cell_6t
Xbit_r220_c17 bl[17] br[17] wl[220] vdd gnd cell_6t
Xbit_r221_c17 bl[17] br[17] wl[221] vdd gnd cell_6t
Xbit_r222_c17 bl[17] br[17] wl[222] vdd gnd cell_6t
Xbit_r223_c17 bl[17] br[17] wl[223] vdd gnd cell_6t
Xbit_r224_c17 bl[17] br[17] wl[224] vdd gnd cell_6t
Xbit_r225_c17 bl[17] br[17] wl[225] vdd gnd cell_6t
Xbit_r226_c17 bl[17] br[17] wl[226] vdd gnd cell_6t
Xbit_r227_c17 bl[17] br[17] wl[227] vdd gnd cell_6t
Xbit_r228_c17 bl[17] br[17] wl[228] vdd gnd cell_6t
Xbit_r229_c17 bl[17] br[17] wl[229] vdd gnd cell_6t
Xbit_r230_c17 bl[17] br[17] wl[230] vdd gnd cell_6t
Xbit_r231_c17 bl[17] br[17] wl[231] vdd gnd cell_6t
Xbit_r232_c17 bl[17] br[17] wl[232] vdd gnd cell_6t
Xbit_r233_c17 bl[17] br[17] wl[233] vdd gnd cell_6t
Xbit_r234_c17 bl[17] br[17] wl[234] vdd gnd cell_6t
Xbit_r235_c17 bl[17] br[17] wl[235] vdd gnd cell_6t
Xbit_r236_c17 bl[17] br[17] wl[236] vdd gnd cell_6t
Xbit_r237_c17 bl[17] br[17] wl[237] vdd gnd cell_6t
Xbit_r238_c17 bl[17] br[17] wl[238] vdd gnd cell_6t
Xbit_r239_c17 bl[17] br[17] wl[239] vdd gnd cell_6t
Xbit_r240_c17 bl[17] br[17] wl[240] vdd gnd cell_6t
Xbit_r241_c17 bl[17] br[17] wl[241] vdd gnd cell_6t
Xbit_r242_c17 bl[17] br[17] wl[242] vdd gnd cell_6t
Xbit_r243_c17 bl[17] br[17] wl[243] vdd gnd cell_6t
Xbit_r244_c17 bl[17] br[17] wl[244] vdd gnd cell_6t
Xbit_r245_c17 bl[17] br[17] wl[245] vdd gnd cell_6t
Xbit_r246_c17 bl[17] br[17] wl[246] vdd gnd cell_6t
Xbit_r247_c17 bl[17] br[17] wl[247] vdd gnd cell_6t
Xbit_r248_c17 bl[17] br[17] wl[248] vdd gnd cell_6t
Xbit_r249_c17 bl[17] br[17] wl[249] vdd gnd cell_6t
Xbit_r250_c17 bl[17] br[17] wl[250] vdd gnd cell_6t
Xbit_r251_c17 bl[17] br[17] wl[251] vdd gnd cell_6t
Xbit_r252_c17 bl[17] br[17] wl[252] vdd gnd cell_6t
Xbit_r253_c17 bl[17] br[17] wl[253] vdd gnd cell_6t
Xbit_r254_c17 bl[17] br[17] wl[254] vdd gnd cell_6t
Xbit_r255_c17 bl[17] br[17] wl[255] vdd gnd cell_6t
Xbit_r256_c17 bl[17] br[17] wl[256] vdd gnd cell_6t
Xbit_r257_c17 bl[17] br[17] wl[257] vdd gnd cell_6t
Xbit_r258_c17 bl[17] br[17] wl[258] vdd gnd cell_6t
Xbit_r259_c17 bl[17] br[17] wl[259] vdd gnd cell_6t
Xbit_r260_c17 bl[17] br[17] wl[260] vdd gnd cell_6t
Xbit_r261_c17 bl[17] br[17] wl[261] vdd gnd cell_6t
Xbit_r262_c17 bl[17] br[17] wl[262] vdd gnd cell_6t
Xbit_r263_c17 bl[17] br[17] wl[263] vdd gnd cell_6t
Xbit_r264_c17 bl[17] br[17] wl[264] vdd gnd cell_6t
Xbit_r265_c17 bl[17] br[17] wl[265] vdd gnd cell_6t
Xbit_r266_c17 bl[17] br[17] wl[266] vdd gnd cell_6t
Xbit_r267_c17 bl[17] br[17] wl[267] vdd gnd cell_6t
Xbit_r268_c17 bl[17] br[17] wl[268] vdd gnd cell_6t
Xbit_r269_c17 bl[17] br[17] wl[269] vdd gnd cell_6t
Xbit_r270_c17 bl[17] br[17] wl[270] vdd gnd cell_6t
Xbit_r271_c17 bl[17] br[17] wl[271] vdd gnd cell_6t
Xbit_r272_c17 bl[17] br[17] wl[272] vdd gnd cell_6t
Xbit_r273_c17 bl[17] br[17] wl[273] vdd gnd cell_6t
Xbit_r274_c17 bl[17] br[17] wl[274] vdd gnd cell_6t
Xbit_r275_c17 bl[17] br[17] wl[275] vdd gnd cell_6t
Xbit_r276_c17 bl[17] br[17] wl[276] vdd gnd cell_6t
Xbit_r277_c17 bl[17] br[17] wl[277] vdd gnd cell_6t
Xbit_r278_c17 bl[17] br[17] wl[278] vdd gnd cell_6t
Xbit_r279_c17 bl[17] br[17] wl[279] vdd gnd cell_6t
Xbit_r280_c17 bl[17] br[17] wl[280] vdd gnd cell_6t
Xbit_r281_c17 bl[17] br[17] wl[281] vdd gnd cell_6t
Xbit_r282_c17 bl[17] br[17] wl[282] vdd gnd cell_6t
Xbit_r283_c17 bl[17] br[17] wl[283] vdd gnd cell_6t
Xbit_r284_c17 bl[17] br[17] wl[284] vdd gnd cell_6t
Xbit_r285_c17 bl[17] br[17] wl[285] vdd gnd cell_6t
Xbit_r286_c17 bl[17] br[17] wl[286] vdd gnd cell_6t
Xbit_r287_c17 bl[17] br[17] wl[287] vdd gnd cell_6t
Xbit_r288_c17 bl[17] br[17] wl[288] vdd gnd cell_6t
Xbit_r289_c17 bl[17] br[17] wl[289] vdd gnd cell_6t
Xbit_r290_c17 bl[17] br[17] wl[290] vdd gnd cell_6t
Xbit_r291_c17 bl[17] br[17] wl[291] vdd gnd cell_6t
Xbit_r292_c17 bl[17] br[17] wl[292] vdd gnd cell_6t
Xbit_r293_c17 bl[17] br[17] wl[293] vdd gnd cell_6t
Xbit_r294_c17 bl[17] br[17] wl[294] vdd gnd cell_6t
Xbit_r295_c17 bl[17] br[17] wl[295] vdd gnd cell_6t
Xbit_r296_c17 bl[17] br[17] wl[296] vdd gnd cell_6t
Xbit_r297_c17 bl[17] br[17] wl[297] vdd gnd cell_6t
Xbit_r298_c17 bl[17] br[17] wl[298] vdd gnd cell_6t
Xbit_r299_c17 bl[17] br[17] wl[299] vdd gnd cell_6t
Xbit_r300_c17 bl[17] br[17] wl[300] vdd gnd cell_6t
Xbit_r301_c17 bl[17] br[17] wl[301] vdd gnd cell_6t
Xbit_r302_c17 bl[17] br[17] wl[302] vdd gnd cell_6t
Xbit_r303_c17 bl[17] br[17] wl[303] vdd gnd cell_6t
Xbit_r304_c17 bl[17] br[17] wl[304] vdd gnd cell_6t
Xbit_r305_c17 bl[17] br[17] wl[305] vdd gnd cell_6t
Xbit_r306_c17 bl[17] br[17] wl[306] vdd gnd cell_6t
Xbit_r307_c17 bl[17] br[17] wl[307] vdd gnd cell_6t
Xbit_r308_c17 bl[17] br[17] wl[308] vdd gnd cell_6t
Xbit_r309_c17 bl[17] br[17] wl[309] vdd gnd cell_6t
Xbit_r310_c17 bl[17] br[17] wl[310] vdd gnd cell_6t
Xbit_r311_c17 bl[17] br[17] wl[311] vdd gnd cell_6t
Xbit_r312_c17 bl[17] br[17] wl[312] vdd gnd cell_6t
Xbit_r313_c17 bl[17] br[17] wl[313] vdd gnd cell_6t
Xbit_r314_c17 bl[17] br[17] wl[314] vdd gnd cell_6t
Xbit_r315_c17 bl[17] br[17] wl[315] vdd gnd cell_6t
Xbit_r316_c17 bl[17] br[17] wl[316] vdd gnd cell_6t
Xbit_r317_c17 bl[17] br[17] wl[317] vdd gnd cell_6t
Xbit_r318_c17 bl[17] br[17] wl[318] vdd gnd cell_6t
Xbit_r319_c17 bl[17] br[17] wl[319] vdd gnd cell_6t
Xbit_r320_c17 bl[17] br[17] wl[320] vdd gnd cell_6t
Xbit_r321_c17 bl[17] br[17] wl[321] vdd gnd cell_6t
Xbit_r322_c17 bl[17] br[17] wl[322] vdd gnd cell_6t
Xbit_r323_c17 bl[17] br[17] wl[323] vdd gnd cell_6t
Xbit_r324_c17 bl[17] br[17] wl[324] vdd gnd cell_6t
Xbit_r325_c17 bl[17] br[17] wl[325] vdd gnd cell_6t
Xbit_r326_c17 bl[17] br[17] wl[326] vdd gnd cell_6t
Xbit_r327_c17 bl[17] br[17] wl[327] vdd gnd cell_6t
Xbit_r328_c17 bl[17] br[17] wl[328] vdd gnd cell_6t
Xbit_r329_c17 bl[17] br[17] wl[329] vdd gnd cell_6t
Xbit_r330_c17 bl[17] br[17] wl[330] vdd gnd cell_6t
Xbit_r331_c17 bl[17] br[17] wl[331] vdd gnd cell_6t
Xbit_r332_c17 bl[17] br[17] wl[332] vdd gnd cell_6t
Xbit_r333_c17 bl[17] br[17] wl[333] vdd gnd cell_6t
Xbit_r334_c17 bl[17] br[17] wl[334] vdd gnd cell_6t
Xbit_r335_c17 bl[17] br[17] wl[335] vdd gnd cell_6t
Xbit_r336_c17 bl[17] br[17] wl[336] vdd gnd cell_6t
Xbit_r337_c17 bl[17] br[17] wl[337] vdd gnd cell_6t
Xbit_r338_c17 bl[17] br[17] wl[338] vdd gnd cell_6t
Xbit_r339_c17 bl[17] br[17] wl[339] vdd gnd cell_6t
Xbit_r340_c17 bl[17] br[17] wl[340] vdd gnd cell_6t
Xbit_r341_c17 bl[17] br[17] wl[341] vdd gnd cell_6t
Xbit_r342_c17 bl[17] br[17] wl[342] vdd gnd cell_6t
Xbit_r343_c17 bl[17] br[17] wl[343] vdd gnd cell_6t
Xbit_r344_c17 bl[17] br[17] wl[344] vdd gnd cell_6t
Xbit_r345_c17 bl[17] br[17] wl[345] vdd gnd cell_6t
Xbit_r346_c17 bl[17] br[17] wl[346] vdd gnd cell_6t
Xbit_r347_c17 bl[17] br[17] wl[347] vdd gnd cell_6t
Xbit_r348_c17 bl[17] br[17] wl[348] vdd gnd cell_6t
Xbit_r349_c17 bl[17] br[17] wl[349] vdd gnd cell_6t
Xbit_r350_c17 bl[17] br[17] wl[350] vdd gnd cell_6t
Xbit_r351_c17 bl[17] br[17] wl[351] vdd gnd cell_6t
Xbit_r352_c17 bl[17] br[17] wl[352] vdd gnd cell_6t
Xbit_r353_c17 bl[17] br[17] wl[353] vdd gnd cell_6t
Xbit_r354_c17 bl[17] br[17] wl[354] vdd gnd cell_6t
Xbit_r355_c17 bl[17] br[17] wl[355] vdd gnd cell_6t
Xbit_r356_c17 bl[17] br[17] wl[356] vdd gnd cell_6t
Xbit_r357_c17 bl[17] br[17] wl[357] vdd gnd cell_6t
Xbit_r358_c17 bl[17] br[17] wl[358] vdd gnd cell_6t
Xbit_r359_c17 bl[17] br[17] wl[359] vdd gnd cell_6t
Xbit_r360_c17 bl[17] br[17] wl[360] vdd gnd cell_6t
Xbit_r361_c17 bl[17] br[17] wl[361] vdd gnd cell_6t
Xbit_r362_c17 bl[17] br[17] wl[362] vdd gnd cell_6t
Xbit_r363_c17 bl[17] br[17] wl[363] vdd gnd cell_6t
Xbit_r364_c17 bl[17] br[17] wl[364] vdd gnd cell_6t
Xbit_r365_c17 bl[17] br[17] wl[365] vdd gnd cell_6t
Xbit_r366_c17 bl[17] br[17] wl[366] vdd gnd cell_6t
Xbit_r367_c17 bl[17] br[17] wl[367] vdd gnd cell_6t
Xbit_r368_c17 bl[17] br[17] wl[368] vdd gnd cell_6t
Xbit_r369_c17 bl[17] br[17] wl[369] vdd gnd cell_6t
Xbit_r370_c17 bl[17] br[17] wl[370] vdd gnd cell_6t
Xbit_r371_c17 bl[17] br[17] wl[371] vdd gnd cell_6t
Xbit_r372_c17 bl[17] br[17] wl[372] vdd gnd cell_6t
Xbit_r373_c17 bl[17] br[17] wl[373] vdd gnd cell_6t
Xbit_r374_c17 bl[17] br[17] wl[374] vdd gnd cell_6t
Xbit_r375_c17 bl[17] br[17] wl[375] vdd gnd cell_6t
Xbit_r376_c17 bl[17] br[17] wl[376] vdd gnd cell_6t
Xbit_r377_c17 bl[17] br[17] wl[377] vdd gnd cell_6t
Xbit_r378_c17 bl[17] br[17] wl[378] vdd gnd cell_6t
Xbit_r379_c17 bl[17] br[17] wl[379] vdd gnd cell_6t
Xbit_r380_c17 bl[17] br[17] wl[380] vdd gnd cell_6t
Xbit_r381_c17 bl[17] br[17] wl[381] vdd gnd cell_6t
Xbit_r382_c17 bl[17] br[17] wl[382] vdd gnd cell_6t
Xbit_r383_c17 bl[17] br[17] wl[383] vdd gnd cell_6t
Xbit_r384_c17 bl[17] br[17] wl[384] vdd gnd cell_6t
Xbit_r385_c17 bl[17] br[17] wl[385] vdd gnd cell_6t
Xbit_r386_c17 bl[17] br[17] wl[386] vdd gnd cell_6t
Xbit_r387_c17 bl[17] br[17] wl[387] vdd gnd cell_6t
Xbit_r388_c17 bl[17] br[17] wl[388] vdd gnd cell_6t
Xbit_r389_c17 bl[17] br[17] wl[389] vdd gnd cell_6t
Xbit_r390_c17 bl[17] br[17] wl[390] vdd gnd cell_6t
Xbit_r391_c17 bl[17] br[17] wl[391] vdd gnd cell_6t
Xbit_r392_c17 bl[17] br[17] wl[392] vdd gnd cell_6t
Xbit_r393_c17 bl[17] br[17] wl[393] vdd gnd cell_6t
Xbit_r394_c17 bl[17] br[17] wl[394] vdd gnd cell_6t
Xbit_r395_c17 bl[17] br[17] wl[395] vdd gnd cell_6t
Xbit_r396_c17 bl[17] br[17] wl[396] vdd gnd cell_6t
Xbit_r397_c17 bl[17] br[17] wl[397] vdd gnd cell_6t
Xbit_r398_c17 bl[17] br[17] wl[398] vdd gnd cell_6t
Xbit_r399_c17 bl[17] br[17] wl[399] vdd gnd cell_6t
Xbit_r400_c17 bl[17] br[17] wl[400] vdd gnd cell_6t
Xbit_r401_c17 bl[17] br[17] wl[401] vdd gnd cell_6t
Xbit_r402_c17 bl[17] br[17] wl[402] vdd gnd cell_6t
Xbit_r403_c17 bl[17] br[17] wl[403] vdd gnd cell_6t
Xbit_r404_c17 bl[17] br[17] wl[404] vdd gnd cell_6t
Xbit_r405_c17 bl[17] br[17] wl[405] vdd gnd cell_6t
Xbit_r406_c17 bl[17] br[17] wl[406] vdd gnd cell_6t
Xbit_r407_c17 bl[17] br[17] wl[407] vdd gnd cell_6t
Xbit_r408_c17 bl[17] br[17] wl[408] vdd gnd cell_6t
Xbit_r409_c17 bl[17] br[17] wl[409] vdd gnd cell_6t
Xbit_r410_c17 bl[17] br[17] wl[410] vdd gnd cell_6t
Xbit_r411_c17 bl[17] br[17] wl[411] vdd gnd cell_6t
Xbit_r412_c17 bl[17] br[17] wl[412] vdd gnd cell_6t
Xbit_r413_c17 bl[17] br[17] wl[413] vdd gnd cell_6t
Xbit_r414_c17 bl[17] br[17] wl[414] vdd gnd cell_6t
Xbit_r415_c17 bl[17] br[17] wl[415] vdd gnd cell_6t
Xbit_r416_c17 bl[17] br[17] wl[416] vdd gnd cell_6t
Xbit_r417_c17 bl[17] br[17] wl[417] vdd gnd cell_6t
Xbit_r418_c17 bl[17] br[17] wl[418] vdd gnd cell_6t
Xbit_r419_c17 bl[17] br[17] wl[419] vdd gnd cell_6t
Xbit_r420_c17 bl[17] br[17] wl[420] vdd gnd cell_6t
Xbit_r421_c17 bl[17] br[17] wl[421] vdd gnd cell_6t
Xbit_r422_c17 bl[17] br[17] wl[422] vdd gnd cell_6t
Xbit_r423_c17 bl[17] br[17] wl[423] vdd gnd cell_6t
Xbit_r424_c17 bl[17] br[17] wl[424] vdd gnd cell_6t
Xbit_r425_c17 bl[17] br[17] wl[425] vdd gnd cell_6t
Xbit_r426_c17 bl[17] br[17] wl[426] vdd gnd cell_6t
Xbit_r427_c17 bl[17] br[17] wl[427] vdd gnd cell_6t
Xbit_r428_c17 bl[17] br[17] wl[428] vdd gnd cell_6t
Xbit_r429_c17 bl[17] br[17] wl[429] vdd gnd cell_6t
Xbit_r430_c17 bl[17] br[17] wl[430] vdd gnd cell_6t
Xbit_r431_c17 bl[17] br[17] wl[431] vdd gnd cell_6t
Xbit_r432_c17 bl[17] br[17] wl[432] vdd gnd cell_6t
Xbit_r433_c17 bl[17] br[17] wl[433] vdd gnd cell_6t
Xbit_r434_c17 bl[17] br[17] wl[434] vdd gnd cell_6t
Xbit_r435_c17 bl[17] br[17] wl[435] vdd gnd cell_6t
Xbit_r436_c17 bl[17] br[17] wl[436] vdd gnd cell_6t
Xbit_r437_c17 bl[17] br[17] wl[437] vdd gnd cell_6t
Xbit_r438_c17 bl[17] br[17] wl[438] vdd gnd cell_6t
Xbit_r439_c17 bl[17] br[17] wl[439] vdd gnd cell_6t
Xbit_r440_c17 bl[17] br[17] wl[440] vdd gnd cell_6t
Xbit_r441_c17 bl[17] br[17] wl[441] vdd gnd cell_6t
Xbit_r442_c17 bl[17] br[17] wl[442] vdd gnd cell_6t
Xbit_r443_c17 bl[17] br[17] wl[443] vdd gnd cell_6t
Xbit_r444_c17 bl[17] br[17] wl[444] vdd gnd cell_6t
Xbit_r445_c17 bl[17] br[17] wl[445] vdd gnd cell_6t
Xbit_r446_c17 bl[17] br[17] wl[446] vdd gnd cell_6t
Xbit_r447_c17 bl[17] br[17] wl[447] vdd gnd cell_6t
Xbit_r448_c17 bl[17] br[17] wl[448] vdd gnd cell_6t
Xbit_r449_c17 bl[17] br[17] wl[449] vdd gnd cell_6t
Xbit_r450_c17 bl[17] br[17] wl[450] vdd gnd cell_6t
Xbit_r451_c17 bl[17] br[17] wl[451] vdd gnd cell_6t
Xbit_r452_c17 bl[17] br[17] wl[452] vdd gnd cell_6t
Xbit_r453_c17 bl[17] br[17] wl[453] vdd gnd cell_6t
Xbit_r454_c17 bl[17] br[17] wl[454] vdd gnd cell_6t
Xbit_r455_c17 bl[17] br[17] wl[455] vdd gnd cell_6t
Xbit_r456_c17 bl[17] br[17] wl[456] vdd gnd cell_6t
Xbit_r457_c17 bl[17] br[17] wl[457] vdd gnd cell_6t
Xbit_r458_c17 bl[17] br[17] wl[458] vdd gnd cell_6t
Xbit_r459_c17 bl[17] br[17] wl[459] vdd gnd cell_6t
Xbit_r460_c17 bl[17] br[17] wl[460] vdd gnd cell_6t
Xbit_r461_c17 bl[17] br[17] wl[461] vdd gnd cell_6t
Xbit_r462_c17 bl[17] br[17] wl[462] vdd gnd cell_6t
Xbit_r463_c17 bl[17] br[17] wl[463] vdd gnd cell_6t
Xbit_r464_c17 bl[17] br[17] wl[464] vdd gnd cell_6t
Xbit_r465_c17 bl[17] br[17] wl[465] vdd gnd cell_6t
Xbit_r466_c17 bl[17] br[17] wl[466] vdd gnd cell_6t
Xbit_r467_c17 bl[17] br[17] wl[467] vdd gnd cell_6t
Xbit_r468_c17 bl[17] br[17] wl[468] vdd gnd cell_6t
Xbit_r469_c17 bl[17] br[17] wl[469] vdd gnd cell_6t
Xbit_r470_c17 bl[17] br[17] wl[470] vdd gnd cell_6t
Xbit_r471_c17 bl[17] br[17] wl[471] vdd gnd cell_6t
Xbit_r472_c17 bl[17] br[17] wl[472] vdd gnd cell_6t
Xbit_r473_c17 bl[17] br[17] wl[473] vdd gnd cell_6t
Xbit_r474_c17 bl[17] br[17] wl[474] vdd gnd cell_6t
Xbit_r475_c17 bl[17] br[17] wl[475] vdd gnd cell_6t
Xbit_r476_c17 bl[17] br[17] wl[476] vdd gnd cell_6t
Xbit_r477_c17 bl[17] br[17] wl[477] vdd gnd cell_6t
Xbit_r478_c17 bl[17] br[17] wl[478] vdd gnd cell_6t
Xbit_r479_c17 bl[17] br[17] wl[479] vdd gnd cell_6t
Xbit_r480_c17 bl[17] br[17] wl[480] vdd gnd cell_6t
Xbit_r481_c17 bl[17] br[17] wl[481] vdd gnd cell_6t
Xbit_r482_c17 bl[17] br[17] wl[482] vdd gnd cell_6t
Xbit_r483_c17 bl[17] br[17] wl[483] vdd gnd cell_6t
Xbit_r484_c17 bl[17] br[17] wl[484] vdd gnd cell_6t
Xbit_r485_c17 bl[17] br[17] wl[485] vdd gnd cell_6t
Xbit_r486_c17 bl[17] br[17] wl[486] vdd gnd cell_6t
Xbit_r487_c17 bl[17] br[17] wl[487] vdd gnd cell_6t
Xbit_r488_c17 bl[17] br[17] wl[488] vdd gnd cell_6t
Xbit_r489_c17 bl[17] br[17] wl[489] vdd gnd cell_6t
Xbit_r490_c17 bl[17] br[17] wl[490] vdd gnd cell_6t
Xbit_r491_c17 bl[17] br[17] wl[491] vdd gnd cell_6t
Xbit_r492_c17 bl[17] br[17] wl[492] vdd gnd cell_6t
Xbit_r493_c17 bl[17] br[17] wl[493] vdd gnd cell_6t
Xbit_r494_c17 bl[17] br[17] wl[494] vdd gnd cell_6t
Xbit_r495_c17 bl[17] br[17] wl[495] vdd gnd cell_6t
Xbit_r496_c17 bl[17] br[17] wl[496] vdd gnd cell_6t
Xbit_r497_c17 bl[17] br[17] wl[497] vdd gnd cell_6t
Xbit_r498_c17 bl[17] br[17] wl[498] vdd gnd cell_6t
Xbit_r499_c17 bl[17] br[17] wl[499] vdd gnd cell_6t
Xbit_r500_c17 bl[17] br[17] wl[500] vdd gnd cell_6t
Xbit_r501_c17 bl[17] br[17] wl[501] vdd gnd cell_6t
Xbit_r502_c17 bl[17] br[17] wl[502] vdd gnd cell_6t
Xbit_r503_c17 bl[17] br[17] wl[503] vdd gnd cell_6t
Xbit_r504_c17 bl[17] br[17] wl[504] vdd gnd cell_6t
Xbit_r505_c17 bl[17] br[17] wl[505] vdd gnd cell_6t
Xbit_r506_c17 bl[17] br[17] wl[506] vdd gnd cell_6t
Xbit_r507_c17 bl[17] br[17] wl[507] vdd gnd cell_6t
Xbit_r508_c17 bl[17] br[17] wl[508] vdd gnd cell_6t
Xbit_r509_c17 bl[17] br[17] wl[509] vdd gnd cell_6t
Xbit_r510_c17 bl[17] br[17] wl[510] vdd gnd cell_6t
Xbit_r511_c17 bl[17] br[17] wl[511] vdd gnd cell_6t
Xbit_r0_c18 bl[18] br[18] wl[0] vdd gnd cell_6t
Xbit_r1_c18 bl[18] br[18] wl[1] vdd gnd cell_6t
Xbit_r2_c18 bl[18] br[18] wl[2] vdd gnd cell_6t
Xbit_r3_c18 bl[18] br[18] wl[3] vdd gnd cell_6t
Xbit_r4_c18 bl[18] br[18] wl[4] vdd gnd cell_6t
Xbit_r5_c18 bl[18] br[18] wl[5] vdd gnd cell_6t
Xbit_r6_c18 bl[18] br[18] wl[6] vdd gnd cell_6t
Xbit_r7_c18 bl[18] br[18] wl[7] vdd gnd cell_6t
Xbit_r8_c18 bl[18] br[18] wl[8] vdd gnd cell_6t
Xbit_r9_c18 bl[18] br[18] wl[9] vdd gnd cell_6t
Xbit_r10_c18 bl[18] br[18] wl[10] vdd gnd cell_6t
Xbit_r11_c18 bl[18] br[18] wl[11] vdd gnd cell_6t
Xbit_r12_c18 bl[18] br[18] wl[12] vdd gnd cell_6t
Xbit_r13_c18 bl[18] br[18] wl[13] vdd gnd cell_6t
Xbit_r14_c18 bl[18] br[18] wl[14] vdd gnd cell_6t
Xbit_r15_c18 bl[18] br[18] wl[15] vdd gnd cell_6t
Xbit_r16_c18 bl[18] br[18] wl[16] vdd gnd cell_6t
Xbit_r17_c18 bl[18] br[18] wl[17] vdd gnd cell_6t
Xbit_r18_c18 bl[18] br[18] wl[18] vdd gnd cell_6t
Xbit_r19_c18 bl[18] br[18] wl[19] vdd gnd cell_6t
Xbit_r20_c18 bl[18] br[18] wl[20] vdd gnd cell_6t
Xbit_r21_c18 bl[18] br[18] wl[21] vdd gnd cell_6t
Xbit_r22_c18 bl[18] br[18] wl[22] vdd gnd cell_6t
Xbit_r23_c18 bl[18] br[18] wl[23] vdd gnd cell_6t
Xbit_r24_c18 bl[18] br[18] wl[24] vdd gnd cell_6t
Xbit_r25_c18 bl[18] br[18] wl[25] vdd gnd cell_6t
Xbit_r26_c18 bl[18] br[18] wl[26] vdd gnd cell_6t
Xbit_r27_c18 bl[18] br[18] wl[27] vdd gnd cell_6t
Xbit_r28_c18 bl[18] br[18] wl[28] vdd gnd cell_6t
Xbit_r29_c18 bl[18] br[18] wl[29] vdd gnd cell_6t
Xbit_r30_c18 bl[18] br[18] wl[30] vdd gnd cell_6t
Xbit_r31_c18 bl[18] br[18] wl[31] vdd gnd cell_6t
Xbit_r32_c18 bl[18] br[18] wl[32] vdd gnd cell_6t
Xbit_r33_c18 bl[18] br[18] wl[33] vdd gnd cell_6t
Xbit_r34_c18 bl[18] br[18] wl[34] vdd gnd cell_6t
Xbit_r35_c18 bl[18] br[18] wl[35] vdd gnd cell_6t
Xbit_r36_c18 bl[18] br[18] wl[36] vdd gnd cell_6t
Xbit_r37_c18 bl[18] br[18] wl[37] vdd gnd cell_6t
Xbit_r38_c18 bl[18] br[18] wl[38] vdd gnd cell_6t
Xbit_r39_c18 bl[18] br[18] wl[39] vdd gnd cell_6t
Xbit_r40_c18 bl[18] br[18] wl[40] vdd gnd cell_6t
Xbit_r41_c18 bl[18] br[18] wl[41] vdd gnd cell_6t
Xbit_r42_c18 bl[18] br[18] wl[42] vdd gnd cell_6t
Xbit_r43_c18 bl[18] br[18] wl[43] vdd gnd cell_6t
Xbit_r44_c18 bl[18] br[18] wl[44] vdd gnd cell_6t
Xbit_r45_c18 bl[18] br[18] wl[45] vdd gnd cell_6t
Xbit_r46_c18 bl[18] br[18] wl[46] vdd gnd cell_6t
Xbit_r47_c18 bl[18] br[18] wl[47] vdd gnd cell_6t
Xbit_r48_c18 bl[18] br[18] wl[48] vdd gnd cell_6t
Xbit_r49_c18 bl[18] br[18] wl[49] vdd gnd cell_6t
Xbit_r50_c18 bl[18] br[18] wl[50] vdd gnd cell_6t
Xbit_r51_c18 bl[18] br[18] wl[51] vdd gnd cell_6t
Xbit_r52_c18 bl[18] br[18] wl[52] vdd gnd cell_6t
Xbit_r53_c18 bl[18] br[18] wl[53] vdd gnd cell_6t
Xbit_r54_c18 bl[18] br[18] wl[54] vdd gnd cell_6t
Xbit_r55_c18 bl[18] br[18] wl[55] vdd gnd cell_6t
Xbit_r56_c18 bl[18] br[18] wl[56] vdd gnd cell_6t
Xbit_r57_c18 bl[18] br[18] wl[57] vdd gnd cell_6t
Xbit_r58_c18 bl[18] br[18] wl[58] vdd gnd cell_6t
Xbit_r59_c18 bl[18] br[18] wl[59] vdd gnd cell_6t
Xbit_r60_c18 bl[18] br[18] wl[60] vdd gnd cell_6t
Xbit_r61_c18 bl[18] br[18] wl[61] vdd gnd cell_6t
Xbit_r62_c18 bl[18] br[18] wl[62] vdd gnd cell_6t
Xbit_r63_c18 bl[18] br[18] wl[63] vdd gnd cell_6t
Xbit_r64_c18 bl[18] br[18] wl[64] vdd gnd cell_6t
Xbit_r65_c18 bl[18] br[18] wl[65] vdd gnd cell_6t
Xbit_r66_c18 bl[18] br[18] wl[66] vdd gnd cell_6t
Xbit_r67_c18 bl[18] br[18] wl[67] vdd gnd cell_6t
Xbit_r68_c18 bl[18] br[18] wl[68] vdd gnd cell_6t
Xbit_r69_c18 bl[18] br[18] wl[69] vdd gnd cell_6t
Xbit_r70_c18 bl[18] br[18] wl[70] vdd gnd cell_6t
Xbit_r71_c18 bl[18] br[18] wl[71] vdd gnd cell_6t
Xbit_r72_c18 bl[18] br[18] wl[72] vdd gnd cell_6t
Xbit_r73_c18 bl[18] br[18] wl[73] vdd gnd cell_6t
Xbit_r74_c18 bl[18] br[18] wl[74] vdd gnd cell_6t
Xbit_r75_c18 bl[18] br[18] wl[75] vdd gnd cell_6t
Xbit_r76_c18 bl[18] br[18] wl[76] vdd gnd cell_6t
Xbit_r77_c18 bl[18] br[18] wl[77] vdd gnd cell_6t
Xbit_r78_c18 bl[18] br[18] wl[78] vdd gnd cell_6t
Xbit_r79_c18 bl[18] br[18] wl[79] vdd gnd cell_6t
Xbit_r80_c18 bl[18] br[18] wl[80] vdd gnd cell_6t
Xbit_r81_c18 bl[18] br[18] wl[81] vdd gnd cell_6t
Xbit_r82_c18 bl[18] br[18] wl[82] vdd gnd cell_6t
Xbit_r83_c18 bl[18] br[18] wl[83] vdd gnd cell_6t
Xbit_r84_c18 bl[18] br[18] wl[84] vdd gnd cell_6t
Xbit_r85_c18 bl[18] br[18] wl[85] vdd gnd cell_6t
Xbit_r86_c18 bl[18] br[18] wl[86] vdd gnd cell_6t
Xbit_r87_c18 bl[18] br[18] wl[87] vdd gnd cell_6t
Xbit_r88_c18 bl[18] br[18] wl[88] vdd gnd cell_6t
Xbit_r89_c18 bl[18] br[18] wl[89] vdd gnd cell_6t
Xbit_r90_c18 bl[18] br[18] wl[90] vdd gnd cell_6t
Xbit_r91_c18 bl[18] br[18] wl[91] vdd gnd cell_6t
Xbit_r92_c18 bl[18] br[18] wl[92] vdd gnd cell_6t
Xbit_r93_c18 bl[18] br[18] wl[93] vdd gnd cell_6t
Xbit_r94_c18 bl[18] br[18] wl[94] vdd gnd cell_6t
Xbit_r95_c18 bl[18] br[18] wl[95] vdd gnd cell_6t
Xbit_r96_c18 bl[18] br[18] wl[96] vdd gnd cell_6t
Xbit_r97_c18 bl[18] br[18] wl[97] vdd gnd cell_6t
Xbit_r98_c18 bl[18] br[18] wl[98] vdd gnd cell_6t
Xbit_r99_c18 bl[18] br[18] wl[99] vdd gnd cell_6t
Xbit_r100_c18 bl[18] br[18] wl[100] vdd gnd cell_6t
Xbit_r101_c18 bl[18] br[18] wl[101] vdd gnd cell_6t
Xbit_r102_c18 bl[18] br[18] wl[102] vdd gnd cell_6t
Xbit_r103_c18 bl[18] br[18] wl[103] vdd gnd cell_6t
Xbit_r104_c18 bl[18] br[18] wl[104] vdd gnd cell_6t
Xbit_r105_c18 bl[18] br[18] wl[105] vdd gnd cell_6t
Xbit_r106_c18 bl[18] br[18] wl[106] vdd gnd cell_6t
Xbit_r107_c18 bl[18] br[18] wl[107] vdd gnd cell_6t
Xbit_r108_c18 bl[18] br[18] wl[108] vdd gnd cell_6t
Xbit_r109_c18 bl[18] br[18] wl[109] vdd gnd cell_6t
Xbit_r110_c18 bl[18] br[18] wl[110] vdd gnd cell_6t
Xbit_r111_c18 bl[18] br[18] wl[111] vdd gnd cell_6t
Xbit_r112_c18 bl[18] br[18] wl[112] vdd gnd cell_6t
Xbit_r113_c18 bl[18] br[18] wl[113] vdd gnd cell_6t
Xbit_r114_c18 bl[18] br[18] wl[114] vdd gnd cell_6t
Xbit_r115_c18 bl[18] br[18] wl[115] vdd gnd cell_6t
Xbit_r116_c18 bl[18] br[18] wl[116] vdd gnd cell_6t
Xbit_r117_c18 bl[18] br[18] wl[117] vdd gnd cell_6t
Xbit_r118_c18 bl[18] br[18] wl[118] vdd gnd cell_6t
Xbit_r119_c18 bl[18] br[18] wl[119] vdd gnd cell_6t
Xbit_r120_c18 bl[18] br[18] wl[120] vdd gnd cell_6t
Xbit_r121_c18 bl[18] br[18] wl[121] vdd gnd cell_6t
Xbit_r122_c18 bl[18] br[18] wl[122] vdd gnd cell_6t
Xbit_r123_c18 bl[18] br[18] wl[123] vdd gnd cell_6t
Xbit_r124_c18 bl[18] br[18] wl[124] vdd gnd cell_6t
Xbit_r125_c18 bl[18] br[18] wl[125] vdd gnd cell_6t
Xbit_r126_c18 bl[18] br[18] wl[126] vdd gnd cell_6t
Xbit_r127_c18 bl[18] br[18] wl[127] vdd gnd cell_6t
Xbit_r128_c18 bl[18] br[18] wl[128] vdd gnd cell_6t
Xbit_r129_c18 bl[18] br[18] wl[129] vdd gnd cell_6t
Xbit_r130_c18 bl[18] br[18] wl[130] vdd gnd cell_6t
Xbit_r131_c18 bl[18] br[18] wl[131] vdd gnd cell_6t
Xbit_r132_c18 bl[18] br[18] wl[132] vdd gnd cell_6t
Xbit_r133_c18 bl[18] br[18] wl[133] vdd gnd cell_6t
Xbit_r134_c18 bl[18] br[18] wl[134] vdd gnd cell_6t
Xbit_r135_c18 bl[18] br[18] wl[135] vdd gnd cell_6t
Xbit_r136_c18 bl[18] br[18] wl[136] vdd gnd cell_6t
Xbit_r137_c18 bl[18] br[18] wl[137] vdd gnd cell_6t
Xbit_r138_c18 bl[18] br[18] wl[138] vdd gnd cell_6t
Xbit_r139_c18 bl[18] br[18] wl[139] vdd gnd cell_6t
Xbit_r140_c18 bl[18] br[18] wl[140] vdd gnd cell_6t
Xbit_r141_c18 bl[18] br[18] wl[141] vdd gnd cell_6t
Xbit_r142_c18 bl[18] br[18] wl[142] vdd gnd cell_6t
Xbit_r143_c18 bl[18] br[18] wl[143] vdd gnd cell_6t
Xbit_r144_c18 bl[18] br[18] wl[144] vdd gnd cell_6t
Xbit_r145_c18 bl[18] br[18] wl[145] vdd gnd cell_6t
Xbit_r146_c18 bl[18] br[18] wl[146] vdd gnd cell_6t
Xbit_r147_c18 bl[18] br[18] wl[147] vdd gnd cell_6t
Xbit_r148_c18 bl[18] br[18] wl[148] vdd gnd cell_6t
Xbit_r149_c18 bl[18] br[18] wl[149] vdd gnd cell_6t
Xbit_r150_c18 bl[18] br[18] wl[150] vdd gnd cell_6t
Xbit_r151_c18 bl[18] br[18] wl[151] vdd gnd cell_6t
Xbit_r152_c18 bl[18] br[18] wl[152] vdd gnd cell_6t
Xbit_r153_c18 bl[18] br[18] wl[153] vdd gnd cell_6t
Xbit_r154_c18 bl[18] br[18] wl[154] vdd gnd cell_6t
Xbit_r155_c18 bl[18] br[18] wl[155] vdd gnd cell_6t
Xbit_r156_c18 bl[18] br[18] wl[156] vdd gnd cell_6t
Xbit_r157_c18 bl[18] br[18] wl[157] vdd gnd cell_6t
Xbit_r158_c18 bl[18] br[18] wl[158] vdd gnd cell_6t
Xbit_r159_c18 bl[18] br[18] wl[159] vdd gnd cell_6t
Xbit_r160_c18 bl[18] br[18] wl[160] vdd gnd cell_6t
Xbit_r161_c18 bl[18] br[18] wl[161] vdd gnd cell_6t
Xbit_r162_c18 bl[18] br[18] wl[162] vdd gnd cell_6t
Xbit_r163_c18 bl[18] br[18] wl[163] vdd gnd cell_6t
Xbit_r164_c18 bl[18] br[18] wl[164] vdd gnd cell_6t
Xbit_r165_c18 bl[18] br[18] wl[165] vdd gnd cell_6t
Xbit_r166_c18 bl[18] br[18] wl[166] vdd gnd cell_6t
Xbit_r167_c18 bl[18] br[18] wl[167] vdd gnd cell_6t
Xbit_r168_c18 bl[18] br[18] wl[168] vdd gnd cell_6t
Xbit_r169_c18 bl[18] br[18] wl[169] vdd gnd cell_6t
Xbit_r170_c18 bl[18] br[18] wl[170] vdd gnd cell_6t
Xbit_r171_c18 bl[18] br[18] wl[171] vdd gnd cell_6t
Xbit_r172_c18 bl[18] br[18] wl[172] vdd gnd cell_6t
Xbit_r173_c18 bl[18] br[18] wl[173] vdd gnd cell_6t
Xbit_r174_c18 bl[18] br[18] wl[174] vdd gnd cell_6t
Xbit_r175_c18 bl[18] br[18] wl[175] vdd gnd cell_6t
Xbit_r176_c18 bl[18] br[18] wl[176] vdd gnd cell_6t
Xbit_r177_c18 bl[18] br[18] wl[177] vdd gnd cell_6t
Xbit_r178_c18 bl[18] br[18] wl[178] vdd gnd cell_6t
Xbit_r179_c18 bl[18] br[18] wl[179] vdd gnd cell_6t
Xbit_r180_c18 bl[18] br[18] wl[180] vdd gnd cell_6t
Xbit_r181_c18 bl[18] br[18] wl[181] vdd gnd cell_6t
Xbit_r182_c18 bl[18] br[18] wl[182] vdd gnd cell_6t
Xbit_r183_c18 bl[18] br[18] wl[183] vdd gnd cell_6t
Xbit_r184_c18 bl[18] br[18] wl[184] vdd gnd cell_6t
Xbit_r185_c18 bl[18] br[18] wl[185] vdd gnd cell_6t
Xbit_r186_c18 bl[18] br[18] wl[186] vdd gnd cell_6t
Xbit_r187_c18 bl[18] br[18] wl[187] vdd gnd cell_6t
Xbit_r188_c18 bl[18] br[18] wl[188] vdd gnd cell_6t
Xbit_r189_c18 bl[18] br[18] wl[189] vdd gnd cell_6t
Xbit_r190_c18 bl[18] br[18] wl[190] vdd gnd cell_6t
Xbit_r191_c18 bl[18] br[18] wl[191] vdd gnd cell_6t
Xbit_r192_c18 bl[18] br[18] wl[192] vdd gnd cell_6t
Xbit_r193_c18 bl[18] br[18] wl[193] vdd gnd cell_6t
Xbit_r194_c18 bl[18] br[18] wl[194] vdd gnd cell_6t
Xbit_r195_c18 bl[18] br[18] wl[195] vdd gnd cell_6t
Xbit_r196_c18 bl[18] br[18] wl[196] vdd gnd cell_6t
Xbit_r197_c18 bl[18] br[18] wl[197] vdd gnd cell_6t
Xbit_r198_c18 bl[18] br[18] wl[198] vdd gnd cell_6t
Xbit_r199_c18 bl[18] br[18] wl[199] vdd gnd cell_6t
Xbit_r200_c18 bl[18] br[18] wl[200] vdd gnd cell_6t
Xbit_r201_c18 bl[18] br[18] wl[201] vdd gnd cell_6t
Xbit_r202_c18 bl[18] br[18] wl[202] vdd gnd cell_6t
Xbit_r203_c18 bl[18] br[18] wl[203] vdd gnd cell_6t
Xbit_r204_c18 bl[18] br[18] wl[204] vdd gnd cell_6t
Xbit_r205_c18 bl[18] br[18] wl[205] vdd gnd cell_6t
Xbit_r206_c18 bl[18] br[18] wl[206] vdd gnd cell_6t
Xbit_r207_c18 bl[18] br[18] wl[207] vdd gnd cell_6t
Xbit_r208_c18 bl[18] br[18] wl[208] vdd gnd cell_6t
Xbit_r209_c18 bl[18] br[18] wl[209] vdd gnd cell_6t
Xbit_r210_c18 bl[18] br[18] wl[210] vdd gnd cell_6t
Xbit_r211_c18 bl[18] br[18] wl[211] vdd gnd cell_6t
Xbit_r212_c18 bl[18] br[18] wl[212] vdd gnd cell_6t
Xbit_r213_c18 bl[18] br[18] wl[213] vdd gnd cell_6t
Xbit_r214_c18 bl[18] br[18] wl[214] vdd gnd cell_6t
Xbit_r215_c18 bl[18] br[18] wl[215] vdd gnd cell_6t
Xbit_r216_c18 bl[18] br[18] wl[216] vdd gnd cell_6t
Xbit_r217_c18 bl[18] br[18] wl[217] vdd gnd cell_6t
Xbit_r218_c18 bl[18] br[18] wl[218] vdd gnd cell_6t
Xbit_r219_c18 bl[18] br[18] wl[219] vdd gnd cell_6t
Xbit_r220_c18 bl[18] br[18] wl[220] vdd gnd cell_6t
Xbit_r221_c18 bl[18] br[18] wl[221] vdd gnd cell_6t
Xbit_r222_c18 bl[18] br[18] wl[222] vdd gnd cell_6t
Xbit_r223_c18 bl[18] br[18] wl[223] vdd gnd cell_6t
Xbit_r224_c18 bl[18] br[18] wl[224] vdd gnd cell_6t
Xbit_r225_c18 bl[18] br[18] wl[225] vdd gnd cell_6t
Xbit_r226_c18 bl[18] br[18] wl[226] vdd gnd cell_6t
Xbit_r227_c18 bl[18] br[18] wl[227] vdd gnd cell_6t
Xbit_r228_c18 bl[18] br[18] wl[228] vdd gnd cell_6t
Xbit_r229_c18 bl[18] br[18] wl[229] vdd gnd cell_6t
Xbit_r230_c18 bl[18] br[18] wl[230] vdd gnd cell_6t
Xbit_r231_c18 bl[18] br[18] wl[231] vdd gnd cell_6t
Xbit_r232_c18 bl[18] br[18] wl[232] vdd gnd cell_6t
Xbit_r233_c18 bl[18] br[18] wl[233] vdd gnd cell_6t
Xbit_r234_c18 bl[18] br[18] wl[234] vdd gnd cell_6t
Xbit_r235_c18 bl[18] br[18] wl[235] vdd gnd cell_6t
Xbit_r236_c18 bl[18] br[18] wl[236] vdd gnd cell_6t
Xbit_r237_c18 bl[18] br[18] wl[237] vdd gnd cell_6t
Xbit_r238_c18 bl[18] br[18] wl[238] vdd gnd cell_6t
Xbit_r239_c18 bl[18] br[18] wl[239] vdd gnd cell_6t
Xbit_r240_c18 bl[18] br[18] wl[240] vdd gnd cell_6t
Xbit_r241_c18 bl[18] br[18] wl[241] vdd gnd cell_6t
Xbit_r242_c18 bl[18] br[18] wl[242] vdd gnd cell_6t
Xbit_r243_c18 bl[18] br[18] wl[243] vdd gnd cell_6t
Xbit_r244_c18 bl[18] br[18] wl[244] vdd gnd cell_6t
Xbit_r245_c18 bl[18] br[18] wl[245] vdd gnd cell_6t
Xbit_r246_c18 bl[18] br[18] wl[246] vdd gnd cell_6t
Xbit_r247_c18 bl[18] br[18] wl[247] vdd gnd cell_6t
Xbit_r248_c18 bl[18] br[18] wl[248] vdd gnd cell_6t
Xbit_r249_c18 bl[18] br[18] wl[249] vdd gnd cell_6t
Xbit_r250_c18 bl[18] br[18] wl[250] vdd gnd cell_6t
Xbit_r251_c18 bl[18] br[18] wl[251] vdd gnd cell_6t
Xbit_r252_c18 bl[18] br[18] wl[252] vdd gnd cell_6t
Xbit_r253_c18 bl[18] br[18] wl[253] vdd gnd cell_6t
Xbit_r254_c18 bl[18] br[18] wl[254] vdd gnd cell_6t
Xbit_r255_c18 bl[18] br[18] wl[255] vdd gnd cell_6t
Xbit_r256_c18 bl[18] br[18] wl[256] vdd gnd cell_6t
Xbit_r257_c18 bl[18] br[18] wl[257] vdd gnd cell_6t
Xbit_r258_c18 bl[18] br[18] wl[258] vdd gnd cell_6t
Xbit_r259_c18 bl[18] br[18] wl[259] vdd gnd cell_6t
Xbit_r260_c18 bl[18] br[18] wl[260] vdd gnd cell_6t
Xbit_r261_c18 bl[18] br[18] wl[261] vdd gnd cell_6t
Xbit_r262_c18 bl[18] br[18] wl[262] vdd gnd cell_6t
Xbit_r263_c18 bl[18] br[18] wl[263] vdd gnd cell_6t
Xbit_r264_c18 bl[18] br[18] wl[264] vdd gnd cell_6t
Xbit_r265_c18 bl[18] br[18] wl[265] vdd gnd cell_6t
Xbit_r266_c18 bl[18] br[18] wl[266] vdd gnd cell_6t
Xbit_r267_c18 bl[18] br[18] wl[267] vdd gnd cell_6t
Xbit_r268_c18 bl[18] br[18] wl[268] vdd gnd cell_6t
Xbit_r269_c18 bl[18] br[18] wl[269] vdd gnd cell_6t
Xbit_r270_c18 bl[18] br[18] wl[270] vdd gnd cell_6t
Xbit_r271_c18 bl[18] br[18] wl[271] vdd gnd cell_6t
Xbit_r272_c18 bl[18] br[18] wl[272] vdd gnd cell_6t
Xbit_r273_c18 bl[18] br[18] wl[273] vdd gnd cell_6t
Xbit_r274_c18 bl[18] br[18] wl[274] vdd gnd cell_6t
Xbit_r275_c18 bl[18] br[18] wl[275] vdd gnd cell_6t
Xbit_r276_c18 bl[18] br[18] wl[276] vdd gnd cell_6t
Xbit_r277_c18 bl[18] br[18] wl[277] vdd gnd cell_6t
Xbit_r278_c18 bl[18] br[18] wl[278] vdd gnd cell_6t
Xbit_r279_c18 bl[18] br[18] wl[279] vdd gnd cell_6t
Xbit_r280_c18 bl[18] br[18] wl[280] vdd gnd cell_6t
Xbit_r281_c18 bl[18] br[18] wl[281] vdd gnd cell_6t
Xbit_r282_c18 bl[18] br[18] wl[282] vdd gnd cell_6t
Xbit_r283_c18 bl[18] br[18] wl[283] vdd gnd cell_6t
Xbit_r284_c18 bl[18] br[18] wl[284] vdd gnd cell_6t
Xbit_r285_c18 bl[18] br[18] wl[285] vdd gnd cell_6t
Xbit_r286_c18 bl[18] br[18] wl[286] vdd gnd cell_6t
Xbit_r287_c18 bl[18] br[18] wl[287] vdd gnd cell_6t
Xbit_r288_c18 bl[18] br[18] wl[288] vdd gnd cell_6t
Xbit_r289_c18 bl[18] br[18] wl[289] vdd gnd cell_6t
Xbit_r290_c18 bl[18] br[18] wl[290] vdd gnd cell_6t
Xbit_r291_c18 bl[18] br[18] wl[291] vdd gnd cell_6t
Xbit_r292_c18 bl[18] br[18] wl[292] vdd gnd cell_6t
Xbit_r293_c18 bl[18] br[18] wl[293] vdd gnd cell_6t
Xbit_r294_c18 bl[18] br[18] wl[294] vdd gnd cell_6t
Xbit_r295_c18 bl[18] br[18] wl[295] vdd gnd cell_6t
Xbit_r296_c18 bl[18] br[18] wl[296] vdd gnd cell_6t
Xbit_r297_c18 bl[18] br[18] wl[297] vdd gnd cell_6t
Xbit_r298_c18 bl[18] br[18] wl[298] vdd gnd cell_6t
Xbit_r299_c18 bl[18] br[18] wl[299] vdd gnd cell_6t
Xbit_r300_c18 bl[18] br[18] wl[300] vdd gnd cell_6t
Xbit_r301_c18 bl[18] br[18] wl[301] vdd gnd cell_6t
Xbit_r302_c18 bl[18] br[18] wl[302] vdd gnd cell_6t
Xbit_r303_c18 bl[18] br[18] wl[303] vdd gnd cell_6t
Xbit_r304_c18 bl[18] br[18] wl[304] vdd gnd cell_6t
Xbit_r305_c18 bl[18] br[18] wl[305] vdd gnd cell_6t
Xbit_r306_c18 bl[18] br[18] wl[306] vdd gnd cell_6t
Xbit_r307_c18 bl[18] br[18] wl[307] vdd gnd cell_6t
Xbit_r308_c18 bl[18] br[18] wl[308] vdd gnd cell_6t
Xbit_r309_c18 bl[18] br[18] wl[309] vdd gnd cell_6t
Xbit_r310_c18 bl[18] br[18] wl[310] vdd gnd cell_6t
Xbit_r311_c18 bl[18] br[18] wl[311] vdd gnd cell_6t
Xbit_r312_c18 bl[18] br[18] wl[312] vdd gnd cell_6t
Xbit_r313_c18 bl[18] br[18] wl[313] vdd gnd cell_6t
Xbit_r314_c18 bl[18] br[18] wl[314] vdd gnd cell_6t
Xbit_r315_c18 bl[18] br[18] wl[315] vdd gnd cell_6t
Xbit_r316_c18 bl[18] br[18] wl[316] vdd gnd cell_6t
Xbit_r317_c18 bl[18] br[18] wl[317] vdd gnd cell_6t
Xbit_r318_c18 bl[18] br[18] wl[318] vdd gnd cell_6t
Xbit_r319_c18 bl[18] br[18] wl[319] vdd gnd cell_6t
Xbit_r320_c18 bl[18] br[18] wl[320] vdd gnd cell_6t
Xbit_r321_c18 bl[18] br[18] wl[321] vdd gnd cell_6t
Xbit_r322_c18 bl[18] br[18] wl[322] vdd gnd cell_6t
Xbit_r323_c18 bl[18] br[18] wl[323] vdd gnd cell_6t
Xbit_r324_c18 bl[18] br[18] wl[324] vdd gnd cell_6t
Xbit_r325_c18 bl[18] br[18] wl[325] vdd gnd cell_6t
Xbit_r326_c18 bl[18] br[18] wl[326] vdd gnd cell_6t
Xbit_r327_c18 bl[18] br[18] wl[327] vdd gnd cell_6t
Xbit_r328_c18 bl[18] br[18] wl[328] vdd gnd cell_6t
Xbit_r329_c18 bl[18] br[18] wl[329] vdd gnd cell_6t
Xbit_r330_c18 bl[18] br[18] wl[330] vdd gnd cell_6t
Xbit_r331_c18 bl[18] br[18] wl[331] vdd gnd cell_6t
Xbit_r332_c18 bl[18] br[18] wl[332] vdd gnd cell_6t
Xbit_r333_c18 bl[18] br[18] wl[333] vdd gnd cell_6t
Xbit_r334_c18 bl[18] br[18] wl[334] vdd gnd cell_6t
Xbit_r335_c18 bl[18] br[18] wl[335] vdd gnd cell_6t
Xbit_r336_c18 bl[18] br[18] wl[336] vdd gnd cell_6t
Xbit_r337_c18 bl[18] br[18] wl[337] vdd gnd cell_6t
Xbit_r338_c18 bl[18] br[18] wl[338] vdd gnd cell_6t
Xbit_r339_c18 bl[18] br[18] wl[339] vdd gnd cell_6t
Xbit_r340_c18 bl[18] br[18] wl[340] vdd gnd cell_6t
Xbit_r341_c18 bl[18] br[18] wl[341] vdd gnd cell_6t
Xbit_r342_c18 bl[18] br[18] wl[342] vdd gnd cell_6t
Xbit_r343_c18 bl[18] br[18] wl[343] vdd gnd cell_6t
Xbit_r344_c18 bl[18] br[18] wl[344] vdd gnd cell_6t
Xbit_r345_c18 bl[18] br[18] wl[345] vdd gnd cell_6t
Xbit_r346_c18 bl[18] br[18] wl[346] vdd gnd cell_6t
Xbit_r347_c18 bl[18] br[18] wl[347] vdd gnd cell_6t
Xbit_r348_c18 bl[18] br[18] wl[348] vdd gnd cell_6t
Xbit_r349_c18 bl[18] br[18] wl[349] vdd gnd cell_6t
Xbit_r350_c18 bl[18] br[18] wl[350] vdd gnd cell_6t
Xbit_r351_c18 bl[18] br[18] wl[351] vdd gnd cell_6t
Xbit_r352_c18 bl[18] br[18] wl[352] vdd gnd cell_6t
Xbit_r353_c18 bl[18] br[18] wl[353] vdd gnd cell_6t
Xbit_r354_c18 bl[18] br[18] wl[354] vdd gnd cell_6t
Xbit_r355_c18 bl[18] br[18] wl[355] vdd gnd cell_6t
Xbit_r356_c18 bl[18] br[18] wl[356] vdd gnd cell_6t
Xbit_r357_c18 bl[18] br[18] wl[357] vdd gnd cell_6t
Xbit_r358_c18 bl[18] br[18] wl[358] vdd gnd cell_6t
Xbit_r359_c18 bl[18] br[18] wl[359] vdd gnd cell_6t
Xbit_r360_c18 bl[18] br[18] wl[360] vdd gnd cell_6t
Xbit_r361_c18 bl[18] br[18] wl[361] vdd gnd cell_6t
Xbit_r362_c18 bl[18] br[18] wl[362] vdd gnd cell_6t
Xbit_r363_c18 bl[18] br[18] wl[363] vdd gnd cell_6t
Xbit_r364_c18 bl[18] br[18] wl[364] vdd gnd cell_6t
Xbit_r365_c18 bl[18] br[18] wl[365] vdd gnd cell_6t
Xbit_r366_c18 bl[18] br[18] wl[366] vdd gnd cell_6t
Xbit_r367_c18 bl[18] br[18] wl[367] vdd gnd cell_6t
Xbit_r368_c18 bl[18] br[18] wl[368] vdd gnd cell_6t
Xbit_r369_c18 bl[18] br[18] wl[369] vdd gnd cell_6t
Xbit_r370_c18 bl[18] br[18] wl[370] vdd gnd cell_6t
Xbit_r371_c18 bl[18] br[18] wl[371] vdd gnd cell_6t
Xbit_r372_c18 bl[18] br[18] wl[372] vdd gnd cell_6t
Xbit_r373_c18 bl[18] br[18] wl[373] vdd gnd cell_6t
Xbit_r374_c18 bl[18] br[18] wl[374] vdd gnd cell_6t
Xbit_r375_c18 bl[18] br[18] wl[375] vdd gnd cell_6t
Xbit_r376_c18 bl[18] br[18] wl[376] vdd gnd cell_6t
Xbit_r377_c18 bl[18] br[18] wl[377] vdd gnd cell_6t
Xbit_r378_c18 bl[18] br[18] wl[378] vdd gnd cell_6t
Xbit_r379_c18 bl[18] br[18] wl[379] vdd gnd cell_6t
Xbit_r380_c18 bl[18] br[18] wl[380] vdd gnd cell_6t
Xbit_r381_c18 bl[18] br[18] wl[381] vdd gnd cell_6t
Xbit_r382_c18 bl[18] br[18] wl[382] vdd gnd cell_6t
Xbit_r383_c18 bl[18] br[18] wl[383] vdd gnd cell_6t
Xbit_r384_c18 bl[18] br[18] wl[384] vdd gnd cell_6t
Xbit_r385_c18 bl[18] br[18] wl[385] vdd gnd cell_6t
Xbit_r386_c18 bl[18] br[18] wl[386] vdd gnd cell_6t
Xbit_r387_c18 bl[18] br[18] wl[387] vdd gnd cell_6t
Xbit_r388_c18 bl[18] br[18] wl[388] vdd gnd cell_6t
Xbit_r389_c18 bl[18] br[18] wl[389] vdd gnd cell_6t
Xbit_r390_c18 bl[18] br[18] wl[390] vdd gnd cell_6t
Xbit_r391_c18 bl[18] br[18] wl[391] vdd gnd cell_6t
Xbit_r392_c18 bl[18] br[18] wl[392] vdd gnd cell_6t
Xbit_r393_c18 bl[18] br[18] wl[393] vdd gnd cell_6t
Xbit_r394_c18 bl[18] br[18] wl[394] vdd gnd cell_6t
Xbit_r395_c18 bl[18] br[18] wl[395] vdd gnd cell_6t
Xbit_r396_c18 bl[18] br[18] wl[396] vdd gnd cell_6t
Xbit_r397_c18 bl[18] br[18] wl[397] vdd gnd cell_6t
Xbit_r398_c18 bl[18] br[18] wl[398] vdd gnd cell_6t
Xbit_r399_c18 bl[18] br[18] wl[399] vdd gnd cell_6t
Xbit_r400_c18 bl[18] br[18] wl[400] vdd gnd cell_6t
Xbit_r401_c18 bl[18] br[18] wl[401] vdd gnd cell_6t
Xbit_r402_c18 bl[18] br[18] wl[402] vdd gnd cell_6t
Xbit_r403_c18 bl[18] br[18] wl[403] vdd gnd cell_6t
Xbit_r404_c18 bl[18] br[18] wl[404] vdd gnd cell_6t
Xbit_r405_c18 bl[18] br[18] wl[405] vdd gnd cell_6t
Xbit_r406_c18 bl[18] br[18] wl[406] vdd gnd cell_6t
Xbit_r407_c18 bl[18] br[18] wl[407] vdd gnd cell_6t
Xbit_r408_c18 bl[18] br[18] wl[408] vdd gnd cell_6t
Xbit_r409_c18 bl[18] br[18] wl[409] vdd gnd cell_6t
Xbit_r410_c18 bl[18] br[18] wl[410] vdd gnd cell_6t
Xbit_r411_c18 bl[18] br[18] wl[411] vdd gnd cell_6t
Xbit_r412_c18 bl[18] br[18] wl[412] vdd gnd cell_6t
Xbit_r413_c18 bl[18] br[18] wl[413] vdd gnd cell_6t
Xbit_r414_c18 bl[18] br[18] wl[414] vdd gnd cell_6t
Xbit_r415_c18 bl[18] br[18] wl[415] vdd gnd cell_6t
Xbit_r416_c18 bl[18] br[18] wl[416] vdd gnd cell_6t
Xbit_r417_c18 bl[18] br[18] wl[417] vdd gnd cell_6t
Xbit_r418_c18 bl[18] br[18] wl[418] vdd gnd cell_6t
Xbit_r419_c18 bl[18] br[18] wl[419] vdd gnd cell_6t
Xbit_r420_c18 bl[18] br[18] wl[420] vdd gnd cell_6t
Xbit_r421_c18 bl[18] br[18] wl[421] vdd gnd cell_6t
Xbit_r422_c18 bl[18] br[18] wl[422] vdd gnd cell_6t
Xbit_r423_c18 bl[18] br[18] wl[423] vdd gnd cell_6t
Xbit_r424_c18 bl[18] br[18] wl[424] vdd gnd cell_6t
Xbit_r425_c18 bl[18] br[18] wl[425] vdd gnd cell_6t
Xbit_r426_c18 bl[18] br[18] wl[426] vdd gnd cell_6t
Xbit_r427_c18 bl[18] br[18] wl[427] vdd gnd cell_6t
Xbit_r428_c18 bl[18] br[18] wl[428] vdd gnd cell_6t
Xbit_r429_c18 bl[18] br[18] wl[429] vdd gnd cell_6t
Xbit_r430_c18 bl[18] br[18] wl[430] vdd gnd cell_6t
Xbit_r431_c18 bl[18] br[18] wl[431] vdd gnd cell_6t
Xbit_r432_c18 bl[18] br[18] wl[432] vdd gnd cell_6t
Xbit_r433_c18 bl[18] br[18] wl[433] vdd gnd cell_6t
Xbit_r434_c18 bl[18] br[18] wl[434] vdd gnd cell_6t
Xbit_r435_c18 bl[18] br[18] wl[435] vdd gnd cell_6t
Xbit_r436_c18 bl[18] br[18] wl[436] vdd gnd cell_6t
Xbit_r437_c18 bl[18] br[18] wl[437] vdd gnd cell_6t
Xbit_r438_c18 bl[18] br[18] wl[438] vdd gnd cell_6t
Xbit_r439_c18 bl[18] br[18] wl[439] vdd gnd cell_6t
Xbit_r440_c18 bl[18] br[18] wl[440] vdd gnd cell_6t
Xbit_r441_c18 bl[18] br[18] wl[441] vdd gnd cell_6t
Xbit_r442_c18 bl[18] br[18] wl[442] vdd gnd cell_6t
Xbit_r443_c18 bl[18] br[18] wl[443] vdd gnd cell_6t
Xbit_r444_c18 bl[18] br[18] wl[444] vdd gnd cell_6t
Xbit_r445_c18 bl[18] br[18] wl[445] vdd gnd cell_6t
Xbit_r446_c18 bl[18] br[18] wl[446] vdd gnd cell_6t
Xbit_r447_c18 bl[18] br[18] wl[447] vdd gnd cell_6t
Xbit_r448_c18 bl[18] br[18] wl[448] vdd gnd cell_6t
Xbit_r449_c18 bl[18] br[18] wl[449] vdd gnd cell_6t
Xbit_r450_c18 bl[18] br[18] wl[450] vdd gnd cell_6t
Xbit_r451_c18 bl[18] br[18] wl[451] vdd gnd cell_6t
Xbit_r452_c18 bl[18] br[18] wl[452] vdd gnd cell_6t
Xbit_r453_c18 bl[18] br[18] wl[453] vdd gnd cell_6t
Xbit_r454_c18 bl[18] br[18] wl[454] vdd gnd cell_6t
Xbit_r455_c18 bl[18] br[18] wl[455] vdd gnd cell_6t
Xbit_r456_c18 bl[18] br[18] wl[456] vdd gnd cell_6t
Xbit_r457_c18 bl[18] br[18] wl[457] vdd gnd cell_6t
Xbit_r458_c18 bl[18] br[18] wl[458] vdd gnd cell_6t
Xbit_r459_c18 bl[18] br[18] wl[459] vdd gnd cell_6t
Xbit_r460_c18 bl[18] br[18] wl[460] vdd gnd cell_6t
Xbit_r461_c18 bl[18] br[18] wl[461] vdd gnd cell_6t
Xbit_r462_c18 bl[18] br[18] wl[462] vdd gnd cell_6t
Xbit_r463_c18 bl[18] br[18] wl[463] vdd gnd cell_6t
Xbit_r464_c18 bl[18] br[18] wl[464] vdd gnd cell_6t
Xbit_r465_c18 bl[18] br[18] wl[465] vdd gnd cell_6t
Xbit_r466_c18 bl[18] br[18] wl[466] vdd gnd cell_6t
Xbit_r467_c18 bl[18] br[18] wl[467] vdd gnd cell_6t
Xbit_r468_c18 bl[18] br[18] wl[468] vdd gnd cell_6t
Xbit_r469_c18 bl[18] br[18] wl[469] vdd gnd cell_6t
Xbit_r470_c18 bl[18] br[18] wl[470] vdd gnd cell_6t
Xbit_r471_c18 bl[18] br[18] wl[471] vdd gnd cell_6t
Xbit_r472_c18 bl[18] br[18] wl[472] vdd gnd cell_6t
Xbit_r473_c18 bl[18] br[18] wl[473] vdd gnd cell_6t
Xbit_r474_c18 bl[18] br[18] wl[474] vdd gnd cell_6t
Xbit_r475_c18 bl[18] br[18] wl[475] vdd gnd cell_6t
Xbit_r476_c18 bl[18] br[18] wl[476] vdd gnd cell_6t
Xbit_r477_c18 bl[18] br[18] wl[477] vdd gnd cell_6t
Xbit_r478_c18 bl[18] br[18] wl[478] vdd gnd cell_6t
Xbit_r479_c18 bl[18] br[18] wl[479] vdd gnd cell_6t
Xbit_r480_c18 bl[18] br[18] wl[480] vdd gnd cell_6t
Xbit_r481_c18 bl[18] br[18] wl[481] vdd gnd cell_6t
Xbit_r482_c18 bl[18] br[18] wl[482] vdd gnd cell_6t
Xbit_r483_c18 bl[18] br[18] wl[483] vdd gnd cell_6t
Xbit_r484_c18 bl[18] br[18] wl[484] vdd gnd cell_6t
Xbit_r485_c18 bl[18] br[18] wl[485] vdd gnd cell_6t
Xbit_r486_c18 bl[18] br[18] wl[486] vdd gnd cell_6t
Xbit_r487_c18 bl[18] br[18] wl[487] vdd gnd cell_6t
Xbit_r488_c18 bl[18] br[18] wl[488] vdd gnd cell_6t
Xbit_r489_c18 bl[18] br[18] wl[489] vdd gnd cell_6t
Xbit_r490_c18 bl[18] br[18] wl[490] vdd gnd cell_6t
Xbit_r491_c18 bl[18] br[18] wl[491] vdd gnd cell_6t
Xbit_r492_c18 bl[18] br[18] wl[492] vdd gnd cell_6t
Xbit_r493_c18 bl[18] br[18] wl[493] vdd gnd cell_6t
Xbit_r494_c18 bl[18] br[18] wl[494] vdd gnd cell_6t
Xbit_r495_c18 bl[18] br[18] wl[495] vdd gnd cell_6t
Xbit_r496_c18 bl[18] br[18] wl[496] vdd gnd cell_6t
Xbit_r497_c18 bl[18] br[18] wl[497] vdd gnd cell_6t
Xbit_r498_c18 bl[18] br[18] wl[498] vdd gnd cell_6t
Xbit_r499_c18 bl[18] br[18] wl[499] vdd gnd cell_6t
Xbit_r500_c18 bl[18] br[18] wl[500] vdd gnd cell_6t
Xbit_r501_c18 bl[18] br[18] wl[501] vdd gnd cell_6t
Xbit_r502_c18 bl[18] br[18] wl[502] vdd gnd cell_6t
Xbit_r503_c18 bl[18] br[18] wl[503] vdd gnd cell_6t
Xbit_r504_c18 bl[18] br[18] wl[504] vdd gnd cell_6t
Xbit_r505_c18 bl[18] br[18] wl[505] vdd gnd cell_6t
Xbit_r506_c18 bl[18] br[18] wl[506] vdd gnd cell_6t
Xbit_r507_c18 bl[18] br[18] wl[507] vdd gnd cell_6t
Xbit_r508_c18 bl[18] br[18] wl[508] vdd gnd cell_6t
Xbit_r509_c18 bl[18] br[18] wl[509] vdd gnd cell_6t
Xbit_r510_c18 bl[18] br[18] wl[510] vdd gnd cell_6t
Xbit_r511_c18 bl[18] br[18] wl[511] vdd gnd cell_6t
Xbit_r0_c19 bl[19] br[19] wl[0] vdd gnd cell_6t
Xbit_r1_c19 bl[19] br[19] wl[1] vdd gnd cell_6t
Xbit_r2_c19 bl[19] br[19] wl[2] vdd gnd cell_6t
Xbit_r3_c19 bl[19] br[19] wl[3] vdd gnd cell_6t
Xbit_r4_c19 bl[19] br[19] wl[4] vdd gnd cell_6t
Xbit_r5_c19 bl[19] br[19] wl[5] vdd gnd cell_6t
Xbit_r6_c19 bl[19] br[19] wl[6] vdd gnd cell_6t
Xbit_r7_c19 bl[19] br[19] wl[7] vdd gnd cell_6t
Xbit_r8_c19 bl[19] br[19] wl[8] vdd gnd cell_6t
Xbit_r9_c19 bl[19] br[19] wl[9] vdd gnd cell_6t
Xbit_r10_c19 bl[19] br[19] wl[10] vdd gnd cell_6t
Xbit_r11_c19 bl[19] br[19] wl[11] vdd gnd cell_6t
Xbit_r12_c19 bl[19] br[19] wl[12] vdd gnd cell_6t
Xbit_r13_c19 bl[19] br[19] wl[13] vdd gnd cell_6t
Xbit_r14_c19 bl[19] br[19] wl[14] vdd gnd cell_6t
Xbit_r15_c19 bl[19] br[19] wl[15] vdd gnd cell_6t
Xbit_r16_c19 bl[19] br[19] wl[16] vdd gnd cell_6t
Xbit_r17_c19 bl[19] br[19] wl[17] vdd gnd cell_6t
Xbit_r18_c19 bl[19] br[19] wl[18] vdd gnd cell_6t
Xbit_r19_c19 bl[19] br[19] wl[19] vdd gnd cell_6t
Xbit_r20_c19 bl[19] br[19] wl[20] vdd gnd cell_6t
Xbit_r21_c19 bl[19] br[19] wl[21] vdd gnd cell_6t
Xbit_r22_c19 bl[19] br[19] wl[22] vdd gnd cell_6t
Xbit_r23_c19 bl[19] br[19] wl[23] vdd gnd cell_6t
Xbit_r24_c19 bl[19] br[19] wl[24] vdd gnd cell_6t
Xbit_r25_c19 bl[19] br[19] wl[25] vdd gnd cell_6t
Xbit_r26_c19 bl[19] br[19] wl[26] vdd gnd cell_6t
Xbit_r27_c19 bl[19] br[19] wl[27] vdd gnd cell_6t
Xbit_r28_c19 bl[19] br[19] wl[28] vdd gnd cell_6t
Xbit_r29_c19 bl[19] br[19] wl[29] vdd gnd cell_6t
Xbit_r30_c19 bl[19] br[19] wl[30] vdd gnd cell_6t
Xbit_r31_c19 bl[19] br[19] wl[31] vdd gnd cell_6t
Xbit_r32_c19 bl[19] br[19] wl[32] vdd gnd cell_6t
Xbit_r33_c19 bl[19] br[19] wl[33] vdd gnd cell_6t
Xbit_r34_c19 bl[19] br[19] wl[34] vdd gnd cell_6t
Xbit_r35_c19 bl[19] br[19] wl[35] vdd gnd cell_6t
Xbit_r36_c19 bl[19] br[19] wl[36] vdd gnd cell_6t
Xbit_r37_c19 bl[19] br[19] wl[37] vdd gnd cell_6t
Xbit_r38_c19 bl[19] br[19] wl[38] vdd gnd cell_6t
Xbit_r39_c19 bl[19] br[19] wl[39] vdd gnd cell_6t
Xbit_r40_c19 bl[19] br[19] wl[40] vdd gnd cell_6t
Xbit_r41_c19 bl[19] br[19] wl[41] vdd gnd cell_6t
Xbit_r42_c19 bl[19] br[19] wl[42] vdd gnd cell_6t
Xbit_r43_c19 bl[19] br[19] wl[43] vdd gnd cell_6t
Xbit_r44_c19 bl[19] br[19] wl[44] vdd gnd cell_6t
Xbit_r45_c19 bl[19] br[19] wl[45] vdd gnd cell_6t
Xbit_r46_c19 bl[19] br[19] wl[46] vdd gnd cell_6t
Xbit_r47_c19 bl[19] br[19] wl[47] vdd gnd cell_6t
Xbit_r48_c19 bl[19] br[19] wl[48] vdd gnd cell_6t
Xbit_r49_c19 bl[19] br[19] wl[49] vdd gnd cell_6t
Xbit_r50_c19 bl[19] br[19] wl[50] vdd gnd cell_6t
Xbit_r51_c19 bl[19] br[19] wl[51] vdd gnd cell_6t
Xbit_r52_c19 bl[19] br[19] wl[52] vdd gnd cell_6t
Xbit_r53_c19 bl[19] br[19] wl[53] vdd gnd cell_6t
Xbit_r54_c19 bl[19] br[19] wl[54] vdd gnd cell_6t
Xbit_r55_c19 bl[19] br[19] wl[55] vdd gnd cell_6t
Xbit_r56_c19 bl[19] br[19] wl[56] vdd gnd cell_6t
Xbit_r57_c19 bl[19] br[19] wl[57] vdd gnd cell_6t
Xbit_r58_c19 bl[19] br[19] wl[58] vdd gnd cell_6t
Xbit_r59_c19 bl[19] br[19] wl[59] vdd gnd cell_6t
Xbit_r60_c19 bl[19] br[19] wl[60] vdd gnd cell_6t
Xbit_r61_c19 bl[19] br[19] wl[61] vdd gnd cell_6t
Xbit_r62_c19 bl[19] br[19] wl[62] vdd gnd cell_6t
Xbit_r63_c19 bl[19] br[19] wl[63] vdd gnd cell_6t
Xbit_r64_c19 bl[19] br[19] wl[64] vdd gnd cell_6t
Xbit_r65_c19 bl[19] br[19] wl[65] vdd gnd cell_6t
Xbit_r66_c19 bl[19] br[19] wl[66] vdd gnd cell_6t
Xbit_r67_c19 bl[19] br[19] wl[67] vdd gnd cell_6t
Xbit_r68_c19 bl[19] br[19] wl[68] vdd gnd cell_6t
Xbit_r69_c19 bl[19] br[19] wl[69] vdd gnd cell_6t
Xbit_r70_c19 bl[19] br[19] wl[70] vdd gnd cell_6t
Xbit_r71_c19 bl[19] br[19] wl[71] vdd gnd cell_6t
Xbit_r72_c19 bl[19] br[19] wl[72] vdd gnd cell_6t
Xbit_r73_c19 bl[19] br[19] wl[73] vdd gnd cell_6t
Xbit_r74_c19 bl[19] br[19] wl[74] vdd gnd cell_6t
Xbit_r75_c19 bl[19] br[19] wl[75] vdd gnd cell_6t
Xbit_r76_c19 bl[19] br[19] wl[76] vdd gnd cell_6t
Xbit_r77_c19 bl[19] br[19] wl[77] vdd gnd cell_6t
Xbit_r78_c19 bl[19] br[19] wl[78] vdd gnd cell_6t
Xbit_r79_c19 bl[19] br[19] wl[79] vdd gnd cell_6t
Xbit_r80_c19 bl[19] br[19] wl[80] vdd gnd cell_6t
Xbit_r81_c19 bl[19] br[19] wl[81] vdd gnd cell_6t
Xbit_r82_c19 bl[19] br[19] wl[82] vdd gnd cell_6t
Xbit_r83_c19 bl[19] br[19] wl[83] vdd gnd cell_6t
Xbit_r84_c19 bl[19] br[19] wl[84] vdd gnd cell_6t
Xbit_r85_c19 bl[19] br[19] wl[85] vdd gnd cell_6t
Xbit_r86_c19 bl[19] br[19] wl[86] vdd gnd cell_6t
Xbit_r87_c19 bl[19] br[19] wl[87] vdd gnd cell_6t
Xbit_r88_c19 bl[19] br[19] wl[88] vdd gnd cell_6t
Xbit_r89_c19 bl[19] br[19] wl[89] vdd gnd cell_6t
Xbit_r90_c19 bl[19] br[19] wl[90] vdd gnd cell_6t
Xbit_r91_c19 bl[19] br[19] wl[91] vdd gnd cell_6t
Xbit_r92_c19 bl[19] br[19] wl[92] vdd gnd cell_6t
Xbit_r93_c19 bl[19] br[19] wl[93] vdd gnd cell_6t
Xbit_r94_c19 bl[19] br[19] wl[94] vdd gnd cell_6t
Xbit_r95_c19 bl[19] br[19] wl[95] vdd gnd cell_6t
Xbit_r96_c19 bl[19] br[19] wl[96] vdd gnd cell_6t
Xbit_r97_c19 bl[19] br[19] wl[97] vdd gnd cell_6t
Xbit_r98_c19 bl[19] br[19] wl[98] vdd gnd cell_6t
Xbit_r99_c19 bl[19] br[19] wl[99] vdd gnd cell_6t
Xbit_r100_c19 bl[19] br[19] wl[100] vdd gnd cell_6t
Xbit_r101_c19 bl[19] br[19] wl[101] vdd gnd cell_6t
Xbit_r102_c19 bl[19] br[19] wl[102] vdd gnd cell_6t
Xbit_r103_c19 bl[19] br[19] wl[103] vdd gnd cell_6t
Xbit_r104_c19 bl[19] br[19] wl[104] vdd gnd cell_6t
Xbit_r105_c19 bl[19] br[19] wl[105] vdd gnd cell_6t
Xbit_r106_c19 bl[19] br[19] wl[106] vdd gnd cell_6t
Xbit_r107_c19 bl[19] br[19] wl[107] vdd gnd cell_6t
Xbit_r108_c19 bl[19] br[19] wl[108] vdd gnd cell_6t
Xbit_r109_c19 bl[19] br[19] wl[109] vdd gnd cell_6t
Xbit_r110_c19 bl[19] br[19] wl[110] vdd gnd cell_6t
Xbit_r111_c19 bl[19] br[19] wl[111] vdd gnd cell_6t
Xbit_r112_c19 bl[19] br[19] wl[112] vdd gnd cell_6t
Xbit_r113_c19 bl[19] br[19] wl[113] vdd gnd cell_6t
Xbit_r114_c19 bl[19] br[19] wl[114] vdd gnd cell_6t
Xbit_r115_c19 bl[19] br[19] wl[115] vdd gnd cell_6t
Xbit_r116_c19 bl[19] br[19] wl[116] vdd gnd cell_6t
Xbit_r117_c19 bl[19] br[19] wl[117] vdd gnd cell_6t
Xbit_r118_c19 bl[19] br[19] wl[118] vdd gnd cell_6t
Xbit_r119_c19 bl[19] br[19] wl[119] vdd gnd cell_6t
Xbit_r120_c19 bl[19] br[19] wl[120] vdd gnd cell_6t
Xbit_r121_c19 bl[19] br[19] wl[121] vdd gnd cell_6t
Xbit_r122_c19 bl[19] br[19] wl[122] vdd gnd cell_6t
Xbit_r123_c19 bl[19] br[19] wl[123] vdd gnd cell_6t
Xbit_r124_c19 bl[19] br[19] wl[124] vdd gnd cell_6t
Xbit_r125_c19 bl[19] br[19] wl[125] vdd gnd cell_6t
Xbit_r126_c19 bl[19] br[19] wl[126] vdd gnd cell_6t
Xbit_r127_c19 bl[19] br[19] wl[127] vdd gnd cell_6t
Xbit_r128_c19 bl[19] br[19] wl[128] vdd gnd cell_6t
Xbit_r129_c19 bl[19] br[19] wl[129] vdd gnd cell_6t
Xbit_r130_c19 bl[19] br[19] wl[130] vdd gnd cell_6t
Xbit_r131_c19 bl[19] br[19] wl[131] vdd gnd cell_6t
Xbit_r132_c19 bl[19] br[19] wl[132] vdd gnd cell_6t
Xbit_r133_c19 bl[19] br[19] wl[133] vdd gnd cell_6t
Xbit_r134_c19 bl[19] br[19] wl[134] vdd gnd cell_6t
Xbit_r135_c19 bl[19] br[19] wl[135] vdd gnd cell_6t
Xbit_r136_c19 bl[19] br[19] wl[136] vdd gnd cell_6t
Xbit_r137_c19 bl[19] br[19] wl[137] vdd gnd cell_6t
Xbit_r138_c19 bl[19] br[19] wl[138] vdd gnd cell_6t
Xbit_r139_c19 bl[19] br[19] wl[139] vdd gnd cell_6t
Xbit_r140_c19 bl[19] br[19] wl[140] vdd gnd cell_6t
Xbit_r141_c19 bl[19] br[19] wl[141] vdd gnd cell_6t
Xbit_r142_c19 bl[19] br[19] wl[142] vdd gnd cell_6t
Xbit_r143_c19 bl[19] br[19] wl[143] vdd gnd cell_6t
Xbit_r144_c19 bl[19] br[19] wl[144] vdd gnd cell_6t
Xbit_r145_c19 bl[19] br[19] wl[145] vdd gnd cell_6t
Xbit_r146_c19 bl[19] br[19] wl[146] vdd gnd cell_6t
Xbit_r147_c19 bl[19] br[19] wl[147] vdd gnd cell_6t
Xbit_r148_c19 bl[19] br[19] wl[148] vdd gnd cell_6t
Xbit_r149_c19 bl[19] br[19] wl[149] vdd gnd cell_6t
Xbit_r150_c19 bl[19] br[19] wl[150] vdd gnd cell_6t
Xbit_r151_c19 bl[19] br[19] wl[151] vdd gnd cell_6t
Xbit_r152_c19 bl[19] br[19] wl[152] vdd gnd cell_6t
Xbit_r153_c19 bl[19] br[19] wl[153] vdd gnd cell_6t
Xbit_r154_c19 bl[19] br[19] wl[154] vdd gnd cell_6t
Xbit_r155_c19 bl[19] br[19] wl[155] vdd gnd cell_6t
Xbit_r156_c19 bl[19] br[19] wl[156] vdd gnd cell_6t
Xbit_r157_c19 bl[19] br[19] wl[157] vdd gnd cell_6t
Xbit_r158_c19 bl[19] br[19] wl[158] vdd gnd cell_6t
Xbit_r159_c19 bl[19] br[19] wl[159] vdd gnd cell_6t
Xbit_r160_c19 bl[19] br[19] wl[160] vdd gnd cell_6t
Xbit_r161_c19 bl[19] br[19] wl[161] vdd gnd cell_6t
Xbit_r162_c19 bl[19] br[19] wl[162] vdd gnd cell_6t
Xbit_r163_c19 bl[19] br[19] wl[163] vdd gnd cell_6t
Xbit_r164_c19 bl[19] br[19] wl[164] vdd gnd cell_6t
Xbit_r165_c19 bl[19] br[19] wl[165] vdd gnd cell_6t
Xbit_r166_c19 bl[19] br[19] wl[166] vdd gnd cell_6t
Xbit_r167_c19 bl[19] br[19] wl[167] vdd gnd cell_6t
Xbit_r168_c19 bl[19] br[19] wl[168] vdd gnd cell_6t
Xbit_r169_c19 bl[19] br[19] wl[169] vdd gnd cell_6t
Xbit_r170_c19 bl[19] br[19] wl[170] vdd gnd cell_6t
Xbit_r171_c19 bl[19] br[19] wl[171] vdd gnd cell_6t
Xbit_r172_c19 bl[19] br[19] wl[172] vdd gnd cell_6t
Xbit_r173_c19 bl[19] br[19] wl[173] vdd gnd cell_6t
Xbit_r174_c19 bl[19] br[19] wl[174] vdd gnd cell_6t
Xbit_r175_c19 bl[19] br[19] wl[175] vdd gnd cell_6t
Xbit_r176_c19 bl[19] br[19] wl[176] vdd gnd cell_6t
Xbit_r177_c19 bl[19] br[19] wl[177] vdd gnd cell_6t
Xbit_r178_c19 bl[19] br[19] wl[178] vdd gnd cell_6t
Xbit_r179_c19 bl[19] br[19] wl[179] vdd gnd cell_6t
Xbit_r180_c19 bl[19] br[19] wl[180] vdd gnd cell_6t
Xbit_r181_c19 bl[19] br[19] wl[181] vdd gnd cell_6t
Xbit_r182_c19 bl[19] br[19] wl[182] vdd gnd cell_6t
Xbit_r183_c19 bl[19] br[19] wl[183] vdd gnd cell_6t
Xbit_r184_c19 bl[19] br[19] wl[184] vdd gnd cell_6t
Xbit_r185_c19 bl[19] br[19] wl[185] vdd gnd cell_6t
Xbit_r186_c19 bl[19] br[19] wl[186] vdd gnd cell_6t
Xbit_r187_c19 bl[19] br[19] wl[187] vdd gnd cell_6t
Xbit_r188_c19 bl[19] br[19] wl[188] vdd gnd cell_6t
Xbit_r189_c19 bl[19] br[19] wl[189] vdd gnd cell_6t
Xbit_r190_c19 bl[19] br[19] wl[190] vdd gnd cell_6t
Xbit_r191_c19 bl[19] br[19] wl[191] vdd gnd cell_6t
Xbit_r192_c19 bl[19] br[19] wl[192] vdd gnd cell_6t
Xbit_r193_c19 bl[19] br[19] wl[193] vdd gnd cell_6t
Xbit_r194_c19 bl[19] br[19] wl[194] vdd gnd cell_6t
Xbit_r195_c19 bl[19] br[19] wl[195] vdd gnd cell_6t
Xbit_r196_c19 bl[19] br[19] wl[196] vdd gnd cell_6t
Xbit_r197_c19 bl[19] br[19] wl[197] vdd gnd cell_6t
Xbit_r198_c19 bl[19] br[19] wl[198] vdd gnd cell_6t
Xbit_r199_c19 bl[19] br[19] wl[199] vdd gnd cell_6t
Xbit_r200_c19 bl[19] br[19] wl[200] vdd gnd cell_6t
Xbit_r201_c19 bl[19] br[19] wl[201] vdd gnd cell_6t
Xbit_r202_c19 bl[19] br[19] wl[202] vdd gnd cell_6t
Xbit_r203_c19 bl[19] br[19] wl[203] vdd gnd cell_6t
Xbit_r204_c19 bl[19] br[19] wl[204] vdd gnd cell_6t
Xbit_r205_c19 bl[19] br[19] wl[205] vdd gnd cell_6t
Xbit_r206_c19 bl[19] br[19] wl[206] vdd gnd cell_6t
Xbit_r207_c19 bl[19] br[19] wl[207] vdd gnd cell_6t
Xbit_r208_c19 bl[19] br[19] wl[208] vdd gnd cell_6t
Xbit_r209_c19 bl[19] br[19] wl[209] vdd gnd cell_6t
Xbit_r210_c19 bl[19] br[19] wl[210] vdd gnd cell_6t
Xbit_r211_c19 bl[19] br[19] wl[211] vdd gnd cell_6t
Xbit_r212_c19 bl[19] br[19] wl[212] vdd gnd cell_6t
Xbit_r213_c19 bl[19] br[19] wl[213] vdd gnd cell_6t
Xbit_r214_c19 bl[19] br[19] wl[214] vdd gnd cell_6t
Xbit_r215_c19 bl[19] br[19] wl[215] vdd gnd cell_6t
Xbit_r216_c19 bl[19] br[19] wl[216] vdd gnd cell_6t
Xbit_r217_c19 bl[19] br[19] wl[217] vdd gnd cell_6t
Xbit_r218_c19 bl[19] br[19] wl[218] vdd gnd cell_6t
Xbit_r219_c19 bl[19] br[19] wl[219] vdd gnd cell_6t
Xbit_r220_c19 bl[19] br[19] wl[220] vdd gnd cell_6t
Xbit_r221_c19 bl[19] br[19] wl[221] vdd gnd cell_6t
Xbit_r222_c19 bl[19] br[19] wl[222] vdd gnd cell_6t
Xbit_r223_c19 bl[19] br[19] wl[223] vdd gnd cell_6t
Xbit_r224_c19 bl[19] br[19] wl[224] vdd gnd cell_6t
Xbit_r225_c19 bl[19] br[19] wl[225] vdd gnd cell_6t
Xbit_r226_c19 bl[19] br[19] wl[226] vdd gnd cell_6t
Xbit_r227_c19 bl[19] br[19] wl[227] vdd gnd cell_6t
Xbit_r228_c19 bl[19] br[19] wl[228] vdd gnd cell_6t
Xbit_r229_c19 bl[19] br[19] wl[229] vdd gnd cell_6t
Xbit_r230_c19 bl[19] br[19] wl[230] vdd gnd cell_6t
Xbit_r231_c19 bl[19] br[19] wl[231] vdd gnd cell_6t
Xbit_r232_c19 bl[19] br[19] wl[232] vdd gnd cell_6t
Xbit_r233_c19 bl[19] br[19] wl[233] vdd gnd cell_6t
Xbit_r234_c19 bl[19] br[19] wl[234] vdd gnd cell_6t
Xbit_r235_c19 bl[19] br[19] wl[235] vdd gnd cell_6t
Xbit_r236_c19 bl[19] br[19] wl[236] vdd gnd cell_6t
Xbit_r237_c19 bl[19] br[19] wl[237] vdd gnd cell_6t
Xbit_r238_c19 bl[19] br[19] wl[238] vdd gnd cell_6t
Xbit_r239_c19 bl[19] br[19] wl[239] vdd gnd cell_6t
Xbit_r240_c19 bl[19] br[19] wl[240] vdd gnd cell_6t
Xbit_r241_c19 bl[19] br[19] wl[241] vdd gnd cell_6t
Xbit_r242_c19 bl[19] br[19] wl[242] vdd gnd cell_6t
Xbit_r243_c19 bl[19] br[19] wl[243] vdd gnd cell_6t
Xbit_r244_c19 bl[19] br[19] wl[244] vdd gnd cell_6t
Xbit_r245_c19 bl[19] br[19] wl[245] vdd gnd cell_6t
Xbit_r246_c19 bl[19] br[19] wl[246] vdd gnd cell_6t
Xbit_r247_c19 bl[19] br[19] wl[247] vdd gnd cell_6t
Xbit_r248_c19 bl[19] br[19] wl[248] vdd gnd cell_6t
Xbit_r249_c19 bl[19] br[19] wl[249] vdd gnd cell_6t
Xbit_r250_c19 bl[19] br[19] wl[250] vdd gnd cell_6t
Xbit_r251_c19 bl[19] br[19] wl[251] vdd gnd cell_6t
Xbit_r252_c19 bl[19] br[19] wl[252] vdd gnd cell_6t
Xbit_r253_c19 bl[19] br[19] wl[253] vdd gnd cell_6t
Xbit_r254_c19 bl[19] br[19] wl[254] vdd gnd cell_6t
Xbit_r255_c19 bl[19] br[19] wl[255] vdd gnd cell_6t
Xbit_r256_c19 bl[19] br[19] wl[256] vdd gnd cell_6t
Xbit_r257_c19 bl[19] br[19] wl[257] vdd gnd cell_6t
Xbit_r258_c19 bl[19] br[19] wl[258] vdd gnd cell_6t
Xbit_r259_c19 bl[19] br[19] wl[259] vdd gnd cell_6t
Xbit_r260_c19 bl[19] br[19] wl[260] vdd gnd cell_6t
Xbit_r261_c19 bl[19] br[19] wl[261] vdd gnd cell_6t
Xbit_r262_c19 bl[19] br[19] wl[262] vdd gnd cell_6t
Xbit_r263_c19 bl[19] br[19] wl[263] vdd gnd cell_6t
Xbit_r264_c19 bl[19] br[19] wl[264] vdd gnd cell_6t
Xbit_r265_c19 bl[19] br[19] wl[265] vdd gnd cell_6t
Xbit_r266_c19 bl[19] br[19] wl[266] vdd gnd cell_6t
Xbit_r267_c19 bl[19] br[19] wl[267] vdd gnd cell_6t
Xbit_r268_c19 bl[19] br[19] wl[268] vdd gnd cell_6t
Xbit_r269_c19 bl[19] br[19] wl[269] vdd gnd cell_6t
Xbit_r270_c19 bl[19] br[19] wl[270] vdd gnd cell_6t
Xbit_r271_c19 bl[19] br[19] wl[271] vdd gnd cell_6t
Xbit_r272_c19 bl[19] br[19] wl[272] vdd gnd cell_6t
Xbit_r273_c19 bl[19] br[19] wl[273] vdd gnd cell_6t
Xbit_r274_c19 bl[19] br[19] wl[274] vdd gnd cell_6t
Xbit_r275_c19 bl[19] br[19] wl[275] vdd gnd cell_6t
Xbit_r276_c19 bl[19] br[19] wl[276] vdd gnd cell_6t
Xbit_r277_c19 bl[19] br[19] wl[277] vdd gnd cell_6t
Xbit_r278_c19 bl[19] br[19] wl[278] vdd gnd cell_6t
Xbit_r279_c19 bl[19] br[19] wl[279] vdd gnd cell_6t
Xbit_r280_c19 bl[19] br[19] wl[280] vdd gnd cell_6t
Xbit_r281_c19 bl[19] br[19] wl[281] vdd gnd cell_6t
Xbit_r282_c19 bl[19] br[19] wl[282] vdd gnd cell_6t
Xbit_r283_c19 bl[19] br[19] wl[283] vdd gnd cell_6t
Xbit_r284_c19 bl[19] br[19] wl[284] vdd gnd cell_6t
Xbit_r285_c19 bl[19] br[19] wl[285] vdd gnd cell_6t
Xbit_r286_c19 bl[19] br[19] wl[286] vdd gnd cell_6t
Xbit_r287_c19 bl[19] br[19] wl[287] vdd gnd cell_6t
Xbit_r288_c19 bl[19] br[19] wl[288] vdd gnd cell_6t
Xbit_r289_c19 bl[19] br[19] wl[289] vdd gnd cell_6t
Xbit_r290_c19 bl[19] br[19] wl[290] vdd gnd cell_6t
Xbit_r291_c19 bl[19] br[19] wl[291] vdd gnd cell_6t
Xbit_r292_c19 bl[19] br[19] wl[292] vdd gnd cell_6t
Xbit_r293_c19 bl[19] br[19] wl[293] vdd gnd cell_6t
Xbit_r294_c19 bl[19] br[19] wl[294] vdd gnd cell_6t
Xbit_r295_c19 bl[19] br[19] wl[295] vdd gnd cell_6t
Xbit_r296_c19 bl[19] br[19] wl[296] vdd gnd cell_6t
Xbit_r297_c19 bl[19] br[19] wl[297] vdd gnd cell_6t
Xbit_r298_c19 bl[19] br[19] wl[298] vdd gnd cell_6t
Xbit_r299_c19 bl[19] br[19] wl[299] vdd gnd cell_6t
Xbit_r300_c19 bl[19] br[19] wl[300] vdd gnd cell_6t
Xbit_r301_c19 bl[19] br[19] wl[301] vdd gnd cell_6t
Xbit_r302_c19 bl[19] br[19] wl[302] vdd gnd cell_6t
Xbit_r303_c19 bl[19] br[19] wl[303] vdd gnd cell_6t
Xbit_r304_c19 bl[19] br[19] wl[304] vdd gnd cell_6t
Xbit_r305_c19 bl[19] br[19] wl[305] vdd gnd cell_6t
Xbit_r306_c19 bl[19] br[19] wl[306] vdd gnd cell_6t
Xbit_r307_c19 bl[19] br[19] wl[307] vdd gnd cell_6t
Xbit_r308_c19 bl[19] br[19] wl[308] vdd gnd cell_6t
Xbit_r309_c19 bl[19] br[19] wl[309] vdd gnd cell_6t
Xbit_r310_c19 bl[19] br[19] wl[310] vdd gnd cell_6t
Xbit_r311_c19 bl[19] br[19] wl[311] vdd gnd cell_6t
Xbit_r312_c19 bl[19] br[19] wl[312] vdd gnd cell_6t
Xbit_r313_c19 bl[19] br[19] wl[313] vdd gnd cell_6t
Xbit_r314_c19 bl[19] br[19] wl[314] vdd gnd cell_6t
Xbit_r315_c19 bl[19] br[19] wl[315] vdd gnd cell_6t
Xbit_r316_c19 bl[19] br[19] wl[316] vdd gnd cell_6t
Xbit_r317_c19 bl[19] br[19] wl[317] vdd gnd cell_6t
Xbit_r318_c19 bl[19] br[19] wl[318] vdd gnd cell_6t
Xbit_r319_c19 bl[19] br[19] wl[319] vdd gnd cell_6t
Xbit_r320_c19 bl[19] br[19] wl[320] vdd gnd cell_6t
Xbit_r321_c19 bl[19] br[19] wl[321] vdd gnd cell_6t
Xbit_r322_c19 bl[19] br[19] wl[322] vdd gnd cell_6t
Xbit_r323_c19 bl[19] br[19] wl[323] vdd gnd cell_6t
Xbit_r324_c19 bl[19] br[19] wl[324] vdd gnd cell_6t
Xbit_r325_c19 bl[19] br[19] wl[325] vdd gnd cell_6t
Xbit_r326_c19 bl[19] br[19] wl[326] vdd gnd cell_6t
Xbit_r327_c19 bl[19] br[19] wl[327] vdd gnd cell_6t
Xbit_r328_c19 bl[19] br[19] wl[328] vdd gnd cell_6t
Xbit_r329_c19 bl[19] br[19] wl[329] vdd gnd cell_6t
Xbit_r330_c19 bl[19] br[19] wl[330] vdd gnd cell_6t
Xbit_r331_c19 bl[19] br[19] wl[331] vdd gnd cell_6t
Xbit_r332_c19 bl[19] br[19] wl[332] vdd gnd cell_6t
Xbit_r333_c19 bl[19] br[19] wl[333] vdd gnd cell_6t
Xbit_r334_c19 bl[19] br[19] wl[334] vdd gnd cell_6t
Xbit_r335_c19 bl[19] br[19] wl[335] vdd gnd cell_6t
Xbit_r336_c19 bl[19] br[19] wl[336] vdd gnd cell_6t
Xbit_r337_c19 bl[19] br[19] wl[337] vdd gnd cell_6t
Xbit_r338_c19 bl[19] br[19] wl[338] vdd gnd cell_6t
Xbit_r339_c19 bl[19] br[19] wl[339] vdd gnd cell_6t
Xbit_r340_c19 bl[19] br[19] wl[340] vdd gnd cell_6t
Xbit_r341_c19 bl[19] br[19] wl[341] vdd gnd cell_6t
Xbit_r342_c19 bl[19] br[19] wl[342] vdd gnd cell_6t
Xbit_r343_c19 bl[19] br[19] wl[343] vdd gnd cell_6t
Xbit_r344_c19 bl[19] br[19] wl[344] vdd gnd cell_6t
Xbit_r345_c19 bl[19] br[19] wl[345] vdd gnd cell_6t
Xbit_r346_c19 bl[19] br[19] wl[346] vdd gnd cell_6t
Xbit_r347_c19 bl[19] br[19] wl[347] vdd gnd cell_6t
Xbit_r348_c19 bl[19] br[19] wl[348] vdd gnd cell_6t
Xbit_r349_c19 bl[19] br[19] wl[349] vdd gnd cell_6t
Xbit_r350_c19 bl[19] br[19] wl[350] vdd gnd cell_6t
Xbit_r351_c19 bl[19] br[19] wl[351] vdd gnd cell_6t
Xbit_r352_c19 bl[19] br[19] wl[352] vdd gnd cell_6t
Xbit_r353_c19 bl[19] br[19] wl[353] vdd gnd cell_6t
Xbit_r354_c19 bl[19] br[19] wl[354] vdd gnd cell_6t
Xbit_r355_c19 bl[19] br[19] wl[355] vdd gnd cell_6t
Xbit_r356_c19 bl[19] br[19] wl[356] vdd gnd cell_6t
Xbit_r357_c19 bl[19] br[19] wl[357] vdd gnd cell_6t
Xbit_r358_c19 bl[19] br[19] wl[358] vdd gnd cell_6t
Xbit_r359_c19 bl[19] br[19] wl[359] vdd gnd cell_6t
Xbit_r360_c19 bl[19] br[19] wl[360] vdd gnd cell_6t
Xbit_r361_c19 bl[19] br[19] wl[361] vdd gnd cell_6t
Xbit_r362_c19 bl[19] br[19] wl[362] vdd gnd cell_6t
Xbit_r363_c19 bl[19] br[19] wl[363] vdd gnd cell_6t
Xbit_r364_c19 bl[19] br[19] wl[364] vdd gnd cell_6t
Xbit_r365_c19 bl[19] br[19] wl[365] vdd gnd cell_6t
Xbit_r366_c19 bl[19] br[19] wl[366] vdd gnd cell_6t
Xbit_r367_c19 bl[19] br[19] wl[367] vdd gnd cell_6t
Xbit_r368_c19 bl[19] br[19] wl[368] vdd gnd cell_6t
Xbit_r369_c19 bl[19] br[19] wl[369] vdd gnd cell_6t
Xbit_r370_c19 bl[19] br[19] wl[370] vdd gnd cell_6t
Xbit_r371_c19 bl[19] br[19] wl[371] vdd gnd cell_6t
Xbit_r372_c19 bl[19] br[19] wl[372] vdd gnd cell_6t
Xbit_r373_c19 bl[19] br[19] wl[373] vdd gnd cell_6t
Xbit_r374_c19 bl[19] br[19] wl[374] vdd gnd cell_6t
Xbit_r375_c19 bl[19] br[19] wl[375] vdd gnd cell_6t
Xbit_r376_c19 bl[19] br[19] wl[376] vdd gnd cell_6t
Xbit_r377_c19 bl[19] br[19] wl[377] vdd gnd cell_6t
Xbit_r378_c19 bl[19] br[19] wl[378] vdd gnd cell_6t
Xbit_r379_c19 bl[19] br[19] wl[379] vdd gnd cell_6t
Xbit_r380_c19 bl[19] br[19] wl[380] vdd gnd cell_6t
Xbit_r381_c19 bl[19] br[19] wl[381] vdd gnd cell_6t
Xbit_r382_c19 bl[19] br[19] wl[382] vdd gnd cell_6t
Xbit_r383_c19 bl[19] br[19] wl[383] vdd gnd cell_6t
Xbit_r384_c19 bl[19] br[19] wl[384] vdd gnd cell_6t
Xbit_r385_c19 bl[19] br[19] wl[385] vdd gnd cell_6t
Xbit_r386_c19 bl[19] br[19] wl[386] vdd gnd cell_6t
Xbit_r387_c19 bl[19] br[19] wl[387] vdd gnd cell_6t
Xbit_r388_c19 bl[19] br[19] wl[388] vdd gnd cell_6t
Xbit_r389_c19 bl[19] br[19] wl[389] vdd gnd cell_6t
Xbit_r390_c19 bl[19] br[19] wl[390] vdd gnd cell_6t
Xbit_r391_c19 bl[19] br[19] wl[391] vdd gnd cell_6t
Xbit_r392_c19 bl[19] br[19] wl[392] vdd gnd cell_6t
Xbit_r393_c19 bl[19] br[19] wl[393] vdd gnd cell_6t
Xbit_r394_c19 bl[19] br[19] wl[394] vdd gnd cell_6t
Xbit_r395_c19 bl[19] br[19] wl[395] vdd gnd cell_6t
Xbit_r396_c19 bl[19] br[19] wl[396] vdd gnd cell_6t
Xbit_r397_c19 bl[19] br[19] wl[397] vdd gnd cell_6t
Xbit_r398_c19 bl[19] br[19] wl[398] vdd gnd cell_6t
Xbit_r399_c19 bl[19] br[19] wl[399] vdd gnd cell_6t
Xbit_r400_c19 bl[19] br[19] wl[400] vdd gnd cell_6t
Xbit_r401_c19 bl[19] br[19] wl[401] vdd gnd cell_6t
Xbit_r402_c19 bl[19] br[19] wl[402] vdd gnd cell_6t
Xbit_r403_c19 bl[19] br[19] wl[403] vdd gnd cell_6t
Xbit_r404_c19 bl[19] br[19] wl[404] vdd gnd cell_6t
Xbit_r405_c19 bl[19] br[19] wl[405] vdd gnd cell_6t
Xbit_r406_c19 bl[19] br[19] wl[406] vdd gnd cell_6t
Xbit_r407_c19 bl[19] br[19] wl[407] vdd gnd cell_6t
Xbit_r408_c19 bl[19] br[19] wl[408] vdd gnd cell_6t
Xbit_r409_c19 bl[19] br[19] wl[409] vdd gnd cell_6t
Xbit_r410_c19 bl[19] br[19] wl[410] vdd gnd cell_6t
Xbit_r411_c19 bl[19] br[19] wl[411] vdd gnd cell_6t
Xbit_r412_c19 bl[19] br[19] wl[412] vdd gnd cell_6t
Xbit_r413_c19 bl[19] br[19] wl[413] vdd gnd cell_6t
Xbit_r414_c19 bl[19] br[19] wl[414] vdd gnd cell_6t
Xbit_r415_c19 bl[19] br[19] wl[415] vdd gnd cell_6t
Xbit_r416_c19 bl[19] br[19] wl[416] vdd gnd cell_6t
Xbit_r417_c19 bl[19] br[19] wl[417] vdd gnd cell_6t
Xbit_r418_c19 bl[19] br[19] wl[418] vdd gnd cell_6t
Xbit_r419_c19 bl[19] br[19] wl[419] vdd gnd cell_6t
Xbit_r420_c19 bl[19] br[19] wl[420] vdd gnd cell_6t
Xbit_r421_c19 bl[19] br[19] wl[421] vdd gnd cell_6t
Xbit_r422_c19 bl[19] br[19] wl[422] vdd gnd cell_6t
Xbit_r423_c19 bl[19] br[19] wl[423] vdd gnd cell_6t
Xbit_r424_c19 bl[19] br[19] wl[424] vdd gnd cell_6t
Xbit_r425_c19 bl[19] br[19] wl[425] vdd gnd cell_6t
Xbit_r426_c19 bl[19] br[19] wl[426] vdd gnd cell_6t
Xbit_r427_c19 bl[19] br[19] wl[427] vdd gnd cell_6t
Xbit_r428_c19 bl[19] br[19] wl[428] vdd gnd cell_6t
Xbit_r429_c19 bl[19] br[19] wl[429] vdd gnd cell_6t
Xbit_r430_c19 bl[19] br[19] wl[430] vdd gnd cell_6t
Xbit_r431_c19 bl[19] br[19] wl[431] vdd gnd cell_6t
Xbit_r432_c19 bl[19] br[19] wl[432] vdd gnd cell_6t
Xbit_r433_c19 bl[19] br[19] wl[433] vdd gnd cell_6t
Xbit_r434_c19 bl[19] br[19] wl[434] vdd gnd cell_6t
Xbit_r435_c19 bl[19] br[19] wl[435] vdd gnd cell_6t
Xbit_r436_c19 bl[19] br[19] wl[436] vdd gnd cell_6t
Xbit_r437_c19 bl[19] br[19] wl[437] vdd gnd cell_6t
Xbit_r438_c19 bl[19] br[19] wl[438] vdd gnd cell_6t
Xbit_r439_c19 bl[19] br[19] wl[439] vdd gnd cell_6t
Xbit_r440_c19 bl[19] br[19] wl[440] vdd gnd cell_6t
Xbit_r441_c19 bl[19] br[19] wl[441] vdd gnd cell_6t
Xbit_r442_c19 bl[19] br[19] wl[442] vdd gnd cell_6t
Xbit_r443_c19 bl[19] br[19] wl[443] vdd gnd cell_6t
Xbit_r444_c19 bl[19] br[19] wl[444] vdd gnd cell_6t
Xbit_r445_c19 bl[19] br[19] wl[445] vdd gnd cell_6t
Xbit_r446_c19 bl[19] br[19] wl[446] vdd gnd cell_6t
Xbit_r447_c19 bl[19] br[19] wl[447] vdd gnd cell_6t
Xbit_r448_c19 bl[19] br[19] wl[448] vdd gnd cell_6t
Xbit_r449_c19 bl[19] br[19] wl[449] vdd gnd cell_6t
Xbit_r450_c19 bl[19] br[19] wl[450] vdd gnd cell_6t
Xbit_r451_c19 bl[19] br[19] wl[451] vdd gnd cell_6t
Xbit_r452_c19 bl[19] br[19] wl[452] vdd gnd cell_6t
Xbit_r453_c19 bl[19] br[19] wl[453] vdd gnd cell_6t
Xbit_r454_c19 bl[19] br[19] wl[454] vdd gnd cell_6t
Xbit_r455_c19 bl[19] br[19] wl[455] vdd gnd cell_6t
Xbit_r456_c19 bl[19] br[19] wl[456] vdd gnd cell_6t
Xbit_r457_c19 bl[19] br[19] wl[457] vdd gnd cell_6t
Xbit_r458_c19 bl[19] br[19] wl[458] vdd gnd cell_6t
Xbit_r459_c19 bl[19] br[19] wl[459] vdd gnd cell_6t
Xbit_r460_c19 bl[19] br[19] wl[460] vdd gnd cell_6t
Xbit_r461_c19 bl[19] br[19] wl[461] vdd gnd cell_6t
Xbit_r462_c19 bl[19] br[19] wl[462] vdd gnd cell_6t
Xbit_r463_c19 bl[19] br[19] wl[463] vdd gnd cell_6t
Xbit_r464_c19 bl[19] br[19] wl[464] vdd gnd cell_6t
Xbit_r465_c19 bl[19] br[19] wl[465] vdd gnd cell_6t
Xbit_r466_c19 bl[19] br[19] wl[466] vdd gnd cell_6t
Xbit_r467_c19 bl[19] br[19] wl[467] vdd gnd cell_6t
Xbit_r468_c19 bl[19] br[19] wl[468] vdd gnd cell_6t
Xbit_r469_c19 bl[19] br[19] wl[469] vdd gnd cell_6t
Xbit_r470_c19 bl[19] br[19] wl[470] vdd gnd cell_6t
Xbit_r471_c19 bl[19] br[19] wl[471] vdd gnd cell_6t
Xbit_r472_c19 bl[19] br[19] wl[472] vdd gnd cell_6t
Xbit_r473_c19 bl[19] br[19] wl[473] vdd gnd cell_6t
Xbit_r474_c19 bl[19] br[19] wl[474] vdd gnd cell_6t
Xbit_r475_c19 bl[19] br[19] wl[475] vdd gnd cell_6t
Xbit_r476_c19 bl[19] br[19] wl[476] vdd gnd cell_6t
Xbit_r477_c19 bl[19] br[19] wl[477] vdd gnd cell_6t
Xbit_r478_c19 bl[19] br[19] wl[478] vdd gnd cell_6t
Xbit_r479_c19 bl[19] br[19] wl[479] vdd gnd cell_6t
Xbit_r480_c19 bl[19] br[19] wl[480] vdd gnd cell_6t
Xbit_r481_c19 bl[19] br[19] wl[481] vdd gnd cell_6t
Xbit_r482_c19 bl[19] br[19] wl[482] vdd gnd cell_6t
Xbit_r483_c19 bl[19] br[19] wl[483] vdd gnd cell_6t
Xbit_r484_c19 bl[19] br[19] wl[484] vdd gnd cell_6t
Xbit_r485_c19 bl[19] br[19] wl[485] vdd gnd cell_6t
Xbit_r486_c19 bl[19] br[19] wl[486] vdd gnd cell_6t
Xbit_r487_c19 bl[19] br[19] wl[487] vdd gnd cell_6t
Xbit_r488_c19 bl[19] br[19] wl[488] vdd gnd cell_6t
Xbit_r489_c19 bl[19] br[19] wl[489] vdd gnd cell_6t
Xbit_r490_c19 bl[19] br[19] wl[490] vdd gnd cell_6t
Xbit_r491_c19 bl[19] br[19] wl[491] vdd gnd cell_6t
Xbit_r492_c19 bl[19] br[19] wl[492] vdd gnd cell_6t
Xbit_r493_c19 bl[19] br[19] wl[493] vdd gnd cell_6t
Xbit_r494_c19 bl[19] br[19] wl[494] vdd gnd cell_6t
Xbit_r495_c19 bl[19] br[19] wl[495] vdd gnd cell_6t
Xbit_r496_c19 bl[19] br[19] wl[496] vdd gnd cell_6t
Xbit_r497_c19 bl[19] br[19] wl[497] vdd gnd cell_6t
Xbit_r498_c19 bl[19] br[19] wl[498] vdd gnd cell_6t
Xbit_r499_c19 bl[19] br[19] wl[499] vdd gnd cell_6t
Xbit_r500_c19 bl[19] br[19] wl[500] vdd gnd cell_6t
Xbit_r501_c19 bl[19] br[19] wl[501] vdd gnd cell_6t
Xbit_r502_c19 bl[19] br[19] wl[502] vdd gnd cell_6t
Xbit_r503_c19 bl[19] br[19] wl[503] vdd gnd cell_6t
Xbit_r504_c19 bl[19] br[19] wl[504] vdd gnd cell_6t
Xbit_r505_c19 bl[19] br[19] wl[505] vdd gnd cell_6t
Xbit_r506_c19 bl[19] br[19] wl[506] vdd gnd cell_6t
Xbit_r507_c19 bl[19] br[19] wl[507] vdd gnd cell_6t
Xbit_r508_c19 bl[19] br[19] wl[508] vdd gnd cell_6t
Xbit_r509_c19 bl[19] br[19] wl[509] vdd gnd cell_6t
Xbit_r510_c19 bl[19] br[19] wl[510] vdd gnd cell_6t
Xbit_r511_c19 bl[19] br[19] wl[511] vdd gnd cell_6t
Xbit_r0_c20 bl[20] br[20] wl[0] vdd gnd cell_6t
Xbit_r1_c20 bl[20] br[20] wl[1] vdd gnd cell_6t
Xbit_r2_c20 bl[20] br[20] wl[2] vdd gnd cell_6t
Xbit_r3_c20 bl[20] br[20] wl[3] vdd gnd cell_6t
Xbit_r4_c20 bl[20] br[20] wl[4] vdd gnd cell_6t
Xbit_r5_c20 bl[20] br[20] wl[5] vdd gnd cell_6t
Xbit_r6_c20 bl[20] br[20] wl[6] vdd gnd cell_6t
Xbit_r7_c20 bl[20] br[20] wl[7] vdd gnd cell_6t
Xbit_r8_c20 bl[20] br[20] wl[8] vdd gnd cell_6t
Xbit_r9_c20 bl[20] br[20] wl[9] vdd gnd cell_6t
Xbit_r10_c20 bl[20] br[20] wl[10] vdd gnd cell_6t
Xbit_r11_c20 bl[20] br[20] wl[11] vdd gnd cell_6t
Xbit_r12_c20 bl[20] br[20] wl[12] vdd gnd cell_6t
Xbit_r13_c20 bl[20] br[20] wl[13] vdd gnd cell_6t
Xbit_r14_c20 bl[20] br[20] wl[14] vdd gnd cell_6t
Xbit_r15_c20 bl[20] br[20] wl[15] vdd gnd cell_6t
Xbit_r16_c20 bl[20] br[20] wl[16] vdd gnd cell_6t
Xbit_r17_c20 bl[20] br[20] wl[17] vdd gnd cell_6t
Xbit_r18_c20 bl[20] br[20] wl[18] vdd gnd cell_6t
Xbit_r19_c20 bl[20] br[20] wl[19] vdd gnd cell_6t
Xbit_r20_c20 bl[20] br[20] wl[20] vdd gnd cell_6t
Xbit_r21_c20 bl[20] br[20] wl[21] vdd gnd cell_6t
Xbit_r22_c20 bl[20] br[20] wl[22] vdd gnd cell_6t
Xbit_r23_c20 bl[20] br[20] wl[23] vdd gnd cell_6t
Xbit_r24_c20 bl[20] br[20] wl[24] vdd gnd cell_6t
Xbit_r25_c20 bl[20] br[20] wl[25] vdd gnd cell_6t
Xbit_r26_c20 bl[20] br[20] wl[26] vdd gnd cell_6t
Xbit_r27_c20 bl[20] br[20] wl[27] vdd gnd cell_6t
Xbit_r28_c20 bl[20] br[20] wl[28] vdd gnd cell_6t
Xbit_r29_c20 bl[20] br[20] wl[29] vdd gnd cell_6t
Xbit_r30_c20 bl[20] br[20] wl[30] vdd gnd cell_6t
Xbit_r31_c20 bl[20] br[20] wl[31] vdd gnd cell_6t
Xbit_r32_c20 bl[20] br[20] wl[32] vdd gnd cell_6t
Xbit_r33_c20 bl[20] br[20] wl[33] vdd gnd cell_6t
Xbit_r34_c20 bl[20] br[20] wl[34] vdd gnd cell_6t
Xbit_r35_c20 bl[20] br[20] wl[35] vdd gnd cell_6t
Xbit_r36_c20 bl[20] br[20] wl[36] vdd gnd cell_6t
Xbit_r37_c20 bl[20] br[20] wl[37] vdd gnd cell_6t
Xbit_r38_c20 bl[20] br[20] wl[38] vdd gnd cell_6t
Xbit_r39_c20 bl[20] br[20] wl[39] vdd gnd cell_6t
Xbit_r40_c20 bl[20] br[20] wl[40] vdd gnd cell_6t
Xbit_r41_c20 bl[20] br[20] wl[41] vdd gnd cell_6t
Xbit_r42_c20 bl[20] br[20] wl[42] vdd gnd cell_6t
Xbit_r43_c20 bl[20] br[20] wl[43] vdd gnd cell_6t
Xbit_r44_c20 bl[20] br[20] wl[44] vdd gnd cell_6t
Xbit_r45_c20 bl[20] br[20] wl[45] vdd gnd cell_6t
Xbit_r46_c20 bl[20] br[20] wl[46] vdd gnd cell_6t
Xbit_r47_c20 bl[20] br[20] wl[47] vdd gnd cell_6t
Xbit_r48_c20 bl[20] br[20] wl[48] vdd gnd cell_6t
Xbit_r49_c20 bl[20] br[20] wl[49] vdd gnd cell_6t
Xbit_r50_c20 bl[20] br[20] wl[50] vdd gnd cell_6t
Xbit_r51_c20 bl[20] br[20] wl[51] vdd gnd cell_6t
Xbit_r52_c20 bl[20] br[20] wl[52] vdd gnd cell_6t
Xbit_r53_c20 bl[20] br[20] wl[53] vdd gnd cell_6t
Xbit_r54_c20 bl[20] br[20] wl[54] vdd gnd cell_6t
Xbit_r55_c20 bl[20] br[20] wl[55] vdd gnd cell_6t
Xbit_r56_c20 bl[20] br[20] wl[56] vdd gnd cell_6t
Xbit_r57_c20 bl[20] br[20] wl[57] vdd gnd cell_6t
Xbit_r58_c20 bl[20] br[20] wl[58] vdd gnd cell_6t
Xbit_r59_c20 bl[20] br[20] wl[59] vdd gnd cell_6t
Xbit_r60_c20 bl[20] br[20] wl[60] vdd gnd cell_6t
Xbit_r61_c20 bl[20] br[20] wl[61] vdd gnd cell_6t
Xbit_r62_c20 bl[20] br[20] wl[62] vdd gnd cell_6t
Xbit_r63_c20 bl[20] br[20] wl[63] vdd gnd cell_6t
Xbit_r64_c20 bl[20] br[20] wl[64] vdd gnd cell_6t
Xbit_r65_c20 bl[20] br[20] wl[65] vdd gnd cell_6t
Xbit_r66_c20 bl[20] br[20] wl[66] vdd gnd cell_6t
Xbit_r67_c20 bl[20] br[20] wl[67] vdd gnd cell_6t
Xbit_r68_c20 bl[20] br[20] wl[68] vdd gnd cell_6t
Xbit_r69_c20 bl[20] br[20] wl[69] vdd gnd cell_6t
Xbit_r70_c20 bl[20] br[20] wl[70] vdd gnd cell_6t
Xbit_r71_c20 bl[20] br[20] wl[71] vdd gnd cell_6t
Xbit_r72_c20 bl[20] br[20] wl[72] vdd gnd cell_6t
Xbit_r73_c20 bl[20] br[20] wl[73] vdd gnd cell_6t
Xbit_r74_c20 bl[20] br[20] wl[74] vdd gnd cell_6t
Xbit_r75_c20 bl[20] br[20] wl[75] vdd gnd cell_6t
Xbit_r76_c20 bl[20] br[20] wl[76] vdd gnd cell_6t
Xbit_r77_c20 bl[20] br[20] wl[77] vdd gnd cell_6t
Xbit_r78_c20 bl[20] br[20] wl[78] vdd gnd cell_6t
Xbit_r79_c20 bl[20] br[20] wl[79] vdd gnd cell_6t
Xbit_r80_c20 bl[20] br[20] wl[80] vdd gnd cell_6t
Xbit_r81_c20 bl[20] br[20] wl[81] vdd gnd cell_6t
Xbit_r82_c20 bl[20] br[20] wl[82] vdd gnd cell_6t
Xbit_r83_c20 bl[20] br[20] wl[83] vdd gnd cell_6t
Xbit_r84_c20 bl[20] br[20] wl[84] vdd gnd cell_6t
Xbit_r85_c20 bl[20] br[20] wl[85] vdd gnd cell_6t
Xbit_r86_c20 bl[20] br[20] wl[86] vdd gnd cell_6t
Xbit_r87_c20 bl[20] br[20] wl[87] vdd gnd cell_6t
Xbit_r88_c20 bl[20] br[20] wl[88] vdd gnd cell_6t
Xbit_r89_c20 bl[20] br[20] wl[89] vdd gnd cell_6t
Xbit_r90_c20 bl[20] br[20] wl[90] vdd gnd cell_6t
Xbit_r91_c20 bl[20] br[20] wl[91] vdd gnd cell_6t
Xbit_r92_c20 bl[20] br[20] wl[92] vdd gnd cell_6t
Xbit_r93_c20 bl[20] br[20] wl[93] vdd gnd cell_6t
Xbit_r94_c20 bl[20] br[20] wl[94] vdd gnd cell_6t
Xbit_r95_c20 bl[20] br[20] wl[95] vdd gnd cell_6t
Xbit_r96_c20 bl[20] br[20] wl[96] vdd gnd cell_6t
Xbit_r97_c20 bl[20] br[20] wl[97] vdd gnd cell_6t
Xbit_r98_c20 bl[20] br[20] wl[98] vdd gnd cell_6t
Xbit_r99_c20 bl[20] br[20] wl[99] vdd gnd cell_6t
Xbit_r100_c20 bl[20] br[20] wl[100] vdd gnd cell_6t
Xbit_r101_c20 bl[20] br[20] wl[101] vdd gnd cell_6t
Xbit_r102_c20 bl[20] br[20] wl[102] vdd gnd cell_6t
Xbit_r103_c20 bl[20] br[20] wl[103] vdd gnd cell_6t
Xbit_r104_c20 bl[20] br[20] wl[104] vdd gnd cell_6t
Xbit_r105_c20 bl[20] br[20] wl[105] vdd gnd cell_6t
Xbit_r106_c20 bl[20] br[20] wl[106] vdd gnd cell_6t
Xbit_r107_c20 bl[20] br[20] wl[107] vdd gnd cell_6t
Xbit_r108_c20 bl[20] br[20] wl[108] vdd gnd cell_6t
Xbit_r109_c20 bl[20] br[20] wl[109] vdd gnd cell_6t
Xbit_r110_c20 bl[20] br[20] wl[110] vdd gnd cell_6t
Xbit_r111_c20 bl[20] br[20] wl[111] vdd gnd cell_6t
Xbit_r112_c20 bl[20] br[20] wl[112] vdd gnd cell_6t
Xbit_r113_c20 bl[20] br[20] wl[113] vdd gnd cell_6t
Xbit_r114_c20 bl[20] br[20] wl[114] vdd gnd cell_6t
Xbit_r115_c20 bl[20] br[20] wl[115] vdd gnd cell_6t
Xbit_r116_c20 bl[20] br[20] wl[116] vdd gnd cell_6t
Xbit_r117_c20 bl[20] br[20] wl[117] vdd gnd cell_6t
Xbit_r118_c20 bl[20] br[20] wl[118] vdd gnd cell_6t
Xbit_r119_c20 bl[20] br[20] wl[119] vdd gnd cell_6t
Xbit_r120_c20 bl[20] br[20] wl[120] vdd gnd cell_6t
Xbit_r121_c20 bl[20] br[20] wl[121] vdd gnd cell_6t
Xbit_r122_c20 bl[20] br[20] wl[122] vdd gnd cell_6t
Xbit_r123_c20 bl[20] br[20] wl[123] vdd gnd cell_6t
Xbit_r124_c20 bl[20] br[20] wl[124] vdd gnd cell_6t
Xbit_r125_c20 bl[20] br[20] wl[125] vdd gnd cell_6t
Xbit_r126_c20 bl[20] br[20] wl[126] vdd gnd cell_6t
Xbit_r127_c20 bl[20] br[20] wl[127] vdd gnd cell_6t
Xbit_r128_c20 bl[20] br[20] wl[128] vdd gnd cell_6t
Xbit_r129_c20 bl[20] br[20] wl[129] vdd gnd cell_6t
Xbit_r130_c20 bl[20] br[20] wl[130] vdd gnd cell_6t
Xbit_r131_c20 bl[20] br[20] wl[131] vdd gnd cell_6t
Xbit_r132_c20 bl[20] br[20] wl[132] vdd gnd cell_6t
Xbit_r133_c20 bl[20] br[20] wl[133] vdd gnd cell_6t
Xbit_r134_c20 bl[20] br[20] wl[134] vdd gnd cell_6t
Xbit_r135_c20 bl[20] br[20] wl[135] vdd gnd cell_6t
Xbit_r136_c20 bl[20] br[20] wl[136] vdd gnd cell_6t
Xbit_r137_c20 bl[20] br[20] wl[137] vdd gnd cell_6t
Xbit_r138_c20 bl[20] br[20] wl[138] vdd gnd cell_6t
Xbit_r139_c20 bl[20] br[20] wl[139] vdd gnd cell_6t
Xbit_r140_c20 bl[20] br[20] wl[140] vdd gnd cell_6t
Xbit_r141_c20 bl[20] br[20] wl[141] vdd gnd cell_6t
Xbit_r142_c20 bl[20] br[20] wl[142] vdd gnd cell_6t
Xbit_r143_c20 bl[20] br[20] wl[143] vdd gnd cell_6t
Xbit_r144_c20 bl[20] br[20] wl[144] vdd gnd cell_6t
Xbit_r145_c20 bl[20] br[20] wl[145] vdd gnd cell_6t
Xbit_r146_c20 bl[20] br[20] wl[146] vdd gnd cell_6t
Xbit_r147_c20 bl[20] br[20] wl[147] vdd gnd cell_6t
Xbit_r148_c20 bl[20] br[20] wl[148] vdd gnd cell_6t
Xbit_r149_c20 bl[20] br[20] wl[149] vdd gnd cell_6t
Xbit_r150_c20 bl[20] br[20] wl[150] vdd gnd cell_6t
Xbit_r151_c20 bl[20] br[20] wl[151] vdd gnd cell_6t
Xbit_r152_c20 bl[20] br[20] wl[152] vdd gnd cell_6t
Xbit_r153_c20 bl[20] br[20] wl[153] vdd gnd cell_6t
Xbit_r154_c20 bl[20] br[20] wl[154] vdd gnd cell_6t
Xbit_r155_c20 bl[20] br[20] wl[155] vdd gnd cell_6t
Xbit_r156_c20 bl[20] br[20] wl[156] vdd gnd cell_6t
Xbit_r157_c20 bl[20] br[20] wl[157] vdd gnd cell_6t
Xbit_r158_c20 bl[20] br[20] wl[158] vdd gnd cell_6t
Xbit_r159_c20 bl[20] br[20] wl[159] vdd gnd cell_6t
Xbit_r160_c20 bl[20] br[20] wl[160] vdd gnd cell_6t
Xbit_r161_c20 bl[20] br[20] wl[161] vdd gnd cell_6t
Xbit_r162_c20 bl[20] br[20] wl[162] vdd gnd cell_6t
Xbit_r163_c20 bl[20] br[20] wl[163] vdd gnd cell_6t
Xbit_r164_c20 bl[20] br[20] wl[164] vdd gnd cell_6t
Xbit_r165_c20 bl[20] br[20] wl[165] vdd gnd cell_6t
Xbit_r166_c20 bl[20] br[20] wl[166] vdd gnd cell_6t
Xbit_r167_c20 bl[20] br[20] wl[167] vdd gnd cell_6t
Xbit_r168_c20 bl[20] br[20] wl[168] vdd gnd cell_6t
Xbit_r169_c20 bl[20] br[20] wl[169] vdd gnd cell_6t
Xbit_r170_c20 bl[20] br[20] wl[170] vdd gnd cell_6t
Xbit_r171_c20 bl[20] br[20] wl[171] vdd gnd cell_6t
Xbit_r172_c20 bl[20] br[20] wl[172] vdd gnd cell_6t
Xbit_r173_c20 bl[20] br[20] wl[173] vdd gnd cell_6t
Xbit_r174_c20 bl[20] br[20] wl[174] vdd gnd cell_6t
Xbit_r175_c20 bl[20] br[20] wl[175] vdd gnd cell_6t
Xbit_r176_c20 bl[20] br[20] wl[176] vdd gnd cell_6t
Xbit_r177_c20 bl[20] br[20] wl[177] vdd gnd cell_6t
Xbit_r178_c20 bl[20] br[20] wl[178] vdd gnd cell_6t
Xbit_r179_c20 bl[20] br[20] wl[179] vdd gnd cell_6t
Xbit_r180_c20 bl[20] br[20] wl[180] vdd gnd cell_6t
Xbit_r181_c20 bl[20] br[20] wl[181] vdd gnd cell_6t
Xbit_r182_c20 bl[20] br[20] wl[182] vdd gnd cell_6t
Xbit_r183_c20 bl[20] br[20] wl[183] vdd gnd cell_6t
Xbit_r184_c20 bl[20] br[20] wl[184] vdd gnd cell_6t
Xbit_r185_c20 bl[20] br[20] wl[185] vdd gnd cell_6t
Xbit_r186_c20 bl[20] br[20] wl[186] vdd gnd cell_6t
Xbit_r187_c20 bl[20] br[20] wl[187] vdd gnd cell_6t
Xbit_r188_c20 bl[20] br[20] wl[188] vdd gnd cell_6t
Xbit_r189_c20 bl[20] br[20] wl[189] vdd gnd cell_6t
Xbit_r190_c20 bl[20] br[20] wl[190] vdd gnd cell_6t
Xbit_r191_c20 bl[20] br[20] wl[191] vdd gnd cell_6t
Xbit_r192_c20 bl[20] br[20] wl[192] vdd gnd cell_6t
Xbit_r193_c20 bl[20] br[20] wl[193] vdd gnd cell_6t
Xbit_r194_c20 bl[20] br[20] wl[194] vdd gnd cell_6t
Xbit_r195_c20 bl[20] br[20] wl[195] vdd gnd cell_6t
Xbit_r196_c20 bl[20] br[20] wl[196] vdd gnd cell_6t
Xbit_r197_c20 bl[20] br[20] wl[197] vdd gnd cell_6t
Xbit_r198_c20 bl[20] br[20] wl[198] vdd gnd cell_6t
Xbit_r199_c20 bl[20] br[20] wl[199] vdd gnd cell_6t
Xbit_r200_c20 bl[20] br[20] wl[200] vdd gnd cell_6t
Xbit_r201_c20 bl[20] br[20] wl[201] vdd gnd cell_6t
Xbit_r202_c20 bl[20] br[20] wl[202] vdd gnd cell_6t
Xbit_r203_c20 bl[20] br[20] wl[203] vdd gnd cell_6t
Xbit_r204_c20 bl[20] br[20] wl[204] vdd gnd cell_6t
Xbit_r205_c20 bl[20] br[20] wl[205] vdd gnd cell_6t
Xbit_r206_c20 bl[20] br[20] wl[206] vdd gnd cell_6t
Xbit_r207_c20 bl[20] br[20] wl[207] vdd gnd cell_6t
Xbit_r208_c20 bl[20] br[20] wl[208] vdd gnd cell_6t
Xbit_r209_c20 bl[20] br[20] wl[209] vdd gnd cell_6t
Xbit_r210_c20 bl[20] br[20] wl[210] vdd gnd cell_6t
Xbit_r211_c20 bl[20] br[20] wl[211] vdd gnd cell_6t
Xbit_r212_c20 bl[20] br[20] wl[212] vdd gnd cell_6t
Xbit_r213_c20 bl[20] br[20] wl[213] vdd gnd cell_6t
Xbit_r214_c20 bl[20] br[20] wl[214] vdd gnd cell_6t
Xbit_r215_c20 bl[20] br[20] wl[215] vdd gnd cell_6t
Xbit_r216_c20 bl[20] br[20] wl[216] vdd gnd cell_6t
Xbit_r217_c20 bl[20] br[20] wl[217] vdd gnd cell_6t
Xbit_r218_c20 bl[20] br[20] wl[218] vdd gnd cell_6t
Xbit_r219_c20 bl[20] br[20] wl[219] vdd gnd cell_6t
Xbit_r220_c20 bl[20] br[20] wl[220] vdd gnd cell_6t
Xbit_r221_c20 bl[20] br[20] wl[221] vdd gnd cell_6t
Xbit_r222_c20 bl[20] br[20] wl[222] vdd gnd cell_6t
Xbit_r223_c20 bl[20] br[20] wl[223] vdd gnd cell_6t
Xbit_r224_c20 bl[20] br[20] wl[224] vdd gnd cell_6t
Xbit_r225_c20 bl[20] br[20] wl[225] vdd gnd cell_6t
Xbit_r226_c20 bl[20] br[20] wl[226] vdd gnd cell_6t
Xbit_r227_c20 bl[20] br[20] wl[227] vdd gnd cell_6t
Xbit_r228_c20 bl[20] br[20] wl[228] vdd gnd cell_6t
Xbit_r229_c20 bl[20] br[20] wl[229] vdd gnd cell_6t
Xbit_r230_c20 bl[20] br[20] wl[230] vdd gnd cell_6t
Xbit_r231_c20 bl[20] br[20] wl[231] vdd gnd cell_6t
Xbit_r232_c20 bl[20] br[20] wl[232] vdd gnd cell_6t
Xbit_r233_c20 bl[20] br[20] wl[233] vdd gnd cell_6t
Xbit_r234_c20 bl[20] br[20] wl[234] vdd gnd cell_6t
Xbit_r235_c20 bl[20] br[20] wl[235] vdd gnd cell_6t
Xbit_r236_c20 bl[20] br[20] wl[236] vdd gnd cell_6t
Xbit_r237_c20 bl[20] br[20] wl[237] vdd gnd cell_6t
Xbit_r238_c20 bl[20] br[20] wl[238] vdd gnd cell_6t
Xbit_r239_c20 bl[20] br[20] wl[239] vdd gnd cell_6t
Xbit_r240_c20 bl[20] br[20] wl[240] vdd gnd cell_6t
Xbit_r241_c20 bl[20] br[20] wl[241] vdd gnd cell_6t
Xbit_r242_c20 bl[20] br[20] wl[242] vdd gnd cell_6t
Xbit_r243_c20 bl[20] br[20] wl[243] vdd gnd cell_6t
Xbit_r244_c20 bl[20] br[20] wl[244] vdd gnd cell_6t
Xbit_r245_c20 bl[20] br[20] wl[245] vdd gnd cell_6t
Xbit_r246_c20 bl[20] br[20] wl[246] vdd gnd cell_6t
Xbit_r247_c20 bl[20] br[20] wl[247] vdd gnd cell_6t
Xbit_r248_c20 bl[20] br[20] wl[248] vdd gnd cell_6t
Xbit_r249_c20 bl[20] br[20] wl[249] vdd gnd cell_6t
Xbit_r250_c20 bl[20] br[20] wl[250] vdd gnd cell_6t
Xbit_r251_c20 bl[20] br[20] wl[251] vdd gnd cell_6t
Xbit_r252_c20 bl[20] br[20] wl[252] vdd gnd cell_6t
Xbit_r253_c20 bl[20] br[20] wl[253] vdd gnd cell_6t
Xbit_r254_c20 bl[20] br[20] wl[254] vdd gnd cell_6t
Xbit_r255_c20 bl[20] br[20] wl[255] vdd gnd cell_6t
Xbit_r256_c20 bl[20] br[20] wl[256] vdd gnd cell_6t
Xbit_r257_c20 bl[20] br[20] wl[257] vdd gnd cell_6t
Xbit_r258_c20 bl[20] br[20] wl[258] vdd gnd cell_6t
Xbit_r259_c20 bl[20] br[20] wl[259] vdd gnd cell_6t
Xbit_r260_c20 bl[20] br[20] wl[260] vdd gnd cell_6t
Xbit_r261_c20 bl[20] br[20] wl[261] vdd gnd cell_6t
Xbit_r262_c20 bl[20] br[20] wl[262] vdd gnd cell_6t
Xbit_r263_c20 bl[20] br[20] wl[263] vdd gnd cell_6t
Xbit_r264_c20 bl[20] br[20] wl[264] vdd gnd cell_6t
Xbit_r265_c20 bl[20] br[20] wl[265] vdd gnd cell_6t
Xbit_r266_c20 bl[20] br[20] wl[266] vdd gnd cell_6t
Xbit_r267_c20 bl[20] br[20] wl[267] vdd gnd cell_6t
Xbit_r268_c20 bl[20] br[20] wl[268] vdd gnd cell_6t
Xbit_r269_c20 bl[20] br[20] wl[269] vdd gnd cell_6t
Xbit_r270_c20 bl[20] br[20] wl[270] vdd gnd cell_6t
Xbit_r271_c20 bl[20] br[20] wl[271] vdd gnd cell_6t
Xbit_r272_c20 bl[20] br[20] wl[272] vdd gnd cell_6t
Xbit_r273_c20 bl[20] br[20] wl[273] vdd gnd cell_6t
Xbit_r274_c20 bl[20] br[20] wl[274] vdd gnd cell_6t
Xbit_r275_c20 bl[20] br[20] wl[275] vdd gnd cell_6t
Xbit_r276_c20 bl[20] br[20] wl[276] vdd gnd cell_6t
Xbit_r277_c20 bl[20] br[20] wl[277] vdd gnd cell_6t
Xbit_r278_c20 bl[20] br[20] wl[278] vdd gnd cell_6t
Xbit_r279_c20 bl[20] br[20] wl[279] vdd gnd cell_6t
Xbit_r280_c20 bl[20] br[20] wl[280] vdd gnd cell_6t
Xbit_r281_c20 bl[20] br[20] wl[281] vdd gnd cell_6t
Xbit_r282_c20 bl[20] br[20] wl[282] vdd gnd cell_6t
Xbit_r283_c20 bl[20] br[20] wl[283] vdd gnd cell_6t
Xbit_r284_c20 bl[20] br[20] wl[284] vdd gnd cell_6t
Xbit_r285_c20 bl[20] br[20] wl[285] vdd gnd cell_6t
Xbit_r286_c20 bl[20] br[20] wl[286] vdd gnd cell_6t
Xbit_r287_c20 bl[20] br[20] wl[287] vdd gnd cell_6t
Xbit_r288_c20 bl[20] br[20] wl[288] vdd gnd cell_6t
Xbit_r289_c20 bl[20] br[20] wl[289] vdd gnd cell_6t
Xbit_r290_c20 bl[20] br[20] wl[290] vdd gnd cell_6t
Xbit_r291_c20 bl[20] br[20] wl[291] vdd gnd cell_6t
Xbit_r292_c20 bl[20] br[20] wl[292] vdd gnd cell_6t
Xbit_r293_c20 bl[20] br[20] wl[293] vdd gnd cell_6t
Xbit_r294_c20 bl[20] br[20] wl[294] vdd gnd cell_6t
Xbit_r295_c20 bl[20] br[20] wl[295] vdd gnd cell_6t
Xbit_r296_c20 bl[20] br[20] wl[296] vdd gnd cell_6t
Xbit_r297_c20 bl[20] br[20] wl[297] vdd gnd cell_6t
Xbit_r298_c20 bl[20] br[20] wl[298] vdd gnd cell_6t
Xbit_r299_c20 bl[20] br[20] wl[299] vdd gnd cell_6t
Xbit_r300_c20 bl[20] br[20] wl[300] vdd gnd cell_6t
Xbit_r301_c20 bl[20] br[20] wl[301] vdd gnd cell_6t
Xbit_r302_c20 bl[20] br[20] wl[302] vdd gnd cell_6t
Xbit_r303_c20 bl[20] br[20] wl[303] vdd gnd cell_6t
Xbit_r304_c20 bl[20] br[20] wl[304] vdd gnd cell_6t
Xbit_r305_c20 bl[20] br[20] wl[305] vdd gnd cell_6t
Xbit_r306_c20 bl[20] br[20] wl[306] vdd gnd cell_6t
Xbit_r307_c20 bl[20] br[20] wl[307] vdd gnd cell_6t
Xbit_r308_c20 bl[20] br[20] wl[308] vdd gnd cell_6t
Xbit_r309_c20 bl[20] br[20] wl[309] vdd gnd cell_6t
Xbit_r310_c20 bl[20] br[20] wl[310] vdd gnd cell_6t
Xbit_r311_c20 bl[20] br[20] wl[311] vdd gnd cell_6t
Xbit_r312_c20 bl[20] br[20] wl[312] vdd gnd cell_6t
Xbit_r313_c20 bl[20] br[20] wl[313] vdd gnd cell_6t
Xbit_r314_c20 bl[20] br[20] wl[314] vdd gnd cell_6t
Xbit_r315_c20 bl[20] br[20] wl[315] vdd gnd cell_6t
Xbit_r316_c20 bl[20] br[20] wl[316] vdd gnd cell_6t
Xbit_r317_c20 bl[20] br[20] wl[317] vdd gnd cell_6t
Xbit_r318_c20 bl[20] br[20] wl[318] vdd gnd cell_6t
Xbit_r319_c20 bl[20] br[20] wl[319] vdd gnd cell_6t
Xbit_r320_c20 bl[20] br[20] wl[320] vdd gnd cell_6t
Xbit_r321_c20 bl[20] br[20] wl[321] vdd gnd cell_6t
Xbit_r322_c20 bl[20] br[20] wl[322] vdd gnd cell_6t
Xbit_r323_c20 bl[20] br[20] wl[323] vdd gnd cell_6t
Xbit_r324_c20 bl[20] br[20] wl[324] vdd gnd cell_6t
Xbit_r325_c20 bl[20] br[20] wl[325] vdd gnd cell_6t
Xbit_r326_c20 bl[20] br[20] wl[326] vdd gnd cell_6t
Xbit_r327_c20 bl[20] br[20] wl[327] vdd gnd cell_6t
Xbit_r328_c20 bl[20] br[20] wl[328] vdd gnd cell_6t
Xbit_r329_c20 bl[20] br[20] wl[329] vdd gnd cell_6t
Xbit_r330_c20 bl[20] br[20] wl[330] vdd gnd cell_6t
Xbit_r331_c20 bl[20] br[20] wl[331] vdd gnd cell_6t
Xbit_r332_c20 bl[20] br[20] wl[332] vdd gnd cell_6t
Xbit_r333_c20 bl[20] br[20] wl[333] vdd gnd cell_6t
Xbit_r334_c20 bl[20] br[20] wl[334] vdd gnd cell_6t
Xbit_r335_c20 bl[20] br[20] wl[335] vdd gnd cell_6t
Xbit_r336_c20 bl[20] br[20] wl[336] vdd gnd cell_6t
Xbit_r337_c20 bl[20] br[20] wl[337] vdd gnd cell_6t
Xbit_r338_c20 bl[20] br[20] wl[338] vdd gnd cell_6t
Xbit_r339_c20 bl[20] br[20] wl[339] vdd gnd cell_6t
Xbit_r340_c20 bl[20] br[20] wl[340] vdd gnd cell_6t
Xbit_r341_c20 bl[20] br[20] wl[341] vdd gnd cell_6t
Xbit_r342_c20 bl[20] br[20] wl[342] vdd gnd cell_6t
Xbit_r343_c20 bl[20] br[20] wl[343] vdd gnd cell_6t
Xbit_r344_c20 bl[20] br[20] wl[344] vdd gnd cell_6t
Xbit_r345_c20 bl[20] br[20] wl[345] vdd gnd cell_6t
Xbit_r346_c20 bl[20] br[20] wl[346] vdd gnd cell_6t
Xbit_r347_c20 bl[20] br[20] wl[347] vdd gnd cell_6t
Xbit_r348_c20 bl[20] br[20] wl[348] vdd gnd cell_6t
Xbit_r349_c20 bl[20] br[20] wl[349] vdd gnd cell_6t
Xbit_r350_c20 bl[20] br[20] wl[350] vdd gnd cell_6t
Xbit_r351_c20 bl[20] br[20] wl[351] vdd gnd cell_6t
Xbit_r352_c20 bl[20] br[20] wl[352] vdd gnd cell_6t
Xbit_r353_c20 bl[20] br[20] wl[353] vdd gnd cell_6t
Xbit_r354_c20 bl[20] br[20] wl[354] vdd gnd cell_6t
Xbit_r355_c20 bl[20] br[20] wl[355] vdd gnd cell_6t
Xbit_r356_c20 bl[20] br[20] wl[356] vdd gnd cell_6t
Xbit_r357_c20 bl[20] br[20] wl[357] vdd gnd cell_6t
Xbit_r358_c20 bl[20] br[20] wl[358] vdd gnd cell_6t
Xbit_r359_c20 bl[20] br[20] wl[359] vdd gnd cell_6t
Xbit_r360_c20 bl[20] br[20] wl[360] vdd gnd cell_6t
Xbit_r361_c20 bl[20] br[20] wl[361] vdd gnd cell_6t
Xbit_r362_c20 bl[20] br[20] wl[362] vdd gnd cell_6t
Xbit_r363_c20 bl[20] br[20] wl[363] vdd gnd cell_6t
Xbit_r364_c20 bl[20] br[20] wl[364] vdd gnd cell_6t
Xbit_r365_c20 bl[20] br[20] wl[365] vdd gnd cell_6t
Xbit_r366_c20 bl[20] br[20] wl[366] vdd gnd cell_6t
Xbit_r367_c20 bl[20] br[20] wl[367] vdd gnd cell_6t
Xbit_r368_c20 bl[20] br[20] wl[368] vdd gnd cell_6t
Xbit_r369_c20 bl[20] br[20] wl[369] vdd gnd cell_6t
Xbit_r370_c20 bl[20] br[20] wl[370] vdd gnd cell_6t
Xbit_r371_c20 bl[20] br[20] wl[371] vdd gnd cell_6t
Xbit_r372_c20 bl[20] br[20] wl[372] vdd gnd cell_6t
Xbit_r373_c20 bl[20] br[20] wl[373] vdd gnd cell_6t
Xbit_r374_c20 bl[20] br[20] wl[374] vdd gnd cell_6t
Xbit_r375_c20 bl[20] br[20] wl[375] vdd gnd cell_6t
Xbit_r376_c20 bl[20] br[20] wl[376] vdd gnd cell_6t
Xbit_r377_c20 bl[20] br[20] wl[377] vdd gnd cell_6t
Xbit_r378_c20 bl[20] br[20] wl[378] vdd gnd cell_6t
Xbit_r379_c20 bl[20] br[20] wl[379] vdd gnd cell_6t
Xbit_r380_c20 bl[20] br[20] wl[380] vdd gnd cell_6t
Xbit_r381_c20 bl[20] br[20] wl[381] vdd gnd cell_6t
Xbit_r382_c20 bl[20] br[20] wl[382] vdd gnd cell_6t
Xbit_r383_c20 bl[20] br[20] wl[383] vdd gnd cell_6t
Xbit_r384_c20 bl[20] br[20] wl[384] vdd gnd cell_6t
Xbit_r385_c20 bl[20] br[20] wl[385] vdd gnd cell_6t
Xbit_r386_c20 bl[20] br[20] wl[386] vdd gnd cell_6t
Xbit_r387_c20 bl[20] br[20] wl[387] vdd gnd cell_6t
Xbit_r388_c20 bl[20] br[20] wl[388] vdd gnd cell_6t
Xbit_r389_c20 bl[20] br[20] wl[389] vdd gnd cell_6t
Xbit_r390_c20 bl[20] br[20] wl[390] vdd gnd cell_6t
Xbit_r391_c20 bl[20] br[20] wl[391] vdd gnd cell_6t
Xbit_r392_c20 bl[20] br[20] wl[392] vdd gnd cell_6t
Xbit_r393_c20 bl[20] br[20] wl[393] vdd gnd cell_6t
Xbit_r394_c20 bl[20] br[20] wl[394] vdd gnd cell_6t
Xbit_r395_c20 bl[20] br[20] wl[395] vdd gnd cell_6t
Xbit_r396_c20 bl[20] br[20] wl[396] vdd gnd cell_6t
Xbit_r397_c20 bl[20] br[20] wl[397] vdd gnd cell_6t
Xbit_r398_c20 bl[20] br[20] wl[398] vdd gnd cell_6t
Xbit_r399_c20 bl[20] br[20] wl[399] vdd gnd cell_6t
Xbit_r400_c20 bl[20] br[20] wl[400] vdd gnd cell_6t
Xbit_r401_c20 bl[20] br[20] wl[401] vdd gnd cell_6t
Xbit_r402_c20 bl[20] br[20] wl[402] vdd gnd cell_6t
Xbit_r403_c20 bl[20] br[20] wl[403] vdd gnd cell_6t
Xbit_r404_c20 bl[20] br[20] wl[404] vdd gnd cell_6t
Xbit_r405_c20 bl[20] br[20] wl[405] vdd gnd cell_6t
Xbit_r406_c20 bl[20] br[20] wl[406] vdd gnd cell_6t
Xbit_r407_c20 bl[20] br[20] wl[407] vdd gnd cell_6t
Xbit_r408_c20 bl[20] br[20] wl[408] vdd gnd cell_6t
Xbit_r409_c20 bl[20] br[20] wl[409] vdd gnd cell_6t
Xbit_r410_c20 bl[20] br[20] wl[410] vdd gnd cell_6t
Xbit_r411_c20 bl[20] br[20] wl[411] vdd gnd cell_6t
Xbit_r412_c20 bl[20] br[20] wl[412] vdd gnd cell_6t
Xbit_r413_c20 bl[20] br[20] wl[413] vdd gnd cell_6t
Xbit_r414_c20 bl[20] br[20] wl[414] vdd gnd cell_6t
Xbit_r415_c20 bl[20] br[20] wl[415] vdd gnd cell_6t
Xbit_r416_c20 bl[20] br[20] wl[416] vdd gnd cell_6t
Xbit_r417_c20 bl[20] br[20] wl[417] vdd gnd cell_6t
Xbit_r418_c20 bl[20] br[20] wl[418] vdd gnd cell_6t
Xbit_r419_c20 bl[20] br[20] wl[419] vdd gnd cell_6t
Xbit_r420_c20 bl[20] br[20] wl[420] vdd gnd cell_6t
Xbit_r421_c20 bl[20] br[20] wl[421] vdd gnd cell_6t
Xbit_r422_c20 bl[20] br[20] wl[422] vdd gnd cell_6t
Xbit_r423_c20 bl[20] br[20] wl[423] vdd gnd cell_6t
Xbit_r424_c20 bl[20] br[20] wl[424] vdd gnd cell_6t
Xbit_r425_c20 bl[20] br[20] wl[425] vdd gnd cell_6t
Xbit_r426_c20 bl[20] br[20] wl[426] vdd gnd cell_6t
Xbit_r427_c20 bl[20] br[20] wl[427] vdd gnd cell_6t
Xbit_r428_c20 bl[20] br[20] wl[428] vdd gnd cell_6t
Xbit_r429_c20 bl[20] br[20] wl[429] vdd gnd cell_6t
Xbit_r430_c20 bl[20] br[20] wl[430] vdd gnd cell_6t
Xbit_r431_c20 bl[20] br[20] wl[431] vdd gnd cell_6t
Xbit_r432_c20 bl[20] br[20] wl[432] vdd gnd cell_6t
Xbit_r433_c20 bl[20] br[20] wl[433] vdd gnd cell_6t
Xbit_r434_c20 bl[20] br[20] wl[434] vdd gnd cell_6t
Xbit_r435_c20 bl[20] br[20] wl[435] vdd gnd cell_6t
Xbit_r436_c20 bl[20] br[20] wl[436] vdd gnd cell_6t
Xbit_r437_c20 bl[20] br[20] wl[437] vdd gnd cell_6t
Xbit_r438_c20 bl[20] br[20] wl[438] vdd gnd cell_6t
Xbit_r439_c20 bl[20] br[20] wl[439] vdd gnd cell_6t
Xbit_r440_c20 bl[20] br[20] wl[440] vdd gnd cell_6t
Xbit_r441_c20 bl[20] br[20] wl[441] vdd gnd cell_6t
Xbit_r442_c20 bl[20] br[20] wl[442] vdd gnd cell_6t
Xbit_r443_c20 bl[20] br[20] wl[443] vdd gnd cell_6t
Xbit_r444_c20 bl[20] br[20] wl[444] vdd gnd cell_6t
Xbit_r445_c20 bl[20] br[20] wl[445] vdd gnd cell_6t
Xbit_r446_c20 bl[20] br[20] wl[446] vdd gnd cell_6t
Xbit_r447_c20 bl[20] br[20] wl[447] vdd gnd cell_6t
Xbit_r448_c20 bl[20] br[20] wl[448] vdd gnd cell_6t
Xbit_r449_c20 bl[20] br[20] wl[449] vdd gnd cell_6t
Xbit_r450_c20 bl[20] br[20] wl[450] vdd gnd cell_6t
Xbit_r451_c20 bl[20] br[20] wl[451] vdd gnd cell_6t
Xbit_r452_c20 bl[20] br[20] wl[452] vdd gnd cell_6t
Xbit_r453_c20 bl[20] br[20] wl[453] vdd gnd cell_6t
Xbit_r454_c20 bl[20] br[20] wl[454] vdd gnd cell_6t
Xbit_r455_c20 bl[20] br[20] wl[455] vdd gnd cell_6t
Xbit_r456_c20 bl[20] br[20] wl[456] vdd gnd cell_6t
Xbit_r457_c20 bl[20] br[20] wl[457] vdd gnd cell_6t
Xbit_r458_c20 bl[20] br[20] wl[458] vdd gnd cell_6t
Xbit_r459_c20 bl[20] br[20] wl[459] vdd gnd cell_6t
Xbit_r460_c20 bl[20] br[20] wl[460] vdd gnd cell_6t
Xbit_r461_c20 bl[20] br[20] wl[461] vdd gnd cell_6t
Xbit_r462_c20 bl[20] br[20] wl[462] vdd gnd cell_6t
Xbit_r463_c20 bl[20] br[20] wl[463] vdd gnd cell_6t
Xbit_r464_c20 bl[20] br[20] wl[464] vdd gnd cell_6t
Xbit_r465_c20 bl[20] br[20] wl[465] vdd gnd cell_6t
Xbit_r466_c20 bl[20] br[20] wl[466] vdd gnd cell_6t
Xbit_r467_c20 bl[20] br[20] wl[467] vdd gnd cell_6t
Xbit_r468_c20 bl[20] br[20] wl[468] vdd gnd cell_6t
Xbit_r469_c20 bl[20] br[20] wl[469] vdd gnd cell_6t
Xbit_r470_c20 bl[20] br[20] wl[470] vdd gnd cell_6t
Xbit_r471_c20 bl[20] br[20] wl[471] vdd gnd cell_6t
Xbit_r472_c20 bl[20] br[20] wl[472] vdd gnd cell_6t
Xbit_r473_c20 bl[20] br[20] wl[473] vdd gnd cell_6t
Xbit_r474_c20 bl[20] br[20] wl[474] vdd gnd cell_6t
Xbit_r475_c20 bl[20] br[20] wl[475] vdd gnd cell_6t
Xbit_r476_c20 bl[20] br[20] wl[476] vdd gnd cell_6t
Xbit_r477_c20 bl[20] br[20] wl[477] vdd gnd cell_6t
Xbit_r478_c20 bl[20] br[20] wl[478] vdd gnd cell_6t
Xbit_r479_c20 bl[20] br[20] wl[479] vdd gnd cell_6t
Xbit_r480_c20 bl[20] br[20] wl[480] vdd gnd cell_6t
Xbit_r481_c20 bl[20] br[20] wl[481] vdd gnd cell_6t
Xbit_r482_c20 bl[20] br[20] wl[482] vdd gnd cell_6t
Xbit_r483_c20 bl[20] br[20] wl[483] vdd gnd cell_6t
Xbit_r484_c20 bl[20] br[20] wl[484] vdd gnd cell_6t
Xbit_r485_c20 bl[20] br[20] wl[485] vdd gnd cell_6t
Xbit_r486_c20 bl[20] br[20] wl[486] vdd gnd cell_6t
Xbit_r487_c20 bl[20] br[20] wl[487] vdd gnd cell_6t
Xbit_r488_c20 bl[20] br[20] wl[488] vdd gnd cell_6t
Xbit_r489_c20 bl[20] br[20] wl[489] vdd gnd cell_6t
Xbit_r490_c20 bl[20] br[20] wl[490] vdd gnd cell_6t
Xbit_r491_c20 bl[20] br[20] wl[491] vdd gnd cell_6t
Xbit_r492_c20 bl[20] br[20] wl[492] vdd gnd cell_6t
Xbit_r493_c20 bl[20] br[20] wl[493] vdd gnd cell_6t
Xbit_r494_c20 bl[20] br[20] wl[494] vdd gnd cell_6t
Xbit_r495_c20 bl[20] br[20] wl[495] vdd gnd cell_6t
Xbit_r496_c20 bl[20] br[20] wl[496] vdd gnd cell_6t
Xbit_r497_c20 bl[20] br[20] wl[497] vdd gnd cell_6t
Xbit_r498_c20 bl[20] br[20] wl[498] vdd gnd cell_6t
Xbit_r499_c20 bl[20] br[20] wl[499] vdd gnd cell_6t
Xbit_r500_c20 bl[20] br[20] wl[500] vdd gnd cell_6t
Xbit_r501_c20 bl[20] br[20] wl[501] vdd gnd cell_6t
Xbit_r502_c20 bl[20] br[20] wl[502] vdd gnd cell_6t
Xbit_r503_c20 bl[20] br[20] wl[503] vdd gnd cell_6t
Xbit_r504_c20 bl[20] br[20] wl[504] vdd gnd cell_6t
Xbit_r505_c20 bl[20] br[20] wl[505] vdd gnd cell_6t
Xbit_r506_c20 bl[20] br[20] wl[506] vdd gnd cell_6t
Xbit_r507_c20 bl[20] br[20] wl[507] vdd gnd cell_6t
Xbit_r508_c20 bl[20] br[20] wl[508] vdd gnd cell_6t
Xbit_r509_c20 bl[20] br[20] wl[509] vdd gnd cell_6t
Xbit_r510_c20 bl[20] br[20] wl[510] vdd gnd cell_6t
Xbit_r511_c20 bl[20] br[20] wl[511] vdd gnd cell_6t
Xbit_r0_c21 bl[21] br[21] wl[0] vdd gnd cell_6t
Xbit_r1_c21 bl[21] br[21] wl[1] vdd gnd cell_6t
Xbit_r2_c21 bl[21] br[21] wl[2] vdd gnd cell_6t
Xbit_r3_c21 bl[21] br[21] wl[3] vdd gnd cell_6t
Xbit_r4_c21 bl[21] br[21] wl[4] vdd gnd cell_6t
Xbit_r5_c21 bl[21] br[21] wl[5] vdd gnd cell_6t
Xbit_r6_c21 bl[21] br[21] wl[6] vdd gnd cell_6t
Xbit_r7_c21 bl[21] br[21] wl[7] vdd gnd cell_6t
Xbit_r8_c21 bl[21] br[21] wl[8] vdd gnd cell_6t
Xbit_r9_c21 bl[21] br[21] wl[9] vdd gnd cell_6t
Xbit_r10_c21 bl[21] br[21] wl[10] vdd gnd cell_6t
Xbit_r11_c21 bl[21] br[21] wl[11] vdd gnd cell_6t
Xbit_r12_c21 bl[21] br[21] wl[12] vdd gnd cell_6t
Xbit_r13_c21 bl[21] br[21] wl[13] vdd gnd cell_6t
Xbit_r14_c21 bl[21] br[21] wl[14] vdd gnd cell_6t
Xbit_r15_c21 bl[21] br[21] wl[15] vdd gnd cell_6t
Xbit_r16_c21 bl[21] br[21] wl[16] vdd gnd cell_6t
Xbit_r17_c21 bl[21] br[21] wl[17] vdd gnd cell_6t
Xbit_r18_c21 bl[21] br[21] wl[18] vdd gnd cell_6t
Xbit_r19_c21 bl[21] br[21] wl[19] vdd gnd cell_6t
Xbit_r20_c21 bl[21] br[21] wl[20] vdd gnd cell_6t
Xbit_r21_c21 bl[21] br[21] wl[21] vdd gnd cell_6t
Xbit_r22_c21 bl[21] br[21] wl[22] vdd gnd cell_6t
Xbit_r23_c21 bl[21] br[21] wl[23] vdd gnd cell_6t
Xbit_r24_c21 bl[21] br[21] wl[24] vdd gnd cell_6t
Xbit_r25_c21 bl[21] br[21] wl[25] vdd gnd cell_6t
Xbit_r26_c21 bl[21] br[21] wl[26] vdd gnd cell_6t
Xbit_r27_c21 bl[21] br[21] wl[27] vdd gnd cell_6t
Xbit_r28_c21 bl[21] br[21] wl[28] vdd gnd cell_6t
Xbit_r29_c21 bl[21] br[21] wl[29] vdd gnd cell_6t
Xbit_r30_c21 bl[21] br[21] wl[30] vdd gnd cell_6t
Xbit_r31_c21 bl[21] br[21] wl[31] vdd gnd cell_6t
Xbit_r32_c21 bl[21] br[21] wl[32] vdd gnd cell_6t
Xbit_r33_c21 bl[21] br[21] wl[33] vdd gnd cell_6t
Xbit_r34_c21 bl[21] br[21] wl[34] vdd gnd cell_6t
Xbit_r35_c21 bl[21] br[21] wl[35] vdd gnd cell_6t
Xbit_r36_c21 bl[21] br[21] wl[36] vdd gnd cell_6t
Xbit_r37_c21 bl[21] br[21] wl[37] vdd gnd cell_6t
Xbit_r38_c21 bl[21] br[21] wl[38] vdd gnd cell_6t
Xbit_r39_c21 bl[21] br[21] wl[39] vdd gnd cell_6t
Xbit_r40_c21 bl[21] br[21] wl[40] vdd gnd cell_6t
Xbit_r41_c21 bl[21] br[21] wl[41] vdd gnd cell_6t
Xbit_r42_c21 bl[21] br[21] wl[42] vdd gnd cell_6t
Xbit_r43_c21 bl[21] br[21] wl[43] vdd gnd cell_6t
Xbit_r44_c21 bl[21] br[21] wl[44] vdd gnd cell_6t
Xbit_r45_c21 bl[21] br[21] wl[45] vdd gnd cell_6t
Xbit_r46_c21 bl[21] br[21] wl[46] vdd gnd cell_6t
Xbit_r47_c21 bl[21] br[21] wl[47] vdd gnd cell_6t
Xbit_r48_c21 bl[21] br[21] wl[48] vdd gnd cell_6t
Xbit_r49_c21 bl[21] br[21] wl[49] vdd gnd cell_6t
Xbit_r50_c21 bl[21] br[21] wl[50] vdd gnd cell_6t
Xbit_r51_c21 bl[21] br[21] wl[51] vdd gnd cell_6t
Xbit_r52_c21 bl[21] br[21] wl[52] vdd gnd cell_6t
Xbit_r53_c21 bl[21] br[21] wl[53] vdd gnd cell_6t
Xbit_r54_c21 bl[21] br[21] wl[54] vdd gnd cell_6t
Xbit_r55_c21 bl[21] br[21] wl[55] vdd gnd cell_6t
Xbit_r56_c21 bl[21] br[21] wl[56] vdd gnd cell_6t
Xbit_r57_c21 bl[21] br[21] wl[57] vdd gnd cell_6t
Xbit_r58_c21 bl[21] br[21] wl[58] vdd gnd cell_6t
Xbit_r59_c21 bl[21] br[21] wl[59] vdd gnd cell_6t
Xbit_r60_c21 bl[21] br[21] wl[60] vdd gnd cell_6t
Xbit_r61_c21 bl[21] br[21] wl[61] vdd gnd cell_6t
Xbit_r62_c21 bl[21] br[21] wl[62] vdd gnd cell_6t
Xbit_r63_c21 bl[21] br[21] wl[63] vdd gnd cell_6t
Xbit_r64_c21 bl[21] br[21] wl[64] vdd gnd cell_6t
Xbit_r65_c21 bl[21] br[21] wl[65] vdd gnd cell_6t
Xbit_r66_c21 bl[21] br[21] wl[66] vdd gnd cell_6t
Xbit_r67_c21 bl[21] br[21] wl[67] vdd gnd cell_6t
Xbit_r68_c21 bl[21] br[21] wl[68] vdd gnd cell_6t
Xbit_r69_c21 bl[21] br[21] wl[69] vdd gnd cell_6t
Xbit_r70_c21 bl[21] br[21] wl[70] vdd gnd cell_6t
Xbit_r71_c21 bl[21] br[21] wl[71] vdd gnd cell_6t
Xbit_r72_c21 bl[21] br[21] wl[72] vdd gnd cell_6t
Xbit_r73_c21 bl[21] br[21] wl[73] vdd gnd cell_6t
Xbit_r74_c21 bl[21] br[21] wl[74] vdd gnd cell_6t
Xbit_r75_c21 bl[21] br[21] wl[75] vdd gnd cell_6t
Xbit_r76_c21 bl[21] br[21] wl[76] vdd gnd cell_6t
Xbit_r77_c21 bl[21] br[21] wl[77] vdd gnd cell_6t
Xbit_r78_c21 bl[21] br[21] wl[78] vdd gnd cell_6t
Xbit_r79_c21 bl[21] br[21] wl[79] vdd gnd cell_6t
Xbit_r80_c21 bl[21] br[21] wl[80] vdd gnd cell_6t
Xbit_r81_c21 bl[21] br[21] wl[81] vdd gnd cell_6t
Xbit_r82_c21 bl[21] br[21] wl[82] vdd gnd cell_6t
Xbit_r83_c21 bl[21] br[21] wl[83] vdd gnd cell_6t
Xbit_r84_c21 bl[21] br[21] wl[84] vdd gnd cell_6t
Xbit_r85_c21 bl[21] br[21] wl[85] vdd gnd cell_6t
Xbit_r86_c21 bl[21] br[21] wl[86] vdd gnd cell_6t
Xbit_r87_c21 bl[21] br[21] wl[87] vdd gnd cell_6t
Xbit_r88_c21 bl[21] br[21] wl[88] vdd gnd cell_6t
Xbit_r89_c21 bl[21] br[21] wl[89] vdd gnd cell_6t
Xbit_r90_c21 bl[21] br[21] wl[90] vdd gnd cell_6t
Xbit_r91_c21 bl[21] br[21] wl[91] vdd gnd cell_6t
Xbit_r92_c21 bl[21] br[21] wl[92] vdd gnd cell_6t
Xbit_r93_c21 bl[21] br[21] wl[93] vdd gnd cell_6t
Xbit_r94_c21 bl[21] br[21] wl[94] vdd gnd cell_6t
Xbit_r95_c21 bl[21] br[21] wl[95] vdd gnd cell_6t
Xbit_r96_c21 bl[21] br[21] wl[96] vdd gnd cell_6t
Xbit_r97_c21 bl[21] br[21] wl[97] vdd gnd cell_6t
Xbit_r98_c21 bl[21] br[21] wl[98] vdd gnd cell_6t
Xbit_r99_c21 bl[21] br[21] wl[99] vdd gnd cell_6t
Xbit_r100_c21 bl[21] br[21] wl[100] vdd gnd cell_6t
Xbit_r101_c21 bl[21] br[21] wl[101] vdd gnd cell_6t
Xbit_r102_c21 bl[21] br[21] wl[102] vdd gnd cell_6t
Xbit_r103_c21 bl[21] br[21] wl[103] vdd gnd cell_6t
Xbit_r104_c21 bl[21] br[21] wl[104] vdd gnd cell_6t
Xbit_r105_c21 bl[21] br[21] wl[105] vdd gnd cell_6t
Xbit_r106_c21 bl[21] br[21] wl[106] vdd gnd cell_6t
Xbit_r107_c21 bl[21] br[21] wl[107] vdd gnd cell_6t
Xbit_r108_c21 bl[21] br[21] wl[108] vdd gnd cell_6t
Xbit_r109_c21 bl[21] br[21] wl[109] vdd gnd cell_6t
Xbit_r110_c21 bl[21] br[21] wl[110] vdd gnd cell_6t
Xbit_r111_c21 bl[21] br[21] wl[111] vdd gnd cell_6t
Xbit_r112_c21 bl[21] br[21] wl[112] vdd gnd cell_6t
Xbit_r113_c21 bl[21] br[21] wl[113] vdd gnd cell_6t
Xbit_r114_c21 bl[21] br[21] wl[114] vdd gnd cell_6t
Xbit_r115_c21 bl[21] br[21] wl[115] vdd gnd cell_6t
Xbit_r116_c21 bl[21] br[21] wl[116] vdd gnd cell_6t
Xbit_r117_c21 bl[21] br[21] wl[117] vdd gnd cell_6t
Xbit_r118_c21 bl[21] br[21] wl[118] vdd gnd cell_6t
Xbit_r119_c21 bl[21] br[21] wl[119] vdd gnd cell_6t
Xbit_r120_c21 bl[21] br[21] wl[120] vdd gnd cell_6t
Xbit_r121_c21 bl[21] br[21] wl[121] vdd gnd cell_6t
Xbit_r122_c21 bl[21] br[21] wl[122] vdd gnd cell_6t
Xbit_r123_c21 bl[21] br[21] wl[123] vdd gnd cell_6t
Xbit_r124_c21 bl[21] br[21] wl[124] vdd gnd cell_6t
Xbit_r125_c21 bl[21] br[21] wl[125] vdd gnd cell_6t
Xbit_r126_c21 bl[21] br[21] wl[126] vdd gnd cell_6t
Xbit_r127_c21 bl[21] br[21] wl[127] vdd gnd cell_6t
Xbit_r128_c21 bl[21] br[21] wl[128] vdd gnd cell_6t
Xbit_r129_c21 bl[21] br[21] wl[129] vdd gnd cell_6t
Xbit_r130_c21 bl[21] br[21] wl[130] vdd gnd cell_6t
Xbit_r131_c21 bl[21] br[21] wl[131] vdd gnd cell_6t
Xbit_r132_c21 bl[21] br[21] wl[132] vdd gnd cell_6t
Xbit_r133_c21 bl[21] br[21] wl[133] vdd gnd cell_6t
Xbit_r134_c21 bl[21] br[21] wl[134] vdd gnd cell_6t
Xbit_r135_c21 bl[21] br[21] wl[135] vdd gnd cell_6t
Xbit_r136_c21 bl[21] br[21] wl[136] vdd gnd cell_6t
Xbit_r137_c21 bl[21] br[21] wl[137] vdd gnd cell_6t
Xbit_r138_c21 bl[21] br[21] wl[138] vdd gnd cell_6t
Xbit_r139_c21 bl[21] br[21] wl[139] vdd gnd cell_6t
Xbit_r140_c21 bl[21] br[21] wl[140] vdd gnd cell_6t
Xbit_r141_c21 bl[21] br[21] wl[141] vdd gnd cell_6t
Xbit_r142_c21 bl[21] br[21] wl[142] vdd gnd cell_6t
Xbit_r143_c21 bl[21] br[21] wl[143] vdd gnd cell_6t
Xbit_r144_c21 bl[21] br[21] wl[144] vdd gnd cell_6t
Xbit_r145_c21 bl[21] br[21] wl[145] vdd gnd cell_6t
Xbit_r146_c21 bl[21] br[21] wl[146] vdd gnd cell_6t
Xbit_r147_c21 bl[21] br[21] wl[147] vdd gnd cell_6t
Xbit_r148_c21 bl[21] br[21] wl[148] vdd gnd cell_6t
Xbit_r149_c21 bl[21] br[21] wl[149] vdd gnd cell_6t
Xbit_r150_c21 bl[21] br[21] wl[150] vdd gnd cell_6t
Xbit_r151_c21 bl[21] br[21] wl[151] vdd gnd cell_6t
Xbit_r152_c21 bl[21] br[21] wl[152] vdd gnd cell_6t
Xbit_r153_c21 bl[21] br[21] wl[153] vdd gnd cell_6t
Xbit_r154_c21 bl[21] br[21] wl[154] vdd gnd cell_6t
Xbit_r155_c21 bl[21] br[21] wl[155] vdd gnd cell_6t
Xbit_r156_c21 bl[21] br[21] wl[156] vdd gnd cell_6t
Xbit_r157_c21 bl[21] br[21] wl[157] vdd gnd cell_6t
Xbit_r158_c21 bl[21] br[21] wl[158] vdd gnd cell_6t
Xbit_r159_c21 bl[21] br[21] wl[159] vdd gnd cell_6t
Xbit_r160_c21 bl[21] br[21] wl[160] vdd gnd cell_6t
Xbit_r161_c21 bl[21] br[21] wl[161] vdd gnd cell_6t
Xbit_r162_c21 bl[21] br[21] wl[162] vdd gnd cell_6t
Xbit_r163_c21 bl[21] br[21] wl[163] vdd gnd cell_6t
Xbit_r164_c21 bl[21] br[21] wl[164] vdd gnd cell_6t
Xbit_r165_c21 bl[21] br[21] wl[165] vdd gnd cell_6t
Xbit_r166_c21 bl[21] br[21] wl[166] vdd gnd cell_6t
Xbit_r167_c21 bl[21] br[21] wl[167] vdd gnd cell_6t
Xbit_r168_c21 bl[21] br[21] wl[168] vdd gnd cell_6t
Xbit_r169_c21 bl[21] br[21] wl[169] vdd gnd cell_6t
Xbit_r170_c21 bl[21] br[21] wl[170] vdd gnd cell_6t
Xbit_r171_c21 bl[21] br[21] wl[171] vdd gnd cell_6t
Xbit_r172_c21 bl[21] br[21] wl[172] vdd gnd cell_6t
Xbit_r173_c21 bl[21] br[21] wl[173] vdd gnd cell_6t
Xbit_r174_c21 bl[21] br[21] wl[174] vdd gnd cell_6t
Xbit_r175_c21 bl[21] br[21] wl[175] vdd gnd cell_6t
Xbit_r176_c21 bl[21] br[21] wl[176] vdd gnd cell_6t
Xbit_r177_c21 bl[21] br[21] wl[177] vdd gnd cell_6t
Xbit_r178_c21 bl[21] br[21] wl[178] vdd gnd cell_6t
Xbit_r179_c21 bl[21] br[21] wl[179] vdd gnd cell_6t
Xbit_r180_c21 bl[21] br[21] wl[180] vdd gnd cell_6t
Xbit_r181_c21 bl[21] br[21] wl[181] vdd gnd cell_6t
Xbit_r182_c21 bl[21] br[21] wl[182] vdd gnd cell_6t
Xbit_r183_c21 bl[21] br[21] wl[183] vdd gnd cell_6t
Xbit_r184_c21 bl[21] br[21] wl[184] vdd gnd cell_6t
Xbit_r185_c21 bl[21] br[21] wl[185] vdd gnd cell_6t
Xbit_r186_c21 bl[21] br[21] wl[186] vdd gnd cell_6t
Xbit_r187_c21 bl[21] br[21] wl[187] vdd gnd cell_6t
Xbit_r188_c21 bl[21] br[21] wl[188] vdd gnd cell_6t
Xbit_r189_c21 bl[21] br[21] wl[189] vdd gnd cell_6t
Xbit_r190_c21 bl[21] br[21] wl[190] vdd gnd cell_6t
Xbit_r191_c21 bl[21] br[21] wl[191] vdd gnd cell_6t
Xbit_r192_c21 bl[21] br[21] wl[192] vdd gnd cell_6t
Xbit_r193_c21 bl[21] br[21] wl[193] vdd gnd cell_6t
Xbit_r194_c21 bl[21] br[21] wl[194] vdd gnd cell_6t
Xbit_r195_c21 bl[21] br[21] wl[195] vdd gnd cell_6t
Xbit_r196_c21 bl[21] br[21] wl[196] vdd gnd cell_6t
Xbit_r197_c21 bl[21] br[21] wl[197] vdd gnd cell_6t
Xbit_r198_c21 bl[21] br[21] wl[198] vdd gnd cell_6t
Xbit_r199_c21 bl[21] br[21] wl[199] vdd gnd cell_6t
Xbit_r200_c21 bl[21] br[21] wl[200] vdd gnd cell_6t
Xbit_r201_c21 bl[21] br[21] wl[201] vdd gnd cell_6t
Xbit_r202_c21 bl[21] br[21] wl[202] vdd gnd cell_6t
Xbit_r203_c21 bl[21] br[21] wl[203] vdd gnd cell_6t
Xbit_r204_c21 bl[21] br[21] wl[204] vdd gnd cell_6t
Xbit_r205_c21 bl[21] br[21] wl[205] vdd gnd cell_6t
Xbit_r206_c21 bl[21] br[21] wl[206] vdd gnd cell_6t
Xbit_r207_c21 bl[21] br[21] wl[207] vdd gnd cell_6t
Xbit_r208_c21 bl[21] br[21] wl[208] vdd gnd cell_6t
Xbit_r209_c21 bl[21] br[21] wl[209] vdd gnd cell_6t
Xbit_r210_c21 bl[21] br[21] wl[210] vdd gnd cell_6t
Xbit_r211_c21 bl[21] br[21] wl[211] vdd gnd cell_6t
Xbit_r212_c21 bl[21] br[21] wl[212] vdd gnd cell_6t
Xbit_r213_c21 bl[21] br[21] wl[213] vdd gnd cell_6t
Xbit_r214_c21 bl[21] br[21] wl[214] vdd gnd cell_6t
Xbit_r215_c21 bl[21] br[21] wl[215] vdd gnd cell_6t
Xbit_r216_c21 bl[21] br[21] wl[216] vdd gnd cell_6t
Xbit_r217_c21 bl[21] br[21] wl[217] vdd gnd cell_6t
Xbit_r218_c21 bl[21] br[21] wl[218] vdd gnd cell_6t
Xbit_r219_c21 bl[21] br[21] wl[219] vdd gnd cell_6t
Xbit_r220_c21 bl[21] br[21] wl[220] vdd gnd cell_6t
Xbit_r221_c21 bl[21] br[21] wl[221] vdd gnd cell_6t
Xbit_r222_c21 bl[21] br[21] wl[222] vdd gnd cell_6t
Xbit_r223_c21 bl[21] br[21] wl[223] vdd gnd cell_6t
Xbit_r224_c21 bl[21] br[21] wl[224] vdd gnd cell_6t
Xbit_r225_c21 bl[21] br[21] wl[225] vdd gnd cell_6t
Xbit_r226_c21 bl[21] br[21] wl[226] vdd gnd cell_6t
Xbit_r227_c21 bl[21] br[21] wl[227] vdd gnd cell_6t
Xbit_r228_c21 bl[21] br[21] wl[228] vdd gnd cell_6t
Xbit_r229_c21 bl[21] br[21] wl[229] vdd gnd cell_6t
Xbit_r230_c21 bl[21] br[21] wl[230] vdd gnd cell_6t
Xbit_r231_c21 bl[21] br[21] wl[231] vdd gnd cell_6t
Xbit_r232_c21 bl[21] br[21] wl[232] vdd gnd cell_6t
Xbit_r233_c21 bl[21] br[21] wl[233] vdd gnd cell_6t
Xbit_r234_c21 bl[21] br[21] wl[234] vdd gnd cell_6t
Xbit_r235_c21 bl[21] br[21] wl[235] vdd gnd cell_6t
Xbit_r236_c21 bl[21] br[21] wl[236] vdd gnd cell_6t
Xbit_r237_c21 bl[21] br[21] wl[237] vdd gnd cell_6t
Xbit_r238_c21 bl[21] br[21] wl[238] vdd gnd cell_6t
Xbit_r239_c21 bl[21] br[21] wl[239] vdd gnd cell_6t
Xbit_r240_c21 bl[21] br[21] wl[240] vdd gnd cell_6t
Xbit_r241_c21 bl[21] br[21] wl[241] vdd gnd cell_6t
Xbit_r242_c21 bl[21] br[21] wl[242] vdd gnd cell_6t
Xbit_r243_c21 bl[21] br[21] wl[243] vdd gnd cell_6t
Xbit_r244_c21 bl[21] br[21] wl[244] vdd gnd cell_6t
Xbit_r245_c21 bl[21] br[21] wl[245] vdd gnd cell_6t
Xbit_r246_c21 bl[21] br[21] wl[246] vdd gnd cell_6t
Xbit_r247_c21 bl[21] br[21] wl[247] vdd gnd cell_6t
Xbit_r248_c21 bl[21] br[21] wl[248] vdd gnd cell_6t
Xbit_r249_c21 bl[21] br[21] wl[249] vdd gnd cell_6t
Xbit_r250_c21 bl[21] br[21] wl[250] vdd gnd cell_6t
Xbit_r251_c21 bl[21] br[21] wl[251] vdd gnd cell_6t
Xbit_r252_c21 bl[21] br[21] wl[252] vdd gnd cell_6t
Xbit_r253_c21 bl[21] br[21] wl[253] vdd gnd cell_6t
Xbit_r254_c21 bl[21] br[21] wl[254] vdd gnd cell_6t
Xbit_r255_c21 bl[21] br[21] wl[255] vdd gnd cell_6t
Xbit_r256_c21 bl[21] br[21] wl[256] vdd gnd cell_6t
Xbit_r257_c21 bl[21] br[21] wl[257] vdd gnd cell_6t
Xbit_r258_c21 bl[21] br[21] wl[258] vdd gnd cell_6t
Xbit_r259_c21 bl[21] br[21] wl[259] vdd gnd cell_6t
Xbit_r260_c21 bl[21] br[21] wl[260] vdd gnd cell_6t
Xbit_r261_c21 bl[21] br[21] wl[261] vdd gnd cell_6t
Xbit_r262_c21 bl[21] br[21] wl[262] vdd gnd cell_6t
Xbit_r263_c21 bl[21] br[21] wl[263] vdd gnd cell_6t
Xbit_r264_c21 bl[21] br[21] wl[264] vdd gnd cell_6t
Xbit_r265_c21 bl[21] br[21] wl[265] vdd gnd cell_6t
Xbit_r266_c21 bl[21] br[21] wl[266] vdd gnd cell_6t
Xbit_r267_c21 bl[21] br[21] wl[267] vdd gnd cell_6t
Xbit_r268_c21 bl[21] br[21] wl[268] vdd gnd cell_6t
Xbit_r269_c21 bl[21] br[21] wl[269] vdd gnd cell_6t
Xbit_r270_c21 bl[21] br[21] wl[270] vdd gnd cell_6t
Xbit_r271_c21 bl[21] br[21] wl[271] vdd gnd cell_6t
Xbit_r272_c21 bl[21] br[21] wl[272] vdd gnd cell_6t
Xbit_r273_c21 bl[21] br[21] wl[273] vdd gnd cell_6t
Xbit_r274_c21 bl[21] br[21] wl[274] vdd gnd cell_6t
Xbit_r275_c21 bl[21] br[21] wl[275] vdd gnd cell_6t
Xbit_r276_c21 bl[21] br[21] wl[276] vdd gnd cell_6t
Xbit_r277_c21 bl[21] br[21] wl[277] vdd gnd cell_6t
Xbit_r278_c21 bl[21] br[21] wl[278] vdd gnd cell_6t
Xbit_r279_c21 bl[21] br[21] wl[279] vdd gnd cell_6t
Xbit_r280_c21 bl[21] br[21] wl[280] vdd gnd cell_6t
Xbit_r281_c21 bl[21] br[21] wl[281] vdd gnd cell_6t
Xbit_r282_c21 bl[21] br[21] wl[282] vdd gnd cell_6t
Xbit_r283_c21 bl[21] br[21] wl[283] vdd gnd cell_6t
Xbit_r284_c21 bl[21] br[21] wl[284] vdd gnd cell_6t
Xbit_r285_c21 bl[21] br[21] wl[285] vdd gnd cell_6t
Xbit_r286_c21 bl[21] br[21] wl[286] vdd gnd cell_6t
Xbit_r287_c21 bl[21] br[21] wl[287] vdd gnd cell_6t
Xbit_r288_c21 bl[21] br[21] wl[288] vdd gnd cell_6t
Xbit_r289_c21 bl[21] br[21] wl[289] vdd gnd cell_6t
Xbit_r290_c21 bl[21] br[21] wl[290] vdd gnd cell_6t
Xbit_r291_c21 bl[21] br[21] wl[291] vdd gnd cell_6t
Xbit_r292_c21 bl[21] br[21] wl[292] vdd gnd cell_6t
Xbit_r293_c21 bl[21] br[21] wl[293] vdd gnd cell_6t
Xbit_r294_c21 bl[21] br[21] wl[294] vdd gnd cell_6t
Xbit_r295_c21 bl[21] br[21] wl[295] vdd gnd cell_6t
Xbit_r296_c21 bl[21] br[21] wl[296] vdd gnd cell_6t
Xbit_r297_c21 bl[21] br[21] wl[297] vdd gnd cell_6t
Xbit_r298_c21 bl[21] br[21] wl[298] vdd gnd cell_6t
Xbit_r299_c21 bl[21] br[21] wl[299] vdd gnd cell_6t
Xbit_r300_c21 bl[21] br[21] wl[300] vdd gnd cell_6t
Xbit_r301_c21 bl[21] br[21] wl[301] vdd gnd cell_6t
Xbit_r302_c21 bl[21] br[21] wl[302] vdd gnd cell_6t
Xbit_r303_c21 bl[21] br[21] wl[303] vdd gnd cell_6t
Xbit_r304_c21 bl[21] br[21] wl[304] vdd gnd cell_6t
Xbit_r305_c21 bl[21] br[21] wl[305] vdd gnd cell_6t
Xbit_r306_c21 bl[21] br[21] wl[306] vdd gnd cell_6t
Xbit_r307_c21 bl[21] br[21] wl[307] vdd gnd cell_6t
Xbit_r308_c21 bl[21] br[21] wl[308] vdd gnd cell_6t
Xbit_r309_c21 bl[21] br[21] wl[309] vdd gnd cell_6t
Xbit_r310_c21 bl[21] br[21] wl[310] vdd gnd cell_6t
Xbit_r311_c21 bl[21] br[21] wl[311] vdd gnd cell_6t
Xbit_r312_c21 bl[21] br[21] wl[312] vdd gnd cell_6t
Xbit_r313_c21 bl[21] br[21] wl[313] vdd gnd cell_6t
Xbit_r314_c21 bl[21] br[21] wl[314] vdd gnd cell_6t
Xbit_r315_c21 bl[21] br[21] wl[315] vdd gnd cell_6t
Xbit_r316_c21 bl[21] br[21] wl[316] vdd gnd cell_6t
Xbit_r317_c21 bl[21] br[21] wl[317] vdd gnd cell_6t
Xbit_r318_c21 bl[21] br[21] wl[318] vdd gnd cell_6t
Xbit_r319_c21 bl[21] br[21] wl[319] vdd gnd cell_6t
Xbit_r320_c21 bl[21] br[21] wl[320] vdd gnd cell_6t
Xbit_r321_c21 bl[21] br[21] wl[321] vdd gnd cell_6t
Xbit_r322_c21 bl[21] br[21] wl[322] vdd gnd cell_6t
Xbit_r323_c21 bl[21] br[21] wl[323] vdd gnd cell_6t
Xbit_r324_c21 bl[21] br[21] wl[324] vdd gnd cell_6t
Xbit_r325_c21 bl[21] br[21] wl[325] vdd gnd cell_6t
Xbit_r326_c21 bl[21] br[21] wl[326] vdd gnd cell_6t
Xbit_r327_c21 bl[21] br[21] wl[327] vdd gnd cell_6t
Xbit_r328_c21 bl[21] br[21] wl[328] vdd gnd cell_6t
Xbit_r329_c21 bl[21] br[21] wl[329] vdd gnd cell_6t
Xbit_r330_c21 bl[21] br[21] wl[330] vdd gnd cell_6t
Xbit_r331_c21 bl[21] br[21] wl[331] vdd gnd cell_6t
Xbit_r332_c21 bl[21] br[21] wl[332] vdd gnd cell_6t
Xbit_r333_c21 bl[21] br[21] wl[333] vdd gnd cell_6t
Xbit_r334_c21 bl[21] br[21] wl[334] vdd gnd cell_6t
Xbit_r335_c21 bl[21] br[21] wl[335] vdd gnd cell_6t
Xbit_r336_c21 bl[21] br[21] wl[336] vdd gnd cell_6t
Xbit_r337_c21 bl[21] br[21] wl[337] vdd gnd cell_6t
Xbit_r338_c21 bl[21] br[21] wl[338] vdd gnd cell_6t
Xbit_r339_c21 bl[21] br[21] wl[339] vdd gnd cell_6t
Xbit_r340_c21 bl[21] br[21] wl[340] vdd gnd cell_6t
Xbit_r341_c21 bl[21] br[21] wl[341] vdd gnd cell_6t
Xbit_r342_c21 bl[21] br[21] wl[342] vdd gnd cell_6t
Xbit_r343_c21 bl[21] br[21] wl[343] vdd gnd cell_6t
Xbit_r344_c21 bl[21] br[21] wl[344] vdd gnd cell_6t
Xbit_r345_c21 bl[21] br[21] wl[345] vdd gnd cell_6t
Xbit_r346_c21 bl[21] br[21] wl[346] vdd gnd cell_6t
Xbit_r347_c21 bl[21] br[21] wl[347] vdd gnd cell_6t
Xbit_r348_c21 bl[21] br[21] wl[348] vdd gnd cell_6t
Xbit_r349_c21 bl[21] br[21] wl[349] vdd gnd cell_6t
Xbit_r350_c21 bl[21] br[21] wl[350] vdd gnd cell_6t
Xbit_r351_c21 bl[21] br[21] wl[351] vdd gnd cell_6t
Xbit_r352_c21 bl[21] br[21] wl[352] vdd gnd cell_6t
Xbit_r353_c21 bl[21] br[21] wl[353] vdd gnd cell_6t
Xbit_r354_c21 bl[21] br[21] wl[354] vdd gnd cell_6t
Xbit_r355_c21 bl[21] br[21] wl[355] vdd gnd cell_6t
Xbit_r356_c21 bl[21] br[21] wl[356] vdd gnd cell_6t
Xbit_r357_c21 bl[21] br[21] wl[357] vdd gnd cell_6t
Xbit_r358_c21 bl[21] br[21] wl[358] vdd gnd cell_6t
Xbit_r359_c21 bl[21] br[21] wl[359] vdd gnd cell_6t
Xbit_r360_c21 bl[21] br[21] wl[360] vdd gnd cell_6t
Xbit_r361_c21 bl[21] br[21] wl[361] vdd gnd cell_6t
Xbit_r362_c21 bl[21] br[21] wl[362] vdd gnd cell_6t
Xbit_r363_c21 bl[21] br[21] wl[363] vdd gnd cell_6t
Xbit_r364_c21 bl[21] br[21] wl[364] vdd gnd cell_6t
Xbit_r365_c21 bl[21] br[21] wl[365] vdd gnd cell_6t
Xbit_r366_c21 bl[21] br[21] wl[366] vdd gnd cell_6t
Xbit_r367_c21 bl[21] br[21] wl[367] vdd gnd cell_6t
Xbit_r368_c21 bl[21] br[21] wl[368] vdd gnd cell_6t
Xbit_r369_c21 bl[21] br[21] wl[369] vdd gnd cell_6t
Xbit_r370_c21 bl[21] br[21] wl[370] vdd gnd cell_6t
Xbit_r371_c21 bl[21] br[21] wl[371] vdd gnd cell_6t
Xbit_r372_c21 bl[21] br[21] wl[372] vdd gnd cell_6t
Xbit_r373_c21 bl[21] br[21] wl[373] vdd gnd cell_6t
Xbit_r374_c21 bl[21] br[21] wl[374] vdd gnd cell_6t
Xbit_r375_c21 bl[21] br[21] wl[375] vdd gnd cell_6t
Xbit_r376_c21 bl[21] br[21] wl[376] vdd gnd cell_6t
Xbit_r377_c21 bl[21] br[21] wl[377] vdd gnd cell_6t
Xbit_r378_c21 bl[21] br[21] wl[378] vdd gnd cell_6t
Xbit_r379_c21 bl[21] br[21] wl[379] vdd gnd cell_6t
Xbit_r380_c21 bl[21] br[21] wl[380] vdd gnd cell_6t
Xbit_r381_c21 bl[21] br[21] wl[381] vdd gnd cell_6t
Xbit_r382_c21 bl[21] br[21] wl[382] vdd gnd cell_6t
Xbit_r383_c21 bl[21] br[21] wl[383] vdd gnd cell_6t
Xbit_r384_c21 bl[21] br[21] wl[384] vdd gnd cell_6t
Xbit_r385_c21 bl[21] br[21] wl[385] vdd gnd cell_6t
Xbit_r386_c21 bl[21] br[21] wl[386] vdd gnd cell_6t
Xbit_r387_c21 bl[21] br[21] wl[387] vdd gnd cell_6t
Xbit_r388_c21 bl[21] br[21] wl[388] vdd gnd cell_6t
Xbit_r389_c21 bl[21] br[21] wl[389] vdd gnd cell_6t
Xbit_r390_c21 bl[21] br[21] wl[390] vdd gnd cell_6t
Xbit_r391_c21 bl[21] br[21] wl[391] vdd gnd cell_6t
Xbit_r392_c21 bl[21] br[21] wl[392] vdd gnd cell_6t
Xbit_r393_c21 bl[21] br[21] wl[393] vdd gnd cell_6t
Xbit_r394_c21 bl[21] br[21] wl[394] vdd gnd cell_6t
Xbit_r395_c21 bl[21] br[21] wl[395] vdd gnd cell_6t
Xbit_r396_c21 bl[21] br[21] wl[396] vdd gnd cell_6t
Xbit_r397_c21 bl[21] br[21] wl[397] vdd gnd cell_6t
Xbit_r398_c21 bl[21] br[21] wl[398] vdd gnd cell_6t
Xbit_r399_c21 bl[21] br[21] wl[399] vdd gnd cell_6t
Xbit_r400_c21 bl[21] br[21] wl[400] vdd gnd cell_6t
Xbit_r401_c21 bl[21] br[21] wl[401] vdd gnd cell_6t
Xbit_r402_c21 bl[21] br[21] wl[402] vdd gnd cell_6t
Xbit_r403_c21 bl[21] br[21] wl[403] vdd gnd cell_6t
Xbit_r404_c21 bl[21] br[21] wl[404] vdd gnd cell_6t
Xbit_r405_c21 bl[21] br[21] wl[405] vdd gnd cell_6t
Xbit_r406_c21 bl[21] br[21] wl[406] vdd gnd cell_6t
Xbit_r407_c21 bl[21] br[21] wl[407] vdd gnd cell_6t
Xbit_r408_c21 bl[21] br[21] wl[408] vdd gnd cell_6t
Xbit_r409_c21 bl[21] br[21] wl[409] vdd gnd cell_6t
Xbit_r410_c21 bl[21] br[21] wl[410] vdd gnd cell_6t
Xbit_r411_c21 bl[21] br[21] wl[411] vdd gnd cell_6t
Xbit_r412_c21 bl[21] br[21] wl[412] vdd gnd cell_6t
Xbit_r413_c21 bl[21] br[21] wl[413] vdd gnd cell_6t
Xbit_r414_c21 bl[21] br[21] wl[414] vdd gnd cell_6t
Xbit_r415_c21 bl[21] br[21] wl[415] vdd gnd cell_6t
Xbit_r416_c21 bl[21] br[21] wl[416] vdd gnd cell_6t
Xbit_r417_c21 bl[21] br[21] wl[417] vdd gnd cell_6t
Xbit_r418_c21 bl[21] br[21] wl[418] vdd gnd cell_6t
Xbit_r419_c21 bl[21] br[21] wl[419] vdd gnd cell_6t
Xbit_r420_c21 bl[21] br[21] wl[420] vdd gnd cell_6t
Xbit_r421_c21 bl[21] br[21] wl[421] vdd gnd cell_6t
Xbit_r422_c21 bl[21] br[21] wl[422] vdd gnd cell_6t
Xbit_r423_c21 bl[21] br[21] wl[423] vdd gnd cell_6t
Xbit_r424_c21 bl[21] br[21] wl[424] vdd gnd cell_6t
Xbit_r425_c21 bl[21] br[21] wl[425] vdd gnd cell_6t
Xbit_r426_c21 bl[21] br[21] wl[426] vdd gnd cell_6t
Xbit_r427_c21 bl[21] br[21] wl[427] vdd gnd cell_6t
Xbit_r428_c21 bl[21] br[21] wl[428] vdd gnd cell_6t
Xbit_r429_c21 bl[21] br[21] wl[429] vdd gnd cell_6t
Xbit_r430_c21 bl[21] br[21] wl[430] vdd gnd cell_6t
Xbit_r431_c21 bl[21] br[21] wl[431] vdd gnd cell_6t
Xbit_r432_c21 bl[21] br[21] wl[432] vdd gnd cell_6t
Xbit_r433_c21 bl[21] br[21] wl[433] vdd gnd cell_6t
Xbit_r434_c21 bl[21] br[21] wl[434] vdd gnd cell_6t
Xbit_r435_c21 bl[21] br[21] wl[435] vdd gnd cell_6t
Xbit_r436_c21 bl[21] br[21] wl[436] vdd gnd cell_6t
Xbit_r437_c21 bl[21] br[21] wl[437] vdd gnd cell_6t
Xbit_r438_c21 bl[21] br[21] wl[438] vdd gnd cell_6t
Xbit_r439_c21 bl[21] br[21] wl[439] vdd gnd cell_6t
Xbit_r440_c21 bl[21] br[21] wl[440] vdd gnd cell_6t
Xbit_r441_c21 bl[21] br[21] wl[441] vdd gnd cell_6t
Xbit_r442_c21 bl[21] br[21] wl[442] vdd gnd cell_6t
Xbit_r443_c21 bl[21] br[21] wl[443] vdd gnd cell_6t
Xbit_r444_c21 bl[21] br[21] wl[444] vdd gnd cell_6t
Xbit_r445_c21 bl[21] br[21] wl[445] vdd gnd cell_6t
Xbit_r446_c21 bl[21] br[21] wl[446] vdd gnd cell_6t
Xbit_r447_c21 bl[21] br[21] wl[447] vdd gnd cell_6t
Xbit_r448_c21 bl[21] br[21] wl[448] vdd gnd cell_6t
Xbit_r449_c21 bl[21] br[21] wl[449] vdd gnd cell_6t
Xbit_r450_c21 bl[21] br[21] wl[450] vdd gnd cell_6t
Xbit_r451_c21 bl[21] br[21] wl[451] vdd gnd cell_6t
Xbit_r452_c21 bl[21] br[21] wl[452] vdd gnd cell_6t
Xbit_r453_c21 bl[21] br[21] wl[453] vdd gnd cell_6t
Xbit_r454_c21 bl[21] br[21] wl[454] vdd gnd cell_6t
Xbit_r455_c21 bl[21] br[21] wl[455] vdd gnd cell_6t
Xbit_r456_c21 bl[21] br[21] wl[456] vdd gnd cell_6t
Xbit_r457_c21 bl[21] br[21] wl[457] vdd gnd cell_6t
Xbit_r458_c21 bl[21] br[21] wl[458] vdd gnd cell_6t
Xbit_r459_c21 bl[21] br[21] wl[459] vdd gnd cell_6t
Xbit_r460_c21 bl[21] br[21] wl[460] vdd gnd cell_6t
Xbit_r461_c21 bl[21] br[21] wl[461] vdd gnd cell_6t
Xbit_r462_c21 bl[21] br[21] wl[462] vdd gnd cell_6t
Xbit_r463_c21 bl[21] br[21] wl[463] vdd gnd cell_6t
Xbit_r464_c21 bl[21] br[21] wl[464] vdd gnd cell_6t
Xbit_r465_c21 bl[21] br[21] wl[465] vdd gnd cell_6t
Xbit_r466_c21 bl[21] br[21] wl[466] vdd gnd cell_6t
Xbit_r467_c21 bl[21] br[21] wl[467] vdd gnd cell_6t
Xbit_r468_c21 bl[21] br[21] wl[468] vdd gnd cell_6t
Xbit_r469_c21 bl[21] br[21] wl[469] vdd gnd cell_6t
Xbit_r470_c21 bl[21] br[21] wl[470] vdd gnd cell_6t
Xbit_r471_c21 bl[21] br[21] wl[471] vdd gnd cell_6t
Xbit_r472_c21 bl[21] br[21] wl[472] vdd gnd cell_6t
Xbit_r473_c21 bl[21] br[21] wl[473] vdd gnd cell_6t
Xbit_r474_c21 bl[21] br[21] wl[474] vdd gnd cell_6t
Xbit_r475_c21 bl[21] br[21] wl[475] vdd gnd cell_6t
Xbit_r476_c21 bl[21] br[21] wl[476] vdd gnd cell_6t
Xbit_r477_c21 bl[21] br[21] wl[477] vdd gnd cell_6t
Xbit_r478_c21 bl[21] br[21] wl[478] vdd gnd cell_6t
Xbit_r479_c21 bl[21] br[21] wl[479] vdd gnd cell_6t
Xbit_r480_c21 bl[21] br[21] wl[480] vdd gnd cell_6t
Xbit_r481_c21 bl[21] br[21] wl[481] vdd gnd cell_6t
Xbit_r482_c21 bl[21] br[21] wl[482] vdd gnd cell_6t
Xbit_r483_c21 bl[21] br[21] wl[483] vdd gnd cell_6t
Xbit_r484_c21 bl[21] br[21] wl[484] vdd gnd cell_6t
Xbit_r485_c21 bl[21] br[21] wl[485] vdd gnd cell_6t
Xbit_r486_c21 bl[21] br[21] wl[486] vdd gnd cell_6t
Xbit_r487_c21 bl[21] br[21] wl[487] vdd gnd cell_6t
Xbit_r488_c21 bl[21] br[21] wl[488] vdd gnd cell_6t
Xbit_r489_c21 bl[21] br[21] wl[489] vdd gnd cell_6t
Xbit_r490_c21 bl[21] br[21] wl[490] vdd gnd cell_6t
Xbit_r491_c21 bl[21] br[21] wl[491] vdd gnd cell_6t
Xbit_r492_c21 bl[21] br[21] wl[492] vdd gnd cell_6t
Xbit_r493_c21 bl[21] br[21] wl[493] vdd gnd cell_6t
Xbit_r494_c21 bl[21] br[21] wl[494] vdd gnd cell_6t
Xbit_r495_c21 bl[21] br[21] wl[495] vdd gnd cell_6t
Xbit_r496_c21 bl[21] br[21] wl[496] vdd gnd cell_6t
Xbit_r497_c21 bl[21] br[21] wl[497] vdd gnd cell_6t
Xbit_r498_c21 bl[21] br[21] wl[498] vdd gnd cell_6t
Xbit_r499_c21 bl[21] br[21] wl[499] vdd gnd cell_6t
Xbit_r500_c21 bl[21] br[21] wl[500] vdd gnd cell_6t
Xbit_r501_c21 bl[21] br[21] wl[501] vdd gnd cell_6t
Xbit_r502_c21 bl[21] br[21] wl[502] vdd gnd cell_6t
Xbit_r503_c21 bl[21] br[21] wl[503] vdd gnd cell_6t
Xbit_r504_c21 bl[21] br[21] wl[504] vdd gnd cell_6t
Xbit_r505_c21 bl[21] br[21] wl[505] vdd gnd cell_6t
Xbit_r506_c21 bl[21] br[21] wl[506] vdd gnd cell_6t
Xbit_r507_c21 bl[21] br[21] wl[507] vdd gnd cell_6t
Xbit_r508_c21 bl[21] br[21] wl[508] vdd gnd cell_6t
Xbit_r509_c21 bl[21] br[21] wl[509] vdd gnd cell_6t
Xbit_r510_c21 bl[21] br[21] wl[510] vdd gnd cell_6t
Xbit_r511_c21 bl[21] br[21] wl[511] vdd gnd cell_6t
Xbit_r0_c22 bl[22] br[22] wl[0] vdd gnd cell_6t
Xbit_r1_c22 bl[22] br[22] wl[1] vdd gnd cell_6t
Xbit_r2_c22 bl[22] br[22] wl[2] vdd gnd cell_6t
Xbit_r3_c22 bl[22] br[22] wl[3] vdd gnd cell_6t
Xbit_r4_c22 bl[22] br[22] wl[4] vdd gnd cell_6t
Xbit_r5_c22 bl[22] br[22] wl[5] vdd gnd cell_6t
Xbit_r6_c22 bl[22] br[22] wl[6] vdd gnd cell_6t
Xbit_r7_c22 bl[22] br[22] wl[7] vdd gnd cell_6t
Xbit_r8_c22 bl[22] br[22] wl[8] vdd gnd cell_6t
Xbit_r9_c22 bl[22] br[22] wl[9] vdd gnd cell_6t
Xbit_r10_c22 bl[22] br[22] wl[10] vdd gnd cell_6t
Xbit_r11_c22 bl[22] br[22] wl[11] vdd gnd cell_6t
Xbit_r12_c22 bl[22] br[22] wl[12] vdd gnd cell_6t
Xbit_r13_c22 bl[22] br[22] wl[13] vdd gnd cell_6t
Xbit_r14_c22 bl[22] br[22] wl[14] vdd gnd cell_6t
Xbit_r15_c22 bl[22] br[22] wl[15] vdd gnd cell_6t
Xbit_r16_c22 bl[22] br[22] wl[16] vdd gnd cell_6t
Xbit_r17_c22 bl[22] br[22] wl[17] vdd gnd cell_6t
Xbit_r18_c22 bl[22] br[22] wl[18] vdd gnd cell_6t
Xbit_r19_c22 bl[22] br[22] wl[19] vdd gnd cell_6t
Xbit_r20_c22 bl[22] br[22] wl[20] vdd gnd cell_6t
Xbit_r21_c22 bl[22] br[22] wl[21] vdd gnd cell_6t
Xbit_r22_c22 bl[22] br[22] wl[22] vdd gnd cell_6t
Xbit_r23_c22 bl[22] br[22] wl[23] vdd gnd cell_6t
Xbit_r24_c22 bl[22] br[22] wl[24] vdd gnd cell_6t
Xbit_r25_c22 bl[22] br[22] wl[25] vdd gnd cell_6t
Xbit_r26_c22 bl[22] br[22] wl[26] vdd gnd cell_6t
Xbit_r27_c22 bl[22] br[22] wl[27] vdd gnd cell_6t
Xbit_r28_c22 bl[22] br[22] wl[28] vdd gnd cell_6t
Xbit_r29_c22 bl[22] br[22] wl[29] vdd gnd cell_6t
Xbit_r30_c22 bl[22] br[22] wl[30] vdd gnd cell_6t
Xbit_r31_c22 bl[22] br[22] wl[31] vdd gnd cell_6t
Xbit_r32_c22 bl[22] br[22] wl[32] vdd gnd cell_6t
Xbit_r33_c22 bl[22] br[22] wl[33] vdd gnd cell_6t
Xbit_r34_c22 bl[22] br[22] wl[34] vdd gnd cell_6t
Xbit_r35_c22 bl[22] br[22] wl[35] vdd gnd cell_6t
Xbit_r36_c22 bl[22] br[22] wl[36] vdd gnd cell_6t
Xbit_r37_c22 bl[22] br[22] wl[37] vdd gnd cell_6t
Xbit_r38_c22 bl[22] br[22] wl[38] vdd gnd cell_6t
Xbit_r39_c22 bl[22] br[22] wl[39] vdd gnd cell_6t
Xbit_r40_c22 bl[22] br[22] wl[40] vdd gnd cell_6t
Xbit_r41_c22 bl[22] br[22] wl[41] vdd gnd cell_6t
Xbit_r42_c22 bl[22] br[22] wl[42] vdd gnd cell_6t
Xbit_r43_c22 bl[22] br[22] wl[43] vdd gnd cell_6t
Xbit_r44_c22 bl[22] br[22] wl[44] vdd gnd cell_6t
Xbit_r45_c22 bl[22] br[22] wl[45] vdd gnd cell_6t
Xbit_r46_c22 bl[22] br[22] wl[46] vdd gnd cell_6t
Xbit_r47_c22 bl[22] br[22] wl[47] vdd gnd cell_6t
Xbit_r48_c22 bl[22] br[22] wl[48] vdd gnd cell_6t
Xbit_r49_c22 bl[22] br[22] wl[49] vdd gnd cell_6t
Xbit_r50_c22 bl[22] br[22] wl[50] vdd gnd cell_6t
Xbit_r51_c22 bl[22] br[22] wl[51] vdd gnd cell_6t
Xbit_r52_c22 bl[22] br[22] wl[52] vdd gnd cell_6t
Xbit_r53_c22 bl[22] br[22] wl[53] vdd gnd cell_6t
Xbit_r54_c22 bl[22] br[22] wl[54] vdd gnd cell_6t
Xbit_r55_c22 bl[22] br[22] wl[55] vdd gnd cell_6t
Xbit_r56_c22 bl[22] br[22] wl[56] vdd gnd cell_6t
Xbit_r57_c22 bl[22] br[22] wl[57] vdd gnd cell_6t
Xbit_r58_c22 bl[22] br[22] wl[58] vdd gnd cell_6t
Xbit_r59_c22 bl[22] br[22] wl[59] vdd gnd cell_6t
Xbit_r60_c22 bl[22] br[22] wl[60] vdd gnd cell_6t
Xbit_r61_c22 bl[22] br[22] wl[61] vdd gnd cell_6t
Xbit_r62_c22 bl[22] br[22] wl[62] vdd gnd cell_6t
Xbit_r63_c22 bl[22] br[22] wl[63] vdd gnd cell_6t
Xbit_r64_c22 bl[22] br[22] wl[64] vdd gnd cell_6t
Xbit_r65_c22 bl[22] br[22] wl[65] vdd gnd cell_6t
Xbit_r66_c22 bl[22] br[22] wl[66] vdd gnd cell_6t
Xbit_r67_c22 bl[22] br[22] wl[67] vdd gnd cell_6t
Xbit_r68_c22 bl[22] br[22] wl[68] vdd gnd cell_6t
Xbit_r69_c22 bl[22] br[22] wl[69] vdd gnd cell_6t
Xbit_r70_c22 bl[22] br[22] wl[70] vdd gnd cell_6t
Xbit_r71_c22 bl[22] br[22] wl[71] vdd gnd cell_6t
Xbit_r72_c22 bl[22] br[22] wl[72] vdd gnd cell_6t
Xbit_r73_c22 bl[22] br[22] wl[73] vdd gnd cell_6t
Xbit_r74_c22 bl[22] br[22] wl[74] vdd gnd cell_6t
Xbit_r75_c22 bl[22] br[22] wl[75] vdd gnd cell_6t
Xbit_r76_c22 bl[22] br[22] wl[76] vdd gnd cell_6t
Xbit_r77_c22 bl[22] br[22] wl[77] vdd gnd cell_6t
Xbit_r78_c22 bl[22] br[22] wl[78] vdd gnd cell_6t
Xbit_r79_c22 bl[22] br[22] wl[79] vdd gnd cell_6t
Xbit_r80_c22 bl[22] br[22] wl[80] vdd gnd cell_6t
Xbit_r81_c22 bl[22] br[22] wl[81] vdd gnd cell_6t
Xbit_r82_c22 bl[22] br[22] wl[82] vdd gnd cell_6t
Xbit_r83_c22 bl[22] br[22] wl[83] vdd gnd cell_6t
Xbit_r84_c22 bl[22] br[22] wl[84] vdd gnd cell_6t
Xbit_r85_c22 bl[22] br[22] wl[85] vdd gnd cell_6t
Xbit_r86_c22 bl[22] br[22] wl[86] vdd gnd cell_6t
Xbit_r87_c22 bl[22] br[22] wl[87] vdd gnd cell_6t
Xbit_r88_c22 bl[22] br[22] wl[88] vdd gnd cell_6t
Xbit_r89_c22 bl[22] br[22] wl[89] vdd gnd cell_6t
Xbit_r90_c22 bl[22] br[22] wl[90] vdd gnd cell_6t
Xbit_r91_c22 bl[22] br[22] wl[91] vdd gnd cell_6t
Xbit_r92_c22 bl[22] br[22] wl[92] vdd gnd cell_6t
Xbit_r93_c22 bl[22] br[22] wl[93] vdd gnd cell_6t
Xbit_r94_c22 bl[22] br[22] wl[94] vdd gnd cell_6t
Xbit_r95_c22 bl[22] br[22] wl[95] vdd gnd cell_6t
Xbit_r96_c22 bl[22] br[22] wl[96] vdd gnd cell_6t
Xbit_r97_c22 bl[22] br[22] wl[97] vdd gnd cell_6t
Xbit_r98_c22 bl[22] br[22] wl[98] vdd gnd cell_6t
Xbit_r99_c22 bl[22] br[22] wl[99] vdd gnd cell_6t
Xbit_r100_c22 bl[22] br[22] wl[100] vdd gnd cell_6t
Xbit_r101_c22 bl[22] br[22] wl[101] vdd gnd cell_6t
Xbit_r102_c22 bl[22] br[22] wl[102] vdd gnd cell_6t
Xbit_r103_c22 bl[22] br[22] wl[103] vdd gnd cell_6t
Xbit_r104_c22 bl[22] br[22] wl[104] vdd gnd cell_6t
Xbit_r105_c22 bl[22] br[22] wl[105] vdd gnd cell_6t
Xbit_r106_c22 bl[22] br[22] wl[106] vdd gnd cell_6t
Xbit_r107_c22 bl[22] br[22] wl[107] vdd gnd cell_6t
Xbit_r108_c22 bl[22] br[22] wl[108] vdd gnd cell_6t
Xbit_r109_c22 bl[22] br[22] wl[109] vdd gnd cell_6t
Xbit_r110_c22 bl[22] br[22] wl[110] vdd gnd cell_6t
Xbit_r111_c22 bl[22] br[22] wl[111] vdd gnd cell_6t
Xbit_r112_c22 bl[22] br[22] wl[112] vdd gnd cell_6t
Xbit_r113_c22 bl[22] br[22] wl[113] vdd gnd cell_6t
Xbit_r114_c22 bl[22] br[22] wl[114] vdd gnd cell_6t
Xbit_r115_c22 bl[22] br[22] wl[115] vdd gnd cell_6t
Xbit_r116_c22 bl[22] br[22] wl[116] vdd gnd cell_6t
Xbit_r117_c22 bl[22] br[22] wl[117] vdd gnd cell_6t
Xbit_r118_c22 bl[22] br[22] wl[118] vdd gnd cell_6t
Xbit_r119_c22 bl[22] br[22] wl[119] vdd gnd cell_6t
Xbit_r120_c22 bl[22] br[22] wl[120] vdd gnd cell_6t
Xbit_r121_c22 bl[22] br[22] wl[121] vdd gnd cell_6t
Xbit_r122_c22 bl[22] br[22] wl[122] vdd gnd cell_6t
Xbit_r123_c22 bl[22] br[22] wl[123] vdd gnd cell_6t
Xbit_r124_c22 bl[22] br[22] wl[124] vdd gnd cell_6t
Xbit_r125_c22 bl[22] br[22] wl[125] vdd gnd cell_6t
Xbit_r126_c22 bl[22] br[22] wl[126] vdd gnd cell_6t
Xbit_r127_c22 bl[22] br[22] wl[127] vdd gnd cell_6t
Xbit_r128_c22 bl[22] br[22] wl[128] vdd gnd cell_6t
Xbit_r129_c22 bl[22] br[22] wl[129] vdd gnd cell_6t
Xbit_r130_c22 bl[22] br[22] wl[130] vdd gnd cell_6t
Xbit_r131_c22 bl[22] br[22] wl[131] vdd gnd cell_6t
Xbit_r132_c22 bl[22] br[22] wl[132] vdd gnd cell_6t
Xbit_r133_c22 bl[22] br[22] wl[133] vdd gnd cell_6t
Xbit_r134_c22 bl[22] br[22] wl[134] vdd gnd cell_6t
Xbit_r135_c22 bl[22] br[22] wl[135] vdd gnd cell_6t
Xbit_r136_c22 bl[22] br[22] wl[136] vdd gnd cell_6t
Xbit_r137_c22 bl[22] br[22] wl[137] vdd gnd cell_6t
Xbit_r138_c22 bl[22] br[22] wl[138] vdd gnd cell_6t
Xbit_r139_c22 bl[22] br[22] wl[139] vdd gnd cell_6t
Xbit_r140_c22 bl[22] br[22] wl[140] vdd gnd cell_6t
Xbit_r141_c22 bl[22] br[22] wl[141] vdd gnd cell_6t
Xbit_r142_c22 bl[22] br[22] wl[142] vdd gnd cell_6t
Xbit_r143_c22 bl[22] br[22] wl[143] vdd gnd cell_6t
Xbit_r144_c22 bl[22] br[22] wl[144] vdd gnd cell_6t
Xbit_r145_c22 bl[22] br[22] wl[145] vdd gnd cell_6t
Xbit_r146_c22 bl[22] br[22] wl[146] vdd gnd cell_6t
Xbit_r147_c22 bl[22] br[22] wl[147] vdd gnd cell_6t
Xbit_r148_c22 bl[22] br[22] wl[148] vdd gnd cell_6t
Xbit_r149_c22 bl[22] br[22] wl[149] vdd gnd cell_6t
Xbit_r150_c22 bl[22] br[22] wl[150] vdd gnd cell_6t
Xbit_r151_c22 bl[22] br[22] wl[151] vdd gnd cell_6t
Xbit_r152_c22 bl[22] br[22] wl[152] vdd gnd cell_6t
Xbit_r153_c22 bl[22] br[22] wl[153] vdd gnd cell_6t
Xbit_r154_c22 bl[22] br[22] wl[154] vdd gnd cell_6t
Xbit_r155_c22 bl[22] br[22] wl[155] vdd gnd cell_6t
Xbit_r156_c22 bl[22] br[22] wl[156] vdd gnd cell_6t
Xbit_r157_c22 bl[22] br[22] wl[157] vdd gnd cell_6t
Xbit_r158_c22 bl[22] br[22] wl[158] vdd gnd cell_6t
Xbit_r159_c22 bl[22] br[22] wl[159] vdd gnd cell_6t
Xbit_r160_c22 bl[22] br[22] wl[160] vdd gnd cell_6t
Xbit_r161_c22 bl[22] br[22] wl[161] vdd gnd cell_6t
Xbit_r162_c22 bl[22] br[22] wl[162] vdd gnd cell_6t
Xbit_r163_c22 bl[22] br[22] wl[163] vdd gnd cell_6t
Xbit_r164_c22 bl[22] br[22] wl[164] vdd gnd cell_6t
Xbit_r165_c22 bl[22] br[22] wl[165] vdd gnd cell_6t
Xbit_r166_c22 bl[22] br[22] wl[166] vdd gnd cell_6t
Xbit_r167_c22 bl[22] br[22] wl[167] vdd gnd cell_6t
Xbit_r168_c22 bl[22] br[22] wl[168] vdd gnd cell_6t
Xbit_r169_c22 bl[22] br[22] wl[169] vdd gnd cell_6t
Xbit_r170_c22 bl[22] br[22] wl[170] vdd gnd cell_6t
Xbit_r171_c22 bl[22] br[22] wl[171] vdd gnd cell_6t
Xbit_r172_c22 bl[22] br[22] wl[172] vdd gnd cell_6t
Xbit_r173_c22 bl[22] br[22] wl[173] vdd gnd cell_6t
Xbit_r174_c22 bl[22] br[22] wl[174] vdd gnd cell_6t
Xbit_r175_c22 bl[22] br[22] wl[175] vdd gnd cell_6t
Xbit_r176_c22 bl[22] br[22] wl[176] vdd gnd cell_6t
Xbit_r177_c22 bl[22] br[22] wl[177] vdd gnd cell_6t
Xbit_r178_c22 bl[22] br[22] wl[178] vdd gnd cell_6t
Xbit_r179_c22 bl[22] br[22] wl[179] vdd gnd cell_6t
Xbit_r180_c22 bl[22] br[22] wl[180] vdd gnd cell_6t
Xbit_r181_c22 bl[22] br[22] wl[181] vdd gnd cell_6t
Xbit_r182_c22 bl[22] br[22] wl[182] vdd gnd cell_6t
Xbit_r183_c22 bl[22] br[22] wl[183] vdd gnd cell_6t
Xbit_r184_c22 bl[22] br[22] wl[184] vdd gnd cell_6t
Xbit_r185_c22 bl[22] br[22] wl[185] vdd gnd cell_6t
Xbit_r186_c22 bl[22] br[22] wl[186] vdd gnd cell_6t
Xbit_r187_c22 bl[22] br[22] wl[187] vdd gnd cell_6t
Xbit_r188_c22 bl[22] br[22] wl[188] vdd gnd cell_6t
Xbit_r189_c22 bl[22] br[22] wl[189] vdd gnd cell_6t
Xbit_r190_c22 bl[22] br[22] wl[190] vdd gnd cell_6t
Xbit_r191_c22 bl[22] br[22] wl[191] vdd gnd cell_6t
Xbit_r192_c22 bl[22] br[22] wl[192] vdd gnd cell_6t
Xbit_r193_c22 bl[22] br[22] wl[193] vdd gnd cell_6t
Xbit_r194_c22 bl[22] br[22] wl[194] vdd gnd cell_6t
Xbit_r195_c22 bl[22] br[22] wl[195] vdd gnd cell_6t
Xbit_r196_c22 bl[22] br[22] wl[196] vdd gnd cell_6t
Xbit_r197_c22 bl[22] br[22] wl[197] vdd gnd cell_6t
Xbit_r198_c22 bl[22] br[22] wl[198] vdd gnd cell_6t
Xbit_r199_c22 bl[22] br[22] wl[199] vdd gnd cell_6t
Xbit_r200_c22 bl[22] br[22] wl[200] vdd gnd cell_6t
Xbit_r201_c22 bl[22] br[22] wl[201] vdd gnd cell_6t
Xbit_r202_c22 bl[22] br[22] wl[202] vdd gnd cell_6t
Xbit_r203_c22 bl[22] br[22] wl[203] vdd gnd cell_6t
Xbit_r204_c22 bl[22] br[22] wl[204] vdd gnd cell_6t
Xbit_r205_c22 bl[22] br[22] wl[205] vdd gnd cell_6t
Xbit_r206_c22 bl[22] br[22] wl[206] vdd gnd cell_6t
Xbit_r207_c22 bl[22] br[22] wl[207] vdd gnd cell_6t
Xbit_r208_c22 bl[22] br[22] wl[208] vdd gnd cell_6t
Xbit_r209_c22 bl[22] br[22] wl[209] vdd gnd cell_6t
Xbit_r210_c22 bl[22] br[22] wl[210] vdd gnd cell_6t
Xbit_r211_c22 bl[22] br[22] wl[211] vdd gnd cell_6t
Xbit_r212_c22 bl[22] br[22] wl[212] vdd gnd cell_6t
Xbit_r213_c22 bl[22] br[22] wl[213] vdd gnd cell_6t
Xbit_r214_c22 bl[22] br[22] wl[214] vdd gnd cell_6t
Xbit_r215_c22 bl[22] br[22] wl[215] vdd gnd cell_6t
Xbit_r216_c22 bl[22] br[22] wl[216] vdd gnd cell_6t
Xbit_r217_c22 bl[22] br[22] wl[217] vdd gnd cell_6t
Xbit_r218_c22 bl[22] br[22] wl[218] vdd gnd cell_6t
Xbit_r219_c22 bl[22] br[22] wl[219] vdd gnd cell_6t
Xbit_r220_c22 bl[22] br[22] wl[220] vdd gnd cell_6t
Xbit_r221_c22 bl[22] br[22] wl[221] vdd gnd cell_6t
Xbit_r222_c22 bl[22] br[22] wl[222] vdd gnd cell_6t
Xbit_r223_c22 bl[22] br[22] wl[223] vdd gnd cell_6t
Xbit_r224_c22 bl[22] br[22] wl[224] vdd gnd cell_6t
Xbit_r225_c22 bl[22] br[22] wl[225] vdd gnd cell_6t
Xbit_r226_c22 bl[22] br[22] wl[226] vdd gnd cell_6t
Xbit_r227_c22 bl[22] br[22] wl[227] vdd gnd cell_6t
Xbit_r228_c22 bl[22] br[22] wl[228] vdd gnd cell_6t
Xbit_r229_c22 bl[22] br[22] wl[229] vdd gnd cell_6t
Xbit_r230_c22 bl[22] br[22] wl[230] vdd gnd cell_6t
Xbit_r231_c22 bl[22] br[22] wl[231] vdd gnd cell_6t
Xbit_r232_c22 bl[22] br[22] wl[232] vdd gnd cell_6t
Xbit_r233_c22 bl[22] br[22] wl[233] vdd gnd cell_6t
Xbit_r234_c22 bl[22] br[22] wl[234] vdd gnd cell_6t
Xbit_r235_c22 bl[22] br[22] wl[235] vdd gnd cell_6t
Xbit_r236_c22 bl[22] br[22] wl[236] vdd gnd cell_6t
Xbit_r237_c22 bl[22] br[22] wl[237] vdd gnd cell_6t
Xbit_r238_c22 bl[22] br[22] wl[238] vdd gnd cell_6t
Xbit_r239_c22 bl[22] br[22] wl[239] vdd gnd cell_6t
Xbit_r240_c22 bl[22] br[22] wl[240] vdd gnd cell_6t
Xbit_r241_c22 bl[22] br[22] wl[241] vdd gnd cell_6t
Xbit_r242_c22 bl[22] br[22] wl[242] vdd gnd cell_6t
Xbit_r243_c22 bl[22] br[22] wl[243] vdd gnd cell_6t
Xbit_r244_c22 bl[22] br[22] wl[244] vdd gnd cell_6t
Xbit_r245_c22 bl[22] br[22] wl[245] vdd gnd cell_6t
Xbit_r246_c22 bl[22] br[22] wl[246] vdd gnd cell_6t
Xbit_r247_c22 bl[22] br[22] wl[247] vdd gnd cell_6t
Xbit_r248_c22 bl[22] br[22] wl[248] vdd gnd cell_6t
Xbit_r249_c22 bl[22] br[22] wl[249] vdd gnd cell_6t
Xbit_r250_c22 bl[22] br[22] wl[250] vdd gnd cell_6t
Xbit_r251_c22 bl[22] br[22] wl[251] vdd gnd cell_6t
Xbit_r252_c22 bl[22] br[22] wl[252] vdd gnd cell_6t
Xbit_r253_c22 bl[22] br[22] wl[253] vdd gnd cell_6t
Xbit_r254_c22 bl[22] br[22] wl[254] vdd gnd cell_6t
Xbit_r255_c22 bl[22] br[22] wl[255] vdd gnd cell_6t
Xbit_r256_c22 bl[22] br[22] wl[256] vdd gnd cell_6t
Xbit_r257_c22 bl[22] br[22] wl[257] vdd gnd cell_6t
Xbit_r258_c22 bl[22] br[22] wl[258] vdd gnd cell_6t
Xbit_r259_c22 bl[22] br[22] wl[259] vdd gnd cell_6t
Xbit_r260_c22 bl[22] br[22] wl[260] vdd gnd cell_6t
Xbit_r261_c22 bl[22] br[22] wl[261] vdd gnd cell_6t
Xbit_r262_c22 bl[22] br[22] wl[262] vdd gnd cell_6t
Xbit_r263_c22 bl[22] br[22] wl[263] vdd gnd cell_6t
Xbit_r264_c22 bl[22] br[22] wl[264] vdd gnd cell_6t
Xbit_r265_c22 bl[22] br[22] wl[265] vdd gnd cell_6t
Xbit_r266_c22 bl[22] br[22] wl[266] vdd gnd cell_6t
Xbit_r267_c22 bl[22] br[22] wl[267] vdd gnd cell_6t
Xbit_r268_c22 bl[22] br[22] wl[268] vdd gnd cell_6t
Xbit_r269_c22 bl[22] br[22] wl[269] vdd gnd cell_6t
Xbit_r270_c22 bl[22] br[22] wl[270] vdd gnd cell_6t
Xbit_r271_c22 bl[22] br[22] wl[271] vdd gnd cell_6t
Xbit_r272_c22 bl[22] br[22] wl[272] vdd gnd cell_6t
Xbit_r273_c22 bl[22] br[22] wl[273] vdd gnd cell_6t
Xbit_r274_c22 bl[22] br[22] wl[274] vdd gnd cell_6t
Xbit_r275_c22 bl[22] br[22] wl[275] vdd gnd cell_6t
Xbit_r276_c22 bl[22] br[22] wl[276] vdd gnd cell_6t
Xbit_r277_c22 bl[22] br[22] wl[277] vdd gnd cell_6t
Xbit_r278_c22 bl[22] br[22] wl[278] vdd gnd cell_6t
Xbit_r279_c22 bl[22] br[22] wl[279] vdd gnd cell_6t
Xbit_r280_c22 bl[22] br[22] wl[280] vdd gnd cell_6t
Xbit_r281_c22 bl[22] br[22] wl[281] vdd gnd cell_6t
Xbit_r282_c22 bl[22] br[22] wl[282] vdd gnd cell_6t
Xbit_r283_c22 bl[22] br[22] wl[283] vdd gnd cell_6t
Xbit_r284_c22 bl[22] br[22] wl[284] vdd gnd cell_6t
Xbit_r285_c22 bl[22] br[22] wl[285] vdd gnd cell_6t
Xbit_r286_c22 bl[22] br[22] wl[286] vdd gnd cell_6t
Xbit_r287_c22 bl[22] br[22] wl[287] vdd gnd cell_6t
Xbit_r288_c22 bl[22] br[22] wl[288] vdd gnd cell_6t
Xbit_r289_c22 bl[22] br[22] wl[289] vdd gnd cell_6t
Xbit_r290_c22 bl[22] br[22] wl[290] vdd gnd cell_6t
Xbit_r291_c22 bl[22] br[22] wl[291] vdd gnd cell_6t
Xbit_r292_c22 bl[22] br[22] wl[292] vdd gnd cell_6t
Xbit_r293_c22 bl[22] br[22] wl[293] vdd gnd cell_6t
Xbit_r294_c22 bl[22] br[22] wl[294] vdd gnd cell_6t
Xbit_r295_c22 bl[22] br[22] wl[295] vdd gnd cell_6t
Xbit_r296_c22 bl[22] br[22] wl[296] vdd gnd cell_6t
Xbit_r297_c22 bl[22] br[22] wl[297] vdd gnd cell_6t
Xbit_r298_c22 bl[22] br[22] wl[298] vdd gnd cell_6t
Xbit_r299_c22 bl[22] br[22] wl[299] vdd gnd cell_6t
Xbit_r300_c22 bl[22] br[22] wl[300] vdd gnd cell_6t
Xbit_r301_c22 bl[22] br[22] wl[301] vdd gnd cell_6t
Xbit_r302_c22 bl[22] br[22] wl[302] vdd gnd cell_6t
Xbit_r303_c22 bl[22] br[22] wl[303] vdd gnd cell_6t
Xbit_r304_c22 bl[22] br[22] wl[304] vdd gnd cell_6t
Xbit_r305_c22 bl[22] br[22] wl[305] vdd gnd cell_6t
Xbit_r306_c22 bl[22] br[22] wl[306] vdd gnd cell_6t
Xbit_r307_c22 bl[22] br[22] wl[307] vdd gnd cell_6t
Xbit_r308_c22 bl[22] br[22] wl[308] vdd gnd cell_6t
Xbit_r309_c22 bl[22] br[22] wl[309] vdd gnd cell_6t
Xbit_r310_c22 bl[22] br[22] wl[310] vdd gnd cell_6t
Xbit_r311_c22 bl[22] br[22] wl[311] vdd gnd cell_6t
Xbit_r312_c22 bl[22] br[22] wl[312] vdd gnd cell_6t
Xbit_r313_c22 bl[22] br[22] wl[313] vdd gnd cell_6t
Xbit_r314_c22 bl[22] br[22] wl[314] vdd gnd cell_6t
Xbit_r315_c22 bl[22] br[22] wl[315] vdd gnd cell_6t
Xbit_r316_c22 bl[22] br[22] wl[316] vdd gnd cell_6t
Xbit_r317_c22 bl[22] br[22] wl[317] vdd gnd cell_6t
Xbit_r318_c22 bl[22] br[22] wl[318] vdd gnd cell_6t
Xbit_r319_c22 bl[22] br[22] wl[319] vdd gnd cell_6t
Xbit_r320_c22 bl[22] br[22] wl[320] vdd gnd cell_6t
Xbit_r321_c22 bl[22] br[22] wl[321] vdd gnd cell_6t
Xbit_r322_c22 bl[22] br[22] wl[322] vdd gnd cell_6t
Xbit_r323_c22 bl[22] br[22] wl[323] vdd gnd cell_6t
Xbit_r324_c22 bl[22] br[22] wl[324] vdd gnd cell_6t
Xbit_r325_c22 bl[22] br[22] wl[325] vdd gnd cell_6t
Xbit_r326_c22 bl[22] br[22] wl[326] vdd gnd cell_6t
Xbit_r327_c22 bl[22] br[22] wl[327] vdd gnd cell_6t
Xbit_r328_c22 bl[22] br[22] wl[328] vdd gnd cell_6t
Xbit_r329_c22 bl[22] br[22] wl[329] vdd gnd cell_6t
Xbit_r330_c22 bl[22] br[22] wl[330] vdd gnd cell_6t
Xbit_r331_c22 bl[22] br[22] wl[331] vdd gnd cell_6t
Xbit_r332_c22 bl[22] br[22] wl[332] vdd gnd cell_6t
Xbit_r333_c22 bl[22] br[22] wl[333] vdd gnd cell_6t
Xbit_r334_c22 bl[22] br[22] wl[334] vdd gnd cell_6t
Xbit_r335_c22 bl[22] br[22] wl[335] vdd gnd cell_6t
Xbit_r336_c22 bl[22] br[22] wl[336] vdd gnd cell_6t
Xbit_r337_c22 bl[22] br[22] wl[337] vdd gnd cell_6t
Xbit_r338_c22 bl[22] br[22] wl[338] vdd gnd cell_6t
Xbit_r339_c22 bl[22] br[22] wl[339] vdd gnd cell_6t
Xbit_r340_c22 bl[22] br[22] wl[340] vdd gnd cell_6t
Xbit_r341_c22 bl[22] br[22] wl[341] vdd gnd cell_6t
Xbit_r342_c22 bl[22] br[22] wl[342] vdd gnd cell_6t
Xbit_r343_c22 bl[22] br[22] wl[343] vdd gnd cell_6t
Xbit_r344_c22 bl[22] br[22] wl[344] vdd gnd cell_6t
Xbit_r345_c22 bl[22] br[22] wl[345] vdd gnd cell_6t
Xbit_r346_c22 bl[22] br[22] wl[346] vdd gnd cell_6t
Xbit_r347_c22 bl[22] br[22] wl[347] vdd gnd cell_6t
Xbit_r348_c22 bl[22] br[22] wl[348] vdd gnd cell_6t
Xbit_r349_c22 bl[22] br[22] wl[349] vdd gnd cell_6t
Xbit_r350_c22 bl[22] br[22] wl[350] vdd gnd cell_6t
Xbit_r351_c22 bl[22] br[22] wl[351] vdd gnd cell_6t
Xbit_r352_c22 bl[22] br[22] wl[352] vdd gnd cell_6t
Xbit_r353_c22 bl[22] br[22] wl[353] vdd gnd cell_6t
Xbit_r354_c22 bl[22] br[22] wl[354] vdd gnd cell_6t
Xbit_r355_c22 bl[22] br[22] wl[355] vdd gnd cell_6t
Xbit_r356_c22 bl[22] br[22] wl[356] vdd gnd cell_6t
Xbit_r357_c22 bl[22] br[22] wl[357] vdd gnd cell_6t
Xbit_r358_c22 bl[22] br[22] wl[358] vdd gnd cell_6t
Xbit_r359_c22 bl[22] br[22] wl[359] vdd gnd cell_6t
Xbit_r360_c22 bl[22] br[22] wl[360] vdd gnd cell_6t
Xbit_r361_c22 bl[22] br[22] wl[361] vdd gnd cell_6t
Xbit_r362_c22 bl[22] br[22] wl[362] vdd gnd cell_6t
Xbit_r363_c22 bl[22] br[22] wl[363] vdd gnd cell_6t
Xbit_r364_c22 bl[22] br[22] wl[364] vdd gnd cell_6t
Xbit_r365_c22 bl[22] br[22] wl[365] vdd gnd cell_6t
Xbit_r366_c22 bl[22] br[22] wl[366] vdd gnd cell_6t
Xbit_r367_c22 bl[22] br[22] wl[367] vdd gnd cell_6t
Xbit_r368_c22 bl[22] br[22] wl[368] vdd gnd cell_6t
Xbit_r369_c22 bl[22] br[22] wl[369] vdd gnd cell_6t
Xbit_r370_c22 bl[22] br[22] wl[370] vdd gnd cell_6t
Xbit_r371_c22 bl[22] br[22] wl[371] vdd gnd cell_6t
Xbit_r372_c22 bl[22] br[22] wl[372] vdd gnd cell_6t
Xbit_r373_c22 bl[22] br[22] wl[373] vdd gnd cell_6t
Xbit_r374_c22 bl[22] br[22] wl[374] vdd gnd cell_6t
Xbit_r375_c22 bl[22] br[22] wl[375] vdd gnd cell_6t
Xbit_r376_c22 bl[22] br[22] wl[376] vdd gnd cell_6t
Xbit_r377_c22 bl[22] br[22] wl[377] vdd gnd cell_6t
Xbit_r378_c22 bl[22] br[22] wl[378] vdd gnd cell_6t
Xbit_r379_c22 bl[22] br[22] wl[379] vdd gnd cell_6t
Xbit_r380_c22 bl[22] br[22] wl[380] vdd gnd cell_6t
Xbit_r381_c22 bl[22] br[22] wl[381] vdd gnd cell_6t
Xbit_r382_c22 bl[22] br[22] wl[382] vdd gnd cell_6t
Xbit_r383_c22 bl[22] br[22] wl[383] vdd gnd cell_6t
Xbit_r384_c22 bl[22] br[22] wl[384] vdd gnd cell_6t
Xbit_r385_c22 bl[22] br[22] wl[385] vdd gnd cell_6t
Xbit_r386_c22 bl[22] br[22] wl[386] vdd gnd cell_6t
Xbit_r387_c22 bl[22] br[22] wl[387] vdd gnd cell_6t
Xbit_r388_c22 bl[22] br[22] wl[388] vdd gnd cell_6t
Xbit_r389_c22 bl[22] br[22] wl[389] vdd gnd cell_6t
Xbit_r390_c22 bl[22] br[22] wl[390] vdd gnd cell_6t
Xbit_r391_c22 bl[22] br[22] wl[391] vdd gnd cell_6t
Xbit_r392_c22 bl[22] br[22] wl[392] vdd gnd cell_6t
Xbit_r393_c22 bl[22] br[22] wl[393] vdd gnd cell_6t
Xbit_r394_c22 bl[22] br[22] wl[394] vdd gnd cell_6t
Xbit_r395_c22 bl[22] br[22] wl[395] vdd gnd cell_6t
Xbit_r396_c22 bl[22] br[22] wl[396] vdd gnd cell_6t
Xbit_r397_c22 bl[22] br[22] wl[397] vdd gnd cell_6t
Xbit_r398_c22 bl[22] br[22] wl[398] vdd gnd cell_6t
Xbit_r399_c22 bl[22] br[22] wl[399] vdd gnd cell_6t
Xbit_r400_c22 bl[22] br[22] wl[400] vdd gnd cell_6t
Xbit_r401_c22 bl[22] br[22] wl[401] vdd gnd cell_6t
Xbit_r402_c22 bl[22] br[22] wl[402] vdd gnd cell_6t
Xbit_r403_c22 bl[22] br[22] wl[403] vdd gnd cell_6t
Xbit_r404_c22 bl[22] br[22] wl[404] vdd gnd cell_6t
Xbit_r405_c22 bl[22] br[22] wl[405] vdd gnd cell_6t
Xbit_r406_c22 bl[22] br[22] wl[406] vdd gnd cell_6t
Xbit_r407_c22 bl[22] br[22] wl[407] vdd gnd cell_6t
Xbit_r408_c22 bl[22] br[22] wl[408] vdd gnd cell_6t
Xbit_r409_c22 bl[22] br[22] wl[409] vdd gnd cell_6t
Xbit_r410_c22 bl[22] br[22] wl[410] vdd gnd cell_6t
Xbit_r411_c22 bl[22] br[22] wl[411] vdd gnd cell_6t
Xbit_r412_c22 bl[22] br[22] wl[412] vdd gnd cell_6t
Xbit_r413_c22 bl[22] br[22] wl[413] vdd gnd cell_6t
Xbit_r414_c22 bl[22] br[22] wl[414] vdd gnd cell_6t
Xbit_r415_c22 bl[22] br[22] wl[415] vdd gnd cell_6t
Xbit_r416_c22 bl[22] br[22] wl[416] vdd gnd cell_6t
Xbit_r417_c22 bl[22] br[22] wl[417] vdd gnd cell_6t
Xbit_r418_c22 bl[22] br[22] wl[418] vdd gnd cell_6t
Xbit_r419_c22 bl[22] br[22] wl[419] vdd gnd cell_6t
Xbit_r420_c22 bl[22] br[22] wl[420] vdd gnd cell_6t
Xbit_r421_c22 bl[22] br[22] wl[421] vdd gnd cell_6t
Xbit_r422_c22 bl[22] br[22] wl[422] vdd gnd cell_6t
Xbit_r423_c22 bl[22] br[22] wl[423] vdd gnd cell_6t
Xbit_r424_c22 bl[22] br[22] wl[424] vdd gnd cell_6t
Xbit_r425_c22 bl[22] br[22] wl[425] vdd gnd cell_6t
Xbit_r426_c22 bl[22] br[22] wl[426] vdd gnd cell_6t
Xbit_r427_c22 bl[22] br[22] wl[427] vdd gnd cell_6t
Xbit_r428_c22 bl[22] br[22] wl[428] vdd gnd cell_6t
Xbit_r429_c22 bl[22] br[22] wl[429] vdd gnd cell_6t
Xbit_r430_c22 bl[22] br[22] wl[430] vdd gnd cell_6t
Xbit_r431_c22 bl[22] br[22] wl[431] vdd gnd cell_6t
Xbit_r432_c22 bl[22] br[22] wl[432] vdd gnd cell_6t
Xbit_r433_c22 bl[22] br[22] wl[433] vdd gnd cell_6t
Xbit_r434_c22 bl[22] br[22] wl[434] vdd gnd cell_6t
Xbit_r435_c22 bl[22] br[22] wl[435] vdd gnd cell_6t
Xbit_r436_c22 bl[22] br[22] wl[436] vdd gnd cell_6t
Xbit_r437_c22 bl[22] br[22] wl[437] vdd gnd cell_6t
Xbit_r438_c22 bl[22] br[22] wl[438] vdd gnd cell_6t
Xbit_r439_c22 bl[22] br[22] wl[439] vdd gnd cell_6t
Xbit_r440_c22 bl[22] br[22] wl[440] vdd gnd cell_6t
Xbit_r441_c22 bl[22] br[22] wl[441] vdd gnd cell_6t
Xbit_r442_c22 bl[22] br[22] wl[442] vdd gnd cell_6t
Xbit_r443_c22 bl[22] br[22] wl[443] vdd gnd cell_6t
Xbit_r444_c22 bl[22] br[22] wl[444] vdd gnd cell_6t
Xbit_r445_c22 bl[22] br[22] wl[445] vdd gnd cell_6t
Xbit_r446_c22 bl[22] br[22] wl[446] vdd gnd cell_6t
Xbit_r447_c22 bl[22] br[22] wl[447] vdd gnd cell_6t
Xbit_r448_c22 bl[22] br[22] wl[448] vdd gnd cell_6t
Xbit_r449_c22 bl[22] br[22] wl[449] vdd gnd cell_6t
Xbit_r450_c22 bl[22] br[22] wl[450] vdd gnd cell_6t
Xbit_r451_c22 bl[22] br[22] wl[451] vdd gnd cell_6t
Xbit_r452_c22 bl[22] br[22] wl[452] vdd gnd cell_6t
Xbit_r453_c22 bl[22] br[22] wl[453] vdd gnd cell_6t
Xbit_r454_c22 bl[22] br[22] wl[454] vdd gnd cell_6t
Xbit_r455_c22 bl[22] br[22] wl[455] vdd gnd cell_6t
Xbit_r456_c22 bl[22] br[22] wl[456] vdd gnd cell_6t
Xbit_r457_c22 bl[22] br[22] wl[457] vdd gnd cell_6t
Xbit_r458_c22 bl[22] br[22] wl[458] vdd gnd cell_6t
Xbit_r459_c22 bl[22] br[22] wl[459] vdd gnd cell_6t
Xbit_r460_c22 bl[22] br[22] wl[460] vdd gnd cell_6t
Xbit_r461_c22 bl[22] br[22] wl[461] vdd gnd cell_6t
Xbit_r462_c22 bl[22] br[22] wl[462] vdd gnd cell_6t
Xbit_r463_c22 bl[22] br[22] wl[463] vdd gnd cell_6t
Xbit_r464_c22 bl[22] br[22] wl[464] vdd gnd cell_6t
Xbit_r465_c22 bl[22] br[22] wl[465] vdd gnd cell_6t
Xbit_r466_c22 bl[22] br[22] wl[466] vdd gnd cell_6t
Xbit_r467_c22 bl[22] br[22] wl[467] vdd gnd cell_6t
Xbit_r468_c22 bl[22] br[22] wl[468] vdd gnd cell_6t
Xbit_r469_c22 bl[22] br[22] wl[469] vdd gnd cell_6t
Xbit_r470_c22 bl[22] br[22] wl[470] vdd gnd cell_6t
Xbit_r471_c22 bl[22] br[22] wl[471] vdd gnd cell_6t
Xbit_r472_c22 bl[22] br[22] wl[472] vdd gnd cell_6t
Xbit_r473_c22 bl[22] br[22] wl[473] vdd gnd cell_6t
Xbit_r474_c22 bl[22] br[22] wl[474] vdd gnd cell_6t
Xbit_r475_c22 bl[22] br[22] wl[475] vdd gnd cell_6t
Xbit_r476_c22 bl[22] br[22] wl[476] vdd gnd cell_6t
Xbit_r477_c22 bl[22] br[22] wl[477] vdd gnd cell_6t
Xbit_r478_c22 bl[22] br[22] wl[478] vdd gnd cell_6t
Xbit_r479_c22 bl[22] br[22] wl[479] vdd gnd cell_6t
Xbit_r480_c22 bl[22] br[22] wl[480] vdd gnd cell_6t
Xbit_r481_c22 bl[22] br[22] wl[481] vdd gnd cell_6t
Xbit_r482_c22 bl[22] br[22] wl[482] vdd gnd cell_6t
Xbit_r483_c22 bl[22] br[22] wl[483] vdd gnd cell_6t
Xbit_r484_c22 bl[22] br[22] wl[484] vdd gnd cell_6t
Xbit_r485_c22 bl[22] br[22] wl[485] vdd gnd cell_6t
Xbit_r486_c22 bl[22] br[22] wl[486] vdd gnd cell_6t
Xbit_r487_c22 bl[22] br[22] wl[487] vdd gnd cell_6t
Xbit_r488_c22 bl[22] br[22] wl[488] vdd gnd cell_6t
Xbit_r489_c22 bl[22] br[22] wl[489] vdd gnd cell_6t
Xbit_r490_c22 bl[22] br[22] wl[490] vdd gnd cell_6t
Xbit_r491_c22 bl[22] br[22] wl[491] vdd gnd cell_6t
Xbit_r492_c22 bl[22] br[22] wl[492] vdd gnd cell_6t
Xbit_r493_c22 bl[22] br[22] wl[493] vdd gnd cell_6t
Xbit_r494_c22 bl[22] br[22] wl[494] vdd gnd cell_6t
Xbit_r495_c22 bl[22] br[22] wl[495] vdd gnd cell_6t
Xbit_r496_c22 bl[22] br[22] wl[496] vdd gnd cell_6t
Xbit_r497_c22 bl[22] br[22] wl[497] vdd gnd cell_6t
Xbit_r498_c22 bl[22] br[22] wl[498] vdd gnd cell_6t
Xbit_r499_c22 bl[22] br[22] wl[499] vdd gnd cell_6t
Xbit_r500_c22 bl[22] br[22] wl[500] vdd gnd cell_6t
Xbit_r501_c22 bl[22] br[22] wl[501] vdd gnd cell_6t
Xbit_r502_c22 bl[22] br[22] wl[502] vdd gnd cell_6t
Xbit_r503_c22 bl[22] br[22] wl[503] vdd gnd cell_6t
Xbit_r504_c22 bl[22] br[22] wl[504] vdd gnd cell_6t
Xbit_r505_c22 bl[22] br[22] wl[505] vdd gnd cell_6t
Xbit_r506_c22 bl[22] br[22] wl[506] vdd gnd cell_6t
Xbit_r507_c22 bl[22] br[22] wl[507] vdd gnd cell_6t
Xbit_r508_c22 bl[22] br[22] wl[508] vdd gnd cell_6t
Xbit_r509_c22 bl[22] br[22] wl[509] vdd gnd cell_6t
Xbit_r510_c22 bl[22] br[22] wl[510] vdd gnd cell_6t
Xbit_r511_c22 bl[22] br[22] wl[511] vdd gnd cell_6t
Xbit_r0_c23 bl[23] br[23] wl[0] vdd gnd cell_6t
Xbit_r1_c23 bl[23] br[23] wl[1] vdd gnd cell_6t
Xbit_r2_c23 bl[23] br[23] wl[2] vdd gnd cell_6t
Xbit_r3_c23 bl[23] br[23] wl[3] vdd gnd cell_6t
Xbit_r4_c23 bl[23] br[23] wl[4] vdd gnd cell_6t
Xbit_r5_c23 bl[23] br[23] wl[5] vdd gnd cell_6t
Xbit_r6_c23 bl[23] br[23] wl[6] vdd gnd cell_6t
Xbit_r7_c23 bl[23] br[23] wl[7] vdd gnd cell_6t
Xbit_r8_c23 bl[23] br[23] wl[8] vdd gnd cell_6t
Xbit_r9_c23 bl[23] br[23] wl[9] vdd gnd cell_6t
Xbit_r10_c23 bl[23] br[23] wl[10] vdd gnd cell_6t
Xbit_r11_c23 bl[23] br[23] wl[11] vdd gnd cell_6t
Xbit_r12_c23 bl[23] br[23] wl[12] vdd gnd cell_6t
Xbit_r13_c23 bl[23] br[23] wl[13] vdd gnd cell_6t
Xbit_r14_c23 bl[23] br[23] wl[14] vdd gnd cell_6t
Xbit_r15_c23 bl[23] br[23] wl[15] vdd gnd cell_6t
Xbit_r16_c23 bl[23] br[23] wl[16] vdd gnd cell_6t
Xbit_r17_c23 bl[23] br[23] wl[17] vdd gnd cell_6t
Xbit_r18_c23 bl[23] br[23] wl[18] vdd gnd cell_6t
Xbit_r19_c23 bl[23] br[23] wl[19] vdd gnd cell_6t
Xbit_r20_c23 bl[23] br[23] wl[20] vdd gnd cell_6t
Xbit_r21_c23 bl[23] br[23] wl[21] vdd gnd cell_6t
Xbit_r22_c23 bl[23] br[23] wl[22] vdd gnd cell_6t
Xbit_r23_c23 bl[23] br[23] wl[23] vdd gnd cell_6t
Xbit_r24_c23 bl[23] br[23] wl[24] vdd gnd cell_6t
Xbit_r25_c23 bl[23] br[23] wl[25] vdd gnd cell_6t
Xbit_r26_c23 bl[23] br[23] wl[26] vdd gnd cell_6t
Xbit_r27_c23 bl[23] br[23] wl[27] vdd gnd cell_6t
Xbit_r28_c23 bl[23] br[23] wl[28] vdd gnd cell_6t
Xbit_r29_c23 bl[23] br[23] wl[29] vdd gnd cell_6t
Xbit_r30_c23 bl[23] br[23] wl[30] vdd gnd cell_6t
Xbit_r31_c23 bl[23] br[23] wl[31] vdd gnd cell_6t
Xbit_r32_c23 bl[23] br[23] wl[32] vdd gnd cell_6t
Xbit_r33_c23 bl[23] br[23] wl[33] vdd gnd cell_6t
Xbit_r34_c23 bl[23] br[23] wl[34] vdd gnd cell_6t
Xbit_r35_c23 bl[23] br[23] wl[35] vdd gnd cell_6t
Xbit_r36_c23 bl[23] br[23] wl[36] vdd gnd cell_6t
Xbit_r37_c23 bl[23] br[23] wl[37] vdd gnd cell_6t
Xbit_r38_c23 bl[23] br[23] wl[38] vdd gnd cell_6t
Xbit_r39_c23 bl[23] br[23] wl[39] vdd gnd cell_6t
Xbit_r40_c23 bl[23] br[23] wl[40] vdd gnd cell_6t
Xbit_r41_c23 bl[23] br[23] wl[41] vdd gnd cell_6t
Xbit_r42_c23 bl[23] br[23] wl[42] vdd gnd cell_6t
Xbit_r43_c23 bl[23] br[23] wl[43] vdd gnd cell_6t
Xbit_r44_c23 bl[23] br[23] wl[44] vdd gnd cell_6t
Xbit_r45_c23 bl[23] br[23] wl[45] vdd gnd cell_6t
Xbit_r46_c23 bl[23] br[23] wl[46] vdd gnd cell_6t
Xbit_r47_c23 bl[23] br[23] wl[47] vdd gnd cell_6t
Xbit_r48_c23 bl[23] br[23] wl[48] vdd gnd cell_6t
Xbit_r49_c23 bl[23] br[23] wl[49] vdd gnd cell_6t
Xbit_r50_c23 bl[23] br[23] wl[50] vdd gnd cell_6t
Xbit_r51_c23 bl[23] br[23] wl[51] vdd gnd cell_6t
Xbit_r52_c23 bl[23] br[23] wl[52] vdd gnd cell_6t
Xbit_r53_c23 bl[23] br[23] wl[53] vdd gnd cell_6t
Xbit_r54_c23 bl[23] br[23] wl[54] vdd gnd cell_6t
Xbit_r55_c23 bl[23] br[23] wl[55] vdd gnd cell_6t
Xbit_r56_c23 bl[23] br[23] wl[56] vdd gnd cell_6t
Xbit_r57_c23 bl[23] br[23] wl[57] vdd gnd cell_6t
Xbit_r58_c23 bl[23] br[23] wl[58] vdd gnd cell_6t
Xbit_r59_c23 bl[23] br[23] wl[59] vdd gnd cell_6t
Xbit_r60_c23 bl[23] br[23] wl[60] vdd gnd cell_6t
Xbit_r61_c23 bl[23] br[23] wl[61] vdd gnd cell_6t
Xbit_r62_c23 bl[23] br[23] wl[62] vdd gnd cell_6t
Xbit_r63_c23 bl[23] br[23] wl[63] vdd gnd cell_6t
Xbit_r64_c23 bl[23] br[23] wl[64] vdd gnd cell_6t
Xbit_r65_c23 bl[23] br[23] wl[65] vdd gnd cell_6t
Xbit_r66_c23 bl[23] br[23] wl[66] vdd gnd cell_6t
Xbit_r67_c23 bl[23] br[23] wl[67] vdd gnd cell_6t
Xbit_r68_c23 bl[23] br[23] wl[68] vdd gnd cell_6t
Xbit_r69_c23 bl[23] br[23] wl[69] vdd gnd cell_6t
Xbit_r70_c23 bl[23] br[23] wl[70] vdd gnd cell_6t
Xbit_r71_c23 bl[23] br[23] wl[71] vdd gnd cell_6t
Xbit_r72_c23 bl[23] br[23] wl[72] vdd gnd cell_6t
Xbit_r73_c23 bl[23] br[23] wl[73] vdd gnd cell_6t
Xbit_r74_c23 bl[23] br[23] wl[74] vdd gnd cell_6t
Xbit_r75_c23 bl[23] br[23] wl[75] vdd gnd cell_6t
Xbit_r76_c23 bl[23] br[23] wl[76] vdd gnd cell_6t
Xbit_r77_c23 bl[23] br[23] wl[77] vdd gnd cell_6t
Xbit_r78_c23 bl[23] br[23] wl[78] vdd gnd cell_6t
Xbit_r79_c23 bl[23] br[23] wl[79] vdd gnd cell_6t
Xbit_r80_c23 bl[23] br[23] wl[80] vdd gnd cell_6t
Xbit_r81_c23 bl[23] br[23] wl[81] vdd gnd cell_6t
Xbit_r82_c23 bl[23] br[23] wl[82] vdd gnd cell_6t
Xbit_r83_c23 bl[23] br[23] wl[83] vdd gnd cell_6t
Xbit_r84_c23 bl[23] br[23] wl[84] vdd gnd cell_6t
Xbit_r85_c23 bl[23] br[23] wl[85] vdd gnd cell_6t
Xbit_r86_c23 bl[23] br[23] wl[86] vdd gnd cell_6t
Xbit_r87_c23 bl[23] br[23] wl[87] vdd gnd cell_6t
Xbit_r88_c23 bl[23] br[23] wl[88] vdd gnd cell_6t
Xbit_r89_c23 bl[23] br[23] wl[89] vdd gnd cell_6t
Xbit_r90_c23 bl[23] br[23] wl[90] vdd gnd cell_6t
Xbit_r91_c23 bl[23] br[23] wl[91] vdd gnd cell_6t
Xbit_r92_c23 bl[23] br[23] wl[92] vdd gnd cell_6t
Xbit_r93_c23 bl[23] br[23] wl[93] vdd gnd cell_6t
Xbit_r94_c23 bl[23] br[23] wl[94] vdd gnd cell_6t
Xbit_r95_c23 bl[23] br[23] wl[95] vdd gnd cell_6t
Xbit_r96_c23 bl[23] br[23] wl[96] vdd gnd cell_6t
Xbit_r97_c23 bl[23] br[23] wl[97] vdd gnd cell_6t
Xbit_r98_c23 bl[23] br[23] wl[98] vdd gnd cell_6t
Xbit_r99_c23 bl[23] br[23] wl[99] vdd gnd cell_6t
Xbit_r100_c23 bl[23] br[23] wl[100] vdd gnd cell_6t
Xbit_r101_c23 bl[23] br[23] wl[101] vdd gnd cell_6t
Xbit_r102_c23 bl[23] br[23] wl[102] vdd gnd cell_6t
Xbit_r103_c23 bl[23] br[23] wl[103] vdd gnd cell_6t
Xbit_r104_c23 bl[23] br[23] wl[104] vdd gnd cell_6t
Xbit_r105_c23 bl[23] br[23] wl[105] vdd gnd cell_6t
Xbit_r106_c23 bl[23] br[23] wl[106] vdd gnd cell_6t
Xbit_r107_c23 bl[23] br[23] wl[107] vdd gnd cell_6t
Xbit_r108_c23 bl[23] br[23] wl[108] vdd gnd cell_6t
Xbit_r109_c23 bl[23] br[23] wl[109] vdd gnd cell_6t
Xbit_r110_c23 bl[23] br[23] wl[110] vdd gnd cell_6t
Xbit_r111_c23 bl[23] br[23] wl[111] vdd gnd cell_6t
Xbit_r112_c23 bl[23] br[23] wl[112] vdd gnd cell_6t
Xbit_r113_c23 bl[23] br[23] wl[113] vdd gnd cell_6t
Xbit_r114_c23 bl[23] br[23] wl[114] vdd gnd cell_6t
Xbit_r115_c23 bl[23] br[23] wl[115] vdd gnd cell_6t
Xbit_r116_c23 bl[23] br[23] wl[116] vdd gnd cell_6t
Xbit_r117_c23 bl[23] br[23] wl[117] vdd gnd cell_6t
Xbit_r118_c23 bl[23] br[23] wl[118] vdd gnd cell_6t
Xbit_r119_c23 bl[23] br[23] wl[119] vdd gnd cell_6t
Xbit_r120_c23 bl[23] br[23] wl[120] vdd gnd cell_6t
Xbit_r121_c23 bl[23] br[23] wl[121] vdd gnd cell_6t
Xbit_r122_c23 bl[23] br[23] wl[122] vdd gnd cell_6t
Xbit_r123_c23 bl[23] br[23] wl[123] vdd gnd cell_6t
Xbit_r124_c23 bl[23] br[23] wl[124] vdd gnd cell_6t
Xbit_r125_c23 bl[23] br[23] wl[125] vdd gnd cell_6t
Xbit_r126_c23 bl[23] br[23] wl[126] vdd gnd cell_6t
Xbit_r127_c23 bl[23] br[23] wl[127] vdd gnd cell_6t
Xbit_r128_c23 bl[23] br[23] wl[128] vdd gnd cell_6t
Xbit_r129_c23 bl[23] br[23] wl[129] vdd gnd cell_6t
Xbit_r130_c23 bl[23] br[23] wl[130] vdd gnd cell_6t
Xbit_r131_c23 bl[23] br[23] wl[131] vdd gnd cell_6t
Xbit_r132_c23 bl[23] br[23] wl[132] vdd gnd cell_6t
Xbit_r133_c23 bl[23] br[23] wl[133] vdd gnd cell_6t
Xbit_r134_c23 bl[23] br[23] wl[134] vdd gnd cell_6t
Xbit_r135_c23 bl[23] br[23] wl[135] vdd gnd cell_6t
Xbit_r136_c23 bl[23] br[23] wl[136] vdd gnd cell_6t
Xbit_r137_c23 bl[23] br[23] wl[137] vdd gnd cell_6t
Xbit_r138_c23 bl[23] br[23] wl[138] vdd gnd cell_6t
Xbit_r139_c23 bl[23] br[23] wl[139] vdd gnd cell_6t
Xbit_r140_c23 bl[23] br[23] wl[140] vdd gnd cell_6t
Xbit_r141_c23 bl[23] br[23] wl[141] vdd gnd cell_6t
Xbit_r142_c23 bl[23] br[23] wl[142] vdd gnd cell_6t
Xbit_r143_c23 bl[23] br[23] wl[143] vdd gnd cell_6t
Xbit_r144_c23 bl[23] br[23] wl[144] vdd gnd cell_6t
Xbit_r145_c23 bl[23] br[23] wl[145] vdd gnd cell_6t
Xbit_r146_c23 bl[23] br[23] wl[146] vdd gnd cell_6t
Xbit_r147_c23 bl[23] br[23] wl[147] vdd gnd cell_6t
Xbit_r148_c23 bl[23] br[23] wl[148] vdd gnd cell_6t
Xbit_r149_c23 bl[23] br[23] wl[149] vdd gnd cell_6t
Xbit_r150_c23 bl[23] br[23] wl[150] vdd gnd cell_6t
Xbit_r151_c23 bl[23] br[23] wl[151] vdd gnd cell_6t
Xbit_r152_c23 bl[23] br[23] wl[152] vdd gnd cell_6t
Xbit_r153_c23 bl[23] br[23] wl[153] vdd gnd cell_6t
Xbit_r154_c23 bl[23] br[23] wl[154] vdd gnd cell_6t
Xbit_r155_c23 bl[23] br[23] wl[155] vdd gnd cell_6t
Xbit_r156_c23 bl[23] br[23] wl[156] vdd gnd cell_6t
Xbit_r157_c23 bl[23] br[23] wl[157] vdd gnd cell_6t
Xbit_r158_c23 bl[23] br[23] wl[158] vdd gnd cell_6t
Xbit_r159_c23 bl[23] br[23] wl[159] vdd gnd cell_6t
Xbit_r160_c23 bl[23] br[23] wl[160] vdd gnd cell_6t
Xbit_r161_c23 bl[23] br[23] wl[161] vdd gnd cell_6t
Xbit_r162_c23 bl[23] br[23] wl[162] vdd gnd cell_6t
Xbit_r163_c23 bl[23] br[23] wl[163] vdd gnd cell_6t
Xbit_r164_c23 bl[23] br[23] wl[164] vdd gnd cell_6t
Xbit_r165_c23 bl[23] br[23] wl[165] vdd gnd cell_6t
Xbit_r166_c23 bl[23] br[23] wl[166] vdd gnd cell_6t
Xbit_r167_c23 bl[23] br[23] wl[167] vdd gnd cell_6t
Xbit_r168_c23 bl[23] br[23] wl[168] vdd gnd cell_6t
Xbit_r169_c23 bl[23] br[23] wl[169] vdd gnd cell_6t
Xbit_r170_c23 bl[23] br[23] wl[170] vdd gnd cell_6t
Xbit_r171_c23 bl[23] br[23] wl[171] vdd gnd cell_6t
Xbit_r172_c23 bl[23] br[23] wl[172] vdd gnd cell_6t
Xbit_r173_c23 bl[23] br[23] wl[173] vdd gnd cell_6t
Xbit_r174_c23 bl[23] br[23] wl[174] vdd gnd cell_6t
Xbit_r175_c23 bl[23] br[23] wl[175] vdd gnd cell_6t
Xbit_r176_c23 bl[23] br[23] wl[176] vdd gnd cell_6t
Xbit_r177_c23 bl[23] br[23] wl[177] vdd gnd cell_6t
Xbit_r178_c23 bl[23] br[23] wl[178] vdd gnd cell_6t
Xbit_r179_c23 bl[23] br[23] wl[179] vdd gnd cell_6t
Xbit_r180_c23 bl[23] br[23] wl[180] vdd gnd cell_6t
Xbit_r181_c23 bl[23] br[23] wl[181] vdd gnd cell_6t
Xbit_r182_c23 bl[23] br[23] wl[182] vdd gnd cell_6t
Xbit_r183_c23 bl[23] br[23] wl[183] vdd gnd cell_6t
Xbit_r184_c23 bl[23] br[23] wl[184] vdd gnd cell_6t
Xbit_r185_c23 bl[23] br[23] wl[185] vdd gnd cell_6t
Xbit_r186_c23 bl[23] br[23] wl[186] vdd gnd cell_6t
Xbit_r187_c23 bl[23] br[23] wl[187] vdd gnd cell_6t
Xbit_r188_c23 bl[23] br[23] wl[188] vdd gnd cell_6t
Xbit_r189_c23 bl[23] br[23] wl[189] vdd gnd cell_6t
Xbit_r190_c23 bl[23] br[23] wl[190] vdd gnd cell_6t
Xbit_r191_c23 bl[23] br[23] wl[191] vdd gnd cell_6t
Xbit_r192_c23 bl[23] br[23] wl[192] vdd gnd cell_6t
Xbit_r193_c23 bl[23] br[23] wl[193] vdd gnd cell_6t
Xbit_r194_c23 bl[23] br[23] wl[194] vdd gnd cell_6t
Xbit_r195_c23 bl[23] br[23] wl[195] vdd gnd cell_6t
Xbit_r196_c23 bl[23] br[23] wl[196] vdd gnd cell_6t
Xbit_r197_c23 bl[23] br[23] wl[197] vdd gnd cell_6t
Xbit_r198_c23 bl[23] br[23] wl[198] vdd gnd cell_6t
Xbit_r199_c23 bl[23] br[23] wl[199] vdd gnd cell_6t
Xbit_r200_c23 bl[23] br[23] wl[200] vdd gnd cell_6t
Xbit_r201_c23 bl[23] br[23] wl[201] vdd gnd cell_6t
Xbit_r202_c23 bl[23] br[23] wl[202] vdd gnd cell_6t
Xbit_r203_c23 bl[23] br[23] wl[203] vdd gnd cell_6t
Xbit_r204_c23 bl[23] br[23] wl[204] vdd gnd cell_6t
Xbit_r205_c23 bl[23] br[23] wl[205] vdd gnd cell_6t
Xbit_r206_c23 bl[23] br[23] wl[206] vdd gnd cell_6t
Xbit_r207_c23 bl[23] br[23] wl[207] vdd gnd cell_6t
Xbit_r208_c23 bl[23] br[23] wl[208] vdd gnd cell_6t
Xbit_r209_c23 bl[23] br[23] wl[209] vdd gnd cell_6t
Xbit_r210_c23 bl[23] br[23] wl[210] vdd gnd cell_6t
Xbit_r211_c23 bl[23] br[23] wl[211] vdd gnd cell_6t
Xbit_r212_c23 bl[23] br[23] wl[212] vdd gnd cell_6t
Xbit_r213_c23 bl[23] br[23] wl[213] vdd gnd cell_6t
Xbit_r214_c23 bl[23] br[23] wl[214] vdd gnd cell_6t
Xbit_r215_c23 bl[23] br[23] wl[215] vdd gnd cell_6t
Xbit_r216_c23 bl[23] br[23] wl[216] vdd gnd cell_6t
Xbit_r217_c23 bl[23] br[23] wl[217] vdd gnd cell_6t
Xbit_r218_c23 bl[23] br[23] wl[218] vdd gnd cell_6t
Xbit_r219_c23 bl[23] br[23] wl[219] vdd gnd cell_6t
Xbit_r220_c23 bl[23] br[23] wl[220] vdd gnd cell_6t
Xbit_r221_c23 bl[23] br[23] wl[221] vdd gnd cell_6t
Xbit_r222_c23 bl[23] br[23] wl[222] vdd gnd cell_6t
Xbit_r223_c23 bl[23] br[23] wl[223] vdd gnd cell_6t
Xbit_r224_c23 bl[23] br[23] wl[224] vdd gnd cell_6t
Xbit_r225_c23 bl[23] br[23] wl[225] vdd gnd cell_6t
Xbit_r226_c23 bl[23] br[23] wl[226] vdd gnd cell_6t
Xbit_r227_c23 bl[23] br[23] wl[227] vdd gnd cell_6t
Xbit_r228_c23 bl[23] br[23] wl[228] vdd gnd cell_6t
Xbit_r229_c23 bl[23] br[23] wl[229] vdd gnd cell_6t
Xbit_r230_c23 bl[23] br[23] wl[230] vdd gnd cell_6t
Xbit_r231_c23 bl[23] br[23] wl[231] vdd gnd cell_6t
Xbit_r232_c23 bl[23] br[23] wl[232] vdd gnd cell_6t
Xbit_r233_c23 bl[23] br[23] wl[233] vdd gnd cell_6t
Xbit_r234_c23 bl[23] br[23] wl[234] vdd gnd cell_6t
Xbit_r235_c23 bl[23] br[23] wl[235] vdd gnd cell_6t
Xbit_r236_c23 bl[23] br[23] wl[236] vdd gnd cell_6t
Xbit_r237_c23 bl[23] br[23] wl[237] vdd gnd cell_6t
Xbit_r238_c23 bl[23] br[23] wl[238] vdd gnd cell_6t
Xbit_r239_c23 bl[23] br[23] wl[239] vdd gnd cell_6t
Xbit_r240_c23 bl[23] br[23] wl[240] vdd gnd cell_6t
Xbit_r241_c23 bl[23] br[23] wl[241] vdd gnd cell_6t
Xbit_r242_c23 bl[23] br[23] wl[242] vdd gnd cell_6t
Xbit_r243_c23 bl[23] br[23] wl[243] vdd gnd cell_6t
Xbit_r244_c23 bl[23] br[23] wl[244] vdd gnd cell_6t
Xbit_r245_c23 bl[23] br[23] wl[245] vdd gnd cell_6t
Xbit_r246_c23 bl[23] br[23] wl[246] vdd gnd cell_6t
Xbit_r247_c23 bl[23] br[23] wl[247] vdd gnd cell_6t
Xbit_r248_c23 bl[23] br[23] wl[248] vdd gnd cell_6t
Xbit_r249_c23 bl[23] br[23] wl[249] vdd gnd cell_6t
Xbit_r250_c23 bl[23] br[23] wl[250] vdd gnd cell_6t
Xbit_r251_c23 bl[23] br[23] wl[251] vdd gnd cell_6t
Xbit_r252_c23 bl[23] br[23] wl[252] vdd gnd cell_6t
Xbit_r253_c23 bl[23] br[23] wl[253] vdd gnd cell_6t
Xbit_r254_c23 bl[23] br[23] wl[254] vdd gnd cell_6t
Xbit_r255_c23 bl[23] br[23] wl[255] vdd gnd cell_6t
Xbit_r256_c23 bl[23] br[23] wl[256] vdd gnd cell_6t
Xbit_r257_c23 bl[23] br[23] wl[257] vdd gnd cell_6t
Xbit_r258_c23 bl[23] br[23] wl[258] vdd gnd cell_6t
Xbit_r259_c23 bl[23] br[23] wl[259] vdd gnd cell_6t
Xbit_r260_c23 bl[23] br[23] wl[260] vdd gnd cell_6t
Xbit_r261_c23 bl[23] br[23] wl[261] vdd gnd cell_6t
Xbit_r262_c23 bl[23] br[23] wl[262] vdd gnd cell_6t
Xbit_r263_c23 bl[23] br[23] wl[263] vdd gnd cell_6t
Xbit_r264_c23 bl[23] br[23] wl[264] vdd gnd cell_6t
Xbit_r265_c23 bl[23] br[23] wl[265] vdd gnd cell_6t
Xbit_r266_c23 bl[23] br[23] wl[266] vdd gnd cell_6t
Xbit_r267_c23 bl[23] br[23] wl[267] vdd gnd cell_6t
Xbit_r268_c23 bl[23] br[23] wl[268] vdd gnd cell_6t
Xbit_r269_c23 bl[23] br[23] wl[269] vdd gnd cell_6t
Xbit_r270_c23 bl[23] br[23] wl[270] vdd gnd cell_6t
Xbit_r271_c23 bl[23] br[23] wl[271] vdd gnd cell_6t
Xbit_r272_c23 bl[23] br[23] wl[272] vdd gnd cell_6t
Xbit_r273_c23 bl[23] br[23] wl[273] vdd gnd cell_6t
Xbit_r274_c23 bl[23] br[23] wl[274] vdd gnd cell_6t
Xbit_r275_c23 bl[23] br[23] wl[275] vdd gnd cell_6t
Xbit_r276_c23 bl[23] br[23] wl[276] vdd gnd cell_6t
Xbit_r277_c23 bl[23] br[23] wl[277] vdd gnd cell_6t
Xbit_r278_c23 bl[23] br[23] wl[278] vdd gnd cell_6t
Xbit_r279_c23 bl[23] br[23] wl[279] vdd gnd cell_6t
Xbit_r280_c23 bl[23] br[23] wl[280] vdd gnd cell_6t
Xbit_r281_c23 bl[23] br[23] wl[281] vdd gnd cell_6t
Xbit_r282_c23 bl[23] br[23] wl[282] vdd gnd cell_6t
Xbit_r283_c23 bl[23] br[23] wl[283] vdd gnd cell_6t
Xbit_r284_c23 bl[23] br[23] wl[284] vdd gnd cell_6t
Xbit_r285_c23 bl[23] br[23] wl[285] vdd gnd cell_6t
Xbit_r286_c23 bl[23] br[23] wl[286] vdd gnd cell_6t
Xbit_r287_c23 bl[23] br[23] wl[287] vdd gnd cell_6t
Xbit_r288_c23 bl[23] br[23] wl[288] vdd gnd cell_6t
Xbit_r289_c23 bl[23] br[23] wl[289] vdd gnd cell_6t
Xbit_r290_c23 bl[23] br[23] wl[290] vdd gnd cell_6t
Xbit_r291_c23 bl[23] br[23] wl[291] vdd gnd cell_6t
Xbit_r292_c23 bl[23] br[23] wl[292] vdd gnd cell_6t
Xbit_r293_c23 bl[23] br[23] wl[293] vdd gnd cell_6t
Xbit_r294_c23 bl[23] br[23] wl[294] vdd gnd cell_6t
Xbit_r295_c23 bl[23] br[23] wl[295] vdd gnd cell_6t
Xbit_r296_c23 bl[23] br[23] wl[296] vdd gnd cell_6t
Xbit_r297_c23 bl[23] br[23] wl[297] vdd gnd cell_6t
Xbit_r298_c23 bl[23] br[23] wl[298] vdd gnd cell_6t
Xbit_r299_c23 bl[23] br[23] wl[299] vdd gnd cell_6t
Xbit_r300_c23 bl[23] br[23] wl[300] vdd gnd cell_6t
Xbit_r301_c23 bl[23] br[23] wl[301] vdd gnd cell_6t
Xbit_r302_c23 bl[23] br[23] wl[302] vdd gnd cell_6t
Xbit_r303_c23 bl[23] br[23] wl[303] vdd gnd cell_6t
Xbit_r304_c23 bl[23] br[23] wl[304] vdd gnd cell_6t
Xbit_r305_c23 bl[23] br[23] wl[305] vdd gnd cell_6t
Xbit_r306_c23 bl[23] br[23] wl[306] vdd gnd cell_6t
Xbit_r307_c23 bl[23] br[23] wl[307] vdd gnd cell_6t
Xbit_r308_c23 bl[23] br[23] wl[308] vdd gnd cell_6t
Xbit_r309_c23 bl[23] br[23] wl[309] vdd gnd cell_6t
Xbit_r310_c23 bl[23] br[23] wl[310] vdd gnd cell_6t
Xbit_r311_c23 bl[23] br[23] wl[311] vdd gnd cell_6t
Xbit_r312_c23 bl[23] br[23] wl[312] vdd gnd cell_6t
Xbit_r313_c23 bl[23] br[23] wl[313] vdd gnd cell_6t
Xbit_r314_c23 bl[23] br[23] wl[314] vdd gnd cell_6t
Xbit_r315_c23 bl[23] br[23] wl[315] vdd gnd cell_6t
Xbit_r316_c23 bl[23] br[23] wl[316] vdd gnd cell_6t
Xbit_r317_c23 bl[23] br[23] wl[317] vdd gnd cell_6t
Xbit_r318_c23 bl[23] br[23] wl[318] vdd gnd cell_6t
Xbit_r319_c23 bl[23] br[23] wl[319] vdd gnd cell_6t
Xbit_r320_c23 bl[23] br[23] wl[320] vdd gnd cell_6t
Xbit_r321_c23 bl[23] br[23] wl[321] vdd gnd cell_6t
Xbit_r322_c23 bl[23] br[23] wl[322] vdd gnd cell_6t
Xbit_r323_c23 bl[23] br[23] wl[323] vdd gnd cell_6t
Xbit_r324_c23 bl[23] br[23] wl[324] vdd gnd cell_6t
Xbit_r325_c23 bl[23] br[23] wl[325] vdd gnd cell_6t
Xbit_r326_c23 bl[23] br[23] wl[326] vdd gnd cell_6t
Xbit_r327_c23 bl[23] br[23] wl[327] vdd gnd cell_6t
Xbit_r328_c23 bl[23] br[23] wl[328] vdd gnd cell_6t
Xbit_r329_c23 bl[23] br[23] wl[329] vdd gnd cell_6t
Xbit_r330_c23 bl[23] br[23] wl[330] vdd gnd cell_6t
Xbit_r331_c23 bl[23] br[23] wl[331] vdd gnd cell_6t
Xbit_r332_c23 bl[23] br[23] wl[332] vdd gnd cell_6t
Xbit_r333_c23 bl[23] br[23] wl[333] vdd gnd cell_6t
Xbit_r334_c23 bl[23] br[23] wl[334] vdd gnd cell_6t
Xbit_r335_c23 bl[23] br[23] wl[335] vdd gnd cell_6t
Xbit_r336_c23 bl[23] br[23] wl[336] vdd gnd cell_6t
Xbit_r337_c23 bl[23] br[23] wl[337] vdd gnd cell_6t
Xbit_r338_c23 bl[23] br[23] wl[338] vdd gnd cell_6t
Xbit_r339_c23 bl[23] br[23] wl[339] vdd gnd cell_6t
Xbit_r340_c23 bl[23] br[23] wl[340] vdd gnd cell_6t
Xbit_r341_c23 bl[23] br[23] wl[341] vdd gnd cell_6t
Xbit_r342_c23 bl[23] br[23] wl[342] vdd gnd cell_6t
Xbit_r343_c23 bl[23] br[23] wl[343] vdd gnd cell_6t
Xbit_r344_c23 bl[23] br[23] wl[344] vdd gnd cell_6t
Xbit_r345_c23 bl[23] br[23] wl[345] vdd gnd cell_6t
Xbit_r346_c23 bl[23] br[23] wl[346] vdd gnd cell_6t
Xbit_r347_c23 bl[23] br[23] wl[347] vdd gnd cell_6t
Xbit_r348_c23 bl[23] br[23] wl[348] vdd gnd cell_6t
Xbit_r349_c23 bl[23] br[23] wl[349] vdd gnd cell_6t
Xbit_r350_c23 bl[23] br[23] wl[350] vdd gnd cell_6t
Xbit_r351_c23 bl[23] br[23] wl[351] vdd gnd cell_6t
Xbit_r352_c23 bl[23] br[23] wl[352] vdd gnd cell_6t
Xbit_r353_c23 bl[23] br[23] wl[353] vdd gnd cell_6t
Xbit_r354_c23 bl[23] br[23] wl[354] vdd gnd cell_6t
Xbit_r355_c23 bl[23] br[23] wl[355] vdd gnd cell_6t
Xbit_r356_c23 bl[23] br[23] wl[356] vdd gnd cell_6t
Xbit_r357_c23 bl[23] br[23] wl[357] vdd gnd cell_6t
Xbit_r358_c23 bl[23] br[23] wl[358] vdd gnd cell_6t
Xbit_r359_c23 bl[23] br[23] wl[359] vdd gnd cell_6t
Xbit_r360_c23 bl[23] br[23] wl[360] vdd gnd cell_6t
Xbit_r361_c23 bl[23] br[23] wl[361] vdd gnd cell_6t
Xbit_r362_c23 bl[23] br[23] wl[362] vdd gnd cell_6t
Xbit_r363_c23 bl[23] br[23] wl[363] vdd gnd cell_6t
Xbit_r364_c23 bl[23] br[23] wl[364] vdd gnd cell_6t
Xbit_r365_c23 bl[23] br[23] wl[365] vdd gnd cell_6t
Xbit_r366_c23 bl[23] br[23] wl[366] vdd gnd cell_6t
Xbit_r367_c23 bl[23] br[23] wl[367] vdd gnd cell_6t
Xbit_r368_c23 bl[23] br[23] wl[368] vdd gnd cell_6t
Xbit_r369_c23 bl[23] br[23] wl[369] vdd gnd cell_6t
Xbit_r370_c23 bl[23] br[23] wl[370] vdd gnd cell_6t
Xbit_r371_c23 bl[23] br[23] wl[371] vdd gnd cell_6t
Xbit_r372_c23 bl[23] br[23] wl[372] vdd gnd cell_6t
Xbit_r373_c23 bl[23] br[23] wl[373] vdd gnd cell_6t
Xbit_r374_c23 bl[23] br[23] wl[374] vdd gnd cell_6t
Xbit_r375_c23 bl[23] br[23] wl[375] vdd gnd cell_6t
Xbit_r376_c23 bl[23] br[23] wl[376] vdd gnd cell_6t
Xbit_r377_c23 bl[23] br[23] wl[377] vdd gnd cell_6t
Xbit_r378_c23 bl[23] br[23] wl[378] vdd gnd cell_6t
Xbit_r379_c23 bl[23] br[23] wl[379] vdd gnd cell_6t
Xbit_r380_c23 bl[23] br[23] wl[380] vdd gnd cell_6t
Xbit_r381_c23 bl[23] br[23] wl[381] vdd gnd cell_6t
Xbit_r382_c23 bl[23] br[23] wl[382] vdd gnd cell_6t
Xbit_r383_c23 bl[23] br[23] wl[383] vdd gnd cell_6t
Xbit_r384_c23 bl[23] br[23] wl[384] vdd gnd cell_6t
Xbit_r385_c23 bl[23] br[23] wl[385] vdd gnd cell_6t
Xbit_r386_c23 bl[23] br[23] wl[386] vdd gnd cell_6t
Xbit_r387_c23 bl[23] br[23] wl[387] vdd gnd cell_6t
Xbit_r388_c23 bl[23] br[23] wl[388] vdd gnd cell_6t
Xbit_r389_c23 bl[23] br[23] wl[389] vdd gnd cell_6t
Xbit_r390_c23 bl[23] br[23] wl[390] vdd gnd cell_6t
Xbit_r391_c23 bl[23] br[23] wl[391] vdd gnd cell_6t
Xbit_r392_c23 bl[23] br[23] wl[392] vdd gnd cell_6t
Xbit_r393_c23 bl[23] br[23] wl[393] vdd gnd cell_6t
Xbit_r394_c23 bl[23] br[23] wl[394] vdd gnd cell_6t
Xbit_r395_c23 bl[23] br[23] wl[395] vdd gnd cell_6t
Xbit_r396_c23 bl[23] br[23] wl[396] vdd gnd cell_6t
Xbit_r397_c23 bl[23] br[23] wl[397] vdd gnd cell_6t
Xbit_r398_c23 bl[23] br[23] wl[398] vdd gnd cell_6t
Xbit_r399_c23 bl[23] br[23] wl[399] vdd gnd cell_6t
Xbit_r400_c23 bl[23] br[23] wl[400] vdd gnd cell_6t
Xbit_r401_c23 bl[23] br[23] wl[401] vdd gnd cell_6t
Xbit_r402_c23 bl[23] br[23] wl[402] vdd gnd cell_6t
Xbit_r403_c23 bl[23] br[23] wl[403] vdd gnd cell_6t
Xbit_r404_c23 bl[23] br[23] wl[404] vdd gnd cell_6t
Xbit_r405_c23 bl[23] br[23] wl[405] vdd gnd cell_6t
Xbit_r406_c23 bl[23] br[23] wl[406] vdd gnd cell_6t
Xbit_r407_c23 bl[23] br[23] wl[407] vdd gnd cell_6t
Xbit_r408_c23 bl[23] br[23] wl[408] vdd gnd cell_6t
Xbit_r409_c23 bl[23] br[23] wl[409] vdd gnd cell_6t
Xbit_r410_c23 bl[23] br[23] wl[410] vdd gnd cell_6t
Xbit_r411_c23 bl[23] br[23] wl[411] vdd gnd cell_6t
Xbit_r412_c23 bl[23] br[23] wl[412] vdd gnd cell_6t
Xbit_r413_c23 bl[23] br[23] wl[413] vdd gnd cell_6t
Xbit_r414_c23 bl[23] br[23] wl[414] vdd gnd cell_6t
Xbit_r415_c23 bl[23] br[23] wl[415] vdd gnd cell_6t
Xbit_r416_c23 bl[23] br[23] wl[416] vdd gnd cell_6t
Xbit_r417_c23 bl[23] br[23] wl[417] vdd gnd cell_6t
Xbit_r418_c23 bl[23] br[23] wl[418] vdd gnd cell_6t
Xbit_r419_c23 bl[23] br[23] wl[419] vdd gnd cell_6t
Xbit_r420_c23 bl[23] br[23] wl[420] vdd gnd cell_6t
Xbit_r421_c23 bl[23] br[23] wl[421] vdd gnd cell_6t
Xbit_r422_c23 bl[23] br[23] wl[422] vdd gnd cell_6t
Xbit_r423_c23 bl[23] br[23] wl[423] vdd gnd cell_6t
Xbit_r424_c23 bl[23] br[23] wl[424] vdd gnd cell_6t
Xbit_r425_c23 bl[23] br[23] wl[425] vdd gnd cell_6t
Xbit_r426_c23 bl[23] br[23] wl[426] vdd gnd cell_6t
Xbit_r427_c23 bl[23] br[23] wl[427] vdd gnd cell_6t
Xbit_r428_c23 bl[23] br[23] wl[428] vdd gnd cell_6t
Xbit_r429_c23 bl[23] br[23] wl[429] vdd gnd cell_6t
Xbit_r430_c23 bl[23] br[23] wl[430] vdd gnd cell_6t
Xbit_r431_c23 bl[23] br[23] wl[431] vdd gnd cell_6t
Xbit_r432_c23 bl[23] br[23] wl[432] vdd gnd cell_6t
Xbit_r433_c23 bl[23] br[23] wl[433] vdd gnd cell_6t
Xbit_r434_c23 bl[23] br[23] wl[434] vdd gnd cell_6t
Xbit_r435_c23 bl[23] br[23] wl[435] vdd gnd cell_6t
Xbit_r436_c23 bl[23] br[23] wl[436] vdd gnd cell_6t
Xbit_r437_c23 bl[23] br[23] wl[437] vdd gnd cell_6t
Xbit_r438_c23 bl[23] br[23] wl[438] vdd gnd cell_6t
Xbit_r439_c23 bl[23] br[23] wl[439] vdd gnd cell_6t
Xbit_r440_c23 bl[23] br[23] wl[440] vdd gnd cell_6t
Xbit_r441_c23 bl[23] br[23] wl[441] vdd gnd cell_6t
Xbit_r442_c23 bl[23] br[23] wl[442] vdd gnd cell_6t
Xbit_r443_c23 bl[23] br[23] wl[443] vdd gnd cell_6t
Xbit_r444_c23 bl[23] br[23] wl[444] vdd gnd cell_6t
Xbit_r445_c23 bl[23] br[23] wl[445] vdd gnd cell_6t
Xbit_r446_c23 bl[23] br[23] wl[446] vdd gnd cell_6t
Xbit_r447_c23 bl[23] br[23] wl[447] vdd gnd cell_6t
Xbit_r448_c23 bl[23] br[23] wl[448] vdd gnd cell_6t
Xbit_r449_c23 bl[23] br[23] wl[449] vdd gnd cell_6t
Xbit_r450_c23 bl[23] br[23] wl[450] vdd gnd cell_6t
Xbit_r451_c23 bl[23] br[23] wl[451] vdd gnd cell_6t
Xbit_r452_c23 bl[23] br[23] wl[452] vdd gnd cell_6t
Xbit_r453_c23 bl[23] br[23] wl[453] vdd gnd cell_6t
Xbit_r454_c23 bl[23] br[23] wl[454] vdd gnd cell_6t
Xbit_r455_c23 bl[23] br[23] wl[455] vdd gnd cell_6t
Xbit_r456_c23 bl[23] br[23] wl[456] vdd gnd cell_6t
Xbit_r457_c23 bl[23] br[23] wl[457] vdd gnd cell_6t
Xbit_r458_c23 bl[23] br[23] wl[458] vdd gnd cell_6t
Xbit_r459_c23 bl[23] br[23] wl[459] vdd gnd cell_6t
Xbit_r460_c23 bl[23] br[23] wl[460] vdd gnd cell_6t
Xbit_r461_c23 bl[23] br[23] wl[461] vdd gnd cell_6t
Xbit_r462_c23 bl[23] br[23] wl[462] vdd gnd cell_6t
Xbit_r463_c23 bl[23] br[23] wl[463] vdd gnd cell_6t
Xbit_r464_c23 bl[23] br[23] wl[464] vdd gnd cell_6t
Xbit_r465_c23 bl[23] br[23] wl[465] vdd gnd cell_6t
Xbit_r466_c23 bl[23] br[23] wl[466] vdd gnd cell_6t
Xbit_r467_c23 bl[23] br[23] wl[467] vdd gnd cell_6t
Xbit_r468_c23 bl[23] br[23] wl[468] vdd gnd cell_6t
Xbit_r469_c23 bl[23] br[23] wl[469] vdd gnd cell_6t
Xbit_r470_c23 bl[23] br[23] wl[470] vdd gnd cell_6t
Xbit_r471_c23 bl[23] br[23] wl[471] vdd gnd cell_6t
Xbit_r472_c23 bl[23] br[23] wl[472] vdd gnd cell_6t
Xbit_r473_c23 bl[23] br[23] wl[473] vdd gnd cell_6t
Xbit_r474_c23 bl[23] br[23] wl[474] vdd gnd cell_6t
Xbit_r475_c23 bl[23] br[23] wl[475] vdd gnd cell_6t
Xbit_r476_c23 bl[23] br[23] wl[476] vdd gnd cell_6t
Xbit_r477_c23 bl[23] br[23] wl[477] vdd gnd cell_6t
Xbit_r478_c23 bl[23] br[23] wl[478] vdd gnd cell_6t
Xbit_r479_c23 bl[23] br[23] wl[479] vdd gnd cell_6t
Xbit_r480_c23 bl[23] br[23] wl[480] vdd gnd cell_6t
Xbit_r481_c23 bl[23] br[23] wl[481] vdd gnd cell_6t
Xbit_r482_c23 bl[23] br[23] wl[482] vdd gnd cell_6t
Xbit_r483_c23 bl[23] br[23] wl[483] vdd gnd cell_6t
Xbit_r484_c23 bl[23] br[23] wl[484] vdd gnd cell_6t
Xbit_r485_c23 bl[23] br[23] wl[485] vdd gnd cell_6t
Xbit_r486_c23 bl[23] br[23] wl[486] vdd gnd cell_6t
Xbit_r487_c23 bl[23] br[23] wl[487] vdd gnd cell_6t
Xbit_r488_c23 bl[23] br[23] wl[488] vdd gnd cell_6t
Xbit_r489_c23 bl[23] br[23] wl[489] vdd gnd cell_6t
Xbit_r490_c23 bl[23] br[23] wl[490] vdd gnd cell_6t
Xbit_r491_c23 bl[23] br[23] wl[491] vdd gnd cell_6t
Xbit_r492_c23 bl[23] br[23] wl[492] vdd gnd cell_6t
Xbit_r493_c23 bl[23] br[23] wl[493] vdd gnd cell_6t
Xbit_r494_c23 bl[23] br[23] wl[494] vdd gnd cell_6t
Xbit_r495_c23 bl[23] br[23] wl[495] vdd gnd cell_6t
Xbit_r496_c23 bl[23] br[23] wl[496] vdd gnd cell_6t
Xbit_r497_c23 bl[23] br[23] wl[497] vdd gnd cell_6t
Xbit_r498_c23 bl[23] br[23] wl[498] vdd gnd cell_6t
Xbit_r499_c23 bl[23] br[23] wl[499] vdd gnd cell_6t
Xbit_r500_c23 bl[23] br[23] wl[500] vdd gnd cell_6t
Xbit_r501_c23 bl[23] br[23] wl[501] vdd gnd cell_6t
Xbit_r502_c23 bl[23] br[23] wl[502] vdd gnd cell_6t
Xbit_r503_c23 bl[23] br[23] wl[503] vdd gnd cell_6t
Xbit_r504_c23 bl[23] br[23] wl[504] vdd gnd cell_6t
Xbit_r505_c23 bl[23] br[23] wl[505] vdd gnd cell_6t
Xbit_r506_c23 bl[23] br[23] wl[506] vdd gnd cell_6t
Xbit_r507_c23 bl[23] br[23] wl[507] vdd gnd cell_6t
Xbit_r508_c23 bl[23] br[23] wl[508] vdd gnd cell_6t
Xbit_r509_c23 bl[23] br[23] wl[509] vdd gnd cell_6t
Xbit_r510_c23 bl[23] br[23] wl[510] vdd gnd cell_6t
Xbit_r511_c23 bl[23] br[23] wl[511] vdd gnd cell_6t
Xbit_r0_c24 bl[24] br[24] wl[0] vdd gnd cell_6t
Xbit_r1_c24 bl[24] br[24] wl[1] vdd gnd cell_6t
Xbit_r2_c24 bl[24] br[24] wl[2] vdd gnd cell_6t
Xbit_r3_c24 bl[24] br[24] wl[3] vdd gnd cell_6t
Xbit_r4_c24 bl[24] br[24] wl[4] vdd gnd cell_6t
Xbit_r5_c24 bl[24] br[24] wl[5] vdd gnd cell_6t
Xbit_r6_c24 bl[24] br[24] wl[6] vdd gnd cell_6t
Xbit_r7_c24 bl[24] br[24] wl[7] vdd gnd cell_6t
Xbit_r8_c24 bl[24] br[24] wl[8] vdd gnd cell_6t
Xbit_r9_c24 bl[24] br[24] wl[9] vdd gnd cell_6t
Xbit_r10_c24 bl[24] br[24] wl[10] vdd gnd cell_6t
Xbit_r11_c24 bl[24] br[24] wl[11] vdd gnd cell_6t
Xbit_r12_c24 bl[24] br[24] wl[12] vdd gnd cell_6t
Xbit_r13_c24 bl[24] br[24] wl[13] vdd gnd cell_6t
Xbit_r14_c24 bl[24] br[24] wl[14] vdd gnd cell_6t
Xbit_r15_c24 bl[24] br[24] wl[15] vdd gnd cell_6t
Xbit_r16_c24 bl[24] br[24] wl[16] vdd gnd cell_6t
Xbit_r17_c24 bl[24] br[24] wl[17] vdd gnd cell_6t
Xbit_r18_c24 bl[24] br[24] wl[18] vdd gnd cell_6t
Xbit_r19_c24 bl[24] br[24] wl[19] vdd gnd cell_6t
Xbit_r20_c24 bl[24] br[24] wl[20] vdd gnd cell_6t
Xbit_r21_c24 bl[24] br[24] wl[21] vdd gnd cell_6t
Xbit_r22_c24 bl[24] br[24] wl[22] vdd gnd cell_6t
Xbit_r23_c24 bl[24] br[24] wl[23] vdd gnd cell_6t
Xbit_r24_c24 bl[24] br[24] wl[24] vdd gnd cell_6t
Xbit_r25_c24 bl[24] br[24] wl[25] vdd gnd cell_6t
Xbit_r26_c24 bl[24] br[24] wl[26] vdd gnd cell_6t
Xbit_r27_c24 bl[24] br[24] wl[27] vdd gnd cell_6t
Xbit_r28_c24 bl[24] br[24] wl[28] vdd gnd cell_6t
Xbit_r29_c24 bl[24] br[24] wl[29] vdd gnd cell_6t
Xbit_r30_c24 bl[24] br[24] wl[30] vdd gnd cell_6t
Xbit_r31_c24 bl[24] br[24] wl[31] vdd gnd cell_6t
Xbit_r32_c24 bl[24] br[24] wl[32] vdd gnd cell_6t
Xbit_r33_c24 bl[24] br[24] wl[33] vdd gnd cell_6t
Xbit_r34_c24 bl[24] br[24] wl[34] vdd gnd cell_6t
Xbit_r35_c24 bl[24] br[24] wl[35] vdd gnd cell_6t
Xbit_r36_c24 bl[24] br[24] wl[36] vdd gnd cell_6t
Xbit_r37_c24 bl[24] br[24] wl[37] vdd gnd cell_6t
Xbit_r38_c24 bl[24] br[24] wl[38] vdd gnd cell_6t
Xbit_r39_c24 bl[24] br[24] wl[39] vdd gnd cell_6t
Xbit_r40_c24 bl[24] br[24] wl[40] vdd gnd cell_6t
Xbit_r41_c24 bl[24] br[24] wl[41] vdd gnd cell_6t
Xbit_r42_c24 bl[24] br[24] wl[42] vdd gnd cell_6t
Xbit_r43_c24 bl[24] br[24] wl[43] vdd gnd cell_6t
Xbit_r44_c24 bl[24] br[24] wl[44] vdd gnd cell_6t
Xbit_r45_c24 bl[24] br[24] wl[45] vdd gnd cell_6t
Xbit_r46_c24 bl[24] br[24] wl[46] vdd gnd cell_6t
Xbit_r47_c24 bl[24] br[24] wl[47] vdd gnd cell_6t
Xbit_r48_c24 bl[24] br[24] wl[48] vdd gnd cell_6t
Xbit_r49_c24 bl[24] br[24] wl[49] vdd gnd cell_6t
Xbit_r50_c24 bl[24] br[24] wl[50] vdd gnd cell_6t
Xbit_r51_c24 bl[24] br[24] wl[51] vdd gnd cell_6t
Xbit_r52_c24 bl[24] br[24] wl[52] vdd gnd cell_6t
Xbit_r53_c24 bl[24] br[24] wl[53] vdd gnd cell_6t
Xbit_r54_c24 bl[24] br[24] wl[54] vdd gnd cell_6t
Xbit_r55_c24 bl[24] br[24] wl[55] vdd gnd cell_6t
Xbit_r56_c24 bl[24] br[24] wl[56] vdd gnd cell_6t
Xbit_r57_c24 bl[24] br[24] wl[57] vdd gnd cell_6t
Xbit_r58_c24 bl[24] br[24] wl[58] vdd gnd cell_6t
Xbit_r59_c24 bl[24] br[24] wl[59] vdd gnd cell_6t
Xbit_r60_c24 bl[24] br[24] wl[60] vdd gnd cell_6t
Xbit_r61_c24 bl[24] br[24] wl[61] vdd gnd cell_6t
Xbit_r62_c24 bl[24] br[24] wl[62] vdd gnd cell_6t
Xbit_r63_c24 bl[24] br[24] wl[63] vdd gnd cell_6t
Xbit_r64_c24 bl[24] br[24] wl[64] vdd gnd cell_6t
Xbit_r65_c24 bl[24] br[24] wl[65] vdd gnd cell_6t
Xbit_r66_c24 bl[24] br[24] wl[66] vdd gnd cell_6t
Xbit_r67_c24 bl[24] br[24] wl[67] vdd gnd cell_6t
Xbit_r68_c24 bl[24] br[24] wl[68] vdd gnd cell_6t
Xbit_r69_c24 bl[24] br[24] wl[69] vdd gnd cell_6t
Xbit_r70_c24 bl[24] br[24] wl[70] vdd gnd cell_6t
Xbit_r71_c24 bl[24] br[24] wl[71] vdd gnd cell_6t
Xbit_r72_c24 bl[24] br[24] wl[72] vdd gnd cell_6t
Xbit_r73_c24 bl[24] br[24] wl[73] vdd gnd cell_6t
Xbit_r74_c24 bl[24] br[24] wl[74] vdd gnd cell_6t
Xbit_r75_c24 bl[24] br[24] wl[75] vdd gnd cell_6t
Xbit_r76_c24 bl[24] br[24] wl[76] vdd gnd cell_6t
Xbit_r77_c24 bl[24] br[24] wl[77] vdd gnd cell_6t
Xbit_r78_c24 bl[24] br[24] wl[78] vdd gnd cell_6t
Xbit_r79_c24 bl[24] br[24] wl[79] vdd gnd cell_6t
Xbit_r80_c24 bl[24] br[24] wl[80] vdd gnd cell_6t
Xbit_r81_c24 bl[24] br[24] wl[81] vdd gnd cell_6t
Xbit_r82_c24 bl[24] br[24] wl[82] vdd gnd cell_6t
Xbit_r83_c24 bl[24] br[24] wl[83] vdd gnd cell_6t
Xbit_r84_c24 bl[24] br[24] wl[84] vdd gnd cell_6t
Xbit_r85_c24 bl[24] br[24] wl[85] vdd gnd cell_6t
Xbit_r86_c24 bl[24] br[24] wl[86] vdd gnd cell_6t
Xbit_r87_c24 bl[24] br[24] wl[87] vdd gnd cell_6t
Xbit_r88_c24 bl[24] br[24] wl[88] vdd gnd cell_6t
Xbit_r89_c24 bl[24] br[24] wl[89] vdd gnd cell_6t
Xbit_r90_c24 bl[24] br[24] wl[90] vdd gnd cell_6t
Xbit_r91_c24 bl[24] br[24] wl[91] vdd gnd cell_6t
Xbit_r92_c24 bl[24] br[24] wl[92] vdd gnd cell_6t
Xbit_r93_c24 bl[24] br[24] wl[93] vdd gnd cell_6t
Xbit_r94_c24 bl[24] br[24] wl[94] vdd gnd cell_6t
Xbit_r95_c24 bl[24] br[24] wl[95] vdd gnd cell_6t
Xbit_r96_c24 bl[24] br[24] wl[96] vdd gnd cell_6t
Xbit_r97_c24 bl[24] br[24] wl[97] vdd gnd cell_6t
Xbit_r98_c24 bl[24] br[24] wl[98] vdd gnd cell_6t
Xbit_r99_c24 bl[24] br[24] wl[99] vdd gnd cell_6t
Xbit_r100_c24 bl[24] br[24] wl[100] vdd gnd cell_6t
Xbit_r101_c24 bl[24] br[24] wl[101] vdd gnd cell_6t
Xbit_r102_c24 bl[24] br[24] wl[102] vdd gnd cell_6t
Xbit_r103_c24 bl[24] br[24] wl[103] vdd gnd cell_6t
Xbit_r104_c24 bl[24] br[24] wl[104] vdd gnd cell_6t
Xbit_r105_c24 bl[24] br[24] wl[105] vdd gnd cell_6t
Xbit_r106_c24 bl[24] br[24] wl[106] vdd gnd cell_6t
Xbit_r107_c24 bl[24] br[24] wl[107] vdd gnd cell_6t
Xbit_r108_c24 bl[24] br[24] wl[108] vdd gnd cell_6t
Xbit_r109_c24 bl[24] br[24] wl[109] vdd gnd cell_6t
Xbit_r110_c24 bl[24] br[24] wl[110] vdd gnd cell_6t
Xbit_r111_c24 bl[24] br[24] wl[111] vdd gnd cell_6t
Xbit_r112_c24 bl[24] br[24] wl[112] vdd gnd cell_6t
Xbit_r113_c24 bl[24] br[24] wl[113] vdd gnd cell_6t
Xbit_r114_c24 bl[24] br[24] wl[114] vdd gnd cell_6t
Xbit_r115_c24 bl[24] br[24] wl[115] vdd gnd cell_6t
Xbit_r116_c24 bl[24] br[24] wl[116] vdd gnd cell_6t
Xbit_r117_c24 bl[24] br[24] wl[117] vdd gnd cell_6t
Xbit_r118_c24 bl[24] br[24] wl[118] vdd gnd cell_6t
Xbit_r119_c24 bl[24] br[24] wl[119] vdd gnd cell_6t
Xbit_r120_c24 bl[24] br[24] wl[120] vdd gnd cell_6t
Xbit_r121_c24 bl[24] br[24] wl[121] vdd gnd cell_6t
Xbit_r122_c24 bl[24] br[24] wl[122] vdd gnd cell_6t
Xbit_r123_c24 bl[24] br[24] wl[123] vdd gnd cell_6t
Xbit_r124_c24 bl[24] br[24] wl[124] vdd gnd cell_6t
Xbit_r125_c24 bl[24] br[24] wl[125] vdd gnd cell_6t
Xbit_r126_c24 bl[24] br[24] wl[126] vdd gnd cell_6t
Xbit_r127_c24 bl[24] br[24] wl[127] vdd gnd cell_6t
Xbit_r128_c24 bl[24] br[24] wl[128] vdd gnd cell_6t
Xbit_r129_c24 bl[24] br[24] wl[129] vdd gnd cell_6t
Xbit_r130_c24 bl[24] br[24] wl[130] vdd gnd cell_6t
Xbit_r131_c24 bl[24] br[24] wl[131] vdd gnd cell_6t
Xbit_r132_c24 bl[24] br[24] wl[132] vdd gnd cell_6t
Xbit_r133_c24 bl[24] br[24] wl[133] vdd gnd cell_6t
Xbit_r134_c24 bl[24] br[24] wl[134] vdd gnd cell_6t
Xbit_r135_c24 bl[24] br[24] wl[135] vdd gnd cell_6t
Xbit_r136_c24 bl[24] br[24] wl[136] vdd gnd cell_6t
Xbit_r137_c24 bl[24] br[24] wl[137] vdd gnd cell_6t
Xbit_r138_c24 bl[24] br[24] wl[138] vdd gnd cell_6t
Xbit_r139_c24 bl[24] br[24] wl[139] vdd gnd cell_6t
Xbit_r140_c24 bl[24] br[24] wl[140] vdd gnd cell_6t
Xbit_r141_c24 bl[24] br[24] wl[141] vdd gnd cell_6t
Xbit_r142_c24 bl[24] br[24] wl[142] vdd gnd cell_6t
Xbit_r143_c24 bl[24] br[24] wl[143] vdd gnd cell_6t
Xbit_r144_c24 bl[24] br[24] wl[144] vdd gnd cell_6t
Xbit_r145_c24 bl[24] br[24] wl[145] vdd gnd cell_6t
Xbit_r146_c24 bl[24] br[24] wl[146] vdd gnd cell_6t
Xbit_r147_c24 bl[24] br[24] wl[147] vdd gnd cell_6t
Xbit_r148_c24 bl[24] br[24] wl[148] vdd gnd cell_6t
Xbit_r149_c24 bl[24] br[24] wl[149] vdd gnd cell_6t
Xbit_r150_c24 bl[24] br[24] wl[150] vdd gnd cell_6t
Xbit_r151_c24 bl[24] br[24] wl[151] vdd gnd cell_6t
Xbit_r152_c24 bl[24] br[24] wl[152] vdd gnd cell_6t
Xbit_r153_c24 bl[24] br[24] wl[153] vdd gnd cell_6t
Xbit_r154_c24 bl[24] br[24] wl[154] vdd gnd cell_6t
Xbit_r155_c24 bl[24] br[24] wl[155] vdd gnd cell_6t
Xbit_r156_c24 bl[24] br[24] wl[156] vdd gnd cell_6t
Xbit_r157_c24 bl[24] br[24] wl[157] vdd gnd cell_6t
Xbit_r158_c24 bl[24] br[24] wl[158] vdd gnd cell_6t
Xbit_r159_c24 bl[24] br[24] wl[159] vdd gnd cell_6t
Xbit_r160_c24 bl[24] br[24] wl[160] vdd gnd cell_6t
Xbit_r161_c24 bl[24] br[24] wl[161] vdd gnd cell_6t
Xbit_r162_c24 bl[24] br[24] wl[162] vdd gnd cell_6t
Xbit_r163_c24 bl[24] br[24] wl[163] vdd gnd cell_6t
Xbit_r164_c24 bl[24] br[24] wl[164] vdd gnd cell_6t
Xbit_r165_c24 bl[24] br[24] wl[165] vdd gnd cell_6t
Xbit_r166_c24 bl[24] br[24] wl[166] vdd gnd cell_6t
Xbit_r167_c24 bl[24] br[24] wl[167] vdd gnd cell_6t
Xbit_r168_c24 bl[24] br[24] wl[168] vdd gnd cell_6t
Xbit_r169_c24 bl[24] br[24] wl[169] vdd gnd cell_6t
Xbit_r170_c24 bl[24] br[24] wl[170] vdd gnd cell_6t
Xbit_r171_c24 bl[24] br[24] wl[171] vdd gnd cell_6t
Xbit_r172_c24 bl[24] br[24] wl[172] vdd gnd cell_6t
Xbit_r173_c24 bl[24] br[24] wl[173] vdd gnd cell_6t
Xbit_r174_c24 bl[24] br[24] wl[174] vdd gnd cell_6t
Xbit_r175_c24 bl[24] br[24] wl[175] vdd gnd cell_6t
Xbit_r176_c24 bl[24] br[24] wl[176] vdd gnd cell_6t
Xbit_r177_c24 bl[24] br[24] wl[177] vdd gnd cell_6t
Xbit_r178_c24 bl[24] br[24] wl[178] vdd gnd cell_6t
Xbit_r179_c24 bl[24] br[24] wl[179] vdd gnd cell_6t
Xbit_r180_c24 bl[24] br[24] wl[180] vdd gnd cell_6t
Xbit_r181_c24 bl[24] br[24] wl[181] vdd gnd cell_6t
Xbit_r182_c24 bl[24] br[24] wl[182] vdd gnd cell_6t
Xbit_r183_c24 bl[24] br[24] wl[183] vdd gnd cell_6t
Xbit_r184_c24 bl[24] br[24] wl[184] vdd gnd cell_6t
Xbit_r185_c24 bl[24] br[24] wl[185] vdd gnd cell_6t
Xbit_r186_c24 bl[24] br[24] wl[186] vdd gnd cell_6t
Xbit_r187_c24 bl[24] br[24] wl[187] vdd gnd cell_6t
Xbit_r188_c24 bl[24] br[24] wl[188] vdd gnd cell_6t
Xbit_r189_c24 bl[24] br[24] wl[189] vdd gnd cell_6t
Xbit_r190_c24 bl[24] br[24] wl[190] vdd gnd cell_6t
Xbit_r191_c24 bl[24] br[24] wl[191] vdd gnd cell_6t
Xbit_r192_c24 bl[24] br[24] wl[192] vdd gnd cell_6t
Xbit_r193_c24 bl[24] br[24] wl[193] vdd gnd cell_6t
Xbit_r194_c24 bl[24] br[24] wl[194] vdd gnd cell_6t
Xbit_r195_c24 bl[24] br[24] wl[195] vdd gnd cell_6t
Xbit_r196_c24 bl[24] br[24] wl[196] vdd gnd cell_6t
Xbit_r197_c24 bl[24] br[24] wl[197] vdd gnd cell_6t
Xbit_r198_c24 bl[24] br[24] wl[198] vdd gnd cell_6t
Xbit_r199_c24 bl[24] br[24] wl[199] vdd gnd cell_6t
Xbit_r200_c24 bl[24] br[24] wl[200] vdd gnd cell_6t
Xbit_r201_c24 bl[24] br[24] wl[201] vdd gnd cell_6t
Xbit_r202_c24 bl[24] br[24] wl[202] vdd gnd cell_6t
Xbit_r203_c24 bl[24] br[24] wl[203] vdd gnd cell_6t
Xbit_r204_c24 bl[24] br[24] wl[204] vdd gnd cell_6t
Xbit_r205_c24 bl[24] br[24] wl[205] vdd gnd cell_6t
Xbit_r206_c24 bl[24] br[24] wl[206] vdd gnd cell_6t
Xbit_r207_c24 bl[24] br[24] wl[207] vdd gnd cell_6t
Xbit_r208_c24 bl[24] br[24] wl[208] vdd gnd cell_6t
Xbit_r209_c24 bl[24] br[24] wl[209] vdd gnd cell_6t
Xbit_r210_c24 bl[24] br[24] wl[210] vdd gnd cell_6t
Xbit_r211_c24 bl[24] br[24] wl[211] vdd gnd cell_6t
Xbit_r212_c24 bl[24] br[24] wl[212] vdd gnd cell_6t
Xbit_r213_c24 bl[24] br[24] wl[213] vdd gnd cell_6t
Xbit_r214_c24 bl[24] br[24] wl[214] vdd gnd cell_6t
Xbit_r215_c24 bl[24] br[24] wl[215] vdd gnd cell_6t
Xbit_r216_c24 bl[24] br[24] wl[216] vdd gnd cell_6t
Xbit_r217_c24 bl[24] br[24] wl[217] vdd gnd cell_6t
Xbit_r218_c24 bl[24] br[24] wl[218] vdd gnd cell_6t
Xbit_r219_c24 bl[24] br[24] wl[219] vdd gnd cell_6t
Xbit_r220_c24 bl[24] br[24] wl[220] vdd gnd cell_6t
Xbit_r221_c24 bl[24] br[24] wl[221] vdd gnd cell_6t
Xbit_r222_c24 bl[24] br[24] wl[222] vdd gnd cell_6t
Xbit_r223_c24 bl[24] br[24] wl[223] vdd gnd cell_6t
Xbit_r224_c24 bl[24] br[24] wl[224] vdd gnd cell_6t
Xbit_r225_c24 bl[24] br[24] wl[225] vdd gnd cell_6t
Xbit_r226_c24 bl[24] br[24] wl[226] vdd gnd cell_6t
Xbit_r227_c24 bl[24] br[24] wl[227] vdd gnd cell_6t
Xbit_r228_c24 bl[24] br[24] wl[228] vdd gnd cell_6t
Xbit_r229_c24 bl[24] br[24] wl[229] vdd gnd cell_6t
Xbit_r230_c24 bl[24] br[24] wl[230] vdd gnd cell_6t
Xbit_r231_c24 bl[24] br[24] wl[231] vdd gnd cell_6t
Xbit_r232_c24 bl[24] br[24] wl[232] vdd gnd cell_6t
Xbit_r233_c24 bl[24] br[24] wl[233] vdd gnd cell_6t
Xbit_r234_c24 bl[24] br[24] wl[234] vdd gnd cell_6t
Xbit_r235_c24 bl[24] br[24] wl[235] vdd gnd cell_6t
Xbit_r236_c24 bl[24] br[24] wl[236] vdd gnd cell_6t
Xbit_r237_c24 bl[24] br[24] wl[237] vdd gnd cell_6t
Xbit_r238_c24 bl[24] br[24] wl[238] vdd gnd cell_6t
Xbit_r239_c24 bl[24] br[24] wl[239] vdd gnd cell_6t
Xbit_r240_c24 bl[24] br[24] wl[240] vdd gnd cell_6t
Xbit_r241_c24 bl[24] br[24] wl[241] vdd gnd cell_6t
Xbit_r242_c24 bl[24] br[24] wl[242] vdd gnd cell_6t
Xbit_r243_c24 bl[24] br[24] wl[243] vdd gnd cell_6t
Xbit_r244_c24 bl[24] br[24] wl[244] vdd gnd cell_6t
Xbit_r245_c24 bl[24] br[24] wl[245] vdd gnd cell_6t
Xbit_r246_c24 bl[24] br[24] wl[246] vdd gnd cell_6t
Xbit_r247_c24 bl[24] br[24] wl[247] vdd gnd cell_6t
Xbit_r248_c24 bl[24] br[24] wl[248] vdd gnd cell_6t
Xbit_r249_c24 bl[24] br[24] wl[249] vdd gnd cell_6t
Xbit_r250_c24 bl[24] br[24] wl[250] vdd gnd cell_6t
Xbit_r251_c24 bl[24] br[24] wl[251] vdd gnd cell_6t
Xbit_r252_c24 bl[24] br[24] wl[252] vdd gnd cell_6t
Xbit_r253_c24 bl[24] br[24] wl[253] vdd gnd cell_6t
Xbit_r254_c24 bl[24] br[24] wl[254] vdd gnd cell_6t
Xbit_r255_c24 bl[24] br[24] wl[255] vdd gnd cell_6t
Xbit_r256_c24 bl[24] br[24] wl[256] vdd gnd cell_6t
Xbit_r257_c24 bl[24] br[24] wl[257] vdd gnd cell_6t
Xbit_r258_c24 bl[24] br[24] wl[258] vdd gnd cell_6t
Xbit_r259_c24 bl[24] br[24] wl[259] vdd gnd cell_6t
Xbit_r260_c24 bl[24] br[24] wl[260] vdd gnd cell_6t
Xbit_r261_c24 bl[24] br[24] wl[261] vdd gnd cell_6t
Xbit_r262_c24 bl[24] br[24] wl[262] vdd gnd cell_6t
Xbit_r263_c24 bl[24] br[24] wl[263] vdd gnd cell_6t
Xbit_r264_c24 bl[24] br[24] wl[264] vdd gnd cell_6t
Xbit_r265_c24 bl[24] br[24] wl[265] vdd gnd cell_6t
Xbit_r266_c24 bl[24] br[24] wl[266] vdd gnd cell_6t
Xbit_r267_c24 bl[24] br[24] wl[267] vdd gnd cell_6t
Xbit_r268_c24 bl[24] br[24] wl[268] vdd gnd cell_6t
Xbit_r269_c24 bl[24] br[24] wl[269] vdd gnd cell_6t
Xbit_r270_c24 bl[24] br[24] wl[270] vdd gnd cell_6t
Xbit_r271_c24 bl[24] br[24] wl[271] vdd gnd cell_6t
Xbit_r272_c24 bl[24] br[24] wl[272] vdd gnd cell_6t
Xbit_r273_c24 bl[24] br[24] wl[273] vdd gnd cell_6t
Xbit_r274_c24 bl[24] br[24] wl[274] vdd gnd cell_6t
Xbit_r275_c24 bl[24] br[24] wl[275] vdd gnd cell_6t
Xbit_r276_c24 bl[24] br[24] wl[276] vdd gnd cell_6t
Xbit_r277_c24 bl[24] br[24] wl[277] vdd gnd cell_6t
Xbit_r278_c24 bl[24] br[24] wl[278] vdd gnd cell_6t
Xbit_r279_c24 bl[24] br[24] wl[279] vdd gnd cell_6t
Xbit_r280_c24 bl[24] br[24] wl[280] vdd gnd cell_6t
Xbit_r281_c24 bl[24] br[24] wl[281] vdd gnd cell_6t
Xbit_r282_c24 bl[24] br[24] wl[282] vdd gnd cell_6t
Xbit_r283_c24 bl[24] br[24] wl[283] vdd gnd cell_6t
Xbit_r284_c24 bl[24] br[24] wl[284] vdd gnd cell_6t
Xbit_r285_c24 bl[24] br[24] wl[285] vdd gnd cell_6t
Xbit_r286_c24 bl[24] br[24] wl[286] vdd gnd cell_6t
Xbit_r287_c24 bl[24] br[24] wl[287] vdd gnd cell_6t
Xbit_r288_c24 bl[24] br[24] wl[288] vdd gnd cell_6t
Xbit_r289_c24 bl[24] br[24] wl[289] vdd gnd cell_6t
Xbit_r290_c24 bl[24] br[24] wl[290] vdd gnd cell_6t
Xbit_r291_c24 bl[24] br[24] wl[291] vdd gnd cell_6t
Xbit_r292_c24 bl[24] br[24] wl[292] vdd gnd cell_6t
Xbit_r293_c24 bl[24] br[24] wl[293] vdd gnd cell_6t
Xbit_r294_c24 bl[24] br[24] wl[294] vdd gnd cell_6t
Xbit_r295_c24 bl[24] br[24] wl[295] vdd gnd cell_6t
Xbit_r296_c24 bl[24] br[24] wl[296] vdd gnd cell_6t
Xbit_r297_c24 bl[24] br[24] wl[297] vdd gnd cell_6t
Xbit_r298_c24 bl[24] br[24] wl[298] vdd gnd cell_6t
Xbit_r299_c24 bl[24] br[24] wl[299] vdd gnd cell_6t
Xbit_r300_c24 bl[24] br[24] wl[300] vdd gnd cell_6t
Xbit_r301_c24 bl[24] br[24] wl[301] vdd gnd cell_6t
Xbit_r302_c24 bl[24] br[24] wl[302] vdd gnd cell_6t
Xbit_r303_c24 bl[24] br[24] wl[303] vdd gnd cell_6t
Xbit_r304_c24 bl[24] br[24] wl[304] vdd gnd cell_6t
Xbit_r305_c24 bl[24] br[24] wl[305] vdd gnd cell_6t
Xbit_r306_c24 bl[24] br[24] wl[306] vdd gnd cell_6t
Xbit_r307_c24 bl[24] br[24] wl[307] vdd gnd cell_6t
Xbit_r308_c24 bl[24] br[24] wl[308] vdd gnd cell_6t
Xbit_r309_c24 bl[24] br[24] wl[309] vdd gnd cell_6t
Xbit_r310_c24 bl[24] br[24] wl[310] vdd gnd cell_6t
Xbit_r311_c24 bl[24] br[24] wl[311] vdd gnd cell_6t
Xbit_r312_c24 bl[24] br[24] wl[312] vdd gnd cell_6t
Xbit_r313_c24 bl[24] br[24] wl[313] vdd gnd cell_6t
Xbit_r314_c24 bl[24] br[24] wl[314] vdd gnd cell_6t
Xbit_r315_c24 bl[24] br[24] wl[315] vdd gnd cell_6t
Xbit_r316_c24 bl[24] br[24] wl[316] vdd gnd cell_6t
Xbit_r317_c24 bl[24] br[24] wl[317] vdd gnd cell_6t
Xbit_r318_c24 bl[24] br[24] wl[318] vdd gnd cell_6t
Xbit_r319_c24 bl[24] br[24] wl[319] vdd gnd cell_6t
Xbit_r320_c24 bl[24] br[24] wl[320] vdd gnd cell_6t
Xbit_r321_c24 bl[24] br[24] wl[321] vdd gnd cell_6t
Xbit_r322_c24 bl[24] br[24] wl[322] vdd gnd cell_6t
Xbit_r323_c24 bl[24] br[24] wl[323] vdd gnd cell_6t
Xbit_r324_c24 bl[24] br[24] wl[324] vdd gnd cell_6t
Xbit_r325_c24 bl[24] br[24] wl[325] vdd gnd cell_6t
Xbit_r326_c24 bl[24] br[24] wl[326] vdd gnd cell_6t
Xbit_r327_c24 bl[24] br[24] wl[327] vdd gnd cell_6t
Xbit_r328_c24 bl[24] br[24] wl[328] vdd gnd cell_6t
Xbit_r329_c24 bl[24] br[24] wl[329] vdd gnd cell_6t
Xbit_r330_c24 bl[24] br[24] wl[330] vdd gnd cell_6t
Xbit_r331_c24 bl[24] br[24] wl[331] vdd gnd cell_6t
Xbit_r332_c24 bl[24] br[24] wl[332] vdd gnd cell_6t
Xbit_r333_c24 bl[24] br[24] wl[333] vdd gnd cell_6t
Xbit_r334_c24 bl[24] br[24] wl[334] vdd gnd cell_6t
Xbit_r335_c24 bl[24] br[24] wl[335] vdd gnd cell_6t
Xbit_r336_c24 bl[24] br[24] wl[336] vdd gnd cell_6t
Xbit_r337_c24 bl[24] br[24] wl[337] vdd gnd cell_6t
Xbit_r338_c24 bl[24] br[24] wl[338] vdd gnd cell_6t
Xbit_r339_c24 bl[24] br[24] wl[339] vdd gnd cell_6t
Xbit_r340_c24 bl[24] br[24] wl[340] vdd gnd cell_6t
Xbit_r341_c24 bl[24] br[24] wl[341] vdd gnd cell_6t
Xbit_r342_c24 bl[24] br[24] wl[342] vdd gnd cell_6t
Xbit_r343_c24 bl[24] br[24] wl[343] vdd gnd cell_6t
Xbit_r344_c24 bl[24] br[24] wl[344] vdd gnd cell_6t
Xbit_r345_c24 bl[24] br[24] wl[345] vdd gnd cell_6t
Xbit_r346_c24 bl[24] br[24] wl[346] vdd gnd cell_6t
Xbit_r347_c24 bl[24] br[24] wl[347] vdd gnd cell_6t
Xbit_r348_c24 bl[24] br[24] wl[348] vdd gnd cell_6t
Xbit_r349_c24 bl[24] br[24] wl[349] vdd gnd cell_6t
Xbit_r350_c24 bl[24] br[24] wl[350] vdd gnd cell_6t
Xbit_r351_c24 bl[24] br[24] wl[351] vdd gnd cell_6t
Xbit_r352_c24 bl[24] br[24] wl[352] vdd gnd cell_6t
Xbit_r353_c24 bl[24] br[24] wl[353] vdd gnd cell_6t
Xbit_r354_c24 bl[24] br[24] wl[354] vdd gnd cell_6t
Xbit_r355_c24 bl[24] br[24] wl[355] vdd gnd cell_6t
Xbit_r356_c24 bl[24] br[24] wl[356] vdd gnd cell_6t
Xbit_r357_c24 bl[24] br[24] wl[357] vdd gnd cell_6t
Xbit_r358_c24 bl[24] br[24] wl[358] vdd gnd cell_6t
Xbit_r359_c24 bl[24] br[24] wl[359] vdd gnd cell_6t
Xbit_r360_c24 bl[24] br[24] wl[360] vdd gnd cell_6t
Xbit_r361_c24 bl[24] br[24] wl[361] vdd gnd cell_6t
Xbit_r362_c24 bl[24] br[24] wl[362] vdd gnd cell_6t
Xbit_r363_c24 bl[24] br[24] wl[363] vdd gnd cell_6t
Xbit_r364_c24 bl[24] br[24] wl[364] vdd gnd cell_6t
Xbit_r365_c24 bl[24] br[24] wl[365] vdd gnd cell_6t
Xbit_r366_c24 bl[24] br[24] wl[366] vdd gnd cell_6t
Xbit_r367_c24 bl[24] br[24] wl[367] vdd gnd cell_6t
Xbit_r368_c24 bl[24] br[24] wl[368] vdd gnd cell_6t
Xbit_r369_c24 bl[24] br[24] wl[369] vdd gnd cell_6t
Xbit_r370_c24 bl[24] br[24] wl[370] vdd gnd cell_6t
Xbit_r371_c24 bl[24] br[24] wl[371] vdd gnd cell_6t
Xbit_r372_c24 bl[24] br[24] wl[372] vdd gnd cell_6t
Xbit_r373_c24 bl[24] br[24] wl[373] vdd gnd cell_6t
Xbit_r374_c24 bl[24] br[24] wl[374] vdd gnd cell_6t
Xbit_r375_c24 bl[24] br[24] wl[375] vdd gnd cell_6t
Xbit_r376_c24 bl[24] br[24] wl[376] vdd gnd cell_6t
Xbit_r377_c24 bl[24] br[24] wl[377] vdd gnd cell_6t
Xbit_r378_c24 bl[24] br[24] wl[378] vdd gnd cell_6t
Xbit_r379_c24 bl[24] br[24] wl[379] vdd gnd cell_6t
Xbit_r380_c24 bl[24] br[24] wl[380] vdd gnd cell_6t
Xbit_r381_c24 bl[24] br[24] wl[381] vdd gnd cell_6t
Xbit_r382_c24 bl[24] br[24] wl[382] vdd gnd cell_6t
Xbit_r383_c24 bl[24] br[24] wl[383] vdd gnd cell_6t
Xbit_r384_c24 bl[24] br[24] wl[384] vdd gnd cell_6t
Xbit_r385_c24 bl[24] br[24] wl[385] vdd gnd cell_6t
Xbit_r386_c24 bl[24] br[24] wl[386] vdd gnd cell_6t
Xbit_r387_c24 bl[24] br[24] wl[387] vdd gnd cell_6t
Xbit_r388_c24 bl[24] br[24] wl[388] vdd gnd cell_6t
Xbit_r389_c24 bl[24] br[24] wl[389] vdd gnd cell_6t
Xbit_r390_c24 bl[24] br[24] wl[390] vdd gnd cell_6t
Xbit_r391_c24 bl[24] br[24] wl[391] vdd gnd cell_6t
Xbit_r392_c24 bl[24] br[24] wl[392] vdd gnd cell_6t
Xbit_r393_c24 bl[24] br[24] wl[393] vdd gnd cell_6t
Xbit_r394_c24 bl[24] br[24] wl[394] vdd gnd cell_6t
Xbit_r395_c24 bl[24] br[24] wl[395] vdd gnd cell_6t
Xbit_r396_c24 bl[24] br[24] wl[396] vdd gnd cell_6t
Xbit_r397_c24 bl[24] br[24] wl[397] vdd gnd cell_6t
Xbit_r398_c24 bl[24] br[24] wl[398] vdd gnd cell_6t
Xbit_r399_c24 bl[24] br[24] wl[399] vdd gnd cell_6t
Xbit_r400_c24 bl[24] br[24] wl[400] vdd gnd cell_6t
Xbit_r401_c24 bl[24] br[24] wl[401] vdd gnd cell_6t
Xbit_r402_c24 bl[24] br[24] wl[402] vdd gnd cell_6t
Xbit_r403_c24 bl[24] br[24] wl[403] vdd gnd cell_6t
Xbit_r404_c24 bl[24] br[24] wl[404] vdd gnd cell_6t
Xbit_r405_c24 bl[24] br[24] wl[405] vdd gnd cell_6t
Xbit_r406_c24 bl[24] br[24] wl[406] vdd gnd cell_6t
Xbit_r407_c24 bl[24] br[24] wl[407] vdd gnd cell_6t
Xbit_r408_c24 bl[24] br[24] wl[408] vdd gnd cell_6t
Xbit_r409_c24 bl[24] br[24] wl[409] vdd gnd cell_6t
Xbit_r410_c24 bl[24] br[24] wl[410] vdd gnd cell_6t
Xbit_r411_c24 bl[24] br[24] wl[411] vdd gnd cell_6t
Xbit_r412_c24 bl[24] br[24] wl[412] vdd gnd cell_6t
Xbit_r413_c24 bl[24] br[24] wl[413] vdd gnd cell_6t
Xbit_r414_c24 bl[24] br[24] wl[414] vdd gnd cell_6t
Xbit_r415_c24 bl[24] br[24] wl[415] vdd gnd cell_6t
Xbit_r416_c24 bl[24] br[24] wl[416] vdd gnd cell_6t
Xbit_r417_c24 bl[24] br[24] wl[417] vdd gnd cell_6t
Xbit_r418_c24 bl[24] br[24] wl[418] vdd gnd cell_6t
Xbit_r419_c24 bl[24] br[24] wl[419] vdd gnd cell_6t
Xbit_r420_c24 bl[24] br[24] wl[420] vdd gnd cell_6t
Xbit_r421_c24 bl[24] br[24] wl[421] vdd gnd cell_6t
Xbit_r422_c24 bl[24] br[24] wl[422] vdd gnd cell_6t
Xbit_r423_c24 bl[24] br[24] wl[423] vdd gnd cell_6t
Xbit_r424_c24 bl[24] br[24] wl[424] vdd gnd cell_6t
Xbit_r425_c24 bl[24] br[24] wl[425] vdd gnd cell_6t
Xbit_r426_c24 bl[24] br[24] wl[426] vdd gnd cell_6t
Xbit_r427_c24 bl[24] br[24] wl[427] vdd gnd cell_6t
Xbit_r428_c24 bl[24] br[24] wl[428] vdd gnd cell_6t
Xbit_r429_c24 bl[24] br[24] wl[429] vdd gnd cell_6t
Xbit_r430_c24 bl[24] br[24] wl[430] vdd gnd cell_6t
Xbit_r431_c24 bl[24] br[24] wl[431] vdd gnd cell_6t
Xbit_r432_c24 bl[24] br[24] wl[432] vdd gnd cell_6t
Xbit_r433_c24 bl[24] br[24] wl[433] vdd gnd cell_6t
Xbit_r434_c24 bl[24] br[24] wl[434] vdd gnd cell_6t
Xbit_r435_c24 bl[24] br[24] wl[435] vdd gnd cell_6t
Xbit_r436_c24 bl[24] br[24] wl[436] vdd gnd cell_6t
Xbit_r437_c24 bl[24] br[24] wl[437] vdd gnd cell_6t
Xbit_r438_c24 bl[24] br[24] wl[438] vdd gnd cell_6t
Xbit_r439_c24 bl[24] br[24] wl[439] vdd gnd cell_6t
Xbit_r440_c24 bl[24] br[24] wl[440] vdd gnd cell_6t
Xbit_r441_c24 bl[24] br[24] wl[441] vdd gnd cell_6t
Xbit_r442_c24 bl[24] br[24] wl[442] vdd gnd cell_6t
Xbit_r443_c24 bl[24] br[24] wl[443] vdd gnd cell_6t
Xbit_r444_c24 bl[24] br[24] wl[444] vdd gnd cell_6t
Xbit_r445_c24 bl[24] br[24] wl[445] vdd gnd cell_6t
Xbit_r446_c24 bl[24] br[24] wl[446] vdd gnd cell_6t
Xbit_r447_c24 bl[24] br[24] wl[447] vdd gnd cell_6t
Xbit_r448_c24 bl[24] br[24] wl[448] vdd gnd cell_6t
Xbit_r449_c24 bl[24] br[24] wl[449] vdd gnd cell_6t
Xbit_r450_c24 bl[24] br[24] wl[450] vdd gnd cell_6t
Xbit_r451_c24 bl[24] br[24] wl[451] vdd gnd cell_6t
Xbit_r452_c24 bl[24] br[24] wl[452] vdd gnd cell_6t
Xbit_r453_c24 bl[24] br[24] wl[453] vdd gnd cell_6t
Xbit_r454_c24 bl[24] br[24] wl[454] vdd gnd cell_6t
Xbit_r455_c24 bl[24] br[24] wl[455] vdd gnd cell_6t
Xbit_r456_c24 bl[24] br[24] wl[456] vdd gnd cell_6t
Xbit_r457_c24 bl[24] br[24] wl[457] vdd gnd cell_6t
Xbit_r458_c24 bl[24] br[24] wl[458] vdd gnd cell_6t
Xbit_r459_c24 bl[24] br[24] wl[459] vdd gnd cell_6t
Xbit_r460_c24 bl[24] br[24] wl[460] vdd gnd cell_6t
Xbit_r461_c24 bl[24] br[24] wl[461] vdd gnd cell_6t
Xbit_r462_c24 bl[24] br[24] wl[462] vdd gnd cell_6t
Xbit_r463_c24 bl[24] br[24] wl[463] vdd gnd cell_6t
Xbit_r464_c24 bl[24] br[24] wl[464] vdd gnd cell_6t
Xbit_r465_c24 bl[24] br[24] wl[465] vdd gnd cell_6t
Xbit_r466_c24 bl[24] br[24] wl[466] vdd gnd cell_6t
Xbit_r467_c24 bl[24] br[24] wl[467] vdd gnd cell_6t
Xbit_r468_c24 bl[24] br[24] wl[468] vdd gnd cell_6t
Xbit_r469_c24 bl[24] br[24] wl[469] vdd gnd cell_6t
Xbit_r470_c24 bl[24] br[24] wl[470] vdd gnd cell_6t
Xbit_r471_c24 bl[24] br[24] wl[471] vdd gnd cell_6t
Xbit_r472_c24 bl[24] br[24] wl[472] vdd gnd cell_6t
Xbit_r473_c24 bl[24] br[24] wl[473] vdd gnd cell_6t
Xbit_r474_c24 bl[24] br[24] wl[474] vdd gnd cell_6t
Xbit_r475_c24 bl[24] br[24] wl[475] vdd gnd cell_6t
Xbit_r476_c24 bl[24] br[24] wl[476] vdd gnd cell_6t
Xbit_r477_c24 bl[24] br[24] wl[477] vdd gnd cell_6t
Xbit_r478_c24 bl[24] br[24] wl[478] vdd gnd cell_6t
Xbit_r479_c24 bl[24] br[24] wl[479] vdd gnd cell_6t
Xbit_r480_c24 bl[24] br[24] wl[480] vdd gnd cell_6t
Xbit_r481_c24 bl[24] br[24] wl[481] vdd gnd cell_6t
Xbit_r482_c24 bl[24] br[24] wl[482] vdd gnd cell_6t
Xbit_r483_c24 bl[24] br[24] wl[483] vdd gnd cell_6t
Xbit_r484_c24 bl[24] br[24] wl[484] vdd gnd cell_6t
Xbit_r485_c24 bl[24] br[24] wl[485] vdd gnd cell_6t
Xbit_r486_c24 bl[24] br[24] wl[486] vdd gnd cell_6t
Xbit_r487_c24 bl[24] br[24] wl[487] vdd gnd cell_6t
Xbit_r488_c24 bl[24] br[24] wl[488] vdd gnd cell_6t
Xbit_r489_c24 bl[24] br[24] wl[489] vdd gnd cell_6t
Xbit_r490_c24 bl[24] br[24] wl[490] vdd gnd cell_6t
Xbit_r491_c24 bl[24] br[24] wl[491] vdd gnd cell_6t
Xbit_r492_c24 bl[24] br[24] wl[492] vdd gnd cell_6t
Xbit_r493_c24 bl[24] br[24] wl[493] vdd gnd cell_6t
Xbit_r494_c24 bl[24] br[24] wl[494] vdd gnd cell_6t
Xbit_r495_c24 bl[24] br[24] wl[495] vdd gnd cell_6t
Xbit_r496_c24 bl[24] br[24] wl[496] vdd gnd cell_6t
Xbit_r497_c24 bl[24] br[24] wl[497] vdd gnd cell_6t
Xbit_r498_c24 bl[24] br[24] wl[498] vdd gnd cell_6t
Xbit_r499_c24 bl[24] br[24] wl[499] vdd gnd cell_6t
Xbit_r500_c24 bl[24] br[24] wl[500] vdd gnd cell_6t
Xbit_r501_c24 bl[24] br[24] wl[501] vdd gnd cell_6t
Xbit_r502_c24 bl[24] br[24] wl[502] vdd gnd cell_6t
Xbit_r503_c24 bl[24] br[24] wl[503] vdd gnd cell_6t
Xbit_r504_c24 bl[24] br[24] wl[504] vdd gnd cell_6t
Xbit_r505_c24 bl[24] br[24] wl[505] vdd gnd cell_6t
Xbit_r506_c24 bl[24] br[24] wl[506] vdd gnd cell_6t
Xbit_r507_c24 bl[24] br[24] wl[507] vdd gnd cell_6t
Xbit_r508_c24 bl[24] br[24] wl[508] vdd gnd cell_6t
Xbit_r509_c24 bl[24] br[24] wl[509] vdd gnd cell_6t
Xbit_r510_c24 bl[24] br[24] wl[510] vdd gnd cell_6t
Xbit_r511_c24 bl[24] br[24] wl[511] vdd gnd cell_6t
Xbit_r0_c25 bl[25] br[25] wl[0] vdd gnd cell_6t
Xbit_r1_c25 bl[25] br[25] wl[1] vdd gnd cell_6t
Xbit_r2_c25 bl[25] br[25] wl[2] vdd gnd cell_6t
Xbit_r3_c25 bl[25] br[25] wl[3] vdd gnd cell_6t
Xbit_r4_c25 bl[25] br[25] wl[4] vdd gnd cell_6t
Xbit_r5_c25 bl[25] br[25] wl[5] vdd gnd cell_6t
Xbit_r6_c25 bl[25] br[25] wl[6] vdd gnd cell_6t
Xbit_r7_c25 bl[25] br[25] wl[7] vdd gnd cell_6t
Xbit_r8_c25 bl[25] br[25] wl[8] vdd gnd cell_6t
Xbit_r9_c25 bl[25] br[25] wl[9] vdd gnd cell_6t
Xbit_r10_c25 bl[25] br[25] wl[10] vdd gnd cell_6t
Xbit_r11_c25 bl[25] br[25] wl[11] vdd gnd cell_6t
Xbit_r12_c25 bl[25] br[25] wl[12] vdd gnd cell_6t
Xbit_r13_c25 bl[25] br[25] wl[13] vdd gnd cell_6t
Xbit_r14_c25 bl[25] br[25] wl[14] vdd gnd cell_6t
Xbit_r15_c25 bl[25] br[25] wl[15] vdd gnd cell_6t
Xbit_r16_c25 bl[25] br[25] wl[16] vdd gnd cell_6t
Xbit_r17_c25 bl[25] br[25] wl[17] vdd gnd cell_6t
Xbit_r18_c25 bl[25] br[25] wl[18] vdd gnd cell_6t
Xbit_r19_c25 bl[25] br[25] wl[19] vdd gnd cell_6t
Xbit_r20_c25 bl[25] br[25] wl[20] vdd gnd cell_6t
Xbit_r21_c25 bl[25] br[25] wl[21] vdd gnd cell_6t
Xbit_r22_c25 bl[25] br[25] wl[22] vdd gnd cell_6t
Xbit_r23_c25 bl[25] br[25] wl[23] vdd gnd cell_6t
Xbit_r24_c25 bl[25] br[25] wl[24] vdd gnd cell_6t
Xbit_r25_c25 bl[25] br[25] wl[25] vdd gnd cell_6t
Xbit_r26_c25 bl[25] br[25] wl[26] vdd gnd cell_6t
Xbit_r27_c25 bl[25] br[25] wl[27] vdd gnd cell_6t
Xbit_r28_c25 bl[25] br[25] wl[28] vdd gnd cell_6t
Xbit_r29_c25 bl[25] br[25] wl[29] vdd gnd cell_6t
Xbit_r30_c25 bl[25] br[25] wl[30] vdd gnd cell_6t
Xbit_r31_c25 bl[25] br[25] wl[31] vdd gnd cell_6t
Xbit_r32_c25 bl[25] br[25] wl[32] vdd gnd cell_6t
Xbit_r33_c25 bl[25] br[25] wl[33] vdd gnd cell_6t
Xbit_r34_c25 bl[25] br[25] wl[34] vdd gnd cell_6t
Xbit_r35_c25 bl[25] br[25] wl[35] vdd gnd cell_6t
Xbit_r36_c25 bl[25] br[25] wl[36] vdd gnd cell_6t
Xbit_r37_c25 bl[25] br[25] wl[37] vdd gnd cell_6t
Xbit_r38_c25 bl[25] br[25] wl[38] vdd gnd cell_6t
Xbit_r39_c25 bl[25] br[25] wl[39] vdd gnd cell_6t
Xbit_r40_c25 bl[25] br[25] wl[40] vdd gnd cell_6t
Xbit_r41_c25 bl[25] br[25] wl[41] vdd gnd cell_6t
Xbit_r42_c25 bl[25] br[25] wl[42] vdd gnd cell_6t
Xbit_r43_c25 bl[25] br[25] wl[43] vdd gnd cell_6t
Xbit_r44_c25 bl[25] br[25] wl[44] vdd gnd cell_6t
Xbit_r45_c25 bl[25] br[25] wl[45] vdd gnd cell_6t
Xbit_r46_c25 bl[25] br[25] wl[46] vdd gnd cell_6t
Xbit_r47_c25 bl[25] br[25] wl[47] vdd gnd cell_6t
Xbit_r48_c25 bl[25] br[25] wl[48] vdd gnd cell_6t
Xbit_r49_c25 bl[25] br[25] wl[49] vdd gnd cell_6t
Xbit_r50_c25 bl[25] br[25] wl[50] vdd gnd cell_6t
Xbit_r51_c25 bl[25] br[25] wl[51] vdd gnd cell_6t
Xbit_r52_c25 bl[25] br[25] wl[52] vdd gnd cell_6t
Xbit_r53_c25 bl[25] br[25] wl[53] vdd gnd cell_6t
Xbit_r54_c25 bl[25] br[25] wl[54] vdd gnd cell_6t
Xbit_r55_c25 bl[25] br[25] wl[55] vdd gnd cell_6t
Xbit_r56_c25 bl[25] br[25] wl[56] vdd gnd cell_6t
Xbit_r57_c25 bl[25] br[25] wl[57] vdd gnd cell_6t
Xbit_r58_c25 bl[25] br[25] wl[58] vdd gnd cell_6t
Xbit_r59_c25 bl[25] br[25] wl[59] vdd gnd cell_6t
Xbit_r60_c25 bl[25] br[25] wl[60] vdd gnd cell_6t
Xbit_r61_c25 bl[25] br[25] wl[61] vdd gnd cell_6t
Xbit_r62_c25 bl[25] br[25] wl[62] vdd gnd cell_6t
Xbit_r63_c25 bl[25] br[25] wl[63] vdd gnd cell_6t
Xbit_r64_c25 bl[25] br[25] wl[64] vdd gnd cell_6t
Xbit_r65_c25 bl[25] br[25] wl[65] vdd gnd cell_6t
Xbit_r66_c25 bl[25] br[25] wl[66] vdd gnd cell_6t
Xbit_r67_c25 bl[25] br[25] wl[67] vdd gnd cell_6t
Xbit_r68_c25 bl[25] br[25] wl[68] vdd gnd cell_6t
Xbit_r69_c25 bl[25] br[25] wl[69] vdd gnd cell_6t
Xbit_r70_c25 bl[25] br[25] wl[70] vdd gnd cell_6t
Xbit_r71_c25 bl[25] br[25] wl[71] vdd gnd cell_6t
Xbit_r72_c25 bl[25] br[25] wl[72] vdd gnd cell_6t
Xbit_r73_c25 bl[25] br[25] wl[73] vdd gnd cell_6t
Xbit_r74_c25 bl[25] br[25] wl[74] vdd gnd cell_6t
Xbit_r75_c25 bl[25] br[25] wl[75] vdd gnd cell_6t
Xbit_r76_c25 bl[25] br[25] wl[76] vdd gnd cell_6t
Xbit_r77_c25 bl[25] br[25] wl[77] vdd gnd cell_6t
Xbit_r78_c25 bl[25] br[25] wl[78] vdd gnd cell_6t
Xbit_r79_c25 bl[25] br[25] wl[79] vdd gnd cell_6t
Xbit_r80_c25 bl[25] br[25] wl[80] vdd gnd cell_6t
Xbit_r81_c25 bl[25] br[25] wl[81] vdd gnd cell_6t
Xbit_r82_c25 bl[25] br[25] wl[82] vdd gnd cell_6t
Xbit_r83_c25 bl[25] br[25] wl[83] vdd gnd cell_6t
Xbit_r84_c25 bl[25] br[25] wl[84] vdd gnd cell_6t
Xbit_r85_c25 bl[25] br[25] wl[85] vdd gnd cell_6t
Xbit_r86_c25 bl[25] br[25] wl[86] vdd gnd cell_6t
Xbit_r87_c25 bl[25] br[25] wl[87] vdd gnd cell_6t
Xbit_r88_c25 bl[25] br[25] wl[88] vdd gnd cell_6t
Xbit_r89_c25 bl[25] br[25] wl[89] vdd gnd cell_6t
Xbit_r90_c25 bl[25] br[25] wl[90] vdd gnd cell_6t
Xbit_r91_c25 bl[25] br[25] wl[91] vdd gnd cell_6t
Xbit_r92_c25 bl[25] br[25] wl[92] vdd gnd cell_6t
Xbit_r93_c25 bl[25] br[25] wl[93] vdd gnd cell_6t
Xbit_r94_c25 bl[25] br[25] wl[94] vdd gnd cell_6t
Xbit_r95_c25 bl[25] br[25] wl[95] vdd gnd cell_6t
Xbit_r96_c25 bl[25] br[25] wl[96] vdd gnd cell_6t
Xbit_r97_c25 bl[25] br[25] wl[97] vdd gnd cell_6t
Xbit_r98_c25 bl[25] br[25] wl[98] vdd gnd cell_6t
Xbit_r99_c25 bl[25] br[25] wl[99] vdd gnd cell_6t
Xbit_r100_c25 bl[25] br[25] wl[100] vdd gnd cell_6t
Xbit_r101_c25 bl[25] br[25] wl[101] vdd gnd cell_6t
Xbit_r102_c25 bl[25] br[25] wl[102] vdd gnd cell_6t
Xbit_r103_c25 bl[25] br[25] wl[103] vdd gnd cell_6t
Xbit_r104_c25 bl[25] br[25] wl[104] vdd gnd cell_6t
Xbit_r105_c25 bl[25] br[25] wl[105] vdd gnd cell_6t
Xbit_r106_c25 bl[25] br[25] wl[106] vdd gnd cell_6t
Xbit_r107_c25 bl[25] br[25] wl[107] vdd gnd cell_6t
Xbit_r108_c25 bl[25] br[25] wl[108] vdd gnd cell_6t
Xbit_r109_c25 bl[25] br[25] wl[109] vdd gnd cell_6t
Xbit_r110_c25 bl[25] br[25] wl[110] vdd gnd cell_6t
Xbit_r111_c25 bl[25] br[25] wl[111] vdd gnd cell_6t
Xbit_r112_c25 bl[25] br[25] wl[112] vdd gnd cell_6t
Xbit_r113_c25 bl[25] br[25] wl[113] vdd gnd cell_6t
Xbit_r114_c25 bl[25] br[25] wl[114] vdd gnd cell_6t
Xbit_r115_c25 bl[25] br[25] wl[115] vdd gnd cell_6t
Xbit_r116_c25 bl[25] br[25] wl[116] vdd gnd cell_6t
Xbit_r117_c25 bl[25] br[25] wl[117] vdd gnd cell_6t
Xbit_r118_c25 bl[25] br[25] wl[118] vdd gnd cell_6t
Xbit_r119_c25 bl[25] br[25] wl[119] vdd gnd cell_6t
Xbit_r120_c25 bl[25] br[25] wl[120] vdd gnd cell_6t
Xbit_r121_c25 bl[25] br[25] wl[121] vdd gnd cell_6t
Xbit_r122_c25 bl[25] br[25] wl[122] vdd gnd cell_6t
Xbit_r123_c25 bl[25] br[25] wl[123] vdd gnd cell_6t
Xbit_r124_c25 bl[25] br[25] wl[124] vdd gnd cell_6t
Xbit_r125_c25 bl[25] br[25] wl[125] vdd gnd cell_6t
Xbit_r126_c25 bl[25] br[25] wl[126] vdd gnd cell_6t
Xbit_r127_c25 bl[25] br[25] wl[127] vdd gnd cell_6t
Xbit_r128_c25 bl[25] br[25] wl[128] vdd gnd cell_6t
Xbit_r129_c25 bl[25] br[25] wl[129] vdd gnd cell_6t
Xbit_r130_c25 bl[25] br[25] wl[130] vdd gnd cell_6t
Xbit_r131_c25 bl[25] br[25] wl[131] vdd gnd cell_6t
Xbit_r132_c25 bl[25] br[25] wl[132] vdd gnd cell_6t
Xbit_r133_c25 bl[25] br[25] wl[133] vdd gnd cell_6t
Xbit_r134_c25 bl[25] br[25] wl[134] vdd gnd cell_6t
Xbit_r135_c25 bl[25] br[25] wl[135] vdd gnd cell_6t
Xbit_r136_c25 bl[25] br[25] wl[136] vdd gnd cell_6t
Xbit_r137_c25 bl[25] br[25] wl[137] vdd gnd cell_6t
Xbit_r138_c25 bl[25] br[25] wl[138] vdd gnd cell_6t
Xbit_r139_c25 bl[25] br[25] wl[139] vdd gnd cell_6t
Xbit_r140_c25 bl[25] br[25] wl[140] vdd gnd cell_6t
Xbit_r141_c25 bl[25] br[25] wl[141] vdd gnd cell_6t
Xbit_r142_c25 bl[25] br[25] wl[142] vdd gnd cell_6t
Xbit_r143_c25 bl[25] br[25] wl[143] vdd gnd cell_6t
Xbit_r144_c25 bl[25] br[25] wl[144] vdd gnd cell_6t
Xbit_r145_c25 bl[25] br[25] wl[145] vdd gnd cell_6t
Xbit_r146_c25 bl[25] br[25] wl[146] vdd gnd cell_6t
Xbit_r147_c25 bl[25] br[25] wl[147] vdd gnd cell_6t
Xbit_r148_c25 bl[25] br[25] wl[148] vdd gnd cell_6t
Xbit_r149_c25 bl[25] br[25] wl[149] vdd gnd cell_6t
Xbit_r150_c25 bl[25] br[25] wl[150] vdd gnd cell_6t
Xbit_r151_c25 bl[25] br[25] wl[151] vdd gnd cell_6t
Xbit_r152_c25 bl[25] br[25] wl[152] vdd gnd cell_6t
Xbit_r153_c25 bl[25] br[25] wl[153] vdd gnd cell_6t
Xbit_r154_c25 bl[25] br[25] wl[154] vdd gnd cell_6t
Xbit_r155_c25 bl[25] br[25] wl[155] vdd gnd cell_6t
Xbit_r156_c25 bl[25] br[25] wl[156] vdd gnd cell_6t
Xbit_r157_c25 bl[25] br[25] wl[157] vdd gnd cell_6t
Xbit_r158_c25 bl[25] br[25] wl[158] vdd gnd cell_6t
Xbit_r159_c25 bl[25] br[25] wl[159] vdd gnd cell_6t
Xbit_r160_c25 bl[25] br[25] wl[160] vdd gnd cell_6t
Xbit_r161_c25 bl[25] br[25] wl[161] vdd gnd cell_6t
Xbit_r162_c25 bl[25] br[25] wl[162] vdd gnd cell_6t
Xbit_r163_c25 bl[25] br[25] wl[163] vdd gnd cell_6t
Xbit_r164_c25 bl[25] br[25] wl[164] vdd gnd cell_6t
Xbit_r165_c25 bl[25] br[25] wl[165] vdd gnd cell_6t
Xbit_r166_c25 bl[25] br[25] wl[166] vdd gnd cell_6t
Xbit_r167_c25 bl[25] br[25] wl[167] vdd gnd cell_6t
Xbit_r168_c25 bl[25] br[25] wl[168] vdd gnd cell_6t
Xbit_r169_c25 bl[25] br[25] wl[169] vdd gnd cell_6t
Xbit_r170_c25 bl[25] br[25] wl[170] vdd gnd cell_6t
Xbit_r171_c25 bl[25] br[25] wl[171] vdd gnd cell_6t
Xbit_r172_c25 bl[25] br[25] wl[172] vdd gnd cell_6t
Xbit_r173_c25 bl[25] br[25] wl[173] vdd gnd cell_6t
Xbit_r174_c25 bl[25] br[25] wl[174] vdd gnd cell_6t
Xbit_r175_c25 bl[25] br[25] wl[175] vdd gnd cell_6t
Xbit_r176_c25 bl[25] br[25] wl[176] vdd gnd cell_6t
Xbit_r177_c25 bl[25] br[25] wl[177] vdd gnd cell_6t
Xbit_r178_c25 bl[25] br[25] wl[178] vdd gnd cell_6t
Xbit_r179_c25 bl[25] br[25] wl[179] vdd gnd cell_6t
Xbit_r180_c25 bl[25] br[25] wl[180] vdd gnd cell_6t
Xbit_r181_c25 bl[25] br[25] wl[181] vdd gnd cell_6t
Xbit_r182_c25 bl[25] br[25] wl[182] vdd gnd cell_6t
Xbit_r183_c25 bl[25] br[25] wl[183] vdd gnd cell_6t
Xbit_r184_c25 bl[25] br[25] wl[184] vdd gnd cell_6t
Xbit_r185_c25 bl[25] br[25] wl[185] vdd gnd cell_6t
Xbit_r186_c25 bl[25] br[25] wl[186] vdd gnd cell_6t
Xbit_r187_c25 bl[25] br[25] wl[187] vdd gnd cell_6t
Xbit_r188_c25 bl[25] br[25] wl[188] vdd gnd cell_6t
Xbit_r189_c25 bl[25] br[25] wl[189] vdd gnd cell_6t
Xbit_r190_c25 bl[25] br[25] wl[190] vdd gnd cell_6t
Xbit_r191_c25 bl[25] br[25] wl[191] vdd gnd cell_6t
Xbit_r192_c25 bl[25] br[25] wl[192] vdd gnd cell_6t
Xbit_r193_c25 bl[25] br[25] wl[193] vdd gnd cell_6t
Xbit_r194_c25 bl[25] br[25] wl[194] vdd gnd cell_6t
Xbit_r195_c25 bl[25] br[25] wl[195] vdd gnd cell_6t
Xbit_r196_c25 bl[25] br[25] wl[196] vdd gnd cell_6t
Xbit_r197_c25 bl[25] br[25] wl[197] vdd gnd cell_6t
Xbit_r198_c25 bl[25] br[25] wl[198] vdd gnd cell_6t
Xbit_r199_c25 bl[25] br[25] wl[199] vdd gnd cell_6t
Xbit_r200_c25 bl[25] br[25] wl[200] vdd gnd cell_6t
Xbit_r201_c25 bl[25] br[25] wl[201] vdd gnd cell_6t
Xbit_r202_c25 bl[25] br[25] wl[202] vdd gnd cell_6t
Xbit_r203_c25 bl[25] br[25] wl[203] vdd gnd cell_6t
Xbit_r204_c25 bl[25] br[25] wl[204] vdd gnd cell_6t
Xbit_r205_c25 bl[25] br[25] wl[205] vdd gnd cell_6t
Xbit_r206_c25 bl[25] br[25] wl[206] vdd gnd cell_6t
Xbit_r207_c25 bl[25] br[25] wl[207] vdd gnd cell_6t
Xbit_r208_c25 bl[25] br[25] wl[208] vdd gnd cell_6t
Xbit_r209_c25 bl[25] br[25] wl[209] vdd gnd cell_6t
Xbit_r210_c25 bl[25] br[25] wl[210] vdd gnd cell_6t
Xbit_r211_c25 bl[25] br[25] wl[211] vdd gnd cell_6t
Xbit_r212_c25 bl[25] br[25] wl[212] vdd gnd cell_6t
Xbit_r213_c25 bl[25] br[25] wl[213] vdd gnd cell_6t
Xbit_r214_c25 bl[25] br[25] wl[214] vdd gnd cell_6t
Xbit_r215_c25 bl[25] br[25] wl[215] vdd gnd cell_6t
Xbit_r216_c25 bl[25] br[25] wl[216] vdd gnd cell_6t
Xbit_r217_c25 bl[25] br[25] wl[217] vdd gnd cell_6t
Xbit_r218_c25 bl[25] br[25] wl[218] vdd gnd cell_6t
Xbit_r219_c25 bl[25] br[25] wl[219] vdd gnd cell_6t
Xbit_r220_c25 bl[25] br[25] wl[220] vdd gnd cell_6t
Xbit_r221_c25 bl[25] br[25] wl[221] vdd gnd cell_6t
Xbit_r222_c25 bl[25] br[25] wl[222] vdd gnd cell_6t
Xbit_r223_c25 bl[25] br[25] wl[223] vdd gnd cell_6t
Xbit_r224_c25 bl[25] br[25] wl[224] vdd gnd cell_6t
Xbit_r225_c25 bl[25] br[25] wl[225] vdd gnd cell_6t
Xbit_r226_c25 bl[25] br[25] wl[226] vdd gnd cell_6t
Xbit_r227_c25 bl[25] br[25] wl[227] vdd gnd cell_6t
Xbit_r228_c25 bl[25] br[25] wl[228] vdd gnd cell_6t
Xbit_r229_c25 bl[25] br[25] wl[229] vdd gnd cell_6t
Xbit_r230_c25 bl[25] br[25] wl[230] vdd gnd cell_6t
Xbit_r231_c25 bl[25] br[25] wl[231] vdd gnd cell_6t
Xbit_r232_c25 bl[25] br[25] wl[232] vdd gnd cell_6t
Xbit_r233_c25 bl[25] br[25] wl[233] vdd gnd cell_6t
Xbit_r234_c25 bl[25] br[25] wl[234] vdd gnd cell_6t
Xbit_r235_c25 bl[25] br[25] wl[235] vdd gnd cell_6t
Xbit_r236_c25 bl[25] br[25] wl[236] vdd gnd cell_6t
Xbit_r237_c25 bl[25] br[25] wl[237] vdd gnd cell_6t
Xbit_r238_c25 bl[25] br[25] wl[238] vdd gnd cell_6t
Xbit_r239_c25 bl[25] br[25] wl[239] vdd gnd cell_6t
Xbit_r240_c25 bl[25] br[25] wl[240] vdd gnd cell_6t
Xbit_r241_c25 bl[25] br[25] wl[241] vdd gnd cell_6t
Xbit_r242_c25 bl[25] br[25] wl[242] vdd gnd cell_6t
Xbit_r243_c25 bl[25] br[25] wl[243] vdd gnd cell_6t
Xbit_r244_c25 bl[25] br[25] wl[244] vdd gnd cell_6t
Xbit_r245_c25 bl[25] br[25] wl[245] vdd gnd cell_6t
Xbit_r246_c25 bl[25] br[25] wl[246] vdd gnd cell_6t
Xbit_r247_c25 bl[25] br[25] wl[247] vdd gnd cell_6t
Xbit_r248_c25 bl[25] br[25] wl[248] vdd gnd cell_6t
Xbit_r249_c25 bl[25] br[25] wl[249] vdd gnd cell_6t
Xbit_r250_c25 bl[25] br[25] wl[250] vdd gnd cell_6t
Xbit_r251_c25 bl[25] br[25] wl[251] vdd gnd cell_6t
Xbit_r252_c25 bl[25] br[25] wl[252] vdd gnd cell_6t
Xbit_r253_c25 bl[25] br[25] wl[253] vdd gnd cell_6t
Xbit_r254_c25 bl[25] br[25] wl[254] vdd gnd cell_6t
Xbit_r255_c25 bl[25] br[25] wl[255] vdd gnd cell_6t
Xbit_r256_c25 bl[25] br[25] wl[256] vdd gnd cell_6t
Xbit_r257_c25 bl[25] br[25] wl[257] vdd gnd cell_6t
Xbit_r258_c25 bl[25] br[25] wl[258] vdd gnd cell_6t
Xbit_r259_c25 bl[25] br[25] wl[259] vdd gnd cell_6t
Xbit_r260_c25 bl[25] br[25] wl[260] vdd gnd cell_6t
Xbit_r261_c25 bl[25] br[25] wl[261] vdd gnd cell_6t
Xbit_r262_c25 bl[25] br[25] wl[262] vdd gnd cell_6t
Xbit_r263_c25 bl[25] br[25] wl[263] vdd gnd cell_6t
Xbit_r264_c25 bl[25] br[25] wl[264] vdd gnd cell_6t
Xbit_r265_c25 bl[25] br[25] wl[265] vdd gnd cell_6t
Xbit_r266_c25 bl[25] br[25] wl[266] vdd gnd cell_6t
Xbit_r267_c25 bl[25] br[25] wl[267] vdd gnd cell_6t
Xbit_r268_c25 bl[25] br[25] wl[268] vdd gnd cell_6t
Xbit_r269_c25 bl[25] br[25] wl[269] vdd gnd cell_6t
Xbit_r270_c25 bl[25] br[25] wl[270] vdd gnd cell_6t
Xbit_r271_c25 bl[25] br[25] wl[271] vdd gnd cell_6t
Xbit_r272_c25 bl[25] br[25] wl[272] vdd gnd cell_6t
Xbit_r273_c25 bl[25] br[25] wl[273] vdd gnd cell_6t
Xbit_r274_c25 bl[25] br[25] wl[274] vdd gnd cell_6t
Xbit_r275_c25 bl[25] br[25] wl[275] vdd gnd cell_6t
Xbit_r276_c25 bl[25] br[25] wl[276] vdd gnd cell_6t
Xbit_r277_c25 bl[25] br[25] wl[277] vdd gnd cell_6t
Xbit_r278_c25 bl[25] br[25] wl[278] vdd gnd cell_6t
Xbit_r279_c25 bl[25] br[25] wl[279] vdd gnd cell_6t
Xbit_r280_c25 bl[25] br[25] wl[280] vdd gnd cell_6t
Xbit_r281_c25 bl[25] br[25] wl[281] vdd gnd cell_6t
Xbit_r282_c25 bl[25] br[25] wl[282] vdd gnd cell_6t
Xbit_r283_c25 bl[25] br[25] wl[283] vdd gnd cell_6t
Xbit_r284_c25 bl[25] br[25] wl[284] vdd gnd cell_6t
Xbit_r285_c25 bl[25] br[25] wl[285] vdd gnd cell_6t
Xbit_r286_c25 bl[25] br[25] wl[286] vdd gnd cell_6t
Xbit_r287_c25 bl[25] br[25] wl[287] vdd gnd cell_6t
Xbit_r288_c25 bl[25] br[25] wl[288] vdd gnd cell_6t
Xbit_r289_c25 bl[25] br[25] wl[289] vdd gnd cell_6t
Xbit_r290_c25 bl[25] br[25] wl[290] vdd gnd cell_6t
Xbit_r291_c25 bl[25] br[25] wl[291] vdd gnd cell_6t
Xbit_r292_c25 bl[25] br[25] wl[292] vdd gnd cell_6t
Xbit_r293_c25 bl[25] br[25] wl[293] vdd gnd cell_6t
Xbit_r294_c25 bl[25] br[25] wl[294] vdd gnd cell_6t
Xbit_r295_c25 bl[25] br[25] wl[295] vdd gnd cell_6t
Xbit_r296_c25 bl[25] br[25] wl[296] vdd gnd cell_6t
Xbit_r297_c25 bl[25] br[25] wl[297] vdd gnd cell_6t
Xbit_r298_c25 bl[25] br[25] wl[298] vdd gnd cell_6t
Xbit_r299_c25 bl[25] br[25] wl[299] vdd gnd cell_6t
Xbit_r300_c25 bl[25] br[25] wl[300] vdd gnd cell_6t
Xbit_r301_c25 bl[25] br[25] wl[301] vdd gnd cell_6t
Xbit_r302_c25 bl[25] br[25] wl[302] vdd gnd cell_6t
Xbit_r303_c25 bl[25] br[25] wl[303] vdd gnd cell_6t
Xbit_r304_c25 bl[25] br[25] wl[304] vdd gnd cell_6t
Xbit_r305_c25 bl[25] br[25] wl[305] vdd gnd cell_6t
Xbit_r306_c25 bl[25] br[25] wl[306] vdd gnd cell_6t
Xbit_r307_c25 bl[25] br[25] wl[307] vdd gnd cell_6t
Xbit_r308_c25 bl[25] br[25] wl[308] vdd gnd cell_6t
Xbit_r309_c25 bl[25] br[25] wl[309] vdd gnd cell_6t
Xbit_r310_c25 bl[25] br[25] wl[310] vdd gnd cell_6t
Xbit_r311_c25 bl[25] br[25] wl[311] vdd gnd cell_6t
Xbit_r312_c25 bl[25] br[25] wl[312] vdd gnd cell_6t
Xbit_r313_c25 bl[25] br[25] wl[313] vdd gnd cell_6t
Xbit_r314_c25 bl[25] br[25] wl[314] vdd gnd cell_6t
Xbit_r315_c25 bl[25] br[25] wl[315] vdd gnd cell_6t
Xbit_r316_c25 bl[25] br[25] wl[316] vdd gnd cell_6t
Xbit_r317_c25 bl[25] br[25] wl[317] vdd gnd cell_6t
Xbit_r318_c25 bl[25] br[25] wl[318] vdd gnd cell_6t
Xbit_r319_c25 bl[25] br[25] wl[319] vdd gnd cell_6t
Xbit_r320_c25 bl[25] br[25] wl[320] vdd gnd cell_6t
Xbit_r321_c25 bl[25] br[25] wl[321] vdd gnd cell_6t
Xbit_r322_c25 bl[25] br[25] wl[322] vdd gnd cell_6t
Xbit_r323_c25 bl[25] br[25] wl[323] vdd gnd cell_6t
Xbit_r324_c25 bl[25] br[25] wl[324] vdd gnd cell_6t
Xbit_r325_c25 bl[25] br[25] wl[325] vdd gnd cell_6t
Xbit_r326_c25 bl[25] br[25] wl[326] vdd gnd cell_6t
Xbit_r327_c25 bl[25] br[25] wl[327] vdd gnd cell_6t
Xbit_r328_c25 bl[25] br[25] wl[328] vdd gnd cell_6t
Xbit_r329_c25 bl[25] br[25] wl[329] vdd gnd cell_6t
Xbit_r330_c25 bl[25] br[25] wl[330] vdd gnd cell_6t
Xbit_r331_c25 bl[25] br[25] wl[331] vdd gnd cell_6t
Xbit_r332_c25 bl[25] br[25] wl[332] vdd gnd cell_6t
Xbit_r333_c25 bl[25] br[25] wl[333] vdd gnd cell_6t
Xbit_r334_c25 bl[25] br[25] wl[334] vdd gnd cell_6t
Xbit_r335_c25 bl[25] br[25] wl[335] vdd gnd cell_6t
Xbit_r336_c25 bl[25] br[25] wl[336] vdd gnd cell_6t
Xbit_r337_c25 bl[25] br[25] wl[337] vdd gnd cell_6t
Xbit_r338_c25 bl[25] br[25] wl[338] vdd gnd cell_6t
Xbit_r339_c25 bl[25] br[25] wl[339] vdd gnd cell_6t
Xbit_r340_c25 bl[25] br[25] wl[340] vdd gnd cell_6t
Xbit_r341_c25 bl[25] br[25] wl[341] vdd gnd cell_6t
Xbit_r342_c25 bl[25] br[25] wl[342] vdd gnd cell_6t
Xbit_r343_c25 bl[25] br[25] wl[343] vdd gnd cell_6t
Xbit_r344_c25 bl[25] br[25] wl[344] vdd gnd cell_6t
Xbit_r345_c25 bl[25] br[25] wl[345] vdd gnd cell_6t
Xbit_r346_c25 bl[25] br[25] wl[346] vdd gnd cell_6t
Xbit_r347_c25 bl[25] br[25] wl[347] vdd gnd cell_6t
Xbit_r348_c25 bl[25] br[25] wl[348] vdd gnd cell_6t
Xbit_r349_c25 bl[25] br[25] wl[349] vdd gnd cell_6t
Xbit_r350_c25 bl[25] br[25] wl[350] vdd gnd cell_6t
Xbit_r351_c25 bl[25] br[25] wl[351] vdd gnd cell_6t
Xbit_r352_c25 bl[25] br[25] wl[352] vdd gnd cell_6t
Xbit_r353_c25 bl[25] br[25] wl[353] vdd gnd cell_6t
Xbit_r354_c25 bl[25] br[25] wl[354] vdd gnd cell_6t
Xbit_r355_c25 bl[25] br[25] wl[355] vdd gnd cell_6t
Xbit_r356_c25 bl[25] br[25] wl[356] vdd gnd cell_6t
Xbit_r357_c25 bl[25] br[25] wl[357] vdd gnd cell_6t
Xbit_r358_c25 bl[25] br[25] wl[358] vdd gnd cell_6t
Xbit_r359_c25 bl[25] br[25] wl[359] vdd gnd cell_6t
Xbit_r360_c25 bl[25] br[25] wl[360] vdd gnd cell_6t
Xbit_r361_c25 bl[25] br[25] wl[361] vdd gnd cell_6t
Xbit_r362_c25 bl[25] br[25] wl[362] vdd gnd cell_6t
Xbit_r363_c25 bl[25] br[25] wl[363] vdd gnd cell_6t
Xbit_r364_c25 bl[25] br[25] wl[364] vdd gnd cell_6t
Xbit_r365_c25 bl[25] br[25] wl[365] vdd gnd cell_6t
Xbit_r366_c25 bl[25] br[25] wl[366] vdd gnd cell_6t
Xbit_r367_c25 bl[25] br[25] wl[367] vdd gnd cell_6t
Xbit_r368_c25 bl[25] br[25] wl[368] vdd gnd cell_6t
Xbit_r369_c25 bl[25] br[25] wl[369] vdd gnd cell_6t
Xbit_r370_c25 bl[25] br[25] wl[370] vdd gnd cell_6t
Xbit_r371_c25 bl[25] br[25] wl[371] vdd gnd cell_6t
Xbit_r372_c25 bl[25] br[25] wl[372] vdd gnd cell_6t
Xbit_r373_c25 bl[25] br[25] wl[373] vdd gnd cell_6t
Xbit_r374_c25 bl[25] br[25] wl[374] vdd gnd cell_6t
Xbit_r375_c25 bl[25] br[25] wl[375] vdd gnd cell_6t
Xbit_r376_c25 bl[25] br[25] wl[376] vdd gnd cell_6t
Xbit_r377_c25 bl[25] br[25] wl[377] vdd gnd cell_6t
Xbit_r378_c25 bl[25] br[25] wl[378] vdd gnd cell_6t
Xbit_r379_c25 bl[25] br[25] wl[379] vdd gnd cell_6t
Xbit_r380_c25 bl[25] br[25] wl[380] vdd gnd cell_6t
Xbit_r381_c25 bl[25] br[25] wl[381] vdd gnd cell_6t
Xbit_r382_c25 bl[25] br[25] wl[382] vdd gnd cell_6t
Xbit_r383_c25 bl[25] br[25] wl[383] vdd gnd cell_6t
Xbit_r384_c25 bl[25] br[25] wl[384] vdd gnd cell_6t
Xbit_r385_c25 bl[25] br[25] wl[385] vdd gnd cell_6t
Xbit_r386_c25 bl[25] br[25] wl[386] vdd gnd cell_6t
Xbit_r387_c25 bl[25] br[25] wl[387] vdd gnd cell_6t
Xbit_r388_c25 bl[25] br[25] wl[388] vdd gnd cell_6t
Xbit_r389_c25 bl[25] br[25] wl[389] vdd gnd cell_6t
Xbit_r390_c25 bl[25] br[25] wl[390] vdd gnd cell_6t
Xbit_r391_c25 bl[25] br[25] wl[391] vdd gnd cell_6t
Xbit_r392_c25 bl[25] br[25] wl[392] vdd gnd cell_6t
Xbit_r393_c25 bl[25] br[25] wl[393] vdd gnd cell_6t
Xbit_r394_c25 bl[25] br[25] wl[394] vdd gnd cell_6t
Xbit_r395_c25 bl[25] br[25] wl[395] vdd gnd cell_6t
Xbit_r396_c25 bl[25] br[25] wl[396] vdd gnd cell_6t
Xbit_r397_c25 bl[25] br[25] wl[397] vdd gnd cell_6t
Xbit_r398_c25 bl[25] br[25] wl[398] vdd gnd cell_6t
Xbit_r399_c25 bl[25] br[25] wl[399] vdd gnd cell_6t
Xbit_r400_c25 bl[25] br[25] wl[400] vdd gnd cell_6t
Xbit_r401_c25 bl[25] br[25] wl[401] vdd gnd cell_6t
Xbit_r402_c25 bl[25] br[25] wl[402] vdd gnd cell_6t
Xbit_r403_c25 bl[25] br[25] wl[403] vdd gnd cell_6t
Xbit_r404_c25 bl[25] br[25] wl[404] vdd gnd cell_6t
Xbit_r405_c25 bl[25] br[25] wl[405] vdd gnd cell_6t
Xbit_r406_c25 bl[25] br[25] wl[406] vdd gnd cell_6t
Xbit_r407_c25 bl[25] br[25] wl[407] vdd gnd cell_6t
Xbit_r408_c25 bl[25] br[25] wl[408] vdd gnd cell_6t
Xbit_r409_c25 bl[25] br[25] wl[409] vdd gnd cell_6t
Xbit_r410_c25 bl[25] br[25] wl[410] vdd gnd cell_6t
Xbit_r411_c25 bl[25] br[25] wl[411] vdd gnd cell_6t
Xbit_r412_c25 bl[25] br[25] wl[412] vdd gnd cell_6t
Xbit_r413_c25 bl[25] br[25] wl[413] vdd gnd cell_6t
Xbit_r414_c25 bl[25] br[25] wl[414] vdd gnd cell_6t
Xbit_r415_c25 bl[25] br[25] wl[415] vdd gnd cell_6t
Xbit_r416_c25 bl[25] br[25] wl[416] vdd gnd cell_6t
Xbit_r417_c25 bl[25] br[25] wl[417] vdd gnd cell_6t
Xbit_r418_c25 bl[25] br[25] wl[418] vdd gnd cell_6t
Xbit_r419_c25 bl[25] br[25] wl[419] vdd gnd cell_6t
Xbit_r420_c25 bl[25] br[25] wl[420] vdd gnd cell_6t
Xbit_r421_c25 bl[25] br[25] wl[421] vdd gnd cell_6t
Xbit_r422_c25 bl[25] br[25] wl[422] vdd gnd cell_6t
Xbit_r423_c25 bl[25] br[25] wl[423] vdd gnd cell_6t
Xbit_r424_c25 bl[25] br[25] wl[424] vdd gnd cell_6t
Xbit_r425_c25 bl[25] br[25] wl[425] vdd gnd cell_6t
Xbit_r426_c25 bl[25] br[25] wl[426] vdd gnd cell_6t
Xbit_r427_c25 bl[25] br[25] wl[427] vdd gnd cell_6t
Xbit_r428_c25 bl[25] br[25] wl[428] vdd gnd cell_6t
Xbit_r429_c25 bl[25] br[25] wl[429] vdd gnd cell_6t
Xbit_r430_c25 bl[25] br[25] wl[430] vdd gnd cell_6t
Xbit_r431_c25 bl[25] br[25] wl[431] vdd gnd cell_6t
Xbit_r432_c25 bl[25] br[25] wl[432] vdd gnd cell_6t
Xbit_r433_c25 bl[25] br[25] wl[433] vdd gnd cell_6t
Xbit_r434_c25 bl[25] br[25] wl[434] vdd gnd cell_6t
Xbit_r435_c25 bl[25] br[25] wl[435] vdd gnd cell_6t
Xbit_r436_c25 bl[25] br[25] wl[436] vdd gnd cell_6t
Xbit_r437_c25 bl[25] br[25] wl[437] vdd gnd cell_6t
Xbit_r438_c25 bl[25] br[25] wl[438] vdd gnd cell_6t
Xbit_r439_c25 bl[25] br[25] wl[439] vdd gnd cell_6t
Xbit_r440_c25 bl[25] br[25] wl[440] vdd gnd cell_6t
Xbit_r441_c25 bl[25] br[25] wl[441] vdd gnd cell_6t
Xbit_r442_c25 bl[25] br[25] wl[442] vdd gnd cell_6t
Xbit_r443_c25 bl[25] br[25] wl[443] vdd gnd cell_6t
Xbit_r444_c25 bl[25] br[25] wl[444] vdd gnd cell_6t
Xbit_r445_c25 bl[25] br[25] wl[445] vdd gnd cell_6t
Xbit_r446_c25 bl[25] br[25] wl[446] vdd gnd cell_6t
Xbit_r447_c25 bl[25] br[25] wl[447] vdd gnd cell_6t
Xbit_r448_c25 bl[25] br[25] wl[448] vdd gnd cell_6t
Xbit_r449_c25 bl[25] br[25] wl[449] vdd gnd cell_6t
Xbit_r450_c25 bl[25] br[25] wl[450] vdd gnd cell_6t
Xbit_r451_c25 bl[25] br[25] wl[451] vdd gnd cell_6t
Xbit_r452_c25 bl[25] br[25] wl[452] vdd gnd cell_6t
Xbit_r453_c25 bl[25] br[25] wl[453] vdd gnd cell_6t
Xbit_r454_c25 bl[25] br[25] wl[454] vdd gnd cell_6t
Xbit_r455_c25 bl[25] br[25] wl[455] vdd gnd cell_6t
Xbit_r456_c25 bl[25] br[25] wl[456] vdd gnd cell_6t
Xbit_r457_c25 bl[25] br[25] wl[457] vdd gnd cell_6t
Xbit_r458_c25 bl[25] br[25] wl[458] vdd gnd cell_6t
Xbit_r459_c25 bl[25] br[25] wl[459] vdd gnd cell_6t
Xbit_r460_c25 bl[25] br[25] wl[460] vdd gnd cell_6t
Xbit_r461_c25 bl[25] br[25] wl[461] vdd gnd cell_6t
Xbit_r462_c25 bl[25] br[25] wl[462] vdd gnd cell_6t
Xbit_r463_c25 bl[25] br[25] wl[463] vdd gnd cell_6t
Xbit_r464_c25 bl[25] br[25] wl[464] vdd gnd cell_6t
Xbit_r465_c25 bl[25] br[25] wl[465] vdd gnd cell_6t
Xbit_r466_c25 bl[25] br[25] wl[466] vdd gnd cell_6t
Xbit_r467_c25 bl[25] br[25] wl[467] vdd gnd cell_6t
Xbit_r468_c25 bl[25] br[25] wl[468] vdd gnd cell_6t
Xbit_r469_c25 bl[25] br[25] wl[469] vdd gnd cell_6t
Xbit_r470_c25 bl[25] br[25] wl[470] vdd gnd cell_6t
Xbit_r471_c25 bl[25] br[25] wl[471] vdd gnd cell_6t
Xbit_r472_c25 bl[25] br[25] wl[472] vdd gnd cell_6t
Xbit_r473_c25 bl[25] br[25] wl[473] vdd gnd cell_6t
Xbit_r474_c25 bl[25] br[25] wl[474] vdd gnd cell_6t
Xbit_r475_c25 bl[25] br[25] wl[475] vdd gnd cell_6t
Xbit_r476_c25 bl[25] br[25] wl[476] vdd gnd cell_6t
Xbit_r477_c25 bl[25] br[25] wl[477] vdd gnd cell_6t
Xbit_r478_c25 bl[25] br[25] wl[478] vdd gnd cell_6t
Xbit_r479_c25 bl[25] br[25] wl[479] vdd gnd cell_6t
Xbit_r480_c25 bl[25] br[25] wl[480] vdd gnd cell_6t
Xbit_r481_c25 bl[25] br[25] wl[481] vdd gnd cell_6t
Xbit_r482_c25 bl[25] br[25] wl[482] vdd gnd cell_6t
Xbit_r483_c25 bl[25] br[25] wl[483] vdd gnd cell_6t
Xbit_r484_c25 bl[25] br[25] wl[484] vdd gnd cell_6t
Xbit_r485_c25 bl[25] br[25] wl[485] vdd gnd cell_6t
Xbit_r486_c25 bl[25] br[25] wl[486] vdd gnd cell_6t
Xbit_r487_c25 bl[25] br[25] wl[487] vdd gnd cell_6t
Xbit_r488_c25 bl[25] br[25] wl[488] vdd gnd cell_6t
Xbit_r489_c25 bl[25] br[25] wl[489] vdd gnd cell_6t
Xbit_r490_c25 bl[25] br[25] wl[490] vdd gnd cell_6t
Xbit_r491_c25 bl[25] br[25] wl[491] vdd gnd cell_6t
Xbit_r492_c25 bl[25] br[25] wl[492] vdd gnd cell_6t
Xbit_r493_c25 bl[25] br[25] wl[493] vdd gnd cell_6t
Xbit_r494_c25 bl[25] br[25] wl[494] vdd gnd cell_6t
Xbit_r495_c25 bl[25] br[25] wl[495] vdd gnd cell_6t
Xbit_r496_c25 bl[25] br[25] wl[496] vdd gnd cell_6t
Xbit_r497_c25 bl[25] br[25] wl[497] vdd gnd cell_6t
Xbit_r498_c25 bl[25] br[25] wl[498] vdd gnd cell_6t
Xbit_r499_c25 bl[25] br[25] wl[499] vdd gnd cell_6t
Xbit_r500_c25 bl[25] br[25] wl[500] vdd gnd cell_6t
Xbit_r501_c25 bl[25] br[25] wl[501] vdd gnd cell_6t
Xbit_r502_c25 bl[25] br[25] wl[502] vdd gnd cell_6t
Xbit_r503_c25 bl[25] br[25] wl[503] vdd gnd cell_6t
Xbit_r504_c25 bl[25] br[25] wl[504] vdd gnd cell_6t
Xbit_r505_c25 bl[25] br[25] wl[505] vdd gnd cell_6t
Xbit_r506_c25 bl[25] br[25] wl[506] vdd gnd cell_6t
Xbit_r507_c25 bl[25] br[25] wl[507] vdd gnd cell_6t
Xbit_r508_c25 bl[25] br[25] wl[508] vdd gnd cell_6t
Xbit_r509_c25 bl[25] br[25] wl[509] vdd gnd cell_6t
Xbit_r510_c25 bl[25] br[25] wl[510] vdd gnd cell_6t
Xbit_r511_c25 bl[25] br[25] wl[511] vdd gnd cell_6t
Xbit_r0_c26 bl[26] br[26] wl[0] vdd gnd cell_6t
Xbit_r1_c26 bl[26] br[26] wl[1] vdd gnd cell_6t
Xbit_r2_c26 bl[26] br[26] wl[2] vdd gnd cell_6t
Xbit_r3_c26 bl[26] br[26] wl[3] vdd gnd cell_6t
Xbit_r4_c26 bl[26] br[26] wl[4] vdd gnd cell_6t
Xbit_r5_c26 bl[26] br[26] wl[5] vdd gnd cell_6t
Xbit_r6_c26 bl[26] br[26] wl[6] vdd gnd cell_6t
Xbit_r7_c26 bl[26] br[26] wl[7] vdd gnd cell_6t
Xbit_r8_c26 bl[26] br[26] wl[8] vdd gnd cell_6t
Xbit_r9_c26 bl[26] br[26] wl[9] vdd gnd cell_6t
Xbit_r10_c26 bl[26] br[26] wl[10] vdd gnd cell_6t
Xbit_r11_c26 bl[26] br[26] wl[11] vdd gnd cell_6t
Xbit_r12_c26 bl[26] br[26] wl[12] vdd gnd cell_6t
Xbit_r13_c26 bl[26] br[26] wl[13] vdd gnd cell_6t
Xbit_r14_c26 bl[26] br[26] wl[14] vdd gnd cell_6t
Xbit_r15_c26 bl[26] br[26] wl[15] vdd gnd cell_6t
Xbit_r16_c26 bl[26] br[26] wl[16] vdd gnd cell_6t
Xbit_r17_c26 bl[26] br[26] wl[17] vdd gnd cell_6t
Xbit_r18_c26 bl[26] br[26] wl[18] vdd gnd cell_6t
Xbit_r19_c26 bl[26] br[26] wl[19] vdd gnd cell_6t
Xbit_r20_c26 bl[26] br[26] wl[20] vdd gnd cell_6t
Xbit_r21_c26 bl[26] br[26] wl[21] vdd gnd cell_6t
Xbit_r22_c26 bl[26] br[26] wl[22] vdd gnd cell_6t
Xbit_r23_c26 bl[26] br[26] wl[23] vdd gnd cell_6t
Xbit_r24_c26 bl[26] br[26] wl[24] vdd gnd cell_6t
Xbit_r25_c26 bl[26] br[26] wl[25] vdd gnd cell_6t
Xbit_r26_c26 bl[26] br[26] wl[26] vdd gnd cell_6t
Xbit_r27_c26 bl[26] br[26] wl[27] vdd gnd cell_6t
Xbit_r28_c26 bl[26] br[26] wl[28] vdd gnd cell_6t
Xbit_r29_c26 bl[26] br[26] wl[29] vdd gnd cell_6t
Xbit_r30_c26 bl[26] br[26] wl[30] vdd gnd cell_6t
Xbit_r31_c26 bl[26] br[26] wl[31] vdd gnd cell_6t
Xbit_r32_c26 bl[26] br[26] wl[32] vdd gnd cell_6t
Xbit_r33_c26 bl[26] br[26] wl[33] vdd gnd cell_6t
Xbit_r34_c26 bl[26] br[26] wl[34] vdd gnd cell_6t
Xbit_r35_c26 bl[26] br[26] wl[35] vdd gnd cell_6t
Xbit_r36_c26 bl[26] br[26] wl[36] vdd gnd cell_6t
Xbit_r37_c26 bl[26] br[26] wl[37] vdd gnd cell_6t
Xbit_r38_c26 bl[26] br[26] wl[38] vdd gnd cell_6t
Xbit_r39_c26 bl[26] br[26] wl[39] vdd gnd cell_6t
Xbit_r40_c26 bl[26] br[26] wl[40] vdd gnd cell_6t
Xbit_r41_c26 bl[26] br[26] wl[41] vdd gnd cell_6t
Xbit_r42_c26 bl[26] br[26] wl[42] vdd gnd cell_6t
Xbit_r43_c26 bl[26] br[26] wl[43] vdd gnd cell_6t
Xbit_r44_c26 bl[26] br[26] wl[44] vdd gnd cell_6t
Xbit_r45_c26 bl[26] br[26] wl[45] vdd gnd cell_6t
Xbit_r46_c26 bl[26] br[26] wl[46] vdd gnd cell_6t
Xbit_r47_c26 bl[26] br[26] wl[47] vdd gnd cell_6t
Xbit_r48_c26 bl[26] br[26] wl[48] vdd gnd cell_6t
Xbit_r49_c26 bl[26] br[26] wl[49] vdd gnd cell_6t
Xbit_r50_c26 bl[26] br[26] wl[50] vdd gnd cell_6t
Xbit_r51_c26 bl[26] br[26] wl[51] vdd gnd cell_6t
Xbit_r52_c26 bl[26] br[26] wl[52] vdd gnd cell_6t
Xbit_r53_c26 bl[26] br[26] wl[53] vdd gnd cell_6t
Xbit_r54_c26 bl[26] br[26] wl[54] vdd gnd cell_6t
Xbit_r55_c26 bl[26] br[26] wl[55] vdd gnd cell_6t
Xbit_r56_c26 bl[26] br[26] wl[56] vdd gnd cell_6t
Xbit_r57_c26 bl[26] br[26] wl[57] vdd gnd cell_6t
Xbit_r58_c26 bl[26] br[26] wl[58] vdd gnd cell_6t
Xbit_r59_c26 bl[26] br[26] wl[59] vdd gnd cell_6t
Xbit_r60_c26 bl[26] br[26] wl[60] vdd gnd cell_6t
Xbit_r61_c26 bl[26] br[26] wl[61] vdd gnd cell_6t
Xbit_r62_c26 bl[26] br[26] wl[62] vdd gnd cell_6t
Xbit_r63_c26 bl[26] br[26] wl[63] vdd gnd cell_6t
Xbit_r64_c26 bl[26] br[26] wl[64] vdd gnd cell_6t
Xbit_r65_c26 bl[26] br[26] wl[65] vdd gnd cell_6t
Xbit_r66_c26 bl[26] br[26] wl[66] vdd gnd cell_6t
Xbit_r67_c26 bl[26] br[26] wl[67] vdd gnd cell_6t
Xbit_r68_c26 bl[26] br[26] wl[68] vdd gnd cell_6t
Xbit_r69_c26 bl[26] br[26] wl[69] vdd gnd cell_6t
Xbit_r70_c26 bl[26] br[26] wl[70] vdd gnd cell_6t
Xbit_r71_c26 bl[26] br[26] wl[71] vdd gnd cell_6t
Xbit_r72_c26 bl[26] br[26] wl[72] vdd gnd cell_6t
Xbit_r73_c26 bl[26] br[26] wl[73] vdd gnd cell_6t
Xbit_r74_c26 bl[26] br[26] wl[74] vdd gnd cell_6t
Xbit_r75_c26 bl[26] br[26] wl[75] vdd gnd cell_6t
Xbit_r76_c26 bl[26] br[26] wl[76] vdd gnd cell_6t
Xbit_r77_c26 bl[26] br[26] wl[77] vdd gnd cell_6t
Xbit_r78_c26 bl[26] br[26] wl[78] vdd gnd cell_6t
Xbit_r79_c26 bl[26] br[26] wl[79] vdd gnd cell_6t
Xbit_r80_c26 bl[26] br[26] wl[80] vdd gnd cell_6t
Xbit_r81_c26 bl[26] br[26] wl[81] vdd gnd cell_6t
Xbit_r82_c26 bl[26] br[26] wl[82] vdd gnd cell_6t
Xbit_r83_c26 bl[26] br[26] wl[83] vdd gnd cell_6t
Xbit_r84_c26 bl[26] br[26] wl[84] vdd gnd cell_6t
Xbit_r85_c26 bl[26] br[26] wl[85] vdd gnd cell_6t
Xbit_r86_c26 bl[26] br[26] wl[86] vdd gnd cell_6t
Xbit_r87_c26 bl[26] br[26] wl[87] vdd gnd cell_6t
Xbit_r88_c26 bl[26] br[26] wl[88] vdd gnd cell_6t
Xbit_r89_c26 bl[26] br[26] wl[89] vdd gnd cell_6t
Xbit_r90_c26 bl[26] br[26] wl[90] vdd gnd cell_6t
Xbit_r91_c26 bl[26] br[26] wl[91] vdd gnd cell_6t
Xbit_r92_c26 bl[26] br[26] wl[92] vdd gnd cell_6t
Xbit_r93_c26 bl[26] br[26] wl[93] vdd gnd cell_6t
Xbit_r94_c26 bl[26] br[26] wl[94] vdd gnd cell_6t
Xbit_r95_c26 bl[26] br[26] wl[95] vdd gnd cell_6t
Xbit_r96_c26 bl[26] br[26] wl[96] vdd gnd cell_6t
Xbit_r97_c26 bl[26] br[26] wl[97] vdd gnd cell_6t
Xbit_r98_c26 bl[26] br[26] wl[98] vdd gnd cell_6t
Xbit_r99_c26 bl[26] br[26] wl[99] vdd gnd cell_6t
Xbit_r100_c26 bl[26] br[26] wl[100] vdd gnd cell_6t
Xbit_r101_c26 bl[26] br[26] wl[101] vdd gnd cell_6t
Xbit_r102_c26 bl[26] br[26] wl[102] vdd gnd cell_6t
Xbit_r103_c26 bl[26] br[26] wl[103] vdd gnd cell_6t
Xbit_r104_c26 bl[26] br[26] wl[104] vdd gnd cell_6t
Xbit_r105_c26 bl[26] br[26] wl[105] vdd gnd cell_6t
Xbit_r106_c26 bl[26] br[26] wl[106] vdd gnd cell_6t
Xbit_r107_c26 bl[26] br[26] wl[107] vdd gnd cell_6t
Xbit_r108_c26 bl[26] br[26] wl[108] vdd gnd cell_6t
Xbit_r109_c26 bl[26] br[26] wl[109] vdd gnd cell_6t
Xbit_r110_c26 bl[26] br[26] wl[110] vdd gnd cell_6t
Xbit_r111_c26 bl[26] br[26] wl[111] vdd gnd cell_6t
Xbit_r112_c26 bl[26] br[26] wl[112] vdd gnd cell_6t
Xbit_r113_c26 bl[26] br[26] wl[113] vdd gnd cell_6t
Xbit_r114_c26 bl[26] br[26] wl[114] vdd gnd cell_6t
Xbit_r115_c26 bl[26] br[26] wl[115] vdd gnd cell_6t
Xbit_r116_c26 bl[26] br[26] wl[116] vdd gnd cell_6t
Xbit_r117_c26 bl[26] br[26] wl[117] vdd gnd cell_6t
Xbit_r118_c26 bl[26] br[26] wl[118] vdd gnd cell_6t
Xbit_r119_c26 bl[26] br[26] wl[119] vdd gnd cell_6t
Xbit_r120_c26 bl[26] br[26] wl[120] vdd gnd cell_6t
Xbit_r121_c26 bl[26] br[26] wl[121] vdd gnd cell_6t
Xbit_r122_c26 bl[26] br[26] wl[122] vdd gnd cell_6t
Xbit_r123_c26 bl[26] br[26] wl[123] vdd gnd cell_6t
Xbit_r124_c26 bl[26] br[26] wl[124] vdd gnd cell_6t
Xbit_r125_c26 bl[26] br[26] wl[125] vdd gnd cell_6t
Xbit_r126_c26 bl[26] br[26] wl[126] vdd gnd cell_6t
Xbit_r127_c26 bl[26] br[26] wl[127] vdd gnd cell_6t
Xbit_r128_c26 bl[26] br[26] wl[128] vdd gnd cell_6t
Xbit_r129_c26 bl[26] br[26] wl[129] vdd gnd cell_6t
Xbit_r130_c26 bl[26] br[26] wl[130] vdd gnd cell_6t
Xbit_r131_c26 bl[26] br[26] wl[131] vdd gnd cell_6t
Xbit_r132_c26 bl[26] br[26] wl[132] vdd gnd cell_6t
Xbit_r133_c26 bl[26] br[26] wl[133] vdd gnd cell_6t
Xbit_r134_c26 bl[26] br[26] wl[134] vdd gnd cell_6t
Xbit_r135_c26 bl[26] br[26] wl[135] vdd gnd cell_6t
Xbit_r136_c26 bl[26] br[26] wl[136] vdd gnd cell_6t
Xbit_r137_c26 bl[26] br[26] wl[137] vdd gnd cell_6t
Xbit_r138_c26 bl[26] br[26] wl[138] vdd gnd cell_6t
Xbit_r139_c26 bl[26] br[26] wl[139] vdd gnd cell_6t
Xbit_r140_c26 bl[26] br[26] wl[140] vdd gnd cell_6t
Xbit_r141_c26 bl[26] br[26] wl[141] vdd gnd cell_6t
Xbit_r142_c26 bl[26] br[26] wl[142] vdd gnd cell_6t
Xbit_r143_c26 bl[26] br[26] wl[143] vdd gnd cell_6t
Xbit_r144_c26 bl[26] br[26] wl[144] vdd gnd cell_6t
Xbit_r145_c26 bl[26] br[26] wl[145] vdd gnd cell_6t
Xbit_r146_c26 bl[26] br[26] wl[146] vdd gnd cell_6t
Xbit_r147_c26 bl[26] br[26] wl[147] vdd gnd cell_6t
Xbit_r148_c26 bl[26] br[26] wl[148] vdd gnd cell_6t
Xbit_r149_c26 bl[26] br[26] wl[149] vdd gnd cell_6t
Xbit_r150_c26 bl[26] br[26] wl[150] vdd gnd cell_6t
Xbit_r151_c26 bl[26] br[26] wl[151] vdd gnd cell_6t
Xbit_r152_c26 bl[26] br[26] wl[152] vdd gnd cell_6t
Xbit_r153_c26 bl[26] br[26] wl[153] vdd gnd cell_6t
Xbit_r154_c26 bl[26] br[26] wl[154] vdd gnd cell_6t
Xbit_r155_c26 bl[26] br[26] wl[155] vdd gnd cell_6t
Xbit_r156_c26 bl[26] br[26] wl[156] vdd gnd cell_6t
Xbit_r157_c26 bl[26] br[26] wl[157] vdd gnd cell_6t
Xbit_r158_c26 bl[26] br[26] wl[158] vdd gnd cell_6t
Xbit_r159_c26 bl[26] br[26] wl[159] vdd gnd cell_6t
Xbit_r160_c26 bl[26] br[26] wl[160] vdd gnd cell_6t
Xbit_r161_c26 bl[26] br[26] wl[161] vdd gnd cell_6t
Xbit_r162_c26 bl[26] br[26] wl[162] vdd gnd cell_6t
Xbit_r163_c26 bl[26] br[26] wl[163] vdd gnd cell_6t
Xbit_r164_c26 bl[26] br[26] wl[164] vdd gnd cell_6t
Xbit_r165_c26 bl[26] br[26] wl[165] vdd gnd cell_6t
Xbit_r166_c26 bl[26] br[26] wl[166] vdd gnd cell_6t
Xbit_r167_c26 bl[26] br[26] wl[167] vdd gnd cell_6t
Xbit_r168_c26 bl[26] br[26] wl[168] vdd gnd cell_6t
Xbit_r169_c26 bl[26] br[26] wl[169] vdd gnd cell_6t
Xbit_r170_c26 bl[26] br[26] wl[170] vdd gnd cell_6t
Xbit_r171_c26 bl[26] br[26] wl[171] vdd gnd cell_6t
Xbit_r172_c26 bl[26] br[26] wl[172] vdd gnd cell_6t
Xbit_r173_c26 bl[26] br[26] wl[173] vdd gnd cell_6t
Xbit_r174_c26 bl[26] br[26] wl[174] vdd gnd cell_6t
Xbit_r175_c26 bl[26] br[26] wl[175] vdd gnd cell_6t
Xbit_r176_c26 bl[26] br[26] wl[176] vdd gnd cell_6t
Xbit_r177_c26 bl[26] br[26] wl[177] vdd gnd cell_6t
Xbit_r178_c26 bl[26] br[26] wl[178] vdd gnd cell_6t
Xbit_r179_c26 bl[26] br[26] wl[179] vdd gnd cell_6t
Xbit_r180_c26 bl[26] br[26] wl[180] vdd gnd cell_6t
Xbit_r181_c26 bl[26] br[26] wl[181] vdd gnd cell_6t
Xbit_r182_c26 bl[26] br[26] wl[182] vdd gnd cell_6t
Xbit_r183_c26 bl[26] br[26] wl[183] vdd gnd cell_6t
Xbit_r184_c26 bl[26] br[26] wl[184] vdd gnd cell_6t
Xbit_r185_c26 bl[26] br[26] wl[185] vdd gnd cell_6t
Xbit_r186_c26 bl[26] br[26] wl[186] vdd gnd cell_6t
Xbit_r187_c26 bl[26] br[26] wl[187] vdd gnd cell_6t
Xbit_r188_c26 bl[26] br[26] wl[188] vdd gnd cell_6t
Xbit_r189_c26 bl[26] br[26] wl[189] vdd gnd cell_6t
Xbit_r190_c26 bl[26] br[26] wl[190] vdd gnd cell_6t
Xbit_r191_c26 bl[26] br[26] wl[191] vdd gnd cell_6t
Xbit_r192_c26 bl[26] br[26] wl[192] vdd gnd cell_6t
Xbit_r193_c26 bl[26] br[26] wl[193] vdd gnd cell_6t
Xbit_r194_c26 bl[26] br[26] wl[194] vdd gnd cell_6t
Xbit_r195_c26 bl[26] br[26] wl[195] vdd gnd cell_6t
Xbit_r196_c26 bl[26] br[26] wl[196] vdd gnd cell_6t
Xbit_r197_c26 bl[26] br[26] wl[197] vdd gnd cell_6t
Xbit_r198_c26 bl[26] br[26] wl[198] vdd gnd cell_6t
Xbit_r199_c26 bl[26] br[26] wl[199] vdd gnd cell_6t
Xbit_r200_c26 bl[26] br[26] wl[200] vdd gnd cell_6t
Xbit_r201_c26 bl[26] br[26] wl[201] vdd gnd cell_6t
Xbit_r202_c26 bl[26] br[26] wl[202] vdd gnd cell_6t
Xbit_r203_c26 bl[26] br[26] wl[203] vdd gnd cell_6t
Xbit_r204_c26 bl[26] br[26] wl[204] vdd gnd cell_6t
Xbit_r205_c26 bl[26] br[26] wl[205] vdd gnd cell_6t
Xbit_r206_c26 bl[26] br[26] wl[206] vdd gnd cell_6t
Xbit_r207_c26 bl[26] br[26] wl[207] vdd gnd cell_6t
Xbit_r208_c26 bl[26] br[26] wl[208] vdd gnd cell_6t
Xbit_r209_c26 bl[26] br[26] wl[209] vdd gnd cell_6t
Xbit_r210_c26 bl[26] br[26] wl[210] vdd gnd cell_6t
Xbit_r211_c26 bl[26] br[26] wl[211] vdd gnd cell_6t
Xbit_r212_c26 bl[26] br[26] wl[212] vdd gnd cell_6t
Xbit_r213_c26 bl[26] br[26] wl[213] vdd gnd cell_6t
Xbit_r214_c26 bl[26] br[26] wl[214] vdd gnd cell_6t
Xbit_r215_c26 bl[26] br[26] wl[215] vdd gnd cell_6t
Xbit_r216_c26 bl[26] br[26] wl[216] vdd gnd cell_6t
Xbit_r217_c26 bl[26] br[26] wl[217] vdd gnd cell_6t
Xbit_r218_c26 bl[26] br[26] wl[218] vdd gnd cell_6t
Xbit_r219_c26 bl[26] br[26] wl[219] vdd gnd cell_6t
Xbit_r220_c26 bl[26] br[26] wl[220] vdd gnd cell_6t
Xbit_r221_c26 bl[26] br[26] wl[221] vdd gnd cell_6t
Xbit_r222_c26 bl[26] br[26] wl[222] vdd gnd cell_6t
Xbit_r223_c26 bl[26] br[26] wl[223] vdd gnd cell_6t
Xbit_r224_c26 bl[26] br[26] wl[224] vdd gnd cell_6t
Xbit_r225_c26 bl[26] br[26] wl[225] vdd gnd cell_6t
Xbit_r226_c26 bl[26] br[26] wl[226] vdd gnd cell_6t
Xbit_r227_c26 bl[26] br[26] wl[227] vdd gnd cell_6t
Xbit_r228_c26 bl[26] br[26] wl[228] vdd gnd cell_6t
Xbit_r229_c26 bl[26] br[26] wl[229] vdd gnd cell_6t
Xbit_r230_c26 bl[26] br[26] wl[230] vdd gnd cell_6t
Xbit_r231_c26 bl[26] br[26] wl[231] vdd gnd cell_6t
Xbit_r232_c26 bl[26] br[26] wl[232] vdd gnd cell_6t
Xbit_r233_c26 bl[26] br[26] wl[233] vdd gnd cell_6t
Xbit_r234_c26 bl[26] br[26] wl[234] vdd gnd cell_6t
Xbit_r235_c26 bl[26] br[26] wl[235] vdd gnd cell_6t
Xbit_r236_c26 bl[26] br[26] wl[236] vdd gnd cell_6t
Xbit_r237_c26 bl[26] br[26] wl[237] vdd gnd cell_6t
Xbit_r238_c26 bl[26] br[26] wl[238] vdd gnd cell_6t
Xbit_r239_c26 bl[26] br[26] wl[239] vdd gnd cell_6t
Xbit_r240_c26 bl[26] br[26] wl[240] vdd gnd cell_6t
Xbit_r241_c26 bl[26] br[26] wl[241] vdd gnd cell_6t
Xbit_r242_c26 bl[26] br[26] wl[242] vdd gnd cell_6t
Xbit_r243_c26 bl[26] br[26] wl[243] vdd gnd cell_6t
Xbit_r244_c26 bl[26] br[26] wl[244] vdd gnd cell_6t
Xbit_r245_c26 bl[26] br[26] wl[245] vdd gnd cell_6t
Xbit_r246_c26 bl[26] br[26] wl[246] vdd gnd cell_6t
Xbit_r247_c26 bl[26] br[26] wl[247] vdd gnd cell_6t
Xbit_r248_c26 bl[26] br[26] wl[248] vdd gnd cell_6t
Xbit_r249_c26 bl[26] br[26] wl[249] vdd gnd cell_6t
Xbit_r250_c26 bl[26] br[26] wl[250] vdd gnd cell_6t
Xbit_r251_c26 bl[26] br[26] wl[251] vdd gnd cell_6t
Xbit_r252_c26 bl[26] br[26] wl[252] vdd gnd cell_6t
Xbit_r253_c26 bl[26] br[26] wl[253] vdd gnd cell_6t
Xbit_r254_c26 bl[26] br[26] wl[254] vdd gnd cell_6t
Xbit_r255_c26 bl[26] br[26] wl[255] vdd gnd cell_6t
Xbit_r256_c26 bl[26] br[26] wl[256] vdd gnd cell_6t
Xbit_r257_c26 bl[26] br[26] wl[257] vdd gnd cell_6t
Xbit_r258_c26 bl[26] br[26] wl[258] vdd gnd cell_6t
Xbit_r259_c26 bl[26] br[26] wl[259] vdd gnd cell_6t
Xbit_r260_c26 bl[26] br[26] wl[260] vdd gnd cell_6t
Xbit_r261_c26 bl[26] br[26] wl[261] vdd gnd cell_6t
Xbit_r262_c26 bl[26] br[26] wl[262] vdd gnd cell_6t
Xbit_r263_c26 bl[26] br[26] wl[263] vdd gnd cell_6t
Xbit_r264_c26 bl[26] br[26] wl[264] vdd gnd cell_6t
Xbit_r265_c26 bl[26] br[26] wl[265] vdd gnd cell_6t
Xbit_r266_c26 bl[26] br[26] wl[266] vdd gnd cell_6t
Xbit_r267_c26 bl[26] br[26] wl[267] vdd gnd cell_6t
Xbit_r268_c26 bl[26] br[26] wl[268] vdd gnd cell_6t
Xbit_r269_c26 bl[26] br[26] wl[269] vdd gnd cell_6t
Xbit_r270_c26 bl[26] br[26] wl[270] vdd gnd cell_6t
Xbit_r271_c26 bl[26] br[26] wl[271] vdd gnd cell_6t
Xbit_r272_c26 bl[26] br[26] wl[272] vdd gnd cell_6t
Xbit_r273_c26 bl[26] br[26] wl[273] vdd gnd cell_6t
Xbit_r274_c26 bl[26] br[26] wl[274] vdd gnd cell_6t
Xbit_r275_c26 bl[26] br[26] wl[275] vdd gnd cell_6t
Xbit_r276_c26 bl[26] br[26] wl[276] vdd gnd cell_6t
Xbit_r277_c26 bl[26] br[26] wl[277] vdd gnd cell_6t
Xbit_r278_c26 bl[26] br[26] wl[278] vdd gnd cell_6t
Xbit_r279_c26 bl[26] br[26] wl[279] vdd gnd cell_6t
Xbit_r280_c26 bl[26] br[26] wl[280] vdd gnd cell_6t
Xbit_r281_c26 bl[26] br[26] wl[281] vdd gnd cell_6t
Xbit_r282_c26 bl[26] br[26] wl[282] vdd gnd cell_6t
Xbit_r283_c26 bl[26] br[26] wl[283] vdd gnd cell_6t
Xbit_r284_c26 bl[26] br[26] wl[284] vdd gnd cell_6t
Xbit_r285_c26 bl[26] br[26] wl[285] vdd gnd cell_6t
Xbit_r286_c26 bl[26] br[26] wl[286] vdd gnd cell_6t
Xbit_r287_c26 bl[26] br[26] wl[287] vdd gnd cell_6t
Xbit_r288_c26 bl[26] br[26] wl[288] vdd gnd cell_6t
Xbit_r289_c26 bl[26] br[26] wl[289] vdd gnd cell_6t
Xbit_r290_c26 bl[26] br[26] wl[290] vdd gnd cell_6t
Xbit_r291_c26 bl[26] br[26] wl[291] vdd gnd cell_6t
Xbit_r292_c26 bl[26] br[26] wl[292] vdd gnd cell_6t
Xbit_r293_c26 bl[26] br[26] wl[293] vdd gnd cell_6t
Xbit_r294_c26 bl[26] br[26] wl[294] vdd gnd cell_6t
Xbit_r295_c26 bl[26] br[26] wl[295] vdd gnd cell_6t
Xbit_r296_c26 bl[26] br[26] wl[296] vdd gnd cell_6t
Xbit_r297_c26 bl[26] br[26] wl[297] vdd gnd cell_6t
Xbit_r298_c26 bl[26] br[26] wl[298] vdd gnd cell_6t
Xbit_r299_c26 bl[26] br[26] wl[299] vdd gnd cell_6t
Xbit_r300_c26 bl[26] br[26] wl[300] vdd gnd cell_6t
Xbit_r301_c26 bl[26] br[26] wl[301] vdd gnd cell_6t
Xbit_r302_c26 bl[26] br[26] wl[302] vdd gnd cell_6t
Xbit_r303_c26 bl[26] br[26] wl[303] vdd gnd cell_6t
Xbit_r304_c26 bl[26] br[26] wl[304] vdd gnd cell_6t
Xbit_r305_c26 bl[26] br[26] wl[305] vdd gnd cell_6t
Xbit_r306_c26 bl[26] br[26] wl[306] vdd gnd cell_6t
Xbit_r307_c26 bl[26] br[26] wl[307] vdd gnd cell_6t
Xbit_r308_c26 bl[26] br[26] wl[308] vdd gnd cell_6t
Xbit_r309_c26 bl[26] br[26] wl[309] vdd gnd cell_6t
Xbit_r310_c26 bl[26] br[26] wl[310] vdd gnd cell_6t
Xbit_r311_c26 bl[26] br[26] wl[311] vdd gnd cell_6t
Xbit_r312_c26 bl[26] br[26] wl[312] vdd gnd cell_6t
Xbit_r313_c26 bl[26] br[26] wl[313] vdd gnd cell_6t
Xbit_r314_c26 bl[26] br[26] wl[314] vdd gnd cell_6t
Xbit_r315_c26 bl[26] br[26] wl[315] vdd gnd cell_6t
Xbit_r316_c26 bl[26] br[26] wl[316] vdd gnd cell_6t
Xbit_r317_c26 bl[26] br[26] wl[317] vdd gnd cell_6t
Xbit_r318_c26 bl[26] br[26] wl[318] vdd gnd cell_6t
Xbit_r319_c26 bl[26] br[26] wl[319] vdd gnd cell_6t
Xbit_r320_c26 bl[26] br[26] wl[320] vdd gnd cell_6t
Xbit_r321_c26 bl[26] br[26] wl[321] vdd gnd cell_6t
Xbit_r322_c26 bl[26] br[26] wl[322] vdd gnd cell_6t
Xbit_r323_c26 bl[26] br[26] wl[323] vdd gnd cell_6t
Xbit_r324_c26 bl[26] br[26] wl[324] vdd gnd cell_6t
Xbit_r325_c26 bl[26] br[26] wl[325] vdd gnd cell_6t
Xbit_r326_c26 bl[26] br[26] wl[326] vdd gnd cell_6t
Xbit_r327_c26 bl[26] br[26] wl[327] vdd gnd cell_6t
Xbit_r328_c26 bl[26] br[26] wl[328] vdd gnd cell_6t
Xbit_r329_c26 bl[26] br[26] wl[329] vdd gnd cell_6t
Xbit_r330_c26 bl[26] br[26] wl[330] vdd gnd cell_6t
Xbit_r331_c26 bl[26] br[26] wl[331] vdd gnd cell_6t
Xbit_r332_c26 bl[26] br[26] wl[332] vdd gnd cell_6t
Xbit_r333_c26 bl[26] br[26] wl[333] vdd gnd cell_6t
Xbit_r334_c26 bl[26] br[26] wl[334] vdd gnd cell_6t
Xbit_r335_c26 bl[26] br[26] wl[335] vdd gnd cell_6t
Xbit_r336_c26 bl[26] br[26] wl[336] vdd gnd cell_6t
Xbit_r337_c26 bl[26] br[26] wl[337] vdd gnd cell_6t
Xbit_r338_c26 bl[26] br[26] wl[338] vdd gnd cell_6t
Xbit_r339_c26 bl[26] br[26] wl[339] vdd gnd cell_6t
Xbit_r340_c26 bl[26] br[26] wl[340] vdd gnd cell_6t
Xbit_r341_c26 bl[26] br[26] wl[341] vdd gnd cell_6t
Xbit_r342_c26 bl[26] br[26] wl[342] vdd gnd cell_6t
Xbit_r343_c26 bl[26] br[26] wl[343] vdd gnd cell_6t
Xbit_r344_c26 bl[26] br[26] wl[344] vdd gnd cell_6t
Xbit_r345_c26 bl[26] br[26] wl[345] vdd gnd cell_6t
Xbit_r346_c26 bl[26] br[26] wl[346] vdd gnd cell_6t
Xbit_r347_c26 bl[26] br[26] wl[347] vdd gnd cell_6t
Xbit_r348_c26 bl[26] br[26] wl[348] vdd gnd cell_6t
Xbit_r349_c26 bl[26] br[26] wl[349] vdd gnd cell_6t
Xbit_r350_c26 bl[26] br[26] wl[350] vdd gnd cell_6t
Xbit_r351_c26 bl[26] br[26] wl[351] vdd gnd cell_6t
Xbit_r352_c26 bl[26] br[26] wl[352] vdd gnd cell_6t
Xbit_r353_c26 bl[26] br[26] wl[353] vdd gnd cell_6t
Xbit_r354_c26 bl[26] br[26] wl[354] vdd gnd cell_6t
Xbit_r355_c26 bl[26] br[26] wl[355] vdd gnd cell_6t
Xbit_r356_c26 bl[26] br[26] wl[356] vdd gnd cell_6t
Xbit_r357_c26 bl[26] br[26] wl[357] vdd gnd cell_6t
Xbit_r358_c26 bl[26] br[26] wl[358] vdd gnd cell_6t
Xbit_r359_c26 bl[26] br[26] wl[359] vdd gnd cell_6t
Xbit_r360_c26 bl[26] br[26] wl[360] vdd gnd cell_6t
Xbit_r361_c26 bl[26] br[26] wl[361] vdd gnd cell_6t
Xbit_r362_c26 bl[26] br[26] wl[362] vdd gnd cell_6t
Xbit_r363_c26 bl[26] br[26] wl[363] vdd gnd cell_6t
Xbit_r364_c26 bl[26] br[26] wl[364] vdd gnd cell_6t
Xbit_r365_c26 bl[26] br[26] wl[365] vdd gnd cell_6t
Xbit_r366_c26 bl[26] br[26] wl[366] vdd gnd cell_6t
Xbit_r367_c26 bl[26] br[26] wl[367] vdd gnd cell_6t
Xbit_r368_c26 bl[26] br[26] wl[368] vdd gnd cell_6t
Xbit_r369_c26 bl[26] br[26] wl[369] vdd gnd cell_6t
Xbit_r370_c26 bl[26] br[26] wl[370] vdd gnd cell_6t
Xbit_r371_c26 bl[26] br[26] wl[371] vdd gnd cell_6t
Xbit_r372_c26 bl[26] br[26] wl[372] vdd gnd cell_6t
Xbit_r373_c26 bl[26] br[26] wl[373] vdd gnd cell_6t
Xbit_r374_c26 bl[26] br[26] wl[374] vdd gnd cell_6t
Xbit_r375_c26 bl[26] br[26] wl[375] vdd gnd cell_6t
Xbit_r376_c26 bl[26] br[26] wl[376] vdd gnd cell_6t
Xbit_r377_c26 bl[26] br[26] wl[377] vdd gnd cell_6t
Xbit_r378_c26 bl[26] br[26] wl[378] vdd gnd cell_6t
Xbit_r379_c26 bl[26] br[26] wl[379] vdd gnd cell_6t
Xbit_r380_c26 bl[26] br[26] wl[380] vdd gnd cell_6t
Xbit_r381_c26 bl[26] br[26] wl[381] vdd gnd cell_6t
Xbit_r382_c26 bl[26] br[26] wl[382] vdd gnd cell_6t
Xbit_r383_c26 bl[26] br[26] wl[383] vdd gnd cell_6t
Xbit_r384_c26 bl[26] br[26] wl[384] vdd gnd cell_6t
Xbit_r385_c26 bl[26] br[26] wl[385] vdd gnd cell_6t
Xbit_r386_c26 bl[26] br[26] wl[386] vdd gnd cell_6t
Xbit_r387_c26 bl[26] br[26] wl[387] vdd gnd cell_6t
Xbit_r388_c26 bl[26] br[26] wl[388] vdd gnd cell_6t
Xbit_r389_c26 bl[26] br[26] wl[389] vdd gnd cell_6t
Xbit_r390_c26 bl[26] br[26] wl[390] vdd gnd cell_6t
Xbit_r391_c26 bl[26] br[26] wl[391] vdd gnd cell_6t
Xbit_r392_c26 bl[26] br[26] wl[392] vdd gnd cell_6t
Xbit_r393_c26 bl[26] br[26] wl[393] vdd gnd cell_6t
Xbit_r394_c26 bl[26] br[26] wl[394] vdd gnd cell_6t
Xbit_r395_c26 bl[26] br[26] wl[395] vdd gnd cell_6t
Xbit_r396_c26 bl[26] br[26] wl[396] vdd gnd cell_6t
Xbit_r397_c26 bl[26] br[26] wl[397] vdd gnd cell_6t
Xbit_r398_c26 bl[26] br[26] wl[398] vdd gnd cell_6t
Xbit_r399_c26 bl[26] br[26] wl[399] vdd gnd cell_6t
Xbit_r400_c26 bl[26] br[26] wl[400] vdd gnd cell_6t
Xbit_r401_c26 bl[26] br[26] wl[401] vdd gnd cell_6t
Xbit_r402_c26 bl[26] br[26] wl[402] vdd gnd cell_6t
Xbit_r403_c26 bl[26] br[26] wl[403] vdd gnd cell_6t
Xbit_r404_c26 bl[26] br[26] wl[404] vdd gnd cell_6t
Xbit_r405_c26 bl[26] br[26] wl[405] vdd gnd cell_6t
Xbit_r406_c26 bl[26] br[26] wl[406] vdd gnd cell_6t
Xbit_r407_c26 bl[26] br[26] wl[407] vdd gnd cell_6t
Xbit_r408_c26 bl[26] br[26] wl[408] vdd gnd cell_6t
Xbit_r409_c26 bl[26] br[26] wl[409] vdd gnd cell_6t
Xbit_r410_c26 bl[26] br[26] wl[410] vdd gnd cell_6t
Xbit_r411_c26 bl[26] br[26] wl[411] vdd gnd cell_6t
Xbit_r412_c26 bl[26] br[26] wl[412] vdd gnd cell_6t
Xbit_r413_c26 bl[26] br[26] wl[413] vdd gnd cell_6t
Xbit_r414_c26 bl[26] br[26] wl[414] vdd gnd cell_6t
Xbit_r415_c26 bl[26] br[26] wl[415] vdd gnd cell_6t
Xbit_r416_c26 bl[26] br[26] wl[416] vdd gnd cell_6t
Xbit_r417_c26 bl[26] br[26] wl[417] vdd gnd cell_6t
Xbit_r418_c26 bl[26] br[26] wl[418] vdd gnd cell_6t
Xbit_r419_c26 bl[26] br[26] wl[419] vdd gnd cell_6t
Xbit_r420_c26 bl[26] br[26] wl[420] vdd gnd cell_6t
Xbit_r421_c26 bl[26] br[26] wl[421] vdd gnd cell_6t
Xbit_r422_c26 bl[26] br[26] wl[422] vdd gnd cell_6t
Xbit_r423_c26 bl[26] br[26] wl[423] vdd gnd cell_6t
Xbit_r424_c26 bl[26] br[26] wl[424] vdd gnd cell_6t
Xbit_r425_c26 bl[26] br[26] wl[425] vdd gnd cell_6t
Xbit_r426_c26 bl[26] br[26] wl[426] vdd gnd cell_6t
Xbit_r427_c26 bl[26] br[26] wl[427] vdd gnd cell_6t
Xbit_r428_c26 bl[26] br[26] wl[428] vdd gnd cell_6t
Xbit_r429_c26 bl[26] br[26] wl[429] vdd gnd cell_6t
Xbit_r430_c26 bl[26] br[26] wl[430] vdd gnd cell_6t
Xbit_r431_c26 bl[26] br[26] wl[431] vdd gnd cell_6t
Xbit_r432_c26 bl[26] br[26] wl[432] vdd gnd cell_6t
Xbit_r433_c26 bl[26] br[26] wl[433] vdd gnd cell_6t
Xbit_r434_c26 bl[26] br[26] wl[434] vdd gnd cell_6t
Xbit_r435_c26 bl[26] br[26] wl[435] vdd gnd cell_6t
Xbit_r436_c26 bl[26] br[26] wl[436] vdd gnd cell_6t
Xbit_r437_c26 bl[26] br[26] wl[437] vdd gnd cell_6t
Xbit_r438_c26 bl[26] br[26] wl[438] vdd gnd cell_6t
Xbit_r439_c26 bl[26] br[26] wl[439] vdd gnd cell_6t
Xbit_r440_c26 bl[26] br[26] wl[440] vdd gnd cell_6t
Xbit_r441_c26 bl[26] br[26] wl[441] vdd gnd cell_6t
Xbit_r442_c26 bl[26] br[26] wl[442] vdd gnd cell_6t
Xbit_r443_c26 bl[26] br[26] wl[443] vdd gnd cell_6t
Xbit_r444_c26 bl[26] br[26] wl[444] vdd gnd cell_6t
Xbit_r445_c26 bl[26] br[26] wl[445] vdd gnd cell_6t
Xbit_r446_c26 bl[26] br[26] wl[446] vdd gnd cell_6t
Xbit_r447_c26 bl[26] br[26] wl[447] vdd gnd cell_6t
Xbit_r448_c26 bl[26] br[26] wl[448] vdd gnd cell_6t
Xbit_r449_c26 bl[26] br[26] wl[449] vdd gnd cell_6t
Xbit_r450_c26 bl[26] br[26] wl[450] vdd gnd cell_6t
Xbit_r451_c26 bl[26] br[26] wl[451] vdd gnd cell_6t
Xbit_r452_c26 bl[26] br[26] wl[452] vdd gnd cell_6t
Xbit_r453_c26 bl[26] br[26] wl[453] vdd gnd cell_6t
Xbit_r454_c26 bl[26] br[26] wl[454] vdd gnd cell_6t
Xbit_r455_c26 bl[26] br[26] wl[455] vdd gnd cell_6t
Xbit_r456_c26 bl[26] br[26] wl[456] vdd gnd cell_6t
Xbit_r457_c26 bl[26] br[26] wl[457] vdd gnd cell_6t
Xbit_r458_c26 bl[26] br[26] wl[458] vdd gnd cell_6t
Xbit_r459_c26 bl[26] br[26] wl[459] vdd gnd cell_6t
Xbit_r460_c26 bl[26] br[26] wl[460] vdd gnd cell_6t
Xbit_r461_c26 bl[26] br[26] wl[461] vdd gnd cell_6t
Xbit_r462_c26 bl[26] br[26] wl[462] vdd gnd cell_6t
Xbit_r463_c26 bl[26] br[26] wl[463] vdd gnd cell_6t
Xbit_r464_c26 bl[26] br[26] wl[464] vdd gnd cell_6t
Xbit_r465_c26 bl[26] br[26] wl[465] vdd gnd cell_6t
Xbit_r466_c26 bl[26] br[26] wl[466] vdd gnd cell_6t
Xbit_r467_c26 bl[26] br[26] wl[467] vdd gnd cell_6t
Xbit_r468_c26 bl[26] br[26] wl[468] vdd gnd cell_6t
Xbit_r469_c26 bl[26] br[26] wl[469] vdd gnd cell_6t
Xbit_r470_c26 bl[26] br[26] wl[470] vdd gnd cell_6t
Xbit_r471_c26 bl[26] br[26] wl[471] vdd gnd cell_6t
Xbit_r472_c26 bl[26] br[26] wl[472] vdd gnd cell_6t
Xbit_r473_c26 bl[26] br[26] wl[473] vdd gnd cell_6t
Xbit_r474_c26 bl[26] br[26] wl[474] vdd gnd cell_6t
Xbit_r475_c26 bl[26] br[26] wl[475] vdd gnd cell_6t
Xbit_r476_c26 bl[26] br[26] wl[476] vdd gnd cell_6t
Xbit_r477_c26 bl[26] br[26] wl[477] vdd gnd cell_6t
Xbit_r478_c26 bl[26] br[26] wl[478] vdd gnd cell_6t
Xbit_r479_c26 bl[26] br[26] wl[479] vdd gnd cell_6t
Xbit_r480_c26 bl[26] br[26] wl[480] vdd gnd cell_6t
Xbit_r481_c26 bl[26] br[26] wl[481] vdd gnd cell_6t
Xbit_r482_c26 bl[26] br[26] wl[482] vdd gnd cell_6t
Xbit_r483_c26 bl[26] br[26] wl[483] vdd gnd cell_6t
Xbit_r484_c26 bl[26] br[26] wl[484] vdd gnd cell_6t
Xbit_r485_c26 bl[26] br[26] wl[485] vdd gnd cell_6t
Xbit_r486_c26 bl[26] br[26] wl[486] vdd gnd cell_6t
Xbit_r487_c26 bl[26] br[26] wl[487] vdd gnd cell_6t
Xbit_r488_c26 bl[26] br[26] wl[488] vdd gnd cell_6t
Xbit_r489_c26 bl[26] br[26] wl[489] vdd gnd cell_6t
Xbit_r490_c26 bl[26] br[26] wl[490] vdd gnd cell_6t
Xbit_r491_c26 bl[26] br[26] wl[491] vdd gnd cell_6t
Xbit_r492_c26 bl[26] br[26] wl[492] vdd gnd cell_6t
Xbit_r493_c26 bl[26] br[26] wl[493] vdd gnd cell_6t
Xbit_r494_c26 bl[26] br[26] wl[494] vdd gnd cell_6t
Xbit_r495_c26 bl[26] br[26] wl[495] vdd gnd cell_6t
Xbit_r496_c26 bl[26] br[26] wl[496] vdd gnd cell_6t
Xbit_r497_c26 bl[26] br[26] wl[497] vdd gnd cell_6t
Xbit_r498_c26 bl[26] br[26] wl[498] vdd gnd cell_6t
Xbit_r499_c26 bl[26] br[26] wl[499] vdd gnd cell_6t
Xbit_r500_c26 bl[26] br[26] wl[500] vdd gnd cell_6t
Xbit_r501_c26 bl[26] br[26] wl[501] vdd gnd cell_6t
Xbit_r502_c26 bl[26] br[26] wl[502] vdd gnd cell_6t
Xbit_r503_c26 bl[26] br[26] wl[503] vdd gnd cell_6t
Xbit_r504_c26 bl[26] br[26] wl[504] vdd gnd cell_6t
Xbit_r505_c26 bl[26] br[26] wl[505] vdd gnd cell_6t
Xbit_r506_c26 bl[26] br[26] wl[506] vdd gnd cell_6t
Xbit_r507_c26 bl[26] br[26] wl[507] vdd gnd cell_6t
Xbit_r508_c26 bl[26] br[26] wl[508] vdd gnd cell_6t
Xbit_r509_c26 bl[26] br[26] wl[509] vdd gnd cell_6t
Xbit_r510_c26 bl[26] br[26] wl[510] vdd gnd cell_6t
Xbit_r511_c26 bl[26] br[26] wl[511] vdd gnd cell_6t
Xbit_r0_c27 bl[27] br[27] wl[0] vdd gnd cell_6t
Xbit_r1_c27 bl[27] br[27] wl[1] vdd gnd cell_6t
Xbit_r2_c27 bl[27] br[27] wl[2] vdd gnd cell_6t
Xbit_r3_c27 bl[27] br[27] wl[3] vdd gnd cell_6t
Xbit_r4_c27 bl[27] br[27] wl[4] vdd gnd cell_6t
Xbit_r5_c27 bl[27] br[27] wl[5] vdd gnd cell_6t
Xbit_r6_c27 bl[27] br[27] wl[6] vdd gnd cell_6t
Xbit_r7_c27 bl[27] br[27] wl[7] vdd gnd cell_6t
Xbit_r8_c27 bl[27] br[27] wl[8] vdd gnd cell_6t
Xbit_r9_c27 bl[27] br[27] wl[9] vdd gnd cell_6t
Xbit_r10_c27 bl[27] br[27] wl[10] vdd gnd cell_6t
Xbit_r11_c27 bl[27] br[27] wl[11] vdd gnd cell_6t
Xbit_r12_c27 bl[27] br[27] wl[12] vdd gnd cell_6t
Xbit_r13_c27 bl[27] br[27] wl[13] vdd gnd cell_6t
Xbit_r14_c27 bl[27] br[27] wl[14] vdd gnd cell_6t
Xbit_r15_c27 bl[27] br[27] wl[15] vdd gnd cell_6t
Xbit_r16_c27 bl[27] br[27] wl[16] vdd gnd cell_6t
Xbit_r17_c27 bl[27] br[27] wl[17] vdd gnd cell_6t
Xbit_r18_c27 bl[27] br[27] wl[18] vdd gnd cell_6t
Xbit_r19_c27 bl[27] br[27] wl[19] vdd gnd cell_6t
Xbit_r20_c27 bl[27] br[27] wl[20] vdd gnd cell_6t
Xbit_r21_c27 bl[27] br[27] wl[21] vdd gnd cell_6t
Xbit_r22_c27 bl[27] br[27] wl[22] vdd gnd cell_6t
Xbit_r23_c27 bl[27] br[27] wl[23] vdd gnd cell_6t
Xbit_r24_c27 bl[27] br[27] wl[24] vdd gnd cell_6t
Xbit_r25_c27 bl[27] br[27] wl[25] vdd gnd cell_6t
Xbit_r26_c27 bl[27] br[27] wl[26] vdd gnd cell_6t
Xbit_r27_c27 bl[27] br[27] wl[27] vdd gnd cell_6t
Xbit_r28_c27 bl[27] br[27] wl[28] vdd gnd cell_6t
Xbit_r29_c27 bl[27] br[27] wl[29] vdd gnd cell_6t
Xbit_r30_c27 bl[27] br[27] wl[30] vdd gnd cell_6t
Xbit_r31_c27 bl[27] br[27] wl[31] vdd gnd cell_6t
Xbit_r32_c27 bl[27] br[27] wl[32] vdd gnd cell_6t
Xbit_r33_c27 bl[27] br[27] wl[33] vdd gnd cell_6t
Xbit_r34_c27 bl[27] br[27] wl[34] vdd gnd cell_6t
Xbit_r35_c27 bl[27] br[27] wl[35] vdd gnd cell_6t
Xbit_r36_c27 bl[27] br[27] wl[36] vdd gnd cell_6t
Xbit_r37_c27 bl[27] br[27] wl[37] vdd gnd cell_6t
Xbit_r38_c27 bl[27] br[27] wl[38] vdd gnd cell_6t
Xbit_r39_c27 bl[27] br[27] wl[39] vdd gnd cell_6t
Xbit_r40_c27 bl[27] br[27] wl[40] vdd gnd cell_6t
Xbit_r41_c27 bl[27] br[27] wl[41] vdd gnd cell_6t
Xbit_r42_c27 bl[27] br[27] wl[42] vdd gnd cell_6t
Xbit_r43_c27 bl[27] br[27] wl[43] vdd gnd cell_6t
Xbit_r44_c27 bl[27] br[27] wl[44] vdd gnd cell_6t
Xbit_r45_c27 bl[27] br[27] wl[45] vdd gnd cell_6t
Xbit_r46_c27 bl[27] br[27] wl[46] vdd gnd cell_6t
Xbit_r47_c27 bl[27] br[27] wl[47] vdd gnd cell_6t
Xbit_r48_c27 bl[27] br[27] wl[48] vdd gnd cell_6t
Xbit_r49_c27 bl[27] br[27] wl[49] vdd gnd cell_6t
Xbit_r50_c27 bl[27] br[27] wl[50] vdd gnd cell_6t
Xbit_r51_c27 bl[27] br[27] wl[51] vdd gnd cell_6t
Xbit_r52_c27 bl[27] br[27] wl[52] vdd gnd cell_6t
Xbit_r53_c27 bl[27] br[27] wl[53] vdd gnd cell_6t
Xbit_r54_c27 bl[27] br[27] wl[54] vdd gnd cell_6t
Xbit_r55_c27 bl[27] br[27] wl[55] vdd gnd cell_6t
Xbit_r56_c27 bl[27] br[27] wl[56] vdd gnd cell_6t
Xbit_r57_c27 bl[27] br[27] wl[57] vdd gnd cell_6t
Xbit_r58_c27 bl[27] br[27] wl[58] vdd gnd cell_6t
Xbit_r59_c27 bl[27] br[27] wl[59] vdd gnd cell_6t
Xbit_r60_c27 bl[27] br[27] wl[60] vdd gnd cell_6t
Xbit_r61_c27 bl[27] br[27] wl[61] vdd gnd cell_6t
Xbit_r62_c27 bl[27] br[27] wl[62] vdd gnd cell_6t
Xbit_r63_c27 bl[27] br[27] wl[63] vdd gnd cell_6t
Xbit_r64_c27 bl[27] br[27] wl[64] vdd gnd cell_6t
Xbit_r65_c27 bl[27] br[27] wl[65] vdd gnd cell_6t
Xbit_r66_c27 bl[27] br[27] wl[66] vdd gnd cell_6t
Xbit_r67_c27 bl[27] br[27] wl[67] vdd gnd cell_6t
Xbit_r68_c27 bl[27] br[27] wl[68] vdd gnd cell_6t
Xbit_r69_c27 bl[27] br[27] wl[69] vdd gnd cell_6t
Xbit_r70_c27 bl[27] br[27] wl[70] vdd gnd cell_6t
Xbit_r71_c27 bl[27] br[27] wl[71] vdd gnd cell_6t
Xbit_r72_c27 bl[27] br[27] wl[72] vdd gnd cell_6t
Xbit_r73_c27 bl[27] br[27] wl[73] vdd gnd cell_6t
Xbit_r74_c27 bl[27] br[27] wl[74] vdd gnd cell_6t
Xbit_r75_c27 bl[27] br[27] wl[75] vdd gnd cell_6t
Xbit_r76_c27 bl[27] br[27] wl[76] vdd gnd cell_6t
Xbit_r77_c27 bl[27] br[27] wl[77] vdd gnd cell_6t
Xbit_r78_c27 bl[27] br[27] wl[78] vdd gnd cell_6t
Xbit_r79_c27 bl[27] br[27] wl[79] vdd gnd cell_6t
Xbit_r80_c27 bl[27] br[27] wl[80] vdd gnd cell_6t
Xbit_r81_c27 bl[27] br[27] wl[81] vdd gnd cell_6t
Xbit_r82_c27 bl[27] br[27] wl[82] vdd gnd cell_6t
Xbit_r83_c27 bl[27] br[27] wl[83] vdd gnd cell_6t
Xbit_r84_c27 bl[27] br[27] wl[84] vdd gnd cell_6t
Xbit_r85_c27 bl[27] br[27] wl[85] vdd gnd cell_6t
Xbit_r86_c27 bl[27] br[27] wl[86] vdd gnd cell_6t
Xbit_r87_c27 bl[27] br[27] wl[87] vdd gnd cell_6t
Xbit_r88_c27 bl[27] br[27] wl[88] vdd gnd cell_6t
Xbit_r89_c27 bl[27] br[27] wl[89] vdd gnd cell_6t
Xbit_r90_c27 bl[27] br[27] wl[90] vdd gnd cell_6t
Xbit_r91_c27 bl[27] br[27] wl[91] vdd gnd cell_6t
Xbit_r92_c27 bl[27] br[27] wl[92] vdd gnd cell_6t
Xbit_r93_c27 bl[27] br[27] wl[93] vdd gnd cell_6t
Xbit_r94_c27 bl[27] br[27] wl[94] vdd gnd cell_6t
Xbit_r95_c27 bl[27] br[27] wl[95] vdd gnd cell_6t
Xbit_r96_c27 bl[27] br[27] wl[96] vdd gnd cell_6t
Xbit_r97_c27 bl[27] br[27] wl[97] vdd gnd cell_6t
Xbit_r98_c27 bl[27] br[27] wl[98] vdd gnd cell_6t
Xbit_r99_c27 bl[27] br[27] wl[99] vdd gnd cell_6t
Xbit_r100_c27 bl[27] br[27] wl[100] vdd gnd cell_6t
Xbit_r101_c27 bl[27] br[27] wl[101] vdd gnd cell_6t
Xbit_r102_c27 bl[27] br[27] wl[102] vdd gnd cell_6t
Xbit_r103_c27 bl[27] br[27] wl[103] vdd gnd cell_6t
Xbit_r104_c27 bl[27] br[27] wl[104] vdd gnd cell_6t
Xbit_r105_c27 bl[27] br[27] wl[105] vdd gnd cell_6t
Xbit_r106_c27 bl[27] br[27] wl[106] vdd gnd cell_6t
Xbit_r107_c27 bl[27] br[27] wl[107] vdd gnd cell_6t
Xbit_r108_c27 bl[27] br[27] wl[108] vdd gnd cell_6t
Xbit_r109_c27 bl[27] br[27] wl[109] vdd gnd cell_6t
Xbit_r110_c27 bl[27] br[27] wl[110] vdd gnd cell_6t
Xbit_r111_c27 bl[27] br[27] wl[111] vdd gnd cell_6t
Xbit_r112_c27 bl[27] br[27] wl[112] vdd gnd cell_6t
Xbit_r113_c27 bl[27] br[27] wl[113] vdd gnd cell_6t
Xbit_r114_c27 bl[27] br[27] wl[114] vdd gnd cell_6t
Xbit_r115_c27 bl[27] br[27] wl[115] vdd gnd cell_6t
Xbit_r116_c27 bl[27] br[27] wl[116] vdd gnd cell_6t
Xbit_r117_c27 bl[27] br[27] wl[117] vdd gnd cell_6t
Xbit_r118_c27 bl[27] br[27] wl[118] vdd gnd cell_6t
Xbit_r119_c27 bl[27] br[27] wl[119] vdd gnd cell_6t
Xbit_r120_c27 bl[27] br[27] wl[120] vdd gnd cell_6t
Xbit_r121_c27 bl[27] br[27] wl[121] vdd gnd cell_6t
Xbit_r122_c27 bl[27] br[27] wl[122] vdd gnd cell_6t
Xbit_r123_c27 bl[27] br[27] wl[123] vdd gnd cell_6t
Xbit_r124_c27 bl[27] br[27] wl[124] vdd gnd cell_6t
Xbit_r125_c27 bl[27] br[27] wl[125] vdd gnd cell_6t
Xbit_r126_c27 bl[27] br[27] wl[126] vdd gnd cell_6t
Xbit_r127_c27 bl[27] br[27] wl[127] vdd gnd cell_6t
Xbit_r128_c27 bl[27] br[27] wl[128] vdd gnd cell_6t
Xbit_r129_c27 bl[27] br[27] wl[129] vdd gnd cell_6t
Xbit_r130_c27 bl[27] br[27] wl[130] vdd gnd cell_6t
Xbit_r131_c27 bl[27] br[27] wl[131] vdd gnd cell_6t
Xbit_r132_c27 bl[27] br[27] wl[132] vdd gnd cell_6t
Xbit_r133_c27 bl[27] br[27] wl[133] vdd gnd cell_6t
Xbit_r134_c27 bl[27] br[27] wl[134] vdd gnd cell_6t
Xbit_r135_c27 bl[27] br[27] wl[135] vdd gnd cell_6t
Xbit_r136_c27 bl[27] br[27] wl[136] vdd gnd cell_6t
Xbit_r137_c27 bl[27] br[27] wl[137] vdd gnd cell_6t
Xbit_r138_c27 bl[27] br[27] wl[138] vdd gnd cell_6t
Xbit_r139_c27 bl[27] br[27] wl[139] vdd gnd cell_6t
Xbit_r140_c27 bl[27] br[27] wl[140] vdd gnd cell_6t
Xbit_r141_c27 bl[27] br[27] wl[141] vdd gnd cell_6t
Xbit_r142_c27 bl[27] br[27] wl[142] vdd gnd cell_6t
Xbit_r143_c27 bl[27] br[27] wl[143] vdd gnd cell_6t
Xbit_r144_c27 bl[27] br[27] wl[144] vdd gnd cell_6t
Xbit_r145_c27 bl[27] br[27] wl[145] vdd gnd cell_6t
Xbit_r146_c27 bl[27] br[27] wl[146] vdd gnd cell_6t
Xbit_r147_c27 bl[27] br[27] wl[147] vdd gnd cell_6t
Xbit_r148_c27 bl[27] br[27] wl[148] vdd gnd cell_6t
Xbit_r149_c27 bl[27] br[27] wl[149] vdd gnd cell_6t
Xbit_r150_c27 bl[27] br[27] wl[150] vdd gnd cell_6t
Xbit_r151_c27 bl[27] br[27] wl[151] vdd gnd cell_6t
Xbit_r152_c27 bl[27] br[27] wl[152] vdd gnd cell_6t
Xbit_r153_c27 bl[27] br[27] wl[153] vdd gnd cell_6t
Xbit_r154_c27 bl[27] br[27] wl[154] vdd gnd cell_6t
Xbit_r155_c27 bl[27] br[27] wl[155] vdd gnd cell_6t
Xbit_r156_c27 bl[27] br[27] wl[156] vdd gnd cell_6t
Xbit_r157_c27 bl[27] br[27] wl[157] vdd gnd cell_6t
Xbit_r158_c27 bl[27] br[27] wl[158] vdd gnd cell_6t
Xbit_r159_c27 bl[27] br[27] wl[159] vdd gnd cell_6t
Xbit_r160_c27 bl[27] br[27] wl[160] vdd gnd cell_6t
Xbit_r161_c27 bl[27] br[27] wl[161] vdd gnd cell_6t
Xbit_r162_c27 bl[27] br[27] wl[162] vdd gnd cell_6t
Xbit_r163_c27 bl[27] br[27] wl[163] vdd gnd cell_6t
Xbit_r164_c27 bl[27] br[27] wl[164] vdd gnd cell_6t
Xbit_r165_c27 bl[27] br[27] wl[165] vdd gnd cell_6t
Xbit_r166_c27 bl[27] br[27] wl[166] vdd gnd cell_6t
Xbit_r167_c27 bl[27] br[27] wl[167] vdd gnd cell_6t
Xbit_r168_c27 bl[27] br[27] wl[168] vdd gnd cell_6t
Xbit_r169_c27 bl[27] br[27] wl[169] vdd gnd cell_6t
Xbit_r170_c27 bl[27] br[27] wl[170] vdd gnd cell_6t
Xbit_r171_c27 bl[27] br[27] wl[171] vdd gnd cell_6t
Xbit_r172_c27 bl[27] br[27] wl[172] vdd gnd cell_6t
Xbit_r173_c27 bl[27] br[27] wl[173] vdd gnd cell_6t
Xbit_r174_c27 bl[27] br[27] wl[174] vdd gnd cell_6t
Xbit_r175_c27 bl[27] br[27] wl[175] vdd gnd cell_6t
Xbit_r176_c27 bl[27] br[27] wl[176] vdd gnd cell_6t
Xbit_r177_c27 bl[27] br[27] wl[177] vdd gnd cell_6t
Xbit_r178_c27 bl[27] br[27] wl[178] vdd gnd cell_6t
Xbit_r179_c27 bl[27] br[27] wl[179] vdd gnd cell_6t
Xbit_r180_c27 bl[27] br[27] wl[180] vdd gnd cell_6t
Xbit_r181_c27 bl[27] br[27] wl[181] vdd gnd cell_6t
Xbit_r182_c27 bl[27] br[27] wl[182] vdd gnd cell_6t
Xbit_r183_c27 bl[27] br[27] wl[183] vdd gnd cell_6t
Xbit_r184_c27 bl[27] br[27] wl[184] vdd gnd cell_6t
Xbit_r185_c27 bl[27] br[27] wl[185] vdd gnd cell_6t
Xbit_r186_c27 bl[27] br[27] wl[186] vdd gnd cell_6t
Xbit_r187_c27 bl[27] br[27] wl[187] vdd gnd cell_6t
Xbit_r188_c27 bl[27] br[27] wl[188] vdd gnd cell_6t
Xbit_r189_c27 bl[27] br[27] wl[189] vdd gnd cell_6t
Xbit_r190_c27 bl[27] br[27] wl[190] vdd gnd cell_6t
Xbit_r191_c27 bl[27] br[27] wl[191] vdd gnd cell_6t
Xbit_r192_c27 bl[27] br[27] wl[192] vdd gnd cell_6t
Xbit_r193_c27 bl[27] br[27] wl[193] vdd gnd cell_6t
Xbit_r194_c27 bl[27] br[27] wl[194] vdd gnd cell_6t
Xbit_r195_c27 bl[27] br[27] wl[195] vdd gnd cell_6t
Xbit_r196_c27 bl[27] br[27] wl[196] vdd gnd cell_6t
Xbit_r197_c27 bl[27] br[27] wl[197] vdd gnd cell_6t
Xbit_r198_c27 bl[27] br[27] wl[198] vdd gnd cell_6t
Xbit_r199_c27 bl[27] br[27] wl[199] vdd gnd cell_6t
Xbit_r200_c27 bl[27] br[27] wl[200] vdd gnd cell_6t
Xbit_r201_c27 bl[27] br[27] wl[201] vdd gnd cell_6t
Xbit_r202_c27 bl[27] br[27] wl[202] vdd gnd cell_6t
Xbit_r203_c27 bl[27] br[27] wl[203] vdd gnd cell_6t
Xbit_r204_c27 bl[27] br[27] wl[204] vdd gnd cell_6t
Xbit_r205_c27 bl[27] br[27] wl[205] vdd gnd cell_6t
Xbit_r206_c27 bl[27] br[27] wl[206] vdd gnd cell_6t
Xbit_r207_c27 bl[27] br[27] wl[207] vdd gnd cell_6t
Xbit_r208_c27 bl[27] br[27] wl[208] vdd gnd cell_6t
Xbit_r209_c27 bl[27] br[27] wl[209] vdd gnd cell_6t
Xbit_r210_c27 bl[27] br[27] wl[210] vdd gnd cell_6t
Xbit_r211_c27 bl[27] br[27] wl[211] vdd gnd cell_6t
Xbit_r212_c27 bl[27] br[27] wl[212] vdd gnd cell_6t
Xbit_r213_c27 bl[27] br[27] wl[213] vdd gnd cell_6t
Xbit_r214_c27 bl[27] br[27] wl[214] vdd gnd cell_6t
Xbit_r215_c27 bl[27] br[27] wl[215] vdd gnd cell_6t
Xbit_r216_c27 bl[27] br[27] wl[216] vdd gnd cell_6t
Xbit_r217_c27 bl[27] br[27] wl[217] vdd gnd cell_6t
Xbit_r218_c27 bl[27] br[27] wl[218] vdd gnd cell_6t
Xbit_r219_c27 bl[27] br[27] wl[219] vdd gnd cell_6t
Xbit_r220_c27 bl[27] br[27] wl[220] vdd gnd cell_6t
Xbit_r221_c27 bl[27] br[27] wl[221] vdd gnd cell_6t
Xbit_r222_c27 bl[27] br[27] wl[222] vdd gnd cell_6t
Xbit_r223_c27 bl[27] br[27] wl[223] vdd gnd cell_6t
Xbit_r224_c27 bl[27] br[27] wl[224] vdd gnd cell_6t
Xbit_r225_c27 bl[27] br[27] wl[225] vdd gnd cell_6t
Xbit_r226_c27 bl[27] br[27] wl[226] vdd gnd cell_6t
Xbit_r227_c27 bl[27] br[27] wl[227] vdd gnd cell_6t
Xbit_r228_c27 bl[27] br[27] wl[228] vdd gnd cell_6t
Xbit_r229_c27 bl[27] br[27] wl[229] vdd gnd cell_6t
Xbit_r230_c27 bl[27] br[27] wl[230] vdd gnd cell_6t
Xbit_r231_c27 bl[27] br[27] wl[231] vdd gnd cell_6t
Xbit_r232_c27 bl[27] br[27] wl[232] vdd gnd cell_6t
Xbit_r233_c27 bl[27] br[27] wl[233] vdd gnd cell_6t
Xbit_r234_c27 bl[27] br[27] wl[234] vdd gnd cell_6t
Xbit_r235_c27 bl[27] br[27] wl[235] vdd gnd cell_6t
Xbit_r236_c27 bl[27] br[27] wl[236] vdd gnd cell_6t
Xbit_r237_c27 bl[27] br[27] wl[237] vdd gnd cell_6t
Xbit_r238_c27 bl[27] br[27] wl[238] vdd gnd cell_6t
Xbit_r239_c27 bl[27] br[27] wl[239] vdd gnd cell_6t
Xbit_r240_c27 bl[27] br[27] wl[240] vdd gnd cell_6t
Xbit_r241_c27 bl[27] br[27] wl[241] vdd gnd cell_6t
Xbit_r242_c27 bl[27] br[27] wl[242] vdd gnd cell_6t
Xbit_r243_c27 bl[27] br[27] wl[243] vdd gnd cell_6t
Xbit_r244_c27 bl[27] br[27] wl[244] vdd gnd cell_6t
Xbit_r245_c27 bl[27] br[27] wl[245] vdd gnd cell_6t
Xbit_r246_c27 bl[27] br[27] wl[246] vdd gnd cell_6t
Xbit_r247_c27 bl[27] br[27] wl[247] vdd gnd cell_6t
Xbit_r248_c27 bl[27] br[27] wl[248] vdd gnd cell_6t
Xbit_r249_c27 bl[27] br[27] wl[249] vdd gnd cell_6t
Xbit_r250_c27 bl[27] br[27] wl[250] vdd gnd cell_6t
Xbit_r251_c27 bl[27] br[27] wl[251] vdd gnd cell_6t
Xbit_r252_c27 bl[27] br[27] wl[252] vdd gnd cell_6t
Xbit_r253_c27 bl[27] br[27] wl[253] vdd gnd cell_6t
Xbit_r254_c27 bl[27] br[27] wl[254] vdd gnd cell_6t
Xbit_r255_c27 bl[27] br[27] wl[255] vdd gnd cell_6t
Xbit_r256_c27 bl[27] br[27] wl[256] vdd gnd cell_6t
Xbit_r257_c27 bl[27] br[27] wl[257] vdd gnd cell_6t
Xbit_r258_c27 bl[27] br[27] wl[258] vdd gnd cell_6t
Xbit_r259_c27 bl[27] br[27] wl[259] vdd gnd cell_6t
Xbit_r260_c27 bl[27] br[27] wl[260] vdd gnd cell_6t
Xbit_r261_c27 bl[27] br[27] wl[261] vdd gnd cell_6t
Xbit_r262_c27 bl[27] br[27] wl[262] vdd gnd cell_6t
Xbit_r263_c27 bl[27] br[27] wl[263] vdd gnd cell_6t
Xbit_r264_c27 bl[27] br[27] wl[264] vdd gnd cell_6t
Xbit_r265_c27 bl[27] br[27] wl[265] vdd gnd cell_6t
Xbit_r266_c27 bl[27] br[27] wl[266] vdd gnd cell_6t
Xbit_r267_c27 bl[27] br[27] wl[267] vdd gnd cell_6t
Xbit_r268_c27 bl[27] br[27] wl[268] vdd gnd cell_6t
Xbit_r269_c27 bl[27] br[27] wl[269] vdd gnd cell_6t
Xbit_r270_c27 bl[27] br[27] wl[270] vdd gnd cell_6t
Xbit_r271_c27 bl[27] br[27] wl[271] vdd gnd cell_6t
Xbit_r272_c27 bl[27] br[27] wl[272] vdd gnd cell_6t
Xbit_r273_c27 bl[27] br[27] wl[273] vdd gnd cell_6t
Xbit_r274_c27 bl[27] br[27] wl[274] vdd gnd cell_6t
Xbit_r275_c27 bl[27] br[27] wl[275] vdd gnd cell_6t
Xbit_r276_c27 bl[27] br[27] wl[276] vdd gnd cell_6t
Xbit_r277_c27 bl[27] br[27] wl[277] vdd gnd cell_6t
Xbit_r278_c27 bl[27] br[27] wl[278] vdd gnd cell_6t
Xbit_r279_c27 bl[27] br[27] wl[279] vdd gnd cell_6t
Xbit_r280_c27 bl[27] br[27] wl[280] vdd gnd cell_6t
Xbit_r281_c27 bl[27] br[27] wl[281] vdd gnd cell_6t
Xbit_r282_c27 bl[27] br[27] wl[282] vdd gnd cell_6t
Xbit_r283_c27 bl[27] br[27] wl[283] vdd gnd cell_6t
Xbit_r284_c27 bl[27] br[27] wl[284] vdd gnd cell_6t
Xbit_r285_c27 bl[27] br[27] wl[285] vdd gnd cell_6t
Xbit_r286_c27 bl[27] br[27] wl[286] vdd gnd cell_6t
Xbit_r287_c27 bl[27] br[27] wl[287] vdd gnd cell_6t
Xbit_r288_c27 bl[27] br[27] wl[288] vdd gnd cell_6t
Xbit_r289_c27 bl[27] br[27] wl[289] vdd gnd cell_6t
Xbit_r290_c27 bl[27] br[27] wl[290] vdd gnd cell_6t
Xbit_r291_c27 bl[27] br[27] wl[291] vdd gnd cell_6t
Xbit_r292_c27 bl[27] br[27] wl[292] vdd gnd cell_6t
Xbit_r293_c27 bl[27] br[27] wl[293] vdd gnd cell_6t
Xbit_r294_c27 bl[27] br[27] wl[294] vdd gnd cell_6t
Xbit_r295_c27 bl[27] br[27] wl[295] vdd gnd cell_6t
Xbit_r296_c27 bl[27] br[27] wl[296] vdd gnd cell_6t
Xbit_r297_c27 bl[27] br[27] wl[297] vdd gnd cell_6t
Xbit_r298_c27 bl[27] br[27] wl[298] vdd gnd cell_6t
Xbit_r299_c27 bl[27] br[27] wl[299] vdd gnd cell_6t
Xbit_r300_c27 bl[27] br[27] wl[300] vdd gnd cell_6t
Xbit_r301_c27 bl[27] br[27] wl[301] vdd gnd cell_6t
Xbit_r302_c27 bl[27] br[27] wl[302] vdd gnd cell_6t
Xbit_r303_c27 bl[27] br[27] wl[303] vdd gnd cell_6t
Xbit_r304_c27 bl[27] br[27] wl[304] vdd gnd cell_6t
Xbit_r305_c27 bl[27] br[27] wl[305] vdd gnd cell_6t
Xbit_r306_c27 bl[27] br[27] wl[306] vdd gnd cell_6t
Xbit_r307_c27 bl[27] br[27] wl[307] vdd gnd cell_6t
Xbit_r308_c27 bl[27] br[27] wl[308] vdd gnd cell_6t
Xbit_r309_c27 bl[27] br[27] wl[309] vdd gnd cell_6t
Xbit_r310_c27 bl[27] br[27] wl[310] vdd gnd cell_6t
Xbit_r311_c27 bl[27] br[27] wl[311] vdd gnd cell_6t
Xbit_r312_c27 bl[27] br[27] wl[312] vdd gnd cell_6t
Xbit_r313_c27 bl[27] br[27] wl[313] vdd gnd cell_6t
Xbit_r314_c27 bl[27] br[27] wl[314] vdd gnd cell_6t
Xbit_r315_c27 bl[27] br[27] wl[315] vdd gnd cell_6t
Xbit_r316_c27 bl[27] br[27] wl[316] vdd gnd cell_6t
Xbit_r317_c27 bl[27] br[27] wl[317] vdd gnd cell_6t
Xbit_r318_c27 bl[27] br[27] wl[318] vdd gnd cell_6t
Xbit_r319_c27 bl[27] br[27] wl[319] vdd gnd cell_6t
Xbit_r320_c27 bl[27] br[27] wl[320] vdd gnd cell_6t
Xbit_r321_c27 bl[27] br[27] wl[321] vdd gnd cell_6t
Xbit_r322_c27 bl[27] br[27] wl[322] vdd gnd cell_6t
Xbit_r323_c27 bl[27] br[27] wl[323] vdd gnd cell_6t
Xbit_r324_c27 bl[27] br[27] wl[324] vdd gnd cell_6t
Xbit_r325_c27 bl[27] br[27] wl[325] vdd gnd cell_6t
Xbit_r326_c27 bl[27] br[27] wl[326] vdd gnd cell_6t
Xbit_r327_c27 bl[27] br[27] wl[327] vdd gnd cell_6t
Xbit_r328_c27 bl[27] br[27] wl[328] vdd gnd cell_6t
Xbit_r329_c27 bl[27] br[27] wl[329] vdd gnd cell_6t
Xbit_r330_c27 bl[27] br[27] wl[330] vdd gnd cell_6t
Xbit_r331_c27 bl[27] br[27] wl[331] vdd gnd cell_6t
Xbit_r332_c27 bl[27] br[27] wl[332] vdd gnd cell_6t
Xbit_r333_c27 bl[27] br[27] wl[333] vdd gnd cell_6t
Xbit_r334_c27 bl[27] br[27] wl[334] vdd gnd cell_6t
Xbit_r335_c27 bl[27] br[27] wl[335] vdd gnd cell_6t
Xbit_r336_c27 bl[27] br[27] wl[336] vdd gnd cell_6t
Xbit_r337_c27 bl[27] br[27] wl[337] vdd gnd cell_6t
Xbit_r338_c27 bl[27] br[27] wl[338] vdd gnd cell_6t
Xbit_r339_c27 bl[27] br[27] wl[339] vdd gnd cell_6t
Xbit_r340_c27 bl[27] br[27] wl[340] vdd gnd cell_6t
Xbit_r341_c27 bl[27] br[27] wl[341] vdd gnd cell_6t
Xbit_r342_c27 bl[27] br[27] wl[342] vdd gnd cell_6t
Xbit_r343_c27 bl[27] br[27] wl[343] vdd gnd cell_6t
Xbit_r344_c27 bl[27] br[27] wl[344] vdd gnd cell_6t
Xbit_r345_c27 bl[27] br[27] wl[345] vdd gnd cell_6t
Xbit_r346_c27 bl[27] br[27] wl[346] vdd gnd cell_6t
Xbit_r347_c27 bl[27] br[27] wl[347] vdd gnd cell_6t
Xbit_r348_c27 bl[27] br[27] wl[348] vdd gnd cell_6t
Xbit_r349_c27 bl[27] br[27] wl[349] vdd gnd cell_6t
Xbit_r350_c27 bl[27] br[27] wl[350] vdd gnd cell_6t
Xbit_r351_c27 bl[27] br[27] wl[351] vdd gnd cell_6t
Xbit_r352_c27 bl[27] br[27] wl[352] vdd gnd cell_6t
Xbit_r353_c27 bl[27] br[27] wl[353] vdd gnd cell_6t
Xbit_r354_c27 bl[27] br[27] wl[354] vdd gnd cell_6t
Xbit_r355_c27 bl[27] br[27] wl[355] vdd gnd cell_6t
Xbit_r356_c27 bl[27] br[27] wl[356] vdd gnd cell_6t
Xbit_r357_c27 bl[27] br[27] wl[357] vdd gnd cell_6t
Xbit_r358_c27 bl[27] br[27] wl[358] vdd gnd cell_6t
Xbit_r359_c27 bl[27] br[27] wl[359] vdd gnd cell_6t
Xbit_r360_c27 bl[27] br[27] wl[360] vdd gnd cell_6t
Xbit_r361_c27 bl[27] br[27] wl[361] vdd gnd cell_6t
Xbit_r362_c27 bl[27] br[27] wl[362] vdd gnd cell_6t
Xbit_r363_c27 bl[27] br[27] wl[363] vdd gnd cell_6t
Xbit_r364_c27 bl[27] br[27] wl[364] vdd gnd cell_6t
Xbit_r365_c27 bl[27] br[27] wl[365] vdd gnd cell_6t
Xbit_r366_c27 bl[27] br[27] wl[366] vdd gnd cell_6t
Xbit_r367_c27 bl[27] br[27] wl[367] vdd gnd cell_6t
Xbit_r368_c27 bl[27] br[27] wl[368] vdd gnd cell_6t
Xbit_r369_c27 bl[27] br[27] wl[369] vdd gnd cell_6t
Xbit_r370_c27 bl[27] br[27] wl[370] vdd gnd cell_6t
Xbit_r371_c27 bl[27] br[27] wl[371] vdd gnd cell_6t
Xbit_r372_c27 bl[27] br[27] wl[372] vdd gnd cell_6t
Xbit_r373_c27 bl[27] br[27] wl[373] vdd gnd cell_6t
Xbit_r374_c27 bl[27] br[27] wl[374] vdd gnd cell_6t
Xbit_r375_c27 bl[27] br[27] wl[375] vdd gnd cell_6t
Xbit_r376_c27 bl[27] br[27] wl[376] vdd gnd cell_6t
Xbit_r377_c27 bl[27] br[27] wl[377] vdd gnd cell_6t
Xbit_r378_c27 bl[27] br[27] wl[378] vdd gnd cell_6t
Xbit_r379_c27 bl[27] br[27] wl[379] vdd gnd cell_6t
Xbit_r380_c27 bl[27] br[27] wl[380] vdd gnd cell_6t
Xbit_r381_c27 bl[27] br[27] wl[381] vdd gnd cell_6t
Xbit_r382_c27 bl[27] br[27] wl[382] vdd gnd cell_6t
Xbit_r383_c27 bl[27] br[27] wl[383] vdd gnd cell_6t
Xbit_r384_c27 bl[27] br[27] wl[384] vdd gnd cell_6t
Xbit_r385_c27 bl[27] br[27] wl[385] vdd gnd cell_6t
Xbit_r386_c27 bl[27] br[27] wl[386] vdd gnd cell_6t
Xbit_r387_c27 bl[27] br[27] wl[387] vdd gnd cell_6t
Xbit_r388_c27 bl[27] br[27] wl[388] vdd gnd cell_6t
Xbit_r389_c27 bl[27] br[27] wl[389] vdd gnd cell_6t
Xbit_r390_c27 bl[27] br[27] wl[390] vdd gnd cell_6t
Xbit_r391_c27 bl[27] br[27] wl[391] vdd gnd cell_6t
Xbit_r392_c27 bl[27] br[27] wl[392] vdd gnd cell_6t
Xbit_r393_c27 bl[27] br[27] wl[393] vdd gnd cell_6t
Xbit_r394_c27 bl[27] br[27] wl[394] vdd gnd cell_6t
Xbit_r395_c27 bl[27] br[27] wl[395] vdd gnd cell_6t
Xbit_r396_c27 bl[27] br[27] wl[396] vdd gnd cell_6t
Xbit_r397_c27 bl[27] br[27] wl[397] vdd gnd cell_6t
Xbit_r398_c27 bl[27] br[27] wl[398] vdd gnd cell_6t
Xbit_r399_c27 bl[27] br[27] wl[399] vdd gnd cell_6t
Xbit_r400_c27 bl[27] br[27] wl[400] vdd gnd cell_6t
Xbit_r401_c27 bl[27] br[27] wl[401] vdd gnd cell_6t
Xbit_r402_c27 bl[27] br[27] wl[402] vdd gnd cell_6t
Xbit_r403_c27 bl[27] br[27] wl[403] vdd gnd cell_6t
Xbit_r404_c27 bl[27] br[27] wl[404] vdd gnd cell_6t
Xbit_r405_c27 bl[27] br[27] wl[405] vdd gnd cell_6t
Xbit_r406_c27 bl[27] br[27] wl[406] vdd gnd cell_6t
Xbit_r407_c27 bl[27] br[27] wl[407] vdd gnd cell_6t
Xbit_r408_c27 bl[27] br[27] wl[408] vdd gnd cell_6t
Xbit_r409_c27 bl[27] br[27] wl[409] vdd gnd cell_6t
Xbit_r410_c27 bl[27] br[27] wl[410] vdd gnd cell_6t
Xbit_r411_c27 bl[27] br[27] wl[411] vdd gnd cell_6t
Xbit_r412_c27 bl[27] br[27] wl[412] vdd gnd cell_6t
Xbit_r413_c27 bl[27] br[27] wl[413] vdd gnd cell_6t
Xbit_r414_c27 bl[27] br[27] wl[414] vdd gnd cell_6t
Xbit_r415_c27 bl[27] br[27] wl[415] vdd gnd cell_6t
Xbit_r416_c27 bl[27] br[27] wl[416] vdd gnd cell_6t
Xbit_r417_c27 bl[27] br[27] wl[417] vdd gnd cell_6t
Xbit_r418_c27 bl[27] br[27] wl[418] vdd gnd cell_6t
Xbit_r419_c27 bl[27] br[27] wl[419] vdd gnd cell_6t
Xbit_r420_c27 bl[27] br[27] wl[420] vdd gnd cell_6t
Xbit_r421_c27 bl[27] br[27] wl[421] vdd gnd cell_6t
Xbit_r422_c27 bl[27] br[27] wl[422] vdd gnd cell_6t
Xbit_r423_c27 bl[27] br[27] wl[423] vdd gnd cell_6t
Xbit_r424_c27 bl[27] br[27] wl[424] vdd gnd cell_6t
Xbit_r425_c27 bl[27] br[27] wl[425] vdd gnd cell_6t
Xbit_r426_c27 bl[27] br[27] wl[426] vdd gnd cell_6t
Xbit_r427_c27 bl[27] br[27] wl[427] vdd gnd cell_6t
Xbit_r428_c27 bl[27] br[27] wl[428] vdd gnd cell_6t
Xbit_r429_c27 bl[27] br[27] wl[429] vdd gnd cell_6t
Xbit_r430_c27 bl[27] br[27] wl[430] vdd gnd cell_6t
Xbit_r431_c27 bl[27] br[27] wl[431] vdd gnd cell_6t
Xbit_r432_c27 bl[27] br[27] wl[432] vdd gnd cell_6t
Xbit_r433_c27 bl[27] br[27] wl[433] vdd gnd cell_6t
Xbit_r434_c27 bl[27] br[27] wl[434] vdd gnd cell_6t
Xbit_r435_c27 bl[27] br[27] wl[435] vdd gnd cell_6t
Xbit_r436_c27 bl[27] br[27] wl[436] vdd gnd cell_6t
Xbit_r437_c27 bl[27] br[27] wl[437] vdd gnd cell_6t
Xbit_r438_c27 bl[27] br[27] wl[438] vdd gnd cell_6t
Xbit_r439_c27 bl[27] br[27] wl[439] vdd gnd cell_6t
Xbit_r440_c27 bl[27] br[27] wl[440] vdd gnd cell_6t
Xbit_r441_c27 bl[27] br[27] wl[441] vdd gnd cell_6t
Xbit_r442_c27 bl[27] br[27] wl[442] vdd gnd cell_6t
Xbit_r443_c27 bl[27] br[27] wl[443] vdd gnd cell_6t
Xbit_r444_c27 bl[27] br[27] wl[444] vdd gnd cell_6t
Xbit_r445_c27 bl[27] br[27] wl[445] vdd gnd cell_6t
Xbit_r446_c27 bl[27] br[27] wl[446] vdd gnd cell_6t
Xbit_r447_c27 bl[27] br[27] wl[447] vdd gnd cell_6t
Xbit_r448_c27 bl[27] br[27] wl[448] vdd gnd cell_6t
Xbit_r449_c27 bl[27] br[27] wl[449] vdd gnd cell_6t
Xbit_r450_c27 bl[27] br[27] wl[450] vdd gnd cell_6t
Xbit_r451_c27 bl[27] br[27] wl[451] vdd gnd cell_6t
Xbit_r452_c27 bl[27] br[27] wl[452] vdd gnd cell_6t
Xbit_r453_c27 bl[27] br[27] wl[453] vdd gnd cell_6t
Xbit_r454_c27 bl[27] br[27] wl[454] vdd gnd cell_6t
Xbit_r455_c27 bl[27] br[27] wl[455] vdd gnd cell_6t
Xbit_r456_c27 bl[27] br[27] wl[456] vdd gnd cell_6t
Xbit_r457_c27 bl[27] br[27] wl[457] vdd gnd cell_6t
Xbit_r458_c27 bl[27] br[27] wl[458] vdd gnd cell_6t
Xbit_r459_c27 bl[27] br[27] wl[459] vdd gnd cell_6t
Xbit_r460_c27 bl[27] br[27] wl[460] vdd gnd cell_6t
Xbit_r461_c27 bl[27] br[27] wl[461] vdd gnd cell_6t
Xbit_r462_c27 bl[27] br[27] wl[462] vdd gnd cell_6t
Xbit_r463_c27 bl[27] br[27] wl[463] vdd gnd cell_6t
Xbit_r464_c27 bl[27] br[27] wl[464] vdd gnd cell_6t
Xbit_r465_c27 bl[27] br[27] wl[465] vdd gnd cell_6t
Xbit_r466_c27 bl[27] br[27] wl[466] vdd gnd cell_6t
Xbit_r467_c27 bl[27] br[27] wl[467] vdd gnd cell_6t
Xbit_r468_c27 bl[27] br[27] wl[468] vdd gnd cell_6t
Xbit_r469_c27 bl[27] br[27] wl[469] vdd gnd cell_6t
Xbit_r470_c27 bl[27] br[27] wl[470] vdd gnd cell_6t
Xbit_r471_c27 bl[27] br[27] wl[471] vdd gnd cell_6t
Xbit_r472_c27 bl[27] br[27] wl[472] vdd gnd cell_6t
Xbit_r473_c27 bl[27] br[27] wl[473] vdd gnd cell_6t
Xbit_r474_c27 bl[27] br[27] wl[474] vdd gnd cell_6t
Xbit_r475_c27 bl[27] br[27] wl[475] vdd gnd cell_6t
Xbit_r476_c27 bl[27] br[27] wl[476] vdd gnd cell_6t
Xbit_r477_c27 bl[27] br[27] wl[477] vdd gnd cell_6t
Xbit_r478_c27 bl[27] br[27] wl[478] vdd gnd cell_6t
Xbit_r479_c27 bl[27] br[27] wl[479] vdd gnd cell_6t
Xbit_r480_c27 bl[27] br[27] wl[480] vdd gnd cell_6t
Xbit_r481_c27 bl[27] br[27] wl[481] vdd gnd cell_6t
Xbit_r482_c27 bl[27] br[27] wl[482] vdd gnd cell_6t
Xbit_r483_c27 bl[27] br[27] wl[483] vdd gnd cell_6t
Xbit_r484_c27 bl[27] br[27] wl[484] vdd gnd cell_6t
Xbit_r485_c27 bl[27] br[27] wl[485] vdd gnd cell_6t
Xbit_r486_c27 bl[27] br[27] wl[486] vdd gnd cell_6t
Xbit_r487_c27 bl[27] br[27] wl[487] vdd gnd cell_6t
Xbit_r488_c27 bl[27] br[27] wl[488] vdd gnd cell_6t
Xbit_r489_c27 bl[27] br[27] wl[489] vdd gnd cell_6t
Xbit_r490_c27 bl[27] br[27] wl[490] vdd gnd cell_6t
Xbit_r491_c27 bl[27] br[27] wl[491] vdd gnd cell_6t
Xbit_r492_c27 bl[27] br[27] wl[492] vdd gnd cell_6t
Xbit_r493_c27 bl[27] br[27] wl[493] vdd gnd cell_6t
Xbit_r494_c27 bl[27] br[27] wl[494] vdd gnd cell_6t
Xbit_r495_c27 bl[27] br[27] wl[495] vdd gnd cell_6t
Xbit_r496_c27 bl[27] br[27] wl[496] vdd gnd cell_6t
Xbit_r497_c27 bl[27] br[27] wl[497] vdd gnd cell_6t
Xbit_r498_c27 bl[27] br[27] wl[498] vdd gnd cell_6t
Xbit_r499_c27 bl[27] br[27] wl[499] vdd gnd cell_6t
Xbit_r500_c27 bl[27] br[27] wl[500] vdd gnd cell_6t
Xbit_r501_c27 bl[27] br[27] wl[501] vdd gnd cell_6t
Xbit_r502_c27 bl[27] br[27] wl[502] vdd gnd cell_6t
Xbit_r503_c27 bl[27] br[27] wl[503] vdd gnd cell_6t
Xbit_r504_c27 bl[27] br[27] wl[504] vdd gnd cell_6t
Xbit_r505_c27 bl[27] br[27] wl[505] vdd gnd cell_6t
Xbit_r506_c27 bl[27] br[27] wl[506] vdd gnd cell_6t
Xbit_r507_c27 bl[27] br[27] wl[507] vdd gnd cell_6t
Xbit_r508_c27 bl[27] br[27] wl[508] vdd gnd cell_6t
Xbit_r509_c27 bl[27] br[27] wl[509] vdd gnd cell_6t
Xbit_r510_c27 bl[27] br[27] wl[510] vdd gnd cell_6t
Xbit_r511_c27 bl[27] br[27] wl[511] vdd gnd cell_6t
Xbit_r0_c28 bl[28] br[28] wl[0] vdd gnd cell_6t
Xbit_r1_c28 bl[28] br[28] wl[1] vdd gnd cell_6t
Xbit_r2_c28 bl[28] br[28] wl[2] vdd gnd cell_6t
Xbit_r3_c28 bl[28] br[28] wl[3] vdd gnd cell_6t
Xbit_r4_c28 bl[28] br[28] wl[4] vdd gnd cell_6t
Xbit_r5_c28 bl[28] br[28] wl[5] vdd gnd cell_6t
Xbit_r6_c28 bl[28] br[28] wl[6] vdd gnd cell_6t
Xbit_r7_c28 bl[28] br[28] wl[7] vdd gnd cell_6t
Xbit_r8_c28 bl[28] br[28] wl[8] vdd gnd cell_6t
Xbit_r9_c28 bl[28] br[28] wl[9] vdd gnd cell_6t
Xbit_r10_c28 bl[28] br[28] wl[10] vdd gnd cell_6t
Xbit_r11_c28 bl[28] br[28] wl[11] vdd gnd cell_6t
Xbit_r12_c28 bl[28] br[28] wl[12] vdd gnd cell_6t
Xbit_r13_c28 bl[28] br[28] wl[13] vdd gnd cell_6t
Xbit_r14_c28 bl[28] br[28] wl[14] vdd gnd cell_6t
Xbit_r15_c28 bl[28] br[28] wl[15] vdd gnd cell_6t
Xbit_r16_c28 bl[28] br[28] wl[16] vdd gnd cell_6t
Xbit_r17_c28 bl[28] br[28] wl[17] vdd gnd cell_6t
Xbit_r18_c28 bl[28] br[28] wl[18] vdd gnd cell_6t
Xbit_r19_c28 bl[28] br[28] wl[19] vdd gnd cell_6t
Xbit_r20_c28 bl[28] br[28] wl[20] vdd gnd cell_6t
Xbit_r21_c28 bl[28] br[28] wl[21] vdd gnd cell_6t
Xbit_r22_c28 bl[28] br[28] wl[22] vdd gnd cell_6t
Xbit_r23_c28 bl[28] br[28] wl[23] vdd gnd cell_6t
Xbit_r24_c28 bl[28] br[28] wl[24] vdd gnd cell_6t
Xbit_r25_c28 bl[28] br[28] wl[25] vdd gnd cell_6t
Xbit_r26_c28 bl[28] br[28] wl[26] vdd gnd cell_6t
Xbit_r27_c28 bl[28] br[28] wl[27] vdd gnd cell_6t
Xbit_r28_c28 bl[28] br[28] wl[28] vdd gnd cell_6t
Xbit_r29_c28 bl[28] br[28] wl[29] vdd gnd cell_6t
Xbit_r30_c28 bl[28] br[28] wl[30] vdd gnd cell_6t
Xbit_r31_c28 bl[28] br[28] wl[31] vdd gnd cell_6t
Xbit_r32_c28 bl[28] br[28] wl[32] vdd gnd cell_6t
Xbit_r33_c28 bl[28] br[28] wl[33] vdd gnd cell_6t
Xbit_r34_c28 bl[28] br[28] wl[34] vdd gnd cell_6t
Xbit_r35_c28 bl[28] br[28] wl[35] vdd gnd cell_6t
Xbit_r36_c28 bl[28] br[28] wl[36] vdd gnd cell_6t
Xbit_r37_c28 bl[28] br[28] wl[37] vdd gnd cell_6t
Xbit_r38_c28 bl[28] br[28] wl[38] vdd gnd cell_6t
Xbit_r39_c28 bl[28] br[28] wl[39] vdd gnd cell_6t
Xbit_r40_c28 bl[28] br[28] wl[40] vdd gnd cell_6t
Xbit_r41_c28 bl[28] br[28] wl[41] vdd gnd cell_6t
Xbit_r42_c28 bl[28] br[28] wl[42] vdd gnd cell_6t
Xbit_r43_c28 bl[28] br[28] wl[43] vdd gnd cell_6t
Xbit_r44_c28 bl[28] br[28] wl[44] vdd gnd cell_6t
Xbit_r45_c28 bl[28] br[28] wl[45] vdd gnd cell_6t
Xbit_r46_c28 bl[28] br[28] wl[46] vdd gnd cell_6t
Xbit_r47_c28 bl[28] br[28] wl[47] vdd gnd cell_6t
Xbit_r48_c28 bl[28] br[28] wl[48] vdd gnd cell_6t
Xbit_r49_c28 bl[28] br[28] wl[49] vdd gnd cell_6t
Xbit_r50_c28 bl[28] br[28] wl[50] vdd gnd cell_6t
Xbit_r51_c28 bl[28] br[28] wl[51] vdd gnd cell_6t
Xbit_r52_c28 bl[28] br[28] wl[52] vdd gnd cell_6t
Xbit_r53_c28 bl[28] br[28] wl[53] vdd gnd cell_6t
Xbit_r54_c28 bl[28] br[28] wl[54] vdd gnd cell_6t
Xbit_r55_c28 bl[28] br[28] wl[55] vdd gnd cell_6t
Xbit_r56_c28 bl[28] br[28] wl[56] vdd gnd cell_6t
Xbit_r57_c28 bl[28] br[28] wl[57] vdd gnd cell_6t
Xbit_r58_c28 bl[28] br[28] wl[58] vdd gnd cell_6t
Xbit_r59_c28 bl[28] br[28] wl[59] vdd gnd cell_6t
Xbit_r60_c28 bl[28] br[28] wl[60] vdd gnd cell_6t
Xbit_r61_c28 bl[28] br[28] wl[61] vdd gnd cell_6t
Xbit_r62_c28 bl[28] br[28] wl[62] vdd gnd cell_6t
Xbit_r63_c28 bl[28] br[28] wl[63] vdd gnd cell_6t
Xbit_r64_c28 bl[28] br[28] wl[64] vdd gnd cell_6t
Xbit_r65_c28 bl[28] br[28] wl[65] vdd gnd cell_6t
Xbit_r66_c28 bl[28] br[28] wl[66] vdd gnd cell_6t
Xbit_r67_c28 bl[28] br[28] wl[67] vdd gnd cell_6t
Xbit_r68_c28 bl[28] br[28] wl[68] vdd gnd cell_6t
Xbit_r69_c28 bl[28] br[28] wl[69] vdd gnd cell_6t
Xbit_r70_c28 bl[28] br[28] wl[70] vdd gnd cell_6t
Xbit_r71_c28 bl[28] br[28] wl[71] vdd gnd cell_6t
Xbit_r72_c28 bl[28] br[28] wl[72] vdd gnd cell_6t
Xbit_r73_c28 bl[28] br[28] wl[73] vdd gnd cell_6t
Xbit_r74_c28 bl[28] br[28] wl[74] vdd gnd cell_6t
Xbit_r75_c28 bl[28] br[28] wl[75] vdd gnd cell_6t
Xbit_r76_c28 bl[28] br[28] wl[76] vdd gnd cell_6t
Xbit_r77_c28 bl[28] br[28] wl[77] vdd gnd cell_6t
Xbit_r78_c28 bl[28] br[28] wl[78] vdd gnd cell_6t
Xbit_r79_c28 bl[28] br[28] wl[79] vdd gnd cell_6t
Xbit_r80_c28 bl[28] br[28] wl[80] vdd gnd cell_6t
Xbit_r81_c28 bl[28] br[28] wl[81] vdd gnd cell_6t
Xbit_r82_c28 bl[28] br[28] wl[82] vdd gnd cell_6t
Xbit_r83_c28 bl[28] br[28] wl[83] vdd gnd cell_6t
Xbit_r84_c28 bl[28] br[28] wl[84] vdd gnd cell_6t
Xbit_r85_c28 bl[28] br[28] wl[85] vdd gnd cell_6t
Xbit_r86_c28 bl[28] br[28] wl[86] vdd gnd cell_6t
Xbit_r87_c28 bl[28] br[28] wl[87] vdd gnd cell_6t
Xbit_r88_c28 bl[28] br[28] wl[88] vdd gnd cell_6t
Xbit_r89_c28 bl[28] br[28] wl[89] vdd gnd cell_6t
Xbit_r90_c28 bl[28] br[28] wl[90] vdd gnd cell_6t
Xbit_r91_c28 bl[28] br[28] wl[91] vdd gnd cell_6t
Xbit_r92_c28 bl[28] br[28] wl[92] vdd gnd cell_6t
Xbit_r93_c28 bl[28] br[28] wl[93] vdd gnd cell_6t
Xbit_r94_c28 bl[28] br[28] wl[94] vdd gnd cell_6t
Xbit_r95_c28 bl[28] br[28] wl[95] vdd gnd cell_6t
Xbit_r96_c28 bl[28] br[28] wl[96] vdd gnd cell_6t
Xbit_r97_c28 bl[28] br[28] wl[97] vdd gnd cell_6t
Xbit_r98_c28 bl[28] br[28] wl[98] vdd gnd cell_6t
Xbit_r99_c28 bl[28] br[28] wl[99] vdd gnd cell_6t
Xbit_r100_c28 bl[28] br[28] wl[100] vdd gnd cell_6t
Xbit_r101_c28 bl[28] br[28] wl[101] vdd gnd cell_6t
Xbit_r102_c28 bl[28] br[28] wl[102] vdd gnd cell_6t
Xbit_r103_c28 bl[28] br[28] wl[103] vdd gnd cell_6t
Xbit_r104_c28 bl[28] br[28] wl[104] vdd gnd cell_6t
Xbit_r105_c28 bl[28] br[28] wl[105] vdd gnd cell_6t
Xbit_r106_c28 bl[28] br[28] wl[106] vdd gnd cell_6t
Xbit_r107_c28 bl[28] br[28] wl[107] vdd gnd cell_6t
Xbit_r108_c28 bl[28] br[28] wl[108] vdd gnd cell_6t
Xbit_r109_c28 bl[28] br[28] wl[109] vdd gnd cell_6t
Xbit_r110_c28 bl[28] br[28] wl[110] vdd gnd cell_6t
Xbit_r111_c28 bl[28] br[28] wl[111] vdd gnd cell_6t
Xbit_r112_c28 bl[28] br[28] wl[112] vdd gnd cell_6t
Xbit_r113_c28 bl[28] br[28] wl[113] vdd gnd cell_6t
Xbit_r114_c28 bl[28] br[28] wl[114] vdd gnd cell_6t
Xbit_r115_c28 bl[28] br[28] wl[115] vdd gnd cell_6t
Xbit_r116_c28 bl[28] br[28] wl[116] vdd gnd cell_6t
Xbit_r117_c28 bl[28] br[28] wl[117] vdd gnd cell_6t
Xbit_r118_c28 bl[28] br[28] wl[118] vdd gnd cell_6t
Xbit_r119_c28 bl[28] br[28] wl[119] vdd gnd cell_6t
Xbit_r120_c28 bl[28] br[28] wl[120] vdd gnd cell_6t
Xbit_r121_c28 bl[28] br[28] wl[121] vdd gnd cell_6t
Xbit_r122_c28 bl[28] br[28] wl[122] vdd gnd cell_6t
Xbit_r123_c28 bl[28] br[28] wl[123] vdd gnd cell_6t
Xbit_r124_c28 bl[28] br[28] wl[124] vdd gnd cell_6t
Xbit_r125_c28 bl[28] br[28] wl[125] vdd gnd cell_6t
Xbit_r126_c28 bl[28] br[28] wl[126] vdd gnd cell_6t
Xbit_r127_c28 bl[28] br[28] wl[127] vdd gnd cell_6t
Xbit_r128_c28 bl[28] br[28] wl[128] vdd gnd cell_6t
Xbit_r129_c28 bl[28] br[28] wl[129] vdd gnd cell_6t
Xbit_r130_c28 bl[28] br[28] wl[130] vdd gnd cell_6t
Xbit_r131_c28 bl[28] br[28] wl[131] vdd gnd cell_6t
Xbit_r132_c28 bl[28] br[28] wl[132] vdd gnd cell_6t
Xbit_r133_c28 bl[28] br[28] wl[133] vdd gnd cell_6t
Xbit_r134_c28 bl[28] br[28] wl[134] vdd gnd cell_6t
Xbit_r135_c28 bl[28] br[28] wl[135] vdd gnd cell_6t
Xbit_r136_c28 bl[28] br[28] wl[136] vdd gnd cell_6t
Xbit_r137_c28 bl[28] br[28] wl[137] vdd gnd cell_6t
Xbit_r138_c28 bl[28] br[28] wl[138] vdd gnd cell_6t
Xbit_r139_c28 bl[28] br[28] wl[139] vdd gnd cell_6t
Xbit_r140_c28 bl[28] br[28] wl[140] vdd gnd cell_6t
Xbit_r141_c28 bl[28] br[28] wl[141] vdd gnd cell_6t
Xbit_r142_c28 bl[28] br[28] wl[142] vdd gnd cell_6t
Xbit_r143_c28 bl[28] br[28] wl[143] vdd gnd cell_6t
Xbit_r144_c28 bl[28] br[28] wl[144] vdd gnd cell_6t
Xbit_r145_c28 bl[28] br[28] wl[145] vdd gnd cell_6t
Xbit_r146_c28 bl[28] br[28] wl[146] vdd gnd cell_6t
Xbit_r147_c28 bl[28] br[28] wl[147] vdd gnd cell_6t
Xbit_r148_c28 bl[28] br[28] wl[148] vdd gnd cell_6t
Xbit_r149_c28 bl[28] br[28] wl[149] vdd gnd cell_6t
Xbit_r150_c28 bl[28] br[28] wl[150] vdd gnd cell_6t
Xbit_r151_c28 bl[28] br[28] wl[151] vdd gnd cell_6t
Xbit_r152_c28 bl[28] br[28] wl[152] vdd gnd cell_6t
Xbit_r153_c28 bl[28] br[28] wl[153] vdd gnd cell_6t
Xbit_r154_c28 bl[28] br[28] wl[154] vdd gnd cell_6t
Xbit_r155_c28 bl[28] br[28] wl[155] vdd gnd cell_6t
Xbit_r156_c28 bl[28] br[28] wl[156] vdd gnd cell_6t
Xbit_r157_c28 bl[28] br[28] wl[157] vdd gnd cell_6t
Xbit_r158_c28 bl[28] br[28] wl[158] vdd gnd cell_6t
Xbit_r159_c28 bl[28] br[28] wl[159] vdd gnd cell_6t
Xbit_r160_c28 bl[28] br[28] wl[160] vdd gnd cell_6t
Xbit_r161_c28 bl[28] br[28] wl[161] vdd gnd cell_6t
Xbit_r162_c28 bl[28] br[28] wl[162] vdd gnd cell_6t
Xbit_r163_c28 bl[28] br[28] wl[163] vdd gnd cell_6t
Xbit_r164_c28 bl[28] br[28] wl[164] vdd gnd cell_6t
Xbit_r165_c28 bl[28] br[28] wl[165] vdd gnd cell_6t
Xbit_r166_c28 bl[28] br[28] wl[166] vdd gnd cell_6t
Xbit_r167_c28 bl[28] br[28] wl[167] vdd gnd cell_6t
Xbit_r168_c28 bl[28] br[28] wl[168] vdd gnd cell_6t
Xbit_r169_c28 bl[28] br[28] wl[169] vdd gnd cell_6t
Xbit_r170_c28 bl[28] br[28] wl[170] vdd gnd cell_6t
Xbit_r171_c28 bl[28] br[28] wl[171] vdd gnd cell_6t
Xbit_r172_c28 bl[28] br[28] wl[172] vdd gnd cell_6t
Xbit_r173_c28 bl[28] br[28] wl[173] vdd gnd cell_6t
Xbit_r174_c28 bl[28] br[28] wl[174] vdd gnd cell_6t
Xbit_r175_c28 bl[28] br[28] wl[175] vdd gnd cell_6t
Xbit_r176_c28 bl[28] br[28] wl[176] vdd gnd cell_6t
Xbit_r177_c28 bl[28] br[28] wl[177] vdd gnd cell_6t
Xbit_r178_c28 bl[28] br[28] wl[178] vdd gnd cell_6t
Xbit_r179_c28 bl[28] br[28] wl[179] vdd gnd cell_6t
Xbit_r180_c28 bl[28] br[28] wl[180] vdd gnd cell_6t
Xbit_r181_c28 bl[28] br[28] wl[181] vdd gnd cell_6t
Xbit_r182_c28 bl[28] br[28] wl[182] vdd gnd cell_6t
Xbit_r183_c28 bl[28] br[28] wl[183] vdd gnd cell_6t
Xbit_r184_c28 bl[28] br[28] wl[184] vdd gnd cell_6t
Xbit_r185_c28 bl[28] br[28] wl[185] vdd gnd cell_6t
Xbit_r186_c28 bl[28] br[28] wl[186] vdd gnd cell_6t
Xbit_r187_c28 bl[28] br[28] wl[187] vdd gnd cell_6t
Xbit_r188_c28 bl[28] br[28] wl[188] vdd gnd cell_6t
Xbit_r189_c28 bl[28] br[28] wl[189] vdd gnd cell_6t
Xbit_r190_c28 bl[28] br[28] wl[190] vdd gnd cell_6t
Xbit_r191_c28 bl[28] br[28] wl[191] vdd gnd cell_6t
Xbit_r192_c28 bl[28] br[28] wl[192] vdd gnd cell_6t
Xbit_r193_c28 bl[28] br[28] wl[193] vdd gnd cell_6t
Xbit_r194_c28 bl[28] br[28] wl[194] vdd gnd cell_6t
Xbit_r195_c28 bl[28] br[28] wl[195] vdd gnd cell_6t
Xbit_r196_c28 bl[28] br[28] wl[196] vdd gnd cell_6t
Xbit_r197_c28 bl[28] br[28] wl[197] vdd gnd cell_6t
Xbit_r198_c28 bl[28] br[28] wl[198] vdd gnd cell_6t
Xbit_r199_c28 bl[28] br[28] wl[199] vdd gnd cell_6t
Xbit_r200_c28 bl[28] br[28] wl[200] vdd gnd cell_6t
Xbit_r201_c28 bl[28] br[28] wl[201] vdd gnd cell_6t
Xbit_r202_c28 bl[28] br[28] wl[202] vdd gnd cell_6t
Xbit_r203_c28 bl[28] br[28] wl[203] vdd gnd cell_6t
Xbit_r204_c28 bl[28] br[28] wl[204] vdd gnd cell_6t
Xbit_r205_c28 bl[28] br[28] wl[205] vdd gnd cell_6t
Xbit_r206_c28 bl[28] br[28] wl[206] vdd gnd cell_6t
Xbit_r207_c28 bl[28] br[28] wl[207] vdd gnd cell_6t
Xbit_r208_c28 bl[28] br[28] wl[208] vdd gnd cell_6t
Xbit_r209_c28 bl[28] br[28] wl[209] vdd gnd cell_6t
Xbit_r210_c28 bl[28] br[28] wl[210] vdd gnd cell_6t
Xbit_r211_c28 bl[28] br[28] wl[211] vdd gnd cell_6t
Xbit_r212_c28 bl[28] br[28] wl[212] vdd gnd cell_6t
Xbit_r213_c28 bl[28] br[28] wl[213] vdd gnd cell_6t
Xbit_r214_c28 bl[28] br[28] wl[214] vdd gnd cell_6t
Xbit_r215_c28 bl[28] br[28] wl[215] vdd gnd cell_6t
Xbit_r216_c28 bl[28] br[28] wl[216] vdd gnd cell_6t
Xbit_r217_c28 bl[28] br[28] wl[217] vdd gnd cell_6t
Xbit_r218_c28 bl[28] br[28] wl[218] vdd gnd cell_6t
Xbit_r219_c28 bl[28] br[28] wl[219] vdd gnd cell_6t
Xbit_r220_c28 bl[28] br[28] wl[220] vdd gnd cell_6t
Xbit_r221_c28 bl[28] br[28] wl[221] vdd gnd cell_6t
Xbit_r222_c28 bl[28] br[28] wl[222] vdd gnd cell_6t
Xbit_r223_c28 bl[28] br[28] wl[223] vdd gnd cell_6t
Xbit_r224_c28 bl[28] br[28] wl[224] vdd gnd cell_6t
Xbit_r225_c28 bl[28] br[28] wl[225] vdd gnd cell_6t
Xbit_r226_c28 bl[28] br[28] wl[226] vdd gnd cell_6t
Xbit_r227_c28 bl[28] br[28] wl[227] vdd gnd cell_6t
Xbit_r228_c28 bl[28] br[28] wl[228] vdd gnd cell_6t
Xbit_r229_c28 bl[28] br[28] wl[229] vdd gnd cell_6t
Xbit_r230_c28 bl[28] br[28] wl[230] vdd gnd cell_6t
Xbit_r231_c28 bl[28] br[28] wl[231] vdd gnd cell_6t
Xbit_r232_c28 bl[28] br[28] wl[232] vdd gnd cell_6t
Xbit_r233_c28 bl[28] br[28] wl[233] vdd gnd cell_6t
Xbit_r234_c28 bl[28] br[28] wl[234] vdd gnd cell_6t
Xbit_r235_c28 bl[28] br[28] wl[235] vdd gnd cell_6t
Xbit_r236_c28 bl[28] br[28] wl[236] vdd gnd cell_6t
Xbit_r237_c28 bl[28] br[28] wl[237] vdd gnd cell_6t
Xbit_r238_c28 bl[28] br[28] wl[238] vdd gnd cell_6t
Xbit_r239_c28 bl[28] br[28] wl[239] vdd gnd cell_6t
Xbit_r240_c28 bl[28] br[28] wl[240] vdd gnd cell_6t
Xbit_r241_c28 bl[28] br[28] wl[241] vdd gnd cell_6t
Xbit_r242_c28 bl[28] br[28] wl[242] vdd gnd cell_6t
Xbit_r243_c28 bl[28] br[28] wl[243] vdd gnd cell_6t
Xbit_r244_c28 bl[28] br[28] wl[244] vdd gnd cell_6t
Xbit_r245_c28 bl[28] br[28] wl[245] vdd gnd cell_6t
Xbit_r246_c28 bl[28] br[28] wl[246] vdd gnd cell_6t
Xbit_r247_c28 bl[28] br[28] wl[247] vdd gnd cell_6t
Xbit_r248_c28 bl[28] br[28] wl[248] vdd gnd cell_6t
Xbit_r249_c28 bl[28] br[28] wl[249] vdd gnd cell_6t
Xbit_r250_c28 bl[28] br[28] wl[250] vdd gnd cell_6t
Xbit_r251_c28 bl[28] br[28] wl[251] vdd gnd cell_6t
Xbit_r252_c28 bl[28] br[28] wl[252] vdd gnd cell_6t
Xbit_r253_c28 bl[28] br[28] wl[253] vdd gnd cell_6t
Xbit_r254_c28 bl[28] br[28] wl[254] vdd gnd cell_6t
Xbit_r255_c28 bl[28] br[28] wl[255] vdd gnd cell_6t
Xbit_r256_c28 bl[28] br[28] wl[256] vdd gnd cell_6t
Xbit_r257_c28 bl[28] br[28] wl[257] vdd gnd cell_6t
Xbit_r258_c28 bl[28] br[28] wl[258] vdd gnd cell_6t
Xbit_r259_c28 bl[28] br[28] wl[259] vdd gnd cell_6t
Xbit_r260_c28 bl[28] br[28] wl[260] vdd gnd cell_6t
Xbit_r261_c28 bl[28] br[28] wl[261] vdd gnd cell_6t
Xbit_r262_c28 bl[28] br[28] wl[262] vdd gnd cell_6t
Xbit_r263_c28 bl[28] br[28] wl[263] vdd gnd cell_6t
Xbit_r264_c28 bl[28] br[28] wl[264] vdd gnd cell_6t
Xbit_r265_c28 bl[28] br[28] wl[265] vdd gnd cell_6t
Xbit_r266_c28 bl[28] br[28] wl[266] vdd gnd cell_6t
Xbit_r267_c28 bl[28] br[28] wl[267] vdd gnd cell_6t
Xbit_r268_c28 bl[28] br[28] wl[268] vdd gnd cell_6t
Xbit_r269_c28 bl[28] br[28] wl[269] vdd gnd cell_6t
Xbit_r270_c28 bl[28] br[28] wl[270] vdd gnd cell_6t
Xbit_r271_c28 bl[28] br[28] wl[271] vdd gnd cell_6t
Xbit_r272_c28 bl[28] br[28] wl[272] vdd gnd cell_6t
Xbit_r273_c28 bl[28] br[28] wl[273] vdd gnd cell_6t
Xbit_r274_c28 bl[28] br[28] wl[274] vdd gnd cell_6t
Xbit_r275_c28 bl[28] br[28] wl[275] vdd gnd cell_6t
Xbit_r276_c28 bl[28] br[28] wl[276] vdd gnd cell_6t
Xbit_r277_c28 bl[28] br[28] wl[277] vdd gnd cell_6t
Xbit_r278_c28 bl[28] br[28] wl[278] vdd gnd cell_6t
Xbit_r279_c28 bl[28] br[28] wl[279] vdd gnd cell_6t
Xbit_r280_c28 bl[28] br[28] wl[280] vdd gnd cell_6t
Xbit_r281_c28 bl[28] br[28] wl[281] vdd gnd cell_6t
Xbit_r282_c28 bl[28] br[28] wl[282] vdd gnd cell_6t
Xbit_r283_c28 bl[28] br[28] wl[283] vdd gnd cell_6t
Xbit_r284_c28 bl[28] br[28] wl[284] vdd gnd cell_6t
Xbit_r285_c28 bl[28] br[28] wl[285] vdd gnd cell_6t
Xbit_r286_c28 bl[28] br[28] wl[286] vdd gnd cell_6t
Xbit_r287_c28 bl[28] br[28] wl[287] vdd gnd cell_6t
Xbit_r288_c28 bl[28] br[28] wl[288] vdd gnd cell_6t
Xbit_r289_c28 bl[28] br[28] wl[289] vdd gnd cell_6t
Xbit_r290_c28 bl[28] br[28] wl[290] vdd gnd cell_6t
Xbit_r291_c28 bl[28] br[28] wl[291] vdd gnd cell_6t
Xbit_r292_c28 bl[28] br[28] wl[292] vdd gnd cell_6t
Xbit_r293_c28 bl[28] br[28] wl[293] vdd gnd cell_6t
Xbit_r294_c28 bl[28] br[28] wl[294] vdd gnd cell_6t
Xbit_r295_c28 bl[28] br[28] wl[295] vdd gnd cell_6t
Xbit_r296_c28 bl[28] br[28] wl[296] vdd gnd cell_6t
Xbit_r297_c28 bl[28] br[28] wl[297] vdd gnd cell_6t
Xbit_r298_c28 bl[28] br[28] wl[298] vdd gnd cell_6t
Xbit_r299_c28 bl[28] br[28] wl[299] vdd gnd cell_6t
Xbit_r300_c28 bl[28] br[28] wl[300] vdd gnd cell_6t
Xbit_r301_c28 bl[28] br[28] wl[301] vdd gnd cell_6t
Xbit_r302_c28 bl[28] br[28] wl[302] vdd gnd cell_6t
Xbit_r303_c28 bl[28] br[28] wl[303] vdd gnd cell_6t
Xbit_r304_c28 bl[28] br[28] wl[304] vdd gnd cell_6t
Xbit_r305_c28 bl[28] br[28] wl[305] vdd gnd cell_6t
Xbit_r306_c28 bl[28] br[28] wl[306] vdd gnd cell_6t
Xbit_r307_c28 bl[28] br[28] wl[307] vdd gnd cell_6t
Xbit_r308_c28 bl[28] br[28] wl[308] vdd gnd cell_6t
Xbit_r309_c28 bl[28] br[28] wl[309] vdd gnd cell_6t
Xbit_r310_c28 bl[28] br[28] wl[310] vdd gnd cell_6t
Xbit_r311_c28 bl[28] br[28] wl[311] vdd gnd cell_6t
Xbit_r312_c28 bl[28] br[28] wl[312] vdd gnd cell_6t
Xbit_r313_c28 bl[28] br[28] wl[313] vdd gnd cell_6t
Xbit_r314_c28 bl[28] br[28] wl[314] vdd gnd cell_6t
Xbit_r315_c28 bl[28] br[28] wl[315] vdd gnd cell_6t
Xbit_r316_c28 bl[28] br[28] wl[316] vdd gnd cell_6t
Xbit_r317_c28 bl[28] br[28] wl[317] vdd gnd cell_6t
Xbit_r318_c28 bl[28] br[28] wl[318] vdd gnd cell_6t
Xbit_r319_c28 bl[28] br[28] wl[319] vdd gnd cell_6t
Xbit_r320_c28 bl[28] br[28] wl[320] vdd gnd cell_6t
Xbit_r321_c28 bl[28] br[28] wl[321] vdd gnd cell_6t
Xbit_r322_c28 bl[28] br[28] wl[322] vdd gnd cell_6t
Xbit_r323_c28 bl[28] br[28] wl[323] vdd gnd cell_6t
Xbit_r324_c28 bl[28] br[28] wl[324] vdd gnd cell_6t
Xbit_r325_c28 bl[28] br[28] wl[325] vdd gnd cell_6t
Xbit_r326_c28 bl[28] br[28] wl[326] vdd gnd cell_6t
Xbit_r327_c28 bl[28] br[28] wl[327] vdd gnd cell_6t
Xbit_r328_c28 bl[28] br[28] wl[328] vdd gnd cell_6t
Xbit_r329_c28 bl[28] br[28] wl[329] vdd gnd cell_6t
Xbit_r330_c28 bl[28] br[28] wl[330] vdd gnd cell_6t
Xbit_r331_c28 bl[28] br[28] wl[331] vdd gnd cell_6t
Xbit_r332_c28 bl[28] br[28] wl[332] vdd gnd cell_6t
Xbit_r333_c28 bl[28] br[28] wl[333] vdd gnd cell_6t
Xbit_r334_c28 bl[28] br[28] wl[334] vdd gnd cell_6t
Xbit_r335_c28 bl[28] br[28] wl[335] vdd gnd cell_6t
Xbit_r336_c28 bl[28] br[28] wl[336] vdd gnd cell_6t
Xbit_r337_c28 bl[28] br[28] wl[337] vdd gnd cell_6t
Xbit_r338_c28 bl[28] br[28] wl[338] vdd gnd cell_6t
Xbit_r339_c28 bl[28] br[28] wl[339] vdd gnd cell_6t
Xbit_r340_c28 bl[28] br[28] wl[340] vdd gnd cell_6t
Xbit_r341_c28 bl[28] br[28] wl[341] vdd gnd cell_6t
Xbit_r342_c28 bl[28] br[28] wl[342] vdd gnd cell_6t
Xbit_r343_c28 bl[28] br[28] wl[343] vdd gnd cell_6t
Xbit_r344_c28 bl[28] br[28] wl[344] vdd gnd cell_6t
Xbit_r345_c28 bl[28] br[28] wl[345] vdd gnd cell_6t
Xbit_r346_c28 bl[28] br[28] wl[346] vdd gnd cell_6t
Xbit_r347_c28 bl[28] br[28] wl[347] vdd gnd cell_6t
Xbit_r348_c28 bl[28] br[28] wl[348] vdd gnd cell_6t
Xbit_r349_c28 bl[28] br[28] wl[349] vdd gnd cell_6t
Xbit_r350_c28 bl[28] br[28] wl[350] vdd gnd cell_6t
Xbit_r351_c28 bl[28] br[28] wl[351] vdd gnd cell_6t
Xbit_r352_c28 bl[28] br[28] wl[352] vdd gnd cell_6t
Xbit_r353_c28 bl[28] br[28] wl[353] vdd gnd cell_6t
Xbit_r354_c28 bl[28] br[28] wl[354] vdd gnd cell_6t
Xbit_r355_c28 bl[28] br[28] wl[355] vdd gnd cell_6t
Xbit_r356_c28 bl[28] br[28] wl[356] vdd gnd cell_6t
Xbit_r357_c28 bl[28] br[28] wl[357] vdd gnd cell_6t
Xbit_r358_c28 bl[28] br[28] wl[358] vdd gnd cell_6t
Xbit_r359_c28 bl[28] br[28] wl[359] vdd gnd cell_6t
Xbit_r360_c28 bl[28] br[28] wl[360] vdd gnd cell_6t
Xbit_r361_c28 bl[28] br[28] wl[361] vdd gnd cell_6t
Xbit_r362_c28 bl[28] br[28] wl[362] vdd gnd cell_6t
Xbit_r363_c28 bl[28] br[28] wl[363] vdd gnd cell_6t
Xbit_r364_c28 bl[28] br[28] wl[364] vdd gnd cell_6t
Xbit_r365_c28 bl[28] br[28] wl[365] vdd gnd cell_6t
Xbit_r366_c28 bl[28] br[28] wl[366] vdd gnd cell_6t
Xbit_r367_c28 bl[28] br[28] wl[367] vdd gnd cell_6t
Xbit_r368_c28 bl[28] br[28] wl[368] vdd gnd cell_6t
Xbit_r369_c28 bl[28] br[28] wl[369] vdd gnd cell_6t
Xbit_r370_c28 bl[28] br[28] wl[370] vdd gnd cell_6t
Xbit_r371_c28 bl[28] br[28] wl[371] vdd gnd cell_6t
Xbit_r372_c28 bl[28] br[28] wl[372] vdd gnd cell_6t
Xbit_r373_c28 bl[28] br[28] wl[373] vdd gnd cell_6t
Xbit_r374_c28 bl[28] br[28] wl[374] vdd gnd cell_6t
Xbit_r375_c28 bl[28] br[28] wl[375] vdd gnd cell_6t
Xbit_r376_c28 bl[28] br[28] wl[376] vdd gnd cell_6t
Xbit_r377_c28 bl[28] br[28] wl[377] vdd gnd cell_6t
Xbit_r378_c28 bl[28] br[28] wl[378] vdd gnd cell_6t
Xbit_r379_c28 bl[28] br[28] wl[379] vdd gnd cell_6t
Xbit_r380_c28 bl[28] br[28] wl[380] vdd gnd cell_6t
Xbit_r381_c28 bl[28] br[28] wl[381] vdd gnd cell_6t
Xbit_r382_c28 bl[28] br[28] wl[382] vdd gnd cell_6t
Xbit_r383_c28 bl[28] br[28] wl[383] vdd gnd cell_6t
Xbit_r384_c28 bl[28] br[28] wl[384] vdd gnd cell_6t
Xbit_r385_c28 bl[28] br[28] wl[385] vdd gnd cell_6t
Xbit_r386_c28 bl[28] br[28] wl[386] vdd gnd cell_6t
Xbit_r387_c28 bl[28] br[28] wl[387] vdd gnd cell_6t
Xbit_r388_c28 bl[28] br[28] wl[388] vdd gnd cell_6t
Xbit_r389_c28 bl[28] br[28] wl[389] vdd gnd cell_6t
Xbit_r390_c28 bl[28] br[28] wl[390] vdd gnd cell_6t
Xbit_r391_c28 bl[28] br[28] wl[391] vdd gnd cell_6t
Xbit_r392_c28 bl[28] br[28] wl[392] vdd gnd cell_6t
Xbit_r393_c28 bl[28] br[28] wl[393] vdd gnd cell_6t
Xbit_r394_c28 bl[28] br[28] wl[394] vdd gnd cell_6t
Xbit_r395_c28 bl[28] br[28] wl[395] vdd gnd cell_6t
Xbit_r396_c28 bl[28] br[28] wl[396] vdd gnd cell_6t
Xbit_r397_c28 bl[28] br[28] wl[397] vdd gnd cell_6t
Xbit_r398_c28 bl[28] br[28] wl[398] vdd gnd cell_6t
Xbit_r399_c28 bl[28] br[28] wl[399] vdd gnd cell_6t
Xbit_r400_c28 bl[28] br[28] wl[400] vdd gnd cell_6t
Xbit_r401_c28 bl[28] br[28] wl[401] vdd gnd cell_6t
Xbit_r402_c28 bl[28] br[28] wl[402] vdd gnd cell_6t
Xbit_r403_c28 bl[28] br[28] wl[403] vdd gnd cell_6t
Xbit_r404_c28 bl[28] br[28] wl[404] vdd gnd cell_6t
Xbit_r405_c28 bl[28] br[28] wl[405] vdd gnd cell_6t
Xbit_r406_c28 bl[28] br[28] wl[406] vdd gnd cell_6t
Xbit_r407_c28 bl[28] br[28] wl[407] vdd gnd cell_6t
Xbit_r408_c28 bl[28] br[28] wl[408] vdd gnd cell_6t
Xbit_r409_c28 bl[28] br[28] wl[409] vdd gnd cell_6t
Xbit_r410_c28 bl[28] br[28] wl[410] vdd gnd cell_6t
Xbit_r411_c28 bl[28] br[28] wl[411] vdd gnd cell_6t
Xbit_r412_c28 bl[28] br[28] wl[412] vdd gnd cell_6t
Xbit_r413_c28 bl[28] br[28] wl[413] vdd gnd cell_6t
Xbit_r414_c28 bl[28] br[28] wl[414] vdd gnd cell_6t
Xbit_r415_c28 bl[28] br[28] wl[415] vdd gnd cell_6t
Xbit_r416_c28 bl[28] br[28] wl[416] vdd gnd cell_6t
Xbit_r417_c28 bl[28] br[28] wl[417] vdd gnd cell_6t
Xbit_r418_c28 bl[28] br[28] wl[418] vdd gnd cell_6t
Xbit_r419_c28 bl[28] br[28] wl[419] vdd gnd cell_6t
Xbit_r420_c28 bl[28] br[28] wl[420] vdd gnd cell_6t
Xbit_r421_c28 bl[28] br[28] wl[421] vdd gnd cell_6t
Xbit_r422_c28 bl[28] br[28] wl[422] vdd gnd cell_6t
Xbit_r423_c28 bl[28] br[28] wl[423] vdd gnd cell_6t
Xbit_r424_c28 bl[28] br[28] wl[424] vdd gnd cell_6t
Xbit_r425_c28 bl[28] br[28] wl[425] vdd gnd cell_6t
Xbit_r426_c28 bl[28] br[28] wl[426] vdd gnd cell_6t
Xbit_r427_c28 bl[28] br[28] wl[427] vdd gnd cell_6t
Xbit_r428_c28 bl[28] br[28] wl[428] vdd gnd cell_6t
Xbit_r429_c28 bl[28] br[28] wl[429] vdd gnd cell_6t
Xbit_r430_c28 bl[28] br[28] wl[430] vdd gnd cell_6t
Xbit_r431_c28 bl[28] br[28] wl[431] vdd gnd cell_6t
Xbit_r432_c28 bl[28] br[28] wl[432] vdd gnd cell_6t
Xbit_r433_c28 bl[28] br[28] wl[433] vdd gnd cell_6t
Xbit_r434_c28 bl[28] br[28] wl[434] vdd gnd cell_6t
Xbit_r435_c28 bl[28] br[28] wl[435] vdd gnd cell_6t
Xbit_r436_c28 bl[28] br[28] wl[436] vdd gnd cell_6t
Xbit_r437_c28 bl[28] br[28] wl[437] vdd gnd cell_6t
Xbit_r438_c28 bl[28] br[28] wl[438] vdd gnd cell_6t
Xbit_r439_c28 bl[28] br[28] wl[439] vdd gnd cell_6t
Xbit_r440_c28 bl[28] br[28] wl[440] vdd gnd cell_6t
Xbit_r441_c28 bl[28] br[28] wl[441] vdd gnd cell_6t
Xbit_r442_c28 bl[28] br[28] wl[442] vdd gnd cell_6t
Xbit_r443_c28 bl[28] br[28] wl[443] vdd gnd cell_6t
Xbit_r444_c28 bl[28] br[28] wl[444] vdd gnd cell_6t
Xbit_r445_c28 bl[28] br[28] wl[445] vdd gnd cell_6t
Xbit_r446_c28 bl[28] br[28] wl[446] vdd gnd cell_6t
Xbit_r447_c28 bl[28] br[28] wl[447] vdd gnd cell_6t
Xbit_r448_c28 bl[28] br[28] wl[448] vdd gnd cell_6t
Xbit_r449_c28 bl[28] br[28] wl[449] vdd gnd cell_6t
Xbit_r450_c28 bl[28] br[28] wl[450] vdd gnd cell_6t
Xbit_r451_c28 bl[28] br[28] wl[451] vdd gnd cell_6t
Xbit_r452_c28 bl[28] br[28] wl[452] vdd gnd cell_6t
Xbit_r453_c28 bl[28] br[28] wl[453] vdd gnd cell_6t
Xbit_r454_c28 bl[28] br[28] wl[454] vdd gnd cell_6t
Xbit_r455_c28 bl[28] br[28] wl[455] vdd gnd cell_6t
Xbit_r456_c28 bl[28] br[28] wl[456] vdd gnd cell_6t
Xbit_r457_c28 bl[28] br[28] wl[457] vdd gnd cell_6t
Xbit_r458_c28 bl[28] br[28] wl[458] vdd gnd cell_6t
Xbit_r459_c28 bl[28] br[28] wl[459] vdd gnd cell_6t
Xbit_r460_c28 bl[28] br[28] wl[460] vdd gnd cell_6t
Xbit_r461_c28 bl[28] br[28] wl[461] vdd gnd cell_6t
Xbit_r462_c28 bl[28] br[28] wl[462] vdd gnd cell_6t
Xbit_r463_c28 bl[28] br[28] wl[463] vdd gnd cell_6t
Xbit_r464_c28 bl[28] br[28] wl[464] vdd gnd cell_6t
Xbit_r465_c28 bl[28] br[28] wl[465] vdd gnd cell_6t
Xbit_r466_c28 bl[28] br[28] wl[466] vdd gnd cell_6t
Xbit_r467_c28 bl[28] br[28] wl[467] vdd gnd cell_6t
Xbit_r468_c28 bl[28] br[28] wl[468] vdd gnd cell_6t
Xbit_r469_c28 bl[28] br[28] wl[469] vdd gnd cell_6t
Xbit_r470_c28 bl[28] br[28] wl[470] vdd gnd cell_6t
Xbit_r471_c28 bl[28] br[28] wl[471] vdd gnd cell_6t
Xbit_r472_c28 bl[28] br[28] wl[472] vdd gnd cell_6t
Xbit_r473_c28 bl[28] br[28] wl[473] vdd gnd cell_6t
Xbit_r474_c28 bl[28] br[28] wl[474] vdd gnd cell_6t
Xbit_r475_c28 bl[28] br[28] wl[475] vdd gnd cell_6t
Xbit_r476_c28 bl[28] br[28] wl[476] vdd gnd cell_6t
Xbit_r477_c28 bl[28] br[28] wl[477] vdd gnd cell_6t
Xbit_r478_c28 bl[28] br[28] wl[478] vdd gnd cell_6t
Xbit_r479_c28 bl[28] br[28] wl[479] vdd gnd cell_6t
Xbit_r480_c28 bl[28] br[28] wl[480] vdd gnd cell_6t
Xbit_r481_c28 bl[28] br[28] wl[481] vdd gnd cell_6t
Xbit_r482_c28 bl[28] br[28] wl[482] vdd gnd cell_6t
Xbit_r483_c28 bl[28] br[28] wl[483] vdd gnd cell_6t
Xbit_r484_c28 bl[28] br[28] wl[484] vdd gnd cell_6t
Xbit_r485_c28 bl[28] br[28] wl[485] vdd gnd cell_6t
Xbit_r486_c28 bl[28] br[28] wl[486] vdd gnd cell_6t
Xbit_r487_c28 bl[28] br[28] wl[487] vdd gnd cell_6t
Xbit_r488_c28 bl[28] br[28] wl[488] vdd gnd cell_6t
Xbit_r489_c28 bl[28] br[28] wl[489] vdd gnd cell_6t
Xbit_r490_c28 bl[28] br[28] wl[490] vdd gnd cell_6t
Xbit_r491_c28 bl[28] br[28] wl[491] vdd gnd cell_6t
Xbit_r492_c28 bl[28] br[28] wl[492] vdd gnd cell_6t
Xbit_r493_c28 bl[28] br[28] wl[493] vdd gnd cell_6t
Xbit_r494_c28 bl[28] br[28] wl[494] vdd gnd cell_6t
Xbit_r495_c28 bl[28] br[28] wl[495] vdd gnd cell_6t
Xbit_r496_c28 bl[28] br[28] wl[496] vdd gnd cell_6t
Xbit_r497_c28 bl[28] br[28] wl[497] vdd gnd cell_6t
Xbit_r498_c28 bl[28] br[28] wl[498] vdd gnd cell_6t
Xbit_r499_c28 bl[28] br[28] wl[499] vdd gnd cell_6t
Xbit_r500_c28 bl[28] br[28] wl[500] vdd gnd cell_6t
Xbit_r501_c28 bl[28] br[28] wl[501] vdd gnd cell_6t
Xbit_r502_c28 bl[28] br[28] wl[502] vdd gnd cell_6t
Xbit_r503_c28 bl[28] br[28] wl[503] vdd gnd cell_6t
Xbit_r504_c28 bl[28] br[28] wl[504] vdd gnd cell_6t
Xbit_r505_c28 bl[28] br[28] wl[505] vdd gnd cell_6t
Xbit_r506_c28 bl[28] br[28] wl[506] vdd gnd cell_6t
Xbit_r507_c28 bl[28] br[28] wl[507] vdd gnd cell_6t
Xbit_r508_c28 bl[28] br[28] wl[508] vdd gnd cell_6t
Xbit_r509_c28 bl[28] br[28] wl[509] vdd gnd cell_6t
Xbit_r510_c28 bl[28] br[28] wl[510] vdd gnd cell_6t
Xbit_r511_c28 bl[28] br[28] wl[511] vdd gnd cell_6t
Xbit_r0_c29 bl[29] br[29] wl[0] vdd gnd cell_6t
Xbit_r1_c29 bl[29] br[29] wl[1] vdd gnd cell_6t
Xbit_r2_c29 bl[29] br[29] wl[2] vdd gnd cell_6t
Xbit_r3_c29 bl[29] br[29] wl[3] vdd gnd cell_6t
Xbit_r4_c29 bl[29] br[29] wl[4] vdd gnd cell_6t
Xbit_r5_c29 bl[29] br[29] wl[5] vdd gnd cell_6t
Xbit_r6_c29 bl[29] br[29] wl[6] vdd gnd cell_6t
Xbit_r7_c29 bl[29] br[29] wl[7] vdd gnd cell_6t
Xbit_r8_c29 bl[29] br[29] wl[8] vdd gnd cell_6t
Xbit_r9_c29 bl[29] br[29] wl[9] vdd gnd cell_6t
Xbit_r10_c29 bl[29] br[29] wl[10] vdd gnd cell_6t
Xbit_r11_c29 bl[29] br[29] wl[11] vdd gnd cell_6t
Xbit_r12_c29 bl[29] br[29] wl[12] vdd gnd cell_6t
Xbit_r13_c29 bl[29] br[29] wl[13] vdd gnd cell_6t
Xbit_r14_c29 bl[29] br[29] wl[14] vdd gnd cell_6t
Xbit_r15_c29 bl[29] br[29] wl[15] vdd gnd cell_6t
Xbit_r16_c29 bl[29] br[29] wl[16] vdd gnd cell_6t
Xbit_r17_c29 bl[29] br[29] wl[17] vdd gnd cell_6t
Xbit_r18_c29 bl[29] br[29] wl[18] vdd gnd cell_6t
Xbit_r19_c29 bl[29] br[29] wl[19] vdd gnd cell_6t
Xbit_r20_c29 bl[29] br[29] wl[20] vdd gnd cell_6t
Xbit_r21_c29 bl[29] br[29] wl[21] vdd gnd cell_6t
Xbit_r22_c29 bl[29] br[29] wl[22] vdd gnd cell_6t
Xbit_r23_c29 bl[29] br[29] wl[23] vdd gnd cell_6t
Xbit_r24_c29 bl[29] br[29] wl[24] vdd gnd cell_6t
Xbit_r25_c29 bl[29] br[29] wl[25] vdd gnd cell_6t
Xbit_r26_c29 bl[29] br[29] wl[26] vdd gnd cell_6t
Xbit_r27_c29 bl[29] br[29] wl[27] vdd gnd cell_6t
Xbit_r28_c29 bl[29] br[29] wl[28] vdd gnd cell_6t
Xbit_r29_c29 bl[29] br[29] wl[29] vdd gnd cell_6t
Xbit_r30_c29 bl[29] br[29] wl[30] vdd gnd cell_6t
Xbit_r31_c29 bl[29] br[29] wl[31] vdd gnd cell_6t
Xbit_r32_c29 bl[29] br[29] wl[32] vdd gnd cell_6t
Xbit_r33_c29 bl[29] br[29] wl[33] vdd gnd cell_6t
Xbit_r34_c29 bl[29] br[29] wl[34] vdd gnd cell_6t
Xbit_r35_c29 bl[29] br[29] wl[35] vdd gnd cell_6t
Xbit_r36_c29 bl[29] br[29] wl[36] vdd gnd cell_6t
Xbit_r37_c29 bl[29] br[29] wl[37] vdd gnd cell_6t
Xbit_r38_c29 bl[29] br[29] wl[38] vdd gnd cell_6t
Xbit_r39_c29 bl[29] br[29] wl[39] vdd gnd cell_6t
Xbit_r40_c29 bl[29] br[29] wl[40] vdd gnd cell_6t
Xbit_r41_c29 bl[29] br[29] wl[41] vdd gnd cell_6t
Xbit_r42_c29 bl[29] br[29] wl[42] vdd gnd cell_6t
Xbit_r43_c29 bl[29] br[29] wl[43] vdd gnd cell_6t
Xbit_r44_c29 bl[29] br[29] wl[44] vdd gnd cell_6t
Xbit_r45_c29 bl[29] br[29] wl[45] vdd gnd cell_6t
Xbit_r46_c29 bl[29] br[29] wl[46] vdd gnd cell_6t
Xbit_r47_c29 bl[29] br[29] wl[47] vdd gnd cell_6t
Xbit_r48_c29 bl[29] br[29] wl[48] vdd gnd cell_6t
Xbit_r49_c29 bl[29] br[29] wl[49] vdd gnd cell_6t
Xbit_r50_c29 bl[29] br[29] wl[50] vdd gnd cell_6t
Xbit_r51_c29 bl[29] br[29] wl[51] vdd gnd cell_6t
Xbit_r52_c29 bl[29] br[29] wl[52] vdd gnd cell_6t
Xbit_r53_c29 bl[29] br[29] wl[53] vdd gnd cell_6t
Xbit_r54_c29 bl[29] br[29] wl[54] vdd gnd cell_6t
Xbit_r55_c29 bl[29] br[29] wl[55] vdd gnd cell_6t
Xbit_r56_c29 bl[29] br[29] wl[56] vdd gnd cell_6t
Xbit_r57_c29 bl[29] br[29] wl[57] vdd gnd cell_6t
Xbit_r58_c29 bl[29] br[29] wl[58] vdd gnd cell_6t
Xbit_r59_c29 bl[29] br[29] wl[59] vdd gnd cell_6t
Xbit_r60_c29 bl[29] br[29] wl[60] vdd gnd cell_6t
Xbit_r61_c29 bl[29] br[29] wl[61] vdd gnd cell_6t
Xbit_r62_c29 bl[29] br[29] wl[62] vdd gnd cell_6t
Xbit_r63_c29 bl[29] br[29] wl[63] vdd gnd cell_6t
Xbit_r64_c29 bl[29] br[29] wl[64] vdd gnd cell_6t
Xbit_r65_c29 bl[29] br[29] wl[65] vdd gnd cell_6t
Xbit_r66_c29 bl[29] br[29] wl[66] vdd gnd cell_6t
Xbit_r67_c29 bl[29] br[29] wl[67] vdd gnd cell_6t
Xbit_r68_c29 bl[29] br[29] wl[68] vdd gnd cell_6t
Xbit_r69_c29 bl[29] br[29] wl[69] vdd gnd cell_6t
Xbit_r70_c29 bl[29] br[29] wl[70] vdd gnd cell_6t
Xbit_r71_c29 bl[29] br[29] wl[71] vdd gnd cell_6t
Xbit_r72_c29 bl[29] br[29] wl[72] vdd gnd cell_6t
Xbit_r73_c29 bl[29] br[29] wl[73] vdd gnd cell_6t
Xbit_r74_c29 bl[29] br[29] wl[74] vdd gnd cell_6t
Xbit_r75_c29 bl[29] br[29] wl[75] vdd gnd cell_6t
Xbit_r76_c29 bl[29] br[29] wl[76] vdd gnd cell_6t
Xbit_r77_c29 bl[29] br[29] wl[77] vdd gnd cell_6t
Xbit_r78_c29 bl[29] br[29] wl[78] vdd gnd cell_6t
Xbit_r79_c29 bl[29] br[29] wl[79] vdd gnd cell_6t
Xbit_r80_c29 bl[29] br[29] wl[80] vdd gnd cell_6t
Xbit_r81_c29 bl[29] br[29] wl[81] vdd gnd cell_6t
Xbit_r82_c29 bl[29] br[29] wl[82] vdd gnd cell_6t
Xbit_r83_c29 bl[29] br[29] wl[83] vdd gnd cell_6t
Xbit_r84_c29 bl[29] br[29] wl[84] vdd gnd cell_6t
Xbit_r85_c29 bl[29] br[29] wl[85] vdd gnd cell_6t
Xbit_r86_c29 bl[29] br[29] wl[86] vdd gnd cell_6t
Xbit_r87_c29 bl[29] br[29] wl[87] vdd gnd cell_6t
Xbit_r88_c29 bl[29] br[29] wl[88] vdd gnd cell_6t
Xbit_r89_c29 bl[29] br[29] wl[89] vdd gnd cell_6t
Xbit_r90_c29 bl[29] br[29] wl[90] vdd gnd cell_6t
Xbit_r91_c29 bl[29] br[29] wl[91] vdd gnd cell_6t
Xbit_r92_c29 bl[29] br[29] wl[92] vdd gnd cell_6t
Xbit_r93_c29 bl[29] br[29] wl[93] vdd gnd cell_6t
Xbit_r94_c29 bl[29] br[29] wl[94] vdd gnd cell_6t
Xbit_r95_c29 bl[29] br[29] wl[95] vdd gnd cell_6t
Xbit_r96_c29 bl[29] br[29] wl[96] vdd gnd cell_6t
Xbit_r97_c29 bl[29] br[29] wl[97] vdd gnd cell_6t
Xbit_r98_c29 bl[29] br[29] wl[98] vdd gnd cell_6t
Xbit_r99_c29 bl[29] br[29] wl[99] vdd gnd cell_6t
Xbit_r100_c29 bl[29] br[29] wl[100] vdd gnd cell_6t
Xbit_r101_c29 bl[29] br[29] wl[101] vdd gnd cell_6t
Xbit_r102_c29 bl[29] br[29] wl[102] vdd gnd cell_6t
Xbit_r103_c29 bl[29] br[29] wl[103] vdd gnd cell_6t
Xbit_r104_c29 bl[29] br[29] wl[104] vdd gnd cell_6t
Xbit_r105_c29 bl[29] br[29] wl[105] vdd gnd cell_6t
Xbit_r106_c29 bl[29] br[29] wl[106] vdd gnd cell_6t
Xbit_r107_c29 bl[29] br[29] wl[107] vdd gnd cell_6t
Xbit_r108_c29 bl[29] br[29] wl[108] vdd gnd cell_6t
Xbit_r109_c29 bl[29] br[29] wl[109] vdd gnd cell_6t
Xbit_r110_c29 bl[29] br[29] wl[110] vdd gnd cell_6t
Xbit_r111_c29 bl[29] br[29] wl[111] vdd gnd cell_6t
Xbit_r112_c29 bl[29] br[29] wl[112] vdd gnd cell_6t
Xbit_r113_c29 bl[29] br[29] wl[113] vdd gnd cell_6t
Xbit_r114_c29 bl[29] br[29] wl[114] vdd gnd cell_6t
Xbit_r115_c29 bl[29] br[29] wl[115] vdd gnd cell_6t
Xbit_r116_c29 bl[29] br[29] wl[116] vdd gnd cell_6t
Xbit_r117_c29 bl[29] br[29] wl[117] vdd gnd cell_6t
Xbit_r118_c29 bl[29] br[29] wl[118] vdd gnd cell_6t
Xbit_r119_c29 bl[29] br[29] wl[119] vdd gnd cell_6t
Xbit_r120_c29 bl[29] br[29] wl[120] vdd gnd cell_6t
Xbit_r121_c29 bl[29] br[29] wl[121] vdd gnd cell_6t
Xbit_r122_c29 bl[29] br[29] wl[122] vdd gnd cell_6t
Xbit_r123_c29 bl[29] br[29] wl[123] vdd gnd cell_6t
Xbit_r124_c29 bl[29] br[29] wl[124] vdd gnd cell_6t
Xbit_r125_c29 bl[29] br[29] wl[125] vdd gnd cell_6t
Xbit_r126_c29 bl[29] br[29] wl[126] vdd gnd cell_6t
Xbit_r127_c29 bl[29] br[29] wl[127] vdd gnd cell_6t
Xbit_r128_c29 bl[29] br[29] wl[128] vdd gnd cell_6t
Xbit_r129_c29 bl[29] br[29] wl[129] vdd gnd cell_6t
Xbit_r130_c29 bl[29] br[29] wl[130] vdd gnd cell_6t
Xbit_r131_c29 bl[29] br[29] wl[131] vdd gnd cell_6t
Xbit_r132_c29 bl[29] br[29] wl[132] vdd gnd cell_6t
Xbit_r133_c29 bl[29] br[29] wl[133] vdd gnd cell_6t
Xbit_r134_c29 bl[29] br[29] wl[134] vdd gnd cell_6t
Xbit_r135_c29 bl[29] br[29] wl[135] vdd gnd cell_6t
Xbit_r136_c29 bl[29] br[29] wl[136] vdd gnd cell_6t
Xbit_r137_c29 bl[29] br[29] wl[137] vdd gnd cell_6t
Xbit_r138_c29 bl[29] br[29] wl[138] vdd gnd cell_6t
Xbit_r139_c29 bl[29] br[29] wl[139] vdd gnd cell_6t
Xbit_r140_c29 bl[29] br[29] wl[140] vdd gnd cell_6t
Xbit_r141_c29 bl[29] br[29] wl[141] vdd gnd cell_6t
Xbit_r142_c29 bl[29] br[29] wl[142] vdd gnd cell_6t
Xbit_r143_c29 bl[29] br[29] wl[143] vdd gnd cell_6t
Xbit_r144_c29 bl[29] br[29] wl[144] vdd gnd cell_6t
Xbit_r145_c29 bl[29] br[29] wl[145] vdd gnd cell_6t
Xbit_r146_c29 bl[29] br[29] wl[146] vdd gnd cell_6t
Xbit_r147_c29 bl[29] br[29] wl[147] vdd gnd cell_6t
Xbit_r148_c29 bl[29] br[29] wl[148] vdd gnd cell_6t
Xbit_r149_c29 bl[29] br[29] wl[149] vdd gnd cell_6t
Xbit_r150_c29 bl[29] br[29] wl[150] vdd gnd cell_6t
Xbit_r151_c29 bl[29] br[29] wl[151] vdd gnd cell_6t
Xbit_r152_c29 bl[29] br[29] wl[152] vdd gnd cell_6t
Xbit_r153_c29 bl[29] br[29] wl[153] vdd gnd cell_6t
Xbit_r154_c29 bl[29] br[29] wl[154] vdd gnd cell_6t
Xbit_r155_c29 bl[29] br[29] wl[155] vdd gnd cell_6t
Xbit_r156_c29 bl[29] br[29] wl[156] vdd gnd cell_6t
Xbit_r157_c29 bl[29] br[29] wl[157] vdd gnd cell_6t
Xbit_r158_c29 bl[29] br[29] wl[158] vdd gnd cell_6t
Xbit_r159_c29 bl[29] br[29] wl[159] vdd gnd cell_6t
Xbit_r160_c29 bl[29] br[29] wl[160] vdd gnd cell_6t
Xbit_r161_c29 bl[29] br[29] wl[161] vdd gnd cell_6t
Xbit_r162_c29 bl[29] br[29] wl[162] vdd gnd cell_6t
Xbit_r163_c29 bl[29] br[29] wl[163] vdd gnd cell_6t
Xbit_r164_c29 bl[29] br[29] wl[164] vdd gnd cell_6t
Xbit_r165_c29 bl[29] br[29] wl[165] vdd gnd cell_6t
Xbit_r166_c29 bl[29] br[29] wl[166] vdd gnd cell_6t
Xbit_r167_c29 bl[29] br[29] wl[167] vdd gnd cell_6t
Xbit_r168_c29 bl[29] br[29] wl[168] vdd gnd cell_6t
Xbit_r169_c29 bl[29] br[29] wl[169] vdd gnd cell_6t
Xbit_r170_c29 bl[29] br[29] wl[170] vdd gnd cell_6t
Xbit_r171_c29 bl[29] br[29] wl[171] vdd gnd cell_6t
Xbit_r172_c29 bl[29] br[29] wl[172] vdd gnd cell_6t
Xbit_r173_c29 bl[29] br[29] wl[173] vdd gnd cell_6t
Xbit_r174_c29 bl[29] br[29] wl[174] vdd gnd cell_6t
Xbit_r175_c29 bl[29] br[29] wl[175] vdd gnd cell_6t
Xbit_r176_c29 bl[29] br[29] wl[176] vdd gnd cell_6t
Xbit_r177_c29 bl[29] br[29] wl[177] vdd gnd cell_6t
Xbit_r178_c29 bl[29] br[29] wl[178] vdd gnd cell_6t
Xbit_r179_c29 bl[29] br[29] wl[179] vdd gnd cell_6t
Xbit_r180_c29 bl[29] br[29] wl[180] vdd gnd cell_6t
Xbit_r181_c29 bl[29] br[29] wl[181] vdd gnd cell_6t
Xbit_r182_c29 bl[29] br[29] wl[182] vdd gnd cell_6t
Xbit_r183_c29 bl[29] br[29] wl[183] vdd gnd cell_6t
Xbit_r184_c29 bl[29] br[29] wl[184] vdd gnd cell_6t
Xbit_r185_c29 bl[29] br[29] wl[185] vdd gnd cell_6t
Xbit_r186_c29 bl[29] br[29] wl[186] vdd gnd cell_6t
Xbit_r187_c29 bl[29] br[29] wl[187] vdd gnd cell_6t
Xbit_r188_c29 bl[29] br[29] wl[188] vdd gnd cell_6t
Xbit_r189_c29 bl[29] br[29] wl[189] vdd gnd cell_6t
Xbit_r190_c29 bl[29] br[29] wl[190] vdd gnd cell_6t
Xbit_r191_c29 bl[29] br[29] wl[191] vdd gnd cell_6t
Xbit_r192_c29 bl[29] br[29] wl[192] vdd gnd cell_6t
Xbit_r193_c29 bl[29] br[29] wl[193] vdd gnd cell_6t
Xbit_r194_c29 bl[29] br[29] wl[194] vdd gnd cell_6t
Xbit_r195_c29 bl[29] br[29] wl[195] vdd gnd cell_6t
Xbit_r196_c29 bl[29] br[29] wl[196] vdd gnd cell_6t
Xbit_r197_c29 bl[29] br[29] wl[197] vdd gnd cell_6t
Xbit_r198_c29 bl[29] br[29] wl[198] vdd gnd cell_6t
Xbit_r199_c29 bl[29] br[29] wl[199] vdd gnd cell_6t
Xbit_r200_c29 bl[29] br[29] wl[200] vdd gnd cell_6t
Xbit_r201_c29 bl[29] br[29] wl[201] vdd gnd cell_6t
Xbit_r202_c29 bl[29] br[29] wl[202] vdd gnd cell_6t
Xbit_r203_c29 bl[29] br[29] wl[203] vdd gnd cell_6t
Xbit_r204_c29 bl[29] br[29] wl[204] vdd gnd cell_6t
Xbit_r205_c29 bl[29] br[29] wl[205] vdd gnd cell_6t
Xbit_r206_c29 bl[29] br[29] wl[206] vdd gnd cell_6t
Xbit_r207_c29 bl[29] br[29] wl[207] vdd gnd cell_6t
Xbit_r208_c29 bl[29] br[29] wl[208] vdd gnd cell_6t
Xbit_r209_c29 bl[29] br[29] wl[209] vdd gnd cell_6t
Xbit_r210_c29 bl[29] br[29] wl[210] vdd gnd cell_6t
Xbit_r211_c29 bl[29] br[29] wl[211] vdd gnd cell_6t
Xbit_r212_c29 bl[29] br[29] wl[212] vdd gnd cell_6t
Xbit_r213_c29 bl[29] br[29] wl[213] vdd gnd cell_6t
Xbit_r214_c29 bl[29] br[29] wl[214] vdd gnd cell_6t
Xbit_r215_c29 bl[29] br[29] wl[215] vdd gnd cell_6t
Xbit_r216_c29 bl[29] br[29] wl[216] vdd gnd cell_6t
Xbit_r217_c29 bl[29] br[29] wl[217] vdd gnd cell_6t
Xbit_r218_c29 bl[29] br[29] wl[218] vdd gnd cell_6t
Xbit_r219_c29 bl[29] br[29] wl[219] vdd gnd cell_6t
Xbit_r220_c29 bl[29] br[29] wl[220] vdd gnd cell_6t
Xbit_r221_c29 bl[29] br[29] wl[221] vdd gnd cell_6t
Xbit_r222_c29 bl[29] br[29] wl[222] vdd gnd cell_6t
Xbit_r223_c29 bl[29] br[29] wl[223] vdd gnd cell_6t
Xbit_r224_c29 bl[29] br[29] wl[224] vdd gnd cell_6t
Xbit_r225_c29 bl[29] br[29] wl[225] vdd gnd cell_6t
Xbit_r226_c29 bl[29] br[29] wl[226] vdd gnd cell_6t
Xbit_r227_c29 bl[29] br[29] wl[227] vdd gnd cell_6t
Xbit_r228_c29 bl[29] br[29] wl[228] vdd gnd cell_6t
Xbit_r229_c29 bl[29] br[29] wl[229] vdd gnd cell_6t
Xbit_r230_c29 bl[29] br[29] wl[230] vdd gnd cell_6t
Xbit_r231_c29 bl[29] br[29] wl[231] vdd gnd cell_6t
Xbit_r232_c29 bl[29] br[29] wl[232] vdd gnd cell_6t
Xbit_r233_c29 bl[29] br[29] wl[233] vdd gnd cell_6t
Xbit_r234_c29 bl[29] br[29] wl[234] vdd gnd cell_6t
Xbit_r235_c29 bl[29] br[29] wl[235] vdd gnd cell_6t
Xbit_r236_c29 bl[29] br[29] wl[236] vdd gnd cell_6t
Xbit_r237_c29 bl[29] br[29] wl[237] vdd gnd cell_6t
Xbit_r238_c29 bl[29] br[29] wl[238] vdd gnd cell_6t
Xbit_r239_c29 bl[29] br[29] wl[239] vdd gnd cell_6t
Xbit_r240_c29 bl[29] br[29] wl[240] vdd gnd cell_6t
Xbit_r241_c29 bl[29] br[29] wl[241] vdd gnd cell_6t
Xbit_r242_c29 bl[29] br[29] wl[242] vdd gnd cell_6t
Xbit_r243_c29 bl[29] br[29] wl[243] vdd gnd cell_6t
Xbit_r244_c29 bl[29] br[29] wl[244] vdd gnd cell_6t
Xbit_r245_c29 bl[29] br[29] wl[245] vdd gnd cell_6t
Xbit_r246_c29 bl[29] br[29] wl[246] vdd gnd cell_6t
Xbit_r247_c29 bl[29] br[29] wl[247] vdd gnd cell_6t
Xbit_r248_c29 bl[29] br[29] wl[248] vdd gnd cell_6t
Xbit_r249_c29 bl[29] br[29] wl[249] vdd gnd cell_6t
Xbit_r250_c29 bl[29] br[29] wl[250] vdd gnd cell_6t
Xbit_r251_c29 bl[29] br[29] wl[251] vdd gnd cell_6t
Xbit_r252_c29 bl[29] br[29] wl[252] vdd gnd cell_6t
Xbit_r253_c29 bl[29] br[29] wl[253] vdd gnd cell_6t
Xbit_r254_c29 bl[29] br[29] wl[254] vdd gnd cell_6t
Xbit_r255_c29 bl[29] br[29] wl[255] vdd gnd cell_6t
Xbit_r256_c29 bl[29] br[29] wl[256] vdd gnd cell_6t
Xbit_r257_c29 bl[29] br[29] wl[257] vdd gnd cell_6t
Xbit_r258_c29 bl[29] br[29] wl[258] vdd gnd cell_6t
Xbit_r259_c29 bl[29] br[29] wl[259] vdd gnd cell_6t
Xbit_r260_c29 bl[29] br[29] wl[260] vdd gnd cell_6t
Xbit_r261_c29 bl[29] br[29] wl[261] vdd gnd cell_6t
Xbit_r262_c29 bl[29] br[29] wl[262] vdd gnd cell_6t
Xbit_r263_c29 bl[29] br[29] wl[263] vdd gnd cell_6t
Xbit_r264_c29 bl[29] br[29] wl[264] vdd gnd cell_6t
Xbit_r265_c29 bl[29] br[29] wl[265] vdd gnd cell_6t
Xbit_r266_c29 bl[29] br[29] wl[266] vdd gnd cell_6t
Xbit_r267_c29 bl[29] br[29] wl[267] vdd gnd cell_6t
Xbit_r268_c29 bl[29] br[29] wl[268] vdd gnd cell_6t
Xbit_r269_c29 bl[29] br[29] wl[269] vdd gnd cell_6t
Xbit_r270_c29 bl[29] br[29] wl[270] vdd gnd cell_6t
Xbit_r271_c29 bl[29] br[29] wl[271] vdd gnd cell_6t
Xbit_r272_c29 bl[29] br[29] wl[272] vdd gnd cell_6t
Xbit_r273_c29 bl[29] br[29] wl[273] vdd gnd cell_6t
Xbit_r274_c29 bl[29] br[29] wl[274] vdd gnd cell_6t
Xbit_r275_c29 bl[29] br[29] wl[275] vdd gnd cell_6t
Xbit_r276_c29 bl[29] br[29] wl[276] vdd gnd cell_6t
Xbit_r277_c29 bl[29] br[29] wl[277] vdd gnd cell_6t
Xbit_r278_c29 bl[29] br[29] wl[278] vdd gnd cell_6t
Xbit_r279_c29 bl[29] br[29] wl[279] vdd gnd cell_6t
Xbit_r280_c29 bl[29] br[29] wl[280] vdd gnd cell_6t
Xbit_r281_c29 bl[29] br[29] wl[281] vdd gnd cell_6t
Xbit_r282_c29 bl[29] br[29] wl[282] vdd gnd cell_6t
Xbit_r283_c29 bl[29] br[29] wl[283] vdd gnd cell_6t
Xbit_r284_c29 bl[29] br[29] wl[284] vdd gnd cell_6t
Xbit_r285_c29 bl[29] br[29] wl[285] vdd gnd cell_6t
Xbit_r286_c29 bl[29] br[29] wl[286] vdd gnd cell_6t
Xbit_r287_c29 bl[29] br[29] wl[287] vdd gnd cell_6t
Xbit_r288_c29 bl[29] br[29] wl[288] vdd gnd cell_6t
Xbit_r289_c29 bl[29] br[29] wl[289] vdd gnd cell_6t
Xbit_r290_c29 bl[29] br[29] wl[290] vdd gnd cell_6t
Xbit_r291_c29 bl[29] br[29] wl[291] vdd gnd cell_6t
Xbit_r292_c29 bl[29] br[29] wl[292] vdd gnd cell_6t
Xbit_r293_c29 bl[29] br[29] wl[293] vdd gnd cell_6t
Xbit_r294_c29 bl[29] br[29] wl[294] vdd gnd cell_6t
Xbit_r295_c29 bl[29] br[29] wl[295] vdd gnd cell_6t
Xbit_r296_c29 bl[29] br[29] wl[296] vdd gnd cell_6t
Xbit_r297_c29 bl[29] br[29] wl[297] vdd gnd cell_6t
Xbit_r298_c29 bl[29] br[29] wl[298] vdd gnd cell_6t
Xbit_r299_c29 bl[29] br[29] wl[299] vdd gnd cell_6t
Xbit_r300_c29 bl[29] br[29] wl[300] vdd gnd cell_6t
Xbit_r301_c29 bl[29] br[29] wl[301] vdd gnd cell_6t
Xbit_r302_c29 bl[29] br[29] wl[302] vdd gnd cell_6t
Xbit_r303_c29 bl[29] br[29] wl[303] vdd gnd cell_6t
Xbit_r304_c29 bl[29] br[29] wl[304] vdd gnd cell_6t
Xbit_r305_c29 bl[29] br[29] wl[305] vdd gnd cell_6t
Xbit_r306_c29 bl[29] br[29] wl[306] vdd gnd cell_6t
Xbit_r307_c29 bl[29] br[29] wl[307] vdd gnd cell_6t
Xbit_r308_c29 bl[29] br[29] wl[308] vdd gnd cell_6t
Xbit_r309_c29 bl[29] br[29] wl[309] vdd gnd cell_6t
Xbit_r310_c29 bl[29] br[29] wl[310] vdd gnd cell_6t
Xbit_r311_c29 bl[29] br[29] wl[311] vdd gnd cell_6t
Xbit_r312_c29 bl[29] br[29] wl[312] vdd gnd cell_6t
Xbit_r313_c29 bl[29] br[29] wl[313] vdd gnd cell_6t
Xbit_r314_c29 bl[29] br[29] wl[314] vdd gnd cell_6t
Xbit_r315_c29 bl[29] br[29] wl[315] vdd gnd cell_6t
Xbit_r316_c29 bl[29] br[29] wl[316] vdd gnd cell_6t
Xbit_r317_c29 bl[29] br[29] wl[317] vdd gnd cell_6t
Xbit_r318_c29 bl[29] br[29] wl[318] vdd gnd cell_6t
Xbit_r319_c29 bl[29] br[29] wl[319] vdd gnd cell_6t
Xbit_r320_c29 bl[29] br[29] wl[320] vdd gnd cell_6t
Xbit_r321_c29 bl[29] br[29] wl[321] vdd gnd cell_6t
Xbit_r322_c29 bl[29] br[29] wl[322] vdd gnd cell_6t
Xbit_r323_c29 bl[29] br[29] wl[323] vdd gnd cell_6t
Xbit_r324_c29 bl[29] br[29] wl[324] vdd gnd cell_6t
Xbit_r325_c29 bl[29] br[29] wl[325] vdd gnd cell_6t
Xbit_r326_c29 bl[29] br[29] wl[326] vdd gnd cell_6t
Xbit_r327_c29 bl[29] br[29] wl[327] vdd gnd cell_6t
Xbit_r328_c29 bl[29] br[29] wl[328] vdd gnd cell_6t
Xbit_r329_c29 bl[29] br[29] wl[329] vdd gnd cell_6t
Xbit_r330_c29 bl[29] br[29] wl[330] vdd gnd cell_6t
Xbit_r331_c29 bl[29] br[29] wl[331] vdd gnd cell_6t
Xbit_r332_c29 bl[29] br[29] wl[332] vdd gnd cell_6t
Xbit_r333_c29 bl[29] br[29] wl[333] vdd gnd cell_6t
Xbit_r334_c29 bl[29] br[29] wl[334] vdd gnd cell_6t
Xbit_r335_c29 bl[29] br[29] wl[335] vdd gnd cell_6t
Xbit_r336_c29 bl[29] br[29] wl[336] vdd gnd cell_6t
Xbit_r337_c29 bl[29] br[29] wl[337] vdd gnd cell_6t
Xbit_r338_c29 bl[29] br[29] wl[338] vdd gnd cell_6t
Xbit_r339_c29 bl[29] br[29] wl[339] vdd gnd cell_6t
Xbit_r340_c29 bl[29] br[29] wl[340] vdd gnd cell_6t
Xbit_r341_c29 bl[29] br[29] wl[341] vdd gnd cell_6t
Xbit_r342_c29 bl[29] br[29] wl[342] vdd gnd cell_6t
Xbit_r343_c29 bl[29] br[29] wl[343] vdd gnd cell_6t
Xbit_r344_c29 bl[29] br[29] wl[344] vdd gnd cell_6t
Xbit_r345_c29 bl[29] br[29] wl[345] vdd gnd cell_6t
Xbit_r346_c29 bl[29] br[29] wl[346] vdd gnd cell_6t
Xbit_r347_c29 bl[29] br[29] wl[347] vdd gnd cell_6t
Xbit_r348_c29 bl[29] br[29] wl[348] vdd gnd cell_6t
Xbit_r349_c29 bl[29] br[29] wl[349] vdd gnd cell_6t
Xbit_r350_c29 bl[29] br[29] wl[350] vdd gnd cell_6t
Xbit_r351_c29 bl[29] br[29] wl[351] vdd gnd cell_6t
Xbit_r352_c29 bl[29] br[29] wl[352] vdd gnd cell_6t
Xbit_r353_c29 bl[29] br[29] wl[353] vdd gnd cell_6t
Xbit_r354_c29 bl[29] br[29] wl[354] vdd gnd cell_6t
Xbit_r355_c29 bl[29] br[29] wl[355] vdd gnd cell_6t
Xbit_r356_c29 bl[29] br[29] wl[356] vdd gnd cell_6t
Xbit_r357_c29 bl[29] br[29] wl[357] vdd gnd cell_6t
Xbit_r358_c29 bl[29] br[29] wl[358] vdd gnd cell_6t
Xbit_r359_c29 bl[29] br[29] wl[359] vdd gnd cell_6t
Xbit_r360_c29 bl[29] br[29] wl[360] vdd gnd cell_6t
Xbit_r361_c29 bl[29] br[29] wl[361] vdd gnd cell_6t
Xbit_r362_c29 bl[29] br[29] wl[362] vdd gnd cell_6t
Xbit_r363_c29 bl[29] br[29] wl[363] vdd gnd cell_6t
Xbit_r364_c29 bl[29] br[29] wl[364] vdd gnd cell_6t
Xbit_r365_c29 bl[29] br[29] wl[365] vdd gnd cell_6t
Xbit_r366_c29 bl[29] br[29] wl[366] vdd gnd cell_6t
Xbit_r367_c29 bl[29] br[29] wl[367] vdd gnd cell_6t
Xbit_r368_c29 bl[29] br[29] wl[368] vdd gnd cell_6t
Xbit_r369_c29 bl[29] br[29] wl[369] vdd gnd cell_6t
Xbit_r370_c29 bl[29] br[29] wl[370] vdd gnd cell_6t
Xbit_r371_c29 bl[29] br[29] wl[371] vdd gnd cell_6t
Xbit_r372_c29 bl[29] br[29] wl[372] vdd gnd cell_6t
Xbit_r373_c29 bl[29] br[29] wl[373] vdd gnd cell_6t
Xbit_r374_c29 bl[29] br[29] wl[374] vdd gnd cell_6t
Xbit_r375_c29 bl[29] br[29] wl[375] vdd gnd cell_6t
Xbit_r376_c29 bl[29] br[29] wl[376] vdd gnd cell_6t
Xbit_r377_c29 bl[29] br[29] wl[377] vdd gnd cell_6t
Xbit_r378_c29 bl[29] br[29] wl[378] vdd gnd cell_6t
Xbit_r379_c29 bl[29] br[29] wl[379] vdd gnd cell_6t
Xbit_r380_c29 bl[29] br[29] wl[380] vdd gnd cell_6t
Xbit_r381_c29 bl[29] br[29] wl[381] vdd gnd cell_6t
Xbit_r382_c29 bl[29] br[29] wl[382] vdd gnd cell_6t
Xbit_r383_c29 bl[29] br[29] wl[383] vdd gnd cell_6t
Xbit_r384_c29 bl[29] br[29] wl[384] vdd gnd cell_6t
Xbit_r385_c29 bl[29] br[29] wl[385] vdd gnd cell_6t
Xbit_r386_c29 bl[29] br[29] wl[386] vdd gnd cell_6t
Xbit_r387_c29 bl[29] br[29] wl[387] vdd gnd cell_6t
Xbit_r388_c29 bl[29] br[29] wl[388] vdd gnd cell_6t
Xbit_r389_c29 bl[29] br[29] wl[389] vdd gnd cell_6t
Xbit_r390_c29 bl[29] br[29] wl[390] vdd gnd cell_6t
Xbit_r391_c29 bl[29] br[29] wl[391] vdd gnd cell_6t
Xbit_r392_c29 bl[29] br[29] wl[392] vdd gnd cell_6t
Xbit_r393_c29 bl[29] br[29] wl[393] vdd gnd cell_6t
Xbit_r394_c29 bl[29] br[29] wl[394] vdd gnd cell_6t
Xbit_r395_c29 bl[29] br[29] wl[395] vdd gnd cell_6t
Xbit_r396_c29 bl[29] br[29] wl[396] vdd gnd cell_6t
Xbit_r397_c29 bl[29] br[29] wl[397] vdd gnd cell_6t
Xbit_r398_c29 bl[29] br[29] wl[398] vdd gnd cell_6t
Xbit_r399_c29 bl[29] br[29] wl[399] vdd gnd cell_6t
Xbit_r400_c29 bl[29] br[29] wl[400] vdd gnd cell_6t
Xbit_r401_c29 bl[29] br[29] wl[401] vdd gnd cell_6t
Xbit_r402_c29 bl[29] br[29] wl[402] vdd gnd cell_6t
Xbit_r403_c29 bl[29] br[29] wl[403] vdd gnd cell_6t
Xbit_r404_c29 bl[29] br[29] wl[404] vdd gnd cell_6t
Xbit_r405_c29 bl[29] br[29] wl[405] vdd gnd cell_6t
Xbit_r406_c29 bl[29] br[29] wl[406] vdd gnd cell_6t
Xbit_r407_c29 bl[29] br[29] wl[407] vdd gnd cell_6t
Xbit_r408_c29 bl[29] br[29] wl[408] vdd gnd cell_6t
Xbit_r409_c29 bl[29] br[29] wl[409] vdd gnd cell_6t
Xbit_r410_c29 bl[29] br[29] wl[410] vdd gnd cell_6t
Xbit_r411_c29 bl[29] br[29] wl[411] vdd gnd cell_6t
Xbit_r412_c29 bl[29] br[29] wl[412] vdd gnd cell_6t
Xbit_r413_c29 bl[29] br[29] wl[413] vdd gnd cell_6t
Xbit_r414_c29 bl[29] br[29] wl[414] vdd gnd cell_6t
Xbit_r415_c29 bl[29] br[29] wl[415] vdd gnd cell_6t
Xbit_r416_c29 bl[29] br[29] wl[416] vdd gnd cell_6t
Xbit_r417_c29 bl[29] br[29] wl[417] vdd gnd cell_6t
Xbit_r418_c29 bl[29] br[29] wl[418] vdd gnd cell_6t
Xbit_r419_c29 bl[29] br[29] wl[419] vdd gnd cell_6t
Xbit_r420_c29 bl[29] br[29] wl[420] vdd gnd cell_6t
Xbit_r421_c29 bl[29] br[29] wl[421] vdd gnd cell_6t
Xbit_r422_c29 bl[29] br[29] wl[422] vdd gnd cell_6t
Xbit_r423_c29 bl[29] br[29] wl[423] vdd gnd cell_6t
Xbit_r424_c29 bl[29] br[29] wl[424] vdd gnd cell_6t
Xbit_r425_c29 bl[29] br[29] wl[425] vdd gnd cell_6t
Xbit_r426_c29 bl[29] br[29] wl[426] vdd gnd cell_6t
Xbit_r427_c29 bl[29] br[29] wl[427] vdd gnd cell_6t
Xbit_r428_c29 bl[29] br[29] wl[428] vdd gnd cell_6t
Xbit_r429_c29 bl[29] br[29] wl[429] vdd gnd cell_6t
Xbit_r430_c29 bl[29] br[29] wl[430] vdd gnd cell_6t
Xbit_r431_c29 bl[29] br[29] wl[431] vdd gnd cell_6t
Xbit_r432_c29 bl[29] br[29] wl[432] vdd gnd cell_6t
Xbit_r433_c29 bl[29] br[29] wl[433] vdd gnd cell_6t
Xbit_r434_c29 bl[29] br[29] wl[434] vdd gnd cell_6t
Xbit_r435_c29 bl[29] br[29] wl[435] vdd gnd cell_6t
Xbit_r436_c29 bl[29] br[29] wl[436] vdd gnd cell_6t
Xbit_r437_c29 bl[29] br[29] wl[437] vdd gnd cell_6t
Xbit_r438_c29 bl[29] br[29] wl[438] vdd gnd cell_6t
Xbit_r439_c29 bl[29] br[29] wl[439] vdd gnd cell_6t
Xbit_r440_c29 bl[29] br[29] wl[440] vdd gnd cell_6t
Xbit_r441_c29 bl[29] br[29] wl[441] vdd gnd cell_6t
Xbit_r442_c29 bl[29] br[29] wl[442] vdd gnd cell_6t
Xbit_r443_c29 bl[29] br[29] wl[443] vdd gnd cell_6t
Xbit_r444_c29 bl[29] br[29] wl[444] vdd gnd cell_6t
Xbit_r445_c29 bl[29] br[29] wl[445] vdd gnd cell_6t
Xbit_r446_c29 bl[29] br[29] wl[446] vdd gnd cell_6t
Xbit_r447_c29 bl[29] br[29] wl[447] vdd gnd cell_6t
Xbit_r448_c29 bl[29] br[29] wl[448] vdd gnd cell_6t
Xbit_r449_c29 bl[29] br[29] wl[449] vdd gnd cell_6t
Xbit_r450_c29 bl[29] br[29] wl[450] vdd gnd cell_6t
Xbit_r451_c29 bl[29] br[29] wl[451] vdd gnd cell_6t
Xbit_r452_c29 bl[29] br[29] wl[452] vdd gnd cell_6t
Xbit_r453_c29 bl[29] br[29] wl[453] vdd gnd cell_6t
Xbit_r454_c29 bl[29] br[29] wl[454] vdd gnd cell_6t
Xbit_r455_c29 bl[29] br[29] wl[455] vdd gnd cell_6t
Xbit_r456_c29 bl[29] br[29] wl[456] vdd gnd cell_6t
Xbit_r457_c29 bl[29] br[29] wl[457] vdd gnd cell_6t
Xbit_r458_c29 bl[29] br[29] wl[458] vdd gnd cell_6t
Xbit_r459_c29 bl[29] br[29] wl[459] vdd gnd cell_6t
Xbit_r460_c29 bl[29] br[29] wl[460] vdd gnd cell_6t
Xbit_r461_c29 bl[29] br[29] wl[461] vdd gnd cell_6t
Xbit_r462_c29 bl[29] br[29] wl[462] vdd gnd cell_6t
Xbit_r463_c29 bl[29] br[29] wl[463] vdd gnd cell_6t
Xbit_r464_c29 bl[29] br[29] wl[464] vdd gnd cell_6t
Xbit_r465_c29 bl[29] br[29] wl[465] vdd gnd cell_6t
Xbit_r466_c29 bl[29] br[29] wl[466] vdd gnd cell_6t
Xbit_r467_c29 bl[29] br[29] wl[467] vdd gnd cell_6t
Xbit_r468_c29 bl[29] br[29] wl[468] vdd gnd cell_6t
Xbit_r469_c29 bl[29] br[29] wl[469] vdd gnd cell_6t
Xbit_r470_c29 bl[29] br[29] wl[470] vdd gnd cell_6t
Xbit_r471_c29 bl[29] br[29] wl[471] vdd gnd cell_6t
Xbit_r472_c29 bl[29] br[29] wl[472] vdd gnd cell_6t
Xbit_r473_c29 bl[29] br[29] wl[473] vdd gnd cell_6t
Xbit_r474_c29 bl[29] br[29] wl[474] vdd gnd cell_6t
Xbit_r475_c29 bl[29] br[29] wl[475] vdd gnd cell_6t
Xbit_r476_c29 bl[29] br[29] wl[476] vdd gnd cell_6t
Xbit_r477_c29 bl[29] br[29] wl[477] vdd gnd cell_6t
Xbit_r478_c29 bl[29] br[29] wl[478] vdd gnd cell_6t
Xbit_r479_c29 bl[29] br[29] wl[479] vdd gnd cell_6t
Xbit_r480_c29 bl[29] br[29] wl[480] vdd gnd cell_6t
Xbit_r481_c29 bl[29] br[29] wl[481] vdd gnd cell_6t
Xbit_r482_c29 bl[29] br[29] wl[482] vdd gnd cell_6t
Xbit_r483_c29 bl[29] br[29] wl[483] vdd gnd cell_6t
Xbit_r484_c29 bl[29] br[29] wl[484] vdd gnd cell_6t
Xbit_r485_c29 bl[29] br[29] wl[485] vdd gnd cell_6t
Xbit_r486_c29 bl[29] br[29] wl[486] vdd gnd cell_6t
Xbit_r487_c29 bl[29] br[29] wl[487] vdd gnd cell_6t
Xbit_r488_c29 bl[29] br[29] wl[488] vdd gnd cell_6t
Xbit_r489_c29 bl[29] br[29] wl[489] vdd gnd cell_6t
Xbit_r490_c29 bl[29] br[29] wl[490] vdd gnd cell_6t
Xbit_r491_c29 bl[29] br[29] wl[491] vdd gnd cell_6t
Xbit_r492_c29 bl[29] br[29] wl[492] vdd gnd cell_6t
Xbit_r493_c29 bl[29] br[29] wl[493] vdd gnd cell_6t
Xbit_r494_c29 bl[29] br[29] wl[494] vdd gnd cell_6t
Xbit_r495_c29 bl[29] br[29] wl[495] vdd gnd cell_6t
Xbit_r496_c29 bl[29] br[29] wl[496] vdd gnd cell_6t
Xbit_r497_c29 bl[29] br[29] wl[497] vdd gnd cell_6t
Xbit_r498_c29 bl[29] br[29] wl[498] vdd gnd cell_6t
Xbit_r499_c29 bl[29] br[29] wl[499] vdd gnd cell_6t
Xbit_r500_c29 bl[29] br[29] wl[500] vdd gnd cell_6t
Xbit_r501_c29 bl[29] br[29] wl[501] vdd gnd cell_6t
Xbit_r502_c29 bl[29] br[29] wl[502] vdd gnd cell_6t
Xbit_r503_c29 bl[29] br[29] wl[503] vdd gnd cell_6t
Xbit_r504_c29 bl[29] br[29] wl[504] vdd gnd cell_6t
Xbit_r505_c29 bl[29] br[29] wl[505] vdd gnd cell_6t
Xbit_r506_c29 bl[29] br[29] wl[506] vdd gnd cell_6t
Xbit_r507_c29 bl[29] br[29] wl[507] vdd gnd cell_6t
Xbit_r508_c29 bl[29] br[29] wl[508] vdd gnd cell_6t
Xbit_r509_c29 bl[29] br[29] wl[509] vdd gnd cell_6t
Xbit_r510_c29 bl[29] br[29] wl[510] vdd gnd cell_6t
Xbit_r511_c29 bl[29] br[29] wl[511] vdd gnd cell_6t
Xbit_r0_c30 bl[30] br[30] wl[0] vdd gnd cell_6t
Xbit_r1_c30 bl[30] br[30] wl[1] vdd gnd cell_6t
Xbit_r2_c30 bl[30] br[30] wl[2] vdd gnd cell_6t
Xbit_r3_c30 bl[30] br[30] wl[3] vdd gnd cell_6t
Xbit_r4_c30 bl[30] br[30] wl[4] vdd gnd cell_6t
Xbit_r5_c30 bl[30] br[30] wl[5] vdd gnd cell_6t
Xbit_r6_c30 bl[30] br[30] wl[6] vdd gnd cell_6t
Xbit_r7_c30 bl[30] br[30] wl[7] vdd gnd cell_6t
Xbit_r8_c30 bl[30] br[30] wl[8] vdd gnd cell_6t
Xbit_r9_c30 bl[30] br[30] wl[9] vdd gnd cell_6t
Xbit_r10_c30 bl[30] br[30] wl[10] vdd gnd cell_6t
Xbit_r11_c30 bl[30] br[30] wl[11] vdd gnd cell_6t
Xbit_r12_c30 bl[30] br[30] wl[12] vdd gnd cell_6t
Xbit_r13_c30 bl[30] br[30] wl[13] vdd gnd cell_6t
Xbit_r14_c30 bl[30] br[30] wl[14] vdd gnd cell_6t
Xbit_r15_c30 bl[30] br[30] wl[15] vdd gnd cell_6t
Xbit_r16_c30 bl[30] br[30] wl[16] vdd gnd cell_6t
Xbit_r17_c30 bl[30] br[30] wl[17] vdd gnd cell_6t
Xbit_r18_c30 bl[30] br[30] wl[18] vdd gnd cell_6t
Xbit_r19_c30 bl[30] br[30] wl[19] vdd gnd cell_6t
Xbit_r20_c30 bl[30] br[30] wl[20] vdd gnd cell_6t
Xbit_r21_c30 bl[30] br[30] wl[21] vdd gnd cell_6t
Xbit_r22_c30 bl[30] br[30] wl[22] vdd gnd cell_6t
Xbit_r23_c30 bl[30] br[30] wl[23] vdd gnd cell_6t
Xbit_r24_c30 bl[30] br[30] wl[24] vdd gnd cell_6t
Xbit_r25_c30 bl[30] br[30] wl[25] vdd gnd cell_6t
Xbit_r26_c30 bl[30] br[30] wl[26] vdd gnd cell_6t
Xbit_r27_c30 bl[30] br[30] wl[27] vdd gnd cell_6t
Xbit_r28_c30 bl[30] br[30] wl[28] vdd gnd cell_6t
Xbit_r29_c30 bl[30] br[30] wl[29] vdd gnd cell_6t
Xbit_r30_c30 bl[30] br[30] wl[30] vdd gnd cell_6t
Xbit_r31_c30 bl[30] br[30] wl[31] vdd gnd cell_6t
Xbit_r32_c30 bl[30] br[30] wl[32] vdd gnd cell_6t
Xbit_r33_c30 bl[30] br[30] wl[33] vdd gnd cell_6t
Xbit_r34_c30 bl[30] br[30] wl[34] vdd gnd cell_6t
Xbit_r35_c30 bl[30] br[30] wl[35] vdd gnd cell_6t
Xbit_r36_c30 bl[30] br[30] wl[36] vdd gnd cell_6t
Xbit_r37_c30 bl[30] br[30] wl[37] vdd gnd cell_6t
Xbit_r38_c30 bl[30] br[30] wl[38] vdd gnd cell_6t
Xbit_r39_c30 bl[30] br[30] wl[39] vdd gnd cell_6t
Xbit_r40_c30 bl[30] br[30] wl[40] vdd gnd cell_6t
Xbit_r41_c30 bl[30] br[30] wl[41] vdd gnd cell_6t
Xbit_r42_c30 bl[30] br[30] wl[42] vdd gnd cell_6t
Xbit_r43_c30 bl[30] br[30] wl[43] vdd gnd cell_6t
Xbit_r44_c30 bl[30] br[30] wl[44] vdd gnd cell_6t
Xbit_r45_c30 bl[30] br[30] wl[45] vdd gnd cell_6t
Xbit_r46_c30 bl[30] br[30] wl[46] vdd gnd cell_6t
Xbit_r47_c30 bl[30] br[30] wl[47] vdd gnd cell_6t
Xbit_r48_c30 bl[30] br[30] wl[48] vdd gnd cell_6t
Xbit_r49_c30 bl[30] br[30] wl[49] vdd gnd cell_6t
Xbit_r50_c30 bl[30] br[30] wl[50] vdd gnd cell_6t
Xbit_r51_c30 bl[30] br[30] wl[51] vdd gnd cell_6t
Xbit_r52_c30 bl[30] br[30] wl[52] vdd gnd cell_6t
Xbit_r53_c30 bl[30] br[30] wl[53] vdd gnd cell_6t
Xbit_r54_c30 bl[30] br[30] wl[54] vdd gnd cell_6t
Xbit_r55_c30 bl[30] br[30] wl[55] vdd gnd cell_6t
Xbit_r56_c30 bl[30] br[30] wl[56] vdd gnd cell_6t
Xbit_r57_c30 bl[30] br[30] wl[57] vdd gnd cell_6t
Xbit_r58_c30 bl[30] br[30] wl[58] vdd gnd cell_6t
Xbit_r59_c30 bl[30] br[30] wl[59] vdd gnd cell_6t
Xbit_r60_c30 bl[30] br[30] wl[60] vdd gnd cell_6t
Xbit_r61_c30 bl[30] br[30] wl[61] vdd gnd cell_6t
Xbit_r62_c30 bl[30] br[30] wl[62] vdd gnd cell_6t
Xbit_r63_c30 bl[30] br[30] wl[63] vdd gnd cell_6t
Xbit_r64_c30 bl[30] br[30] wl[64] vdd gnd cell_6t
Xbit_r65_c30 bl[30] br[30] wl[65] vdd gnd cell_6t
Xbit_r66_c30 bl[30] br[30] wl[66] vdd gnd cell_6t
Xbit_r67_c30 bl[30] br[30] wl[67] vdd gnd cell_6t
Xbit_r68_c30 bl[30] br[30] wl[68] vdd gnd cell_6t
Xbit_r69_c30 bl[30] br[30] wl[69] vdd gnd cell_6t
Xbit_r70_c30 bl[30] br[30] wl[70] vdd gnd cell_6t
Xbit_r71_c30 bl[30] br[30] wl[71] vdd gnd cell_6t
Xbit_r72_c30 bl[30] br[30] wl[72] vdd gnd cell_6t
Xbit_r73_c30 bl[30] br[30] wl[73] vdd gnd cell_6t
Xbit_r74_c30 bl[30] br[30] wl[74] vdd gnd cell_6t
Xbit_r75_c30 bl[30] br[30] wl[75] vdd gnd cell_6t
Xbit_r76_c30 bl[30] br[30] wl[76] vdd gnd cell_6t
Xbit_r77_c30 bl[30] br[30] wl[77] vdd gnd cell_6t
Xbit_r78_c30 bl[30] br[30] wl[78] vdd gnd cell_6t
Xbit_r79_c30 bl[30] br[30] wl[79] vdd gnd cell_6t
Xbit_r80_c30 bl[30] br[30] wl[80] vdd gnd cell_6t
Xbit_r81_c30 bl[30] br[30] wl[81] vdd gnd cell_6t
Xbit_r82_c30 bl[30] br[30] wl[82] vdd gnd cell_6t
Xbit_r83_c30 bl[30] br[30] wl[83] vdd gnd cell_6t
Xbit_r84_c30 bl[30] br[30] wl[84] vdd gnd cell_6t
Xbit_r85_c30 bl[30] br[30] wl[85] vdd gnd cell_6t
Xbit_r86_c30 bl[30] br[30] wl[86] vdd gnd cell_6t
Xbit_r87_c30 bl[30] br[30] wl[87] vdd gnd cell_6t
Xbit_r88_c30 bl[30] br[30] wl[88] vdd gnd cell_6t
Xbit_r89_c30 bl[30] br[30] wl[89] vdd gnd cell_6t
Xbit_r90_c30 bl[30] br[30] wl[90] vdd gnd cell_6t
Xbit_r91_c30 bl[30] br[30] wl[91] vdd gnd cell_6t
Xbit_r92_c30 bl[30] br[30] wl[92] vdd gnd cell_6t
Xbit_r93_c30 bl[30] br[30] wl[93] vdd gnd cell_6t
Xbit_r94_c30 bl[30] br[30] wl[94] vdd gnd cell_6t
Xbit_r95_c30 bl[30] br[30] wl[95] vdd gnd cell_6t
Xbit_r96_c30 bl[30] br[30] wl[96] vdd gnd cell_6t
Xbit_r97_c30 bl[30] br[30] wl[97] vdd gnd cell_6t
Xbit_r98_c30 bl[30] br[30] wl[98] vdd gnd cell_6t
Xbit_r99_c30 bl[30] br[30] wl[99] vdd gnd cell_6t
Xbit_r100_c30 bl[30] br[30] wl[100] vdd gnd cell_6t
Xbit_r101_c30 bl[30] br[30] wl[101] vdd gnd cell_6t
Xbit_r102_c30 bl[30] br[30] wl[102] vdd gnd cell_6t
Xbit_r103_c30 bl[30] br[30] wl[103] vdd gnd cell_6t
Xbit_r104_c30 bl[30] br[30] wl[104] vdd gnd cell_6t
Xbit_r105_c30 bl[30] br[30] wl[105] vdd gnd cell_6t
Xbit_r106_c30 bl[30] br[30] wl[106] vdd gnd cell_6t
Xbit_r107_c30 bl[30] br[30] wl[107] vdd gnd cell_6t
Xbit_r108_c30 bl[30] br[30] wl[108] vdd gnd cell_6t
Xbit_r109_c30 bl[30] br[30] wl[109] vdd gnd cell_6t
Xbit_r110_c30 bl[30] br[30] wl[110] vdd gnd cell_6t
Xbit_r111_c30 bl[30] br[30] wl[111] vdd gnd cell_6t
Xbit_r112_c30 bl[30] br[30] wl[112] vdd gnd cell_6t
Xbit_r113_c30 bl[30] br[30] wl[113] vdd gnd cell_6t
Xbit_r114_c30 bl[30] br[30] wl[114] vdd gnd cell_6t
Xbit_r115_c30 bl[30] br[30] wl[115] vdd gnd cell_6t
Xbit_r116_c30 bl[30] br[30] wl[116] vdd gnd cell_6t
Xbit_r117_c30 bl[30] br[30] wl[117] vdd gnd cell_6t
Xbit_r118_c30 bl[30] br[30] wl[118] vdd gnd cell_6t
Xbit_r119_c30 bl[30] br[30] wl[119] vdd gnd cell_6t
Xbit_r120_c30 bl[30] br[30] wl[120] vdd gnd cell_6t
Xbit_r121_c30 bl[30] br[30] wl[121] vdd gnd cell_6t
Xbit_r122_c30 bl[30] br[30] wl[122] vdd gnd cell_6t
Xbit_r123_c30 bl[30] br[30] wl[123] vdd gnd cell_6t
Xbit_r124_c30 bl[30] br[30] wl[124] vdd gnd cell_6t
Xbit_r125_c30 bl[30] br[30] wl[125] vdd gnd cell_6t
Xbit_r126_c30 bl[30] br[30] wl[126] vdd gnd cell_6t
Xbit_r127_c30 bl[30] br[30] wl[127] vdd gnd cell_6t
Xbit_r128_c30 bl[30] br[30] wl[128] vdd gnd cell_6t
Xbit_r129_c30 bl[30] br[30] wl[129] vdd gnd cell_6t
Xbit_r130_c30 bl[30] br[30] wl[130] vdd gnd cell_6t
Xbit_r131_c30 bl[30] br[30] wl[131] vdd gnd cell_6t
Xbit_r132_c30 bl[30] br[30] wl[132] vdd gnd cell_6t
Xbit_r133_c30 bl[30] br[30] wl[133] vdd gnd cell_6t
Xbit_r134_c30 bl[30] br[30] wl[134] vdd gnd cell_6t
Xbit_r135_c30 bl[30] br[30] wl[135] vdd gnd cell_6t
Xbit_r136_c30 bl[30] br[30] wl[136] vdd gnd cell_6t
Xbit_r137_c30 bl[30] br[30] wl[137] vdd gnd cell_6t
Xbit_r138_c30 bl[30] br[30] wl[138] vdd gnd cell_6t
Xbit_r139_c30 bl[30] br[30] wl[139] vdd gnd cell_6t
Xbit_r140_c30 bl[30] br[30] wl[140] vdd gnd cell_6t
Xbit_r141_c30 bl[30] br[30] wl[141] vdd gnd cell_6t
Xbit_r142_c30 bl[30] br[30] wl[142] vdd gnd cell_6t
Xbit_r143_c30 bl[30] br[30] wl[143] vdd gnd cell_6t
Xbit_r144_c30 bl[30] br[30] wl[144] vdd gnd cell_6t
Xbit_r145_c30 bl[30] br[30] wl[145] vdd gnd cell_6t
Xbit_r146_c30 bl[30] br[30] wl[146] vdd gnd cell_6t
Xbit_r147_c30 bl[30] br[30] wl[147] vdd gnd cell_6t
Xbit_r148_c30 bl[30] br[30] wl[148] vdd gnd cell_6t
Xbit_r149_c30 bl[30] br[30] wl[149] vdd gnd cell_6t
Xbit_r150_c30 bl[30] br[30] wl[150] vdd gnd cell_6t
Xbit_r151_c30 bl[30] br[30] wl[151] vdd gnd cell_6t
Xbit_r152_c30 bl[30] br[30] wl[152] vdd gnd cell_6t
Xbit_r153_c30 bl[30] br[30] wl[153] vdd gnd cell_6t
Xbit_r154_c30 bl[30] br[30] wl[154] vdd gnd cell_6t
Xbit_r155_c30 bl[30] br[30] wl[155] vdd gnd cell_6t
Xbit_r156_c30 bl[30] br[30] wl[156] vdd gnd cell_6t
Xbit_r157_c30 bl[30] br[30] wl[157] vdd gnd cell_6t
Xbit_r158_c30 bl[30] br[30] wl[158] vdd gnd cell_6t
Xbit_r159_c30 bl[30] br[30] wl[159] vdd gnd cell_6t
Xbit_r160_c30 bl[30] br[30] wl[160] vdd gnd cell_6t
Xbit_r161_c30 bl[30] br[30] wl[161] vdd gnd cell_6t
Xbit_r162_c30 bl[30] br[30] wl[162] vdd gnd cell_6t
Xbit_r163_c30 bl[30] br[30] wl[163] vdd gnd cell_6t
Xbit_r164_c30 bl[30] br[30] wl[164] vdd gnd cell_6t
Xbit_r165_c30 bl[30] br[30] wl[165] vdd gnd cell_6t
Xbit_r166_c30 bl[30] br[30] wl[166] vdd gnd cell_6t
Xbit_r167_c30 bl[30] br[30] wl[167] vdd gnd cell_6t
Xbit_r168_c30 bl[30] br[30] wl[168] vdd gnd cell_6t
Xbit_r169_c30 bl[30] br[30] wl[169] vdd gnd cell_6t
Xbit_r170_c30 bl[30] br[30] wl[170] vdd gnd cell_6t
Xbit_r171_c30 bl[30] br[30] wl[171] vdd gnd cell_6t
Xbit_r172_c30 bl[30] br[30] wl[172] vdd gnd cell_6t
Xbit_r173_c30 bl[30] br[30] wl[173] vdd gnd cell_6t
Xbit_r174_c30 bl[30] br[30] wl[174] vdd gnd cell_6t
Xbit_r175_c30 bl[30] br[30] wl[175] vdd gnd cell_6t
Xbit_r176_c30 bl[30] br[30] wl[176] vdd gnd cell_6t
Xbit_r177_c30 bl[30] br[30] wl[177] vdd gnd cell_6t
Xbit_r178_c30 bl[30] br[30] wl[178] vdd gnd cell_6t
Xbit_r179_c30 bl[30] br[30] wl[179] vdd gnd cell_6t
Xbit_r180_c30 bl[30] br[30] wl[180] vdd gnd cell_6t
Xbit_r181_c30 bl[30] br[30] wl[181] vdd gnd cell_6t
Xbit_r182_c30 bl[30] br[30] wl[182] vdd gnd cell_6t
Xbit_r183_c30 bl[30] br[30] wl[183] vdd gnd cell_6t
Xbit_r184_c30 bl[30] br[30] wl[184] vdd gnd cell_6t
Xbit_r185_c30 bl[30] br[30] wl[185] vdd gnd cell_6t
Xbit_r186_c30 bl[30] br[30] wl[186] vdd gnd cell_6t
Xbit_r187_c30 bl[30] br[30] wl[187] vdd gnd cell_6t
Xbit_r188_c30 bl[30] br[30] wl[188] vdd gnd cell_6t
Xbit_r189_c30 bl[30] br[30] wl[189] vdd gnd cell_6t
Xbit_r190_c30 bl[30] br[30] wl[190] vdd gnd cell_6t
Xbit_r191_c30 bl[30] br[30] wl[191] vdd gnd cell_6t
Xbit_r192_c30 bl[30] br[30] wl[192] vdd gnd cell_6t
Xbit_r193_c30 bl[30] br[30] wl[193] vdd gnd cell_6t
Xbit_r194_c30 bl[30] br[30] wl[194] vdd gnd cell_6t
Xbit_r195_c30 bl[30] br[30] wl[195] vdd gnd cell_6t
Xbit_r196_c30 bl[30] br[30] wl[196] vdd gnd cell_6t
Xbit_r197_c30 bl[30] br[30] wl[197] vdd gnd cell_6t
Xbit_r198_c30 bl[30] br[30] wl[198] vdd gnd cell_6t
Xbit_r199_c30 bl[30] br[30] wl[199] vdd gnd cell_6t
Xbit_r200_c30 bl[30] br[30] wl[200] vdd gnd cell_6t
Xbit_r201_c30 bl[30] br[30] wl[201] vdd gnd cell_6t
Xbit_r202_c30 bl[30] br[30] wl[202] vdd gnd cell_6t
Xbit_r203_c30 bl[30] br[30] wl[203] vdd gnd cell_6t
Xbit_r204_c30 bl[30] br[30] wl[204] vdd gnd cell_6t
Xbit_r205_c30 bl[30] br[30] wl[205] vdd gnd cell_6t
Xbit_r206_c30 bl[30] br[30] wl[206] vdd gnd cell_6t
Xbit_r207_c30 bl[30] br[30] wl[207] vdd gnd cell_6t
Xbit_r208_c30 bl[30] br[30] wl[208] vdd gnd cell_6t
Xbit_r209_c30 bl[30] br[30] wl[209] vdd gnd cell_6t
Xbit_r210_c30 bl[30] br[30] wl[210] vdd gnd cell_6t
Xbit_r211_c30 bl[30] br[30] wl[211] vdd gnd cell_6t
Xbit_r212_c30 bl[30] br[30] wl[212] vdd gnd cell_6t
Xbit_r213_c30 bl[30] br[30] wl[213] vdd gnd cell_6t
Xbit_r214_c30 bl[30] br[30] wl[214] vdd gnd cell_6t
Xbit_r215_c30 bl[30] br[30] wl[215] vdd gnd cell_6t
Xbit_r216_c30 bl[30] br[30] wl[216] vdd gnd cell_6t
Xbit_r217_c30 bl[30] br[30] wl[217] vdd gnd cell_6t
Xbit_r218_c30 bl[30] br[30] wl[218] vdd gnd cell_6t
Xbit_r219_c30 bl[30] br[30] wl[219] vdd gnd cell_6t
Xbit_r220_c30 bl[30] br[30] wl[220] vdd gnd cell_6t
Xbit_r221_c30 bl[30] br[30] wl[221] vdd gnd cell_6t
Xbit_r222_c30 bl[30] br[30] wl[222] vdd gnd cell_6t
Xbit_r223_c30 bl[30] br[30] wl[223] vdd gnd cell_6t
Xbit_r224_c30 bl[30] br[30] wl[224] vdd gnd cell_6t
Xbit_r225_c30 bl[30] br[30] wl[225] vdd gnd cell_6t
Xbit_r226_c30 bl[30] br[30] wl[226] vdd gnd cell_6t
Xbit_r227_c30 bl[30] br[30] wl[227] vdd gnd cell_6t
Xbit_r228_c30 bl[30] br[30] wl[228] vdd gnd cell_6t
Xbit_r229_c30 bl[30] br[30] wl[229] vdd gnd cell_6t
Xbit_r230_c30 bl[30] br[30] wl[230] vdd gnd cell_6t
Xbit_r231_c30 bl[30] br[30] wl[231] vdd gnd cell_6t
Xbit_r232_c30 bl[30] br[30] wl[232] vdd gnd cell_6t
Xbit_r233_c30 bl[30] br[30] wl[233] vdd gnd cell_6t
Xbit_r234_c30 bl[30] br[30] wl[234] vdd gnd cell_6t
Xbit_r235_c30 bl[30] br[30] wl[235] vdd gnd cell_6t
Xbit_r236_c30 bl[30] br[30] wl[236] vdd gnd cell_6t
Xbit_r237_c30 bl[30] br[30] wl[237] vdd gnd cell_6t
Xbit_r238_c30 bl[30] br[30] wl[238] vdd gnd cell_6t
Xbit_r239_c30 bl[30] br[30] wl[239] vdd gnd cell_6t
Xbit_r240_c30 bl[30] br[30] wl[240] vdd gnd cell_6t
Xbit_r241_c30 bl[30] br[30] wl[241] vdd gnd cell_6t
Xbit_r242_c30 bl[30] br[30] wl[242] vdd gnd cell_6t
Xbit_r243_c30 bl[30] br[30] wl[243] vdd gnd cell_6t
Xbit_r244_c30 bl[30] br[30] wl[244] vdd gnd cell_6t
Xbit_r245_c30 bl[30] br[30] wl[245] vdd gnd cell_6t
Xbit_r246_c30 bl[30] br[30] wl[246] vdd gnd cell_6t
Xbit_r247_c30 bl[30] br[30] wl[247] vdd gnd cell_6t
Xbit_r248_c30 bl[30] br[30] wl[248] vdd gnd cell_6t
Xbit_r249_c30 bl[30] br[30] wl[249] vdd gnd cell_6t
Xbit_r250_c30 bl[30] br[30] wl[250] vdd gnd cell_6t
Xbit_r251_c30 bl[30] br[30] wl[251] vdd gnd cell_6t
Xbit_r252_c30 bl[30] br[30] wl[252] vdd gnd cell_6t
Xbit_r253_c30 bl[30] br[30] wl[253] vdd gnd cell_6t
Xbit_r254_c30 bl[30] br[30] wl[254] vdd gnd cell_6t
Xbit_r255_c30 bl[30] br[30] wl[255] vdd gnd cell_6t
Xbit_r256_c30 bl[30] br[30] wl[256] vdd gnd cell_6t
Xbit_r257_c30 bl[30] br[30] wl[257] vdd gnd cell_6t
Xbit_r258_c30 bl[30] br[30] wl[258] vdd gnd cell_6t
Xbit_r259_c30 bl[30] br[30] wl[259] vdd gnd cell_6t
Xbit_r260_c30 bl[30] br[30] wl[260] vdd gnd cell_6t
Xbit_r261_c30 bl[30] br[30] wl[261] vdd gnd cell_6t
Xbit_r262_c30 bl[30] br[30] wl[262] vdd gnd cell_6t
Xbit_r263_c30 bl[30] br[30] wl[263] vdd gnd cell_6t
Xbit_r264_c30 bl[30] br[30] wl[264] vdd gnd cell_6t
Xbit_r265_c30 bl[30] br[30] wl[265] vdd gnd cell_6t
Xbit_r266_c30 bl[30] br[30] wl[266] vdd gnd cell_6t
Xbit_r267_c30 bl[30] br[30] wl[267] vdd gnd cell_6t
Xbit_r268_c30 bl[30] br[30] wl[268] vdd gnd cell_6t
Xbit_r269_c30 bl[30] br[30] wl[269] vdd gnd cell_6t
Xbit_r270_c30 bl[30] br[30] wl[270] vdd gnd cell_6t
Xbit_r271_c30 bl[30] br[30] wl[271] vdd gnd cell_6t
Xbit_r272_c30 bl[30] br[30] wl[272] vdd gnd cell_6t
Xbit_r273_c30 bl[30] br[30] wl[273] vdd gnd cell_6t
Xbit_r274_c30 bl[30] br[30] wl[274] vdd gnd cell_6t
Xbit_r275_c30 bl[30] br[30] wl[275] vdd gnd cell_6t
Xbit_r276_c30 bl[30] br[30] wl[276] vdd gnd cell_6t
Xbit_r277_c30 bl[30] br[30] wl[277] vdd gnd cell_6t
Xbit_r278_c30 bl[30] br[30] wl[278] vdd gnd cell_6t
Xbit_r279_c30 bl[30] br[30] wl[279] vdd gnd cell_6t
Xbit_r280_c30 bl[30] br[30] wl[280] vdd gnd cell_6t
Xbit_r281_c30 bl[30] br[30] wl[281] vdd gnd cell_6t
Xbit_r282_c30 bl[30] br[30] wl[282] vdd gnd cell_6t
Xbit_r283_c30 bl[30] br[30] wl[283] vdd gnd cell_6t
Xbit_r284_c30 bl[30] br[30] wl[284] vdd gnd cell_6t
Xbit_r285_c30 bl[30] br[30] wl[285] vdd gnd cell_6t
Xbit_r286_c30 bl[30] br[30] wl[286] vdd gnd cell_6t
Xbit_r287_c30 bl[30] br[30] wl[287] vdd gnd cell_6t
Xbit_r288_c30 bl[30] br[30] wl[288] vdd gnd cell_6t
Xbit_r289_c30 bl[30] br[30] wl[289] vdd gnd cell_6t
Xbit_r290_c30 bl[30] br[30] wl[290] vdd gnd cell_6t
Xbit_r291_c30 bl[30] br[30] wl[291] vdd gnd cell_6t
Xbit_r292_c30 bl[30] br[30] wl[292] vdd gnd cell_6t
Xbit_r293_c30 bl[30] br[30] wl[293] vdd gnd cell_6t
Xbit_r294_c30 bl[30] br[30] wl[294] vdd gnd cell_6t
Xbit_r295_c30 bl[30] br[30] wl[295] vdd gnd cell_6t
Xbit_r296_c30 bl[30] br[30] wl[296] vdd gnd cell_6t
Xbit_r297_c30 bl[30] br[30] wl[297] vdd gnd cell_6t
Xbit_r298_c30 bl[30] br[30] wl[298] vdd gnd cell_6t
Xbit_r299_c30 bl[30] br[30] wl[299] vdd gnd cell_6t
Xbit_r300_c30 bl[30] br[30] wl[300] vdd gnd cell_6t
Xbit_r301_c30 bl[30] br[30] wl[301] vdd gnd cell_6t
Xbit_r302_c30 bl[30] br[30] wl[302] vdd gnd cell_6t
Xbit_r303_c30 bl[30] br[30] wl[303] vdd gnd cell_6t
Xbit_r304_c30 bl[30] br[30] wl[304] vdd gnd cell_6t
Xbit_r305_c30 bl[30] br[30] wl[305] vdd gnd cell_6t
Xbit_r306_c30 bl[30] br[30] wl[306] vdd gnd cell_6t
Xbit_r307_c30 bl[30] br[30] wl[307] vdd gnd cell_6t
Xbit_r308_c30 bl[30] br[30] wl[308] vdd gnd cell_6t
Xbit_r309_c30 bl[30] br[30] wl[309] vdd gnd cell_6t
Xbit_r310_c30 bl[30] br[30] wl[310] vdd gnd cell_6t
Xbit_r311_c30 bl[30] br[30] wl[311] vdd gnd cell_6t
Xbit_r312_c30 bl[30] br[30] wl[312] vdd gnd cell_6t
Xbit_r313_c30 bl[30] br[30] wl[313] vdd gnd cell_6t
Xbit_r314_c30 bl[30] br[30] wl[314] vdd gnd cell_6t
Xbit_r315_c30 bl[30] br[30] wl[315] vdd gnd cell_6t
Xbit_r316_c30 bl[30] br[30] wl[316] vdd gnd cell_6t
Xbit_r317_c30 bl[30] br[30] wl[317] vdd gnd cell_6t
Xbit_r318_c30 bl[30] br[30] wl[318] vdd gnd cell_6t
Xbit_r319_c30 bl[30] br[30] wl[319] vdd gnd cell_6t
Xbit_r320_c30 bl[30] br[30] wl[320] vdd gnd cell_6t
Xbit_r321_c30 bl[30] br[30] wl[321] vdd gnd cell_6t
Xbit_r322_c30 bl[30] br[30] wl[322] vdd gnd cell_6t
Xbit_r323_c30 bl[30] br[30] wl[323] vdd gnd cell_6t
Xbit_r324_c30 bl[30] br[30] wl[324] vdd gnd cell_6t
Xbit_r325_c30 bl[30] br[30] wl[325] vdd gnd cell_6t
Xbit_r326_c30 bl[30] br[30] wl[326] vdd gnd cell_6t
Xbit_r327_c30 bl[30] br[30] wl[327] vdd gnd cell_6t
Xbit_r328_c30 bl[30] br[30] wl[328] vdd gnd cell_6t
Xbit_r329_c30 bl[30] br[30] wl[329] vdd gnd cell_6t
Xbit_r330_c30 bl[30] br[30] wl[330] vdd gnd cell_6t
Xbit_r331_c30 bl[30] br[30] wl[331] vdd gnd cell_6t
Xbit_r332_c30 bl[30] br[30] wl[332] vdd gnd cell_6t
Xbit_r333_c30 bl[30] br[30] wl[333] vdd gnd cell_6t
Xbit_r334_c30 bl[30] br[30] wl[334] vdd gnd cell_6t
Xbit_r335_c30 bl[30] br[30] wl[335] vdd gnd cell_6t
Xbit_r336_c30 bl[30] br[30] wl[336] vdd gnd cell_6t
Xbit_r337_c30 bl[30] br[30] wl[337] vdd gnd cell_6t
Xbit_r338_c30 bl[30] br[30] wl[338] vdd gnd cell_6t
Xbit_r339_c30 bl[30] br[30] wl[339] vdd gnd cell_6t
Xbit_r340_c30 bl[30] br[30] wl[340] vdd gnd cell_6t
Xbit_r341_c30 bl[30] br[30] wl[341] vdd gnd cell_6t
Xbit_r342_c30 bl[30] br[30] wl[342] vdd gnd cell_6t
Xbit_r343_c30 bl[30] br[30] wl[343] vdd gnd cell_6t
Xbit_r344_c30 bl[30] br[30] wl[344] vdd gnd cell_6t
Xbit_r345_c30 bl[30] br[30] wl[345] vdd gnd cell_6t
Xbit_r346_c30 bl[30] br[30] wl[346] vdd gnd cell_6t
Xbit_r347_c30 bl[30] br[30] wl[347] vdd gnd cell_6t
Xbit_r348_c30 bl[30] br[30] wl[348] vdd gnd cell_6t
Xbit_r349_c30 bl[30] br[30] wl[349] vdd gnd cell_6t
Xbit_r350_c30 bl[30] br[30] wl[350] vdd gnd cell_6t
Xbit_r351_c30 bl[30] br[30] wl[351] vdd gnd cell_6t
Xbit_r352_c30 bl[30] br[30] wl[352] vdd gnd cell_6t
Xbit_r353_c30 bl[30] br[30] wl[353] vdd gnd cell_6t
Xbit_r354_c30 bl[30] br[30] wl[354] vdd gnd cell_6t
Xbit_r355_c30 bl[30] br[30] wl[355] vdd gnd cell_6t
Xbit_r356_c30 bl[30] br[30] wl[356] vdd gnd cell_6t
Xbit_r357_c30 bl[30] br[30] wl[357] vdd gnd cell_6t
Xbit_r358_c30 bl[30] br[30] wl[358] vdd gnd cell_6t
Xbit_r359_c30 bl[30] br[30] wl[359] vdd gnd cell_6t
Xbit_r360_c30 bl[30] br[30] wl[360] vdd gnd cell_6t
Xbit_r361_c30 bl[30] br[30] wl[361] vdd gnd cell_6t
Xbit_r362_c30 bl[30] br[30] wl[362] vdd gnd cell_6t
Xbit_r363_c30 bl[30] br[30] wl[363] vdd gnd cell_6t
Xbit_r364_c30 bl[30] br[30] wl[364] vdd gnd cell_6t
Xbit_r365_c30 bl[30] br[30] wl[365] vdd gnd cell_6t
Xbit_r366_c30 bl[30] br[30] wl[366] vdd gnd cell_6t
Xbit_r367_c30 bl[30] br[30] wl[367] vdd gnd cell_6t
Xbit_r368_c30 bl[30] br[30] wl[368] vdd gnd cell_6t
Xbit_r369_c30 bl[30] br[30] wl[369] vdd gnd cell_6t
Xbit_r370_c30 bl[30] br[30] wl[370] vdd gnd cell_6t
Xbit_r371_c30 bl[30] br[30] wl[371] vdd gnd cell_6t
Xbit_r372_c30 bl[30] br[30] wl[372] vdd gnd cell_6t
Xbit_r373_c30 bl[30] br[30] wl[373] vdd gnd cell_6t
Xbit_r374_c30 bl[30] br[30] wl[374] vdd gnd cell_6t
Xbit_r375_c30 bl[30] br[30] wl[375] vdd gnd cell_6t
Xbit_r376_c30 bl[30] br[30] wl[376] vdd gnd cell_6t
Xbit_r377_c30 bl[30] br[30] wl[377] vdd gnd cell_6t
Xbit_r378_c30 bl[30] br[30] wl[378] vdd gnd cell_6t
Xbit_r379_c30 bl[30] br[30] wl[379] vdd gnd cell_6t
Xbit_r380_c30 bl[30] br[30] wl[380] vdd gnd cell_6t
Xbit_r381_c30 bl[30] br[30] wl[381] vdd gnd cell_6t
Xbit_r382_c30 bl[30] br[30] wl[382] vdd gnd cell_6t
Xbit_r383_c30 bl[30] br[30] wl[383] vdd gnd cell_6t
Xbit_r384_c30 bl[30] br[30] wl[384] vdd gnd cell_6t
Xbit_r385_c30 bl[30] br[30] wl[385] vdd gnd cell_6t
Xbit_r386_c30 bl[30] br[30] wl[386] vdd gnd cell_6t
Xbit_r387_c30 bl[30] br[30] wl[387] vdd gnd cell_6t
Xbit_r388_c30 bl[30] br[30] wl[388] vdd gnd cell_6t
Xbit_r389_c30 bl[30] br[30] wl[389] vdd gnd cell_6t
Xbit_r390_c30 bl[30] br[30] wl[390] vdd gnd cell_6t
Xbit_r391_c30 bl[30] br[30] wl[391] vdd gnd cell_6t
Xbit_r392_c30 bl[30] br[30] wl[392] vdd gnd cell_6t
Xbit_r393_c30 bl[30] br[30] wl[393] vdd gnd cell_6t
Xbit_r394_c30 bl[30] br[30] wl[394] vdd gnd cell_6t
Xbit_r395_c30 bl[30] br[30] wl[395] vdd gnd cell_6t
Xbit_r396_c30 bl[30] br[30] wl[396] vdd gnd cell_6t
Xbit_r397_c30 bl[30] br[30] wl[397] vdd gnd cell_6t
Xbit_r398_c30 bl[30] br[30] wl[398] vdd gnd cell_6t
Xbit_r399_c30 bl[30] br[30] wl[399] vdd gnd cell_6t
Xbit_r400_c30 bl[30] br[30] wl[400] vdd gnd cell_6t
Xbit_r401_c30 bl[30] br[30] wl[401] vdd gnd cell_6t
Xbit_r402_c30 bl[30] br[30] wl[402] vdd gnd cell_6t
Xbit_r403_c30 bl[30] br[30] wl[403] vdd gnd cell_6t
Xbit_r404_c30 bl[30] br[30] wl[404] vdd gnd cell_6t
Xbit_r405_c30 bl[30] br[30] wl[405] vdd gnd cell_6t
Xbit_r406_c30 bl[30] br[30] wl[406] vdd gnd cell_6t
Xbit_r407_c30 bl[30] br[30] wl[407] vdd gnd cell_6t
Xbit_r408_c30 bl[30] br[30] wl[408] vdd gnd cell_6t
Xbit_r409_c30 bl[30] br[30] wl[409] vdd gnd cell_6t
Xbit_r410_c30 bl[30] br[30] wl[410] vdd gnd cell_6t
Xbit_r411_c30 bl[30] br[30] wl[411] vdd gnd cell_6t
Xbit_r412_c30 bl[30] br[30] wl[412] vdd gnd cell_6t
Xbit_r413_c30 bl[30] br[30] wl[413] vdd gnd cell_6t
Xbit_r414_c30 bl[30] br[30] wl[414] vdd gnd cell_6t
Xbit_r415_c30 bl[30] br[30] wl[415] vdd gnd cell_6t
Xbit_r416_c30 bl[30] br[30] wl[416] vdd gnd cell_6t
Xbit_r417_c30 bl[30] br[30] wl[417] vdd gnd cell_6t
Xbit_r418_c30 bl[30] br[30] wl[418] vdd gnd cell_6t
Xbit_r419_c30 bl[30] br[30] wl[419] vdd gnd cell_6t
Xbit_r420_c30 bl[30] br[30] wl[420] vdd gnd cell_6t
Xbit_r421_c30 bl[30] br[30] wl[421] vdd gnd cell_6t
Xbit_r422_c30 bl[30] br[30] wl[422] vdd gnd cell_6t
Xbit_r423_c30 bl[30] br[30] wl[423] vdd gnd cell_6t
Xbit_r424_c30 bl[30] br[30] wl[424] vdd gnd cell_6t
Xbit_r425_c30 bl[30] br[30] wl[425] vdd gnd cell_6t
Xbit_r426_c30 bl[30] br[30] wl[426] vdd gnd cell_6t
Xbit_r427_c30 bl[30] br[30] wl[427] vdd gnd cell_6t
Xbit_r428_c30 bl[30] br[30] wl[428] vdd gnd cell_6t
Xbit_r429_c30 bl[30] br[30] wl[429] vdd gnd cell_6t
Xbit_r430_c30 bl[30] br[30] wl[430] vdd gnd cell_6t
Xbit_r431_c30 bl[30] br[30] wl[431] vdd gnd cell_6t
Xbit_r432_c30 bl[30] br[30] wl[432] vdd gnd cell_6t
Xbit_r433_c30 bl[30] br[30] wl[433] vdd gnd cell_6t
Xbit_r434_c30 bl[30] br[30] wl[434] vdd gnd cell_6t
Xbit_r435_c30 bl[30] br[30] wl[435] vdd gnd cell_6t
Xbit_r436_c30 bl[30] br[30] wl[436] vdd gnd cell_6t
Xbit_r437_c30 bl[30] br[30] wl[437] vdd gnd cell_6t
Xbit_r438_c30 bl[30] br[30] wl[438] vdd gnd cell_6t
Xbit_r439_c30 bl[30] br[30] wl[439] vdd gnd cell_6t
Xbit_r440_c30 bl[30] br[30] wl[440] vdd gnd cell_6t
Xbit_r441_c30 bl[30] br[30] wl[441] vdd gnd cell_6t
Xbit_r442_c30 bl[30] br[30] wl[442] vdd gnd cell_6t
Xbit_r443_c30 bl[30] br[30] wl[443] vdd gnd cell_6t
Xbit_r444_c30 bl[30] br[30] wl[444] vdd gnd cell_6t
Xbit_r445_c30 bl[30] br[30] wl[445] vdd gnd cell_6t
Xbit_r446_c30 bl[30] br[30] wl[446] vdd gnd cell_6t
Xbit_r447_c30 bl[30] br[30] wl[447] vdd gnd cell_6t
Xbit_r448_c30 bl[30] br[30] wl[448] vdd gnd cell_6t
Xbit_r449_c30 bl[30] br[30] wl[449] vdd gnd cell_6t
Xbit_r450_c30 bl[30] br[30] wl[450] vdd gnd cell_6t
Xbit_r451_c30 bl[30] br[30] wl[451] vdd gnd cell_6t
Xbit_r452_c30 bl[30] br[30] wl[452] vdd gnd cell_6t
Xbit_r453_c30 bl[30] br[30] wl[453] vdd gnd cell_6t
Xbit_r454_c30 bl[30] br[30] wl[454] vdd gnd cell_6t
Xbit_r455_c30 bl[30] br[30] wl[455] vdd gnd cell_6t
Xbit_r456_c30 bl[30] br[30] wl[456] vdd gnd cell_6t
Xbit_r457_c30 bl[30] br[30] wl[457] vdd gnd cell_6t
Xbit_r458_c30 bl[30] br[30] wl[458] vdd gnd cell_6t
Xbit_r459_c30 bl[30] br[30] wl[459] vdd gnd cell_6t
Xbit_r460_c30 bl[30] br[30] wl[460] vdd gnd cell_6t
Xbit_r461_c30 bl[30] br[30] wl[461] vdd gnd cell_6t
Xbit_r462_c30 bl[30] br[30] wl[462] vdd gnd cell_6t
Xbit_r463_c30 bl[30] br[30] wl[463] vdd gnd cell_6t
Xbit_r464_c30 bl[30] br[30] wl[464] vdd gnd cell_6t
Xbit_r465_c30 bl[30] br[30] wl[465] vdd gnd cell_6t
Xbit_r466_c30 bl[30] br[30] wl[466] vdd gnd cell_6t
Xbit_r467_c30 bl[30] br[30] wl[467] vdd gnd cell_6t
Xbit_r468_c30 bl[30] br[30] wl[468] vdd gnd cell_6t
Xbit_r469_c30 bl[30] br[30] wl[469] vdd gnd cell_6t
Xbit_r470_c30 bl[30] br[30] wl[470] vdd gnd cell_6t
Xbit_r471_c30 bl[30] br[30] wl[471] vdd gnd cell_6t
Xbit_r472_c30 bl[30] br[30] wl[472] vdd gnd cell_6t
Xbit_r473_c30 bl[30] br[30] wl[473] vdd gnd cell_6t
Xbit_r474_c30 bl[30] br[30] wl[474] vdd gnd cell_6t
Xbit_r475_c30 bl[30] br[30] wl[475] vdd gnd cell_6t
Xbit_r476_c30 bl[30] br[30] wl[476] vdd gnd cell_6t
Xbit_r477_c30 bl[30] br[30] wl[477] vdd gnd cell_6t
Xbit_r478_c30 bl[30] br[30] wl[478] vdd gnd cell_6t
Xbit_r479_c30 bl[30] br[30] wl[479] vdd gnd cell_6t
Xbit_r480_c30 bl[30] br[30] wl[480] vdd gnd cell_6t
Xbit_r481_c30 bl[30] br[30] wl[481] vdd gnd cell_6t
Xbit_r482_c30 bl[30] br[30] wl[482] vdd gnd cell_6t
Xbit_r483_c30 bl[30] br[30] wl[483] vdd gnd cell_6t
Xbit_r484_c30 bl[30] br[30] wl[484] vdd gnd cell_6t
Xbit_r485_c30 bl[30] br[30] wl[485] vdd gnd cell_6t
Xbit_r486_c30 bl[30] br[30] wl[486] vdd gnd cell_6t
Xbit_r487_c30 bl[30] br[30] wl[487] vdd gnd cell_6t
Xbit_r488_c30 bl[30] br[30] wl[488] vdd gnd cell_6t
Xbit_r489_c30 bl[30] br[30] wl[489] vdd gnd cell_6t
Xbit_r490_c30 bl[30] br[30] wl[490] vdd gnd cell_6t
Xbit_r491_c30 bl[30] br[30] wl[491] vdd gnd cell_6t
Xbit_r492_c30 bl[30] br[30] wl[492] vdd gnd cell_6t
Xbit_r493_c30 bl[30] br[30] wl[493] vdd gnd cell_6t
Xbit_r494_c30 bl[30] br[30] wl[494] vdd gnd cell_6t
Xbit_r495_c30 bl[30] br[30] wl[495] vdd gnd cell_6t
Xbit_r496_c30 bl[30] br[30] wl[496] vdd gnd cell_6t
Xbit_r497_c30 bl[30] br[30] wl[497] vdd gnd cell_6t
Xbit_r498_c30 bl[30] br[30] wl[498] vdd gnd cell_6t
Xbit_r499_c30 bl[30] br[30] wl[499] vdd gnd cell_6t
Xbit_r500_c30 bl[30] br[30] wl[500] vdd gnd cell_6t
Xbit_r501_c30 bl[30] br[30] wl[501] vdd gnd cell_6t
Xbit_r502_c30 bl[30] br[30] wl[502] vdd gnd cell_6t
Xbit_r503_c30 bl[30] br[30] wl[503] vdd gnd cell_6t
Xbit_r504_c30 bl[30] br[30] wl[504] vdd gnd cell_6t
Xbit_r505_c30 bl[30] br[30] wl[505] vdd gnd cell_6t
Xbit_r506_c30 bl[30] br[30] wl[506] vdd gnd cell_6t
Xbit_r507_c30 bl[30] br[30] wl[507] vdd gnd cell_6t
Xbit_r508_c30 bl[30] br[30] wl[508] vdd gnd cell_6t
Xbit_r509_c30 bl[30] br[30] wl[509] vdd gnd cell_6t
Xbit_r510_c30 bl[30] br[30] wl[510] vdd gnd cell_6t
Xbit_r511_c30 bl[30] br[30] wl[511] vdd gnd cell_6t
Xbit_r0_c31 bl[31] br[31] wl[0] vdd gnd cell_6t
Xbit_r1_c31 bl[31] br[31] wl[1] vdd gnd cell_6t
Xbit_r2_c31 bl[31] br[31] wl[2] vdd gnd cell_6t
Xbit_r3_c31 bl[31] br[31] wl[3] vdd gnd cell_6t
Xbit_r4_c31 bl[31] br[31] wl[4] vdd gnd cell_6t
Xbit_r5_c31 bl[31] br[31] wl[5] vdd gnd cell_6t
Xbit_r6_c31 bl[31] br[31] wl[6] vdd gnd cell_6t
Xbit_r7_c31 bl[31] br[31] wl[7] vdd gnd cell_6t
Xbit_r8_c31 bl[31] br[31] wl[8] vdd gnd cell_6t
Xbit_r9_c31 bl[31] br[31] wl[9] vdd gnd cell_6t
Xbit_r10_c31 bl[31] br[31] wl[10] vdd gnd cell_6t
Xbit_r11_c31 bl[31] br[31] wl[11] vdd gnd cell_6t
Xbit_r12_c31 bl[31] br[31] wl[12] vdd gnd cell_6t
Xbit_r13_c31 bl[31] br[31] wl[13] vdd gnd cell_6t
Xbit_r14_c31 bl[31] br[31] wl[14] vdd gnd cell_6t
Xbit_r15_c31 bl[31] br[31] wl[15] vdd gnd cell_6t
Xbit_r16_c31 bl[31] br[31] wl[16] vdd gnd cell_6t
Xbit_r17_c31 bl[31] br[31] wl[17] vdd gnd cell_6t
Xbit_r18_c31 bl[31] br[31] wl[18] vdd gnd cell_6t
Xbit_r19_c31 bl[31] br[31] wl[19] vdd gnd cell_6t
Xbit_r20_c31 bl[31] br[31] wl[20] vdd gnd cell_6t
Xbit_r21_c31 bl[31] br[31] wl[21] vdd gnd cell_6t
Xbit_r22_c31 bl[31] br[31] wl[22] vdd gnd cell_6t
Xbit_r23_c31 bl[31] br[31] wl[23] vdd gnd cell_6t
Xbit_r24_c31 bl[31] br[31] wl[24] vdd gnd cell_6t
Xbit_r25_c31 bl[31] br[31] wl[25] vdd gnd cell_6t
Xbit_r26_c31 bl[31] br[31] wl[26] vdd gnd cell_6t
Xbit_r27_c31 bl[31] br[31] wl[27] vdd gnd cell_6t
Xbit_r28_c31 bl[31] br[31] wl[28] vdd gnd cell_6t
Xbit_r29_c31 bl[31] br[31] wl[29] vdd gnd cell_6t
Xbit_r30_c31 bl[31] br[31] wl[30] vdd gnd cell_6t
Xbit_r31_c31 bl[31] br[31] wl[31] vdd gnd cell_6t
Xbit_r32_c31 bl[31] br[31] wl[32] vdd gnd cell_6t
Xbit_r33_c31 bl[31] br[31] wl[33] vdd gnd cell_6t
Xbit_r34_c31 bl[31] br[31] wl[34] vdd gnd cell_6t
Xbit_r35_c31 bl[31] br[31] wl[35] vdd gnd cell_6t
Xbit_r36_c31 bl[31] br[31] wl[36] vdd gnd cell_6t
Xbit_r37_c31 bl[31] br[31] wl[37] vdd gnd cell_6t
Xbit_r38_c31 bl[31] br[31] wl[38] vdd gnd cell_6t
Xbit_r39_c31 bl[31] br[31] wl[39] vdd gnd cell_6t
Xbit_r40_c31 bl[31] br[31] wl[40] vdd gnd cell_6t
Xbit_r41_c31 bl[31] br[31] wl[41] vdd gnd cell_6t
Xbit_r42_c31 bl[31] br[31] wl[42] vdd gnd cell_6t
Xbit_r43_c31 bl[31] br[31] wl[43] vdd gnd cell_6t
Xbit_r44_c31 bl[31] br[31] wl[44] vdd gnd cell_6t
Xbit_r45_c31 bl[31] br[31] wl[45] vdd gnd cell_6t
Xbit_r46_c31 bl[31] br[31] wl[46] vdd gnd cell_6t
Xbit_r47_c31 bl[31] br[31] wl[47] vdd gnd cell_6t
Xbit_r48_c31 bl[31] br[31] wl[48] vdd gnd cell_6t
Xbit_r49_c31 bl[31] br[31] wl[49] vdd gnd cell_6t
Xbit_r50_c31 bl[31] br[31] wl[50] vdd gnd cell_6t
Xbit_r51_c31 bl[31] br[31] wl[51] vdd gnd cell_6t
Xbit_r52_c31 bl[31] br[31] wl[52] vdd gnd cell_6t
Xbit_r53_c31 bl[31] br[31] wl[53] vdd gnd cell_6t
Xbit_r54_c31 bl[31] br[31] wl[54] vdd gnd cell_6t
Xbit_r55_c31 bl[31] br[31] wl[55] vdd gnd cell_6t
Xbit_r56_c31 bl[31] br[31] wl[56] vdd gnd cell_6t
Xbit_r57_c31 bl[31] br[31] wl[57] vdd gnd cell_6t
Xbit_r58_c31 bl[31] br[31] wl[58] vdd gnd cell_6t
Xbit_r59_c31 bl[31] br[31] wl[59] vdd gnd cell_6t
Xbit_r60_c31 bl[31] br[31] wl[60] vdd gnd cell_6t
Xbit_r61_c31 bl[31] br[31] wl[61] vdd gnd cell_6t
Xbit_r62_c31 bl[31] br[31] wl[62] vdd gnd cell_6t
Xbit_r63_c31 bl[31] br[31] wl[63] vdd gnd cell_6t
Xbit_r64_c31 bl[31] br[31] wl[64] vdd gnd cell_6t
Xbit_r65_c31 bl[31] br[31] wl[65] vdd gnd cell_6t
Xbit_r66_c31 bl[31] br[31] wl[66] vdd gnd cell_6t
Xbit_r67_c31 bl[31] br[31] wl[67] vdd gnd cell_6t
Xbit_r68_c31 bl[31] br[31] wl[68] vdd gnd cell_6t
Xbit_r69_c31 bl[31] br[31] wl[69] vdd gnd cell_6t
Xbit_r70_c31 bl[31] br[31] wl[70] vdd gnd cell_6t
Xbit_r71_c31 bl[31] br[31] wl[71] vdd gnd cell_6t
Xbit_r72_c31 bl[31] br[31] wl[72] vdd gnd cell_6t
Xbit_r73_c31 bl[31] br[31] wl[73] vdd gnd cell_6t
Xbit_r74_c31 bl[31] br[31] wl[74] vdd gnd cell_6t
Xbit_r75_c31 bl[31] br[31] wl[75] vdd gnd cell_6t
Xbit_r76_c31 bl[31] br[31] wl[76] vdd gnd cell_6t
Xbit_r77_c31 bl[31] br[31] wl[77] vdd gnd cell_6t
Xbit_r78_c31 bl[31] br[31] wl[78] vdd gnd cell_6t
Xbit_r79_c31 bl[31] br[31] wl[79] vdd gnd cell_6t
Xbit_r80_c31 bl[31] br[31] wl[80] vdd gnd cell_6t
Xbit_r81_c31 bl[31] br[31] wl[81] vdd gnd cell_6t
Xbit_r82_c31 bl[31] br[31] wl[82] vdd gnd cell_6t
Xbit_r83_c31 bl[31] br[31] wl[83] vdd gnd cell_6t
Xbit_r84_c31 bl[31] br[31] wl[84] vdd gnd cell_6t
Xbit_r85_c31 bl[31] br[31] wl[85] vdd gnd cell_6t
Xbit_r86_c31 bl[31] br[31] wl[86] vdd gnd cell_6t
Xbit_r87_c31 bl[31] br[31] wl[87] vdd gnd cell_6t
Xbit_r88_c31 bl[31] br[31] wl[88] vdd gnd cell_6t
Xbit_r89_c31 bl[31] br[31] wl[89] vdd gnd cell_6t
Xbit_r90_c31 bl[31] br[31] wl[90] vdd gnd cell_6t
Xbit_r91_c31 bl[31] br[31] wl[91] vdd gnd cell_6t
Xbit_r92_c31 bl[31] br[31] wl[92] vdd gnd cell_6t
Xbit_r93_c31 bl[31] br[31] wl[93] vdd gnd cell_6t
Xbit_r94_c31 bl[31] br[31] wl[94] vdd gnd cell_6t
Xbit_r95_c31 bl[31] br[31] wl[95] vdd gnd cell_6t
Xbit_r96_c31 bl[31] br[31] wl[96] vdd gnd cell_6t
Xbit_r97_c31 bl[31] br[31] wl[97] vdd gnd cell_6t
Xbit_r98_c31 bl[31] br[31] wl[98] vdd gnd cell_6t
Xbit_r99_c31 bl[31] br[31] wl[99] vdd gnd cell_6t
Xbit_r100_c31 bl[31] br[31] wl[100] vdd gnd cell_6t
Xbit_r101_c31 bl[31] br[31] wl[101] vdd gnd cell_6t
Xbit_r102_c31 bl[31] br[31] wl[102] vdd gnd cell_6t
Xbit_r103_c31 bl[31] br[31] wl[103] vdd gnd cell_6t
Xbit_r104_c31 bl[31] br[31] wl[104] vdd gnd cell_6t
Xbit_r105_c31 bl[31] br[31] wl[105] vdd gnd cell_6t
Xbit_r106_c31 bl[31] br[31] wl[106] vdd gnd cell_6t
Xbit_r107_c31 bl[31] br[31] wl[107] vdd gnd cell_6t
Xbit_r108_c31 bl[31] br[31] wl[108] vdd gnd cell_6t
Xbit_r109_c31 bl[31] br[31] wl[109] vdd gnd cell_6t
Xbit_r110_c31 bl[31] br[31] wl[110] vdd gnd cell_6t
Xbit_r111_c31 bl[31] br[31] wl[111] vdd gnd cell_6t
Xbit_r112_c31 bl[31] br[31] wl[112] vdd gnd cell_6t
Xbit_r113_c31 bl[31] br[31] wl[113] vdd gnd cell_6t
Xbit_r114_c31 bl[31] br[31] wl[114] vdd gnd cell_6t
Xbit_r115_c31 bl[31] br[31] wl[115] vdd gnd cell_6t
Xbit_r116_c31 bl[31] br[31] wl[116] vdd gnd cell_6t
Xbit_r117_c31 bl[31] br[31] wl[117] vdd gnd cell_6t
Xbit_r118_c31 bl[31] br[31] wl[118] vdd gnd cell_6t
Xbit_r119_c31 bl[31] br[31] wl[119] vdd gnd cell_6t
Xbit_r120_c31 bl[31] br[31] wl[120] vdd gnd cell_6t
Xbit_r121_c31 bl[31] br[31] wl[121] vdd gnd cell_6t
Xbit_r122_c31 bl[31] br[31] wl[122] vdd gnd cell_6t
Xbit_r123_c31 bl[31] br[31] wl[123] vdd gnd cell_6t
Xbit_r124_c31 bl[31] br[31] wl[124] vdd gnd cell_6t
Xbit_r125_c31 bl[31] br[31] wl[125] vdd gnd cell_6t
Xbit_r126_c31 bl[31] br[31] wl[126] vdd gnd cell_6t
Xbit_r127_c31 bl[31] br[31] wl[127] vdd gnd cell_6t
Xbit_r128_c31 bl[31] br[31] wl[128] vdd gnd cell_6t
Xbit_r129_c31 bl[31] br[31] wl[129] vdd gnd cell_6t
Xbit_r130_c31 bl[31] br[31] wl[130] vdd gnd cell_6t
Xbit_r131_c31 bl[31] br[31] wl[131] vdd gnd cell_6t
Xbit_r132_c31 bl[31] br[31] wl[132] vdd gnd cell_6t
Xbit_r133_c31 bl[31] br[31] wl[133] vdd gnd cell_6t
Xbit_r134_c31 bl[31] br[31] wl[134] vdd gnd cell_6t
Xbit_r135_c31 bl[31] br[31] wl[135] vdd gnd cell_6t
Xbit_r136_c31 bl[31] br[31] wl[136] vdd gnd cell_6t
Xbit_r137_c31 bl[31] br[31] wl[137] vdd gnd cell_6t
Xbit_r138_c31 bl[31] br[31] wl[138] vdd gnd cell_6t
Xbit_r139_c31 bl[31] br[31] wl[139] vdd gnd cell_6t
Xbit_r140_c31 bl[31] br[31] wl[140] vdd gnd cell_6t
Xbit_r141_c31 bl[31] br[31] wl[141] vdd gnd cell_6t
Xbit_r142_c31 bl[31] br[31] wl[142] vdd gnd cell_6t
Xbit_r143_c31 bl[31] br[31] wl[143] vdd gnd cell_6t
Xbit_r144_c31 bl[31] br[31] wl[144] vdd gnd cell_6t
Xbit_r145_c31 bl[31] br[31] wl[145] vdd gnd cell_6t
Xbit_r146_c31 bl[31] br[31] wl[146] vdd gnd cell_6t
Xbit_r147_c31 bl[31] br[31] wl[147] vdd gnd cell_6t
Xbit_r148_c31 bl[31] br[31] wl[148] vdd gnd cell_6t
Xbit_r149_c31 bl[31] br[31] wl[149] vdd gnd cell_6t
Xbit_r150_c31 bl[31] br[31] wl[150] vdd gnd cell_6t
Xbit_r151_c31 bl[31] br[31] wl[151] vdd gnd cell_6t
Xbit_r152_c31 bl[31] br[31] wl[152] vdd gnd cell_6t
Xbit_r153_c31 bl[31] br[31] wl[153] vdd gnd cell_6t
Xbit_r154_c31 bl[31] br[31] wl[154] vdd gnd cell_6t
Xbit_r155_c31 bl[31] br[31] wl[155] vdd gnd cell_6t
Xbit_r156_c31 bl[31] br[31] wl[156] vdd gnd cell_6t
Xbit_r157_c31 bl[31] br[31] wl[157] vdd gnd cell_6t
Xbit_r158_c31 bl[31] br[31] wl[158] vdd gnd cell_6t
Xbit_r159_c31 bl[31] br[31] wl[159] vdd gnd cell_6t
Xbit_r160_c31 bl[31] br[31] wl[160] vdd gnd cell_6t
Xbit_r161_c31 bl[31] br[31] wl[161] vdd gnd cell_6t
Xbit_r162_c31 bl[31] br[31] wl[162] vdd gnd cell_6t
Xbit_r163_c31 bl[31] br[31] wl[163] vdd gnd cell_6t
Xbit_r164_c31 bl[31] br[31] wl[164] vdd gnd cell_6t
Xbit_r165_c31 bl[31] br[31] wl[165] vdd gnd cell_6t
Xbit_r166_c31 bl[31] br[31] wl[166] vdd gnd cell_6t
Xbit_r167_c31 bl[31] br[31] wl[167] vdd gnd cell_6t
Xbit_r168_c31 bl[31] br[31] wl[168] vdd gnd cell_6t
Xbit_r169_c31 bl[31] br[31] wl[169] vdd gnd cell_6t
Xbit_r170_c31 bl[31] br[31] wl[170] vdd gnd cell_6t
Xbit_r171_c31 bl[31] br[31] wl[171] vdd gnd cell_6t
Xbit_r172_c31 bl[31] br[31] wl[172] vdd gnd cell_6t
Xbit_r173_c31 bl[31] br[31] wl[173] vdd gnd cell_6t
Xbit_r174_c31 bl[31] br[31] wl[174] vdd gnd cell_6t
Xbit_r175_c31 bl[31] br[31] wl[175] vdd gnd cell_6t
Xbit_r176_c31 bl[31] br[31] wl[176] vdd gnd cell_6t
Xbit_r177_c31 bl[31] br[31] wl[177] vdd gnd cell_6t
Xbit_r178_c31 bl[31] br[31] wl[178] vdd gnd cell_6t
Xbit_r179_c31 bl[31] br[31] wl[179] vdd gnd cell_6t
Xbit_r180_c31 bl[31] br[31] wl[180] vdd gnd cell_6t
Xbit_r181_c31 bl[31] br[31] wl[181] vdd gnd cell_6t
Xbit_r182_c31 bl[31] br[31] wl[182] vdd gnd cell_6t
Xbit_r183_c31 bl[31] br[31] wl[183] vdd gnd cell_6t
Xbit_r184_c31 bl[31] br[31] wl[184] vdd gnd cell_6t
Xbit_r185_c31 bl[31] br[31] wl[185] vdd gnd cell_6t
Xbit_r186_c31 bl[31] br[31] wl[186] vdd gnd cell_6t
Xbit_r187_c31 bl[31] br[31] wl[187] vdd gnd cell_6t
Xbit_r188_c31 bl[31] br[31] wl[188] vdd gnd cell_6t
Xbit_r189_c31 bl[31] br[31] wl[189] vdd gnd cell_6t
Xbit_r190_c31 bl[31] br[31] wl[190] vdd gnd cell_6t
Xbit_r191_c31 bl[31] br[31] wl[191] vdd gnd cell_6t
Xbit_r192_c31 bl[31] br[31] wl[192] vdd gnd cell_6t
Xbit_r193_c31 bl[31] br[31] wl[193] vdd gnd cell_6t
Xbit_r194_c31 bl[31] br[31] wl[194] vdd gnd cell_6t
Xbit_r195_c31 bl[31] br[31] wl[195] vdd gnd cell_6t
Xbit_r196_c31 bl[31] br[31] wl[196] vdd gnd cell_6t
Xbit_r197_c31 bl[31] br[31] wl[197] vdd gnd cell_6t
Xbit_r198_c31 bl[31] br[31] wl[198] vdd gnd cell_6t
Xbit_r199_c31 bl[31] br[31] wl[199] vdd gnd cell_6t
Xbit_r200_c31 bl[31] br[31] wl[200] vdd gnd cell_6t
Xbit_r201_c31 bl[31] br[31] wl[201] vdd gnd cell_6t
Xbit_r202_c31 bl[31] br[31] wl[202] vdd gnd cell_6t
Xbit_r203_c31 bl[31] br[31] wl[203] vdd gnd cell_6t
Xbit_r204_c31 bl[31] br[31] wl[204] vdd gnd cell_6t
Xbit_r205_c31 bl[31] br[31] wl[205] vdd gnd cell_6t
Xbit_r206_c31 bl[31] br[31] wl[206] vdd gnd cell_6t
Xbit_r207_c31 bl[31] br[31] wl[207] vdd gnd cell_6t
Xbit_r208_c31 bl[31] br[31] wl[208] vdd gnd cell_6t
Xbit_r209_c31 bl[31] br[31] wl[209] vdd gnd cell_6t
Xbit_r210_c31 bl[31] br[31] wl[210] vdd gnd cell_6t
Xbit_r211_c31 bl[31] br[31] wl[211] vdd gnd cell_6t
Xbit_r212_c31 bl[31] br[31] wl[212] vdd gnd cell_6t
Xbit_r213_c31 bl[31] br[31] wl[213] vdd gnd cell_6t
Xbit_r214_c31 bl[31] br[31] wl[214] vdd gnd cell_6t
Xbit_r215_c31 bl[31] br[31] wl[215] vdd gnd cell_6t
Xbit_r216_c31 bl[31] br[31] wl[216] vdd gnd cell_6t
Xbit_r217_c31 bl[31] br[31] wl[217] vdd gnd cell_6t
Xbit_r218_c31 bl[31] br[31] wl[218] vdd gnd cell_6t
Xbit_r219_c31 bl[31] br[31] wl[219] vdd gnd cell_6t
Xbit_r220_c31 bl[31] br[31] wl[220] vdd gnd cell_6t
Xbit_r221_c31 bl[31] br[31] wl[221] vdd gnd cell_6t
Xbit_r222_c31 bl[31] br[31] wl[222] vdd gnd cell_6t
Xbit_r223_c31 bl[31] br[31] wl[223] vdd gnd cell_6t
Xbit_r224_c31 bl[31] br[31] wl[224] vdd gnd cell_6t
Xbit_r225_c31 bl[31] br[31] wl[225] vdd gnd cell_6t
Xbit_r226_c31 bl[31] br[31] wl[226] vdd gnd cell_6t
Xbit_r227_c31 bl[31] br[31] wl[227] vdd gnd cell_6t
Xbit_r228_c31 bl[31] br[31] wl[228] vdd gnd cell_6t
Xbit_r229_c31 bl[31] br[31] wl[229] vdd gnd cell_6t
Xbit_r230_c31 bl[31] br[31] wl[230] vdd gnd cell_6t
Xbit_r231_c31 bl[31] br[31] wl[231] vdd gnd cell_6t
Xbit_r232_c31 bl[31] br[31] wl[232] vdd gnd cell_6t
Xbit_r233_c31 bl[31] br[31] wl[233] vdd gnd cell_6t
Xbit_r234_c31 bl[31] br[31] wl[234] vdd gnd cell_6t
Xbit_r235_c31 bl[31] br[31] wl[235] vdd gnd cell_6t
Xbit_r236_c31 bl[31] br[31] wl[236] vdd gnd cell_6t
Xbit_r237_c31 bl[31] br[31] wl[237] vdd gnd cell_6t
Xbit_r238_c31 bl[31] br[31] wl[238] vdd gnd cell_6t
Xbit_r239_c31 bl[31] br[31] wl[239] vdd gnd cell_6t
Xbit_r240_c31 bl[31] br[31] wl[240] vdd gnd cell_6t
Xbit_r241_c31 bl[31] br[31] wl[241] vdd gnd cell_6t
Xbit_r242_c31 bl[31] br[31] wl[242] vdd gnd cell_6t
Xbit_r243_c31 bl[31] br[31] wl[243] vdd gnd cell_6t
Xbit_r244_c31 bl[31] br[31] wl[244] vdd gnd cell_6t
Xbit_r245_c31 bl[31] br[31] wl[245] vdd gnd cell_6t
Xbit_r246_c31 bl[31] br[31] wl[246] vdd gnd cell_6t
Xbit_r247_c31 bl[31] br[31] wl[247] vdd gnd cell_6t
Xbit_r248_c31 bl[31] br[31] wl[248] vdd gnd cell_6t
Xbit_r249_c31 bl[31] br[31] wl[249] vdd gnd cell_6t
Xbit_r250_c31 bl[31] br[31] wl[250] vdd gnd cell_6t
Xbit_r251_c31 bl[31] br[31] wl[251] vdd gnd cell_6t
Xbit_r252_c31 bl[31] br[31] wl[252] vdd gnd cell_6t
Xbit_r253_c31 bl[31] br[31] wl[253] vdd gnd cell_6t
Xbit_r254_c31 bl[31] br[31] wl[254] vdd gnd cell_6t
Xbit_r255_c31 bl[31] br[31] wl[255] vdd gnd cell_6t
Xbit_r256_c31 bl[31] br[31] wl[256] vdd gnd cell_6t
Xbit_r257_c31 bl[31] br[31] wl[257] vdd gnd cell_6t
Xbit_r258_c31 bl[31] br[31] wl[258] vdd gnd cell_6t
Xbit_r259_c31 bl[31] br[31] wl[259] vdd gnd cell_6t
Xbit_r260_c31 bl[31] br[31] wl[260] vdd gnd cell_6t
Xbit_r261_c31 bl[31] br[31] wl[261] vdd gnd cell_6t
Xbit_r262_c31 bl[31] br[31] wl[262] vdd gnd cell_6t
Xbit_r263_c31 bl[31] br[31] wl[263] vdd gnd cell_6t
Xbit_r264_c31 bl[31] br[31] wl[264] vdd gnd cell_6t
Xbit_r265_c31 bl[31] br[31] wl[265] vdd gnd cell_6t
Xbit_r266_c31 bl[31] br[31] wl[266] vdd gnd cell_6t
Xbit_r267_c31 bl[31] br[31] wl[267] vdd gnd cell_6t
Xbit_r268_c31 bl[31] br[31] wl[268] vdd gnd cell_6t
Xbit_r269_c31 bl[31] br[31] wl[269] vdd gnd cell_6t
Xbit_r270_c31 bl[31] br[31] wl[270] vdd gnd cell_6t
Xbit_r271_c31 bl[31] br[31] wl[271] vdd gnd cell_6t
Xbit_r272_c31 bl[31] br[31] wl[272] vdd gnd cell_6t
Xbit_r273_c31 bl[31] br[31] wl[273] vdd gnd cell_6t
Xbit_r274_c31 bl[31] br[31] wl[274] vdd gnd cell_6t
Xbit_r275_c31 bl[31] br[31] wl[275] vdd gnd cell_6t
Xbit_r276_c31 bl[31] br[31] wl[276] vdd gnd cell_6t
Xbit_r277_c31 bl[31] br[31] wl[277] vdd gnd cell_6t
Xbit_r278_c31 bl[31] br[31] wl[278] vdd gnd cell_6t
Xbit_r279_c31 bl[31] br[31] wl[279] vdd gnd cell_6t
Xbit_r280_c31 bl[31] br[31] wl[280] vdd gnd cell_6t
Xbit_r281_c31 bl[31] br[31] wl[281] vdd gnd cell_6t
Xbit_r282_c31 bl[31] br[31] wl[282] vdd gnd cell_6t
Xbit_r283_c31 bl[31] br[31] wl[283] vdd gnd cell_6t
Xbit_r284_c31 bl[31] br[31] wl[284] vdd gnd cell_6t
Xbit_r285_c31 bl[31] br[31] wl[285] vdd gnd cell_6t
Xbit_r286_c31 bl[31] br[31] wl[286] vdd gnd cell_6t
Xbit_r287_c31 bl[31] br[31] wl[287] vdd gnd cell_6t
Xbit_r288_c31 bl[31] br[31] wl[288] vdd gnd cell_6t
Xbit_r289_c31 bl[31] br[31] wl[289] vdd gnd cell_6t
Xbit_r290_c31 bl[31] br[31] wl[290] vdd gnd cell_6t
Xbit_r291_c31 bl[31] br[31] wl[291] vdd gnd cell_6t
Xbit_r292_c31 bl[31] br[31] wl[292] vdd gnd cell_6t
Xbit_r293_c31 bl[31] br[31] wl[293] vdd gnd cell_6t
Xbit_r294_c31 bl[31] br[31] wl[294] vdd gnd cell_6t
Xbit_r295_c31 bl[31] br[31] wl[295] vdd gnd cell_6t
Xbit_r296_c31 bl[31] br[31] wl[296] vdd gnd cell_6t
Xbit_r297_c31 bl[31] br[31] wl[297] vdd gnd cell_6t
Xbit_r298_c31 bl[31] br[31] wl[298] vdd gnd cell_6t
Xbit_r299_c31 bl[31] br[31] wl[299] vdd gnd cell_6t
Xbit_r300_c31 bl[31] br[31] wl[300] vdd gnd cell_6t
Xbit_r301_c31 bl[31] br[31] wl[301] vdd gnd cell_6t
Xbit_r302_c31 bl[31] br[31] wl[302] vdd gnd cell_6t
Xbit_r303_c31 bl[31] br[31] wl[303] vdd gnd cell_6t
Xbit_r304_c31 bl[31] br[31] wl[304] vdd gnd cell_6t
Xbit_r305_c31 bl[31] br[31] wl[305] vdd gnd cell_6t
Xbit_r306_c31 bl[31] br[31] wl[306] vdd gnd cell_6t
Xbit_r307_c31 bl[31] br[31] wl[307] vdd gnd cell_6t
Xbit_r308_c31 bl[31] br[31] wl[308] vdd gnd cell_6t
Xbit_r309_c31 bl[31] br[31] wl[309] vdd gnd cell_6t
Xbit_r310_c31 bl[31] br[31] wl[310] vdd gnd cell_6t
Xbit_r311_c31 bl[31] br[31] wl[311] vdd gnd cell_6t
Xbit_r312_c31 bl[31] br[31] wl[312] vdd gnd cell_6t
Xbit_r313_c31 bl[31] br[31] wl[313] vdd gnd cell_6t
Xbit_r314_c31 bl[31] br[31] wl[314] vdd gnd cell_6t
Xbit_r315_c31 bl[31] br[31] wl[315] vdd gnd cell_6t
Xbit_r316_c31 bl[31] br[31] wl[316] vdd gnd cell_6t
Xbit_r317_c31 bl[31] br[31] wl[317] vdd gnd cell_6t
Xbit_r318_c31 bl[31] br[31] wl[318] vdd gnd cell_6t
Xbit_r319_c31 bl[31] br[31] wl[319] vdd gnd cell_6t
Xbit_r320_c31 bl[31] br[31] wl[320] vdd gnd cell_6t
Xbit_r321_c31 bl[31] br[31] wl[321] vdd gnd cell_6t
Xbit_r322_c31 bl[31] br[31] wl[322] vdd gnd cell_6t
Xbit_r323_c31 bl[31] br[31] wl[323] vdd gnd cell_6t
Xbit_r324_c31 bl[31] br[31] wl[324] vdd gnd cell_6t
Xbit_r325_c31 bl[31] br[31] wl[325] vdd gnd cell_6t
Xbit_r326_c31 bl[31] br[31] wl[326] vdd gnd cell_6t
Xbit_r327_c31 bl[31] br[31] wl[327] vdd gnd cell_6t
Xbit_r328_c31 bl[31] br[31] wl[328] vdd gnd cell_6t
Xbit_r329_c31 bl[31] br[31] wl[329] vdd gnd cell_6t
Xbit_r330_c31 bl[31] br[31] wl[330] vdd gnd cell_6t
Xbit_r331_c31 bl[31] br[31] wl[331] vdd gnd cell_6t
Xbit_r332_c31 bl[31] br[31] wl[332] vdd gnd cell_6t
Xbit_r333_c31 bl[31] br[31] wl[333] vdd gnd cell_6t
Xbit_r334_c31 bl[31] br[31] wl[334] vdd gnd cell_6t
Xbit_r335_c31 bl[31] br[31] wl[335] vdd gnd cell_6t
Xbit_r336_c31 bl[31] br[31] wl[336] vdd gnd cell_6t
Xbit_r337_c31 bl[31] br[31] wl[337] vdd gnd cell_6t
Xbit_r338_c31 bl[31] br[31] wl[338] vdd gnd cell_6t
Xbit_r339_c31 bl[31] br[31] wl[339] vdd gnd cell_6t
Xbit_r340_c31 bl[31] br[31] wl[340] vdd gnd cell_6t
Xbit_r341_c31 bl[31] br[31] wl[341] vdd gnd cell_6t
Xbit_r342_c31 bl[31] br[31] wl[342] vdd gnd cell_6t
Xbit_r343_c31 bl[31] br[31] wl[343] vdd gnd cell_6t
Xbit_r344_c31 bl[31] br[31] wl[344] vdd gnd cell_6t
Xbit_r345_c31 bl[31] br[31] wl[345] vdd gnd cell_6t
Xbit_r346_c31 bl[31] br[31] wl[346] vdd gnd cell_6t
Xbit_r347_c31 bl[31] br[31] wl[347] vdd gnd cell_6t
Xbit_r348_c31 bl[31] br[31] wl[348] vdd gnd cell_6t
Xbit_r349_c31 bl[31] br[31] wl[349] vdd gnd cell_6t
Xbit_r350_c31 bl[31] br[31] wl[350] vdd gnd cell_6t
Xbit_r351_c31 bl[31] br[31] wl[351] vdd gnd cell_6t
Xbit_r352_c31 bl[31] br[31] wl[352] vdd gnd cell_6t
Xbit_r353_c31 bl[31] br[31] wl[353] vdd gnd cell_6t
Xbit_r354_c31 bl[31] br[31] wl[354] vdd gnd cell_6t
Xbit_r355_c31 bl[31] br[31] wl[355] vdd gnd cell_6t
Xbit_r356_c31 bl[31] br[31] wl[356] vdd gnd cell_6t
Xbit_r357_c31 bl[31] br[31] wl[357] vdd gnd cell_6t
Xbit_r358_c31 bl[31] br[31] wl[358] vdd gnd cell_6t
Xbit_r359_c31 bl[31] br[31] wl[359] vdd gnd cell_6t
Xbit_r360_c31 bl[31] br[31] wl[360] vdd gnd cell_6t
Xbit_r361_c31 bl[31] br[31] wl[361] vdd gnd cell_6t
Xbit_r362_c31 bl[31] br[31] wl[362] vdd gnd cell_6t
Xbit_r363_c31 bl[31] br[31] wl[363] vdd gnd cell_6t
Xbit_r364_c31 bl[31] br[31] wl[364] vdd gnd cell_6t
Xbit_r365_c31 bl[31] br[31] wl[365] vdd gnd cell_6t
Xbit_r366_c31 bl[31] br[31] wl[366] vdd gnd cell_6t
Xbit_r367_c31 bl[31] br[31] wl[367] vdd gnd cell_6t
Xbit_r368_c31 bl[31] br[31] wl[368] vdd gnd cell_6t
Xbit_r369_c31 bl[31] br[31] wl[369] vdd gnd cell_6t
Xbit_r370_c31 bl[31] br[31] wl[370] vdd gnd cell_6t
Xbit_r371_c31 bl[31] br[31] wl[371] vdd gnd cell_6t
Xbit_r372_c31 bl[31] br[31] wl[372] vdd gnd cell_6t
Xbit_r373_c31 bl[31] br[31] wl[373] vdd gnd cell_6t
Xbit_r374_c31 bl[31] br[31] wl[374] vdd gnd cell_6t
Xbit_r375_c31 bl[31] br[31] wl[375] vdd gnd cell_6t
Xbit_r376_c31 bl[31] br[31] wl[376] vdd gnd cell_6t
Xbit_r377_c31 bl[31] br[31] wl[377] vdd gnd cell_6t
Xbit_r378_c31 bl[31] br[31] wl[378] vdd gnd cell_6t
Xbit_r379_c31 bl[31] br[31] wl[379] vdd gnd cell_6t
Xbit_r380_c31 bl[31] br[31] wl[380] vdd gnd cell_6t
Xbit_r381_c31 bl[31] br[31] wl[381] vdd gnd cell_6t
Xbit_r382_c31 bl[31] br[31] wl[382] vdd gnd cell_6t
Xbit_r383_c31 bl[31] br[31] wl[383] vdd gnd cell_6t
Xbit_r384_c31 bl[31] br[31] wl[384] vdd gnd cell_6t
Xbit_r385_c31 bl[31] br[31] wl[385] vdd gnd cell_6t
Xbit_r386_c31 bl[31] br[31] wl[386] vdd gnd cell_6t
Xbit_r387_c31 bl[31] br[31] wl[387] vdd gnd cell_6t
Xbit_r388_c31 bl[31] br[31] wl[388] vdd gnd cell_6t
Xbit_r389_c31 bl[31] br[31] wl[389] vdd gnd cell_6t
Xbit_r390_c31 bl[31] br[31] wl[390] vdd gnd cell_6t
Xbit_r391_c31 bl[31] br[31] wl[391] vdd gnd cell_6t
Xbit_r392_c31 bl[31] br[31] wl[392] vdd gnd cell_6t
Xbit_r393_c31 bl[31] br[31] wl[393] vdd gnd cell_6t
Xbit_r394_c31 bl[31] br[31] wl[394] vdd gnd cell_6t
Xbit_r395_c31 bl[31] br[31] wl[395] vdd gnd cell_6t
Xbit_r396_c31 bl[31] br[31] wl[396] vdd gnd cell_6t
Xbit_r397_c31 bl[31] br[31] wl[397] vdd gnd cell_6t
Xbit_r398_c31 bl[31] br[31] wl[398] vdd gnd cell_6t
Xbit_r399_c31 bl[31] br[31] wl[399] vdd gnd cell_6t
Xbit_r400_c31 bl[31] br[31] wl[400] vdd gnd cell_6t
Xbit_r401_c31 bl[31] br[31] wl[401] vdd gnd cell_6t
Xbit_r402_c31 bl[31] br[31] wl[402] vdd gnd cell_6t
Xbit_r403_c31 bl[31] br[31] wl[403] vdd gnd cell_6t
Xbit_r404_c31 bl[31] br[31] wl[404] vdd gnd cell_6t
Xbit_r405_c31 bl[31] br[31] wl[405] vdd gnd cell_6t
Xbit_r406_c31 bl[31] br[31] wl[406] vdd gnd cell_6t
Xbit_r407_c31 bl[31] br[31] wl[407] vdd gnd cell_6t
Xbit_r408_c31 bl[31] br[31] wl[408] vdd gnd cell_6t
Xbit_r409_c31 bl[31] br[31] wl[409] vdd gnd cell_6t
Xbit_r410_c31 bl[31] br[31] wl[410] vdd gnd cell_6t
Xbit_r411_c31 bl[31] br[31] wl[411] vdd gnd cell_6t
Xbit_r412_c31 bl[31] br[31] wl[412] vdd gnd cell_6t
Xbit_r413_c31 bl[31] br[31] wl[413] vdd gnd cell_6t
Xbit_r414_c31 bl[31] br[31] wl[414] vdd gnd cell_6t
Xbit_r415_c31 bl[31] br[31] wl[415] vdd gnd cell_6t
Xbit_r416_c31 bl[31] br[31] wl[416] vdd gnd cell_6t
Xbit_r417_c31 bl[31] br[31] wl[417] vdd gnd cell_6t
Xbit_r418_c31 bl[31] br[31] wl[418] vdd gnd cell_6t
Xbit_r419_c31 bl[31] br[31] wl[419] vdd gnd cell_6t
Xbit_r420_c31 bl[31] br[31] wl[420] vdd gnd cell_6t
Xbit_r421_c31 bl[31] br[31] wl[421] vdd gnd cell_6t
Xbit_r422_c31 bl[31] br[31] wl[422] vdd gnd cell_6t
Xbit_r423_c31 bl[31] br[31] wl[423] vdd gnd cell_6t
Xbit_r424_c31 bl[31] br[31] wl[424] vdd gnd cell_6t
Xbit_r425_c31 bl[31] br[31] wl[425] vdd gnd cell_6t
Xbit_r426_c31 bl[31] br[31] wl[426] vdd gnd cell_6t
Xbit_r427_c31 bl[31] br[31] wl[427] vdd gnd cell_6t
Xbit_r428_c31 bl[31] br[31] wl[428] vdd gnd cell_6t
Xbit_r429_c31 bl[31] br[31] wl[429] vdd gnd cell_6t
Xbit_r430_c31 bl[31] br[31] wl[430] vdd gnd cell_6t
Xbit_r431_c31 bl[31] br[31] wl[431] vdd gnd cell_6t
Xbit_r432_c31 bl[31] br[31] wl[432] vdd gnd cell_6t
Xbit_r433_c31 bl[31] br[31] wl[433] vdd gnd cell_6t
Xbit_r434_c31 bl[31] br[31] wl[434] vdd gnd cell_6t
Xbit_r435_c31 bl[31] br[31] wl[435] vdd gnd cell_6t
Xbit_r436_c31 bl[31] br[31] wl[436] vdd gnd cell_6t
Xbit_r437_c31 bl[31] br[31] wl[437] vdd gnd cell_6t
Xbit_r438_c31 bl[31] br[31] wl[438] vdd gnd cell_6t
Xbit_r439_c31 bl[31] br[31] wl[439] vdd gnd cell_6t
Xbit_r440_c31 bl[31] br[31] wl[440] vdd gnd cell_6t
Xbit_r441_c31 bl[31] br[31] wl[441] vdd gnd cell_6t
Xbit_r442_c31 bl[31] br[31] wl[442] vdd gnd cell_6t
Xbit_r443_c31 bl[31] br[31] wl[443] vdd gnd cell_6t
Xbit_r444_c31 bl[31] br[31] wl[444] vdd gnd cell_6t
Xbit_r445_c31 bl[31] br[31] wl[445] vdd gnd cell_6t
Xbit_r446_c31 bl[31] br[31] wl[446] vdd gnd cell_6t
Xbit_r447_c31 bl[31] br[31] wl[447] vdd gnd cell_6t
Xbit_r448_c31 bl[31] br[31] wl[448] vdd gnd cell_6t
Xbit_r449_c31 bl[31] br[31] wl[449] vdd gnd cell_6t
Xbit_r450_c31 bl[31] br[31] wl[450] vdd gnd cell_6t
Xbit_r451_c31 bl[31] br[31] wl[451] vdd gnd cell_6t
Xbit_r452_c31 bl[31] br[31] wl[452] vdd gnd cell_6t
Xbit_r453_c31 bl[31] br[31] wl[453] vdd gnd cell_6t
Xbit_r454_c31 bl[31] br[31] wl[454] vdd gnd cell_6t
Xbit_r455_c31 bl[31] br[31] wl[455] vdd gnd cell_6t
Xbit_r456_c31 bl[31] br[31] wl[456] vdd gnd cell_6t
Xbit_r457_c31 bl[31] br[31] wl[457] vdd gnd cell_6t
Xbit_r458_c31 bl[31] br[31] wl[458] vdd gnd cell_6t
Xbit_r459_c31 bl[31] br[31] wl[459] vdd gnd cell_6t
Xbit_r460_c31 bl[31] br[31] wl[460] vdd gnd cell_6t
Xbit_r461_c31 bl[31] br[31] wl[461] vdd gnd cell_6t
Xbit_r462_c31 bl[31] br[31] wl[462] vdd gnd cell_6t
Xbit_r463_c31 bl[31] br[31] wl[463] vdd gnd cell_6t
Xbit_r464_c31 bl[31] br[31] wl[464] vdd gnd cell_6t
Xbit_r465_c31 bl[31] br[31] wl[465] vdd gnd cell_6t
Xbit_r466_c31 bl[31] br[31] wl[466] vdd gnd cell_6t
Xbit_r467_c31 bl[31] br[31] wl[467] vdd gnd cell_6t
Xbit_r468_c31 bl[31] br[31] wl[468] vdd gnd cell_6t
Xbit_r469_c31 bl[31] br[31] wl[469] vdd gnd cell_6t
Xbit_r470_c31 bl[31] br[31] wl[470] vdd gnd cell_6t
Xbit_r471_c31 bl[31] br[31] wl[471] vdd gnd cell_6t
Xbit_r472_c31 bl[31] br[31] wl[472] vdd gnd cell_6t
Xbit_r473_c31 bl[31] br[31] wl[473] vdd gnd cell_6t
Xbit_r474_c31 bl[31] br[31] wl[474] vdd gnd cell_6t
Xbit_r475_c31 bl[31] br[31] wl[475] vdd gnd cell_6t
Xbit_r476_c31 bl[31] br[31] wl[476] vdd gnd cell_6t
Xbit_r477_c31 bl[31] br[31] wl[477] vdd gnd cell_6t
Xbit_r478_c31 bl[31] br[31] wl[478] vdd gnd cell_6t
Xbit_r479_c31 bl[31] br[31] wl[479] vdd gnd cell_6t
Xbit_r480_c31 bl[31] br[31] wl[480] vdd gnd cell_6t
Xbit_r481_c31 bl[31] br[31] wl[481] vdd gnd cell_6t
Xbit_r482_c31 bl[31] br[31] wl[482] vdd gnd cell_6t
Xbit_r483_c31 bl[31] br[31] wl[483] vdd gnd cell_6t
Xbit_r484_c31 bl[31] br[31] wl[484] vdd gnd cell_6t
Xbit_r485_c31 bl[31] br[31] wl[485] vdd gnd cell_6t
Xbit_r486_c31 bl[31] br[31] wl[486] vdd gnd cell_6t
Xbit_r487_c31 bl[31] br[31] wl[487] vdd gnd cell_6t
Xbit_r488_c31 bl[31] br[31] wl[488] vdd gnd cell_6t
Xbit_r489_c31 bl[31] br[31] wl[489] vdd gnd cell_6t
Xbit_r490_c31 bl[31] br[31] wl[490] vdd gnd cell_6t
Xbit_r491_c31 bl[31] br[31] wl[491] vdd gnd cell_6t
Xbit_r492_c31 bl[31] br[31] wl[492] vdd gnd cell_6t
Xbit_r493_c31 bl[31] br[31] wl[493] vdd gnd cell_6t
Xbit_r494_c31 bl[31] br[31] wl[494] vdd gnd cell_6t
Xbit_r495_c31 bl[31] br[31] wl[495] vdd gnd cell_6t
Xbit_r496_c31 bl[31] br[31] wl[496] vdd gnd cell_6t
Xbit_r497_c31 bl[31] br[31] wl[497] vdd gnd cell_6t
Xbit_r498_c31 bl[31] br[31] wl[498] vdd gnd cell_6t
Xbit_r499_c31 bl[31] br[31] wl[499] vdd gnd cell_6t
Xbit_r500_c31 bl[31] br[31] wl[500] vdd gnd cell_6t
Xbit_r501_c31 bl[31] br[31] wl[501] vdd gnd cell_6t
Xbit_r502_c31 bl[31] br[31] wl[502] vdd gnd cell_6t
Xbit_r503_c31 bl[31] br[31] wl[503] vdd gnd cell_6t
Xbit_r504_c31 bl[31] br[31] wl[504] vdd gnd cell_6t
Xbit_r505_c31 bl[31] br[31] wl[505] vdd gnd cell_6t
Xbit_r506_c31 bl[31] br[31] wl[506] vdd gnd cell_6t
Xbit_r507_c31 bl[31] br[31] wl[507] vdd gnd cell_6t
Xbit_r508_c31 bl[31] br[31] wl[508] vdd gnd cell_6t
Xbit_r509_c31 bl[31] br[31] wl[509] vdd gnd cell_6t
Xbit_r510_c31 bl[31] br[31] wl[510] vdd gnd cell_6t
Xbit_r511_c31 bl[31] br[31] wl[511] vdd gnd cell_6t
Xbit_r0_c32 bl[32] br[32] wl[0] vdd gnd cell_6t
Xbit_r1_c32 bl[32] br[32] wl[1] vdd gnd cell_6t
Xbit_r2_c32 bl[32] br[32] wl[2] vdd gnd cell_6t
Xbit_r3_c32 bl[32] br[32] wl[3] vdd gnd cell_6t
Xbit_r4_c32 bl[32] br[32] wl[4] vdd gnd cell_6t
Xbit_r5_c32 bl[32] br[32] wl[5] vdd gnd cell_6t
Xbit_r6_c32 bl[32] br[32] wl[6] vdd gnd cell_6t
Xbit_r7_c32 bl[32] br[32] wl[7] vdd gnd cell_6t
Xbit_r8_c32 bl[32] br[32] wl[8] vdd gnd cell_6t
Xbit_r9_c32 bl[32] br[32] wl[9] vdd gnd cell_6t
Xbit_r10_c32 bl[32] br[32] wl[10] vdd gnd cell_6t
Xbit_r11_c32 bl[32] br[32] wl[11] vdd gnd cell_6t
Xbit_r12_c32 bl[32] br[32] wl[12] vdd gnd cell_6t
Xbit_r13_c32 bl[32] br[32] wl[13] vdd gnd cell_6t
Xbit_r14_c32 bl[32] br[32] wl[14] vdd gnd cell_6t
Xbit_r15_c32 bl[32] br[32] wl[15] vdd gnd cell_6t
Xbit_r16_c32 bl[32] br[32] wl[16] vdd gnd cell_6t
Xbit_r17_c32 bl[32] br[32] wl[17] vdd gnd cell_6t
Xbit_r18_c32 bl[32] br[32] wl[18] vdd gnd cell_6t
Xbit_r19_c32 bl[32] br[32] wl[19] vdd gnd cell_6t
Xbit_r20_c32 bl[32] br[32] wl[20] vdd gnd cell_6t
Xbit_r21_c32 bl[32] br[32] wl[21] vdd gnd cell_6t
Xbit_r22_c32 bl[32] br[32] wl[22] vdd gnd cell_6t
Xbit_r23_c32 bl[32] br[32] wl[23] vdd gnd cell_6t
Xbit_r24_c32 bl[32] br[32] wl[24] vdd gnd cell_6t
Xbit_r25_c32 bl[32] br[32] wl[25] vdd gnd cell_6t
Xbit_r26_c32 bl[32] br[32] wl[26] vdd gnd cell_6t
Xbit_r27_c32 bl[32] br[32] wl[27] vdd gnd cell_6t
Xbit_r28_c32 bl[32] br[32] wl[28] vdd gnd cell_6t
Xbit_r29_c32 bl[32] br[32] wl[29] vdd gnd cell_6t
Xbit_r30_c32 bl[32] br[32] wl[30] vdd gnd cell_6t
Xbit_r31_c32 bl[32] br[32] wl[31] vdd gnd cell_6t
Xbit_r32_c32 bl[32] br[32] wl[32] vdd gnd cell_6t
Xbit_r33_c32 bl[32] br[32] wl[33] vdd gnd cell_6t
Xbit_r34_c32 bl[32] br[32] wl[34] vdd gnd cell_6t
Xbit_r35_c32 bl[32] br[32] wl[35] vdd gnd cell_6t
Xbit_r36_c32 bl[32] br[32] wl[36] vdd gnd cell_6t
Xbit_r37_c32 bl[32] br[32] wl[37] vdd gnd cell_6t
Xbit_r38_c32 bl[32] br[32] wl[38] vdd gnd cell_6t
Xbit_r39_c32 bl[32] br[32] wl[39] vdd gnd cell_6t
Xbit_r40_c32 bl[32] br[32] wl[40] vdd gnd cell_6t
Xbit_r41_c32 bl[32] br[32] wl[41] vdd gnd cell_6t
Xbit_r42_c32 bl[32] br[32] wl[42] vdd gnd cell_6t
Xbit_r43_c32 bl[32] br[32] wl[43] vdd gnd cell_6t
Xbit_r44_c32 bl[32] br[32] wl[44] vdd gnd cell_6t
Xbit_r45_c32 bl[32] br[32] wl[45] vdd gnd cell_6t
Xbit_r46_c32 bl[32] br[32] wl[46] vdd gnd cell_6t
Xbit_r47_c32 bl[32] br[32] wl[47] vdd gnd cell_6t
Xbit_r48_c32 bl[32] br[32] wl[48] vdd gnd cell_6t
Xbit_r49_c32 bl[32] br[32] wl[49] vdd gnd cell_6t
Xbit_r50_c32 bl[32] br[32] wl[50] vdd gnd cell_6t
Xbit_r51_c32 bl[32] br[32] wl[51] vdd gnd cell_6t
Xbit_r52_c32 bl[32] br[32] wl[52] vdd gnd cell_6t
Xbit_r53_c32 bl[32] br[32] wl[53] vdd gnd cell_6t
Xbit_r54_c32 bl[32] br[32] wl[54] vdd gnd cell_6t
Xbit_r55_c32 bl[32] br[32] wl[55] vdd gnd cell_6t
Xbit_r56_c32 bl[32] br[32] wl[56] vdd gnd cell_6t
Xbit_r57_c32 bl[32] br[32] wl[57] vdd gnd cell_6t
Xbit_r58_c32 bl[32] br[32] wl[58] vdd gnd cell_6t
Xbit_r59_c32 bl[32] br[32] wl[59] vdd gnd cell_6t
Xbit_r60_c32 bl[32] br[32] wl[60] vdd gnd cell_6t
Xbit_r61_c32 bl[32] br[32] wl[61] vdd gnd cell_6t
Xbit_r62_c32 bl[32] br[32] wl[62] vdd gnd cell_6t
Xbit_r63_c32 bl[32] br[32] wl[63] vdd gnd cell_6t
Xbit_r64_c32 bl[32] br[32] wl[64] vdd gnd cell_6t
Xbit_r65_c32 bl[32] br[32] wl[65] vdd gnd cell_6t
Xbit_r66_c32 bl[32] br[32] wl[66] vdd gnd cell_6t
Xbit_r67_c32 bl[32] br[32] wl[67] vdd gnd cell_6t
Xbit_r68_c32 bl[32] br[32] wl[68] vdd gnd cell_6t
Xbit_r69_c32 bl[32] br[32] wl[69] vdd gnd cell_6t
Xbit_r70_c32 bl[32] br[32] wl[70] vdd gnd cell_6t
Xbit_r71_c32 bl[32] br[32] wl[71] vdd gnd cell_6t
Xbit_r72_c32 bl[32] br[32] wl[72] vdd gnd cell_6t
Xbit_r73_c32 bl[32] br[32] wl[73] vdd gnd cell_6t
Xbit_r74_c32 bl[32] br[32] wl[74] vdd gnd cell_6t
Xbit_r75_c32 bl[32] br[32] wl[75] vdd gnd cell_6t
Xbit_r76_c32 bl[32] br[32] wl[76] vdd gnd cell_6t
Xbit_r77_c32 bl[32] br[32] wl[77] vdd gnd cell_6t
Xbit_r78_c32 bl[32] br[32] wl[78] vdd gnd cell_6t
Xbit_r79_c32 bl[32] br[32] wl[79] vdd gnd cell_6t
Xbit_r80_c32 bl[32] br[32] wl[80] vdd gnd cell_6t
Xbit_r81_c32 bl[32] br[32] wl[81] vdd gnd cell_6t
Xbit_r82_c32 bl[32] br[32] wl[82] vdd gnd cell_6t
Xbit_r83_c32 bl[32] br[32] wl[83] vdd gnd cell_6t
Xbit_r84_c32 bl[32] br[32] wl[84] vdd gnd cell_6t
Xbit_r85_c32 bl[32] br[32] wl[85] vdd gnd cell_6t
Xbit_r86_c32 bl[32] br[32] wl[86] vdd gnd cell_6t
Xbit_r87_c32 bl[32] br[32] wl[87] vdd gnd cell_6t
Xbit_r88_c32 bl[32] br[32] wl[88] vdd gnd cell_6t
Xbit_r89_c32 bl[32] br[32] wl[89] vdd gnd cell_6t
Xbit_r90_c32 bl[32] br[32] wl[90] vdd gnd cell_6t
Xbit_r91_c32 bl[32] br[32] wl[91] vdd gnd cell_6t
Xbit_r92_c32 bl[32] br[32] wl[92] vdd gnd cell_6t
Xbit_r93_c32 bl[32] br[32] wl[93] vdd gnd cell_6t
Xbit_r94_c32 bl[32] br[32] wl[94] vdd gnd cell_6t
Xbit_r95_c32 bl[32] br[32] wl[95] vdd gnd cell_6t
Xbit_r96_c32 bl[32] br[32] wl[96] vdd gnd cell_6t
Xbit_r97_c32 bl[32] br[32] wl[97] vdd gnd cell_6t
Xbit_r98_c32 bl[32] br[32] wl[98] vdd gnd cell_6t
Xbit_r99_c32 bl[32] br[32] wl[99] vdd gnd cell_6t
Xbit_r100_c32 bl[32] br[32] wl[100] vdd gnd cell_6t
Xbit_r101_c32 bl[32] br[32] wl[101] vdd gnd cell_6t
Xbit_r102_c32 bl[32] br[32] wl[102] vdd gnd cell_6t
Xbit_r103_c32 bl[32] br[32] wl[103] vdd gnd cell_6t
Xbit_r104_c32 bl[32] br[32] wl[104] vdd gnd cell_6t
Xbit_r105_c32 bl[32] br[32] wl[105] vdd gnd cell_6t
Xbit_r106_c32 bl[32] br[32] wl[106] vdd gnd cell_6t
Xbit_r107_c32 bl[32] br[32] wl[107] vdd gnd cell_6t
Xbit_r108_c32 bl[32] br[32] wl[108] vdd gnd cell_6t
Xbit_r109_c32 bl[32] br[32] wl[109] vdd gnd cell_6t
Xbit_r110_c32 bl[32] br[32] wl[110] vdd gnd cell_6t
Xbit_r111_c32 bl[32] br[32] wl[111] vdd gnd cell_6t
Xbit_r112_c32 bl[32] br[32] wl[112] vdd gnd cell_6t
Xbit_r113_c32 bl[32] br[32] wl[113] vdd gnd cell_6t
Xbit_r114_c32 bl[32] br[32] wl[114] vdd gnd cell_6t
Xbit_r115_c32 bl[32] br[32] wl[115] vdd gnd cell_6t
Xbit_r116_c32 bl[32] br[32] wl[116] vdd gnd cell_6t
Xbit_r117_c32 bl[32] br[32] wl[117] vdd gnd cell_6t
Xbit_r118_c32 bl[32] br[32] wl[118] vdd gnd cell_6t
Xbit_r119_c32 bl[32] br[32] wl[119] vdd gnd cell_6t
Xbit_r120_c32 bl[32] br[32] wl[120] vdd gnd cell_6t
Xbit_r121_c32 bl[32] br[32] wl[121] vdd gnd cell_6t
Xbit_r122_c32 bl[32] br[32] wl[122] vdd gnd cell_6t
Xbit_r123_c32 bl[32] br[32] wl[123] vdd gnd cell_6t
Xbit_r124_c32 bl[32] br[32] wl[124] vdd gnd cell_6t
Xbit_r125_c32 bl[32] br[32] wl[125] vdd gnd cell_6t
Xbit_r126_c32 bl[32] br[32] wl[126] vdd gnd cell_6t
Xbit_r127_c32 bl[32] br[32] wl[127] vdd gnd cell_6t
Xbit_r128_c32 bl[32] br[32] wl[128] vdd gnd cell_6t
Xbit_r129_c32 bl[32] br[32] wl[129] vdd gnd cell_6t
Xbit_r130_c32 bl[32] br[32] wl[130] vdd gnd cell_6t
Xbit_r131_c32 bl[32] br[32] wl[131] vdd gnd cell_6t
Xbit_r132_c32 bl[32] br[32] wl[132] vdd gnd cell_6t
Xbit_r133_c32 bl[32] br[32] wl[133] vdd gnd cell_6t
Xbit_r134_c32 bl[32] br[32] wl[134] vdd gnd cell_6t
Xbit_r135_c32 bl[32] br[32] wl[135] vdd gnd cell_6t
Xbit_r136_c32 bl[32] br[32] wl[136] vdd gnd cell_6t
Xbit_r137_c32 bl[32] br[32] wl[137] vdd gnd cell_6t
Xbit_r138_c32 bl[32] br[32] wl[138] vdd gnd cell_6t
Xbit_r139_c32 bl[32] br[32] wl[139] vdd gnd cell_6t
Xbit_r140_c32 bl[32] br[32] wl[140] vdd gnd cell_6t
Xbit_r141_c32 bl[32] br[32] wl[141] vdd gnd cell_6t
Xbit_r142_c32 bl[32] br[32] wl[142] vdd gnd cell_6t
Xbit_r143_c32 bl[32] br[32] wl[143] vdd gnd cell_6t
Xbit_r144_c32 bl[32] br[32] wl[144] vdd gnd cell_6t
Xbit_r145_c32 bl[32] br[32] wl[145] vdd gnd cell_6t
Xbit_r146_c32 bl[32] br[32] wl[146] vdd gnd cell_6t
Xbit_r147_c32 bl[32] br[32] wl[147] vdd gnd cell_6t
Xbit_r148_c32 bl[32] br[32] wl[148] vdd gnd cell_6t
Xbit_r149_c32 bl[32] br[32] wl[149] vdd gnd cell_6t
Xbit_r150_c32 bl[32] br[32] wl[150] vdd gnd cell_6t
Xbit_r151_c32 bl[32] br[32] wl[151] vdd gnd cell_6t
Xbit_r152_c32 bl[32] br[32] wl[152] vdd gnd cell_6t
Xbit_r153_c32 bl[32] br[32] wl[153] vdd gnd cell_6t
Xbit_r154_c32 bl[32] br[32] wl[154] vdd gnd cell_6t
Xbit_r155_c32 bl[32] br[32] wl[155] vdd gnd cell_6t
Xbit_r156_c32 bl[32] br[32] wl[156] vdd gnd cell_6t
Xbit_r157_c32 bl[32] br[32] wl[157] vdd gnd cell_6t
Xbit_r158_c32 bl[32] br[32] wl[158] vdd gnd cell_6t
Xbit_r159_c32 bl[32] br[32] wl[159] vdd gnd cell_6t
Xbit_r160_c32 bl[32] br[32] wl[160] vdd gnd cell_6t
Xbit_r161_c32 bl[32] br[32] wl[161] vdd gnd cell_6t
Xbit_r162_c32 bl[32] br[32] wl[162] vdd gnd cell_6t
Xbit_r163_c32 bl[32] br[32] wl[163] vdd gnd cell_6t
Xbit_r164_c32 bl[32] br[32] wl[164] vdd gnd cell_6t
Xbit_r165_c32 bl[32] br[32] wl[165] vdd gnd cell_6t
Xbit_r166_c32 bl[32] br[32] wl[166] vdd gnd cell_6t
Xbit_r167_c32 bl[32] br[32] wl[167] vdd gnd cell_6t
Xbit_r168_c32 bl[32] br[32] wl[168] vdd gnd cell_6t
Xbit_r169_c32 bl[32] br[32] wl[169] vdd gnd cell_6t
Xbit_r170_c32 bl[32] br[32] wl[170] vdd gnd cell_6t
Xbit_r171_c32 bl[32] br[32] wl[171] vdd gnd cell_6t
Xbit_r172_c32 bl[32] br[32] wl[172] vdd gnd cell_6t
Xbit_r173_c32 bl[32] br[32] wl[173] vdd gnd cell_6t
Xbit_r174_c32 bl[32] br[32] wl[174] vdd gnd cell_6t
Xbit_r175_c32 bl[32] br[32] wl[175] vdd gnd cell_6t
Xbit_r176_c32 bl[32] br[32] wl[176] vdd gnd cell_6t
Xbit_r177_c32 bl[32] br[32] wl[177] vdd gnd cell_6t
Xbit_r178_c32 bl[32] br[32] wl[178] vdd gnd cell_6t
Xbit_r179_c32 bl[32] br[32] wl[179] vdd gnd cell_6t
Xbit_r180_c32 bl[32] br[32] wl[180] vdd gnd cell_6t
Xbit_r181_c32 bl[32] br[32] wl[181] vdd gnd cell_6t
Xbit_r182_c32 bl[32] br[32] wl[182] vdd gnd cell_6t
Xbit_r183_c32 bl[32] br[32] wl[183] vdd gnd cell_6t
Xbit_r184_c32 bl[32] br[32] wl[184] vdd gnd cell_6t
Xbit_r185_c32 bl[32] br[32] wl[185] vdd gnd cell_6t
Xbit_r186_c32 bl[32] br[32] wl[186] vdd gnd cell_6t
Xbit_r187_c32 bl[32] br[32] wl[187] vdd gnd cell_6t
Xbit_r188_c32 bl[32] br[32] wl[188] vdd gnd cell_6t
Xbit_r189_c32 bl[32] br[32] wl[189] vdd gnd cell_6t
Xbit_r190_c32 bl[32] br[32] wl[190] vdd gnd cell_6t
Xbit_r191_c32 bl[32] br[32] wl[191] vdd gnd cell_6t
Xbit_r192_c32 bl[32] br[32] wl[192] vdd gnd cell_6t
Xbit_r193_c32 bl[32] br[32] wl[193] vdd gnd cell_6t
Xbit_r194_c32 bl[32] br[32] wl[194] vdd gnd cell_6t
Xbit_r195_c32 bl[32] br[32] wl[195] vdd gnd cell_6t
Xbit_r196_c32 bl[32] br[32] wl[196] vdd gnd cell_6t
Xbit_r197_c32 bl[32] br[32] wl[197] vdd gnd cell_6t
Xbit_r198_c32 bl[32] br[32] wl[198] vdd gnd cell_6t
Xbit_r199_c32 bl[32] br[32] wl[199] vdd gnd cell_6t
Xbit_r200_c32 bl[32] br[32] wl[200] vdd gnd cell_6t
Xbit_r201_c32 bl[32] br[32] wl[201] vdd gnd cell_6t
Xbit_r202_c32 bl[32] br[32] wl[202] vdd gnd cell_6t
Xbit_r203_c32 bl[32] br[32] wl[203] vdd gnd cell_6t
Xbit_r204_c32 bl[32] br[32] wl[204] vdd gnd cell_6t
Xbit_r205_c32 bl[32] br[32] wl[205] vdd gnd cell_6t
Xbit_r206_c32 bl[32] br[32] wl[206] vdd gnd cell_6t
Xbit_r207_c32 bl[32] br[32] wl[207] vdd gnd cell_6t
Xbit_r208_c32 bl[32] br[32] wl[208] vdd gnd cell_6t
Xbit_r209_c32 bl[32] br[32] wl[209] vdd gnd cell_6t
Xbit_r210_c32 bl[32] br[32] wl[210] vdd gnd cell_6t
Xbit_r211_c32 bl[32] br[32] wl[211] vdd gnd cell_6t
Xbit_r212_c32 bl[32] br[32] wl[212] vdd gnd cell_6t
Xbit_r213_c32 bl[32] br[32] wl[213] vdd gnd cell_6t
Xbit_r214_c32 bl[32] br[32] wl[214] vdd gnd cell_6t
Xbit_r215_c32 bl[32] br[32] wl[215] vdd gnd cell_6t
Xbit_r216_c32 bl[32] br[32] wl[216] vdd gnd cell_6t
Xbit_r217_c32 bl[32] br[32] wl[217] vdd gnd cell_6t
Xbit_r218_c32 bl[32] br[32] wl[218] vdd gnd cell_6t
Xbit_r219_c32 bl[32] br[32] wl[219] vdd gnd cell_6t
Xbit_r220_c32 bl[32] br[32] wl[220] vdd gnd cell_6t
Xbit_r221_c32 bl[32] br[32] wl[221] vdd gnd cell_6t
Xbit_r222_c32 bl[32] br[32] wl[222] vdd gnd cell_6t
Xbit_r223_c32 bl[32] br[32] wl[223] vdd gnd cell_6t
Xbit_r224_c32 bl[32] br[32] wl[224] vdd gnd cell_6t
Xbit_r225_c32 bl[32] br[32] wl[225] vdd gnd cell_6t
Xbit_r226_c32 bl[32] br[32] wl[226] vdd gnd cell_6t
Xbit_r227_c32 bl[32] br[32] wl[227] vdd gnd cell_6t
Xbit_r228_c32 bl[32] br[32] wl[228] vdd gnd cell_6t
Xbit_r229_c32 bl[32] br[32] wl[229] vdd gnd cell_6t
Xbit_r230_c32 bl[32] br[32] wl[230] vdd gnd cell_6t
Xbit_r231_c32 bl[32] br[32] wl[231] vdd gnd cell_6t
Xbit_r232_c32 bl[32] br[32] wl[232] vdd gnd cell_6t
Xbit_r233_c32 bl[32] br[32] wl[233] vdd gnd cell_6t
Xbit_r234_c32 bl[32] br[32] wl[234] vdd gnd cell_6t
Xbit_r235_c32 bl[32] br[32] wl[235] vdd gnd cell_6t
Xbit_r236_c32 bl[32] br[32] wl[236] vdd gnd cell_6t
Xbit_r237_c32 bl[32] br[32] wl[237] vdd gnd cell_6t
Xbit_r238_c32 bl[32] br[32] wl[238] vdd gnd cell_6t
Xbit_r239_c32 bl[32] br[32] wl[239] vdd gnd cell_6t
Xbit_r240_c32 bl[32] br[32] wl[240] vdd gnd cell_6t
Xbit_r241_c32 bl[32] br[32] wl[241] vdd gnd cell_6t
Xbit_r242_c32 bl[32] br[32] wl[242] vdd gnd cell_6t
Xbit_r243_c32 bl[32] br[32] wl[243] vdd gnd cell_6t
Xbit_r244_c32 bl[32] br[32] wl[244] vdd gnd cell_6t
Xbit_r245_c32 bl[32] br[32] wl[245] vdd gnd cell_6t
Xbit_r246_c32 bl[32] br[32] wl[246] vdd gnd cell_6t
Xbit_r247_c32 bl[32] br[32] wl[247] vdd gnd cell_6t
Xbit_r248_c32 bl[32] br[32] wl[248] vdd gnd cell_6t
Xbit_r249_c32 bl[32] br[32] wl[249] vdd gnd cell_6t
Xbit_r250_c32 bl[32] br[32] wl[250] vdd gnd cell_6t
Xbit_r251_c32 bl[32] br[32] wl[251] vdd gnd cell_6t
Xbit_r252_c32 bl[32] br[32] wl[252] vdd gnd cell_6t
Xbit_r253_c32 bl[32] br[32] wl[253] vdd gnd cell_6t
Xbit_r254_c32 bl[32] br[32] wl[254] vdd gnd cell_6t
Xbit_r255_c32 bl[32] br[32] wl[255] vdd gnd cell_6t
Xbit_r256_c32 bl[32] br[32] wl[256] vdd gnd cell_6t
Xbit_r257_c32 bl[32] br[32] wl[257] vdd gnd cell_6t
Xbit_r258_c32 bl[32] br[32] wl[258] vdd gnd cell_6t
Xbit_r259_c32 bl[32] br[32] wl[259] vdd gnd cell_6t
Xbit_r260_c32 bl[32] br[32] wl[260] vdd gnd cell_6t
Xbit_r261_c32 bl[32] br[32] wl[261] vdd gnd cell_6t
Xbit_r262_c32 bl[32] br[32] wl[262] vdd gnd cell_6t
Xbit_r263_c32 bl[32] br[32] wl[263] vdd gnd cell_6t
Xbit_r264_c32 bl[32] br[32] wl[264] vdd gnd cell_6t
Xbit_r265_c32 bl[32] br[32] wl[265] vdd gnd cell_6t
Xbit_r266_c32 bl[32] br[32] wl[266] vdd gnd cell_6t
Xbit_r267_c32 bl[32] br[32] wl[267] vdd gnd cell_6t
Xbit_r268_c32 bl[32] br[32] wl[268] vdd gnd cell_6t
Xbit_r269_c32 bl[32] br[32] wl[269] vdd gnd cell_6t
Xbit_r270_c32 bl[32] br[32] wl[270] vdd gnd cell_6t
Xbit_r271_c32 bl[32] br[32] wl[271] vdd gnd cell_6t
Xbit_r272_c32 bl[32] br[32] wl[272] vdd gnd cell_6t
Xbit_r273_c32 bl[32] br[32] wl[273] vdd gnd cell_6t
Xbit_r274_c32 bl[32] br[32] wl[274] vdd gnd cell_6t
Xbit_r275_c32 bl[32] br[32] wl[275] vdd gnd cell_6t
Xbit_r276_c32 bl[32] br[32] wl[276] vdd gnd cell_6t
Xbit_r277_c32 bl[32] br[32] wl[277] vdd gnd cell_6t
Xbit_r278_c32 bl[32] br[32] wl[278] vdd gnd cell_6t
Xbit_r279_c32 bl[32] br[32] wl[279] vdd gnd cell_6t
Xbit_r280_c32 bl[32] br[32] wl[280] vdd gnd cell_6t
Xbit_r281_c32 bl[32] br[32] wl[281] vdd gnd cell_6t
Xbit_r282_c32 bl[32] br[32] wl[282] vdd gnd cell_6t
Xbit_r283_c32 bl[32] br[32] wl[283] vdd gnd cell_6t
Xbit_r284_c32 bl[32] br[32] wl[284] vdd gnd cell_6t
Xbit_r285_c32 bl[32] br[32] wl[285] vdd gnd cell_6t
Xbit_r286_c32 bl[32] br[32] wl[286] vdd gnd cell_6t
Xbit_r287_c32 bl[32] br[32] wl[287] vdd gnd cell_6t
Xbit_r288_c32 bl[32] br[32] wl[288] vdd gnd cell_6t
Xbit_r289_c32 bl[32] br[32] wl[289] vdd gnd cell_6t
Xbit_r290_c32 bl[32] br[32] wl[290] vdd gnd cell_6t
Xbit_r291_c32 bl[32] br[32] wl[291] vdd gnd cell_6t
Xbit_r292_c32 bl[32] br[32] wl[292] vdd gnd cell_6t
Xbit_r293_c32 bl[32] br[32] wl[293] vdd gnd cell_6t
Xbit_r294_c32 bl[32] br[32] wl[294] vdd gnd cell_6t
Xbit_r295_c32 bl[32] br[32] wl[295] vdd gnd cell_6t
Xbit_r296_c32 bl[32] br[32] wl[296] vdd gnd cell_6t
Xbit_r297_c32 bl[32] br[32] wl[297] vdd gnd cell_6t
Xbit_r298_c32 bl[32] br[32] wl[298] vdd gnd cell_6t
Xbit_r299_c32 bl[32] br[32] wl[299] vdd gnd cell_6t
Xbit_r300_c32 bl[32] br[32] wl[300] vdd gnd cell_6t
Xbit_r301_c32 bl[32] br[32] wl[301] vdd gnd cell_6t
Xbit_r302_c32 bl[32] br[32] wl[302] vdd gnd cell_6t
Xbit_r303_c32 bl[32] br[32] wl[303] vdd gnd cell_6t
Xbit_r304_c32 bl[32] br[32] wl[304] vdd gnd cell_6t
Xbit_r305_c32 bl[32] br[32] wl[305] vdd gnd cell_6t
Xbit_r306_c32 bl[32] br[32] wl[306] vdd gnd cell_6t
Xbit_r307_c32 bl[32] br[32] wl[307] vdd gnd cell_6t
Xbit_r308_c32 bl[32] br[32] wl[308] vdd gnd cell_6t
Xbit_r309_c32 bl[32] br[32] wl[309] vdd gnd cell_6t
Xbit_r310_c32 bl[32] br[32] wl[310] vdd gnd cell_6t
Xbit_r311_c32 bl[32] br[32] wl[311] vdd gnd cell_6t
Xbit_r312_c32 bl[32] br[32] wl[312] vdd gnd cell_6t
Xbit_r313_c32 bl[32] br[32] wl[313] vdd gnd cell_6t
Xbit_r314_c32 bl[32] br[32] wl[314] vdd gnd cell_6t
Xbit_r315_c32 bl[32] br[32] wl[315] vdd gnd cell_6t
Xbit_r316_c32 bl[32] br[32] wl[316] vdd gnd cell_6t
Xbit_r317_c32 bl[32] br[32] wl[317] vdd gnd cell_6t
Xbit_r318_c32 bl[32] br[32] wl[318] vdd gnd cell_6t
Xbit_r319_c32 bl[32] br[32] wl[319] vdd gnd cell_6t
Xbit_r320_c32 bl[32] br[32] wl[320] vdd gnd cell_6t
Xbit_r321_c32 bl[32] br[32] wl[321] vdd gnd cell_6t
Xbit_r322_c32 bl[32] br[32] wl[322] vdd gnd cell_6t
Xbit_r323_c32 bl[32] br[32] wl[323] vdd gnd cell_6t
Xbit_r324_c32 bl[32] br[32] wl[324] vdd gnd cell_6t
Xbit_r325_c32 bl[32] br[32] wl[325] vdd gnd cell_6t
Xbit_r326_c32 bl[32] br[32] wl[326] vdd gnd cell_6t
Xbit_r327_c32 bl[32] br[32] wl[327] vdd gnd cell_6t
Xbit_r328_c32 bl[32] br[32] wl[328] vdd gnd cell_6t
Xbit_r329_c32 bl[32] br[32] wl[329] vdd gnd cell_6t
Xbit_r330_c32 bl[32] br[32] wl[330] vdd gnd cell_6t
Xbit_r331_c32 bl[32] br[32] wl[331] vdd gnd cell_6t
Xbit_r332_c32 bl[32] br[32] wl[332] vdd gnd cell_6t
Xbit_r333_c32 bl[32] br[32] wl[333] vdd gnd cell_6t
Xbit_r334_c32 bl[32] br[32] wl[334] vdd gnd cell_6t
Xbit_r335_c32 bl[32] br[32] wl[335] vdd gnd cell_6t
Xbit_r336_c32 bl[32] br[32] wl[336] vdd gnd cell_6t
Xbit_r337_c32 bl[32] br[32] wl[337] vdd gnd cell_6t
Xbit_r338_c32 bl[32] br[32] wl[338] vdd gnd cell_6t
Xbit_r339_c32 bl[32] br[32] wl[339] vdd gnd cell_6t
Xbit_r340_c32 bl[32] br[32] wl[340] vdd gnd cell_6t
Xbit_r341_c32 bl[32] br[32] wl[341] vdd gnd cell_6t
Xbit_r342_c32 bl[32] br[32] wl[342] vdd gnd cell_6t
Xbit_r343_c32 bl[32] br[32] wl[343] vdd gnd cell_6t
Xbit_r344_c32 bl[32] br[32] wl[344] vdd gnd cell_6t
Xbit_r345_c32 bl[32] br[32] wl[345] vdd gnd cell_6t
Xbit_r346_c32 bl[32] br[32] wl[346] vdd gnd cell_6t
Xbit_r347_c32 bl[32] br[32] wl[347] vdd gnd cell_6t
Xbit_r348_c32 bl[32] br[32] wl[348] vdd gnd cell_6t
Xbit_r349_c32 bl[32] br[32] wl[349] vdd gnd cell_6t
Xbit_r350_c32 bl[32] br[32] wl[350] vdd gnd cell_6t
Xbit_r351_c32 bl[32] br[32] wl[351] vdd gnd cell_6t
Xbit_r352_c32 bl[32] br[32] wl[352] vdd gnd cell_6t
Xbit_r353_c32 bl[32] br[32] wl[353] vdd gnd cell_6t
Xbit_r354_c32 bl[32] br[32] wl[354] vdd gnd cell_6t
Xbit_r355_c32 bl[32] br[32] wl[355] vdd gnd cell_6t
Xbit_r356_c32 bl[32] br[32] wl[356] vdd gnd cell_6t
Xbit_r357_c32 bl[32] br[32] wl[357] vdd gnd cell_6t
Xbit_r358_c32 bl[32] br[32] wl[358] vdd gnd cell_6t
Xbit_r359_c32 bl[32] br[32] wl[359] vdd gnd cell_6t
Xbit_r360_c32 bl[32] br[32] wl[360] vdd gnd cell_6t
Xbit_r361_c32 bl[32] br[32] wl[361] vdd gnd cell_6t
Xbit_r362_c32 bl[32] br[32] wl[362] vdd gnd cell_6t
Xbit_r363_c32 bl[32] br[32] wl[363] vdd gnd cell_6t
Xbit_r364_c32 bl[32] br[32] wl[364] vdd gnd cell_6t
Xbit_r365_c32 bl[32] br[32] wl[365] vdd gnd cell_6t
Xbit_r366_c32 bl[32] br[32] wl[366] vdd gnd cell_6t
Xbit_r367_c32 bl[32] br[32] wl[367] vdd gnd cell_6t
Xbit_r368_c32 bl[32] br[32] wl[368] vdd gnd cell_6t
Xbit_r369_c32 bl[32] br[32] wl[369] vdd gnd cell_6t
Xbit_r370_c32 bl[32] br[32] wl[370] vdd gnd cell_6t
Xbit_r371_c32 bl[32] br[32] wl[371] vdd gnd cell_6t
Xbit_r372_c32 bl[32] br[32] wl[372] vdd gnd cell_6t
Xbit_r373_c32 bl[32] br[32] wl[373] vdd gnd cell_6t
Xbit_r374_c32 bl[32] br[32] wl[374] vdd gnd cell_6t
Xbit_r375_c32 bl[32] br[32] wl[375] vdd gnd cell_6t
Xbit_r376_c32 bl[32] br[32] wl[376] vdd gnd cell_6t
Xbit_r377_c32 bl[32] br[32] wl[377] vdd gnd cell_6t
Xbit_r378_c32 bl[32] br[32] wl[378] vdd gnd cell_6t
Xbit_r379_c32 bl[32] br[32] wl[379] vdd gnd cell_6t
Xbit_r380_c32 bl[32] br[32] wl[380] vdd gnd cell_6t
Xbit_r381_c32 bl[32] br[32] wl[381] vdd gnd cell_6t
Xbit_r382_c32 bl[32] br[32] wl[382] vdd gnd cell_6t
Xbit_r383_c32 bl[32] br[32] wl[383] vdd gnd cell_6t
Xbit_r384_c32 bl[32] br[32] wl[384] vdd gnd cell_6t
Xbit_r385_c32 bl[32] br[32] wl[385] vdd gnd cell_6t
Xbit_r386_c32 bl[32] br[32] wl[386] vdd gnd cell_6t
Xbit_r387_c32 bl[32] br[32] wl[387] vdd gnd cell_6t
Xbit_r388_c32 bl[32] br[32] wl[388] vdd gnd cell_6t
Xbit_r389_c32 bl[32] br[32] wl[389] vdd gnd cell_6t
Xbit_r390_c32 bl[32] br[32] wl[390] vdd gnd cell_6t
Xbit_r391_c32 bl[32] br[32] wl[391] vdd gnd cell_6t
Xbit_r392_c32 bl[32] br[32] wl[392] vdd gnd cell_6t
Xbit_r393_c32 bl[32] br[32] wl[393] vdd gnd cell_6t
Xbit_r394_c32 bl[32] br[32] wl[394] vdd gnd cell_6t
Xbit_r395_c32 bl[32] br[32] wl[395] vdd gnd cell_6t
Xbit_r396_c32 bl[32] br[32] wl[396] vdd gnd cell_6t
Xbit_r397_c32 bl[32] br[32] wl[397] vdd gnd cell_6t
Xbit_r398_c32 bl[32] br[32] wl[398] vdd gnd cell_6t
Xbit_r399_c32 bl[32] br[32] wl[399] vdd gnd cell_6t
Xbit_r400_c32 bl[32] br[32] wl[400] vdd gnd cell_6t
Xbit_r401_c32 bl[32] br[32] wl[401] vdd gnd cell_6t
Xbit_r402_c32 bl[32] br[32] wl[402] vdd gnd cell_6t
Xbit_r403_c32 bl[32] br[32] wl[403] vdd gnd cell_6t
Xbit_r404_c32 bl[32] br[32] wl[404] vdd gnd cell_6t
Xbit_r405_c32 bl[32] br[32] wl[405] vdd gnd cell_6t
Xbit_r406_c32 bl[32] br[32] wl[406] vdd gnd cell_6t
Xbit_r407_c32 bl[32] br[32] wl[407] vdd gnd cell_6t
Xbit_r408_c32 bl[32] br[32] wl[408] vdd gnd cell_6t
Xbit_r409_c32 bl[32] br[32] wl[409] vdd gnd cell_6t
Xbit_r410_c32 bl[32] br[32] wl[410] vdd gnd cell_6t
Xbit_r411_c32 bl[32] br[32] wl[411] vdd gnd cell_6t
Xbit_r412_c32 bl[32] br[32] wl[412] vdd gnd cell_6t
Xbit_r413_c32 bl[32] br[32] wl[413] vdd gnd cell_6t
Xbit_r414_c32 bl[32] br[32] wl[414] vdd gnd cell_6t
Xbit_r415_c32 bl[32] br[32] wl[415] vdd gnd cell_6t
Xbit_r416_c32 bl[32] br[32] wl[416] vdd gnd cell_6t
Xbit_r417_c32 bl[32] br[32] wl[417] vdd gnd cell_6t
Xbit_r418_c32 bl[32] br[32] wl[418] vdd gnd cell_6t
Xbit_r419_c32 bl[32] br[32] wl[419] vdd gnd cell_6t
Xbit_r420_c32 bl[32] br[32] wl[420] vdd gnd cell_6t
Xbit_r421_c32 bl[32] br[32] wl[421] vdd gnd cell_6t
Xbit_r422_c32 bl[32] br[32] wl[422] vdd gnd cell_6t
Xbit_r423_c32 bl[32] br[32] wl[423] vdd gnd cell_6t
Xbit_r424_c32 bl[32] br[32] wl[424] vdd gnd cell_6t
Xbit_r425_c32 bl[32] br[32] wl[425] vdd gnd cell_6t
Xbit_r426_c32 bl[32] br[32] wl[426] vdd gnd cell_6t
Xbit_r427_c32 bl[32] br[32] wl[427] vdd gnd cell_6t
Xbit_r428_c32 bl[32] br[32] wl[428] vdd gnd cell_6t
Xbit_r429_c32 bl[32] br[32] wl[429] vdd gnd cell_6t
Xbit_r430_c32 bl[32] br[32] wl[430] vdd gnd cell_6t
Xbit_r431_c32 bl[32] br[32] wl[431] vdd gnd cell_6t
Xbit_r432_c32 bl[32] br[32] wl[432] vdd gnd cell_6t
Xbit_r433_c32 bl[32] br[32] wl[433] vdd gnd cell_6t
Xbit_r434_c32 bl[32] br[32] wl[434] vdd gnd cell_6t
Xbit_r435_c32 bl[32] br[32] wl[435] vdd gnd cell_6t
Xbit_r436_c32 bl[32] br[32] wl[436] vdd gnd cell_6t
Xbit_r437_c32 bl[32] br[32] wl[437] vdd gnd cell_6t
Xbit_r438_c32 bl[32] br[32] wl[438] vdd gnd cell_6t
Xbit_r439_c32 bl[32] br[32] wl[439] vdd gnd cell_6t
Xbit_r440_c32 bl[32] br[32] wl[440] vdd gnd cell_6t
Xbit_r441_c32 bl[32] br[32] wl[441] vdd gnd cell_6t
Xbit_r442_c32 bl[32] br[32] wl[442] vdd gnd cell_6t
Xbit_r443_c32 bl[32] br[32] wl[443] vdd gnd cell_6t
Xbit_r444_c32 bl[32] br[32] wl[444] vdd gnd cell_6t
Xbit_r445_c32 bl[32] br[32] wl[445] vdd gnd cell_6t
Xbit_r446_c32 bl[32] br[32] wl[446] vdd gnd cell_6t
Xbit_r447_c32 bl[32] br[32] wl[447] vdd gnd cell_6t
Xbit_r448_c32 bl[32] br[32] wl[448] vdd gnd cell_6t
Xbit_r449_c32 bl[32] br[32] wl[449] vdd gnd cell_6t
Xbit_r450_c32 bl[32] br[32] wl[450] vdd gnd cell_6t
Xbit_r451_c32 bl[32] br[32] wl[451] vdd gnd cell_6t
Xbit_r452_c32 bl[32] br[32] wl[452] vdd gnd cell_6t
Xbit_r453_c32 bl[32] br[32] wl[453] vdd gnd cell_6t
Xbit_r454_c32 bl[32] br[32] wl[454] vdd gnd cell_6t
Xbit_r455_c32 bl[32] br[32] wl[455] vdd gnd cell_6t
Xbit_r456_c32 bl[32] br[32] wl[456] vdd gnd cell_6t
Xbit_r457_c32 bl[32] br[32] wl[457] vdd gnd cell_6t
Xbit_r458_c32 bl[32] br[32] wl[458] vdd gnd cell_6t
Xbit_r459_c32 bl[32] br[32] wl[459] vdd gnd cell_6t
Xbit_r460_c32 bl[32] br[32] wl[460] vdd gnd cell_6t
Xbit_r461_c32 bl[32] br[32] wl[461] vdd gnd cell_6t
Xbit_r462_c32 bl[32] br[32] wl[462] vdd gnd cell_6t
Xbit_r463_c32 bl[32] br[32] wl[463] vdd gnd cell_6t
Xbit_r464_c32 bl[32] br[32] wl[464] vdd gnd cell_6t
Xbit_r465_c32 bl[32] br[32] wl[465] vdd gnd cell_6t
Xbit_r466_c32 bl[32] br[32] wl[466] vdd gnd cell_6t
Xbit_r467_c32 bl[32] br[32] wl[467] vdd gnd cell_6t
Xbit_r468_c32 bl[32] br[32] wl[468] vdd gnd cell_6t
Xbit_r469_c32 bl[32] br[32] wl[469] vdd gnd cell_6t
Xbit_r470_c32 bl[32] br[32] wl[470] vdd gnd cell_6t
Xbit_r471_c32 bl[32] br[32] wl[471] vdd gnd cell_6t
Xbit_r472_c32 bl[32] br[32] wl[472] vdd gnd cell_6t
Xbit_r473_c32 bl[32] br[32] wl[473] vdd gnd cell_6t
Xbit_r474_c32 bl[32] br[32] wl[474] vdd gnd cell_6t
Xbit_r475_c32 bl[32] br[32] wl[475] vdd gnd cell_6t
Xbit_r476_c32 bl[32] br[32] wl[476] vdd gnd cell_6t
Xbit_r477_c32 bl[32] br[32] wl[477] vdd gnd cell_6t
Xbit_r478_c32 bl[32] br[32] wl[478] vdd gnd cell_6t
Xbit_r479_c32 bl[32] br[32] wl[479] vdd gnd cell_6t
Xbit_r480_c32 bl[32] br[32] wl[480] vdd gnd cell_6t
Xbit_r481_c32 bl[32] br[32] wl[481] vdd gnd cell_6t
Xbit_r482_c32 bl[32] br[32] wl[482] vdd gnd cell_6t
Xbit_r483_c32 bl[32] br[32] wl[483] vdd gnd cell_6t
Xbit_r484_c32 bl[32] br[32] wl[484] vdd gnd cell_6t
Xbit_r485_c32 bl[32] br[32] wl[485] vdd gnd cell_6t
Xbit_r486_c32 bl[32] br[32] wl[486] vdd gnd cell_6t
Xbit_r487_c32 bl[32] br[32] wl[487] vdd gnd cell_6t
Xbit_r488_c32 bl[32] br[32] wl[488] vdd gnd cell_6t
Xbit_r489_c32 bl[32] br[32] wl[489] vdd gnd cell_6t
Xbit_r490_c32 bl[32] br[32] wl[490] vdd gnd cell_6t
Xbit_r491_c32 bl[32] br[32] wl[491] vdd gnd cell_6t
Xbit_r492_c32 bl[32] br[32] wl[492] vdd gnd cell_6t
Xbit_r493_c32 bl[32] br[32] wl[493] vdd gnd cell_6t
Xbit_r494_c32 bl[32] br[32] wl[494] vdd gnd cell_6t
Xbit_r495_c32 bl[32] br[32] wl[495] vdd gnd cell_6t
Xbit_r496_c32 bl[32] br[32] wl[496] vdd gnd cell_6t
Xbit_r497_c32 bl[32] br[32] wl[497] vdd gnd cell_6t
Xbit_r498_c32 bl[32] br[32] wl[498] vdd gnd cell_6t
Xbit_r499_c32 bl[32] br[32] wl[499] vdd gnd cell_6t
Xbit_r500_c32 bl[32] br[32] wl[500] vdd gnd cell_6t
Xbit_r501_c32 bl[32] br[32] wl[501] vdd gnd cell_6t
Xbit_r502_c32 bl[32] br[32] wl[502] vdd gnd cell_6t
Xbit_r503_c32 bl[32] br[32] wl[503] vdd gnd cell_6t
Xbit_r504_c32 bl[32] br[32] wl[504] vdd gnd cell_6t
Xbit_r505_c32 bl[32] br[32] wl[505] vdd gnd cell_6t
Xbit_r506_c32 bl[32] br[32] wl[506] vdd gnd cell_6t
Xbit_r507_c32 bl[32] br[32] wl[507] vdd gnd cell_6t
Xbit_r508_c32 bl[32] br[32] wl[508] vdd gnd cell_6t
Xbit_r509_c32 bl[32] br[32] wl[509] vdd gnd cell_6t
Xbit_r510_c32 bl[32] br[32] wl[510] vdd gnd cell_6t
Xbit_r511_c32 bl[32] br[32] wl[511] vdd gnd cell_6t
Xbit_r0_c33 bl[33] br[33] wl[0] vdd gnd cell_6t
Xbit_r1_c33 bl[33] br[33] wl[1] vdd gnd cell_6t
Xbit_r2_c33 bl[33] br[33] wl[2] vdd gnd cell_6t
Xbit_r3_c33 bl[33] br[33] wl[3] vdd gnd cell_6t
Xbit_r4_c33 bl[33] br[33] wl[4] vdd gnd cell_6t
Xbit_r5_c33 bl[33] br[33] wl[5] vdd gnd cell_6t
Xbit_r6_c33 bl[33] br[33] wl[6] vdd gnd cell_6t
Xbit_r7_c33 bl[33] br[33] wl[7] vdd gnd cell_6t
Xbit_r8_c33 bl[33] br[33] wl[8] vdd gnd cell_6t
Xbit_r9_c33 bl[33] br[33] wl[9] vdd gnd cell_6t
Xbit_r10_c33 bl[33] br[33] wl[10] vdd gnd cell_6t
Xbit_r11_c33 bl[33] br[33] wl[11] vdd gnd cell_6t
Xbit_r12_c33 bl[33] br[33] wl[12] vdd gnd cell_6t
Xbit_r13_c33 bl[33] br[33] wl[13] vdd gnd cell_6t
Xbit_r14_c33 bl[33] br[33] wl[14] vdd gnd cell_6t
Xbit_r15_c33 bl[33] br[33] wl[15] vdd gnd cell_6t
Xbit_r16_c33 bl[33] br[33] wl[16] vdd gnd cell_6t
Xbit_r17_c33 bl[33] br[33] wl[17] vdd gnd cell_6t
Xbit_r18_c33 bl[33] br[33] wl[18] vdd gnd cell_6t
Xbit_r19_c33 bl[33] br[33] wl[19] vdd gnd cell_6t
Xbit_r20_c33 bl[33] br[33] wl[20] vdd gnd cell_6t
Xbit_r21_c33 bl[33] br[33] wl[21] vdd gnd cell_6t
Xbit_r22_c33 bl[33] br[33] wl[22] vdd gnd cell_6t
Xbit_r23_c33 bl[33] br[33] wl[23] vdd gnd cell_6t
Xbit_r24_c33 bl[33] br[33] wl[24] vdd gnd cell_6t
Xbit_r25_c33 bl[33] br[33] wl[25] vdd gnd cell_6t
Xbit_r26_c33 bl[33] br[33] wl[26] vdd gnd cell_6t
Xbit_r27_c33 bl[33] br[33] wl[27] vdd gnd cell_6t
Xbit_r28_c33 bl[33] br[33] wl[28] vdd gnd cell_6t
Xbit_r29_c33 bl[33] br[33] wl[29] vdd gnd cell_6t
Xbit_r30_c33 bl[33] br[33] wl[30] vdd gnd cell_6t
Xbit_r31_c33 bl[33] br[33] wl[31] vdd gnd cell_6t
Xbit_r32_c33 bl[33] br[33] wl[32] vdd gnd cell_6t
Xbit_r33_c33 bl[33] br[33] wl[33] vdd gnd cell_6t
Xbit_r34_c33 bl[33] br[33] wl[34] vdd gnd cell_6t
Xbit_r35_c33 bl[33] br[33] wl[35] vdd gnd cell_6t
Xbit_r36_c33 bl[33] br[33] wl[36] vdd gnd cell_6t
Xbit_r37_c33 bl[33] br[33] wl[37] vdd gnd cell_6t
Xbit_r38_c33 bl[33] br[33] wl[38] vdd gnd cell_6t
Xbit_r39_c33 bl[33] br[33] wl[39] vdd gnd cell_6t
Xbit_r40_c33 bl[33] br[33] wl[40] vdd gnd cell_6t
Xbit_r41_c33 bl[33] br[33] wl[41] vdd gnd cell_6t
Xbit_r42_c33 bl[33] br[33] wl[42] vdd gnd cell_6t
Xbit_r43_c33 bl[33] br[33] wl[43] vdd gnd cell_6t
Xbit_r44_c33 bl[33] br[33] wl[44] vdd gnd cell_6t
Xbit_r45_c33 bl[33] br[33] wl[45] vdd gnd cell_6t
Xbit_r46_c33 bl[33] br[33] wl[46] vdd gnd cell_6t
Xbit_r47_c33 bl[33] br[33] wl[47] vdd gnd cell_6t
Xbit_r48_c33 bl[33] br[33] wl[48] vdd gnd cell_6t
Xbit_r49_c33 bl[33] br[33] wl[49] vdd gnd cell_6t
Xbit_r50_c33 bl[33] br[33] wl[50] vdd gnd cell_6t
Xbit_r51_c33 bl[33] br[33] wl[51] vdd gnd cell_6t
Xbit_r52_c33 bl[33] br[33] wl[52] vdd gnd cell_6t
Xbit_r53_c33 bl[33] br[33] wl[53] vdd gnd cell_6t
Xbit_r54_c33 bl[33] br[33] wl[54] vdd gnd cell_6t
Xbit_r55_c33 bl[33] br[33] wl[55] vdd gnd cell_6t
Xbit_r56_c33 bl[33] br[33] wl[56] vdd gnd cell_6t
Xbit_r57_c33 bl[33] br[33] wl[57] vdd gnd cell_6t
Xbit_r58_c33 bl[33] br[33] wl[58] vdd gnd cell_6t
Xbit_r59_c33 bl[33] br[33] wl[59] vdd gnd cell_6t
Xbit_r60_c33 bl[33] br[33] wl[60] vdd gnd cell_6t
Xbit_r61_c33 bl[33] br[33] wl[61] vdd gnd cell_6t
Xbit_r62_c33 bl[33] br[33] wl[62] vdd gnd cell_6t
Xbit_r63_c33 bl[33] br[33] wl[63] vdd gnd cell_6t
Xbit_r64_c33 bl[33] br[33] wl[64] vdd gnd cell_6t
Xbit_r65_c33 bl[33] br[33] wl[65] vdd gnd cell_6t
Xbit_r66_c33 bl[33] br[33] wl[66] vdd gnd cell_6t
Xbit_r67_c33 bl[33] br[33] wl[67] vdd gnd cell_6t
Xbit_r68_c33 bl[33] br[33] wl[68] vdd gnd cell_6t
Xbit_r69_c33 bl[33] br[33] wl[69] vdd gnd cell_6t
Xbit_r70_c33 bl[33] br[33] wl[70] vdd gnd cell_6t
Xbit_r71_c33 bl[33] br[33] wl[71] vdd gnd cell_6t
Xbit_r72_c33 bl[33] br[33] wl[72] vdd gnd cell_6t
Xbit_r73_c33 bl[33] br[33] wl[73] vdd gnd cell_6t
Xbit_r74_c33 bl[33] br[33] wl[74] vdd gnd cell_6t
Xbit_r75_c33 bl[33] br[33] wl[75] vdd gnd cell_6t
Xbit_r76_c33 bl[33] br[33] wl[76] vdd gnd cell_6t
Xbit_r77_c33 bl[33] br[33] wl[77] vdd gnd cell_6t
Xbit_r78_c33 bl[33] br[33] wl[78] vdd gnd cell_6t
Xbit_r79_c33 bl[33] br[33] wl[79] vdd gnd cell_6t
Xbit_r80_c33 bl[33] br[33] wl[80] vdd gnd cell_6t
Xbit_r81_c33 bl[33] br[33] wl[81] vdd gnd cell_6t
Xbit_r82_c33 bl[33] br[33] wl[82] vdd gnd cell_6t
Xbit_r83_c33 bl[33] br[33] wl[83] vdd gnd cell_6t
Xbit_r84_c33 bl[33] br[33] wl[84] vdd gnd cell_6t
Xbit_r85_c33 bl[33] br[33] wl[85] vdd gnd cell_6t
Xbit_r86_c33 bl[33] br[33] wl[86] vdd gnd cell_6t
Xbit_r87_c33 bl[33] br[33] wl[87] vdd gnd cell_6t
Xbit_r88_c33 bl[33] br[33] wl[88] vdd gnd cell_6t
Xbit_r89_c33 bl[33] br[33] wl[89] vdd gnd cell_6t
Xbit_r90_c33 bl[33] br[33] wl[90] vdd gnd cell_6t
Xbit_r91_c33 bl[33] br[33] wl[91] vdd gnd cell_6t
Xbit_r92_c33 bl[33] br[33] wl[92] vdd gnd cell_6t
Xbit_r93_c33 bl[33] br[33] wl[93] vdd gnd cell_6t
Xbit_r94_c33 bl[33] br[33] wl[94] vdd gnd cell_6t
Xbit_r95_c33 bl[33] br[33] wl[95] vdd gnd cell_6t
Xbit_r96_c33 bl[33] br[33] wl[96] vdd gnd cell_6t
Xbit_r97_c33 bl[33] br[33] wl[97] vdd gnd cell_6t
Xbit_r98_c33 bl[33] br[33] wl[98] vdd gnd cell_6t
Xbit_r99_c33 bl[33] br[33] wl[99] vdd gnd cell_6t
Xbit_r100_c33 bl[33] br[33] wl[100] vdd gnd cell_6t
Xbit_r101_c33 bl[33] br[33] wl[101] vdd gnd cell_6t
Xbit_r102_c33 bl[33] br[33] wl[102] vdd gnd cell_6t
Xbit_r103_c33 bl[33] br[33] wl[103] vdd gnd cell_6t
Xbit_r104_c33 bl[33] br[33] wl[104] vdd gnd cell_6t
Xbit_r105_c33 bl[33] br[33] wl[105] vdd gnd cell_6t
Xbit_r106_c33 bl[33] br[33] wl[106] vdd gnd cell_6t
Xbit_r107_c33 bl[33] br[33] wl[107] vdd gnd cell_6t
Xbit_r108_c33 bl[33] br[33] wl[108] vdd gnd cell_6t
Xbit_r109_c33 bl[33] br[33] wl[109] vdd gnd cell_6t
Xbit_r110_c33 bl[33] br[33] wl[110] vdd gnd cell_6t
Xbit_r111_c33 bl[33] br[33] wl[111] vdd gnd cell_6t
Xbit_r112_c33 bl[33] br[33] wl[112] vdd gnd cell_6t
Xbit_r113_c33 bl[33] br[33] wl[113] vdd gnd cell_6t
Xbit_r114_c33 bl[33] br[33] wl[114] vdd gnd cell_6t
Xbit_r115_c33 bl[33] br[33] wl[115] vdd gnd cell_6t
Xbit_r116_c33 bl[33] br[33] wl[116] vdd gnd cell_6t
Xbit_r117_c33 bl[33] br[33] wl[117] vdd gnd cell_6t
Xbit_r118_c33 bl[33] br[33] wl[118] vdd gnd cell_6t
Xbit_r119_c33 bl[33] br[33] wl[119] vdd gnd cell_6t
Xbit_r120_c33 bl[33] br[33] wl[120] vdd gnd cell_6t
Xbit_r121_c33 bl[33] br[33] wl[121] vdd gnd cell_6t
Xbit_r122_c33 bl[33] br[33] wl[122] vdd gnd cell_6t
Xbit_r123_c33 bl[33] br[33] wl[123] vdd gnd cell_6t
Xbit_r124_c33 bl[33] br[33] wl[124] vdd gnd cell_6t
Xbit_r125_c33 bl[33] br[33] wl[125] vdd gnd cell_6t
Xbit_r126_c33 bl[33] br[33] wl[126] vdd gnd cell_6t
Xbit_r127_c33 bl[33] br[33] wl[127] vdd gnd cell_6t
Xbit_r128_c33 bl[33] br[33] wl[128] vdd gnd cell_6t
Xbit_r129_c33 bl[33] br[33] wl[129] vdd gnd cell_6t
Xbit_r130_c33 bl[33] br[33] wl[130] vdd gnd cell_6t
Xbit_r131_c33 bl[33] br[33] wl[131] vdd gnd cell_6t
Xbit_r132_c33 bl[33] br[33] wl[132] vdd gnd cell_6t
Xbit_r133_c33 bl[33] br[33] wl[133] vdd gnd cell_6t
Xbit_r134_c33 bl[33] br[33] wl[134] vdd gnd cell_6t
Xbit_r135_c33 bl[33] br[33] wl[135] vdd gnd cell_6t
Xbit_r136_c33 bl[33] br[33] wl[136] vdd gnd cell_6t
Xbit_r137_c33 bl[33] br[33] wl[137] vdd gnd cell_6t
Xbit_r138_c33 bl[33] br[33] wl[138] vdd gnd cell_6t
Xbit_r139_c33 bl[33] br[33] wl[139] vdd gnd cell_6t
Xbit_r140_c33 bl[33] br[33] wl[140] vdd gnd cell_6t
Xbit_r141_c33 bl[33] br[33] wl[141] vdd gnd cell_6t
Xbit_r142_c33 bl[33] br[33] wl[142] vdd gnd cell_6t
Xbit_r143_c33 bl[33] br[33] wl[143] vdd gnd cell_6t
Xbit_r144_c33 bl[33] br[33] wl[144] vdd gnd cell_6t
Xbit_r145_c33 bl[33] br[33] wl[145] vdd gnd cell_6t
Xbit_r146_c33 bl[33] br[33] wl[146] vdd gnd cell_6t
Xbit_r147_c33 bl[33] br[33] wl[147] vdd gnd cell_6t
Xbit_r148_c33 bl[33] br[33] wl[148] vdd gnd cell_6t
Xbit_r149_c33 bl[33] br[33] wl[149] vdd gnd cell_6t
Xbit_r150_c33 bl[33] br[33] wl[150] vdd gnd cell_6t
Xbit_r151_c33 bl[33] br[33] wl[151] vdd gnd cell_6t
Xbit_r152_c33 bl[33] br[33] wl[152] vdd gnd cell_6t
Xbit_r153_c33 bl[33] br[33] wl[153] vdd gnd cell_6t
Xbit_r154_c33 bl[33] br[33] wl[154] vdd gnd cell_6t
Xbit_r155_c33 bl[33] br[33] wl[155] vdd gnd cell_6t
Xbit_r156_c33 bl[33] br[33] wl[156] vdd gnd cell_6t
Xbit_r157_c33 bl[33] br[33] wl[157] vdd gnd cell_6t
Xbit_r158_c33 bl[33] br[33] wl[158] vdd gnd cell_6t
Xbit_r159_c33 bl[33] br[33] wl[159] vdd gnd cell_6t
Xbit_r160_c33 bl[33] br[33] wl[160] vdd gnd cell_6t
Xbit_r161_c33 bl[33] br[33] wl[161] vdd gnd cell_6t
Xbit_r162_c33 bl[33] br[33] wl[162] vdd gnd cell_6t
Xbit_r163_c33 bl[33] br[33] wl[163] vdd gnd cell_6t
Xbit_r164_c33 bl[33] br[33] wl[164] vdd gnd cell_6t
Xbit_r165_c33 bl[33] br[33] wl[165] vdd gnd cell_6t
Xbit_r166_c33 bl[33] br[33] wl[166] vdd gnd cell_6t
Xbit_r167_c33 bl[33] br[33] wl[167] vdd gnd cell_6t
Xbit_r168_c33 bl[33] br[33] wl[168] vdd gnd cell_6t
Xbit_r169_c33 bl[33] br[33] wl[169] vdd gnd cell_6t
Xbit_r170_c33 bl[33] br[33] wl[170] vdd gnd cell_6t
Xbit_r171_c33 bl[33] br[33] wl[171] vdd gnd cell_6t
Xbit_r172_c33 bl[33] br[33] wl[172] vdd gnd cell_6t
Xbit_r173_c33 bl[33] br[33] wl[173] vdd gnd cell_6t
Xbit_r174_c33 bl[33] br[33] wl[174] vdd gnd cell_6t
Xbit_r175_c33 bl[33] br[33] wl[175] vdd gnd cell_6t
Xbit_r176_c33 bl[33] br[33] wl[176] vdd gnd cell_6t
Xbit_r177_c33 bl[33] br[33] wl[177] vdd gnd cell_6t
Xbit_r178_c33 bl[33] br[33] wl[178] vdd gnd cell_6t
Xbit_r179_c33 bl[33] br[33] wl[179] vdd gnd cell_6t
Xbit_r180_c33 bl[33] br[33] wl[180] vdd gnd cell_6t
Xbit_r181_c33 bl[33] br[33] wl[181] vdd gnd cell_6t
Xbit_r182_c33 bl[33] br[33] wl[182] vdd gnd cell_6t
Xbit_r183_c33 bl[33] br[33] wl[183] vdd gnd cell_6t
Xbit_r184_c33 bl[33] br[33] wl[184] vdd gnd cell_6t
Xbit_r185_c33 bl[33] br[33] wl[185] vdd gnd cell_6t
Xbit_r186_c33 bl[33] br[33] wl[186] vdd gnd cell_6t
Xbit_r187_c33 bl[33] br[33] wl[187] vdd gnd cell_6t
Xbit_r188_c33 bl[33] br[33] wl[188] vdd gnd cell_6t
Xbit_r189_c33 bl[33] br[33] wl[189] vdd gnd cell_6t
Xbit_r190_c33 bl[33] br[33] wl[190] vdd gnd cell_6t
Xbit_r191_c33 bl[33] br[33] wl[191] vdd gnd cell_6t
Xbit_r192_c33 bl[33] br[33] wl[192] vdd gnd cell_6t
Xbit_r193_c33 bl[33] br[33] wl[193] vdd gnd cell_6t
Xbit_r194_c33 bl[33] br[33] wl[194] vdd gnd cell_6t
Xbit_r195_c33 bl[33] br[33] wl[195] vdd gnd cell_6t
Xbit_r196_c33 bl[33] br[33] wl[196] vdd gnd cell_6t
Xbit_r197_c33 bl[33] br[33] wl[197] vdd gnd cell_6t
Xbit_r198_c33 bl[33] br[33] wl[198] vdd gnd cell_6t
Xbit_r199_c33 bl[33] br[33] wl[199] vdd gnd cell_6t
Xbit_r200_c33 bl[33] br[33] wl[200] vdd gnd cell_6t
Xbit_r201_c33 bl[33] br[33] wl[201] vdd gnd cell_6t
Xbit_r202_c33 bl[33] br[33] wl[202] vdd gnd cell_6t
Xbit_r203_c33 bl[33] br[33] wl[203] vdd gnd cell_6t
Xbit_r204_c33 bl[33] br[33] wl[204] vdd gnd cell_6t
Xbit_r205_c33 bl[33] br[33] wl[205] vdd gnd cell_6t
Xbit_r206_c33 bl[33] br[33] wl[206] vdd gnd cell_6t
Xbit_r207_c33 bl[33] br[33] wl[207] vdd gnd cell_6t
Xbit_r208_c33 bl[33] br[33] wl[208] vdd gnd cell_6t
Xbit_r209_c33 bl[33] br[33] wl[209] vdd gnd cell_6t
Xbit_r210_c33 bl[33] br[33] wl[210] vdd gnd cell_6t
Xbit_r211_c33 bl[33] br[33] wl[211] vdd gnd cell_6t
Xbit_r212_c33 bl[33] br[33] wl[212] vdd gnd cell_6t
Xbit_r213_c33 bl[33] br[33] wl[213] vdd gnd cell_6t
Xbit_r214_c33 bl[33] br[33] wl[214] vdd gnd cell_6t
Xbit_r215_c33 bl[33] br[33] wl[215] vdd gnd cell_6t
Xbit_r216_c33 bl[33] br[33] wl[216] vdd gnd cell_6t
Xbit_r217_c33 bl[33] br[33] wl[217] vdd gnd cell_6t
Xbit_r218_c33 bl[33] br[33] wl[218] vdd gnd cell_6t
Xbit_r219_c33 bl[33] br[33] wl[219] vdd gnd cell_6t
Xbit_r220_c33 bl[33] br[33] wl[220] vdd gnd cell_6t
Xbit_r221_c33 bl[33] br[33] wl[221] vdd gnd cell_6t
Xbit_r222_c33 bl[33] br[33] wl[222] vdd gnd cell_6t
Xbit_r223_c33 bl[33] br[33] wl[223] vdd gnd cell_6t
Xbit_r224_c33 bl[33] br[33] wl[224] vdd gnd cell_6t
Xbit_r225_c33 bl[33] br[33] wl[225] vdd gnd cell_6t
Xbit_r226_c33 bl[33] br[33] wl[226] vdd gnd cell_6t
Xbit_r227_c33 bl[33] br[33] wl[227] vdd gnd cell_6t
Xbit_r228_c33 bl[33] br[33] wl[228] vdd gnd cell_6t
Xbit_r229_c33 bl[33] br[33] wl[229] vdd gnd cell_6t
Xbit_r230_c33 bl[33] br[33] wl[230] vdd gnd cell_6t
Xbit_r231_c33 bl[33] br[33] wl[231] vdd gnd cell_6t
Xbit_r232_c33 bl[33] br[33] wl[232] vdd gnd cell_6t
Xbit_r233_c33 bl[33] br[33] wl[233] vdd gnd cell_6t
Xbit_r234_c33 bl[33] br[33] wl[234] vdd gnd cell_6t
Xbit_r235_c33 bl[33] br[33] wl[235] vdd gnd cell_6t
Xbit_r236_c33 bl[33] br[33] wl[236] vdd gnd cell_6t
Xbit_r237_c33 bl[33] br[33] wl[237] vdd gnd cell_6t
Xbit_r238_c33 bl[33] br[33] wl[238] vdd gnd cell_6t
Xbit_r239_c33 bl[33] br[33] wl[239] vdd gnd cell_6t
Xbit_r240_c33 bl[33] br[33] wl[240] vdd gnd cell_6t
Xbit_r241_c33 bl[33] br[33] wl[241] vdd gnd cell_6t
Xbit_r242_c33 bl[33] br[33] wl[242] vdd gnd cell_6t
Xbit_r243_c33 bl[33] br[33] wl[243] vdd gnd cell_6t
Xbit_r244_c33 bl[33] br[33] wl[244] vdd gnd cell_6t
Xbit_r245_c33 bl[33] br[33] wl[245] vdd gnd cell_6t
Xbit_r246_c33 bl[33] br[33] wl[246] vdd gnd cell_6t
Xbit_r247_c33 bl[33] br[33] wl[247] vdd gnd cell_6t
Xbit_r248_c33 bl[33] br[33] wl[248] vdd gnd cell_6t
Xbit_r249_c33 bl[33] br[33] wl[249] vdd gnd cell_6t
Xbit_r250_c33 bl[33] br[33] wl[250] vdd gnd cell_6t
Xbit_r251_c33 bl[33] br[33] wl[251] vdd gnd cell_6t
Xbit_r252_c33 bl[33] br[33] wl[252] vdd gnd cell_6t
Xbit_r253_c33 bl[33] br[33] wl[253] vdd gnd cell_6t
Xbit_r254_c33 bl[33] br[33] wl[254] vdd gnd cell_6t
Xbit_r255_c33 bl[33] br[33] wl[255] vdd gnd cell_6t
Xbit_r256_c33 bl[33] br[33] wl[256] vdd gnd cell_6t
Xbit_r257_c33 bl[33] br[33] wl[257] vdd gnd cell_6t
Xbit_r258_c33 bl[33] br[33] wl[258] vdd gnd cell_6t
Xbit_r259_c33 bl[33] br[33] wl[259] vdd gnd cell_6t
Xbit_r260_c33 bl[33] br[33] wl[260] vdd gnd cell_6t
Xbit_r261_c33 bl[33] br[33] wl[261] vdd gnd cell_6t
Xbit_r262_c33 bl[33] br[33] wl[262] vdd gnd cell_6t
Xbit_r263_c33 bl[33] br[33] wl[263] vdd gnd cell_6t
Xbit_r264_c33 bl[33] br[33] wl[264] vdd gnd cell_6t
Xbit_r265_c33 bl[33] br[33] wl[265] vdd gnd cell_6t
Xbit_r266_c33 bl[33] br[33] wl[266] vdd gnd cell_6t
Xbit_r267_c33 bl[33] br[33] wl[267] vdd gnd cell_6t
Xbit_r268_c33 bl[33] br[33] wl[268] vdd gnd cell_6t
Xbit_r269_c33 bl[33] br[33] wl[269] vdd gnd cell_6t
Xbit_r270_c33 bl[33] br[33] wl[270] vdd gnd cell_6t
Xbit_r271_c33 bl[33] br[33] wl[271] vdd gnd cell_6t
Xbit_r272_c33 bl[33] br[33] wl[272] vdd gnd cell_6t
Xbit_r273_c33 bl[33] br[33] wl[273] vdd gnd cell_6t
Xbit_r274_c33 bl[33] br[33] wl[274] vdd gnd cell_6t
Xbit_r275_c33 bl[33] br[33] wl[275] vdd gnd cell_6t
Xbit_r276_c33 bl[33] br[33] wl[276] vdd gnd cell_6t
Xbit_r277_c33 bl[33] br[33] wl[277] vdd gnd cell_6t
Xbit_r278_c33 bl[33] br[33] wl[278] vdd gnd cell_6t
Xbit_r279_c33 bl[33] br[33] wl[279] vdd gnd cell_6t
Xbit_r280_c33 bl[33] br[33] wl[280] vdd gnd cell_6t
Xbit_r281_c33 bl[33] br[33] wl[281] vdd gnd cell_6t
Xbit_r282_c33 bl[33] br[33] wl[282] vdd gnd cell_6t
Xbit_r283_c33 bl[33] br[33] wl[283] vdd gnd cell_6t
Xbit_r284_c33 bl[33] br[33] wl[284] vdd gnd cell_6t
Xbit_r285_c33 bl[33] br[33] wl[285] vdd gnd cell_6t
Xbit_r286_c33 bl[33] br[33] wl[286] vdd gnd cell_6t
Xbit_r287_c33 bl[33] br[33] wl[287] vdd gnd cell_6t
Xbit_r288_c33 bl[33] br[33] wl[288] vdd gnd cell_6t
Xbit_r289_c33 bl[33] br[33] wl[289] vdd gnd cell_6t
Xbit_r290_c33 bl[33] br[33] wl[290] vdd gnd cell_6t
Xbit_r291_c33 bl[33] br[33] wl[291] vdd gnd cell_6t
Xbit_r292_c33 bl[33] br[33] wl[292] vdd gnd cell_6t
Xbit_r293_c33 bl[33] br[33] wl[293] vdd gnd cell_6t
Xbit_r294_c33 bl[33] br[33] wl[294] vdd gnd cell_6t
Xbit_r295_c33 bl[33] br[33] wl[295] vdd gnd cell_6t
Xbit_r296_c33 bl[33] br[33] wl[296] vdd gnd cell_6t
Xbit_r297_c33 bl[33] br[33] wl[297] vdd gnd cell_6t
Xbit_r298_c33 bl[33] br[33] wl[298] vdd gnd cell_6t
Xbit_r299_c33 bl[33] br[33] wl[299] vdd gnd cell_6t
Xbit_r300_c33 bl[33] br[33] wl[300] vdd gnd cell_6t
Xbit_r301_c33 bl[33] br[33] wl[301] vdd gnd cell_6t
Xbit_r302_c33 bl[33] br[33] wl[302] vdd gnd cell_6t
Xbit_r303_c33 bl[33] br[33] wl[303] vdd gnd cell_6t
Xbit_r304_c33 bl[33] br[33] wl[304] vdd gnd cell_6t
Xbit_r305_c33 bl[33] br[33] wl[305] vdd gnd cell_6t
Xbit_r306_c33 bl[33] br[33] wl[306] vdd gnd cell_6t
Xbit_r307_c33 bl[33] br[33] wl[307] vdd gnd cell_6t
Xbit_r308_c33 bl[33] br[33] wl[308] vdd gnd cell_6t
Xbit_r309_c33 bl[33] br[33] wl[309] vdd gnd cell_6t
Xbit_r310_c33 bl[33] br[33] wl[310] vdd gnd cell_6t
Xbit_r311_c33 bl[33] br[33] wl[311] vdd gnd cell_6t
Xbit_r312_c33 bl[33] br[33] wl[312] vdd gnd cell_6t
Xbit_r313_c33 bl[33] br[33] wl[313] vdd gnd cell_6t
Xbit_r314_c33 bl[33] br[33] wl[314] vdd gnd cell_6t
Xbit_r315_c33 bl[33] br[33] wl[315] vdd gnd cell_6t
Xbit_r316_c33 bl[33] br[33] wl[316] vdd gnd cell_6t
Xbit_r317_c33 bl[33] br[33] wl[317] vdd gnd cell_6t
Xbit_r318_c33 bl[33] br[33] wl[318] vdd gnd cell_6t
Xbit_r319_c33 bl[33] br[33] wl[319] vdd gnd cell_6t
Xbit_r320_c33 bl[33] br[33] wl[320] vdd gnd cell_6t
Xbit_r321_c33 bl[33] br[33] wl[321] vdd gnd cell_6t
Xbit_r322_c33 bl[33] br[33] wl[322] vdd gnd cell_6t
Xbit_r323_c33 bl[33] br[33] wl[323] vdd gnd cell_6t
Xbit_r324_c33 bl[33] br[33] wl[324] vdd gnd cell_6t
Xbit_r325_c33 bl[33] br[33] wl[325] vdd gnd cell_6t
Xbit_r326_c33 bl[33] br[33] wl[326] vdd gnd cell_6t
Xbit_r327_c33 bl[33] br[33] wl[327] vdd gnd cell_6t
Xbit_r328_c33 bl[33] br[33] wl[328] vdd gnd cell_6t
Xbit_r329_c33 bl[33] br[33] wl[329] vdd gnd cell_6t
Xbit_r330_c33 bl[33] br[33] wl[330] vdd gnd cell_6t
Xbit_r331_c33 bl[33] br[33] wl[331] vdd gnd cell_6t
Xbit_r332_c33 bl[33] br[33] wl[332] vdd gnd cell_6t
Xbit_r333_c33 bl[33] br[33] wl[333] vdd gnd cell_6t
Xbit_r334_c33 bl[33] br[33] wl[334] vdd gnd cell_6t
Xbit_r335_c33 bl[33] br[33] wl[335] vdd gnd cell_6t
Xbit_r336_c33 bl[33] br[33] wl[336] vdd gnd cell_6t
Xbit_r337_c33 bl[33] br[33] wl[337] vdd gnd cell_6t
Xbit_r338_c33 bl[33] br[33] wl[338] vdd gnd cell_6t
Xbit_r339_c33 bl[33] br[33] wl[339] vdd gnd cell_6t
Xbit_r340_c33 bl[33] br[33] wl[340] vdd gnd cell_6t
Xbit_r341_c33 bl[33] br[33] wl[341] vdd gnd cell_6t
Xbit_r342_c33 bl[33] br[33] wl[342] vdd gnd cell_6t
Xbit_r343_c33 bl[33] br[33] wl[343] vdd gnd cell_6t
Xbit_r344_c33 bl[33] br[33] wl[344] vdd gnd cell_6t
Xbit_r345_c33 bl[33] br[33] wl[345] vdd gnd cell_6t
Xbit_r346_c33 bl[33] br[33] wl[346] vdd gnd cell_6t
Xbit_r347_c33 bl[33] br[33] wl[347] vdd gnd cell_6t
Xbit_r348_c33 bl[33] br[33] wl[348] vdd gnd cell_6t
Xbit_r349_c33 bl[33] br[33] wl[349] vdd gnd cell_6t
Xbit_r350_c33 bl[33] br[33] wl[350] vdd gnd cell_6t
Xbit_r351_c33 bl[33] br[33] wl[351] vdd gnd cell_6t
Xbit_r352_c33 bl[33] br[33] wl[352] vdd gnd cell_6t
Xbit_r353_c33 bl[33] br[33] wl[353] vdd gnd cell_6t
Xbit_r354_c33 bl[33] br[33] wl[354] vdd gnd cell_6t
Xbit_r355_c33 bl[33] br[33] wl[355] vdd gnd cell_6t
Xbit_r356_c33 bl[33] br[33] wl[356] vdd gnd cell_6t
Xbit_r357_c33 bl[33] br[33] wl[357] vdd gnd cell_6t
Xbit_r358_c33 bl[33] br[33] wl[358] vdd gnd cell_6t
Xbit_r359_c33 bl[33] br[33] wl[359] vdd gnd cell_6t
Xbit_r360_c33 bl[33] br[33] wl[360] vdd gnd cell_6t
Xbit_r361_c33 bl[33] br[33] wl[361] vdd gnd cell_6t
Xbit_r362_c33 bl[33] br[33] wl[362] vdd gnd cell_6t
Xbit_r363_c33 bl[33] br[33] wl[363] vdd gnd cell_6t
Xbit_r364_c33 bl[33] br[33] wl[364] vdd gnd cell_6t
Xbit_r365_c33 bl[33] br[33] wl[365] vdd gnd cell_6t
Xbit_r366_c33 bl[33] br[33] wl[366] vdd gnd cell_6t
Xbit_r367_c33 bl[33] br[33] wl[367] vdd gnd cell_6t
Xbit_r368_c33 bl[33] br[33] wl[368] vdd gnd cell_6t
Xbit_r369_c33 bl[33] br[33] wl[369] vdd gnd cell_6t
Xbit_r370_c33 bl[33] br[33] wl[370] vdd gnd cell_6t
Xbit_r371_c33 bl[33] br[33] wl[371] vdd gnd cell_6t
Xbit_r372_c33 bl[33] br[33] wl[372] vdd gnd cell_6t
Xbit_r373_c33 bl[33] br[33] wl[373] vdd gnd cell_6t
Xbit_r374_c33 bl[33] br[33] wl[374] vdd gnd cell_6t
Xbit_r375_c33 bl[33] br[33] wl[375] vdd gnd cell_6t
Xbit_r376_c33 bl[33] br[33] wl[376] vdd gnd cell_6t
Xbit_r377_c33 bl[33] br[33] wl[377] vdd gnd cell_6t
Xbit_r378_c33 bl[33] br[33] wl[378] vdd gnd cell_6t
Xbit_r379_c33 bl[33] br[33] wl[379] vdd gnd cell_6t
Xbit_r380_c33 bl[33] br[33] wl[380] vdd gnd cell_6t
Xbit_r381_c33 bl[33] br[33] wl[381] vdd gnd cell_6t
Xbit_r382_c33 bl[33] br[33] wl[382] vdd gnd cell_6t
Xbit_r383_c33 bl[33] br[33] wl[383] vdd gnd cell_6t
Xbit_r384_c33 bl[33] br[33] wl[384] vdd gnd cell_6t
Xbit_r385_c33 bl[33] br[33] wl[385] vdd gnd cell_6t
Xbit_r386_c33 bl[33] br[33] wl[386] vdd gnd cell_6t
Xbit_r387_c33 bl[33] br[33] wl[387] vdd gnd cell_6t
Xbit_r388_c33 bl[33] br[33] wl[388] vdd gnd cell_6t
Xbit_r389_c33 bl[33] br[33] wl[389] vdd gnd cell_6t
Xbit_r390_c33 bl[33] br[33] wl[390] vdd gnd cell_6t
Xbit_r391_c33 bl[33] br[33] wl[391] vdd gnd cell_6t
Xbit_r392_c33 bl[33] br[33] wl[392] vdd gnd cell_6t
Xbit_r393_c33 bl[33] br[33] wl[393] vdd gnd cell_6t
Xbit_r394_c33 bl[33] br[33] wl[394] vdd gnd cell_6t
Xbit_r395_c33 bl[33] br[33] wl[395] vdd gnd cell_6t
Xbit_r396_c33 bl[33] br[33] wl[396] vdd gnd cell_6t
Xbit_r397_c33 bl[33] br[33] wl[397] vdd gnd cell_6t
Xbit_r398_c33 bl[33] br[33] wl[398] vdd gnd cell_6t
Xbit_r399_c33 bl[33] br[33] wl[399] vdd gnd cell_6t
Xbit_r400_c33 bl[33] br[33] wl[400] vdd gnd cell_6t
Xbit_r401_c33 bl[33] br[33] wl[401] vdd gnd cell_6t
Xbit_r402_c33 bl[33] br[33] wl[402] vdd gnd cell_6t
Xbit_r403_c33 bl[33] br[33] wl[403] vdd gnd cell_6t
Xbit_r404_c33 bl[33] br[33] wl[404] vdd gnd cell_6t
Xbit_r405_c33 bl[33] br[33] wl[405] vdd gnd cell_6t
Xbit_r406_c33 bl[33] br[33] wl[406] vdd gnd cell_6t
Xbit_r407_c33 bl[33] br[33] wl[407] vdd gnd cell_6t
Xbit_r408_c33 bl[33] br[33] wl[408] vdd gnd cell_6t
Xbit_r409_c33 bl[33] br[33] wl[409] vdd gnd cell_6t
Xbit_r410_c33 bl[33] br[33] wl[410] vdd gnd cell_6t
Xbit_r411_c33 bl[33] br[33] wl[411] vdd gnd cell_6t
Xbit_r412_c33 bl[33] br[33] wl[412] vdd gnd cell_6t
Xbit_r413_c33 bl[33] br[33] wl[413] vdd gnd cell_6t
Xbit_r414_c33 bl[33] br[33] wl[414] vdd gnd cell_6t
Xbit_r415_c33 bl[33] br[33] wl[415] vdd gnd cell_6t
Xbit_r416_c33 bl[33] br[33] wl[416] vdd gnd cell_6t
Xbit_r417_c33 bl[33] br[33] wl[417] vdd gnd cell_6t
Xbit_r418_c33 bl[33] br[33] wl[418] vdd gnd cell_6t
Xbit_r419_c33 bl[33] br[33] wl[419] vdd gnd cell_6t
Xbit_r420_c33 bl[33] br[33] wl[420] vdd gnd cell_6t
Xbit_r421_c33 bl[33] br[33] wl[421] vdd gnd cell_6t
Xbit_r422_c33 bl[33] br[33] wl[422] vdd gnd cell_6t
Xbit_r423_c33 bl[33] br[33] wl[423] vdd gnd cell_6t
Xbit_r424_c33 bl[33] br[33] wl[424] vdd gnd cell_6t
Xbit_r425_c33 bl[33] br[33] wl[425] vdd gnd cell_6t
Xbit_r426_c33 bl[33] br[33] wl[426] vdd gnd cell_6t
Xbit_r427_c33 bl[33] br[33] wl[427] vdd gnd cell_6t
Xbit_r428_c33 bl[33] br[33] wl[428] vdd gnd cell_6t
Xbit_r429_c33 bl[33] br[33] wl[429] vdd gnd cell_6t
Xbit_r430_c33 bl[33] br[33] wl[430] vdd gnd cell_6t
Xbit_r431_c33 bl[33] br[33] wl[431] vdd gnd cell_6t
Xbit_r432_c33 bl[33] br[33] wl[432] vdd gnd cell_6t
Xbit_r433_c33 bl[33] br[33] wl[433] vdd gnd cell_6t
Xbit_r434_c33 bl[33] br[33] wl[434] vdd gnd cell_6t
Xbit_r435_c33 bl[33] br[33] wl[435] vdd gnd cell_6t
Xbit_r436_c33 bl[33] br[33] wl[436] vdd gnd cell_6t
Xbit_r437_c33 bl[33] br[33] wl[437] vdd gnd cell_6t
Xbit_r438_c33 bl[33] br[33] wl[438] vdd gnd cell_6t
Xbit_r439_c33 bl[33] br[33] wl[439] vdd gnd cell_6t
Xbit_r440_c33 bl[33] br[33] wl[440] vdd gnd cell_6t
Xbit_r441_c33 bl[33] br[33] wl[441] vdd gnd cell_6t
Xbit_r442_c33 bl[33] br[33] wl[442] vdd gnd cell_6t
Xbit_r443_c33 bl[33] br[33] wl[443] vdd gnd cell_6t
Xbit_r444_c33 bl[33] br[33] wl[444] vdd gnd cell_6t
Xbit_r445_c33 bl[33] br[33] wl[445] vdd gnd cell_6t
Xbit_r446_c33 bl[33] br[33] wl[446] vdd gnd cell_6t
Xbit_r447_c33 bl[33] br[33] wl[447] vdd gnd cell_6t
Xbit_r448_c33 bl[33] br[33] wl[448] vdd gnd cell_6t
Xbit_r449_c33 bl[33] br[33] wl[449] vdd gnd cell_6t
Xbit_r450_c33 bl[33] br[33] wl[450] vdd gnd cell_6t
Xbit_r451_c33 bl[33] br[33] wl[451] vdd gnd cell_6t
Xbit_r452_c33 bl[33] br[33] wl[452] vdd gnd cell_6t
Xbit_r453_c33 bl[33] br[33] wl[453] vdd gnd cell_6t
Xbit_r454_c33 bl[33] br[33] wl[454] vdd gnd cell_6t
Xbit_r455_c33 bl[33] br[33] wl[455] vdd gnd cell_6t
Xbit_r456_c33 bl[33] br[33] wl[456] vdd gnd cell_6t
Xbit_r457_c33 bl[33] br[33] wl[457] vdd gnd cell_6t
Xbit_r458_c33 bl[33] br[33] wl[458] vdd gnd cell_6t
Xbit_r459_c33 bl[33] br[33] wl[459] vdd gnd cell_6t
Xbit_r460_c33 bl[33] br[33] wl[460] vdd gnd cell_6t
Xbit_r461_c33 bl[33] br[33] wl[461] vdd gnd cell_6t
Xbit_r462_c33 bl[33] br[33] wl[462] vdd gnd cell_6t
Xbit_r463_c33 bl[33] br[33] wl[463] vdd gnd cell_6t
Xbit_r464_c33 bl[33] br[33] wl[464] vdd gnd cell_6t
Xbit_r465_c33 bl[33] br[33] wl[465] vdd gnd cell_6t
Xbit_r466_c33 bl[33] br[33] wl[466] vdd gnd cell_6t
Xbit_r467_c33 bl[33] br[33] wl[467] vdd gnd cell_6t
Xbit_r468_c33 bl[33] br[33] wl[468] vdd gnd cell_6t
Xbit_r469_c33 bl[33] br[33] wl[469] vdd gnd cell_6t
Xbit_r470_c33 bl[33] br[33] wl[470] vdd gnd cell_6t
Xbit_r471_c33 bl[33] br[33] wl[471] vdd gnd cell_6t
Xbit_r472_c33 bl[33] br[33] wl[472] vdd gnd cell_6t
Xbit_r473_c33 bl[33] br[33] wl[473] vdd gnd cell_6t
Xbit_r474_c33 bl[33] br[33] wl[474] vdd gnd cell_6t
Xbit_r475_c33 bl[33] br[33] wl[475] vdd gnd cell_6t
Xbit_r476_c33 bl[33] br[33] wl[476] vdd gnd cell_6t
Xbit_r477_c33 bl[33] br[33] wl[477] vdd gnd cell_6t
Xbit_r478_c33 bl[33] br[33] wl[478] vdd gnd cell_6t
Xbit_r479_c33 bl[33] br[33] wl[479] vdd gnd cell_6t
Xbit_r480_c33 bl[33] br[33] wl[480] vdd gnd cell_6t
Xbit_r481_c33 bl[33] br[33] wl[481] vdd gnd cell_6t
Xbit_r482_c33 bl[33] br[33] wl[482] vdd gnd cell_6t
Xbit_r483_c33 bl[33] br[33] wl[483] vdd gnd cell_6t
Xbit_r484_c33 bl[33] br[33] wl[484] vdd gnd cell_6t
Xbit_r485_c33 bl[33] br[33] wl[485] vdd gnd cell_6t
Xbit_r486_c33 bl[33] br[33] wl[486] vdd gnd cell_6t
Xbit_r487_c33 bl[33] br[33] wl[487] vdd gnd cell_6t
Xbit_r488_c33 bl[33] br[33] wl[488] vdd gnd cell_6t
Xbit_r489_c33 bl[33] br[33] wl[489] vdd gnd cell_6t
Xbit_r490_c33 bl[33] br[33] wl[490] vdd gnd cell_6t
Xbit_r491_c33 bl[33] br[33] wl[491] vdd gnd cell_6t
Xbit_r492_c33 bl[33] br[33] wl[492] vdd gnd cell_6t
Xbit_r493_c33 bl[33] br[33] wl[493] vdd gnd cell_6t
Xbit_r494_c33 bl[33] br[33] wl[494] vdd gnd cell_6t
Xbit_r495_c33 bl[33] br[33] wl[495] vdd gnd cell_6t
Xbit_r496_c33 bl[33] br[33] wl[496] vdd gnd cell_6t
Xbit_r497_c33 bl[33] br[33] wl[497] vdd gnd cell_6t
Xbit_r498_c33 bl[33] br[33] wl[498] vdd gnd cell_6t
Xbit_r499_c33 bl[33] br[33] wl[499] vdd gnd cell_6t
Xbit_r500_c33 bl[33] br[33] wl[500] vdd gnd cell_6t
Xbit_r501_c33 bl[33] br[33] wl[501] vdd gnd cell_6t
Xbit_r502_c33 bl[33] br[33] wl[502] vdd gnd cell_6t
Xbit_r503_c33 bl[33] br[33] wl[503] vdd gnd cell_6t
Xbit_r504_c33 bl[33] br[33] wl[504] vdd gnd cell_6t
Xbit_r505_c33 bl[33] br[33] wl[505] vdd gnd cell_6t
Xbit_r506_c33 bl[33] br[33] wl[506] vdd gnd cell_6t
Xbit_r507_c33 bl[33] br[33] wl[507] vdd gnd cell_6t
Xbit_r508_c33 bl[33] br[33] wl[508] vdd gnd cell_6t
Xbit_r509_c33 bl[33] br[33] wl[509] vdd gnd cell_6t
Xbit_r510_c33 bl[33] br[33] wl[510] vdd gnd cell_6t
Xbit_r511_c33 bl[33] br[33] wl[511] vdd gnd cell_6t
Xbit_r0_c34 bl[34] br[34] wl[0] vdd gnd cell_6t
Xbit_r1_c34 bl[34] br[34] wl[1] vdd gnd cell_6t
Xbit_r2_c34 bl[34] br[34] wl[2] vdd gnd cell_6t
Xbit_r3_c34 bl[34] br[34] wl[3] vdd gnd cell_6t
Xbit_r4_c34 bl[34] br[34] wl[4] vdd gnd cell_6t
Xbit_r5_c34 bl[34] br[34] wl[5] vdd gnd cell_6t
Xbit_r6_c34 bl[34] br[34] wl[6] vdd gnd cell_6t
Xbit_r7_c34 bl[34] br[34] wl[7] vdd gnd cell_6t
Xbit_r8_c34 bl[34] br[34] wl[8] vdd gnd cell_6t
Xbit_r9_c34 bl[34] br[34] wl[9] vdd gnd cell_6t
Xbit_r10_c34 bl[34] br[34] wl[10] vdd gnd cell_6t
Xbit_r11_c34 bl[34] br[34] wl[11] vdd gnd cell_6t
Xbit_r12_c34 bl[34] br[34] wl[12] vdd gnd cell_6t
Xbit_r13_c34 bl[34] br[34] wl[13] vdd gnd cell_6t
Xbit_r14_c34 bl[34] br[34] wl[14] vdd gnd cell_6t
Xbit_r15_c34 bl[34] br[34] wl[15] vdd gnd cell_6t
Xbit_r16_c34 bl[34] br[34] wl[16] vdd gnd cell_6t
Xbit_r17_c34 bl[34] br[34] wl[17] vdd gnd cell_6t
Xbit_r18_c34 bl[34] br[34] wl[18] vdd gnd cell_6t
Xbit_r19_c34 bl[34] br[34] wl[19] vdd gnd cell_6t
Xbit_r20_c34 bl[34] br[34] wl[20] vdd gnd cell_6t
Xbit_r21_c34 bl[34] br[34] wl[21] vdd gnd cell_6t
Xbit_r22_c34 bl[34] br[34] wl[22] vdd gnd cell_6t
Xbit_r23_c34 bl[34] br[34] wl[23] vdd gnd cell_6t
Xbit_r24_c34 bl[34] br[34] wl[24] vdd gnd cell_6t
Xbit_r25_c34 bl[34] br[34] wl[25] vdd gnd cell_6t
Xbit_r26_c34 bl[34] br[34] wl[26] vdd gnd cell_6t
Xbit_r27_c34 bl[34] br[34] wl[27] vdd gnd cell_6t
Xbit_r28_c34 bl[34] br[34] wl[28] vdd gnd cell_6t
Xbit_r29_c34 bl[34] br[34] wl[29] vdd gnd cell_6t
Xbit_r30_c34 bl[34] br[34] wl[30] vdd gnd cell_6t
Xbit_r31_c34 bl[34] br[34] wl[31] vdd gnd cell_6t
Xbit_r32_c34 bl[34] br[34] wl[32] vdd gnd cell_6t
Xbit_r33_c34 bl[34] br[34] wl[33] vdd gnd cell_6t
Xbit_r34_c34 bl[34] br[34] wl[34] vdd gnd cell_6t
Xbit_r35_c34 bl[34] br[34] wl[35] vdd gnd cell_6t
Xbit_r36_c34 bl[34] br[34] wl[36] vdd gnd cell_6t
Xbit_r37_c34 bl[34] br[34] wl[37] vdd gnd cell_6t
Xbit_r38_c34 bl[34] br[34] wl[38] vdd gnd cell_6t
Xbit_r39_c34 bl[34] br[34] wl[39] vdd gnd cell_6t
Xbit_r40_c34 bl[34] br[34] wl[40] vdd gnd cell_6t
Xbit_r41_c34 bl[34] br[34] wl[41] vdd gnd cell_6t
Xbit_r42_c34 bl[34] br[34] wl[42] vdd gnd cell_6t
Xbit_r43_c34 bl[34] br[34] wl[43] vdd gnd cell_6t
Xbit_r44_c34 bl[34] br[34] wl[44] vdd gnd cell_6t
Xbit_r45_c34 bl[34] br[34] wl[45] vdd gnd cell_6t
Xbit_r46_c34 bl[34] br[34] wl[46] vdd gnd cell_6t
Xbit_r47_c34 bl[34] br[34] wl[47] vdd gnd cell_6t
Xbit_r48_c34 bl[34] br[34] wl[48] vdd gnd cell_6t
Xbit_r49_c34 bl[34] br[34] wl[49] vdd gnd cell_6t
Xbit_r50_c34 bl[34] br[34] wl[50] vdd gnd cell_6t
Xbit_r51_c34 bl[34] br[34] wl[51] vdd gnd cell_6t
Xbit_r52_c34 bl[34] br[34] wl[52] vdd gnd cell_6t
Xbit_r53_c34 bl[34] br[34] wl[53] vdd gnd cell_6t
Xbit_r54_c34 bl[34] br[34] wl[54] vdd gnd cell_6t
Xbit_r55_c34 bl[34] br[34] wl[55] vdd gnd cell_6t
Xbit_r56_c34 bl[34] br[34] wl[56] vdd gnd cell_6t
Xbit_r57_c34 bl[34] br[34] wl[57] vdd gnd cell_6t
Xbit_r58_c34 bl[34] br[34] wl[58] vdd gnd cell_6t
Xbit_r59_c34 bl[34] br[34] wl[59] vdd gnd cell_6t
Xbit_r60_c34 bl[34] br[34] wl[60] vdd gnd cell_6t
Xbit_r61_c34 bl[34] br[34] wl[61] vdd gnd cell_6t
Xbit_r62_c34 bl[34] br[34] wl[62] vdd gnd cell_6t
Xbit_r63_c34 bl[34] br[34] wl[63] vdd gnd cell_6t
Xbit_r64_c34 bl[34] br[34] wl[64] vdd gnd cell_6t
Xbit_r65_c34 bl[34] br[34] wl[65] vdd gnd cell_6t
Xbit_r66_c34 bl[34] br[34] wl[66] vdd gnd cell_6t
Xbit_r67_c34 bl[34] br[34] wl[67] vdd gnd cell_6t
Xbit_r68_c34 bl[34] br[34] wl[68] vdd gnd cell_6t
Xbit_r69_c34 bl[34] br[34] wl[69] vdd gnd cell_6t
Xbit_r70_c34 bl[34] br[34] wl[70] vdd gnd cell_6t
Xbit_r71_c34 bl[34] br[34] wl[71] vdd gnd cell_6t
Xbit_r72_c34 bl[34] br[34] wl[72] vdd gnd cell_6t
Xbit_r73_c34 bl[34] br[34] wl[73] vdd gnd cell_6t
Xbit_r74_c34 bl[34] br[34] wl[74] vdd gnd cell_6t
Xbit_r75_c34 bl[34] br[34] wl[75] vdd gnd cell_6t
Xbit_r76_c34 bl[34] br[34] wl[76] vdd gnd cell_6t
Xbit_r77_c34 bl[34] br[34] wl[77] vdd gnd cell_6t
Xbit_r78_c34 bl[34] br[34] wl[78] vdd gnd cell_6t
Xbit_r79_c34 bl[34] br[34] wl[79] vdd gnd cell_6t
Xbit_r80_c34 bl[34] br[34] wl[80] vdd gnd cell_6t
Xbit_r81_c34 bl[34] br[34] wl[81] vdd gnd cell_6t
Xbit_r82_c34 bl[34] br[34] wl[82] vdd gnd cell_6t
Xbit_r83_c34 bl[34] br[34] wl[83] vdd gnd cell_6t
Xbit_r84_c34 bl[34] br[34] wl[84] vdd gnd cell_6t
Xbit_r85_c34 bl[34] br[34] wl[85] vdd gnd cell_6t
Xbit_r86_c34 bl[34] br[34] wl[86] vdd gnd cell_6t
Xbit_r87_c34 bl[34] br[34] wl[87] vdd gnd cell_6t
Xbit_r88_c34 bl[34] br[34] wl[88] vdd gnd cell_6t
Xbit_r89_c34 bl[34] br[34] wl[89] vdd gnd cell_6t
Xbit_r90_c34 bl[34] br[34] wl[90] vdd gnd cell_6t
Xbit_r91_c34 bl[34] br[34] wl[91] vdd gnd cell_6t
Xbit_r92_c34 bl[34] br[34] wl[92] vdd gnd cell_6t
Xbit_r93_c34 bl[34] br[34] wl[93] vdd gnd cell_6t
Xbit_r94_c34 bl[34] br[34] wl[94] vdd gnd cell_6t
Xbit_r95_c34 bl[34] br[34] wl[95] vdd gnd cell_6t
Xbit_r96_c34 bl[34] br[34] wl[96] vdd gnd cell_6t
Xbit_r97_c34 bl[34] br[34] wl[97] vdd gnd cell_6t
Xbit_r98_c34 bl[34] br[34] wl[98] vdd gnd cell_6t
Xbit_r99_c34 bl[34] br[34] wl[99] vdd gnd cell_6t
Xbit_r100_c34 bl[34] br[34] wl[100] vdd gnd cell_6t
Xbit_r101_c34 bl[34] br[34] wl[101] vdd gnd cell_6t
Xbit_r102_c34 bl[34] br[34] wl[102] vdd gnd cell_6t
Xbit_r103_c34 bl[34] br[34] wl[103] vdd gnd cell_6t
Xbit_r104_c34 bl[34] br[34] wl[104] vdd gnd cell_6t
Xbit_r105_c34 bl[34] br[34] wl[105] vdd gnd cell_6t
Xbit_r106_c34 bl[34] br[34] wl[106] vdd gnd cell_6t
Xbit_r107_c34 bl[34] br[34] wl[107] vdd gnd cell_6t
Xbit_r108_c34 bl[34] br[34] wl[108] vdd gnd cell_6t
Xbit_r109_c34 bl[34] br[34] wl[109] vdd gnd cell_6t
Xbit_r110_c34 bl[34] br[34] wl[110] vdd gnd cell_6t
Xbit_r111_c34 bl[34] br[34] wl[111] vdd gnd cell_6t
Xbit_r112_c34 bl[34] br[34] wl[112] vdd gnd cell_6t
Xbit_r113_c34 bl[34] br[34] wl[113] vdd gnd cell_6t
Xbit_r114_c34 bl[34] br[34] wl[114] vdd gnd cell_6t
Xbit_r115_c34 bl[34] br[34] wl[115] vdd gnd cell_6t
Xbit_r116_c34 bl[34] br[34] wl[116] vdd gnd cell_6t
Xbit_r117_c34 bl[34] br[34] wl[117] vdd gnd cell_6t
Xbit_r118_c34 bl[34] br[34] wl[118] vdd gnd cell_6t
Xbit_r119_c34 bl[34] br[34] wl[119] vdd gnd cell_6t
Xbit_r120_c34 bl[34] br[34] wl[120] vdd gnd cell_6t
Xbit_r121_c34 bl[34] br[34] wl[121] vdd gnd cell_6t
Xbit_r122_c34 bl[34] br[34] wl[122] vdd gnd cell_6t
Xbit_r123_c34 bl[34] br[34] wl[123] vdd gnd cell_6t
Xbit_r124_c34 bl[34] br[34] wl[124] vdd gnd cell_6t
Xbit_r125_c34 bl[34] br[34] wl[125] vdd gnd cell_6t
Xbit_r126_c34 bl[34] br[34] wl[126] vdd gnd cell_6t
Xbit_r127_c34 bl[34] br[34] wl[127] vdd gnd cell_6t
Xbit_r128_c34 bl[34] br[34] wl[128] vdd gnd cell_6t
Xbit_r129_c34 bl[34] br[34] wl[129] vdd gnd cell_6t
Xbit_r130_c34 bl[34] br[34] wl[130] vdd gnd cell_6t
Xbit_r131_c34 bl[34] br[34] wl[131] vdd gnd cell_6t
Xbit_r132_c34 bl[34] br[34] wl[132] vdd gnd cell_6t
Xbit_r133_c34 bl[34] br[34] wl[133] vdd gnd cell_6t
Xbit_r134_c34 bl[34] br[34] wl[134] vdd gnd cell_6t
Xbit_r135_c34 bl[34] br[34] wl[135] vdd gnd cell_6t
Xbit_r136_c34 bl[34] br[34] wl[136] vdd gnd cell_6t
Xbit_r137_c34 bl[34] br[34] wl[137] vdd gnd cell_6t
Xbit_r138_c34 bl[34] br[34] wl[138] vdd gnd cell_6t
Xbit_r139_c34 bl[34] br[34] wl[139] vdd gnd cell_6t
Xbit_r140_c34 bl[34] br[34] wl[140] vdd gnd cell_6t
Xbit_r141_c34 bl[34] br[34] wl[141] vdd gnd cell_6t
Xbit_r142_c34 bl[34] br[34] wl[142] vdd gnd cell_6t
Xbit_r143_c34 bl[34] br[34] wl[143] vdd gnd cell_6t
Xbit_r144_c34 bl[34] br[34] wl[144] vdd gnd cell_6t
Xbit_r145_c34 bl[34] br[34] wl[145] vdd gnd cell_6t
Xbit_r146_c34 bl[34] br[34] wl[146] vdd gnd cell_6t
Xbit_r147_c34 bl[34] br[34] wl[147] vdd gnd cell_6t
Xbit_r148_c34 bl[34] br[34] wl[148] vdd gnd cell_6t
Xbit_r149_c34 bl[34] br[34] wl[149] vdd gnd cell_6t
Xbit_r150_c34 bl[34] br[34] wl[150] vdd gnd cell_6t
Xbit_r151_c34 bl[34] br[34] wl[151] vdd gnd cell_6t
Xbit_r152_c34 bl[34] br[34] wl[152] vdd gnd cell_6t
Xbit_r153_c34 bl[34] br[34] wl[153] vdd gnd cell_6t
Xbit_r154_c34 bl[34] br[34] wl[154] vdd gnd cell_6t
Xbit_r155_c34 bl[34] br[34] wl[155] vdd gnd cell_6t
Xbit_r156_c34 bl[34] br[34] wl[156] vdd gnd cell_6t
Xbit_r157_c34 bl[34] br[34] wl[157] vdd gnd cell_6t
Xbit_r158_c34 bl[34] br[34] wl[158] vdd gnd cell_6t
Xbit_r159_c34 bl[34] br[34] wl[159] vdd gnd cell_6t
Xbit_r160_c34 bl[34] br[34] wl[160] vdd gnd cell_6t
Xbit_r161_c34 bl[34] br[34] wl[161] vdd gnd cell_6t
Xbit_r162_c34 bl[34] br[34] wl[162] vdd gnd cell_6t
Xbit_r163_c34 bl[34] br[34] wl[163] vdd gnd cell_6t
Xbit_r164_c34 bl[34] br[34] wl[164] vdd gnd cell_6t
Xbit_r165_c34 bl[34] br[34] wl[165] vdd gnd cell_6t
Xbit_r166_c34 bl[34] br[34] wl[166] vdd gnd cell_6t
Xbit_r167_c34 bl[34] br[34] wl[167] vdd gnd cell_6t
Xbit_r168_c34 bl[34] br[34] wl[168] vdd gnd cell_6t
Xbit_r169_c34 bl[34] br[34] wl[169] vdd gnd cell_6t
Xbit_r170_c34 bl[34] br[34] wl[170] vdd gnd cell_6t
Xbit_r171_c34 bl[34] br[34] wl[171] vdd gnd cell_6t
Xbit_r172_c34 bl[34] br[34] wl[172] vdd gnd cell_6t
Xbit_r173_c34 bl[34] br[34] wl[173] vdd gnd cell_6t
Xbit_r174_c34 bl[34] br[34] wl[174] vdd gnd cell_6t
Xbit_r175_c34 bl[34] br[34] wl[175] vdd gnd cell_6t
Xbit_r176_c34 bl[34] br[34] wl[176] vdd gnd cell_6t
Xbit_r177_c34 bl[34] br[34] wl[177] vdd gnd cell_6t
Xbit_r178_c34 bl[34] br[34] wl[178] vdd gnd cell_6t
Xbit_r179_c34 bl[34] br[34] wl[179] vdd gnd cell_6t
Xbit_r180_c34 bl[34] br[34] wl[180] vdd gnd cell_6t
Xbit_r181_c34 bl[34] br[34] wl[181] vdd gnd cell_6t
Xbit_r182_c34 bl[34] br[34] wl[182] vdd gnd cell_6t
Xbit_r183_c34 bl[34] br[34] wl[183] vdd gnd cell_6t
Xbit_r184_c34 bl[34] br[34] wl[184] vdd gnd cell_6t
Xbit_r185_c34 bl[34] br[34] wl[185] vdd gnd cell_6t
Xbit_r186_c34 bl[34] br[34] wl[186] vdd gnd cell_6t
Xbit_r187_c34 bl[34] br[34] wl[187] vdd gnd cell_6t
Xbit_r188_c34 bl[34] br[34] wl[188] vdd gnd cell_6t
Xbit_r189_c34 bl[34] br[34] wl[189] vdd gnd cell_6t
Xbit_r190_c34 bl[34] br[34] wl[190] vdd gnd cell_6t
Xbit_r191_c34 bl[34] br[34] wl[191] vdd gnd cell_6t
Xbit_r192_c34 bl[34] br[34] wl[192] vdd gnd cell_6t
Xbit_r193_c34 bl[34] br[34] wl[193] vdd gnd cell_6t
Xbit_r194_c34 bl[34] br[34] wl[194] vdd gnd cell_6t
Xbit_r195_c34 bl[34] br[34] wl[195] vdd gnd cell_6t
Xbit_r196_c34 bl[34] br[34] wl[196] vdd gnd cell_6t
Xbit_r197_c34 bl[34] br[34] wl[197] vdd gnd cell_6t
Xbit_r198_c34 bl[34] br[34] wl[198] vdd gnd cell_6t
Xbit_r199_c34 bl[34] br[34] wl[199] vdd gnd cell_6t
Xbit_r200_c34 bl[34] br[34] wl[200] vdd gnd cell_6t
Xbit_r201_c34 bl[34] br[34] wl[201] vdd gnd cell_6t
Xbit_r202_c34 bl[34] br[34] wl[202] vdd gnd cell_6t
Xbit_r203_c34 bl[34] br[34] wl[203] vdd gnd cell_6t
Xbit_r204_c34 bl[34] br[34] wl[204] vdd gnd cell_6t
Xbit_r205_c34 bl[34] br[34] wl[205] vdd gnd cell_6t
Xbit_r206_c34 bl[34] br[34] wl[206] vdd gnd cell_6t
Xbit_r207_c34 bl[34] br[34] wl[207] vdd gnd cell_6t
Xbit_r208_c34 bl[34] br[34] wl[208] vdd gnd cell_6t
Xbit_r209_c34 bl[34] br[34] wl[209] vdd gnd cell_6t
Xbit_r210_c34 bl[34] br[34] wl[210] vdd gnd cell_6t
Xbit_r211_c34 bl[34] br[34] wl[211] vdd gnd cell_6t
Xbit_r212_c34 bl[34] br[34] wl[212] vdd gnd cell_6t
Xbit_r213_c34 bl[34] br[34] wl[213] vdd gnd cell_6t
Xbit_r214_c34 bl[34] br[34] wl[214] vdd gnd cell_6t
Xbit_r215_c34 bl[34] br[34] wl[215] vdd gnd cell_6t
Xbit_r216_c34 bl[34] br[34] wl[216] vdd gnd cell_6t
Xbit_r217_c34 bl[34] br[34] wl[217] vdd gnd cell_6t
Xbit_r218_c34 bl[34] br[34] wl[218] vdd gnd cell_6t
Xbit_r219_c34 bl[34] br[34] wl[219] vdd gnd cell_6t
Xbit_r220_c34 bl[34] br[34] wl[220] vdd gnd cell_6t
Xbit_r221_c34 bl[34] br[34] wl[221] vdd gnd cell_6t
Xbit_r222_c34 bl[34] br[34] wl[222] vdd gnd cell_6t
Xbit_r223_c34 bl[34] br[34] wl[223] vdd gnd cell_6t
Xbit_r224_c34 bl[34] br[34] wl[224] vdd gnd cell_6t
Xbit_r225_c34 bl[34] br[34] wl[225] vdd gnd cell_6t
Xbit_r226_c34 bl[34] br[34] wl[226] vdd gnd cell_6t
Xbit_r227_c34 bl[34] br[34] wl[227] vdd gnd cell_6t
Xbit_r228_c34 bl[34] br[34] wl[228] vdd gnd cell_6t
Xbit_r229_c34 bl[34] br[34] wl[229] vdd gnd cell_6t
Xbit_r230_c34 bl[34] br[34] wl[230] vdd gnd cell_6t
Xbit_r231_c34 bl[34] br[34] wl[231] vdd gnd cell_6t
Xbit_r232_c34 bl[34] br[34] wl[232] vdd gnd cell_6t
Xbit_r233_c34 bl[34] br[34] wl[233] vdd gnd cell_6t
Xbit_r234_c34 bl[34] br[34] wl[234] vdd gnd cell_6t
Xbit_r235_c34 bl[34] br[34] wl[235] vdd gnd cell_6t
Xbit_r236_c34 bl[34] br[34] wl[236] vdd gnd cell_6t
Xbit_r237_c34 bl[34] br[34] wl[237] vdd gnd cell_6t
Xbit_r238_c34 bl[34] br[34] wl[238] vdd gnd cell_6t
Xbit_r239_c34 bl[34] br[34] wl[239] vdd gnd cell_6t
Xbit_r240_c34 bl[34] br[34] wl[240] vdd gnd cell_6t
Xbit_r241_c34 bl[34] br[34] wl[241] vdd gnd cell_6t
Xbit_r242_c34 bl[34] br[34] wl[242] vdd gnd cell_6t
Xbit_r243_c34 bl[34] br[34] wl[243] vdd gnd cell_6t
Xbit_r244_c34 bl[34] br[34] wl[244] vdd gnd cell_6t
Xbit_r245_c34 bl[34] br[34] wl[245] vdd gnd cell_6t
Xbit_r246_c34 bl[34] br[34] wl[246] vdd gnd cell_6t
Xbit_r247_c34 bl[34] br[34] wl[247] vdd gnd cell_6t
Xbit_r248_c34 bl[34] br[34] wl[248] vdd gnd cell_6t
Xbit_r249_c34 bl[34] br[34] wl[249] vdd gnd cell_6t
Xbit_r250_c34 bl[34] br[34] wl[250] vdd gnd cell_6t
Xbit_r251_c34 bl[34] br[34] wl[251] vdd gnd cell_6t
Xbit_r252_c34 bl[34] br[34] wl[252] vdd gnd cell_6t
Xbit_r253_c34 bl[34] br[34] wl[253] vdd gnd cell_6t
Xbit_r254_c34 bl[34] br[34] wl[254] vdd gnd cell_6t
Xbit_r255_c34 bl[34] br[34] wl[255] vdd gnd cell_6t
Xbit_r256_c34 bl[34] br[34] wl[256] vdd gnd cell_6t
Xbit_r257_c34 bl[34] br[34] wl[257] vdd gnd cell_6t
Xbit_r258_c34 bl[34] br[34] wl[258] vdd gnd cell_6t
Xbit_r259_c34 bl[34] br[34] wl[259] vdd gnd cell_6t
Xbit_r260_c34 bl[34] br[34] wl[260] vdd gnd cell_6t
Xbit_r261_c34 bl[34] br[34] wl[261] vdd gnd cell_6t
Xbit_r262_c34 bl[34] br[34] wl[262] vdd gnd cell_6t
Xbit_r263_c34 bl[34] br[34] wl[263] vdd gnd cell_6t
Xbit_r264_c34 bl[34] br[34] wl[264] vdd gnd cell_6t
Xbit_r265_c34 bl[34] br[34] wl[265] vdd gnd cell_6t
Xbit_r266_c34 bl[34] br[34] wl[266] vdd gnd cell_6t
Xbit_r267_c34 bl[34] br[34] wl[267] vdd gnd cell_6t
Xbit_r268_c34 bl[34] br[34] wl[268] vdd gnd cell_6t
Xbit_r269_c34 bl[34] br[34] wl[269] vdd gnd cell_6t
Xbit_r270_c34 bl[34] br[34] wl[270] vdd gnd cell_6t
Xbit_r271_c34 bl[34] br[34] wl[271] vdd gnd cell_6t
Xbit_r272_c34 bl[34] br[34] wl[272] vdd gnd cell_6t
Xbit_r273_c34 bl[34] br[34] wl[273] vdd gnd cell_6t
Xbit_r274_c34 bl[34] br[34] wl[274] vdd gnd cell_6t
Xbit_r275_c34 bl[34] br[34] wl[275] vdd gnd cell_6t
Xbit_r276_c34 bl[34] br[34] wl[276] vdd gnd cell_6t
Xbit_r277_c34 bl[34] br[34] wl[277] vdd gnd cell_6t
Xbit_r278_c34 bl[34] br[34] wl[278] vdd gnd cell_6t
Xbit_r279_c34 bl[34] br[34] wl[279] vdd gnd cell_6t
Xbit_r280_c34 bl[34] br[34] wl[280] vdd gnd cell_6t
Xbit_r281_c34 bl[34] br[34] wl[281] vdd gnd cell_6t
Xbit_r282_c34 bl[34] br[34] wl[282] vdd gnd cell_6t
Xbit_r283_c34 bl[34] br[34] wl[283] vdd gnd cell_6t
Xbit_r284_c34 bl[34] br[34] wl[284] vdd gnd cell_6t
Xbit_r285_c34 bl[34] br[34] wl[285] vdd gnd cell_6t
Xbit_r286_c34 bl[34] br[34] wl[286] vdd gnd cell_6t
Xbit_r287_c34 bl[34] br[34] wl[287] vdd gnd cell_6t
Xbit_r288_c34 bl[34] br[34] wl[288] vdd gnd cell_6t
Xbit_r289_c34 bl[34] br[34] wl[289] vdd gnd cell_6t
Xbit_r290_c34 bl[34] br[34] wl[290] vdd gnd cell_6t
Xbit_r291_c34 bl[34] br[34] wl[291] vdd gnd cell_6t
Xbit_r292_c34 bl[34] br[34] wl[292] vdd gnd cell_6t
Xbit_r293_c34 bl[34] br[34] wl[293] vdd gnd cell_6t
Xbit_r294_c34 bl[34] br[34] wl[294] vdd gnd cell_6t
Xbit_r295_c34 bl[34] br[34] wl[295] vdd gnd cell_6t
Xbit_r296_c34 bl[34] br[34] wl[296] vdd gnd cell_6t
Xbit_r297_c34 bl[34] br[34] wl[297] vdd gnd cell_6t
Xbit_r298_c34 bl[34] br[34] wl[298] vdd gnd cell_6t
Xbit_r299_c34 bl[34] br[34] wl[299] vdd gnd cell_6t
Xbit_r300_c34 bl[34] br[34] wl[300] vdd gnd cell_6t
Xbit_r301_c34 bl[34] br[34] wl[301] vdd gnd cell_6t
Xbit_r302_c34 bl[34] br[34] wl[302] vdd gnd cell_6t
Xbit_r303_c34 bl[34] br[34] wl[303] vdd gnd cell_6t
Xbit_r304_c34 bl[34] br[34] wl[304] vdd gnd cell_6t
Xbit_r305_c34 bl[34] br[34] wl[305] vdd gnd cell_6t
Xbit_r306_c34 bl[34] br[34] wl[306] vdd gnd cell_6t
Xbit_r307_c34 bl[34] br[34] wl[307] vdd gnd cell_6t
Xbit_r308_c34 bl[34] br[34] wl[308] vdd gnd cell_6t
Xbit_r309_c34 bl[34] br[34] wl[309] vdd gnd cell_6t
Xbit_r310_c34 bl[34] br[34] wl[310] vdd gnd cell_6t
Xbit_r311_c34 bl[34] br[34] wl[311] vdd gnd cell_6t
Xbit_r312_c34 bl[34] br[34] wl[312] vdd gnd cell_6t
Xbit_r313_c34 bl[34] br[34] wl[313] vdd gnd cell_6t
Xbit_r314_c34 bl[34] br[34] wl[314] vdd gnd cell_6t
Xbit_r315_c34 bl[34] br[34] wl[315] vdd gnd cell_6t
Xbit_r316_c34 bl[34] br[34] wl[316] vdd gnd cell_6t
Xbit_r317_c34 bl[34] br[34] wl[317] vdd gnd cell_6t
Xbit_r318_c34 bl[34] br[34] wl[318] vdd gnd cell_6t
Xbit_r319_c34 bl[34] br[34] wl[319] vdd gnd cell_6t
Xbit_r320_c34 bl[34] br[34] wl[320] vdd gnd cell_6t
Xbit_r321_c34 bl[34] br[34] wl[321] vdd gnd cell_6t
Xbit_r322_c34 bl[34] br[34] wl[322] vdd gnd cell_6t
Xbit_r323_c34 bl[34] br[34] wl[323] vdd gnd cell_6t
Xbit_r324_c34 bl[34] br[34] wl[324] vdd gnd cell_6t
Xbit_r325_c34 bl[34] br[34] wl[325] vdd gnd cell_6t
Xbit_r326_c34 bl[34] br[34] wl[326] vdd gnd cell_6t
Xbit_r327_c34 bl[34] br[34] wl[327] vdd gnd cell_6t
Xbit_r328_c34 bl[34] br[34] wl[328] vdd gnd cell_6t
Xbit_r329_c34 bl[34] br[34] wl[329] vdd gnd cell_6t
Xbit_r330_c34 bl[34] br[34] wl[330] vdd gnd cell_6t
Xbit_r331_c34 bl[34] br[34] wl[331] vdd gnd cell_6t
Xbit_r332_c34 bl[34] br[34] wl[332] vdd gnd cell_6t
Xbit_r333_c34 bl[34] br[34] wl[333] vdd gnd cell_6t
Xbit_r334_c34 bl[34] br[34] wl[334] vdd gnd cell_6t
Xbit_r335_c34 bl[34] br[34] wl[335] vdd gnd cell_6t
Xbit_r336_c34 bl[34] br[34] wl[336] vdd gnd cell_6t
Xbit_r337_c34 bl[34] br[34] wl[337] vdd gnd cell_6t
Xbit_r338_c34 bl[34] br[34] wl[338] vdd gnd cell_6t
Xbit_r339_c34 bl[34] br[34] wl[339] vdd gnd cell_6t
Xbit_r340_c34 bl[34] br[34] wl[340] vdd gnd cell_6t
Xbit_r341_c34 bl[34] br[34] wl[341] vdd gnd cell_6t
Xbit_r342_c34 bl[34] br[34] wl[342] vdd gnd cell_6t
Xbit_r343_c34 bl[34] br[34] wl[343] vdd gnd cell_6t
Xbit_r344_c34 bl[34] br[34] wl[344] vdd gnd cell_6t
Xbit_r345_c34 bl[34] br[34] wl[345] vdd gnd cell_6t
Xbit_r346_c34 bl[34] br[34] wl[346] vdd gnd cell_6t
Xbit_r347_c34 bl[34] br[34] wl[347] vdd gnd cell_6t
Xbit_r348_c34 bl[34] br[34] wl[348] vdd gnd cell_6t
Xbit_r349_c34 bl[34] br[34] wl[349] vdd gnd cell_6t
Xbit_r350_c34 bl[34] br[34] wl[350] vdd gnd cell_6t
Xbit_r351_c34 bl[34] br[34] wl[351] vdd gnd cell_6t
Xbit_r352_c34 bl[34] br[34] wl[352] vdd gnd cell_6t
Xbit_r353_c34 bl[34] br[34] wl[353] vdd gnd cell_6t
Xbit_r354_c34 bl[34] br[34] wl[354] vdd gnd cell_6t
Xbit_r355_c34 bl[34] br[34] wl[355] vdd gnd cell_6t
Xbit_r356_c34 bl[34] br[34] wl[356] vdd gnd cell_6t
Xbit_r357_c34 bl[34] br[34] wl[357] vdd gnd cell_6t
Xbit_r358_c34 bl[34] br[34] wl[358] vdd gnd cell_6t
Xbit_r359_c34 bl[34] br[34] wl[359] vdd gnd cell_6t
Xbit_r360_c34 bl[34] br[34] wl[360] vdd gnd cell_6t
Xbit_r361_c34 bl[34] br[34] wl[361] vdd gnd cell_6t
Xbit_r362_c34 bl[34] br[34] wl[362] vdd gnd cell_6t
Xbit_r363_c34 bl[34] br[34] wl[363] vdd gnd cell_6t
Xbit_r364_c34 bl[34] br[34] wl[364] vdd gnd cell_6t
Xbit_r365_c34 bl[34] br[34] wl[365] vdd gnd cell_6t
Xbit_r366_c34 bl[34] br[34] wl[366] vdd gnd cell_6t
Xbit_r367_c34 bl[34] br[34] wl[367] vdd gnd cell_6t
Xbit_r368_c34 bl[34] br[34] wl[368] vdd gnd cell_6t
Xbit_r369_c34 bl[34] br[34] wl[369] vdd gnd cell_6t
Xbit_r370_c34 bl[34] br[34] wl[370] vdd gnd cell_6t
Xbit_r371_c34 bl[34] br[34] wl[371] vdd gnd cell_6t
Xbit_r372_c34 bl[34] br[34] wl[372] vdd gnd cell_6t
Xbit_r373_c34 bl[34] br[34] wl[373] vdd gnd cell_6t
Xbit_r374_c34 bl[34] br[34] wl[374] vdd gnd cell_6t
Xbit_r375_c34 bl[34] br[34] wl[375] vdd gnd cell_6t
Xbit_r376_c34 bl[34] br[34] wl[376] vdd gnd cell_6t
Xbit_r377_c34 bl[34] br[34] wl[377] vdd gnd cell_6t
Xbit_r378_c34 bl[34] br[34] wl[378] vdd gnd cell_6t
Xbit_r379_c34 bl[34] br[34] wl[379] vdd gnd cell_6t
Xbit_r380_c34 bl[34] br[34] wl[380] vdd gnd cell_6t
Xbit_r381_c34 bl[34] br[34] wl[381] vdd gnd cell_6t
Xbit_r382_c34 bl[34] br[34] wl[382] vdd gnd cell_6t
Xbit_r383_c34 bl[34] br[34] wl[383] vdd gnd cell_6t
Xbit_r384_c34 bl[34] br[34] wl[384] vdd gnd cell_6t
Xbit_r385_c34 bl[34] br[34] wl[385] vdd gnd cell_6t
Xbit_r386_c34 bl[34] br[34] wl[386] vdd gnd cell_6t
Xbit_r387_c34 bl[34] br[34] wl[387] vdd gnd cell_6t
Xbit_r388_c34 bl[34] br[34] wl[388] vdd gnd cell_6t
Xbit_r389_c34 bl[34] br[34] wl[389] vdd gnd cell_6t
Xbit_r390_c34 bl[34] br[34] wl[390] vdd gnd cell_6t
Xbit_r391_c34 bl[34] br[34] wl[391] vdd gnd cell_6t
Xbit_r392_c34 bl[34] br[34] wl[392] vdd gnd cell_6t
Xbit_r393_c34 bl[34] br[34] wl[393] vdd gnd cell_6t
Xbit_r394_c34 bl[34] br[34] wl[394] vdd gnd cell_6t
Xbit_r395_c34 bl[34] br[34] wl[395] vdd gnd cell_6t
Xbit_r396_c34 bl[34] br[34] wl[396] vdd gnd cell_6t
Xbit_r397_c34 bl[34] br[34] wl[397] vdd gnd cell_6t
Xbit_r398_c34 bl[34] br[34] wl[398] vdd gnd cell_6t
Xbit_r399_c34 bl[34] br[34] wl[399] vdd gnd cell_6t
Xbit_r400_c34 bl[34] br[34] wl[400] vdd gnd cell_6t
Xbit_r401_c34 bl[34] br[34] wl[401] vdd gnd cell_6t
Xbit_r402_c34 bl[34] br[34] wl[402] vdd gnd cell_6t
Xbit_r403_c34 bl[34] br[34] wl[403] vdd gnd cell_6t
Xbit_r404_c34 bl[34] br[34] wl[404] vdd gnd cell_6t
Xbit_r405_c34 bl[34] br[34] wl[405] vdd gnd cell_6t
Xbit_r406_c34 bl[34] br[34] wl[406] vdd gnd cell_6t
Xbit_r407_c34 bl[34] br[34] wl[407] vdd gnd cell_6t
Xbit_r408_c34 bl[34] br[34] wl[408] vdd gnd cell_6t
Xbit_r409_c34 bl[34] br[34] wl[409] vdd gnd cell_6t
Xbit_r410_c34 bl[34] br[34] wl[410] vdd gnd cell_6t
Xbit_r411_c34 bl[34] br[34] wl[411] vdd gnd cell_6t
Xbit_r412_c34 bl[34] br[34] wl[412] vdd gnd cell_6t
Xbit_r413_c34 bl[34] br[34] wl[413] vdd gnd cell_6t
Xbit_r414_c34 bl[34] br[34] wl[414] vdd gnd cell_6t
Xbit_r415_c34 bl[34] br[34] wl[415] vdd gnd cell_6t
Xbit_r416_c34 bl[34] br[34] wl[416] vdd gnd cell_6t
Xbit_r417_c34 bl[34] br[34] wl[417] vdd gnd cell_6t
Xbit_r418_c34 bl[34] br[34] wl[418] vdd gnd cell_6t
Xbit_r419_c34 bl[34] br[34] wl[419] vdd gnd cell_6t
Xbit_r420_c34 bl[34] br[34] wl[420] vdd gnd cell_6t
Xbit_r421_c34 bl[34] br[34] wl[421] vdd gnd cell_6t
Xbit_r422_c34 bl[34] br[34] wl[422] vdd gnd cell_6t
Xbit_r423_c34 bl[34] br[34] wl[423] vdd gnd cell_6t
Xbit_r424_c34 bl[34] br[34] wl[424] vdd gnd cell_6t
Xbit_r425_c34 bl[34] br[34] wl[425] vdd gnd cell_6t
Xbit_r426_c34 bl[34] br[34] wl[426] vdd gnd cell_6t
Xbit_r427_c34 bl[34] br[34] wl[427] vdd gnd cell_6t
Xbit_r428_c34 bl[34] br[34] wl[428] vdd gnd cell_6t
Xbit_r429_c34 bl[34] br[34] wl[429] vdd gnd cell_6t
Xbit_r430_c34 bl[34] br[34] wl[430] vdd gnd cell_6t
Xbit_r431_c34 bl[34] br[34] wl[431] vdd gnd cell_6t
Xbit_r432_c34 bl[34] br[34] wl[432] vdd gnd cell_6t
Xbit_r433_c34 bl[34] br[34] wl[433] vdd gnd cell_6t
Xbit_r434_c34 bl[34] br[34] wl[434] vdd gnd cell_6t
Xbit_r435_c34 bl[34] br[34] wl[435] vdd gnd cell_6t
Xbit_r436_c34 bl[34] br[34] wl[436] vdd gnd cell_6t
Xbit_r437_c34 bl[34] br[34] wl[437] vdd gnd cell_6t
Xbit_r438_c34 bl[34] br[34] wl[438] vdd gnd cell_6t
Xbit_r439_c34 bl[34] br[34] wl[439] vdd gnd cell_6t
Xbit_r440_c34 bl[34] br[34] wl[440] vdd gnd cell_6t
Xbit_r441_c34 bl[34] br[34] wl[441] vdd gnd cell_6t
Xbit_r442_c34 bl[34] br[34] wl[442] vdd gnd cell_6t
Xbit_r443_c34 bl[34] br[34] wl[443] vdd gnd cell_6t
Xbit_r444_c34 bl[34] br[34] wl[444] vdd gnd cell_6t
Xbit_r445_c34 bl[34] br[34] wl[445] vdd gnd cell_6t
Xbit_r446_c34 bl[34] br[34] wl[446] vdd gnd cell_6t
Xbit_r447_c34 bl[34] br[34] wl[447] vdd gnd cell_6t
Xbit_r448_c34 bl[34] br[34] wl[448] vdd gnd cell_6t
Xbit_r449_c34 bl[34] br[34] wl[449] vdd gnd cell_6t
Xbit_r450_c34 bl[34] br[34] wl[450] vdd gnd cell_6t
Xbit_r451_c34 bl[34] br[34] wl[451] vdd gnd cell_6t
Xbit_r452_c34 bl[34] br[34] wl[452] vdd gnd cell_6t
Xbit_r453_c34 bl[34] br[34] wl[453] vdd gnd cell_6t
Xbit_r454_c34 bl[34] br[34] wl[454] vdd gnd cell_6t
Xbit_r455_c34 bl[34] br[34] wl[455] vdd gnd cell_6t
Xbit_r456_c34 bl[34] br[34] wl[456] vdd gnd cell_6t
Xbit_r457_c34 bl[34] br[34] wl[457] vdd gnd cell_6t
Xbit_r458_c34 bl[34] br[34] wl[458] vdd gnd cell_6t
Xbit_r459_c34 bl[34] br[34] wl[459] vdd gnd cell_6t
Xbit_r460_c34 bl[34] br[34] wl[460] vdd gnd cell_6t
Xbit_r461_c34 bl[34] br[34] wl[461] vdd gnd cell_6t
Xbit_r462_c34 bl[34] br[34] wl[462] vdd gnd cell_6t
Xbit_r463_c34 bl[34] br[34] wl[463] vdd gnd cell_6t
Xbit_r464_c34 bl[34] br[34] wl[464] vdd gnd cell_6t
Xbit_r465_c34 bl[34] br[34] wl[465] vdd gnd cell_6t
Xbit_r466_c34 bl[34] br[34] wl[466] vdd gnd cell_6t
Xbit_r467_c34 bl[34] br[34] wl[467] vdd gnd cell_6t
Xbit_r468_c34 bl[34] br[34] wl[468] vdd gnd cell_6t
Xbit_r469_c34 bl[34] br[34] wl[469] vdd gnd cell_6t
Xbit_r470_c34 bl[34] br[34] wl[470] vdd gnd cell_6t
Xbit_r471_c34 bl[34] br[34] wl[471] vdd gnd cell_6t
Xbit_r472_c34 bl[34] br[34] wl[472] vdd gnd cell_6t
Xbit_r473_c34 bl[34] br[34] wl[473] vdd gnd cell_6t
Xbit_r474_c34 bl[34] br[34] wl[474] vdd gnd cell_6t
Xbit_r475_c34 bl[34] br[34] wl[475] vdd gnd cell_6t
Xbit_r476_c34 bl[34] br[34] wl[476] vdd gnd cell_6t
Xbit_r477_c34 bl[34] br[34] wl[477] vdd gnd cell_6t
Xbit_r478_c34 bl[34] br[34] wl[478] vdd gnd cell_6t
Xbit_r479_c34 bl[34] br[34] wl[479] vdd gnd cell_6t
Xbit_r480_c34 bl[34] br[34] wl[480] vdd gnd cell_6t
Xbit_r481_c34 bl[34] br[34] wl[481] vdd gnd cell_6t
Xbit_r482_c34 bl[34] br[34] wl[482] vdd gnd cell_6t
Xbit_r483_c34 bl[34] br[34] wl[483] vdd gnd cell_6t
Xbit_r484_c34 bl[34] br[34] wl[484] vdd gnd cell_6t
Xbit_r485_c34 bl[34] br[34] wl[485] vdd gnd cell_6t
Xbit_r486_c34 bl[34] br[34] wl[486] vdd gnd cell_6t
Xbit_r487_c34 bl[34] br[34] wl[487] vdd gnd cell_6t
Xbit_r488_c34 bl[34] br[34] wl[488] vdd gnd cell_6t
Xbit_r489_c34 bl[34] br[34] wl[489] vdd gnd cell_6t
Xbit_r490_c34 bl[34] br[34] wl[490] vdd gnd cell_6t
Xbit_r491_c34 bl[34] br[34] wl[491] vdd gnd cell_6t
Xbit_r492_c34 bl[34] br[34] wl[492] vdd gnd cell_6t
Xbit_r493_c34 bl[34] br[34] wl[493] vdd gnd cell_6t
Xbit_r494_c34 bl[34] br[34] wl[494] vdd gnd cell_6t
Xbit_r495_c34 bl[34] br[34] wl[495] vdd gnd cell_6t
Xbit_r496_c34 bl[34] br[34] wl[496] vdd gnd cell_6t
Xbit_r497_c34 bl[34] br[34] wl[497] vdd gnd cell_6t
Xbit_r498_c34 bl[34] br[34] wl[498] vdd gnd cell_6t
Xbit_r499_c34 bl[34] br[34] wl[499] vdd gnd cell_6t
Xbit_r500_c34 bl[34] br[34] wl[500] vdd gnd cell_6t
Xbit_r501_c34 bl[34] br[34] wl[501] vdd gnd cell_6t
Xbit_r502_c34 bl[34] br[34] wl[502] vdd gnd cell_6t
Xbit_r503_c34 bl[34] br[34] wl[503] vdd gnd cell_6t
Xbit_r504_c34 bl[34] br[34] wl[504] vdd gnd cell_6t
Xbit_r505_c34 bl[34] br[34] wl[505] vdd gnd cell_6t
Xbit_r506_c34 bl[34] br[34] wl[506] vdd gnd cell_6t
Xbit_r507_c34 bl[34] br[34] wl[507] vdd gnd cell_6t
Xbit_r508_c34 bl[34] br[34] wl[508] vdd gnd cell_6t
Xbit_r509_c34 bl[34] br[34] wl[509] vdd gnd cell_6t
Xbit_r510_c34 bl[34] br[34] wl[510] vdd gnd cell_6t
Xbit_r511_c34 bl[34] br[34] wl[511] vdd gnd cell_6t
Xbit_r0_c35 bl[35] br[35] wl[0] vdd gnd cell_6t
Xbit_r1_c35 bl[35] br[35] wl[1] vdd gnd cell_6t
Xbit_r2_c35 bl[35] br[35] wl[2] vdd gnd cell_6t
Xbit_r3_c35 bl[35] br[35] wl[3] vdd gnd cell_6t
Xbit_r4_c35 bl[35] br[35] wl[4] vdd gnd cell_6t
Xbit_r5_c35 bl[35] br[35] wl[5] vdd gnd cell_6t
Xbit_r6_c35 bl[35] br[35] wl[6] vdd gnd cell_6t
Xbit_r7_c35 bl[35] br[35] wl[7] vdd gnd cell_6t
Xbit_r8_c35 bl[35] br[35] wl[8] vdd gnd cell_6t
Xbit_r9_c35 bl[35] br[35] wl[9] vdd gnd cell_6t
Xbit_r10_c35 bl[35] br[35] wl[10] vdd gnd cell_6t
Xbit_r11_c35 bl[35] br[35] wl[11] vdd gnd cell_6t
Xbit_r12_c35 bl[35] br[35] wl[12] vdd gnd cell_6t
Xbit_r13_c35 bl[35] br[35] wl[13] vdd gnd cell_6t
Xbit_r14_c35 bl[35] br[35] wl[14] vdd gnd cell_6t
Xbit_r15_c35 bl[35] br[35] wl[15] vdd gnd cell_6t
Xbit_r16_c35 bl[35] br[35] wl[16] vdd gnd cell_6t
Xbit_r17_c35 bl[35] br[35] wl[17] vdd gnd cell_6t
Xbit_r18_c35 bl[35] br[35] wl[18] vdd gnd cell_6t
Xbit_r19_c35 bl[35] br[35] wl[19] vdd gnd cell_6t
Xbit_r20_c35 bl[35] br[35] wl[20] vdd gnd cell_6t
Xbit_r21_c35 bl[35] br[35] wl[21] vdd gnd cell_6t
Xbit_r22_c35 bl[35] br[35] wl[22] vdd gnd cell_6t
Xbit_r23_c35 bl[35] br[35] wl[23] vdd gnd cell_6t
Xbit_r24_c35 bl[35] br[35] wl[24] vdd gnd cell_6t
Xbit_r25_c35 bl[35] br[35] wl[25] vdd gnd cell_6t
Xbit_r26_c35 bl[35] br[35] wl[26] vdd gnd cell_6t
Xbit_r27_c35 bl[35] br[35] wl[27] vdd gnd cell_6t
Xbit_r28_c35 bl[35] br[35] wl[28] vdd gnd cell_6t
Xbit_r29_c35 bl[35] br[35] wl[29] vdd gnd cell_6t
Xbit_r30_c35 bl[35] br[35] wl[30] vdd gnd cell_6t
Xbit_r31_c35 bl[35] br[35] wl[31] vdd gnd cell_6t
Xbit_r32_c35 bl[35] br[35] wl[32] vdd gnd cell_6t
Xbit_r33_c35 bl[35] br[35] wl[33] vdd gnd cell_6t
Xbit_r34_c35 bl[35] br[35] wl[34] vdd gnd cell_6t
Xbit_r35_c35 bl[35] br[35] wl[35] vdd gnd cell_6t
Xbit_r36_c35 bl[35] br[35] wl[36] vdd gnd cell_6t
Xbit_r37_c35 bl[35] br[35] wl[37] vdd gnd cell_6t
Xbit_r38_c35 bl[35] br[35] wl[38] vdd gnd cell_6t
Xbit_r39_c35 bl[35] br[35] wl[39] vdd gnd cell_6t
Xbit_r40_c35 bl[35] br[35] wl[40] vdd gnd cell_6t
Xbit_r41_c35 bl[35] br[35] wl[41] vdd gnd cell_6t
Xbit_r42_c35 bl[35] br[35] wl[42] vdd gnd cell_6t
Xbit_r43_c35 bl[35] br[35] wl[43] vdd gnd cell_6t
Xbit_r44_c35 bl[35] br[35] wl[44] vdd gnd cell_6t
Xbit_r45_c35 bl[35] br[35] wl[45] vdd gnd cell_6t
Xbit_r46_c35 bl[35] br[35] wl[46] vdd gnd cell_6t
Xbit_r47_c35 bl[35] br[35] wl[47] vdd gnd cell_6t
Xbit_r48_c35 bl[35] br[35] wl[48] vdd gnd cell_6t
Xbit_r49_c35 bl[35] br[35] wl[49] vdd gnd cell_6t
Xbit_r50_c35 bl[35] br[35] wl[50] vdd gnd cell_6t
Xbit_r51_c35 bl[35] br[35] wl[51] vdd gnd cell_6t
Xbit_r52_c35 bl[35] br[35] wl[52] vdd gnd cell_6t
Xbit_r53_c35 bl[35] br[35] wl[53] vdd gnd cell_6t
Xbit_r54_c35 bl[35] br[35] wl[54] vdd gnd cell_6t
Xbit_r55_c35 bl[35] br[35] wl[55] vdd gnd cell_6t
Xbit_r56_c35 bl[35] br[35] wl[56] vdd gnd cell_6t
Xbit_r57_c35 bl[35] br[35] wl[57] vdd gnd cell_6t
Xbit_r58_c35 bl[35] br[35] wl[58] vdd gnd cell_6t
Xbit_r59_c35 bl[35] br[35] wl[59] vdd gnd cell_6t
Xbit_r60_c35 bl[35] br[35] wl[60] vdd gnd cell_6t
Xbit_r61_c35 bl[35] br[35] wl[61] vdd gnd cell_6t
Xbit_r62_c35 bl[35] br[35] wl[62] vdd gnd cell_6t
Xbit_r63_c35 bl[35] br[35] wl[63] vdd gnd cell_6t
Xbit_r64_c35 bl[35] br[35] wl[64] vdd gnd cell_6t
Xbit_r65_c35 bl[35] br[35] wl[65] vdd gnd cell_6t
Xbit_r66_c35 bl[35] br[35] wl[66] vdd gnd cell_6t
Xbit_r67_c35 bl[35] br[35] wl[67] vdd gnd cell_6t
Xbit_r68_c35 bl[35] br[35] wl[68] vdd gnd cell_6t
Xbit_r69_c35 bl[35] br[35] wl[69] vdd gnd cell_6t
Xbit_r70_c35 bl[35] br[35] wl[70] vdd gnd cell_6t
Xbit_r71_c35 bl[35] br[35] wl[71] vdd gnd cell_6t
Xbit_r72_c35 bl[35] br[35] wl[72] vdd gnd cell_6t
Xbit_r73_c35 bl[35] br[35] wl[73] vdd gnd cell_6t
Xbit_r74_c35 bl[35] br[35] wl[74] vdd gnd cell_6t
Xbit_r75_c35 bl[35] br[35] wl[75] vdd gnd cell_6t
Xbit_r76_c35 bl[35] br[35] wl[76] vdd gnd cell_6t
Xbit_r77_c35 bl[35] br[35] wl[77] vdd gnd cell_6t
Xbit_r78_c35 bl[35] br[35] wl[78] vdd gnd cell_6t
Xbit_r79_c35 bl[35] br[35] wl[79] vdd gnd cell_6t
Xbit_r80_c35 bl[35] br[35] wl[80] vdd gnd cell_6t
Xbit_r81_c35 bl[35] br[35] wl[81] vdd gnd cell_6t
Xbit_r82_c35 bl[35] br[35] wl[82] vdd gnd cell_6t
Xbit_r83_c35 bl[35] br[35] wl[83] vdd gnd cell_6t
Xbit_r84_c35 bl[35] br[35] wl[84] vdd gnd cell_6t
Xbit_r85_c35 bl[35] br[35] wl[85] vdd gnd cell_6t
Xbit_r86_c35 bl[35] br[35] wl[86] vdd gnd cell_6t
Xbit_r87_c35 bl[35] br[35] wl[87] vdd gnd cell_6t
Xbit_r88_c35 bl[35] br[35] wl[88] vdd gnd cell_6t
Xbit_r89_c35 bl[35] br[35] wl[89] vdd gnd cell_6t
Xbit_r90_c35 bl[35] br[35] wl[90] vdd gnd cell_6t
Xbit_r91_c35 bl[35] br[35] wl[91] vdd gnd cell_6t
Xbit_r92_c35 bl[35] br[35] wl[92] vdd gnd cell_6t
Xbit_r93_c35 bl[35] br[35] wl[93] vdd gnd cell_6t
Xbit_r94_c35 bl[35] br[35] wl[94] vdd gnd cell_6t
Xbit_r95_c35 bl[35] br[35] wl[95] vdd gnd cell_6t
Xbit_r96_c35 bl[35] br[35] wl[96] vdd gnd cell_6t
Xbit_r97_c35 bl[35] br[35] wl[97] vdd gnd cell_6t
Xbit_r98_c35 bl[35] br[35] wl[98] vdd gnd cell_6t
Xbit_r99_c35 bl[35] br[35] wl[99] vdd gnd cell_6t
Xbit_r100_c35 bl[35] br[35] wl[100] vdd gnd cell_6t
Xbit_r101_c35 bl[35] br[35] wl[101] vdd gnd cell_6t
Xbit_r102_c35 bl[35] br[35] wl[102] vdd gnd cell_6t
Xbit_r103_c35 bl[35] br[35] wl[103] vdd gnd cell_6t
Xbit_r104_c35 bl[35] br[35] wl[104] vdd gnd cell_6t
Xbit_r105_c35 bl[35] br[35] wl[105] vdd gnd cell_6t
Xbit_r106_c35 bl[35] br[35] wl[106] vdd gnd cell_6t
Xbit_r107_c35 bl[35] br[35] wl[107] vdd gnd cell_6t
Xbit_r108_c35 bl[35] br[35] wl[108] vdd gnd cell_6t
Xbit_r109_c35 bl[35] br[35] wl[109] vdd gnd cell_6t
Xbit_r110_c35 bl[35] br[35] wl[110] vdd gnd cell_6t
Xbit_r111_c35 bl[35] br[35] wl[111] vdd gnd cell_6t
Xbit_r112_c35 bl[35] br[35] wl[112] vdd gnd cell_6t
Xbit_r113_c35 bl[35] br[35] wl[113] vdd gnd cell_6t
Xbit_r114_c35 bl[35] br[35] wl[114] vdd gnd cell_6t
Xbit_r115_c35 bl[35] br[35] wl[115] vdd gnd cell_6t
Xbit_r116_c35 bl[35] br[35] wl[116] vdd gnd cell_6t
Xbit_r117_c35 bl[35] br[35] wl[117] vdd gnd cell_6t
Xbit_r118_c35 bl[35] br[35] wl[118] vdd gnd cell_6t
Xbit_r119_c35 bl[35] br[35] wl[119] vdd gnd cell_6t
Xbit_r120_c35 bl[35] br[35] wl[120] vdd gnd cell_6t
Xbit_r121_c35 bl[35] br[35] wl[121] vdd gnd cell_6t
Xbit_r122_c35 bl[35] br[35] wl[122] vdd gnd cell_6t
Xbit_r123_c35 bl[35] br[35] wl[123] vdd gnd cell_6t
Xbit_r124_c35 bl[35] br[35] wl[124] vdd gnd cell_6t
Xbit_r125_c35 bl[35] br[35] wl[125] vdd gnd cell_6t
Xbit_r126_c35 bl[35] br[35] wl[126] vdd gnd cell_6t
Xbit_r127_c35 bl[35] br[35] wl[127] vdd gnd cell_6t
Xbit_r128_c35 bl[35] br[35] wl[128] vdd gnd cell_6t
Xbit_r129_c35 bl[35] br[35] wl[129] vdd gnd cell_6t
Xbit_r130_c35 bl[35] br[35] wl[130] vdd gnd cell_6t
Xbit_r131_c35 bl[35] br[35] wl[131] vdd gnd cell_6t
Xbit_r132_c35 bl[35] br[35] wl[132] vdd gnd cell_6t
Xbit_r133_c35 bl[35] br[35] wl[133] vdd gnd cell_6t
Xbit_r134_c35 bl[35] br[35] wl[134] vdd gnd cell_6t
Xbit_r135_c35 bl[35] br[35] wl[135] vdd gnd cell_6t
Xbit_r136_c35 bl[35] br[35] wl[136] vdd gnd cell_6t
Xbit_r137_c35 bl[35] br[35] wl[137] vdd gnd cell_6t
Xbit_r138_c35 bl[35] br[35] wl[138] vdd gnd cell_6t
Xbit_r139_c35 bl[35] br[35] wl[139] vdd gnd cell_6t
Xbit_r140_c35 bl[35] br[35] wl[140] vdd gnd cell_6t
Xbit_r141_c35 bl[35] br[35] wl[141] vdd gnd cell_6t
Xbit_r142_c35 bl[35] br[35] wl[142] vdd gnd cell_6t
Xbit_r143_c35 bl[35] br[35] wl[143] vdd gnd cell_6t
Xbit_r144_c35 bl[35] br[35] wl[144] vdd gnd cell_6t
Xbit_r145_c35 bl[35] br[35] wl[145] vdd gnd cell_6t
Xbit_r146_c35 bl[35] br[35] wl[146] vdd gnd cell_6t
Xbit_r147_c35 bl[35] br[35] wl[147] vdd gnd cell_6t
Xbit_r148_c35 bl[35] br[35] wl[148] vdd gnd cell_6t
Xbit_r149_c35 bl[35] br[35] wl[149] vdd gnd cell_6t
Xbit_r150_c35 bl[35] br[35] wl[150] vdd gnd cell_6t
Xbit_r151_c35 bl[35] br[35] wl[151] vdd gnd cell_6t
Xbit_r152_c35 bl[35] br[35] wl[152] vdd gnd cell_6t
Xbit_r153_c35 bl[35] br[35] wl[153] vdd gnd cell_6t
Xbit_r154_c35 bl[35] br[35] wl[154] vdd gnd cell_6t
Xbit_r155_c35 bl[35] br[35] wl[155] vdd gnd cell_6t
Xbit_r156_c35 bl[35] br[35] wl[156] vdd gnd cell_6t
Xbit_r157_c35 bl[35] br[35] wl[157] vdd gnd cell_6t
Xbit_r158_c35 bl[35] br[35] wl[158] vdd gnd cell_6t
Xbit_r159_c35 bl[35] br[35] wl[159] vdd gnd cell_6t
Xbit_r160_c35 bl[35] br[35] wl[160] vdd gnd cell_6t
Xbit_r161_c35 bl[35] br[35] wl[161] vdd gnd cell_6t
Xbit_r162_c35 bl[35] br[35] wl[162] vdd gnd cell_6t
Xbit_r163_c35 bl[35] br[35] wl[163] vdd gnd cell_6t
Xbit_r164_c35 bl[35] br[35] wl[164] vdd gnd cell_6t
Xbit_r165_c35 bl[35] br[35] wl[165] vdd gnd cell_6t
Xbit_r166_c35 bl[35] br[35] wl[166] vdd gnd cell_6t
Xbit_r167_c35 bl[35] br[35] wl[167] vdd gnd cell_6t
Xbit_r168_c35 bl[35] br[35] wl[168] vdd gnd cell_6t
Xbit_r169_c35 bl[35] br[35] wl[169] vdd gnd cell_6t
Xbit_r170_c35 bl[35] br[35] wl[170] vdd gnd cell_6t
Xbit_r171_c35 bl[35] br[35] wl[171] vdd gnd cell_6t
Xbit_r172_c35 bl[35] br[35] wl[172] vdd gnd cell_6t
Xbit_r173_c35 bl[35] br[35] wl[173] vdd gnd cell_6t
Xbit_r174_c35 bl[35] br[35] wl[174] vdd gnd cell_6t
Xbit_r175_c35 bl[35] br[35] wl[175] vdd gnd cell_6t
Xbit_r176_c35 bl[35] br[35] wl[176] vdd gnd cell_6t
Xbit_r177_c35 bl[35] br[35] wl[177] vdd gnd cell_6t
Xbit_r178_c35 bl[35] br[35] wl[178] vdd gnd cell_6t
Xbit_r179_c35 bl[35] br[35] wl[179] vdd gnd cell_6t
Xbit_r180_c35 bl[35] br[35] wl[180] vdd gnd cell_6t
Xbit_r181_c35 bl[35] br[35] wl[181] vdd gnd cell_6t
Xbit_r182_c35 bl[35] br[35] wl[182] vdd gnd cell_6t
Xbit_r183_c35 bl[35] br[35] wl[183] vdd gnd cell_6t
Xbit_r184_c35 bl[35] br[35] wl[184] vdd gnd cell_6t
Xbit_r185_c35 bl[35] br[35] wl[185] vdd gnd cell_6t
Xbit_r186_c35 bl[35] br[35] wl[186] vdd gnd cell_6t
Xbit_r187_c35 bl[35] br[35] wl[187] vdd gnd cell_6t
Xbit_r188_c35 bl[35] br[35] wl[188] vdd gnd cell_6t
Xbit_r189_c35 bl[35] br[35] wl[189] vdd gnd cell_6t
Xbit_r190_c35 bl[35] br[35] wl[190] vdd gnd cell_6t
Xbit_r191_c35 bl[35] br[35] wl[191] vdd gnd cell_6t
Xbit_r192_c35 bl[35] br[35] wl[192] vdd gnd cell_6t
Xbit_r193_c35 bl[35] br[35] wl[193] vdd gnd cell_6t
Xbit_r194_c35 bl[35] br[35] wl[194] vdd gnd cell_6t
Xbit_r195_c35 bl[35] br[35] wl[195] vdd gnd cell_6t
Xbit_r196_c35 bl[35] br[35] wl[196] vdd gnd cell_6t
Xbit_r197_c35 bl[35] br[35] wl[197] vdd gnd cell_6t
Xbit_r198_c35 bl[35] br[35] wl[198] vdd gnd cell_6t
Xbit_r199_c35 bl[35] br[35] wl[199] vdd gnd cell_6t
Xbit_r200_c35 bl[35] br[35] wl[200] vdd gnd cell_6t
Xbit_r201_c35 bl[35] br[35] wl[201] vdd gnd cell_6t
Xbit_r202_c35 bl[35] br[35] wl[202] vdd gnd cell_6t
Xbit_r203_c35 bl[35] br[35] wl[203] vdd gnd cell_6t
Xbit_r204_c35 bl[35] br[35] wl[204] vdd gnd cell_6t
Xbit_r205_c35 bl[35] br[35] wl[205] vdd gnd cell_6t
Xbit_r206_c35 bl[35] br[35] wl[206] vdd gnd cell_6t
Xbit_r207_c35 bl[35] br[35] wl[207] vdd gnd cell_6t
Xbit_r208_c35 bl[35] br[35] wl[208] vdd gnd cell_6t
Xbit_r209_c35 bl[35] br[35] wl[209] vdd gnd cell_6t
Xbit_r210_c35 bl[35] br[35] wl[210] vdd gnd cell_6t
Xbit_r211_c35 bl[35] br[35] wl[211] vdd gnd cell_6t
Xbit_r212_c35 bl[35] br[35] wl[212] vdd gnd cell_6t
Xbit_r213_c35 bl[35] br[35] wl[213] vdd gnd cell_6t
Xbit_r214_c35 bl[35] br[35] wl[214] vdd gnd cell_6t
Xbit_r215_c35 bl[35] br[35] wl[215] vdd gnd cell_6t
Xbit_r216_c35 bl[35] br[35] wl[216] vdd gnd cell_6t
Xbit_r217_c35 bl[35] br[35] wl[217] vdd gnd cell_6t
Xbit_r218_c35 bl[35] br[35] wl[218] vdd gnd cell_6t
Xbit_r219_c35 bl[35] br[35] wl[219] vdd gnd cell_6t
Xbit_r220_c35 bl[35] br[35] wl[220] vdd gnd cell_6t
Xbit_r221_c35 bl[35] br[35] wl[221] vdd gnd cell_6t
Xbit_r222_c35 bl[35] br[35] wl[222] vdd gnd cell_6t
Xbit_r223_c35 bl[35] br[35] wl[223] vdd gnd cell_6t
Xbit_r224_c35 bl[35] br[35] wl[224] vdd gnd cell_6t
Xbit_r225_c35 bl[35] br[35] wl[225] vdd gnd cell_6t
Xbit_r226_c35 bl[35] br[35] wl[226] vdd gnd cell_6t
Xbit_r227_c35 bl[35] br[35] wl[227] vdd gnd cell_6t
Xbit_r228_c35 bl[35] br[35] wl[228] vdd gnd cell_6t
Xbit_r229_c35 bl[35] br[35] wl[229] vdd gnd cell_6t
Xbit_r230_c35 bl[35] br[35] wl[230] vdd gnd cell_6t
Xbit_r231_c35 bl[35] br[35] wl[231] vdd gnd cell_6t
Xbit_r232_c35 bl[35] br[35] wl[232] vdd gnd cell_6t
Xbit_r233_c35 bl[35] br[35] wl[233] vdd gnd cell_6t
Xbit_r234_c35 bl[35] br[35] wl[234] vdd gnd cell_6t
Xbit_r235_c35 bl[35] br[35] wl[235] vdd gnd cell_6t
Xbit_r236_c35 bl[35] br[35] wl[236] vdd gnd cell_6t
Xbit_r237_c35 bl[35] br[35] wl[237] vdd gnd cell_6t
Xbit_r238_c35 bl[35] br[35] wl[238] vdd gnd cell_6t
Xbit_r239_c35 bl[35] br[35] wl[239] vdd gnd cell_6t
Xbit_r240_c35 bl[35] br[35] wl[240] vdd gnd cell_6t
Xbit_r241_c35 bl[35] br[35] wl[241] vdd gnd cell_6t
Xbit_r242_c35 bl[35] br[35] wl[242] vdd gnd cell_6t
Xbit_r243_c35 bl[35] br[35] wl[243] vdd gnd cell_6t
Xbit_r244_c35 bl[35] br[35] wl[244] vdd gnd cell_6t
Xbit_r245_c35 bl[35] br[35] wl[245] vdd gnd cell_6t
Xbit_r246_c35 bl[35] br[35] wl[246] vdd gnd cell_6t
Xbit_r247_c35 bl[35] br[35] wl[247] vdd gnd cell_6t
Xbit_r248_c35 bl[35] br[35] wl[248] vdd gnd cell_6t
Xbit_r249_c35 bl[35] br[35] wl[249] vdd gnd cell_6t
Xbit_r250_c35 bl[35] br[35] wl[250] vdd gnd cell_6t
Xbit_r251_c35 bl[35] br[35] wl[251] vdd gnd cell_6t
Xbit_r252_c35 bl[35] br[35] wl[252] vdd gnd cell_6t
Xbit_r253_c35 bl[35] br[35] wl[253] vdd gnd cell_6t
Xbit_r254_c35 bl[35] br[35] wl[254] vdd gnd cell_6t
Xbit_r255_c35 bl[35] br[35] wl[255] vdd gnd cell_6t
Xbit_r256_c35 bl[35] br[35] wl[256] vdd gnd cell_6t
Xbit_r257_c35 bl[35] br[35] wl[257] vdd gnd cell_6t
Xbit_r258_c35 bl[35] br[35] wl[258] vdd gnd cell_6t
Xbit_r259_c35 bl[35] br[35] wl[259] vdd gnd cell_6t
Xbit_r260_c35 bl[35] br[35] wl[260] vdd gnd cell_6t
Xbit_r261_c35 bl[35] br[35] wl[261] vdd gnd cell_6t
Xbit_r262_c35 bl[35] br[35] wl[262] vdd gnd cell_6t
Xbit_r263_c35 bl[35] br[35] wl[263] vdd gnd cell_6t
Xbit_r264_c35 bl[35] br[35] wl[264] vdd gnd cell_6t
Xbit_r265_c35 bl[35] br[35] wl[265] vdd gnd cell_6t
Xbit_r266_c35 bl[35] br[35] wl[266] vdd gnd cell_6t
Xbit_r267_c35 bl[35] br[35] wl[267] vdd gnd cell_6t
Xbit_r268_c35 bl[35] br[35] wl[268] vdd gnd cell_6t
Xbit_r269_c35 bl[35] br[35] wl[269] vdd gnd cell_6t
Xbit_r270_c35 bl[35] br[35] wl[270] vdd gnd cell_6t
Xbit_r271_c35 bl[35] br[35] wl[271] vdd gnd cell_6t
Xbit_r272_c35 bl[35] br[35] wl[272] vdd gnd cell_6t
Xbit_r273_c35 bl[35] br[35] wl[273] vdd gnd cell_6t
Xbit_r274_c35 bl[35] br[35] wl[274] vdd gnd cell_6t
Xbit_r275_c35 bl[35] br[35] wl[275] vdd gnd cell_6t
Xbit_r276_c35 bl[35] br[35] wl[276] vdd gnd cell_6t
Xbit_r277_c35 bl[35] br[35] wl[277] vdd gnd cell_6t
Xbit_r278_c35 bl[35] br[35] wl[278] vdd gnd cell_6t
Xbit_r279_c35 bl[35] br[35] wl[279] vdd gnd cell_6t
Xbit_r280_c35 bl[35] br[35] wl[280] vdd gnd cell_6t
Xbit_r281_c35 bl[35] br[35] wl[281] vdd gnd cell_6t
Xbit_r282_c35 bl[35] br[35] wl[282] vdd gnd cell_6t
Xbit_r283_c35 bl[35] br[35] wl[283] vdd gnd cell_6t
Xbit_r284_c35 bl[35] br[35] wl[284] vdd gnd cell_6t
Xbit_r285_c35 bl[35] br[35] wl[285] vdd gnd cell_6t
Xbit_r286_c35 bl[35] br[35] wl[286] vdd gnd cell_6t
Xbit_r287_c35 bl[35] br[35] wl[287] vdd gnd cell_6t
Xbit_r288_c35 bl[35] br[35] wl[288] vdd gnd cell_6t
Xbit_r289_c35 bl[35] br[35] wl[289] vdd gnd cell_6t
Xbit_r290_c35 bl[35] br[35] wl[290] vdd gnd cell_6t
Xbit_r291_c35 bl[35] br[35] wl[291] vdd gnd cell_6t
Xbit_r292_c35 bl[35] br[35] wl[292] vdd gnd cell_6t
Xbit_r293_c35 bl[35] br[35] wl[293] vdd gnd cell_6t
Xbit_r294_c35 bl[35] br[35] wl[294] vdd gnd cell_6t
Xbit_r295_c35 bl[35] br[35] wl[295] vdd gnd cell_6t
Xbit_r296_c35 bl[35] br[35] wl[296] vdd gnd cell_6t
Xbit_r297_c35 bl[35] br[35] wl[297] vdd gnd cell_6t
Xbit_r298_c35 bl[35] br[35] wl[298] vdd gnd cell_6t
Xbit_r299_c35 bl[35] br[35] wl[299] vdd gnd cell_6t
Xbit_r300_c35 bl[35] br[35] wl[300] vdd gnd cell_6t
Xbit_r301_c35 bl[35] br[35] wl[301] vdd gnd cell_6t
Xbit_r302_c35 bl[35] br[35] wl[302] vdd gnd cell_6t
Xbit_r303_c35 bl[35] br[35] wl[303] vdd gnd cell_6t
Xbit_r304_c35 bl[35] br[35] wl[304] vdd gnd cell_6t
Xbit_r305_c35 bl[35] br[35] wl[305] vdd gnd cell_6t
Xbit_r306_c35 bl[35] br[35] wl[306] vdd gnd cell_6t
Xbit_r307_c35 bl[35] br[35] wl[307] vdd gnd cell_6t
Xbit_r308_c35 bl[35] br[35] wl[308] vdd gnd cell_6t
Xbit_r309_c35 bl[35] br[35] wl[309] vdd gnd cell_6t
Xbit_r310_c35 bl[35] br[35] wl[310] vdd gnd cell_6t
Xbit_r311_c35 bl[35] br[35] wl[311] vdd gnd cell_6t
Xbit_r312_c35 bl[35] br[35] wl[312] vdd gnd cell_6t
Xbit_r313_c35 bl[35] br[35] wl[313] vdd gnd cell_6t
Xbit_r314_c35 bl[35] br[35] wl[314] vdd gnd cell_6t
Xbit_r315_c35 bl[35] br[35] wl[315] vdd gnd cell_6t
Xbit_r316_c35 bl[35] br[35] wl[316] vdd gnd cell_6t
Xbit_r317_c35 bl[35] br[35] wl[317] vdd gnd cell_6t
Xbit_r318_c35 bl[35] br[35] wl[318] vdd gnd cell_6t
Xbit_r319_c35 bl[35] br[35] wl[319] vdd gnd cell_6t
Xbit_r320_c35 bl[35] br[35] wl[320] vdd gnd cell_6t
Xbit_r321_c35 bl[35] br[35] wl[321] vdd gnd cell_6t
Xbit_r322_c35 bl[35] br[35] wl[322] vdd gnd cell_6t
Xbit_r323_c35 bl[35] br[35] wl[323] vdd gnd cell_6t
Xbit_r324_c35 bl[35] br[35] wl[324] vdd gnd cell_6t
Xbit_r325_c35 bl[35] br[35] wl[325] vdd gnd cell_6t
Xbit_r326_c35 bl[35] br[35] wl[326] vdd gnd cell_6t
Xbit_r327_c35 bl[35] br[35] wl[327] vdd gnd cell_6t
Xbit_r328_c35 bl[35] br[35] wl[328] vdd gnd cell_6t
Xbit_r329_c35 bl[35] br[35] wl[329] vdd gnd cell_6t
Xbit_r330_c35 bl[35] br[35] wl[330] vdd gnd cell_6t
Xbit_r331_c35 bl[35] br[35] wl[331] vdd gnd cell_6t
Xbit_r332_c35 bl[35] br[35] wl[332] vdd gnd cell_6t
Xbit_r333_c35 bl[35] br[35] wl[333] vdd gnd cell_6t
Xbit_r334_c35 bl[35] br[35] wl[334] vdd gnd cell_6t
Xbit_r335_c35 bl[35] br[35] wl[335] vdd gnd cell_6t
Xbit_r336_c35 bl[35] br[35] wl[336] vdd gnd cell_6t
Xbit_r337_c35 bl[35] br[35] wl[337] vdd gnd cell_6t
Xbit_r338_c35 bl[35] br[35] wl[338] vdd gnd cell_6t
Xbit_r339_c35 bl[35] br[35] wl[339] vdd gnd cell_6t
Xbit_r340_c35 bl[35] br[35] wl[340] vdd gnd cell_6t
Xbit_r341_c35 bl[35] br[35] wl[341] vdd gnd cell_6t
Xbit_r342_c35 bl[35] br[35] wl[342] vdd gnd cell_6t
Xbit_r343_c35 bl[35] br[35] wl[343] vdd gnd cell_6t
Xbit_r344_c35 bl[35] br[35] wl[344] vdd gnd cell_6t
Xbit_r345_c35 bl[35] br[35] wl[345] vdd gnd cell_6t
Xbit_r346_c35 bl[35] br[35] wl[346] vdd gnd cell_6t
Xbit_r347_c35 bl[35] br[35] wl[347] vdd gnd cell_6t
Xbit_r348_c35 bl[35] br[35] wl[348] vdd gnd cell_6t
Xbit_r349_c35 bl[35] br[35] wl[349] vdd gnd cell_6t
Xbit_r350_c35 bl[35] br[35] wl[350] vdd gnd cell_6t
Xbit_r351_c35 bl[35] br[35] wl[351] vdd gnd cell_6t
Xbit_r352_c35 bl[35] br[35] wl[352] vdd gnd cell_6t
Xbit_r353_c35 bl[35] br[35] wl[353] vdd gnd cell_6t
Xbit_r354_c35 bl[35] br[35] wl[354] vdd gnd cell_6t
Xbit_r355_c35 bl[35] br[35] wl[355] vdd gnd cell_6t
Xbit_r356_c35 bl[35] br[35] wl[356] vdd gnd cell_6t
Xbit_r357_c35 bl[35] br[35] wl[357] vdd gnd cell_6t
Xbit_r358_c35 bl[35] br[35] wl[358] vdd gnd cell_6t
Xbit_r359_c35 bl[35] br[35] wl[359] vdd gnd cell_6t
Xbit_r360_c35 bl[35] br[35] wl[360] vdd gnd cell_6t
Xbit_r361_c35 bl[35] br[35] wl[361] vdd gnd cell_6t
Xbit_r362_c35 bl[35] br[35] wl[362] vdd gnd cell_6t
Xbit_r363_c35 bl[35] br[35] wl[363] vdd gnd cell_6t
Xbit_r364_c35 bl[35] br[35] wl[364] vdd gnd cell_6t
Xbit_r365_c35 bl[35] br[35] wl[365] vdd gnd cell_6t
Xbit_r366_c35 bl[35] br[35] wl[366] vdd gnd cell_6t
Xbit_r367_c35 bl[35] br[35] wl[367] vdd gnd cell_6t
Xbit_r368_c35 bl[35] br[35] wl[368] vdd gnd cell_6t
Xbit_r369_c35 bl[35] br[35] wl[369] vdd gnd cell_6t
Xbit_r370_c35 bl[35] br[35] wl[370] vdd gnd cell_6t
Xbit_r371_c35 bl[35] br[35] wl[371] vdd gnd cell_6t
Xbit_r372_c35 bl[35] br[35] wl[372] vdd gnd cell_6t
Xbit_r373_c35 bl[35] br[35] wl[373] vdd gnd cell_6t
Xbit_r374_c35 bl[35] br[35] wl[374] vdd gnd cell_6t
Xbit_r375_c35 bl[35] br[35] wl[375] vdd gnd cell_6t
Xbit_r376_c35 bl[35] br[35] wl[376] vdd gnd cell_6t
Xbit_r377_c35 bl[35] br[35] wl[377] vdd gnd cell_6t
Xbit_r378_c35 bl[35] br[35] wl[378] vdd gnd cell_6t
Xbit_r379_c35 bl[35] br[35] wl[379] vdd gnd cell_6t
Xbit_r380_c35 bl[35] br[35] wl[380] vdd gnd cell_6t
Xbit_r381_c35 bl[35] br[35] wl[381] vdd gnd cell_6t
Xbit_r382_c35 bl[35] br[35] wl[382] vdd gnd cell_6t
Xbit_r383_c35 bl[35] br[35] wl[383] vdd gnd cell_6t
Xbit_r384_c35 bl[35] br[35] wl[384] vdd gnd cell_6t
Xbit_r385_c35 bl[35] br[35] wl[385] vdd gnd cell_6t
Xbit_r386_c35 bl[35] br[35] wl[386] vdd gnd cell_6t
Xbit_r387_c35 bl[35] br[35] wl[387] vdd gnd cell_6t
Xbit_r388_c35 bl[35] br[35] wl[388] vdd gnd cell_6t
Xbit_r389_c35 bl[35] br[35] wl[389] vdd gnd cell_6t
Xbit_r390_c35 bl[35] br[35] wl[390] vdd gnd cell_6t
Xbit_r391_c35 bl[35] br[35] wl[391] vdd gnd cell_6t
Xbit_r392_c35 bl[35] br[35] wl[392] vdd gnd cell_6t
Xbit_r393_c35 bl[35] br[35] wl[393] vdd gnd cell_6t
Xbit_r394_c35 bl[35] br[35] wl[394] vdd gnd cell_6t
Xbit_r395_c35 bl[35] br[35] wl[395] vdd gnd cell_6t
Xbit_r396_c35 bl[35] br[35] wl[396] vdd gnd cell_6t
Xbit_r397_c35 bl[35] br[35] wl[397] vdd gnd cell_6t
Xbit_r398_c35 bl[35] br[35] wl[398] vdd gnd cell_6t
Xbit_r399_c35 bl[35] br[35] wl[399] vdd gnd cell_6t
Xbit_r400_c35 bl[35] br[35] wl[400] vdd gnd cell_6t
Xbit_r401_c35 bl[35] br[35] wl[401] vdd gnd cell_6t
Xbit_r402_c35 bl[35] br[35] wl[402] vdd gnd cell_6t
Xbit_r403_c35 bl[35] br[35] wl[403] vdd gnd cell_6t
Xbit_r404_c35 bl[35] br[35] wl[404] vdd gnd cell_6t
Xbit_r405_c35 bl[35] br[35] wl[405] vdd gnd cell_6t
Xbit_r406_c35 bl[35] br[35] wl[406] vdd gnd cell_6t
Xbit_r407_c35 bl[35] br[35] wl[407] vdd gnd cell_6t
Xbit_r408_c35 bl[35] br[35] wl[408] vdd gnd cell_6t
Xbit_r409_c35 bl[35] br[35] wl[409] vdd gnd cell_6t
Xbit_r410_c35 bl[35] br[35] wl[410] vdd gnd cell_6t
Xbit_r411_c35 bl[35] br[35] wl[411] vdd gnd cell_6t
Xbit_r412_c35 bl[35] br[35] wl[412] vdd gnd cell_6t
Xbit_r413_c35 bl[35] br[35] wl[413] vdd gnd cell_6t
Xbit_r414_c35 bl[35] br[35] wl[414] vdd gnd cell_6t
Xbit_r415_c35 bl[35] br[35] wl[415] vdd gnd cell_6t
Xbit_r416_c35 bl[35] br[35] wl[416] vdd gnd cell_6t
Xbit_r417_c35 bl[35] br[35] wl[417] vdd gnd cell_6t
Xbit_r418_c35 bl[35] br[35] wl[418] vdd gnd cell_6t
Xbit_r419_c35 bl[35] br[35] wl[419] vdd gnd cell_6t
Xbit_r420_c35 bl[35] br[35] wl[420] vdd gnd cell_6t
Xbit_r421_c35 bl[35] br[35] wl[421] vdd gnd cell_6t
Xbit_r422_c35 bl[35] br[35] wl[422] vdd gnd cell_6t
Xbit_r423_c35 bl[35] br[35] wl[423] vdd gnd cell_6t
Xbit_r424_c35 bl[35] br[35] wl[424] vdd gnd cell_6t
Xbit_r425_c35 bl[35] br[35] wl[425] vdd gnd cell_6t
Xbit_r426_c35 bl[35] br[35] wl[426] vdd gnd cell_6t
Xbit_r427_c35 bl[35] br[35] wl[427] vdd gnd cell_6t
Xbit_r428_c35 bl[35] br[35] wl[428] vdd gnd cell_6t
Xbit_r429_c35 bl[35] br[35] wl[429] vdd gnd cell_6t
Xbit_r430_c35 bl[35] br[35] wl[430] vdd gnd cell_6t
Xbit_r431_c35 bl[35] br[35] wl[431] vdd gnd cell_6t
Xbit_r432_c35 bl[35] br[35] wl[432] vdd gnd cell_6t
Xbit_r433_c35 bl[35] br[35] wl[433] vdd gnd cell_6t
Xbit_r434_c35 bl[35] br[35] wl[434] vdd gnd cell_6t
Xbit_r435_c35 bl[35] br[35] wl[435] vdd gnd cell_6t
Xbit_r436_c35 bl[35] br[35] wl[436] vdd gnd cell_6t
Xbit_r437_c35 bl[35] br[35] wl[437] vdd gnd cell_6t
Xbit_r438_c35 bl[35] br[35] wl[438] vdd gnd cell_6t
Xbit_r439_c35 bl[35] br[35] wl[439] vdd gnd cell_6t
Xbit_r440_c35 bl[35] br[35] wl[440] vdd gnd cell_6t
Xbit_r441_c35 bl[35] br[35] wl[441] vdd gnd cell_6t
Xbit_r442_c35 bl[35] br[35] wl[442] vdd gnd cell_6t
Xbit_r443_c35 bl[35] br[35] wl[443] vdd gnd cell_6t
Xbit_r444_c35 bl[35] br[35] wl[444] vdd gnd cell_6t
Xbit_r445_c35 bl[35] br[35] wl[445] vdd gnd cell_6t
Xbit_r446_c35 bl[35] br[35] wl[446] vdd gnd cell_6t
Xbit_r447_c35 bl[35] br[35] wl[447] vdd gnd cell_6t
Xbit_r448_c35 bl[35] br[35] wl[448] vdd gnd cell_6t
Xbit_r449_c35 bl[35] br[35] wl[449] vdd gnd cell_6t
Xbit_r450_c35 bl[35] br[35] wl[450] vdd gnd cell_6t
Xbit_r451_c35 bl[35] br[35] wl[451] vdd gnd cell_6t
Xbit_r452_c35 bl[35] br[35] wl[452] vdd gnd cell_6t
Xbit_r453_c35 bl[35] br[35] wl[453] vdd gnd cell_6t
Xbit_r454_c35 bl[35] br[35] wl[454] vdd gnd cell_6t
Xbit_r455_c35 bl[35] br[35] wl[455] vdd gnd cell_6t
Xbit_r456_c35 bl[35] br[35] wl[456] vdd gnd cell_6t
Xbit_r457_c35 bl[35] br[35] wl[457] vdd gnd cell_6t
Xbit_r458_c35 bl[35] br[35] wl[458] vdd gnd cell_6t
Xbit_r459_c35 bl[35] br[35] wl[459] vdd gnd cell_6t
Xbit_r460_c35 bl[35] br[35] wl[460] vdd gnd cell_6t
Xbit_r461_c35 bl[35] br[35] wl[461] vdd gnd cell_6t
Xbit_r462_c35 bl[35] br[35] wl[462] vdd gnd cell_6t
Xbit_r463_c35 bl[35] br[35] wl[463] vdd gnd cell_6t
Xbit_r464_c35 bl[35] br[35] wl[464] vdd gnd cell_6t
Xbit_r465_c35 bl[35] br[35] wl[465] vdd gnd cell_6t
Xbit_r466_c35 bl[35] br[35] wl[466] vdd gnd cell_6t
Xbit_r467_c35 bl[35] br[35] wl[467] vdd gnd cell_6t
Xbit_r468_c35 bl[35] br[35] wl[468] vdd gnd cell_6t
Xbit_r469_c35 bl[35] br[35] wl[469] vdd gnd cell_6t
Xbit_r470_c35 bl[35] br[35] wl[470] vdd gnd cell_6t
Xbit_r471_c35 bl[35] br[35] wl[471] vdd gnd cell_6t
Xbit_r472_c35 bl[35] br[35] wl[472] vdd gnd cell_6t
Xbit_r473_c35 bl[35] br[35] wl[473] vdd gnd cell_6t
Xbit_r474_c35 bl[35] br[35] wl[474] vdd gnd cell_6t
Xbit_r475_c35 bl[35] br[35] wl[475] vdd gnd cell_6t
Xbit_r476_c35 bl[35] br[35] wl[476] vdd gnd cell_6t
Xbit_r477_c35 bl[35] br[35] wl[477] vdd gnd cell_6t
Xbit_r478_c35 bl[35] br[35] wl[478] vdd gnd cell_6t
Xbit_r479_c35 bl[35] br[35] wl[479] vdd gnd cell_6t
Xbit_r480_c35 bl[35] br[35] wl[480] vdd gnd cell_6t
Xbit_r481_c35 bl[35] br[35] wl[481] vdd gnd cell_6t
Xbit_r482_c35 bl[35] br[35] wl[482] vdd gnd cell_6t
Xbit_r483_c35 bl[35] br[35] wl[483] vdd gnd cell_6t
Xbit_r484_c35 bl[35] br[35] wl[484] vdd gnd cell_6t
Xbit_r485_c35 bl[35] br[35] wl[485] vdd gnd cell_6t
Xbit_r486_c35 bl[35] br[35] wl[486] vdd gnd cell_6t
Xbit_r487_c35 bl[35] br[35] wl[487] vdd gnd cell_6t
Xbit_r488_c35 bl[35] br[35] wl[488] vdd gnd cell_6t
Xbit_r489_c35 bl[35] br[35] wl[489] vdd gnd cell_6t
Xbit_r490_c35 bl[35] br[35] wl[490] vdd gnd cell_6t
Xbit_r491_c35 bl[35] br[35] wl[491] vdd gnd cell_6t
Xbit_r492_c35 bl[35] br[35] wl[492] vdd gnd cell_6t
Xbit_r493_c35 bl[35] br[35] wl[493] vdd gnd cell_6t
Xbit_r494_c35 bl[35] br[35] wl[494] vdd gnd cell_6t
Xbit_r495_c35 bl[35] br[35] wl[495] vdd gnd cell_6t
Xbit_r496_c35 bl[35] br[35] wl[496] vdd gnd cell_6t
Xbit_r497_c35 bl[35] br[35] wl[497] vdd gnd cell_6t
Xbit_r498_c35 bl[35] br[35] wl[498] vdd gnd cell_6t
Xbit_r499_c35 bl[35] br[35] wl[499] vdd gnd cell_6t
Xbit_r500_c35 bl[35] br[35] wl[500] vdd gnd cell_6t
Xbit_r501_c35 bl[35] br[35] wl[501] vdd gnd cell_6t
Xbit_r502_c35 bl[35] br[35] wl[502] vdd gnd cell_6t
Xbit_r503_c35 bl[35] br[35] wl[503] vdd gnd cell_6t
Xbit_r504_c35 bl[35] br[35] wl[504] vdd gnd cell_6t
Xbit_r505_c35 bl[35] br[35] wl[505] vdd gnd cell_6t
Xbit_r506_c35 bl[35] br[35] wl[506] vdd gnd cell_6t
Xbit_r507_c35 bl[35] br[35] wl[507] vdd gnd cell_6t
Xbit_r508_c35 bl[35] br[35] wl[508] vdd gnd cell_6t
Xbit_r509_c35 bl[35] br[35] wl[509] vdd gnd cell_6t
Xbit_r510_c35 bl[35] br[35] wl[510] vdd gnd cell_6t
Xbit_r511_c35 bl[35] br[35] wl[511] vdd gnd cell_6t
Xbit_r0_c36 bl[36] br[36] wl[0] vdd gnd cell_6t
Xbit_r1_c36 bl[36] br[36] wl[1] vdd gnd cell_6t
Xbit_r2_c36 bl[36] br[36] wl[2] vdd gnd cell_6t
Xbit_r3_c36 bl[36] br[36] wl[3] vdd gnd cell_6t
Xbit_r4_c36 bl[36] br[36] wl[4] vdd gnd cell_6t
Xbit_r5_c36 bl[36] br[36] wl[5] vdd gnd cell_6t
Xbit_r6_c36 bl[36] br[36] wl[6] vdd gnd cell_6t
Xbit_r7_c36 bl[36] br[36] wl[7] vdd gnd cell_6t
Xbit_r8_c36 bl[36] br[36] wl[8] vdd gnd cell_6t
Xbit_r9_c36 bl[36] br[36] wl[9] vdd gnd cell_6t
Xbit_r10_c36 bl[36] br[36] wl[10] vdd gnd cell_6t
Xbit_r11_c36 bl[36] br[36] wl[11] vdd gnd cell_6t
Xbit_r12_c36 bl[36] br[36] wl[12] vdd gnd cell_6t
Xbit_r13_c36 bl[36] br[36] wl[13] vdd gnd cell_6t
Xbit_r14_c36 bl[36] br[36] wl[14] vdd gnd cell_6t
Xbit_r15_c36 bl[36] br[36] wl[15] vdd gnd cell_6t
Xbit_r16_c36 bl[36] br[36] wl[16] vdd gnd cell_6t
Xbit_r17_c36 bl[36] br[36] wl[17] vdd gnd cell_6t
Xbit_r18_c36 bl[36] br[36] wl[18] vdd gnd cell_6t
Xbit_r19_c36 bl[36] br[36] wl[19] vdd gnd cell_6t
Xbit_r20_c36 bl[36] br[36] wl[20] vdd gnd cell_6t
Xbit_r21_c36 bl[36] br[36] wl[21] vdd gnd cell_6t
Xbit_r22_c36 bl[36] br[36] wl[22] vdd gnd cell_6t
Xbit_r23_c36 bl[36] br[36] wl[23] vdd gnd cell_6t
Xbit_r24_c36 bl[36] br[36] wl[24] vdd gnd cell_6t
Xbit_r25_c36 bl[36] br[36] wl[25] vdd gnd cell_6t
Xbit_r26_c36 bl[36] br[36] wl[26] vdd gnd cell_6t
Xbit_r27_c36 bl[36] br[36] wl[27] vdd gnd cell_6t
Xbit_r28_c36 bl[36] br[36] wl[28] vdd gnd cell_6t
Xbit_r29_c36 bl[36] br[36] wl[29] vdd gnd cell_6t
Xbit_r30_c36 bl[36] br[36] wl[30] vdd gnd cell_6t
Xbit_r31_c36 bl[36] br[36] wl[31] vdd gnd cell_6t
Xbit_r32_c36 bl[36] br[36] wl[32] vdd gnd cell_6t
Xbit_r33_c36 bl[36] br[36] wl[33] vdd gnd cell_6t
Xbit_r34_c36 bl[36] br[36] wl[34] vdd gnd cell_6t
Xbit_r35_c36 bl[36] br[36] wl[35] vdd gnd cell_6t
Xbit_r36_c36 bl[36] br[36] wl[36] vdd gnd cell_6t
Xbit_r37_c36 bl[36] br[36] wl[37] vdd gnd cell_6t
Xbit_r38_c36 bl[36] br[36] wl[38] vdd gnd cell_6t
Xbit_r39_c36 bl[36] br[36] wl[39] vdd gnd cell_6t
Xbit_r40_c36 bl[36] br[36] wl[40] vdd gnd cell_6t
Xbit_r41_c36 bl[36] br[36] wl[41] vdd gnd cell_6t
Xbit_r42_c36 bl[36] br[36] wl[42] vdd gnd cell_6t
Xbit_r43_c36 bl[36] br[36] wl[43] vdd gnd cell_6t
Xbit_r44_c36 bl[36] br[36] wl[44] vdd gnd cell_6t
Xbit_r45_c36 bl[36] br[36] wl[45] vdd gnd cell_6t
Xbit_r46_c36 bl[36] br[36] wl[46] vdd gnd cell_6t
Xbit_r47_c36 bl[36] br[36] wl[47] vdd gnd cell_6t
Xbit_r48_c36 bl[36] br[36] wl[48] vdd gnd cell_6t
Xbit_r49_c36 bl[36] br[36] wl[49] vdd gnd cell_6t
Xbit_r50_c36 bl[36] br[36] wl[50] vdd gnd cell_6t
Xbit_r51_c36 bl[36] br[36] wl[51] vdd gnd cell_6t
Xbit_r52_c36 bl[36] br[36] wl[52] vdd gnd cell_6t
Xbit_r53_c36 bl[36] br[36] wl[53] vdd gnd cell_6t
Xbit_r54_c36 bl[36] br[36] wl[54] vdd gnd cell_6t
Xbit_r55_c36 bl[36] br[36] wl[55] vdd gnd cell_6t
Xbit_r56_c36 bl[36] br[36] wl[56] vdd gnd cell_6t
Xbit_r57_c36 bl[36] br[36] wl[57] vdd gnd cell_6t
Xbit_r58_c36 bl[36] br[36] wl[58] vdd gnd cell_6t
Xbit_r59_c36 bl[36] br[36] wl[59] vdd gnd cell_6t
Xbit_r60_c36 bl[36] br[36] wl[60] vdd gnd cell_6t
Xbit_r61_c36 bl[36] br[36] wl[61] vdd gnd cell_6t
Xbit_r62_c36 bl[36] br[36] wl[62] vdd gnd cell_6t
Xbit_r63_c36 bl[36] br[36] wl[63] vdd gnd cell_6t
Xbit_r64_c36 bl[36] br[36] wl[64] vdd gnd cell_6t
Xbit_r65_c36 bl[36] br[36] wl[65] vdd gnd cell_6t
Xbit_r66_c36 bl[36] br[36] wl[66] vdd gnd cell_6t
Xbit_r67_c36 bl[36] br[36] wl[67] vdd gnd cell_6t
Xbit_r68_c36 bl[36] br[36] wl[68] vdd gnd cell_6t
Xbit_r69_c36 bl[36] br[36] wl[69] vdd gnd cell_6t
Xbit_r70_c36 bl[36] br[36] wl[70] vdd gnd cell_6t
Xbit_r71_c36 bl[36] br[36] wl[71] vdd gnd cell_6t
Xbit_r72_c36 bl[36] br[36] wl[72] vdd gnd cell_6t
Xbit_r73_c36 bl[36] br[36] wl[73] vdd gnd cell_6t
Xbit_r74_c36 bl[36] br[36] wl[74] vdd gnd cell_6t
Xbit_r75_c36 bl[36] br[36] wl[75] vdd gnd cell_6t
Xbit_r76_c36 bl[36] br[36] wl[76] vdd gnd cell_6t
Xbit_r77_c36 bl[36] br[36] wl[77] vdd gnd cell_6t
Xbit_r78_c36 bl[36] br[36] wl[78] vdd gnd cell_6t
Xbit_r79_c36 bl[36] br[36] wl[79] vdd gnd cell_6t
Xbit_r80_c36 bl[36] br[36] wl[80] vdd gnd cell_6t
Xbit_r81_c36 bl[36] br[36] wl[81] vdd gnd cell_6t
Xbit_r82_c36 bl[36] br[36] wl[82] vdd gnd cell_6t
Xbit_r83_c36 bl[36] br[36] wl[83] vdd gnd cell_6t
Xbit_r84_c36 bl[36] br[36] wl[84] vdd gnd cell_6t
Xbit_r85_c36 bl[36] br[36] wl[85] vdd gnd cell_6t
Xbit_r86_c36 bl[36] br[36] wl[86] vdd gnd cell_6t
Xbit_r87_c36 bl[36] br[36] wl[87] vdd gnd cell_6t
Xbit_r88_c36 bl[36] br[36] wl[88] vdd gnd cell_6t
Xbit_r89_c36 bl[36] br[36] wl[89] vdd gnd cell_6t
Xbit_r90_c36 bl[36] br[36] wl[90] vdd gnd cell_6t
Xbit_r91_c36 bl[36] br[36] wl[91] vdd gnd cell_6t
Xbit_r92_c36 bl[36] br[36] wl[92] vdd gnd cell_6t
Xbit_r93_c36 bl[36] br[36] wl[93] vdd gnd cell_6t
Xbit_r94_c36 bl[36] br[36] wl[94] vdd gnd cell_6t
Xbit_r95_c36 bl[36] br[36] wl[95] vdd gnd cell_6t
Xbit_r96_c36 bl[36] br[36] wl[96] vdd gnd cell_6t
Xbit_r97_c36 bl[36] br[36] wl[97] vdd gnd cell_6t
Xbit_r98_c36 bl[36] br[36] wl[98] vdd gnd cell_6t
Xbit_r99_c36 bl[36] br[36] wl[99] vdd gnd cell_6t
Xbit_r100_c36 bl[36] br[36] wl[100] vdd gnd cell_6t
Xbit_r101_c36 bl[36] br[36] wl[101] vdd gnd cell_6t
Xbit_r102_c36 bl[36] br[36] wl[102] vdd gnd cell_6t
Xbit_r103_c36 bl[36] br[36] wl[103] vdd gnd cell_6t
Xbit_r104_c36 bl[36] br[36] wl[104] vdd gnd cell_6t
Xbit_r105_c36 bl[36] br[36] wl[105] vdd gnd cell_6t
Xbit_r106_c36 bl[36] br[36] wl[106] vdd gnd cell_6t
Xbit_r107_c36 bl[36] br[36] wl[107] vdd gnd cell_6t
Xbit_r108_c36 bl[36] br[36] wl[108] vdd gnd cell_6t
Xbit_r109_c36 bl[36] br[36] wl[109] vdd gnd cell_6t
Xbit_r110_c36 bl[36] br[36] wl[110] vdd gnd cell_6t
Xbit_r111_c36 bl[36] br[36] wl[111] vdd gnd cell_6t
Xbit_r112_c36 bl[36] br[36] wl[112] vdd gnd cell_6t
Xbit_r113_c36 bl[36] br[36] wl[113] vdd gnd cell_6t
Xbit_r114_c36 bl[36] br[36] wl[114] vdd gnd cell_6t
Xbit_r115_c36 bl[36] br[36] wl[115] vdd gnd cell_6t
Xbit_r116_c36 bl[36] br[36] wl[116] vdd gnd cell_6t
Xbit_r117_c36 bl[36] br[36] wl[117] vdd gnd cell_6t
Xbit_r118_c36 bl[36] br[36] wl[118] vdd gnd cell_6t
Xbit_r119_c36 bl[36] br[36] wl[119] vdd gnd cell_6t
Xbit_r120_c36 bl[36] br[36] wl[120] vdd gnd cell_6t
Xbit_r121_c36 bl[36] br[36] wl[121] vdd gnd cell_6t
Xbit_r122_c36 bl[36] br[36] wl[122] vdd gnd cell_6t
Xbit_r123_c36 bl[36] br[36] wl[123] vdd gnd cell_6t
Xbit_r124_c36 bl[36] br[36] wl[124] vdd gnd cell_6t
Xbit_r125_c36 bl[36] br[36] wl[125] vdd gnd cell_6t
Xbit_r126_c36 bl[36] br[36] wl[126] vdd gnd cell_6t
Xbit_r127_c36 bl[36] br[36] wl[127] vdd gnd cell_6t
Xbit_r128_c36 bl[36] br[36] wl[128] vdd gnd cell_6t
Xbit_r129_c36 bl[36] br[36] wl[129] vdd gnd cell_6t
Xbit_r130_c36 bl[36] br[36] wl[130] vdd gnd cell_6t
Xbit_r131_c36 bl[36] br[36] wl[131] vdd gnd cell_6t
Xbit_r132_c36 bl[36] br[36] wl[132] vdd gnd cell_6t
Xbit_r133_c36 bl[36] br[36] wl[133] vdd gnd cell_6t
Xbit_r134_c36 bl[36] br[36] wl[134] vdd gnd cell_6t
Xbit_r135_c36 bl[36] br[36] wl[135] vdd gnd cell_6t
Xbit_r136_c36 bl[36] br[36] wl[136] vdd gnd cell_6t
Xbit_r137_c36 bl[36] br[36] wl[137] vdd gnd cell_6t
Xbit_r138_c36 bl[36] br[36] wl[138] vdd gnd cell_6t
Xbit_r139_c36 bl[36] br[36] wl[139] vdd gnd cell_6t
Xbit_r140_c36 bl[36] br[36] wl[140] vdd gnd cell_6t
Xbit_r141_c36 bl[36] br[36] wl[141] vdd gnd cell_6t
Xbit_r142_c36 bl[36] br[36] wl[142] vdd gnd cell_6t
Xbit_r143_c36 bl[36] br[36] wl[143] vdd gnd cell_6t
Xbit_r144_c36 bl[36] br[36] wl[144] vdd gnd cell_6t
Xbit_r145_c36 bl[36] br[36] wl[145] vdd gnd cell_6t
Xbit_r146_c36 bl[36] br[36] wl[146] vdd gnd cell_6t
Xbit_r147_c36 bl[36] br[36] wl[147] vdd gnd cell_6t
Xbit_r148_c36 bl[36] br[36] wl[148] vdd gnd cell_6t
Xbit_r149_c36 bl[36] br[36] wl[149] vdd gnd cell_6t
Xbit_r150_c36 bl[36] br[36] wl[150] vdd gnd cell_6t
Xbit_r151_c36 bl[36] br[36] wl[151] vdd gnd cell_6t
Xbit_r152_c36 bl[36] br[36] wl[152] vdd gnd cell_6t
Xbit_r153_c36 bl[36] br[36] wl[153] vdd gnd cell_6t
Xbit_r154_c36 bl[36] br[36] wl[154] vdd gnd cell_6t
Xbit_r155_c36 bl[36] br[36] wl[155] vdd gnd cell_6t
Xbit_r156_c36 bl[36] br[36] wl[156] vdd gnd cell_6t
Xbit_r157_c36 bl[36] br[36] wl[157] vdd gnd cell_6t
Xbit_r158_c36 bl[36] br[36] wl[158] vdd gnd cell_6t
Xbit_r159_c36 bl[36] br[36] wl[159] vdd gnd cell_6t
Xbit_r160_c36 bl[36] br[36] wl[160] vdd gnd cell_6t
Xbit_r161_c36 bl[36] br[36] wl[161] vdd gnd cell_6t
Xbit_r162_c36 bl[36] br[36] wl[162] vdd gnd cell_6t
Xbit_r163_c36 bl[36] br[36] wl[163] vdd gnd cell_6t
Xbit_r164_c36 bl[36] br[36] wl[164] vdd gnd cell_6t
Xbit_r165_c36 bl[36] br[36] wl[165] vdd gnd cell_6t
Xbit_r166_c36 bl[36] br[36] wl[166] vdd gnd cell_6t
Xbit_r167_c36 bl[36] br[36] wl[167] vdd gnd cell_6t
Xbit_r168_c36 bl[36] br[36] wl[168] vdd gnd cell_6t
Xbit_r169_c36 bl[36] br[36] wl[169] vdd gnd cell_6t
Xbit_r170_c36 bl[36] br[36] wl[170] vdd gnd cell_6t
Xbit_r171_c36 bl[36] br[36] wl[171] vdd gnd cell_6t
Xbit_r172_c36 bl[36] br[36] wl[172] vdd gnd cell_6t
Xbit_r173_c36 bl[36] br[36] wl[173] vdd gnd cell_6t
Xbit_r174_c36 bl[36] br[36] wl[174] vdd gnd cell_6t
Xbit_r175_c36 bl[36] br[36] wl[175] vdd gnd cell_6t
Xbit_r176_c36 bl[36] br[36] wl[176] vdd gnd cell_6t
Xbit_r177_c36 bl[36] br[36] wl[177] vdd gnd cell_6t
Xbit_r178_c36 bl[36] br[36] wl[178] vdd gnd cell_6t
Xbit_r179_c36 bl[36] br[36] wl[179] vdd gnd cell_6t
Xbit_r180_c36 bl[36] br[36] wl[180] vdd gnd cell_6t
Xbit_r181_c36 bl[36] br[36] wl[181] vdd gnd cell_6t
Xbit_r182_c36 bl[36] br[36] wl[182] vdd gnd cell_6t
Xbit_r183_c36 bl[36] br[36] wl[183] vdd gnd cell_6t
Xbit_r184_c36 bl[36] br[36] wl[184] vdd gnd cell_6t
Xbit_r185_c36 bl[36] br[36] wl[185] vdd gnd cell_6t
Xbit_r186_c36 bl[36] br[36] wl[186] vdd gnd cell_6t
Xbit_r187_c36 bl[36] br[36] wl[187] vdd gnd cell_6t
Xbit_r188_c36 bl[36] br[36] wl[188] vdd gnd cell_6t
Xbit_r189_c36 bl[36] br[36] wl[189] vdd gnd cell_6t
Xbit_r190_c36 bl[36] br[36] wl[190] vdd gnd cell_6t
Xbit_r191_c36 bl[36] br[36] wl[191] vdd gnd cell_6t
Xbit_r192_c36 bl[36] br[36] wl[192] vdd gnd cell_6t
Xbit_r193_c36 bl[36] br[36] wl[193] vdd gnd cell_6t
Xbit_r194_c36 bl[36] br[36] wl[194] vdd gnd cell_6t
Xbit_r195_c36 bl[36] br[36] wl[195] vdd gnd cell_6t
Xbit_r196_c36 bl[36] br[36] wl[196] vdd gnd cell_6t
Xbit_r197_c36 bl[36] br[36] wl[197] vdd gnd cell_6t
Xbit_r198_c36 bl[36] br[36] wl[198] vdd gnd cell_6t
Xbit_r199_c36 bl[36] br[36] wl[199] vdd gnd cell_6t
Xbit_r200_c36 bl[36] br[36] wl[200] vdd gnd cell_6t
Xbit_r201_c36 bl[36] br[36] wl[201] vdd gnd cell_6t
Xbit_r202_c36 bl[36] br[36] wl[202] vdd gnd cell_6t
Xbit_r203_c36 bl[36] br[36] wl[203] vdd gnd cell_6t
Xbit_r204_c36 bl[36] br[36] wl[204] vdd gnd cell_6t
Xbit_r205_c36 bl[36] br[36] wl[205] vdd gnd cell_6t
Xbit_r206_c36 bl[36] br[36] wl[206] vdd gnd cell_6t
Xbit_r207_c36 bl[36] br[36] wl[207] vdd gnd cell_6t
Xbit_r208_c36 bl[36] br[36] wl[208] vdd gnd cell_6t
Xbit_r209_c36 bl[36] br[36] wl[209] vdd gnd cell_6t
Xbit_r210_c36 bl[36] br[36] wl[210] vdd gnd cell_6t
Xbit_r211_c36 bl[36] br[36] wl[211] vdd gnd cell_6t
Xbit_r212_c36 bl[36] br[36] wl[212] vdd gnd cell_6t
Xbit_r213_c36 bl[36] br[36] wl[213] vdd gnd cell_6t
Xbit_r214_c36 bl[36] br[36] wl[214] vdd gnd cell_6t
Xbit_r215_c36 bl[36] br[36] wl[215] vdd gnd cell_6t
Xbit_r216_c36 bl[36] br[36] wl[216] vdd gnd cell_6t
Xbit_r217_c36 bl[36] br[36] wl[217] vdd gnd cell_6t
Xbit_r218_c36 bl[36] br[36] wl[218] vdd gnd cell_6t
Xbit_r219_c36 bl[36] br[36] wl[219] vdd gnd cell_6t
Xbit_r220_c36 bl[36] br[36] wl[220] vdd gnd cell_6t
Xbit_r221_c36 bl[36] br[36] wl[221] vdd gnd cell_6t
Xbit_r222_c36 bl[36] br[36] wl[222] vdd gnd cell_6t
Xbit_r223_c36 bl[36] br[36] wl[223] vdd gnd cell_6t
Xbit_r224_c36 bl[36] br[36] wl[224] vdd gnd cell_6t
Xbit_r225_c36 bl[36] br[36] wl[225] vdd gnd cell_6t
Xbit_r226_c36 bl[36] br[36] wl[226] vdd gnd cell_6t
Xbit_r227_c36 bl[36] br[36] wl[227] vdd gnd cell_6t
Xbit_r228_c36 bl[36] br[36] wl[228] vdd gnd cell_6t
Xbit_r229_c36 bl[36] br[36] wl[229] vdd gnd cell_6t
Xbit_r230_c36 bl[36] br[36] wl[230] vdd gnd cell_6t
Xbit_r231_c36 bl[36] br[36] wl[231] vdd gnd cell_6t
Xbit_r232_c36 bl[36] br[36] wl[232] vdd gnd cell_6t
Xbit_r233_c36 bl[36] br[36] wl[233] vdd gnd cell_6t
Xbit_r234_c36 bl[36] br[36] wl[234] vdd gnd cell_6t
Xbit_r235_c36 bl[36] br[36] wl[235] vdd gnd cell_6t
Xbit_r236_c36 bl[36] br[36] wl[236] vdd gnd cell_6t
Xbit_r237_c36 bl[36] br[36] wl[237] vdd gnd cell_6t
Xbit_r238_c36 bl[36] br[36] wl[238] vdd gnd cell_6t
Xbit_r239_c36 bl[36] br[36] wl[239] vdd gnd cell_6t
Xbit_r240_c36 bl[36] br[36] wl[240] vdd gnd cell_6t
Xbit_r241_c36 bl[36] br[36] wl[241] vdd gnd cell_6t
Xbit_r242_c36 bl[36] br[36] wl[242] vdd gnd cell_6t
Xbit_r243_c36 bl[36] br[36] wl[243] vdd gnd cell_6t
Xbit_r244_c36 bl[36] br[36] wl[244] vdd gnd cell_6t
Xbit_r245_c36 bl[36] br[36] wl[245] vdd gnd cell_6t
Xbit_r246_c36 bl[36] br[36] wl[246] vdd gnd cell_6t
Xbit_r247_c36 bl[36] br[36] wl[247] vdd gnd cell_6t
Xbit_r248_c36 bl[36] br[36] wl[248] vdd gnd cell_6t
Xbit_r249_c36 bl[36] br[36] wl[249] vdd gnd cell_6t
Xbit_r250_c36 bl[36] br[36] wl[250] vdd gnd cell_6t
Xbit_r251_c36 bl[36] br[36] wl[251] vdd gnd cell_6t
Xbit_r252_c36 bl[36] br[36] wl[252] vdd gnd cell_6t
Xbit_r253_c36 bl[36] br[36] wl[253] vdd gnd cell_6t
Xbit_r254_c36 bl[36] br[36] wl[254] vdd gnd cell_6t
Xbit_r255_c36 bl[36] br[36] wl[255] vdd gnd cell_6t
Xbit_r256_c36 bl[36] br[36] wl[256] vdd gnd cell_6t
Xbit_r257_c36 bl[36] br[36] wl[257] vdd gnd cell_6t
Xbit_r258_c36 bl[36] br[36] wl[258] vdd gnd cell_6t
Xbit_r259_c36 bl[36] br[36] wl[259] vdd gnd cell_6t
Xbit_r260_c36 bl[36] br[36] wl[260] vdd gnd cell_6t
Xbit_r261_c36 bl[36] br[36] wl[261] vdd gnd cell_6t
Xbit_r262_c36 bl[36] br[36] wl[262] vdd gnd cell_6t
Xbit_r263_c36 bl[36] br[36] wl[263] vdd gnd cell_6t
Xbit_r264_c36 bl[36] br[36] wl[264] vdd gnd cell_6t
Xbit_r265_c36 bl[36] br[36] wl[265] vdd gnd cell_6t
Xbit_r266_c36 bl[36] br[36] wl[266] vdd gnd cell_6t
Xbit_r267_c36 bl[36] br[36] wl[267] vdd gnd cell_6t
Xbit_r268_c36 bl[36] br[36] wl[268] vdd gnd cell_6t
Xbit_r269_c36 bl[36] br[36] wl[269] vdd gnd cell_6t
Xbit_r270_c36 bl[36] br[36] wl[270] vdd gnd cell_6t
Xbit_r271_c36 bl[36] br[36] wl[271] vdd gnd cell_6t
Xbit_r272_c36 bl[36] br[36] wl[272] vdd gnd cell_6t
Xbit_r273_c36 bl[36] br[36] wl[273] vdd gnd cell_6t
Xbit_r274_c36 bl[36] br[36] wl[274] vdd gnd cell_6t
Xbit_r275_c36 bl[36] br[36] wl[275] vdd gnd cell_6t
Xbit_r276_c36 bl[36] br[36] wl[276] vdd gnd cell_6t
Xbit_r277_c36 bl[36] br[36] wl[277] vdd gnd cell_6t
Xbit_r278_c36 bl[36] br[36] wl[278] vdd gnd cell_6t
Xbit_r279_c36 bl[36] br[36] wl[279] vdd gnd cell_6t
Xbit_r280_c36 bl[36] br[36] wl[280] vdd gnd cell_6t
Xbit_r281_c36 bl[36] br[36] wl[281] vdd gnd cell_6t
Xbit_r282_c36 bl[36] br[36] wl[282] vdd gnd cell_6t
Xbit_r283_c36 bl[36] br[36] wl[283] vdd gnd cell_6t
Xbit_r284_c36 bl[36] br[36] wl[284] vdd gnd cell_6t
Xbit_r285_c36 bl[36] br[36] wl[285] vdd gnd cell_6t
Xbit_r286_c36 bl[36] br[36] wl[286] vdd gnd cell_6t
Xbit_r287_c36 bl[36] br[36] wl[287] vdd gnd cell_6t
Xbit_r288_c36 bl[36] br[36] wl[288] vdd gnd cell_6t
Xbit_r289_c36 bl[36] br[36] wl[289] vdd gnd cell_6t
Xbit_r290_c36 bl[36] br[36] wl[290] vdd gnd cell_6t
Xbit_r291_c36 bl[36] br[36] wl[291] vdd gnd cell_6t
Xbit_r292_c36 bl[36] br[36] wl[292] vdd gnd cell_6t
Xbit_r293_c36 bl[36] br[36] wl[293] vdd gnd cell_6t
Xbit_r294_c36 bl[36] br[36] wl[294] vdd gnd cell_6t
Xbit_r295_c36 bl[36] br[36] wl[295] vdd gnd cell_6t
Xbit_r296_c36 bl[36] br[36] wl[296] vdd gnd cell_6t
Xbit_r297_c36 bl[36] br[36] wl[297] vdd gnd cell_6t
Xbit_r298_c36 bl[36] br[36] wl[298] vdd gnd cell_6t
Xbit_r299_c36 bl[36] br[36] wl[299] vdd gnd cell_6t
Xbit_r300_c36 bl[36] br[36] wl[300] vdd gnd cell_6t
Xbit_r301_c36 bl[36] br[36] wl[301] vdd gnd cell_6t
Xbit_r302_c36 bl[36] br[36] wl[302] vdd gnd cell_6t
Xbit_r303_c36 bl[36] br[36] wl[303] vdd gnd cell_6t
Xbit_r304_c36 bl[36] br[36] wl[304] vdd gnd cell_6t
Xbit_r305_c36 bl[36] br[36] wl[305] vdd gnd cell_6t
Xbit_r306_c36 bl[36] br[36] wl[306] vdd gnd cell_6t
Xbit_r307_c36 bl[36] br[36] wl[307] vdd gnd cell_6t
Xbit_r308_c36 bl[36] br[36] wl[308] vdd gnd cell_6t
Xbit_r309_c36 bl[36] br[36] wl[309] vdd gnd cell_6t
Xbit_r310_c36 bl[36] br[36] wl[310] vdd gnd cell_6t
Xbit_r311_c36 bl[36] br[36] wl[311] vdd gnd cell_6t
Xbit_r312_c36 bl[36] br[36] wl[312] vdd gnd cell_6t
Xbit_r313_c36 bl[36] br[36] wl[313] vdd gnd cell_6t
Xbit_r314_c36 bl[36] br[36] wl[314] vdd gnd cell_6t
Xbit_r315_c36 bl[36] br[36] wl[315] vdd gnd cell_6t
Xbit_r316_c36 bl[36] br[36] wl[316] vdd gnd cell_6t
Xbit_r317_c36 bl[36] br[36] wl[317] vdd gnd cell_6t
Xbit_r318_c36 bl[36] br[36] wl[318] vdd gnd cell_6t
Xbit_r319_c36 bl[36] br[36] wl[319] vdd gnd cell_6t
Xbit_r320_c36 bl[36] br[36] wl[320] vdd gnd cell_6t
Xbit_r321_c36 bl[36] br[36] wl[321] vdd gnd cell_6t
Xbit_r322_c36 bl[36] br[36] wl[322] vdd gnd cell_6t
Xbit_r323_c36 bl[36] br[36] wl[323] vdd gnd cell_6t
Xbit_r324_c36 bl[36] br[36] wl[324] vdd gnd cell_6t
Xbit_r325_c36 bl[36] br[36] wl[325] vdd gnd cell_6t
Xbit_r326_c36 bl[36] br[36] wl[326] vdd gnd cell_6t
Xbit_r327_c36 bl[36] br[36] wl[327] vdd gnd cell_6t
Xbit_r328_c36 bl[36] br[36] wl[328] vdd gnd cell_6t
Xbit_r329_c36 bl[36] br[36] wl[329] vdd gnd cell_6t
Xbit_r330_c36 bl[36] br[36] wl[330] vdd gnd cell_6t
Xbit_r331_c36 bl[36] br[36] wl[331] vdd gnd cell_6t
Xbit_r332_c36 bl[36] br[36] wl[332] vdd gnd cell_6t
Xbit_r333_c36 bl[36] br[36] wl[333] vdd gnd cell_6t
Xbit_r334_c36 bl[36] br[36] wl[334] vdd gnd cell_6t
Xbit_r335_c36 bl[36] br[36] wl[335] vdd gnd cell_6t
Xbit_r336_c36 bl[36] br[36] wl[336] vdd gnd cell_6t
Xbit_r337_c36 bl[36] br[36] wl[337] vdd gnd cell_6t
Xbit_r338_c36 bl[36] br[36] wl[338] vdd gnd cell_6t
Xbit_r339_c36 bl[36] br[36] wl[339] vdd gnd cell_6t
Xbit_r340_c36 bl[36] br[36] wl[340] vdd gnd cell_6t
Xbit_r341_c36 bl[36] br[36] wl[341] vdd gnd cell_6t
Xbit_r342_c36 bl[36] br[36] wl[342] vdd gnd cell_6t
Xbit_r343_c36 bl[36] br[36] wl[343] vdd gnd cell_6t
Xbit_r344_c36 bl[36] br[36] wl[344] vdd gnd cell_6t
Xbit_r345_c36 bl[36] br[36] wl[345] vdd gnd cell_6t
Xbit_r346_c36 bl[36] br[36] wl[346] vdd gnd cell_6t
Xbit_r347_c36 bl[36] br[36] wl[347] vdd gnd cell_6t
Xbit_r348_c36 bl[36] br[36] wl[348] vdd gnd cell_6t
Xbit_r349_c36 bl[36] br[36] wl[349] vdd gnd cell_6t
Xbit_r350_c36 bl[36] br[36] wl[350] vdd gnd cell_6t
Xbit_r351_c36 bl[36] br[36] wl[351] vdd gnd cell_6t
Xbit_r352_c36 bl[36] br[36] wl[352] vdd gnd cell_6t
Xbit_r353_c36 bl[36] br[36] wl[353] vdd gnd cell_6t
Xbit_r354_c36 bl[36] br[36] wl[354] vdd gnd cell_6t
Xbit_r355_c36 bl[36] br[36] wl[355] vdd gnd cell_6t
Xbit_r356_c36 bl[36] br[36] wl[356] vdd gnd cell_6t
Xbit_r357_c36 bl[36] br[36] wl[357] vdd gnd cell_6t
Xbit_r358_c36 bl[36] br[36] wl[358] vdd gnd cell_6t
Xbit_r359_c36 bl[36] br[36] wl[359] vdd gnd cell_6t
Xbit_r360_c36 bl[36] br[36] wl[360] vdd gnd cell_6t
Xbit_r361_c36 bl[36] br[36] wl[361] vdd gnd cell_6t
Xbit_r362_c36 bl[36] br[36] wl[362] vdd gnd cell_6t
Xbit_r363_c36 bl[36] br[36] wl[363] vdd gnd cell_6t
Xbit_r364_c36 bl[36] br[36] wl[364] vdd gnd cell_6t
Xbit_r365_c36 bl[36] br[36] wl[365] vdd gnd cell_6t
Xbit_r366_c36 bl[36] br[36] wl[366] vdd gnd cell_6t
Xbit_r367_c36 bl[36] br[36] wl[367] vdd gnd cell_6t
Xbit_r368_c36 bl[36] br[36] wl[368] vdd gnd cell_6t
Xbit_r369_c36 bl[36] br[36] wl[369] vdd gnd cell_6t
Xbit_r370_c36 bl[36] br[36] wl[370] vdd gnd cell_6t
Xbit_r371_c36 bl[36] br[36] wl[371] vdd gnd cell_6t
Xbit_r372_c36 bl[36] br[36] wl[372] vdd gnd cell_6t
Xbit_r373_c36 bl[36] br[36] wl[373] vdd gnd cell_6t
Xbit_r374_c36 bl[36] br[36] wl[374] vdd gnd cell_6t
Xbit_r375_c36 bl[36] br[36] wl[375] vdd gnd cell_6t
Xbit_r376_c36 bl[36] br[36] wl[376] vdd gnd cell_6t
Xbit_r377_c36 bl[36] br[36] wl[377] vdd gnd cell_6t
Xbit_r378_c36 bl[36] br[36] wl[378] vdd gnd cell_6t
Xbit_r379_c36 bl[36] br[36] wl[379] vdd gnd cell_6t
Xbit_r380_c36 bl[36] br[36] wl[380] vdd gnd cell_6t
Xbit_r381_c36 bl[36] br[36] wl[381] vdd gnd cell_6t
Xbit_r382_c36 bl[36] br[36] wl[382] vdd gnd cell_6t
Xbit_r383_c36 bl[36] br[36] wl[383] vdd gnd cell_6t
Xbit_r384_c36 bl[36] br[36] wl[384] vdd gnd cell_6t
Xbit_r385_c36 bl[36] br[36] wl[385] vdd gnd cell_6t
Xbit_r386_c36 bl[36] br[36] wl[386] vdd gnd cell_6t
Xbit_r387_c36 bl[36] br[36] wl[387] vdd gnd cell_6t
Xbit_r388_c36 bl[36] br[36] wl[388] vdd gnd cell_6t
Xbit_r389_c36 bl[36] br[36] wl[389] vdd gnd cell_6t
Xbit_r390_c36 bl[36] br[36] wl[390] vdd gnd cell_6t
Xbit_r391_c36 bl[36] br[36] wl[391] vdd gnd cell_6t
Xbit_r392_c36 bl[36] br[36] wl[392] vdd gnd cell_6t
Xbit_r393_c36 bl[36] br[36] wl[393] vdd gnd cell_6t
Xbit_r394_c36 bl[36] br[36] wl[394] vdd gnd cell_6t
Xbit_r395_c36 bl[36] br[36] wl[395] vdd gnd cell_6t
Xbit_r396_c36 bl[36] br[36] wl[396] vdd gnd cell_6t
Xbit_r397_c36 bl[36] br[36] wl[397] vdd gnd cell_6t
Xbit_r398_c36 bl[36] br[36] wl[398] vdd gnd cell_6t
Xbit_r399_c36 bl[36] br[36] wl[399] vdd gnd cell_6t
Xbit_r400_c36 bl[36] br[36] wl[400] vdd gnd cell_6t
Xbit_r401_c36 bl[36] br[36] wl[401] vdd gnd cell_6t
Xbit_r402_c36 bl[36] br[36] wl[402] vdd gnd cell_6t
Xbit_r403_c36 bl[36] br[36] wl[403] vdd gnd cell_6t
Xbit_r404_c36 bl[36] br[36] wl[404] vdd gnd cell_6t
Xbit_r405_c36 bl[36] br[36] wl[405] vdd gnd cell_6t
Xbit_r406_c36 bl[36] br[36] wl[406] vdd gnd cell_6t
Xbit_r407_c36 bl[36] br[36] wl[407] vdd gnd cell_6t
Xbit_r408_c36 bl[36] br[36] wl[408] vdd gnd cell_6t
Xbit_r409_c36 bl[36] br[36] wl[409] vdd gnd cell_6t
Xbit_r410_c36 bl[36] br[36] wl[410] vdd gnd cell_6t
Xbit_r411_c36 bl[36] br[36] wl[411] vdd gnd cell_6t
Xbit_r412_c36 bl[36] br[36] wl[412] vdd gnd cell_6t
Xbit_r413_c36 bl[36] br[36] wl[413] vdd gnd cell_6t
Xbit_r414_c36 bl[36] br[36] wl[414] vdd gnd cell_6t
Xbit_r415_c36 bl[36] br[36] wl[415] vdd gnd cell_6t
Xbit_r416_c36 bl[36] br[36] wl[416] vdd gnd cell_6t
Xbit_r417_c36 bl[36] br[36] wl[417] vdd gnd cell_6t
Xbit_r418_c36 bl[36] br[36] wl[418] vdd gnd cell_6t
Xbit_r419_c36 bl[36] br[36] wl[419] vdd gnd cell_6t
Xbit_r420_c36 bl[36] br[36] wl[420] vdd gnd cell_6t
Xbit_r421_c36 bl[36] br[36] wl[421] vdd gnd cell_6t
Xbit_r422_c36 bl[36] br[36] wl[422] vdd gnd cell_6t
Xbit_r423_c36 bl[36] br[36] wl[423] vdd gnd cell_6t
Xbit_r424_c36 bl[36] br[36] wl[424] vdd gnd cell_6t
Xbit_r425_c36 bl[36] br[36] wl[425] vdd gnd cell_6t
Xbit_r426_c36 bl[36] br[36] wl[426] vdd gnd cell_6t
Xbit_r427_c36 bl[36] br[36] wl[427] vdd gnd cell_6t
Xbit_r428_c36 bl[36] br[36] wl[428] vdd gnd cell_6t
Xbit_r429_c36 bl[36] br[36] wl[429] vdd gnd cell_6t
Xbit_r430_c36 bl[36] br[36] wl[430] vdd gnd cell_6t
Xbit_r431_c36 bl[36] br[36] wl[431] vdd gnd cell_6t
Xbit_r432_c36 bl[36] br[36] wl[432] vdd gnd cell_6t
Xbit_r433_c36 bl[36] br[36] wl[433] vdd gnd cell_6t
Xbit_r434_c36 bl[36] br[36] wl[434] vdd gnd cell_6t
Xbit_r435_c36 bl[36] br[36] wl[435] vdd gnd cell_6t
Xbit_r436_c36 bl[36] br[36] wl[436] vdd gnd cell_6t
Xbit_r437_c36 bl[36] br[36] wl[437] vdd gnd cell_6t
Xbit_r438_c36 bl[36] br[36] wl[438] vdd gnd cell_6t
Xbit_r439_c36 bl[36] br[36] wl[439] vdd gnd cell_6t
Xbit_r440_c36 bl[36] br[36] wl[440] vdd gnd cell_6t
Xbit_r441_c36 bl[36] br[36] wl[441] vdd gnd cell_6t
Xbit_r442_c36 bl[36] br[36] wl[442] vdd gnd cell_6t
Xbit_r443_c36 bl[36] br[36] wl[443] vdd gnd cell_6t
Xbit_r444_c36 bl[36] br[36] wl[444] vdd gnd cell_6t
Xbit_r445_c36 bl[36] br[36] wl[445] vdd gnd cell_6t
Xbit_r446_c36 bl[36] br[36] wl[446] vdd gnd cell_6t
Xbit_r447_c36 bl[36] br[36] wl[447] vdd gnd cell_6t
Xbit_r448_c36 bl[36] br[36] wl[448] vdd gnd cell_6t
Xbit_r449_c36 bl[36] br[36] wl[449] vdd gnd cell_6t
Xbit_r450_c36 bl[36] br[36] wl[450] vdd gnd cell_6t
Xbit_r451_c36 bl[36] br[36] wl[451] vdd gnd cell_6t
Xbit_r452_c36 bl[36] br[36] wl[452] vdd gnd cell_6t
Xbit_r453_c36 bl[36] br[36] wl[453] vdd gnd cell_6t
Xbit_r454_c36 bl[36] br[36] wl[454] vdd gnd cell_6t
Xbit_r455_c36 bl[36] br[36] wl[455] vdd gnd cell_6t
Xbit_r456_c36 bl[36] br[36] wl[456] vdd gnd cell_6t
Xbit_r457_c36 bl[36] br[36] wl[457] vdd gnd cell_6t
Xbit_r458_c36 bl[36] br[36] wl[458] vdd gnd cell_6t
Xbit_r459_c36 bl[36] br[36] wl[459] vdd gnd cell_6t
Xbit_r460_c36 bl[36] br[36] wl[460] vdd gnd cell_6t
Xbit_r461_c36 bl[36] br[36] wl[461] vdd gnd cell_6t
Xbit_r462_c36 bl[36] br[36] wl[462] vdd gnd cell_6t
Xbit_r463_c36 bl[36] br[36] wl[463] vdd gnd cell_6t
Xbit_r464_c36 bl[36] br[36] wl[464] vdd gnd cell_6t
Xbit_r465_c36 bl[36] br[36] wl[465] vdd gnd cell_6t
Xbit_r466_c36 bl[36] br[36] wl[466] vdd gnd cell_6t
Xbit_r467_c36 bl[36] br[36] wl[467] vdd gnd cell_6t
Xbit_r468_c36 bl[36] br[36] wl[468] vdd gnd cell_6t
Xbit_r469_c36 bl[36] br[36] wl[469] vdd gnd cell_6t
Xbit_r470_c36 bl[36] br[36] wl[470] vdd gnd cell_6t
Xbit_r471_c36 bl[36] br[36] wl[471] vdd gnd cell_6t
Xbit_r472_c36 bl[36] br[36] wl[472] vdd gnd cell_6t
Xbit_r473_c36 bl[36] br[36] wl[473] vdd gnd cell_6t
Xbit_r474_c36 bl[36] br[36] wl[474] vdd gnd cell_6t
Xbit_r475_c36 bl[36] br[36] wl[475] vdd gnd cell_6t
Xbit_r476_c36 bl[36] br[36] wl[476] vdd gnd cell_6t
Xbit_r477_c36 bl[36] br[36] wl[477] vdd gnd cell_6t
Xbit_r478_c36 bl[36] br[36] wl[478] vdd gnd cell_6t
Xbit_r479_c36 bl[36] br[36] wl[479] vdd gnd cell_6t
Xbit_r480_c36 bl[36] br[36] wl[480] vdd gnd cell_6t
Xbit_r481_c36 bl[36] br[36] wl[481] vdd gnd cell_6t
Xbit_r482_c36 bl[36] br[36] wl[482] vdd gnd cell_6t
Xbit_r483_c36 bl[36] br[36] wl[483] vdd gnd cell_6t
Xbit_r484_c36 bl[36] br[36] wl[484] vdd gnd cell_6t
Xbit_r485_c36 bl[36] br[36] wl[485] vdd gnd cell_6t
Xbit_r486_c36 bl[36] br[36] wl[486] vdd gnd cell_6t
Xbit_r487_c36 bl[36] br[36] wl[487] vdd gnd cell_6t
Xbit_r488_c36 bl[36] br[36] wl[488] vdd gnd cell_6t
Xbit_r489_c36 bl[36] br[36] wl[489] vdd gnd cell_6t
Xbit_r490_c36 bl[36] br[36] wl[490] vdd gnd cell_6t
Xbit_r491_c36 bl[36] br[36] wl[491] vdd gnd cell_6t
Xbit_r492_c36 bl[36] br[36] wl[492] vdd gnd cell_6t
Xbit_r493_c36 bl[36] br[36] wl[493] vdd gnd cell_6t
Xbit_r494_c36 bl[36] br[36] wl[494] vdd gnd cell_6t
Xbit_r495_c36 bl[36] br[36] wl[495] vdd gnd cell_6t
Xbit_r496_c36 bl[36] br[36] wl[496] vdd gnd cell_6t
Xbit_r497_c36 bl[36] br[36] wl[497] vdd gnd cell_6t
Xbit_r498_c36 bl[36] br[36] wl[498] vdd gnd cell_6t
Xbit_r499_c36 bl[36] br[36] wl[499] vdd gnd cell_6t
Xbit_r500_c36 bl[36] br[36] wl[500] vdd gnd cell_6t
Xbit_r501_c36 bl[36] br[36] wl[501] vdd gnd cell_6t
Xbit_r502_c36 bl[36] br[36] wl[502] vdd gnd cell_6t
Xbit_r503_c36 bl[36] br[36] wl[503] vdd gnd cell_6t
Xbit_r504_c36 bl[36] br[36] wl[504] vdd gnd cell_6t
Xbit_r505_c36 bl[36] br[36] wl[505] vdd gnd cell_6t
Xbit_r506_c36 bl[36] br[36] wl[506] vdd gnd cell_6t
Xbit_r507_c36 bl[36] br[36] wl[507] vdd gnd cell_6t
Xbit_r508_c36 bl[36] br[36] wl[508] vdd gnd cell_6t
Xbit_r509_c36 bl[36] br[36] wl[509] vdd gnd cell_6t
Xbit_r510_c36 bl[36] br[36] wl[510] vdd gnd cell_6t
Xbit_r511_c36 bl[36] br[36] wl[511] vdd gnd cell_6t
Xbit_r0_c37 bl[37] br[37] wl[0] vdd gnd cell_6t
Xbit_r1_c37 bl[37] br[37] wl[1] vdd gnd cell_6t
Xbit_r2_c37 bl[37] br[37] wl[2] vdd gnd cell_6t
Xbit_r3_c37 bl[37] br[37] wl[3] vdd gnd cell_6t
Xbit_r4_c37 bl[37] br[37] wl[4] vdd gnd cell_6t
Xbit_r5_c37 bl[37] br[37] wl[5] vdd gnd cell_6t
Xbit_r6_c37 bl[37] br[37] wl[6] vdd gnd cell_6t
Xbit_r7_c37 bl[37] br[37] wl[7] vdd gnd cell_6t
Xbit_r8_c37 bl[37] br[37] wl[8] vdd gnd cell_6t
Xbit_r9_c37 bl[37] br[37] wl[9] vdd gnd cell_6t
Xbit_r10_c37 bl[37] br[37] wl[10] vdd gnd cell_6t
Xbit_r11_c37 bl[37] br[37] wl[11] vdd gnd cell_6t
Xbit_r12_c37 bl[37] br[37] wl[12] vdd gnd cell_6t
Xbit_r13_c37 bl[37] br[37] wl[13] vdd gnd cell_6t
Xbit_r14_c37 bl[37] br[37] wl[14] vdd gnd cell_6t
Xbit_r15_c37 bl[37] br[37] wl[15] vdd gnd cell_6t
Xbit_r16_c37 bl[37] br[37] wl[16] vdd gnd cell_6t
Xbit_r17_c37 bl[37] br[37] wl[17] vdd gnd cell_6t
Xbit_r18_c37 bl[37] br[37] wl[18] vdd gnd cell_6t
Xbit_r19_c37 bl[37] br[37] wl[19] vdd gnd cell_6t
Xbit_r20_c37 bl[37] br[37] wl[20] vdd gnd cell_6t
Xbit_r21_c37 bl[37] br[37] wl[21] vdd gnd cell_6t
Xbit_r22_c37 bl[37] br[37] wl[22] vdd gnd cell_6t
Xbit_r23_c37 bl[37] br[37] wl[23] vdd gnd cell_6t
Xbit_r24_c37 bl[37] br[37] wl[24] vdd gnd cell_6t
Xbit_r25_c37 bl[37] br[37] wl[25] vdd gnd cell_6t
Xbit_r26_c37 bl[37] br[37] wl[26] vdd gnd cell_6t
Xbit_r27_c37 bl[37] br[37] wl[27] vdd gnd cell_6t
Xbit_r28_c37 bl[37] br[37] wl[28] vdd gnd cell_6t
Xbit_r29_c37 bl[37] br[37] wl[29] vdd gnd cell_6t
Xbit_r30_c37 bl[37] br[37] wl[30] vdd gnd cell_6t
Xbit_r31_c37 bl[37] br[37] wl[31] vdd gnd cell_6t
Xbit_r32_c37 bl[37] br[37] wl[32] vdd gnd cell_6t
Xbit_r33_c37 bl[37] br[37] wl[33] vdd gnd cell_6t
Xbit_r34_c37 bl[37] br[37] wl[34] vdd gnd cell_6t
Xbit_r35_c37 bl[37] br[37] wl[35] vdd gnd cell_6t
Xbit_r36_c37 bl[37] br[37] wl[36] vdd gnd cell_6t
Xbit_r37_c37 bl[37] br[37] wl[37] vdd gnd cell_6t
Xbit_r38_c37 bl[37] br[37] wl[38] vdd gnd cell_6t
Xbit_r39_c37 bl[37] br[37] wl[39] vdd gnd cell_6t
Xbit_r40_c37 bl[37] br[37] wl[40] vdd gnd cell_6t
Xbit_r41_c37 bl[37] br[37] wl[41] vdd gnd cell_6t
Xbit_r42_c37 bl[37] br[37] wl[42] vdd gnd cell_6t
Xbit_r43_c37 bl[37] br[37] wl[43] vdd gnd cell_6t
Xbit_r44_c37 bl[37] br[37] wl[44] vdd gnd cell_6t
Xbit_r45_c37 bl[37] br[37] wl[45] vdd gnd cell_6t
Xbit_r46_c37 bl[37] br[37] wl[46] vdd gnd cell_6t
Xbit_r47_c37 bl[37] br[37] wl[47] vdd gnd cell_6t
Xbit_r48_c37 bl[37] br[37] wl[48] vdd gnd cell_6t
Xbit_r49_c37 bl[37] br[37] wl[49] vdd gnd cell_6t
Xbit_r50_c37 bl[37] br[37] wl[50] vdd gnd cell_6t
Xbit_r51_c37 bl[37] br[37] wl[51] vdd gnd cell_6t
Xbit_r52_c37 bl[37] br[37] wl[52] vdd gnd cell_6t
Xbit_r53_c37 bl[37] br[37] wl[53] vdd gnd cell_6t
Xbit_r54_c37 bl[37] br[37] wl[54] vdd gnd cell_6t
Xbit_r55_c37 bl[37] br[37] wl[55] vdd gnd cell_6t
Xbit_r56_c37 bl[37] br[37] wl[56] vdd gnd cell_6t
Xbit_r57_c37 bl[37] br[37] wl[57] vdd gnd cell_6t
Xbit_r58_c37 bl[37] br[37] wl[58] vdd gnd cell_6t
Xbit_r59_c37 bl[37] br[37] wl[59] vdd gnd cell_6t
Xbit_r60_c37 bl[37] br[37] wl[60] vdd gnd cell_6t
Xbit_r61_c37 bl[37] br[37] wl[61] vdd gnd cell_6t
Xbit_r62_c37 bl[37] br[37] wl[62] vdd gnd cell_6t
Xbit_r63_c37 bl[37] br[37] wl[63] vdd gnd cell_6t
Xbit_r64_c37 bl[37] br[37] wl[64] vdd gnd cell_6t
Xbit_r65_c37 bl[37] br[37] wl[65] vdd gnd cell_6t
Xbit_r66_c37 bl[37] br[37] wl[66] vdd gnd cell_6t
Xbit_r67_c37 bl[37] br[37] wl[67] vdd gnd cell_6t
Xbit_r68_c37 bl[37] br[37] wl[68] vdd gnd cell_6t
Xbit_r69_c37 bl[37] br[37] wl[69] vdd gnd cell_6t
Xbit_r70_c37 bl[37] br[37] wl[70] vdd gnd cell_6t
Xbit_r71_c37 bl[37] br[37] wl[71] vdd gnd cell_6t
Xbit_r72_c37 bl[37] br[37] wl[72] vdd gnd cell_6t
Xbit_r73_c37 bl[37] br[37] wl[73] vdd gnd cell_6t
Xbit_r74_c37 bl[37] br[37] wl[74] vdd gnd cell_6t
Xbit_r75_c37 bl[37] br[37] wl[75] vdd gnd cell_6t
Xbit_r76_c37 bl[37] br[37] wl[76] vdd gnd cell_6t
Xbit_r77_c37 bl[37] br[37] wl[77] vdd gnd cell_6t
Xbit_r78_c37 bl[37] br[37] wl[78] vdd gnd cell_6t
Xbit_r79_c37 bl[37] br[37] wl[79] vdd gnd cell_6t
Xbit_r80_c37 bl[37] br[37] wl[80] vdd gnd cell_6t
Xbit_r81_c37 bl[37] br[37] wl[81] vdd gnd cell_6t
Xbit_r82_c37 bl[37] br[37] wl[82] vdd gnd cell_6t
Xbit_r83_c37 bl[37] br[37] wl[83] vdd gnd cell_6t
Xbit_r84_c37 bl[37] br[37] wl[84] vdd gnd cell_6t
Xbit_r85_c37 bl[37] br[37] wl[85] vdd gnd cell_6t
Xbit_r86_c37 bl[37] br[37] wl[86] vdd gnd cell_6t
Xbit_r87_c37 bl[37] br[37] wl[87] vdd gnd cell_6t
Xbit_r88_c37 bl[37] br[37] wl[88] vdd gnd cell_6t
Xbit_r89_c37 bl[37] br[37] wl[89] vdd gnd cell_6t
Xbit_r90_c37 bl[37] br[37] wl[90] vdd gnd cell_6t
Xbit_r91_c37 bl[37] br[37] wl[91] vdd gnd cell_6t
Xbit_r92_c37 bl[37] br[37] wl[92] vdd gnd cell_6t
Xbit_r93_c37 bl[37] br[37] wl[93] vdd gnd cell_6t
Xbit_r94_c37 bl[37] br[37] wl[94] vdd gnd cell_6t
Xbit_r95_c37 bl[37] br[37] wl[95] vdd gnd cell_6t
Xbit_r96_c37 bl[37] br[37] wl[96] vdd gnd cell_6t
Xbit_r97_c37 bl[37] br[37] wl[97] vdd gnd cell_6t
Xbit_r98_c37 bl[37] br[37] wl[98] vdd gnd cell_6t
Xbit_r99_c37 bl[37] br[37] wl[99] vdd gnd cell_6t
Xbit_r100_c37 bl[37] br[37] wl[100] vdd gnd cell_6t
Xbit_r101_c37 bl[37] br[37] wl[101] vdd gnd cell_6t
Xbit_r102_c37 bl[37] br[37] wl[102] vdd gnd cell_6t
Xbit_r103_c37 bl[37] br[37] wl[103] vdd gnd cell_6t
Xbit_r104_c37 bl[37] br[37] wl[104] vdd gnd cell_6t
Xbit_r105_c37 bl[37] br[37] wl[105] vdd gnd cell_6t
Xbit_r106_c37 bl[37] br[37] wl[106] vdd gnd cell_6t
Xbit_r107_c37 bl[37] br[37] wl[107] vdd gnd cell_6t
Xbit_r108_c37 bl[37] br[37] wl[108] vdd gnd cell_6t
Xbit_r109_c37 bl[37] br[37] wl[109] vdd gnd cell_6t
Xbit_r110_c37 bl[37] br[37] wl[110] vdd gnd cell_6t
Xbit_r111_c37 bl[37] br[37] wl[111] vdd gnd cell_6t
Xbit_r112_c37 bl[37] br[37] wl[112] vdd gnd cell_6t
Xbit_r113_c37 bl[37] br[37] wl[113] vdd gnd cell_6t
Xbit_r114_c37 bl[37] br[37] wl[114] vdd gnd cell_6t
Xbit_r115_c37 bl[37] br[37] wl[115] vdd gnd cell_6t
Xbit_r116_c37 bl[37] br[37] wl[116] vdd gnd cell_6t
Xbit_r117_c37 bl[37] br[37] wl[117] vdd gnd cell_6t
Xbit_r118_c37 bl[37] br[37] wl[118] vdd gnd cell_6t
Xbit_r119_c37 bl[37] br[37] wl[119] vdd gnd cell_6t
Xbit_r120_c37 bl[37] br[37] wl[120] vdd gnd cell_6t
Xbit_r121_c37 bl[37] br[37] wl[121] vdd gnd cell_6t
Xbit_r122_c37 bl[37] br[37] wl[122] vdd gnd cell_6t
Xbit_r123_c37 bl[37] br[37] wl[123] vdd gnd cell_6t
Xbit_r124_c37 bl[37] br[37] wl[124] vdd gnd cell_6t
Xbit_r125_c37 bl[37] br[37] wl[125] vdd gnd cell_6t
Xbit_r126_c37 bl[37] br[37] wl[126] vdd gnd cell_6t
Xbit_r127_c37 bl[37] br[37] wl[127] vdd gnd cell_6t
Xbit_r128_c37 bl[37] br[37] wl[128] vdd gnd cell_6t
Xbit_r129_c37 bl[37] br[37] wl[129] vdd gnd cell_6t
Xbit_r130_c37 bl[37] br[37] wl[130] vdd gnd cell_6t
Xbit_r131_c37 bl[37] br[37] wl[131] vdd gnd cell_6t
Xbit_r132_c37 bl[37] br[37] wl[132] vdd gnd cell_6t
Xbit_r133_c37 bl[37] br[37] wl[133] vdd gnd cell_6t
Xbit_r134_c37 bl[37] br[37] wl[134] vdd gnd cell_6t
Xbit_r135_c37 bl[37] br[37] wl[135] vdd gnd cell_6t
Xbit_r136_c37 bl[37] br[37] wl[136] vdd gnd cell_6t
Xbit_r137_c37 bl[37] br[37] wl[137] vdd gnd cell_6t
Xbit_r138_c37 bl[37] br[37] wl[138] vdd gnd cell_6t
Xbit_r139_c37 bl[37] br[37] wl[139] vdd gnd cell_6t
Xbit_r140_c37 bl[37] br[37] wl[140] vdd gnd cell_6t
Xbit_r141_c37 bl[37] br[37] wl[141] vdd gnd cell_6t
Xbit_r142_c37 bl[37] br[37] wl[142] vdd gnd cell_6t
Xbit_r143_c37 bl[37] br[37] wl[143] vdd gnd cell_6t
Xbit_r144_c37 bl[37] br[37] wl[144] vdd gnd cell_6t
Xbit_r145_c37 bl[37] br[37] wl[145] vdd gnd cell_6t
Xbit_r146_c37 bl[37] br[37] wl[146] vdd gnd cell_6t
Xbit_r147_c37 bl[37] br[37] wl[147] vdd gnd cell_6t
Xbit_r148_c37 bl[37] br[37] wl[148] vdd gnd cell_6t
Xbit_r149_c37 bl[37] br[37] wl[149] vdd gnd cell_6t
Xbit_r150_c37 bl[37] br[37] wl[150] vdd gnd cell_6t
Xbit_r151_c37 bl[37] br[37] wl[151] vdd gnd cell_6t
Xbit_r152_c37 bl[37] br[37] wl[152] vdd gnd cell_6t
Xbit_r153_c37 bl[37] br[37] wl[153] vdd gnd cell_6t
Xbit_r154_c37 bl[37] br[37] wl[154] vdd gnd cell_6t
Xbit_r155_c37 bl[37] br[37] wl[155] vdd gnd cell_6t
Xbit_r156_c37 bl[37] br[37] wl[156] vdd gnd cell_6t
Xbit_r157_c37 bl[37] br[37] wl[157] vdd gnd cell_6t
Xbit_r158_c37 bl[37] br[37] wl[158] vdd gnd cell_6t
Xbit_r159_c37 bl[37] br[37] wl[159] vdd gnd cell_6t
Xbit_r160_c37 bl[37] br[37] wl[160] vdd gnd cell_6t
Xbit_r161_c37 bl[37] br[37] wl[161] vdd gnd cell_6t
Xbit_r162_c37 bl[37] br[37] wl[162] vdd gnd cell_6t
Xbit_r163_c37 bl[37] br[37] wl[163] vdd gnd cell_6t
Xbit_r164_c37 bl[37] br[37] wl[164] vdd gnd cell_6t
Xbit_r165_c37 bl[37] br[37] wl[165] vdd gnd cell_6t
Xbit_r166_c37 bl[37] br[37] wl[166] vdd gnd cell_6t
Xbit_r167_c37 bl[37] br[37] wl[167] vdd gnd cell_6t
Xbit_r168_c37 bl[37] br[37] wl[168] vdd gnd cell_6t
Xbit_r169_c37 bl[37] br[37] wl[169] vdd gnd cell_6t
Xbit_r170_c37 bl[37] br[37] wl[170] vdd gnd cell_6t
Xbit_r171_c37 bl[37] br[37] wl[171] vdd gnd cell_6t
Xbit_r172_c37 bl[37] br[37] wl[172] vdd gnd cell_6t
Xbit_r173_c37 bl[37] br[37] wl[173] vdd gnd cell_6t
Xbit_r174_c37 bl[37] br[37] wl[174] vdd gnd cell_6t
Xbit_r175_c37 bl[37] br[37] wl[175] vdd gnd cell_6t
Xbit_r176_c37 bl[37] br[37] wl[176] vdd gnd cell_6t
Xbit_r177_c37 bl[37] br[37] wl[177] vdd gnd cell_6t
Xbit_r178_c37 bl[37] br[37] wl[178] vdd gnd cell_6t
Xbit_r179_c37 bl[37] br[37] wl[179] vdd gnd cell_6t
Xbit_r180_c37 bl[37] br[37] wl[180] vdd gnd cell_6t
Xbit_r181_c37 bl[37] br[37] wl[181] vdd gnd cell_6t
Xbit_r182_c37 bl[37] br[37] wl[182] vdd gnd cell_6t
Xbit_r183_c37 bl[37] br[37] wl[183] vdd gnd cell_6t
Xbit_r184_c37 bl[37] br[37] wl[184] vdd gnd cell_6t
Xbit_r185_c37 bl[37] br[37] wl[185] vdd gnd cell_6t
Xbit_r186_c37 bl[37] br[37] wl[186] vdd gnd cell_6t
Xbit_r187_c37 bl[37] br[37] wl[187] vdd gnd cell_6t
Xbit_r188_c37 bl[37] br[37] wl[188] vdd gnd cell_6t
Xbit_r189_c37 bl[37] br[37] wl[189] vdd gnd cell_6t
Xbit_r190_c37 bl[37] br[37] wl[190] vdd gnd cell_6t
Xbit_r191_c37 bl[37] br[37] wl[191] vdd gnd cell_6t
Xbit_r192_c37 bl[37] br[37] wl[192] vdd gnd cell_6t
Xbit_r193_c37 bl[37] br[37] wl[193] vdd gnd cell_6t
Xbit_r194_c37 bl[37] br[37] wl[194] vdd gnd cell_6t
Xbit_r195_c37 bl[37] br[37] wl[195] vdd gnd cell_6t
Xbit_r196_c37 bl[37] br[37] wl[196] vdd gnd cell_6t
Xbit_r197_c37 bl[37] br[37] wl[197] vdd gnd cell_6t
Xbit_r198_c37 bl[37] br[37] wl[198] vdd gnd cell_6t
Xbit_r199_c37 bl[37] br[37] wl[199] vdd gnd cell_6t
Xbit_r200_c37 bl[37] br[37] wl[200] vdd gnd cell_6t
Xbit_r201_c37 bl[37] br[37] wl[201] vdd gnd cell_6t
Xbit_r202_c37 bl[37] br[37] wl[202] vdd gnd cell_6t
Xbit_r203_c37 bl[37] br[37] wl[203] vdd gnd cell_6t
Xbit_r204_c37 bl[37] br[37] wl[204] vdd gnd cell_6t
Xbit_r205_c37 bl[37] br[37] wl[205] vdd gnd cell_6t
Xbit_r206_c37 bl[37] br[37] wl[206] vdd gnd cell_6t
Xbit_r207_c37 bl[37] br[37] wl[207] vdd gnd cell_6t
Xbit_r208_c37 bl[37] br[37] wl[208] vdd gnd cell_6t
Xbit_r209_c37 bl[37] br[37] wl[209] vdd gnd cell_6t
Xbit_r210_c37 bl[37] br[37] wl[210] vdd gnd cell_6t
Xbit_r211_c37 bl[37] br[37] wl[211] vdd gnd cell_6t
Xbit_r212_c37 bl[37] br[37] wl[212] vdd gnd cell_6t
Xbit_r213_c37 bl[37] br[37] wl[213] vdd gnd cell_6t
Xbit_r214_c37 bl[37] br[37] wl[214] vdd gnd cell_6t
Xbit_r215_c37 bl[37] br[37] wl[215] vdd gnd cell_6t
Xbit_r216_c37 bl[37] br[37] wl[216] vdd gnd cell_6t
Xbit_r217_c37 bl[37] br[37] wl[217] vdd gnd cell_6t
Xbit_r218_c37 bl[37] br[37] wl[218] vdd gnd cell_6t
Xbit_r219_c37 bl[37] br[37] wl[219] vdd gnd cell_6t
Xbit_r220_c37 bl[37] br[37] wl[220] vdd gnd cell_6t
Xbit_r221_c37 bl[37] br[37] wl[221] vdd gnd cell_6t
Xbit_r222_c37 bl[37] br[37] wl[222] vdd gnd cell_6t
Xbit_r223_c37 bl[37] br[37] wl[223] vdd gnd cell_6t
Xbit_r224_c37 bl[37] br[37] wl[224] vdd gnd cell_6t
Xbit_r225_c37 bl[37] br[37] wl[225] vdd gnd cell_6t
Xbit_r226_c37 bl[37] br[37] wl[226] vdd gnd cell_6t
Xbit_r227_c37 bl[37] br[37] wl[227] vdd gnd cell_6t
Xbit_r228_c37 bl[37] br[37] wl[228] vdd gnd cell_6t
Xbit_r229_c37 bl[37] br[37] wl[229] vdd gnd cell_6t
Xbit_r230_c37 bl[37] br[37] wl[230] vdd gnd cell_6t
Xbit_r231_c37 bl[37] br[37] wl[231] vdd gnd cell_6t
Xbit_r232_c37 bl[37] br[37] wl[232] vdd gnd cell_6t
Xbit_r233_c37 bl[37] br[37] wl[233] vdd gnd cell_6t
Xbit_r234_c37 bl[37] br[37] wl[234] vdd gnd cell_6t
Xbit_r235_c37 bl[37] br[37] wl[235] vdd gnd cell_6t
Xbit_r236_c37 bl[37] br[37] wl[236] vdd gnd cell_6t
Xbit_r237_c37 bl[37] br[37] wl[237] vdd gnd cell_6t
Xbit_r238_c37 bl[37] br[37] wl[238] vdd gnd cell_6t
Xbit_r239_c37 bl[37] br[37] wl[239] vdd gnd cell_6t
Xbit_r240_c37 bl[37] br[37] wl[240] vdd gnd cell_6t
Xbit_r241_c37 bl[37] br[37] wl[241] vdd gnd cell_6t
Xbit_r242_c37 bl[37] br[37] wl[242] vdd gnd cell_6t
Xbit_r243_c37 bl[37] br[37] wl[243] vdd gnd cell_6t
Xbit_r244_c37 bl[37] br[37] wl[244] vdd gnd cell_6t
Xbit_r245_c37 bl[37] br[37] wl[245] vdd gnd cell_6t
Xbit_r246_c37 bl[37] br[37] wl[246] vdd gnd cell_6t
Xbit_r247_c37 bl[37] br[37] wl[247] vdd gnd cell_6t
Xbit_r248_c37 bl[37] br[37] wl[248] vdd gnd cell_6t
Xbit_r249_c37 bl[37] br[37] wl[249] vdd gnd cell_6t
Xbit_r250_c37 bl[37] br[37] wl[250] vdd gnd cell_6t
Xbit_r251_c37 bl[37] br[37] wl[251] vdd gnd cell_6t
Xbit_r252_c37 bl[37] br[37] wl[252] vdd gnd cell_6t
Xbit_r253_c37 bl[37] br[37] wl[253] vdd gnd cell_6t
Xbit_r254_c37 bl[37] br[37] wl[254] vdd gnd cell_6t
Xbit_r255_c37 bl[37] br[37] wl[255] vdd gnd cell_6t
Xbit_r256_c37 bl[37] br[37] wl[256] vdd gnd cell_6t
Xbit_r257_c37 bl[37] br[37] wl[257] vdd gnd cell_6t
Xbit_r258_c37 bl[37] br[37] wl[258] vdd gnd cell_6t
Xbit_r259_c37 bl[37] br[37] wl[259] vdd gnd cell_6t
Xbit_r260_c37 bl[37] br[37] wl[260] vdd gnd cell_6t
Xbit_r261_c37 bl[37] br[37] wl[261] vdd gnd cell_6t
Xbit_r262_c37 bl[37] br[37] wl[262] vdd gnd cell_6t
Xbit_r263_c37 bl[37] br[37] wl[263] vdd gnd cell_6t
Xbit_r264_c37 bl[37] br[37] wl[264] vdd gnd cell_6t
Xbit_r265_c37 bl[37] br[37] wl[265] vdd gnd cell_6t
Xbit_r266_c37 bl[37] br[37] wl[266] vdd gnd cell_6t
Xbit_r267_c37 bl[37] br[37] wl[267] vdd gnd cell_6t
Xbit_r268_c37 bl[37] br[37] wl[268] vdd gnd cell_6t
Xbit_r269_c37 bl[37] br[37] wl[269] vdd gnd cell_6t
Xbit_r270_c37 bl[37] br[37] wl[270] vdd gnd cell_6t
Xbit_r271_c37 bl[37] br[37] wl[271] vdd gnd cell_6t
Xbit_r272_c37 bl[37] br[37] wl[272] vdd gnd cell_6t
Xbit_r273_c37 bl[37] br[37] wl[273] vdd gnd cell_6t
Xbit_r274_c37 bl[37] br[37] wl[274] vdd gnd cell_6t
Xbit_r275_c37 bl[37] br[37] wl[275] vdd gnd cell_6t
Xbit_r276_c37 bl[37] br[37] wl[276] vdd gnd cell_6t
Xbit_r277_c37 bl[37] br[37] wl[277] vdd gnd cell_6t
Xbit_r278_c37 bl[37] br[37] wl[278] vdd gnd cell_6t
Xbit_r279_c37 bl[37] br[37] wl[279] vdd gnd cell_6t
Xbit_r280_c37 bl[37] br[37] wl[280] vdd gnd cell_6t
Xbit_r281_c37 bl[37] br[37] wl[281] vdd gnd cell_6t
Xbit_r282_c37 bl[37] br[37] wl[282] vdd gnd cell_6t
Xbit_r283_c37 bl[37] br[37] wl[283] vdd gnd cell_6t
Xbit_r284_c37 bl[37] br[37] wl[284] vdd gnd cell_6t
Xbit_r285_c37 bl[37] br[37] wl[285] vdd gnd cell_6t
Xbit_r286_c37 bl[37] br[37] wl[286] vdd gnd cell_6t
Xbit_r287_c37 bl[37] br[37] wl[287] vdd gnd cell_6t
Xbit_r288_c37 bl[37] br[37] wl[288] vdd gnd cell_6t
Xbit_r289_c37 bl[37] br[37] wl[289] vdd gnd cell_6t
Xbit_r290_c37 bl[37] br[37] wl[290] vdd gnd cell_6t
Xbit_r291_c37 bl[37] br[37] wl[291] vdd gnd cell_6t
Xbit_r292_c37 bl[37] br[37] wl[292] vdd gnd cell_6t
Xbit_r293_c37 bl[37] br[37] wl[293] vdd gnd cell_6t
Xbit_r294_c37 bl[37] br[37] wl[294] vdd gnd cell_6t
Xbit_r295_c37 bl[37] br[37] wl[295] vdd gnd cell_6t
Xbit_r296_c37 bl[37] br[37] wl[296] vdd gnd cell_6t
Xbit_r297_c37 bl[37] br[37] wl[297] vdd gnd cell_6t
Xbit_r298_c37 bl[37] br[37] wl[298] vdd gnd cell_6t
Xbit_r299_c37 bl[37] br[37] wl[299] vdd gnd cell_6t
Xbit_r300_c37 bl[37] br[37] wl[300] vdd gnd cell_6t
Xbit_r301_c37 bl[37] br[37] wl[301] vdd gnd cell_6t
Xbit_r302_c37 bl[37] br[37] wl[302] vdd gnd cell_6t
Xbit_r303_c37 bl[37] br[37] wl[303] vdd gnd cell_6t
Xbit_r304_c37 bl[37] br[37] wl[304] vdd gnd cell_6t
Xbit_r305_c37 bl[37] br[37] wl[305] vdd gnd cell_6t
Xbit_r306_c37 bl[37] br[37] wl[306] vdd gnd cell_6t
Xbit_r307_c37 bl[37] br[37] wl[307] vdd gnd cell_6t
Xbit_r308_c37 bl[37] br[37] wl[308] vdd gnd cell_6t
Xbit_r309_c37 bl[37] br[37] wl[309] vdd gnd cell_6t
Xbit_r310_c37 bl[37] br[37] wl[310] vdd gnd cell_6t
Xbit_r311_c37 bl[37] br[37] wl[311] vdd gnd cell_6t
Xbit_r312_c37 bl[37] br[37] wl[312] vdd gnd cell_6t
Xbit_r313_c37 bl[37] br[37] wl[313] vdd gnd cell_6t
Xbit_r314_c37 bl[37] br[37] wl[314] vdd gnd cell_6t
Xbit_r315_c37 bl[37] br[37] wl[315] vdd gnd cell_6t
Xbit_r316_c37 bl[37] br[37] wl[316] vdd gnd cell_6t
Xbit_r317_c37 bl[37] br[37] wl[317] vdd gnd cell_6t
Xbit_r318_c37 bl[37] br[37] wl[318] vdd gnd cell_6t
Xbit_r319_c37 bl[37] br[37] wl[319] vdd gnd cell_6t
Xbit_r320_c37 bl[37] br[37] wl[320] vdd gnd cell_6t
Xbit_r321_c37 bl[37] br[37] wl[321] vdd gnd cell_6t
Xbit_r322_c37 bl[37] br[37] wl[322] vdd gnd cell_6t
Xbit_r323_c37 bl[37] br[37] wl[323] vdd gnd cell_6t
Xbit_r324_c37 bl[37] br[37] wl[324] vdd gnd cell_6t
Xbit_r325_c37 bl[37] br[37] wl[325] vdd gnd cell_6t
Xbit_r326_c37 bl[37] br[37] wl[326] vdd gnd cell_6t
Xbit_r327_c37 bl[37] br[37] wl[327] vdd gnd cell_6t
Xbit_r328_c37 bl[37] br[37] wl[328] vdd gnd cell_6t
Xbit_r329_c37 bl[37] br[37] wl[329] vdd gnd cell_6t
Xbit_r330_c37 bl[37] br[37] wl[330] vdd gnd cell_6t
Xbit_r331_c37 bl[37] br[37] wl[331] vdd gnd cell_6t
Xbit_r332_c37 bl[37] br[37] wl[332] vdd gnd cell_6t
Xbit_r333_c37 bl[37] br[37] wl[333] vdd gnd cell_6t
Xbit_r334_c37 bl[37] br[37] wl[334] vdd gnd cell_6t
Xbit_r335_c37 bl[37] br[37] wl[335] vdd gnd cell_6t
Xbit_r336_c37 bl[37] br[37] wl[336] vdd gnd cell_6t
Xbit_r337_c37 bl[37] br[37] wl[337] vdd gnd cell_6t
Xbit_r338_c37 bl[37] br[37] wl[338] vdd gnd cell_6t
Xbit_r339_c37 bl[37] br[37] wl[339] vdd gnd cell_6t
Xbit_r340_c37 bl[37] br[37] wl[340] vdd gnd cell_6t
Xbit_r341_c37 bl[37] br[37] wl[341] vdd gnd cell_6t
Xbit_r342_c37 bl[37] br[37] wl[342] vdd gnd cell_6t
Xbit_r343_c37 bl[37] br[37] wl[343] vdd gnd cell_6t
Xbit_r344_c37 bl[37] br[37] wl[344] vdd gnd cell_6t
Xbit_r345_c37 bl[37] br[37] wl[345] vdd gnd cell_6t
Xbit_r346_c37 bl[37] br[37] wl[346] vdd gnd cell_6t
Xbit_r347_c37 bl[37] br[37] wl[347] vdd gnd cell_6t
Xbit_r348_c37 bl[37] br[37] wl[348] vdd gnd cell_6t
Xbit_r349_c37 bl[37] br[37] wl[349] vdd gnd cell_6t
Xbit_r350_c37 bl[37] br[37] wl[350] vdd gnd cell_6t
Xbit_r351_c37 bl[37] br[37] wl[351] vdd gnd cell_6t
Xbit_r352_c37 bl[37] br[37] wl[352] vdd gnd cell_6t
Xbit_r353_c37 bl[37] br[37] wl[353] vdd gnd cell_6t
Xbit_r354_c37 bl[37] br[37] wl[354] vdd gnd cell_6t
Xbit_r355_c37 bl[37] br[37] wl[355] vdd gnd cell_6t
Xbit_r356_c37 bl[37] br[37] wl[356] vdd gnd cell_6t
Xbit_r357_c37 bl[37] br[37] wl[357] vdd gnd cell_6t
Xbit_r358_c37 bl[37] br[37] wl[358] vdd gnd cell_6t
Xbit_r359_c37 bl[37] br[37] wl[359] vdd gnd cell_6t
Xbit_r360_c37 bl[37] br[37] wl[360] vdd gnd cell_6t
Xbit_r361_c37 bl[37] br[37] wl[361] vdd gnd cell_6t
Xbit_r362_c37 bl[37] br[37] wl[362] vdd gnd cell_6t
Xbit_r363_c37 bl[37] br[37] wl[363] vdd gnd cell_6t
Xbit_r364_c37 bl[37] br[37] wl[364] vdd gnd cell_6t
Xbit_r365_c37 bl[37] br[37] wl[365] vdd gnd cell_6t
Xbit_r366_c37 bl[37] br[37] wl[366] vdd gnd cell_6t
Xbit_r367_c37 bl[37] br[37] wl[367] vdd gnd cell_6t
Xbit_r368_c37 bl[37] br[37] wl[368] vdd gnd cell_6t
Xbit_r369_c37 bl[37] br[37] wl[369] vdd gnd cell_6t
Xbit_r370_c37 bl[37] br[37] wl[370] vdd gnd cell_6t
Xbit_r371_c37 bl[37] br[37] wl[371] vdd gnd cell_6t
Xbit_r372_c37 bl[37] br[37] wl[372] vdd gnd cell_6t
Xbit_r373_c37 bl[37] br[37] wl[373] vdd gnd cell_6t
Xbit_r374_c37 bl[37] br[37] wl[374] vdd gnd cell_6t
Xbit_r375_c37 bl[37] br[37] wl[375] vdd gnd cell_6t
Xbit_r376_c37 bl[37] br[37] wl[376] vdd gnd cell_6t
Xbit_r377_c37 bl[37] br[37] wl[377] vdd gnd cell_6t
Xbit_r378_c37 bl[37] br[37] wl[378] vdd gnd cell_6t
Xbit_r379_c37 bl[37] br[37] wl[379] vdd gnd cell_6t
Xbit_r380_c37 bl[37] br[37] wl[380] vdd gnd cell_6t
Xbit_r381_c37 bl[37] br[37] wl[381] vdd gnd cell_6t
Xbit_r382_c37 bl[37] br[37] wl[382] vdd gnd cell_6t
Xbit_r383_c37 bl[37] br[37] wl[383] vdd gnd cell_6t
Xbit_r384_c37 bl[37] br[37] wl[384] vdd gnd cell_6t
Xbit_r385_c37 bl[37] br[37] wl[385] vdd gnd cell_6t
Xbit_r386_c37 bl[37] br[37] wl[386] vdd gnd cell_6t
Xbit_r387_c37 bl[37] br[37] wl[387] vdd gnd cell_6t
Xbit_r388_c37 bl[37] br[37] wl[388] vdd gnd cell_6t
Xbit_r389_c37 bl[37] br[37] wl[389] vdd gnd cell_6t
Xbit_r390_c37 bl[37] br[37] wl[390] vdd gnd cell_6t
Xbit_r391_c37 bl[37] br[37] wl[391] vdd gnd cell_6t
Xbit_r392_c37 bl[37] br[37] wl[392] vdd gnd cell_6t
Xbit_r393_c37 bl[37] br[37] wl[393] vdd gnd cell_6t
Xbit_r394_c37 bl[37] br[37] wl[394] vdd gnd cell_6t
Xbit_r395_c37 bl[37] br[37] wl[395] vdd gnd cell_6t
Xbit_r396_c37 bl[37] br[37] wl[396] vdd gnd cell_6t
Xbit_r397_c37 bl[37] br[37] wl[397] vdd gnd cell_6t
Xbit_r398_c37 bl[37] br[37] wl[398] vdd gnd cell_6t
Xbit_r399_c37 bl[37] br[37] wl[399] vdd gnd cell_6t
Xbit_r400_c37 bl[37] br[37] wl[400] vdd gnd cell_6t
Xbit_r401_c37 bl[37] br[37] wl[401] vdd gnd cell_6t
Xbit_r402_c37 bl[37] br[37] wl[402] vdd gnd cell_6t
Xbit_r403_c37 bl[37] br[37] wl[403] vdd gnd cell_6t
Xbit_r404_c37 bl[37] br[37] wl[404] vdd gnd cell_6t
Xbit_r405_c37 bl[37] br[37] wl[405] vdd gnd cell_6t
Xbit_r406_c37 bl[37] br[37] wl[406] vdd gnd cell_6t
Xbit_r407_c37 bl[37] br[37] wl[407] vdd gnd cell_6t
Xbit_r408_c37 bl[37] br[37] wl[408] vdd gnd cell_6t
Xbit_r409_c37 bl[37] br[37] wl[409] vdd gnd cell_6t
Xbit_r410_c37 bl[37] br[37] wl[410] vdd gnd cell_6t
Xbit_r411_c37 bl[37] br[37] wl[411] vdd gnd cell_6t
Xbit_r412_c37 bl[37] br[37] wl[412] vdd gnd cell_6t
Xbit_r413_c37 bl[37] br[37] wl[413] vdd gnd cell_6t
Xbit_r414_c37 bl[37] br[37] wl[414] vdd gnd cell_6t
Xbit_r415_c37 bl[37] br[37] wl[415] vdd gnd cell_6t
Xbit_r416_c37 bl[37] br[37] wl[416] vdd gnd cell_6t
Xbit_r417_c37 bl[37] br[37] wl[417] vdd gnd cell_6t
Xbit_r418_c37 bl[37] br[37] wl[418] vdd gnd cell_6t
Xbit_r419_c37 bl[37] br[37] wl[419] vdd gnd cell_6t
Xbit_r420_c37 bl[37] br[37] wl[420] vdd gnd cell_6t
Xbit_r421_c37 bl[37] br[37] wl[421] vdd gnd cell_6t
Xbit_r422_c37 bl[37] br[37] wl[422] vdd gnd cell_6t
Xbit_r423_c37 bl[37] br[37] wl[423] vdd gnd cell_6t
Xbit_r424_c37 bl[37] br[37] wl[424] vdd gnd cell_6t
Xbit_r425_c37 bl[37] br[37] wl[425] vdd gnd cell_6t
Xbit_r426_c37 bl[37] br[37] wl[426] vdd gnd cell_6t
Xbit_r427_c37 bl[37] br[37] wl[427] vdd gnd cell_6t
Xbit_r428_c37 bl[37] br[37] wl[428] vdd gnd cell_6t
Xbit_r429_c37 bl[37] br[37] wl[429] vdd gnd cell_6t
Xbit_r430_c37 bl[37] br[37] wl[430] vdd gnd cell_6t
Xbit_r431_c37 bl[37] br[37] wl[431] vdd gnd cell_6t
Xbit_r432_c37 bl[37] br[37] wl[432] vdd gnd cell_6t
Xbit_r433_c37 bl[37] br[37] wl[433] vdd gnd cell_6t
Xbit_r434_c37 bl[37] br[37] wl[434] vdd gnd cell_6t
Xbit_r435_c37 bl[37] br[37] wl[435] vdd gnd cell_6t
Xbit_r436_c37 bl[37] br[37] wl[436] vdd gnd cell_6t
Xbit_r437_c37 bl[37] br[37] wl[437] vdd gnd cell_6t
Xbit_r438_c37 bl[37] br[37] wl[438] vdd gnd cell_6t
Xbit_r439_c37 bl[37] br[37] wl[439] vdd gnd cell_6t
Xbit_r440_c37 bl[37] br[37] wl[440] vdd gnd cell_6t
Xbit_r441_c37 bl[37] br[37] wl[441] vdd gnd cell_6t
Xbit_r442_c37 bl[37] br[37] wl[442] vdd gnd cell_6t
Xbit_r443_c37 bl[37] br[37] wl[443] vdd gnd cell_6t
Xbit_r444_c37 bl[37] br[37] wl[444] vdd gnd cell_6t
Xbit_r445_c37 bl[37] br[37] wl[445] vdd gnd cell_6t
Xbit_r446_c37 bl[37] br[37] wl[446] vdd gnd cell_6t
Xbit_r447_c37 bl[37] br[37] wl[447] vdd gnd cell_6t
Xbit_r448_c37 bl[37] br[37] wl[448] vdd gnd cell_6t
Xbit_r449_c37 bl[37] br[37] wl[449] vdd gnd cell_6t
Xbit_r450_c37 bl[37] br[37] wl[450] vdd gnd cell_6t
Xbit_r451_c37 bl[37] br[37] wl[451] vdd gnd cell_6t
Xbit_r452_c37 bl[37] br[37] wl[452] vdd gnd cell_6t
Xbit_r453_c37 bl[37] br[37] wl[453] vdd gnd cell_6t
Xbit_r454_c37 bl[37] br[37] wl[454] vdd gnd cell_6t
Xbit_r455_c37 bl[37] br[37] wl[455] vdd gnd cell_6t
Xbit_r456_c37 bl[37] br[37] wl[456] vdd gnd cell_6t
Xbit_r457_c37 bl[37] br[37] wl[457] vdd gnd cell_6t
Xbit_r458_c37 bl[37] br[37] wl[458] vdd gnd cell_6t
Xbit_r459_c37 bl[37] br[37] wl[459] vdd gnd cell_6t
Xbit_r460_c37 bl[37] br[37] wl[460] vdd gnd cell_6t
Xbit_r461_c37 bl[37] br[37] wl[461] vdd gnd cell_6t
Xbit_r462_c37 bl[37] br[37] wl[462] vdd gnd cell_6t
Xbit_r463_c37 bl[37] br[37] wl[463] vdd gnd cell_6t
Xbit_r464_c37 bl[37] br[37] wl[464] vdd gnd cell_6t
Xbit_r465_c37 bl[37] br[37] wl[465] vdd gnd cell_6t
Xbit_r466_c37 bl[37] br[37] wl[466] vdd gnd cell_6t
Xbit_r467_c37 bl[37] br[37] wl[467] vdd gnd cell_6t
Xbit_r468_c37 bl[37] br[37] wl[468] vdd gnd cell_6t
Xbit_r469_c37 bl[37] br[37] wl[469] vdd gnd cell_6t
Xbit_r470_c37 bl[37] br[37] wl[470] vdd gnd cell_6t
Xbit_r471_c37 bl[37] br[37] wl[471] vdd gnd cell_6t
Xbit_r472_c37 bl[37] br[37] wl[472] vdd gnd cell_6t
Xbit_r473_c37 bl[37] br[37] wl[473] vdd gnd cell_6t
Xbit_r474_c37 bl[37] br[37] wl[474] vdd gnd cell_6t
Xbit_r475_c37 bl[37] br[37] wl[475] vdd gnd cell_6t
Xbit_r476_c37 bl[37] br[37] wl[476] vdd gnd cell_6t
Xbit_r477_c37 bl[37] br[37] wl[477] vdd gnd cell_6t
Xbit_r478_c37 bl[37] br[37] wl[478] vdd gnd cell_6t
Xbit_r479_c37 bl[37] br[37] wl[479] vdd gnd cell_6t
Xbit_r480_c37 bl[37] br[37] wl[480] vdd gnd cell_6t
Xbit_r481_c37 bl[37] br[37] wl[481] vdd gnd cell_6t
Xbit_r482_c37 bl[37] br[37] wl[482] vdd gnd cell_6t
Xbit_r483_c37 bl[37] br[37] wl[483] vdd gnd cell_6t
Xbit_r484_c37 bl[37] br[37] wl[484] vdd gnd cell_6t
Xbit_r485_c37 bl[37] br[37] wl[485] vdd gnd cell_6t
Xbit_r486_c37 bl[37] br[37] wl[486] vdd gnd cell_6t
Xbit_r487_c37 bl[37] br[37] wl[487] vdd gnd cell_6t
Xbit_r488_c37 bl[37] br[37] wl[488] vdd gnd cell_6t
Xbit_r489_c37 bl[37] br[37] wl[489] vdd gnd cell_6t
Xbit_r490_c37 bl[37] br[37] wl[490] vdd gnd cell_6t
Xbit_r491_c37 bl[37] br[37] wl[491] vdd gnd cell_6t
Xbit_r492_c37 bl[37] br[37] wl[492] vdd gnd cell_6t
Xbit_r493_c37 bl[37] br[37] wl[493] vdd gnd cell_6t
Xbit_r494_c37 bl[37] br[37] wl[494] vdd gnd cell_6t
Xbit_r495_c37 bl[37] br[37] wl[495] vdd gnd cell_6t
Xbit_r496_c37 bl[37] br[37] wl[496] vdd gnd cell_6t
Xbit_r497_c37 bl[37] br[37] wl[497] vdd gnd cell_6t
Xbit_r498_c37 bl[37] br[37] wl[498] vdd gnd cell_6t
Xbit_r499_c37 bl[37] br[37] wl[499] vdd gnd cell_6t
Xbit_r500_c37 bl[37] br[37] wl[500] vdd gnd cell_6t
Xbit_r501_c37 bl[37] br[37] wl[501] vdd gnd cell_6t
Xbit_r502_c37 bl[37] br[37] wl[502] vdd gnd cell_6t
Xbit_r503_c37 bl[37] br[37] wl[503] vdd gnd cell_6t
Xbit_r504_c37 bl[37] br[37] wl[504] vdd gnd cell_6t
Xbit_r505_c37 bl[37] br[37] wl[505] vdd gnd cell_6t
Xbit_r506_c37 bl[37] br[37] wl[506] vdd gnd cell_6t
Xbit_r507_c37 bl[37] br[37] wl[507] vdd gnd cell_6t
Xbit_r508_c37 bl[37] br[37] wl[508] vdd gnd cell_6t
Xbit_r509_c37 bl[37] br[37] wl[509] vdd gnd cell_6t
Xbit_r510_c37 bl[37] br[37] wl[510] vdd gnd cell_6t
Xbit_r511_c37 bl[37] br[37] wl[511] vdd gnd cell_6t
Xbit_r0_c38 bl[38] br[38] wl[0] vdd gnd cell_6t
Xbit_r1_c38 bl[38] br[38] wl[1] vdd gnd cell_6t
Xbit_r2_c38 bl[38] br[38] wl[2] vdd gnd cell_6t
Xbit_r3_c38 bl[38] br[38] wl[3] vdd gnd cell_6t
Xbit_r4_c38 bl[38] br[38] wl[4] vdd gnd cell_6t
Xbit_r5_c38 bl[38] br[38] wl[5] vdd gnd cell_6t
Xbit_r6_c38 bl[38] br[38] wl[6] vdd gnd cell_6t
Xbit_r7_c38 bl[38] br[38] wl[7] vdd gnd cell_6t
Xbit_r8_c38 bl[38] br[38] wl[8] vdd gnd cell_6t
Xbit_r9_c38 bl[38] br[38] wl[9] vdd gnd cell_6t
Xbit_r10_c38 bl[38] br[38] wl[10] vdd gnd cell_6t
Xbit_r11_c38 bl[38] br[38] wl[11] vdd gnd cell_6t
Xbit_r12_c38 bl[38] br[38] wl[12] vdd gnd cell_6t
Xbit_r13_c38 bl[38] br[38] wl[13] vdd gnd cell_6t
Xbit_r14_c38 bl[38] br[38] wl[14] vdd gnd cell_6t
Xbit_r15_c38 bl[38] br[38] wl[15] vdd gnd cell_6t
Xbit_r16_c38 bl[38] br[38] wl[16] vdd gnd cell_6t
Xbit_r17_c38 bl[38] br[38] wl[17] vdd gnd cell_6t
Xbit_r18_c38 bl[38] br[38] wl[18] vdd gnd cell_6t
Xbit_r19_c38 bl[38] br[38] wl[19] vdd gnd cell_6t
Xbit_r20_c38 bl[38] br[38] wl[20] vdd gnd cell_6t
Xbit_r21_c38 bl[38] br[38] wl[21] vdd gnd cell_6t
Xbit_r22_c38 bl[38] br[38] wl[22] vdd gnd cell_6t
Xbit_r23_c38 bl[38] br[38] wl[23] vdd gnd cell_6t
Xbit_r24_c38 bl[38] br[38] wl[24] vdd gnd cell_6t
Xbit_r25_c38 bl[38] br[38] wl[25] vdd gnd cell_6t
Xbit_r26_c38 bl[38] br[38] wl[26] vdd gnd cell_6t
Xbit_r27_c38 bl[38] br[38] wl[27] vdd gnd cell_6t
Xbit_r28_c38 bl[38] br[38] wl[28] vdd gnd cell_6t
Xbit_r29_c38 bl[38] br[38] wl[29] vdd gnd cell_6t
Xbit_r30_c38 bl[38] br[38] wl[30] vdd gnd cell_6t
Xbit_r31_c38 bl[38] br[38] wl[31] vdd gnd cell_6t
Xbit_r32_c38 bl[38] br[38] wl[32] vdd gnd cell_6t
Xbit_r33_c38 bl[38] br[38] wl[33] vdd gnd cell_6t
Xbit_r34_c38 bl[38] br[38] wl[34] vdd gnd cell_6t
Xbit_r35_c38 bl[38] br[38] wl[35] vdd gnd cell_6t
Xbit_r36_c38 bl[38] br[38] wl[36] vdd gnd cell_6t
Xbit_r37_c38 bl[38] br[38] wl[37] vdd gnd cell_6t
Xbit_r38_c38 bl[38] br[38] wl[38] vdd gnd cell_6t
Xbit_r39_c38 bl[38] br[38] wl[39] vdd gnd cell_6t
Xbit_r40_c38 bl[38] br[38] wl[40] vdd gnd cell_6t
Xbit_r41_c38 bl[38] br[38] wl[41] vdd gnd cell_6t
Xbit_r42_c38 bl[38] br[38] wl[42] vdd gnd cell_6t
Xbit_r43_c38 bl[38] br[38] wl[43] vdd gnd cell_6t
Xbit_r44_c38 bl[38] br[38] wl[44] vdd gnd cell_6t
Xbit_r45_c38 bl[38] br[38] wl[45] vdd gnd cell_6t
Xbit_r46_c38 bl[38] br[38] wl[46] vdd gnd cell_6t
Xbit_r47_c38 bl[38] br[38] wl[47] vdd gnd cell_6t
Xbit_r48_c38 bl[38] br[38] wl[48] vdd gnd cell_6t
Xbit_r49_c38 bl[38] br[38] wl[49] vdd gnd cell_6t
Xbit_r50_c38 bl[38] br[38] wl[50] vdd gnd cell_6t
Xbit_r51_c38 bl[38] br[38] wl[51] vdd gnd cell_6t
Xbit_r52_c38 bl[38] br[38] wl[52] vdd gnd cell_6t
Xbit_r53_c38 bl[38] br[38] wl[53] vdd gnd cell_6t
Xbit_r54_c38 bl[38] br[38] wl[54] vdd gnd cell_6t
Xbit_r55_c38 bl[38] br[38] wl[55] vdd gnd cell_6t
Xbit_r56_c38 bl[38] br[38] wl[56] vdd gnd cell_6t
Xbit_r57_c38 bl[38] br[38] wl[57] vdd gnd cell_6t
Xbit_r58_c38 bl[38] br[38] wl[58] vdd gnd cell_6t
Xbit_r59_c38 bl[38] br[38] wl[59] vdd gnd cell_6t
Xbit_r60_c38 bl[38] br[38] wl[60] vdd gnd cell_6t
Xbit_r61_c38 bl[38] br[38] wl[61] vdd gnd cell_6t
Xbit_r62_c38 bl[38] br[38] wl[62] vdd gnd cell_6t
Xbit_r63_c38 bl[38] br[38] wl[63] vdd gnd cell_6t
Xbit_r64_c38 bl[38] br[38] wl[64] vdd gnd cell_6t
Xbit_r65_c38 bl[38] br[38] wl[65] vdd gnd cell_6t
Xbit_r66_c38 bl[38] br[38] wl[66] vdd gnd cell_6t
Xbit_r67_c38 bl[38] br[38] wl[67] vdd gnd cell_6t
Xbit_r68_c38 bl[38] br[38] wl[68] vdd gnd cell_6t
Xbit_r69_c38 bl[38] br[38] wl[69] vdd gnd cell_6t
Xbit_r70_c38 bl[38] br[38] wl[70] vdd gnd cell_6t
Xbit_r71_c38 bl[38] br[38] wl[71] vdd gnd cell_6t
Xbit_r72_c38 bl[38] br[38] wl[72] vdd gnd cell_6t
Xbit_r73_c38 bl[38] br[38] wl[73] vdd gnd cell_6t
Xbit_r74_c38 bl[38] br[38] wl[74] vdd gnd cell_6t
Xbit_r75_c38 bl[38] br[38] wl[75] vdd gnd cell_6t
Xbit_r76_c38 bl[38] br[38] wl[76] vdd gnd cell_6t
Xbit_r77_c38 bl[38] br[38] wl[77] vdd gnd cell_6t
Xbit_r78_c38 bl[38] br[38] wl[78] vdd gnd cell_6t
Xbit_r79_c38 bl[38] br[38] wl[79] vdd gnd cell_6t
Xbit_r80_c38 bl[38] br[38] wl[80] vdd gnd cell_6t
Xbit_r81_c38 bl[38] br[38] wl[81] vdd gnd cell_6t
Xbit_r82_c38 bl[38] br[38] wl[82] vdd gnd cell_6t
Xbit_r83_c38 bl[38] br[38] wl[83] vdd gnd cell_6t
Xbit_r84_c38 bl[38] br[38] wl[84] vdd gnd cell_6t
Xbit_r85_c38 bl[38] br[38] wl[85] vdd gnd cell_6t
Xbit_r86_c38 bl[38] br[38] wl[86] vdd gnd cell_6t
Xbit_r87_c38 bl[38] br[38] wl[87] vdd gnd cell_6t
Xbit_r88_c38 bl[38] br[38] wl[88] vdd gnd cell_6t
Xbit_r89_c38 bl[38] br[38] wl[89] vdd gnd cell_6t
Xbit_r90_c38 bl[38] br[38] wl[90] vdd gnd cell_6t
Xbit_r91_c38 bl[38] br[38] wl[91] vdd gnd cell_6t
Xbit_r92_c38 bl[38] br[38] wl[92] vdd gnd cell_6t
Xbit_r93_c38 bl[38] br[38] wl[93] vdd gnd cell_6t
Xbit_r94_c38 bl[38] br[38] wl[94] vdd gnd cell_6t
Xbit_r95_c38 bl[38] br[38] wl[95] vdd gnd cell_6t
Xbit_r96_c38 bl[38] br[38] wl[96] vdd gnd cell_6t
Xbit_r97_c38 bl[38] br[38] wl[97] vdd gnd cell_6t
Xbit_r98_c38 bl[38] br[38] wl[98] vdd gnd cell_6t
Xbit_r99_c38 bl[38] br[38] wl[99] vdd gnd cell_6t
Xbit_r100_c38 bl[38] br[38] wl[100] vdd gnd cell_6t
Xbit_r101_c38 bl[38] br[38] wl[101] vdd gnd cell_6t
Xbit_r102_c38 bl[38] br[38] wl[102] vdd gnd cell_6t
Xbit_r103_c38 bl[38] br[38] wl[103] vdd gnd cell_6t
Xbit_r104_c38 bl[38] br[38] wl[104] vdd gnd cell_6t
Xbit_r105_c38 bl[38] br[38] wl[105] vdd gnd cell_6t
Xbit_r106_c38 bl[38] br[38] wl[106] vdd gnd cell_6t
Xbit_r107_c38 bl[38] br[38] wl[107] vdd gnd cell_6t
Xbit_r108_c38 bl[38] br[38] wl[108] vdd gnd cell_6t
Xbit_r109_c38 bl[38] br[38] wl[109] vdd gnd cell_6t
Xbit_r110_c38 bl[38] br[38] wl[110] vdd gnd cell_6t
Xbit_r111_c38 bl[38] br[38] wl[111] vdd gnd cell_6t
Xbit_r112_c38 bl[38] br[38] wl[112] vdd gnd cell_6t
Xbit_r113_c38 bl[38] br[38] wl[113] vdd gnd cell_6t
Xbit_r114_c38 bl[38] br[38] wl[114] vdd gnd cell_6t
Xbit_r115_c38 bl[38] br[38] wl[115] vdd gnd cell_6t
Xbit_r116_c38 bl[38] br[38] wl[116] vdd gnd cell_6t
Xbit_r117_c38 bl[38] br[38] wl[117] vdd gnd cell_6t
Xbit_r118_c38 bl[38] br[38] wl[118] vdd gnd cell_6t
Xbit_r119_c38 bl[38] br[38] wl[119] vdd gnd cell_6t
Xbit_r120_c38 bl[38] br[38] wl[120] vdd gnd cell_6t
Xbit_r121_c38 bl[38] br[38] wl[121] vdd gnd cell_6t
Xbit_r122_c38 bl[38] br[38] wl[122] vdd gnd cell_6t
Xbit_r123_c38 bl[38] br[38] wl[123] vdd gnd cell_6t
Xbit_r124_c38 bl[38] br[38] wl[124] vdd gnd cell_6t
Xbit_r125_c38 bl[38] br[38] wl[125] vdd gnd cell_6t
Xbit_r126_c38 bl[38] br[38] wl[126] vdd gnd cell_6t
Xbit_r127_c38 bl[38] br[38] wl[127] vdd gnd cell_6t
Xbit_r128_c38 bl[38] br[38] wl[128] vdd gnd cell_6t
Xbit_r129_c38 bl[38] br[38] wl[129] vdd gnd cell_6t
Xbit_r130_c38 bl[38] br[38] wl[130] vdd gnd cell_6t
Xbit_r131_c38 bl[38] br[38] wl[131] vdd gnd cell_6t
Xbit_r132_c38 bl[38] br[38] wl[132] vdd gnd cell_6t
Xbit_r133_c38 bl[38] br[38] wl[133] vdd gnd cell_6t
Xbit_r134_c38 bl[38] br[38] wl[134] vdd gnd cell_6t
Xbit_r135_c38 bl[38] br[38] wl[135] vdd gnd cell_6t
Xbit_r136_c38 bl[38] br[38] wl[136] vdd gnd cell_6t
Xbit_r137_c38 bl[38] br[38] wl[137] vdd gnd cell_6t
Xbit_r138_c38 bl[38] br[38] wl[138] vdd gnd cell_6t
Xbit_r139_c38 bl[38] br[38] wl[139] vdd gnd cell_6t
Xbit_r140_c38 bl[38] br[38] wl[140] vdd gnd cell_6t
Xbit_r141_c38 bl[38] br[38] wl[141] vdd gnd cell_6t
Xbit_r142_c38 bl[38] br[38] wl[142] vdd gnd cell_6t
Xbit_r143_c38 bl[38] br[38] wl[143] vdd gnd cell_6t
Xbit_r144_c38 bl[38] br[38] wl[144] vdd gnd cell_6t
Xbit_r145_c38 bl[38] br[38] wl[145] vdd gnd cell_6t
Xbit_r146_c38 bl[38] br[38] wl[146] vdd gnd cell_6t
Xbit_r147_c38 bl[38] br[38] wl[147] vdd gnd cell_6t
Xbit_r148_c38 bl[38] br[38] wl[148] vdd gnd cell_6t
Xbit_r149_c38 bl[38] br[38] wl[149] vdd gnd cell_6t
Xbit_r150_c38 bl[38] br[38] wl[150] vdd gnd cell_6t
Xbit_r151_c38 bl[38] br[38] wl[151] vdd gnd cell_6t
Xbit_r152_c38 bl[38] br[38] wl[152] vdd gnd cell_6t
Xbit_r153_c38 bl[38] br[38] wl[153] vdd gnd cell_6t
Xbit_r154_c38 bl[38] br[38] wl[154] vdd gnd cell_6t
Xbit_r155_c38 bl[38] br[38] wl[155] vdd gnd cell_6t
Xbit_r156_c38 bl[38] br[38] wl[156] vdd gnd cell_6t
Xbit_r157_c38 bl[38] br[38] wl[157] vdd gnd cell_6t
Xbit_r158_c38 bl[38] br[38] wl[158] vdd gnd cell_6t
Xbit_r159_c38 bl[38] br[38] wl[159] vdd gnd cell_6t
Xbit_r160_c38 bl[38] br[38] wl[160] vdd gnd cell_6t
Xbit_r161_c38 bl[38] br[38] wl[161] vdd gnd cell_6t
Xbit_r162_c38 bl[38] br[38] wl[162] vdd gnd cell_6t
Xbit_r163_c38 bl[38] br[38] wl[163] vdd gnd cell_6t
Xbit_r164_c38 bl[38] br[38] wl[164] vdd gnd cell_6t
Xbit_r165_c38 bl[38] br[38] wl[165] vdd gnd cell_6t
Xbit_r166_c38 bl[38] br[38] wl[166] vdd gnd cell_6t
Xbit_r167_c38 bl[38] br[38] wl[167] vdd gnd cell_6t
Xbit_r168_c38 bl[38] br[38] wl[168] vdd gnd cell_6t
Xbit_r169_c38 bl[38] br[38] wl[169] vdd gnd cell_6t
Xbit_r170_c38 bl[38] br[38] wl[170] vdd gnd cell_6t
Xbit_r171_c38 bl[38] br[38] wl[171] vdd gnd cell_6t
Xbit_r172_c38 bl[38] br[38] wl[172] vdd gnd cell_6t
Xbit_r173_c38 bl[38] br[38] wl[173] vdd gnd cell_6t
Xbit_r174_c38 bl[38] br[38] wl[174] vdd gnd cell_6t
Xbit_r175_c38 bl[38] br[38] wl[175] vdd gnd cell_6t
Xbit_r176_c38 bl[38] br[38] wl[176] vdd gnd cell_6t
Xbit_r177_c38 bl[38] br[38] wl[177] vdd gnd cell_6t
Xbit_r178_c38 bl[38] br[38] wl[178] vdd gnd cell_6t
Xbit_r179_c38 bl[38] br[38] wl[179] vdd gnd cell_6t
Xbit_r180_c38 bl[38] br[38] wl[180] vdd gnd cell_6t
Xbit_r181_c38 bl[38] br[38] wl[181] vdd gnd cell_6t
Xbit_r182_c38 bl[38] br[38] wl[182] vdd gnd cell_6t
Xbit_r183_c38 bl[38] br[38] wl[183] vdd gnd cell_6t
Xbit_r184_c38 bl[38] br[38] wl[184] vdd gnd cell_6t
Xbit_r185_c38 bl[38] br[38] wl[185] vdd gnd cell_6t
Xbit_r186_c38 bl[38] br[38] wl[186] vdd gnd cell_6t
Xbit_r187_c38 bl[38] br[38] wl[187] vdd gnd cell_6t
Xbit_r188_c38 bl[38] br[38] wl[188] vdd gnd cell_6t
Xbit_r189_c38 bl[38] br[38] wl[189] vdd gnd cell_6t
Xbit_r190_c38 bl[38] br[38] wl[190] vdd gnd cell_6t
Xbit_r191_c38 bl[38] br[38] wl[191] vdd gnd cell_6t
Xbit_r192_c38 bl[38] br[38] wl[192] vdd gnd cell_6t
Xbit_r193_c38 bl[38] br[38] wl[193] vdd gnd cell_6t
Xbit_r194_c38 bl[38] br[38] wl[194] vdd gnd cell_6t
Xbit_r195_c38 bl[38] br[38] wl[195] vdd gnd cell_6t
Xbit_r196_c38 bl[38] br[38] wl[196] vdd gnd cell_6t
Xbit_r197_c38 bl[38] br[38] wl[197] vdd gnd cell_6t
Xbit_r198_c38 bl[38] br[38] wl[198] vdd gnd cell_6t
Xbit_r199_c38 bl[38] br[38] wl[199] vdd gnd cell_6t
Xbit_r200_c38 bl[38] br[38] wl[200] vdd gnd cell_6t
Xbit_r201_c38 bl[38] br[38] wl[201] vdd gnd cell_6t
Xbit_r202_c38 bl[38] br[38] wl[202] vdd gnd cell_6t
Xbit_r203_c38 bl[38] br[38] wl[203] vdd gnd cell_6t
Xbit_r204_c38 bl[38] br[38] wl[204] vdd gnd cell_6t
Xbit_r205_c38 bl[38] br[38] wl[205] vdd gnd cell_6t
Xbit_r206_c38 bl[38] br[38] wl[206] vdd gnd cell_6t
Xbit_r207_c38 bl[38] br[38] wl[207] vdd gnd cell_6t
Xbit_r208_c38 bl[38] br[38] wl[208] vdd gnd cell_6t
Xbit_r209_c38 bl[38] br[38] wl[209] vdd gnd cell_6t
Xbit_r210_c38 bl[38] br[38] wl[210] vdd gnd cell_6t
Xbit_r211_c38 bl[38] br[38] wl[211] vdd gnd cell_6t
Xbit_r212_c38 bl[38] br[38] wl[212] vdd gnd cell_6t
Xbit_r213_c38 bl[38] br[38] wl[213] vdd gnd cell_6t
Xbit_r214_c38 bl[38] br[38] wl[214] vdd gnd cell_6t
Xbit_r215_c38 bl[38] br[38] wl[215] vdd gnd cell_6t
Xbit_r216_c38 bl[38] br[38] wl[216] vdd gnd cell_6t
Xbit_r217_c38 bl[38] br[38] wl[217] vdd gnd cell_6t
Xbit_r218_c38 bl[38] br[38] wl[218] vdd gnd cell_6t
Xbit_r219_c38 bl[38] br[38] wl[219] vdd gnd cell_6t
Xbit_r220_c38 bl[38] br[38] wl[220] vdd gnd cell_6t
Xbit_r221_c38 bl[38] br[38] wl[221] vdd gnd cell_6t
Xbit_r222_c38 bl[38] br[38] wl[222] vdd gnd cell_6t
Xbit_r223_c38 bl[38] br[38] wl[223] vdd gnd cell_6t
Xbit_r224_c38 bl[38] br[38] wl[224] vdd gnd cell_6t
Xbit_r225_c38 bl[38] br[38] wl[225] vdd gnd cell_6t
Xbit_r226_c38 bl[38] br[38] wl[226] vdd gnd cell_6t
Xbit_r227_c38 bl[38] br[38] wl[227] vdd gnd cell_6t
Xbit_r228_c38 bl[38] br[38] wl[228] vdd gnd cell_6t
Xbit_r229_c38 bl[38] br[38] wl[229] vdd gnd cell_6t
Xbit_r230_c38 bl[38] br[38] wl[230] vdd gnd cell_6t
Xbit_r231_c38 bl[38] br[38] wl[231] vdd gnd cell_6t
Xbit_r232_c38 bl[38] br[38] wl[232] vdd gnd cell_6t
Xbit_r233_c38 bl[38] br[38] wl[233] vdd gnd cell_6t
Xbit_r234_c38 bl[38] br[38] wl[234] vdd gnd cell_6t
Xbit_r235_c38 bl[38] br[38] wl[235] vdd gnd cell_6t
Xbit_r236_c38 bl[38] br[38] wl[236] vdd gnd cell_6t
Xbit_r237_c38 bl[38] br[38] wl[237] vdd gnd cell_6t
Xbit_r238_c38 bl[38] br[38] wl[238] vdd gnd cell_6t
Xbit_r239_c38 bl[38] br[38] wl[239] vdd gnd cell_6t
Xbit_r240_c38 bl[38] br[38] wl[240] vdd gnd cell_6t
Xbit_r241_c38 bl[38] br[38] wl[241] vdd gnd cell_6t
Xbit_r242_c38 bl[38] br[38] wl[242] vdd gnd cell_6t
Xbit_r243_c38 bl[38] br[38] wl[243] vdd gnd cell_6t
Xbit_r244_c38 bl[38] br[38] wl[244] vdd gnd cell_6t
Xbit_r245_c38 bl[38] br[38] wl[245] vdd gnd cell_6t
Xbit_r246_c38 bl[38] br[38] wl[246] vdd gnd cell_6t
Xbit_r247_c38 bl[38] br[38] wl[247] vdd gnd cell_6t
Xbit_r248_c38 bl[38] br[38] wl[248] vdd gnd cell_6t
Xbit_r249_c38 bl[38] br[38] wl[249] vdd gnd cell_6t
Xbit_r250_c38 bl[38] br[38] wl[250] vdd gnd cell_6t
Xbit_r251_c38 bl[38] br[38] wl[251] vdd gnd cell_6t
Xbit_r252_c38 bl[38] br[38] wl[252] vdd gnd cell_6t
Xbit_r253_c38 bl[38] br[38] wl[253] vdd gnd cell_6t
Xbit_r254_c38 bl[38] br[38] wl[254] vdd gnd cell_6t
Xbit_r255_c38 bl[38] br[38] wl[255] vdd gnd cell_6t
Xbit_r256_c38 bl[38] br[38] wl[256] vdd gnd cell_6t
Xbit_r257_c38 bl[38] br[38] wl[257] vdd gnd cell_6t
Xbit_r258_c38 bl[38] br[38] wl[258] vdd gnd cell_6t
Xbit_r259_c38 bl[38] br[38] wl[259] vdd gnd cell_6t
Xbit_r260_c38 bl[38] br[38] wl[260] vdd gnd cell_6t
Xbit_r261_c38 bl[38] br[38] wl[261] vdd gnd cell_6t
Xbit_r262_c38 bl[38] br[38] wl[262] vdd gnd cell_6t
Xbit_r263_c38 bl[38] br[38] wl[263] vdd gnd cell_6t
Xbit_r264_c38 bl[38] br[38] wl[264] vdd gnd cell_6t
Xbit_r265_c38 bl[38] br[38] wl[265] vdd gnd cell_6t
Xbit_r266_c38 bl[38] br[38] wl[266] vdd gnd cell_6t
Xbit_r267_c38 bl[38] br[38] wl[267] vdd gnd cell_6t
Xbit_r268_c38 bl[38] br[38] wl[268] vdd gnd cell_6t
Xbit_r269_c38 bl[38] br[38] wl[269] vdd gnd cell_6t
Xbit_r270_c38 bl[38] br[38] wl[270] vdd gnd cell_6t
Xbit_r271_c38 bl[38] br[38] wl[271] vdd gnd cell_6t
Xbit_r272_c38 bl[38] br[38] wl[272] vdd gnd cell_6t
Xbit_r273_c38 bl[38] br[38] wl[273] vdd gnd cell_6t
Xbit_r274_c38 bl[38] br[38] wl[274] vdd gnd cell_6t
Xbit_r275_c38 bl[38] br[38] wl[275] vdd gnd cell_6t
Xbit_r276_c38 bl[38] br[38] wl[276] vdd gnd cell_6t
Xbit_r277_c38 bl[38] br[38] wl[277] vdd gnd cell_6t
Xbit_r278_c38 bl[38] br[38] wl[278] vdd gnd cell_6t
Xbit_r279_c38 bl[38] br[38] wl[279] vdd gnd cell_6t
Xbit_r280_c38 bl[38] br[38] wl[280] vdd gnd cell_6t
Xbit_r281_c38 bl[38] br[38] wl[281] vdd gnd cell_6t
Xbit_r282_c38 bl[38] br[38] wl[282] vdd gnd cell_6t
Xbit_r283_c38 bl[38] br[38] wl[283] vdd gnd cell_6t
Xbit_r284_c38 bl[38] br[38] wl[284] vdd gnd cell_6t
Xbit_r285_c38 bl[38] br[38] wl[285] vdd gnd cell_6t
Xbit_r286_c38 bl[38] br[38] wl[286] vdd gnd cell_6t
Xbit_r287_c38 bl[38] br[38] wl[287] vdd gnd cell_6t
Xbit_r288_c38 bl[38] br[38] wl[288] vdd gnd cell_6t
Xbit_r289_c38 bl[38] br[38] wl[289] vdd gnd cell_6t
Xbit_r290_c38 bl[38] br[38] wl[290] vdd gnd cell_6t
Xbit_r291_c38 bl[38] br[38] wl[291] vdd gnd cell_6t
Xbit_r292_c38 bl[38] br[38] wl[292] vdd gnd cell_6t
Xbit_r293_c38 bl[38] br[38] wl[293] vdd gnd cell_6t
Xbit_r294_c38 bl[38] br[38] wl[294] vdd gnd cell_6t
Xbit_r295_c38 bl[38] br[38] wl[295] vdd gnd cell_6t
Xbit_r296_c38 bl[38] br[38] wl[296] vdd gnd cell_6t
Xbit_r297_c38 bl[38] br[38] wl[297] vdd gnd cell_6t
Xbit_r298_c38 bl[38] br[38] wl[298] vdd gnd cell_6t
Xbit_r299_c38 bl[38] br[38] wl[299] vdd gnd cell_6t
Xbit_r300_c38 bl[38] br[38] wl[300] vdd gnd cell_6t
Xbit_r301_c38 bl[38] br[38] wl[301] vdd gnd cell_6t
Xbit_r302_c38 bl[38] br[38] wl[302] vdd gnd cell_6t
Xbit_r303_c38 bl[38] br[38] wl[303] vdd gnd cell_6t
Xbit_r304_c38 bl[38] br[38] wl[304] vdd gnd cell_6t
Xbit_r305_c38 bl[38] br[38] wl[305] vdd gnd cell_6t
Xbit_r306_c38 bl[38] br[38] wl[306] vdd gnd cell_6t
Xbit_r307_c38 bl[38] br[38] wl[307] vdd gnd cell_6t
Xbit_r308_c38 bl[38] br[38] wl[308] vdd gnd cell_6t
Xbit_r309_c38 bl[38] br[38] wl[309] vdd gnd cell_6t
Xbit_r310_c38 bl[38] br[38] wl[310] vdd gnd cell_6t
Xbit_r311_c38 bl[38] br[38] wl[311] vdd gnd cell_6t
Xbit_r312_c38 bl[38] br[38] wl[312] vdd gnd cell_6t
Xbit_r313_c38 bl[38] br[38] wl[313] vdd gnd cell_6t
Xbit_r314_c38 bl[38] br[38] wl[314] vdd gnd cell_6t
Xbit_r315_c38 bl[38] br[38] wl[315] vdd gnd cell_6t
Xbit_r316_c38 bl[38] br[38] wl[316] vdd gnd cell_6t
Xbit_r317_c38 bl[38] br[38] wl[317] vdd gnd cell_6t
Xbit_r318_c38 bl[38] br[38] wl[318] vdd gnd cell_6t
Xbit_r319_c38 bl[38] br[38] wl[319] vdd gnd cell_6t
Xbit_r320_c38 bl[38] br[38] wl[320] vdd gnd cell_6t
Xbit_r321_c38 bl[38] br[38] wl[321] vdd gnd cell_6t
Xbit_r322_c38 bl[38] br[38] wl[322] vdd gnd cell_6t
Xbit_r323_c38 bl[38] br[38] wl[323] vdd gnd cell_6t
Xbit_r324_c38 bl[38] br[38] wl[324] vdd gnd cell_6t
Xbit_r325_c38 bl[38] br[38] wl[325] vdd gnd cell_6t
Xbit_r326_c38 bl[38] br[38] wl[326] vdd gnd cell_6t
Xbit_r327_c38 bl[38] br[38] wl[327] vdd gnd cell_6t
Xbit_r328_c38 bl[38] br[38] wl[328] vdd gnd cell_6t
Xbit_r329_c38 bl[38] br[38] wl[329] vdd gnd cell_6t
Xbit_r330_c38 bl[38] br[38] wl[330] vdd gnd cell_6t
Xbit_r331_c38 bl[38] br[38] wl[331] vdd gnd cell_6t
Xbit_r332_c38 bl[38] br[38] wl[332] vdd gnd cell_6t
Xbit_r333_c38 bl[38] br[38] wl[333] vdd gnd cell_6t
Xbit_r334_c38 bl[38] br[38] wl[334] vdd gnd cell_6t
Xbit_r335_c38 bl[38] br[38] wl[335] vdd gnd cell_6t
Xbit_r336_c38 bl[38] br[38] wl[336] vdd gnd cell_6t
Xbit_r337_c38 bl[38] br[38] wl[337] vdd gnd cell_6t
Xbit_r338_c38 bl[38] br[38] wl[338] vdd gnd cell_6t
Xbit_r339_c38 bl[38] br[38] wl[339] vdd gnd cell_6t
Xbit_r340_c38 bl[38] br[38] wl[340] vdd gnd cell_6t
Xbit_r341_c38 bl[38] br[38] wl[341] vdd gnd cell_6t
Xbit_r342_c38 bl[38] br[38] wl[342] vdd gnd cell_6t
Xbit_r343_c38 bl[38] br[38] wl[343] vdd gnd cell_6t
Xbit_r344_c38 bl[38] br[38] wl[344] vdd gnd cell_6t
Xbit_r345_c38 bl[38] br[38] wl[345] vdd gnd cell_6t
Xbit_r346_c38 bl[38] br[38] wl[346] vdd gnd cell_6t
Xbit_r347_c38 bl[38] br[38] wl[347] vdd gnd cell_6t
Xbit_r348_c38 bl[38] br[38] wl[348] vdd gnd cell_6t
Xbit_r349_c38 bl[38] br[38] wl[349] vdd gnd cell_6t
Xbit_r350_c38 bl[38] br[38] wl[350] vdd gnd cell_6t
Xbit_r351_c38 bl[38] br[38] wl[351] vdd gnd cell_6t
Xbit_r352_c38 bl[38] br[38] wl[352] vdd gnd cell_6t
Xbit_r353_c38 bl[38] br[38] wl[353] vdd gnd cell_6t
Xbit_r354_c38 bl[38] br[38] wl[354] vdd gnd cell_6t
Xbit_r355_c38 bl[38] br[38] wl[355] vdd gnd cell_6t
Xbit_r356_c38 bl[38] br[38] wl[356] vdd gnd cell_6t
Xbit_r357_c38 bl[38] br[38] wl[357] vdd gnd cell_6t
Xbit_r358_c38 bl[38] br[38] wl[358] vdd gnd cell_6t
Xbit_r359_c38 bl[38] br[38] wl[359] vdd gnd cell_6t
Xbit_r360_c38 bl[38] br[38] wl[360] vdd gnd cell_6t
Xbit_r361_c38 bl[38] br[38] wl[361] vdd gnd cell_6t
Xbit_r362_c38 bl[38] br[38] wl[362] vdd gnd cell_6t
Xbit_r363_c38 bl[38] br[38] wl[363] vdd gnd cell_6t
Xbit_r364_c38 bl[38] br[38] wl[364] vdd gnd cell_6t
Xbit_r365_c38 bl[38] br[38] wl[365] vdd gnd cell_6t
Xbit_r366_c38 bl[38] br[38] wl[366] vdd gnd cell_6t
Xbit_r367_c38 bl[38] br[38] wl[367] vdd gnd cell_6t
Xbit_r368_c38 bl[38] br[38] wl[368] vdd gnd cell_6t
Xbit_r369_c38 bl[38] br[38] wl[369] vdd gnd cell_6t
Xbit_r370_c38 bl[38] br[38] wl[370] vdd gnd cell_6t
Xbit_r371_c38 bl[38] br[38] wl[371] vdd gnd cell_6t
Xbit_r372_c38 bl[38] br[38] wl[372] vdd gnd cell_6t
Xbit_r373_c38 bl[38] br[38] wl[373] vdd gnd cell_6t
Xbit_r374_c38 bl[38] br[38] wl[374] vdd gnd cell_6t
Xbit_r375_c38 bl[38] br[38] wl[375] vdd gnd cell_6t
Xbit_r376_c38 bl[38] br[38] wl[376] vdd gnd cell_6t
Xbit_r377_c38 bl[38] br[38] wl[377] vdd gnd cell_6t
Xbit_r378_c38 bl[38] br[38] wl[378] vdd gnd cell_6t
Xbit_r379_c38 bl[38] br[38] wl[379] vdd gnd cell_6t
Xbit_r380_c38 bl[38] br[38] wl[380] vdd gnd cell_6t
Xbit_r381_c38 bl[38] br[38] wl[381] vdd gnd cell_6t
Xbit_r382_c38 bl[38] br[38] wl[382] vdd gnd cell_6t
Xbit_r383_c38 bl[38] br[38] wl[383] vdd gnd cell_6t
Xbit_r384_c38 bl[38] br[38] wl[384] vdd gnd cell_6t
Xbit_r385_c38 bl[38] br[38] wl[385] vdd gnd cell_6t
Xbit_r386_c38 bl[38] br[38] wl[386] vdd gnd cell_6t
Xbit_r387_c38 bl[38] br[38] wl[387] vdd gnd cell_6t
Xbit_r388_c38 bl[38] br[38] wl[388] vdd gnd cell_6t
Xbit_r389_c38 bl[38] br[38] wl[389] vdd gnd cell_6t
Xbit_r390_c38 bl[38] br[38] wl[390] vdd gnd cell_6t
Xbit_r391_c38 bl[38] br[38] wl[391] vdd gnd cell_6t
Xbit_r392_c38 bl[38] br[38] wl[392] vdd gnd cell_6t
Xbit_r393_c38 bl[38] br[38] wl[393] vdd gnd cell_6t
Xbit_r394_c38 bl[38] br[38] wl[394] vdd gnd cell_6t
Xbit_r395_c38 bl[38] br[38] wl[395] vdd gnd cell_6t
Xbit_r396_c38 bl[38] br[38] wl[396] vdd gnd cell_6t
Xbit_r397_c38 bl[38] br[38] wl[397] vdd gnd cell_6t
Xbit_r398_c38 bl[38] br[38] wl[398] vdd gnd cell_6t
Xbit_r399_c38 bl[38] br[38] wl[399] vdd gnd cell_6t
Xbit_r400_c38 bl[38] br[38] wl[400] vdd gnd cell_6t
Xbit_r401_c38 bl[38] br[38] wl[401] vdd gnd cell_6t
Xbit_r402_c38 bl[38] br[38] wl[402] vdd gnd cell_6t
Xbit_r403_c38 bl[38] br[38] wl[403] vdd gnd cell_6t
Xbit_r404_c38 bl[38] br[38] wl[404] vdd gnd cell_6t
Xbit_r405_c38 bl[38] br[38] wl[405] vdd gnd cell_6t
Xbit_r406_c38 bl[38] br[38] wl[406] vdd gnd cell_6t
Xbit_r407_c38 bl[38] br[38] wl[407] vdd gnd cell_6t
Xbit_r408_c38 bl[38] br[38] wl[408] vdd gnd cell_6t
Xbit_r409_c38 bl[38] br[38] wl[409] vdd gnd cell_6t
Xbit_r410_c38 bl[38] br[38] wl[410] vdd gnd cell_6t
Xbit_r411_c38 bl[38] br[38] wl[411] vdd gnd cell_6t
Xbit_r412_c38 bl[38] br[38] wl[412] vdd gnd cell_6t
Xbit_r413_c38 bl[38] br[38] wl[413] vdd gnd cell_6t
Xbit_r414_c38 bl[38] br[38] wl[414] vdd gnd cell_6t
Xbit_r415_c38 bl[38] br[38] wl[415] vdd gnd cell_6t
Xbit_r416_c38 bl[38] br[38] wl[416] vdd gnd cell_6t
Xbit_r417_c38 bl[38] br[38] wl[417] vdd gnd cell_6t
Xbit_r418_c38 bl[38] br[38] wl[418] vdd gnd cell_6t
Xbit_r419_c38 bl[38] br[38] wl[419] vdd gnd cell_6t
Xbit_r420_c38 bl[38] br[38] wl[420] vdd gnd cell_6t
Xbit_r421_c38 bl[38] br[38] wl[421] vdd gnd cell_6t
Xbit_r422_c38 bl[38] br[38] wl[422] vdd gnd cell_6t
Xbit_r423_c38 bl[38] br[38] wl[423] vdd gnd cell_6t
Xbit_r424_c38 bl[38] br[38] wl[424] vdd gnd cell_6t
Xbit_r425_c38 bl[38] br[38] wl[425] vdd gnd cell_6t
Xbit_r426_c38 bl[38] br[38] wl[426] vdd gnd cell_6t
Xbit_r427_c38 bl[38] br[38] wl[427] vdd gnd cell_6t
Xbit_r428_c38 bl[38] br[38] wl[428] vdd gnd cell_6t
Xbit_r429_c38 bl[38] br[38] wl[429] vdd gnd cell_6t
Xbit_r430_c38 bl[38] br[38] wl[430] vdd gnd cell_6t
Xbit_r431_c38 bl[38] br[38] wl[431] vdd gnd cell_6t
Xbit_r432_c38 bl[38] br[38] wl[432] vdd gnd cell_6t
Xbit_r433_c38 bl[38] br[38] wl[433] vdd gnd cell_6t
Xbit_r434_c38 bl[38] br[38] wl[434] vdd gnd cell_6t
Xbit_r435_c38 bl[38] br[38] wl[435] vdd gnd cell_6t
Xbit_r436_c38 bl[38] br[38] wl[436] vdd gnd cell_6t
Xbit_r437_c38 bl[38] br[38] wl[437] vdd gnd cell_6t
Xbit_r438_c38 bl[38] br[38] wl[438] vdd gnd cell_6t
Xbit_r439_c38 bl[38] br[38] wl[439] vdd gnd cell_6t
Xbit_r440_c38 bl[38] br[38] wl[440] vdd gnd cell_6t
Xbit_r441_c38 bl[38] br[38] wl[441] vdd gnd cell_6t
Xbit_r442_c38 bl[38] br[38] wl[442] vdd gnd cell_6t
Xbit_r443_c38 bl[38] br[38] wl[443] vdd gnd cell_6t
Xbit_r444_c38 bl[38] br[38] wl[444] vdd gnd cell_6t
Xbit_r445_c38 bl[38] br[38] wl[445] vdd gnd cell_6t
Xbit_r446_c38 bl[38] br[38] wl[446] vdd gnd cell_6t
Xbit_r447_c38 bl[38] br[38] wl[447] vdd gnd cell_6t
Xbit_r448_c38 bl[38] br[38] wl[448] vdd gnd cell_6t
Xbit_r449_c38 bl[38] br[38] wl[449] vdd gnd cell_6t
Xbit_r450_c38 bl[38] br[38] wl[450] vdd gnd cell_6t
Xbit_r451_c38 bl[38] br[38] wl[451] vdd gnd cell_6t
Xbit_r452_c38 bl[38] br[38] wl[452] vdd gnd cell_6t
Xbit_r453_c38 bl[38] br[38] wl[453] vdd gnd cell_6t
Xbit_r454_c38 bl[38] br[38] wl[454] vdd gnd cell_6t
Xbit_r455_c38 bl[38] br[38] wl[455] vdd gnd cell_6t
Xbit_r456_c38 bl[38] br[38] wl[456] vdd gnd cell_6t
Xbit_r457_c38 bl[38] br[38] wl[457] vdd gnd cell_6t
Xbit_r458_c38 bl[38] br[38] wl[458] vdd gnd cell_6t
Xbit_r459_c38 bl[38] br[38] wl[459] vdd gnd cell_6t
Xbit_r460_c38 bl[38] br[38] wl[460] vdd gnd cell_6t
Xbit_r461_c38 bl[38] br[38] wl[461] vdd gnd cell_6t
Xbit_r462_c38 bl[38] br[38] wl[462] vdd gnd cell_6t
Xbit_r463_c38 bl[38] br[38] wl[463] vdd gnd cell_6t
Xbit_r464_c38 bl[38] br[38] wl[464] vdd gnd cell_6t
Xbit_r465_c38 bl[38] br[38] wl[465] vdd gnd cell_6t
Xbit_r466_c38 bl[38] br[38] wl[466] vdd gnd cell_6t
Xbit_r467_c38 bl[38] br[38] wl[467] vdd gnd cell_6t
Xbit_r468_c38 bl[38] br[38] wl[468] vdd gnd cell_6t
Xbit_r469_c38 bl[38] br[38] wl[469] vdd gnd cell_6t
Xbit_r470_c38 bl[38] br[38] wl[470] vdd gnd cell_6t
Xbit_r471_c38 bl[38] br[38] wl[471] vdd gnd cell_6t
Xbit_r472_c38 bl[38] br[38] wl[472] vdd gnd cell_6t
Xbit_r473_c38 bl[38] br[38] wl[473] vdd gnd cell_6t
Xbit_r474_c38 bl[38] br[38] wl[474] vdd gnd cell_6t
Xbit_r475_c38 bl[38] br[38] wl[475] vdd gnd cell_6t
Xbit_r476_c38 bl[38] br[38] wl[476] vdd gnd cell_6t
Xbit_r477_c38 bl[38] br[38] wl[477] vdd gnd cell_6t
Xbit_r478_c38 bl[38] br[38] wl[478] vdd gnd cell_6t
Xbit_r479_c38 bl[38] br[38] wl[479] vdd gnd cell_6t
Xbit_r480_c38 bl[38] br[38] wl[480] vdd gnd cell_6t
Xbit_r481_c38 bl[38] br[38] wl[481] vdd gnd cell_6t
Xbit_r482_c38 bl[38] br[38] wl[482] vdd gnd cell_6t
Xbit_r483_c38 bl[38] br[38] wl[483] vdd gnd cell_6t
Xbit_r484_c38 bl[38] br[38] wl[484] vdd gnd cell_6t
Xbit_r485_c38 bl[38] br[38] wl[485] vdd gnd cell_6t
Xbit_r486_c38 bl[38] br[38] wl[486] vdd gnd cell_6t
Xbit_r487_c38 bl[38] br[38] wl[487] vdd gnd cell_6t
Xbit_r488_c38 bl[38] br[38] wl[488] vdd gnd cell_6t
Xbit_r489_c38 bl[38] br[38] wl[489] vdd gnd cell_6t
Xbit_r490_c38 bl[38] br[38] wl[490] vdd gnd cell_6t
Xbit_r491_c38 bl[38] br[38] wl[491] vdd gnd cell_6t
Xbit_r492_c38 bl[38] br[38] wl[492] vdd gnd cell_6t
Xbit_r493_c38 bl[38] br[38] wl[493] vdd gnd cell_6t
Xbit_r494_c38 bl[38] br[38] wl[494] vdd gnd cell_6t
Xbit_r495_c38 bl[38] br[38] wl[495] vdd gnd cell_6t
Xbit_r496_c38 bl[38] br[38] wl[496] vdd gnd cell_6t
Xbit_r497_c38 bl[38] br[38] wl[497] vdd gnd cell_6t
Xbit_r498_c38 bl[38] br[38] wl[498] vdd gnd cell_6t
Xbit_r499_c38 bl[38] br[38] wl[499] vdd gnd cell_6t
Xbit_r500_c38 bl[38] br[38] wl[500] vdd gnd cell_6t
Xbit_r501_c38 bl[38] br[38] wl[501] vdd gnd cell_6t
Xbit_r502_c38 bl[38] br[38] wl[502] vdd gnd cell_6t
Xbit_r503_c38 bl[38] br[38] wl[503] vdd gnd cell_6t
Xbit_r504_c38 bl[38] br[38] wl[504] vdd gnd cell_6t
Xbit_r505_c38 bl[38] br[38] wl[505] vdd gnd cell_6t
Xbit_r506_c38 bl[38] br[38] wl[506] vdd gnd cell_6t
Xbit_r507_c38 bl[38] br[38] wl[507] vdd gnd cell_6t
Xbit_r508_c38 bl[38] br[38] wl[508] vdd gnd cell_6t
Xbit_r509_c38 bl[38] br[38] wl[509] vdd gnd cell_6t
Xbit_r510_c38 bl[38] br[38] wl[510] vdd gnd cell_6t
Xbit_r511_c38 bl[38] br[38] wl[511] vdd gnd cell_6t
Xbit_r0_c39 bl[39] br[39] wl[0] vdd gnd cell_6t
Xbit_r1_c39 bl[39] br[39] wl[1] vdd gnd cell_6t
Xbit_r2_c39 bl[39] br[39] wl[2] vdd gnd cell_6t
Xbit_r3_c39 bl[39] br[39] wl[3] vdd gnd cell_6t
Xbit_r4_c39 bl[39] br[39] wl[4] vdd gnd cell_6t
Xbit_r5_c39 bl[39] br[39] wl[5] vdd gnd cell_6t
Xbit_r6_c39 bl[39] br[39] wl[6] vdd gnd cell_6t
Xbit_r7_c39 bl[39] br[39] wl[7] vdd gnd cell_6t
Xbit_r8_c39 bl[39] br[39] wl[8] vdd gnd cell_6t
Xbit_r9_c39 bl[39] br[39] wl[9] vdd gnd cell_6t
Xbit_r10_c39 bl[39] br[39] wl[10] vdd gnd cell_6t
Xbit_r11_c39 bl[39] br[39] wl[11] vdd gnd cell_6t
Xbit_r12_c39 bl[39] br[39] wl[12] vdd gnd cell_6t
Xbit_r13_c39 bl[39] br[39] wl[13] vdd gnd cell_6t
Xbit_r14_c39 bl[39] br[39] wl[14] vdd gnd cell_6t
Xbit_r15_c39 bl[39] br[39] wl[15] vdd gnd cell_6t
Xbit_r16_c39 bl[39] br[39] wl[16] vdd gnd cell_6t
Xbit_r17_c39 bl[39] br[39] wl[17] vdd gnd cell_6t
Xbit_r18_c39 bl[39] br[39] wl[18] vdd gnd cell_6t
Xbit_r19_c39 bl[39] br[39] wl[19] vdd gnd cell_6t
Xbit_r20_c39 bl[39] br[39] wl[20] vdd gnd cell_6t
Xbit_r21_c39 bl[39] br[39] wl[21] vdd gnd cell_6t
Xbit_r22_c39 bl[39] br[39] wl[22] vdd gnd cell_6t
Xbit_r23_c39 bl[39] br[39] wl[23] vdd gnd cell_6t
Xbit_r24_c39 bl[39] br[39] wl[24] vdd gnd cell_6t
Xbit_r25_c39 bl[39] br[39] wl[25] vdd gnd cell_6t
Xbit_r26_c39 bl[39] br[39] wl[26] vdd gnd cell_6t
Xbit_r27_c39 bl[39] br[39] wl[27] vdd gnd cell_6t
Xbit_r28_c39 bl[39] br[39] wl[28] vdd gnd cell_6t
Xbit_r29_c39 bl[39] br[39] wl[29] vdd gnd cell_6t
Xbit_r30_c39 bl[39] br[39] wl[30] vdd gnd cell_6t
Xbit_r31_c39 bl[39] br[39] wl[31] vdd gnd cell_6t
Xbit_r32_c39 bl[39] br[39] wl[32] vdd gnd cell_6t
Xbit_r33_c39 bl[39] br[39] wl[33] vdd gnd cell_6t
Xbit_r34_c39 bl[39] br[39] wl[34] vdd gnd cell_6t
Xbit_r35_c39 bl[39] br[39] wl[35] vdd gnd cell_6t
Xbit_r36_c39 bl[39] br[39] wl[36] vdd gnd cell_6t
Xbit_r37_c39 bl[39] br[39] wl[37] vdd gnd cell_6t
Xbit_r38_c39 bl[39] br[39] wl[38] vdd gnd cell_6t
Xbit_r39_c39 bl[39] br[39] wl[39] vdd gnd cell_6t
Xbit_r40_c39 bl[39] br[39] wl[40] vdd gnd cell_6t
Xbit_r41_c39 bl[39] br[39] wl[41] vdd gnd cell_6t
Xbit_r42_c39 bl[39] br[39] wl[42] vdd gnd cell_6t
Xbit_r43_c39 bl[39] br[39] wl[43] vdd gnd cell_6t
Xbit_r44_c39 bl[39] br[39] wl[44] vdd gnd cell_6t
Xbit_r45_c39 bl[39] br[39] wl[45] vdd gnd cell_6t
Xbit_r46_c39 bl[39] br[39] wl[46] vdd gnd cell_6t
Xbit_r47_c39 bl[39] br[39] wl[47] vdd gnd cell_6t
Xbit_r48_c39 bl[39] br[39] wl[48] vdd gnd cell_6t
Xbit_r49_c39 bl[39] br[39] wl[49] vdd gnd cell_6t
Xbit_r50_c39 bl[39] br[39] wl[50] vdd gnd cell_6t
Xbit_r51_c39 bl[39] br[39] wl[51] vdd gnd cell_6t
Xbit_r52_c39 bl[39] br[39] wl[52] vdd gnd cell_6t
Xbit_r53_c39 bl[39] br[39] wl[53] vdd gnd cell_6t
Xbit_r54_c39 bl[39] br[39] wl[54] vdd gnd cell_6t
Xbit_r55_c39 bl[39] br[39] wl[55] vdd gnd cell_6t
Xbit_r56_c39 bl[39] br[39] wl[56] vdd gnd cell_6t
Xbit_r57_c39 bl[39] br[39] wl[57] vdd gnd cell_6t
Xbit_r58_c39 bl[39] br[39] wl[58] vdd gnd cell_6t
Xbit_r59_c39 bl[39] br[39] wl[59] vdd gnd cell_6t
Xbit_r60_c39 bl[39] br[39] wl[60] vdd gnd cell_6t
Xbit_r61_c39 bl[39] br[39] wl[61] vdd gnd cell_6t
Xbit_r62_c39 bl[39] br[39] wl[62] vdd gnd cell_6t
Xbit_r63_c39 bl[39] br[39] wl[63] vdd gnd cell_6t
Xbit_r64_c39 bl[39] br[39] wl[64] vdd gnd cell_6t
Xbit_r65_c39 bl[39] br[39] wl[65] vdd gnd cell_6t
Xbit_r66_c39 bl[39] br[39] wl[66] vdd gnd cell_6t
Xbit_r67_c39 bl[39] br[39] wl[67] vdd gnd cell_6t
Xbit_r68_c39 bl[39] br[39] wl[68] vdd gnd cell_6t
Xbit_r69_c39 bl[39] br[39] wl[69] vdd gnd cell_6t
Xbit_r70_c39 bl[39] br[39] wl[70] vdd gnd cell_6t
Xbit_r71_c39 bl[39] br[39] wl[71] vdd gnd cell_6t
Xbit_r72_c39 bl[39] br[39] wl[72] vdd gnd cell_6t
Xbit_r73_c39 bl[39] br[39] wl[73] vdd gnd cell_6t
Xbit_r74_c39 bl[39] br[39] wl[74] vdd gnd cell_6t
Xbit_r75_c39 bl[39] br[39] wl[75] vdd gnd cell_6t
Xbit_r76_c39 bl[39] br[39] wl[76] vdd gnd cell_6t
Xbit_r77_c39 bl[39] br[39] wl[77] vdd gnd cell_6t
Xbit_r78_c39 bl[39] br[39] wl[78] vdd gnd cell_6t
Xbit_r79_c39 bl[39] br[39] wl[79] vdd gnd cell_6t
Xbit_r80_c39 bl[39] br[39] wl[80] vdd gnd cell_6t
Xbit_r81_c39 bl[39] br[39] wl[81] vdd gnd cell_6t
Xbit_r82_c39 bl[39] br[39] wl[82] vdd gnd cell_6t
Xbit_r83_c39 bl[39] br[39] wl[83] vdd gnd cell_6t
Xbit_r84_c39 bl[39] br[39] wl[84] vdd gnd cell_6t
Xbit_r85_c39 bl[39] br[39] wl[85] vdd gnd cell_6t
Xbit_r86_c39 bl[39] br[39] wl[86] vdd gnd cell_6t
Xbit_r87_c39 bl[39] br[39] wl[87] vdd gnd cell_6t
Xbit_r88_c39 bl[39] br[39] wl[88] vdd gnd cell_6t
Xbit_r89_c39 bl[39] br[39] wl[89] vdd gnd cell_6t
Xbit_r90_c39 bl[39] br[39] wl[90] vdd gnd cell_6t
Xbit_r91_c39 bl[39] br[39] wl[91] vdd gnd cell_6t
Xbit_r92_c39 bl[39] br[39] wl[92] vdd gnd cell_6t
Xbit_r93_c39 bl[39] br[39] wl[93] vdd gnd cell_6t
Xbit_r94_c39 bl[39] br[39] wl[94] vdd gnd cell_6t
Xbit_r95_c39 bl[39] br[39] wl[95] vdd gnd cell_6t
Xbit_r96_c39 bl[39] br[39] wl[96] vdd gnd cell_6t
Xbit_r97_c39 bl[39] br[39] wl[97] vdd gnd cell_6t
Xbit_r98_c39 bl[39] br[39] wl[98] vdd gnd cell_6t
Xbit_r99_c39 bl[39] br[39] wl[99] vdd gnd cell_6t
Xbit_r100_c39 bl[39] br[39] wl[100] vdd gnd cell_6t
Xbit_r101_c39 bl[39] br[39] wl[101] vdd gnd cell_6t
Xbit_r102_c39 bl[39] br[39] wl[102] vdd gnd cell_6t
Xbit_r103_c39 bl[39] br[39] wl[103] vdd gnd cell_6t
Xbit_r104_c39 bl[39] br[39] wl[104] vdd gnd cell_6t
Xbit_r105_c39 bl[39] br[39] wl[105] vdd gnd cell_6t
Xbit_r106_c39 bl[39] br[39] wl[106] vdd gnd cell_6t
Xbit_r107_c39 bl[39] br[39] wl[107] vdd gnd cell_6t
Xbit_r108_c39 bl[39] br[39] wl[108] vdd gnd cell_6t
Xbit_r109_c39 bl[39] br[39] wl[109] vdd gnd cell_6t
Xbit_r110_c39 bl[39] br[39] wl[110] vdd gnd cell_6t
Xbit_r111_c39 bl[39] br[39] wl[111] vdd gnd cell_6t
Xbit_r112_c39 bl[39] br[39] wl[112] vdd gnd cell_6t
Xbit_r113_c39 bl[39] br[39] wl[113] vdd gnd cell_6t
Xbit_r114_c39 bl[39] br[39] wl[114] vdd gnd cell_6t
Xbit_r115_c39 bl[39] br[39] wl[115] vdd gnd cell_6t
Xbit_r116_c39 bl[39] br[39] wl[116] vdd gnd cell_6t
Xbit_r117_c39 bl[39] br[39] wl[117] vdd gnd cell_6t
Xbit_r118_c39 bl[39] br[39] wl[118] vdd gnd cell_6t
Xbit_r119_c39 bl[39] br[39] wl[119] vdd gnd cell_6t
Xbit_r120_c39 bl[39] br[39] wl[120] vdd gnd cell_6t
Xbit_r121_c39 bl[39] br[39] wl[121] vdd gnd cell_6t
Xbit_r122_c39 bl[39] br[39] wl[122] vdd gnd cell_6t
Xbit_r123_c39 bl[39] br[39] wl[123] vdd gnd cell_6t
Xbit_r124_c39 bl[39] br[39] wl[124] vdd gnd cell_6t
Xbit_r125_c39 bl[39] br[39] wl[125] vdd gnd cell_6t
Xbit_r126_c39 bl[39] br[39] wl[126] vdd gnd cell_6t
Xbit_r127_c39 bl[39] br[39] wl[127] vdd gnd cell_6t
Xbit_r128_c39 bl[39] br[39] wl[128] vdd gnd cell_6t
Xbit_r129_c39 bl[39] br[39] wl[129] vdd gnd cell_6t
Xbit_r130_c39 bl[39] br[39] wl[130] vdd gnd cell_6t
Xbit_r131_c39 bl[39] br[39] wl[131] vdd gnd cell_6t
Xbit_r132_c39 bl[39] br[39] wl[132] vdd gnd cell_6t
Xbit_r133_c39 bl[39] br[39] wl[133] vdd gnd cell_6t
Xbit_r134_c39 bl[39] br[39] wl[134] vdd gnd cell_6t
Xbit_r135_c39 bl[39] br[39] wl[135] vdd gnd cell_6t
Xbit_r136_c39 bl[39] br[39] wl[136] vdd gnd cell_6t
Xbit_r137_c39 bl[39] br[39] wl[137] vdd gnd cell_6t
Xbit_r138_c39 bl[39] br[39] wl[138] vdd gnd cell_6t
Xbit_r139_c39 bl[39] br[39] wl[139] vdd gnd cell_6t
Xbit_r140_c39 bl[39] br[39] wl[140] vdd gnd cell_6t
Xbit_r141_c39 bl[39] br[39] wl[141] vdd gnd cell_6t
Xbit_r142_c39 bl[39] br[39] wl[142] vdd gnd cell_6t
Xbit_r143_c39 bl[39] br[39] wl[143] vdd gnd cell_6t
Xbit_r144_c39 bl[39] br[39] wl[144] vdd gnd cell_6t
Xbit_r145_c39 bl[39] br[39] wl[145] vdd gnd cell_6t
Xbit_r146_c39 bl[39] br[39] wl[146] vdd gnd cell_6t
Xbit_r147_c39 bl[39] br[39] wl[147] vdd gnd cell_6t
Xbit_r148_c39 bl[39] br[39] wl[148] vdd gnd cell_6t
Xbit_r149_c39 bl[39] br[39] wl[149] vdd gnd cell_6t
Xbit_r150_c39 bl[39] br[39] wl[150] vdd gnd cell_6t
Xbit_r151_c39 bl[39] br[39] wl[151] vdd gnd cell_6t
Xbit_r152_c39 bl[39] br[39] wl[152] vdd gnd cell_6t
Xbit_r153_c39 bl[39] br[39] wl[153] vdd gnd cell_6t
Xbit_r154_c39 bl[39] br[39] wl[154] vdd gnd cell_6t
Xbit_r155_c39 bl[39] br[39] wl[155] vdd gnd cell_6t
Xbit_r156_c39 bl[39] br[39] wl[156] vdd gnd cell_6t
Xbit_r157_c39 bl[39] br[39] wl[157] vdd gnd cell_6t
Xbit_r158_c39 bl[39] br[39] wl[158] vdd gnd cell_6t
Xbit_r159_c39 bl[39] br[39] wl[159] vdd gnd cell_6t
Xbit_r160_c39 bl[39] br[39] wl[160] vdd gnd cell_6t
Xbit_r161_c39 bl[39] br[39] wl[161] vdd gnd cell_6t
Xbit_r162_c39 bl[39] br[39] wl[162] vdd gnd cell_6t
Xbit_r163_c39 bl[39] br[39] wl[163] vdd gnd cell_6t
Xbit_r164_c39 bl[39] br[39] wl[164] vdd gnd cell_6t
Xbit_r165_c39 bl[39] br[39] wl[165] vdd gnd cell_6t
Xbit_r166_c39 bl[39] br[39] wl[166] vdd gnd cell_6t
Xbit_r167_c39 bl[39] br[39] wl[167] vdd gnd cell_6t
Xbit_r168_c39 bl[39] br[39] wl[168] vdd gnd cell_6t
Xbit_r169_c39 bl[39] br[39] wl[169] vdd gnd cell_6t
Xbit_r170_c39 bl[39] br[39] wl[170] vdd gnd cell_6t
Xbit_r171_c39 bl[39] br[39] wl[171] vdd gnd cell_6t
Xbit_r172_c39 bl[39] br[39] wl[172] vdd gnd cell_6t
Xbit_r173_c39 bl[39] br[39] wl[173] vdd gnd cell_6t
Xbit_r174_c39 bl[39] br[39] wl[174] vdd gnd cell_6t
Xbit_r175_c39 bl[39] br[39] wl[175] vdd gnd cell_6t
Xbit_r176_c39 bl[39] br[39] wl[176] vdd gnd cell_6t
Xbit_r177_c39 bl[39] br[39] wl[177] vdd gnd cell_6t
Xbit_r178_c39 bl[39] br[39] wl[178] vdd gnd cell_6t
Xbit_r179_c39 bl[39] br[39] wl[179] vdd gnd cell_6t
Xbit_r180_c39 bl[39] br[39] wl[180] vdd gnd cell_6t
Xbit_r181_c39 bl[39] br[39] wl[181] vdd gnd cell_6t
Xbit_r182_c39 bl[39] br[39] wl[182] vdd gnd cell_6t
Xbit_r183_c39 bl[39] br[39] wl[183] vdd gnd cell_6t
Xbit_r184_c39 bl[39] br[39] wl[184] vdd gnd cell_6t
Xbit_r185_c39 bl[39] br[39] wl[185] vdd gnd cell_6t
Xbit_r186_c39 bl[39] br[39] wl[186] vdd gnd cell_6t
Xbit_r187_c39 bl[39] br[39] wl[187] vdd gnd cell_6t
Xbit_r188_c39 bl[39] br[39] wl[188] vdd gnd cell_6t
Xbit_r189_c39 bl[39] br[39] wl[189] vdd gnd cell_6t
Xbit_r190_c39 bl[39] br[39] wl[190] vdd gnd cell_6t
Xbit_r191_c39 bl[39] br[39] wl[191] vdd gnd cell_6t
Xbit_r192_c39 bl[39] br[39] wl[192] vdd gnd cell_6t
Xbit_r193_c39 bl[39] br[39] wl[193] vdd gnd cell_6t
Xbit_r194_c39 bl[39] br[39] wl[194] vdd gnd cell_6t
Xbit_r195_c39 bl[39] br[39] wl[195] vdd gnd cell_6t
Xbit_r196_c39 bl[39] br[39] wl[196] vdd gnd cell_6t
Xbit_r197_c39 bl[39] br[39] wl[197] vdd gnd cell_6t
Xbit_r198_c39 bl[39] br[39] wl[198] vdd gnd cell_6t
Xbit_r199_c39 bl[39] br[39] wl[199] vdd gnd cell_6t
Xbit_r200_c39 bl[39] br[39] wl[200] vdd gnd cell_6t
Xbit_r201_c39 bl[39] br[39] wl[201] vdd gnd cell_6t
Xbit_r202_c39 bl[39] br[39] wl[202] vdd gnd cell_6t
Xbit_r203_c39 bl[39] br[39] wl[203] vdd gnd cell_6t
Xbit_r204_c39 bl[39] br[39] wl[204] vdd gnd cell_6t
Xbit_r205_c39 bl[39] br[39] wl[205] vdd gnd cell_6t
Xbit_r206_c39 bl[39] br[39] wl[206] vdd gnd cell_6t
Xbit_r207_c39 bl[39] br[39] wl[207] vdd gnd cell_6t
Xbit_r208_c39 bl[39] br[39] wl[208] vdd gnd cell_6t
Xbit_r209_c39 bl[39] br[39] wl[209] vdd gnd cell_6t
Xbit_r210_c39 bl[39] br[39] wl[210] vdd gnd cell_6t
Xbit_r211_c39 bl[39] br[39] wl[211] vdd gnd cell_6t
Xbit_r212_c39 bl[39] br[39] wl[212] vdd gnd cell_6t
Xbit_r213_c39 bl[39] br[39] wl[213] vdd gnd cell_6t
Xbit_r214_c39 bl[39] br[39] wl[214] vdd gnd cell_6t
Xbit_r215_c39 bl[39] br[39] wl[215] vdd gnd cell_6t
Xbit_r216_c39 bl[39] br[39] wl[216] vdd gnd cell_6t
Xbit_r217_c39 bl[39] br[39] wl[217] vdd gnd cell_6t
Xbit_r218_c39 bl[39] br[39] wl[218] vdd gnd cell_6t
Xbit_r219_c39 bl[39] br[39] wl[219] vdd gnd cell_6t
Xbit_r220_c39 bl[39] br[39] wl[220] vdd gnd cell_6t
Xbit_r221_c39 bl[39] br[39] wl[221] vdd gnd cell_6t
Xbit_r222_c39 bl[39] br[39] wl[222] vdd gnd cell_6t
Xbit_r223_c39 bl[39] br[39] wl[223] vdd gnd cell_6t
Xbit_r224_c39 bl[39] br[39] wl[224] vdd gnd cell_6t
Xbit_r225_c39 bl[39] br[39] wl[225] vdd gnd cell_6t
Xbit_r226_c39 bl[39] br[39] wl[226] vdd gnd cell_6t
Xbit_r227_c39 bl[39] br[39] wl[227] vdd gnd cell_6t
Xbit_r228_c39 bl[39] br[39] wl[228] vdd gnd cell_6t
Xbit_r229_c39 bl[39] br[39] wl[229] vdd gnd cell_6t
Xbit_r230_c39 bl[39] br[39] wl[230] vdd gnd cell_6t
Xbit_r231_c39 bl[39] br[39] wl[231] vdd gnd cell_6t
Xbit_r232_c39 bl[39] br[39] wl[232] vdd gnd cell_6t
Xbit_r233_c39 bl[39] br[39] wl[233] vdd gnd cell_6t
Xbit_r234_c39 bl[39] br[39] wl[234] vdd gnd cell_6t
Xbit_r235_c39 bl[39] br[39] wl[235] vdd gnd cell_6t
Xbit_r236_c39 bl[39] br[39] wl[236] vdd gnd cell_6t
Xbit_r237_c39 bl[39] br[39] wl[237] vdd gnd cell_6t
Xbit_r238_c39 bl[39] br[39] wl[238] vdd gnd cell_6t
Xbit_r239_c39 bl[39] br[39] wl[239] vdd gnd cell_6t
Xbit_r240_c39 bl[39] br[39] wl[240] vdd gnd cell_6t
Xbit_r241_c39 bl[39] br[39] wl[241] vdd gnd cell_6t
Xbit_r242_c39 bl[39] br[39] wl[242] vdd gnd cell_6t
Xbit_r243_c39 bl[39] br[39] wl[243] vdd gnd cell_6t
Xbit_r244_c39 bl[39] br[39] wl[244] vdd gnd cell_6t
Xbit_r245_c39 bl[39] br[39] wl[245] vdd gnd cell_6t
Xbit_r246_c39 bl[39] br[39] wl[246] vdd gnd cell_6t
Xbit_r247_c39 bl[39] br[39] wl[247] vdd gnd cell_6t
Xbit_r248_c39 bl[39] br[39] wl[248] vdd gnd cell_6t
Xbit_r249_c39 bl[39] br[39] wl[249] vdd gnd cell_6t
Xbit_r250_c39 bl[39] br[39] wl[250] vdd gnd cell_6t
Xbit_r251_c39 bl[39] br[39] wl[251] vdd gnd cell_6t
Xbit_r252_c39 bl[39] br[39] wl[252] vdd gnd cell_6t
Xbit_r253_c39 bl[39] br[39] wl[253] vdd gnd cell_6t
Xbit_r254_c39 bl[39] br[39] wl[254] vdd gnd cell_6t
Xbit_r255_c39 bl[39] br[39] wl[255] vdd gnd cell_6t
Xbit_r256_c39 bl[39] br[39] wl[256] vdd gnd cell_6t
Xbit_r257_c39 bl[39] br[39] wl[257] vdd gnd cell_6t
Xbit_r258_c39 bl[39] br[39] wl[258] vdd gnd cell_6t
Xbit_r259_c39 bl[39] br[39] wl[259] vdd gnd cell_6t
Xbit_r260_c39 bl[39] br[39] wl[260] vdd gnd cell_6t
Xbit_r261_c39 bl[39] br[39] wl[261] vdd gnd cell_6t
Xbit_r262_c39 bl[39] br[39] wl[262] vdd gnd cell_6t
Xbit_r263_c39 bl[39] br[39] wl[263] vdd gnd cell_6t
Xbit_r264_c39 bl[39] br[39] wl[264] vdd gnd cell_6t
Xbit_r265_c39 bl[39] br[39] wl[265] vdd gnd cell_6t
Xbit_r266_c39 bl[39] br[39] wl[266] vdd gnd cell_6t
Xbit_r267_c39 bl[39] br[39] wl[267] vdd gnd cell_6t
Xbit_r268_c39 bl[39] br[39] wl[268] vdd gnd cell_6t
Xbit_r269_c39 bl[39] br[39] wl[269] vdd gnd cell_6t
Xbit_r270_c39 bl[39] br[39] wl[270] vdd gnd cell_6t
Xbit_r271_c39 bl[39] br[39] wl[271] vdd gnd cell_6t
Xbit_r272_c39 bl[39] br[39] wl[272] vdd gnd cell_6t
Xbit_r273_c39 bl[39] br[39] wl[273] vdd gnd cell_6t
Xbit_r274_c39 bl[39] br[39] wl[274] vdd gnd cell_6t
Xbit_r275_c39 bl[39] br[39] wl[275] vdd gnd cell_6t
Xbit_r276_c39 bl[39] br[39] wl[276] vdd gnd cell_6t
Xbit_r277_c39 bl[39] br[39] wl[277] vdd gnd cell_6t
Xbit_r278_c39 bl[39] br[39] wl[278] vdd gnd cell_6t
Xbit_r279_c39 bl[39] br[39] wl[279] vdd gnd cell_6t
Xbit_r280_c39 bl[39] br[39] wl[280] vdd gnd cell_6t
Xbit_r281_c39 bl[39] br[39] wl[281] vdd gnd cell_6t
Xbit_r282_c39 bl[39] br[39] wl[282] vdd gnd cell_6t
Xbit_r283_c39 bl[39] br[39] wl[283] vdd gnd cell_6t
Xbit_r284_c39 bl[39] br[39] wl[284] vdd gnd cell_6t
Xbit_r285_c39 bl[39] br[39] wl[285] vdd gnd cell_6t
Xbit_r286_c39 bl[39] br[39] wl[286] vdd gnd cell_6t
Xbit_r287_c39 bl[39] br[39] wl[287] vdd gnd cell_6t
Xbit_r288_c39 bl[39] br[39] wl[288] vdd gnd cell_6t
Xbit_r289_c39 bl[39] br[39] wl[289] vdd gnd cell_6t
Xbit_r290_c39 bl[39] br[39] wl[290] vdd gnd cell_6t
Xbit_r291_c39 bl[39] br[39] wl[291] vdd gnd cell_6t
Xbit_r292_c39 bl[39] br[39] wl[292] vdd gnd cell_6t
Xbit_r293_c39 bl[39] br[39] wl[293] vdd gnd cell_6t
Xbit_r294_c39 bl[39] br[39] wl[294] vdd gnd cell_6t
Xbit_r295_c39 bl[39] br[39] wl[295] vdd gnd cell_6t
Xbit_r296_c39 bl[39] br[39] wl[296] vdd gnd cell_6t
Xbit_r297_c39 bl[39] br[39] wl[297] vdd gnd cell_6t
Xbit_r298_c39 bl[39] br[39] wl[298] vdd gnd cell_6t
Xbit_r299_c39 bl[39] br[39] wl[299] vdd gnd cell_6t
Xbit_r300_c39 bl[39] br[39] wl[300] vdd gnd cell_6t
Xbit_r301_c39 bl[39] br[39] wl[301] vdd gnd cell_6t
Xbit_r302_c39 bl[39] br[39] wl[302] vdd gnd cell_6t
Xbit_r303_c39 bl[39] br[39] wl[303] vdd gnd cell_6t
Xbit_r304_c39 bl[39] br[39] wl[304] vdd gnd cell_6t
Xbit_r305_c39 bl[39] br[39] wl[305] vdd gnd cell_6t
Xbit_r306_c39 bl[39] br[39] wl[306] vdd gnd cell_6t
Xbit_r307_c39 bl[39] br[39] wl[307] vdd gnd cell_6t
Xbit_r308_c39 bl[39] br[39] wl[308] vdd gnd cell_6t
Xbit_r309_c39 bl[39] br[39] wl[309] vdd gnd cell_6t
Xbit_r310_c39 bl[39] br[39] wl[310] vdd gnd cell_6t
Xbit_r311_c39 bl[39] br[39] wl[311] vdd gnd cell_6t
Xbit_r312_c39 bl[39] br[39] wl[312] vdd gnd cell_6t
Xbit_r313_c39 bl[39] br[39] wl[313] vdd gnd cell_6t
Xbit_r314_c39 bl[39] br[39] wl[314] vdd gnd cell_6t
Xbit_r315_c39 bl[39] br[39] wl[315] vdd gnd cell_6t
Xbit_r316_c39 bl[39] br[39] wl[316] vdd gnd cell_6t
Xbit_r317_c39 bl[39] br[39] wl[317] vdd gnd cell_6t
Xbit_r318_c39 bl[39] br[39] wl[318] vdd gnd cell_6t
Xbit_r319_c39 bl[39] br[39] wl[319] vdd gnd cell_6t
Xbit_r320_c39 bl[39] br[39] wl[320] vdd gnd cell_6t
Xbit_r321_c39 bl[39] br[39] wl[321] vdd gnd cell_6t
Xbit_r322_c39 bl[39] br[39] wl[322] vdd gnd cell_6t
Xbit_r323_c39 bl[39] br[39] wl[323] vdd gnd cell_6t
Xbit_r324_c39 bl[39] br[39] wl[324] vdd gnd cell_6t
Xbit_r325_c39 bl[39] br[39] wl[325] vdd gnd cell_6t
Xbit_r326_c39 bl[39] br[39] wl[326] vdd gnd cell_6t
Xbit_r327_c39 bl[39] br[39] wl[327] vdd gnd cell_6t
Xbit_r328_c39 bl[39] br[39] wl[328] vdd gnd cell_6t
Xbit_r329_c39 bl[39] br[39] wl[329] vdd gnd cell_6t
Xbit_r330_c39 bl[39] br[39] wl[330] vdd gnd cell_6t
Xbit_r331_c39 bl[39] br[39] wl[331] vdd gnd cell_6t
Xbit_r332_c39 bl[39] br[39] wl[332] vdd gnd cell_6t
Xbit_r333_c39 bl[39] br[39] wl[333] vdd gnd cell_6t
Xbit_r334_c39 bl[39] br[39] wl[334] vdd gnd cell_6t
Xbit_r335_c39 bl[39] br[39] wl[335] vdd gnd cell_6t
Xbit_r336_c39 bl[39] br[39] wl[336] vdd gnd cell_6t
Xbit_r337_c39 bl[39] br[39] wl[337] vdd gnd cell_6t
Xbit_r338_c39 bl[39] br[39] wl[338] vdd gnd cell_6t
Xbit_r339_c39 bl[39] br[39] wl[339] vdd gnd cell_6t
Xbit_r340_c39 bl[39] br[39] wl[340] vdd gnd cell_6t
Xbit_r341_c39 bl[39] br[39] wl[341] vdd gnd cell_6t
Xbit_r342_c39 bl[39] br[39] wl[342] vdd gnd cell_6t
Xbit_r343_c39 bl[39] br[39] wl[343] vdd gnd cell_6t
Xbit_r344_c39 bl[39] br[39] wl[344] vdd gnd cell_6t
Xbit_r345_c39 bl[39] br[39] wl[345] vdd gnd cell_6t
Xbit_r346_c39 bl[39] br[39] wl[346] vdd gnd cell_6t
Xbit_r347_c39 bl[39] br[39] wl[347] vdd gnd cell_6t
Xbit_r348_c39 bl[39] br[39] wl[348] vdd gnd cell_6t
Xbit_r349_c39 bl[39] br[39] wl[349] vdd gnd cell_6t
Xbit_r350_c39 bl[39] br[39] wl[350] vdd gnd cell_6t
Xbit_r351_c39 bl[39] br[39] wl[351] vdd gnd cell_6t
Xbit_r352_c39 bl[39] br[39] wl[352] vdd gnd cell_6t
Xbit_r353_c39 bl[39] br[39] wl[353] vdd gnd cell_6t
Xbit_r354_c39 bl[39] br[39] wl[354] vdd gnd cell_6t
Xbit_r355_c39 bl[39] br[39] wl[355] vdd gnd cell_6t
Xbit_r356_c39 bl[39] br[39] wl[356] vdd gnd cell_6t
Xbit_r357_c39 bl[39] br[39] wl[357] vdd gnd cell_6t
Xbit_r358_c39 bl[39] br[39] wl[358] vdd gnd cell_6t
Xbit_r359_c39 bl[39] br[39] wl[359] vdd gnd cell_6t
Xbit_r360_c39 bl[39] br[39] wl[360] vdd gnd cell_6t
Xbit_r361_c39 bl[39] br[39] wl[361] vdd gnd cell_6t
Xbit_r362_c39 bl[39] br[39] wl[362] vdd gnd cell_6t
Xbit_r363_c39 bl[39] br[39] wl[363] vdd gnd cell_6t
Xbit_r364_c39 bl[39] br[39] wl[364] vdd gnd cell_6t
Xbit_r365_c39 bl[39] br[39] wl[365] vdd gnd cell_6t
Xbit_r366_c39 bl[39] br[39] wl[366] vdd gnd cell_6t
Xbit_r367_c39 bl[39] br[39] wl[367] vdd gnd cell_6t
Xbit_r368_c39 bl[39] br[39] wl[368] vdd gnd cell_6t
Xbit_r369_c39 bl[39] br[39] wl[369] vdd gnd cell_6t
Xbit_r370_c39 bl[39] br[39] wl[370] vdd gnd cell_6t
Xbit_r371_c39 bl[39] br[39] wl[371] vdd gnd cell_6t
Xbit_r372_c39 bl[39] br[39] wl[372] vdd gnd cell_6t
Xbit_r373_c39 bl[39] br[39] wl[373] vdd gnd cell_6t
Xbit_r374_c39 bl[39] br[39] wl[374] vdd gnd cell_6t
Xbit_r375_c39 bl[39] br[39] wl[375] vdd gnd cell_6t
Xbit_r376_c39 bl[39] br[39] wl[376] vdd gnd cell_6t
Xbit_r377_c39 bl[39] br[39] wl[377] vdd gnd cell_6t
Xbit_r378_c39 bl[39] br[39] wl[378] vdd gnd cell_6t
Xbit_r379_c39 bl[39] br[39] wl[379] vdd gnd cell_6t
Xbit_r380_c39 bl[39] br[39] wl[380] vdd gnd cell_6t
Xbit_r381_c39 bl[39] br[39] wl[381] vdd gnd cell_6t
Xbit_r382_c39 bl[39] br[39] wl[382] vdd gnd cell_6t
Xbit_r383_c39 bl[39] br[39] wl[383] vdd gnd cell_6t
Xbit_r384_c39 bl[39] br[39] wl[384] vdd gnd cell_6t
Xbit_r385_c39 bl[39] br[39] wl[385] vdd gnd cell_6t
Xbit_r386_c39 bl[39] br[39] wl[386] vdd gnd cell_6t
Xbit_r387_c39 bl[39] br[39] wl[387] vdd gnd cell_6t
Xbit_r388_c39 bl[39] br[39] wl[388] vdd gnd cell_6t
Xbit_r389_c39 bl[39] br[39] wl[389] vdd gnd cell_6t
Xbit_r390_c39 bl[39] br[39] wl[390] vdd gnd cell_6t
Xbit_r391_c39 bl[39] br[39] wl[391] vdd gnd cell_6t
Xbit_r392_c39 bl[39] br[39] wl[392] vdd gnd cell_6t
Xbit_r393_c39 bl[39] br[39] wl[393] vdd gnd cell_6t
Xbit_r394_c39 bl[39] br[39] wl[394] vdd gnd cell_6t
Xbit_r395_c39 bl[39] br[39] wl[395] vdd gnd cell_6t
Xbit_r396_c39 bl[39] br[39] wl[396] vdd gnd cell_6t
Xbit_r397_c39 bl[39] br[39] wl[397] vdd gnd cell_6t
Xbit_r398_c39 bl[39] br[39] wl[398] vdd gnd cell_6t
Xbit_r399_c39 bl[39] br[39] wl[399] vdd gnd cell_6t
Xbit_r400_c39 bl[39] br[39] wl[400] vdd gnd cell_6t
Xbit_r401_c39 bl[39] br[39] wl[401] vdd gnd cell_6t
Xbit_r402_c39 bl[39] br[39] wl[402] vdd gnd cell_6t
Xbit_r403_c39 bl[39] br[39] wl[403] vdd gnd cell_6t
Xbit_r404_c39 bl[39] br[39] wl[404] vdd gnd cell_6t
Xbit_r405_c39 bl[39] br[39] wl[405] vdd gnd cell_6t
Xbit_r406_c39 bl[39] br[39] wl[406] vdd gnd cell_6t
Xbit_r407_c39 bl[39] br[39] wl[407] vdd gnd cell_6t
Xbit_r408_c39 bl[39] br[39] wl[408] vdd gnd cell_6t
Xbit_r409_c39 bl[39] br[39] wl[409] vdd gnd cell_6t
Xbit_r410_c39 bl[39] br[39] wl[410] vdd gnd cell_6t
Xbit_r411_c39 bl[39] br[39] wl[411] vdd gnd cell_6t
Xbit_r412_c39 bl[39] br[39] wl[412] vdd gnd cell_6t
Xbit_r413_c39 bl[39] br[39] wl[413] vdd gnd cell_6t
Xbit_r414_c39 bl[39] br[39] wl[414] vdd gnd cell_6t
Xbit_r415_c39 bl[39] br[39] wl[415] vdd gnd cell_6t
Xbit_r416_c39 bl[39] br[39] wl[416] vdd gnd cell_6t
Xbit_r417_c39 bl[39] br[39] wl[417] vdd gnd cell_6t
Xbit_r418_c39 bl[39] br[39] wl[418] vdd gnd cell_6t
Xbit_r419_c39 bl[39] br[39] wl[419] vdd gnd cell_6t
Xbit_r420_c39 bl[39] br[39] wl[420] vdd gnd cell_6t
Xbit_r421_c39 bl[39] br[39] wl[421] vdd gnd cell_6t
Xbit_r422_c39 bl[39] br[39] wl[422] vdd gnd cell_6t
Xbit_r423_c39 bl[39] br[39] wl[423] vdd gnd cell_6t
Xbit_r424_c39 bl[39] br[39] wl[424] vdd gnd cell_6t
Xbit_r425_c39 bl[39] br[39] wl[425] vdd gnd cell_6t
Xbit_r426_c39 bl[39] br[39] wl[426] vdd gnd cell_6t
Xbit_r427_c39 bl[39] br[39] wl[427] vdd gnd cell_6t
Xbit_r428_c39 bl[39] br[39] wl[428] vdd gnd cell_6t
Xbit_r429_c39 bl[39] br[39] wl[429] vdd gnd cell_6t
Xbit_r430_c39 bl[39] br[39] wl[430] vdd gnd cell_6t
Xbit_r431_c39 bl[39] br[39] wl[431] vdd gnd cell_6t
Xbit_r432_c39 bl[39] br[39] wl[432] vdd gnd cell_6t
Xbit_r433_c39 bl[39] br[39] wl[433] vdd gnd cell_6t
Xbit_r434_c39 bl[39] br[39] wl[434] vdd gnd cell_6t
Xbit_r435_c39 bl[39] br[39] wl[435] vdd gnd cell_6t
Xbit_r436_c39 bl[39] br[39] wl[436] vdd gnd cell_6t
Xbit_r437_c39 bl[39] br[39] wl[437] vdd gnd cell_6t
Xbit_r438_c39 bl[39] br[39] wl[438] vdd gnd cell_6t
Xbit_r439_c39 bl[39] br[39] wl[439] vdd gnd cell_6t
Xbit_r440_c39 bl[39] br[39] wl[440] vdd gnd cell_6t
Xbit_r441_c39 bl[39] br[39] wl[441] vdd gnd cell_6t
Xbit_r442_c39 bl[39] br[39] wl[442] vdd gnd cell_6t
Xbit_r443_c39 bl[39] br[39] wl[443] vdd gnd cell_6t
Xbit_r444_c39 bl[39] br[39] wl[444] vdd gnd cell_6t
Xbit_r445_c39 bl[39] br[39] wl[445] vdd gnd cell_6t
Xbit_r446_c39 bl[39] br[39] wl[446] vdd gnd cell_6t
Xbit_r447_c39 bl[39] br[39] wl[447] vdd gnd cell_6t
Xbit_r448_c39 bl[39] br[39] wl[448] vdd gnd cell_6t
Xbit_r449_c39 bl[39] br[39] wl[449] vdd gnd cell_6t
Xbit_r450_c39 bl[39] br[39] wl[450] vdd gnd cell_6t
Xbit_r451_c39 bl[39] br[39] wl[451] vdd gnd cell_6t
Xbit_r452_c39 bl[39] br[39] wl[452] vdd gnd cell_6t
Xbit_r453_c39 bl[39] br[39] wl[453] vdd gnd cell_6t
Xbit_r454_c39 bl[39] br[39] wl[454] vdd gnd cell_6t
Xbit_r455_c39 bl[39] br[39] wl[455] vdd gnd cell_6t
Xbit_r456_c39 bl[39] br[39] wl[456] vdd gnd cell_6t
Xbit_r457_c39 bl[39] br[39] wl[457] vdd gnd cell_6t
Xbit_r458_c39 bl[39] br[39] wl[458] vdd gnd cell_6t
Xbit_r459_c39 bl[39] br[39] wl[459] vdd gnd cell_6t
Xbit_r460_c39 bl[39] br[39] wl[460] vdd gnd cell_6t
Xbit_r461_c39 bl[39] br[39] wl[461] vdd gnd cell_6t
Xbit_r462_c39 bl[39] br[39] wl[462] vdd gnd cell_6t
Xbit_r463_c39 bl[39] br[39] wl[463] vdd gnd cell_6t
Xbit_r464_c39 bl[39] br[39] wl[464] vdd gnd cell_6t
Xbit_r465_c39 bl[39] br[39] wl[465] vdd gnd cell_6t
Xbit_r466_c39 bl[39] br[39] wl[466] vdd gnd cell_6t
Xbit_r467_c39 bl[39] br[39] wl[467] vdd gnd cell_6t
Xbit_r468_c39 bl[39] br[39] wl[468] vdd gnd cell_6t
Xbit_r469_c39 bl[39] br[39] wl[469] vdd gnd cell_6t
Xbit_r470_c39 bl[39] br[39] wl[470] vdd gnd cell_6t
Xbit_r471_c39 bl[39] br[39] wl[471] vdd gnd cell_6t
Xbit_r472_c39 bl[39] br[39] wl[472] vdd gnd cell_6t
Xbit_r473_c39 bl[39] br[39] wl[473] vdd gnd cell_6t
Xbit_r474_c39 bl[39] br[39] wl[474] vdd gnd cell_6t
Xbit_r475_c39 bl[39] br[39] wl[475] vdd gnd cell_6t
Xbit_r476_c39 bl[39] br[39] wl[476] vdd gnd cell_6t
Xbit_r477_c39 bl[39] br[39] wl[477] vdd gnd cell_6t
Xbit_r478_c39 bl[39] br[39] wl[478] vdd gnd cell_6t
Xbit_r479_c39 bl[39] br[39] wl[479] vdd gnd cell_6t
Xbit_r480_c39 bl[39] br[39] wl[480] vdd gnd cell_6t
Xbit_r481_c39 bl[39] br[39] wl[481] vdd gnd cell_6t
Xbit_r482_c39 bl[39] br[39] wl[482] vdd gnd cell_6t
Xbit_r483_c39 bl[39] br[39] wl[483] vdd gnd cell_6t
Xbit_r484_c39 bl[39] br[39] wl[484] vdd gnd cell_6t
Xbit_r485_c39 bl[39] br[39] wl[485] vdd gnd cell_6t
Xbit_r486_c39 bl[39] br[39] wl[486] vdd gnd cell_6t
Xbit_r487_c39 bl[39] br[39] wl[487] vdd gnd cell_6t
Xbit_r488_c39 bl[39] br[39] wl[488] vdd gnd cell_6t
Xbit_r489_c39 bl[39] br[39] wl[489] vdd gnd cell_6t
Xbit_r490_c39 bl[39] br[39] wl[490] vdd gnd cell_6t
Xbit_r491_c39 bl[39] br[39] wl[491] vdd gnd cell_6t
Xbit_r492_c39 bl[39] br[39] wl[492] vdd gnd cell_6t
Xbit_r493_c39 bl[39] br[39] wl[493] vdd gnd cell_6t
Xbit_r494_c39 bl[39] br[39] wl[494] vdd gnd cell_6t
Xbit_r495_c39 bl[39] br[39] wl[495] vdd gnd cell_6t
Xbit_r496_c39 bl[39] br[39] wl[496] vdd gnd cell_6t
Xbit_r497_c39 bl[39] br[39] wl[497] vdd gnd cell_6t
Xbit_r498_c39 bl[39] br[39] wl[498] vdd gnd cell_6t
Xbit_r499_c39 bl[39] br[39] wl[499] vdd gnd cell_6t
Xbit_r500_c39 bl[39] br[39] wl[500] vdd gnd cell_6t
Xbit_r501_c39 bl[39] br[39] wl[501] vdd gnd cell_6t
Xbit_r502_c39 bl[39] br[39] wl[502] vdd gnd cell_6t
Xbit_r503_c39 bl[39] br[39] wl[503] vdd gnd cell_6t
Xbit_r504_c39 bl[39] br[39] wl[504] vdd gnd cell_6t
Xbit_r505_c39 bl[39] br[39] wl[505] vdd gnd cell_6t
Xbit_r506_c39 bl[39] br[39] wl[506] vdd gnd cell_6t
Xbit_r507_c39 bl[39] br[39] wl[507] vdd gnd cell_6t
Xbit_r508_c39 bl[39] br[39] wl[508] vdd gnd cell_6t
Xbit_r509_c39 bl[39] br[39] wl[509] vdd gnd cell_6t
Xbit_r510_c39 bl[39] br[39] wl[510] vdd gnd cell_6t
Xbit_r511_c39 bl[39] br[39] wl[511] vdd gnd cell_6t
Xbit_r0_c40 bl[40] br[40] wl[0] vdd gnd cell_6t
Xbit_r1_c40 bl[40] br[40] wl[1] vdd gnd cell_6t
Xbit_r2_c40 bl[40] br[40] wl[2] vdd gnd cell_6t
Xbit_r3_c40 bl[40] br[40] wl[3] vdd gnd cell_6t
Xbit_r4_c40 bl[40] br[40] wl[4] vdd gnd cell_6t
Xbit_r5_c40 bl[40] br[40] wl[5] vdd gnd cell_6t
Xbit_r6_c40 bl[40] br[40] wl[6] vdd gnd cell_6t
Xbit_r7_c40 bl[40] br[40] wl[7] vdd gnd cell_6t
Xbit_r8_c40 bl[40] br[40] wl[8] vdd gnd cell_6t
Xbit_r9_c40 bl[40] br[40] wl[9] vdd gnd cell_6t
Xbit_r10_c40 bl[40] br[40] wl[10] vdd gnd cell_6t
Xbit_r11_c40 bl[40] br[40] wl[11] vdd gnd cell_6t
Xbit_r12_c40 bl[40] br[40] wl[12] vdd gnd cell_6t
Xbit_r13_c40 bl[40] br[40] wl[13] vdd gnd cell_6t
Xbit_r14_c40 bl[40] br[40] wl[14] vdd gnd cell_6t
Xbit_r15_c40 bl[40] br[40] wl[15] vdd gnd cell_6t
Xbit_r16_c40 bl[40] br[40] wl[16] vdd gnd cell_6t
Xbit_r17_c40 bl[40] br[40] wl[17] vdd gnd cell_6t
Xbit_r18_c40 bl[40] br[40] wl[18] vdd gnd cell_6t
Xbit_r19_c40 bl[40] br[40] wl[19] vdd gnd cell_6t
Xbit_r20_c40 bl[40] br[40] wl[20] vdd gnd cell_6t
Xbit_r21_c40 bl[40] br[40] wl[21] vdd gnd cell_6t
Xbit_r22_c40 bl[40] br[40] wl[22] vdd gnd cell_6t
Xbit_r23_c40 bl[40] br[40] wl[23] vdd gnd cell_6t
Xbit_r24_c40 bl[40] br[40] wl[24] vdd gnd cell_6t
Xbit_r25_c40 bl[40] br[40] wl[25] vdd gnd cell_6t
Xbit_r26_c40 bl[40] br[40] wl[26] vdd gnd cell_6t
Xbit_r27_c40 bl[40] br[40] wl[27] vdd gnd cell_6t
Xbit_r28_c40 bl[40] br[40] wl[28] vdd gnd cell_6t
Xbit_r29_c40 bl[40] br[40] wl[29] vdd gnd cell_6t
Xbit_r30_c40 bl[40] br[40] wl[30] vdd gnd cell_6t
Xbit_r31_c40 bl[40] br[40] wl[31] vdd gnd cell_6t
Xbit_r32_c40 bl[40] br[40] wl[32] vdd gnd cell_6t
Xbit_r33_c40 bl[40] br[40] wl[33] vdd gnd cell_6t
Xbit_r34_c40 bl[40] br[40] wl[34] vdd gnd cell_6t
Xbit_r35_c40 bl[40] br[40] wl[35] vdd gnd cell_6t
Xbit_r36_c40 bl[40] br[40] wl[36] vdd gnd cell_6t
Xbit_r37_c40 bl[40] br[40] wl[37] vdd gnd cell_6t
Xbit_r38_c40 bl[40] br[40] wl[38] vdd gnd cell_6t
Xbit_r39_c40 bl[40] br[40] wl[39] vdd gnd cell_6t
Xbit_r40_c40 bl[40] br[40] wl[40] vdd gnd cell_6t
Xbit_r41_c40 bl[40] br[40] wl[41] vdd gnd cell_6t
Xbit_r42_c40 bl[40] br[40] wl[42] vdd gnd cell_6t
Xbit_r43_c40 bl[40] br[40] wl[43] vdd gnd cell_6t
Xbit_r44_c40 bl[40] br[40] wl[44] vdd gnd cell_6t
Xbit_r45_c40 bl[40] br[40] wl[45] vdd gnd cell_6t
Xbit_r46_c40 bl[40] br[40] wl[46] vdd gnd cell_6t
Xbit_r47_c40 bl[40] br[40] wl[47] vdd gnd cell_6t
Xbit_r48_c40 bl[40] br[40] wl[48] vdd gnd cell_6t
Xbit_r49_c40 bl[40] br[40] wl[49] vdd gnd cell_6t
Xbit_r50_c40 bl[40] br[40] wl[50] vdd gnd cell_6t
Xbit_r51_c40 bl[40] br[40] wl[51] vdd gnd cell_6t
Xbit_r52_c40 bl[40] br[40] wl[52] vdd gnd cell_6t
Xbit_r53_c40 bl[40] br[40] wl[53] vdd gnd cell_6t
Xbit_r54_c40 bl[40] br[40] wl[54] vdd gnd cell_6t
Xbit_r55_c40 bl[40] br[40] wl[55] vdd gnd cell_6t
Xbit_r56_c40 bl[40] br[40] wl[56] vdd gnd cell_6t
Xbit_r57_c40 bl[40] br[40] wl[57] vdd gnd cell_6t
Xbit_r58_c40 bl[40] br[40] wl[58] vdd gnd cell_6t
Xbit_r59_c40 bl[40] br[40] wl[59] vdd gnd cell_6t
Xbit_r60_c40 bl[40] br[40] wl[60] vdd gnd cell_6t
Xbit_r61_c40 bl[40] br[40] wl[61] vdd gnd cell_6t
Xbit_r62_c40 bl[40] br[40] wl[62] vdd gnd cell_6t
Xbit_r63_c40 bl[40] br[40] wl[63] vdd gnd cell_6t
Xbit_r64_c40 bl[40] br[40] wl[64] vdd gnd cell_6t
Xbit_r65_c40 bl[40] br[40] wl[65] vdd gnd cell_6t
Xbit_r66_c40 bl[40] br[40] wl[66] vdd gnd cell_6t
Xbit_r67_c40 bl[40] br[40] wl[67] vdd gnd cell_6t
Xbit_r68_c40 bl[40] br[40] wl[68] vdd gnd cell_6t
Xbit_r69_c40 bl[40] br[40] wl[69] vdd gnd cell_6t
Xbit_r70_c40 bl[40] br[40] wl[70] vdd gnd cell_6t
Xbit_r71_c40 bl[40] br[40] wl[71] vdd gnd cell_6t
Xbit_r72_c40 bl[40] br[40] wl[72] vdd gnd cell_6t
Xbit_r73_c40 bl[40] br[40] wl[73] vdd gnd cell_6t
Xbit_r74_c40 bl[40] br[40] wl[74] vdd gnd cell_6t
Xbit_r75_c40 bl[40] br[40] wl[75] vdd gnd cell_6t
Xbit_r76_c40 bl[40] br[40] wl[76] vdd gnd cell_6t
Xbit_r77_c40 bl[40] br[40] wl[77] vdd gnd cell_6t
Xbit_r78_c40 bl[40] br[40] wl[78] vdd gnd cell_6t
Xbit_r79_c40 bl[40] br[40] wl[79] vdd gnd cell_6t
Xbit_r80_c40 bl[40] br[40] wl[80] vdd gnd cell_6t
Xbit_r81_c40 bl[40] br[40] wl[81] vdd gnd cell_6t
Xbit_r82_c40 bl[40] br[40] wl[82] vdd gnd cell_6t
Xbit_r83_c40 bl[40] br[40] wl[83] vdd gnd cell_6t
Xbit_r84_c40 bl[40] br[40] wl[84] vdd gnd cell_6t
Xbit_r85_c40 bl[40] br[40] wl[85] vdd gnd cell_6t
Xbit_r86_c40 bl[40] br[40] wl[86] vdd gnd cell_6t
Xbit_r87_c40 bl[40] br[40] wl[87] vdd gnd cell_6t
Xbit_r88_c40 bl[40] br[40] wl[88] vdd gnd cell_6t
Xbit_r89_c40 bl[40] br[40] wl[89] vdd gnd cell_6t
Xbit_r90_c40 bl[40] br[40] wl[90] vdd gnd cell_6t
Xbit_r91_c40 bl[40] br[40] wl[91] vdd gnd cell_6t
Xbit_r92_c40 bl[40] br[40] wl[92] vdd gnd cell_6t
Xbit_r93_c40 bl[40] br[40] wl[93] vdd gnd cell_6t
Xbit_r94_c40 bl[40] br[40] wl[94] vdd gnd cell_6t
Xbit_r95_c40 bl[40] br[40] wl[95] vdd gnd cell_6t
Xbit_r96_c40 bl[40] br[40] wl[96] vdd gnd cell_6t
Xbit_r97_c40 bl[40] br[40] wl[97] vdd gnd cell_6t
Xbit_r98_c40 bl[40] br[40] wl[98] vdd gnd cell_6t
Xbit_r99_c40 bl[40] br[40] wl[99] vdd gnd cell_6t
Xbit_r100_c40 bl[40] br[40] wl[100] vdd gnd cell_6t
Xbit_r101_c40 bl[40] br[40] wl[101] vdd gnd cell_6t
Xbit_r102_c40 bl[40] br[40] wl[102] vdd gnd cell_6t
Xbit_r103_c40 bl[40] br[40] wl[103] vdd gnd cell_6t
Xbit_r104_c40 bl[40] br[40] wl[104] vdd gnd cell_6t
Xbit_r105_c40 bl[40] br[40] wl[105] vdd gnd cell_6t
Xbit_r106_c40 bl[40] br[40] wl[106] vdd gnd cell_6t
Xbit_r107_c40 bl[40] br[40] wl[107] vdd gnd cell_6t
Xbit_r108_c40 bl[40] br[40] wl[108] vdd gnd cell_6t
Xbit_r109_c40 bl[40] br[40] wl[109] vdd gnd cell_6t
Xbit_r110_c40 bl[40] br[40] wl[110] vdd gnd cell_6t
Xbit_r111_c40 bl[40] br[40] wl[111] vdd gnd cell_6t
Xbit_r112_c40 bl[40] br[40] wl[112] vdd gnd cell_6t
Xbit_r113_c40 bl[40] br[40] wl[113] vdd gnd cell_6t
Xbit_r114_c40 bl[40] br[40] wl[114] vdd gnd cell_6t
Xbit_r115_c40 bl[40] br[40] wl[115] vdd gnd cell_6t
Xbit_r116_c40 bl[40] br[40] wl[116] vdd gnd cell_6t
Xbit_r117_c40 bl[40] br[40] wl[117] vdd gnd cell_6t
Xbit_r118_c40 bl[40] br[40] wl[118] vdd gnd cell_6t
Xbit_r119_c40 bl[40] br[40] wl[119] vdd gnd cell_6t
Xbit_r120_c40 bl[40] br[40] wl[120] vdd gnd cell_6t
Xbit_r121_c40 bl[40] br[40] wl[121] vdd gnd cell_6t
Xbit_r122_c40 bl[40] br[40] wl[122] vdd gnd cell_6t
Xbit_r123_c40 bl[40] br[40] wl[123] vdd gnd cell_6t
Xbit_r124_c40 bl[40] br[40] wl[124] vdd gnd cell_6t
Xbit_r125_c40 bl[40] br[40] wl[125] vdd gnd cell_6t
Xbit_r126_c40 bl[40] br[40] wl[126] vdd gnd cell_6t
Xbit_r127_c40 bl[40] br[40] wl[127] vdd gnd cell_6t
Xbit_r128_c40 bl[40] br[40] wl[128] vdd gnd cell_6t
Xbit_r129_c40 bl[40] br[40] wl[129] vdd gnd cell_6t
Xbit_r130_c40 bl[40] br[40] wl[130] vdd gnd cell_6t
Xbit_r131_c40 bl[40] br[40] wl[131] vdd gnd cell_6t
Xbit_r132_c40 bl[40] br[40] wl[132] vdd gnd cell_6t
Xbit_r133_c40 bl[40] br[40] wl[133] vdd gnd cell_6t
Xbit_r134_c40 bl[40] br[40] wl[134] vdd gnd cell_6t
Xbit_r135_c40 bl[40] br[40] wl[135] vdd gnd cell_6t
Xbit_r136_c40 bl[40] br[40] wl[136] vdd gnd cell_6t
Xbit_r137_c40 bl[40] br[40] wl[137] vdd gnd cell_6t
Xbit_r138_c40 bl[40] br[40] wl[138] vdd gnd cell_6t
Xbit_r139_c40 bl[40] br[40] wl[139] vdd gnd cell_6t
Xbit_r140_c40 bl[40] br[40] wl[140] vdd gnd cell_6t
Xbit_r141_c40 bl[40] br[40] wl[141] vdd gnd cell_6t
Xbit_r142_c40 bl[40] br[40] wl[142] vdd gnd cell_6t
Xbit_r143_c40 bl[40] br[40] wl[143] vdd gnd cell_6t
Xbit_r144_c40 bl[40] br[40] wl[144] vdd gnd cell_6t
Xbit_r145_c40 bl[40] br[40] wl[145] vdd gnd cell_6t
Xbit_r146_c40 bl[40] br[40] wl[146] vdd gnd cell_6t
Xbit_r147_c40 bl[40] br[40] wl[147] vdd gnd cell_6t
Xbit_r148_c40 bl[40] br[40] wl[148] vdd gnd cell_6t
Xbit_r149_c40 bl[40] br[40] wl[149] vdd gnd cell_6t
Xbit_r150_c40 bl[40] br[40] wl[150] vdd gnd cell_6t
Xbit_r151_c40 bl[40] br[40] wl[151] vdd gnd cell_6t
Xbit_r152_c40 bl[40] br[40] wl[152] vdd gnd cell_6t
Xbit_r153_c40 bl[40] br[40] wl[153] vdd gnd cell_6t
Xbit_r154_c40 bl[40] br[40] wl[154] vdd gnd cell_6t
Xbit_r155_c40 bl[40] br[40] wl[155] vdd gnd cell_6t
Xbit_r156_c40 bl[40] br[40] wl[156] vdd gnd cell_6t
Xbit_r157_c40 bl[40] br[40] wl[157] vdd gnd cell_6t
Xbit_r158_c40 bl[40] br[40] wl[158] vdd gnd cell_6t
Xbit_r159_c40 bl[40] br[40] wl[159] vdd gnd cell_6t
Xbit_r160_c40 bl[40] br[40] wl[160] vdd gnd cell_6t
Xbit_r161_c40 bl[40] br[40] wl[161] vdd gnd cell_6t
Xbit_r162_c40 bl[40] br[40] wl[162] vdd gnd cell_6t
Xbit_r163_c40 bl[40] br[40] wl[163] vdd gnd cell_6t
Xbit_r164_c40 bl[40] br[40] wl[164] vdd gnd cell_6t
Xbit_r165_c40 bl[40] br[40] wl[165] vdd gnd cell_6t
Xbit_r166_c40 bl[40] br[40] wl[166] vdd gnd cell_6t
Xbit_r167_c40 bl[40] br[40] wl[167] vdd gnd cell_6t
Xbit_r168_c40 bl[40] br[40] wl[168] vdd gnd cell_6t
Xbit_r169_c40 bl[40] br[40] wl[169] vdd gnd cell_6t
Xbit_r170_c40 bl[40] br[40] wl[170] vdd gnd cell_6t
Xbit_r171_c40 bl[40] br[40] wl[171] vdd gnd cell_6t
Xbit_r172_c40 bl[40] br[40] wl[172] vdd gnd cell_6t
Xbit_r173_c40 bl[40] br[40] wl[173] vdd gnd cell_6t
Xbit_r174_c40 bl[40] br[40] wl[174] vdd gnd cell_6t
Xbit_r175_c40 bl[40] br[40] wl[175] vdd gnd cell_6t
Xbit_r176_c40 bl[40] br[40] wl[176] vdd gnd cell_6t
Xbit_r177_c40 bl[40] br[40] wl[177] vdd gnd cell_6t
Xbit_r178_c40 bl[40] br[40] wl[178] vdd gnd cell_6t
Xbit_r179_c40 bl[40] br[40] wl[179] vdd gnd cell_6t
Xbit_r180_c40 bl[40] br[40] wl[180] vdd gnd cell_6t
Xbit_r181_c40 bl[40] br[40] wl[181] vdd gnd cell_6t
Xbit_r182_c40 bl[40] br[40] wl[182] vdd gnd cell_6t
Xbit_r183_c40 bl[40] br[40] wl[183] vdd gnd cell_6t
Xbit_r184_c40 bl[40] br[40] wl[184] vdd gnd cell_6t
Xbit_r185_c40 bl[40] br[40] wl[185] vdd gnd cell_6t
Xbit_r186_c40 bl[40] br[40] wl[186] vdd gnd cell_6t
Xbit_r187_c40 bl[40] br[40] wl[187] vdd gnd cell_6t
Xbit_r188_c40 bl[40] br[40] wl[188] vdd gnd cell_6t
Xbit_r189_c40 bl[40] br[40] wl[189] vdd gnd cell_6t
Xbit_r190_c40 bl[40] br[40] wl[190] vdd gnd cell_6t
Xbit_r191_c40 bl[40] br[40] wl[191] vdd gnd cell_6t
Xbit_r192_c40 bl[40] br[40] wl[192] vdd gnd cell_6t
Xbit_r193_c40 bl[40] br[40] wl[193] vdd gnd cell_6t
Xbit_r194_c40 bl[40] br[40] wl[194] vdd gnd cell_6t
Xbit_r195_c40 bl[40] br[40] wl[195] vdd gnd cell_6t
Xbit_r196_c40 bl[40] br[40] wl[196] vdd gnd cell_6t
Xbit_r197_c40 bl[40] br[40] wl[197] vdd gnd cell_6t
Xbit_r198_c40 bl[40] br[40] wl[198] vdd gnd cell_6t
Xbit_r199_c40 bl[40] br[40] wl[199] vdd gnd cell_6t
Xbit_r200_c40 bl[40] br[40] wl[200] vdd gnd cell_6t
Xbit_r201_c40 bl[40] br[40] wl[201] vdd gnd cell_6t
Xbit_r202_c40 bl[40] br[40] wl[202] vdd gnd cell_6t
Xbit_r203_c40 bl[40] br[40] wl[203] vdd gnd cell_6t
Xbit_r204_c40 bl[40] br[40] wl[204] vdd gnd cell_6t
Xbit_r205_c40 bl[40] br[40] wl[205] vdd gnd cell_6t
Xbit_r206_c40 bl[40] br[40] wl[206] vdd gnd cell_6t
Xbit_r207_c40 bl[40] br[40] wl[207] vdd gnd cell_6t
Xbit_r208_c40 bl[40] br[40] wl[208] vdd gnd cell_6t
Xbit_r209_c40 bl[40] br[40] wl[209] vdd gnd cell_6t
Xbit_r210_c40 bl[40] br[40] wl[210] vdd gnd cell_6t
Xbit_r211_c40 bl[40] br[40] wl[211] vdd gnd cell_6t
Xbit_r212_c40 bl[40] br[40] wl[212] vdd gnd cell_6t
Xbit_r213_c40 bl[40] br[40] wl[213] vdd gnd cell_6t
Xbit_r214_c40 bl[40] br[40] wl[214] vdd gnd cell_6t
Xbit_r215_c40 bl[40] br[40] wl[215] vdd gnd cell_6t
Xbit_r216_c40 bl[40] br[40] wl[216] vdd gnd cell_6t
Xbit_r217_c40 bl[40] br[40] wl[217] vdd gnd cell_6t
Xbit_r218_c40 bl[40] br[40] wl[218] vdd gnd cell_6t
Xbit_r219_c40 bl[40] br[40] wl[219] vdd gnd cell_6t
Xbit_r220_c40 bl[40] br[40] wl[220] vdd gnd cell_6t
Xbit_r221_c40 bl[40] br[40] wl[221] vdd gnd cell_6t
Xbit_r222_c40 bl[40] br[40] wl[222] vdd gnd cell_6t
Xbit_r223_c40 bl[40] br[40] wl[223] vdd gnd cell_6t
Xbit_r224_c40 bl[40] br[40] wl[224] vdd gnd cell_6t
Xbit_r225_c40 bl[40] br[40] wl[225] vdd gnd cell_6t
Xbit_r226_c40 bl[40] br[40] wl[226] vdd gnd cell_6t
Xbit_r227_c40 bl[40] br[40] wl[227] vdd gnd cell_6t
Xbit_r228_c40 bl[40] br[40] wl[228] vdd gnd cell_6t
Xbit_r229_c40 bl[40] br[40] wl[229] vdd gnd cell_6t
Xbit_r230_c40 bl[40] br[40] wl[230] vdd gnd cell_6t
Xbit_r231_c40 bl[40] br[40] wl[231] vdd gnd cell_6t
Xbit_r232_c40 bl[40] br[40] wl[232] vdd gnd cell_6t
Xbit_r233_c40 bl[40] br[40] wl[233] vdd gnd cell_6t
Xbit_r234_c40 bl[40] br[40] wl[234] vdd gnd cell_6t
Xbit_r235_c40 bl[40] br[40] wl[235] vdd gnd cell_6t
Xbit_r236_c40 bl[40] br[40] wl[236] vdd gnd cell_6t
Xbit_r237_c40 bl[40] br[40] wl[237] vdd gnd cell_6t
Xbit_r238_c40 bl[40] br[40] wl[238] vdd gnd cell_6t
Xbit_r239_c40 bl[40] br[40] wl[239] vdd gnd cell_6t
Xbit_r240_c40 bl[40] br[40] wl[240] vdd gnd cell_6t
Xbit_r241_c40 bl[40] br[40] wl[241] vdd gnd cell_6t
Xbit_r242_c40 bl[40] br[40] wl[242] vdd gnd cell_6t
Xbit_r243_c40 bl[40] br[40] wl[243] vdd gnd cell_6t
Xbit_r244_c40 bl[40] br[40] wl[244] vdd gnd cell_6t
Xbit_r245_c40 bl[40] br[40] wl[245] vdd gnd cell_6t
Xbit_r246_c40 bl[40] br[40] wl[246] vdd gnd cell_6t
Xbit_r247_c40 bl[40] br[40] wl[247] vdd gnd cell_6t
Xbit_r248_c40 bl[40] br[40] wl[248] vdd gnd cell_6t
Xbit_r249_c40 bl[40] br[40] wl[249] vdd gnd cell_6t
Xbit_r250_c40 bl[40] br[40] wl[250] vdd gnd cell_6t
Xbit_r251_c40 bl[40] br[40] wl[251] vdd gnd cell_6t
Xbit_r252_c40 bl[40] br[40] wl[252] vdd gnd cell_6t
Xbit_r253_c40 bl[40] br[40] wl[253] vdd gnd cell_6t
Xbit_r254_c40 bl[40] br[40] wl[254] vdd gnd cell_6t
Xbit_r255_c40 bl[40] br[40] wl[255] vdd gnd cell_6t
Xbit_r256_c40 bl[40] br[40] wl[256] vdd gnd cell_6t
Xbit_r257_c40 bl[40] br[40] wl[257] vdd gnd cell_6t
Xbit_r258_c40 bl[40] br[40] wl[258] vdd gnd cell_6t
Xbit_r259_c40 bl[40] br[40] wl[259] vdd gnd cell_6t
Xbit_r260_c40 bl[40] br[40] wl[260] vdd gnd cell_6t
Xbit_r261_c40 bl[40] br[40] wl[261] vdd gnd cell_6t
Xbit_r262_c40 bl[40] br[40] wl[262] vdd gnd cell_6t
Xbit_r263_c40 bl[40] br[40] wl[263] vdd gnd cell_6t
Xbit_r264_c40 bl[40] br[40] wl[264] vdd gnd cell_6t
Xbit_r265_c40 bl[40] br[40] wl[265] vdd gnd cell_6t
Xbit_r266_c40 bl[40] br[40] wl[266] vdd gnd cell_6t
Xbit_r267_c40 bl[40] br[40] wl[267] vdd gnd cell_6t
Xbit_r268_c40 bl[40] br[40] wl[268] vdd gnd cell_6t
Xbit_r269_c40 bl[40] br[40] wl[269] vdd gnd cell_6t
Xbit_r270_c40 bl[40] br[40] wl[270] vdd gnd cell_6t
Xbit_r271_c40 bl[40] br[40] wl[271] vdd gnd cell_6t
Xbit_r272_c40 bl[40] br[40] wl[272] vdd gnd cell_6t
Xbit_r273_c40 bl[40] br[40] wl[273] vdd gnd cell_6t
Xbit_r274_c40 bl[40] br[40] wl[274] vdd gnd cell_6t
Xbit_r275_c40 bl[40] br[40] wl[275] vdd gnd cell_6t
Xbit_r276_c40 bl[40] br[40] wl[276] vdd gnd cell_6t
Xbit_r277_c40 bl[40] br[40] wl[277] vdd gnd cell_6t
Xbit_r278_c40 bl[40] br[40] wl[278] vdd gnd cell_6t
Xbit_r279_c40 bl[40] br[40] wl[279] vdd gnd cell_6t
Xbit_r280_c40 bl[40] br[40] wl[280] vdd gnd cell_6t
Xbit_r281_c40 bl[40] br[40] wl[281] vdd gnd cell_6t
Xbit_r282_c40 bl[40] br[40] wl[282] vdd gnd cell_6t
Xbit_r283_c40 bl[40] br[40] wl[283] vdd gnd cell_6t
Xbit_r284_c40 bl[40] br[40] wl[284] vdd gnd cell_6t
Xbit_r285_c40 bl[40] br[40] wl[285] vdd gnd cell_6t
Xbit_r286_c40 bl[40] br[40] wl[286] vdd gnd cell_6t
Xbit_r287_c40 bl[40] br[40] wl[287] vdd gnd cell_6t
Xbit_r288_c40 bl[40] br[40] wl[288] vdd gnd cell_6t
Xbit_r289_c40 bl[40] br[40] wl[289] vdd gnd cell_6t
Xbit_r290_c40 bl[40] br[40] wl[290] vdd gnd cell_6t
Xbit_r291_c40 bl[40] br[40] wl[291] vdd gnd cell_6t
Xbit_r292_c40 bl[40] br[40] wl[292] vdd gnd cell_6t
Xbit_r293_c40 bl[40] br[40] wl[293] vdd gnd cell_6t
Xbit_r294_c40 bl[40] br[40] wl[294] vdd gnd cell_6t
Xbit_r295_c40 bl[40] br[40] wl[295] vdd gnd cell_6t
Xbit_r296_c40 bl[40] br[40] wl[296] vdd gnd cell_6t
Xbit_r297_c40 bl[40] br[40] wl[297] vdd gnd cell_6t
Xbit_r298_c40 bl[40] br[40] wl[298] vdd gnd cell_6t
Xbit_r299_c40 bl[40] br[40] wl[299] vdd gnd cell_6t
Xbit_r300_c40 bl[40] br[40] wl[300] vdd gnd cell_6t
Xbit_r301_c40 bl[40] br[40] wl[301] vdd gnd cell_6t
Xbit_r302_c40 bl[40] br[40] wl[302] vdd gnd cell_6t
Xbit_r303_c40 bl[40] br[40] wl[303] vdd gnd cell_6t
Xbit_r304_c40 bl[40] br[40] wl[304] vdd gnd cell_6t
Xbit_r305_c40 bl[40] br[40] wl[305] vdd gnd cell_6t
Xbit_r306_c40 bl[40] br[40] wl[306] vdd gnd cell_6t
Xbit_r307_c40 bl[40] br[40] wl[307] vdd gnd cell_6t
Xbit_r308_c40 bl[40] br[40] wl[308] vdd gnd cell_6t
Xbit_r309_c40 bl[40] br[40] wl[309] vdd gnd cell_6t
Xbit_r310_c40 bl[40] br[40] wl[310] vdd gnd cell_6t
Xbit_r311_c40 bl[40] br[40] wl[311] vdd gnd cell_6t
Xbit_r312_c40 bl[40] br[40] wl[312] vdd gnd cell_6t
Xbit_r313_c40 bl[40] br[40] wl[313] vdd gnd cell_6t
Xbit_r314_c40 bl[40] br[40] wl[314] vdd gnd cell_6t
Xbit_r315_c40 bl[40] br[40] wl[315] vdd gnd cell_6t
Xbit_r316_c40 bl[40] br[40] wl[316] vdd gnd cell_6t
Xbit_r317_c40 bl[40] br[40] wl[317] vdd gnd cell_6t
Xbit_r318_c40 bl[40] br[40] wl[318] vdd gnd cell_6t
Xbit_r319_c40 bl[40] br[40] wl[319] vdd gnd cell_6t
Xbit_r320_c40 bl[40] br[40] wl[320] vdd gnd cell_6t
Xbit_r321_c40 bl[40] br[40] wl[321] vdd gnd cell_6t
Xbit_r322_c40 bl[40] br[40] wl[322] vdd gnd cell_6t
Xbit_r323_c40 bl[40] br[40] wl[323] vdd gnd cell_6t
Xbit_r324_c40 bl[40] br[40] wl[324] vdd gnd cell_6t
Xbit_r325_c40 bl[40] br[40] wl[325] vdd gnd cell_6t
Xbit_r326_c40 bl[40] br[40] wl[326] vdd gnd cell_6t
Xbit_r327_c40 bl[40] br[40] wl[327] vdd gnd cell_6t
Xbit_r328_c40 bl[40] br[40] wl[328] vdd gnd cell_6t
Xbit_r329_c40 bl[40] br[40] wl[329] vdd gnd cell_6t
Xbit_r330_c40 bl[40] br[40] wl[330] vdd gnd cell_6t
Xbit_r331_c40 bl[40] br[40] wl[331] vdd gnd cell_6t
Xbit_r332_c40 bl[40] br[40] wl[332] vdd gnd cell_6t
Xbit_r333_c40 bl[40] br[40] wl[333] vdd gnd cell_6t
Xbit_r334_c40 bl[40] br[40] wl[334] vdd gnd cell_6t
Xbit_r335_c40 bl[40] br[40] wl[335] vdd gnd cell_6t
Xbit_r336_c40 bl[40] br[40] wl[336] vdd gnd cell_6t
Xbit_r337_c40 bl[40] br[40] wl[337] vdd gnd cell_6t
Xbit_r338_c40 bl[40] br[40] wl[338] vdd gnd cell_6t
Xbit_r339_c40 bl[40] br[40] wl[339] vdd gnd cell_6t
Xbit_r340_c40 bl[40] br[40] wl[340] vdd gnd cell_6t
Xbit_r341_c40 bl[40] br[40] wl[341] vdd gnd cell_6t
Xbit_r342_c40 bl[40] br[40] wl[342] vdd gnd cell_6t
Xbit_r343_c40 bl[40] br[40] wl[343] vdd gnd cell_6t
Xbit_r344_c40 bl[40] br[40] wl[344] vdd gnd cell_6t
Xbit_r345_c40 bl[40] br[40] wl[345] vdd gnd cell_6t
Xbit_r346_c40 bl[40] br[40] wl[346] vdd gnd cell_6t
Xbit_r347_c40 bl[40] br[40] wl[347] vdd gnd cell_6t
Xbit_r348_c40 bl[40] br[40] wl[348] vdd gnd cell_6t
Xbit_r349_c40 bl[40] br[40] wl[349] vdd gnd cell_6t
Xbit_r350_c40 bl[40] br[40] wl[350] vdd gnd cell_6t
Xbit_r351_c40 bl[40] br[40] wl[351] vdd gnd cell_6t
Xbit_r352_c40 bl[40] br[40] wl[352] vdd gnd cell_6t
Xbit_r353_c40 bl[40] br[40] wl[353] vdd gnd cell_6t
Xbit_r354_c40 bl[40] br[40] wl[354] vdd gnd cell_6t
Xbit_r355_c40 bl[40] br[40] wl[355] vdd gnd cell_6t
Xbit_r356_c40 bl[40] br[40] wl[356] vdd gnd cell_6t
Xbit_r357_c40 bl[40] br[40] wl[357] vdd gnd cell_6t
Xbit_r358_c40 bl[40] br[40] wl[358] vdd gnd cell_6t
Xbit_r359_c40 bl[40] br[40] wl[359] vdd gnd cell_6t
Xbit_r360_c40 bl[40] br[40] wl[360] vdd gnd cell_6t
Xbit_r361_c40 bl[40] br[40] wl[361] vdd gnd cell_6t
Xbit_r362_c40 bl[40] br[40] wl[362] vdd gnd cell_6t
Xbit_r363_c40 bl[40] br[40] wl[363] vdd gnd cell_6t
Xbit_r364_c40 bl[40] br[40] wl[364] vdd gnd cell_6t
Xbit_r365_c40 bl[40] br[40] wl[365] vdd gnd cell_6t
Xbit_r366_c40 bl[40] br[40] wl[366] vdd gnd cell_6t
Xbit_r367_c40 bl[40] br[40] wl[367] vdd gnd cell_6t
Xbit_r368_c40 bl[40] br[40] wl[368] vdd gnd cell_6t
Xbit_r369_c40 bl[40] br[40] wl[369] vdd gnd cell_6t
Xbit_r370_c40 bl[40] br[40] wl[370] vdd gnd cell_6t
Xbit_r371_c40 bl[40] br[40] wl[371] vdd gnd cell_6t
Xbit_r372_c40 bl[40] br[40] wl[372] vdd gnd cell_6t
Xbit_r373_c40 bl[40] br[40] wl[373] vdd gnd cell_6t
Xbit_r374_c40 bl[40] br[40] wl[374] vdd gnd cell_6t
Xbit_r375_c40 bl[40] br[40] wl[375] vdd gnd cell_6t
Xbit_r376_c40 bl[40] br[40] wl[376] vdd gnd cell_6t
Xbit_r377_c40 bl[40] br[40] wl[377] vdd gnd cell_6t
Xbit_r378_c40 bl[40] br[40] wl[378] vdd gnd cell_6t
Xbit_r379_c40 bl[40] br[40] wl[379] vdd gnd cell_6t
Xbit_r380_c40 bl[40] br[40] wl[380] vdd gnd cell_6t
Xbit_r381_c40 bl[40] br[40] wl[381] vdd gnd cell_6t
Xbit_r382_c40 bl[40] br[40] wl[382] vdd gnd cell_6t
Xbit_r383_c40 bl[40] br[40] wl[383] vdd gnd cell_6t
Xbit_r384_c40 bl[40] br[40] wl[384] vdd gnd cell_6t
Xbit_r385_c40 bl[40] br[40] wl[385] vdd gnd cell_6t
Xbit_r386_c40 bl[40] br[40] wl[386] vdd gnd cell_6t
Xbit_r387_c40 bl[40] br[40] wl[387] vdd gnd cell_6t
Xbit_r388_c40 bl[40] br[40] wl[388] vdd gnd cell_6t
Xbit_r389_c40 bl[40] br[40] wl[389] vdd gnd cell_6t
Xbit_r390_c40 bl[40] br[40] wl[390] vdd gnd cell_6t
Xbit_r391_c40 bl[40] br[40] wl[391] vdd gnd cell_6t
Xbit_r392_c40 bl[40] br[40] wl[392] vdd gnd cell_6t
Xbit_r393_c40 bl[40] br[40] wl[393] vdd gnd cell_6t
Xbit_r394_c40 bl[40] br[40] wl[394] vdd gnd cell_6t
Xbit_r395_c40 bl[40] br[40] wl[395] vdd gnd cell_6t
Xbit_r396_c40 bl[40] br[40] wl[396] vdd gnd cell_6t
Xbit_r397_c40 bl[40] br[40] wl[397] vdd gnd cell_6t
Xbit_r398_c40 bl[40] br[40] wl[398] vdd gnd cell_6t
Xbit_r399_c40 bl[40] br[40] wl[399] vdd gnd cell_6t
Xbit_r400_c40 bl[40] br[40] wl[400] vdd gnd cell_6t
Xbit_r401_c40 bl[40] br[40] wl[401] vdd gnd cell_6t
Xbit_r402_c40 bl[40] br[40] wl[402] vdd gnd cell_6t
Xbit_r403_c40 bl[40] br[40] wl[403] vdd gnd cell_6t
Xbit_r404_c40 bl[40] br[40] wl[404] vdd gnd cell_6t
Xbit_r405_c40 bl[40] br[40] wl[405] vdd gnd cell_6t
Xbit_r406_c40 bl[40] br[40] wl[406] vdd gnd cell_6t
Xbit_r407_c40 bl[40] br[40] wl[407] vdd gnd cell_6t
Xbit_r408_c40 bl[40] br[40] wl[408] vdd gnd cell_6t
Xbit_r409_c40 bl[40] br[40] wl[409] vdd gnd cell_6t
Xbit_r410_c40 bl[40] br[40] wl[410] vdd gnd cell_6t
Xbit_r411_c40 bl[40] br[40] wl[411] vdd gnd cell_6t
Xbit_r412_c40 bl[40] br[40] wl[412] vdd gnd cell_6t
Xbit_r413_c40 bl[40] br[40] wl[413] vdd gnd cell_6t
Xbit_r414_c40 bl[40] br[40] wl[414] vdd gnd cell_6t
Xbit_r415_c40 bl[40] br[40] wl[415] vdd gnd cell_6t
Xbit_r416_c40 bl[40] br[40] wl[416] vdd gnd cell_6t
Xbit_r417_c40 bl[40] br[40] wl[417] vdd gnd cell_6t
Xbit_r418_c40 bl[40] br[40] wl[418] vdd gnd cell_6t
Xbit_r419_c40 bl[40] br[40] wl[419] vdd gnd cell_6t
Xbit_r420_c40 bl[40] br[40] wl[420] vdd gnd cell_6t
Xbit_r421_c40 bl[40] br[40] wl[421] vdd gnd cell_6t
Xbit_r422_c40 bl[40] br[40] wl[422] vdd gnd cell_6t
Xbit_r423_c40 bl[40] br[40] wl[423] vdd gnd cell_6t
Xbit_r424_c40 bl[40] br[40] wl[424] vdd gnd cell_6t
Xbit_r425_c40 bl[40] br[40] wl[425] vdd gnd cell_6t
Xbit_r426_c40 bl[40] br[40] wl[426] vdd gnd cell_6t
Xbit_r427_c40 bl[40] br[40] wl[427] vdd gnd cell_6t
Xbit_r428_c40 bl[40] br[40] wl[428] vdd gnd cell_6t
Xbit_r429_c40 bl[40] br[40] wl[429] vdd gnd cell_6t
Xbit_r430_c40 bl[40] br[40] wl[430] vdd gnd cell_6t
Xbit_r431_c40 bl[40] br[40] wl[431] vdd gnd cell_6t
Xbit_r432_c40 bl[40] br[40] wl[432] vdd gnd cell_6t
Xbit_r433_c40 bl[40] br[40] wl[433] vdd gnd cell_6t
Xbit_r434_c40 bl[40] br[40] wl[434] vdd gnd cell_6t
Xbit_r435_c40 bl[40] br[40] wl[435] vdd gnd cell_6t
Xbit_r436_c40 bl[40] br[40] wl[436] vdd gnd cell_6t
Xbit_r437_c40 bl[40] br[40] wl[437] vdd gnd cell_6t
Xbit_r438_c40 bl[40] br[40] wl[438] vdd gnd cell_6t
Xbit_r439_c40 bl[40] br[40] wl[439] vdd gnd cell_6t
Xbit_r440_c40 bl[40] br[40] wl[440] vdd gnd cell_6t
Xbit_r441_c40 bl[40] br[40] wl[441] vdd gnd cell_6t
Xbit_r442_c40 bl[40] br[40] wl[442] vdd gnd cell_6t
Xbit_r443_c40 bl[40] br[40] wl[443] vdd gnd cell_6t
Xbit_r444_c40 bl[40] br[40] wl[444] vdd gnd cell_6t
Xbit_r445_c40 bl[40] br[40] wl[445] vdd gnd cell_6t
Xbit_r446_c40 bl[40] br[40] wl[446] vdd gnd cell_6t
Xbit_r447_c40 bl[40] br[40] wl[447] vdd gnd cell_6t
Xbit_r448_c40 bl[40] br[40] wl[448] vdd gnd cell_6t
Xbit_r449_c40 bl[40] br[40] wl[449] vdd gnd cell_6t
Xbit_r450_c40 bl[40] br[40] wl[450] vdd gnd cell_6t
Xbit_r451_c40 bl[40] br[40] wl[451] vdd gnd cell_6t
Xbit_r452_c40 bl[40] br[40] wl[452] vdd gnd cell_6t
Xbit_r453_c40 bl[40] br[40] wl[453] vdd gnd cell_6t
Xbit_r454_c40 bl[40] br[40] wl[454] vdd gnd cell_6t
Xbit_r455_c40 bl[40] br[40] wl[455] vdd gnd cell_6t
Xbit_r456_c40 bl[40] br[40] wl[456] vdd gnd cell_6t
Xbit_r457_c40 bl[40] br[40] wl[457] vdd gnd cell_6t
Xbit_r458_c40 bl[40] br[40] wl[458] vdd gnd cell_6t
Xbit_r459_c40 bl[40] br[40] wl[459] vdd gnd cell_6t
Xbit_r460_c40 bl[40] br[40] wl[460] vdd gnd cell_6t
Xbit_r461_c40 bl[40] br[40] wl[461] vdd gnd cell_6t
Xbit_r462_c40 bl[40] br[40] wl[462] vdd gnd cell_6t
Xbit_r463_c40 bl[40] br[40] wl[463] vdd gnd cell_6t
Xbit_r464_c40 bl[40] br[40] wl[464] vdd gnd cell_6t
Xbit_r465_c40 bl[40] br[40] wl[465] vdd gnd cell_6t
Xbit_r466_c40 bl[40] br[40] wl[466] vdd gnd cell_6t
Xbit_r467_c40 bl[40] br[40] wl[467] vdd gnd cell_6t
Xbit_r468_c40 bl[40] br[40] wl[468] vdd gnd cell_6t
Xbit_r469_c40 bl[40] br[40] wl[469] vdd gnd cell_6t
Xbit_r470_c40 bl[40] br[40] wl[470] vdd gnd cell_6t
Xbit_r471_c40 bl[40] br[40] wl[471] vdd gnd cell_6t
Xbit_r472_c40 bl[40] br[40] wl[472] vdd gnd cell_6t
Xbit_r473_c40 bl[40] br[40] wl[473] vdd gnd cell_6t
Xbit_r474_c40 bl[40] br[40] wl[474] vdd gnd cell_6t
Xbit_r475_c40 bl[40] br[40] wl[475] vdd gnd cell_6t
Xbit_r476_c40 bl[40] br[40] wl[476] vdd gnd cell_6t
Xbit_r477_c40 bl[40] br[40] wl[477] vdd gnd cell_6t
Xbit_r478_c40 bl[40] br[40] wl[478] vdd gnd cell_6t
Xbit_r479_c40 bl[40] br[40] wl[479] vdd gnd cell_6t
Xbit_r480_c40 bl[40] br[40] wl[480] vdd gnd cell_6t
Xbit_r481_c40 bl[40] br[40] wl[481] vdd gnd cell_6t
Xbit_r482_c40 bl[40] br[40] wl[482] vdd gnd cell_6t
Xbit_r483_c40 bl[40] br[40] wl[483] vdd gnd cell_6t
Xbit_r484_c40 bl[40] br[40] wl[484] vdd gnd cell_6t
Xbit_r485_c40 bl[40] br[40] wl[485] vdd gnd cell_6t
Xbit_r486_c40 bl[40] br[40] wl[486] vdd gnd cell_6t
Xbit_r487_c40 bl[40] br[40] wl[487] vdd gnd cell_6t
Xbit_r488_c40 bl[40] br[40] wl[488] vdd gnd cell_6t
Xbit_r489_c40 bl[40] br[40] wl[489] vdd gnd cell_6t
Xbit_r490_c40 bl[40] br[40] wl[490] vdd gnd cell_6t
Xbit_r491_c40 bl[40] br[40] wl[491] vdd gnd cell_6t
Xbit_r492_c40 bl[40] br[40] wl[492] vdd gnd cell_6t
Xbit_r493_c40 bl[40] br[40] wl[493] vdd gnd cell_6t
Xbit_r494_c40 bl[40] br[40] wl[494] vdd gnd cell_6t
Xbit_r495_c40 bl[40] br[40] wl[495] vdd gnd cell_6t
Xbit_r496_c40 bl[40] br[40] wl[496] vdd gnd cell_6t
Xbit_r497_c40 bl[40] br[40] wl[497] vdd gnd cell_6t
Xbit_r498_c40 bl[40] br[40] wl[498] vdd gnd cell_6t
Xbit_r499_c40 bl[40] br[40] wl[499] vdd gnd cell_6t
Xbit_r500_c40 bl[40] br[40] wl[500] vdd gnd cell_6t
Xbit_r501_c40 bl[40] br[40] wl[501] vdd gnd cell_6t
Xbit_r502_c40 bl[40] br[40] wl[502] vdd gnd cell_6t
Xbit_r503_c40 bl[40] br[40] wl[503] vdd gnd cell_6t
Xbit_r504_c40 bl[40] br[40] wl[504] vdd gnd cell_6t
Xbit_r505_c40 bl[40] br[40] wl[505] vdd gnd cell_6t
Xbit_r506_c40 bl[40] br[40] wl[506] vdd gnd cell_6t
Xbit_r507_c40 bl[40] br[40] wl[507] vdd gnd cell_6t
Xbit_r508_c40 bl[40] br[40] wl[508] vdd gnd cell_6t
Xbit_r509_c40 bl[40] br[40] wl[509] vdd gnd cell_6t
Xbit_r510_c40 bl[40] br[40] wl[510] vdd gnd cell_6t
Xbit_r511_c40 bl[40] br[40] wl[511] vdd gnd cell_6t
Xbit_r0_c41 bl[41] br[41] wl[0] vdd gnd cell_6t
Xbit_r1_c41 bl[41] br[41] wl[1] vdd gnd cell_6t
Xbit_r2_c41 bl[41] br[41] wl[2] vdd gnd cell_6t
Xbit_r3_c41 bl[41] br[41] wl[3] vdd gnd cell_6t
Xbit_r4_c41 bl[41] br[41] wl[4] vdd gnd cell_6t
Xbit_r5_c41 bl[41] br[41] wl[5] vdd gnd cell_6t
Xbit_r6_c41 bl[41] br[41] wl[6] vdd gnd cell_6t
Xbit_r7_c41 bl[41] br[41] wl[7] vdd gnd cell_6t
Xbit_r8_c41 bl[41] br[41] wl[8] vdd gnd cell_6t
Xbit_r9_c41 bl[41] br[41] wl[9] vdd gnd cell_6t
Xbit_r10_c41 bl[41] br[41] wl[10] vdd gnd cell_6t
Xbit_r11_c41 bl[41] br[41] wl[11] vdd gnd cell_6t
Xbit_r12_c41 bl[41] br[41] wl[12] vdd gnd cell_6t
Xbit_r13_c41 bl[41] br[41] wl[13] vdd gnd cell_6t
Xbit_r14_c41 bl[41] br[41] wl[14] vdd gnd cell_6t
Xbit_r15_c41 bl[41] br[41] wl[15] vdd gnd cell_6t
Xbit_r16_c41 bl[41] br[41] wl[16] vdd gnd cell_6t
Xbit_r17_c41 bl[41] br[41] wl[17] vdd gnd cell_6t
Xbit_r18_c41 bl[41] br[41] wl[18] vdd gnd cell_6t
Xbit_r19_c41 bl[41] br[41] wl[19] vdd gnd cell_6t
Xbit_r20_c41 bl[41] br[41] wl[20] vdd gnd cell_6t
Xbit_r21_c41 bl[41] br[41] wl[21] vdd gnd cell_6t
Xbit_r22_c41 bl[41] br[41] wl[22] vdd gnd cell_6t
Xbit_r23_c41 bl[41] br[41] wl[23] vdd gnd cell_6t
Xbit_r24_c41 bl[41] br[41] wl[24] vdd gnd cell_6t
Xbit_r25_c41 bl[41] br[41] wl[25] vdd gnd cell_6t
Xbit_r26_c41 bl[41] br[41] wl[26] vdd gnd cell_6t
Xbit_r27_c41 bl[41] br[41] wl[27] vdd gnd cell_6t
Xbit_r28_c41 bl[41] br[41] wl[28] vdd gnd cell_6t
Xbit_r29_c41 bl[41] br[41] wl[29] vdd gnd cell_6t
Xbit_r30_c41 bl[41] br[41] wl[30] vdd gnd cell_6t
Xbit_r31_c41 bl[41] br[41] wl[31] vdd gnd cell_6t
Xbit_r32_c41 bl[41] br[41] wl[32] vdd gnd cell_6t
Xbit_r33_c41 bl[41] br[41] wl[33] vdd gnd cell_6t
Xbit_r34_c41 bl[41] br[41] wl[34] vdd gnd cell_6t
Xbit_r35_c41 bl[41] br[41] wl[35] vdd gnd cell_6t
Xbit_r36_c41 bl[41] br[41] wl[36] vdd gnd cell_6t
Xbit_r37_c41 bl[41] br[41] wl[37] vdd gnd cell_6t
Xbit_r38_c41 bl[41] br[41] wl[38] vdd gnd cell_6t
Xbit_r39_c41 bl[41] br[41] wl[39] vdd gnd cell_6t
Xbit_r40_c41 bl[41] br[41] wl[40] vdd gnd cell_6t
Xbit_r41_c41 bl[41] br[41] wl[41] vdd gnd cell_6t
Xbit_r42_c41 bl[41] br[41] wl[42] vdd gnd cell_6t
Xbit_r43_c41 bl[41] br[41] wl[43] vdd gnd cell_6t
Xbit_r44_c41 bl[41] br[41] wl[44] vdd gnd cell_6t
Xbit_r45_c41 bl[41] br[41] wl[45] vdd gnd cell_6t
Xbit_r46_c41 bl[41] br[41] wl[46] vdd gnd cell_6t
Xbit_r47_c41 bl[41] br[41] wl[47] vdd gnd cell_6t
Xbit_r48_c41 bl[41] br[41] wl[48] vdd gnd cell_6t
Xbit_r49_c41 bl[41] br[41] wl[49] vdd gnd cell_6t
Xbit_r50_c41 bl[41] br[41] wl[50] vdd gnd cell_6t
Xbit_r51_c41 bl[41] br[41] wl[51] vdd gnd cell_6t
Xbit_r52_c41 bl[41] br[41] wl[52] vdd gnd cell_6t
Xbit_r53_c41 bl[41] br[41] wl[53] vdd gnd cell_6t
Xbit_r54_c41 bl[41] br[41] wl[54] vdd gnd cell_6t
Xbit_r55_c41 bl[41] br[41] wl[55] vdd gnd cell_6t
Xbit_r56_c41 bl[41] br[41] wl[56] vdd gnd cell_6t
Xbit_r57_c41 bl[41] br[41] wl[57] vdd gnd cell_6t
Xbit_r58_c41 bl[41] br[41] wl[58] vdd gnd cell_6t
Xbit_r59_c41 bl[41] br[41] wl[59] vdd gnd cell_6t
Xbit_r60_c41 bl[41] br[41] wl[60] vdd gnd cell_6t
Xbit_r61_c41 bl[41] br[41] wl[61] vdd gnd cell_6t
Xbit_r62_c41 bl[41] br[41] wl[62] vdd gnd cell_6t
Xbit_r63_c41 bl[41] br[41] wl[63] vdd gnd cell_6t
Xbit_r64_c41 bl[41] br[41] wl[64] vdd gnd cell_6t
Xbit_r65_c41 bl[41] br[41] wl[65] vdd gnd cell_6t
Xbit_r66_c41 bl[41] br[41] wl[66] vdd gnd cell_6t
Xbit_r67_c41 bl[41] br[41] wl[67] vdd gnd cell_6t
Xbit_r68_c41 bl[41] br[41] wl[68] vdd gnd cell_6t
Xbit_r69_c41 bl[41] br[41] wl[69] vdd gnd cell_6t
Xbit_r70_c41 bl[41] br[41] wl[70] vdd gnd cell_6t
Xbit_r71_c41 bl[41] br[41] wl[71] vdd gnd cell_6t
Xbit_r72_c41 bl[41] br[41] wl[72] vdd gnd cell_6t
Xbit_r73_c41 bl[41] br[41] wl[73] vdd gnd cell_6t
Xbit_r74_c41 bl[41] br[41] wl[74] vdd gnd cell_6t
Xbit_r75_c41 bl[41] br[41] wl[75] vdd gnd cell_6t
Xbit_r76_c41 bl[41] br[41] wl[76] vdd gnd cell_6t
Xbit_r77_c41 bl[41] br[41] wl[77] vdd gnd cell_6t
Xbit_r78_c41 bl[41] br[41] wl[78] vdd gnd cell_6t
Xbit_r79_c41 bl[41] br[41] wl[79] vdd gnd cell_6t
Xbit_r80_c41 bl[41] br[41] wl[80] vdd gnd cell_6t
Xbit_r81_c41 bl[41] br[41] wl[81] vdd gnd cell_6t
Xbit_r82_c41 bl[41] br[41] wl[82] vdd gnd cell_6t
Xbit_r83_c41 bl[41] br[41] wl[83] vdd gnd cell_6t
Xbit_r84_c41 bl[41] br[41] wl[84] vdd gnd cell_6t
Xbit_r85_c41 bl[41] br[41] wl[85] vdd gnd cell_6t
Xbit_r86_c41 bl[41] br[41] wl[86] vdd gnd cell_6t
Xbit_r87_c41 bl[41] br[41] wl[87] vdd gnd cell_6t
Xbit_r88_c41 bl[41] br[41] wl[88] vdd gnd cell_6t
Xbit_r89_c41 bl[41] br[41] wl[89] vdd gnd cell_6t
Xbit_r90_c41 bl[41] br[41] wl[90] vdd gnd cell_6t
Xbit_r91_c41 bl[41] br[41] wl[91] vdd gnd cell_6t
Xbit_r92_c41 bl[41] br[41] wl[92] vdd gnd cell_6t
Xbit_r93_c41 bl[41] br[41] wl[93] vdd gnd cell_6t
Xbit_r94_c41 bl[41] br[41] wl[94] vdd gnd cell_6t
Xbit_r95_c41 bl[41] br[41] wl[95] vdd gnd cell_6t
Xbit_r96_c41 bl[41] br[41] wl[96] vdd gnd cell_6t
Xbit_r97_c41 bl[41] br[41] wl[97] vdd gnd cell_6t
Xbit_r98_c41 bl[41] br[41] wl[98] vdd gnd cell_6t
Xbit_r99_c41 bl[41] br[41] wl[99] vdd gnd cell_6t
Xbit_r100_c41 bl[41] br[41] wl[100] vdd gnd cell_6t
Xbit_r101_c41 bl[41] br[41] wl[101] vdd gnd cell_6t
Xbit_r102_c41 bl[41] br[41] wl[102] vdd gnd cell_6t
Xbit_r103_c41 bl[41] br[41] wl[103] vdd gnd cell_6t
Xbit_r104_c41 bl[41] br[41] wl[104] vdd gnd cell_6t
Xbit_r105_c41 bl[41] br[41] wl[105] vdd gnd cell_6t
Xbit_r106_c41 bl[41] br[41] wl[106] vdd gnd cell_6t
Xbit_r107_c41 bl[41] br[41] wl[107] vdd gnd cell_6t
Xbit_r108_c41 bl[41] br[41] wl[108] vdd gnd cell_6t
Xbit_r109_c41 bl[41] br[41] wl[109] vdd gnd cell_6t
Xbit_r110_c41 bl[41] br[41] wl[110] vdd gnd cell_6t
Xbit_r111_c41 bl[41] br[41] wl[111] vdd gnd cell_6t
Xbit_r112_c41 bl[41] br[41] wl[112] vdd gnd cell_6t
Xbit_r113_c41 bl[41] br[41] wl[113] vdd gnd cell_6t
Xbit_r114_c41 bl[41] br[41] wl[114] vdd gnd cell_6t
Xbit_r115_c41 bl[41] br[41] wl[115] vdd gnd cell_6t
Xbit_r116_c41 bl[41] br[41] wl[116] vdd gnd cell_6t
Xbit_r117_c41 bl[41] br[41] wl[117] vdd gnd cell_6t
Xbit_r118_c41 bl[41] br[41] wl[118] vdd gnd cell_6t
Xbit_r119_c41 bl[41] br[41] wl[119] vdd gnd cell_6t
Xbit_r120_c41 bl[41] br[41] wl[120] vdd gnd cell_6t
Xbit_r121_c41 bl[41] br[41] wl[121] vdd gnd cell_6t
Xbit_r122_c41 bl[41] br[41] wl[122] vdd gnd cell_6t
Xbit_r123_c41 bl[41] br[41] wl[123] vdd gnd cell_6t
Xbit_r124_c41 bl[41] br[41] wl[124] vdd gnd cell_6t
Xbit_r125_c41 bl[41] br[41] wl[125] vdd gnd cell_6t
Xbit_r126_c41 bl[41] br[41] wl[126] vdd gnd cell_6t
Xbit_r127_c41 bl[41] br[41] wl[127] vdd gnd cell_6t
Xbit_r128_c41 bl[41] br[41] wl[128] vdd gnd cell_6t
Xbit_r129_c41 bl[41] br[41] wl[129] vdd gnd cell_6t
Xbit_r130_c41 bl[41] br[41] wl[130] vdd gnd cell_6t
Xbit_r131_c41 bl[41] br[41] wl[131] vdd gnd cell_6t
Xbit_r132_c41 bl[41] br[41] wl[132] vdd gnd cell_6t
Xbit_r133_c41 bl[41] br[41] wl[133] vdd gnd cell_6t
Xbit_r134_c41 bl[41] br[41] wl[134] vdd gnd cell_6t
Xbit_r135_c41 bl[41] br[41] wl[135] vdd gnd cell_6t
Xbit_r136_c41 bl[41] br[41] wl[136] vdd gnd cell_6t
Xbit_r137_c41 bl[41] br[41] wl[137] vdd gnd cell_6t
Xbit_r138_c41 bl[41] br[41] wl[138] vdd gnd cell_6t
Xbit_r139_c41 bl[41] br[41] wl[139] vdd gnd cell_6t
Xbit_r140_c41 bl[41] br[41] wl[140] vdd gnd cell_6t
Xbit_r141_c41 bl[41] br[41] wl[141] vdd gnd cell_6t
Xbit_r142_c41 bl[41] br[41] wl[142] vdd gnd cell_6t
Xbit_r143_c41 bl[41] br[41] wl[143] vdd gnd cell_6t
Xbit_r144_c41 bl[41] br[41] wl[144] vdd gnd cell_6t
Xbit_r145_c41 bl[41] br[41] wl[145] vdd gnd cell_6t
Xbit_r146_c41 bl[41] br[41] wl[146] vdd gnd cell_6t
Xbit_r147_c41 bl[41] br[41] wl[147] vdd gnd cell_6t
Xbit_r148_c41 bl[41] br[41] wl[148] vdd gnd cell_6t
Xbit_r149_c41 bl[41] br[41] wl[149] vdd gnd cell_6t
Xbit_r150_c41 bl[41] br[41] wl[150] vdd gnd cell_6t
Xbit_r151_c41 bl[41] br[41] wl[151] vdd gnd cell_6t
Xbit_r152_c41 bl[41] br[41] wl[152] vdd gnd cell_6t
Xbit_r153_c41 bl[41] br[41] wl[153] vdd gnd cell_6t
Xbit_r154_c41 bl[41] br[41] wl[154] vdd gnd cell_6t
Xbit_r155_c41 bl[41] br[41] wl[155] vdd gnd cell_6t
Xbit_r156_c41 bl[41] br[41] wl[156] vdd gnd cell_6t
Xbit_r157_c41 bl[41] br[41] wl[157] vdd gnd cell_6t
Xbit_r158_c41 bl[41] br[41] wl[158] vdd gnd cell_6t
Xbit_r159_c41 bl[41] br[41] wl[159] vdd gnd cell_6t
Xbit_r160_c41 bl[41] br[41] wl[160] vdd gnd cell_6t
Xbit_r161_c41 bl[41] br[41] wl[161] vdd gnd cell_6t
Xbit_r162_c41 bl[41] br[41] wl[162] vdd gnd cell_6t
Xbit_r163_c41 bl[41] br[41] wl[163] vdd gnd cell_6t
Xbit_r164_c41 bl[41] br[41] wl[164] vdd gnd cell_6t
Xbit_r165_c41 bl[41] br[41] wl[165] vdd gnd cell_6t
Xbit_r166_c41 bl[41] br[41] wl[166] vdd gnd cell_6t
Xbit_r167_c41 bl[41] br[41] wl[167] vdd gnd cell_6t
Xbit_r168_c41 bl[41] br[41] wl[168] vdd gnd cell_6t
Xbit_r169_c41 bl[41] br[41] wl[169] vdd gnd cell_6t
Xbit_r170_c41 bl[41] br[41] wl[170] vdd gnd cell_6t
Xbit_r171_c41 bl[41] br[41] wl[171] vdd gnd cell_6t
Xbit_r172_c41 bl[41] br[41] wl[172] vdd gnd cell_6t
Xbit_r173_c41 bl[41] br[41] wl[173] vdd gnd cell_6t
Xbit_r174_c41 bl[41] br[41] wl[174] vdd gnd cell_6t
Xbit_r175_c41 bl[41] br[41] wl[175] vdd gnd cell_6t
Xbit_r176_c41 bl[41] br[41] wl[176] vdd gnd cell_6t
Xbit_r177_c41 bl[41] br[41] wl[177] vdd gnd cell_6t
Xbit_r178_c41 bl[41] br[41] wl[178] vdd gnd cell_6t
Xbit_r179_c41 bl[41] br[41] wl[179] vdd gnd cell_6t
Xbit_r180_c41 bl[41] br[41] wl[180] vdd gnd cell_6t
Xbit_r181_c41 bl[41] br[41] wl[181] vdd gnd cell_6t
Xbit_r182_c41 bl[41] br[41] wl[182] vdd gnd cell_6t
Xbit_r183_c41 bl[41] br[41] wl[183] vdd gnd cell_6t
Xbit_r184_c41 bl[41] br[41] wl[184] vdd gnd cell_6t
Xbit_r185_c41 bl[41] br[41] wl[185] vdd gnd cell_6t
Xbit_r186_c41 bl[41] br[41] wl[186] vdd gnd cell_6t
Xbit_r187_c41 bl[41] br[41] wl[187] vdd gnd cell_6t
Xbit_r188_c41 bl[41] br[41] wl[188] vdd gnd cell_6t
Xbit_r189_c41 bl[41] br[41] wl[189] vdd gnd cell_6t
Xbit_r190_c41 bl[41] br[41] wl[190] vdd gnd cell_6t
Xbit_r191_c41 bl[41] br[41] wl[191] vdd gnd cell_6t
Xbit_r192_c41 bl[41] br[41] wl[192] vdd gnd cell_6t
Xbit_r193_c41 bl[41] br[41] wl[193] vdd gnd cell_6t
Xbit_r194_c41 bl[41] br[41] wl[194] vdd gnd cell_6t
Xbit_r195_c41 bl[41] br[41] wl[195] vdd gnd cell_6t
Xbit_r196_c41 bl[41] br[41] wl[196] vdd gnd cell_6t
Xbit_r197_c41 bl[41] br[41] wl[197] vdd gnd cell_6t
Xbit_r198_c41 bl[41] br[41] wl[198] vdd gnd cell_6t
Xbit_r199_c41 bl[41] br[41] wl[199] vdd gnd cell_6t
Xbit_r200_c41 bl[41] br[41] wl[200] vdd gnd cell_6t
Xbit_r201_c41 bl[41] br[41] wl[201] vdd gnd cell_6t
Xbit_r202_c41 bl[41] br[41] wl[202] vdd gnd cell_6t
Xbit_r203_c41 bl[41] br[41] wl[203] vdd gnd cell_6t
Xbit_r204_c41 bl[41] br[41] wl[204] vdd gnd cell_6t
Xbit_r205_c41 bl[41] br[41] wl[205] vdd gnd cell_6t
Xbit_r206_c41 bl[41] br[41] wl[206] vdd gnd cell_6t
Xbit_r207_c41 bl[41] br[41] wl[207] vdd gnd cell_6t
Xbit_r208_c41 bl[41] br[41] wl[208] vdd gnd cell_6t
Xbit_r209_c41 bl[41] br[41] wl[209] vdd gnd cell_6t
Xbit_r210_c41 bl[41] br[41] wl[210] vdd gnd cell_6t
Xbit_r211_c41 bl[41] br[41] wl[211] vdd gnd cell_6t
Xbit_r212_c41 bl[41] br[41] wl[212] vdd gnd cell_6t
Xbit_r213_c41 bl[41] br[41] wl[213] vdd gnd cell_6t
Xbit_r214_c41 bl[41] br[41] wl[214] vdd gnd cell_6t
Xbit_r215_c41 bl[41] br[41] wl[215] vdd gnd cell_6t
Xbit_r216_c41 bl[41] br[41] wl[216] vdd gnd cell_6t
Xbit_r217_c41 bl[41] br[41] wl[217] vdd gnd cell_6t
Xbit_r218_c41 bl[41] br[41] wl[218] vdd gnd cell_6t
Xbit_r219_c41 bl[41] br[41] wl[219] vdd gnd cell_6t
Xbit_r220_c41 bl[41] br[41] wl[220] vdd gnd cell_6t
Xbit_r221_c41 bl[41] br[41] wl[221] vdd gnd cell_6t
Xbit_r222_c41 bl[41] br[41] wl[222] vdd gnd cell_6t
Xbit_r223_c41 bl[41] br[41] wl[223] vdd gnd cell_6t
Xbit_r224_c41 bl[41] br[41] wl[224] vdd gnd cell_6t
Xbit_r225_c41 bl[41] br[41] wl[225] vdd gnd cell_6t
Xbit_r226_c41 bl[41] br[41] wl[226] vdd gnd cell_6t
Xbit_r227_c41 bl[41] br[41] wl[227] vdd gnd cell_6t
Xbit_r228_c41 bl[41] br[41] wl[228] vdd gnd cell_6t
Xbit_r229_c41 bl[41] br[41] wl[229] vdd gnd cell_6t
Xbit_r230_c41 bl[41] br[41] wl[230] vdd gnd cell_6t
Xbit_r231_c41 bl[41] br[41] wl[231] vdd gnd cell_6t
Xbit_r232_c41 bl[41] br[41] wl[232] vdd gnd cell_6t
Xbit_r233_c41 bl[41] br[41] wl[233] vdd gnd cell_6t
Xbit_r234_c41 bl[41] br[41] wl[234] vdd gnd cell_6t
Xbit_r235_c41 bl[41] br[41] wl[235] vdd gnd cell_6t
Xbit_r236_c41 bl[41] br[41] wl[236] vdd gnd cell_6t
Xbit_r237_c41 bl[41] br[41] wl[237] vdd gnd cell_6t
Xbit_r238_c41 bl[41] br[41] wl[238] vdd gnd cell_6t
Xbit_r239_c41 bl[41] br[41] wl[239] vdd gnd cell_6t
Xbit_r240_c41 bl[41] br[41] wl[240] vdd gnd cell_6t
Xbit_r241_c41 bl[41] br[41] wl[241] vdd gnd cell_6t
Xbit_r242_c41 bl[41] br[41] wl[242] vdd gnd cell_6t
Xbit_r243_c41 bl[41] br[41] wl[243] vdd gnd cell_6t
Xbit_r244_c41 bl[41] br[41] wl[244] vdd gnd cell_6t
Xbit_r245_c41 bl[41] br[41] wl[245] vdd gnd cell_6t
Xbit_r246_c41 bl[41] br[41] wl[246] vdd gnd cell_6t
Xbit_r247_c41 bl[41] br[41] wl[247] vdd gnd cell_6t
Xbit_r248_c41 bl[41] br[41] wl[248] vdd gnd cell_6t
Xbit_r249_c41 bl[41] br[41] wl[249] vdd gnd cell_6t
Xbit_r250_c41 bl[41] br[41] wl[250] vdd gnd cell_6t
Xbit_r251_c41 bl[41] br[41] wl[251] vdd gnd cell_6t
Xbit_r252_c41 bl[41] br[41] wl[252] vdd gnd cell_6t
Xbit_r253_c41 bl[41] br[41] wl[253] vdd gnd cell_6t
Xbit_r254_c41 bl[41] br[41] wl[254] vdd gnd cell_6t
Xbit_r255_c41 bl[41] br[41] wl[255] vdd gnd cell_6t
Xbit_r256_c41 bl[41] br[41] wl[256] vdd gnd cell_6t
Xbit_r257_c41 bl[41] br[41] wl[257] vdd gnd cell_6t
Xbit_r258_c41 bl[41] br[41] wl[258] vdd gnd cell_6t
Xbit_r259_c41 bl[41] br[41] wl[259] vdd gnd cell_6t
Xbit_r260_c41 bl[41] br[41] wl[260] vdd gnd cell_6t
Xbit_r261_c41 bl[41] br[41] wl[261] vdd gnd cell_6t
Xbit_r262_c41 bl[41] br[41] wl[262] vdd gnd cell_6t
Xbit_r263_c41 bl[41] br[41] wl[263] vdd gnd cell_6t
Xbit_r264_c41 bl[41] br[41] wl[264] vdd gnd cell_6t
Xbit_r265_c41 bl[41] br[41] wl[265] vdd gnd cell_6t
Xbit_r266_c41 bl[41] br[41] wl[266] vdd gnd cell_6t
Xbit_r267_c41 bl[41] br[41] wl[267] vdd gnd cell_6t
Xbit_r268_c41 bl[41] br[41] wl[268] vdd gnd cell_6t
Xbit_r269_c41 bl[41] br[41] wl[269] vdd gnd cell_6t
Xbit_r270_c41 bl[41] br[41] wl[270] vdd gnd cell_6t
Xbit_r271_c41 bl[41] br[41] wl[271] vdd gnd cell_6t
Xbit_r272_c41 bl[41] br[41] wl[272] vdd gnd cell_6t
Xbit_r273_c41 bl[41] br[41] wl[273] vdd gnd cell_6t
Xbit_r274_c41 bl[41] br[41] wl[274] vdd gnd cell_6t
Xbit_r275_c41 bl[41] br[41] wl[275] vdd gnd cell_6t
Xbit_r276_c41 bl[41] br[41] wl[276] vdd gnd cell_6t
Xbit_r277_c41 bl[41] br[41] wl[277] vdd gnd cell_6t
Xbit_r278_c41 bl[41] br[41] wl[278] vdd gnd cell_6t
Xbit_r279_c41 bl[41] br[41] wl[279] vdd gnd cell_6t
Xbit_r280_c41 bl[41] br[41] wl[280] vdd gnd cell_6t
Xbit_r281_c41 bl[41] br[41] wl[281] vdd gnd cell_6t
Xbit_r282_c41 bl[41] br[41] wl[282] vdd gnd cell_6t
Xbit_r283_c41 bl[41] br[41] wl[283] vdd gnd cell_6t
Xbit_r284_c41 bl[41] br[41] wl[284] vdd gnd cell_6t
Xbit_r285_c41 bl[41] br[41] wl[285] vdd gnd cell_6t
Xbit_r286_c41 bl[41] br[41] wl[286] vdd gnd cell_6t
Xbit_r287_c41 bl[41] br[41] wl[287] vdd gnd cell_6t
Xbit_r288_c41 bl[41] br[41] wl[288] vdd gnd cell_6t
Xbit_r289_c41 bl[41] br[41] wl[289] vdd gnd cell_6t
Xbit_r290_c41 bl[41] br[41] wl[290] vdd gnd cell_6t
Xbit_r291_c41 bl[41] br[41] wl[291] vdd gnd cell_6t
Xbit_r292_c41 bl[41] br[41] wl[292] vdd gnd cell_6t
Xbit_r293_c41 bl[41] br[41] wl[293] vdd gnd cell_6t
Xbit_r294_c41 bl[41] br[41] wl[294] vdd gnd cell_6t
Xbit_r295_c41 bl[41] br[41] wl[295] vdd gnd cell_6t
Xbit_r296_c41 bl[41] br[41] wl[296] vdd gnd cell_6t
Xbit_r297_c41 bl[41] br[41] wl[297] vdd gnd cell_6t
Xbit_r298_c41 bl[41] br[41] wl[298] vdd gnd cell_6t
Xbit_r299_c41 bl[41] br[41] wl[299] vdd gnd cell_6t
Xbit_r300_c41 bl[41] br[41] wl[300] vdd gnd cell_6t
Xbit_r301_c41 bl[41] br[41] wl[301] vdd gnd cell_6t
Xbit_r302_c41 bl[41] br[41] wl[302] vdd gnd cell_6t
Xbit_r303_c41 bl[41] br[41] wl[303] vdd gnd cell_6t
Xbit_r304_c41 bl[41] br[41] wl[304] vdd gnd cell_6t
Xbit_r305_c41 bl[41] br[41] wl[305] vdd gnd cell_6t
Xbit_r306_c41 bl[41] br[41] wl[306] vdd gnd cell_6t
Xbit_r307_c41 bl[41] br[41] wl[307] vdd gnd cell_6t
Xbit_r308_c41 bl[41] br[41] wl[308] vdd gnd cell_6t
Xbit_r309_c41 bl[41] br[41] wl[309] vdd gnd cell_6t
Xbit_r310_c41 bl[41] br[41] wl[310] vdd gnd cell_6t
Xbit_r311_c41 bl[41] br[41] wl[311] vdd gnd cell_6t
Xbit_r312_c41 bl[41] br[41] wl[312] vdd gnd cell_6t
Xbit_r313_c41 bl[41] br[41] wl[313] vdd gnd cell_6t
Xbit_r314_c41 bl[41] br[41] wl[314] vdd gnd cell_6t
Xbit_r315_c41 bl[41] br[41] wl[315] vdd gnd cell_6t
Xbit_r316_c41 bl[41] br[41] wl[316] vdd gnd cell_6t
Xbit_r317_c41 bl[41] br[41] wl[317] vdd gnd cell_6t
Xbit_r318_c41 bl[41] br[41] wl[318] vdd gnd cell_6t
Xbit_r319_c41 bl[41] br[41] wl[319] vdd gnd cell_6t
Xbit_r320_c41 bl[41] br[41] wl[320] vdd gnd cell_6t
Xbit_r321_c41 bl[41] br[41] wl[321] vdd gnd cell_6t
Xbit_r322_c41 bl[41] br[41] wl[322] vdd gnd cell_6t
Xbit_r323_c41 bl[41] br[41] wl[323] vdd gnd cell_6t
Xbit_r324_c41 bl[41] br[41] wl[324] vdd gnd cell_6t
Xbit_r325_c41 bl[41] br[41] wl[325] vdd gnd cell_6t
Xbit_r326_c41 bl[41] br[41] wl[326] vdd gnd cell_6t
Xbit_r327_c41 bl[41] br[41] wl[327] vdd gnd cell_6t
Xbit_r328_c41 bl[41] br[41] wl[328] vdd gnd cell_6t
Xbit_r329_c41 bl[41] br[41] wl[329] vdd gnd cell_6t
Xbit_r330_c41 bl[41] br[41] wl[330] vdd gnd cell_6t
Xbit_r331_c41 bl[41] br[41] wl[331] vdd gnd cell_6t
Xbit_r332_c41 bl[41] br[41] wl[332] vdd gnd cell_6t
Xbit_r333_c41 bl[41] br[41] wl[333] vdd gnd cell_6t
Xbit_r334_c41 bl[41] br[41] wl[334] vdd gnd cell_6t
Xbit_r335_c41 bl[41] br[41] wl[335] vdd gnd cell_6t
Xbit_r336_c41 bl[41] br[41] wl[336] vdd gnd cell_6t
Xbit_r337_c41 bl[41] br[41] wl[337] vdd gnd cell_6t
Xbit_r338_c41 bl[41] br[41] wl[338] vdd gnd cell_6t
Xbit_r339_c41 bl[41] br[41] wl[339] vdd gnd cell_6t
Xbit_r340_c41 bl[41] br[41] wl[340] vdd gnd cell_6t
Xbit_r341_c41 bl[41] br[41] wl[341] vdd gnd cell_6t
Xbit_r342_c41 bl[41] br[41] wl[342] vdd gnd cell_6t
Xbit_r343_c41 bl[41] br[41] wl[343] vdd gnd cell_6t
Xbit_r344_c41 bl[41] br[41] wl[344] vdd gnd cell_6t
Xbit_r345_c41 bl[41] br[41] wl[345] vdd gnd cell_6t
Xbit_r346_c41 bl[41] br[41] wl[346] vdd gnd cell_6t
Xbit_r347_c41 bl[41] br[41] wl[347] vdd gnd cell_6t
Xbit_r348_c41 bl[41] br[41] wl[348] vdd gnd cell_6t
Xbit_r349_c41 bl[41] br[41] wl[349] vdd gnd cell_6t
Xbit_r350_c41 bl[41] br[41] wl[350] vdd gnd cell_6t
Xbit_r351_c41 bl[41] br[41] wl[351] vdd gnd cell_6t
Xbit_r352_c41 bl[41] br[41] wl[352] vdd gnd cell_6t
Xbit_r353_c41 bl[41] br[41] wl[353] vdd gnd cell_6t
Xbit_r354_c41 bl[41] br[41] wl[354] vdd gnd cell_6t
Xbit_r355_c41 bl[41] br[41] wl[355] vdd gnd cell_6t
Xbit_r356_c41 bl[41] br[41] wl[356] vdd gnd cell_6t
Xbit_r357_c41 bl[41] br[41] wl[357] vdd gnd cell_6t
Xbit_r358_c41 bl[41] br[41] wl[358] vdd gnd cell_6t
Xbit_r359_c41 bl[41] br[41] wl[359] vdd gnd cell_6t
Xbit_r360_c41 bl[41] br[41] wl[360] vdd gnd cell_6t
Xbit_r361_c41 bl[41] br[41] wl[361] vdd gnd cell_6t
Xbit_r362_c41 bl[41] br[41] wl[362] vdd gnd cell_6t
Xbit_r363_c41 bl[41] br[41] wl[363] vdd gnd cell_6t
Xbit_r364_c41 bl[41] br[41] wl[364] vdd gnd cell_6t
Xbit_r365_c41 bl[41] br[41] wl[365] vdd gnd cell_6t
Xbit_r366_c41 bl[41] br[41] wl[366] vdd gnd cell_6t
Xbit_r367_c41 bl[41] br[41] wl[367] vdd gnd cell_6t
Xbit_r368_c41 bl[41] br[41] wl[368] vdd gnd cell_6t
Xbit_r369_c41 bl[41] br[41] wl[369] vdd gnd cell_6t
Xbit_r370_c41 bl[41] br[41] wl[370] vdd gnd cell_6t
Xbit_r371_c41 bl[41] br[41] wl[371] vdd gnd cell_6t
Xbit_r372_c41 bl[41] br[41] wl[372] vdd gnd cell_6t
Xbit_r373_c41 bl[41] br[41] wl[373] vdd gnd cell_6t
Xbit_r374_c41 bl[41] br[41] wl[374] vdd gnd cell_6t
Xbit_r375_c41 bl[41] br[41] wl[375] vdd gnd cell_6t
Xbit_r376_c41 bl[41] br[41] wl[376] vdd gnd cell_6t
Xbit_r377_c41 bl[41] br[41] wl[377] vdd gnd cell_6t
Xbit_r378_c41 bl[41] br[41] wl[378] vdd gnd cell_6t
Xbit_r379_c41 bl[41] br[41] wl[379] vdd gnd cell_6t
Xbit_r380_c41 bl[41] br[41] wl[380] vdd gnd cell_6t
Xbit_r381_c41 bl[41] br[41] wl[381] vdd gnd cell_6t
Xbit_r382_c41 bl[41] br[41] wl[382] vdd gnd cell_6t
Xbit_r383_c41 bl[41] br[41] wl[383] vdd gnd cell_6t
Xbit_r384_c41 bl[41] br[41] wl[384] vdd gnd cell_6t
Xbit_r385_c41 bl[41] br[41] wl[385] vdd gnd cell_6t
Xbit_r386_c41 bl[41] br[41] wl[386] vdd gnd cell_6t
Xbit_r387_c41 bl[41] br[41] wl[387] vdd gnd cell_6t
Xbit_r388_c41 bl[41] br[41] wl[388] vdd gnd cell_6t
Xbit_r389_c41 bl[41] br[41] wl[389] vdd gnd cell_6t
Xbit_r390_c41 bl[41] br[41] wl[390] vdd gnd cell_6t
Xbit_r391_c41 bl[41] br[41] wl[391] vdd gnd cell_6t
Xbit_r392_c41 bl[41] br[41] wl[392] vdd gnd cell_6t
Xbit_r393_c41 bl[41] br[41] wl[393] vdd gnd cell_6t
Xbit_r394_c41 bl[41] br[41] wl[394] vdd gnd cell_6t
Xbit_r395_c41 bl[41] br[41] wl[395] vdd gnd cell_6t
Xbit_r396_c41 bl[41] br[41] wl[396] vdd gnd cell_6t
Xbit_r397_c41 bl[41] br[41] wl[397] vdd gnd cell_6t
Xbit_r398_c41 bl[41] br[41] wl[398] vdd gnd cell_6t
Xbit_r399_c41 bl[41] br[41] wl[399] vdd gnd cell_6t
Xbit_r400_c41 bl[41] br[41] wl[400] vdd gnd cell_6t
Xbit_r401_c41 bl[41] br[41] wl[401] vdd gnd cell_6t
Xbit_r402_c41 bl[41] br[41] wl[402] vdd gnd cell_6t
Xbit_r403_c41 bl[41] br[41] wl[403] vdd gnd cell_6t
Xbit_r404_c41 bl[41] br[41] wl[404] vdd gnd cell_6t
Xbit_r405_c41 bl[41] br[41] wl[405] vdd gnd cell_6t
Xbit_r406_c41 bl[41] br[41] wl[406] vdd gnd cell_6t
Xbit_r407_c41 bl[41] br[41] wl[407] vdd gnd cell_6t
Xbit_r408_c41 bl[41] br[41] wl[408] vdd gnd cell_6t
Xbit_r409_c41 bl[41] br[41] wl[409] vdd gnd cell_6t
Xbit_r410_c41 bl[41] br[41] wl[410] vdd gnd cell_6t
Xbit_r411_c41 bl[41] br[41] wl[411] vdd gnd cell_6t
Xbit_r412_c41 bl[41] br[41] wl[412] vdd gnd cell_6t
Xbit_r413_c41 bl[41] br[41] wl[413] vdd gnd cell_6t
Xbit_r414_c41 bl[41] br[41] wl[414] vdd gnd cell_6t
Xbit_r415_c41 bl[41] br[41] wl[415] vdd gnd cell_6t
Xbit_r416_c41 bl[41] br[41] wl[416] vdd gnd cell_6t
Xbit_r417_c41 bl[41] br[41] wl[417] vdd gnd cell_6t
Xbit_r418_c41 bl[41] br[41] wl[418] vdd gnd cell_6t
Xbit_r419_c41 bl[41] br[41] wl[419] vdd gnd cell_6t
Xbit_r420_c41 bl[41] br[41] wl[420] vdd gnd cell_6t
Xbit_r421_c41 bl[41] br[41] wl[421] vdd gnd cell_6t
Xbit_r422_c41 bl[41] br[41] wl[422] vdd gnd cell_6t
Xbit_r423_c41 bl[41] br[41] wl[423] vdd gnd cell_6t
Xbit_r424_c41 bl[41] br[41] wl[424] vdd gnd cell_6t
Xbit_r425_c41 bl[41] br[41] wl[425] vdd gnd cell_6t
Xbit_r426_c41 bl[41] br[41] wl[426] vdd gnd cell_6t
Xbit_r427_c41 bl[41] br[41] wl[427] vdd gnd cell_6t
Xbit_r428_c41 bl[41] br[41] wl[428] vdd gnd cell_6t
Xbit_r429_c41 bl[41] br[41] wl[429] vdd gnd cell_6t
Xbit_r430_c41 bl[41] br[41] wl[430] vdd gnd cell_6t
Xbit_r431_c41 bl[41] br[41] wl[431] vdd gnd cell_6t
Xbit_r432_c41 bl[41] br[41] wl[432] vdd gnd cell_6t
Xbit_r433_c41 bl[41] br[41] wl[433] vdd gnd cell_6t
Xbit_r434_c41 bl[41] br[41] wl[434] vdd gnd cell_6t
Xbit_r435_c41 bl[41] br[41] wl[435] vdd gnd cell_6t
Xbit_r436_c41 bl[41] br[41] wl[436] vdd gnd cell_6t
Xbit_r437_c41 bl[41] br[41] wl[437] vdd gnd cell_6t
Xbit_r438_c41 bl[41] br[41] wl[438] vdd gnd cell_6t
Xbit_r439_c41 bl[41] br[41] wl[439] vdd gnd cell_6t
Xbit_r440_c41 bl[41] br[41] wl[440] vdd gnd cell_6t
Xbit_r441_c41 bl[41] br[41] wl[441] vdd gnd cell_6t
Xbit_r442_c41 bl[41] br[41] wl[442] vdd gnd cell_6t
Xbit_r443_c41 bl[41] br[41] wl[443] vdd gnd cell_6t
Xbit_r444_c41 bl[41] br[41] wl[444] vdd gnd cell_6t
Xbit_r445_c41 bl[41] br[41] wl[445] vdd gnd cell_6t
Xbit_r446_c41 bl[41] br[41] wl[446] vdd gnd cell_6t
Xbit_r447_c41 bl[41] br[41] wl[447] vdd gnd cell_6t
Xbit_r448_c41 bl[41] br[41] wl[448] vdd gnd cell_6t
Xbit_r449_c41 bl[41] br[41] wl[449] vdd gnd cell_6t
Xbit_r450_c41 bl[41] br[41] wl[450] vdd gnd cell_6t
Xbit_r451_c41 bl[41] br[41] wl[451] vdd gnd cell_6t
Xbit_r452_c41 bl[41] br[41] wl[452] vdd gnd cell_6t
Xbit_r453_c41 bl[41] br[41] wl[453] vdd gnd cell_6t
Xbit_r454_c41 bl[41] br[41] wl[454] vdd gnd cell_6t
Xbit_r455_c41 bl[41] br[41] wl[455] vdd gnd cell_6t
Xbit_r456_c41 bl[41] br[41] wl[456] vdd gnd cell_6t
Xbit_r457_c41 bl[41] br[41] wl[457] vdd gnd cell_6t
Xbit_r458_c41 bl[41] br[41] wl[458] vdd gnd cell_6t
Xbit_r459_c41 bl[41] br[41] wl[459] vdd gnd cell_6t
Xbit_r460_c41 bl[41] br[41] wl[460] vdd gnd cell_6t
Xbit_r461_c41 bl[41] br[41] wl[461] vdd gnd cell_6t
Xbit_r462_c41 bl[41] br[41] wl[462] vdd gnd cell_6t
Xbit_r463_c41 bl[41] br[41] wl[463] vdd gnd cell_6t
Xbit_r464_c41 bl[41] br[41] wl[464] vdd gnd cell_6t
Xbit_r465_c41 bl[41] br[41] wl[465] vdd gnd cell_6t
Xbit_r466_c41 bl[41] br[41] wl[466] vdd gnd cell_6t
Xbit_r467_c41 bl[41] br[41] wl[467] vdd gnd cell_6t
Xbit_r468_c41 bl[41] br[41] wl[468] vdd gnd cell_6t
Xbit_r469_c41 bl[41] br[41] wl[469] vdd gnd cell_6t
Xbit_r470_c41 bl[41] br[41] wl[470] vdd gnd cell_6t
Xbit_r471_c41 bl[41] br[41] wl[471] vdd gnd cell_6t
Xbit_r472_c41 bl[41] br[41] wl[472] vdd gnd cell_6t
Xbit_r473_c41 bl[41] br[41] wl[473] vdd gnd cell_6t
Xbit_r474_c41 bl[41] br[41] wl[474] vdd gnd cell_6t
Xbit_r475_c41 bl[41] br[41] wl[475] vdd gnd cell_6t
Xbit_r476_c41 bl[41] br[41] wl[476] vdd gnd cell_6t
Xbit_r477_c41 bl[41] br[41] wl[477] vdd gnd cell_6t
Xbit_r478_c41 bl[41] br[41] wl[478] vdd gnd cell_6t
Xbit_r479_c41 bl[41] br[41] wl[479] vdd gnd cell_6t
Xbit_r480_c41 bl[41] br[41] wl[480] vdd gnd cell_6t
Xbit_r481_c41 bl[41] br[41] wl[481] vdd gnd cell_6t
Xbit_r482_c41 bl[41] br[41] wl[482] vdd gnd cell_6t
Xbit_r483_c41 bl[41] br[41] wl[483] vdd gnd cell_6t
Xbit_r484_c41 bl[41] br[41] wl[484] vdd gnd cell_6t
Xbit_r485_c41 bl[41] br[41] wl[485] vdd gnd cell_6t
Xbit_r486_c41 bl[41] br[41] wl[486] vdd gnd cell_6t
Xbit_r487_c41 bl[41] br[41] wl[487] vdd gnd cell_6t
Xbit_r488_c41 bl[41] br[41] wl[488] vdd gnd cell_6t
Xbit_r489_c41 bl[41] br[41] wl[489] vdd gnd cell_6t
Xbit_r490_c41 bl[41] br[41] wl[490] vdd gnd cell_6t
Xbit_r491_c41 bl[41] br[41] wl[491] vdd gnd cell_6t
Xbit_r492_c41 bl[41] br[41] wl[492] vdd gnd cell_6t
Xbit_r493_c41 bl[41] br[41] wl[493] vdd gnd cell_6t
Xbit_r494_c41 bl[41] br[41] wl[494] vdd gnd cell_6t
Xbit_r495_c41 bl[41] br[41] wl[495] vdd gnd cell_6t
Xbit_r496_c41 bl[41] br[41] wl[496] vdd gnd cell_6t
Xbit_r497_c41 bl[41] br[41] wl[497] vdd gnd cell_6t
Xbit_r498_c41 bl[41] br[41] wl[498] vdd gnd cell_6t
Xbit_r499_c41 bl[41] br[41] wl[499] vdd gnd cell_6t
Xbit_r500_c41 bl[41] br[41] wl[500] vdd gnd cell_6t
Xbit_r501_c41 bl[41] br[41] wl[501] vdd gnd cell_6t
Xbit_r502_c41 bl[41] br[41] wl[502] vdd gnd cell_6t
Xbit_r503_c41 bl[41] br[41] wl[503] vdd gnd cell_6t
Xbit_r504_c41 bl[41] br[41] wl[504] vdd gnd cell_6t
Xbit_r505_c41 bl[41] br[41] wl[505] vdd gnd cell_6t
Xbit_r506_c41 bl[41] br[41] wl[506] vdd gnd cell_6t
Xbit_r507_c41 bl[41] br[41] wl[507] vdd gnd cell_6t
Xbit_r508_c41 bl[41] br[41] wl[508] vdd gnd cell_6t
Xbit_r509_c41 bl[41] br[41] wl[509] vdd gnd cell_6t
Xbit_r510_c41 bl[41] br[41] wl[510] vdd gnd cell_6t
Xbit_r511_c41 bl[41] br[41] wl[511] vdd gnd cell_6t
Xbit_r0_c42 bl[42] br[42] wl[0] vdd gnd cell_6t
Xbit_r1_c42 bl[42] br[42] wl[1] vdd gnd cell_6t
Xbit_r2_c42 bl[42] br[42] wl[2] vdd gnd cell_6t
Xbit_r3_c42 bl[42] br[42] wl[3] vdd gnd cell_6t
Xbit_r4_c42 bl[42] br[42] wl[4] vdd gnd cell_6t
Xbit_r5_c42 bl[42] br[42] wl[5] vdd gnd cell_6t
Xbit_r6_c42 bl[42] br[42] wl[6] vdd gnd cell_6t
Xbit_r7_c42 bl[42] br[42] wl[7] vdd gnd cell_6t
Xbit_r8_c42 bl[42] br[42] wl[8] vdd gnd cell_6t
Xbit_r9_c42 bl[42] br[42] wl[9] vdd gnd cell_6t
Xbit_r10_c42 bl[42] br[42] wl[10] vdd gnd cell_6t
Xbit_r11_c42 bl[42] br[42] wl[11] vdd gnd cell_6t
Xbit_r12_c42 bl[42] br[42] wl[12] vdd gnd cell_6t
Xbit_r13_c42 bl[42] br[42] wl[13] vdd gnd cell_6t
Xbit_r14_c42 bl[42] br[42] wl[14] vdd gnd cell_6t
Xbit_r15_c42 bl[42] br[42] wl[15] vdd gnd cell_6t
Xbit_r16_c42 bl[42] br[42] wl[16] vdd gnd cell_6t
Xbit_r17_c42 bl[42] br[42] wl[17] vdd gnd cell_6t
Xbit_r18_c42 bl[42] br[42] wl[18] vdd gnd cell_6t
Xbit_r19_c42 bl[42] br[42] wl[19] vdd gnd cell_6t
Xbit_r20_c42 bl[42] br[42] wl[20] vdd gnd cell_6t
Xbit_r21_c42 bl[42] br[42] wl[21] vdd gnd cell_6t
Xbit_r22_c42 bl[42] br[42] wl[22] vdd gnd cell_6t
Xbit_r23_c42 bl[42] br[42] wl[23] vdd gnd cell_6t
Xbit_r24_c42 bl[42] br[42] wl[24] vdd gnd cell_6t
Xbit_r25_c42 bl[42] br[42] wl[25] vdd gnd cell_6t
Xbit_r26_c42 bl[42] br[42] wl[26] vdd gnd cell_6t
Xbit_r27_c42 bl[42] br[42] wl[27] vdd gnd cell_6t
Xbit_r28_c42 bl[42] br[42] wl[28] vdd gnd cell_6t
Xbit_r29_c42 bl[42] br[42] wl[29] vdd gnd cell_6t
Xbit_r30_c42 bl[42] br[42] wl[30] vdd gnd cell_6t
Xbit_r31_c42 bl[42] br[42] wl[31] vdd gnd cell_6t
Xbit_r32_c42 bl[42] br[42] wl[32] vdd gnd cell_6t
Xbit_r33_c42 bl[42] br[42] wl[33] vdd gnd cell_6t
Xbit_r34_c42 bl[42] br[42] wl[34] vdd gnd cell_6t
Xbit_r35_c42 bl[42] br[42] wl[35] vdd gnd cell_6t
Xbit_r36_c42 bl[42] br[42] wl[36] vdd gnd cell_6t
Xbit_r37_c42 bl[42] br[42] wl[37] vdd gnd cell_6t
Xbit_r38_c42 bl[42] br[42] wl[38] vdd gnd cell_6t
Xbit_r39_c42 bl[42] br[42] wl[39] vdd gnd cell_6t
Xbit_r40_c42 bl[42] br[42] wl[40] vdd gnd cell_6t
Xbit_r41_c42 bl[42] br[42] wl[41] vdd gnd cell_6t
Xbit_r42_c42 bl[42] br[42] wl[42] vdd gnd cell_6t
Xbit_r43_c42 bl[42] br[42] wl[43] vdd gnd cell_6t
Xbit_r44_c42 bl[42] br[42] wl[44] vdd gnd cell_6t
Xbit_r45_c42 bl[42] br[42] wl[45] vdd gnd cell_6t
Xbit_r46_c42 bl[42] br[42] wl[46] vdd gnd cell_6t
Xbit_r47_c42 bl[42] br[42] wl[47] vdd gnd cell_6t
Xbit_r48_c42 bl[42] br[42] wl[48] vdd gnd cell_6t
Xbit_r49_c42 bl[42] br[42] wl[49] vdd gnd cell_6t
Xbit_r50_c42 bl[42] br[42] wl[50] vdd gnd cell_6t
Xbit_r51_c42 bl[42] br[42] wl[51] vdd gnd cell_6t
Xbit_r52_c42 bl[42] br[42] wl[52] vdd gnd cell_6t
Xbit_r53_c42 bl[42] br[42] wl[53] vdd gnd cell_6t
Xbit_r54_c42 bl[42] br[42] wl[54] vdd gnd cell_6t
Xbit_r55_c42 bl[42] br[42] wl[55] vdd gnd cell_6t
Xbit_r56_c42 bl[42] br[42] wl[56] vdd gnd cell_6t
Xbit_r57_c42 bl[42] br[42] wl[57] vdd gnd cell_6t
Xbit_r58_c42 bl[42] br[42] wl[58] vdd gnd cell_6t
Xbit_r59_c42 bl[42] br[42] wl[59] vdd gnd cell_6t
Xbit_r60_c42 bl[42] br[42] wl[60] vdd gnd cell_6t
Xbit_r61_c42 bl[42] br[42] wl[61] vdd gnd cell_6t
Xbit_r62_c42 bl[42] br[42] wl[62] vdd gnd cell_6t
Xbit_r63_c42 bl[42] br[42] wl[63] vdd gnd cell_6t
Xbit_r64_c42 bl[42] br[42] wl[64] vdd gnd cell_6t
Xbit_r65_c42 bl[42] br[42] wl[65] vdd gnd cell_6t
Xbit_r66_c42 bl[42] br[42] wl[66] vdd gnd cell_6t
Xbit_r67_c42 bl[42] br[42] wl[67] vdd gnd cell_6t
Xbit_r68_c42 bl[42] br[42] wl[68] vdd gnd cell_6t
Xbit_r69_c42 bl[42] br[42] wl[69] vdd gnd cell_6t
Xbit_r70_c42 bl[42] br[42] wl[70] vdd gnd cell_6t
Xbit_r71_c42 bl[42] br[42] wl[71] vdd gnd cell_6t
Xbit_r72_c42 bl[42] br[42] wl[72] vdd gnd cell_6t
Xbit_r73_c42 bl[42] br[42] wl[73] vdd gnd cell_6t
Xbit_r74_c42 bl[42] br[42] wl[74] vdd gnd cell_6t
Xbit_r75_c42 bl[42] br[42] wl[75] vdd gnd cell_6t
Xbit_r76_c42 bl[42] br[42] wl[76] vdd gnd cell_6t
Xbit_r77_c42 bl[42] br[42] wl[77] vdd gnd cell_6t
Xbit_r78_c42 bl[42] br[42] wl[78] vdd gnd cell_6t
Xbit_r79_c42 bl[42] br[42] wl[79] vdd gnd cell_6t
Xbit_r80_c42 bl[42] br[42] wl[80] vdd gnd cell_6t
Xbit_r81_c42 bl[42] br[42] wl[81] vdd gnd cell_6t
Xbit_r82_c42 bl[42] br[42] wl[82] vdd gnd cell_6t
Xbit_r83_c42 bl[42] br[42] wl[83] vdd gnd cell_6t
Xbit_r84_c42 bl[42] br[42] wl[84] vdd gnd cell_6t
Xbit_r85_c42 bl[42] br[42] wl[85] vdd gnd cell_6t
Xbit_r86_c42 bl[42] br[42] wl[86] vdd gnd cell_6t
Xbit_r87_c42 bl[42] br[42] wl[87] vdd gnd cell_6t
Xbit_r88_c42 bl[42] br[42] wl[88] vdd gnd cell_6t
Xbit_r89_c42 bl[42] br[42] wl[89] vdd gnd cell_6t
Xbit_r90_c42 bl[42] br[42] wl[90] vdd gnd cell_6t
Xbit_r91_c42 bl[42] br[42] wl[91] vdd gnd cell_6t
Xbit_r92_c42 bl[42] br[42] wl[92] vdd gnd cell_6t
Xbit_r93_c42 bl[42] br[42] wl[93] vdd gnd cell_6t
Xbit_r94_c42 bl[42] br[42] wl[94] vdd gnd cell_6t
Xbit_r95_c42 bl[42] br[42] wl[95] vdd gnd cell_6t
Xbit_r96_c42 bl[42] br[42] wl[96] vdd gnd cell_6t
Xbit_r97_c42 bl[42] br[42] wl[97] vdd gnd cell_6t
Xbit_r98_c42 bl[42] br[42] wl[98] vdd gnd cell_6t
Xbit_r99_c42 bl[42] br[42] wl[99] vdd gnd cell_6t
Xbit_r100_c42 bl[42] br[42] wl[100] vdd gnd cell_6t
Xbit_r101_c42 bl[42] br[42] wl[101] vdd gnd cell_6t
Xbit_r102_c42 bl[42] br[42] wl[102] vdd gnd cell_6t
Xbit_r103_c42 bl[42] br[42] wl[103] vdd gnd cell_6t
Xbit_r104_c42 bl[42] br[42] wl[104] vdd gnd cell_6t
Xbit_r105_c42 bl[42] br[42] wl[105] vdd gnd cell_6t
Xbit_r106_c42 bl[42] br[42] wl[106] vdd gnd cell_6t
Xbit_r107_c42 bl[42] br[42] wl[107] vdd gnd cell_6t
Xbit_r108_c42 bl[42] br[42] wl[108] vdd gnd cell_6t
Xbit_r109_c42 bl[42] br[42] wl[109] vdd gnd cell_6t
Xbit_r110_c42 bl[42] br[42] wl[110] vdd gnd cell_6t
Xbit_r111_c42 bl[42] br[42] wl[111] vdd gnd cell_6t
Xbit_r112_c42 bl[42] br[42] wl[112] vdd gnd cell_6t
Xbit_r113_c42 bl[42] br[42] wl[113] vdd gnd cell_6t
Xbit_r114_c42 bl[42] br[42] wl[114] vdd gnd cell_6t
Xbit_r115_c42 bl[42] br[42] wl[115] vdd gnd cell_6t
Xbit_r116_c42 bl[42] br[42] wl[116] vdd gnd cell_6t
Xbit_r117_c42 bl[42] br[42] wl[117] vdd gnd cell_6t
Xbit_r118_c42 bl[42] br[42] wl[118] vdd gnd cell_6t
Xbit_r119_c42 bl[42] br[42] wl[119] vdd gnd cell_6t
Xbit_r120_c42 bl[42] br[42] wl[120] vdd gnd cell_6t
Xbit_r121_c42 bl[42] br[42] wl[121] vdd gnd cell_6t
Xbit_r122_c42 bl[42] br[42] wl[122] vdd gnd cell_6t
Xbit_r123_c42 bl[42] br[42] wl[123] vdd gnd cell_6t
Xbit_r124_c42 bl[42] br[42] wl[124] vdd gnd cell_6t
Xbit_r125_c42 bl[42] br[42] wl[125] vdd gnd cell_6t
Xbit_r126_c42 bl[42] br[42] wl[126] vdd gnd cell_6t
Xbit_r127_c42 bl[42] br[42] wl[127] vdd gnd cell_6t
Xbit_r128_c42 bl[42] br[42] wl[128] vdd gnd cell_6t
Xbit_r129_c42 bl[42] br[42] wl[129] vdd gnd cell_6t
Xbit_r130_c42 bl[42] br[42] wl[130] vdd gnd cell_6t
Xbit_r131_c42 bl[42] br[42] wl[131] vdd gnd cell_6t
Xbit_r132_c42 bl[42] br[42] wl[132] vdd gnd cell_6t
Xbit_r133_c42 bl[42] br[42] wl[133] vdd gnd cell_6t
Xbit_r134_c42 bl[42] br[42] wl[134] vdd gnd cell_6t
Xbit_r135_c42 bl[42] br[42] wl[135] vdd gnd cell_6t
Xbit_r136_c42 bl[42] br[42] wl[136] vdd gnd cell_6t
Xbit_r137_c42 bl[42] br[42] wl[137] vdd gnd cell_6t
Xbit_r138_c42 bl[42] br[42] wl[138] vdd gnd cell_6t
Xbit_r139_c42 bl[42] br[42] wl[139] vdd gnd cell_6t
Xbit_r140_c42 bl[42] br[42] wl[140] vdd gnd cell_6t
Xbit_r141_c42 bl[42] br[42] wl[141] vdd gnd cell_6t
Xbit_r142_c42 bl[42] br[42] wl[142] vdd gnd cell_6t
Xbit_r143_c42 bl[42] br[42] wl[143] vdd gnd cell_6t
Xbit_r144_c42 bl[42] br[42] wl[144] vdd gnd cell_6t
Xbit_r145_c42 bl[42] br[42] wl[145] vdd gnd cell_6t
Xbit_r146_c42 bl[42] br[42] wl[146] vdd gnd cell_6t
Xbit_r147_c42 bl[42] br[42] wl[147] vdd gnd cell_6t
Xbit_r148_c42 bl[42] br[42] wl[148] vdd gnd cell_6t
Xbit_r149_c42 bl[42] br[42] wl[149] vdd gnd cell_6t
Xbit_r150_c42 bl[42] br[42] wl[150] vdd gnd cell_6t
Xbit_r151_c42 bl[42] br[42] wl[151] vdd gnd cell_6t
Xbit_r152_c42 bl[42] br[42] wl[152] vdd gnd cell_6t
Xbit_r153_c42 bl[42] br[42] wl[153] vdd gnd cell_6t
Xbit_r154_c42 bl[42] br[42] wl[154] vdd gnd cell_6t
Xbit_r155_c42 bl[42] br[42] wl[155] vdd gnd cell_6t
Xbit_r156_c42 bl[42] br[42] wl[156] vdd gnd cell_6t
Xbit_r157_c42 bl[42] br[42] wl[157] vdd gnd cell_6t
Xbit_r158_c42 bl[42] br[42] wl[158] vdd gnd cell_6t
Xbit_r159_c42 bl[42] br[42] wl[159] vdd gnd cell_6t
Xbit_r160_c42 bl[42] br[42] wl[160] vdd gnd cell_6t
Xbit_r161_c42 bl[42] br[42] wl[161] vdd gnd cell_6t
Xbit_r162_c42 bl[42] br[42] wl[162] vdd gnd cell_6t
Xbit_r163_c42 bl[42] br[42] wl[163] vdd gnd cell_6t
Xbit_r164_c42 bl[42] br[42] wl[164] vdd gnd cell_6t
Xbit_r165_c42 bl[42] br[42] wl[165] vdd gnd cell_6t
Xbit_r166_c42 bl[42] br[42] wl[166] vdd gnd cell_6t
Xbit_r167_c42 bl[42] br[42] wl[167] vdd gnd cell_6t
Xbit_r168_c42 bl[42] br[42] wl[168] vdd gnd cell_6t
Xbit_r169_c42 bl[42] br[42] wl[169] vdd gnd cell_6t
Xbit_r170_c42 bl[42] br[42] wl[170] vdd gnd cell_6t
Xbit_r171_c42 bl[42] br[42] wl[171] vdd gnd cell_6t
Xbit_r172_c42 bl[42] br[42] wl[172] vdd gnd cell_6t
Xbit_r173_c42 bl[42] br[42] wl[173] vdd gnd cell_6t
Xbit_r174_c42 bl[42] br[42] wl[174] vdd gnd cell_6t
Xbit_r175_c42 bl[42] br[42] wl[175] vdd gnd cell_6t
Xbit_r176_c42 bl[42] br[42] wl[176] vdd gnd cell_6t
Xbit_r177_c42 bl[42] br[42] wl[177] vdd gnd cell_6t
Xbit_r178_c42 bl[42] br[42] wl[178] vdd gnd cell_6t
Xbit_r179_c42 bl[42] br[42] wl[179] vdd gnd cell_6t
Xbit_r180_c42 bl[42] br[42] wl[180] vdd gnd cell_6t
Xbit_r181_c42 bl[42] br[42] wl[181] vdd gnd cell_6t
Xbit_r182_c42 bl[42] br[42] wl[182] vdd gnd cell_6t
Xbit_r183_c42 bl[42] br[42] wl[183] vdd gnd cell_6t
Xbit_r184_c42 bl[42] br[42] wl[184] vdd gnd cell_6t
Xbit_r185_c42 bl[42] br[42] wl[185] vdd gnd cell_6t
Xbit_r186_c42 bl[42] br[42] wl[186] vdd gnd cell_6t
Xbit_r187_c42 bl[42] br[42] wl[187] vdd gnd cell_6t
Xbit_r188_c42 bl[42] br[42] wl[188] vdd gnd cell_6t
Xbit_r189_c42 bl[42] br[42] wl[189] vdd gnd cell_6t
Xbit_r190_c42 bl[42] br[42] wl[190] vdd gnd cell_6t
Xbit_r191_c42 bl[42] br[42] wl[191] vdd gnd cell_6t
Xbit_r192_c42 bl[42] br[42] wl[192] vdd gnd cell_6t
Xbit_r193_c42 bl[42] br[42] wl[193] vdd gnd cell_6t
Xbit_r194_c42 bl[42] br[42] wl[194] vdd gnd cell_6t
Xbit_r195_c42 bl[42] br[42] wl[195] vdd gnd cell_6t
Xbit_r196_c42 bl[42] br[42] wl[196] vdd gnd cell_6t
Xbit_r197_c42 bl[42] br[42] wl[197] vdd gnd cell_6t
Xbit_r198_c42 bl[42] br[42] wl[198] vdd gnd cell_6t
Xbit_r199_c42 bl[42] br[42] wl[199] vdd gnd cell_6t
Xbit_r200_c42 bl[42] br[42] wl[200] vdd gnd cell_6t
Xbit_r201_c42 bl[42] br[42] wl[201] vdd gnd cell_6t
Xbit_r202_c42 bl[42] br[42] wl[202] vdd gnd cell_6t
Xbit_r203_c42 bl[42] br[42] wl[203] vdd gnd cell_6t
Xbit_r204_c42 bl[42] br[42] wl[204] vdd gnd cell_6t
Xbit_r205_c42 bl[42] br[42] wl[205] vdd gnd cell_6t
Xbit_r206_c42 bl[42] br[42] wl[206] vdd gnd cell_6t
Xbit_r207_c42 bl[42] br[42] wl[207] vdd gnd cell_6t
Xbit_r208_c42 bl[42] br[42] wl[208] vdd gnd cell_6t
Xbit_r209_c42 bl[42] br[42] wl[209] vdd gnd cell_6t
Xbit_r210_c42 bl[42] br[42] wl[210] vdd gnd cell_6t
Xbit_r211_c42 bl[42] br[42] wl[211] vdd gnd cell_6t
Xbit_r212_c42 bl[42] br[42] wl[212] vdd gnd cell_6t
Xbit_r213_c42 bl[42] br[42] wl[213] vdd gnd cell_6t
Xbit_r214_c42 bl[42] br[42] wl[214] vdd gnd cell_6t
Xbit_r215_c42 bl[42] br[42] wl[215] vdd gnd cell_6t
Xbit_r216_c42 bl[42] br[42] wl[216] vdd gnd cell_6t
Xbit_r217_c42 bl[42] br[42] wl[217] vdd gnd cell_6t
Xbit_r218_c42 bl[42] br[42] wl[218] vdd gnd cell_6t
Xbit_r219_c42 bl[42] br[42] wl[219] vdd gnd cell_6t
Xbit_r220_c42 bl[42] br[42] wl[220] vdd gnd cell_6t
Xbit_r221_c42 bl[42] br[42] wl[221] vdd gnd cell_6t
Xbit_r222_c42 bl[42] br[42] wl[222] vdd gnd cell_6t
Xbit_r223_c42 bl[42] br[42] wl[223] vdd gnd cell_6t
Xbit_r224_c42 bl[42] br[42] wl[224] vdd gnd cell_6t
Xbit_r225_c42 bl[42] br[42] wl[225] vdd gnd cell_6t
Xbit_r226_c42 bl[42] br[42] wl[226] vdd gnd cell_6t
Xbit_r227_c42 bl[42] br[42] wl[227] vdd gnd cell_6t
Xbit_r228_c42 bl[42] br[42] wl[228] vdd gnd cell_6t
Xbit_r229_c42 bl[42] br[42] wl[229] vdd gnd cell_6t
Xbit_r230_c42 bl[42] br[42] wl[230] vdd gnd cell_6t
Xbit_r231_c42 bl[42] br[42] wl[231] vdd gnd cell_6t
Xbit_r232_c42 bl[42] br[42] wl[232] vdd gnd cell_6t
Xbit_r233_c42 bl[42] br[42] wl[233] vdd gnd cell_6t
Xbit_r234_c42 bl[42] br[42] wl[234] vdd gnd cell_6t
Xbit_r235_c42 bl[42] br[42] wl[235] vdd gnd cell_6t
Xbit_r236_c42 bl[42] br[42] wl[236] vdd gnd cell_6t
Xbit_r237_c42 bl[42] br[42] wl[237] vdd gnd cell_6t
Xbit_r238_c42 bl[42] br[42] wl[238] vdd gnd cell_6t
Xbit_r239_c42 bl[42] br[42] wl[239] vdd gnd cell_6t
Xbit_r240_c42 bl[42] br[42] wl[240] vdd gnd cell_6t
Xbit_r241_c42 bl[42] br[42] wl[241] vdd gnd cell_6t
Xbit_r242_c42 bl[42] br[42] wl[242] vdd gnd cell_6t
Xbit_r243_c42 bl[42] br[42] wl[243] vdd gnd cell_6t
Xbit_r244_c42 bl[42] br[42] wl[244] vdd gnd cell_6t
Xbit_r245_c42 bl[42] br[42] wl[245] vdd gnd cell_6t
Xbit_r246_c42 bl[42] br[42] wl[246] vdd gnd cell_6t
Xbit_r247_c42 bl[42] br[42] wl[247] vdd gnd cell_6t
Xbit_r248_c42 bl[42] br[42] wl[248] vdd gnd cell_6t
Xbit_r249_c42 bl[42] br[42] wl[249] vdd gnd cell_6t
Xbit_r250_c42 bl[42] br[42] wl[250] vdd gnd cell_6t
Xbit_r251_c42 bl[42] br[42] wl[251] vdd gnd cell_6t
Xbit_r252_c42 bl[42] br[42] wl[252] vdd gnd cell_6t
Xbit_r253_c42 bl[42] br[42] wl[253] vdd gnd cell_6t
Xbit_r254_c42 bl[42] br[42] wl[254] vdd gnd cell_6t
Xbit_r255_c42 bl[42] br[42] wl[255] vdd gnd cell_6t
Xbit_r256_c42 bl[42] br[42] wl[256] vdd gnd cell_6t
Xbit_r257_c42 bl[42] br[42] wl[257] vdd gnd cell_6t
Xbit_r258_c42 bl[42] br[42] wl[258] vdd gnd cell_6t
Xbit_r259_c42 bl[42] br[42] wl[259] vdd gnd cell_6t
Xbit_r260_c42 bl[42] br[42] wl[260] vdd gnd cell_6t
Xbit_r261_c42 bl[42] br[42] wl[261] vdd gnd cell_6t
Xbit_r262_c42 bl[42] br[42] wl[262] vdd gnd cell_6t
Xbit_r263_c42 bl[42] br[42] wl[263] vdd gnd cell_6t
Xbit_r264_c42 bl[42] br[42] wl[264] vdd gnd cell_6t
Xbit_r265_c42 bl[42] br[42] wl[265] vdd gnd cell_6t
Xbit_r266_c42 bl[42] br[42] wl[266] vdd gnd cell_6t
Xbit_r267_c42 bl[42] br[42] wl[267] vdd gnd cell_6t
Xbit_r268_c42 bl[42] br[42] wl[268] vdd gnd cell_6t
Xbit_r269_c42 bl[42] br[42] wl[269] vdd gnd cell_6t
Xbit_r270_c42 bl[42] br[42] wl[270] vdd gnd cell_6t
Xbit_r271_c42 bl[42] br[42] wl[271] vdd gnd cell_6t
Xbit_r272_c42 bl[42] br[42] wl[272] vdd gnd cell_6t
Xbit_r273_c42 bl[42] br[42] wl[273] vdd gnd cell_6t
Xbit_r274_c42 bl[42] br[42] wl[274] vdd gnd cell_6t
Xbit_r275_c42 bl[42] br[42] wl[275] vdd gnd cell_6t
Xbit_r276_c42 bl[42] br[42] wl[276] vdd gnd cell_6t
Xbit_r277_c42 bl[42] br[42] wl[277] vdd gnd cell_6t
Xbit_r278_c42 bl[42] br[42] wl[278] vdd gnd cell_6t
Xbit_r279_c42 bl[42] br[42] wl[279] vdd gnd cell_6t
Xbit_r280_c42 bl[42] br[42] wl[280] vdd gnd cell_6t
Xbit_r281_c42 bl[42] br[42] wl[281] vdd gnd cell_6t
Xbit_r282_c42 bl[42] br[42] wl[282] vdd gnd cell_6t
Xbit_r283_c42 bl[42] br[42] wl[283] vdd gnd cell_6t
Xbit_r284_c42 bl[42] br[42] wl[284] vdd gnd cell_6t
Xbit_r285_c42 bl[42] br[42] wl[285] vdd gnd cell_6t
Xbit_r286_c42 bl[42] br[42] wl[286] vdd gnd cell_6t
Xbit_r287_c42 bl[42] br[42] wl[287] vdd gnd cell_6t
Xbit_r288_c42 bl[42] br[42] wl[288] vdd gnd cell_6t
Xbit_r289_c42 bl[42] br[42] wl[289] vdd gnd cell_6t
Xbit_r290_c42 bl[42] br[42] wl[290] vdd gnd cell_6t
Xbit_r291_c42 bl[42] br[42] wl[291] vdd gnd cell_6t
Xbit_r292_c42 bl[42] br[42] wl[292] vdd gnd cell_6t
Xbit_r293_c42 bl[42] br[42] wl[293] vdd gnd cell_6t
Xbit_r294_c42 bl[42] br[42] wl[294] vdd gnd cell_6t
Xbit_r295_c42 bl[42] br[42] wl[295] vdd gnd cell_6t
Xbit_r296_c42 bl[42] br[42] wl[296] vdd gnd cell_6t
Xbit_r297_c42 bl[42] br[42] wl[297] vdd gnd cell_6t
Xbit_r298_c42 bl[42] br[42] wl[298] vdd gnd cell_6t
Xbit_r299_c42 bl[42] br[42] wl[299] vdd gnd cell_6t
Xbit_r300_c42 bl[42] br[42] wl[300] vdd gnd cell_6t
Xbit_r301_c42 bl[42] br[42] wl[301] vdd gnd cell_6t
Xbit_r302_c42 bl[42] br[42] wl[302] vdd gnd cell_6t
Xbit_r303_c42 bl[42] br[42] wl[303] vdd gnd cell_6t
Xbit_r304_c42 bl[42] br[42] wl[304] vdd gnd cell_6t
Xbit_r305_c42 bl[42] br[42] wl[305] vdd gnd cell_6t
Xbit_r306_c42 bl[42] br[42] wl[306] vdd gnd cell_6t
Xbit_r307_c42 bl[42] br[42] wl[307] vdd gnd cell_6t
Xbit_r308_c42 bl[42] br[42] wl[308] vdd gnd cell_6t
Xbit_r309_c42 bl[42] br[42] wl[309] vdd gnd cell_6t
Xbit_r310_c42 bl[42] br[42] wl[310] vdd gnd cell_6t
Xbit_r311_c42 bl[42] br[42] wl[311] vdd gnd cell_6t
Xbit_r312_c42 bl[42] br[42] wl[312] vdd gnd cell_6t
Xbit_r313_c42 bl[42] br[42] wl[313] vdd gnd cell_6t
Xbit_r314_c42 bl[42] br[42] wl[314] vdd gnd cell_6t
Xbit_r315_c42 bl[42] br[42] wl[315] vdd gnd cell_6t
Xbit_r316_c42 bl[42] br[42] wl[316] vdd gnd cell_6t
Xbit_r317_c42 bl[42] br[42] wl[317] vdd gnd cell_6t
Xbit_r318_c42 bl[42] br[42] wl[318] vdd gnd cell_6t
Xbit_r319_c42 bl[42] br[42] wl[319] vdd gnd cell_6t
Xbit_r320_c42 bl[42] br[42] wl[320] vdd gnd cell_6t
Xbit_r321_c42 bl[42] br[42] wl[321] vdd gnd cell_6t
Xbit_r322_c42 bl[42] br[42] wl[322] vdd gnd cell_6t
Xbit_r323_c42 bl[42] br[42] wl[323] vdd gnd cell_6t
Xbit_r324_c42 bl[42] br[42] wl[324] vdd gnd cell_6t
Xbit_r325_c42 bl[42] br[42] wl[325] vdd gnd cell_6t
Xbit_r326_c42 bl[42] br[42] wl[326] vdd gnd cell_6t
Xbit_r327_c42 bl[42] br[42] wl[327] vdd gnd cell_6t
Xbit_r328_c42 bl[42] br[42] wl[328] vdd gnd cell_6t
Xbit_r329_c42 bl[42] br[42] wl[329] vdd gnd cell_6t
Xbit_r330_c42 bl[42] br[42] wl[330] vdd gnd cell_6t
Xbit_r331_c42 bl[42] br[42] wl[331] vdd gnd cell_6t
Xbit_r332_c42 bl[42] br[42] wl[332] vdd gnd cell_6t
Xbit_r333_c42 bl[42] br[42] wl[333] vdd gnd cell_6t
Xbit_r334_c42 bl[42] br[42] wl[334] vdd gnd cell_6t
Xbit_r335_c42 bl[42] br[42] wl[335] vdd gnd cell_6t
Xbit_r336_c42 bl[42] br[42] wl[336] vdd gnd cell_6t
Xbit_r337_c42 bl[42] br[42] wl[337] vdd gnd cell_6t
Xbit_r338_c42 bl[42] br[42] wl[338] vdd gnd cell_6t
Xbit_r339_c42 bl[42] br[42] wl[339] vdd gnd cell_6t
Xbit_r340_c42 bl[42] br[42] wl[340] vdd gnd cell_6t
Xbit_r341_c42 bl[42] br[42] wl[341] vdd gnd cell_6t
Xbit_r342_c42 bl[42] br[42] wl[342] vdd gnd cell_6t
Xbit_r343_c42 bl[42] br[42] wl[343] vdd gnd cell_6t
Xbit_r344_c42 bl[42] br[42] wl[344] vdd gnd cell_6t
Xbit_r345_c42 bl[42] br[42] wl[345] vdd gnd cell_6t
Xbit_r346_c42 bl[42] br[42] wl[346] vdd gnd cell_6t
Xbit_r347_c42 bl[42] br[42] wl[347] vdd gnd cell_6t
Xbit_r348_c42 bl[42] br[42] wl[348] vdd gnd cell_6t
Xbit_r349_c42 bl[42] br[42] wl[349] vdd gnd cell_6t
Xbit_r350_c42 bl[42] br[42] wl[350] vdd gnd cell_6t
Xbit_r351_c42 bl[42] br[42] wl[351] vdd gnd cell_6t
Xbit_r352_c42 bl[42] br[42] wl[352] vdd gnd cell_6t
Xbit_r353_c42 bl[42] br[42] wl[353] vdd gnd cell_6t
Xbit_r354_c42 bl[42] br[42] wl[354] vdd gnd cell_6t
Xbit_r355_c42 bl[42] br[42] wl[355] vdd gnd cell_6t
Xbit_r356_c42 bl[42] br[42] wl[356] vdd gnd cell_6t
Xbit_r357_c42 bl[42] br[42] wl[357] vdd gnd cell_6t
Xbit_r358_c42 bl[42] br[42] wl[358] vdd gnd cell_6t
Xbit_r359_c42 bl[42] br[42] wl[359] vdd gnd cell_6t
Xbit_r360_c42 bl[42] br[42] wl[360] vdd gnd cell_6t
Xbit_r361_c42 bl[42] br[42] wl[361] vdd gnd cell_6t
Xbit_r362_c42 bl[42] br[42] wl[362] vdd gnd cell_6t
Xbit_r363_c42 bl[42] br[42] wl[363] vdd gnd cell_6t
Xbit_r364_c42 bl[42] br[42] wl[364] vdd gnd cell_6t
Xbit_r365_c42 bl[42] br[42] wl[365] vdd gnd cell_6t
Xbit_r366_c42 bl[42] br[42] wl[366] vdd gnd cell_6t
Xbit_r367_c42 bl[42] br[42] wl[367] vdd gnd cell_6t
Xbit_r368_c42 bl[42] br[42] wl[368] vdd gnd cell_6t
Xbit_r369_c42 bl[42] br[42] wl[369] vdd gnd cell_6t
Xbit_r370_c42 bl[42] br[42] wl[370] vdd gnd cell_6t
Xbit_r371_c42 bl[42] br[42] wl[371] vdd gnd cell_6t
Xbit_r372_c42 bl[42] br[42] wl[372] vdd gnd cell_6t
Xbit_r373_c42 bl[42] br[42] wl[373] vdd gnd cell_6t
Xbit_r374_c42 bl[42] br[42] wl[374] vdd gnd cell_6t
Xbit_r375_c42 bl[42] br[42] wl[375] vdd gnd cell_6t
Xbit_r376_c42 bl[42] br[42] wl[376] vdd gnd cell_6t
Xbit_r377_c42 bl[42] br[42] wl[377] vdd gnd cell_6t
Xbit_r378_c42 bl[42] br[42] wl[378] vdd gnd cell_6t
Xbit_r379_c42 bl[42] br[42] wl[379] vdd gnd cell_6t
Xbit_r380_c42 bl[42] br[42] wl[380] vdd gnd cell_6t
Xbit_r381_c42 bl[42] br[42] wl[381] vdd gnd cell_6t
Xbit_r382_c42 bl[42] br[42] wl[382] vdd gnd cell_6t
Xbit_r383_c42 bl[42] br[42] wl[383] vdd gnd cell_6t
Xbit_r384_c42 bl[42] br[42] wl[384] vdd gnd cell_6t
Xbit_r385_c42 bl[42] br[42] wl[385] vdd gnd cell_6t
Xbit_r386_c42 bl[42] br[42] wl[386] vdd gnd cell_6t
Xbit_r387_c42 bl[42] br[42] wl[387] vdd gnd cell_6t
Xbit_r388_c42 bl[42] br[42] wl[388] vdd gnd cell_6t
Xbit_r389_c42 bl[42] br[42] wl[389] vdd gnd cell_6t
Xbit_r390_c42 bl[42] br[42] wl[390] vdd gnd cell_6t
Xbit_r391_c42 bl[42] br[42] wl[391] vdd gnd cell_6t
Xbit_r392_c42 bl[42] br[42] wl[392] vdd gnd cell_6t
Xbit_r393_c42 bl[42] br[42] wl[393] vdd gnd cell_6t
Xbit_r394_c42 bl[42] br[42] wl[394] vdd gnd cell_6t
Xbit_r395_c42 bl[42] br[42] wl[395] vdd gnd cell_6t
Xbit_r396_c42 bl[42] br[42] wl[396] vdd gnd cell_6t
Xbit_r397_c42 bl[42] br[42] wl[397] vdd gnd cell_6t
Xbit_r398_c42 bl[42] br[42] wl[398] vdd gnd cell_6t
Xbit_r399_c42 bl[42] br[42] wl[399] vdd gnd cell_6t
Xbit_r400_c42 bl[42] br[42] wl[400] vdd gnd cell_6t
Xbit_r401_c42 bl[42] br[42] wl[401] vdd gnd cell_6t
Xbit_r402_c42 bl[42] br[42] wl[402] vdd gnd cell_6t
Xbit_r403_c42 bl[42] br[42] wl[403] vdd gnd cell_6t
Xbit_r404_c42 bl[42] br[42] wl[404] vdd gnd cell_6t
Xbit_r405_c42 bl[42] br[42] wl[405] vdd gnd cell_6t
Xbit_r406_c42 bl[42] br[42] wl[406] vdd gnd cell_6t
Xbit_r407_c42 bl[42] br[42] wl[407] vdd gnd cell_6t
Xbit_r408_c42 bl[42] br[42] wl[408] vdd gnd cell_6t
Xbit_r409_c42 bl[42] br[42] wl[409] vdd gnd cell_6t
Xbit_r410_c42 bl[42] br[42] wl[410] vdd gnd cell_6t
Xbit_r411_c42 bl[42] br[42] wl[411] vdd gnd cell_6t
Xbit_r412_c42 bl[42] br[42] wl[412] vdd gnd cell_6t
Xbit_r413_c42 bl[42] br[42] wl[413] vdd gnd cell_6t
Xbit_r414_c42 bl[42] br[42] wl[414] vdd gnd cell_6t
Xbit_r415_c42 bl[42] br[42] wl[415] vdd gnd cell_6t
Xbit_r416_c42 bl[42] br[42] wl[416] vdd gnd cell_6t
Xbit_r417_c42 bl[42] br[42] wl[417] vdd gnd cell_6t
Xbit_r418_c42 bl[42] br[42] wl[418] vdd gnd cell_6t
Xbit_r419_c42 bl[42] br[42] wl[419] vdd gnd cell_6t
Xbit_r420_c42 bl[42] br[42] wl[420] vdd gnd cell_6t
Xbit_r421_c42 bl[42] br[42] wl[421] vdd gnd cell_6t
Xbit_r422_c42 bl[42] br[42] wl[422] vdd gnd cell_6t
Xbit_r423_c42 bl[42] br[42] wl[423] vdd gnd cell_6t
Xbit_r424_c42 bl[42] br[42] wl[424] vdd gnd cell_6t
Xbit_r425_c42 bl[42] br[42] wl[425] vdd gnd cell_6t
Xbit_r426_c42 bl[42] br[42] wl[426] vdd gnd cell_6t
Xbit_r427_c42 bl[42] br[42] wl[427] vdd gnd cell_6t
Xbit_r428_c42 bl[42] br[42] wl[428] vdd gnd cell_6t
Xbit_r429_c42 bl[42] br[42] wl[429] vdd gnd cell_6t
Xbit_r430_c42 bl[42] br[42] wl[430] vdd gnd cell_6t
Xbit_r431_c42 bl[42] br[42] wl[431] vdd gnd cell_6t
Xbit_r432_c42 bl[42] br[42] wl[432] vdd gnd cell_6t
Xbit_r433_c42 bl[42] br[42] wl[433] vdd gnd cell_6t
Xbit_r434_c42 bl[42] br[42] wl[434] vdd gnd cell_6t
Xbit_r435_c42 bl[42] br[42] wl[435] vdd gnd cell_6t
Xbit_r436_c42 bl[42] br[42] wl[436] vdd gnd cell_6t
Xbit_r437_c42 bl[42] br[42] wl[437] vdd gnd cell_6t
Xbit_r438_c42 bl[42] br[42] wl[438] vdd gnd cell_6t
Xbit_r439_c42 bl[42] br[42] wl[439] vdd gnd cell_6t
Xbit_r440_c42 bl[42] br[42] wl[440] vdd gnd cell_6t
Xbit_r441_c42 bl[42] br[42] wl[441] vdd gnd cell_6t
Xbit_r442_c42 bl[42] br[42] wl[442] vdd gnd cell_6t
Xbit_r443_c42 bl[42] br[42] wl[443] vdd gnd cell_6t
Xbit_r444_c42 bl[42] br[42] wl[444] vdd gnd cell_6t
Xbit_r445_c42 bl[42] br[42] wl[445] vdd gnd cell_6t
Xbit_r446_c42 bl[42] br[42] wl[446] vdd gnd cell_6t
Xbit_r447_c42 bl[42] br[42] wl[447] vdd gnd cell_6t
Xbit_r448_c42 bl[42] br[42] wl[448] vdd gnd cell_6t
Xbit_r449_c42 bl[42] br[42] wl[449] vdd gnd cell_6t
Xbit_r450_c42 bl[42] br[42] wl[450] vdd gnd cell_6t
Xbit_r451_c42 bl[42] br[42] wl[451] vdd gnd cell_6t
Xbit_r452_c42 bl[42] br[42] wl[452] vdd gnd cell_6t
Xbit_r453_c42 bl[42] br[42] wl[453] vdd gnd cell_6t
Xbit_r454_c42 bl[42] br[42] wl[454] vdd gnd cell_6t
Xbit_r455_c42 bl[42] br[42] wl[455] vdd gnd cell_6t
Xbit_r456_c42 bl[42] br[42] wl[456] vdd gnd cell_6t
Xbit_r457_c42 bl[42] br[42] wl[457] vdd gnd cell_6t
Xbit_r458_c42 bl[42] br[42] wl[458] vdd gnd cell_6t
Xbit_r459_c42 bl[42] br[42] wl[459] vdd gnd cell_6t
Xbit_r460_c42 bl[42] br[42] wl[460] vdd gnd cell_6t
Xbit_r461_c42 bl[42] br[42] wl[461] vdd gnd cell_6t
Xbit_r462_c42 bl[42] br[42] wl[462] vdd gnd cell_6t
Xbit_r463_c42 bl[42] br[42] wl[463] vdd gnd cell_6t
Xbit_r464_c42 bl[42] br[42] wl[464] vdd gnd cell_6t
Xbit_r465_c42 bl[42] br[42] wl[465] vdd gnd cell_6t
Xbit_r466_c42 bl[42] br[42] wl[466] vdd gnd cell_6t
Xbit_r467_c42 bl[42] br[42] wl[467] vdd gnd cell_6t
Xbit_r468_c42 bl[42] br[42] wl[468] vdd gnd cell_6t
Xbit_r469_c42 bl[42] br[42] wl[469] vdd gnd cell_6t
Xbit_r470_c42 bl[42] br[42] wl[470] vdd gnd cell_6t
Xbit_r471_c42 bl[42] br[42] wl[471] vdd gnd cell_6t
Xbit_r472_c42 bl[42] br[42] wl[472] vdd gnd cell_6t
Xbit_r473_c42 bl[42] br[42] wl[473] vdd gnd cell_6t
Xbit_r474_c42 bl[42] br[42] wl[474] vdd gnd cell_6t
Xbit_r475_c42 bl[42] br[42] wl[475] vdd gnd cell_6t
Xbit_r476_c42 bl[42] br[42] wl[476] vdd gnd cell_6t
Xbit_r477_c42 bl[42] br[42] wl[477] vdd gnd cell_6t
Xbit_r478_c42 bl[42] br[42] wl[478] vdd gnd cell_6t
Xbit_r479_c42 bl[42] br[42] wl[479] vdd gnd cell_6t
Xbit_r480_c42 bl[42] br[42] wl[480] vdd gnd cell_6t
Xbit_r481_c42 bl[42] br[42] wl[481] vdd gnd cell_6t
Xbit_r482_c42 bl[42] br[42] wl[482] vdd gnd cell_6t
Xbit_r483_c42 bl[42] br[42] wl[483] vdd gnd cell_6t
Xbit_r484_c42 bl[42] br[42] wl[484] vdd gnd cell_6t
Xbit_r485_c42 bl[42] br[42] wl[485] vdd gnd cell_6t
Xbit_r486_c42 bl[42] br[42] wl[486] vdd gnd cell_6t
Xbit_r487_c42 bl[42] br[42] wl[487] vdd gnd cell_6t
Xbit_r488_c42 bl[42] br[42] wl[488] vdd gnd cell_6t
Xbit_r489_c42 bl[42] br[42] wl[489] vdd gnd cell_6t
Xbit_r490_c42 bl[42] br[42] wl[490] vdd gnd cell_6t
Xbit_r491_c42 bl[42] br[42] wl[491] vdd gnd cell_6t
Xbit_r492_c42 bl[42] br[42] wl[492] vdd gnd cell_6t
Xbit_r493_c42 bl[42] br[42] wl[493] vdd gnd cell_6t
Xbit_r494_c42 bl[42] br[42] wl[494] vdd gnd cell_6t
Xbit_r495_c42 bl[42] br[42] wl[495] vdd gnd cell_6t
Xbit_r496_c42 bl[42] br[42] wl[496] vdd gnd cell_6t
Xbit_r497_c42 bl[42] br[42] wl[497] vdd gnd cell_6t
Xbit_r498_c42 bl[42] br[42] wl[498] vdd gnd cell_6t
Xbit_r499_c42 bl[42] br[42] wl[499] vdd gnd cell_6t
Xbit_r500_c42 bl[42] br[42] wl[500] vdd gnd cell_6t
Xbit_r501_c42 bl[42] br[42] wl[501] vdd gnd cell_6t
Xbit_r502_c42 bl[42] br[42] wl[502] vdd gnd cell_6t
Xbit_r503_c42 bl[42] br[42] wl[503] vdd gnd cell_6t
Xbit_r504_c42 bl[42] br[42] wl[504] vdd gnd cell_6t
Xbit_r505_c42 bl[42] br[42] wl[505] vdd gnd cell_6t
Xbit_r506_c42 bl[42] br[42] wl[506] vdd gnd cell_6t
Xbit_r507_c42 bl[42] br[42] wl[507] vdd gnd cell_6t
Xbit_r508_c42 bl[42] br[42] wl[508] vdd gnd cell_6t
Xbit_r509_c42 bl[42] br[42] wl[509] vdd gnd cell_6t
Xbit_r510_c42 bl[42] br[42] wl[510] vdd gnd cell_6t
Xbit_r511_c42 bl[42] br[42] wl[511] vdd gnd cell_6t
Xbit_r0_c43 bl[43] br[43] wl[0] vdd gnd cell_6t
Xbit_r1_c43 bl[43] br[43] wl[1] vdd gnd cell_6t
Xbit_r2_c43 bl[43] br[43] wl[2] vdd gnd cell_6t
Xbit_r3_c43 bl[43] br[43] wl[3] vdd gnd cell_6t
Xbit_r4_c43 bl[43] br[43] wl[4] vdd gnd cell_6t
Xbit_r5_c43 bl[43] br[43] wl[5] vdd gnd cell_6t
Xbit_r6_c43 bl[43] br[43] wl[6] vdd gnd cell_6t
Xbit_r7_c43 bl[43] br[43] wl[7] vdd gnd cell_6t
Xbit_r8_c43 bl[43] br[43] wl[8] vdd gnd cell_6t
Xbit_r9_c43 bl[43] br[43] wl[9] vdd gnd cell_6t
Xbit_r10_c43 bl[43] br[43] wl[10] vdd gnd cell_6t
Xbit_r11_c43 bl[43] br[43] wl[11] vdd gnd cell_6t
Xbit_r12_c43 bl[43] br[43] wl[12] vdd gnd cell_6t
Xbit_r13_c43 bl[43] br[43] wl[13] vdd gnd cell_6t
Xbit_r14_c43 bl[43] br[43] wl[14] vdd gnd cell_6t
Xbit_r15_c43 bl[43] br[43] wl[15] vdd gnd cell_6t
Xbit_r16_c43 bl[43] br[43] wl[16] vdd gnd cell_6t
Xbit_r17_c43 bl[43] br[43] wl[17] vdd gnd cell_6t
Xbit_r18_c43 bl[43] br[43] wl[18] vdd gnd cell_6t
Xbit_r19_c43 bl[43] br[43] wl[19] vdd gnd cell_6t
Xbit_r20_c43 bl[43] br[43] wl[20] vdd gnd cell_6t
Xbit_r21_c43 bl[43] br[43] wl[21] vdd gnd cell_6t
Xbit_r22_c43 bl[43] br[43] wl[22] vdd gnd cell_6t
Xbit_r23_c43 bl[43] br[43] wl[23] vdd gnd cell_6t
Xbit_r24_c43 bl[43] br[43] wl[24] vdd gnd cell_6t
Xbit_r25_c43 bl[43] br[43] wl[25] vdd gnd cell_6t
Xbit_r26_c43 bl[43] br[43] wl[26] vdd gnd cell_6t
Xbit_r27_c43 bl[43] br[43] wl[27] vdd gnd cell_6t
Xbit_r28_c43 bl[43] br[43] wl[28] vdd gnd cell_6t
Xbit_r29_c43 bl[43] br[43] wl[29] vdd gnd cell_6t
Xbit_r30_c43 bl[43] br[43] wl[30] vdd gnd cell_6t
Xbit_r31_c43 bl[43] br[43] wl[31] vdd gnd cell_6t
Xbit_r32_c43 bl[43] br[43] wl[32] vdd gnd cell_6t
Xbit_r33_c43 bl[43] br[43] wl[33] vdd gnd cell_6t
Xbit_r34_c43 bl[43] br[43] wl[34] vdd gnd cell_6t
Xbit_r35_c43 bl[43] br[43] wl[35] vdd gnd cell_6t
Xbit_r36_c43 bl[43] br[43] wl[36] vdd gnd cell_6t
Xbit_r37_c43 bl[43] br[43] wl[37] vdd gnd cell_6t
Xbit_r38_c43 bl[43] br[43] wl[38] vdd gnd cell_6t
Xbit_r39_c43 bl[43] br[43] wl[39] vdd gnd cell_6t
Xbit_r40_c43 bl[43] br[43] wl[40] vdd gnd cell_6t
Xbit_r41_c43 bl[43] br[43] wl[41] vdd gnd cell_6t
Xbit_r42_c43 bl[43] br[43] wl[42] vdd gnd cell_6t
Xbit_r43_c43 bl[43] br[43] wl[43] vdd gnd cell_6t
Xbit_r44_c43 bl[43] br[43] wl[44] vdd gnd cell_6t
Xbit_r45_c43 bl[43] br[43] wl[45] vdd gnd cell_6t
Xbit_r46_c43 bl[43] br[43] wl[46] vdd gnd cell_6t
Xbit_r47_c43 bl[43] br[43] wl[47] vdd gnd cell_6t
Xbit_r48_c43 bl[43] br[43] wl[48] vdd gnd cell_6t
Xbit_r49_c43 bl[43] br[43] wl[49] vdd gnd cell_6t
Xbit_r50_c43 bl[43] br[43] wl[50] vdd gnd cell_6t
Xbit_r51_c43 bl[43] br[43] wl[51] vdd gnd cell_6t
Xbit_r52_c43 bl[43] br[43] wl[52] vdd gnd cell_6t
Xbit_r53_c43 bl[43] br[43] wl[53] vdd gnd cell_6t
Xbit_r54_c43 bl[43] br[43] wl[54] vdd gnd cell_6t
Xbit_r55_c43 bl[43] br[43] wl[55] vdd gnd cell_6t
Xbit_r56_c43 bl[43] br[43] wl[56] vdd gnd cell_6t
Xbit_r57_c43 bl[43] br[43] wl[57] vdd gnd cell_6t
Xbit_r58_c43 bl[43] br[43] wl[58] vdd gnd cell_6t
Xbit_r59_c43 bl[43] br[43] wl[59] vdd gnd cell_6t
Xbit_r60_c43 bl[43] br[43] wl[60] vdd gnd cell_6t
Xbit_r61_c43 bl[43] br[43] wl[61] vdd gnd cell_6t
Xbit_r62_c43 bl[43] br[43] wl[62] vdd gnd cell_6t
Xbit_r63_c43 bl[43] br[43] wl[63] vdd gnd cell_6t
Xbit_r64_c43 bl[43] br[43] wl[64] vdd gnd cell_6t
Xbit_r65_c43 bl[43] br[43] wl[65] vdd gnd cell_6t
Xbit_r66_c43 bl[43] br[43] wl[66] vdd gnd cell_6t
Xbit_r67_c43 bl[43] br[43] wl[67] vdd gnd cell_6t
Xbit_r68_c43 bl[43] br[43] wl[68] vdd gnd cell_6t
Xbit_r69_c43 bl[43] br[43] wl[69] vdd gnd cell_6t
Xbit_r70_c43 bl[43] br[43] wl[70] vdd gnd cell_6t
Xbit_r71_c43 bl[43] br[43] wl[71] vdd gnd cell_6t
Xbit_r72_c43 bl[43] br[43] wl[72] vdd gnd cell_6t
Xbit_r73_c43 bl[43] br[43] wl[73] vdd gnd cell_6t
Xbit_r74_c43 bl[43] br[43] wl[74] vdd gnd cell_6t
Xbit_r75_c43 bl[43] br[43] wl[75] vdd gnd cell_6t
Xbit_r76_c43 bl[43] br[43] wl[76] vdd gnd cell_6t
Xbit_r77_c43 bl[43] br[43] wl[77] vdd gnd cell_6t
Xbit_r78_c43 bl[43] br[43] wl[78] vdd gnd cell_6t
Xbit_r79_c43 bl[43] br[43] wl[79] vdd gnd cell_6t
Xbit_r80_c43 bl[43] br[43] wl[80] vdd gnd cell_6t
Xbit_r81_c43 bl[43] br[43] wl[81] vdd gnd cell_6t
Xbit_r82_c43 bl[43] br[43] wl[82] vdd gnd cell_6t
Xbit_r83_c43 bl[43] br[43] wl[83] vdd gnd cell_6t
Xbit_r84_c43 bl[43] br[43] wl[84] vdd gnd cell_6t
Xbit_r85_c43 bl[43] br[43] wl[85] vdd gnd cell_6t
Xbit_r86_c43 bl[43] br[43] wl[86] vdd gnd cell_6t
Xbit_r87_c43 bl[43] br[43] wl[87] vdd gnd cell_6t
Xbit_r88_c43 bl[43] br[43] wl[88] vdd gnd cell_6t
Xbit_r89_c43 bl[43] br[43] wl[89] vdd gnd cell_6t
Xbit_r90_c43 bl[43] br[43] wl[90] vdd gnd cell_6t
Xbit_r91_c43 bl[43] br[43] wl[91] vdd gnd cell_6t
Xbit_r92_c43 bl[43] br[43] wl[92] vdd gnd cell_6t
Xbit_r93_c43 bl[43] br[43] wl[93] vdd gnd cell_6t
Xbit_r94_c43 bl[43] br[43] wl[94] vdd gnd cell_6t
Xbit_r95_c43 bl[43] br[43] wl[95] vdd gnd cell_6t
Xbit_r96_c43 bl[43] br[43] wl[96] vdd gnd cell_6t
Xbit_r97_c43 bl[43] br[43] wl[97] vdd gnd cell_6t
Xbit_r98_c43 bl[43] br[43] wl[98] vdd gnd cell_6t
Xbit_r99_c43 bl[43] br[43] wl[99] vdd gnd cell_6t
Xbit_r100_c43 bl[43] br[43] wl[100] vdd gnd cell_6t
Xbit_r101_c43 bl[43] br[43] wl[101] vdd gnd cell_6t
Xbit_r102_c43 bl[43] br[43] wl[102] vdd gnd cell_6t
Xbit_r103_c43 bl[43] br[43] wl[103] vdd gnd cell_6t
Xbit_r104_c43 bl[43] br[43] wl[104] vdd gnd cell_6t
Xbit_r105_c43 bl[43] br[43] wl[105] vdd gnd cell_6t
Xbit_r106_c43 bl[43] br[43] wl[106] vdd gnd cell_6t
Xbit_r107_c43 bl[43] br[43] wl[107] vdd gnd cell_6t
Xbit_r108_c43 bl[43] br[43] wl[108] vdd gnd cell_6t
Xbit_r109_c43 bl[43] br[43] wl[109] vdd gnd cell_6t
Xbit_r110_c43 bl[43] br[43] wl[110] vdd gnd cell_6t
Xbit_r111_c43 bl[43] br[43] wl[111] vdd gnd cell_6t
Xbit_r112_c43 bl[43] br[43] wl[112] vdd gnd cell_6t
Xbit_r113_c43 bl[43] br[43] wl[113] vdd gnd cell_6t
Xbit_r114_c43 bl[43] br[43] wl[114] vdd gnd cell_6t
Xbit_r115_c43 bl[43] br[43] wl[115] vdd gnd cell_6t
Xbit_r116_c43 bl[43] br[43] wl[116] vdd gnd cell_6t
Xbit_r117_c43 bl[43] br[43] wl[117] vdd gnd cell_6t
Xbit_r118_c43 bl[43] br[43] wl[118] vdd gnd cell_6t
Xbit_r119_c43 bl[43] br[43] wl[119] vdd gnd cell_6t
Xbit_r120_c43 bl[43] br[43] wl[120] vdd gnd cell_6t
Xbit_r121_c43 bl[43] br[43] wl[121] vdd gnd cell_6t
Xbit_r122_c43 bl[43] br[43] wl[122] vdd gnd cell_6t
Xbit_r123_c43 bl[43] br[43] wl[123] vdd gnd cell_6t
Xbit_r124_c43 bl[43] br[43] wl[124] vdd gnd cell_6t
Xbit_r125_c43 bl[43] br[43] wl[125] vdd gnd cell_6t
Xbit_r126_c43 bl[43] br[43] wl[126] vdd gnd cell_6t
Xbit_r127_c43 bl[43] br[43] wl[127] vdd gnd cell_6t
Xbit_r128_c43 bl[43] br[43] wl[128] vdd gnd cell_6t
Xbit_r129_c43 bl[43] br[43] wl[129] vdd gnd cell_6t
Xbit_r130_c43 bl[43] br[43] wl[130] vdd gnd cell_6t
Xbit_r131_c43 bl[43] br[43] wl[131] vdd gnd cell_6t
Xbit_r132_c43 bl[43] br[43] wl[132] vdd gnd cell_6t
Xbit_r133_c43 bl[43] br[43] wl[133] vdd gnd cell_6t
Xbit_r134_c43 bl[43] br[43] wl[134] vdd gnd cell_6t
Xbit_r135_c43 bl[43] br[43] wl[135] vdd gnd cell_6t
Xbit_r136_c43 bl[43] br[43] wl[136] vdd gnd cell_6t
Xbit_r137_c43 bl[43] br[43] wl[137] vdd gnd cell_6t
Xbit_r138_c43 bl[43] br[43] wl[138] vdd gnd cell_6t
Xbit_r139_c43 bl[43] br[43] wl[139] vdd gnd cell_6t
Xbit_r140_c43 bl[43] br[43] wl[140] vdd gnd cell_6t
Xbit_r141_c43 bl[43] br[43] wl[141] vdd gnd cell_6t
Xbit_r142_c43 bl[43] br[43] wl[142] vdd gnd cell_6t
Xbit_r143_c43 bl[43] br[43] wl[143] vdd gnd cell_6t
Xbit_r144_c43 bl[43] br[43] wl[144] vdd gnd cell_6t
Xbit_r145_c43 bl[43] br[43] wl[145] vdd gnd cell_6t
Xbit_r146_c43 bl[43] br[43] wl[146] vdd gnd cell_6t
Xbit_r147_c43 bl[43] br[43] wl[147] vdd gnd cell_6t
Xbit_r148_c43 bl[43] br[43] wl[148] vdd gnd cell_6t
Xbit_r149_c43 bl[43] br[43] wl[149] vdd gnd cell_6t
Xbit_r150_c43 bl[43] br[43] wl[150] vdd gnd cell_6t
Xbit_r151_c43 bl[43] br[43] wl[151] vdd gnd cell_6t
Xbit_r152_c43 bl[43] br[43] wl[152] vdd gnd cell_6t
Xbit_r153_c43 bl[43] br[43] wl[153] vdd gnd cell_6t
Xbit_r154_c43 bl[43] br[43] wl[154] vdd gnd cell_6t
Xbit_r155_c43 bl[43] br[43] wl[155] vdd gnd cell_6t
Xbit_r156_c43 bl[43] br[43] wl[156] vdd gnd cell_6t
Xbit_r157_c43 bl[43] br[43] wl[157] vdd gnd cell_6t
Xbit_r158_c43 bl[43] br[43] wl[158] vdd gnd cell_6t
Xbit_r159_c43 bl[43] br[43] wl[159] vdd gnd cell_6t
Xbit_r160_c43 bl[43] br[43] wl[160] vdd gnd cell_6t
Xbit_r161_c43 bl[43] br[43] wl[161] vdd gnd cell_6t
Xbit_r162_c43 bl[43] br[43] wl[162] vdd gnd cell_6t
Xbit_r163_c43 bl[43] br[43] wl[163] vdd gnd cell_6t
Xbit_r164_c43 bl[43] br[43] wl[164] vdd gnd cell_6t
Xbit_r165_c43 bl[43] br[43] wl[165] vdd gnd cell_6t
Xbit_r166_c43 bl[43] br[43] wl[166] vdd gnd cell_6t
Xbit_r167_c43 bl[43] br[43] wl[167] vdd gnd cell_6t
Xbit_r168_c43 bl[43] br[43] wl[168] vdd gnd cell_6t
Xbit_r169_c43 bl[43] br[43] wl[169] vdd gnd cell_6t
Xbit_r170_c43 bl[43] br[43] wl[170] vdd gnd cell_6t
Xbit_r171_c43 bl[43] br[43] wl[171] vdd gnd cell_6t
Xbit_r172_c43 bl[43] br[43] wl[172] vdd gnd cell_6t
Xbit_r173_c43 bl[43] br[43] wl[173] vdd gnd cell_6t
Xbit_r174_c43 bl[43] br[43] wl[174] vdd gnd cell_6t
Xbit_r175_c43 bl[43] br[43] wl[175] vdd gnd cell_6t
Xbit_r176_c43 bl[43] br[43] wl[176] vdd gnd cell_6t
Xbit_r177_c43 bl[43] br[43] wl[177] vdd gnd cell_6t
Xbit_r178_c43 bl[43] br[43] wl[178] vdd gnd cell_6t
Xbit_r179_c43 bl[43] br[43] wl[179] vdd gnd cell_6t
Xbit_r180_c43 bl[43] br[43] wl[180] vdd gnd cell_6t
Xbit_r181_c43 bl[43] br[43] wl[181] vdd gnd cell_6t
Xbit_r182_c43 bl[43] br[43] wl[182] vdd gnd cell_6t
Xbit_r183_c43 bl[43] br[43] wl[183] vdd gnd cell_6t
Xbit_r184_c43 bl[43] br[43] wl[184] vdd gnd cell_6t
Xbit_r185_c43 bl[43] br[43] wl[185] vdd gnd cell_6t
Xbit_r186_c43 bl[43] br[43] wl[186] vdd gnd cell_6t
Xbit_r187_c43 bl[43] br[43] wl[187] vdd gnd cell_6t
Xbit_r188_c43 bl[43] br[43] wl[188] vdd gnd cell_6t
Xbit_r189_c43 bl[43] br[43] wl[189] vdd gnd cell_6t
Xbit_r190_c43 bl[43] br[43] wl[190] vdd gnd cell_6t
Xbit_r191_c43 bl[43] br[43] wl[191] vdd gnd cell_6t
Xbit_r192_c43 bl[43] br[43] wl[192] vdd gnd cell_6t
Xbit_r193_c43 bl[43] br[43] wl[193] vdd gnd cell_6t
Xbit_r194_c43 bl[43] br[43] wl[194] vdd gnd cell_6t
Xbit_r195_c43 bl[43] br[43] wl[195] vdd gnd cell_6t
Xbit_r196_c43 bl[43] br[43] wl[196] vdd gnd cell_6t
Xbit_r197_c43 bl[43] br[43] wl[197] vdd gnd cell_6t
Xbit_r198_c43 bl[43] br[43] wl[198] vdd gnd cell_6t
Xbit_r199_c43 bl[43] br[43] wl[199] vdd gnd cell_6t
Xbit_r200_c43 bl[43] br[43] wl[200] vdd gnd cell_6t
Xbit_r201_c43 bl[43] br[43] wl[201] vdd gnd cell_6t
Xbit_r202_c43 bl[43] br[43] wl[202] vdd gnd cell_6t
Xbit_r203_c43 bl[43] br[43] wl[203] vdd gnd cell_6t
Xbit_r204_c43 bl[43] br[43] wl[204] vdd gnd cell_6t
Xbit_r205_c43 bl[43] br[43] wl[205] vdd gnd cell_6t
Xbit_r206_c43 bl[43] br[43] wl[206] vdd gnd cell_6t
Xbit_r207_c43 bl[43] br[43] wl[207] vdd gnd cell_6t
Xbit_r208_c43 bl[43] br[43] wl[208] vdd gnd cell_6t
Xbit_r209_c43 bl[43] br[43] wl[209] vdd gnd cell_6t
Xbit_r210_c43 bl[43] br[43] wl[210] vdd gnd cell_6t
Xbit_r211_c43 bl[43] br[43] wl[211] vdd gnd cell_6t
Xbit_r212_c43 bl[43] br[43] wl[212] vdd gnd cell_6t
Xbit_r213_c43 bl[43] br[43] wl[213] vdd gnd cell_6t
Xbit_r214_c43 bl[43] br[43] wl[214] vdd gnd cell_6t
Xbit_r215_c43 bl[43] br[43] wl[215] vdd gnd cell_6t
Xbit_r216_c43 bl[43] br[43] wl[216] vdd gnd cell_6t
Xbit_r217_c43 bl[43] br[43] wl[217] vdd gnd cell_6t
Xbit_r218_c43 bl[43] br[43] wl[218] vdd gnd cell_6t
Xbit_r219_c43 bl[43] br[43] wl[219] vdd gnd cell_6t
Xbit_r220_c43 bl[43] br[43] wl[220] vdd gnd cell_6t
Xbit_r221_c43 bl[43] br[43] wl[221] vdd gnd cell_6t
Xbit_r222_c43 bl[43] br[43] wl[222] vdd gnd cell_6t
Xbit_r223_c43 bl[43] br[43] wl[223] vdd gnd cell_6t
Xbit_r224_c43 bl[43] br[43] wl[224] vdd gnd cell_6t
Xbit_r225_c43 bl[43] br[43] wl[225] vdd gnd cell_6t
Xbit_r226_c43 bl[43] br[43] wl[226] vdd gnd cell_6t
Xbit_r227_c43 bl[43] br[43] wl[227] vdd gnd cell_6t
Xbit_r228_c43 bl[43] br[43] wl[228] vdd gnd cell_6t
Xbit_r229_c43 bl[43] br[43] wl[229] vdd gnd cell_6t
Xbit_r230_c43 bl[43] br[43] wl[230] vdd gnd cell_6t
Xbit_r231_c43 bl[43] br[43] wl[231] vdd gnd cell_6t
Xbit_r232_c43 bl[43] br[43] wl[232] vdd gnd cell_6t
Xbit_r233_c43 bl[43] br[43] wl[233] vdd gnd cell_6t
Xbit_r234_c43 bl[43] br[43] wl[234] vdd gnd cell_6t
Xbit_r235_c43 bl[43] br[43] wl[235] vdd gnd cell_6t
Xbit_r236_c43 bl[43] br[43] wl[236] vdd gnd cell_6t
Xbit_r237_c43 bl[43] br[43] wl[237] vdd gnd cell_6t
Xbit_r238_c43 bl[43] br[43] wl[238] vdd gnd cell_6t
Xbit_r239_c43 bl[43] br[43] wl[239] vdd gnd cell_6t
Xbit_r240_c43 bl[43] br[43] wl[240] vdd gnd cell_6t
Xbit_r241_c43 bl[43] br[43] wl[241] vdd gnd cell_6t
Xbit_r242_c43 bl[43] br[43] wl[242] vdd gnd cell_6t
Xbit_r243_c43 bl[43] br[43] wl[243] vdd gnd cell_6t
Xbit_r244_c43 bl[43] br[43] wl[244] vdd gnd cell_6t
Xbit_r245_c43 bl[43] br[43] wl[245] vdd gnd cell_6t
Xbit_r246_c43 bl[43] br[43] wl[246] vdd gnd cell_6t
Xbit_r247_c43 bl[43] br[43] wl[247] vdd gnd cell_6t
Xbit_r248_c43 bl[43] br[43] wl[248] vdd gnd cell_6t
Xbit_r249_c43 bl[43] br[43] wl[249] vdd gnd cell_6t
Xbit_r250_c43 bl[43] br[43] wl[250] vdd gnd cell_6t
Xbit_r251_c43 bl[43] br[43] wl[251] vdd gnd cell_6t
Xbit_r252_c43 bl[43] br[43] wl[252] vdd gnd cell_6t
Xbit_r253_c43 bl[43] br[43] wl[253] vdd gnd cell_6t
Xbit_r254_c43 bl[43] br[43] wl[254] vdd gnd cell_6t
Xbit_r255_c43 bl[43] br[43] wl[255] vdd gnd cell_6t
Xbit_r256_c43 bl[43] br[43] wl[256] vdd gnd cell_6t
Xbit_r257_c43 bl[43] br[43] wl[257] vdd gnd cell_6t
Xbit_r258_c43 bl[43] br[43] wl[258] vdd gnd cell_6t
Xbit_r259_c43 bl[43] br[43] wl[259] vdd gnd cell_6t
Xbit_r260_c43 bl[43] br[43] wl[260] vdd gnd cell_6t
Xbit_r261_c43 bl[43] br[43] wl[261] vdd gnd cell_6t
Xbit_r262_c43 bl[43] br[43] wl[262] vdd gnd cell_6t
Xbit_r263_c43 bl[43] br[43] wl[263] vdd gnd cell_6t
Xbit_r264_c43 bl[43] br[43] wl[264] vdd gnd cell_6t
Xbit_r265_c43 bl[43] br[43] wl[265] vdd gnd cell_6t
Xbit_r266_c43 bl[43] br[43] wl[266] vdd gnd cell_6t
Xbit_r267_c43 bl[43] br[43] wl[267] vdd gnd cell_6t
Xbit_r268_c43 bl[43] br[43] wl[268] vdd gnd cell_6t
Xbit_r269_c43 bl[43] br[43] wl[269] vdd gnd cell_6t
Xbit_r270_c43 bl[43] br[43] wl[270] vdd gnd cell_6t
Xbit_r271_c43 bl[43] br[43] wl[271] vdd gnd cell_6t
Xbit_r272_c43 bl[43] br[43] wl[272] vdd gnd cell_6t
Xbit_r273_c43 bl[43] br[43] wl[273] vdd gnd cell_6t
Xbit_r274_c43 bl[43] br[43] wl[274] vdd gnd cell_6t
Xbit_r275_c43 bl[43] br[43] wl[275] vdd gnd cell_6t
Xbit_r276_c43 bl[43] br[43] wl[276] vdd gnd cell_6t
Xbit_r277_c43 bl[43] br[43] wl[277] vdd gnd cell_6t
Xbit_r278_c43 bl[43] br[43] wl[278] vdd gnd cell_6t
Xbit_r279_c43 bl[43] br[43] wl[279] vdd gnd cell_6t
Xbit_r280_c43 bl[43] br[43] wl[280] vdd gnd cell_6t
Xbit_r281_c43 bl[43] br[43] wl[281] vdd gnd cell_6t
Xbit_r282_c43 bl[43] br[43] wl[282] vdd gnd cell_6t
Xbit_r283_c43 bl[43] br[43] wl[283] vdd gnd cell_6t
Xbit_r284_c43 bl[43] br[43] wl[284] vdd gnd cell_6t
Xbit_r285_c43 bl[43] br[43] wl[285] vdd gnd cell_6t
Xbit_r286_c43 bl[43] br[43] wl[286] vdd gnd cell_6t
Xbit_r287_c43 bl[43] br[43] wl[287] vdd gnd cell_6t
Xbit_r288_c43 bl[43] br[43] wl[288] vdd gnd cell_6t
Xbit_r289_c43 bl[43] br[43] wl[289] vdd gnd cell_6t
Xbit_r290_c43 bl[43] br[43] wl[290] vdd gnd cell_6t
Xbit_r291_c43 bl[43] br[43] wl[291] vdd gnd cell_6t
Xbit_r292_c43 bl[43] br[43] wl[292] vdd gnd cell_6t
Xbit_r293_c43 bl[43] br[43] wl[293] vdd gnd cell_6t
Xbit_r294_c43 bl[43] br[43] wl[294] vdd gnd cell_6t
Xbit_r295_c43 bl[43] br[43] wl[295] vdd gnd cell_6t
Xbit_r296_c43 bl[43] br[43] wl[296] vdd gnd cell_6t
Xbit_r297_c43 bl[43] br[43] wl[297] vdd gnd cell_6t
Xbit_r298_c43 bl[43] br[43] wl[298] vdd gnd cell_6t
Xbit_r299_c43 bl[43] br[43] wl[299] vdd gnd cell_6t
Xbit_r300_c43 bl[43] br[43] wl[300] vdd gnd cell_6t
Xbit_r301_c43 bl[43] br[43] wl[301] vdd gnd cell_6t
Xbit_r302_c43 bl[43] br[43] wl[302] vdd gnd cell_6t
Xbit_r303_c43 bl[43] br[43] wl[303] vdd gnd cell_6t
Xbit_r304_c43 bl[43] br[43] wl[304] vdd gnd cell_6t
Xbit_r305_c43 bl[43] br[43] wl[305] vdd gnd cell_6t
Xbit_r306_c43 bl[43] br[43] wl[306] vdd gnd cell_6t
Xbit_r307_c43 bl[43] br[43] wl[307] vdd gnd cell_6t
Xbit_r308_c43 bl[43] br[43] wl[308] vdd gnd cell_6t
Xbit_r309_c43 bl[43] br[43] wl[309] vdd gnd cell_6t
Xbit_r310_c43 bl[43] br[43] wl[310] vdd gnd cell_6t
Xbit_r311_c43 bl[43] br[43] wl[311] vdd gnd cell_6t
Xbit_r312_c43 bl[43] br[43] wl[312] vdd gnd cell_6t
Xbit_r313_c43 bl[43] br[43] wl[313] vdd gnd cell_6t
Xbit_r314_c43 bl[43] br[43] wl[314] vdd gnd cell_6t
Xbit_r315_c43 bl[43] br[43] wl[315] vdd gnd cell_6t
Xbit_r316_c43 bl[43] br[43] wl[316] vdd gnd cell_6t
Xbit_r317_c43 bl[43] br[43] wl[317] vdd gnd cell_6t
Xbit_r318_c43 bl[43] br[43] wl[318] vdd gnd cell_6t
Xbit_r319_c43 bl[43] br[43] wl[319] vdd gnd cell_6t
Xbit_r320_c43 bl[43] br[43] wl[320] vdd gnd cell_6t
Xbit_r321_c43 bl[43] br[43] wl[321] vdd gnd cell_6t
Xbit_r322_c43 bl[43] br[43] wl[322] vdd gnd cell_6t
Xbit_r323_c43 bl[43] br[43] wl[323] vdd gnd cell_6t
Xbit_r324_c43 bl[43] br[43] wl[324] vdd gnd cell_6t
Xbit_r325_c43 bl[43] br[43] wl[325] vdd gnd cell_6t
Xbit_r326_c43 bl[43] br[43] wl[326] vdd gnd cell_6t
Xbit_r327_c43 bl[43] br[43] wl[327] vdd gnd cell_6t
Xbit_r328_c43 bl[43] br[43] wl[328] vdd gnd cell_6t
Xbit_r329_c43 bl[43] br[43] wl[329] vdd gnd cell_6t
Xbit_r330_c43 bl[43] br[43] wl[330] vdd gnd cell_6t
Xbit_r331_c43 bl[43] br[43] wl[331] vdd gnd cell_6t
Xbit_r332_c43 bl[43] br[43] wl[332] vdd gnd cell_6t
Xbit_r333_c43 bl[43] br[43] wl[333] vdd gnd cell_6t
Xbit_r334_c43 bl[43] br[43] wl[334] vdd gnd cell_6t
Xbit_r335_c43 bl[43] br[43] wl[335] vdd gnd cell_6t
Xbit_r336_c43 bl[43] br[43] wl[336] vdd gnd cell_6t
Xbit_r337_c43 bl[43] br[43] wl[337] vdd gnd cell_6t
Xbit_r338_c43 bl[43] br[43] wl[338] vdd gnd cell_6t
Xbit_r339_c43 bl[43] br[43] wl[339] vdd gnd cell_6t
Xbit_r340_c43 bl[43] br[43] wl[340] vdd gnd cell_6t
Xbit_r341_c43 bl[43] br[43] wl[341] vdd gnd cell_6t
Xbit_r342_c43 bl[43] br[43] wl[342] vdd gnd cell_6t
Xbit_r343_c43 bl[43] br[43] wl[343] vdd gnd cell_6t
Xbit_r344_c43 bl[43] br[43] wl[344] vdd gnd cell_6t
Xbit_r345_c43 bl[43] br[43] wl[345] vdd gnd cell_6t
Xbit_r346_c43 bl[43] br[43] wl[346] vdd gnd cell_6t
Xbit_r347_c43 bl[43] br[43] wl[347] vdd gnd cell_6t
Xbit_r348_c43 bl[43] br[43] wl[348] vdd gnd cell_6t
Xbit_r349_c43 bl[43] br[43] wl[349] vdd gnd cell_6t
Xbit_r350_c43 bl[43] br[43] wl[350] vdd gnd cell_6t
Xbit_r351_c43 bl[43] br[43] wl[351] vdd gnd cell_6t
Xbit_r352_c43 bl[43] br[43] wl[352] vdd gnd cell_6t
Xbit_r353_c43 bl[43] br[43] wl[353] vdd gnd cell_6t
Xbit_r354_c43 bl[43] br[43] wl[354] vdd gnd cell_6t
Xbit_r355_c43 bl[43] br[43] wl[355] vdd gnd cell_6t
Xbit_r356_c43 bl[43] br[43] wl[356] vdd gnd cell_6t
Xbit_r357_c43 bl[43] br[43] wl[357] vdd gnd cell_6t
Xbit_r358_c43 bl[43] br[43] wl[358] vdd gnd cell_6t
Xbit_r359_c43 bl[43] br[43] wl[359] vdd gnd cell_6t
Xbit_r360_c43 bl[43] br[43] wl[360] vdd gnd cell_6t
Xbit_r361_c43 bl[43] br[43] wl[361] vdd gnd cell_6t
Xbit_r362_c43 bl[43] br[43] wl[362] vdd gnd cell_6t
Xbit_r363_c43 bl[43] br[43] wl[363] vdd gnd cell_6t
Xbit_r364_c43 bl[43] br[43] wl[364] vdd gnd cell_6t
Xbit_r365_c43 bl[43] br[43] wl[365] vdd gnd cell_6t
Xbit_r366_c43 bl[43] br[43] wl[366] vdd gnd cell_6t
Xbit_r367_c43 bl[43] br[43] wl[367] vdd gnd cell_6t
Xbit_r368_c43 bl[43] br[43] wl[368] vdd gnd cell_6t
Xbit_r369_c43 bl[43] br[43] wl[369] vdd gnd cell_6t
Xbit_r370_c43 bl[43] br[43] wl[370] vdd gnd cell_6t
Xbit_r371_c43 bl[43] br[43] wl[371] vdd gnd cell_6t
Xbit_r372_c43 bl[43] br[43] wl[372] vdd gnd cell_6t
Xbit_r373_c43 bl[43] br[43] wl[373] vdd gnd cell_6t
Xbit_r374_c43 bl[43] br[43] wl[374] vdd gnd cell_6t
Xbit_r375_c43 bl[43] br[43] wl[375] vdd gnd cell_6t
Xbit_r376_c43 bl[43] br[43] wl[376] vdd gnd cell_6t
Xbit_r377_c43 bl[43] br[43] wl[377] vdd gnd cell_6t
Xbit_r378_c43 bl[43] br[43] wl[378] vdd gnd cell_6t
Xbit_r379_c43 bl[43] br[43] wl[379] vdd gnd cell_6t
Xbit_r380_c43 bl[43] br[43] wl[380] vdd gnd cell_6t
Xbit_r381_c43 bl[43] br[43] wl[381] vdd gnd cell_6t
Xbit_r382_c43 bl[43] br[43] wl[382] vdd gnd cell_6t
Xbit_r383_c43 bl[43] br[43] wl[383] vdd gnd cell_6t
Xbit_r384_c43 bl[43] br[43] wl[384] vdd gnd cell_6t
Xbit_r385_c43 bl[43] br[43] wl[385] vdd gnd cell_6t
Xbit_r386_c43 bl[43] br[43] wl[386] vdd gnd cell_6t
Xbit_r387_c43 bl[43] br[43] wl[387] vdd gnd cell_6t
Xbit_r388_c43 bl[43] br[43] wl[388] vdd gnd cell_6t
Xbit_r389_c43 bl[43] br[43] wl[389] vdd gnd cell_6t
Xbit_r390_c43 bl[43] br[43] wl[390] vdd gnd cell_6t
Xbit_r391_c43 bl[43] br[43] wl[391] vdd gnd cell_6t
Xbit_r392_c43 bl[43] br[43] wl[392] vdd gnd cell_6t
Xbit_r393_c43 bl[43] br[43] wl[393] vdd gnd cell_6t
Xbit_r394_c43 bl[43] br[43] wl[394] vdd gnd cell_6t
Xbit_r395_c43 bl[43] br[43] wl[395] vdd gnd cell_6t
Xbit_r396_c43 bl[43] br[43] wl[396] vdd gnd cell_6t
Xbit_r397_c43 bl[43] br[43] wl[397] vdd gnd cell_6t
Xbit_r398_c43 bl[43] br[43] wl[398] vdd gnd cell_6t
Xbit_r399_c43 bl[43] br[43] wl[399] vdd gnd cell_6t
Xbit_r400_c43 bl[43] br[43] wl[400] vdd gnd cell_6t
Xbit_r401_c43 bl[43] br[43] wl[401] vdd gnd cell_6t
Xbit_r402_c43 bl[43] br[43] wl[402] vdd gnd cell_6t
Xbit_r403_c43 bl[43] br[43] wl[403] vdd gnd cell_6t
Xbit_r404_c43 bl[43] br[43] wl[404] vdd gnd cell_6t
Xbit_r405_c43 bl[43] br[43] wl[405] vdd gnd cell_6t
Xbit_r406_c43 bl[43] br[43] wl[406] vdd gnd cell_6t
Xbit_r407_c43 bl[43] br[43] wl[407] vdd gnd cell_6t
Xbit_r408_c43 bl[43] br[43] wl[408] vdd gnd cell_6t
Xbit_r409_c43 bl[43] br[43] wl[409] vdd gnd cell_6t
Xbit_r410_c43 bl[43] br[43] wl[410] vdd gnd cell_6t
Xbit_r411_c43 bl[43] br[43] wl[411] vdd gnd cell_6t
Xbit_r412_c43 bl[43] br[43] wl[412] vdd gnd cell_6t
Xbit_r413_c43 bl[43] br[43] wl[413] vdd gnd cell_6t
Xbit_r414_c43 bl[43] br[43] wl[414] vdd gnd cell_6t
Xbit_r415_c43 bl[43] br[43] wl[415] vdd gnd cell_6t
Xbit_r416_c43 bl[43] br[43] wl[416] vdd gnd cell_6t
Xbit_r417_c43 bl[43] br[43] wl[417] vdd gnd cell_6t
Xbit_r418_c43 bl[43] br[43] wl[418] vdd gnd cell_6t
Xbit_r419_c43 bl[43] br[43] wl[419] vdd gnd cell_6t
Xbit_r420_c43 bl[43] br[43] wl[420] vdd gnd cell_6t
Xbit_r421_c43 bl[43] br[43] wl[421] vdd gnd cell_6t
Xbit_r422_c43 bl[43] br[43] wl[422] vdd gnd cell_6t
Xbit_r423_c43 bl[43] br[43] wl[423] vdd gnd cell_6t
Xbit_r424_c43 bl[43] br[43] wl[424] vdd gnd cell_6t
Xbit_r425_c43 bl[43] br[43] wl[425] vdd gnd cell_6t
Xbit_r426_c43 bl[43] br[43] wl[426] vdd gnd cell_6t
Xbit_r427_c43 bl[43] br[43] wl[427] vdd gnd cell_6t
Xbit_r428_c43 bl[43] br[43] wl[428] vdd gnd cell_6t
Xbit_r429_c43 bl[43] br[43] wl[429] vdd gnd cell_6t
Xbit_r430_c43 bl[43] br[43] wl[430] vdd gnd cell_6t
Xbit_r431_c43 bl[43] br[43] wl[431] vdd gnd cell_6t
Xbit_r432_c43 bl[43] br[43] wl[432] vdd gnd cell_6t
Xbit_r433_c43 bl[43] br[43] wl[433] vdd gnd cell_6t
Xbit_r434_c43 bl[43] br[43] wl[434] vdd gnd cell_6t
Xbit_r435_c43 bl[43] br[43] wl[435] vdd gnd cell_6t
Xbit_r436_c43 bl[43] br[43] wl[436] vdd gnd cell_6t
Xbit_r437_c43 bl[43] br[43] wl[437] vdd gnd cell_6t
Xbit_r438_c43 bl[43] br[43] wl[438] vdd gnd cell_6t
Xbit_r439_c43 bl[43] br[43] wl[439] vdd gnd cell_6t
Xbit_r440_c43 bl[43] br[43] wl[440] vdd gnd cell_6t
Xbit_r441_c43 bl[43] br[43] wl[441] vdd gnd cell_6t
Xbit_r442_c43 bl[43] br[43] wl[442] vdd gnd cell_6t
Xbit_r443_c43 bl[43] br[43] wl[443] vdd gnd cell_6t
Xbit_r444_c43 bl[43] br[43] wl[444] vdd gnd cell_6t
Xbit_r445_c43 bl[43] br[43] wl[445] vdd gnd cell_6t
Xbit_r446_c43 bl[43] br[43] wl[446] vdd gnd cell_6t
Xbit_r447_c43 bl[43] br[43] wl[447] vdd gnd cell_6t
Xbit_r448_c43 bl[43] br[43] wl[448] vdd gnd cell_6t
Xbit_r449_c43 bl[43] br[43] wl[449] vdd gnd cell_6t
Xbit_r450_c43 bl[43] br[43] wl[450] vdd gnd cell_6t
Xbit_r451_c43 bl[43] br[43] wl[451] vdd gnd cell_6t
Xbit_r452_c43 bl[43] br[43] wl[452] vdd gnd cell_6t
Xbit_r453_c43 bl[43] br[43] wl[453] vdd gnd cell_6t
Xbit_r454_c43 bl[43] br[43] wl[454] vdd gnd cell_6t
Xbit_r455_c43 bl[43] br[43] wl[455] vdd gnd cell_6t
Xbit_r456_c43 bl[43] br[43] wl[456] vdd gnd cell_6t
Xbit_r457_c43 bl[43] br[43] wl[457] vdd gnd cell_6t
Xbit_r458_c43 bl[43] br[43] wl[458] vdd gnd cell_6t
Xbit_r459_c43 bl[43] br[43] wl[459] vdd gnd cell_6t
Xbit_r460_c43 bl[43] br[43] wl[460] vdd gnd cell_6t
Xbit_r461_c43 bl[43] br[43] wl[461] vdd gnd cell_6t
Xbit_r462_c43 bl[43] br[43] wl[462] vdd gnd cell_6t
Xbit_r463_c43 bl[43] br[43] wl[463] vdd gnd cell_6t
Xbit_r464_c43 bl[43] br[43] wl[464] vdd gnd cell_6t
Xbit_r465_c43 bl[43] br[43] wl[465] vdd gnd cell_6t
Xbit_r466_c43 bl[43] br[43] wl[466] vdd gnd cell_6t
Xbit_r467_c43 bl[43] br[43] wl[467] vdd gnd cell_6t
Xbit_r468_c43 bl[43] br[43] wl[468] vdd gnd cell_6t
Xbit_r469_c43 bl[43] br[43] wl[469] vdd gnd cell_6t
Xbit_r470_c43 bl[43] br[43] wl[470] vdd gnd cell_6t
Xbit_r471_c43 bl[43] br[43] wl[471] vdd gnd cell_6t
Xbit_r472_c43 bl[43] br[43] wl[472] vdd gnd cell_6t
Xbit_r473_c43 bl[43] br[43] wl[473] vdd gnd cell_6t
Xbit_r474_c43 bl[43] br[43] wl[474] vdd gnd cell_6t
Xbit_r475_c43 bl[43] br[43] wl[475] vdd gnd cell_6t
Xbit_r476_c43 bl[43] br[43] wl[476] vdd gnd cell_6t
Xbit_r477_c43 bl[43] br[43] wl[477] vdd gnd cell_6t
Xbit_r478_c43 bl[43] br[43] wl[478] vdd gnd cell_6t
Xbit_r479_c43 bl[43] br[43] wl[479] vdd gnd cell_6t
Xbit_r480_c43 bl[43] br[43] wl[480] vdd gnd cell_6t
Xbit_r481_c43 bl[43] br[43] wl[481] vdd gnd cell_6t
Xbit_r482_c43 bl[43] br[43] wl[482] vdd gnd cell_6t
Xbit_r483_c43 bl[43] br[43] wl[483] vdd gnd cell_6t
Xbit_r484_c43 bl[43] br[43] wl[484] vdd gnd cell_6t
Xbit_r485_c43 bl[43] br[43] wl[485] vdd gnd cell_6t
Xbit_r486_c43 bl[43] br[43] wl[486] vdd gnd cell_6t
Xbit_r487_c43 bl[43] br[43] wl[487] vdd gnd cell_6t
Xbit_r488_c43 bl[43] br[43] wl[488] vdd gnd cell_6t
Xbit_r489_c43 bl[43] br[43] wl[489] vdd gnd cell_6t
Xbit_r490_c43 bl[43] br[43] wl[490] vdd gnd cell_6t
Xbit_r491_c43 bl[43] br[43] wl[491] vdd gnd cell_6t
Xbit_r492_c43 bl[43] br[43] wl[492] vdd gnd cell_6t
Xbit_r493_c43 bl[43] br[43] wl[493] vdd gnd cell_6t
Xbit_r494_c43 bl[43] br[43] wl[494] vdd gnd cell_6t
Xbit_r495_c43 bl[43] br[43] wl[495] vdd gnd cell_6t
Xbit_r496_c43 bl[43] br[43] wl[496] vdd gnd cell_6t
Xbit_r497_c43 bl[43] br[43] wl[497] vdd gnd cell_6t
Xbit_r498_c43 bl[43] br[43] wl[498] vdd gnd cell_6t
Xbit_r499_c43 bl[43] br[43] wl[499] vdd gnd cell_6t
Xbit_r500_c43 bl[43] br[43] wl[500] vdd gnd cell_6t
Xbit_r501_c43 bl[43] br[43] wl[501] vdd gnd cell_6t
Xbit_r502_c43 bl[43] br[43] wl[502] vdd gnd cell_6t
Xbit_r503_c43 bl[43] br[43] wl[503] vdd gnd cell_6t
Xbit_r504_c43 bl[43] br[43] wl[504] vdd gnd cell_6t
Xbit_r505_c43 bl[43] br[43] wl[505] vdd gnd cell_6t
Xbit_r506_c43 bl[43] br[43] wl[506] vdd gnd cell_6t
Xbit_r507_c43 bl[43] br[43] wl[507] vdd gnd cell_6t
Xbit_r508_c43 bl[43] br[43] wl[508] vdd gnd cell_6t
Xbit_r509_c43 bl[43] br[43] wl[509] vdd gnd cell_6t
Xbit_r510_c43 bl[43] br[43] wl[510] vdd gnd cell_6t
Xbit_r511_c43 bl[43] br[43] wl[511] vdd gnd cell_6t
Xbit_r0_c44 bl[44] br[44] wl[0] vdd gnd cell_6t
Xbit_r1_c44 bl[44] br[44] wl[1] vdd gnd cell_6t
Xbit_r2_c44 bl[44] br[44] wl[2] vdd gnd cell_6t
Xbit_r3_c44 bl[44] br[44] wl[3] vdd gnd cell_6t
Xbit_r4_c44 bl[44] br[44] wl[4] vdd gnd cell_6t
Xbit_r5_c44 bl[44] br[44] wl[5] vdd gnd cell_6t
Xbit_r6_c44 bl[44] br[44] wl[6] vdd gnd cell_6t
Xbit_r7_c44 bl[44] br[44] wl[7] vdd gnd cell_6t
Xbit_r8_c44 bl[44] br[44] wl[8] vdd gnd cell_6t
Xbit_r9_c44 bl[44] br[44] wl[9] vdd gnd cell_6t
Xbit_r10_c44 bl[44] br[44] wl[10] vdd gnd cell_6t
Xbit_r11_c44 bl[44] br[44] wl[11] vdd gnd cell_6t
Xbit_r12_c44 bl[44] br[44] wl[12] vdd gnd cell_6t
Xbit_r13_c44 bl[44] br[44] wl[13] vdd gnd cell_6t
Xbit_r14_c44 bl[44] br[44] wl[14] vdd gnd cell_6t
Xbit_r15_c44 bl[44] br[44] wl[15] vdd gnd cell_6t
Xbit_r16_c44 bl[44] br[44] wl[16] vdd gnd cell_6t
Xbit_r17_c44 bl[44] br[44] wl[17] vdd gnd cell_6t
Xbit_r18_c44 bl[44] br[44] wl[18] vdd gnd cell_6t
Xbit_r19_c44 bl[44] br[44] wl[19] vdd gnd cell_6t
Xbit_r20_c44 bl[44] br[44] wl[20] vdd gnd cell_6t
Xbit_r21_c44 bl[44] br[44] wl[21] vdd gnd cell_6t
Xbit_r22_c44 bl[44] br[44] wl[22] vdd gnd cell_6t
Xbit_r23_c44 bl[44] br[44] wl[23] vdd gnd cell_6t
Xbit_r24_c44 bl[44] br[44] wl[24] vdd gnd cell_6t
Xbit_r25_c44 bl[44] br[44] wl[25] vdd gnd cell_6t
Xbit_r26_c44 bl[44] br[44] wl[26] vdd gnd cell_6t
Xbit_r27_c44 bl[44] br[44] wl[27] vdd gnd cell_6t
Xbit_r28_c44 bl[44] br[44] wl[28] vdd gnd cell_6t
Xbit_r29_c44 bl[44] br[44] wl[29] vdd gnd cell_6t
Xbit_r30_c44 bl[44] br[44] wl[30] vdd gnd cell_6t
Xbit_r31_c44 bl[44] br[44] wl[31] vdd gnd cell_6t
Xbit_r32_c44 bl[44] br[44] wl[32] vdd gnd cell_6t
Xbit_r33_c44 bl[44] br[44] wl[33] vdd gnd cell_6t
Xbit_r34_c44 bl[44] br[44] wl[34] vdd gnd cell_6t
Xbit_r35_c44 bl[44] br[44] wl[35] vdd gnd cell_6t
Xbit_r36_c44 bl[44] br[44] wl[36] vdd gnd cell_6t
Xbit_r37_c44 bl[44] br[44] wl[37] vdd gnd cell_6t
Xbit_r38_c44 bl[44] br[44] wl[38] vdd gnd cell_6t
Xbit_r39_c44 bl[44] br[44] wl[39] vdd gnd cell_6t
Xbit_r40_c44 bl[44] br[44] wl[40] vdd gnd cell_6t
Xbit_r41_c44 bl[44] br[44] wl[41] vdd gnd cell_6t
Xbit_r42_c44 bl[44] br[44] wl[42] vdd gnd cell_6t
Xbit_r43_c44 bl[44] br[44] wl[43] vdd gnd cell_6t
Xbit_r44_c44 bl[44] br[44] wl[44] vdd gnd cell_6t
Xbit_r45_c44 bl[44] br[44] wl[45] vdd gnd cell_6t
Xbit_r46_c44 bl[44] br[44] wl[46] vdd gnd cell_6t
Xbit_r47_c44 bl[44] br[44] wl[47] vdd gnd cell_6t
Xbit_r48_c44 bl[44] br[44] wl[48] vdd gnd cell_6t
Xbit_r49_c44 bl[44] br[44] wl[49] vdd gnd cell_6t
Xbit_r50_c44 bl[44] br[44] wl[50] vdd gnd cell_6t
Xbit_r51_c44 bl[44] br[44] wl[51] vdd gnd cell_6t
Xbit_r52_c44 bl[44] br[44] wl[52] vdd gnd cell_6t
Xbit_r53_c44 bl[44] br[44] wl[53] vdd gnd cell_6t
Xbit_r54_c44 bl[44] br[44] wl[54] vdd gnd cell_6t
Xbit_r55_c44 bl[44] br[44] wl[55] vdd gnd cell_6t
Xbit_r56_c44 bl[44] br[44] wl[56] vdd gnd cell_6t
Xbit_r57_c44 bl[44] br[44] wl[57] vdd gnd cell_6t
Xbit_r58_c44 bl[44] br[44] wl[58] vdd gnd cell_6t
Xbit_r59_c44 bl[44] br[44] wl[59] vdd gnd cell_6t
Xbit_r60_c44 bl[44] br[44] wl[60] vdd gnd cell_6t
Xbit_r61_c44 bl[44] br[44] wl[61] vdd gnd cell_6t
Xbit_r62_c44 bl[44] br[44] wl[62] vdd gnd cell_6t
Xbit_r63_c44 bl[44] br[44] wl[63] vdd gnd cell_6t
Xbit_r64_c44 bl[44] br[44] wl[64] vdd gnd cell_6t
Xbit_r65_c44 bl[44] br[44] wl[65] vdd gnd cell_6t
Xbit_r66_c44 bl[44] br[44] wl[66] vdd gnd cell_6t
Xbit_r67_c44 bl[44] br[44] wl[67] vdd gnd cell_6t
Xbit_r68_c44 bl[44] br[44] wl[68] vdd gnd cell_6t
Xbit_r69_c44 bl[44] br[44] wl[69] vdd gnd cell_6t
Xbit_r70_c44 bl[44] br[44] wl[70] vdd gnd cell_6t
Xbit_r71_c44 bl[44] br[44] wl[71] vdd gnd cell_6t
Xbit_r72_c44 bl[44] br[44] wl[72] vdd gnd cell_6t
Xbit_r73_c44 bl[44] br[44] wl[73] vdd gnd cell_6t
Xbit_r74_c44 bl[44] br[44] wl[74] vdd gnd cell_6t
Xbit_r75_c44 bl[44] br[44] wl[75] vdd gnd cell_6t
Xbit_r76_c44 bl[44] br[44] wl[76] vdd gnd cell_6t
Xbit_r77_c44 bl[44] br[44] wl[77] vdd gnd cell_6t
Xbit_r78_c44 bl[44] br[44] wl[78] vdd gnd cell_6t
Xbit_r79_c44 bl[44] br[44] wl[79] vdd gnd cell_6t
Xbit_r80_c44 bl[44] br[44] wl[80] vdd gnd cell_6t
Xbit_r81_c44 bl[44] br[44] wl[81] vdd gnd cell_6t
Xbit_r82_c44 bl[44] br[44] wl[82] vdd gnd cell_6t
Xbit_r83_c44 bl[44] br[44] wl[83] vdd gnd cell_6t
Xbit_r84_c44 bl[44] br[44] wl[84] vdd gnd cell_6t
Xbit_r85_c44 bl[44] br[44] wl[85] vdd gnd cell_6t
Xbit_r86_c44 bl[44] br[44] wl[86] vdd gnd cell_6t
Xbit_r87_c44 bl[44] br[44] wl[87] vdd gnd cell_6t
Xbit_r88_c44 bl[44] br[44] wl[88] vdd gnd cell_6t
Xbit_r89_c44 bl[44] br[44] wl[89] vdd gnd cell_6t
Xbit_r90_c44 bl[44] br[44] wl[90] vdd gnd cell_6t
Xbit_r91_c44 bl[44] br[44] wl[91] vdd gnd cell_6t
Xbit_r92_c44 bl[44] br[44] wl[92] vdd gnd cell_6t
Xbit_r93_c44 bl[44] br[44] wl[93] vdd gnd cell_6t
Xbit_r94_c44 bl[44] br[44] wl[94] vdd gnd cell_6t
Xbit_r95_c44 bl[44] br[44] wl[95] vdd gnd cell_6t
Xbit_r96_c44 bl[44] br[44] wl[96] vdd gnd cell_6t
Xbit_r97_c44 bl[44] br[44] wl[97] vdd gnd cell_6t
Xbit_r98_c44 bl[44] br[44] wl[98] vdd gnd cell_6t
Xbit_r99_c44 bl[44] br[44] wl[99] vdd gnd cell_6t
Xbit_r100_c44 bl[44] br[44] wl[100] vdd gnd cell_6t
Xbit_r101_c44 bl[44] br[44] wl[101] vdd gnd cell_6t
Xbit_r102_c44 bl[44] br[44] wl[102] vdd gnd cell_6t
Xbit_r103_c44 bl[44] br[44] wl[103] vdd gnd cell_6t
Xbit_r104_c44 bl[44] br[44] wl[104] vdd gnd cell_6t
Xbit_r105_c44 bl[44] br[44] wl[105] vdd gnd cell_6t
Xbit_r106_c44 bl[44] br[44] wl[106] vdd gnd cell_6t
Xbit_r107_c44 bl[44] br[44] wl[107] vdd gnd cell_6t
Xbit_r108_c44 bl[44] br[44] wl[108] vdd gnd cell_6t
Xbit_r109_c44 bl[44] br[44] wl[109] vdd gnd cell_6t
Xbit_r110_c44 bl[44] br[44] wl[110] vdd gnd cell_6t
Xbit_r111_c44 bl[44] br[44] wl[111] vdd gnd cell_6t
Xbit_r112_c44 bl[44] br[44] wl[112] vdd gnd cell_6t
Xbit_r113_c44 bl[44] br[44] wl[113] vdd gnd cell_6t
Xbit_r114_c44 bl[44] br[44] wl[114] vdd gnd cell_6t
Xbit_r115_c44 bl[44] br[44] wl[115] vdd gnd cell_6t
Xbit_r116_c44 bl[44] br[44] wl[116] vdd gnd cell_6t
Xbit_r117_c44 bl[44] br[44] wl[117] vdd gnd cell_6t
Xbit_r118_c44 bl[44] br[44] wl[118] vdd gnd cell_6t
Xbit_r119_c44 bl[44] br[44] wl[119] vdd gnd cell_6t
Xbit_r120_c44 bl[44] br[44] wl[120] vdd gnd cell_6t
Xbit_r121_c44 bl[44] br[44] wl[121] vdd gnd cell_6t
Xbit_r122_c44 bl[44] br[44] wl[122] vdd gnd cell_6t
Xbit_r123_c44 bl[44] br[44] wl[123] vdd gnd cell_6t
Xbit_r124_c44 bl[44] br[44] wl[124] vdd gnd cell_6t
Xbit_r125_c44 bl[44] br[44] wl[125] vdd gnd cell_6t
Xbit_r126_c44 bl[44] br[44] wl[126] vdd gnd cell_6t
Xbit_r127_c44 bl[44] br[44] wl[127] vdd gnd cell_6t
Xbit_r128_c44 bl[44] br[44] wl[128] vdd gnd cell_6t
Xbit_r129_c44 bl[44] br[44] wl[129] vdd gnd cell_6t
Xbit_r130_c44 bl[44] br[44] wl[130] vdd gnd cell_6t
Xbit_r131_c44 bl[44] br[44] wl[131] vdd gnd cell_6t
Xbit_r132_c44 bl[44] br[44] wl[132] vdd gnd cell_6t
Xbit_r133_c44 bl[44] br[44] wl[133] vdd gnd cell_6t
Xbit_r134_c44 bl[44] br[44] wl[134] vdd gnd cell_6t
Xbit_r135_c44 bl[44] br[44] wl[135] vdd gnd cell_6t
Xbit_r136_c44 bl[44] br[44] wl[136] vdd gnd cell_6t
Xbit_r137_c44 bl[44] br[44] wl[137] vdd gnd cell_6t
Xbit_r138_c44 bl[44] br[44] wl[138] vdd gnd cell_6t
Xbit_r139_c44 bl[44] br[44] wl[139] vdd gnd cell_6t
Xbit_r140_c44 bl[44] br[44] wl[140] vdd gnd cell_6t
Xbit_r141_c44 bl[44] br[44] wl[141] vdd gnd cell_6t
Xbit_r142_c44 bl[44] br[44] wl[142] vdd gnd cell_6t
Xbit_r143_c44 bl[44] br[44] wl[143] vdd gnd cell_6t
Xbit_r144_c44 bl[44] br[44] wl[144] vdd gnd cell_6t
Xbit_r145_c44 bl[44] br[44] wl[145] vdd gnd cell_6t
Xbit_r146_c44 bl[44] br[44] wl[146] vdd gnd cell_6t
Xbit_r147_c44 bl[44] br[44] wl[147] vdd gnd cell_6t
Xbit_r148_c44 bl[44] br[44] wl[148] vdd gnd cell_6t
Xbit_r149_c44 bl[44] br[44] wl[149] vdd gnd cell_6t
Xbit_r150_c44 bl[44] br[44] wl[150] vdd gnd cell_6t
Xbit_r151_c44 bl[44] br[44] wl[151] vdd gnd cell_6t
Xbit_r152_c44 bl[44] br[44] wl[152] vdd gnd cell_6t
Xbit_r153_c44 bl[44] br[44] wl[153] vdd gnd cell_6t
Xbit_r154_c44 bl[44] br[44] wl[154] vdd gnd cell_6t
Xbit_r155_c44 bl[44] br[44] wl[155] vdd gnd cell_6t
Xbit_r156_c44 bl[44] br[44] wl[156] vdd gnd cell_6t
Xbit_r157_c44 bl[44] br[44] wl[157] vdd gnd cell_6t
Xbit_r158_c44 bl[44] br[44] wl[158] vdd gnd cell_6t
Xbit_r159_c44 bl[44] br[44] wl[159] vdd gnd cell_6t
Xbit_r160_c44 bl[44] br[44] wl[160] vdd gnd cell_6t
Xbit_r161_c44 bl[44] br[44] wl[161] vdd gnd cell_6t
Xbit_r162_c44 bl[44] br[44] wl[162] vdd gnd cell_6t
Xbit_r163_c44 bl[44] br[44] wl[163] vdd gnd cell_6t
Xbit_r164_c44 bl[44] br[44] wl[164] vdd gnd cell_6t
Xbit_r165_c44 bl[44] br[44] wl[165] vdd gnd cell_6t
Xbit_r166_c44 bl[44] br[44] wl[166] vdd gnd cell_6t
Xbit_r167_c44 bl[44] br[44] wl[167] vdd gnd cell_6t
Xbit_r168_c44 bl[44] br[44] wl[168] vdd gnd cell_6t
Xbit_r169_c44 bl[44] br[44] wl[169] vdd gnd cell_6t
Xbit_r170_c44 bl[44] br[44] wl[170] vdd gnd cell_6t
Xbit_r171_c44 bl[44] br[44] wl[171] vdd gnd cell_6t
Xbit_r172_c44 bl[44] br[44] wl[172] vdd gnd cell_6t
Xbit_r173_c44 bl[44] br[44] wl[173] vdd gnd cell_6t
Xbit_r174_c44 bl[44] br[44] wl[174] vdd gnd cell_6t
Xbit_r175_c44 bl[44] br[44] wl[175] vdd gnd cell_6t
Xbit_r176_c44 bl[44] br[44] wl[176] vdd gnd cell_6t
Xbit_r177_c44 bl[44] br[44] wl[177] vdd gnd cell_6t
Xbit_r178_c44 bl[44] br[44] wl[178] vdd gnd cell_6t
Xbit_r179_c44 bl[44] br[44] wl[179] vdd gnd cell_6t
Xbit_r180_c44 bl[44] br[44] wl[180] vdd gnd cell_6t
Xbit_r181_c44 bl[44] br[44] wl[181] vdd gnd cell_6t
Xbit_r182_c44 bl[44] br[44] wl[182] vdd gnd cell_6t
Xbit_r183_c44 bl[44] br[44] wl[183] vdd gnd cell_6t
Xbit_r184_c44 bl[44] br[44] wl[184] vdd gnd cell_6t
Xbit_r185_c44 bl[44] br[44] wl[185] vdd gnd cell_6t
Xbit_r186_c44 bl[44] br[44] wl[186] vdd gnd cell_6t
Xbit_r187_c44 bl[44] br[44] wl[187] vdd gnd cell_6t
Xbit_r188_c44 bl[44] br[44] wl[188] vdd gnd cell_6t
Xbit_r189_c44 bl[44] br[44] wl[189] vdd gnd cell_6t
Xbit_r190_c44 bl[44] br[44] wl[190] vdd gnd cell_6t
Xbit_r191_c44 bl[44] br[44] wl[191] vdd gnd cell_6t
Xbit_r192_c44 bl[44] br[44] wl[192] vdd gnd cell_6t
Xbit_r193_c44 bl[44] br[44] wl[193] vdd gnd cell_6t
Xbit_r194_c44 bl[44] br[44] wl[194] vdd gnd cell_6t
Xbit_r195_c44 bl[44] br[44] wl[195] vdd gnd cell_6t
Xbit_r196_c44 bl[44] br[44] wl[196] vdd gnd cell_6t
Xbit_r197_c44 bl[44] br[44] wl[197] vdd gnd cell_6t
Xbit_r198_c44 bl[44] br[44] wl[198] vdd gnd cell_6t
Xbit_r199_c44 bl[44] br[44] wl[199] vdd gnd cell_6t
Xbit_r200_c44 bl[44] br[44] wl[200] vdd gnd cell_6t
Xbit_r201_c44 bl[44] br[44] wl[201] vdd gnd cell_6t
Xbit_r202_c44 bl[44] br[44] wl[202] vdd gnd cell_6t
Xbit_r203_c44 bl[44] br[44] wl[203] vdd gnd cell_6t
Xbit_r204_c44 bl[44] br[44] wl[204] vdd gnd cell_6t
Xbit_r205_c44 bl[44] br[44] wl[205] vdd gnd cell_6t
Xbit_r206_c44 bl[44] br[44] wl[206] vdd gnd cell_6t
Xbit_r207_c44 bl[44] br[44] wl[207] vdd gnd cell_6t
Xbit_r208_c44 bl[44] br[44] wl[208] vdd gnd cell_6t
Xbit_r209_c44 bl[44] br[44] wl[209] vdd gnd cell_6t
Xbit_r210_c44 bl[44] br[44] wl[210] vdd gnd cell_6t
Xbit_r211_c44 bl[44] br[44] wl[211] vdd gnd cell_6t
Xbit_r212_c44 bl[44] br[44] wl[212] vdd gnd cell_6t
Xbit_r213_c44 bl[44] br[44] wl[213] vdd gnd cell_6t
Xbit_r214_c44 bl[44] br[44] wl[214] vdd gnd cell_6t
Xbit_r215_c44 bl[44] br[44] wl[215] vdd gnd cell_6t
Xbit_r216_c44 bl[44] br[44] wl[216] vdd gnd cell_6t
Xbit_r217_c44 bl[44] br[44] wl[217] vdd gnd cell_6t
Xbit_r218_c44 bl[44] br[44] wl[218] vdd gnd cell_6t
Xbit_r219_c44 bl[44] br[44] wl[219] vdd gnd cell_6t
Xbit_r220_c44 bl[44] br[44] wl[220] vdd gnd cell_6t
Xbit_r221_c44 bl[44] br[44] wl[221] vdd gnd cell_6t
Xbit_r222_c44 bl[44] br[44] wl[222] vdd gnd cell_6t
Xbit_r223_c44 bl[44] br[44] wl[223] vdd gnd cell_6t
Xbit_r224_c44 bl[44] br[44] wl[224] vdd gnd cell_6t
Xbit_r225_c44 bl[44] br[44] wl[225] vdd gnd cell_6t
Xbit_r226_c44 bl[44] br[44] wl[226] vdd gnd cell_6t
Xbit_r227_c44 bl[44] br[44] wl[227] vdd gnd cell_6t
Xbit_r228_c44 bl[44] br[44] wl[228] vdd gnd cell_6t
Xbit_r229_c44 bl[44] br[44] wl[229] vdd gnd cell_6t
Xbit_r230_c44 bl[44] br[44] wl[230] vdd gnd cell_6t
Xbit_r231_c44 bl[44] br[44] wl[231] vdd gnd cell_6t
Xbit_r232_c44 bl[44] br[44] wl[232] vdd gnd cell_6t
Xbit_r233_c44 bl[44] br[44] wl[233] vdd gnd cell_6t
Xbit_r234_c44 bl[44] br[44] wl[234] vdd gnd cell_6t
Xbit_r235_c44 bl[44] br[44] wl[235] vdd gnd cell_6t
Xbit_r236_c44 bl[44] br[44] wl[236] vdd gnd cell_6t
Xbit_r237_c44 bl[44] br[44] wl[237] vdd gnd cell_6t
Xbit_r238_c44 bl[44] br[44] wl[238] vdd gnd cell_6t
Xbit_r239_c44 bl[44] br[44] wl[239] vdd gnd cell_6t
Xbit_r240_c44 bl[44] br[44] wl[240] vdd gnd cell_6t
Xbit_r241_c44 bl[44] br[44] wl[241] vdd gnd cell_6t
Xbit_r242_c44 bl[44] br[44] wl[242] vdd gnd cell_6t
Xbit_r243_c44 bl[44] br[44] wl[243] vdd gnd cell_6t
Xbit_r244_c44 bl[44] br[44] wl[244] vdd gnd cell_6t
Xbit_r245_c44 bl[44] br[44] wl[245] vdd gnd cell_6t
Xbit_r246_c44 bl[44] br[44] wl[246] vdd gnd cell_6t
Xbit_r247_c44 bl[44] br[44] wl[247] vdd gnd cell_6t
Xbit_r248_c44 bl[44] br[44] wl[248] vdd gnd cell_6t
Xbit_r249_c44 bl[44] br[44] wl[249] vdd gnd cell_6t
Xbit_r250_c44 bl[44] br[44] wl[250] vdd gnd cell_6t
Xbit_r251_c44 bl[44] br[44] wl[251] vdd gnd cell_6t
Xbit_r252_c44 bl[44] br[44] wl[252] vdd gnd cell_6t
Xbit_r253_c44 bl[44] br[44] wl[253] vdd gnd cell_6t
Xbit_r254_c44 bl[44] br[44] wl[254] vdd gnd cell_6t
Xbit_r255_c44 bl[44] br[44] wl[255] vdd gnd cell_6t
Xbit_r256_c44 bl[44] br[44] wl[256] vdd gnd cell_6t
Xbit_r257_c44 bl[44] br[44] wl[257] vdd gnd cell_6t
Xbit_r258_c44 bl[44] br[44] wl[258] vdd gnd cell_6t
Xbit_r259_c44 bl[44] br[44] wl[259] vdd gnd cell_6t
Xbit_r260_c44 bl[44] br[44] wl[260] vdd gnd cell_6t
Xbit_r261_c44 bl[44] br[44] wl[261] vdd gnd cell_6t
Xbit_r262_c44 bl[44] br[44] wl[262] vdd gnd cell_6t
Xbit_r263_c44 bl[44] br[44] wl[263] vdd gnd cell_6t
Xbit_r264_c44 bl[44] br[44] wl[264] vdd gnd cell_6t
Xbit_r265_c44 bl[44] br[44] wl[265] vdd gnd cell_6t
Xbit_r266_c44 bl[44] br[44] wl[266] vdd gnd cell_6t
Xbit_r267_c44 bl[44] br[44] wl[267] vdd gnd cell_6t
Xbit_r268_c44 bl[44] br[44] wl[268] vdd gnd cell_6t
Xbit_r269_c44 bl[44] br[44] wl[269] vdd gnd cell_6t
Xbit_r270_c44 bl[44] br[44] wl[270] vdd gnd cell_6t
Xbit_r271_c44 bl[44] br[44] wl[271] vdd gnd cell_6t
Xbit_r272_c44 bl[44] br[44] wl[272] vdd gnd cell_6t
Xbit_r273_c44 bl[44] br[44] wl[273] vdd gnd cell_6t
Xbit_r274_c44 bl[44] br[44] wl[274] vdd gnd cell_6t
Xbit_r275_c44 bl[44] br[44] wl[275] vdd gnd cell_6t
Xbit_r276_c44 bl[44] br[44] wl[276] vdd gnd cell_6t
Xbit_r277_c44 bl[44] br[44] wl[277] vdd gnd cell_6t
Xbit_r278_c44 bl[44] br[44] wl[278] vdd gnd cell_6t
Xbit_r279_c44 bl[44] br[44] wl[279] vdd gnd cell_6t
Xbit_r280_c44 bl[44] br[44] wl[280] vdd gnd cell_6t
Xbit_r281_c44 bl[44] br[44] wl[281] vdd gnd cell_6t
Xbit_r282_c44 bl[44] br[44] wl[282] vdd gnd cell_6t
Xbit_r283_c44 bl[44] br[44] wl[283] vdd gnd cell_6t
Xbit_r284_c44 bl[44] br[44] wl[284] vdd gnd cell_6t
Xbit_r285_c44 bl[44] br[44] wl[285] vdd gnd cell_6t
Xbit_r286_c44 bl[44] br[44] wl[286] vdd gnd cell_6t
Xbit_r287_c44 bl[44] br[44] wl[287] vdd gnd cell_6t
Xbit_r288_c44 bl[44] br[44] wl[288] vdd gnd cell_6t
Xbit_r289_c44 bl[44] br[44] wl[289] vdd gnd cell_6t
Xbit_r290_c44 bl[44] br[44] wl[290] vdd gnd cell_6t
Xbit_r291_c44 bl[44] br[44] wl[291] vdd gnd cell_6t
Xbit_r292_c44 bl[44] br[44] wl[292] vdd gnd cell_6t
Xbit_r293_c44 bl[44] br[44] wl[293] vdd gnd cell_6t
Xbit_r294_c44 bl[44] br[44] wl[294] vdd gnd cell_6t
Xbit_r295_c44 bl[44] br[44] wl[295] vdd gnd cell_6t
Xbit_r296_c44 bl[44] br[44] wl[296] vdd gnd cell_6t
Xbit_r297_c44 bl[44] br[44] wl[297] vdd gnd cell_6t
Xbit_r298_c44 bl[44] br[44] wl[298] vdd gnd cell_6t
Xbit_r299_c44 bl[44] br[44] wl[299] vdd gnd cell_6t
Xbit_r300_c44 bl[44] br[44] wl[300] vdd gnd cell_6t
Xbit_r301_c44 bl[44] br[44] wl[301] vdd gnd cell_6t
Xbit_r302_c44 bl[44] br[44] wl[302] vdd gnd cell_6t
Xbit_r303_c44 bl[44] br[44] wl[303] vdd gnd cell_6t
Xbit_r304_c44 bl[44] br[44] wl[304] vdd gnd cell_6t
Xbit_r305_c44 bl[44] br[44] wl[305] vdd gnd cell_6t
Xbit_r306_c44 bl[44] br[44] wl[306] vdd gnd cell_6t
Xbit_r307_c44 bl[44] br[44] wl[307] vdd gnd cell_6t
Xbit_r308_c44 bl[44] br[44] wl[308] vdd gnd cell_6t
Xbit_r309_c44 bl[44] br[44] wl[309] vdd gnd cell_6t
Xbit_r310_c44 bl[44] br[44] wl[310] vdd gnd cell_6t
Xbit_r311_c44 bl[44] br[44] wl[311] vdd gnd cell_6t
Xbit_r312_c44 bl[44] br[44] wl[312] vdd gnd cell_6t
Xbit_r313_c44 bl[44] br[44] wl[313] vdd gnd cell_6t
Xbit_r314_c44 bl[44] br[44] wl[314] vdd gnd cell_6t
Xbit_r315_c44 bl[44] br[44] wl[315] vdd gnd cell_6t
Xbit_r316_c44 bl[44] br[44] wl[316] vdd gnd cell_6t
Xbit_r317_c44 bl[44] br[44] wl[317] vdd gnd cell_6t
Xbit_r318_c44 bl[44] br[44] wl[318] vdd gnd cell_6t
Xbit_r319_c44 bl[44] br[44] wl[319] vdd gnd cell_6t
Xbit_r320_c44 bl[44] br[44] wl[320] vdd gnd cell_6t
Xbit_r321_c44 bl[44] br[44] wl[321] vdd gnd cell_6t
Xbit_r322_c44 bl[44] br[44] wl[322] vdd gnd cell_6t
Xbit_r323_c44 bl[44] br[44] wl[323] vdd gnd cell_6t
Xbit_r324_c44 bl[44] br[44] wl[324] vdd gnd cell_6t
Xbit_r325_c44 bl[44] br[44] wl[325] vdd gnd cell_6t
Xbit_r326_c44 bl[44] br[44] wl[326] vdd gnd cell_6t
Xbit_r327_c44 bl[44] br[44] wl[327] vdd gnd cell_6t
Xbit_r328_c44 bl[44] br[44] wl[328] vdd gnd cell_6t
Xbit_r329_c44 bl[44] br[44] wl[329] vdd gnd cell_6t
Xbit_r330_c44 bl[44] br[44] wl[330] vdd gnd cell_6t
Xbit_r331_c44 bl[44] br[44] wl[331] vdd gnd cell_6t
Xbit_r332_c44 bl[44] br[44] wl[332] vdd gnd cell_6t
Xbit_r333_c44 bl[44] br[44] wl[333] vdd gnd cell_6t
Xbit_r334_c44 bl[44] br[44] wl[334] vdd gnd cell_6t
Xbit_r335_c44 bl[44] br[44] wl[335] vdd gnd cell_6t
Xbit_r336_c44 bl[44] br[44] wl[336] vdd gnd cell_6t
Xbit_r337_c44 bl[44] br[44] wl[337] vdd gnd cell_6t
Xbit_r338_c44 bl[44] br[44] wl[338] vdd gnd cell_6t
Xbit_r339_c44 bl[44] br[44] wl[339] vdd gnd cell_6t
Xbit_r340_c44 bl[44] br[44] wl[340] vdd gnd cell_6t
Xbit_r341_c44 bl[44] br[44] wl[341] vdd gnd cell_6t
Xbit_r342_c44 bl[44] br[44] wl[342] vdd gnd cell_6t
Xbit_r343_c44 bl[44] br[44] wl[343] vdd gnd cell_6t
Xbit_r344_c44 bl[44] br[44] wl[344] vdd gnd cell_6t
Xbit_r345_c44 bl[44] br[44] wl[345] vdd gnd cell_6t
Xbit_r346_c44 bl[44] br[44] wl[346] vdd gnd cell_6t
Xbit_r347_c44 bl[44] br[44] wl[347] vdd gnd cell_6t
Xbit_r348_c44 bl[44] br[44] wl[348] vdd gnd cell_6t
Xbit_r349_c44 bl[44] br[44] wl[349] vdd gnd cell_6t
Xbit_r350_c44 bl[44] br[44] wl[350] vdd gnd cell_6t
Xbit_r351_c44 bl[44] br[44] wl[351] vdd gnd cell_6t
Xbit_r352_c44 bl[44] br[44] wl[352] vdd gnd cell_6t
Xbit_r353_c44 bl[44] br[44] wl[353] vdd gnd cell_6t
Xbit_r354_c44 bl[44] br[44] wl[354] vdd gnd cell_6t
Xbit_r355_c44 bl[44] br[44] wl[355] vdd gnd cell_6t
Xbit_r356_c44 bl[44] br[44] wl[356] vdd gnd cell_6t
Xbit_r357_c44 bl[44] br[44] wl[357] vdd gnd cell_6t
Xbit_r358_c44 bl[44] br[44] wl[358] vdd gnd cell_6t
Xbit_r359_c44 bl[44] br[44] wl[359] vdd gnd cell_6t
Xbit_r360_c44 bl[44] br[44] wl[360] vdd gnd cell_6t
Xbit_r361_c44 bl[44] br[44] wl[361] vdd gnd cell_6t
Xbit_r362_c44 bl[44] br[44] wl[362] vdd gnd cell_6t
Xbit_r363_c44 bl[44] br[44] wl[363] vdd gnd cell_6t
Xbit_r364_c44 bl[44] br[44] wl[364] vdd gnd cell_6t
Xbit_r365_c44 bl[44] br[44] wl[365] vdd gnd cell_6t
Xbit_r366_c44 bl[44] br[44] wl[366] vdd gnd cell_6t
Xbit_r367_c44 bl[44] br[44] wl[367] vdd gnd cell_6t
Xbit_r368_c44 bl[44] br[44] wl[368] vdd gnd cell_6t
Xbit_r369_c44 bl[44] br[44] wl[369] vdd gnd cell_6t
Xbit_r370_c44 bl[44] br[44] wl[370] vdd gnd cell_6t
Xbit_r371_c44 bl[44] br[44] wl[371] vdd gnd cell_6t
Xbit_r372_c44 bl[44] br[44] wl[372] vdd gnd cell_6t
Xbit_r373_c44 bl[44] br[44] wl[373] vdd gnd cell_6t
Xbit_r374_c44 bl[44] br[44] wl[374] vdd gnd cell_6t
Xbit_r375_c44 bl[44] br[44] wl[375] vdd gnd cell_6t
Xbit_r376_c44 bl[44] br[44] wl[376] vdd gnd cell_6t
Xbit_r377_c44 bl[44] br[44] wl[377] vdd gnd cell_6t
Xbit_r378_c44 bl[44] br[44] wl[378] vdd gnd cell_6t
Xbit_r379_c44 bl[44] br[44] wl[379] vdd gnd cell_6t
Xbit_r380_c44 bl[44] br[44] wl[380] vdd gnd cell_6t
Xbit_r381_c44 bl[44] br[44] wl[381] vdd gnd cell_6t
Xbit_r382_c44 bl[44] br[44] wl[382] vdd gnd cell_6t
Xbit_r383_c44 bl[44] br[44] wl[383] vdd gnd cell_6t
Xbit_r384_c44 bl[44] br[44] wl[384] vdd gnd cell_6t
Xbit_r385_c44 bl[44] br[44] wl[385] vdd gnd cell_6t
Xbit_r386_c44 bl[44] br[44] wl[386] vdd gnd cell_6t
Xbit_r387_c44 bl[44] br[44] wl[387] vdd gnd cell_6t
Xbit_r388_c44 bl[44] br[44] wl[388] vdd gnd cell_6t
Xbit_r389_c44 bl[44] br[44] wl[389] vdd gnd cell_6t
Xbit_r390_c44 bl[44] br[44] wl[390] vdd gnd cell_6t
Xbit_r391_c44 bl[44] br[44] wl[391] vdd gnd cell_6t
Xbit_r392_c44 bl[44] br[44] wl[392] vdd gnd cell_6t
Xbit_r393_c44 bl[44] br[44] wl[393] vdd gnd cell_6t
Xbit_r394_c44 bl[44] br[44] wl[394] vdd gnd cell_6t
Xbit_r395_c44 bl[44] br[44] wl[395] vdd gnd cell_6t
Xbit_r396_c44 bl[44] br[44] wl[396] vdd gnd cell_6t
Xbit_r397_c44 bl[44] br[44] wl[397] vdd gnd cell_6t
Xbit_r398_c44 bl[44] br[44] wl[398] vdd gnd cell_6t
Xbit_r399_c44 bl[44] br[44] wl[399] vdd gnd cell_6t
Xbit_r400_c44 bl[44] br[44] wl[400] vdd gnd cell_6t
Xbit_r401_c44 bl[44] br[44] wl[401] vdd gnd cell_6t
Xbit_r402_c44 bl[44] br[44] wl[402] vdd gnd cell_6t
Xbit_r403_c44 bl[44] br[44] wl[403] vdd gnd cell_6t
Xbit_r404_c44 bl[44] br[44] wl[404] vdd gnd cell_6t
Xbit_r405_c44 bl[44] br[44] wl[405] vdd gnd cell_6t
Xbit_r406_c44 bl[44] br[44] wl[406] vdd gnd cell_6t
Xbit_r407_c44 bl[44] br[44] wl[407] vdd gnd cell_6t
Xbit_r408_c44 bl[44] br[44] wl[408] vdd gnd cell_6t
Xbit_r409_c44 bl[44] br[44] wl[409] vdd gnd cell_6t
Xbit_r410_c44 bl[44] br[44] wl[410] vdd gnd cell_6t
Xbit_r411_c44 bl[44] br[44] wl[411] vdd gnd cell_6t
Xbit_r412_c44 bl[44] br[44] wl[412] vdd gnd cell_6t
Xbit_r413_c44 bl[44] br[44] wl[413] vdd gnd cell_6t
Xbit_r414_c44 bl[44] br[44] wl[414] vdd gnd cell_6t
Xbit_r415_c44 bl[44] br[44] wl[415] vdd gnd cell_6t
Xbit_r416_c44 bl[44] br[44] wl[416] vdd gnd cell_6t
Xbit_r417_c44 bl[44] br[44] wl[417] vdd gnd cell_6t
Xbit_r418_c44 bl[44] br[44] wl[418] vdd gnd cell_6t
Xbit_r419_c44 bl[44] br[44] wl[419] vdd gnd cell_6t
Xbit_r420_c44 bl[44] br[44] wl[420] vdd gnd cell_6t
Xbit_r421_c44 bl[44] br[44] wl[421] vdd gnd cell_6t
Xbit_r422_c44 bl[44] br[44] wl[422] vdd gnd cell_6t
Xbit_r423_c44 bl[44] br[44] wl[423] vdd gnd cell_6t
Xbit_r424_c44 bl[44] br[44] wl[424] vdd gnd cell_6t
Xbit_r425_c44 bl[44] br[44] wl[425] vdd gnd cell_6t
Xbit_r426_c44 bl[44] br[44] wl[426] vdd gnd cell_6t
Xbit_r427_c44 bl[44] br[44] wl[427] vdd gnd cell_6t
Xbit_r428_c44 bl[44] br[44] wl[428] vdd gnd cell_6t
Xbit_r429_c44 bl[44] br[44] wl[429] vdd gnd cell_6t
Xbit_r430_c44 bl[44] br[44] wl[430] vdd gnd cell_6t
Xbit_r431_c44 bl[44] br[44] wl[431] vdd gnd cell_6t
Xbit_r432_c44 bl[44] br[44] wl[432] vdd gnd cell_6t
Xbit_r433_c44 bl[44] br[44] wl[433] vdd gnd cell_6t
Xbit_r434_c44 bl[44] br[44] wl[434] vdd gnd cell_6t
Xbit_r435_c44 bl[44] br[44] wl[435] vdd gnd cell_6t
Xbit_r436_c44 bl[44] br[44] wl[436] vdd gnd cell_6t
Xbit_r437_c44 bl[44] br[44] wl[437] vdd gnd cell_6t
Xbit_r438_c44 bl[44] br[44] wl[438] vdd gnd cell_6t
Xbit_r439_c44 bl[44] br[44] wl[439] vdd gnd cell_6t
Xbit_r440_c44 bl[44] br[44] wl[440] vdd gnd cell_6t
Xbit_r441_c44 bl[44] br[44] wl[441] vdd gnd cell_6t
Xbit_r442_c44 bl[44] br[44] wl[442] vdd gnd cell_6t
Xbit_r443_c44 bl[44] br[44] wl[443] vdd gnd cell_6t
Xbit_r444_c44 bl[44] br[44] wl[444] vdd gnd cell_6t
Xbit_r445_c44 bl[44] br[44] wl[445] vdd gnd cell_6t
Xbit_r446_c44 bl[44] br[44] wl[446] vdd gnd cell_6t
Xbit_r447_c44 bl[44] br[44] wl[447] vdd gnd cell_6t
Xbit_r448_c44 bl[44] br[44] wl[448] vdd gnd cell_6t
Xbit_r449_c44 bl[44] br[44] wl[449] vdd gnd cell_6t
Xbit_r450_c44 bl[44] br[44] wl[450] vdd gnd cell_6t
Xbit_r451_c44 bl[44] br[44] wl[451] vdd gnd cell_6t
Xbit_r452_c44 bl[44] br[44] wl[452] vdd gnd cell_6t
Xbit_r453_c44 bl[44] br[44] wl[453] vdd gnd cell_6t
Xbit_r454_c44 bl[44] br[44] wl[454] vdd gnd cell_6t
Xbit_r455_c44 bl[44] br[44] wl[455] vdd gnd cell_6t
Xbit_r456_c44 bl[44] br[44] wl[456] vdd gnd cell_6t
Xbit_r457_c44 bl[44] br[44] wl[457] vdd gnd cell_6t
Xbit_r458_c44 bl[44] br[44] wl[458] vdd gnd cell_6t
Xbit_r459_c44 bl[44] br[44] wl[459] vdd gnd cell_6t
Xbit_r460_c44 bl[44] br[44] wl[460] vdd gnd cell_6t
Xbit_r461_c44 bl[44] br[44] wl[461] vdd gnd cell_6t
Xbit_r462_c44 bl[44] br[44] wl[462] vdd gnd cell_6t
Xbit_r463_c44 bl[44] br[44] wl[463] vdd gnd cell_6t
Xbit_r464_c44 bl[44] br[44] wl[464] vdd gnd cell_6t
Xbit_r465_c44 bl[44] br[44] wl[465] vdd gnd cell_6t
Xbit_r466_c44 bl[44] br[44] wl[466] vdd gnd cell_6t
Xbit_r467_c44 bl[44] br[44] wl[467] vdd gnd cell_6t
Xbit_r468_c44 bl[44] br[44] wl[468] vdd gnd cell_6t
Xbit_r469_c44 bl[44] br[44] wl[469] vdd gnd cell_6t
Xbit_r470_c44 bl[44] br[44] wl[470] vdd gnd cell_6t
Xbit_r471_c44 bl[44] br[44] wl[471] vdd gnd cell_6t
Xbit_r472_c44 bl[44] br[44] wl[472] vdd gnd cell_6t
Xbit_r473_c44 bl[44] br[44] wl[473] vdd gnd cell_6t
Xbit_r474_c44 bl[44] br[44] wl[474] vdd gnd cell_6t
Xbit_r475_c44 bl[44] br[44] wl[475] vdd gnd cell_6t
Xbit_r476_c44 bl[44] br[44] wl[476] vdd gnd cell_6t
Xbit_r477_c44 bl[44] br[44] wl[477] vdd gnd cell_6t
Xbit_r478_c44 bl[44] br[44] wl[478] vdd gnd cell_6t
Xbit_r479_c44 bl[44] br[44] wl[479] vdd gnd cell_6t
Xbit_r480_c44 bl[44] br[44] wl[480] vdd gnd cell_6t
Xbit_r481_c44 bl[44] br[44] wl[481] vdd gnd cell_6t
Xbit_r482_c44 bl[44] br[44] wl[482] vdd gnd cell_6t
Xbit_r483_c44 bl[44] br[44] wl[483] vdd gnd cell_6t
Xbit_r484_c44 bl[44] br[44] wl[484] vdd gnd cell_6t
Xbit_r485_c44 bl[44] br[44] wl[485] vdd gnd cell_6t
Xbit_r486_c44 bl[44] br[44] wl[486] vdd gnd cell_6t
Xbit_r487_c44 bl[44] br[44] wl[487] vdd gnd cell_6t
Xbit_r488_c44 bl[44] br[44] wl[488] vdd gnd cell_6t
Xbit_r489_c44 bl[44] br[44] wl[489] vdd gnd cell_6t
Xbit_r490_c44 bl[44] br[44] wl[490] vdd gnd cell_6t
Xbit_r491_c44 bl[44] br[44] wl[491] vdd gnd cell_6t
Xbit_r492_c44 bl[44] br[44] wl[492] vdd gnd cell_6t
Xbit_r493_c44 bl[44] br[44] wl[493] vdd gnd cell_6t
Xbit_r494_c44 bl[44] br[44] wl[494] vdd gnd cell_6t
Xbit_r495_c44 bl[44] br[44] wl[495] vdd gnd cell_6t
Xbit_r496_c44 bl[44] br[44] wl[496] vdd gnd cell_6t
Xbit_r497_c44 bl[44] br[44] wl[497] vdd gnd cell_6t
Xbit_r498_c44 bl[44] br[44] wl[498] vdd gnd cell_6t
Xbit_r499_c44 bl[44] br[44] wl[499] vdd gnd cell_6t
Xbit_r500_c44 bl[44] br[44] wl[500] vdd gnd cell_6t
Xbit_r501_c44 bl[44] br[44] wl[501] vdd gnd cell_6t
Xbit_r502_c44 bl[44] br[44] wl[502] vdd gnd cell_6t
Xbit_r503_c44 bl[44] br[44] wl[503] vdd gnd cell_6t
Xbit_r504_c44 bl[44] br[44] wl[504] vdd gnd cell_6t
Xbit_r505_c44 bl[44] br[44] wl[505] vdd gnd cell_6t
Xbit_r506_c44 bl[44] br[44] wl[506] vdd gnd cell_6t
Xbit_r507_c44 bl[44] br[44] wl[507] vdd gnd cell_6t
Xbit_r508_c44 bl[44] br[44] wl[508] vdd gnd cell_6t
Xbit_r509_c44 bl[44] br[44] wl[509] vdd gnd cell_6t
Xbit_r510_c44 bl[44] br[44] wl[510] vdd gnd cell_6t
Xbit_r511_c44 bl[44] br[44] wl[511] vdd gnd cell_6t
Xbit_r0_c45 bl[45] br[45] wl[0] vdd gnd cell_6t
Xbit_r1_c45 bl[45] br[45] wl[1] vdd gnd cell_6t
Xbit_r2_c45 bl[45] br[45] wl[2] vdd gnd cell_6t
Xbit_r3_c45 bl[45] br[45] wl[3] vdd gnd cell_6t
Xbit_r4_c45 bl[45] br[45] wl[4] vdd gnd cell_6t
Xbit_r5_c45 bl[45] br[45] wl[5] vdd gnd cell_6t
Xbit_r6_c45 bl[45] br[45] wl[6] vdd gnd cell_6t
Xbit_r7_c45 bl[45] br[45] wl[7] vdd gnd cell_6t
Xbit_r8_c45 bl[45] br[45] wl[8] vdd gnd cell_6t
Xbit_r9_c45 bl[45] br[45] wl[9] vdd gnd cell_6t
Xbit_r10_c45 bl[45] br[45] wl[10] vdd gnd cell_6t
Xbit_r11_c45 bl[45] br[45] wl[11] vdd gnd cell_6t
Xbit_r12_c45 bl[45] br[45] wl[12] vdd gnd cell_6t
Xbit_r13_c45 bl[45] br[45] wl[13] vdd gnd cell_6t
Xbit_r14_c45 bl[45] br[45] wl[14] vdd gnd cell_6t
Xbit_r15_c45 bl[45] br[45] wl[15] vdd gnd cell_6t
Xbit_r16_c45 bl[45] br[45] wl[16] vdd gnd cell_6t
Xbit_r17_c45 bl[45] br[45] wl[17] vdd gnd cell_6t
Xbit_r18_c45 bl[45] br[45] wl[18] vdd gnd cell_6t
Xbit_r19_c45 bl[45] br[45] wl[19] vdd gnd cell_6t
Xbit_r20_c45 bl[45] br[45] wl[20] vdd gnd cell_6t
Xbit_r21_c45 bl[45] br[45] wl[21] vdd gnd cell_6t
Xbit_r22_c45 bl[45] br[45] wl[22] vdd gnd cell_6t
Xbit_r23_c45 bl[45] br[45] wl[23] vdd gnd cell_6t
Xbit_r24_c45 bl[45] br[45] wl[24] vdd gnd cell_6t
Xbit_r25_c45 bl[45] br[45] wl[25] vdd gnd cell_6t
Xbit_r26_c45 bl[45] br[45] wl[26] vdd gnd cell_6t
Xbit_r27_c45 bl[45] br[45] wl[27] vdd gnd cell_6t
Xbit_r28_c45 bl[45] br[45] wl[28] vdd gnd cell_6t
Xbit_r29_c45 bl[45] br[45] wl[29] vdd gnd cell_6t
Xbit_r30_c45 bl[45] br[45] wl[30] vdd gnd cell_6t
Xbit_r31_c45 bl[45] br[45] wl[31] vdd gnd cell_6t
Xbit_r32_c45 bl[45] br[45] wl[32] vdd gnd cell_6t
Xbit_r33_c45 bl[45] br[45] wl[33] vdd gnd cell_6t
Xbit_r34_c45 bl[45] br[45] wl[34] vdd gnd cell_6t
Xbit_r35_c45 bl[45] br[45] wl[35] vdd gnd cell_6t
Xbit_r36_c45 bl[45] br[45] wl[36] vdd gnd cell_6t
Xbit_r37_c45 bl[45] br[45] wl[37] vdd gnd cell_6t
Xbit_r38_c45 bl[45] br[45] wl[38] vdd gnd cell_6t
Xbit_r39_c45 bl[45] br[45] wl[39] vdd gnd cell_6t
Xbit_r40_c45 bl[45] br[45] wl[40] vdd gnd cell_6t
Xbit_r41_c45 bl[45] br[45] wl[41] vdd gnd cell_6t
Xbit_r42_c45 bl[45] br[45] wl[42] vdd gnd cell_6t
Xbit_r43_c45 bl[45] br[45] wl[43] vdd gnd cell_6t
Xbit_r44_c45 bl[45] br[45] wl[44] vdd gnd cell_6t
Xbit_r45_c45 bl[45] br[45] wl[45] vdd gnd cell_6t
Xbit_r46_c45 bl[45] br[45] wl[46] vdd gnd cell_6t
Xbit_r47_c45 bl[45] br[45] wl[47] vdd gnd cell_6t
Xbit_r48_c45 bl[45] br[45] wl[48] vdd gnd cell_6t
Xbit_r49_c45 bl[45] br[45] wl[49] vdd gnd cell_6t
Xbit_r50_c45 bl[45] br[45] wl[50] vdd gnd cell_6t
Xbit_r51_c45 bl[45] br[45] wl[51] vdd gnd cell_6t
Xbit_r52_c45 bl[45] br[45] wl[52] vdd gnd cell_6t
Xbit_r53_c45 bl[45] br[45] wl[53] vdd gnd cell_6t
Xbit_r54_c45 bl[45] br[45] wl[54] vdd gnd cell_6t
Xbit_r55_c45 bl[45] br[45] wl[55] vdd gnd cell_6t
Xbit_r56_c45 bl[45] br[45] wl[56] vdd gnd cell_6t
Xbit_r57_c45 bl[45] br[45] wl[57] vdd gnd cell_6t
Xbit_r58_c45 bl[45] br[45] wl[58] vdd gnd cell_6t
Xbit_r59_c45 bl[45] br[45] wl[59] vdd gnd cell_6t
Xbit_r60_c45 bl[45] br[45] wl[60] vdd gnd cell_6t
Xbit_r61_c45 bl[45] br[45] wl[61] vdd gnd cell_6t
Xbit_r62_c45 bl[45] br[45] wl[62] vdd gnd cell_6t
Xbit_r63_c45 bl[45] br[45] wl[63] vdd gnd cell_6t
Xbit_r64_c45 bl[45] br[45] wl[64] vdd gnd cell_6t
Xbit_r65_c45 bl[45] br[45] wl[65] vdd gnd cell_6t
Xbit_r66_c45 bl[45] br[45] wl[66] vdd gnd cell_6t
Xbit_r67_c45 bl[45] br[45] wl[67] vdd gnd cell_6t
Xbit_r68_c45 bl[45] br[45] wl[68] vdd gnd cell_6t
Xbit_r69_c45 bl[45] br[45] wl[69] vdd gnd cell_6t
Xbit_r70_c45 bl[45] br[45] wl[70] vdd gnd cell_6t
Xbit_r71_c45 bl[45] br[45] wl[71] vdd gnd cell_6t
Xbit_r72_c45 bl[45] br[45] wl[72] vdd gnd cell_6t
Xbit_r73_c45 bl[45] br[45] wl[73] vdd gnd cell_6t
Xbit_r74_c45 bl[45] br[45] wl[74] vdd gnd cell_6t
Xbit_r75_c45 bl[45] br[45] wl[75] vdd gnd cell_6t
Xbit_r76_c45 bl[45] br[45] wl[76] vdd gnd cell_6t
Xbit_r77_c45 bl[45] br[45] wl[77] vdd gnd cell_6t
Xbit_r78_c45 bl[45] br[45] wl[78] vdd gnd cell_6t
Xbit_r79_c45 bl[45] br[45] wl[79] vdd gnd cell_6t
Xbit_r80_c45 bl[45] br[45] wl[80] vdd gnd cell_6t
Xbit_r81_c45 bl[45] br[45] wl[81] vdd gnd cell_6t
Xbit_r82_c45 bl[45] br[45] wl[82] vdd gnd cell_6t
Xbit_r83_c45 bl[45] br[45] wl[83] vdd gnd cell_6t
Xbit_r84_c45 bl[45] br[45] wl[84] vdd gnd cell_6t
Xbit_r85_c45 bl[45] br[45] wl[85] vdd gnd cell_6t
Xbit_r86_c45 bl[45] br[45] wl[86] vdd gnd cell_6t
Xbit_r87_c45 bl[45] br[45] wl[87] vdd gnd cell_6t
Xbit_r88_c45 bl[45] br[45] wl[88] vdd gnd cell_6t
Xbit_r89_c45 bl[45] br[45] wl[89] vdd gnd cell_6t
Xbit_r90_c45 bl[45] br[45] wl[90] vdd gnd cell_6t
Xbit_r91_c45 bl[45] br[45] wl[91] vdd gnd cell_6t
Xbit_r92_c45 bl[45] br[45] wl[92] vdd gnd cell_6t
Xbit_r93_c45 bl[45] br[45] wl[93] vdd gnd cell_6t
Xbit_r94_c45 bl[45] br[45] wl[94] vdd gnd cell_6t
Xbit_r95_c45 bl[45] br[45] wl[95] vdd gnd cell_6t
Xbit_r96_c45 bl[45] br[45] wl[96] vdd gnd cell_6t
Xbit_r97_c45 bl[45] br[45] wl[97] vdd gnd cell_6t
Xbit_r98_c45 bl[45] br[45] wl[98] vdd gnd cell_6t
Xbit_r99_c45 bl[45] br[45] wl[99] vdd gnd cell_6t
Xbit_r100_c45 bl[45] br[45] wl[100] vdd gnd cell_6t
Xbit_r101_c45 bl[45] br[45] wl[101] vdd gnd cell_6t
Xbit_r102_c45 bl[45] br[45] wl[102] vdd gnd cell_6t
Xbit_r103_c45 bl[45] br[45] wl[103] vdd gnd cell_6t
Xbit_r104_c45 bl[45] br[45] wl[104] vdd gnd cell_6t
Xbit_r105_c45 bl[45] br[45] wl[105] vdd gnd cell_6t
Xbit_r106_c45 bl[45] br[45] wl[106] vdd gnd cell_6t
Xbit_r107_c45 bl[45] br[45] wl[107] vdd gnd cell_6t
Xbit_r108_c45 bl[45] br[45] wl[108] vdd gnd cell_6t
Xbit_r109_c45 bl[45] br[45] wl[109] vdd gnd cell_6t
Xbit_r110_c45 bl[45] br[45] wl[110] vdd gnd cell_6t
Xbit_r111_c45 bl[45] br[45] wl[111] vdd gnd cell_6t
Xbit_r112_c45 bl[45] br[45] wl[112] vdd gnd cell_6t
Xbit_r113_c45 bl[45] br[45] wl[113] vdd gnd cell_6t
Xbit_r114_c45 bl[45] br[45] wl[114] vdd gnd cell_6t
Xbit_r115_c45 bl[45] br[45] wl[115] vdd gnd cell_6t
Xbit_r116_c45 bl[45] br[45] wl[116] vdd gnd cell_6t
Xbit_r117_c45 bl[45] br[45] wl[117] vdd gnd cell_6t
Xbit_r118_c45 bl[45] br[45] wl[118] vdd gnd cell_6t
Xbit_r119_c45 bl[45] br[45] wl[119] vdd gnd cell_6t
Xbit_r120_c45 bl[45] br[45] wl[120] vdd gnd cell_6t
Xbit_r121_c45 bl[45] br[45] wl[121] vdd gnd cell_6t
Xbit_r122_c45 bl[45] br[45] wl[122] vdd gnd cell_6t
Xbit_r123_c45 bl[45] br[45] wl[123] vdd gnd cell_6t
Xbit_r124_c45 bl[45] br[45] wl[124] vdd gnd cell_6t
Xbit_r125_c45 bl[45] br[45] wl[125] vdd gnd cell_6t
Xbit_r126_c45 bl[45] br[45] wl[126] vdd gnd cell_6t
Xbit_r127_c45 bl[45] br[45] wl[127] vdd gnd cell_6t
Xbit_r128_c45 bl[45] br[45] wl[128] vdd gnd cell_6t
Xbit_r129_c45 bl[45] br[45] wl[129] vdd gnd cell_6t
Xbit_r130_c45 bl[45] br[45] wl[130] vdd gnd cell_6t
Xbit_r131_c45 bl[45] br[45] wl[131] vdd gnd cell_6t
Xbit_r132_c45 bl[45] br[45] wl[132] vdd gnd cell_6t
Xbit_r133_c45 bl[45] br[45] wl[133] vdd gnd cell_6t
Xbit_r134_c45 bl[45] br[45] wl[134] vdd gnd cell_6t
Xbit_r135_c45 bl[45] br[45] wl[135] vdd gnd cell_6t
Xbit_r136_c45 bl[45] br[45] wl[136] vdd gnd cell_6t
Xbit_r137_c45 bl[45] br[45] wl[137] vdd gnd cell_6t
Xbit_r138_c45 bl[45] br[45] wl[138] vdd gnd cell_6t
Xbit_r139_c45 bl[45] br[45] wl[139] vdd gnd cell_6t
Xbit_r140_c45 bl[45] br[45] wl[140] vdd gnd cell_6t
Xbit_r141_c45 bl[45] br[45] wl[141] vdd gnd cell_6t
Xbit_r142_c45 bl[45] br[45] wl[142] vdd gnd cell_6t
Xbit_r143_c45 bl[45] br[45] wl[143] vdd gnd cell_6t
Xbit_r144_c45 bl[45] br[45] wl[144] vdd gnd cell_6t
Xbit_r145_c45 bl[45] br[45] wl[145] vdd gnd cell_6t
Xbit_r146_c45 bl[45] br[45] wl[146] vdd gnd cell_6t
Xbit_r147_c45 bl[45] br[45] wl[147] vdd gnd cell_6t
Xbit_r148_c45 bl[45] br[45] wl[148] vdd gnd cell_6t
Xbit_r149_c45 bl[45] br[45] wl[149] vdd gnd cell_6t
Xbit_r150_c45 bl[45] br[45] wl[150] vdd gnd cell_6t
Xbit_r151_c45 bl[45] br[45] wl[151] vdd gnd cell_6t
Xbit_r152_c45 bl[45] br[45] wl[152] vdd gnd cell_6t
Xbit_r153_c45 bl[45] br[45] wl[153] vdd gnd cell_6t
Xbit_r154_c45 bl[45] br[45] wl[154] vdd gnd cell_6t
Xbit_r155_c45 bl[45] br[45] wl[155] vdd gnd cell_6t
Xbit_r156_c45 bl[45] br[45] wl[156] vdd gnd cell_6t
Xbit_r157_c45 bl[45] br[45] wl[157] vdd gnd cell_6t
Xbit_r158_c45 bl[45] br[45] wl[158] vdd gnd cell_6t
Xbit_r159_c45 bl[45] br[45] wl[159] vdd gnd cell_6t
Xbit_r160_c45 bl[45] br[45] wl[160] vdd gnd cell_6t
Xbit_r161_c45 bl[45] br[45] wl[161] vdd gnd cell_6t
Xbit_r162_c45 bl[45] br[45] wl[162] vdd gnd cell_6t
Xbit_r163_c45 bl[45] br[45] wl[163] vdd gnd cell_6t
Xbit_r164_c45 bl[45] br[45] wl[164] vdd gnd cell_6t
Xbit_r165_c45 bl[45] br[45] wl[165] vdd gnd cell_6t
Xbit_r166_c45 bl[45] br[45] wl[166] vdd gnd cell_6t
Xbit_r167_c45 bl[45] br[45] wl[167] vdd gnd cell_6t
Xbit_r168_c45 bl[45] br[45] wl[168] vdd gnd cell_6t
Xbit_r169_c45 bl[45] br[45] wl[169] vdd gnd cell_6t
Xbit_r170_c45 bl[45] br[45] wl[170] vdd gnd cell_6t
Xbit_r171_c45 bl[45] br[45] wl[171] vdd gnd cell_6t
Xbit_r172_c45 bl[45] br[45] wl[172] vdd gnd cell_6t
Xbit_r173_c45 bl[45] br[45] wl[173] vdd gnd cell_6t
Xbit_r174_c45 bl[45] br[45] wl[174] vdd gnd cell_6t
Xbit_r175_c45 bl[45] br[45] wl[175] vdd gnd cell_6t
Xbit_r176_c45 bl[45] br[45] wl[176] vdd gnd cell_6t
Xbit_r177_c45 bl[45] br[45] wl[177] vdd gnd cell_6t
Xbit_r178_c45 bl[45] br[45] wl[178] vdd gnd cell_6t
Xbit_r179_c45 bl[45] br[45] wl[179] vdd gnd cell_6t
Xbit_r180_c45 bl[45] br[45] wl[180] vdd gnd cell_6t
Xbit_r181_c45 bl[45] br[45] wl[181] vdd gnd cell_6t
Xbit_r182_c45 bl[45] br[45] wl[182] vdd gnd cell_6t
Xbit_r183_c45 bl[45] br[45] wl[183] vdd gnd cell_6t
Xbit_r184_c45 bl[45] br[45] wl[184] vdd gnd cell_6t
Xbit_r185_c45 bl[45] br[45] wl[185] vdd gnd cell_6t
Xbit_r186_c45 bl[45] br[45] wl[186] vdd gnd cell_6t
Xbit_r187_c45 bl[45] br[45] wl[187] vdd gnd cell_6t
Xbit_r188_c45 bl[45] br[45] wl[188] vdd gnd cell_6t
Xbit_r189_c45 bl[45] br[45] wl[189] vdd gnd cell_6t
Xbit_r190_c45 bl[45] br[45] wl[190] vdd gnd cell_6t
Xbit_r191_c45 bl[45] br[45] wl[191] vdd gnd cell_6t
Xbit_r192_c45 bl[45] br[45] wl[192] vdd gnd cell_6t
Xbit_r193_c45 bl[45] br[45] wl[193] vdd gnd cell_6t
Xbit_r194_c45 bl[45] br[45] wl[194] vdd gnd cell_6t
Xbit_r195_c45 bl[45] br[45] wl[195] vdd gnd cell_6t
Xbit_r196_c45 bl[45] br[45] wl[196] vdd gnd cell_6t
Xbit_r197_c45 bl[45] br[45] wl[197] vdd gnd cell_6t
Xbit_r198_c45 bl[45] br[45] wl[198] vdd gnd cell_6t
Xbit_r199_c45 bl[45] br[45] wl[199] vdd gnd cell_6t
Xbit_r200_c45 bl[45] br[45] wl[200] vdd gnd cell_6t
Xbit_r201_c45 bl[45] br[45] wl[201] vdd gnd cell_6t
Xbit_r202_c45 bl[45] br[45] wl[202] vdd gnd cell_6t
Xbit_r203_c45 bl[45] br[45] wl[203] vdd gnd cell_6t
Xbit_r204_c45 bl[45] br[45] wl[204] vdd gnd cell_6t
Xbit_r205_c45 bl[45] br[45] wl[205] vdd gnd cell_6t
Xbit_r206_c45 bl[45] br[45] wl[206] vdd gnd cell_6t
Xbit_r207_c45 bl[45] br[45] wl[207] vdd gnd cell_6t
Xbit_r208_c45 bl[45] br[45] wl[208] vdd gnd cell_6t
Xbit_r209_c45 bl[45] br[45] wl[209] vdd gnd cell_6t
Xbit_r210_c45 bl[45] br[45] wl[210] vdd gnd cell_6t
Xbit_r211_c45 bl[45] br[45] wl[211] vdd gnd cell_6t
Xbit_r212_c45 bl[45] br[45] wl[212] vdd gnd cell_6t
Xbit_r213_c45 bl[45] br[45] wl[213] vdd gnd cell_6t
Xbit_r214_c45 bl[45] br[45] wl[214] vdd gnd cell_6t
Xbit_r215_c45 bl[45] br[45] wl[215] vdd gnd cell_6t
Xbit_r216_c45 bl[45] br[45] wl[216] vdd gnd cell_6t
Xbit_r217_c45 bl[45] br[45] wl[217] vdd gnd cell_6t
Xbit_r218_c45 bl[45] br[45] wl[218] vdd gnd cell_6t
Xbit_r219_c45 bl[45] br[45] wl[219] vdd gnd cell_6t
Xbit_r220_c45 bl[45] br[45] wl[220] vdd gnd cell_6t
Xbit_r221_c45 bl[45] br[45] wl[221] vdd gnd cell_6t
Xbit_r222_c45 bl[45] br[45] wl[222] vdd gnd cell_6t
Xbit_r223_c45 bl[45] br[45] wl[223] vdd gnd cell_6t
Xbit_r224_c45 bl[45] br[45] wl[224] vdd gnd cell_6t
Xbit_r225_c45 bl[45] br[45] wl[225] vdd gnd cell_6t
Xbit_r226_c45 bl[45] br[45] wl[226] vdd gnd cell_6t
Xbit_r227_c45 bl[45] br[45] wl[227] vdd gnd cell_6t
Xbit_r228_c45 bl[45] br[45] wl[228] vdd gnd cell_6t
Xbit_r229_c45 bl[45] br[45] wl[229] vdd gnd cell_6t
Xbit_r230_c45 bl[45] br[45] wl[230] vdd gnd cell_6t
Xbit_r231_c45 bl[45] br[45] wl[231] vdd gnd cell_6t
Xbit_r232_c45 bl[45] br[45] wl[232] vdd gnd cell_6t
Xbit_r233_c45 bl[45] br[45] wl[233] vdd gnd cell_6t
Xbit_r234_c45 bl[45] br[45] wl[234] vdd gnd cell_6t
Xbit_r235_c45 bl[45] br[45] wl[235] vdd gnd cell_6t
Xbit_r236_c45 bl[45] br[45] wl[236] vdd gnd cell_6t
Xbit_r237_c45 bl[45] br[45] wl[237] vdd gnd cell_6t
Xbit_r238_c45 bl[45] br[45] wl[238] vdd gnd cell_6t
Xbit_r239_c45 bl[45] br[45] wl[239] vdd gnd cell_6t
Xbit_r240_c45 bl[45] br[45] wl[240] vdd gnd cell_6t
Xbit_r241_c45 bl[45] br[45] wl[241] vdd gnd cell_6t
Xbit_r242_c45 bl[45] br[45] wl[242] vdd gnd cell_6t
Xbit_r243_c45 bl[45] br[45] wl[243] vdd gnd cell_6t
Xbit_r244_c45 bl[45] br[45] wl[244] vdd gnd cell_6t
Xbit_r245_c45 bl[45] br[45] wl[245] vdd gnd cell_6t
Xbit_r246_c45 bl[45] br[45] wl[246] vdd gnd cell_6t
Xbit_r247_c45 bl[45] br[45] wl[247] vdd gnd cell_6t
Xbit_r248_c45 bl[45] br[45] wl[248] vdd gnd cell_6t
Xbit_r249_c45 bl[45] br[45] wl[249] vdd gnd cell_6t
Xbit_r250_c45 bl[45] br[45] wl[250] vdd gnd cell_6t
Xbit_r251_c45 bl[45] br[45] wl[251] vdd gnd cell_6t
Xbit_r252_c45 bl[45] br[45] wl[252] vdd gnd cell_6t
Xbit_r253_c45 bl[45] br[45] wl[253] vdd gnd cell_6t
Xbit_r254_c45 bl[45] br[45] wl[254] vdd gnd cell_6t
Xbit_r255_c45 bl[45] br[45] wl[255] vdd gnd cell_6t
Xbit_r256_c45 bl[45] br[45] wl[256] vdd gnd cell_6t
Xbit_r257_c45 bl[45] br[45] wl[257] vdd gnd cell_6t
Xbit_r258_c45 bl[45] br[45] wl[258] vdd gnd cell_6t
Xbit_r259_c45 bl[45] br[45] wl[259] vdd gnd cell_6t
Xbit_r260_c45 bl[45] br[45] wl[260] vdd gnd cell_6t
Xbit_r261_c45 bl[45] br[45] wl[261] vdd gnd cell_6t
Xbit_r262_c45 bl[45] br[45] wl[262] vdd gnd cell_6t
Xbit_r263_c45 bl[45] br[45] wl[263] vdd gnd cell_6t
Xbit_r264_c45 bl[45] br[45] wl[264] vdd gnd cell_6t
Xbit_r265_c45 bl[45] br[45] wl[265] vdd gnd cell_6t
Xbit_r266_c45 bl[45] br[45] wl[266] vdd gnd cell_6t
Xbit_r267_c45 bl[45] br[45] wl[267] vdd gnd cell_6t
Xbit_r268_c45 bl[45] br[45] wl[268] vdd gnd cell_6t
Xbit_r269_c45 bl[45] br[45] wl[269] vdd gnd cell_6t
Xbit_r270_c45 bl[45] br[45] wl[270] vdd gnd cell_6t
Xbit_r271_c45 bl[45] br[45] wl[271] vdd gnd cell_6t
Xbit_r272_c45 bl[45] br[45] wl[272] vdd gnd cell_6t
Xbit_r273_c45 bl[45] br[45] wl[273] vdd gnd cell_6t
Xbit_r274_c45 bl[45] br[45] wl[274] vdd gnd cell_6t
Xbit_r275_c45 bl[45] br[45] wl[275] vdd gnd cell_6t
Xbit_r276_c45 bl[45] br[45] wl[276] vdd gnd cell_6t
Xbit_r277_c45 bl[45] br[45] wl[277] vdd gnd cell_6t
Xbit_r278_c45 bl[45] br[45] wl[278] vdd gnd cell_6t
Xbit_r279_c45 bl[45] br[45] wl[279] vdd gnd cell_6t
Xbit_r280_c45 bl[45] br[45] wl[280] vdd gnd cell_6t
Xbit_r281_c45 bl[45] br[45] wl[281] vdd gnd cell_6t
Xbit_r282_c45 bl[45] br[45] wl[282] vdd gnd cell_6t
Xbit_r283_c45 bl[45] br[45] wl[283] vdd gnd cell_6t
Xbit_r284_c45 bl[45] br[45] wl[284] vdd gnd cell_6t
Xbit_r285_c45 bl[45] br[45] wl[285] vdd gnd cell_6t
Xbit_r286_c45 bl[45] br[45] wl[286] vdd gnd cell_6t
Xbit_r287_c45 bl[45] br[45] wl[287] vdd gnd cell_6t
Xbit_r288_c45 bl[45] br[45] wl[288] vdd gnd cell_6t
Xbit_r289_c45 bl[45] br[45] wl[289] vdd gnd cell_6t
Xbit_r290_c45 bl[45] br[45] wl[290] vdd gnd cell_6t
Xbit_r291_c45 bl[45] br[45] wl[291] vdd gnd cell_6t
Xbit_r292_c45 bl[45] br[45] wl[292] vdd gnd cell_6t
Xbit_r293_c45 bl[45] br[45] wl[293] vdd gnd cell_6t
Xbit_r294_c45 bl[45] br[45] wl[294] vdd gnd cell_6t
Xbit_r295_c45 bl[45] br[45] wl[295] vdd gnd cell_6t
Xbit_r296_c45 bl[45] br[45] wl[296] vdd gnd cell_6t
Xbit_r297_c45 bl[45] br[45] wl[297] vdd gnd cell_6t
Xbit_r298_c45 bl[45] br[45] wl[298] vdd gnd cell_6t
Xbit_r299_c45 bl[45] br[45] wl[299] vdd gnd cell_6t
Xbit_r300_c45 bl[45] br[45] wl[300] vdd gnd cell_6t
Xbit_r301_c45 bl[45] br[45] wl[301] vdd gnd cell_6t
Xbit_r302_c45 bl[45] br[45] wl[302] vdd gnd cell_6t
Xbit_r303_c45 bl[45] br[45] wl[303] vdd gnd cell_6t
Xbit_r304_c45 bl[45] br[45] wl[304] vdd gnd cell_6t
Xbit_r305_c45 bl[45] br[45] wl[305] vdd gnd cell_6t
Xbit_r306_c45 bl[45] br[45] wl[306] vdd gnd cell_6t
Xbit_r307_c45 bl[45] br[45] wl[307] vdd gnd cell_6t
Xbit_r308_c45 bl[45] br[45] wl[308] vdd gnd cell_6t
Xbit_r309_c45 bl[45] br[45] wl[309] vdd gnd cell_6t
Xbit_r310_c45 bl[45] br[45] wl[310] vdd gnd cell_6t
Xbit_r311_c45 bl[45] br[45] wl[311] vdd gnd cell_6t
Xbit_r312_c45 bl[45] br[45] wl[312] vdd gnd cell_6t
Xbit_r313_c45 bl[45] br[45] wl[313] vdd gnd cell_6t
Xbit_r314_c45 bl[45] br[45] wl[314] vdd gnd cell_6t
Xbit_r315_c45 bl[45] br[45] wl[315] vdd gnd cell_6t
Xbit_r316_c45 bl[45] br[45] wl[316] vdd gnd cell_6t
Xbit_r317_c45 bl[45] br[45] wl[317] vdd gnd cell_6t
Xbit_r318_c45 bl[45] br[45] wl[318] vdd gnd cell_6t
Xbit_r319_c45 bl[45] br[45] wl[319] vdd gnd cell_6t
Xbit_r320_c45 bl[45] br[45] wl[320] vdd gnd cell_6t
Xbit_r321_c45 bl[45] br[45] wl[321] vdd gnd cell_6t
Xbit_r322_c45 bl[45] br[45] wl[322] vdd gnd cell_6t
Xbit_r323_c45 bl[45] br[45] wl[323] vdd gnd cell_6t
Xbit_r324_c45 bl[45] br[45] wl[324] vdd gnd cell_6t
Xbit_r325_c45 bl[45] br[45] wl[325] vdd gnd cell_6t
Xbit_r326_c45 bl[45] br[45] wl[326] vdd gnd cell_6t
Xbit_r327_c45 bl[45] br[45] wl[327] vdd gnd cell_6t
Xbit_r328_c45 bl[45] br[45] wl[328] vdd gnd cell_6t
Xbit_r329_c45 bl[45] br[45] wl[329] vdd gnd cell_6t
Xbit_r330_c45 bl[45] br[45] wl[330] vdd gnd cell_6t
Xbit_r331_c45 bl[45] br[45] wl[331] vdd gnd cell_6t
Xbit_r332_c45 bl[45] br[45] wl[332] vdd gnd cell_6t
Xbit_r333_c45 bl[45] br[45] wl[333] vdd gnd cell_6t
Xbit_r334_c45 bl[45] br[45] wl[334] vdd gnd cell_6t
Xbit_r335_c45 bl[45] br[45] wl[335] vdd gnd cell_6t
Xbit_r336_c45 bl[45] br[45] wl[336] vdd gnd cell_6t
Xbit_r337_c45 bl[45] br[45] wl[337] vdd gnd cell_6t
Xbit_r338_c45 bl[45] br[45] wl[338] vdd gnd cell_6t
Xbit_r339_c45 bl[45] br[45] wl[339] vdd gnd cell_6t
Xbit_r340_c45 bl[45] br[45] wl[340] vdd gnd cell_6t
Xbit_r341_c45 bl[45] br[45] wl[341] vdd gnd cell_6t
Xbit_r342_c45 bl[45] br[45] wl[342] vdd gnd cell_6t
Xbit_r343_c45 bl[45] br[45] wl[343] vdd gnd cell_6t
Xbit_r344_c45 bl[45] br[45] wl[344] vdd gnd cell_6t
Xbit_r345_c45 bl[45] br[45] wl[345] vdd gnd cell_6t
Xbit_r346_c45 bl[45] br[45] wl[346] vdd gnd cell_6t
Xbit_r347_c45 bl[45] br[45] wl[347] vdd gnd cell_6t
Xbit_r348_c45 bl[45] br[45] wl[348] vdd gnd cell_6t
Xbit_r349_c45 bl[45] br[45] wl[349] vdd gnd cell_6t
Xbit_r350_c45 bl[45] br[45] wl[350] vdd gnd cell_6t
Xbit_r351_c45 bl[45] br[45] wl[351] vdd gnd cell_6t
Xbit_r352_c45 bl[45] br[45] wl[352] vdd gnd cell_6t
Xbit_r353_c45 bl[45] br[45] wl[353] vdd gnd cell_6t
Xbit_r354_c45 bl[45] br[45] wl[354] vdd gnd cell_6t
Xbit_r355_c45 bl[45] br[45] wl[355] vdd gnd cell_6t
Xbit_r356_c45 bl[45] br[45] wl[356] vdd gnd cell_6t
Xbit_r357_c45 bl[45] br[45] wl[357] vdd gnd cell_6t
Xbit_r358_c45 bl[45] br[45] wl[358] vdd gnd cell_6t
Xbit_r359_c45 bl[45] br[45] wl[359] vdd gnd cell_6t
Xbit_r360_c45 bl[45] br[45] wl[360] vdd gnd cell_6t
Xbit_r361_c45 bl[45] br[45] wl[361] vdd gnd cell_6t
Xbit_r362_c45 bl[45] br[45] wl[362] vdd gnd cell_6t
Xbit_r363_c45 bl[45] br[45] wl[363] vdd gnd cell_6t
Xbit_r364_c45 bl[45] br[45] wl[364] vdd gnd cell_6t
Xbit_r365_c45 bl[45] br[45] wl[365] vdd gnd cell_6t
Xbit_r366_c45 bl[45] br[45] wl[366] vdd gnd cell_6t
Xbit_r367_c45 bl[45] br[45] wl[367] vdd gnd cell_6t
Xbit_r368_c45 bl[45] br[45] wl[368] vdd gnd cell_6t
Xbit_r369_c45 bl[45] br[45] wl[369] vdd gnd cell_6t
Xbit_r370_c45 bl[45] br[45] wl[370] vdd gnd cell_6t
Xbit_r371_c45 bl[45] br[45] wl[371] vdd gnd cell_6t
Xbit_r372_c45 bl[45] br[45] wl[372] vdd gnd cell_6t
Xbit_r373_c45 bl[45] br[45] wl[373] vdd gnd cell_6t
Xbit_r374_c45 bl[45] br[45] wl[374] vdd gnd cell_6t
Xbit_r375_c45 bl[45] br[45] wl[375] vdd gnd cell_6t
Xbit_r376_c45 bl[45] br[45] wl[376] vdd gnd cell_6t
Xbit_r377_c45 bl[45] br[45] wl[377] vdd gnd cell_6t
Xbit_r378_c45 bl[45] br[45] wl[378] vdd gnd cell_6t
Xbit_r379_c45 bl[45] br[45] wl[379] vdd gnd cell_6t
Xbit_r380_c45 bl[45] br[45] wl[380] vdd gnd cell_6t
Xbit_r381_c45 bl[45] br[45] wl[381] vdd gnd cell_6t
Xbit_r382_c45 bl[45] br[45] wl[382] vdd gnd cell_6t
Xbit_r383_c45 bl[45] br[45] wl[383] vdd gnd cell_6t
Xbit_r384_c45 bl[45] br[45] wl[384] vdd gnd cell_6t
Xbit_r385_c45 bl[45] br[45] wl[385] vdd gnd cell_6t
Xbit_r386_c45 bl[45] br[45] wl[386] vdd gnd cell_6t
Xbit_r387_c45 bl[45] br[45] wl[387] vdd gnd cell_6t
Xbit_r388_c45 bl[45] br[45] wl[388] vdd gnd cell_6t
Xbit_r389_c45 bl[45] br[45] wl[389] vdd gnd cell_6t
Xbit_r390_c45 bl[45] br[45] wl[390] vdd gnd cell_6t
Xbit_r391_c45 bl[45] br[45] wl[391] vdd gnd cell_6t
Xbit_r392_c45 bl[45] br[45] wl[392] vdd gnd cell_6t
Xbit_r393_c45 bl[45] br[45] wl[393] vdd gnd cell_6t
Xbit_r394_c45 bl[45] br[45] wl[394] vdd gnd cell_6t
Xbit_r395_c45 bl[45] br[45] wl[395] vdd gnd cell_6t
Xbit_r396_c45 bl[45] br[45] wl[396] vdd gnd cell_6t
Xbit_r397_c45 bl[45] br[45] wl[397] vdd gnd cell_6t
Xbit_r398_c45 bl[45] br[45] wl[398] vdd gnd cell_6t
Xbit_r399_c45 bl[45] br[45] wl[399] vdd gnd cell_6t
Xbit_r400_c45 bl[45] br[45] wl[400] vdd gnd cell_6t
Xbit_r401_c45 bl[45] br[45] wl[401] vdd gnd cell_6t
Xbit_r402_c45 bl[45] br[45] wl[402] vdd gnd cell_6t
Xbit_r403_c45 bl[45] br[45] wl[403] vdd gnd cell_6t
Xbit_r404_c45 bl[45] br[45] wl[404] vdd gnd cell_6t
Xbit_r405_c45 bl[45] br[45] wl[405] vdd gnd cell_6t
Xbit_r406_c45 bl[45] br[45] wl[406] vdd gnd cell_6t
Xbit_r407_c45 bl[45] br[45] wl[407] vdd gnd cell_6t
Xbit_r408_c45 bl[45] br[45] wl[408] vdd gnd cell_6t
Xbit_r409_c45 bl[45] br[45] wl[409] vdd gnd cell_6t
Xbit_r410_c45 bl[45] br[45] wl[410] vdd gnd cell_6t
Xbit_r411_c45 bl[45] br[45] wl[411] vdd gnd cell_6t
Xbit_r412_c45 bl[45] br[45] wl[412] vdd gnd cell_6t
Xbit_r413_c45 bl[45] br[45] wl[413] vdd gnd cell_6t
Xbit_r414_c45 bl[45] br[45] wl[414] vdd gnd cell_6t
Xbit_r415_c45 bl[45] br[45] wl[415] vdd gnd cell_6t
Xbit_r416_c45 bl[45] br[45] wl[416] vdd gnd cell_6t
Xbit_r417_c45 bl[45] br[45] wl[417] vdd gnd cell_6t
Xbit_r418_c45 bl[45] br[45] wl[418] vdd gnd cell_6t
Xbit_r419_c45 bl[45] br[45] wl[419] vdd gnd cell_6t
Xbit_r420_c45 bl[45] br[45] wl[420] vdd gnd cell_6t
Xbit_r421_c45 bl[45] br[45] wl[421] vdd gnd cell_6t
Xbit_r422_c45 bl[45] br[45] wl[422] vdd gnd cell_6t
Xbit_r423_c45 bl[45] br[45] wl[423] vdd gnd cell_6t
Xbit_r424_c45 bl[45] br[45] wl[424] vdd gnd cell_6t
Xbit_r425_c45 bl[45] br[45] wl[425] vdd gnd cell_6t
Xbit_r426_c45 bl[45] br[45] wl[426] vdd gnd cell_6t
Xbit_r427_c45 bl[45] br[45] wl[427] vdd gnd cell_6t
Xbit_r428_c45 bl[45] br[45] wl[428] vdd gnd cell_6t
Xbit_r429_c45 bl[45] br[45] wl[429] vdd gnd cell_6t
Xbit_r430_c45 bl[45] br[45] wl[430] vdd gnd cell_6t
Xbit_r431_c45 bl[45] br[45] wl[431] vdd gnd cell_6t
Xbit_r432_c45 bl[45] br[45] wl[432] vdd gnd cell_6t
Xbit_r433_c45 bl[45] br[45] wl[433] vdd gnd cell_6t
Xbit_r434_c45 bl[45] br[45] wl[434] vdd gnd cell_6t
Xbit_r435_c45 bl[45] br[45] wl[435] vdd gnd cell_6t
Xbit_r436_c45 bl[45] br[45] wl[436] vdd gnd cell_6t
Xbit_r437_c45 bl[45] br[45] wl[437] vdd gnd cell_6t
Xbit_r438_c45 bl[45] br[45] wl[438] vdd gnd cell_6t
Xbit_r439_c45 bl[45] br[45] wl[439] vdd gnd cell_6t
Xbit_r440_c45 bl[45] br[45] wl[440] vdd gnd cell_6t
Xbit_r441_c45 bl[45] br[45] wl[441] vdd gnd cell_6t
Xbit_r442_c45 bl[45] br[45] wl[442] vdd gnd cell_6t
Xbit_r443_c45 bl[45] br[45] wl[443] vdd gnd cell_6t
Xbit_r444_c45 bl[45] br[45] wl[444] vdd gnd cell_6t
Xbit_r445_c45 bl[45] br[45] wl[445] vdd gnd cell_6t
Xbit_r446_c45 bl[45] br[45] wl[446] vdd gnd cell_6t
Xbit_r447_c45 bl[45] br[45] wl[447] vdd gnd cell_6t
Xbit_r448_c45 bl[45] br[45] wl[448] vdd gnd cell_6t
Xbit_r449_c45 bl[45] br[45] wl[449] vdd gnd cell_6t
Xbit_r450_c45 bl[45] br[45] wl[450] vdd gnd cell_6t
Xbit_r451_c45 bl[45] br[45] wl[451] vdd gnd cell_6t
Xbit_r452_c45 bl[45] br[45] wl[452] vdd gnd cell_6t
Xbit_r453_c45 bl[45] br[45] wl[453] vdd gnd cell_6t
Xbit_r454_c45 bl[45] br[45] wl[454] vdd gnd cell_6t
Xbit_r455_c45 bl[45] br[45] wl[455] vdd gnd cell_6t
Xbit_r456_c45 bl[45] br[45] wl[456] vdd gnd cell_6t
Xbit_r457_c45 bl[45] br[45] wl[457] vdd gnd cell_6t
Xbit_r458_c45 bl[45] br[45] wl[458] vdd gnd cell_6t
Xbit_r459_c45 bl[45] br[45] wl[459] vdd gnd cell_6t
Xbit_r460_c45 bl[45] br[45] wl[460] vdd gnd cell_6t
Xbit_r461_c45 bl[45] br[45] wl[461] vdd gnd cell_6t
Xbit_r462_c45 bl[45] br[45] wl[462] vdd gnd cell_6t
Xbit_r463_c45 bl[45] br[45] wl[463] vdd gnd cell_6t
Xbit_r464_c45 bl[45] br[45] wl[464] vdd gnd cell_6t
Xbit_r465_c45 bl[45] br[45] wl[465] vdd gnd cell_6t
Xbit_r466_c45 bl[45] br[45] wl[466] vdd gnd cell_6t
Xbit_r467_c45 bl[45] br[45] wl[467] vdd gnd cell_6t
Xbit_r468_c45 bl[45] br[45] wl[468] vdd gnd cell_6t
Xbit_r469_c45 bl[45] br[45] wl[469] vdd gnd cell_6t
Xbit_r470_c45 bl[45] br[45] wl[470] vdd gnd cell_6t
Xbit_r471_c45 bl[45] br[45] wl[471] vdd gnd cell_6t
Xbit_r472_c45 bl[45] br[45] wl[472] vdd gnd cell_6t
Xbit_r473_c45 bl[45] br[45] wl[473] vdd gnd cell_6t
Xbit_r474_c45 bl[45] br[45] wl[474] vdd gnd cell_6t
Xbit_r475_c45 bl[45] br[45] wl[475] vdd gnd cell_6t
Xbit_r476_c45 bl[45] br[45] wl[476] vdd gnd cell_6t
Xbit_r477_c45 bl[45] br[45] wl[477] vdd gnd cell_6t
Xbit_r478_c45 bl[45] br[45] wl[478] vdd gnd cell_6t
Xbit_r479_c45 bl[45] br[45] wl[479] vdd gnd cell_6t
Xbit_r480_c45 bl[45] br[45] wl[480] vdd gnd cell_6t
Xbit_r481_c45 bl[45] br[45] wl[481] vdd gnd cell_6t
Xbit_r482_c45 bl[45] br[45] wl[482] vdd gnd cell_6t
Xbit_r483_c45 bl[45] br[45] wl[483] vdd gnd cell_6t
Xbit_r484_c45 bl[45] br[45] wl[484] vdd gnd cell_6t
Xbit_r485_c45 bl[45] br[45] wl[485] vdd gnd cell_6t
Xbit_r486_c45 bl[45] br[45] wl[486] vdd gnd cell_6t
Xbit_r487_c45 bl[45] br[45] wl[487] vdd gnd cell_6t
Xbit_r488_c45 bl[45] br[45] wl[488] vdd gnd cell_6t
Xbit_r489_c45 bl[45] br[45] wl[489] vdd gnd cell_6t
Xbit_r490_c45 bl[45] br[45] wl[490] vdd gnd cell_6t
Xbit_r491_c45 bl[45] br[45] wl[491] vdd gnd cell_6t
Xbit_r492_c45 bl[45] br[45] wl[492] vdd gnd cell_6t
Xbit_r493_c45 bl[45] br[45] wl[493] vdd gnd cell_6t
Xbit_r494_c45 bl[45] br[45] wl[494] vdd gnd cell_6t
Xbit_r495_c45 bl[45] br[45] wl[495] vdd gnd cell_6t
Xbit_r496_c45 bl[45] br[45] wl[496] vdd gnd cell_6t
Xbit_r497_c45 bl[45] br[45] wl[497] vdd gnd cell_6t
Xbit_r498_c45 bl[45] br[45] wl[498] vdd gnd cell_6t
Xbit_r499_c45 bl[45] br[45] wl[499] vdd gnd cell_6t
Xbit_r500_c45 bl[45] br[45] wl[500] vdd gnd cell_6t
Xbit_r501_c45 bl[45] br[45] wl[501] vdd gnd cell_6t
Xbit_r502_c45 bl[45] br[45] wl[502] vdd gnd cell_6t
Xbit_r503_c45 bl[45] br[45] wl[503] vdd gnd cell_6t
Xbit_r504_c45 bl[45] br[45] wl[504] vdd gnd cell_6t
Xbit_r505_c45 bl[45] br[45] wl[505] vdd gnd cell_6t
Xbit_r506_c45 bl[45] br[45] wl[506] vdd gnd cell_6t
Xbit_r507_c45 bl[45] br[45] wl[507] vdd gnd cell_6t
Xbit_r508_c45 bl[45] br[45] wl[508] vdd gnd cell_6t
Xbit_r509_c45 bl[45] br[45] wl[509] vdd gnd cell_6t
Xbit_r510_c45 bl[45] br[45] wl[510] vdd gnd cell_6t
Xbit_r511_c45 bl[45] br[45] wl[511] vdd gnd cell_6t
Xbit_r0_c46 bl[46] br[46] wl[0] vdd gnd cell_6t
Xbit_r1_c46 bl[46] br[46] wl[1] vdd gnd cell_6t
Xbit_r2_c46 bl[46] br[46] wl[2] vdd gnd cell_6t
Xbit_r3_c46 bl[46] br[46] wl[3] vdd gnd cell_6t
Xbit_r4_c46 bl[46] br[46] wl[4] vdd gnd cell_6t
Xbit_r5_c46 bl[46] br[46] wl[5] vdd gnd cell_6t
Xbit_r6_c46 bl[46] br[46] wl[6] vdd gnd cell_6t
Xbit_r7_c46 bl[46] br[46] wl[7] vdd gnd cell_6t
Xbit_r8_c46 bl[46] br[46] wl[8] vdd gnd cell_6t
Xbit_r9_c46 bl[46] br[46] wl[9] vdd gnd cell_6t
Xbit_r10_c46 bl[46] br[46] wl[10] vdd gnd cell_6t
Xbit_r11_c46 bl[46] br[46] wl[11] vdd gnd cell_6t
Xbit_r12_c46 bl[46] br[46] wl[12] vdd gnd cell_6t
Xbit_r13_c46 bl[46] br[46] wl[13] vdd gnd cell_6t
Xbit_r14_c46 bl[46] br[46] wl[14] vdd gnd cell_6t
Xbit_r15_c46 bl[46] br[46] wl[15] vdd gnd cell_6t
Xbit_r16_c46 bl[46] br[46] wl[16] vdd gnd cell_6t
Xbit_r17_c46 bl[46] br[46] wl[17] vdd gnd cell_6t
Xbit_r18_c46 bl[46] br[46] wl[18] vdd gnd cell_6t
Xbit_r19_c46 bl[46] br[46] wl[19] vdd gnd cell_6t
Xbit_r20_c46 bl[46] br[46] wl[20] vdd gnd cell_6t
Xbit_r21_c46 bl[46] br[46] wl[21] vdd gnd cell_6t
Xbit_r22_c46 bl[46] br[46] wl[22] vdd gnd cell_6t
Xbit_r23_c46 bl[46] br[46] wl[23] vdd gnd cell_6t
Xbit_r24_c46 bl[46] br[46] wl[24] vdd gnd cell_6t
Xbit_r25_c46 bl[46] br[46] wl[25] vdd gnd cell_6t
Xbit_r26_c46 bl[46] br[46] wl[26] vdd gnd cell_6t
Xbit_r27_c46 bl[46] br[46] wl[27] vdd gnd cell_6t
Xbit_r28_c46 bl[46] br[46] wl[28] vdd gnd cell_6t
Xbit_r29_c46 bl[46] br[46] wl[29] vdd gnd cell_6t
Xbit_r30_c46 bl[46] br[46] wl[30] vdd gnd cell_6t
Xbit_r31_c46 bl[46] br[46] wl[31] vdd gnd cell_6t
Xbit_r32_c46 bl[46] br[46] wl[32] vdd gnd cell_6t
Xbit_r33_c46 bl[46] br[46] wl[33] vdd gnd cell_6t
Xbit_r34_c46 bl[46] br[46] wl[34] vdd gnd cell_6t
Xbit_r35_c46 bl[46] br[46] wl[35] vdd gnd cell_6t
Xbit_r36_c46 bl[46] br[46] wl[36] vdd gnd cell_6t
Xbit_r37_c46 bl[46] br[46] wl[37] vdd gnd cell_6t
Xbit_r38_c46 bl[46] br[46] wl[38] vdd gnd cell_6t
Xbit_r39_c46 bl[46] br[46] wl[39] vdd gnd cell_6t
Xbit_r40_c46 bl[46] br[46] wl[40] vdd gnd cell_6t
Xbit_r41_c46 bl[46] br[46] wl[41] vdd gnd cell_6t
Xbit_r42_c46 bl[46] br[46] wl[42] vdd gnd cell_6t
Xbit_r43_c46 bl[46] br[46] wl[43] vdd gnd cell_6t
Xbit_r44_c46 bl[46] br[46] wl[44] vdd gnd cell_6t
Xbit_r45_c46 bl[46] br[46] wl[45] vdd gnd cell_6t
Xbit_r46_c46 bl[46] br[46] wl[46] vdd gnd cell_6t
Xbit_r47_c46 bl[46] br[46] wl[47] vdd gnd cell_6t
Xbit_r48_c46 bl[46] br[46] wl[48] vdd gnd cell_6t
Xbit_r49_c46 bl[46] br[46] wl[49] vdd gnd cell_6t
Xbit_r50_c46 bl[46] br[46] wl[50] vdd gnd cell_6t
Xbit_r51_c46 bl[46] br[46] wl[51] vdd gnd cell_6t
Xbit_r52_c46 bl[46] br[46] wl[52] vdd gnd cell_6t
Xbit_r53_c46 bl[46] br[46] wl[53] vdd gnd cell_6t
Xbit_r54_c46 bl[46] br[46] wl[54] vdd gnd cell_6t
Xbit_r55_c46 bl[46] br[46] wl[55] vdd gnd cell_6t
Xbit_r56_c46 bl[46] br[46] wl[56] vdd gnd cell_6t
Xbit_r57_c46 bl[46] br[46] wl[57] vdd gnd cell_6t
Xbit_r58_c46 bl[46] br[46] wl[58] vdd gnd cell_6t
Xbit_r59_c46 bl[46] br[46] wl[59] vdd gnd cell_6t
Xbit_r60_c46 bl[46] br[46] wl[60] vdd gnd cell_6t
Xbit_r61_c46 bl[46] br[46] wl[61] vdd gnd cell_6t
Xbit_r62_c46 bl[46] br[46] wl[62] vdd gnd cell_6t
Xbit_r63_c46 bl[46] br[46] wl[63] vdd gnd cell_6t
Xbit_r64_c46 bl[46] br[46] wl[64] vdd gnd cell_6t
Xbit_r65_c46 bl[46] br[46] wl[65] vdd gnd cell_6t
Xbit_r66_c46 bl[46] br[46] wl[66] vdd gnd cell_6t
Xbit_r67_c46 bl[46] br[46] wl[67] vdd gnd cell_6t
Xbit_r68_c46 bl[46] br[46] wl[68] vdd gnd cell_6t
Xbit_r69_c46 bl[46] br[46] wl[69] vdd gnd cell_6t
Xbit_r70_c46 bl[46] br[46] wl[70] vdd gnd cell_6t
Xbit_r71_c46 bl[46] br[46] wl[71] vdd gnd cell_6t
Xbit_r72_c46 bl[46] br[46] wl[72] vdd gnd cell_6t
Xbit_r73_c46 bl[46] br[46] wl[73] vdd gnd cell_6t
Xbit_r74_c46 bl[46] br[46] wl[74] vdd gnd cell_6t
Xbit_r75_c46 bl[46] br[46] wl[75] vdd gnd cell_6t
Xbit_r76_c46 bl[46] br[46] wl[76] vdd gnd cell_6t
Xbit_r77_c46 bl[46] br[46] wl[77] vdd gnd cell_6t
Xbit_r78_c46 bl[46] br[46] wl[78] vdd gnd cell_6t
Xbit_r79_c46 bl[46] br[46] wl[79] vdd gnd cell_6t
Xbit_r80_c46 bl[46] br[46] wl[80] vdd gnd cell_6t
Xbit_r81_c46 bl[46] br[46] wl[81] vdd gnd cell_6t
Xbit_r82_c46 bl[46] br[46] wl[82] vdd gnd cell_6t
Xbit_r83_c46 bl[46] br[46] wl[83] vdd gnd cell_6t
Xbit_r84_c46 bl[46] br[46] wl[84] vdd gnd cell_6t
Xbit_r85_c46 bl[46] br[46] wl[85] vdd gnd cell_6t
Xbit_r86_c46 bl[46] br[46] wl[86] vdd gnd cell_6t
Xbit_r87_c46 bl[46] br[46] wl[87] vdd gnd cell_6t
Xbit_r88_c46 bl[46] br[46] wl[88] vdd gnd cell_6t
Xbit_r89_c46 bl[46] br[46] wl[89] vdd gnd cell_6t
Xbit_r90_c46 bl[46] br[46] wl[90] vdd gnd cell_6t
Xbit_r91_c46 bl[46] br[46] wl[91] vdd gnd cell_6t
Xbit_r92_c46 bl[46] br[46] wl[92] vdd gnd cell_6t
Xbit_r93_c46 bl[46] br[46] wl[93] vdd gnd cell_6t
Xbit_r94_c46 bl[46] br[46] wl[94] vdd gnd cell_6t
Xbit_r95_c46 bl[46] br[46] wl[95] vdd gnd cell_6t
Xbit_r96_c46 bl[46] br[46] wl[96] vdd gnd cell_6t
Xbit_r97_c46 bl[46] br[46] wl[97] vdd gnd cell_6t
Xbit_r98_c46 bl[46] br[46] wl[98] vdd gnd cell_6t
Xbit_r99_c46 bl[46] br[46] wl[99] vdd gnd cell_6t
Xbit_r100_c46 bl[46] br[46] wl[100] vdd gnd cell_6t
Xbit_r101_c46 bl[46] br[46] wl[101] vdd gnd cell_6t
Xbit_r102_c46 bl[46] br[46] wl[102] vdd gnd cell_6t
Xbit_r103_c46 bl[46] br[46] wl[103] vdd gnd cell_6t
Xbit_r104_c46 bl[46] br[46] wl[104] vdd gnd cell_6t
Xbit_r105_c46 bl[46] br[46] wl[105] vdd gnd cell_6t
Xbit_r106_c46 bl[46] br[46] wl[106] vdd gnd cell_6t
Xbit_r107_c46 bl[46] br[46] wl[107] vdd gnd cell_6t
Xbit_r108_c46 bl[46] br[46] wl[108] vdd gnd cell_6t
Xbit_r109_c46 bl[46] br[46] wl[109] vdd gnd cell_6t
Xbit_r110_c46 bl[46] br[46] wl[110] vdd gnd cell_6t
Xbit_r111_c46 bl[46] br[46] wl[111] vdd gnd cell_6t
Xbit_r112_c46 bl[46] br[46] wl[112] vdd gnd cell_6t
Xbit_r113_c46 bl[46] br[46] wl[113] vdd gnd cell_6t
Xbit_r114_c46 bl[46] br[46] wl[114] vdd gnd cell_6t
Xbit_r115_c46 bl[46] br[46] wl[115] vdd gnd cell_6t
Xbit_r116_c46 bl[46] br[46] wl[116] vdd gnd cell_6t
Xbit_r117_c46 bl[46] br[46] wl[117] vdd gnd cell_6t
Xbit_r118_c46 bl[46] br[46] wl[118] vdd gnd cell_6t
Xbit_r119_c46 bl[46] br[46] wl[119] vdd gnd cell_6t
Xbit_r120_c46 bl[46] br[46] wl[120] vdd gnd cell_6t
Xbit_r121_c46 bl[46] br[46] wl[121] vdd gnd cell_6t
Xbit_r122_c46 bl[46] br[46] wl[122] vdd gnd cell_6t
Xbit_r123_c46 bl[46] br[46] wl[123] vdd gnd cell_6t
Xbit_r124_c46 bl[46] br[46] wl[124] vdd gnd cell_6t
Xbit_r125_c46 bl[46] br[46] wl[125] vdd gnd cell_6t
Xbit_r126_c46 bl[46] br[46] wl[126] vdd gnd cell_6t
Xbit_r127_c46 bl[46] br[46] wl[127] vdd gnd cell_6t
Xbit_r128_c46 bl[46] br[46] wl[128] vdd gnd cell_6t
Xbit_r129_c46 bl[46] br[46] wl[129] vdd gnd cell_6t
Xbit_r130_c46 bl[46] br[46] wl[130] vdd gnd cell_6t
Xbit_r131_c46 bl[46] br[46] wl[131] vdd gnd cell_6t
Xbit_r132_c46 bl[46] br[46] wl[132] vdd gnd cell_6t
Xbit_r133_c46 bl[46] br[46] wl[133] vdd gnd cell_6t
Xbit_r134_c46 bl[46] br[46] wl[134] vdd gnd cell_6t
Xbit_r135_c46 bl[46] br[46] wl[135] vdd gnd cell_6t
Xbit_r136_c46 bl[46] br[46] wl[136] vdd gnd cell_6t
Xbit_r137_c46 bl[46] br[46] wl[137] vdd gnd cell_6t
Xbit_r138_c46 bl[46] br[46] wl[138] vdd gnd cell_6t
Xbit_r139_c46 bl[46] br[46] wl[139] vdd gnd cell_6t
Xbit_r140_c46 bl[46] br[46] wl[140] vdd gnd cell_6t
Xbit_r141_c46 bl[46] br[46] wl[141] vdd gnd cell_6t
Xbit_r142_c46 bl[46] br[46] wl[142] vdd gnd cell_6t
Xbit_r143_c46 bl[46] br[46] wl[143] vdd gnd cell_6t
Xbit_r144_c46 bl[46] br[46] wl[144] vdd gnd cell_6t
Xbit_r145_c46 bl[46] br[46] wl[145] vdd gnd cell_6t
Xbit_r146_c46 bl[46] br[46] wl[146] vdd gnd cell_6t
Xbit_r147_c46 bl[46] br[46] wl[147] vdd gnd cell_6t
Xbit_r148_c46 bl[46] br[46] wl[148] vdd gnd cell_6t
Xbit_r149_c46 bl[46] br[46] wl[149] vdd gnd cell_6t
Xbit_r150_c46 bl[46] br[46] wl[150] vdd gnd cell_6t
Xbit_r151_c46 bl[46] br[46] wl[151] vdd gnd cell_6t
Xbit_r152_c46 bl[46] br[46] wl[152] vdd gnd cell_6t
Xbit_r153_c46 bl[46] br[46] wl[153] vdd gnd cell_6t
Xbit_r154_c46 bl[46] br[46] wl[154] vdd gnd cell_6t
Xbit_r155_c46 bl[46] br[46] wl[155] vdd gnd cell_6t
Xbit_r156_c46 bl[46] br[46] wl[156] vdd gnd cell_6t
Xbit_r157_c46 bl[46] br[46] wl[157] vdd gnd cell_6t
Xbit_r158_c46 bl[46] br[46] wl[158] vdd gnd cell_6t
Xbit_r159_c46 bl[46] br[46] wl[159] vdd gnd cell_6t
Xbit_r160_c46 bl[46] br[46] wl[160] vdd gnd cell_6t
Xbit_r161_c46 bl[46] br[46] wl[161] vdd gnd cell_6t
Xbit_r162_c46 bl[46] br[46] wl[162] vdd gnd cell_6t
Xbit_r163_c46 bl[46] br[46] wl[163] vdd gnd cell_6t
Xbit_r164_c46 bl[46] br[46] wl[164] vdd gnd cell_6t
Xbit_r165_c46 bl[46] br[46] wl[165] vdd gnd cell_6t
Xbit_r166_c46 bl[46] br[46] wl[166] vdd gnd cell_6t
Xbit_r167_c46 bl[46] br[46] wl[167] vdd gnd cell_6t
Xbit_r168_c46 bl[46] br[46] wl[168] vdd gnd cell_6t
Xbit_r169_c46 bl[46] br[46] wl[169] vdd gnd cell_6t
Xbit_r170_c46 bl[46] br[46] wl[170] vdd gnd cell_6t
Xbit_r171_c46 bl[46] br[46] wl[171] vdd gnd cell_6t
Xbit_r172_c46 bl[46] br[46] wl[172] vdd gnd cell_6t
Xbit_r173_c46 bl[46] br[46] wl[173] vdd gnd cell_6t
Xbit_r174_c46 bl[46] br[46] wl[174] vdd gnd cell_6t
Xbit_r175_c46 bl[46] br[46] wl[175] vdd gnd cell_6t
Xbit_r176_c46 bl[46] br[46] wl[176] vdd gnd cell_6t
Xbit_r177_c46 bl[46] br[46] wl[177] vdd gnd cell_6t
Xbit_r178_c46 bl[46] br[46] wl[178] vdd gnd cell_6t
Xbit_r179_c46 bl[46] br[46] wl[179] vdd gnd cell_6t
Xbit_r180_c46 bl[46] br[46] wl[180] vdd gnd cell_6t
Xbit_r181_c46 bl[46] br[46] wl[181] vdd gnd cell_6t
Xbit_r182_c46 bl[46] br[46] wl[182] vdd gnd cell_6t
Xbit_r183_c46 bl[46] br[46] wl[183] vdd gnd cell_6t
Xbit_r184_c46 bl[46] br[46] wl[184] vdd gnd cell_6t
Xbit_r185_c46 bl[46] br[46] wl[185] vdd gnd cell_6t
Xbit_r186_c46 bl[46] br[46] wl[186] vdd gnd cell_6t
Xbit_r187_c46 bl[46] br[46] wl[187] vdd gnd cell_6t
Xbit_r188_c46 bl[46] br[46] wl[188] vdd gnd cell_6t
Xbit_r189_c46 bl[46] br[46] wl[189] vdd gnd cell_6t
Xbit_r190_c46 bl[46] br[46] wl[190] vdd gnd cell_6t
Xbit_r191_c46 bl[46] br[46] wl[191] vdd gnd cell_6t
Xbit_r192_c46 bl[46] br[46] wl[192] vdd gnd cell_6t
Xbit_r193_c46 bl[46] br[46] wl[193] vdd gnd cell_6t
Xbit_r194_c46 bl[46] br[46] wl[194] vdd gnd cell_6t
Xbit_r195_c46 bl[46] br[46] wl[195] vdd gnd cell_6t
Xbit_r196_c46 bl[46] br[46] wl[196] vdd gnd cell_6t
Xbit_r197_c46 bl[46] br[46] wl[197] vdd gnd cell_6t
Xbit_r198_c46 bl[46] br[46] wl[198] vdd gnd cell_6t
Xbit_r199_c46 bl[46] br[46] wl[199] vdd gnd cell_6t
Xbit_r200_c46 bl[46] br[46] wl[200] vdd gnd cell_6t
Xbit_r201_c46 bl[46] br[46] wl[201] vdd gnd cell_6t
Xbit_r202_c46 bl[46] br[46] wl[202] vdd gnd cell_6t
Xbit_r203_c46 bl[46] br[46] wl[203] vdd gnd cell_6t
Xbit_r204_c46 bl[46] br[46] wl[204] vdd gnd cell_6t
Xbit_r205_c46 bl[46] br[46] wl[205] vdd gnd cell_6t
Xbit_r206_c46 bl[46] br[46] wl[206] vdd gnd cell_6t
Xbit_r207_c46 bl[46] br[46] wl[207] vdd gnd cell_6t
Xbit_r208_c46 bl[46] br[46] wl[208] vdd gnd cell_6t
Xbit_r209_c46 bl[46] br[46] wl[209] vdd gnd cell_6t
Xbit_r210_c46 bl[46] br[46] wl[210] vdd gnd cell_6t
Xbit_r211_c46 bl[46] br[46] wl[211] vdd gnd cell_6t
Xbit_r212_c46 bl[46] br[46] wl[212] vdd gnd cell_6t
Xbit_r213_c46 bl[46] br[46] wl[213] vdd gnd cell_6t
Xbit_r214_c46 bl[46] br[46] wl[214] vdd gnd cell_6t
Xbit_r215_c46 bl[46] br[46] wl[215] vdd gnd cell_6t
Xbit_r216_c46 bl[46] br[46] wl[216] vdd gnd cell_6t
Xbit_r217_c46 bl[46] br[46] wl[217] vdd gnd cell_6t
Xbit_r218_c46 bl[46] br[46] wl[218] vdd gnd cell_6t
Xbit_r219_c46 bl[46] br[46] wl[219] vdd gnd cell_6t
Xbit_r220_c46 bl[46] br[46] wl[220] vdd gnd cell_6t
Xbit_r221_c46 bl[46] br[46] wl[221] vdd gnd cell_6t
Xbit_r222_c46 bl[46] br[46] wl[222] vdd gnd cell_6t
Xbit_r223_c46 bl[46] br[46] wl[223] vdd gnd cell_6t
Xbit_r224_c46 bl[46] br[46] wl[224] vdd gnd cell_6t
Xbit_r225_c46 bl[46] br[46] wl[225] vdd gnd cell_6t
Xbit_r226_c46 bl[46] br[46] wl[226] vdd gnd cell_6t
Xbit_r227_c46 bl[46] br[46] wl[227] vdd gnd cell_6t
Xbit_r228_c46 bl[46] br[46] wl[228] vdd gnd cell_6t
Xbit_r229_c46 bl[46] br[46] wl[229] vdd gnd cell_6t
Xbit_r230_c46 bl[46] br[46] wl[230] vdd gnd cell_6t
Xbit_r231_c46 bl[46] br[46] wl[231] vdd gnd cell_6t
Xbit_r232_c46 bl[46] br[46] wl[232] vdd gnd cell_6t
Xbit_r233_c46 bl[46] br[46] wl[233] vdd gnd cell_6t
Xbit_r234_c46 bl[46] br[46] wl[234] vdd gnd cell_6t
Xbit_r235_c46 bl[46] br[46] wl[235] vdd gnd cell_6t
Xbit_r236_c46 bl[46] br[46] wl[236] vdd gnd cell_6t
Xbit_r237_c46 bl[46] br[46] wl[237] vdd gnd cell_6t
Xbit_r238_c46 bl[46] br[46] wl[238] vdd gnd cell_6t
Xbit_r239_c46 bl[46] br[46] wl[239] vdd gnd cell_6t
Xbit_r240_c46 bl[46] br[46] wl[240] vdd gnd cell_6t
Xbit_r241_c46 bl[46] br[46] wl[241] vdd gnd cell_6t
Xbit_r242_c46 bl[46] br[46] wl[242] vdd gnd cell_6t
Xbit_r243_c46 bl[46] br[46] wl[243] vdd gnd cell_6t
Xbit_r244_c46 bl[46] br[46] wl[244] vdd gnd cell_6t
Xbit_r245_c46 bl[46] br[46] wl[245] vdd gnd cell_6t
Xbit_r246_c46 bl[46] br[46] wl[246] vdd gnd cell_6t
Xbit_r247_c46 bl[46] br[46] wl[247] vdd gnd cell_6t
Xbit_r248_c46 bl[46] br[46] wl[248] vdd gnd cell_6t
Xbit_r249_c46 bl[46] br[46] wl[249] vdd gnd cell_6t
Xbit_r250_c46 bl[46] br[46] wl[250] vdd gnd cell_6t
Xbit_r251_c46 bl[46] br[46] wl[251] vdd gnd cell_6t
Xbit_r252_c46 bl[46] br[46] wl[252] vdd gnd cell_6t
Xbit_r253_c46 bl[46] br[46] wl[253] vdd gnd cell_6t
Xbit_r254_c46 bl[46] br[46] wl[254] vdd gnd cell_6t
Xbit_r255_c46 bl[46] br[46] wl[255] vdd gnd cell_6t
Xbit_r256_c46 bl[46] br[46] wl[256] vdd gnd cell_6t
Xbit_r257_c46 bl[46] br[46] wl[257] vdd gnd cell_6t
Xbit_r258_c46 bl[46] br[46] wl[258] vdd gnd cell_6t
Xbit_r259_c46 bl[46] br[46] wl[259] vdd gnd cell_6t
Xbit_r260_c46 bl[46] br[46] wl[260] vdd gnd cell_6t
Xbit_r261_c46 bl[46] br[46] wl[261] vdd gnd cell_6t
Xbit_r262_c46 bl[46] br[46] wl[262] vdd gnd cell_6t
Xbit_r263_c46 bl[46] br[46] wl[263] vdd gnd cell_6t
Xbit_r264_c46 bl[46] br[46] wl[264] vdd gnd cell_6t
Xbit_r265_c46 bl[46] br[46] wl[265] vdd gnd cell_6t
Xbit_r266_c46 bl[46] br[46] wl[266] vdd gnd cell_6t
Xbit_r267_c46 bl[46] br[46] wl[267] vdd gnd cell_6t
Xbit_r268_c46 bl[46] br[46] wl[268] vdd gnd cell_6t
Xbit_r269_c46 bl[46] br[46] wl[269] vdd gnd cell_6t
Xbit_r270_c46 bl[46] br[46] wl[270] vdd gnd cell_6t
Xbit_r271_c46 bl[46] br[46] wl[271] vdd gnd cell_6t
Xbit_r272_c46 bl[46] br[46] wl[272] vdd gnd cell_6t
Xbit_r273_c46 bl[46] br[46] wl[273] vdd gnd cell_6t
Xbit_r274_c46 bl[46] br[46] wl[274] vdd gnd cell_6t
Xbit_r275_c46 bl[46] br[46] wl[275] vdd gnd cell_6t
Xbit_r276_c46 bl[46] br[46] wl[276] vdd gnd cell_6t
Xbit_r277_c46 bl[46] br[46] wl[277] vdd gnd cell_6t
Xbit_r278_c46 bl[46] br[46] wl[278] vdd gnd cell_6t
Xbit_r279_c46 bl[46] br[46] wl[279] vdd gnd cell_6t
Xbit_r280_c46 bl[46] br[46] wl[280] vdd gnd cell_6t
Xbit_r281_c46 bl[46] br[46] wl[281] vdd gnd cell_6t
Xbit_r282_c46 bl[46] br[46] wl[282] vdd gnd cell_6t
Xbit_r283_c46 bl[46] br[46] wl[283] vdd gnd cell_6t
Xbit_r284_c46 bl[46] br[46] wl[284] vdd gnd cell_6t
Xbit_r285_c46 bl[46] br[46] wl[285] vdd gnd cell_6t
Xbit_r286_c46 bl[46] br[46] wl[286] vdd gnd cell_6t
Xbit_r287_c46 bl[46] br[46] wl[287] vdd gnd cell_6t
Xbit_r288_c46 bl[46] br[46] wl[288] vdd gnd cell_6t
Xbit_r289_c46 bl[46] br[46] wl[289] vdd gnd cell_6t
Xbit_r290_c46 bl[46] br[46] wl[290] vdd gnd cell_6t
Xbit_r291_c46 bl[46] br[46] wl[291] vdd gnd cell_6t
Xbit_r292_c46 bl[46] br[46] wl[292] vdd gnd cell_6t
Xbit_r293_c46 bl[46] br[46] wl[293] vdd gnd cell_6t
Xbit_r294_c46 bl[46] br[46] wl[294] vdd gnd cell_6t
Xbit_r295_c46 bl[46] br[46] wl[295] vdd gnd cell_6t
Xbit_r296_c46 bl[46] br[46] wl[296] vdd gnd cell_6t
Xbit_r297_c46 bl[46] br[46] wl[297] vdd gnd cell_6t
Xbit_r298_c46 bl[46] br[46] wl[298] vdd gnd cell_6t
Xbit_r299_c46 bl[46] br[46] wl[299] vdd gnd cell_6t
Xbit_r300_c46 bl[46] br[46] wl[300] vdd gnd cell_6t
Xbit_r301_c46 bl[46] br[46] wl[301] vdd gnd cell_6t
Xbit_r302_c46 bl[46] br[46] wl[302] vdd gnd cell_6t
Xbit_r303_c46 bl[46] br[46] wl[303] vdd gnd cell_6t
Xbit_r304_c46 bl[46] br[46] wl[304] vdd gnd cell_6t
Xbit_r305_c46 bl[46] br[46] wl[305] vdd gnd cell_6t
Xbit_r306_c46 bl[46] br[46] wl[306] vdd gnd cell_6t
Xbit_r307_c46 bl[46] br[46] wl[307] vdd gnd cell_6t
Xbit_r308_c46 bl[46] br[46] wl[308] vdd gnd cell_6t
Xbit_r309_c46 bl[46] br[46] wl[309] vdd gnd cell_6t
Xbit_r310_c46 bl[46] br[46] wl[310] vdd gnd cell_6t
Xbit_r311_c46 bl[46] br[46] wl[311] vdd gnd cell_6t
Xbit_r312_c46 bl[46] br[46] wl[312] vdd gnd cell_6t
Xbit_r313_c46 bl[46] br[46] wl[313] vdd gnd cell_6t
Xbit_r314_c46 bl[46] br[46] wl[314] vdd gnd cell_6t
Xbit_r315_c46 bl[46] br[46] wl[315] vdd gnd cell_6t
Xbit_r316_c46 bl[46] br[46] wl[316] vdd gnd cell_6t
Xbit_r317_c46 bl[46] br[46] wl[317] vdd gnd cell_6t
Xbit_r318_c46 bl[46] br[46] wl[318] vdd gnd cell_6t
Xbit_r319_c46 bl[46] br[46] wl[319] vdd gnd cell_6t
Xbit_r320_c46 bl[46] br[46] wl[320] vdd gnd cell_6t
Xbit_r321_c46 bl[46] br[46] wl[321] vdd gnd cell_6t
Xbit_r322_c46 bl[46] br[46] wl[322] vdd gnd cell_6t
Xbit_r323_c46 bl[46] br[46] wl[323] vdd gnd cell_6t
Xbit_r324_c46 bl[46] br[46] wl[324] vdd gnd cell_6t
Xbit_r325_c46 bl[46] br[46] wl[325] vdd gnd cell_6t
Xbit_r326_c46 bl[46] br[46] wl[326] vdd gnd cell_6t
Xbit_r327_c46 bl[46] br[46] wl[327] vdd gnd cell_6t
Xbit_r328_c46 bl[46] br[46] wl[328] vdd gnd cell_6t
Xbit_r329_c46 bl[46] br[46] wl[329] vdd gnd cell_6t
Xbit_r330_c46 bl[46] br[46] wl[330] vdd gnd cell_6t
Xbit_r331_c46 bl[46] br[46] wl[331] vdd gnd cell_6t
Xbit_r332_c46 bl[46] br[46] wl[332] vdd gnd cell_6t
Xbit_r333_c46 bl[46] br[46] wl[333] vdd gnd cell_6t
Xbit_r334_c46 bl[46] br[46] wl[334] vdd gnd cell_6t
Xbit_r335_c46 bl[46] br[46] wl[335] vdd gnd cell_6t
Xbit_r336_c46 bl[46] br[46] wl[336] vdd gnd cell_6t
Xbit_r337_c46 bl[46] br[46] wl[337] vdd gnd cell_6t
Xbit_r338_c46 bl[46] br[46] wl[338] vdd gnd cell_6t
Xbit_r339_c46 bl[46] br[46] wl[339] vdd gnd cell_6t
Xbit_r340_c46 bl[46] br[46] wl[340] vdd gnd cell_6t
Xbit_r341_c46 bl[46] br[46] wl[341] vdd gnd cell_6t
Xbit_r342_c46 bl[46] br[46] wl[342] vdd gnd cell_6t
Xbit_r343_c46 bl[46] br[46] wl[343] vdd gnd cell_6t
Xbit_r344_c46 bl[46] br[46] wl[344] vdd gnd cell_6t
Xbit_r345_c46 bl[46] br[46] wl[345] vdd gnd cell_6t
Xbit_r346_c46 bl[46] br[46] wl[346] vdd gnd cell_6t
Xbit_r347_c46 bl[46] br[46] wl[347] vdd gnd cell_6t
Xbit_r348_c46 bl[46] br[46] wl[348] vdd gnd cell_6t
Xbit_r349_c46 bl[46] br[46] wl[349] vdd gnd cell_6t
Xbit_r350_c46 bl[46] br[46] wl[350] vdd gnd cell_6t
Xbit_r351_c46 bl[46] br[46] wl[351] vdd gnd cell_6t
Xbit_r352_c46 bl[46] br[46] wl[352] vdd gnd cell_6t
Xbit_r353_c46 bl[46] br[46] wl[353] vdd gnd cell_6t
Xbit_r354_c46 bl[46] br[46] wl[354] vdd gnd cell_6t
Xbit_r355_c46 bl[46] br[46] wl[355] vdd gnd cell_6t
Xbit_r356_c46 bl[46] br[46] wl[356] vdd gnd cell_6t
Xbit_r357_c46 bl[46] br[46] wl[357] vdd gnd cell_6t
Xbit_r358_c46 bl[46] br[46] wl[358] vdd gnd cell_6t
Xbit_r359_c46 bl[46] br[46] wl[359] vdd gnd cell_6t
Xbit_r360_c46 bl[46] br[46] wl[360] vdd gnd cell_6t
Xbit_r361_c46 bl[46] br[46] wl[361] vdd gnd cell_6t
Xbit_r362_c46 bl[46] br[46] wl[362] vdd gnd cell_6t
Xbit_r363_c46 bl[46] br[46] wl[363] vdd gnd cell_6t
Xbit_r364_c46 bl[46] br[46] wl[364] vdd gnd cell_6t
Xbit_r365_c46 bl[46] br[46] wl[365] vdd gnd cell_6t
Xbit_r366_c46 bl[46] br[46] wl[366] vdd gnd cell_6t
Xbit_r367_c46 bl[46] br[46] wl[367] vdd gnd cell_6t
Xbit_r368_c46 bl[46] br[46] wl[368] vdd gnd cell_6t
Xbit_r369_c46 bl[46] br[46] wl[369] vdd gnd cell_6t
Xbit_r370_c46 bl[46] br[46] wl[370] vdd gnd cell_6t
Xbit_r371_c46 bl[46] br[46] wl[371] vdd gnd cell_6t
Xbit_r372_c46 bl[46] br[46] wl[372] vdd gnd cell_6t
Xbit_r373_c46 bl[46] br[46] wl[373] vdd gnd cell_6t
Xbit_r374_c46 bl[46] br[46] wl[374] vdd gnd cell_6t
Xbit_r375_c46 bl[46] br[46] wl[375] vdd gnd cell_6t
Xbit_r376_c46 bl[46] br[46] wl[376] vdd gnd cell_6t
Xbit_r377_c46 bl[46] br[46] wl[377] vdd gnd cell_6t
Xbit_r378_c46 bl[46] br[46] wl[378] vdd gnd cell_6t
Xbit_r379_c46 bl[46] br[46] wl[379] vdd gnd cell_6t
Xbit_r380_c46 bl[46] br[46] wl[380] vdd gnd cell_6t
Xbit_r381_c46 bl[46] br[46] wl[381] vdd gnd cell_6t
Xbit_r382_c46 bl[46] br[46] wl[382] vdd gnd cell_6t
Xbit_r383_c46 bl[46] br[46] wl[383] vdd gnd cell_6t
Xbit_r384_c46 bl[46] br[46] wl[384] vdd gnd cell_6t
Xbit_r385_c46 bl[46] br[46] wl[385] vdd gnd cell_6t
Xbit_r386_c46 bl[46] br[46] wl[386] vdd gnd cell_6t
Xbit_r387_c46 bl[46] br[46] wl[387] vdd gnd cell_6t
Xbit_r388_c46 bl[46] br[46] wl[388] vdd gnd cell_6t
Xbit_r389_c46 bl[46] br[46] wl[389] vdd gnd cell_6t
Xbit_r390_c46 bl[46] br[46] wl[390] vdd gnd cell_6t
Xbit_r391_c46 bl[46] br[46] wl[391] vdd gnd cell_6t
Xbit_r392_c46 bl[46] br[46] wl[392] vdd gnd cell_6t
Xbit_r393_c46 bl[46] br[46] wl[393] vdd gnd cell_6t
Xbit_r394_c46 bl[46] br[46] wl[394] vdd gnd cell_6t
Xbit_r395_c46 bl[46] br[46] wl[395] vdd gnd cell_6t
Xbit_r396_c46 bl[46] br[46] wl[396] vdd gnd cell_6t
Xbit_r397_c46 bl[46] br[46] wl[397] vdd gnd cell_6t
Xbit_r398_c46 bl[46] br[46] wl[398] vdd gnd cell_6t
Xbit_r399_c46 bl[46] br[46] wl[399] vdd gnd cell_6t
Xbit_r400_c46 bl[46] br[46] wl[400] vdd gnd cell_6t
Xbit_r401_c46 bl[46] br[46] wl[401] vdd gnd cell_6t
Xbit_r402_c46 bl[46] br[46] wl[402] vdd gnd cell_6t
Xbit_r403_c46 bl[46] br[46] wl[403] vdd gnd cell_6t
Xbit_r404_c46 bl[46] br[46] wl[404] vdd gnd cell_6t
Xbit_r405_c46 bl[46] br[46] wl[405] vdd gnd cell_6t
Xbit_r406_c46 bl[46] br[46] wl[406] vdd gnd cell_6t
Xbit_r407_c46 bl[46] br[46] wl[407] vdd gnd cell_6t
Xbit_r408_c46 bl[46] br[46] wl[408] vdd gnd cell_6t
Xbit_r409_c46 bl[46] br[46] wl[409] vdd gnd cell_6t
Xbit_r410_c46 bl[46] br[46] wl[410] vdd gnd cell_6t
Xbit_r411_c46 bl[46] br[46] wl[411] vdd gnd cell_6t
Xbit_r412_c46 bl[46] br[46] wl[412] vdd gnd cell_6t
Xbit_r413_c46 bl[46] br[46] wl[413] vdd gnd cell_6t
Xbit_r414_c46 bl[46] br[46] wl[414] vdd gnd cell_6t
Xbit_r415_c46 bl[46] br[46] wl[415] vdd gnd cell_6t
Xbit_r416_c46 bl[46] br[46] wl[416] vdd gnd cell_6t
Xbit_r417_c46 bl[46] br[46] wl[417] vdd gnd cell_6t
Xbit_r418_c46 bl[46] br[46] wl[418] vdd gnd cell_6t
Xbit_r419_c46 bl[46] br[46] wl[419] vdd gnd cell_6t
Xbit_r420_c46 bl[46] br[46] wl[420] vdd gnd cell_6t
Xbit_r421_c46 bl[46] br[46] wl[421] vdd gnd cell_6t
Xbit_r422_c46 bl[46] br[46] wl[422] vdd gnd cell_6t
Xbit_r423_c46 bl[46] br[46] wl[423] vdd gnd cell_6t
Xbit_r424_c46 bl[46] br[46] wl[424] vdd gnd cell_6t
Xbit_r425_c46 bl[46] br[46] wl[425] vdd gnd cell_6t
Xbit_r426_c46 bl[46] br[46] wl[426] vdd gnd cell_6t
Xbit_r427_c46 bl[46] br[46] wl[427] vdd gnd cell_6t
Xbit_r428_c46 bl[46] br[46] wl[428] vdd gnd cell_6t
Xbit_r429_c46 bl[46] br[46] wl[429] vdd gnd cell_6t
Xbit_r430_c46 bl[46] br[46] wl[430] vdd gnd cell_6t
Xbit_r431_c46 bl[46] br[46] wl[431] vdd gnd cell_6t
Xbit_r432_c46 bl[46] br[46] wl[432] vdd gnd cell_6t
Xbit_r433_c46 bl[46] br[46] wl[433] vdd gnd cell_6t
Xbit_r434_c46 bl[46] br[46] wl[434] vdd gnd cell_6t
Xbit_r435_c46 bl[46] br[46] wl[435] vdd gnd cell_6t
Xbit_r436_c46 bl[46] br[46] wl[436] vdd gnd cell_6t
Xbit_r437_c46 bl[46] br[46] wl[437] vdd gnd cell_6t
Xbit_r438_c46 bl[46] br[46] wl[438] vdd gnd cell_6t
Xbit_r439_c46 bl[46] br[46] wl[439] vdd gnd cell_6t
Xbit_r440_c46 bl[46] br[46] wl[440] vdd gnd cell_6t
Xbit_r441_c46 bl[46] br[46] wl[441] vdd gnd cell_6t
Xbit_r442_c46 bl[46] br[46] wl[442] vdd gnd cell_6t
Xbit_r443_c46 bl[46] br[46] wl[443] vdd gnd cell_6t
Xbit_r444_c46 bl[46] br[46] wl[444] vdd gnd cell_6t
Xbit_r445_c46 bl[46] br[46] wl[445] vdd gnd cell_6t
Xbit_r446_c46 bl[46] br[46] wl[446] vdd gnd cell_6t
Xbit_r447_c46 bl[46] br[46] wl[447] vdd gnd cell_6t
Xbit_r448_c46 bl[46] br[46] wl[448] vdd gnd cell_6t
Xbit_r449_c46 bl[46] br[46] wl[449] vdd gnd cell_6t
Xbit_r450_c46 bl[46] br[46] wl[450] vdd gnd cell_6t
Xbit_r451_c46 bl[46] br[46] wl[451] vdd gnd cell_6t
Xbit_r452_c46 bl[46] br[46] wl[452] vdd gnd cell_6t
Xbit_r453_c46 bl[46] br[46] wl[453] vdd gnd cell_6t
Xbit_r454_c46 bl[46] br[46] wl[454] vdd gnd cell_6t
Xbit_r455_c46 bl[46] br[46] wl[455] vdd gnd cell_6t
Xbit_r456_c46 bl[46] br[46] wl[456] vdd gnd cell_6t
Xbit_r457_c46 bl[46] br[46] wl[457] vdd gnd cell_6t
Xbit_r458_c46 bl[46] br[46] wl[458] vdd gnd cell_6t
Xbit_r459_c46 bl[46] br[46] wl[459] vdd gnd cell_6t
Xbit_r460_c46 bl[46] br[46] wl[460] vdd gnd cell_6t
Xbit_r461_c46 bl[46] br[46] wl[461] vdd gnd cell_6t
Xbit_r462_c46 bl[46] br[46] wl[462] vdd gnd cell_6t
Xbit_r463_c46 bl[46] br[46] wl[463] vdd gnd cell_6t
Xbit_r464_c46 bl[46] br[46] wl[464] vdd gnd cell_6t
Xbit_r465_c46 bl[46] br[46] wl[465] vdd gnd cell_6t
Xbit_r466_c46 bl[46] br[46] wl[466] vdd gnd cell_6t
Xbit_r467_c46 bl[46] br[46] wl[467] vdd gnd cell_6t
Xbit_r468_c46 bl[46] br[46] wl[468] vdd gnd cell_6t
Xbit_r469_c46 bl[46] br[46] wl[469] vdd gnd cell_6t
Xbit_r470_c46 bl[46] br[46] wl[470] vdd gnd cell_6t
Xbit_r471_c46 bl[46] br[46] wl[471] vdd gnd cell_6t
Xbit_r472_c46 bl[46] br[46] wl[472] vdd gnd cell_6t
Xbit_r473_c46 bl[46] br[46] wl[473] vdd gnd cell_6t
Xbit_r474_c46 bl[46] br[46] wl[474] vdd gnd cell_6t
Xbit_r475_c46 bl[46] br[46] wl[475] vdd gnd cell_6t
Xbit_r476_c46 bl[46] br[46] wl[476] vdd gnd cell_6t
Xbit_r477_c46 bl[46] br[46] wl[477] vdd gnd cell_6t
Xbit_r478_c46 bl[46] br[46] wl[478] vdd gnd cell_6t
Xbit_r479_c46 bl[46] br[46] wl[479] vdd gnd cell_6t
Xbit_r480_c46 bl[46] br[46] wl[480] vdd gnd cell_6t
Xbit_r481_c46 bl[46] br[46] wl[481] vdd gnd cell_6t
Xbit_r482_c46 bl[46] br[46] wl[482] vdd gnd cell_6t
Xbit_r483_c46 bl[46] br[46] wl[483] vdd gnd cell_6t
Xbit_r484_c46 bl[46] br[46] wl[484] vdd gnd cell_6t
Xbit_r485_c46 bl[46] br[46] wl[485] vdd gnd cell_6t
Xbit_r486_c46 bl[46] br[46] wl[486] vdd gnd cell_6t
Xbit_r487_c46 bl[46] br[46] wl[487] vdd gnd cell_6t
Xbit_r488_c46 bl[46] br[46] wl[488] vdd gnd cell_6t
Xbit_r489_c46 bl[46] br[46] wl[489] vdd gnd cell_6t
Xbit_r490_c46 bl[46] br[46] wl[490] vdd gnd cell_6t
Xbit_r491_c46 bl[46] br[46] wl[491] vdd gnd cell_6t
Xbit_r492_c46 bl[46] br[46] wl[492] vdd gnd cell_6t
Xbit_r493_c46 bl[46] br[46] wl[493] vdd gnd cell_6t
Xbit_r494_c46 bl[46] br[46] wl[494] vdd gnd cell_6t
Xbit_r495_c46 bl[46] br[46] wl[495] vdd gnd cell_6t
Xbit_r496_c46 bl[46] br[46] wl[496] vdd gnd cell_6t
Xbit_r497_c46 bl[46] br[46] wl[497] vdd gnd cell_6t
Xbit_r498_c46 bl[46] br[46] wl[498] vdd gnd cell_6t
Xbit_r499_c46 bl[46] br[46] wl[499] vdd gnd cell_6t
Xbit_r500_c46 bl[46] br[46] wl[500] vdd gnd cell_6t
Xbit_r501_c46 bl[46] br[46] wl[501] vdd gnd cell_6t
Xbit_r502_c46 bl[46] br[46] wl[502] vdd gnd cell_6t
Xbit_r503_c46 bl[46] br[46] wl[503] vdd gnd cell_6t
Xbit_r504_c46 bl[46] br[46] wl[504] vdd gnd cell_6t
Xbit_r505_c46 bl[46] br[46] wl[505] vdd gnd cell_6t
Xbit_r506_c46 bl[46] br[46] wl[506] vdd gnd cell_6t
Xbit_r507_c46 bl[46] br[46] wl[507] vdd gnd cell_6t
Xbit_r508_c46 bl[46] br[46] wl[508] vdd gnd cell_6t
Xbit_r509_c46 bl[46] br[46] wl[509] vdd gnd cell_6t
Xbit_r510_c46 bl[46] br[46] wl[510] vdd gnd cell_6t
Xbit_r511_c46 bl[46] br[46] wl[511] vdd gnd cell_6t
Xbit_r0_c47 bl[47] br[47] wl[0] vdd gnd cell_6t
Xbit_r1_c47 bl[47] br[47] wl[1] vdd gnd cell_6t
Xbit_r2_c47 bl[47] br[47] wl[2] vdd gnd cell_6t
Xbit_r3_c47 bl[47] br[47] wl[3] vdd gnd cell_6t
Xbit_r4_c47 bl[47] br[47] wl[4] vdd gnd cell_6t
Xbit_r5_c47 bl[47] br[47] wl[5] vdd gnd cell_6t
Xbit_r6_c47 bl[47] br[47] wl[6] vdd gnd cell_6t
Xbit_r7_c47 bl[47] br[47] wl[7] vdd gnd cell_6t
Xbit_r8_c47 bl[47] br[47] wl[8] vdd gnd cell_6t
Xbit_r9_c47 bl[47] br[47] wl[9] vdd gnd cell_6t
Xbit_r10_c47 bl[47] br[47] wl[10] vdd gnd cell_6t
Xbit_r11_c47 bl[47] br[47] wl[11] vdd gnd cell_6t
Xbit_r12_c47 bl[47] br[47] wl[12] vdd gnd cell_6t
Xbit_r13_c47 bl[47] br[47] wl[13] vdd gnd cell_6t
Xbit_r14_c47 bl[47] br[47] wl[14] vdd gnd cell_6t
Xbit_r15_c47 bl[47] br[47] wl[15] vdd gnd cell_6t
Xbit_r16_c47 bl[47] br[47] wl[16] vdd gnd cell_6t
Xbit_r17_c47 bl[47] br[47] wl[17] vdd gnd cell_6t
Xbit_r18_c47 bl[47] br[47] wl[18] vdd gnd cell_6t
Xbit_r19_c47 bl[47] br[47] wl[19] vdd gnd cell_6t
Xbit_r20_c47 bl[47] br[47] wl[20] vdd gnd cell_6t
Xbit_r21_c47 bl[47] br[47] wl[21] vdd gnd cell_6t
Xbit_r22_c47 bl[47] br[47] wl[22] vdd gnd cell_6t
Xbit_r23_c47 bl[47] br[47] wl[23] vdd gnd cell_6t
Xbit_r24_c47 bl[47] br[47] wl[24] vdd gnd cell_6t
Xbit_r25_c47 bl[47] br[47] wl[25] vdd gnd cell_6t
Xbit_r26_c47 bl[47] br[47] wl[26] vdd gnd cell_6t
Xbit_r27_c47 bl[47] br[47] wl[27] vdd gnd cell_6t
Xbit_r28_c47 bl[47] br[47] wl[28] vdd gnd cell_6t
Xbit_r29_c47 bl[47] br[47] wl[29] vdd gnd cell_6t
Xbit_r30_c47 bl[47] br[47] wl[30] vdd gnd cell_6t
Xbit_r31_c47 bl[47] br[47] wl[31] vdd gnd cell_6t
Xbit_r32_c47 bl[47] br[47] wl[32] vdd gnd cell_6t
Xbit_r33_c47 bl[47] br[47] wl[33] vdd gnd cell_6t
Xbit_r34_c47 bl[47] br[47] wl[34] vdd gnd cell_6t
Xbit_r35_c47 bl[47] br[47] wl[35] vdd gnd cell_6t
Xbit_r36_c47 bl[47] br[47] wl[36] vdd gnd cell_6t
Xbit_r37_c47 bl[47] br[47] wl[37] vdd gnd cell_6t
Xbit_r38_c47 bl[47] br[47] wl[38] vdd gnd cell_6t
Xbit_r39_c47 bl[47] br[47] wl[39] vdd gnd cell_6t
Xbit_r40_c47 bl[47] br[47] wl[40] vdd gnd cell_6t
Xbit_r41_c47 bl[47] br[47] wl[41] vdd gnd cell_6t
Xbit_r42_c47 bl[47] br[47] wl[42] vdd gnd cell_6t
Xbit_r43_c47 bl[47] br[47] wl[43] vdd gnd cell_6t
Xbit_r44_c47 bl[47] br[47] wl[44] vdd gnd cell_6t
Xbit_r45_c47 bl[47] br[47] wl[45] vdd gnd cell_6t
Xbit_r46_c47 bl[47] br[47] wl[46] vdd gnd cell_6t
Xbit_r47_c47 bl[47] br[47] wl[47] vdd gnd cell_6t
Xbit_r48_c47 bl[47] br[47] wl[48] vdd gnd cell_6t
Xbit_r49_c47 bl[47] br[47] wl[49] vdd gnd cell_6t
Xbit_r50_c47 bl[47] br[47] wl[50] vdd gnd cell_6t
Xbit_r51_c47 bl[47] br[47] wl[51] vdd gnd cell_6t
Xbit_r52_c47 bl[47] br[47] wl[52] vdd gnd cell_6t
Xbit_r53_c47 bl[47] br[47] wl[53] vdd gnd cell_6t
Xbit_r54_c47 bl[47] br[47] wl[54] vdd gnd cell_6t
Xbit_r55_c47 bl[47] br[47] wl[55] vdd gnd cell_6t
Xbit_r56_c47 bl[47] br[47] wl[56] vdd gnd cell_6t
Xbit_r57_c47 bl[47] br[47] wl[57] vdd gnd cell_6t
Xbit_r58_c47 bl[47] br[47] wl[58] vdd gnd cell_6t
Xbit_r59_c47 bl[47] br[47] wl[59] vdd gnd cell_6t
Xbit_r60_c47 bl[47] br[47] wl[60] vdd gnd cell_6t
Xbit_r61_c47 bl[47] br[47] wl[61] vdd gnd cell_6t
Xbit_r62_c47 bl[47] br[47] wl[62] vdd gnd cell_6t
Xbit_r63_c47 bl[47] br[47] wl[63] vdd gnd cell_6t
Xbit_r64_c47 bl[47] br[47] wl[64] vdd gnd cell_6t
Xbit_r65_c47 bl[47] br[47] wl[65] vdd gnd cell_6t
Xbit_r66_c47 bl[47] br[47] wl[66] vdd gnd cell_6t
Xbit_r67_c47 bl[47] br[47] wl[67] vdd gnd cell_6t
Xbit_r68_c47 bl[47] br[47] wl[68] vdd gnd cell_6t
Xbit_r69_c47 bl[47] br[47] wl[69] vdd gnd cell_6t
Xbit_r70_c47 bl[47] br[47] wl[70] vdd gnd cell_6t
Xbit_r71_c47 bl[47] br[47] wl[71] vdd gnd cell_6t
Xbit_r72_c47 bl[47] br[47] wl[72] vdd gnd cell_6t
Xbit_r73_c47 bl[47] br[47] wl[73] vdd gnd cell_6t
Xbit_r74_c47 bl[47] br[47] wl[74] vdd gnd cell_6t
Xbit_r75_c47 bl[47] br[47] wl[75] vdd gnd cell_6t
Xbit_r76_c47 bl[47] br[47] wl[76] vdd gnd cell_6t
Xbit_r77_c47 bl[47] br[47] wl[77] vdd gnd cell_6t
Xbit_r78_c47 bl[47] br[47] wl[78] vdd gnd cell_6t
Xbit_r79_c47 bl[47] br[47] wl[79] vdd gnd cell_6t
Xbit_r80_c47 bl[47] br[47] wl[80] vdd gnd cell_6t
Xbit_r81_c47 bl[47] br[47] wl[81] vdd gnd cell_6t
Xbit_r82_c47 bl[47] br[47] wl[82] vdd gnd cell_6t
Xbit_r83_c47 bl[47] br[47] wl[83] vdd gnd cell_6t
Xbit_r84_c47 bl[47] br[47] wl[84] vdd gnd cell_6t
Xbit_r85_c47 bl[47] br[47] wl[85] vdd gnd cell_6t
Xbit_r86_c47 bl[47] br[47] wl[86] vdd gnd cell_6t
Xbit_r87_c47 bl[47] br[47] wl[87] vdd gnd cell_6t
Xbit_r88_c47 bl[47] br[47] wl[88] vdd gnd cell_6t
Xbit_r89_c47 bl[47] br[47] wl[89] vdd gnd cell_6t
Xbit_r90_c47 bl[47] br[47] wl[90] vdd gnd cell_6t
Xbit_r91_c47 bl[47] br[47] wl[91] vdd gnd cell_6t
Xbit_r92_c47 bl[47] br[47] wl[92] vdd gnd cell_6t
Xbit_r93_c47 bl[47] br[47] wl[93] vdd gnd cell_6t
Xbit_r94_c47 bl[47] br[47] wl[94] vdd gnd cell_6t
Xbit_r95_c47 bl[47] br[47] wl[95] vdd gnd cell_6t
Xbit_r96_c47 bl[47] br[47] wl[96] vdd gnd cell_6t
Xbit_r97_c47 bl[47] br[47] wl[97] vdd gnd cell_6t
Xbit_r98_c47 bl[47] br[47] wl[98] vdd gnd cell_6t
Xbit_r99_c47 bl[47] br[47] wl[99] vdd gnd cell_6t
Xbit_r100_c47 bl[47] br[47] wl[100] vdd gnd cell_6t
Xbit_r101_c47 bl[47] br[47] wl[101] vdd gnd cell_6t
Xbit_r102_c47 bl[47] br[47] wl[102] vdd gnd cell_6t
Xbit_r103_c47 bl[47] br[47] wl[103] vdd gnd cell_6t
Xbit_r104_c47 bl[47] br[47] wl[104] vdd gnd cell_6t
Xbit_r105_c47 bl[47] br[47] wl[105] vdd gnd cell_6t
Xbit_r106_c47 bl[47] br[47] wl[106] vdd gnd cell_6t
Xbit_r107_c47 bl[47] br[47] wl[107] vdd gnd cell_6t
Xbit_r108_c47 bl[47] br[47] wl[108] vdd gnd cell_6t
Xbit_r109_c47 bl[47] br[47] wl[109] vdd gnd cell_6t
Xbit_r110_c47 bl[47] br[47] wl[110] vdd gnd cell_6t
Xbit_r111_c47 bl[47] br[47] wl[111] vdd gnd cell_6t
Xbit_r112_c47 bl[47] br[47] wl[112] vdd gnd cell_6t
Xbit_r113_c47 bl[47] br[47] wl[113] vdd gnd cell_6t
Xbit_r114_c47 bl[47] br[47] wl[114] vdd gnd cell_6t
Xbit_r115_c47 bl[47] br[47] wl[115] vdd gnd cell_6t
Xbit_r116_c47 bl[47] br[47] wl[116] vdd gnd cell_6t
Xbit_r117_c47 bl[47] br[47] wl[117] vdd gnd cell_6t
Xbit_r118_c47 bl[47] br[47] wl[118] vdd gnd cell_6t
Xbit_r119_c47 bl[47] br[47] wl[119] vdd gnd cell_6t
Xbit_r120_c47 bl[47] br[47] wl[120] vdd gnd cell_6t
Xbit_r121_c47 bl[47] br[47] wl[121] vdd gnd cell_6t
Xbit_r122_c47 bl[47] br[47] wl[122] vdd gnd cell_6t
Xbit_r123_c47 bl[47] br[47] wl[123] vdd gnd cell_6t
Xbit_r124_c47 bl[47] br[47] wl[124] vdd gnd cell_6t
Xbit_r125_c47 bl[47] br[47] wl[125] vdd gnd cell_6t
Xbit_r126_c47 bl[47] br[47] wl[126] vdd gnd cell_6t
Xbit_r127_c47 bl[47] br[47] wl[127] vdd gnd cell_6t
Xbit_r128_c47 bl[47] br[47] wl[128] vdd gnd cell_6t
Xbit_r129_c47 bl[47] br[47] wl[129] vdd gnd cell_6t
Xbit_r130_c47 bl[47] br[47] wl[130] vdd gnd cell_6t
Xbit_r131_c47 bl[47] br[47] wl[131] vdd gnd cell_6t
Xbit_r132_c47 bl[47] br[47] wl[132] vdd gnd cell_6t
Xbit_r133_c47 bl[47] br[47] wl[133] vdd gnd cell_6t
Xbit_r134_c47 bl[47] br[47] wl[134] vdd gnd cell_6t
Xbit_r135_c47 bl[47] br[47] wl[135] vdd gnd cell_6t
Xbit_r136_c47 bl[47] br[47] wl[136] vdd gnd cell_6t
Xbit_r137_c47 bl[47] br[47] wl[137] vdd gnd cell_6t
Xbit_r138_c47 bl[47] br[47] wl[138] vdd gnd cell_6t
Xbit_r139_c47 bl[47] br[47] wl[139] vdd gnd cell_6t
Xbit_r140_c47 bl[47] br[47] wl[140] vdd gnd cell_6t
Xbit_r141_c47 bl[47] br[47] wl[141] vdd gnd cell_6t
Xbit_r142_c47 bl[47] br[47] wl[142] vdd gnd cell_6t
Xbit_r143_c47 bl[47] br[47] wl[143] vdd gnd cell_6t
Xbit_r144_c47 bl[47] br[47] wl[144] vdd gnd cell_6t
Xbit_r145_c47 bl[47] br[47] wl[145] vdd gnd cell_6t
Xbit_r146_c47 bl[47] br[47] wl[146] vdd gnd cell_6t
Xbit_r147_c47 bl[47] br[47] wl[147] vdd gnd cell_6t
Xbit_r148_c47 bl[47] br[47] wl[148] vdd gnd cell_6t
Xbit_r149_c47 bl[47] br[47] wl[149] vdd gnd cell_6t
Xbit_r150_c47 bl[47] br[47] wl[150] vdd gnd cell_6t
Xbit_r151_c47 bl[47] br[47] wl[151] vdd gnd cell_6t
Xbit_r152_c47 bl[47] br[47] wl[152] vdd gnd cell_6t
Xbit_r153_c47 bl[47] br[47] wl[153] vdd gnd cell_6t
Xbit_r154_c47 bl[47] br[47] wl[154] vdd gnd cell_6t
Xbit_r155_c47 bl[47] br[47] wl[155] vdd gnd cell_6t
Xbit_r156_c47 bl[47] br[47] wl[156] vdd gnd cell_6t
Xbit_r157_c47 bl[47] br[47] wl[157] vdd gnd cell_6t
Xbit_r158_c47 bl[47] br[47] wl[158] vdd gnd cell_6t
Xbit_r159_c47 bl[47] br[47] wl[159] vdd gnd cell_6t
Xbit_r160_c47 bl[47] br[47] wl[160] vdd gnd cell_6t
Xbit_r161_c47 bl[47] br[47] wl[161] vdd gnd cell_6t
Xbit_r162_c47 bl[47] br[47] wl[162] vdd gnd cell_6t
Xbit_r163_c47 bl[47] br[47] wl[163] vdd gnd cell_6t
Xbit_r164_c47 bl[47] br[47] wl[164] vdd gnd cell_6t
Xbit_r165_c47 bl[47] br[47] wl[165] vdd gnd cell_6t
Xbit_r166_c47 bl[47] br[47] wl[166] vdd gnd cell_6t
Xbit_r167_c47 bl[47] br[47] wl[167] vdd gnd cell_6t
Xbit_r168_c47 bl[47] br[47] wl[168] vdd gnd cell_6t
Xbit_r169_c47 bl[47] br[47] wl[169] vdd gnd cell_6t
Xbit_r170_c47 bl[47] br[47] wl[170] vdd gnd cell_6t
Xbit_r171_c47 bl[47] br[47] wl[171] vdd gnd cell_6t
Xbit_r172_c47 bl[47] br[47] wl[172] vdd gnd cell_6t
Xbit_r173_c47 bl[47] br[47] wl[173] vdd gnd cell_6t
Xbit_r174_c47 bl[47] br[47] wl[174] vdd gnd cell_6t
Xbit_r175_c47 bl[47] br[47] wl[175] vdd gnd cell_6t
Xbit_r176_c47 bl[47] br[47] wl[176] vdd gnd cell_6t
Xbit_r177_c47 bl[47] br[47] wl[177] vdd gnd cell_6t
Xbit_r178_c47 bl[47] br[47] wl[178] vdd gnd cell_6t
Xbit_r179_c47 bl[47] br[47] wl[179] vdd gnd cell_6t
Xbit_r180_c47 bl[47] br[47] wl[180] vdd gnd cell_6t
Xbit_r181_c47 bl[47] br[47] wl[181] vdd gnd cell_6t
Xbit_r182_c47 bl[47] br[47] wl[182] vdd gnd cell_6t
Xbit_r183_c47 bl[47] br[47] wl[183] vdd gnd cell_6t
Xbit_r184_c47 bl[47] br[47] wl[184] vdd gnd cell_6t
Xbit_r185_c47 bl[47] br[47] wl[185] vdd gnd cell_6t
Xbit_r186_c47 bl[47] br[47] wl[186] vdd gnd cell_6t
Xbit_r187_c47 bl[47] br[47] wl[187] vdd gnd cell_6t
Xbit_r188_c47 bl[47] br[47] wl[188] vdd gnd cell_6t
Xbit_r189_c47 bl[47] br[47] wl[189] vdd gnd cell_6t
Xbit_r190_c47 bl[47] br[47] wl[190] vdd gnd cell_6t
Xbit_r191_c47 bl[47] br[47] wl[191] vdd gnd cell_6t
Xbit_r192_c47 bl[47] br[47] wl[192] vdd gnd cell_6t
Xbit_r193_c47 bl[47] br[47] wl[193] vdd gnd cell_6t
Xbit_r194_c47 bl[47] br[47] wl[194] vdd gnd cell_6t
Xbit_r195_c47 bl[47] br[47] wl[195] vdd gnd cell_6t
Xbit_r196_c47 bl[47] br[47] wl[196] vdd gnd cell_6t
Xbit_r197_c47 bl[47] br[47] wl[197] vdd gnd cell_6t
Xbit_r198_c47 bl[47] br[47] wl[198] vdd gnd cell_6t
Xbit_r199_c47 bl[47] br[47] wl[199] vdd gnd cell_6t
Xbit_r200_c47 bl[47] br[47] wl[200] vdd gnd cell_6t
Xbit_r201_c47 bl[47] br[47] wl[201] vdd gnd cell_6t
Xbit_r202_c47 bl[47] br[47] wl[202] vdd gnd cell_6t
Xbit_r203_c47 bl[47] br[47] wl[203] vdd gnd cell_6t
Xbit_r204_c47 bl[47] br[47] wl[204] vdd gnd cell_6t
Xbit_r205_c47 bl[47] br[47] wl[205] vdd gnd cell_6t
Xbit_r206_c47 bl[47] br[47] wl[206] vdd gnd cell_6t
Xbit_r207_c47 bl[47] br[47] wl[207] vdd gnd cell_6t
Xbit_r208_c47 bl[47] br[47] wl[208] vdd gnd cell_6t
Xbit_r209_c47 bl[47] br[47] wl[209] vdd gnd cell_6t
Xbit_r210_c47 bl[47] br[47] wl[210] vdd gnd cell_6t
Xbit_r211_c47 bl[47] br[47] wl[211] vdd gnd cell_6t
Xbit_r212_c47 bl[47] br[47] wl[212] vdd gnd cell_6t
Xbit_r213_c47 bl[47] br[47] wl[213] vdd gnd cell_6t
Xbit_r214_c47 bl[47] br[47] wl[214] vdd gnd cell_6t
Xbit_r215_c47 bl[47] br[47] wl[215] vdd gnd cell_6t
Xbit_r216_c47 bl[47] br[47] wl[216] vdd gnd cell_6t
Xbit_r217_c47 bl[47] br[47] wl[217] vdd gnd cell_6t
Xbit_r218_c47 bl[47] br[47] wl[218] vdd gnd cell_6t
Xbit_r219_c47 bl[47] br[47] wl[219] vdd gnd cell_6t
Xbit_r220_c47 bl[47] br[47] wl[220] vdd gnd cell_6t
Xbit_r221_c47 bl[47] br[47] wl[221] vdd gnd cell_6t
Xbit_r222_c47 bl[47] br[47] wl[222] vdd gnd cell_6t
Xbit_r223_c47 bl[47] br[47] wl[223] vdd gnd cell_6t
Xbit_r224_c47 bl[47] br[47] wl[224] vdd gnd cell_6t
Xbit_r225_c47 bl[47] br[47] wl[225] vdd gnd cell_6t
Xbit_r226_c47 bl[47] br[47] wl[226] vdd gnd cell_6t
Xbit_r227_c47 bl[47] br[47] wl[227] vdd gnd cell_6t
Xbit_r228_c47 bl[47] br[47] wl[228] vdd gnd cell_6t
Xbit_r229_c47 bl[47] br[47] wl[229] vdd gnd cell_6t
Xbit_r230_c47 bl[47] br[47] wl[230] vdd gnd cell_6t
Xbit_r231_c47 bl[47] br[47] wl[231] vdd gnd cell_6t
Xbit_r232_c47 bl[47] br[47] wl[232] vdd gnd cell_6t
Xbit_r233_c47 bl[47] br[47] wl[233] vdd gnd cell_6t
Xbit_r234_c47 bl[47] br[47] wl[234] vdd gnd cell_6t
Xbit_r235_c47 bl[47] br[47] wl[235] vdd gnd cell_6t
Xbit_r236_c47 bl[47] br[47] wl[236] vdd gnd cell_6t
Xbit_r237_c47 bl[47] br[47] wl[237] vdd gnd cell_6t
Xbit_r238_c47 bl[47] br[47] wl[238] vdd gnd cell_6t
Xbit_r239_c47 bl[47] br[47] wl[239] vdd gnd cell_6t
Xbit_r240_c47 bl[47] br[47] wl[240] vdd gnd cell_6t
Xbit_r241_c47 bl[47] br[47] wl[241] vdd gnd cell_6t
Xbit_r242_c47 bl[47] br[47] wl[242] vdd gnd cell_6t
Xbit_r243_c47 bl[47] br[47] wl[243] vdd gnd cell_6t
Xbit_r244_c47 bl[47] br[47] wl[244] vdd gnd cell_6t
Xbit_r245_c47 bl[47] br[47] wl[245] vdd gnd cell_6t
Xbit_r246_c47 bl[47] br[47] wl[246] vdd gnd cell_6t
Xbit_r247_c47 bl[47] br[47] wl[247] vdd gnd cell_6t
Xbit_r248_c47 bl[47] br[47] wl[248] vdd gnd cell_6t
Xbit_r249_c47 bl[47] br[47] wl[249] vdd gnd cell_6t
Xbit_r250_c47 bl[47] br[47] wl[250] vdd gnd cell_6t
Xbit_r251_c47 bl[47] br[47] wl[251] vdd gnd cell_6t
Xbit_r252_c47 bl[47] br[47] wl[252] vdd gnd cell_6t
Xbit_r253_c47 bl[47] br[47] wl[253] vdd gnd cell_6t
Xbit_r254_c47 bl[47] br[47] wl[254] vdd gnd cell_6t
Xbit_r255_c47 bl[47] br[47] wl[255] vdd gnd cell_6t
Xbit_r256_c47 bl[47] br[47] wl[256] vdd gnd cell_6t
Xbit_r257_c47 bl[47] br[47] wl[257] vdd gnd cell_6t
Xbit_r258_c47 bl[47] br[47] wl[258] vdd gnd cell_6t
Xbit_r259_c47 bl[47] br[47] wl[259] vdd gnd cell_6t
Xbit_r260_c47 bl[47] br[47] wl[260] vdd gnd cell_6t
Xbit_r261_c47 bl[47] br[47] wl[261] vdd gnd cell_6t
Xbit_r262_c47 bl[47] br[47] wl[262] vdd gnd cell_6t
Xbit_r263_c47 bl[47] br[47] wl[263] vdd gnd cell_6t
Xbit_r264_c47 bl[47] br[47] wl[264] vdd gnd cell_6t
Xbit_r265_c47 bl[47] br[47] wl[265] vdd gnd cell_6t
Xbit_r266_c47 bl[47] br[47] wl[266] vdd gnd cell_6t
Xbit_r267_c47 bl[47] br[47] wl[267] vdd gnd cell_6t
Xbit_r268_c47 bl[47] br[47] wl[268] vdd gnd cell_6t
Xbit_r269_c47 bl[47] br[47] wl[269] vdd gnd cell_6t
Xbit_r270_c47 bl[47] br[47] wl[270] vdd gnd cell_6t
Xbit_r271_c47 bl[47] br[47] wl[271] vdd gnd cell_6t
Xbit_r272_c47 bl[47] br[47] wl[272] vdd gnd cell_6t
Xbit_r273_c47 bl[47] br[47] wl[273] vdd gnd cell_6t
Xbit_r274_c47 bl[47] br[47] wl[274] vdd gnd cell_6t
Xbit_r275_c47 bl[47] br[47] wl[275] vdd gnd cell_6t
Xbit_r276_c47 bl[47] br[47] wl[276] vdd gnd cell_6t
Xbit_r277_c47 bl[47] br[47] wl[277] vdd gnd cell_6t
Xbit_r278_c47 bl[47] br[47] wl[278] vdd gnd cell_6t
Xbit_r279_c47 bl[47] br[47] wl[279] vdd gnd cell_6t
Xbit_r280_c47 bl[47] br[47] wl[280] vdd gnd cell_6t
Xbit_r281_c47 bl[47] br[47] wl[281] vdd gnd cell_6t
Xbit_r282_c47 bl[47] br[47] wl[282] vdd gnd cell_6t
Xbit_r283_c47 bl[47] br[47] wl[283] vdd gnd cell_6t
Xbit_r284_c47 bl[47] br[47] wl[284] vdd gnd cell_6t
Xbit_r285_c47 bl[47] br[47] wl[285] vdd gnd cell_6t
Xbit_r286_c47 bl[47] br[47] wl[286] vdd gnd cell_6t
Xbit_r287_c47 bl[47] br[47] wl[287] vdd gnd cell_6t
Xbit_r288_c47 bl[47] br[47] wl[288] vdd gnd cell_6t
Xbit_r289_c47 bl[47] br[47] wl[289] vdd gnd cell_6t
Xbit_r290_c47 bl[47] br[47] wl[290] vdd gnd cell_6t
Xbit_r291_c47 bl[47] br[47] wl[291] vdd gnd cell_6t
Xbit_r292_c47 bl[47] br[47] wl[292] vdd gnd cell_6t
Xbit_r293_c47 bl[47] br[47] wl[293] vdd gnd cell_6t
Xbit_r294_c47 bl[47] br[47] wl[294] vdd gnd cell_6t
Xbit_r295_c47 bl[47] br[47] wl[295] vdd gnd cell_6t
Xbit_r296_c47 bl[47] br[47] wl[296] vdd gnd cell_6t
Xbit_r297_c47 bl[47] br[47] wl[297] vdd gnd cell_6t
Xbit_r298_c47 bl[47] br[47] wl[298] vdd gnd cell_6t
Xbit_r299_c47 bl[47] br[47] wl[299] vdd gnd cell_6t
Xbit_r300_c47 bl[47] br[47] wl[300] vdd gnd cell_6t
Xbit_r301_c47 bl[47] br[47] wl[301] vdd gnd cell_6t
Xbit_r302_c47 bl[47] br[47] wl[302] vdd gnd cell_6t
Xbit_r303_c47 bl[47] br[47] wl[303] vdd gnd cell_6t
Xbit_r304_c47 bl[47] br[47] wl[304] vdd gnd cell_6t
Xbit_r305_c47 bl[47] br[47] wl[305] vdd gnd cell_6t
Xbit_r306_c47 bl[47] br[47] wl[306] vdd gnd cell_6t
Xbit_r307_c47 bl[47] br[47] wl[307] vdd gnd cell_6t
Xbit_r308_c47 bl[47] br[47] wl[308] vdd gnd cell_6t
Xbit_r309_c47 bl[47] br[47] wl[309] vdd gnd cell_6t
Xbit_r310_c47 bl[47] br[47] wl[310] vdd gnd cell_6t
Xbit_r311_c47 bl[47] br[47] wl[311] vdd gnd cell_6t
Xbit_r312_c47 bl[47] br[47] wl[312] vdd gnd cell_6t
Xbit_r313_c47 bl[47] br[47] wl[313] vdd gnd cell_6t
Xbit_r314_c47 bl[47] br[47] wl[314] vdd gnd cell_6t
Xbit_r315_c47 bl[47] br[47] wl[315] vdd gnd cell_6t
Xbit_r316_c47 bl[47] br[47] wl[316] vdd gnd cell_6t
Xbit_r317_c47 bl[47] br[47] wl[317] vdd gnd cell_6t
Xbit_r318_c47 bl[47] br[47] wl[318] vdd gnd cell_6t
Xbit_r319_c47 bl[47] br[47] wl[319] vdd gnd cell_6t
Xbit_r320_c47 bl[47] br[47] wl[320] vdd gnd cell_6t
Xbit_r321_c47 bl[47] br[47] wl[321] vdd gnd cell_6t
Xbit_r322_c47 bl[47] br[47] wl[322] vdd gnd cell_6t
Xbit_r323_c47 bl[47] br[47] wl[323] vdd gnd cell_6t
Xbit_r324_c47 bl[47] br[47] wl[324] vdd gnd cell_6t
Xbit_r325_c47 bl[47] br[47] wl[325] vdd gnd cell_6t
Xbit_r326_c47 bl[47] br[47] wl[326] vdd gnd cell_6t
Xbit_r327_c47 bl[47] br[47] wl[327] vdd gnd cell_6t
Xbit_r328_c47 bl[47] br[47] wl[328] vdd gnd cell_6t
Xbit_r329_c47 bl[47] br[47] wl[329] vdd gnd cell_6t
Xbit_r330_c47 bl[47] br[47] wl[330] vdd gnd cell_6t
Xbit_r331_c47 bl[47] br[47] wl[331] vdd gnd cell_6t
Xbit_r332_c47 bl[47] br[47] wl[332] vdd gnd cell_6t
Xbit_r333_c47 bl[47] br[47] wl[333] vdd gnd cell_6t
Xbit_r334_c47 bl[47] br[47] wl[334] vdd gnd cell_6t
Xbit_r335_c47 bl[47] br[47] wl[335] vdd gnd cell_6t
Xbit_r336_c47 bl[47] br[47] wl[336] vdd gnd cell_6t
Xbit_r337_c47 bl[47] br[47] wl[337] vdd gnd cell_6t
Xbit_r338_c47 bl[47] br[47] wl[338] vdd gnd cell_6t
Xbit_r339_c47 bl[47] br[47] wl[339] vdd gnd cell_6t
Xbit_r340_c47 bl[47] br[47] wl[340] vdd gnd cell_6t
Xbit_r341_c47 bl[47] br[47] wl[341] vdd gnd cell_6t
Xbit_r342_c47 bl[47] br[47] wl[342] vdd gnd cell_6t
Xbit_r343_c47 bl[47] br[47] wl[343] vdd gnd cell_6t
Xbit_r344_c47 bl[47] br[47] wl[344] vdd gnd cell_6t
Xbit_r345_c47 bl[47] br[47] wl[345] vdd gnd cell_6t
Xbit_r346_c47 bl[47] br[47] wl[346] vdd gnd cell_6t
Xbit_r347_c47 bl[47] br[47] wl[347] vdd gnd cell_6t
Xbit_r348_c47 bl[47] br[47] wl[348] vdd gnd cell_6t
Xbit_r349_c47 bl[47] br[47] wl[349] vdd gnd cell_6t
Xbit_r350_c47 bl[47] br[47] wl[350] vdd gnd cell_6t
Xbit_r351_c47 bl[47] br[47] wl[351] vdd gnd cell_6t
Xbit_r352_c47 bl[47] br[47] wl[352] vdd gnd cell_6t
Xbit_r353_c47 bl[47] br[47] wl[353] vdd gnd cell_6t
Xbit_r354_c47 bl[47] br[47] wl[354] vdd gnd cell_6t
Xbit_r355_c47 bl[47] br[47] wl[355] vdd gnd cell_6t
Xbit_r356_c47 bl[47] br[47] wl[356] vdd gnd cell_6t
Xbit_r357_c47 bl[47] br[47] wl[357] vdd gnd cell_6t
Xbit_r358_c47 bl[47] br[47] wl[358] vdd gnd cell_6t
Xbit_r359_c47 bl[47] br[47] wl[359] vdd gnd cell_6t
Xbit_r360_c47 bl[47] br[47] wl[360] vdd gnd cell_6t
Xbit_r361_c47 bl[47] br[47] wl[361] vdd gnd cell_6t
Xbit_r362_c47 bl[47] br[47] wl[362] vdd gnd cell_6t
Xbit_r363_c47 bl[47] br[47] wl[363] vdd gnd cell_6t
Xbit_r364_c47 bl[47] br[47] wl[364] vdd gnd cell_6t
Xbit_r365_c47 bl[47] br[47] wl[365] vdd gnd cell_6t
Xbit_r366_c47 bl[47] br[47] wl[366] vdd gnd cell_6t
Xbit_r367_c47 bl[47] br[47] wl[367] vdd gnd cell_6t
Xbit_r368_c47 bl[47] br[47] wl[368] vdd gnd cell_6t
Xbit_r369_c47 bl[47] br[47] wl[369] vdd gnd cell_6t
Xbit_r370_c47 bl[47] br[47] wl[370] vdd gnd cell_6t
Xbit_r371_c47 bl[47] br[47] wl[371] vdd gnd cell_6t
Xbit_r372_c47 bl[47] br[47] wl[372] vdd gnd cell_6t
Xbit_r373_c47 bl[47] br[47] wl[373] vdd gnd cell_6t
Xbit_r374_c47 bl[47] br[47] wl[374] vdd gnd cell_6t
Xbit_r375_c47 bl[47] br[47] wl[375] vdd gnd cell_6t
Xbit_r376_c47 bl[47] br[47] wl[376] vdd gnd cell_6t
Xbit_r377_c47 bl[47] br[47] wl[377] vdd gnd cell_6t
Xbit_r378_c47 bl[47] br[47] wl[378] vdd gnd cell_6t
Xbit_r379_c47 bl[47] br[47] wl[379] vdd gnd cell_6t
Xbit_r380_c47 bl[47] br[47] wl[380] vdd gnd cell_6t
Xbit_r381_c47 bl[47] br[47] wl[381] vdd gnd cell_6t
Xbit_r382_c47 bl[47] br[47] wl[382] vdd gnd cell_6t
Xbit_r383_c47 bl[47] br[47] wl[383] vdd gnd cell_6t
Xbit_r384_c47 bl[47] br[47] wl[384] vdd gnd cell_6t
Xbit_r385_c47 bl[47] br[47] wl[385] vdd gnd cell_6t
Xbit_r386_c47 bl[47] br[47] wl[386] vdd gnd cell_6t
Xbit_r387_c47 bl[47] br[47] wl[387] vdd gnd cell_6t
Xbit_r388_c47 bl[47] br[47] wl[388] vdd gnd cell_6t
Xbit_r389_c47 bl[47] br[47] wl[389] vdd gnd cell_6t
Xbit_r390_c47 bl[47] br[47] wl[390] vdd gnd cell_6t
Xbit_r391_c47 bl[47] br[47] wl[391] vdd gnd cell_6t
Xbit_r392_c47 bl[47] br[47] wl[392] vdd gnd cell_6t
Xbit_r393_c47 bl[47] br[47] wl[393] vdd gnd cell_6t
Xbit_r394_c47 bl[47] br[47] wl[394] vdd gnd cell_6t
Xbit_r395_c47 bl[47] br[47] wl[395] vdd gnd cell_6t
Xbit_r396_c47 bl[47] br[47] wl[396] vdd gnd cell_6t
Xbit_r397_c47 bl[47] br[47] wl[397] vdd gnd cell_6t
Xbit_r398_c47 bl[47] br[47] wl[398] vdd gnd cell_6t
Xbit_r399_c47 bl[47] br[47] wl[399] vdd gnd cell_6t
Xbit_r400_c47 bl[47] br[47] wl[400] vdd gnd cell_6t
Xbit_r401_c47 bl[47] br[47] wl[401] vdd gnd cell_6t
Xbit_r402_c47 bl[47] br[47] wl[402] vdd gnd cell_6t
Xbit_r403_c47 bl[47] br[47] wl[403] vdd gnd cell_6t
Xbit_r404_c47 bl[47] br[47] wl[404] vdd gnd cell_6t
Xbit_r405_c47 bl[47] br[47] wl[405] vdd gnd cell_6t
Xbit_r406_c47 bl[47] br[47] wl[406] vdd gnd cell_6t
Xbit_r407_c47 bl[47] br[47] wl[407] vdd gnd cell_6t
Xbit_r408_c47 bl[47] br[47] wl[408] vdd gnd cell_6t
Xbit_r409_c47 bl[47] br[47] wl[409] vdd gnd cell_6t
Xbit_r410_c47 bl[47] br[47] wl[410] vdd gnd cell_6t
Xbit_r411_c47 bl[47] br[47] wl[411] vdd gnd cell_6t
Xbit_r412_c47 bl[47] br[47] wl[412] vdd gnd cell_6t
Xbit_r413_c47 bl[47] br[47] wl[413] vdd gnd cell_6t
Xbit_r414_c47 bl[47] br[47] wl[414] vdd gnd cell_6t
Xbit_r415_c47 bl[47] br[47] wl[415] vdd gnd cell_6t
Xbit_r416_c47 bl[47] br[47] wl[416] vdd gnd cell_6t
Xbit_r417_c47 bl[47] br[47] wl[417] vdd gnd cell_6t
Xbit_r418_c47 bl[47] br[47] wl[418] vdd gnd cell_6t
Xbit_r419_c47 bl[47] br[47] wl[419] vdd gnd cell_6t
Xbit_r420_c47 bl[47] br[47] wl[420] vdd gnd cell_6t
Xbit_r421_c47 bl[47] br[47] wl[421] vdd gnd cell_6t
Xbit_r422_c47 bl[47] br[47] wl[422] vdd gnd cell_6t
Xbit_r423_c47 bl[47] br[47] wl[423] vdd gnd cell_6t
Xbit_r424_c47 bl[47] br[47] wl[424] vdd gnd cell_6t
Xbit_r425_c47 bl[47] br[47] wl[425] vdd gnd cell_6t
Xbit_r426_c47 bl[47] br[47] wl[426] vdd gnd cell_6t
Xbit_r427_c47 bl[47] br[47] wl[427] vdd gnd cell_6t
Xbit_r428_c47 bl[47] br[47] wl[428] vdd gnd cell_6t
Xbit_r429_c47 bl[47] br[47] wl[429] vdd gnd cell_6t
Xbit_r430_c47 bl[47] br[47] wl[430] vdd gnd cell_6t
Xbit_r431_c47 bl[47] br[47] wl[431] vdd gnd cell_6t
Xbit_r432_c47 bl[47] br[47] wl[432] vdd gnd cell_6t
Xbit_r433_c47 bl[47] br[47] wl[433] vdd gnd cell_6t
Xbit_r434_c47 bl[47] br[47] wl[434] vdd gnd cell_6t
Xbit_r435_c47 bl[47] br[47] wl[435] vdd gnd cell_6t
Xbit_r436_c47 bl[47] br[47] wl[436] vdd gnd cell_6t
Xbit_r437_c47 bl[47] br[47] wl[437] vdd gnd cell_6t
Xbit_r438_c47 bl[47] br[47] wl[438] vdd gnd cell_6t
Xbit_r439_c47 bl[47] br[47] wl[439] vdd gnd cell_6t
Xbit_r440_c47 bl[47] br[47] wl[440] vdd gnd cell_6t
Xbit_r441_c47 bl[47] br[47] wl[441] vdd gnd cell_6t
Xbit_r442_c47 bl[47] br[47] wl[442] vdd gnd cell_6t
Xbit_r443_c47 bl[47] br[47] wl[443] vdd gnd cell_6t
Xbit_r444_c47 bl[47] br[47] wl[444] vdd gnd cell_6t
Xbit_r445_c47 bl[47] br[47] wl[445] vdd gnd cell_6t
Xbit_r446_c47 bl[47] br[47] wl[446] vdd gnd cell_6t
Xbit_r447_c47 bl[47] br[47] wl[447] vdd gnd cell_6t
Xbit_r448_c47 bl[47] br[47] wl[448] vdd gnd cell_6t
Xbit_r449_c47 bl[47] br[47] wl[449] vdd gnd cell_6t
Xbit_r450_c47 bl[47] br[47] wl[450] vdd gnd cell_6t
Xbit_r451_c47 bl[47] br[47] wl[451] vdd gnd cell_6t
Xbit_r452_c47 bl[47] br[47] wl[452] vdd gnd cell_6t
Xbit_r453_c47 bl[47] br[47] wl[453] vdd gnd cell_6t
Xbit_r454_c47 bl[47] br[47] wl[454] vdd gnd cell_6t
Xbit_r455_c47 bl[47] br[47] wl[455] vdd gnd cell_6t
Xbit_r456_c47 bl[47] br[47] wl[456] vdd gnd cell_6t
Xbit_r457_c47 bl[47] br[47] wl[457] vdd gnd cell_6t
Xbit_r458_c47 bl[47] br[47] wl[458] vdd gnd cell_6t
Xbit_r459_c47 bl[47] br[47] wl[459] vdd gnd cell_6t
Xbit_r460_c47 bl[47] br[47] wl[460] vdd gnd cell_6t
Xbit_r461_c47 bl[47] br[47] wl[461] vdd gnd cell_6t
Xbit_r462_c47 bl[47] br[47] wl[462] vdd gnd cell_6t
Xbit_r463_c47 bl[47] br[47] wl[463] vdd gnd cell_6t
Xbit_r464_c47 bl[47] br[47] wl[464] vdd gnd cell_6t
Xbit_r465_c47 bl[47] br[47] wl[465] vdd gnd cell_6t
Xbit_r466_c47 bl[47] br[47] wl[466] vdd gnd cell_6t
Xbit_r467_c47 bl[47] br[47] wl[467] vdd gnd cell_6t
Xbit_r468_c47 bl[47] br[47] wl[468] vdd gnd cell_6t
Xbit_r469_c47 bl[47] br[47] wl[469] vdd gnd cell_6t
Xbit_r470_c47 bl[47] br[47] wl[470] vdd gnd cell_6t
Xbit_r471_c47 bl[47] br[47] wl[471] vdd gnd cell_6t
Xbit_r472_c47 bl[47] br[47] wl[472] vdd gnd cell_6t
Xbit_r473_c47 bl[47] br[47] wl[473] vdd gnd cell_6t
Xbit_r474_c47 bl[47] br[47] wl[474] vdd gnd cell_6t
Xbit_r475_c47 bl[47] br[47] wl[475] vdd gnd cell_6t
Xbit_r476_c47 bl[47] br[47] wl[476] vdd gnd cell_6t
Xbit_r477_c47 bl[47] br[47] wl[477] vdd gnd cell_6t
Xbit_r478_c47 bl[47] br[47] wl[478] vdd gnd cell_6t
Xbit_r479_c47 bl[47] br[47] wl[479] vdd gnd cell_6t
Xbit_r480_c47 bl[47] br[47] wl[480] vdd gnd cell_6t
Xbit_r481_c47 bl[47] br[47] wl[481] vdd gnd cell_6t
Xbit_r482_c47 bl[47] br[47] wl[482] vdd gnd cell_6t
Xbit_r483_c47 bl[47] br[47] wl[483] vdd gnd cell_6t
Xbit_r484_c47 bl[47] br[47] wl[484] vdd gnd cell_6t
Xbit_r485_c47 bl[47] br[47] wl[485] vdd gnd cell_6t
Xbit_r486_c47 bl[47] br[47] wl[486] vdd gnd cell_6t
Xbit_r487_c47 bl[47] br[47] wl[487] vdd gnd cell_6t
Xbit_r488_c47 bl[47] br[47] wl[488] vdd gnd cell_6t
Xbit_r489_c47 bl[47] br[47] wl[489] vdd gnd cell_6t
Xbit_r490_c47 bl[47] br[47] wl[490] vdd gnd cell_6t
Xbit_r491_c47 bl[47] br[47] wl[491] vdd gnd cell_6t
Xbit_r492_c47 bl[47] br[47] wl[492] vdd gnd cell_6t
Xbit_r493_c47 bl[47] br[47] wl[493] vdd gnd cell_6t
Xbit_r494_c47 bl[47] br[47] wl[494] vdd gnd cell_6t
Xbit_r495_c47 bl[47] br[47] wl[495] vdd gnd cell_6t
Xbit_r496_c47 bl[47] br[47] wl[496] vdd gnd cell_6t
Xbit_r497_c47 bl[47] br[47] wl[497] vdd gnd cell_6t
Xbit_r498_c47 bl[47] br[47] wl[498] vdd gnd cell_6t
Xbit_r499_c47 bl[47] br[47] wl[499] vdd gnd cell_6t
Xbit_r500_c47 bl[47] br[47] wl[500] vdd gnd cell_6t
Xbit_r501_c47 bl[47] br[47] wl[501] vdd gnd cell_6t
Xbit_r502_c47 bl[47] br[47] wl[502] vdd gnd cell_6t
Xbit_r503_c47 bl[47] br[47] wl[503] vdd gnd cell_6t
Xbit_r504_c47 bl[47] br[47] wl[504] vdd gnd cell_6t
Xbit_r505_c47 bl[47] br[47] wl[505] vdd gnd cell_6t
Xbit_r506_c47 bl[47] br[47] wl[506] vdd gnd cell_6t
Xbit_r507_c47 bl[47] br[47] wl[507] vdd gnd cell_6t
Xbit_r508_c47 bl[47] br[47] wl[508] vdd gnd cell_6t
Xbit_r509_c47 bl[47] br[47] wl[509] vdd gnd cell_6t
Xbit_r510_c47 bl[47] br[47] wl[510] vdd gnd cell_6t
Xbit_r511_c47 bl[47] br[47] wl[511] vdd gnd cell_6t
Xbit_r0_c48 bl[48] br[48] wl[0] vdd gnd cell_6t
Xbit_r1_c48 bl[48] br[48] wl[1] vdd gnd cell_6t
Xbit_r2_c48 bl[48] br[48] wl[2] vdd gnd cell_6t
Xbit_r3_c48 bl[48] br[48] wl[3] vdd gnd cell_6t
Xbit_r4_c48 bl[48] br[48] wl[4] vdd gnd cell_6t
Xbit_r5_c48 bl[48] br[48] wl[5] vdd gnd cell_6t
Xbit_r6_c48 bl[48] br[48] wl[6] vdd gnd cell_6t
Xbit_r7_c48 bl[48] br[48] wl[7] vdd gnd cell_6t
Xbit_r8_c48 bl[48] br[48] wl[8] vdd gnd cell_6t
Xbit_r9_c48 bl[48] br[48] wl[9] vdd gnd cell_6t
Xbit_r10_c48 bl[48] br[48] wl[10] vdd gnd cell_6t
Xbit_r11_c48 bl[48] br[48] wl[11] vdd gnd cell_6t
Xbit_r12_c48 bl[48] br[48] wl[12] vdd gnd cell_6t
Xbit_r13_c48 bl[48] br[48] wl[13] vdd gnd cell_6t
Xbit_r14_c48 bl[48] br[48] wl[14] vdd gnd cell_6t
Xbit_r15_c48 bl[48] br[48] wl[15] vdd gnd cell_6t
Xbit_r16_c48 bl[48] br[48] wl[16] vdd gnd cell_6t
Xbit_r17_c48 bl[48] br[48] wl[17] vdd gnd cell_6t
Xbit_r18_c48 bl[48] br[48] wl[18] vdd gnd cell_6t
Xbit_r19_c48 bl[48] br[48] wl[19] vdd gnd cell_6t
Xbit_r20_c48 bl[48] br[48] wl[20] vdd gnd cell_6t
Xbit_r21_c48 bl[48] br[48] wl[21] vdd gnd cell_6t
Xbit_r22_c48 bl[48] br[48] wl[22] vdd gnd cell_6t
Xbit_r23_c48 bl[48] br[48] wl[23] vdd gnd cell_6t
Xbit_r24_c48 bl[48] br[48] wl[24] vdd gnd cell_6t
Xbit_r25_c48 bl[48] br[48] wl[25] vdd gnd cell_6t
Xbit_r26_c48 bl[48] br[48] wl[26] vdd gnd cell_6t
Xbit_r27_c48 bl[48] br[48] wl[27] vdd gnd cell_6t
Xbit_r28_c48 bl[48] br[48] wl[28] vdd gnd cell_6t
Xbit_r29_c48 bl[48] br[48] wl[29] vdd gnd cell_6t
Xbit_r30_c48 bl[48] br[48] wl[30] vdd gnd cell_6t
Xbit_r31_c48 bl[48] br[48] wl[31] vdd gnd cell_6t
Xbit_r32_c48 bl[48] br[48] wl[32] vdd gnd cell_6t
Xbit_r33_c48 bl[48] br[48] wl[33] vdd gnd cell_6t
Xbit_r34_c48 bl[48] br[48] wl[34] vdd gnd cell_6t
Xbit_r35_c48 bl[48] br[48] wl[35] vdd gnd cell_6t
Xbit_r36_c48 bl[48] br[48] wl[36] vdd gnd cell_6t
Xbit_r37_c48 bl[48] br[48] wl[37] vdd gnd cell_6t
Xbit_r38_c48 bl[48] br[48] wl[38] vdd gnd cell_6t
Xbit_r39_c48 bl[48] br[48] wl[39] vdd gnd cell_6t
Xbit_r40_c48 bl[48] br[48] wl[40] vdd gnd cell_6t
Xbit_r41_c48 bl[48] br[48] wl[41] vdd gnd cell_6t
Xbit_r42_c48 bl[48] br[48] wl[42] vdd gnd cell_6t
Xbit_r43_c48 bl[48] br[48] wl[43] vdd gnd cell_6t
Xbit_r44_c48 bl[48] br[48] wl[44] vdd gnd cell_6t
Xbit_r45_c48 bl[48] br[48] wl[45] vdd gnd cell_6t
Xbit_r46_c48 bl[48] br[48] wl[46] vdd gnd cell_6t
Xbit_r47_c48 bl[48] br[48] wl[47] vdd gnd cell_6t
Xbit_r48_c48 bl[48] br[48] wl[48] vdd gnd cell_6t
Xbit_r49_c48 bl[48] br[48] wl[49] vdd gnd cell_6t
Xbit_r50_c48 bl[48] br[48] wl[50] vdd gnd cell_6t
Xbit_r51_c48 bl[48] br[48] wl[51] vdd gnd cell_6t
Xbit_r52_c48 bl[48] br[48] wl[52] vdd gnd cell_6t
Xbit_r53_c48 bl[48] br[48] wl[53] vdd gnd cell_6t
Xbit_r54_c48 bl[48] br[48] wl[54] vdd gnd cell_6t
Xbit_r55_c48 bl[48] br[48] wl[55] vdd gnd cell_6t
Xbit_r56_c48 bl[48] br[48] wl[56] vdd gnd cell_6t
Xbit_r57_c48 bl[48] br[48] wl[57] vdd gnd cell_6t
Xbit_r58_c48 bl[48] br[48] wl[58] vdd gnd cell_6t
Xbit_r59_c48 bl[48] br[48] wl[59] vdd gnd cell_6t
Xbit_r60_c48 bl[48] br[48] wl[60] vdd gnd cell_6t
Xbit_r61_c48 bl[48] br[48] wl[61] vdd gnd cell_6t
Xbit_r62_c48 bl[48] br[48] wl[62] vdd gnd cell_6t
Xbit_r63_c48 bl[48] br[48] wl[63] vdd gnd cell_6t
Xbit_r64_c48 bl[48] br[48] wl[64] vdd gnd cell_6t
Xbit_r65_c48 bl[48] br[48] wl[65] vdd gnd cell_6t
Xbit_r66_c48 bl[48] br[48] wl[66] vdd gnd cell_6t
Xbit_r67_c48 bl[48] br[48] wl[67] vdd gnd cell_6t
Xbit_r68_c48 bl[48] br[48] wl[68] vdd gnd cell_6t
Xbit_r69_c48 bl[48] br[48] wl[69] vdd gnd cell_6t
Xbit_r70_c48 bl[48] br[48] wl[70] vdd gnd cell_6t
Xbit_r71_c48 bl[48] br[48] wl[71] vdd gnd cell_6t
Xbit_r72_c48 bl[48] br[48] wl[72] vdd gnd cell_6t
Xbit_r73_c48 bl[48] br[48] wl[73] vdd gnd cell_6t
Xbit_r74_c48 bl[48] br[48] wl[74] vdd gnd cell_6t
Xbit_r75_c48 bl[48] br[48] wl[75] vdd gnd cell_6t
Xbit_r76_c48 bl[48] br[48] wl[76] vdd gnd cell_6t
Xbit_r77_c48 bl[48] br[48] wl[77] vdd gnd cell_6t
Xbit_r78_c48 bl[48] br[48] wl[78] vdd gnd cell_6t
Xbit_r79_c48 bl[48] br[48] wl[79] vdd gnd cell_6t
Xbit_r80_c48 bl[48] br[48] wl[80] vdd gnd cell_6t
Xbit_r81_c48 bl[48] br[48] wl[81] vdd gnd cell_6t
Xbit_r82_c48 bl[48] br[48] wl[82] vdd gnd cell_6t
Xbit_r83_c48 bl[48] br[48] wl[83] vdd gnd cell_6t
Xbit_r84_c48 bl[48] br[48] wl[84] vdd gnd cell_6t
Xbit_r85_c48 bl[48] br[48] wl[85] vdd gnd cell_6t
Xbit_r86_c48 bl[48] br[48] wl[86] vdd gnd cell_6t
Xbit_r87_c48 bl[48] br[48] wl[87] vdd gnd cell_6t
Xbit_r88_c48 bl[48] br[48] wl[88] vdd gnd cell_6t
Xbit_r89_c48 bl[48] br[48] wl[89] vdd gnd cell_6t
Xbit_r90_c48 bl[48] br[48] wl[90] vdd gnd cell_6t
Xbit_r91_c48 bl[48] br[48] wl[91] vdd gnd cell_6t
Xbit_r92_c48 bl[48] br[48] wl[92] vdd gnd cell_6t
Xbit_r93_c48 bl[48] br[48] wl[93] vdd gnd cell_6t
Xbit_r94_c48 bl[48] br[48] wl[94] vdd gnd cell_6t
Xbit_r95_c48 bl[48] br[48] wl[95] vdd gnd cell_6t
Xbit_r96_c48 bl[48] br[48] wl[96] vdd gnd cell_6t
Xbit_r97_c48 bl[48] br[48] wl[97] vdd gnd cell_6t
Xbit_r98_c48 bl[48] br[48] wl[98] vdd gnd cell_6t
Xbit_r99_c48 bl[48] br[48] wl[99] vdd gnd cell_6t
Xbit_r100_c48 bl[48] br[48] wl[100] vdd gnd cell_6t
Xbit_r101_c48 bl[48] br[48] wl[101] vdd gnd cell_6t
Xbit_r102_c48 bl[48] br[48] wl[102] vdd gnd cell_6t
Xbit_r103_c48 bl[48] br[48] wl[103] vdd gnd cell_6t
Xbit_r104_c48 bl[48] br[48] wl[104] vdd gnd cell_6t
Xbit_r105_c48 bl[48] br[48] wl[105] vdd gnd cell_6t
Xbit_r106_c48 bl[48] br[48] wl[106] vdd gnd cell_6t
Xbit_r107_c48 bl[48] br[48] wl[107] vdd gnd cell_6t
Xbit_r108_c48 bl[48] br[48] wl[108] vdd gnd cell_6t
Xbit_r109_c48 bl[48] br[48] wl[109] vdd gnd cell_6t
Xbit_r110_c48 bl[48] br[48] wl[110] vdd gnd cell_6t
Xbit_r111_c48 bl[48] br[48] wl[111] vdd gnd cell_6t
Xbit_r112_c48 bl[48] br[48] wl[112] vdd gnd cell_6t
Xbit_r113_c48 bl[48] br[48] wl[113] vdd gnd cell_6t
Xbit_r114_c48 bl[48] br[48] wl[114] vdd gnd cell_6t
Xbit_r115_c48 bl[48] br[48] wl[115] vdd gnd cell_6t
Xbit_r116_c48 bl[48] br[48] wl[116] vdd gnd cell_6t
Xbit_r117_c48 bl[48] br[48] wl[117] vdd gnd cell_6t
Xbit_r118_c48 bl[48] br[48] wl[118] vdd gnd cell_6t
Xbit_r119_c48 bl[48] br[48] wl[119] vdd gnd cell_6t
Xbit_r120_c48 bl[48] br[48] wl[120] vdd gnd cell_6t
Xbit_r121_c48 bl[48] br[48] wl[121] vdd gnd cell_6t
Xbit_r122_c48 bl[48] br[48] wl[122] vdd gnd cell_6t
Xbit_r123_c48 bl[48] br[48] wl[123] vdd gnd cell_6t
Xbit_r124_c48 bl[48] br[48] wl[124] vdd gnd cell_6t
Xbit_r125_c48 bl[48] br[48] wl[125] vdd gnd cell_6t
Xbit_r126_c48 bl[48] br[48] wl[126] vdd gnd cell_6t
Xbit_r127_c48 bl[48] br[48] wl[127] vdd gnd cell_6t
Xbit_r128_c48 bl[48] br[48] wl[128] vdd gnd cell_6t
Xbit_r129_c48 bl[48] br[48] wl[129] vdd gnd cell_6t
Xbit_r130_c48 bl[48] br[48] wl[130] vdd gnd cell_6t
Xbit_r131_c48 bl[48] br[48] wl[131] vdd gnd cell_6t
Xbit_r132_c48 bl[48] br[48] wl[132] vdd gnd cell_6t
Xbit_r133_c48 bl[48] br[48] wl[133] vdd gnd cell_6t
Xbit_r134_c48 bl[48] br[48] wl[134] vdd gnd cell_6t
Xbit_r135_c48 bl[48] br[48] wl[135] vdd gnd cell_6t
Xbit_r136_c48 bl[48] br[48] wl[136] vdd gnd cell_6t
Xbit_r137_c48 bl[48] br[48] wl[137] vdd gnd cell_6t
Xbit_r138_c48 bl[48] br[48] wl[138] vdd gnd cell_6t
Xbit_r139_c48 bl[48] br[48] wl[139] vdd gnd cell_6t
Xbit_r140_c48 bl[48] br[48] wl[140] vdd gnd cell_6t
Xbit_r141_c48 bl[48] br[48] wl[141] vdd gnd cell_6t
Xbit_r142_c48 bl[48] br[48] wl[142] vdd gnd cell_6t
Xbit_r143_c48 bl[48] br[48] wl[143] vdd gnd cell_6t
Xbit_r144_c48 bl[48] br[48] wl[144] vdd gnd cell_6t
Xbit_r145_c48 bl[48] br[48] wl[145] vdd gnd cell_6t
Xbit_r146_c48 bl[48] br[48] wl[146] vdd gnd cell_6t
Xbit_r147_c48 bl[48] br[48] wl[147] vdd gnd cell_6t
Xbit_r148_c48 bl[48] br[48] wl[148] vdd gnd cell_6t
Xbit_r149_c48 bl[48] br[48] wl[149] vdd gnd cell_6t
Xbit_r150_c48 bl[48] br[48] wl[150] vdd gnd cell_6t
Xbit_r151_c48 bl[48] br[48] wl[151] vdd gnd cell_6t
Xbit_r152_c48 bl[48] br[48] wl[152] vdd gnd cell_6t
Xbit_r153_c48 bl[48] br[48] wl[153] vdd gnd cell_6t
Xbit_r154_c48 bl[48] br[48] wl[154] vdd gnd cell_6t
Xbit_r155_c48 bl[48] br[48] wl[155] vdd gnd cell_6t
Xbit_r156_c48 bl[48] br[48] wl[156] vdd gnd cell_6t
Xbit_r157_c48 bl[48] br[48] wl[157] vdd gnd cell_6t
Xbit_r158_c48 bl[48] br[48] wl[158] vdd gnd cell_6t
Xbit_r159_c48 bl[48] br[48] wl[159] vdd gnd cell_6t
Xbit_r160_c48 bl[48] br[48] wl[160] vdd gnd cell_6t
Xbit_r161_c48 bl[48] br[48] wl[161] vdd gnd cell_6t
Xbit_r162_c48 bl[48] br[48] wl[162] vdd gnd cell_6t
Xbit_r163_c48 bl[48] br[48] wl[163] vdd gnd cell_6t
Xbit_r164_c48 bl[48] br[48] wl[164] vdd gnd cell_6t
Xbit_r165_c48 bl[48] br[48] wl[165] vdd gnd cell_6t
Xbit_r166_c48 bl[48] br[48] wl[166] vdd gnd cell_6t
Xbit_r167_c48 bl[48] br[48] wl[167] vdd gnd cell_6t
Xbit_r168_c48 bl[48] br[48] wl[168] vdd gnd cell_6t
Xbit_r169_c48 bl[48] br[48] wl[169] vdd gnd cell_6t
Xbit_r170_c48 bl[48] br[48] wl[170] vdd gnd cell_6t
Xbit_r171_c48 bl[48] br[48] wl[171] vdd gnd cell_6t
Xbit_r172_c48 bl[48] br[48] wl[172] vdd gnd cell_6t
Xbit_r173_c48 bl[48] br[48] wl[173] vdd gnd cell_6t
Xbit_r174_c48 bl[48] br[48] wl[174] vdd gnd cell_6t
Xbit_r175_c48 bl[48] br[48] wl[175] vdd gnd cell_6t
Xbit_r176_c48 bl[48] br[48] wl[176] vdd gnd cell_6t
Xbit_r177_c48 bl[48] br[48] wl[177] vdd gnd cell_6t
Xbit_r178_c48 bl[48] br[48] wl[178] vdd gnd cell_6t
Xbit_r179_c48 bl[48] br[48] wl[179] vdd gnd cell_6t
Xbit_r180_c48 bl[48] br[48] wl[180] vdd gnd cell_6t
Xbit_r181_c48 bl[48] br[48] wl[181] vdd gnd cell_6t
Xbit_r182_c48 bl[48] br[48] wl[182] vdd gnd cell_6t
Xbit_r183_c48 bl[48] br[48] wl[183] vdd gnd cell_6t
Xbit_r184_c48 bl[48] br[48] wl[184] vdd gnd cell_6t
Xbit_r185_c48 bl[48] br[48] wl[185] vdd gnd cell_6t
Xbit_r186_c48 bl[48] br[48] wl[186] vdd gnd cell_6t
Xbit_r187_c48 bl[48] br[48] wl[187] vdd gnd cell_6t
Xbit_r188_c48 bl[48] br[48] wl[188] vdd gnd cell_6t
Xbit_r189_c48 bl[48] br[48] wl[189] vdd gnd cell_6t
Xbit_r190_c48 bl[48] br[48] wl[190] vdd gnd cell_6t
Xbit_r191_c48 bl[48] br[48] wl[191] vdd gnd cell_6t
Xbit_r192_c48 bl[48] br[48] wl[192] vdd gnd cell_6t
Xbit_r193_c48 bl[48] br[48] wl[193] vdd gnd cell_6t
Xbit_r194_c48 bl[48] br[48] wl[194] vdd gnd cell_6t
Xbit_r195_c48 bl[48] br[48] wl[195] vdd gnd cell_6t
Xbit_r196_c48 bl[48] br[48] wl[196] vdd gnd cell_6t
Xbit_r197_c48 bl[48] br[48] wl[197] vdd gnd cell_6t
Xbit_r198_c48 bl[48] br[48] wl[198] vdd gnd cell_6t
Xbit_r199_c48 bl[48] br[48] wl[199] vdd gnd cell_6t
Xbit_r200_c48 bl[48] br[48] wl[200] vdd gnd cell_6t
Xbit_r201_c48 bl[48] br[48] wl[201] vdd gnd cell_6t
Xbit_r202_c48 bl[48] br[48] wl[202] vdd gnd cell_6t
Xbit_r203_c48 bl[48] br[48] wl[203] vdd gnd cell_6t
Xbit_r204_c48 bl[48] br[48] wl[204] vdd gnd cell_6t
Xbit_r205_c48 bl[48] br[48] wl[205] vdd gnd cell_6t
Xbit_r206_c48 bl[48] br[48] wl[206] vdd gnd cell_6t
Xbit_r207_c48 bl[48] br[48] wl[207] vdd gnd cell_6t
Xbit_r208_c48 bl[48] br[48] wl[208] vdd gnd cell_6t
Xbit_r209_c48 bl[48] br[48] wl[209] vdd gnd cell_6t
Xbit_r210_c48 bl[48] br[48] wl[210] vdd gnd cell_6t
Xbit_r211_c48 bl[48] br[48] wl[211] vdd gnd cell_6t
Xbit_r212_c48 bl[48] br[48] wl[212] vdd gnd cell_6t
Xbit_r213_c48 bl[48] br[48] wl[213] vdd gnd cell_6t
Xbit_r214_c48 bl[48] br[48] wl[214] vdd gnd cell_6t
Xbit_r215_c48 bl[48] br[48] wl[215] vdd gnd cell_6t
Xbit_r216_c48 bl[48] br[48] wl[216] vdd gnd cell_6t
Xbit_r217_c48 bl[48] br[48] wl[217] vdd gnd cell_6t
Xbit_r218_c48 bl[48] br[48] wl[218] vdd gnd cell_6t
Xbit_r219_c48 bl[48] br[48] wl[219] vdd gnd cell_6t
Xbit_r220_c48 bl[48] br[48] wl[220] vdd gnd cell_6t
Xbit_r221_c48 bl[48] br[48] wl[221] vdd gnd cell_6t
Xbit_r222_c48 bl[48] br[48] wl[222] vdd gnd cell_6t
Xbit_r223_c48 bl[48] br[48] wl[223] vdd gnd cell_6t
Xbit_r224_c48 bl[48] br[48] wl[224] vdd gnd cell_6t
Xbit_r225_c48 bl[48] br[48] wl[225] vdd gnd cell_6t
Xbit_r226_c48 bl[48] br[48] wl[226] vdd gnd cell_6t
Xbit_r227_c48 bl[48] br[48] wl[227] vdd gnd cell_6t
Xbit_r228_c48 bl[48] br[48] wl[228] vdd gnd cell_6t
Xbit_r229_c48 bl[48] br[48] wl[229] vdd gnd cell_6t
Xbit_r230_c48 bl[48] br[48] wl[230] vdd gnd cell_6t
Xbit_r231_c48 bl[48] br[48] wl[231] vdd gnd cell_6t
Xbit_r232_c48 bl[48] br[48] wl[232] vdd gnd cell_6t
Xbit_r233_c48 bl[48] br[48] wl[233] vdd gnd cell_6t
Xbit_r234_c48 bl[48] br[48] wl[234] vdd gnd cell_6t
Xbit_r235_c48 bl[48] br[48] wl[235] vdd gnd cell_6t
Xbit_r236_c48 bl[48] br[48] wl[236] vdd gnd cell_6t
Xbit_r237_c48 bl[48] br[48] wl[237] vdd gnd cell_6t
Xbit_r238_c48 bl[48] br[48] wl[238] vdd gnd cell_6t
Xbit_r239_c48 bl[48] br[48] wl[239] vdd gnd cell_6t
Xbit_r240_c48 bl[48] br[48] wl[240] vdd gnd cell_6t
Xbit_r241_c48 bl[48] br[48] wl[241] vdd gnd cell_6t
Xbit_r242_c48 bl[48] br[48] wl[242] vdd gnd cell_6t
Xbit_r243_c48 bl[48] br[48] wl[243] vdd gnd cell_6t
Xbit_r244_c48 bl[48] br[48] wl[244] vdd gnd cell_6t
Xbit_r245_c48 bl[48] br[48] wl[245] vdd gnd cell_6t
Xbit_r246_c48 bl[48] br[48] wl[246] vdd gnd cell_6t
Xbit_r247_c48 bl[48] br[48] wl[247] vdd gnd cell_6t
Xbit_r248_c48 bl[48] br[48] wl[248] vdd gnd cell_6t
Xbit_r249_c48 bl[48] br[48] wl[249] vdd gnd cell_6t
Xbit_r250_c48 bl[48] br[48] wl[250] vdd gnd cell_6t
Xbit_r251_c48 bl[48] br[48] wl[251] vdd gnd cell_6t
Xbit_r252_c48 bl[48] br[48] wl[252] vdd gnd cell_6t
Xbit_r253_c48 bl[48] br[48] wl[253] vdd gnd cell_6t
Xbit_r254_c48 bl[48] br[48] wl[254] vdd gnd cell_6t
Xbit_r255_c48 bl[48] br[48] wl[255] vdd gnd cell_6t
Xbit_r256_c48 bl[48] br[48] wl[256] vdd gnd cell_6t
Xbit_r257_c48 bl[48] br[48] wl[257] vdd gnd cell_6t
Xbit_r258_c48 bl[48] br[48] wl[258] vdd gnd cell_6t
Xbit_r259_c48 bl[48] br[48] wl[259] vdd gnd cell_6t
Xbit_r260_c48 bl[48] br[48] wl[260] vdd gnd cell_6t
Xbit_r261_c48 bl[48] br[48] wl[261] vdd gnd cell_6t
Xbit_r262_c48 bl[48] br[48] wl[262] vdd gnd cell_6t
Xbit_r263_c48 bl[48] br[48] wl[263] vdd gnd cell_6t
Xbit_r264_c48 bl[48] br[48] wl[264] vdd gnd cell_6t
Xbit_r265_c48 bl[48] br[48] wl[265] vdd gnd cell_6t
Xbit_r266_c48 bl[48] br[48] wl[266] vdd gnd cell_6t
Xbit_r267_c48 bl[48] br[48] wl[267] vdd gnd cell_6t
Xbit_r268_c48 bl[48] br[48] wl[268] vdd gnd cell_6t
Xbit_r269_c48 bl[48] br[48] wl[269] vdd gnd cell_6t
Xbit_r270_c48 bl[48] br[48] wl[270] vdd gnd cell_6t
Xbit_r271_c48 bl[48] br[48] wl[271] vdd gnd cell_6t
Xbit_r272_c48 bl[48] br[48] wl[272] vdd gnd cell_6t
Xbit_r273_c48 bl[48] br[48] wl[273] vdd gnd cell_6t
Xbit_r274_c48 bl[48] br[48] wl[274] vdd gnd cell_6t
Xbit_r275_c48 bl[48] br[48] wl[275] vdd gnd cell_6t
Xbit_r276_c48 bl[48] br[48] wl[276] vdd gnd cell_6t
Xbit_r277_c48 bl[48] br[48] wl[277] vdd gnd cell_6t
Xbit_r278_c48 bl[48] br[48] wl[278] vdd gnd cell_6t
Xbit_r279_c48 bl[48] br[48] wl[279] vdd gnd cell_6t
Xbit_r280_c48 bl[48] br[48] wl[280] vdd gnd cell_6t
Xbit_r281_c48 bl[48] br[48] wl[281] vdd gnd cell_6t
Xbit_r282_c48 bl[48] br[48] wl[282] vdd gnd cell_6t
Xbit_r283_c48 bl[48] br[48] wl[283] vdd gnd cell_6t
Xbit_r284_c48 bl[48] br[48] wl[284] vdd gnd cell_6t
Xbit_r285_c48 bl[48] br[48] wl[285] vdd gnd cell_6t
Xbit_r286_c48 bl[48] br[48] wl[286] vdd gnd cell_6t
Xbit_r287_c48 bl[48] br[48] wl[287] vdd gnd cell_6t
Xbit_r288_c48 bl[48] br[48] wl[288] vdd gnd cell_6t
Xbit_r289_c48 bl[48] br[48] wl[289] vdd gnd cell_6t
Xbit_r290_c48 bl[48] br[48] wl[290] vdd gnd cell_6t
Xbit_r291_c48 bl[48] br[48] wl[291] vdd gnd cell_6t
Xbit_r292_c48 bl[48] br[48] wl[292] vdd gnd cell_6t
Xbit_r293_c48 bl[48] br[48] wl[293] vdd gnd cell_6t
Xbit_r294_c48 bl[48] br[48] wl[294] vdd gnd cell_6t
Xbit_r295_c48 bl[48] br[48] wl[295] vdd gnd cell_6t
Xbit_r296_c48 bl[48] br[48] wl[296] vdd gnd cell_6t
Xbit_r297_c48 bl[48] br[48] wl[297] vdd gnd cell_6t
Xbit_r298_c48 bl[48] br[48] wl[298] vdd gnd cell_6t
Xbit_r299_c48 bl[48] br[48] wl[299] vdd gnd cell_6t
Xbit_r300_c48 bl[48] br[48] wl[300] vdd gnd cell_6t
Xbit_r301_c48 bl[48] br[48] wl[301] vdd gnd cell_6t
Xbit_r302_c48 bl[48] br[48] wl[302] vdd gnd cell_6t
Xbit_r303_c48 bl[48] br[48] wl[303] vdd gnd cell_6t
Xbit_r304_c48 bl[48] br[48] wl[304] vdd gnd cell_6t
Xbit_r305_c48 bl[48] br[48] wl[305] vdd gnd cell_6t
Xbit_r306_c48 bl[48] br[48] wl[306] vdd gnd cell_6t
Xbit_r307_c48 bl[48] br[48] wl[307] vdd gnd cell_6t
Xbit_r308_c48 bl[48] br[48] wl[308] vdd gnd cell_6t
Xbit_r309_c48 bl[48] br[48] wl[309] vdd gnd cell_6t
Xbit_r310_c48 bl[48] br[48] wl[310] vdd gnd cell_6t
Xbit_r311_c48 bl[48] br[48] wl[311] vdd gnd cell_6t
Xbit_r312_c48 bl[48] br[48] wl[312] vdd gnd cell_6t
Xbit_r313_c48 bl[48] br[48] wl[313] vdd gnd cell_6t
Xbit_r314_c48 bl[48] br[48] wl[314] vdd gnd cell_6t
Xbit_r315_c48 bl[48] br[48] wl[315] vdd gnd cell_6t
Xbit_r316_c48 bl[48] br[48] wl[316] vdd gnd cell_6t
Xbit_r317_c48 bl[48] br[48] wl[317] vdd gnd cell_6t
Xbit_r318_c48 bl[48] br[48] wl[318] vdd gnd cell_6t
Xbit_r319_c48 bl[48] br[48] wl[319] vdd gnd cell_6t
Xbit_r320_c48 bl[48] br[48] wl[320] vdd gnd cell_6t
Xbit_r321_c48 bl[48] br[48] wl[321] vdd gnd cell_6t
Xbit_r322_c48 bl[48] br[48] wl[322] vdd gnd cell_6t
Xbit_r323_c48 bl[48] br[48] wl[323] vdd gnd cell_6t
Xbit_r324_c48 bl[48] br[48] wl[324] vdd gnd cell_6t
Xbit_r325_c48 bl[48] br[48] wl[325] vdd gnd cell_6t
Xbit_r326_c48 bl[48] br[48] wl[326] vdd gnd cell_6t
Xbit_r327_c48 bl[48] br[48] wl[327] vdd gnd cell_6t
Xbit_r328_c48 bl[48] br[48] wl[328] vdd gnd cell_6t
Xbit_r329_c48 bl[48] br[48] wl[329] vdd gnd cell_6t
Xbit_r330_c48 bl[48] br[48] wl[330] vdd gnd cell_6t
Xbit_r331_c48 bl[48] br[48] wl[331] vdd gnd cell_6t
Xbit_r332_c48 bl[48] br[48] wl[332] vdd gnd cell_6t
Xbit_r333_c48 bl[48] br[48] wl[333] vdd gnd cell_6t
Xbit_r334_c48 bl[48] br[48] wl[334] vdd gnd cell_6t
Xbit_r335_c48 bl[48] br[48] wl[335] vdd gnd cell_6t
Xbit_r336_c48 bl[48] br[48] wl[336] vdd gnd cell_6t
Xbit_r337_c48 bl[48] br[48] wl[337] vdd gnd cell_6t
Xbit_r338_c48 bl[48] br[48] wl[338] vdd gnd cell_6t
Xbit_r339_c48 bl[48] br[48] wl[339] vdd gnd cell_6t
Xbit_r340_c48 bl[48] br[48] wl[340] vdd gnd cell_6t
Xbit_r341_c48 bl[48] br[48] wl[341] vdd gnd cell_6t
Xbit_r342_c48 bl[48] br[48] wl[342] vdd gnd cell_6t
Xbit_r343_c48 bl[48] br[48] wl[343] vdd gnd cell_6t
Xbit_r344_c48 bl[48] br[48] wl[344] vdd gnd cell_6t
Xbit_r345_c48 bl[48] br[48] wl[345] vdd gnd cell_6t
Xbit_r346_c48 bl[48] br[48] wl[346] vdd gnd cell_6t
Xbit_r347_c48 bl[48] br[48] wl[347] vdd gnd cell_6t
Xbit_r348_c48 bl[48] br[48] wl[348] vdd gnd cell_6t
Xbit_r349_c48 bl[48] br[48] wl[349] vdd gnd cell_6t
Xbit_r350_c48 bl[48] br[48] wl[350] vdd gnd cell_6t
Xbit_r351_c48 bl[48] br[48] wl[351] vdd gnd cell_6t
Xbit_r352_c48 bl[48] br[48] wl[352] vdd gnd cell_6t
Xbit_r353_c48 bl[48] br[48] wl[353] vdd gnd cell_6t
Xbit_r354_c48 bl[48] br[48] wl[354] vdd gnd cell_6t
Xbit_r355_c48 bl[48] br[48] wl[355] vdd gnd cell_6t
Xbit_r356_c48 bl[48] br[48] wl[356] vdd gnd cell_6t
Xbit_r357_c48 bl[48] br[48] wl[357] vdd gnd cell_6t
Xbit_r358_c48 bl[48] br[48] wl[358] vdd gnd cell_6t
Xbit_r359_c48 bl[48] br[48] wl[359] vdd gnd cell_6t
Xbit_r360_c48 bl[48] br[48] wl[360] vdd gnd cell_6t
Xbit_r361_c48 bl[48] br[48] wl[361] vdd gnd cell_6t
Xbit_r362_c48 bl[48] br[48] wl[362] vdd gnd cell_6t
Xbit_r363_c48 bl[48] br[48] wl[363] vdd gnd cell_6t
Xbit_r364_c48 bl[48] br[48] wl[364] vdd gnd cell_6t
Xbit_r365_c48 bl[48] br[48] wl[365] vdd gnd cell_6t
Xbit_r366_c48 bl[48] br[48] wl[366] vdd gnd cell_6t
Xbit_r367_c48 bl[48] br[48] wl[367] vdd gnd cell_6t
Xbit_r368_c48 bl[48] br[48] wl[368] vdd gnd cell_6t
Xbit_r369_c48 bl[48] br[48] wl[369] vdd gnd cell_6t
Xbit_r370_c48 bl[48] br[48] wl[370] vdd gnd cell_6t
Xbit_r371_c48 bl[48] br[48] wl[371] vdd gnd cell_6t
Xbit_r372_c48 bl[48] br[48] wl[372] vdd gnd cell_6t
Xbit_r373_c48 bl[48] br[48] wl[373] vdd gnd cell_6t
Xbit_r374_c48 bl[48] br[48] wl[374] vdd gnd cell_6t
Xbit_r375_c48 bl[48] br[48] wl[375] vdd gnd cell_6t
Xbit_r376_c48 bl[48] br[48] wl[376] vdd gnd cell_6t
Xbit_r377_c48 bl[48] br[48] wl[377] vdd gnd cell_6t
Xbit_r378_c48 bl[48] br[48] wl[378] vdd gnd cell_6t
Xbit_r379_c48 bl[48] br[48] wl[379] vdd gnd cell_6t
Xbit_r380_c48 bl[48] br[48] wl[380] vdd gnd cell_6t
Xbit_r381_c48 bl[48] br[48] wl[381] vdd gnd cell_6t
Xbit_r382_c48 bl[48] br[48] wl[382] vdd gnd cell_6t
Xbit_r383_c48 bl[48] br[48] wl[383] vdd gnd cell_6t
Xbit_r384_c48 bl[48] br[48] wl[384] vdd gnd cell_6t
Xbit_r385_c48 bl[48] br[48] wl[385] vdd gnd cell_6t
Xbit_r386_c48 bl[48] br[48] wl[386] vdd gnd cell_6t
Xbit_r387_c48 bl[48] br[48] wl[387] vdd gnd cell_6t
Xbit_r388_c48 bl[48] br[48] wl[388] vdd gnd cell_6t
Xbit_r389_c48 bl[48] br[48] wl[389] vdd gnd cell_6t
Xbit_r390_c48 bl[48] br[48] wl[390] vdd gnd cell_6t
Xbit_r391_c48 bl[48] br[48] wl[391] vdd gnd cell_6t
Xbit_r392_c48 bl[48] br[48] wl[392] vdd gnd cell_6t
Xbit_r393_c48 bl[48] br[48] wl[393] vdd gnd cell_6t
Xbit_r394_c48 bl[48] br[48] wl[394] vdd gnd cell_6t
Xbit_r395_c48 bl[48] br[48] wl[395] vdd gnd cell_6t
Xbit_r396_c48 bl[48] br[48] wl[396] vdd gnd cell_6t
Xbit_r397_c48 bl[48] br[48] wl[397] vdd gnd cell_6t
Xbit_r398_c48 bl[48] br[48] wl[398] vdd gnd cell_6t
Xbit_r399_c48 bl[48] br[48] wl[399] vdd gnd cell_6t
Xbit_r400_c48 bl[48] br[48] wl[400] vdd gnd cell_6t
Xbit_r401_c48 bl[48] br[48] wl[401] vdd gnd cell_6t
Xbit_r402_c48 bl[48] br[48] wl[402] vdd gnd cell_6t
Xbit_r403_c48 bl[48] br[48] wl[403] vdd gnd cell_6t
Xbit_r404_c48 bl[48] br[48] wl[404] vdd gnd cell_6t
Xbit_r405_c48 bl[48] br[48] wl[405] vdd gnd cell_6t
Xbit_r406_c48 bl[48] br[48] wl[406] vdd gnd cell_6t
Xbit_r407_c48 bl[48] br[48] wl[407] vdd gnd cell_6t
Xbit_r408_c48 bl[48] br[48] wl[408] vdd gnd cell_6t
Xbit_r409_c48 bl[48] br[48] wl[409] vdd gnd cell_6t
Xbit_r410_c48 bl[48] br[48] wl[410] vdd gnd cell_6t
Xbit_r411_c48 bl[48] br[48] wl[411] vdd gnd cell_6t
Xbit_r412_c48 bl[48] br[48] wl[412] vdd gnd cell_6t
Xbit_r413_c48 bl[48] br[48] wl[413] vdd gnd cell_6t
Xbit_r414_c48 bl[48] br[48] wl[414] vdd gnd cell_6t
Xbit_r415_c48 bl[48] br[48] wl[415] vdd gnd cell_6t
Xbit_r416_c48 bl[48] br[48] wl[416] vdd gnd cell_6t
Xbit_r417_c48 bl[48] br[48] wl[417] vdd gnd cell_6t
Xbit_r418_c48 bl[48] br[48] wl[418] vdd gnd cell_6t
Xbit_r419_c48 bl[48] br[48] wl[419] vdd gnd cell_6t
Xbit_r420_c48 bl[48] br[48] wl[420] vdd gnd cell_6t
Xbit_r421_c48 bl[48] br[48] wl[421] vdd gnd cell_6t
Xbit_r422_c48 bl[48] br[48] wl[422] vdd gnd cell_6t
Xbit_r423_c48 bl[48] br[48] wl[423] vdd gnd cell_6t
Xbit_r424_c48 bl[48] br[48] wl[424] vdd gnd cell_6t
Xbit_r425_c48 bl[48] br[48] wl[425] vdd gnd cell_6t
Xbit_r426_c48 bl[48] br[48] wl[426] vdd gnd cell_6t
Xbit_r427_c48 bl[48] br[48] wl[427] vdd gnd cell_6t
Xbit_r428_c48 bl[48] br[48] wl[428] vdd gnd cell_6t
Xbit_r429_c48 bl[48] br[48] wl[429] vdd gnd cell_6t
Xbit_r430_c48 bl[48] br[48] wl[430] vdd gnd cell_6t
Xbit_r431_c48 bl[48] br[48] wl[431] vdd gnd cell_6t
Xbit_r432_c48 bl[48] br[48] wl[432] vdd gnd cell_6t
Xbit_r433_c48 bl[48] br[48] wl[433] vdd gnd cell_6t
Xbit_r434_c48 bl[48] br[48] wl[434] vdd gnd cell_6t
Xbit_r435_c48 bl[48] br[48] wl[435] vdd gnd cell_6t
Xbit_r436_c48 bl[48] br[48] wl[436] vdd gnd cell_6t
Xbit_r437_c48 bl[48] br[48] wl[437] vdd gnd cell_6t
Xbit_r438_c48 bl[48] br[48] wl[438] vdd gnd cell_6t
Xbit_r439_c48 bl[48] br[48] wl[439] vdd gnd cell_6t
Xbit_r440_c48 bl[48] br[48] wl[440] vdd gnd cell_6t
Xbit_r441_c48 bl[48] br[48] wl[441] vdd gnd cell_6t
Xbit_r442_c48 bl[48] br[48] wl[442] vdd gnd cell_6t
Xbit_r443_c48 bl[48] br[48] wl[443] vdd gnd cell_6t
Xbit_r444_c48 bl[48] br[48] wl[444] vdd gnd cell_6t
Xbit_r445_c48 bl[48] br[48] wl[445] vdd gnd cell_6t
Xbit_r446_c48 bl[48] br[48] wl[446] vdd gnd cell_6t
Xbit_r447_c48 bl[48] br[48] wl[447] vdd gnd cell_6t
Xbit_r448_c48 bl[48] br[48] wl[448] vdd gnd cell_6t
Xbit_r449_c48 bl[48] br[48] wl[449] vdd gnd cell_6t
Xbit_r450_c48 bl[48] br[48] wl[450] vdd gnd cell_6t
Xbit_r451_c48 bl[48] br[48] wl[451] vdd gnd cell_6t
Xbit_r452_c48 bl[48] br[48] wl[452] vdd gnd cell_6t
Xbit_r453_c48 bl[48] br[48] wl[453] vdd gnd cell_6t
Xbit_r454_c48 bl[48] br[48] wl[454] vdd gnd cell_6t
Xbit_r455_c48 bl[48] br[48] wl[455] vdd gnd cell_6t
Xbit_r456_c48 bl[48] br[48] wl[456] vdd gnd cell_6t
Xbit_r457_c48 bl[48] br[48] wl[457] vdd gnd cell_6t
Xbit_r458_c48 bl[48] br[48] wl[458] vdd gnd cell_6t
Xbit_r459_c48 bl[48] br[48] wl[459] vdd gnd cell_6t
Xbit_r460_c48 bl[48] br[48] wl[460] vdd gnd cell_6t
Xbit_r461_c48 bl[48] br[48] wl[461] vdd gnd cell_6t
Xbit_r462_c48 bl[48] br[48] wl[462] vdd gnd cell_6t
Xbit_r463_c48 bl[48] br[48] wl[463] vdd gnd cell_6t
Xbit_r464_c48 bl[48] br[48] wl[464] vdd gnd cell_6t
Xbit_r465_c48 bl[48] br[48] wl[465] vdd gnd cell_6t
Xbit_r466_c48 bl[48] br[48] wl[466] vdd gnd cell_6t
Xbit_r467_c48 bl[48] br[48] wl[467] vdd gnd cell_6t
Xbit_r468_c48 bl[48] br[48] wl[468] vdd gnd cell_6t
Xbit_r469_c48 bl[48] br[48] wl[469] vdd gnd cell_6t
Xbit_r470_c48 bl[48] br[48] wl[470] vdd gnd cell_6t
Xbit_r471_c48 bl[48] br[48] wl[471] vdd gnd cell_6t
Xbit_r472_c48 bl[48] br[48] wl[472] vdd gnd cell_6t
Xbit_r473_c48 bl[48] br[48] wl[473] vdd gnd cell_6t
Xbit_r474_c48 bl[48] br[48] wl[474] vdd gnd cell_6t
Xbit_r475_c48 bl[48] br[48] wl[475] vdd gnd cell_6t
Xbit_r476_c48 bl[48] br[48] wl[476] vdd gnd cell_6t
Xbit_r477_c48 bl[48] br[48] wl[477] vdd gnd cell_6t
Xbit_r478_c48 bl[48] br[48] wl[478] vdd gnd cell_6t
Xbit_r479_c48 bl[48] br[48] wl[479] vdd gnd cell_6t
Xbit_r480_c48 bl[48] br[48] wl[480] vdd gnd cell_6t
Xbit_r481_c48 bl[48] br[48] wl[481] vdd gnd cell_6t
Xbit_r482_c48 bl[48] br[48] wl[482] vdd gnd cell_6t
Xbit_r483_c48 bl[48] br[48] wl[483] vdd gnd cell_6t
Xbit_r484_c48 bl[48] br[48] wl[484] vdd gnd cell_6t
Xbit_r485_c48 bl[48] br[48] wl[485] vdd gnd cell_6t
Xbit_r486_c48 bl[48] br[48] wl[486] vdd gnd cell_6t
Xbit_r487_c48 bl[48] br[48] wl[487] vdd gnd cell_6t
Xbit_r488_c48 bl[48] br[48] wl[488] vdd gnd cell_6t
Xbit_r489_c48 bl[48] br[48] wl[489] vdd gnd cell_6t
Xbit_r490_c48 bl[48] br[48] wl[490] vdd gnd cell_6t
Xbit_r491_c48 bl[48] br[48] wl[491] vdd gnd cell_6t
Xbit_r492_c48 bl[48] br[48] wl[492] vdd gnd cell_6t
Xbit_r493_c48 bl[48] br[48] wl[493] vdd gnd cell_6t
Xbit_r494_c48 bl[48] br[48] wl[494] vdd gnd cell_6t
Xbit_r495_c48 bl[48] br[48] wl[495] vdd gnd cell_6t
Xbit_r496_c48 bl[48] br[48] wl[496] vdd gnd cell_6t
Xbit_r497_c48 bl[48] br[48] wl[497] vdd gnd cell_6t
Xbit_r498_c48 bl[48] br[48] wl[498] vdd gnd cell_6t
Xbit_r499_c48 bl[48] br[48] wl[499] vdd gnd cell_6t
Xbit_r500_c48 bl[48] br[48] wl[500] vdd gnd cell_6t
Xbit_r501_c48 bl[48] br[48] wl[501] vdd gnd cell_6t
Xbit_r502_c48 bl[48] br[48] wl[502] vdd gnd cell_6t
Xbit_r503_c48 bl[48] br[48] wl[503] vdd gnd cell_6t
Xbit_r504_c48 bl[48] br[48] wl[504] vdd gnd cell_6t
Xbit_r505_c48 bl[48] br[48] wl[505] vdd gnd cell_6t
Xbit_r506_c48 bl[48] br[48] wl[506] vdd gnd cell_6t
Xbit_r507_c48 bl[48] br[48] wl[507] vdd gnd cell_6t
Xbit_r508_c48 bl[48] br[48] wl[508] vdd gnd cell_6t
Xbit_r509_c48 bl[48] br[48] wl[509] vdd gnd cell_6t
Xbit_r510_c48 bl[48] br[48] wl[510] vdd gnd cell_6t
Xbit_r511_c48 bl[48] br[48] wl[511] vdd gnd cell_6t
Xbit_r0_c49 bl[49] br[49] wl[0] vdd gnd cell_6t
Xbit_r1_c49 bl[49] br[49] wl[1] vdd gnd cell_6t
Xbit_r2_c49 bl[49] br[49] wl[2] vdd gnd cell_6t
Xbit_r3_c49 bl[49] br[49] wl[3] vdd gnd cell_6t
Xbit_r4_c49 bl[49] br[49] wl[4] vdd gnd cell_6t
Xbit_r5_c49 bl[49] br[49] wl[5] vdd gnd cell_6t
Xbit_r6_c49 bl[49] br[49] wl[6] vdd gnd cell_6t
Xbit_r7_c49 bl[49] br[49] wl[7] vdd gnd cell_6t
Xbit_r8_c49 bl[49] br[49] wl[8] vdd gnd cell_6t
Xbit_r9_c49 bl[49] br[49] wl[9] vdd gnd cell_6t
Xbit_r10_c49 bl[49] br[49] wl[10] vdd gnd cell_6t
Xbit_r11_c49 bl[49] br[49] wl[11] vdd gnd cell_6t
Xbit_r12_c49 bl[49] br[49] wl[12] vdd gnd cell_6t
Xbit_r13_c49 bl[49] br[49] wl[13] vdd gnd cell_6t
Xbit_r14_c49 bl[49] br[49] wl[14] vdd gnd cell_6t
Xbit_r15_c49 bl[49] br[49] wl[15] vdd gnd cell_6t
Xbit_r16_c49 bl[49] br[49] wl[16] vdd gnd cell_6t
Xbit_r17_c49 bl[49] br[49] wl[17] vdd gnd cell_6t
Xbit_r18_c49 bl[49] br[49] wl[18] vdd gnd cell_6t
Xbit_r19_c49 bl[49] br[49] wl[19] vdd gnd cell_6t
Xbit_r20_c49 bl[49] br[49] wl[20] vdd gnd cell_6t
Xbit_r21_c49 bl[49] br[49] wl[21] vdd gnd cell_6t
Xbit_r22_c49 bl[49] br[49] wl[22] vdd gnd cell_6t
Xbit_r23_c49 bl[49] br[49] wl[23] vdd gnd cell_6t
Xbit_r24_c49 bl[49] br[49] wl[24] vdd gnd cell_6t
Xbit_r25_c49 bl[49] br[49] wl[25] vdd gnd cell_6t
Xbit_r26_c49 bl[49] br[49] wl[26] vdd gnd cell_6t
Xbit_r27_c49 bl[49] br[49] wl[27] vdd gnd cell_6t
Xbit_r28_c49 bl[49] br[49] wl[28] vdd gnd cell_6t
Xbit_r29_c49 bl[49] br[49] wl[29] vdd gnd cell_6t
Xbit_r30_c49 bl[49] br[49] wl[30] vdd gnd cell_6t
Xbit_r31_c49 bl[49] br[49] wl[31] vdd gnd cell_6t
Xbit_r32_c49 bl[49] br[49] wl[32] vdd gnd cell_6t
Xbit_r33_c49 bl[49] br[49] wl[33] vdd gnd cell_6t
Xbit_r34_c49 bl[49] br[49] wl[34] vdd gnd cell_6t
Xbit_r35_c49 bl[49] br[49] wl[35] vdd gnd cell_6t
Xbit_r36_c49 bl[49] br[49] wl[36] vdd gnd cell_6t
Xbit_r37_c49 bl[49] br[49] wl[37] vdd gnd cell_6t
Xbit_r38_c49 bl[49] br[49] wl[38] vdd gnd cell_6t
Xbit_r39_c49 bl[49] br[49] wl[39] vdd gnd cell_6t
Xbit_r40_c49 bl[49] br[49] wl[40] vdd gnd cell_6t
Xbit_r41_c49 bl[49] br[49] wl[41] vdd gnd cell_6t
Xbit_r42_c49 bl[49] br[49] wl[42] vdd gnd cell_6t
Xbit_r43_c49 bl[49] br[49] wl[43] vdd gnd cell_6t
Xbit_r44_c49 bl[49] br[49] wl[44] vdd gnd cell_6t
Xbit_r45_c49 bl[49] br[49] wl[45] vdd gnd cell_6t
Xbit_r46_c49 bl[49] br[49] wl[46] vdd gnd cell_6t
Xbit_r47_c49 bl[49] br[49] wl[47] vdd gnd cell_6t
Xbit_r48_c49 bl[49] br[49] wl[48] vdd gnd cell_6t
Xbit_r49_c49 bl[49] br[49] wl[49] vdd gnd cell_6t
Xbit_r50_c49 bl[49] br[49] wl[50] vdd gnd cell_6t
Xbit_r51_c49 bl[49] br[49] wl[51] vdd gnd cell_6t
Xbit_r52_c49 bl[49] br[49] wl[52] vdd gnd cell_6t
Xbit_r53_c49 bl[49] br[49] wl[53] vdd gnd cell_6t
Xbit_r54_c49 bl[49] br[49] wl[54] vdd gnd cell_6t
Xbit_r55_c49 bl[49] br[49] wl[55] vdd gnd cell_6t
Xbit_r56_c49 bl[49] br[49] wl[56] vdd gnd cell_6t
Xbit_r57_c49 bl[49] br[49] wl[57] vdd gnd cell_6t
Xbit_r58_c49 bl[49] br[49] wl[58] vdd gnd cell_6t
Xbit_r59_c49 bl[49] br[49] wl[59] vdd gnd cell_6t
Xbit_r60_c49 bl[49] br[49] wl[60] vdd gnd cell_6t
Xbit_r61_c49 bl[49] br[49] wl[61] vdd gnd cell_6t
Xbit_r62_c49 bl[49] br[49] wl[62] vdd gnd cell_6t
Xbit_r63_c49 bl[49] br[49] wl[63] vdd gnd cell_6t
Xbit_r64_c49 bl[49] br[49] wl[64] vdd gnd cell_6t
Xbit_r65_c49 bl[49] br[49] wl[65] vdd gnd cell_6t
Xbit_r66_c49 bl[49] br[49] wl[66] vdd gnd cell_6t
Xbit_r67_c49 bl[49] br[49] wl[67] vdd gnd cell_6t
Xbit_r68_c49 bl[49] br[49] wl[68] vdd gnd cell_6t
Xbit_r69_c49 bl[49] br[49] wl[69] vdd gnd cell_6t
Xbit_r70_c49 bl[49] br[49] wl[70] vdd gnd cell_6t
Xbit_r71_c49 bl[49] br[49] wl[71] vdd gnd cell_6t
Xbit_r72_c49 bl[49] br[49] wl[72] vdd gnd cell_6t
Xbit_r73_c49 bl[49] br[49] wl[73] vdd gnd cell_6t
Xbit_r74_c49 bl[49] br[49] wl[74] vdd gnd cell_6t
Xbit_r75_c49 bl[49] br[49] wl[75] vdd gnd cell_6t
Xbit_r76_c49 bl[49] br[49] wl[76] vdd gnd cell_6t
Xbit_r77_c49 bl[49] br[49] wl[77] vdd gnd cell_6t
Xbit_r78_c49 bl[49] br[49] wl[78] vdd gnd cell_6t
Xbit_r79_c49 bl[49] br[49] wl[79] vdd gnd cell_6t
Xbit_r80_c49 bl[49] br[49] wl[80] vdd gnd cell_6t
Xbit_r81_c49 bl[49] br[49] wl[81] vdd gnd cell_6t
Xbit_r82_c49 bl[49] br[49] wl[82] vdd gnd cell_6t
Xbit_r83_c49 bl[49] br[49] wl[83] vdd gnd cell_6t
Xbit_r84_c49 bl[49] br[49] wl[84] vdd gnd cell_6t
Xbit_r85_c49 bl[49] br[49] wl[85] vdd gnd cell_6t
Xbit_r86_c49 bl[49] br[49] wl[86] vdd gnd cell_6t
Xbit_r87_c49 bl[49] br[49] wl[87] vdd gnd cell_6t
Xbit_r88_c49 bl[49] br[49] wl[88] vdd gnd cell_6t
Xbit_r89_c49 bl[49] br[49] wl[89] vdd gnd cell_6t
Xbit_r90_c49 bl[49] br[49] wl[90] vdd gnd cell_6t
Xbit_r91_c49 bl[49] br[49] wl[91] vdd gnd cell_6t
Xbit_r92_c49 bl[49] br[49] wl[92] vdd gnd cell_6t
Xbit_r93_c49 bl[49] br[49] wl[93] vdd gnd cell_6t
Xbit_r94_c49 bl[49] br[49] wl[94] vdd gnd cell_6t
Xbit_r95_c49 bl[49] br[49] wl[95] vdd gnd cell_6t
Xbit_r96_c49 bl[49] br[49] wl[96] vdd gnd cell_6t
Xbit_r97_c49 bl[49] br[49] wl[97] vdd gnd cell_6t
Xbit_r98_c49 bl[49] br[49] wl[98] vdd gnd cell_6t
Xbit_r99_c49 bl[49] br[49] wl[99] vdd gnd cell_6t
Xbit_r100_c49 bl[49] br[49] wl[100] vdd gnd cell_6t
Xbit_r101_c49 bl[49] br[49] wl[101] vdd gnd cell_6t
Xbit_r102_c49 bl[49] br[49] wl[102] vdd gnd cell_6t
Xbit_r103_c49 bl[49] br[49] wl[103] vdd gnd cell_6t
Xbit_r104_c49 bl[49] br[49] wl[104] vdd gnd cell_6t
Xbit_r105_c49 bl[49] br[49] wl[105] vdd gnd cell_6t
Xbit_r106_c49 bl[49] br[49] wl[106] vdd gnd cell_6t
Xbit_r107_c49 bl[49] br[49] wl[107] vdd gnd cell_6t
Xbit_r108_c49 bl[49] br[49] wl[108] vdd gnd cell_6t
Xbit_r109_c49 bl[49] br[49] wl[109] vdd gnd cell_6t
Xbit_r110_c49 bl[49] br[49] wl[110] vdd gnd cell_6t
Xbit_r111_c49 bl[49] br[49] wl[111] vdd gnd cell_6t
Xbit_r112_c49 bl[49] br[49] wl[112] vdd gnd cell_6t
Xbit_r113_c49 bl[49] br[49] wl[113] vdd gnd cell_6t
Xbit_r114_c49 bl[49] br[49] wl[114] vdd gnd cell_6t
Xbit_r115_c49 bl[49] br[49] wl[115] vdd gnd cell_6t
Xbit_r116_c49 bl[49] br[49] wl[116] vdd gnd cell_6t
Xbit_r117_c49 bl[49] br[49] wl[117] vdd gnd cell_6t
Xbit_r118_c49 bl[49] br[49] wl[118] vdd gnd cell_6t
Xbit_r119_c49 bl[49] br[49] wl[119] vdd gnd cell_6t
Xbit_r120_c49 bl[49] br[49] wl[120] vdd gnd cell_6t
Xbit_r121_c49 bl[49] br[49] wl[121] vdd gnd cell_6t
Xbit_r122_c49 bl[49] br[49] wl[122] vdd gnd cell_6t
Xbit_r123_c49 bl[49] br[49] wl[123] vdd gnd cell_6t
Xbit_r124_c49 bl[49] br[49] wl[124] vdd gnd cell_6t
Xbit_r125_c49 bl[49] br[49] wl[125] vdd gnd cell_6t
Xbit_r126_c49 bl[49] br[49] wl[126] vdd gnd cell_6t
Xbit_r127_c49 bl[49] br[49] wl[127] vdd gnd cell_6t
Xbit_r128_c49 bl[49] br[49] wl[128] vdd gnd cell_6t
Xbit_r129_c49 bl[49] br[49] wl[129] vdd gnd cell_6t
Xbit_r130_c49 bl[49] br[49] wl[130] vdd gnd cell_6t
Xbit_r131_c49 bl[49] br[49] wl[131] vdd gnd cell_6t
Xbit_r132_c49 bl[49] br[49] wl[132] vdd gnd cell_6t
Xbit_r133_c49 bl[49] br[49] wl[133] vdd gnd cell_6t
Xbit_r134_c49 bl[49] br[49] wl[134] vdd gnd cell_6t
Xbit_r135_c49 bl[49] br[49] wl[135] vdd gnd cell_6t
Xbit_r136_c49 bl[49] br[49] wl[136] vdd gnd cell_6t
Xbit_r137_c49 bl[49] br[49] wl[137] vdd gnd cell_6t
Xbit_r138_c49 bl[49] br[49] wl[138] vdd gnd cell_6t
Xbit_r139_c49 bl[49] br[49] wl[139] vdd gnd cell_6t
Xbit_r140_c49 bl[49] br[49] wl[140] vdd gnd cell_6t
Xbit_r141_c49 bl[49] br[49] wl[141] vdd gnd cell_6t
Xbit_r142_c49 bl[49] br[49] wl[142] vdd gnd cell_6t
Xbit_r143_c49 bl[49] br[49] wl[143] vdd gnd cell_6t
Xbit_r144_c49 bl[49] br[49] wl[144] vdd gnd cell_6t
Xbit_r145_c49 bl[49] br[49] wl[145] vdd gnd cell_6t
Xbit_r146_c49 bl[49] br[49] wl[146] vdd gnd cell_6t
Xbit_r147_c49 bl[49] br[49] wl[147] vdd gnd cell_6t
Xbit_r148_c49 bl[49] br[49] wl[148] vdd gnd cell_6t
Xbit_r149_c49 bl[49] br[49] wl[149] vdd gnd cell_6t
Xbit_r150_c49 bl[49] br[49] wl[150] vdd gnd cell_6t
Xbit_r151_c49 bl[49] br[49] wl[151] vdd gnd cell_6t
Xbit_r152_c49 bl[49] br[49] wl[152] vdd gnd cell_6t
Xbit_r153_c49 bl[49] br[49] wl[153] vdd gnd cell_6t
Xbit_r154_c49 bl[49] br[49] wl[154] vdd gnd cell_6t
Xbit_r155_c49 bl[49] br[49] wl[155] vdd gnd cell_6t
Xbit_r156_c49 bl[49] br[49] wl[156] vdd gnd cell_6t
Xbit_r157_c49 bl[49] br[49] wl[157] vdd gnd cell_6t
Xbit_r158_c49 bl[49] br[49] wl[158] vdd gnd cell_6t
Xbit_r159_c49 bl[49] br[49] wl[159] vdd gnd cell_6t
Xbit_r160_c49 bl[49] br[49] wl[160] vdd gnd cell_6t
Xbit_r161_c49 bl[49] br[49] wl[161] vdd gnd cell_6t
Xbit_r162_c49 bl[49] br[49] wl[162] vdd gnd cell_6t
Xbit_r163_c49 bl[49] br[49] wl[163] vdd gnd cell_6t
Xbit_r164_c49 bl[49] br[49] wl[164] vdd gnd cell_6t
Xbit_r165_c49 bl[49] br[49] wl[165] vdd gnd cell_6t
Xbit_r166_c49 bl[49] br[49] wl[166] vdd gnd cell_6t
Xbit_r167_c49 bl[49] br[49] wl[167] vdd gnd cell_6t
Xbit_r168_c49 bl[49] br[49] wl[168] vdd gnd cell_6t
Xbit_r169_c49 bl[49] br[49] wl[169] vdd gnd cell_6t
Xbit_r170_c49 bl[49] br[49] wl[170] vdd gnd cell_6t
Xbit_r171_c49 bl[49] br[49] wl[171] vdd gnd cell_6t
Xbit_r172_c49 bl[49] br[49] wl[172] vdd gnd cell_6t
Xbit_r173_c49 bl[49] br[49] wl[173] vdd gnd cell_6t
Xbit_r174_c49 bl[49] br[49] wl[174] vdd gnd cell_6t
Xbit_r175_c49 bl[49] br[49] wl[175] vdd gnd cell_6t
Xbit_r176_c49 bl[49] br[49] wl[176] vdd gnd cell_6t
Xbit_r177_c49 bl[49] br[49] wl[177] vdd gnd cell_6t
Xbit_r178_c49 bl[49] br[49] wl[178] vdd gnd cell_6t
Xbit_r179_c49 bl[49] br[49] wl[179] vdd gnd cell_6t
Xbit_r180_c49 bl[49] br[49] wl[180] vdd gnd cell_6t
Xbit_r181_c49 bl[49] br[49] wl[181] vdd gnd cell_6t
Xbit_r182_c49 bl[49] br[49] wl[182] vdd gnd cell_6t
Xbit_r183_c49 bl[49] br[49] wl[183] vdd gnd cell_6t
Xbit_r184_c49 bl[49] br[49] wl[184] vdd gnd cell_6t
Xbit_r185_c49 bl[49] br[49] wl[185] vdd gnd cell_6t
Xbit_r186_c49 bl[49] br[49] wl[186] vdd gnd cell_6t
Xbit_r187_c49 bl[49] br[49] wl[187] vdd gnd cell_6t
Xbit_r188_c49 bl[49] br[49] wl[188] vdd gnd cell_6t
Xbit_r189_c49 bl[49] br[49] wl[189] vdd gnd cell_6t
Xbit_r190_c49 bl[49] br[49] wl[190] vdd gnd cell_6t
Xbit_r191_c49 bl[49] br[49] wl[191] vdd gnd cell_6t
Xbit_r192_c49 bl[49] br[49] wl[192] vdd gnd cell_6t
Xbit_r193_c49 bl[49] br[49] wl[193] vdd gnd cell_6t
Xbit_r194_c49 bl[49] br[49] wl[194] vdd gnd cell_6t
Xbit_r195_c49 bl[49] br[49] wl[195] vdd gnd cell_6t
Xbit_r196_c49 bl[49] br[49] wl[196] vdd gnd cell_6t
Xbit_r197_c49 bl[49] br[49] wl[197] vdd gnd cell_6t
Xbit_r198_c49 bl[49] br[49] wl[198] vdd gnd cell_6t
Xbit_r199_c49 bl[49] br[49] wl[199] vdd gnd cell_6t
Xbit_r200_c49 bl[49] br[49] wl[200] vdd gnd cell_6t
Xbit_r201_c49 bl[49] br[49] wl[201] vdd gnd cell_6t
Xbit_r202_c49 bl[49] br[49] wl[202] vdd gnd cell_6t
Xbit_r203_c49 bl[49] br[49] wl[203] vdd gnd cell_6t
Xbit_r204_c49 bl[49] br[49] wl[204] vdd gnd cell_6t
Xbit_r205_c49 bl[49] br[49] wl[205] vdd gnd cell_6t
Xbit_r206_c49 bl[49] br[49] wl[206] vdd gnd cell_6t
Xbit_r207_c49 bl[49] br[49] wl[207] vdd gnd cell_6t
Xbit_r208_c49 bl[49] br[49] wl[208] vdd gnd cell_6t
Xbit_r209_c49 bl[49] br[49] wl[209] vdd gnd cell_6t
Xbit_r210_c49 bl[49] br[49] wl[210] vdd gnd cell_6t
Xbit_r211_c49 bl[49] br[49] wl[211] vdd gnd cell_6t
Xbit_r212_c49 bl[49] br[49] wl[212] vdd gnd cell_6t
Xbit_r213_c49 bl[49] br[49] wl[213] vdd gnd cell_6t
Xbit_r214_c49 bl[49] br[49] wl[214] vdd gnd cell_6t
Xbit_r215_c49 bl[49] br[49] wl[215] vdd gnd cell_6t
Xbit_r216_c49 bl[49] br[49] wl[216] vdd gnd cell_6t
Xbit_r217_c49 bl[49] br[49] wl[217] vdd gnd cell_6t
Xbit_r218_c49 bl[49] br[49] wl[218] vdd gnd cell_6t
Xbit_r219_c49 bl[49] br[49] wl[219] vdd gnd cell_6t
Xbit_r220_c49 bl[49] br[49] wl[220] vdd gnd cell_6t
Xbit_r221_c49 bl[49] br[49] wl[221] vdd gnd cell_6t
Xbit_r222_c49 bl[49] br[49] wl[222] vdd gnd cell_6t
Xbit_r223_c49 bl[49] br[49] wl[223] vdd gnd cell_6t
Xbit_r224_c49 bl[49] br[49] wl[224] vdd gnd cell_6t
Xbit_r225_c49 bl[49] br[49] wl[225] vdd gnd cell_6t
Xbit_r226_c49 bl[49] br[49] wl[226] vdd gnd cell_6t
Xbit_r227_c49 bl[49] br[49] wl[227] vdd gnd cell_6t
Xbit_r228_c49 bl[49] br[49] wl[228] vdd gnd cell_6t
Xbit_r229_c49 bl[49] br[49] wl[229] vdd gnd cell_6t
Xbit_r230_c49 bl[49] br[49] wl[230] vdd gnd cell_6t
Xbit_r231_c49 bl[49] br[49] wl[231] vdd gnd cell_6t
Xbit_r232_c49 bl[49] br[49] wl[232] vdd gnd cell_6t
Xbit_r233_c49 bl[49] br[49] wl[233] vdd gnd cell_6t
Xbit_r234_c49 bl[49] br[49] wl[234] vdd gnd cell_6t
Xbit_r235_c49 bl[49] br[49] wl[235] vdd gnd cell_6t
Xbit_r236_c49 bl[49] br[49] wl[236] vdd gnd cell_6t
Xbit_r237_c49 bl[49] br[49] wl[237] vdd gnd cell_6t
Xbit_r238_c49 bl[49] br[49] wl[238] vdd gnd cell_6t
Xbit_r239_c49 bl[49] br[49] wl[239] vdd gnd cell_6t
Xbit_r240_c49 bl[49] br[49] wl[240] vdd gnd cell_6t
Xbit_r241_c49 bl[49] br[49] wl[241] vdd gnd cell_6t
Xbit_r242_c49 bl[49] br[49] wl[242] vdd gnd cell_6t
Xbit_r243_c49 bl[49] br[49] wl[243] vdd gnd cell_6t
Xbit_r244_c49 bl[49] br[49] wl[244] vdd gnd cell_6t
Xbit_r245_c49 bl[49] br[49] wl[245] vdd gnd cell_6t
Xbit_r246_c49 bl[49] br[49] wl[246] vdd gnd cell_6t
Xbit_r247_c49 bl[49] br[49] wl[247] vdd gnd cell_6t
Xbit_r248_c49 bl[49] br[49] wl[248] vdd gnd cell_6t
Xbit_r249_c49 bl[49] br[49] wl[249] vdd gnd cell_6t
Xbit_r250_c49 bl[49] br[49] wl[250] vdd gnd cell_6t
Xbit_r251_c49 bl[49] br[49] wl[251] vdd gnd cell_6t
Xbit_r252_c49 bl[49] br[49] wl[252] vdd gnd cell_6t
Xbit_r253_c49 bl[49] br[49] wl[253] vdd gnd cell_6t
Xbit_r254_c49 bl[49] br[49] wl[254] vdd gnd cell_6t
Xbit_r255_c49 bl[49] br[49] wl[255] vdd gnd cell_6t
Xbit_r256_c49 bl[49] br[49] wl[256] vdd gnd cell_6t
Xbit_r257_c49 bl[49] br[49] wl[257] vdd gnd cell_6t
Xbit_r258_c49 bl[49] br[49] wl[258] vdd gnd cell_6t
Xbit_r259_c49 bl[49] br[49] wl[259] vdd gnd cell_6t
Xbit_r260_c49 bl[49] br[49] wl[260] vdd gnd cell_6t
Xbit_r261_c49 bl[49] br[49] wl[261] vdd gnd cell_6t
Xbit_r262_c49 bl[49] br[49] wl[262] vdd gnd cell_6t
Xbit_r263_c49 bl[49] br[49] wl[263] vdd gnd cell_6t
Xbit_r264_c49 bl[49] br[49] wl[264] vdd gnd cell_6t
Xbit_r265_c49 bl[49] br[49] wl[265] vdd gnd cell_6t
Xbit_r266_c49 bl[49] br[49] wl[266] vdd gnd cell_6t
Xbit_r267_c49 bl[49] br[49] wl[267] vdd gnd cell_6t
Xbit_r268_c49 bl[49] br[49] wl[268] vdd gnd cell_6t
Xbit_r269_c49 bl[49] br[49] wl[269] vdd gnd cell_6t
Xbit_r270_c49 bl[49] br[49] wl[270] vdd gnd cell_6t
Xbit_r271_c49 bl[49] br[49] wl[271] vdd gnd cell_6t
Xbit_r272_c49 bl[49] br[49] wl[272] vdd gnd cell_6t
Xbit_r273_c49 bl[49] br[49] wl[273] vdd gnd cell_6t
Xbit_r274_c49 bl[49] br[49] wl[274] vdd gnd cell_6t
Xbit_r275_c49 bl[49] br[49] wl[275] vdd gnd cell_6t
Xbit_r276_c49 bl[49] br[49] wl[276] vdd gnd cell_6t
Xbit_r277_c49 bl[49] br[49] wl[277] vdd gnd cell_6t
Xbit_r278_c49 bl[49] br[49] wl[278] vdd gnd cell_6t
Xbit_r279_c49 bl[49] br[49] wl[279] vdd gnd cell_6t
Xbit_r280_c49 bl[49] br[49] wl[280] vdd gnd cell_6t
Xbit_r281_c49 bl[49] br[49] wl[281] vdd gnd cell_6t
Xbit_r282_c49 bl[49] br[49] wl[282] vdd gnd cell_6t
Xbit_r283_c49 bl[49] br[49] wl[283] vdd gnd cell_6t
Xbit_r284_c49 bl[49] br[49] wl[284] vdd gnd cell_6t
Xbit_r285_c49 bl[49] br[49] wl[285] vdd gnd cell_6t
Xbit_r286_c49 bl[49] br[49] wl[286] vdd gnd cell_6t
Xbit_r287_c49 bl[49] br[49] wl[287] vdd gnd cell_6t
Xbit_r288_c49 bl[49] br[49] wl[288] vdd gnd cell_6t
Xbit_r289_c49 bl[49] br[49] wl[289] vdd gnd cell_6t
Xbit_r290_c49 bl[49] br[49] wl[290] vdd gnd cell_6t
Xbit_r291_c49 bl[49] br[49] wl[291] vdd gnd cell_6t
Xbit_r292_c49 bl[49] br[49] wl[292] vdd gnd cell_6t
Xbit_r293_c49 bl[49] br[49] wl[293] vdd gnd cell_6t
Xbit_r294_c49 bl[49] br[49] wl[294] vdd gnd cell_6t
Xbit_r295_c49 bl[49] br[49] wl[295] vdd gnd cell_6t
Xbit_r296_c49 bl[49] br[49] wl[296] vdd gnd cell_6t
Xbit_r297_c49 bl[49] br[49] wl[297] vdd gnd cell_6t
Xbit_r298_c49 bl[49] br[49] wl[298] vdd gnd cell_6t
Xbit_r299_c49 bl[49] br[49] wl[299] vdd gnd cell_6t
Xbit_r300_c49 bl[49] br[49] wl[300] vdd gnd cell_6t
Xbit_r301_c49 bl[49] br[49] wl[301] vdd gnd cell_6t
Xbit_r302_c49 bl[49] br[49] wl[302] vdd gnd cell_6t
Xbit_r303_c49 bl[49] br[49] wl[303] vdd gnd cell_6t
Xbit_r304_c49 bl[49] br[49] wl[304] vdd gnd cell_6t
Xbit_r305_c49 bl[49] br[49] wl[305] vdd gnd cell_6t
Xbit_r306_c49 bl[49] br[49] wl[306] vdd gnd cell_6t
Xbit_r307_c49 bl[49] br[49] wl[307] vdd gnd cell_6t
Xbit_r308_c49 bl[49] br[49] wl[308] vdd gnd cell_6t
Xbit_r309_c49 bl[49] br[49] wl[309] vdd gnd cell_6t
Xbit_r310_c49 bl[49] br[49] wl[310] vdd gnd cell_6t
Xbit_r311_c49 bl[49] br[49] wl[311] vdd gnd cell_6t
Xbit_r312_c49 bl[49] br[49] wl[312] vdd gnd cell_6t
Xbit_r313_c49 bl[49] br[49] wl[313] vdd gnd cell_6t
Xbit_r314_c49 bl[49] br[49] wl[314] vdd gnd cell_6t
Xbit_r315_c49 bl[49] br[49] wl[315] vdd gnd cell_6t
Xbit_r316_c49 bl[49] br[49] wl[316] vdd gnd cell_6t
Xbit_r317_c49 bl[49] br[49] wl[317] vdd gnd cell_6t
Xbit_r318_c49 bl[49] br[49] wl[318] vdd gnd cell_6t
Xbit_r319_c49 bl[49] br[49] wl[319] vdd gnd cell_6t
Xbit_r320_c49 bl[49] br[49] wl[320] vdd gnd cell_6t
Xbit_r321_c49 bl[49] br[49] wl[321] vdd gnd cell_6t
Xbit_r322_c49 bl[49] br[49] wl[322] vdd gnd cell_6t
Xbit_r323_c49 bl[49] br[49] wl[323] vdd gnd cell_6t
Xbit_r324_c49 bl[49] br[49] wl[324] vdd gnd cell_6t
Xbit_r325_c49 bl[49] br[49] wl[325] vdd gnd cell_6t
Xbit_r326_c49 bl[49] br[49] wl[326] vdd gnd cell_6t
Xbit_r327_c49 bl[49] br[49] wl[327] vdd gnd cell_6t
Xbit_r328_c49 bl[49] br[49] wl[328] vdd gnd cell_6t
Xbit_r329_c49 bl[49] br[49] wl[329] vdd gnd cell_6t
Xbit_r330_c49 bl[49] br[49] wl[330] vdd gnd cell_6t
Xbit_r331_c49 bl[49] br[49] wl[331] vdd gnd cell_6t
Xbit_r332_c49 bl[49] br[49] wl[332] vdd gnd cell_6t
Xbit_r333_c49 bl[49] br[49] wl[333] vdd gnd cell_6t
Xbit_r334_c49 bl[49] br[49] wl[334] vdd gnd cell_6t
Xbit_r335_c49 bl[49] br[49] wl[335] vdd gnd cell_6t
Xbit_r336_c49 bl[49] br[49] wl[336] vdd gnd cell_6t
Xbit_r337_c49 bl[49] br[49] wl[337] vdd gnd cell_6t
Xbit_r338_c49 bl[49] br[49] wl[338] vdd gnd cell_6t
Xbit_r339_c49 bl[49] br[49] wl[339] vdd gnd cell_6t
Xbit_r340_c49 bl[49] br[49] wl[340] vdd gnd cell_6t
Xbit_r341_c49 bl[49] br[49] wl[341] vdd gnd cell_6t
Xbit_r342_c49 bl[49] br[49] wl[342] vdd gnd cell_6t
Xbit_r343_c49 bl[49] br[49] wl[343] vdd gnd cell_6t
Xbit_r344_c49 bl[49] br[49] wl[344] vdd gnd cell_6t
Xbit_r345_c49 bl[49] br[49] wl[345] vdd gnd cell_6t
Xbit_r346_c49 bl[49] br[49] wl[346] vdd gnd cell_6t
Xbit_r347_c49 bl[49] br[49] wl[347] vdd gnd cell_6t
Xbit_r348_c49 bl[49] br[49] wl[348] vdd gnd cell_6t
Xbit_r349_c49 bl[49] br[49] wl[349] vdd gnd cell_6t
Xbit_r350_c49 bl[49] br[49] wl[350] vdd gnd cell_6t
Xbit_r351_c49 bl[49] br[49] wl[351] vdd gnd cell_6t
Xbit_r352_c49 bl[49] br[49] wl[352] vdd gnd cell_6t
Xbit_r353_c49 bl[49] br[49] wl[353] vdd gnd cell_6t
Xbit_r354_c49 bl[49] br[49] wl[354] vdd gnd cell_6t
Xbit_r355_c49 bl[49] br[49] wl[355] vdd gnd cell_6t
Xbit_r356_c49 bl[49] br[49] wl[356] vdd gnd cell_6t
Xbit_r357_c49 bl[49] br[49] wl[357] vdd gnd cell_6t
Xbit_r358_c49 bl[49] br[49] wl[358] vdd gnd cell_6t
Xbit_r359_c49 bl[49] br[49] wl[359] vdd gnd cell_6t
Xbit_r360_c49 bl[49] br[49] wl[360] vdd gnd cell_6t
Xbit_r361_c49 bl[49] br[49] wl[361] vdd gnd cell_6t
Xbit_r362_c49 bl[49] br[49] wl[362] vdd gnd cell_6t
Xbit_r363_c49 bl[49] br[49] wl[363] vdd gnd cell_6t
Xbit_r364_c49 bl[49] br[49] wl[364] vdd gnd cell_6t
Xbit_r365_c49 bl[49] br[49] wl[365] vdd gnd cell_6t
Xbit_r366_c49 bl[49] br[49] wl[366] vdd gnd cell_6t
Xbit_r367_c49 bl[49] br[49] wl[367] vdd gnd cell_6t
Xbit_r368_c49 bl[49] br[49] wl[368] vdd gnd cell_6t
Xbit_r369_c49 bl[49] br[49] wl[369] vdd gnd cell_6t
Xbit_r370_c49 bl[49] br[49] wl[370] vdd gnd cell_6t
Xbit_r371_c49 bl[49] br[49] wl[371] vdd gnd cell_6t
Xbit_r372_c49 bl[49] br[49] wl[372] vdd gnd cell_6t
Xbit_r373_c49 bl[49] br[49] wl[373] vdd gnd cell_6t
Xbit_r374_c49 bl[49] br[49] wl[374] vdd gnd cell_6t
Xbit_r375_c49 bl[49] br[49] wl[375] vdd gnd cell_6t
Xbit_r376_c49 bl[49] br[49] wl[376] vdd gnd cell_6t
Xbit_r377_c49 bl[49] br[49] wl[377] vdd gnd cell_6t
Xbit_r378_c49 bl[49] br[49] wl[378] vdd gnd cell_6t
Xbit_r379_c49 bl[49] br[49] wl[379] vdd gnd cell_6t
Xbit_r380_c49 bl[49] br[49] wl[380] vdd gnd cell_6t
Xbit_r381_c49 bl[49] br[49] wl[381] vdd gnd cell_6t
Xbit_r382_c49 bl[49] br[49] wl[382] vdd gnd cell_6t
Xbit_r383_c49 bl[49] br[49] wl[383] vdd gnd cell_6t
Xbit_r384_c49 bl[49] br[49] wl[384] vdd gnd cell_6t
Xbit_r385_c49 bl[49] br[49] wl[385] vdd gnd cell_6t
Xbit_r386_c49 bl[49] br[49] wl[386] vdd gnd cell_6t
Xbit_r387_c49 bl[49] br[49] wl[387] vdd gnd cell_6t
Xbit_r388_c49 bl[49] br[49] wl[388] vdd gnd cell_6t
Xbit_r389_c49 bl[49] br[49] wl[389] vdd gnd cell_6t
Xbit_r390_c49 bl[49] br[49] wl[390] vdd gnd cell_6t
Xbit_r391_c49 bl[49] br[49] wl[391] vdd gnd cell_6t
Xbit_r392_c49 bl[49] br[49] wl[392] vdd gnd cell_6t
Xbit_r393_c49 bl[49] br[49] wl[393] vdd gnd cell_6t
Xbit_r394_c49 bl[49] br[49] wl[394] vdd gnd cell_6t
Xbit_r395_c49 bl[49] br[49] wl[395] vdd gnd cell_6t
Xbit_r396_c49 bl[49] br[49] wl[396] vdd gnd cell_6t
Xbit_r397_c49 bl[49] br[49] wl[397] vdd gnd cell_6t
Xbit_r398_c49 bl[49] br[49] wl[398] vdd gnd cell_6t
Xbit_r399_c49 bl[49] br[49] wl[399] vdd gnd cell_6t
Xbit_r400_c49 bl[49] br[49] wl[400] vdd gnd cell_6t
Xbit_r401_c49 bl[49] br[49] wl[401] vdd gnd cell_6t
Xbit_r402_c49 bl[49] br[49] wl[402] vdd gnd cell_6t
Xbit_r403_c49 bl[49] br[49] wl[403] vdd gnd cell_6t
Xbit_r404_c49 bl[49] br[49] wl[404] vdd gnd cell_6t
Xbit_r405_c49 bl[49] br[49] wl[405] vdd gnd cell_6t
Xbit_r406_c49 bl[49] br[49] wl[406] vdd gnd cell_6t
Xbit_r407_c49 bl[49] br[49] wl[407] vdd gnd cell_6t
Xbit_r408_c49 bl[49] br[49] wl[408] vdd gnd cell_6t
Xbit_r409_c49 bl[49] br[49] wl[409] vdd gnd cell_6t
Xbit_r410_c49 bl[49] br[49] wl[410] vdd gnd cell_6t
Xbit_r411_c49 bl[49] br[49] wl[411] vdd gnd cell_6t
Xbit_r412_c49 bl[49] br[49] wl[412] vdd gnd cell_6t
Xbit_r413_c49 bl[49] br[49] wl[413] vdd gnd cell_6t
Xbit_r414_c49 bl[49] br[49] wl[414] vdd gnd cell_6t
Xbit_r415_c49 bl[49] br[49] wl[415] vdd gnd cell_6t
Xbit_r416_c49 bl[49] br[49] wl[416] vdd gnd cell_6t
Xbit_r417_c49 bl[49] br[49] wl[417] vdd gnd cell_6t
Xbit_r418_c49 bl[49] br[49] wl[418] vdd gnd cell_6t
Xbit_r419_c49 bl[49] br[49] wl[419] vdd gnd cell_6t
Xbit_r420_c49 bl[49] br[49] wl[420] vdd gnd cell_6t
Xbit_r421_c49 bl[49] br[49] wl[421] vdd gnd cell_6t
Xbit_r422_c49 bl[49] br[49] wl[422] vdd gnd cell_6t
Xbit_r423_c49 bl[49] br[49] wl[423] vdd gnd cell_6t
Xbit_r424_c49 bl[49] br[49] wl[424] vdd gnd cell_6t
Xbit_r425_c49 bl[49] br[49] wl[425] vdd gnd cell_6t
Xbit_r426_c49 bl[49] br[49] wl[426] vdd gnd cell_6t
Xbit_r427_c49 bl[49] br[49] wl[427] vdd gnd cell_6t
Xbit_r428_c49 bl[49] br[49] wl[428] vdd gnd cell_6t
Xbit_r429_c49 bl[49] br[49] wl[429] vdd gnd cell_6t
Xbit_r430_c49 bl[49] br[49] wl[430] vdd gnd cell_6t
Xbit_r431_c49 bl[49] br[49] wl[431] vdd gnd cell_6t
Xbit_r432_c49 bl[49] br[49] wl[432] vdd gnd cell_6t
Xbit_r433_c49 bl[49] br[49] wl[433] vdd gnd cell_6t
Xbit_r434_c49 bl[49] br[49] wl[434] vdd gnd cell_6t
Xbit_r435_c49 bl[49] br[49] wl[435] vdd gnd cell_6t
Xbit_r436_c49 bl[49] br[49] wl[436] vdd gnd cell_6t
Xbit_r437_c49 bl[49] br[49] wl[437] vdd gnd cell_6t
Xbit_r438_c49 bl[49] br[49] wl[438] vdd gnd cell_6t
Xbit_r439_c49 bl[49] br[49] wl[439] vdd gnd cell_6t
Xbit_r440_c49 bl[49] br[49] wl[440] vdd gnd cell_6t
Xbit_r441_c49 bl[49] br[49] wl[441] vdd gnd cell_6t
Xbit_r442_c49 bl[49] br[49] wl[442] vdd gnd cell_6t
Xbit_r443_c49 bl[49] br[49] wl[443] vdd gnd cell_6t
Xbit_r444_c49 bl[49] br[49] wl[444] vdd gnd cell_6t
Xbit_r445_c49 bl[49] br[49] wl[445] vdd gnd cell_6t
Xbit_r446_c49 bl[49] br[49] wl[446] vdd gnd cell_6t
Xbit_r447_c49 bl[49] br[49] wl[447] vdd gnd cell_6t
Xbit_r448_c49 bl[49] br[49] wl[448] vdd gnd cell_6t
Xbit_r449_c49 bl[49] br[49] wl[449] vdd gnd cell_6t
Xbit_r450_c49 bl[49] br[49] wl[450] vdd gnd cell_6t
Xbit_r451_c49 bl[49] br[49] wl[451] vdd gnd cell_6t
Xbit_r452_c49 bl[49] br[49] wl[452] vdd gnd cell_6t
Xbit_r453_c49 bl[49] br[49] wl[453] vdd gnd cell_6t
Xbit_r454_c49 bl[49] br[49] wl[454] vdd gnd cell_6t
Xbit_r455_c49 bl[49] br[49] wl[455] vdd gnd cell_6t
Xbit_r456_c49 bl[49] br[49] wl[456] vdd gnd cell_6t
Xbit_r457_c49 bl[49] br[49] wl[457] vdd gnd cell_6t
Xbit_r458_c49 bl[49] br[49] wl[458] vdd gnd cell_6t
Xbit_r459_c49 bl[49] br[49] wl[459] vdd gnd cell_6t
Xbit_r460_c49 bl[49] br[49] wl[460] vdd gnd cell_6t
Xbit_r461_c49 bl[49] br[49] wl[461] vdd gnd cell_6t
Xbit_r462_c49 bl[49] br[49] wl[462] vdd gnd cell_6t
Xbit_r463_c49 bl[49] br[49] wl[463] vdd gnd cell_6t
Xbit_r464_c49 bl[49] br[49] wl[464] vdd gnd cell_6t
Xbit_r465_c49 bl[49] br[49] wl[465] vdd gnd cell_6t
Xbit_r466_c49 bl[49] br[49] wl[466] vdd gnd cell_6t
Xbit_r467_c49 bl[49] br[49] wl[467] vdd gnd cell_6t
Xbit_r468_c49 bl[49] br[49] wl[468] vdd gnd cell_6t
Xbit_r469_c49 bl[49] br[49] wl[469] vdd gnd cell_6t
Xbit_r470_c49 bl[49] br[49] wl[470] vdd gnd cell_6t
Xbit_r471_c49 bl[49] br[49] wl[471] vdd gnd cell_6t
Xbit_r472_c49 bl[49] br[49] wl[472] vdd gnd cell_6t
Xbit_r473_c49 bl[49] br[49] wl[473] vdd gnd cell_6t
Xbit_r474_c49 bl[49] br[49] wl[474] vdd gnd cell_6t
Xbit_r475_c49 bl[49] br[49] wl[475] vdd gnd cell_6t
Xbit_r476_c49 bl[49] br[49] wl[476] vdd gnd cell_6t
Xbit_r477_c49 bl[49] br[49] wl[477] vdd gnd cell_6t
Xbit_r478_c49 bl[49] br[49] wl[478] vdd gnd cell_6t
Xbit_r479_c49 bl[49] br[49] wl[479] vdd gnd cell_6t
Xbit_r480_c49 bl[49] br[49] wl[480] vdd gnd cell_6t
Xbit_r481_c49 bl[49] br[49] wl[481] vdd gnd cell_6t
Xbit_r482_c49 bl[49] br[49] wl[482] vdd gnd cell_6t
Xbit_r483_c49 bl[49] br[49] wl[483] vdd gnd cell_6t
Xbit_r484_c49 bl[49] br[49] wl[484] vdd gnd cell_6t
Xbit_r485_c49 bl[49] br[49] wl[485] vdd gnd cell_6t
Xbit_r486_c49 bl[49] br[49] wl[486] vdd gnd cell_6t
Xbit_r487_c49 bl[49] br[49] wl[487] vdd gnd cell_6t
Xbit_r488_c49 bl[49] br[49] wl[488] vdd gnd cell_6t
Xbit_r489_c49 bl[49] br[49] wl[489] vdd gnd cell_6t
Xbit_r490_c49 bl[49] br[49] wl[490] vdd gnd cell_6t
Xbit_r491_c49 bl[49] br[49] wl[491] vdd gnd cell_6t
Xbit_r492_c49 bl[49] br[49] wl[492] vdd gnd cell_6t
Xbit_r493_c49 bl[49] br[49] wl[493] vdd gnd cell_6t
Xbit_r494_c49 bl[49] br[49] wl[494] vdd gnd cell_6t
Xbit_r495_c49 bl[49] br[49] wl[495] vdd gnd cell_6t
Xbit_r496_c49 bl[49] br[49] wl[496] vdd gnd cell_6t
Xbit_r497_c49 bl[49] br[49] wl[497] vdd gnd cell_6t
Xbit_r498_c49 bl[49] br[49] wl[498] vdd gnd cell_6t
Xbit_r499_c49 bl[49] br[49] wl[499] vdd gnd cell_6t
Xbit_r500_c49 bl[49] br[49] wl[500] vdd gnd cell_6t
Xbit_r501_c49 bl[49] br[49] wl[501] vdd gnd cell_6t
Xbit_r502_c49 bl[49] br[49] wl[502] vdd gnd cell_6t
Xbit_r503_c49 bl[49] br[49] wl[503] vdd gnd cell_6t
Xbit_r504_c49 bl[49] br[49] wl[504] vdd gnd cell_6t
Xbit_r505_c49 bl[49] br[49] wl[505] vdd gnd cell_6t
Xbit_r506_c49 bl[49] br[49] wl[506] vdd gnd cell_6t
Xbit_r507_c49 bl[49] br[49] wl[507] vdd gnd cell_6t
Xbit_r508_c49 bl[49] br[49] wl[508] vdd gnd cell_6t
Xbit_r509_c49 bl[49] br[49] wl[509] vdd gnd cell_6t
Xbit_r510_c49 bl[49] br[49] wl[510] vdd gnd cell_6t
Xbit_r511_c49 bl[49] br[49] wl[511] vdd gnd cell_6t
Xbit_r0_c50 bl[50] br[50] wl[0] vdd gnd cell_6t
Xbit_r1_c50 bl[50] br[50] wl[1] vdd gnd cell_6t
Xbit_r2_c50 bl[50] br[50] wl[2] vdd gnd cell_6t
Xbit_r3_c50 bl[50] br[50] wl[3] vdd gnd cell_6t
Xbit_r4_c50 bl[50] br[50] wl[4] vdd gnd cell_6t
Xbit_r5_c50 bl[50] br[50] wl[5] vdd gnd cell_6t
Xbit_r6_c50 bl[50] br[50] wl[6] vdd gnd cell_6t
Xbit_r7_c50 bl[50] br[50] wl[7] vdd gnd cell_6t
Xbit_r8_c50 bl[50] br[50] wl[8] vdd gnd cell_6t
Xbit_r9_c50 bl[50] br[50] wl[9] vdd gnd cell_6t
Xbit_r10_c50 bl[50] br[50] wl[10] vdd gnd cell_6t
Xbit_r11_c50 bl[50] br[50] wl[11] vdd gnd cell_6t
Xbit_r12_c50 bl[50] br[50] wl[12] vdd gnd cell_6t
Xbit_r13_c50 bl[50] br[50] wl[13] vdd gnd cell_6t
Xbit_r14_c50 bl[50] br[50] wl[14] vdd gnd cell_6t
Xbit_r15_c50 bl[50] br[50] wl[15] vdd gnd cell_6t
Xbit_r16_c50 bl[50] br[50] wl[16] vdd gnd cell_6t
Xbit_r17_c50 bl[50] br[50] wl[17] vdd gnd cell_6t
Xbit_r18_c50 bl[50] br[50] wl[18] vdd gnd cell_6t
Xbit_r19_c50 bl[50] br[50] wl[19] vdd gnd cell_6t
Xbit_r20_c50 bl[50] br[50] wl[20] vdd gnd cell_6t
Xbit_r21_c50 bl[50] br[50] wl[21] vdd gnd cell_6t
Xbit_r22_c50 bl[50] br[50] wl[22] vdd gnd cell_6t
Xbit_r23_c50 bl[50] br[50] wl[23] vdd gnd cell_6t
Xbit_r24_c50 bl[50] br[50] wl[24] vdd gnd cell_6t
Xbit_r25_c50 bl[50] br[50] wl[25] vdd gnd cell_6t
Xbit_r26_c50 bl[50] br[50] wl[26] vdd gnd cell_6t
Xbit_r27_c50 bl[50] br[50] wl[27] vdd gnd cell_6t
Xbit_r28_c50 bl[50] br[50] wl[28] vdd gnd cell_6t
Xbit_r29_c50 bl[50] br[50] wl[29] vdd gnd cell_6t
Xbit_r30_c50 bl[50] br[50] wl[30] vdd gnd cell_6t
Xbit_r31_c50 bl[50] br[50] wl[31] vdd gnd cell_6t
Xbit_r32_c50 bl[50] br[50] wl[32] vdd gnd cell_6t
Xbit_r33_c50 bl[50] br[50] wl[33] vdd gnd cell_6t
Xbit_r34_c50 bl[50] br[50] wl[34] vdd gnd cell_6t
Xbit_r35_c50 bl[50] br[50] wl[35] vdd gnd cell_6t
Xbit_r36_c50 bl[50] br[50] wl[36] vdd gnd cell_6t
Xbit_r37_c50 bl[50] br[50] wl[37] vdd gnd cell_6t
Xbit_r38_c50 bl[50] br[50] wl[38] vdd gnd cell_6t
Xbit_r39_c50 bl[50] br[50] wl[39] vdd gnd cell_6t
Xbit_r40_c50 bl[50] br[50] wl[40] vdd gnd cell_6t
Xbit_r41_c50 bl[50] br[50] wl[41] vdd gnd cell_6t
Xbit_r42_c50 bl[50] br[50] wl[42] vdd gnd cell_6t
Xbit_r43_c50 bl[50] br[50] wl[43] vdd gnd cell_6t
Xbit_r44_c50 bl[50] br[50] wl[44] vdd gnd cell_6t
Xbit_r45_c50 bl[50] br[50] wl[45] vdd gnd cell_6t
Xbit_r46_c50 bl[50] br[50] wl[46] vdd gnd cell_6t
Xbit_r47_c50 bl[50] br[50] wl[47] vdd gnd cell_6t
Xbit_r48_c50 bl[50] br[50] wl[48] vdd gnd cell_6t
Xbit_r49_c50 bl[50] br[50] wl[49] vdd gnd cell_6t
Xbit_r50_c50 bl[50] br[50] wl[50] vdd gnd cell_6t
Xbit_r51_c50 bl[50] br[50] wl[51] vdd gnd cell_6t
Xbit_r52_c50 bl[50] br[50] wl[52] vdd gnd cell_6t
Xbit_r53_c50 bl[50] br[50] wl[53] vdd gnd cell_6t
Xbit_r54_c50 bl[50] br[50] wl[54] vdd gnd cell_6t
Xbit_r55_c50 bl[50] br[50] wl[55] vdd gnd cell_6t
Xbit_r56_c50 bl[50] br[50] wl[56] vdd gnd cell_6t
Xbit_r57_c50 bl[50] br[50] wl[57] vdd gnd cell_6t
Xbit_r58_c50 bl[50] br[50] wl[58] vdd gnd cell_6t
Xbit_r59_c50 bl[50] br[50] wl[59] vdd gnd cell_6t
Xbit_r60_c50 bl[50] br[50] wl[60] vdd gnd cell_6t
Xbit_r61_c50 bl[50] br[50] wl[61] vdd gnd cell_6t
Xbit_r62_c50 bl[50] br[50] wl[62] vdd gnd cell_6t
Xbit_r63_c50 bl[50] br[50] wl[63] vdd gnd cell_6t
Xbit_r64_c50 bl[50] br[50] wl[64] vdd gnd cell_6t
Xbit_r65_c50 bl[50] br[50] wl[65] vdd gnd cell_6t
Xbit_r66_c50 bl[50] br[50] wl[66] vdd gnd cell_6t
Xbit_r67_c50 bl[50] br[50] wl[67] vdd gnd cell_6t
Xbit_r68_c50 bl[50] br[50] wl[68] vdd gnd cell_6t
Xbit_r69_c50 bl[50] br[50] wl[69] vdd gnd cell_6t
Xbit_r70_c50 bl[50] br[50] wl[70] vdd gnd cell_6t
Xbit_r71_c50 bl[50] br[50] wl[71] vdd gnd cell_6t
Xbit_r72_c50 bl[50] br[50] wl[72] vdd gnd cell_6t
Xbit_r73_c50 bl[50] br[50] wl[73] vdd gnd cell_6t
Xbit_r74_c50 bl[50] br[50] wl[74] vdd gnd cell_6t
Xbit_r75_c50 bl[50] br[50] wl[75] vdd gnd cell_6t
Xbit_r76_c50 bl[50] br[50] wl[76] vdd gnd cell_6t
Xbit_r77_c50 bl[50] br[50] wl[77] vdd gnd cell_6t
Xbit_r78_c50 bl[50] br[50] wl[78] vdd gnd cell_6t
Xbit_r79_c50 bl[50] br[50] wl[79] vdd gnd cell_6t
Xbit_r80_c50 bl[50] br[50] wl[80] vdd gnd cell_6t
Xbit_r81_c50 bl[50] br[50] wl[81] vdd gnd cell_6t
Xbit_r82_c50 bl[50] br[50] wl[82] vdd gnd cell_6t
Xbit_r83_c50 bl[50] br[50] wl[83] vdd gnd cell_6t
Xbit_r84_c50 bl[50] br[50] wl[84] vdd gnd cell_6t
Xbit_r85_c50 bl[50] br[50] wl[85] vdd gnd cell_6t
Xbit_r86_c50 bl[50] br[50] wl[86] vdd gnd cell_6t
Xbit_r87_c50 bl[50] br[50] wl[87] vdd gnd cell_6t
Xbit_r88_c50 bl[50] br[50] wl[88] vdd gnd cell_6t
Xbit_r89_c50 bl[50] br[50] wl[89] vdd gnd cell_6t
Xbit_r90_c50 bl[50] br[50] wl[90] vdd gnd cell_6t
Xbit_r91_c50 bl[50] br[50] wl[91] vdd gnd cell_6t
Xbit_r92_c50 bl[50] br[50] wl[92] vdd gnd cell_6t
Xbit_r93_c50 bl[50] br[50] wl[93] vdd gnd cell_6t
Xbit_r94_c50 bl[50] br[50] wl[94] vdd gnd cell_6t
Xbit_r95_c50 bl[50] br[50] wl[95] vdd gnd cell_6t
Xbit_r96_c50 bl[50] br[50] wl[96] vdd gnd cell_6t
Xbit_r97_c50 bl[50] br[50] wl[97] vdd gnd cell_6t
Xbit_r98_c50 bl[50] br[50] wl[98] vdd gnd cell_6t
Xbit_r99_c50 bl[50] br[50] wl[99] vdd gnd cell_6t
Xbit_r100_c50 bl[50] br[50] wl[100] vdd gnd cell_6t
Xbit_r101_c50 bl[50] br[50] wl[101] vdd gnd cell_6t
Xbit_r102_c50 bl[50] br[50] wl[102] vdd gnd cell_6t
Xbit_r103_c50 bl[50] br[50] wl[103] vdd gnd cell_6t
Xbit_r104_c50 bl[50] br[50] wl[104] vdd gnd cell_6t
Xbit_r105_c50 bl[50] br[50] wl[105] vdd gnd cell_6t
Xbit_r106_c50 bl[50] br[50] wl[106] vdd gnd cell_6t
Xbit_r107_c50 bl[50] br[50] wl[107] vdd gnd cell_6t
Xbit_r108_c50 bl[50] br[50] wl[108] vdd gnd cell_6t
Xbit_r109_c50 bl[50] br[50] wl[109] vdd gnd cell_6t
Xbit_r110_c50 bl[50] br[50] wl[110] vdd gnd cell_6t
Xbit_r111_c50 bl[50] br[50] wl[111] vdd gnd cell_6t
Xbit_r112_c50 bl[50] br[50] wl[112] vdd gnd cell_6t
Xbit_r113_c50 bl[50] br[50] wl[113] vdd gnd cell_6t
Xbit_r114_c50 bl[50] br[50] wl[114] vdd gnd cell_6t
Xbit_r115_c50 bl[50] br[50] wl[115] vdd gnd cell_6t
Xbit_r116_c50 bl[50] br[50] wl[116] vdd gnd cell_6t
Xbit_r117_c50 bl[50] br[50] wl[117] vdd gnd cell_6t
Xbit_r118_c50 bl[50] br[50] wl[118] vdd gnd cell_6t
Xbit_r119_c50 bl[50] br[50] wl[119] vdd gnd cell_6t
Xbit_r120_c50 bl[50] br[50] wl[120] vdd gnd cell_6t
Xbit_r121_c50 bl[50] br[50] wl[121] vdd gnd cell_6t
Xbit_r122_c50 bl[50] br[50] wl[122] vdd gnd cell_6t
Xbit_r123_c50 bl[50] br[50] wl[123] vdd gnd cell_6t
Xbit_r124_c50 bl[50] br[50] wl[124] vdd gnd cell_6t
Xbit_r125_c50 bl[50] br[50] wl[125] vdd gnd cell_6t
Xbit_r126_c50 bl[50] br[50] wl[126] vdd gnd cell_6t
Xbit_r127_c50 bl[50] br[50] wl[127] vdd gnd cell_6t
Xbit_r128_c50 bl[50] br[50] wl[128] vdd gnd cell_6t
Xbit_r129_c50 bl[50] br[50] wl[129] vdd gnd cell_6t
Xbit_r130_c50 bl[50] br[50] wl[130] vdd gnd cell_6t
Xbit_r131_c50 bl[50] br[50] wl[131] vdd gnd cell_6t
Xbit_r132_c50 bl[50] br[50] wl[132] vdd gnd cell_6t
Xbit_r133_c50 bl[50] br[50] wl[133] vdd gnd cell_6t
Xbit_r134_c50 bl[50] br[50] wl[134] vdd gnd cell_6t
Xbit_r135_c50 bl[50] br[50] wl[135] vdd gnd cell_6t
Xbit_r136_c50 bl[50] br[50] wl[136] vdd gnd cell_6t
Xbit_r137_c50 bl[50] br[50] wl[137] vdd gnd cell_6t
Xbit_r138_c50 bl[50] br[50] wl[138] vdd gnd cell_6t
Xbit_r139_c50 bl[50] br[50] wl[139] vdd gnd cell_6t
Xbit_r140_c50 bl[50] br[50] wl[140] vdd gnd cell_6t
Xbit_r141_c50 bl[50] br[50] wl[141] vdd gnd cell_6t
Xbit_r142_c50 bl[50] br[50] wl[142] vdd gnd cell_6t
Xbit_r143_c50 bl[50] br[50] wl[143] vdd gnd cell_6t
Xbit_r144_c50 bl[50] br[50] wl[144] vdd gnd cell_6t
Xbit_r145_c50 bl[50] br[50] wl[145] vdd gnd cell_6t
Xbit_r146_c50 bl[50] br[50] wl[146] vdd gnd cell_6t
Xbit_r147_c50 bl[50] br[50] wl[147] vdd gnd cell_6t
Xbit_r148_c50 bl[50] br[50] wl[148] vdd gnd cell_6t
Xbit_r149_c50 bl[50] br[50] wl[149] vdd gnd cell_6t
Xbit_r150_c50 bl[50] br[50] wl[150] vdd gnd cell_6t
Xbit_r151_c50 bl[50] br[50] wl[151] vdd gnd cell_6t
Xbit_r152_c50 bl[50] br[50] wl[152] vdd gnd cell_6t
Xbit_r153_c50 bl[50] br[50] wl[153] vdd gnd cell_6t
Xbit_r154_c50 bl[50] br[50] wl[154] vdd gnd cell_6t
Xbit_r155_c50 bl[50] br[50] wl[155] vdd gnd cell_6t
Xbit_r156_c50 bl[50] br[50] wl[156] vdd gnd cell_6t
Xbit_r157_c50 bl[50] br[50] wl[157] vdd gnd cell_6t
Xbit_r158_c50 bl[50] br[50] wl[158] vdd gnd cell_6t
Xbit_r159_c50 bl[50] br[50] wl[159] vdd gnd cell_6t
Xbit_r160_c50 bl[50] br[50] wl[160] vdd gnd cell_6t
Xbit_r161_c50 bl[50] br[50] wl[161] vdd gnd cell_6t
Xbit_r162_c50 bl[50] br[50] wl[162] vdd gnd cell_6t
Xbit_r163_c50 bl[50] br[50] wl[163] vdd gnd cell_6t
Xbit_r164_c50 bl[50] br[50] wl[164] vdd gnd cell_6t
Xbit_r165_c50 bl[50] br[50] wl[165] vdd gnd cell_6t
Xbit_r166_c50 bl[50] br[50] wl[166] vdd gnd cell_6t
Xbit_r167_c50 bl[50] br[50] wl[167] vdd gnd cell_6t
Xbit_r168_c50 bl[50] br[50] wl[168] vdd gnd cell_6t
Xbit_r169_c50 bl[50] br[50] wl[169] vdd gnd cell_6t
Xbit_r170_c50 bl[50] br[50] wl[170] vdd gnd cell_6t
Xbit_r171_c50 bl[50] br[50] wl[171] vdd gnd cell_6t
Xbit_r172_c50 bl[50] br[50] wl[172] vdd gnd cell_6t
Xbit_r173_c50 bl[50] br[50] wl[173] vdd gnd cell_6t
Xbit_r174_c50 bl[50] br[50] wl[174] vdd gnd cell_6t
Xbit_r175_c50 bl[50] br[50] wl[175] vdd gnd cell_6t
Xbit_r176_c50 bl[50] br[50] wl[176] vdd gnd cell_6t
Xbit_r177_c50 bl[50] br[50] wl[177] vdd gnd cell_6t
Xbit_r178_c50 bl[50] br[50] wl[178] vdd gnd cell_6t
Xbit_r179_c50 bl[50] br[50] wl[179] vdd gnd cell_6t
Xbit_r180_c50 bl[50] br[50] wl[180] vdd gnd cell_6t
Xbit_r181_c50 bl[50] br[50] wl[181] vdd gnd cell_6t
Xbit_r182_c50 bl[50] br[50] wl[182] vdd gnd cell_6t
Xbit_r183_c50 bl[50] br[50] wl[183] vdd gnd cell_6t
Xbit_r184_c50 bl[50] br[50] wl[184] vdd gnd cell_6t
Xbit_r185_c50 bl[50] br[50] wl[185] vdd gnd cell_6t
Xbit_r186_c50 bl[50] br[50] wl[186] vdd gnd cell_6t
Xbit_r187_c50 bl[50] br[50] wl[187] vdd gnd cell_6t
Xbit_r188_c50 bl[50] br[50] wl[188] vdd gnd cell_6t
Xbit_r189_c50 bl[50] br[50] wl[189] vdd gnd cell_6t
Xbit_r190_c50 bl[50] br[50] wl[190] vdd gnd cell_6t
Xbit_r191_c50 bl[50] br[50] wl[191] vdd gnd cell_6t
Xbit_r192_c50 bl[50] br[50] wl[192] vdd gnd cell_6t
Xbit_r193_c50 bl[50] br[50] wl[193] vdd gnd cell_6t
Xbit_r194_c50 bl[50] br[50] wl[194] vdd gnd cell_6t
Xbit_r195_c50 bl[50] br[50] wl[195] vdd gnd cell_6t
Xbit_r196_c50 bl[50] br[50] wl[196] vdd gnd cell_6t
Xbit_r197_c50 bl[50] br[50] wl[197] vdd gnd cell_6t
Xbit_r198_c50 bl[50] br[50] wl[198] vdd gnd cell_6t
Xbit_r199_c50 bl[50] br[50] wl[199] vdd gnd cell_6t
Xbit_r200_c50 bl[50] br[50] wl[200] vdd gnd cell_6t
Xbit_r201_c50 bl[50] br[50] wl[201] vdd gnd cell_6t
Xbit_r202_c50 bl[50] br[50] wl[202] vdd gnd cell_6t
Xbit_r203_c50 bl[50] br[50] wl[203] vdd gnd cell_6t
Xbit_r204_c50 bl[50] br[50] wl[204] vdd gnd cell_6t
Xbit_r205_c50 bl[50] br[50] wl[205] vdd gnd cell_6t
Xbit_r206_c50 bl[50] br[50] wl[206] vdd gnd cell_6t
Xbit_r207_c50 bl[50] br[50] wl[207] vdd gnd cell_6t
Xbit_r208_c50 bl[50] br[50] wl[208] vdd gnd cell_6t
Xbit_r209_c50 bl[50] br[50] wl[209] vdd gnd cell_6t
Xbit_r210_c50 bl[50] br[50] wl[210] vdd gnd cell_6t
Xbit_r211_c50 bl[50] br[50] wl[211] vdd gnd cell_6t
Xbit_r212_c50 bl[50] br[50] wl[212] vdd gnd cell_6t
Xbit_r213_c50 bl[50] br[50] wl[213] vdd gnd cell_6t
Xbit_r214_c50 bl[50] br[50] wl[214] vdd gnd cell_6t
Xbit_r215_c50 bl[50] br[50] wl[215] vdd gnd cell_6t
Xbit_r216_c50 bl[50] br[50] wl[216] vdd gnd cell_6t
Xbit_r217_c50 bl[50] br[50] wl[217] vdd gnd cell_6t
Xbit_r218_c50 bl[50] br[50] wl[218] vdd gnd cell_6t
Xbit_r219_c50 bl[50] br[50] wl[219] vdd gnd cell_6t
Xbit_r220_c50 bl[50] br[50] wl[220] vdd gnd cell_6t
Xbit_r221_c50 bl[50] br[50] wl[221] vdd gnd cell_6t
Xbit_r222_c50 bl[50] br[50] wl[222] vdd gnd cell_6t
Xbit_r223_c50 bl[50] br[50] wl[223] vdd gnd cell_6t
Xbit_r224_c50 bl[50] br[50] wl[224] vdd gnd cell_6t
Xbit_r225_c50 bl[50] br[50] wl[225] vdd gnd cell_6t
Xbit_r226_c50 bl[50] br[50] wl[226] vdd gnd cell_6t
Xbit_r227_c50 bl[50] br[50] wl[227] vdd gnd cell_6t
Xbit_r228_c50 bl[50] br[50] wl[228] vdd gnd cell_6t
Xbit_r229_c50 bl[50] br[50] wl[229] vdd gnd cell_6t
Xbit_r230_c50 bl[50] br[50] wl[230] vdd gnd cell_6t
Xbit_r231_c50 bl[50] br[50] wl[231] vdd gnd cell_6t
Xbit_r232_c50 bl[50] br[50] wl[232] vdd gnd cell_6t
Xbit_r233_c50 bl[50] br[50] wl[233] vdd gnd cell_6t
Xbit_r234_c50 bl[50] br[50] wl[234] vdd gnd cell_6t
Xbit_r235_c50 bl[50] br[50] wl[235] vdd gnd cell_6t
Xbit_r236_c50 bl[50] br[50] wl[236] vdd gnd cell_6t
Xbit_r237_c50 bl[50] br[50] wl[237] vdd gnd cell_6t
Xbit_r238_c50 bl[50] br[50] wl[238] vdd gnd cell_6t
Xbit_r239_c50 bl[50] br[50] wl[239] vdd gnd cell_6t
Xbit_r240_c50 bl[50] br[50] wl[240] vdd gnd cell_6t
Xbit_r241_c50 bl[50] br[50] wl[241] vdd gnd cell_6t
Xbit_r242_c50 bl[50] br[50] wl[242] vdd gnd cell_6t
Xbit_r243_c50 bl[50] br[50] wl[243] vdd gnd cell_6t
Xbit_r244_c50 bl[50] br[50] wl[244] vdd gnd cell_6t
Xbit_r245_c50 bl[50] br[50] wl[245] vdd gnd cell_6t
Xbit_r246_c50 bl[50] br[50] wl[246] vdd gnd cell_6t
Xbit_r247_c50 bl[50] br[50] wl[247] vdd gnd cell_6t
Xbit_r248_c50 bl[50] br[50] wl[248] vdd gnd cell_6t
Xbit_r249_c50 bl[50] br[50] wl[249] vdd gnd cell_6t
Xbit_r250_c50 bl[50] br[50] wl[250] vdd gnd cell_6t
Xbit_r251_c50 bl[50] br[50] wl[251] vdd gnd cell_6t
Xbit_r252_c50 bl[50] br[50] wl[252] vdd gnd cell_6t
Xbit_r253_c50 bl[50] br[50] wl[253] vdd gnd cell_6t
Xbit_r254_c50 bl[50] br[50] wl[254] vdd gnd cell_6t
Xbit_r255_c50 bl[50] br[50] wl[255] vdd gnd cell_6t
Xbit_r256_c50 bl[50] br[50] wl[256] vdd gnd cell_6t
Xbit_r257_c50 bl[50] br[50] wl[257] vdd gnd cell_6t
Xbit_r258_c50 bl[50] br[50] wl[258] vdd gnd cell_6t
Xbit_r259_c50 bl[50] br[50] wl[259] vdd gnd cell_6t
Xbit_r260_c50 bl[50] br[50] wl[260] vdd gnd cell_6t
Xbit_r261_c50 bl[50] br[50] wl[261] vdd gnd cell_6t
Xbit_r262_c50 bl[50] br[50] wl[262] vdd gnd cell_6t
Xbit_r263_c50 bl[50] br[50] wl[263] vdd gnd cell_6t
Xbit_r264_c50 bl[50] br[50] wl[264] vdd gnd cell_6t
Xbit_r265_c50 bl[50] br[50] wl[265] vdd gnd cell_6t
Xbit_r266_c50 bl[50] br[50] wl[266] vdd gnd cell_6t
Xbit_r267_c50 bl[50] br[50] wl[267] vdd gnd cell_6t
Xbit_r268_c50 bl[50] br[50] wl[268] vdd gnd cell_6t
Xbit_r269_c50 bl[50] br[50] wl[269] vdd gnd cell_6t
Xbit_r270_c50 bl[50] br[50] wl[270] vdd gnd cell_6t
Xbit_r271_c50 bl[50] br[50] wl[271] vdd gnd cell_6t
Xbit_r272_c50 bl[50] br[50] wl[272] vdd gnd cell_6t
Xbit_r273_c50 bl[50] br[50] wl[273] vdd gnd cell_6t
Xbit_r274_c50 bl[50] br[50] wl[274] vdd gnd cell_6t
Xbit_r275_c50 bl[50] br[50] wl[275] vdd gnd cell_6t
Xbit_r276_c50 bl[50] br[50] wl[276] vdd gnd cell_6t
Xbit_r277_c50 bl[50] br[50] wl[277] vdd gnd cell_6t
Xbit_r278_c50 bl[50] br[50] wl[278] vdd gnd cell_6t
Xbit_r279_c50 bl[50] br[50] wl[279] vdd gnd cell_6t
Xbit_r280_c50 bl[50] br[50] wl[280] vdd gnd cell_6t
Xbit_r281_c50 bl[50] br[50] wl[281] vdd gnd cell_6t
Xbit_r282_c50 bl[50] br[50] wl[282] vdd gnd cell_6t
Xbit_r283_c50 bl[50] br[50] wl[283] vdd gnd cell_6t
Xbit_r284_c50 bl[50] br[50] wl[284] vdd gnd cell_6t
Xbit_r285_c50 bl[50] br[50] wl[285] vdd gnd cell_6t
Xbit_r286_c50 bl[50] br[50] wl[286] vdd gnd cell_6t
Xbit_r287_c50 bl[50] br[50] wl[287] vdd gnd cell_6t
Xbit_r288_c50 bl[50] br[50] wl[288] vdd gnd cell_6t
Xbit_r289_c50 bl[50] br[50] wl[289] vdd gnd cell_6t
Xbit_r290_c50 bl[50] br[50] wl[290] vdd gnd cell_6t
Xbit_r291_c50 bl[50] br[50] wl[291] vdd gnd cell_6t
Xbit_r292_c50 bl[50] br[50] wl[292] vdd gnd cell_6t
Xbit_r293_c50 bl[50] br[50] wl[293] vdd gnd cell_6t
Xbit_r294_c50 bl[50] br[50] wl[294] vdd gnd cell_6t
Xbit_r295_c50 bl[50] br[50] wl[295] vdd gnd cell_6t
Xbit_r296_c50 bl[50] br[50] wl[296] vdd gnd cell_6t
Xbit_r297_c50 bl[50] br[50] wl[297] vdd gnd cell_6t
Xbit_r298_c50 bl[50] br[50] wl[298] vdd gnd cell_6t
Xbit_r299_c50 bl[50] br[50] wl[299] vdd gnd cell_6t
Xbit_r300_c50 bl[50] br[50] wl[300] vdd gnd cell_6t
Xbit_r301_c50 bl[50] br[50] wl[301] vdd gnd cell_6t
Xbit_r302_c50 bl[50] br[50] wl[302] vdd gnd cell_6t
Xbit_r303_c50 bl[50] br[50] wl[303] vdd gnd cell_6t
Xbit_r304_c50 bl[50] br[50] wl[304] vdd gnd cell_6t
Xbit_r305_c50 bl[50] br[50] wl[305] vdd gnd cell_6t
Xbit_r306_c50 bl[50] br[50] wl[306] vdd gnd cell_6t
Xbit_r307_c50 bl[50] br[50] wl[307] vdd gnd cell_6t
Xbit_r308_c50 bl[50] br[50] wl[308] vdd gnd cell_6t
Xbit_r309_c50 bl[50] br[50] wl[309] vdd gnd cell_6t
Xbit_r310_c50 bl[50] br[50] wl[310] vdd gnd cell_6t
Xbit_r311_c50 bl[50] br[50] wl[311] vdd gnd cell_6t
Xbit_r312_c50 bl[50] br[50] wl[312] vdd gnd cell_6t
Xbit_r313_c50 bl[50] br[50] wl[313] vdd gnd cell_6t
Xbit_r314_c50 bl[50] br[50] wl[314] vdd gnd cell_6t
Xbit_r315_c50 bl[50] br[50] wl[315] vdd gnd cell_6t
Xbit_r316_c50 bl[50] br[50] wl[316] vdd gnd cell_6t
Xbit_r317_c50 bl[50] br[50] wl[317] vdd gnd cell_6t
Xbit_r318_c50 bl[50] br[50] wl[318] vdd gnd cell_6t
Xbit_r319_c50 bl[50] br[50] wl[319] vdd gnd cell_6t
Xbit_r320_c50 bl[50] br[50] wl[320] vdd gnd cell_6t
Xbit_r321_c50 bl[50] br[50] wl[321] vdd gnd cell_6t
Xbit_r322_c50 bl[50] br[50] wl[322] vdd gnd cell_6t
Xbit_r323_c50 bl[50] br[50] wl[323] vdd gnd cell_6t
Xbit_r324_c50 bl[50] br[50] wl[324] vdd gnd cell_6t
Xbit_r325_c50 bl[50] br[50] wl[325] vdd gnd cell_6t
Xbit_r326_c50 bl[50] br[50] wl[326] vdd gnd cell_6t
Xbit_r327_c50 bl[50] br[50] wl[327] vdd gnd cell_6t
Xbit_r328_c50 bl[50] br[50] wl[328] vdd gnd cell_6t
Xbit_r329_c50 bl[50] br[50] wl[329] vdd gnd cell_6t
Xbit_r330_c50 bl[50] br[50] wl[330] vdd gnd cell_6t
Xbit_r331_c50 bl[50] br[50] wl[331] vdd gnd cell_6t
Xbit_r332_c50 bl[50] br[50] wl[332] vdd gnd cell_6t
Xbit_r333_c50 bl[50] br[50] wl[333] vdd gnd cell_6t
Xbit_r334_c50 bl[50] br[50] wl[334] vdd gnd cell_6t
Xbit_r335_c50 bl[50] br[50] wl[335] vdd gnd cell_6t
Xbit_r336_c50 bl[50] br[50] wl[336] vdd gnd cell_6t
Xbit_r337_c50 bl[50] br[50] wl[337] vdd gnd cell_6t
Xbit_r338_c50 bl[50] br[50] wl[338] vdd gnd cell_6t
Xbit_r339_c50 bl[50] br[50] wl[339] vdd gnd cell_6t
Xbit_r340_c50 bl[50] br[50] wl[340] vdd gnd cell_6t
Xbit_r341_c50 bl[50] br[50] wl[341] vdd gnd cell_6t
Xbit_r342_c50 bl[50] br[50] wl[342] vdd gnd cell_6t
Xbit_r343_c50 bl[50] br[50] wl[343] vdd gnd cell_6t
Xbit_r344_c50 bl[50] br[50] wl[344] vdd gnd cell_6t
Xbit_r345_c50 bl[50] br[50] wl[345] vdd gnd cell_6t
Xbit_r346_c50 bl[50] br[50] wl[346] vdd gnd cell_6t
Xbit_r347_c50 bl[50] br[50] wl[347] vdd gnd cell_6t
Xbit_r348_c50 bl[50] br[50] wl[348] vdd gnd cell_6t
Xbit_r349_c50 bl[50] br[50] wl[349] vdd gnd cell_6t
Xbit_r350_c50 bl[50] br[50] wl[350] vdd gnd cell_6t
Xbit_r351_c50 bl[50] br[50] wl[351] vdd gnd cell_6t
Xbit_r352_c50 bl[50] br[50] wl[352] vdd gnd cell_6t
Xbit_r353_c50 bl[50] br[50] wl[353] vdd gnd cell_6t
Xbit_r354_c50 bl[50] br[50] wl[354] vdd gnd cell_6t
Xbit_r355_c50 bl[50] br[50] wl[355] vdd gnd cell_6t
Xbit_r356_c50 bl[50] br[50] wl[356] vdd gnd cell_6t
Xbit_r357_c50 bl[50] br[50] wl[357] vdd gnd cell_6t
Xbit_r358_c50 bl[50] br[50] wl[358] vdd gnd cell_6t
Xbit_r359_c50 bl[50] br[50] wl[359] vdd gnd cell_6t
Xbit_r360_c50 bl[50] br[50] wl[360] vdd gnd cell_6t
Xbit_r361_c50 bl[50] br[50] wl[361] vdd gnd cell_6t
Xbit_r362_c50 bl[50] br[50] wl[362] vdd gnd cell_6t
Xbit_r363_c50 bl[50] br[50] wl[363] vdd gnd cell_6t
Xbit_r364_c50 bl[50] br[50] wl[364] vdd gnd cell_6t
Xbit_r365_c50 bl[50] br[50] wl[365] vdd gnd cell_6t
Xbit_r366_c50 bl[50] br[50] wl[366] vdd gnd cell_6t
Xbit_r367_c50 bl[50] br[50] wl[367] vdd gnd cell_6t
Xbit_r368_c50 bl[50] br[50] wl[368] vdd gnd cell_6t
Xbit_r369_c50 bl[50] br[50] wl[369] vdd gnd cell_6t
Xbit_r370_c50 bl[50] br[50] wl[370] vdd gnd cell_6t
Xbit_r371_c50 bl[50] br[50] wl[371] vdd gnd cell_6t
Xbit_r372_c50 bl[50] br[50] wl[372] vdd gnd cell_6t
Xbit_r373_c50 bl[50] br[50] wl[373] vdd gnd cell_6t
Xbit_r374_c50 bl[50] br[50] wl[374] vdd gnd cell_6t
Xbit_r375_c50 bl[50] br[50] wl[375] vdd gnd cell_6t
Xbit_r376_c50 bl[50] br[50] wl[376] vdd gnd cell_6t
Xbit_r377_c50 bl[50] br[50] wl[377] vdd gnd cell_6t
Xbit_r378_c50 bl[50] br[50] wl[378] vdd gnd cell_6t
Xbit_r379_c50 bl[50] br[50] wl[379] vdd gnd cell_6t
Xbit_r380_c50 bl[50] br[50] wl[380] vdd gnd cell_6t
Xbit_r381_c50 bl[50] br[50] wl[381] vdd gnd cell_6t
Xbit_r382_c50 bl[50] br[50] wl[382] vdd gnd cell_6t
Xbit_r383_c50 bl[50] br[50] wl[383] vdd gnd cell_6t
Xbit_r384_c50 bl[50] br[50] wl[384] vdd gnd cell_6t
Xbit_r385_c50 bl[50] br[50] wl[385] vdd gnd cell_6t
Xbit_r386_c50 bl[50] br[50] wl[386] vdd gnd cell_6t
Xbit_r387_c50 bl[50] br[50] wl[387] vdd gnd cell_6t
Xbit_r388_c50 bl[50] br[50] wl[388] vdd gnd cell_6t
Xbit_r389_c50 bl[50] br[50] wl[389] vdd gnd cell_6t
Xbit_r390_c50 bl[50] br[50] wl[390] vdd gnd cell_6t
Xbit_r391_c50 bl[50] br[50] wl[391] vdd gnd cell_6t
Xbit_r392_c50 bl[50] br[50] wl[392] vdd gnd cell_6t
Xbit_r393_c50 bl[50] br[50] wl[393] vdd gnd cell_6t
Xbit_r394_c50 bl[50] br[50] wl[394] vdd gnd cell_6t
Xbit_r395_c50 bl[50] br[50] wl[395] vdd gnd cell_6t
Xbit_r396_c50 bl[50] br[50] wl[396] vdd gnd cell_6t
Xbit_r397_c50 bl[50] br[50] wl[397] vdd gnd cell_6t
Xbit_r398_c50 bl[50] br[50] wl[398] vdd gnd cell_6t
Xbit_r399_c50 bl[50] br[50] wl[399] vdd gnd cell_6t
Xbit_r400_c50 bl[50] br[50] wl[400] vdd gnd cell_6t
Xbit_r401_c50 bl[50] br[50] wl[401] vdd gnd cell_6t
Xbit_r402_c50 bl[50] br[50] wl[402] vdd gnd cell_6t
Xbit_r403_c50 bl[50] br[50] wl[403] vdd gnd cell_6t
Xbit_r404_c50 bl[50] br[50] wl[404] vdd gnd cell_6t
Xbit_r405_c50 bl[50] br[50] wl[405] vdd gnd cell_6t
Xbit_r406_c50 bl[50] br[50] wl[406] vdd gnd cell_6t
Xbit_r407_c50 bl[50] br[50] wl[407] vdd gnd cell_6t
Xbit_r408_c50 bl[50] br[50] wl[408] vdd gnd cell_6t
Xbit_r409_c50 bl[50] br[50] wl[409] vdd gnd cell_6t
Xbit_r410_c50 bl[50] br[50] wl[410] vdd gnd cell_6t
Xbit_r411_c50 bl[50] br[50] wl[411] vdd gnd cell_6t
Xbit_r412_c50 bl[50] br[50] wl[412] vdd gnd cell_6t
Xbit_r413_c50 bl[50] br[50] wl[413] vdd gnd cell_6t
Xbit_r414_c50 bl[50] br[50] wl[414] vdd gnd cell_6t
Xbit_r415_c50 bl[50] br[50] wl[415] vdd gnd cell_6t
Xbit_r416_c50 bl[50] br[50] wl[416] vdd gnd cell_6t
Xbit_r417_c50 bl[50] br[50] wl[417] vdd gnd cell_6t
Xbit_r418_c50 bl[50] br[50] wl[418] vdd gnd cell_6t
Xbit_r419_c50 bl[50] br[50] wl[419] vdd gnd cell_6t
Xbit_r420_c50 bl[50] br[50] wl[420] vdd gnd cell_6t
Xbit_r421_c50 bl[50] br[50] wl[421] vdd gnd cell_6t
Xbit_r422_c50 bl[50] br[50] wl[422] vdd gnd cell_6t
Xbit_r423_c50 bl[50] br[50] wl[423] vdd gnd cell_6t
Xbit_r424_c50 bl[50] br[50] wl[424] vdd gnd cell_6t
Xbit_r425_c50 bl[50] br[50] wl[425] vdd gnd cell_6t
Xbit_r426_c50 bl[50] br[50] wl[426] vdd gnd cell_6t
Xbit_r427_c50 bl[50] br[50] wl[427] vdd gnd cell_6t
Xbit_r428_c50 bl[50] br[50] wl[428] vdd gnd cell_6t
Xbit_r429_c50 bl[50] br[50] wl[429] vdd gnd cell_6t
Xbit_r430_c50 bl[50] br[50] wl[430] vdd gnd cell_6t
Xbit_r431_c50 bl[50] br[50] wl[431] vdd gnd cell_6t
Xbit_r432_c50 bl[50] br[50] wl[432] vdd gnd cell_6t
Xbit_r433_c50 bl[50] br[50] wl[433] vdd gnd cell_6t
Xbit_r434_c50 bl[50] br[50] wl[434] vdd gnd cell_6t
Xbit_r435_c50 bl[50] br[50] wl[435] vdd gnd cell_6t
Xbit_r436_c50 bl[50] br[50] wl[436] vdd gnd cell_6t
Xbit_r437_c50 bl[50] br[50] wl[437] vdd gnd cell_6t
Xbit_r438_c50 bl[50] br[50] wl[438] vdd gnd cell_6t
Xbit_r439_c50 bl[50] br[50] wl[439] vdd gnd cell_6t
Xbit_r440_c50 bl[50] br[50] wl[440] vdd gnd cell_6t
Xbit_r441_c50 bl[50] br[50] wl[441] vdd gnd cell_6t
Xbit_r442_c50 bl[50] br[50] wl[442] vdd gnd cell_6t
Xbit_r443_c50 bl[50] br[50] wl[443] vdd gnd cell_6t
Xbit_r444_c50 bl[50] br[50] wl[444] vdd gnd cell_6t
Xbit_r445_c50 bl[50] br[50] wl[445] vdd gnd cell_6t
Xbit_r446_c50 bl[50] br[50] wl[446] vdd gnd cell_6t
Xbit_r447_c50 bl[50] br[50] wl[447] vdd gnd cell_6t
Xbit_r448_c50 bl[50] br[50] wl[448] vdd gnd cell_6t
Xbit_r449_c50 bl[50] br[50] wl[449] vdd gnd cell_6t
Xbit_r450_c50 bl[50] br[50] wl[450] vdd gnd cell_6t
Xbit_r451_c50 bl[50] br[50] wl[451] vdd gnd cell_6t
Xbit_r452_c50 bl[50] br[50] wl[452] vdd gnd cell_6t
Xbit_r453_c50 bl[50] br[50] wl[453] vdd gnd cell_6t
Xbit_r454_c50 bl[50] br[50] wl[454] vdd gnd cell_6t
Xbit_r455_c50 bl[50] br[50] wl[455] vdd gnd cell_6t
Xbit_r456_c50 bl[50] br[50] wl[456] vdd gnd cell_6t
Xbit_r457_c50 bl[50] br[50] wl[457] vdd gnd cell_6t
Xbit_r458_c50 bl[50] br[50] wl[458] vdd gnd cell_6t
Xbit_r459_c50 bl[50] br[50] wl[459] vdd gnd cell_6t
Xbit_r460_c50 bl[50] br[50] wl[460] vdd gnd cell_6t
Xbit_r461_c50 bl[50] br[50] wl[461] vdd gnd cell_6t
Xbit_r462_c50 bl[50] br[50] wl[462] vdd gnd cell_6t
Xbit_r463_c50 bl[50] br[50] wl[463] vdd gnd cell_6t
Xbit_r464_c50 bl[50] br[50] wl[464] vdd gnd cell_6t
Xbit_r465_c50 bl[50] br[50] wl[465] vdd gnd cell_6t
Xbit_r466_c50 bl[50] br[50] wl[466] vdd gnd cell_6t
Xbit_r467_c50 bl[50] br[50] wl[467] vdd gnd cell_6t
Xbit_r468_c50 bl[50] br[50] wl[468] vdd gnd cell_6t
Xbit_r469_c50 bl[50] br[50] wl[469] vdd gnd cell_6t
Xbit_r470_c50 bl[50] br[50] wl[470] vdd gnd cell_6t
Xbit_r471_c50 bl[50] br[50] wl[471] vdd gnd cell_6t
Xbit_r472_c50 bl[50] br[50] wl[472] vdd gnd cell_6t
Xbit_r473_c50 bl[50] br[50] wl[473] vdd gnd cell_6t
Xbit_r474_c50 bl[50] br[50] wl[474] vdd gnd cell_6t
Xbit_r475_c50 bl[50] br[50] wl[475] vdd gnd cell_6t
Xbit_r476_c50 bl[50] br[50] wl[476] vdd gnd cell_6t
Xbit_r477_c50 bl[50] br[50] wl[477] vdd gnd cell_6t
Xbit_r478_c50 bl[50] br[50] wl[478] vdd gnd cell_6t
Xbit_r479_c50 bl[50] br[50] wl[479] vdd gnd cell_6t
Xbit_r480_c50 bl[50] br[50] wl[480] vdd gnd cell_6t
Xbit_r481_c50 bl[50] br[50] wl[481] vdd gnd cell_6t
Xbit_r482_c50 bl[50] br[50] wl[482] vdd gnd cell_6t
Xbit_r483_c50 bl[50] br[50] wl[483] vdd gnd cell_6t
Xbit_r484_c50 bl[50] br[50] wl[484] vdd gnd cell_6t
Xbit_r485_c50 bl[50] br[50] wl[485] vdd gnd cell_6t
Xbit_r486_c50 bl[50] br[50] wl[486] vdd gnd cell_6t
Xbit_r487_c50 bl[50] br[50] wl[487] vdd gnd cell_6t
Xbit_r488_c50 bl[50] br[50] wl[488] vdd gnd cell_6t
Xbit_r489_c50 bl[50] br[50] wl[489] vdd gnd cell_6t
Xbit_r490_c50 bl[50] br[50] wl[490] vdd gnd cell_6t
Xbit_r491_c50 bl[50] br[50] wl[491] vdd gnd cell_6t
Xbit_r492_c50 bl[50] br[50] wl[492] vdd gnd cell_6t
Xbit_r493_c50 bl[50] br[50] wl[493] vdd gnd cell_6t
Xbit_r494_c50 bl[50] br[50] wl[494] vdd gnd cell_6t
Xbit_r495_c50 bl[50] br[50] wl[495] vdd gnd cell_6t
Xbit_r496_c50 bl[50] br[50] wl[496] vdd gnd cell_6t
Xbit_r497_c50 bl[50] br[50] wl[497] vdd gnd cell_6t
Xbit_r498_c50 bl[50] br[50] wl[498] vdd gnd cell_6t
Xbit_r499_c50 bl[50] br[50] wl[499] vdd gnd cell_6t
Xbit_r500_c50 bl[50] br[50] wl[500] vdd gnd cell_6t
Xbit_r501_c50 bl[50] br[50] wl[501] vdd gnd cell_6t
Xbit_r502_c50 bl[50] br[50] wl[502] vdd gnd cell_6t
Xbit_r503_c50 bl[50] br[50] wl[503] vdd gnd cell_6t
Xbit_r504_c50 bl[50] br[50] wl[504] vdd gnd cell_6t
Xbit_r505_c50 bl[50] br[50] wl[505] vdd gnd cell_6t
Xbit_r506_c50 bl[50] br[50] wl[506] vdd gnd cell_6t
Xbit_r507_c50 bl[50] br[50] wl[507] vdd gnd cell_6t
Xbit_r508_c50 bl[50] br[50] wl[508] vdd gnd cell_6t
Xbit_r509_c50 bl[50] br[50] wl[509] vdd gnd cell_6t
Xbit_r510_c50 bl[50] br[50] wl[510] vdd gnd cell_6t
Xbit_r511_c50 bl[50] br[50] wl[511] vdd gnd cell_6t
Xbit_r0_c51 bl[51] br[51] wl[0] vdd gnd cell_6t
Xbit_r1_c51 bl[51] br[51] wl[1] vdd gnd cell_6t
Xbit_r2_c51 bl[51] br[51] wl[2] vdd gnd cell_6t
Xbit_r3_c51 bl[51] br[51] wl[3] vdd gnd cell_6t
Xbit_r4_c51 bl[51] br[51] wl[4] vdd gnd cell_6t
Xbit_r5_c51 bl[51] br[51] wl[5] vdd gnd cell_6t
Xbit_r6_c51 bl[51] br[51] wl[6] vdd gnd cell_6t
Xbit_r7_c51 bl[51] br[51] wl[7] vdd gnd cell_6t
Xbit_r8_c51 bl[51] br[51] wl[8] vdd gnd cell_6t
Xbit_r9_c51 bl[51] br[51] wl[9] vdd gnd cell_6t
Xbit_r10_c51 bl[51] br[51] wl[10] vdd gnd cell_6t
Xbit_r11_c51 bl[51] br[51] wl[11] vdd gnd cell_6t
Xbit_r12_c51 bl[51] br[51] wl[12] vdd gnd cell_6t
Xbit_r13_c51 bl[51] br[51] wl[13] vdd gnd cell_6t
Xbit_r14_c51 bl[51] br[51] wl[14] vdd gnd cell_6t
Xbit_r15_c51 bl[51] br[51] wl[15] vdd gnd cell_6t
Xbit_r16_c51 bl[51] br[51] wl[16] vdd gnd cell_6t
Xbit_r17_c51 bl[51] br[51] wl[17] vdd gnd cell_6t
Xbit_r18_c51 bl[51] br[51] wl[18] vdd gnd cell_6t
Xbit_r19_c51 bl[51] br[51] wl[19] vdd gnd cell_6t
Xbit_r20_c51 bl[51] br[51] wl[20] vdd gnd cell_6t
Xbit_r21_c51 bl[51] br[51] wl[21] vdd gnd cell_6t
Xbit_r22_c51 bl[51] br[51] wl[22] vdd gnd cell_6t
Xbit_r23_c51 bl[51] br[51] wl[23] vdd gnd cell_6t
Xbit_r24_c51 bl[51] br[51] wl[24] vdd gnd cell_6t
Xbit_r25_c51 bl[51] br[51] wl[25] vdd gnd cell_6t
Xbit_r26_c51 bl[51] br[51] wl[26] vdd gnd cell_6t
Xbit_r27_c51 bl[51] br[51] wl[27] vdd gnd cell_6t
Xbit_r28_c51 bl[51] br[51] wl[28] vdd gnd cell_6t
Xbit_r29_c51 bl[51] br[51] wl[29] vdd gnd cell_6t
Xbit_r30_c51 bl[51] br[51] wl[30] vdd gnd cell_6t
Xbit_r31_c51 bl[51] br[51] wl[31] vdd gnd cell_6t
Xbit_r32_c51 bl[51] br[51] wl[32] vdd gnd cell_6t
Xbit_r33_c51 bl[51] br[51] wl[33] vdd gnd cell_6t
Xbit_r34_c51 bl[51] br[51] wl[34] vdd gnd cell_6t
Xbit_r35_c51 bl[51] br[51] wl[35] vdd gnd cell_6t
Xbit_r36_c51 bl[51] br[51] wl[36] vdd gnd cell_6t
Xbit_r37_c51 bl[51] br[51] wl[37] vdd gnd cell_6t
Xbit_r38_c51 bl[51] br[51] wl[38] vdd gnd cell_6t
Xbit_r39_c51 bl[51] br[51] wl[39] vdd gnd cell_6t
Xbit_r40_c51 bl[51] br[51] wl[40] vdd gnd cell_6t
Xbit_r41_c51 bl[51] br[51] wl[41] vdd gnd cell_6t
Xbit_r42_c51 bl[51] br[51] wl[42] vdd gnd cell_6t
Xbit_r43_c51 bl[51] br[51] wl[43] vdd gnd cell_6t
Xbit_r44_c51 bl[51] br[51] wl[44] vdd gnd cell_6t
Xbit_r45_c51 bl[51] br[51] wl[45] vdd gnd cell_6t
Xbit_r46_c51 bl[51] br[51] wl[46] vdd gnd cell_6t
Xbit_r47_c51 bl[51] br[51] wl[47] vdd gnd cell_6t
Xbit_r48_c51 bl[51] br[51] wl[48] vdd gnd cell_6t
Xbit_r49_c51 bl[51] br[51] wl[49] vdd gnd cell_6t
Xbit_r50_c51 bl[51] br[51] wl[50] vdd gnd cell_6t
Xbit_r51_c51 bl[51] br[51] wl[51] vdd gnd cell_6t
Xbit_r52_c51 bl[51] br[51] wl[52] vdd gnd cell_6t
Xbit_r53_c51 bl[51] br[51] wl[53] vdd gnd cell_6t
Xbit_r54_c51 bl[51] br[51] wl[54] vdd gnd cell_6t
Xbit_r55_c51 bl[51] br[51] wl[55] vdd gnd cell_6t
Xbit_r56_c51 bl[51] br[51] wl[56] vdd gnd cell_6t
Xbit_r57_c51 bl[51] br[51] wl[57] vdd gnd cell_6t
Xbit_r58_c51 bl[51] br[51] wl[58] vdd gnd cell_6t
Xbit_r59_c51 bl[51] br[51] wl[59] vdd gnd cell_6t
Xbit_r60_c51 bl[51] br[51] wl[60] vdd gnd cell_6t
Xbit_r61_c51 bl[51] br[51] wl[61] vdd gnd cell_6t
Xbit_r62_c51 bl[51] br[51] wl[62] vdd gnd cell_6t
Xbit_r63_c51 bl[51] br[51] wl[63] vdd gnd cell_6t
Xbit_r64_c51 bl[51] br[51] wl[64] vdd gnd cell_6t
Xbit_r65_c51 bl[51] br[51] wl[65] vdd gnd cell_6t
Xbit_r66_c51 bl[51] br[51] wl[66] vdd gnd cell_6t
Xbit_r67_c51 bl[51] br[51] wl[67] vdd gnd cell_6t
Xbit_r68_c51 bl[51] br[51] wl[68] vdd gnd cell_6t
Xbit_r69_c51 bl[51] br[51] wl[69] vdd gnd cell_6t
Xbit_r70_c51 bl[51] br[51] wl[70] vdd gnd cell_6t
Xbit_r71_c51 bl[51] br[51] wl[71] vdd gnd cell_6t
Xbit_r72_c51 bl[51] br[51] wl[72] vdd gnd cell_6t
Xbit_r73_c51 bl[51] br[51] wl[73] vdd gnd cell_6t
Xbit_r74_c51 bl[51] br[51] wl[74] vdd gnd cell_6t
Xbit_r75_c51 bl[51] br[51] wl[75] vdd gnd cell_6t
Xbit_r76_c51 bl[51] br[51] wl[76] vdd gnd cell_6t
Xbit_r77_c51 bl[51] br[51] wl[77] vdd gnd cell_6t
Xbit_r78_c51 bl[51] br[51] wl[78] vdd gnd cell_6t
Xbit_r79_c51 bl[51] br[51] wl[79] vdd gnd cell_6t
Xbit_r80_c51 bl[51] br[51] wl[80] vdd gnd cell_6t
Xbit_r81_c51 bl[51] br[51] wl[81] vdd gnd cell_6t
Xbit_r82_c51 bl[51] br[51] wl[82] vdd gnd cell_6t
Xbit_r83_c51 bl[51] br[51] wl[83] vdd gnd cell_6t
Xbit_r84_c51 bl[51] br[51] wl[84] vdd gnd cell_6t
Xbit_r85_c51 bl[51] br[51] wl[85] vdd gnd cell_6t
Xbit_r86_c51 bl[51] br[51] wl[86] vdd gnd cell_6t
Xbit_r87_c51 bl[51] br[51] wl[87] vdd gnd cell_6t
Xbit_r88_c51 bl[51] br[51] wl[88] vdd gnd cell_6t
Xbit_r89_c51 bl[51] br[51] wl[89] vdd gnd cell_6t
Xbit_r90_c51 bl[51] br[51] wl[90] vdd gnd cell_6t
Xbit_r91_c51 bl[51] br[51] wl[91] vdd gnd cell_6t
Xbit_r92_c51 bl[51] br[51] wl[92] vdd gnd cell_6t
Xbit_r93_c51 bl[51] br[51] wl[93] vdd gnd cell_6t
Xbit_r94_c51 bl[51] br[51] wl[94] vdd gnd cell_6t
Xbit_r95_c51 bl[51] br[51] wl[95] vdd gnd cell_6t
Xbit_r96_c51 bl[51] br[51] wl[96] vdd gnd cell_6t
Xbit_r97_c51 bl[51] br[51] wl[97] vdd gnd cell_6t
Xbit_r98_c51 bl[51] br[51] wl[98] vdd gnd cell_6t
Xbit_r99_c51 bl[51] br[51] wl[99] vdd gnd cell_6t
Xbit_r100_c51 bl[51] br[51] wl[100] vdd gnd cell_6t
Xbit_r101_c51 bl[51] br[51] wl[101] vdd gnd cell_6t
Xbit_r102_c51 bl[51] br[51] wl[102] vdd gnd cell_6t
Xbit_r103_c51 bl[51] br[51] wl[103] vdd gnd cell_6t
Xbit_r104_c51 bl[51] br[51] wl[104] vdd gnd cell_6t
Xbit_r105_c51 bl[51] br[51] wl[105] vdd gnd cell_6t
Xbit_r106_c51 bl[51] br[51] wl[106] vdd gnd cell_6t
Xbit_r107_c51 bl[51] br[51] wl[107] vdd gnd cell_6t
Xbit_r108_c51 bl[51] br[51] wl[108] vdd gnd cell_6t
Xbit_r109_c51 bl[51] br[51] wl[109] vdd gnd cell_6t
Xbit_r110_c51 bl[51] br[51] wl[110] vdd gnd cell_6t
Xbit_r111_c51 bl[51] br[51] wl[111] vdd gnd cell_6t
Xbit_r112_c51 bl[51] br[51] wl[112] vdd gnd cell_6t
Xbit_r113_c51 bl[51] br[51] wl[113] vdd gnd cell_6t
Xbit_r114_c51 bl[51] br[51] wl[114] vdd gnd cell_6t
Xbit_r115_c51 bl[51] br[51] wl[115] vdd gnd cell_6t
Xbit_r116_c51 bl[51] br[51] wl[116] vdd gnd cell_6t
Xbit_r117_c51 bl[51] br[51] wl[117] vdd gnd cell_6t
Xbit_r118_c51 bl[51] br[51] wl[118] vdd gnd cell_6t
Xbit_r119_c51 bl[51] br[51] wl[119] vdd gnd cell_6t
Xbit_r120_c51 bl[51] br[51] wl[120] vdd gnd cell_6t
Xbit_r121_c51 bl[51] br[51] wl[121] vdd gnd cell_6t
Xbit_r122_c51 bl[51] br[51] wl[122] vdd gnd cell_6t
Xbit_r123_c51 bl[51] br[51] wl[123] vdd gnd cell_6t
Xbit_r124_c51 bl[51] br[51] wl[124] vdd gnd cell_6t
Xbit_r125_c51 bl[51] br[51] wl[125] vdd gnd cell_6t
Xbit_r126_c51 bl[51] br[51] wl[126] vdd gnd cell_6t
Xbit_r127_c51 bl[51] br[51] wl[127] vdd gnd cell_6t
Xbit_r128_c51 bl[51] br[51] wl[128] vdd gnd cell_6t
Xbit_r129_c51 bl[51] br[51] wl[129] vdd gnd cell_6t
Xbit_r130_c51 bl[51] br[51] wl[130] vdd gnd cell_6t
Xbit_r131_c51 bl[51] br[51] wl[131] vdd gnd cell_6t
Xbit_r132_c51 bl[51] br[51] wl[132] vdd gnd cell_6t
Xbit_r133_c51 bl[51] br[51] wl[133] vdd gnd cell_6t
Xbit_r134_c51 bl[51] br[51] wl[134] vdd gnd cell_6t
Xbit_r135_c51 bl[51] br[51] wl[135] vdd gnd cell_6t
Xbit_r136_c51 bl[51] br[51] wl[136] vdd gnd cell_6t
Xbit_r137_c51 bl[51] br[51] wl[137] vdd gnd cell_6t
Xbit_r138_c51 bl[51] br[51] wl[138] vdd gnd cell_6t
Xbit_r139_c51 bl[51] br[51] wl[139] vdd gnd cell_6t
Xbit_r140_c51 bl[51] br[51] wl[140] vdd gnd cell_6t
Xbit_r141_c51 bl[51] br[51] wl[141] vdd gnd cell_6t
Xbit_r142_c51 bl[51] br[51] wl[142] vdd gnd cell_6t
Xbit_r143_c51 bl[51] br[51] wl[143] vdd gnd cell_6t
Xbit_r144_c51 bl[51] br[51] wl[144] vdd gnd cell_6t
Xbit_r145_c51 bl[51] br[51] wl[145] vdd gnd cell_6t
Xbit_r146_c51 bl[51] br[51] wl[146] vdd gnd cell_6t
Xbit_r147_c51 bl[51] br[51] wl[147] vdd gnd cell_6t
Xbit_r148_c51 bl[51] br[51] wl[148] vdd gnd cell_6t
Xbit_r149_c51 bl[51] br[51] wl[149] vdd gnd cell_6t
Xbit_r150_c51 bl[51] br[51] wl[150] vdd gnd cell_6t
Xbit_r151_c51 bl[51] br[51] wl[151] vdd gnd cell_6t
Xbit_r152_c51 bl[51] br[51] wl[152] vdd gnd cell_6t
Xbit_r153_c51 bl[51] br[51] wl[153] vdd gnd cell_6t
Xbit_r154_c51 bl[51] br[51] wl[154] vdd gnd cell_6t
Xbit_r155_c51 bl[51] br[51] wl[155] vdd gnd cell_6t
Xbit_r156_c51 bl[51] br[51] wl[156] vdd gnd cell_6t
Xbit_r157_c51 bl[51] br[51] wl[157] vdd gnd cell_6t
Xbit_r158_c51 bl[51] br[51] wl[158] vdd gnd cell_6t
Xbit_r159_c51 bl[51] br[51] wl[159] vdd gnd cell_6t
Xbit_r160_c51 bl[51] br[51] wl[160] vdd gnd cell_6t
Xbit_r161_c51 bl[51] br[51] wl[161] vdd gnd cell_6t
Xbit_r162_c51 bl[51] br[51] wl[162] vdd gnd cell_6t
Xbit_r163_c51 bl[51] br[51] wl[163] vdd gnd cell_6t
Xbit_r164_c51 bl[51] br[51] wl[164] vdd gnd cell_6t
Xbit_r165_c51 bl[51] br[51] wl[165] vdd gnd cell_6t
Xbit_r166_c51 bl[51] br[51] wl[166] vdd gnd cell_6t
Xbit_r167_c51 bl[51] br[51] wl[167] vdd gnd cell_6t
Xbit_r168_c51 bl[51] br[51] wl[168] vdd gnd cell_6t
Xbit_r169_c51 bl[51] br[51] wl[169] vdd gnd cell_6t
Xbit_r170_c51 bl[51] br[51] wl[170] vdd gnd cell_6t
Xbit_r171_c51 bl[51] br[51] wl[171] vdd gnd cell_6t
Xbit_r172_c51 bl[51] br[51] wl[172] vdd gnd cell_6t
Xbit_r173_c51 bl[51] br[51] wl[173] vdd gnd cell_6t
Xbit_r174_c51 bl[51] br[51] wl[174] vdd gnd cell_6t
Xbit_r175_c51 bl[51] br[51] wl[175] vdd gnd cell_6t
Xbit_r176_c51 bl[51] br[51] wl[176] vdd gnd cell_6t
Xbit_r177_c51 bl[51] br[51] wl[177] vdd gnd cell_6t
Xbit_r178_c51 bl[51] br[51] wl[178] vdd gnd cell_6t
Xbit_r179_c51 bl[51] br[51] wl[179] vdd gnd cell_6t
Xbit_r180_c51 bl[51] br[51] wl[180] vdd gnd cell_6t
Xbit_r181_c51 bl[51] br[51] wl[181] vdd gnd cell_6t
Xbit_r182_c51 bl[51] br[51] wl[182] vdd gnd cell_6t
Xbit_r183_c51 bl[51] br[51] wl[183] vdd gnd cell_6t
Xbit_r184_c51 bl[51] br[51] wl[184] vdd gnd cell_6t
Xbit_r185_c51 bl[51] br[51] wl[185] vdd gnd cell_6t
Xbit_r186_c51 bl[51] br[51] wl[186] vdd gnd cell_6t
Xbit_r187_c51 bl[51] br[51] wl[187] vdd gnd cell_6t
Xbit_r188_c51 bl[51] br[51] wl[188] vdd gnd cell_6t
Xbit_r189_c51 bl[51] br[51] wl[189] vdd gnd cell_6t
Xbit_r190_c51 bl[51] br[51] wl[190] vdd gnd cell_6t
Xbit_r191_c51 bl[51] br[51] wl[191] vdd gnd cell_6t
Xbit_r192_c51 bl[51] br[51] wl[192] vdd gnd cell_6t
Xbit_r193_c51 bl[51] br[51] wl[193] vdd gnd cell_6t
Xbit_r194_c51 bl[51] br[51] wl[194] vdd gnd cell_6t
Xbit_r195_c51 bl[51] br[51] wl[195] vdd gnd cell_6t
Xbit_r196_c51 bl[51] br[51] wl[196] vdd gnd cell_6t
Xbit_r197_c51 bl[51] br[51] wl[197] vdd gnd cell_6t
Xbit_r198_c51 bl[51] br[51] wl[198] vdd gnd cell_6t
Xbit_r199_c51 bl[51] br[51] wl[199] vdd gnd cell_6t
Xbit_r200_c51 bl[51] br[51] wl[200] vdd gnd cell_6t
Xbit_r201_c51 bl[51] br[51] wl[201] vdd gnd cell_6t
Xbit_r202_c51 bl[51] br[51] wl[202] vdd gnd cell_6t
Xbit_r203_c51 bl[51] br[51] wl[203] vdd gnd cell_6t
Xbit_r204_c51 bl[51] br[51] wl[204] vdd gnd cell_6t
Xbit_r205_c51 bl[51] br[51] wl[205] vdd gnd cell_6t
Xbit_r206_c51 bl[51] br[51] wl[206] vdd gnd cell_6t
Xbit_r207_c51 bl[51] br[51] wl[207] vdd gnd cell_6t
Xbit_r208_c51 bl[51] br[51] wl[208] vdd gnd cell_6t
Xbit_r209_c51 bl[51] br[51] wl[209] vdd gnd cell_6t
Xbit_r210_c51 bl[51] br[51] wl[210] vdd gnd cell_6t
Xbit_r211_c51 bl[51] br[51] wl[211] vdd gnd cell_6t
Xbit_r212_c51 bl[51] br[51] wl[212] vdd gnd cell_6t
Xbit_r213_c51 bl[51] br[51] wl[213] vdd gnd cell_6t
Xbit_r214_c51 bl[51] br[51] wl[214] vdd gnd cell_6t
Xbit_r215_c51 bl[51] br[51] wl[215] vdd gnd cell_6t
Xbit_r216_c51 bl[51] br[51] wl[216] vdd gnd cell_6t
Xbit_r217_c51 bl[51] br[51] wl[217] vdd gnd cell_6t
Xbit_r218_c51 bl[51] br[51] wl[218] vdd gnd cell_6t
Xbit_r219_c51 bl[51] br[51] wl[219] vdd gnd cell_6t
Xbit_r220_c51 bl[51] br[51] wl[220] vdd gnd cell_6t
Xbit_r221_c51 bl[51] br[51] wl[221] vdd gnd cell_6t
Xbit_r222_c51 bl[51] br[51] wl[222] vdd gnd cell_6t
Xbit_r223_c51 bl[51] br[51] wl[223] vdd gnd cell_6t
Xbit_r224_c51 bl[51] br[51] wl[224] vdd gnd cell_6t
Xbit_r225_c51 bl[51] br[51] wl[225] vdd gnd cell_6t
Xbit_r226_c51 bl[51] br[51] wl[226] vdd gnd cell_6t
Xbit_r227_c51 bl[51] br[51] wl[227] vdd gnd cell_6t
Xbit_r228_c51 bl[51] br[51] wl[228] vdd gnd cell_6t
Xbit_r229_c51 bl[51] br[51] wl[229] vdd gnd cell_6t
Xbit_r230_c51 bl[51] br[51] wl[230] vdd gnd cell_6t
Xbit_r231_c51 bl[51] br[51] wl[231] vdd gnd cell_6t
Xbit_r232_c51 bl[51] br[51] wl[232] vdd gnd cell_6t
Xbit_r233_c51 bl[51] br[51] wl[233] vdd gnd cell_6t
Xbit_r234_c51 bl[51] br[51] wl[234] vdd gnd cell_6t
Xbit_r235_c51 bl[51] br[51] wl[235] vdd gnd cell_6t
Xbit_r236_c51 bl[51] br[51] wl[236] vdd gnd cell_6t
Xbit_r237_c51 bl[51] br[51] wl[237] vdd gnd cell_6t
Xbit_r238_c51 bl[51] br[51] wl[238] vdd gnd cell_6t
Xbit_r239_c51 bl[51] br[51] wl[239] vdd gnd cell_6t
Xbit_r240_c51 bl[51] br[51] wl[240] vdd gnd cell_6t
Xbit_r241_c51 bl[51] br[51] wl[241] vdd gnd cell_6t
Xbit_r242_c51 bl[51] br[51] wl[242] vdd gnd cell_6t
Xbit_r243_c51 bl[51] br[51] wl[243] vdd gnd cell_6t
Xbit_r244_c51 bl[51] br[51] wl[244] vdd gnd cell_6t
Xbit_r245_c51 bl[51] br[51] wl[245] vdd gnd cell_6t
Xbit_r246_c51 bl[51] br[51] wl[246] vdd gnd cell_6t
Xbit_r247_c51 bl[51] br[51] wl[247] vdd gnd cell_6t
Xbit_r248_c51 bl[51] br[51] wl[248] vdd gnd cell_6t
Xbit_r249_c51 bl[51] br[51] wl[249] vdd gnd cell_6t
Xbit_r250_c51 bl[51] br[51] wl[250] vdd gnd cell_6t
Xbit_r251_c51 bl[51] br[51] wl[251] vdd gnd cell_6t
Xbit_r252_c51 bl[51] br[51] wl[252] vdd gnd cell_6t
Xbit_r253_c51 bl[51] br[51] wl[253] vdd gnd cell_6t
Xbit_r254_c51 bl[51] br[51] wl[254] vdd gnd cell_6t
Xbit_r255_c51 bl[51] br[51] wl[255] vdd gnd cell_6t
Xbit_r256_c51 bl[51] br[51] wl[256] vdd gnd cell_6t
Xbit_r257_c51 bl[51] br[51] wl[257] vdd gnd cell_6t
Xbit_r258_c51 bl[51] br[51] wl[258] vdd gnd cell_6t
Xbit_r259_c51 bl[51] br[51] wl[259] vdd gnd cell_6t
Xbit_r260_c51 bl[51] br[51] wl[260] vdd gnd cell_6t
Xbit_r261_c51 bl[51] br[51] wl[261] vdd gnd cell_6t
Xbit_r262_c51 bl[51] br[51] wl[262] vdd gnd cell_6t
Xbit_r263_c51 bl[51] br[51] wl[263] vdd gnd cell_6t
Xbit_r264_c51 bl[51] br[51] wl[264] vdd gnd cell_6t
Xbit_r265_c51 bl[51] br[51] wl[265] vdd gnd cell_6t
Xbit_r266_c51 bl[51] br[51] wl[266] vdd gnd cell_6t
Xbit_r267_c51 bl[51] br[51] wl[267] vdd gnd cell_6t
Xbit_r268_c51 bl[51] br[51] wl[268] vdd gnd cell_6t
Xbit_r269_c51 bl[51] br[51] wl[269] vdd gnd cell_6t
Xbit_r270_c51 bl[51] br[51] wl[270] vdd gnd cell_6t
Xbit_r271_c51 bl[51] br[51] wl[271] vdd gnd cell_6t
Xbit_r272_c51 bl[51] br[51] wl[272] vdd gnd cell_6t
Xbit_r273_c51 bl[51] br[51] wl[273] vdd gnd cell_6t
Xbit_r274_c51 bl[51] br[51] wl[274] vdd gnd cell_6t
Xbit_r275_c51 bl[51] br[51] wl[275] vdd gnd cell_6t
Xbit_r276_c51 bl[51] br[51] wl[276] vdd gnd cell_6t
Xbit_r277_c51 bl[51] br[51] wl[277] vdd gnd cell_6t
Xbit_r278_c51 bl[51] br[51] wl[278] vdd gnd cell_6t
Xbit_r279_c51 bl[51] br[51] wl[279] vdd gnd cell_6t
Xbit_r280_c51 bl[51] br[51] wl[280] vdd gnd cell_6t
Xbit_r281_c51 bl[51] br[51] wl[281] vdd gnd cell_6t
Xbit_r282_c51 bl[51] br[51] wl[282] vdd gnd cell_6t
Xbit_r283_c51 bl[51] br[51] wl[283] vdd gnd cell_6t
Xbit_r284_c51 bl[51] br[51] wl[284] vdd gnd cell_6t
Xbit_r285_c51 bl[51] br[51] wl[285] vdd gnd cell_6t
Xbit_r286_c51 bl[51] br[51] wl[286] vdd gnd cell_6t
Xbit_r287_c51 bl[51] br[51] wl[287] vdd gnd cell_6t
Xbit_r288_c51 bl[51] br[51] wl[288] vdd gnd cell_6t
Xbit_r289_c51 bl[51] br[51] wl[289] vdd gnd cell_6t
Xbit_r290_c51 bl[51] br[51] wl[290] vdd gnd cell_6t
Xbit_r291_c51 bl[51] br[51] wl[291] vdd gnd cell_6t
Xbit_r292_c51 bl[51] br[51] wl[292] vdd gnd cell_6t
Xbit_r293_c51 bl[51] br[51] wl[293] vdd gnd cell_6t
Xbit_r294_c51 bl[51] br[51] wl[294] vdd gnd cell_6t
Xbit_r295_c51 bl[51] br[51] wl[295] vdd gnd cell_6t
Xbit_r296_c51 bl[51] br[51] wl[296] vdd gnd cell_6t
Xbit_r297_c51 bl[51] br[51] wl[297] vdd gnd cell_6t
Xbit_r298_c51 bl[51] br[51] wl[298] vdd gnd cell_6t
Xbit_r299_c51 bl[51] br[51] wl[299] vdd gnd cell_6t
Xbit_r300_c51 bl[51] br[51] wl[300] vdd gnd cell_6t
Xbit_r301_c51 bl[51] br[51] wl[301] vdd gnd cell_6t
Xbit_r302_c51 bl[51] br[51] wl[302] vdd gnd cell_6t
Xbit_r303_c51 bl[51] br[51] wl[303] vdd gnd cell_6t
Xbit_r304_c51 bl[51] br[51] wl[304] vdd gnd cell_6t
Xbit_r305_c51 bl[51] br[51] wl[305] vdd gnd cell_6t
Xbit_r306_c51 bl[51] br[51] wl[306] vdd gnd cell_6t
Xbit_r307_c51 bl[51] br[51] wl[307] vdd gnd cell_6t
Xbit_r308_c51 bl[51] br[51] wl[308] vdd gnd cell_6t
Xbit_r309_c51 bl[51] br[51] wl[309] vdd gnd cell_6t
Xbit_r310_c51 bl[51] br[51] wl[310] vdd gnd cell_6t
Xbit_r311_c51 bl[51] br[51] wl[311] vdd gnd cell_6t
Xbit_r312_c51 bl[51] br[51] wl[312] vdd gnd cell_6t
Xbit_r313_c51 bl[51] br[51] wl[313] vdd gnd cell_6t
Xbit_r314_c51 bl[51] br[51] wl[314] vdd gnd cell_6t
Xbit_r315_c51 bl[51] br[51] wl[315] vdd gnd cell_6t
Xbit_r316_c51 bl[51] br[51] wl[316] vdd gnd cell_6t
Xbit_r317_c51 bl[51] br[51] wl[317] vdd gnd cell_6t
Xbit_r318_c51 bl[51] br[51] wl[318] vdd gnd cell_6t
Xbit_r319_c51 bl[51] br[51] wl[319] vdd gnd cell_6t
Xbit_r320_c51 bl[51] br[51] wl[320] vdd gnd cell_6t
Xbit_r321_c51 bl[51] br[51] wl[321] vdd gnd cell_6t
Xbit_r322_c51 bl[51] br[51] wl[322] vdd gnd cell_6t
Xbit_r323_c51 bl[51] br[51] wl[323] vdd gnd cell_6t
Xbit_r324_c51 bl[51] br[51] wl[324] vdd gnd cell_6t
Xbit_r325_c51 bl[51] br[51] wl[325] vdd gnd cell_6t
Xbit_r326_c51 bl[51] br[51] wl[326] vdd gnd cell_6t
Xbit_r327_c51 bl[51] br[51] wl[327] vdd gnd cell_6t
Xbit_r328_c51 bl[51] br[51] wl[328] vdd gnd cell_6t
Xbit_r329_c51 bl[51] br[51] wl[329] vdd gnd cell_6t
Xbit_r330_c51 bl[51] br[51] wl[330] vdd gnd cell_6t
Xbit_r331_c51 bl[51] br[51] wl[331] vdd gnd cell_6t
Xbit_r332_c51 bl[51] br[51] wl[332] vdd gnd cell_6t
Xbit_r333_c51 bl[51] br[51] wl[333] vdd gnd cell_6t
Xbit_r334_c51 bl[51] br[51] wl[334] vdd gnd cell_6t
Xbit_r335_c51 bl[51] br[51] wl[335] vdd gnd cell_6t
Xbit_r336_c51 bl[51] br[51] wl[336] vdd gnd cell_6t
Xbit_r337_c51 bl[51] br[51] wl[337] vdd gnd cell_6t
Xbit_r338_c51 bl[51] br[51] wl[338] vdd gnd cell_6t
Xbit_r339_c51 bl[51] br[51] wl[339] vdd gnd cell_6t
Xbit_r340_c51 bl[51] br[51] wl[340] vdd gnd cell_6t
Xbit_r341_c51 bl[51] br[51] wl[341] vdd gnd cell_6t
Xbit_r342_c51 bl[51] br[51] wl[342] vdd gnd cell_6t
Xbit_r343_c51 bl[51] br[51] wl[343] vdd gnd cell_6t
Xbit_r344_c51 bl[51] br[51] wl[344] vdd gnd cell_6t
Xbit_r345_c51 bl[51] br[51] wl[345] vdd gnd cell_6t
Xbit_r346_c51 bl[51] br[51] wl[346] vdd gnd cell_6t
Xbit_r347_c51 bl[51] br[51] wl[347] vdd gnd cell_6t
Xbit_r348_c51 bl[51] br[51] wl[348] vdd gnd cell_6t
Xbit_r349_c51 bl[51] br[51] wl[349] vdd gnd cell_6t
Xbit_r350_c51 bl[51] br[51] wl[350] vdd gnd cell_6t
Xbit_r351_c51 bl[51] br[51] wl[351] vdd gnd cell_6t
Xbit_r352_c51 bl[51] br[51] wl[352] vdd gnd cell_6t
Xbit_r353_c51 bl[51] br[51] wl[353] vdd gnd cell_6t
Xbit_r354_c51 bl[51] br[51] wl[354] vdd gnd cell_6t
Xbit_r355_c51 bl[51] br[51] wl[355] vdd gnd cell_6t
Xbit_r356_c51 bl[51] br[51] wl[356] vdd gnd cell_6t
Xbit_r357_c51 bl[51] br[51] wl[357] vdd gnd cell_6t
Xbit_r358_c51 bl[51] br[51] wl[358] vdd gnd cell_6t
Xbit_r359_c51 bl[51] br[51] wl[359] vdd gnd cell_6t
Xbit_r360_c51 bl[51] br[51] wl[360] vdd gnd cell_6t
Xbit_r361_c51 bl[51] br[51] wl[361] vdd gnd cell_6t
Xbit_r362_c51 bl[51] br[51] wl[362] vdd gnd cell_6t
Xbit_r363_c51 bl[51] br[51] wl[363] vdd gnd cell_6t
Xbit_r364_c51 bl[51] br[51] wl[364] vdd gnd cell_6t
Xbit_r365_c51 bl[51] br[51] wl[365] vdd gnd cell_6t
Xbit_r366_c51 bl[51] br[51] wl[366] vdd gnd cell_6t
Xbit_r367_c51 bl[51] br[51] wl[367] vdd gnd cell_6t
Xbit_r368_c51 bl[51] br[51] wl[368] vdd gnd cell_6t
Xbit_r369_c51 bl[51] br[51] wl[369] vdd gnd cell_6t
Xbit_r370_c51 bl[51] br[51] wl[370] vdd gnd cell_6t
Xbit_r371_c51 bl[51] br[51] wl[371] vdd gnd cell_6t
Xbit_r372_c51 bl[51] br[51] wl[372] vdd gnd cell_6t
Xbit_r373_c51 bl[51] br[51] wl[373] vdd gnd cell_6t
Xbit_r374_c51 bl[51] br[51] wl[374] vdd gnd cell_6t
Xbit_r375_c51 bl[51] br[51] wl[375] vdd gnd cell_6t
Xbit_r376_c51 bl[51] br[51] wl[376] vdd gnd cell_6t
Xbit_r377_c51 bl[51] br[51] wl[377] vdd gnd cell_6t
Xbit_r378_c51 bl[51] br[51] wl[378] vdd gnd cell_6t
Xbit_r379_c51 bl[51] br[51] wl[379] vdd gnd cell_6t
Xbit_r380_c51 bl[51] br[51] wl[380] vdd gnd cell_6t
Xbit_r381_c51 bl[51] br[51] wl[381] vdd gnd cell_6t
Xbit_r382_c51 bl[51] br[51] wl[382] vdd gnd cell_6t
Xbit_r383_c51 bl[51] br[51] wl[383] vdd gnd cell_6t
Xbit_r384_c51 bl[51] br[51] wl[384] vdd gnd cell_6t
Xbit_r385_c51 bl[51] br[51] wl[385] vdd gnd cell_6t
Xbit_r386_c51 bl[51] br[51] wl[386] vdd gnd cell_6t
Xbit_r387_c51 bl[51] br[51] wl[387] vdd gnd cell_6t
Xbit_r388_c51 bl[51] br[51] wl[388] vdd gnd cell_6t
Xbit_r389_c51 bl[51] br[51] wl[389] vdd gnd cell_6t
Xbit_r390_c51 bl[51] br[51] wl[390] vdd gnd cell_6t
Xbit_r391_c51 bl[51] br[51] wl[391] vdd gnd cell_6t
Xbit_r392_c51 bl[51] br[51] wl[392] vdd gnd cell_6t
Xbit_r393_c51 bl[51] br[51] wl[393] vdd gnd cell_6t
Xbit_r394_c51 bl[51] br[51] wl[394] vdd gnd cell_6t
Xbit_r395_c51 bl[51] br[51] wl[395] vdd gnd cell_6t
Xbit_r396_c51 bl[51] br[51] wl[396] vdd gnd cell_6t
Xbit_r397_c51 bl[51] br[51] wl[397] vdd gnd cell_6t
Xbit_r398_c51 bl[51] br[51] wl[398] vdd gnd cell_6t
Xbit_r399_c51 bl[51] br[51] wl[399] vdd gnd cell_6t
Xbit_r400_c51 bl[51] br[51] wl[400] vdd gnd cell_6t
Xbit_r401_c51 bl[51] br[51] wl[401] vdd gnd cell_6t
Xbit_r402_c51 bl[51] br[51] wl[402] vdd gnd cell_6t
Xbit_r403_c51 bl[51] br[51] wl[403] vdd gnd cell_6t
Xbit_r404_c51 bl[51] br[51] wl[404] vdd gnd cell_6t
Xbit_r405_c51 bl[51] br[51] wl[405] vdd gnd cell_6t
Xbit_r406_c51 bl[51] br[51] wl[406] vdd gnd cell_6t
Xbit_r407_c51 bl[51] br[51] wl[407] vdd gnd cell_6t
Xbit_r408_c51 bl[51] br[51] wl[408] vdd gnd cell_6t
Xbit_r409_c51 bl[51] br[51] wl[409] vdd gnd cell_6t
Xbit_r410_c51 bl[51] br[51] wl[410] vdd gnd cell_6t
Xbit_r411_c51 bl[51] br[51] wl[411] vdd gnd cell_6t
Xbit_r412_c51 bl[51] br[51] wl[412] vdd gnd cell_6t
Xbit_r413_c51 bl[51] br[51] wl[413] vdd gnd cell_6t
Xbit_r414_c51 bl[51] br[51] wl[414] vdd gnd cell_6t
Xbit_r415_c51 bl[51] br[51] wl[415] vdd gnd cell_6t
Xbit_r416_c51 bl[51] br[51] wl[416] vdd gnd cell_6t
Xbit_r417_c51 bl[51] br[51] wl[417] vdd gnd cell_6t
Xbit_r418_c51 bl[51] br[51] wl[418] vdd gnd cell_6t
Xbit_r419_c51 bl[51] br[51] wl[419] vdd gnd cell_6t
Xbit_r420_c51 bl[51] br[51] wl[420] vdd gnd cell_6t
Xbit_r421_c51 bl[51] br[51] wl[421] vdd gnd cell_6t
Xbit_r422_c51 bl[51] br[51] wl[422] vdd gnd cell_6t
Xbit_r423_c51 bl[51] br[51] wl[423] vdd gnd cell_6t
Xbit_r424_c51 bl[51] br[51] wl[424] vdd gnd cell_6t
Xbit_r425_c51 bl[51] br[51] wl[425] vdd gnd cell_6t
Xbit_r426_c51 bl[51] br[51] wl[426] vdd gnd cell_6t
Xbit_r427_c51 bl[51] br[51] wl[427] vdd gnd cell_6t
Xbit_r428_c51 bl[51] br[51] wl[428] vdd gnd cell_6t
Xbit_r429_c51 bl[51] br[51] wl[429] vdd gnd cell_6t
Xbit_r430_c51 bl[51] br[51] wl[430] vdd gnd cell_6t
Xbit_r431_c51 bl[51] br[51] wl[431] vdd gnd cell_6t
Xbit_r432_c51 bl[51] br[51] wl[432] vdd gnd cell_6t
Xbit_r433_c51 bl[51] br[51] wl[433] vdd gnd cell_6t
Xbit_r434_c51 bl[51] br[51] wl[434] vdd gnd cell_6t
Xbit_r435_c51 bl[51] br[51] wl[435] vdd gnd cell_6t
Xbit_r436_c51 bl[51] br[51] wl[436] vdd gnd cell_6t
Xbit_r437_c51 bl[51] br[51] wl[437] vdd gnd cell_6t
Xbit_r438_c51 bl[51] br[51] wl[438] vdd gnd cell_6t
Xbit_r439_c51 bl[51] br[51] wl[439] vdd gnd cell_6t
Xbit_r440_c51 bl[51] br[51] wl[440] vdd gnd cell_6t
Xbit_r441_c51 bl[51] br[51] wl[441] vdd gnd cell_6t
Xbit_r442_c51 bl[51] br[51] wl[442] vdd gnd cell_6t
Xbit_r443_c51 bl[51] br[51] wl[443] vdd gnd cell_6t
Xbit_r444_c51 bl[51] br[51] wl[444] vdd gnd cell_6t
Xbit_r445_c51 bl[51] br[51] wl[445] vdd gnd cell_6t
Xbit_r446_c51 bl[51] br[51] wl[446] vdd gnd cell_6t
Xbit_r447_c51 bl[51] br[51] wl[447] vdd gnd cell_6t
Xbit_r448_c51 bl[51] br[51] wl[448] vdd gnd cell_6t
Xbit_r449_c51 bl[51] br[51] wl[449] vdd gnd cell_6t
Xbit_r450_c51 bl[51] br[51] wl[450] vdd gnd cell_6t
Xbit_r451_c51 bl[51] br[51] wl[451] vdd gnd cell_6t
Xbit_r452_c51 bl[51] br[51] wl[452] vdd gnd cell_6t
Xbit_r453_c51 bl[51] br[51] wl[453] vdd gnd cell_6t
Xbit_r454_c51 bl[51] br[51] wl[454] vdd gnd cell_6t
Xbit_r455_c51 bl[51] br[51] wl[455] vdd gnd cell_6t
Xbit_r456_c51 bl[51] br[51] wl[456] vdd gnd cell_6t
Xbit_r457_c51 bl[51] br[51] wl[457] vdd gnd cell_6t
Xbit_r458_c51 bl[51] br[51] wl[458] vdd gnd cell_6t
Xbit_r459_c51 bl[51] br[51] wl[459] vdd gnd cell_6t
Xbit_r460_c51 bl[51] br[51] wl[460] vdd gnd cell_6t
Xbit_r461_c51 bl[51] br[51] wl[461] vdd gnd cell_6t
Xbit_r462_c51 bl[51] br[51] wl[462] vdd gnd cell_6t
Xbit_r463_c51 bl[51] br[51] wl[463] vdd gnd cell_6t
Xbit_r464_c51 bl[51] br[51] wl[464] vdd gnd cell_6t
Xbit_r465_c51 bl[51] br[51] wl[465] vdd gnd cell_6t
Xbit_r466_c51 bl[51] br[51] wl[466] vdd gnd cell_6t
Xbit_r467_c51 bl[51] br[51] wl[467] vdd gnd cell_6t
Xbit_r468_c51 bl[51] br[51] wl[468] vdd gnd cell_6t
Xbit_r469_c51 bl[51] br[51] wl[469] vdd gnd cell_6t
Xbit_r470_c51 bl[51] br[51] wl[470] vdd gnd cell_6t
Xbit_r471_c51 bl[51] br[51] wl[471] vdd gnd cell_6t
Xbit_r472_c51 bl[51] br[51] wl[472] vdd gnd cell_6t
Xbit_r473_c51 bl[51] br[51] wl[473] vdd gnd cell_6t
Xbit_r474_c51 bl[51] br[51] wl[474] vdd gnd cell_6t
Xbit_r475_c51 bl[51] br[51] wl[475] vdd gnd cell_6t
Xbit_r476_c51 bl[51] br[51] wl[476] vdd gnd cell_6t
Xbit_r477_c51 bl[51] br[51] wl[477] vdd gnd cell_6t
Xbit_r478_c51 bl[51] br[51] wl[478] vdd gnd cell_6t
Xbit_r479_c51 bl[51] br[51] wl[479] vdd gnd cell_6t
Xbit_r480_c51 bl[51] br[51] wl[480] vdd gnd cell_6t
Xbit_r481_c51 bl[51] br[51] wl[481] vdd gnd cell_6t
Xbit_r482_c51 bl[51] br[51] wl[482] vdd gnd cell_6t
Xbit_r483_c51 bl[51] br[51] wl[483] vdd gnd cell_6t
Xbit_r484_c51 bl[51] br[51] wl[484] vdd gnd cell_6t
Xbit_r485_c51 bl[51] br[51] wl[485] vdd gnd cell_6t
Xbit_r486_c51 bl[51] br[51] wl[486] vdd gnd cell_6t
Xbit_r487_c51 bl[51] br[51] wl[487] vdd gnd cell_6t
Xbit_r488_c51 bl[51] br[51] wl[488] vdd gnd cell_6t
Xbit_r489_c51 bl[51] br[51] wl[489] vdd gnd cell_6t
Xbit_r490_c51 bl[51] br[51] wl[490] vdd gnd cell_6t
Xbit_r491_c51 bl[51] br[51] wl[491] vdd gnd cell_6t
Xbit_r492_c51 bl[51] br[51] wl[492] vdd gnd cell_6t
Xbit_r493_c51 bl[51] br[51] wl[493] vdd gnd cell_6t
Xbit_r494_c51 bl[51] br[51] wl[494] vdd gnd cell_6t
Xbit_r495_c51 bl[51] br[51] wl[495] vdd gnd cell_6t
Xbit_r496_c51 bl[51] br[51] wl[496] vdd gnd cell_6t
Xbit_r497_c51 bl[51] br[51] wl[497] vdd gnd cell_6t
Xbit_r498_c51 bl[51] br[51] wl[498] vdd gnd cell_6t
Xbit_r499_c51 bl[51] br[51] wl[499] vdd gnd cell_6t
Xbit_r500_c51 bl[51] br[51] wl[500] vdd gnd cell_6t
Xbit_r501_c51 bl[51] br[51] wl[501] vdd gnd cell_6t
Xbit_r502_c51 bl[51] br[51] wl[502] vdd gnd cell_6t
Xbit_r503_c51 bl[51] br[51] wl[503] vdd gnd cell_6t
Xbit_r504_c51 bl[51] br[51] wl[504] vdd gnd cell_6t
Xbit_r505_c51 bl[51] br[51] wl[505] vdd gnd cell_6t
Xbit_r506_c51 bl[51] br[51] wl[506] vdd gnd cell_6t
Xbit_r507_c51 bl[51] br[51] wl[507] vdd gnd cell_6t
Xbit_r508_c51 bl[51] br[51] wl[508] vdd gnd cell_6t
Xbit_r509_c51 bl[51] br[51] wl[509] vdd gnd cell_6t
Xbit_r510_c51 bl[51] br[51] wl[510] vdd gnd cell_6t
Xbit_r511_c51 bl[51] br[51] wl[511] vdd gnd cell_6t
Xbit_r0_c52 bl[52] br[52] wl[0] vdd gnd cell_6t
Xbit_r1_c52 bl[52] br[52] wl[1] vdd gnd cell_6t
Xbit_r2_c52 bl[52] br[52] wl[2] vdd gnd cell_6t
Xbit_r3_c52 bl[52] br[52] wl[3] vdd gnd cell_6t
Xbit_r4_c52 bl[52] br[52] wl[4] vdd gnd cell_6t
Xbit_r5_c52 bl[52] br[52] wl[5] vdd gnd cell_6t
Xbit_r6_c52 bl[52] br[52] wl[6] vdd gnd cell_6t
Xbit_r7_c52 bl[52] br[52] wl[7] vdd gnd cell_6t
Xbit_r8_c52 bl[52] br[52] wl[8] vdd gnd cell_6t
Xbit_r9_c52 bl[52] br[52] wl[9] vdd gnd cell_6t
Xbit_r10_c52 bl[52] br[52] wl[10] vdd gnd cell_6t
Xbit_r11_c52 bl[52] br[52] wl[11] vdd gnd cell_6t
Xbit_r12_c52 bl[52] br[52] wl[12] vdd gnd cell_6t
Xbit_r13_c52 bl[52] br[52] wl[13] vdd gnd cell_6t
Xbit_r14_c52 bl[52] br[52] wl[14] vdd gnd cell_6t
Xbit_r15_c52 bl[52] br[52] wl[15] vdd gnd cell_6t
Xbit_r16_c52 bl[52] br[52] wl[16] vdd gnd cell_6t
Xbit_r17_c52 bl[52] br[52] wl[17] vdd gnd cell_6t
Xbit_r18_c52 bl[52] br[52] wl[18] vdd gnd cell_6t
Xbit_r19_c52 bl[52] br[52] wl[19] vdd gnd cell_6t
Xbit_r20_c52 bl[52] br[52] wl[20] vdd gnd cell_6t
Xbit_r21_c52 bl[52] br[52] wl[21] vdd gnd cell_6t
Xbit_r22_c52 bl[52] br[52] wl[22] vdd gnd cell_6t
Xbit_r23_c52 bl[52] br[52] wl[23] vdd gnd cell_6t
Xbit_r24_c52 bl[52] br[52] wl[24] vdd gnd cell_6t
Xbit_r25_c52 bl[52] br[52] wl[25] vdd gnd cell_6t
Xbit_r26_c52 bl[52] br[52] wl[26] vdd gnd cell_6t
Xbit_r27_c52 bl[52] br[52] wl[27] vdd gnd cell_6t
Xbit_r28_c52 bl[52] br[52] wl[28] vdd gnd cell_6t
Xbit_r29_c52 bl[52] br[52] wl[29] vdd gnd cell_6t
Xbit_r30_c52 bl[52] br[52] wl[30] vdd gnd cell_6t
Xbit_r31_c52 bl[52] br[52] wl[31] vdd gnd cell_6t
Xbit_r32_c52 bl[52] br[52] wl[32] vdd gnd cell_6t
Xbit_r33_c52 bl[52] br[52] wl[33] vdd gnd cell_6t
Xbit_r34_c52 bl[52] br[52] wl[34] vdd gnd cell_6t
Xbit_r35_c52 bl[52] br[52] wl[35] vdd gnd cell_6t
Xbit_r36_c52 bl[52] br[52] wl[36] vdd gnd cell_6t
Xbit_r37_c52 bl[52] br[52] wl[37] vdd gnd cell_6t
Xbit_r38_c52 bl[52] br[52] wl[38] vdd gnd cell_6t
Xbit_r39_c52 bl[52] br[52] wl[39] vdd gnd cell_6t
Xbit_r40_c52 bl[52] br[52] wl[40] vdd gnd cell_6t
Xbit_r41_c52 bl[52] br[52] wl[41] vdd gnd cell_6t
Xbit_r42_c52 bl[52] br[52] wl[42] vdd gnd cell_6t
Xbit_r43_c52 bl[52] br[52] wl[43] vdd gnd cell_6t
Xbit_r44_c52 bl[52] br[52] wl[44] vdd gnd cell_6t
Xbit_r45_c52 bl[52] br[52] wl[45] vdd gnd cell_6t
Xbit_r46_c52 bl[52] br[52] wl[46] vdd gnd cell_6t
Xbit_r47_c52 bl[52] br[52] wl[47] vdd gnd cell_6t
Xbit_r48_c52 bl[52] br[52] wl[48] vdd gnd cell_6t
Xbit_r49_c52 bl[52] br[52] wl[49] vdd gnd cell_6t
Xbit_r50_c52 bl[52] br[52] wl[50] vdd gnd cell_6t
Xbit_r51_c52 bl[52] br[52] wl[51] vdd gnd cell_6t
Xbit_r52_c52 bl[52] br[52] wl[52] vdd gnd cell_6t
Xbit_r53_c52 bl[52] br[52] wl[53] vdd gnd cell_6t
Xbit_r54_c52 bl[52] br[52] wl[54] vdd gnd cell_6t
Xbit_r55_c52 bl[52] br[52] wl[55] vdd gnd cell_6t
Xbit_r56_c52 bl[52] br[52] wl[56] vdd gnd cell_6t
Xbit_r57_c52 bl[52] br[52] wl[57] vdd gnd cell_6t
Xbit_r58_c52 bl[52] br[52] wl[58] vdd gnd cell_6t
Xbit_r59_c52 bl[52] br[52] wl[59] vdd gnd cell_6t
Xbit_r60_c52 bl[52] br[52] wl[60] vdd gnd cell_6t
Xbit_r61_c52 bl[52] br[52] wl[61] vdd gnd cell_6t
Xbit_r62_c52 bl[52] br[52] wl[62] vdd gnd cell_6t
Xbit_r63_c52 bl[52] br[52] wl[63] vdd gnd cell_6t
Xbit_r64_c52 bl[52] br[52] wl[64] vdd gnd cell_6t
Xbit_r65_c52 bl[52] br[52] wl[65] vdd gnd cell_6t
Xbit_r66_c52 bl[52] br[52] wl[66] vdd gnd cell_6t
Xbit_r67_c52 bl[52] br[52] wl[67] vdd gnd cell_6t
Xbit_r68_c52 bl[52] br[52] wl[68] vdd gnd cell_6t
Xbit_r69_c52 bl[52] br[52] wl[69] vdd gnd cell_6t
Xbit_r70_c52 bl[52] br[52] wl[70] vdd gnd cell_6t
Xbit_r71_c52 bl[52] br[52] wl[71] vdd gnd cell_6t
Xbit_r72_c52 bl[52] br[52] wl[72] vdd gnd cell_6t
Xbit_r73_c52 bl[52] br[52] wl[73] vdd gnd cell_6t
Xbit_r74_c52 bl[52] br[52] wl[74] vdd gnd cell_6t
Xbit_r75_c52 bl[52] br[52] wl[75] vdd gnd cell_6t
Xbit_r76_c52 bl[52] br[52] wl[76] vdd gnd cell_6t
Xbit_r77_c52 bl[52] br[52] wl[77] vdd gnd cell_6t
Xbit_r78_c52 bl[52] br[52] wl[78] vdd gnd cell_6t
Xbit_r79_c52 bl[52] br[52] wl[79] vdd gnd cell_6t
Xbit_r80_c52 bl[52] br[52] wl[80] vdd gnd cell_6t
Xbit_r81_c52 bl[52] br[52] wl[81] vdd gnd cell_6t
Xbit_r82_c52 bl[52] br[52] wl[82] vdd gnd cell_6t
Xbit_r83_c52 bl[52] br[52] wl[83] vdd gnd cell_6t
Xbit_r84_c52 bl[52] br[52] wl[84] vdd gnd cell_6t
Xbit_r85_c52 bl[52] br[52] wl[85] vdd gnd cell_6t
Xbit_r86_c52 bl[52] br[52] wl[86] vdd gnd cell_6t
Xbit_r87_c52 bl[52] br[52] wl[87] vdd gnd cell_6t
Xbit_r88_c52 bl[52] br[52] wl[88] vdd gnd cell_6t
Xbit_r89_c52 bl[52] br[52] wl[89] vdd gnd cell_6t
Xbit_r90_c52 bl[52] br[52] wl[90] vdd gnd cell_6t
Xbit_r91_c52 bl[52] br[52] wl[91] vdd gnd cell_6t
Xbit_r92_c52 bl[52] br[52] wl[92] vdd gnd cell_6t
Xbit_r93_c52 bl[52] br[52] wl[93] vdd gnd cell_6t
Xbit_r94_c52 bl[52] br[52] wl[94] vdd gnd cell_6t
Xbit_r95_c52 bl[52] br[52] wl[95] vdd gnd cell_6t
Xbit_r96_c52 bl[52] br[52] wl[96] vdd gnd cell_6t
Xbit_r97_c52 bl[52] br[52] wl[97] vdd gnd cell_6t
Xbit_r98_c52 bl[52] br[52] wl[98] vdd gnd cell_6t
Xbit_r99_c52 bl[52] br[52] wl[99] vdd gnd cell_6t
Xbit_r100_c52 bl[52] br[52] wl[100] vdd gnd cell_6t
Xbit_r101_c52 bl[52] br[52] wl[101] vdd gnd cell_6t
Xbit_r102_c52 bl[52] br[52] wl[102] vdd gnd cell_6t
Xbit_r103_c52 bl[52] br[52] wl[103] vdd gnd cell_6t
Xbit_r104_c52 bl[52] br[52] wl[104] vdd gnd cell_6t
Xbit_r105_c52 bl[52] br[52] wl[105] vdd gnd cell_6t
Xbit_r106_c52 bl[52] br[52] wl[106] vdd gnd cell_6t
Xbit_r107_c52 bl[52] br[52] wl[107] vdd gnd cell_6t
Xbit_r108_c52 bl[52] br[52] wl[108] vdd gnd cell_6t
Xbit_r109_c52 bl[52] br[52] wl[109] vdd gnd cell_6t
Xbit_r110_c52 bl[52] br[52] wl[110] vdd gnd cell_6t
Xbit_r111_c52 bl[52] br[52] wl[111] vdd gnd cell_6t
Xbit_r112_c52 bl[52] br[52] wl[112] vdd gnd cell_6t
Xbit_r113_c52 bl[52] br[52] wl[113] vdd gnd cell_6t
Xbit_r114_c52 bl[52] br[52] wl[114] vdd gnd cell_6t
Xbit_r115_c52 bl[52] br[52] wl[115] vdd gnd cell_6t
Xbit_r116_c52 bl[52] br[52] wl[116] vdd gnd cell_6t
Xbit_r117_c52 bl[52] br[52] wl[117] vdd gnd cell_6t
Xbit_r118_c52 bl[52] br[52] wl[118] vdd gnd cell_6t
Xbit_r119_c52 bl[52] br[52] wl[119] vdd gnd cell_6t
Xbit_r120_c52 bl[52] br[52] wl[120] vdd gnd cell_6t
Xbit_r121_c52 bl[52] br[52] wl[121] vdd gnd cell_6t
Xbit_r122_c52 bl[52] br[52] wl[122] vdd gnd cell_6t
Xbit_r123_c52 bl[52] br[52] wl[123] vdd gnd cell_6t
Xbit_r124_c52 bl[52] br[52] wl[124] vdd gnd cell_6t
Xbit_r125_c52 bl[52] br[52] wl[125] vdd gnd cell_6t
Xbit_r126_c52 bl[52] br[52] wl[126] vdd gnd cell_6t
Xbit_r127_c52 bl[52] br[52] wl[127] vdd gnd cell_6t
Xbit_r128_c52 bl[52] br[52] wl[128] vdd gnd cell_6t
Xbit_r129_c52 bl[52] br[52] wl[129] vdd gnd cell_6t
Xbit_r130_c52 bl[52] br[52] wl[130] vdd gnd cell_6t
Xbit_r131_c52 bl[52] br[52] wl[131] vdd gnd cell_6t
Xbit_r132_c52 bl[52] br[52] wl[132] vdd gnd cell_6t
Xbit_r133_c52 bl[52] br[52] wl[133] vdd gnd cell_6t
Xbit_r134_c52 bl[52] br[52] wl[134] vdd gnd cell_6t
Xbit_r135_c52 bl[52] br[52] wl[135] vdd gnd cell_6t
Xbit_r136_c52 bl[52] br[52] wl[136] vdd gnd cell_6t
Xbit_r137_c52 bl[52] br[52] wl[137] vdd gnd cell_6t
Xbit_r138_c52 bl[52] br[52] wl[138] vdd gnd cell_6t
Xbit_r139_c52 bl[52] br[52] wl[139] vdd gnd cell_6t
Xbit_r140_c52 bl[52] br[52] wl[140] vdd gnd cell_6t
Xbit_r141_c52 bl[52] br[52] wl[141] vdd gnd cell_6t
Xbit_r142_c52 bl[52] br[52] wl[142] vdd gnd cell_6t
Xbit_r143_c52 bl[52] br[52] wl[143] vdd gnd cell_6t
Xbit_r144_c52 bl[52] br[52] wl[144] vdd gnd cell_6t
Xbit_r145_c52 bl[52] br[52] wl[145] vdd gnd cell_6t
Xbit_r146_c52 bl[52] br[52] wl[146] vdd gnd cell_6t
Xbit_r147_c52 bl[52] br[52] wl[147] vdd gnd cell_6t
Xbit_r148_c52 bl[52] br[52] wl[148] vdd gnd cell_6t
Xbit_r149_c52 bl[52] br[52] wl[149] vdd gnd cell_6t
Xbit_r150_c52 bl[52] br[52] wl[150] vdd gnd cell_6t
Xbit_r151_c52 bl[52] br[52] wl[151] vdd gnd cell_6t
Xbit_r152_c52 bl[52] br[52] wl[152] vdd gnd cell_6t
Xbit_r153_c52 bl[52] br[52] wl[153] vdd gnd cell_6t
Xbit_r154_c52 bl[52] br[52] wl[154] vdd gnd cell_6t
Xbit_r155_c52 bl[52] br[52] wl[155] vdd gnd cell_6t
Xbit_r156_c52 bl[52] br[52] wl[156] vdd gnd cell_6t
Xbit_r157_c52 bl[52] br[52] wl[157] vdd gnd cell_6t
Xbit_r158_c52 bl[52] br[52] wl[158] vdd gnd cell_6t
Xbit_r159_c52 bl[52] br[52] wl[159] vdd gnd cell_6t
Xbit_r160_c52 bl[52] br[52] wl[160] vdd gnd cell_6t
Xbit_r161_c52 bl[52] br[52] wl[161] vdd gnd cell_6t
Xbit_r162_c52 bl[52] br[52] wl[162] vdd gnd cell_6t
Xbit_r163_c52 bl[52] br[52] wl[163] vdd gnd cell_6t
Xbit_r164_c52 bl[52] br[52] wl[164] vdd gnd cell_6t
Xbit_r165_c52 bl[52] br[52] wl[165] vdd gnd cell_6t
Xbit_r166_c52 bl[52] br[52] wl[166] vdd gnd cell_6t
Xbit_r167_c52 bl[52] br[52] wl[167] vdd gnd cell_6t
Xbit_r168_c52 bl[52] br[52] wl[168] vdd gnd cell_6t
Xbit_r169_c52 bl[52] br[52] wl[169] vdd gnd cell_6t
Xbit_r170_c52 bl[52] br[52] wl[170] vdd gnd cell_6t
Xbit_r171_c52 bl[52] br[52] wl[171] vdd gnd cell_6t
Xbit_r172_c52 bl[52] br[52] wl[172] vdd gnd cell_6t
Xbit_r173_c52 bl[52] br[52] wl[173] vdd gnd cell_6t
Xbit_r174_c52 bl[52] br[52] wl[174] vdd gnd cell_6t
Xbit_r175_c52 bl[52] br[52] wl[175] vdd gnd cell_6t
Xbit_r176_c52 bl[52] br[52] wl[176] vdd gnd cell_6t
Xbit_r177_c52 bl[52] br[52] wl[177] vdd gnd cell_6t
Xbit_r178_c52 bl[52] br[52] wl[178] vdd gnd cell_6t
Xbit_r179_c52 bl[52] br[52] wl[179] vdd gnd cell_6t
Xbit_r180_c52 bl[52] br[52] wl[180] vdd gnd cell_6t
Xbit_r181_c52 bl[52] br[52] wl[181] vdd gnd cell_6t
Xbit_r182_c52 bl[52] br[52] wl[182] vdd gnd cell_6t
Xbit_r183_c52 bl[52] br[52] wl[183] vdd gnd cell_6t
Xbit_r184_c52 bl[52] br[52] wl[184] vdd gnd cell_6t
Xbit_r185_c52 bl[52] br[52] wl[185] vdd gnd cell_6t
Xbit_r186_c52 bl[52] br[52] wl[186] vdd gnd cell_6t
Xbit_r187_c52 bl[52] br[52] wl[187] vdd gnd cell_6t
Xbit_r188_c52 bl[52] br[52] wl[188] vdd gnd cell_6t
Xbit_r189_c52 bl[52] br[52] wl[189] vdd gnd cell_6t
Xbit_r190_c52 bl[52] br[52] wl[190] vdd gnd cell_6t
Xbit_r191_c52 bl[52] br[52] wl[191] vdd gnd cell_6t
Xbit_r192_c52 bl[52] br[52] wl[192] vdd gnd cell_6t
Xbit_r193_c52 bl[52] br[52] wl[193] vdd gnd cell_6t
Xbit_r194_c52 bl[52] br[52] wl[194] vdd gnd cell_6t
Xbit_r195_c52 bl[52] br[52] wl[195] vdd gnd cell_6t
Xbit_r196_c52 bl[52] br[52] wl[196] vdd gnd cell_6t
Xbit_r197_c52 bl[52] br[52] wl[197] vdd gnd cell_6t
Xbit_r198_c52 bl[52] br[52] wl[198] vdd gnd cell_6t
Xbit_r199_c52 bl[52] br[52] wl[199] vdd gnd cell_6t
Xbit_r200_c52 bl[52] br[52] wl[200] vdd gnd cell_6t
Xbit_r201_c52 bl[52] br[52] wl[201] vdd gnd cell_6t
Xbit_r202_c52 bl[52] br[52] wl[202] vdd gnd cell_6t
Xbit_r203_c52 bl[52] br[52] wl[203] vdd gnd cell_6t
Xbit_r204_c52 bl[52] br[52] wl[204] vdd gnd cell_6t
Xbit_r205_c52 bl[52] br[52] wl[205] vdd gnd cell_6t
Xbit_r206_c52 bl[52] br[52] wl[206] vdd gnd cell_6t
Xbit_r207_c52 bl[52] br[52] wl[207] vdd gnd cell_6t
Xbit_r208_c52 bl[52] br[52] wl[208] vdd gnd cell_6t
Xbit_r209_c52 bl[52] br[52] wl[209] vdd gnd cell_6t
Xbit_r210_c52 bl[52] br[52] wl[210] vdd gnd cell_6t
Xbit_r211_c52 bl[52] br[52] wl[211] vdd gnd cell_6t
Xbit_r212_c52 bl[52] br[52] wl[212] vdd gnd cell_6t
Xbit_r213_c52 bl[52] br[52] wl[213] vdd gnd cell_6t
Xbit_r214_c52 bl[52] br[52] wl[214] vdd gnd cell_6t
Xbit_r215_c52 bl[52] br[52] wl[215] vdd gnd cell_6t
Xbit_r216_c52 bl[52] br[52] wl[216] vdd gnd cell_6t
Xbit_r217_c52 bl[52] br[52] wl[217] vdd gnd cell_6t
Xbit_r218_c52 bl[52] br[52] wl[218] vdd gnd cell_6t
Xbit_r219_c52 bl[52] br[52] wl[219] vdd gnd cell_6t
Xbit_r220_c52 bl[52] br[52] wl[220] vdd gnd cell_6t
Xbit_r221_c52 bl[52] br[52] wl[221] vdd gnd cell_6t
Xbit_r222_c52 bl[52] br[52] wl[222] vdd gnd cell_6t
Xbit_r223_c52 bl[52] br[52] wl[223] vdd gnd cell_6t
Xbit_r224_c52 bl[52] br[52] wl[224] vdd gnd cell_6t
Xbit_r225_c52 bl[52] br[52] wl[225] vdd gnd cell_6t
Xbit_r226_c52 bl[52] br[52] wl[226] vdd gnd cell_6t
Xbit_r227_c52 bl[52] br[52] wl[227] vdd gnd cell_6t
Xbit_r228_c52 bl[52] br[52] wl[228] vdd gnd cell_6t
Xbit_r229_c52 bl[52] br[52] wl[229] vdd gnd cell_6t
Xbit_r230_c52 bl[52] br[52] wl[230] vdd gnd cell_6t
Xbit_r231_c52 bl[52] br[52] wl[231] vdd gnd cell_6t
Xbit_r232_c52 bl[52] br[52] wl[232] vdd gnd cell_6t
Xbit_r233_c52 bl[52] br[52] wl[233] vdd gnd cell_6t
Xbit_r234_c52 bl[52] br[52] wl[234] vdd gnd cell_6t
Xbit_r235_c52 bl[52] br[52] wl[235] vdd gnd cell_6t
Xbit_r236_c52 bl[52] br[52] wl[236] vdd gnd cell_6t
Xbit_r237_c52 bl[52] br[52] wl[237] vdd gnd cell_6t
Xbit_r238_c52 bl[52] br[52] wl[238] vdd gnd cell_6t
Xbit_r239_c52 bl[52] br[52] wl[239] vdd gnd cell_6t
Xbit_r240_c52 bl[52] br[52] wl[240] vdd gnd cell_6t
Xbit_r241_c52 bl[52] br[52] wl[241] vdd gnd cell_6t
Xbit_r242_c52 bl[52] br[52] wl[242] vdd gnd cell_6t
Xbit_r243_c52 bl[52] br[52] wl[243] vdd gnd cell_6t
Xbit_r244_c52 bl[52] br[52] wl[244] vdd gnd cell_6t
Xbit_r245_c52 bl[52] br[52] wl[245] vdd gnd cell_6t
Xbit_r246_c52 bl[52] br[52] wl[246] vdd gnd cell_6t
Xbit_r247_c52 bl[52] br[52] wl[247] vdd gnd cell_6t
Xbit_r248_c52 bl[52] br[52] wl[248] vdd gnd cell_6t
Xbit_r249_c52 bl[52] br[52] wl[249] vdd gnd cell_6t
Xbit_r250_c52 bl[52] br[52] wl[250] vdd gnd cell_6t
Xbit_r251_c52 bl[52] br[52] wl[251] vdd gnd cell_6t
Xbit_r252_c52 bl[52] br[52] wl[252] vdd gnd cell_6t
Xbit_r253_c52 bl[52] br[52] wl[253] vdd gnd cell_6t
Xbit_r254_c52 bl[52] br[52] wl[254] vdd gnd cell_6t
Xbit_r255_c52 bl[52] br[52] wl[255] vdd gnd cell_6t
Xbit_r256_c52 bl[52] br[52] wl[256] vdd gnd cell_6t
Xbit_r257_c52 bl[52] br[52] wl[257] vdd gnd cell_6t
Xbit_r258_c52 bl[52] br[52] wl[258] vdd gnd cell_6t
Xbit_r259_c52 bl[52] br[52] wl[259] vdd gnd cell_6t
Xbit_r260_c52 bl[52] br[52] wl[260] vdd gnd cell_6t
Xbit_r261_c52 bl[52] br[52] wl[261] vdd gnd cell_6t
Xbit_r262_c52 bl[52] br[52] wl[262] vdd gnd cell_6t
Xbit_r263_c52 bl[52] br[52] wl[263] vdd gnd cell_6t
Xbit_r264_c52 bl[52] br[52] wl[264] vdd gnd cell_6t
Xbit_r265_c52 bl[52] br[52] wl[265] vdd gnd cell_6t
Xbit_r266_c52 bl[52] br[52] wl[266] vdd gnd cell_6t
Xbit_r267_c52 bl[52] br[52] wl[267] vdd gnd cell_6t
Xbit_r268_c52 bl[52] br[52] wl[268] vdd gnd cell_6t
Xbit_r269_c52 bl[52] br[52] wl[269] vdd gnd cell_6t
Xbit_r270_c52 bl[52] br[52] wl[270] vdd gnd cell_6t
Xbit_r271_c52 bl[52] br[52] wl[271] vdd gnd cell_6t
Xbit_r272_c52 bl[52] br[52] wl[272] vdd gnd cell_6t
Xbit_r273_c52 bl[52] br[52] wl[273] vdd gnd cell_6t
Xbit_r274_c52 bl[52] br[52] wl[274] vdd gnd cell_6t
Xbit_r275_c52 bl[52] br[52] wl[275] vdd gnd cell_6t
Xbit_r276_c52 bl[52] br[52] wl[276] vdd gnd cell_6t
Xbit_r277_c52 bl[52] br[52] wl[277] vdd gnd cell_6t
Xbit_r278_c52 bl[52] br[52] wl[278] vdd gnd cell_6t
Xbit_r279_c52 bl[52] br[52] wl[279] vdd gnd cell_6t
Xbit_r280_c52 bl[52] br[52] wl[280] vdd gnd cell_6t
Xbit_r281_c52 bl[52] br[52] wl[281] vdd gnd cell_6t
Xbit_r282_c52 bl[52] br[52] wl[282] vdd gnd cell_6t
Xbit_r283_c52 bl[52] br[52] wl[283] vdd gnd cell_6t
Xbit_r284_c52 bl[52] br[52] wl[284] vdd gnd cell_6t
Xbit_r285_c52 bl[52] br[52] wl[285] vdd gnd cell_6t
Xbit_r286_c52 bl[52] br[52] wl[286] vdd gnd cell_6t
Xbit_r287_c52 bl[52] br[52] wl[287] vdd gnd cell_6t
Xbit_r288_c52 bl[52] br[52] wl[288] vdd gnd cell_6t
Xbit_r289_c52 bl[52] br[52] wl[289] vdd gnd cell_6t
Xbit_r290_c52 bl[52] br[52] wl[290] vdd gnd cell_6t
Xbit_r291_c52 bl[52] br[52] wl[291] vdd gnd cell_6t
Xbit_r292_c52 bl[52] br[52] wl[292] vdd gnd cell_6t
Xbit_r293_c52 bl[52] br[52] wl[293] vdd gnd cell_6t
Xbit_r294_c52 bl[52] br[52] wl[294] vdd gnd cell_6t
Xbit_r295_c52 bl[52] br[52] wl[295] vdd gnd cell_6t
Xbit_r296_c52 bl[52] br[52] wl[296] vdd gnd cell_6t
Xbit_r297_c52 bl[52] br[52] wl[297] vdd gnd cell_6t
Xbit_r298_c52 bl[52] br[52] wl[298] vdd gnd cell_6t
Xbit_r299_c52 bl[52] br[52] wl[299] vdd gnd cell_6t
Xbit_r300_c52 bl[52] br[52] wl[300] vdd gnd cell_6t
Xbit_r301_c52 bl[52] br[52] wl[301] vdd gnd cell_6t
Xbit_r302_c52 bl[52] br[52] wl[302] vdd gnd cell_6t
Xbit_r303_c52 bl[52] br[52] wl[303] vdd gnd cell_6t
Xbit_r304_c52 bl[52] br[52] wl[304] vdd gnd cell_6t
Xbit_r305_c52 bl[52] br[52] wl[305] vdd gnd cell_6t
Xbit_r306_c52 bl[52] br[52] wl[306] vdd gnd cell_6t
Xbit_r307_c52 bl[52] br[52] wl[307] vdd gnd cell_6t
Xbit_r308_c52 bl[52] br[52] wl[308] vdd gnd cell_6t
Xbit_r309_c52 bl[52] br[52] wl[309] vdd gnd cell_6t
Xbit_r310_c52 bl[52] br[52] wl[310] vdd gnd cell_6t
Xbit_r311_c52 bl[52] br[52] wl[311] vdd gnd cell_6t
Xbit_r312_c52 bl[52] br[52] wl[312] vdd gnd cell_6t
Xbit_r313_c52 bl[52] br[52] wl[313] vdd gnd cell_6t
Xbit_r314_c52 bl[52] br[52] wl[314] vdd gnd cell_6t
Xbit_r315_c52 bl[52] br[52] wl[315] vdd gnd cell_6t
Xbit_r316_c52 bl[52] br[52] wl[316] vdd gnd cell_6t
Xbit_r317_c52 bl[52] br[52] wl[317] vdd gnd cell_6t
Xbit_r318_c52 bl[52] br[52] wl[318] vdd gnd cell_6t
Xbit_r319_c52 bl[52] br[52] wl[319] vdd gnd cell_6t
Xbit_r320_c52 bl[52] br[52] wl[320] vdd gnd cell_6t
Xbit_r321_c52 bl[52] br[52] wl[321] vdd gnd cell_6t
Xbit_r322_c52 bl[52] br[52] wl[322] vdd gnd cell_6t
Xbit_r323_c52 bl[52] br[52] wl[323] vdd gnd cell_6t
Xbit_r324_c52 bl[52] br[52] wl[324] vdd gnd cell_6t
Xbit_r325_c52 bl[52] br[52] wl[325] vdd gnd cell_6t
Xbit_r326_c52 bl[52] br[52] wl[326] vdd gnd cell_6t
Xbit_r327_c52 bl[52] br[52] wl[327] vdd gnd cell_6t
Xbit_r328_c52 bl[52] br[52] wl[328] vdd gnd cell_6t
Xbit_r329_c52 bl[52] br[52] wl[329] vdd gnd cell_6t
Xbit_r330_c52 bl[52] br[52] wl[330] vdd gnd cell_6t
Xbit_r331_c52 bl[52] br[52] wl[331] vdd gnd cell_6t
Xbit_r332_c52 bl[52] br[52] wl[332] vdd gnd cell_6t
Xbit_r333_c52 bl[52] br[52] wl[333] vdd gnd cell_6t
Xbit_r334_c52 bl[52] br[52] wl[334] vdd gnd cell_6t
Xbit_r335_c52 bl[52] br[52] wl[335] vdd gnd cell_6t
Xbit_r336_c52 bl[52] br[52] wl[336] vdd gnd cell_6t
Xbit_r337_c52 bl[52] br[52] wl[337] vdd gnd cell_6t
Xbit_r338_c52 bl[52] br[52] wl[338] vdd gnd cell_6t
Xbit_r339_c52 bl[52] br[52] wl[339] vdd gnd cell_6t
Xbit_r340_c52 bl[52] br[52] wl[340] vdd gnd cell_6t
Xbit_r341_c52 bl[52] br[52] wl[341] vdd gnd cell_6t
Xbit_r342_c52 bl[52] br[52] wl[342] vdd gnd cell_6t
Xbit_r343_c52 bl[52] br[52] wl[343] vdd gnd cell_6t
Xbit_r344_c52 bl[52] br[52] wl[344] vdd gnd cell_6t
Xbit_r345_c52 bl[52] br[52] wl[345] vdd gnd cell_6t
Xbit_r346_c52 bl[52] br[52] wl[346] vdd gnd cell_6t
Xbit_r347_c52 bl[52] br[52] wl[347] vdd gnd cell_6t
Xbit_r348_c52 bl[52] br[52] wl[348] vdd gnd cell_6t
Xbit_r349_c52 bl[52] br[52] wl[349] vdd gnd cell_6t
Xbit_r350_c52 bl[52] br[52] wl[350] vdd gnd cell_6t
Xbit_r351_c52 bl[52] br[52] wl[351] vdd gnd cell_6t
Xbit_r352_c52 bl[52] br[52] wl[352] vdd gnd cell_6t
Xbit_r353_c52 bl[52] br[52] wl[353] vdd gnd cell_6t
Xbit_r354_c52 bl[52] br[52] wl[354] vdd gnd cell_6t
Xbit_r355_c52 bl[52] br[52] wl[355] vdd gnd cell_6t
Xbit_r356_c52 bl[52] br[52] wl[356] vdd gnd cell_6t
Xbit_r357_c52 bl[52] br[52] wl[357] vdd gnd cell_6t
Xbit_r358_c52 bl[52] br[52] wl[358] vdd gnd cell_6t
Xbit_r359_c52 bl[52] br[52] wl[359] vdd gnd cell_6t
Xbit_r360_c52 bl[52] br[52] wl[360] vdd gnd cell_6t
Xbit_r361_c52 bl[52] br[52] wl[361] vdd gnd cell_6t
Xbit_r362_c52 bl[52] br[52] wl[362] vdd gnd cell_6t
Xbit_r363_c52 bl[52] br[52] wl[363] vdd gnd cell_6t
Xbit_r364_c52 bl[52] br[52] wl[364] vdd gnd cell_6t
Xbit_r365_c52 bl[52] br[52] wl[365] vdd gnd cell_6t
Xbit_r366_c52 bl[52] br[52] wl[366] vdd gnd cell_6t
Xbit_r367_c52 bl[52] br[52] wl[367] vdd gnd cell_6t
Xbit_r368_c52 bl[52] br[52] wl[368] vdd gnd cell_6t
Xbit_r369_c52 bl[52] br[52] wl[369] vdd gnd cell_6t
Xbit_r370_c52 bl[52] br[52] wl[370] vdd gnd cell_6t
Xbit_r371_c52 bl[52] br[52] wl[371] vdd gnd cell_6t
Xbit_r372_c52 bl[52] br[52] wl[372] vdd gnd cell_6t
Xbit_r373_c52 bl[52] br[52] wl[373] vdd gnd cell_6t
Xbit_r374_c52 bl[52] br[52] wl[374] vdd gnd cell_6t
Xbit_r375_c52 bl[52] br[52] wl[375] vdd gnd cell_6t
Xbit_r376_c52 bl[52] br[52] wl[376] vdd gnd cell_6t
Xbit_r377_c52 bl[52] br[52] wl[377] vdd gnd cell_6t
Xbit_r378_c52 bl[52] br[52] wl[378] vdd gnd cell_6t
Xbit_r379_c52 bl[52] br[52] wl[379] vdd gnd cell_6t
Xbit_r380_c52 bl[52] br[52] wl[380] vdd gnd cell_6t
Xbit_r381_c52 bl[52] br[52] wl[381] vdd gnd cell_6t
Xbit_r382_c52 bl[52] br[52] wl[382] vdd gnd cell_6t
Xbit_r383_c52 bl[52] br[52] wl[383] vdd gnd cell_6t
Xbit_r384_c52 bl[52] br[52] wl[384] vdd gnd cell_6t
Xbit_r385_c52 bl[52] br[52] wl[385] vdd gnd cell_6t
Xbit_r386_c52 bl[52] br[52] wl[386] vdd gnd cell_6t
Xbit_r387_c52 bl[52] br[52] wl[387] vdd gnd cell_6t
Xbit_r388_c52 bl[52] br[52] wl[388] vdd gnd cell_6t
Xbit_r389_c52 bl[52] br[52] wl[389] vdd gnd cell_6t
Xbit_r390_c52 bl[52] br[52] wl[390] vdd gnd cell_6t
Xbit_r391_c52 bl[52] br[52] wl[391] vdd gnd cell_6t
Xbit_r392_c52 bl[52] br[52] wl[392] vdd gnd cell_6t
Xbit_r393_c52 bl[52] br[52] wl[393] vdd gnd cell_6t
Xbit_r394_c52 bl[52] br[52] wl[394] vdd gnd cell_6t
Xbit_r395_c52 bl[52] br[52] wl[395] vdd gnd cell_6t
Xbit_r396_c52 bl[52] br[52] wl[396] vdd gnd cell_6t
Xbit_r397_c52 bl[52] br[52] wl[397] vdd gnd cell_6t
Xbit_r398_c52 bl[52] br[52] wl[398] vdd gnd cell_6t
Xbit_r399_c52 bl[52] br[52] wl[399] vdd gnd cell_6t
Xbit_r400_c52 bl[52] br[52] wl[400] vdd gnd cell_6t
Xbit_r401_c52 bl[52] br[52] wl[401] vdd gnd cell_6t
Xbit_r402_c52 bl[52] br[52] wl[402] vdd gnd cell_6t
Xbit_r403_c52 bl[52] br[52] wl[403] vdd gnd cell_6t
Xbit_r404_c52 bl[52] br[52] wl[404] vdd gnd cell_6t
Xbit_r405_c52 bl[52] br[52] wl[405] vdd gnd cell_6t
Xbit_r406_c52 bl[52] br[52] wl[406] vdd gnd cell_6t
Xbit_r407_c52 bl[52] br[52] wl[407] vdd gnd cell_6t
Xbit_r408_c52 bl[52] br[52] wl[408] vdd gnd cell_6t
Xbit_r409_c52 bl[52] br[52] wl[409] vdd gnd cell_6t
Xbit_r410_c52 bl[52] br[52] wl[410] vdd gnd cell_6t
Xbit_r411_c52 bl[52] br[52] wl[411] vdd gnd cell_6t
Xbit_r412_c52 bl[52] br[52] wl[412] vdd gnd cell_6t
Xbit_r413_c52 bl[52] br[52] wl[413] vdd gnd cell_6t
Xbit_r414_c52 bl[52] br[52] wl[414] vdd gnd cell_6t
Xbit_r415_c52 bl[52] br[52] wl[415] vdd gnd cell_6t
Xbit_r416_c52 bl[52] br[52] wl[416] vdd gnd cell_6t
Xbit_r417_c52 bl[52] br[52] wl[417] vdd gnd cell_6t
Xbit_r418_c52 bl[52] br[52] wl[418] vdd gnd cell_6t
Xbit_r419_c52 bl[52] br[52] wl[419] vdd gnd cell_6t
Xbit_r420_c52 bl[52] br[52] wl[420] vdd gnd cell_6t
Xbit_r421_c52 bl[52] br[52] wl[421] vdd gnd cell_6t
Xbit_r422_c52 bl[52] br[52] wl[422] vdd gnd cell_6t
Xbit_r423_c52 bl[52] br[52] wl[423] vdd gnd cell_6t
Xbit_r424_c52 bl[52] br[52] wl[424] vdd gnd cell_6t
Xbit_r425_c52 bl[52] br[52] wl[425] vdd gnd cell_6t
Xbit_r426_c52 bl[52] br[52] wl[426] vdd gnd cell_6t
Xbit_r427_c52 bl[52] br[52] wl[427] vdd gnd cell_6t
Xbit_r428_c52 bl[52] br[52] wl[428] vdd gnd cell_6t
Xbit_r429_c52 bl[52] br[52] wl[429] vdd gnd cell_6t
Xbit_r430_c52 bl[52] br[52] wl[430] vdd gnd cell_6t
Xbit_r431_c52 bl[52] br[52] wl[431] vdd gnd cell_6t
Xbit_r432_c52 bl[52] br[52] wl[432] vdd gnd cell_6t
Xbit_r433_c52 bl[52] br[52] wl[433] vdd gnd cell_6t
Xbit_r434_c52 bl[52] br[52] wl[434] vdd gnd cell_6t
Xbit_r435_c52 bl[52] br[52] wl[435] vdd gnd cell_6t
Xbit_r436_c52 bl[52] br[52] wl[436] vdd gnd cell_6t
Xbit_r437_c52 bl[52] br[52] wl[437] vdd gnd cell_6t
Xbit_r438_c52 bl[52] br[52] wl[438] vdd gnd cell_6t
Xbit_r439_c52 bl[52] br[52] wl[439] vdd gnd cell_6t
Xbit_r440_c52 bl[52] br[52] wl[440] vdd gnd cell_6t
Xbit_r441_c52 bl[52] br[52] wl[441] vdd gnd cell_6t
Xbit_r442_c52 bl[52] br[52] wl[442] vdd gnd cell_6t
Xbit_r443_c52 bl[52] br[52] wl[443] vdd gnd cell_6t
Xbit_r444_c52 bl[52] br[52] wl[444] vdd gnd cell_6t
Xbit_r445_c52 bl[52] br[52] wl[445] vdd gnd cell_6t
Xbit_r446_c52 bl[52] br[52] wl[446] vdd gnd cell_6t
Xbit_r447_c52 bl[52] br[52] wl[447] vdd gnd cell_6t
Xbit_r448_c52 bl[52] br[52] wl[448] vdd gnd cell_6t
Xbit_r449_c52 bl[52] br[52] wl[449] vdd gnd cell_6t
Xbit_r450_c52 bl[52] br[52] wl[450] vdd gnd cell_6t
Xbit_r451_c52 bl[52] br[52] wl[451] vdd gnd cell_6t
Xbit_r452_c52 bl[52] br[52] wl[452] vdd gnd cell_6t
Xbit_r453_c52 bl[52] br[52] wl[453] vdd gnd cell_6t
Xbit_r454_c52 bl[52] br[52] wl[454] vdd gnd cell_6t
Xbit_r455_c52 bl[52] br[52] wl[455] vdd gnd cell_6t
Xbit_r456_c52 bl[52] br[52] wl[456] vdd gnd cell_6t
Xbit_r457_c52 bl[52] br[52] wl[457] vdd gnd cell_6t
Xbit_r458_c52 bl[52] br[52] wl[458] vdd gnd cell_6t
Xbit_r459_c52 bl[52] br[52] wl[459] vdd gnd cell_6t
Xbit_r460_c52 bl[52] br[52] wl[460] vdd gnd cell_6t
Xbit_r461_c52 bl[52] br[52] wl[461] vdd gnd cell_6t
Xbit_r462_c52 bl[52] br[52] wl[462] vdd gnd cell_6t
Xbit_r463_c52 bl[52] br[52] wl[463] vdd gnd cell_6t
Xbit_r464_c52 bl[52] br[52] wl[464] vdd gnd cell_6t
Xbit_r465_c52 bl[52] br[52] wl[465] vdd gnd cell_6t
Xbit_r466_c52 bl[52] br[52] wl[466] vdd gnd cell_6t
Xbit_r467_c52 bl[52] br[52] wl[467] vdd gnd cell_6t
Xbit_r468_c52 bl[52] br[52] wl[468] vdd gnd cell_6t
Xbit_r469_c52 bl[52] br[52] wl[469] vdd gnd cell_6t
Xbit_r470_c52 bl[52] br[52] wl[470] vdd gnd cell_6t
Xbit_r471_c52 bl[52] br[52] wl[471] vdd gnd cell_6t
Xbit_r472_c52 bl[52] br[52] wl[472] vdd gnd cell_6t
Xbit_r473_c52 bl[52] br[52] wl[473] vdd gnd cell_6t
Xbit_r474_c52 bl[52] br[52] wl[474] vdd gnd cell_6t
Xbit_r475_c52 bl[52] br[52] wl[475] vdd gnd cell_6t
Xbit_r476_c52 bl[52] br[52] wl[476] vdd gnd cell_6t
Xbit_r477_c52 bl[52] br[52] wl[477] vdd gnd cell_6t
Xbit_r478_c52 bl[52] br[52] wl[478] vdd gnd cell_6t
Xbit_r479_c52 bl[52] br[52] wl[479] vdd gnd cell_6t
Xbit_r480_c52 bl[52] br[52] wl[480] vdd gnd cell_6t
Xbit_r481_c52 bl[52] br[52] wl[481] vdd gnd cell_6t
Xbit_r482_c52 bl[52] br[52] wl[482] vdd gnd cell_6t
Xbit_r483_c52 bl[52] br[52] wl[483] vdd gnd cell_6t
Xbit_r484_c52 bl[52] br[52] wl[484] vdd gnd cell_6t
Xbit_r485_c52 bl[52] br[52] wl[485] vdd gnd cell_6t
Xbit_r486_c52 bl[52] br[52] wl[486] vdd gnd cell_6t
Xbit_r487_c52 bl[52] br[52] wl[487] vdd gnd cell_6t
Xbit_r488_c52 bl[52] br[52] wl[488] vdd gnd cell_6t
Xbit_r489_c52 bl[52] br[52] wl[489] vdd gnd cell_6t
Xbit_r490_c52 bl[52] br[52] wl[490] vdd gnd cell_6t
Xbit_r491_c52 bl[52] br[52] wl[491] vdd gnd cell_6t
Xbit_r492_c52 bl[52] br[52] wl[492] vdd gnd cell_6t
Xbit_r493_c52 bl[52] br[52] wl[493] vdd gnd cell_6t
Xbit_r494_c52 bl[52] br[52] wl[494] vdd gnd cell_6t
Xbit_r495_c52 bl[52] br[52] wl[495] vdd gnd cell_6t
Xbit_r496_c52 bl[52] br[52] wl[496] vdd gnd cell_6t
Xbit_r497_c52 bl[52] br[52] wl[497] vdd gnd cell_6t
Xbit_r498_c52 bl[52] br[52] wl[498] vdd gnd cell_6t
Xbit_r499_c52 bl[52] br[52] wl[499] vdd gnd cell_6t
Xbit_r500_c52 bl[52] br[52] wl[500] vdd gnd cell_6t
Xbit_r501_c52 bl[52] br[52] wl[501] vdd gnd cell_6t
Xbit_r502_c52 bl[52] br[52] wl[502] vdd gnd cell_6t
Xbit_r503_c52 bl[52] br[52] wl[503] vdd gnd cell_6t
Xbit_r504_c52 bl[52] br[52] wl[504] vdd gnd cell_6t
Xbit_r505_c52 bl[52] br[52] wl[505] vdd gnd cell_6t
Xbit_r506_c52 bl[52] br[52] wl[506] vdd gnd cell_6t
Xbit_r507_c52 bl[52] br[52] wl[507] vdd gnd cell_6t
Xbit_r508_c52 bl[52] br[52] wl[508] vdd gnd cell_6t
Xbit_r509_c52 bl[52] br[52] wl[509] vdd gnd cell_6t
Xbit_r510_c52 bl[52] br[52] wl[510] vdd gnd cell_6t
Xbit_r511_c52 bl[52] br[52] wl[511] vdd gnd cell_6t
Xbit_r0_c53 bl[53] br[53] wl[0] vdd gnd cell_6t
Xbit_r1_c53 bl[53] br[53] wl[1] vdd gnd cell_6t
Xbit_r2_c53 bl[53] br[53] wl[2] vdd gnd cell_6t
Xbit_r3_c53 bl[53] br[53] wl[3] vdd gnd cell_6t
Xbit_r4_c53 bl[53] br[53] wl[4] vdd gnd cell_6t
Xbit_r5_c53 bl[53] br[53] wl[5] vdd gnd cell_6t
Xbit_r6_c53 bl[53] br[53] wl[6] vdd gnd cell_6t
Xbit_r7_c53 bl[53] br[53] wl[7] vdd gnd cell_6t
Xbit_r8_c53 bl[53] br[53] wl[8] vdd gnd cell_6t
Xbit_r9_c53 bl[53] br[53] wl[9] vdd gnd cell_6t
Xbit_r10_c53 bl[53] br[53] wl[10] vdd gnd cell_6t
Xbit_r11_c53 bl[53] br[53] wl[11] vdd gnd cell_6t
Xbit_r12_c53 bl[53] br[53] wl[12] vdd gnd cell_6t
Xbit_r13_c53 bl[53] br[53] wl[13] vdd gnd cell_6t
Xbit_r14_c53 bl[53] br[53] wl[14] vdd gnd cell_6t
Xbit_r15_c53 bl[53] br[53] wl[15] vdd gnd cell_6t
Xbit_r16_c53 bl[53] br[53] wl[16] vdd gnd cell_6t
Xbit_r17_c53 bl[53] br[53] wl[17] vdd gnd cell_6t
Xbit_r18_c53 bl[53] br[53] wl[18] vdd gnd cell_6t
Xbit_r19_c53 bl[53] br[53] wl[19] vdd gnd cell_6t
Xbit_r20_c53 bl[53] br[53] wl[20] vdd gnd cell_6t
Xbit_r21_c53 bl[53] br[53] wl[21] vdd gnd cell_6t
Xbit_r22_c53 bl[53] br[53] wl[22] vdd gnd cell_6t
Xbit_r23_c53 bl[53] br[53] wl[23] vdd gnd cell_6t
Xbit_r24_c53 bl[53] br[53] wl[24] vdd gnd cell_6t
Xbit_r25_c53 bl[53] br[53] wl[25] vdd gnd cell_6t
Xbit_r26_c53 bl[53] br[53] wl[26] vdd gnd cell_6t
Xbit_r27_c53 bl[53] br[53] wl[27] vdd gnd cell_6t
Xbit_r28_c53 bl[53] br[53] wl[28] vdd gnd cell_6t
Xbit_r29_c53 bl[53] br[53] wl[29] vdd gnd cell_6t
Xbit_r30_c53 bl[53] br[53] wl[30] vdd gnd cell_6t
Xbit_r31_c53 bl[53] br[53] wl[31] vdd gnd cell_6t
Xbit_r32_c53 bl[53] br[53] wl[32] vdd gnd cell_6t
Xbit_r33_c53 bl[53] br[53] wl[33] vdd gnd cell_6t
Xbit_r34_c53 bl[53] br[53] wl[34] vdd gnd cell_6t
Xbit_r35_c53 bl[53] br[53] wl[35] vdd gnd cell_6t
Xbit_r36_c53 bl[53] br[53] wl[36] vdd gnd cell_6t
Xbit_r37_c53 bl[53] br[53] wl[37] vdd gnd cell_6t
Xbit_r38_c53 bl[53] br[53] wl[38] vdd gnd cell_6t
Xbit_r39_c53 bl[53] br[53] wl[39] vdd gnd cell_6t
Xbit_r40_c53 bl[53] br[53] wl[40] vdd gnd cell_6t
Xbit_r41_c53 bl[53] br[53] wl[41] vdd gnd cell_6t
Xbit_r42_c53 bl[53] br[53] wl[42] vdd gnd cell_6t
Xbit_r43_c53 bl[53] br[53] wl[43] vdd gnd cell_6t
Xbit_r44_c53 bl[53] br[53] wl[44] vdd gnd cell_6t
Xbit_r45_c53 bl[53] br[53] wl[45] vdd gnd cell_6t
Xbit_r46_c53 bl[53] br[53] wl[46] vdd gnd cell_6t
Xbit_r47_c53 bl[53] br[53] wl[47] vdd gnd cell_6t
Xbit_r48_c53 bl[53] br[53] wl[48] vdd gnd cell_6t
Xbit_r49_c53 bl[53] br[53] wl[49] vdd gnd cell_6t
Xbit_r50_c53 bl[53] br[53] wl[50] vdd gnd cell_6t
Xbit_r51_c53 bl[53] br[53] wl[51] vdd gnd cell_6t
Xbit_r52_c53 bl[53] br[53] wl[52] vdd gnd cell_6t
Xbit_r53_c53 bl[53] br[53] wl[53] vdd gnd cell_6t
Xbit_r54_c53 bl[53] br[53] wl[54] vdd gnd cell_6t
Xbit_r55_c53 bl[53] br[53] wl[55] vdd gnd cell_6t
Xbit_r56_c53 bl[53] br[53] wl[56] vdd gnd cell_6t
Xbit_r57_c53 bl[53] br[53] wl[57] vdd gnd cell_6t
Xbit_r58_c53 bl[53] br[53] wl[58] vdd gnd cell_6t
Xbit_r59_c53 bl[53] br[53] wl[59] vdd gnd cell_6t
Xbit_r60_c53 bl[53] br[53] wl[60] vdd gnd cell_6t
Xbit_r61_c53 bl[53] br[53] wl[61] vdd gnd cell_6t
Xbit_r62_c53 bl[53] br[53] wl[62] vdd gnd cell_6t
Xbit_r63_c53 bl[53] br[53] wl[63] vdd gnd cell_6t
Xbit_r64_c53 bl[53] br[53] wl[64] vdd gnd cell_6t
Xbit_r65_c53 bl[53] br[53] wl[65] vdd gnd cell_6t
Xbit_r66_c53 bl[53] br[53] wl[66] vdd gnd cell_6t
Xbit_r67_c53 bl[53] br[53] wl[67] vdd gnd cell_6t
Xbit_r68_c53 bl[53] br[53] wl[68] vdd gnd cell_6t
Xbit_r69_c53 bl[53] br[53] wl[69] vdd gnd cell_6t
Xbit_r70_c53 bl[53] br[53] wl[70] vdd gnd cell_6t
Xbit_r71_c53 bl[53] br[53] wl[71] vdd gnd cell_6t
Xbit_r72_c53 bl[53] br[53] wl[72] vdd gnd cell_6t
Xbit_r73_c53 bl[53] br[53] wl[73] vdd gnd cell_6t
Xbit_r74_c53 bl[53] br[53] wl[74] vdd gnd cell_6t
Xbit_r75_c53 bl[53] br[53] wl[75] vdd gnd cell_6t
Xbit_r76_c53 bl[53] br[53] wl[76] vdd gnd cell_6t
Xbit_r77_c53 bl[53] br[53] wl[77] vdd gnd cell_6t
Xbit_r78_c53 bl[53] br[53] wl[78] vdd gnd cell_6t
Xbit_r79_c53 bl[53] br[53] wl[79] vdd gnd cell_6t
Xbit_r80_c53 bl[53] br[53] wl[80] vdd gnd cell_6t
Xbit_r81_c53 bl[53] br[53] wl[81] vdd gnd cell_6t
Xbit_r82_c53 bl[53] br[53] wl[82] vdd gnd cell_6t
Xbit_r83_c53 bl[53] br[53] wl[83] vdd gnd cell_6t
Xbit_r84_c53 bl[53] br[53] wl[84] vdd gnd cell_6t
Xbit_r85_c53 bl[53] br[53] wl[85] vdd gnd cell_6t
Xbit_r86_c53 bl[53] br[53] wl[86] vdd gnd cell_6t
Xbit_r87_c53 bl[53] br[53] wl[87] vdd gnd cell_6t
Xbit_r88_c53 bl[53] br[53] wl[88] vdd gnd cell_6t
Xbit_r89_c53 bl[53] br[53] wl[89] vdd gnd cell_6t
Xbit_r90_c53 bl[53] br[53] wl[90] vdd gnd cell_6t
Xbit_r91_c53 bl[53] br[53] wl[91] vdd gnd cell_6t
Xbit_r92_c53 bl[53] br[53] wl[92] vdd gnd cell_6t
Xbit_r93_c53 bl[53] br[53] wl[93] vdd gnd cell_6t
Xbit_r94_c53 bl[53] br[53] wl[94] vdd gnd cell_6t
Xbit_r95_c53 bl[53] br[53] wl[95] vdd gnd cell_6t
Xbit_r96_c53 bl[53] br[53] wl[96] vdd gnd cell_6t
Xbit_r97_c53 bl[53] br[53] wl[97] vdd gnd cell_6t
Xbit_r98_c53 bl[53] br[53] wl[98] vdd gnd cell_6t
Xbit_r99_c53 bl[53] br[53] wl[99] vdd gnd cell_6t
Xbit_r100_c53 bl[53] br[53] wl[100] vdd gnd cell_6t
Xbit_r101_c53 bl[53] br[53] wl[101] vdd gnd cell_6t
Xbit_r102_c53 bl[53] br[53] wl[102] vdd gnd cell_6t
Xbit_r103_c53 bl[53] br[53] wl[103] vdd gnd cell_6t
Xbit_r104_c53 bl[53] br[53] wl[104] vdd gnd cell_6t
Xbit_r105_c53 bl[53] br[53] wl[105] vdd gnd cell_6t
Xbit_r106_c53 bl[53] br[53] wl[106] vdd gnd cell_6t
Xbit_r107_c53 bl[53] br[53] wl[107] vdd gnd cell_6t
Xbit_r108_c53 bl[53] br[53] wl[108] vdd gnd cell_6t
Xbit_r109_c53 bl[53] br[53] wl[109] vdd gnd cell_6t
Xbit_r110_c53 bl[53] br[53] wl[110] vdd gnd cell_6t
Xbit_r111_c53 bl[53] br[53] wl[111] vdd gnd cell_6t
Xbit_r112_c53 bl[53] br[53] wl[112] vdd gnd cell_6t
Xbit_r113_c53 bl[53] br[53] wl[113] vdd gnd cell_6t
Xbit_r114_c53 bl[53] br[53] wl[114] vdd gnd cell_6t
Xbit_r115_c53 bl[53] br[53] wl[115] vdd gnd cell_6t
Xbit_r116_c53 bl[53] br[53] wl[116] vdd gnd cell_6t
Xbit_r117_c53 bl[53] br[53] wl[117] vdd gnd cell_6t
Xbit_r118_c53 bl[53] br[53] wl[118] vdd gnd cell_6t
Xbit_r119_c53 bl[53] br[53] wl[119] vdd gnd cell_6t
Xbit_r120_c53 bl[53] br[53] wl[120] vdd gnd cell_6t
Xbit_r121_c53 bl[53] br[53] wl[121] vdd gnd cell_6t
Xbit_r122_c53 bl[53] br[53] wl[122] vdd gnd cell_6t
Xbit_r123_c53 bl[53] br[53] wl[123] vdd gnd cell_6t
Xbit_r124_c53 bl[53] br[53] wl[124] vdd gnd cell_6t
Xbit_r125_c53 bl[53] br[53] wl[125] vdd gnd cell_6t
Xbit_r126_c53 bl[53] br[53] wl[126] vdd gnd cell_6t
Xbit_r127_c53 bl[53] br[53] wl[127] vdd gnd cell_6t
Xbit_r128_c53 bl[53] br[53] wl[128] vdd gnd cell_6t
Xbit_r129_c53 bl[53] br[53] wl[129] vdd gnd cell_6t
Xbit_r130_c53 bl[53] br[53] wl[130] vdd gnd cell_6t
Xbit_r131_c53 bl[53] br[53] wl[131] vdd gnd cell_6t
Xbit_r132_c53 bl[53] br[53] wl[132] vdd gnd cell_6t
Xbit_r133_c53 bl[53] br[53] wl[133] vdd gnd cell_6t
Xbit_r134_c53 bl[53] br[53] wl[134] vdd gnd cell_6t
Xbit_r135_c53 bl[53] br[53] wl[135] vdd gnd cell_6t
Xbit_r136_c53 bl[53] br[53] wl[136] vdd gnd cell_6t
Xbit_r137_c53 bl[53] br[53] wl[137] vdd gnd cell_6t
Xbit_r138_c53 bl[53] br[53] wl[138] vdd gnd cell_6t
Xbit_r139_c53 bl[53] br[53] wl[139] vdd gnd cell_6t
Xbit_r140_c53 bl[53] br[53] wl[140] vdd gnd cell_6t
Xbit_r141_c53 bl[53] br[53] wl[141] vdd gnd cell_6t
Xbit_r142_c53 bl[53] br[53] wl[142] vdd gnd cell_6t
Xbit_r143_c53 bl[53] br[53] wl[143] vdd gnd cell_6t
Xbit_r144_c53 bl[53] br[53] wl[144] vdd gnd cell_6t
Xbit_r145_c53 bl[53] br[53] wl[145] vdd gnd cell_6t
Xbit_r146_c53 bl[53] br[53] wl[146] vdd gnd cell_6t
Xbit_r147_c53 bl[53] br[53] wl[147] vdd gnd cell_6t
Xbit_r148_c53 bl[53] br[53] wl[148] vdd gnd cell_6t
Xbit_r149_c53 bl[53] br[53] wl[149] vdd gnd cell_6t
Xbit_r150_c53 bl[53] br[53] wl[150] vdd gnd cell_6t
Xbit_r151_c53 bl[53] br[53] wl[151] vdd gnd cell_6t
Xbit_r152_c53 bl[53] br[53] wl[152] vdd gnd cell_6t
Xbit_r153_c53 bl[53] br[53] wl[153] vdd gnd cell_6t
Xbit_r154_c53 bl[53] br[53] wl[154] vdd gnd cell_6t
Xbit_r155_c53 bl[53] br[53] wl[155] vdd gnd cell_6t
Xbit_r156_c53 bl[53] br[53] wl[156] vdd gnd cell_6t
Xbit_r157_c53 bl[53] br[53] wl[157] vdd gnd cell_6t
Xbit_r158_c53 bl[53] br[53] wl[158] vdd gnd cell_6t
Xbit_r159_c53 bl[53] br[53] wl[159] vdd gnd cell_6t
Xbit_r160_c53 bl[53] br[53] wl[160] vdd gnd cell_6t
Xbit_r161_c53 bl[53] br[53] wl[161] vdd gnd cell_6t
Xbit_r162_c53 bl[53] br[53] wl[162] vdd gnd cell_6t
Xbit_r163_c53 bl[53] br[53] wl[163] vdd gnd cell_6t
Xbit_r164_c53 bl[53] br[53] wl[164] vdd gnd cell_6t
Xbit_r165_c53 bl[53] br[53] wl[165] vdd gnd cell_6t
Xbit_r166_c53 bl[53] br[53] wl[166] vdd gnd cell_6t
Xbit_r167_c53 bl[53] br[53] wl[167] vdd gnd cell_6t
Xbit_r168_c53 bl[53] br[53] wl[168] vdd gnd cell_6t
Xbit_r169_c53 bl[53] br[53] wl[169] vdd gnd cell_6t
Xbit_r170_c53 bl[53] br[53] wl[170] vdd gnd cell_6t
Xbit_r171_c53 bl[53] br[53] wl[171] vdd gnd cell_6t
Xbit_r172_c53 bl[53] br[53] wl[172] vdd gnd cell_6t
Xbit_r173_c53 bl[53] br[53] wl[173] vdd gnd cell_6t
Xbit_r174_c53 bl[53] br[53] wl[174] vdd gnd cell_6t
Xbit_r175_c53 bl[53] br[53] wl[175] vdd gnd cell_6t
Xbit_r176_c53 bl[53] br[53] wl[176] vdd gnd cell_6t
Xbit_r177_c53 bl[53] br[53] wl[177] vdd gnd cell_6t
Xbit_r178_c53 bl[53] br[53] wl[178] vdd gnd cell_6t
Xbit_r179_c53 bl[53] br[53] wl[179] vdd gnd cell_6t
Xbit_r180_c53 bl[53] br[53] wl[180] vdd gnd cell_6t
Xbit_r181_c53 bl[53] br[53] wl[181] vdd gnd cell_6t
Xbit_r182_c53 bl[53] br[53] wl[182] vdd gnd cell_6t
Xbit_r183_c53 bl[53] br[53] wl[183] vdd gnd cell_6t
Xbit_r184_c53 bl[53] br[53] wl[184] vdd gnd cell_6t
Xbit_r185_c53 bl[53] br[53] wl[185] vdd gnd cell_6t
Xbit_r186_c53 bl[53] br[53] wl[186] vdd gnd cell_6t
Xbit_r187_c53 bl[53] br[53] wl[187] vdd gnd cell_6t
Xbit_r188_c53 bl[53] br[53] wl[188] vdd gnd cell_6t
Xbit_r189_c53 bl[53] br[53] wl[189] vdd gnd cell_6t
Xbit_r190_c53 bl[53] br[53] wl[190] vdd gnd cell_6t
Xbit_r191_c53 bl[53] br[53] wl[191] vdd gnd cell_6t
Xbit_r192_c53 bl[53] br[53] wl[192] vdd gnd cell_6t
Xbit_r193_c53 bl[53] br[53] wl[193] vdd gnd cell_6t
Xbit_r194_c53 bl[53] br[53] wl[194] vdd gnd cell_6t
Xbit_r195_c53 bl[53] br[53] wl[195] vdd gnd cell_6t
Xbit_r196_c53 bl[53] br[53] wl[196] vdd gnd cell_6t
Xbit_r197_c53 bl[53] br[53] wl[197] vdd gnd cell_6t
Xbit_r198_c53 bl[53] br[53] wl[198] vdd gnd cell_6t
Xbit_r199_c53 bl[53] br[53] wl[199] vdd gnd cell_6t
Xbit_r200_c53 bl[53] br[53] wl[200] vdd gnd cell_6t
Xbit_r201_c53 bl[53] br[53] wl[201] vdd gnd cell_6t
Xbit_r202_c53 bl[53] br[53] wl[202] vdd gnd cell_6t
Xbit_r203_c53 bl[53] br[53] wl[203] vdd gnd cell_6t
Xbit_r204_c53 bl[53] br[53] wl[204] vdd gnd cell_6t
Xbit_r205_c53 bl[53] br[53] wl[205] vdd gnd cell_6t
Xbit_r206_c53 bl[53] br[53] wl[206] vdd gnd cell_6t
Xbit_r207_c53 bl[53] br[53] wl[207] vdd gnd cell_6t
Xbit_r208_c53 bl[53] br[53] wl[208] vdd gnd cell_6t
Xbit_r209_c53 bl[53] br[53] wl[209] vdd gnd cell_6t
Xbit_r210_c53 bl[53] br[53] wl[210] vdd gnd cell_6t
Xbit_r211_c53 bl[53] br[53] wl[211] vdd gnd cell_6t
Xbit_r212_c53 bl[53] br[53] wl[212] vdd gnd cell_6t
Xbit_r213_c53 bl[53] br[53] wl[213] vdd gnd cell_6t
Xbit_r214_c53 bl[53] br[53] wl[214] vdd gnd cell_6t
Xbit_r215_c53 bl[53] br[53] wl[215] vdd gnd cell_6t
Xbit_r216_c53 bl[53] br[53] wl[216] vdd gnd cell_6t
Xbit_r217_c53 bl[53] br[53] wl[217] vdd gnd cell_6t
Xbit_r218_c53 bl[53] br[53] wl[218] vdd gnd cell_6t
Xbit_r219_c53 bl[53] br[53] wl[219] vdd gnd cell_6t
Xbit_r220_c53 bl[53] br[53] wl[220] vdd gnd cell_6t
Xbit_r221_c53 bl[53] br[53] wl[221] vdd gnd cell_6t
Xbit_r222_c53 bl[53] br[53] wl[222] vdd gnd cell_6t
Xbit_r223_c53 bl[53] br[53] wl[223] vdd gnd cell_6t
Xbit_r224_c53 bl[53] br[53] wl[224] vdd gnd cell_6t
Xbit_r225_c53 bl[53] br[53] wl[225] vdd gnd cell_6t
Xbit_r226_c53 bl[53] br[53] wl[226] vdd gnd cell_6t
Xbit_r227_c53 bl[53] br[53] wl[227] vdd gnd cell_6t
Xbit_r228_c53 bl[53] br[53] wl[228] vdd gnd cell_6t
Xbit_r229_c53 bl[53] br[53] wl[229] vdd gnd cell_6t
Xbit_r230_c53 bl[53] br[53] wl[230] vdd gnd cell_6t
Xbit_r231_c53 bl[53] br[53] wl[231] vdd gnd cell_6t
Xbit_r232_c53 bl[53] br[53] wl[232] vdd gnd cell_6t
Xbit_r233_c53 bl[53] br[53] wl[233] vdd gnd cell_6t
Xbit_r234_c53 bl[53] br[53] wl[234] vdd gnd cell_6t
Xbit_r235_c53 bl[53] br[53] wl[235] vdd gnd cell_6t
Xbit_r236_c53 bl[53] br[53] wl[236] vdd gnd cell_6t
Xbit_r237_c53 bl[53] br[53] wl[237] vdd gnd cell_6t
Xbit_r238_c53 bl[53] br[53] wl[238] vdd gnd cell_6t
Xbit_r239_c53 bl[53] br[53] wl[239] vdd gnd cell_6t
Xbit_r240_c53 bl[53] br[53] wl[240] vdd gnd cell_6t
Xbit_r241_c53 bl[53] br[53] wl[241] vdd gnd cell_6t
Xbit_r242_c53 bl[53] br[53] wl[242] vdd gnd cell_6t
Xbit_r243_c53 bl[53] br[53] wl[243] vdd gnd cell_6t
Xbit_r244_c53 bl[53] br[53] wl[244] vdd gnd cell_6t
Xbit_r245_c53 bl[53] br[53] wl[245] vdd gnd cell_6t
Xbit_r246_c53 bl[53] br[53] wl[246] vdd gnd cell_6t
Xbit_r247_c53 bl[53] br[53] wl[247] vdd gnd cell_6t
Xbit_r248_c53 bl[53] br[53] wl[248] vdd gnd cell_6t
Xbit_r249_c53 bl[53] br[53] wl[249] vdd gnd cell_6t
Xbit_r250_c53 bl[53] br[53] wl[250] vdd gnd cell_6t
Xbit_r251_c53 bl[53] br[53] wl[251] vdd gnd cell_6t
Xbit_r252_c53 bl[53] br[53] wl[252] vdd gnd cell_6t
Xbit_r253_c53 bl[53] br[53] wl[253] vdd gnd cell_6t
Xbit_r254_c53 bl[53] br[53] wl[254] vdd gnd cell_6t
Xbit_r255_c53 bl[53] br[53] wl[255] vdd gnd cell_6t
Xbit_r256_c53 bl[53] br[53] wl[256] vdd gnd cell_6t
Xbit_r257_c53 bl[53] br[53] wl[257] vdd gnd cell_6t
Xbit_r258_c53 bl[53] br[53] wl[258] vdd gnd cell_6t
Xbit_r259_c53 bl[53] br[53] wl[259] vdd gnd cell_6t
Xbit_r260_c53 bl[53] br[53] wl[260] vdd gnd cell_6t
Xbit_r261_c53 bl[53] br[53] wl[261] vdd gnd cell_6t
Xbit_r262_c53 bl[53] br[53] wl[262] vdd gnd cell_6t
Xbit_r263_c53 bl[53] br[53] wl[263] vdd gnd cell_6t
Xbit_r264_c53 bl[53] br[53] wl[264] vdd gnd cell_6t
Xbit_r265_c53 bl[53] br[53] wl[265] vdd gnd cell_6t
Xbit_r266_c53 bl[53] br[53] wl[266] vdd gnd cell_6t
Xbit_r267_c53 bl[53] br[53] wl[267] vdd gnd cell_6t
Xbit_r268_c53 bl[53] br[53] wl[268] vdd gnd cell_6t
Xbit_r269_c53 bl[53] br[53] wl[269] vdd gnd cell_6t
Xbit_r270_c53 bl[53] br[53] wl[270] vdd gnd cell_6t
Xbit_r271_c53 bl[53] br[53] wl[271] vdd gnd cell_6t
Xbit_r272_c53 bl[53] br[53] wl[272] vdd gnd cell_6t
Xbit_r273_c53 bl[53] br[53] wl[273] vdd gnd cell_6t
Xbit_r274_c53 bl[53] br[53] wl[274] vdd gnd cell_6t
Xbit_r275_c53 bl[53] br[53] wl[275] vdd gnd cell_6t
Xbit_r276_c53 bl[53] br[53] wl[276] vdd gnd cell_6t
Xbit_r277_c53 bl[53] br[53] wl[277] vdd gnd cell_6t
Xbit_r278_c53 bl[53] br[53] wl[278] vdd gnd cell_6t
Xbit_r279_c53 bl[53] br[53] wl[279] vdd gnd cell_6t
Xbit_r280_c53 bl[53] br[53] wl[280] vdd gnd cell_6t
Xbit_r281_c53 bl[53] br[53] wl[281] vdd gnd cell_6t
Xbit_r282_c53 bl[53] br[53] wl[282] vdd gnd cell_6t
Xbit_r283_c53 bl[53] br[53] wl[283] vdd gnd cell_6t
Xbit_r284_c53 bl[53] br[53] wl[284] vdd gnd cell_6t
Xbit_r285_c53 bl[53] br[53] wl[285] vdd gnd cell_6t
Xbit_r286_c53 bl[53] br[53] wl[286] vdd gnd cell_6t
Xbit_r287_c53 bl[53] br[53] wl[287] vdd gnd cell_6t
Xbit_r288_c53 bl[53] br[53] wl[288] vdd gnd cell_6t
Xbit_r289_c53 bl[53] br[53] wl[289] vdd gnd cell_6t
Xbit_r290_c53 bl[53] br[53] wl[290] vdd gnd cell_6t
Xbit_r291_c53 bl[53] br[53] wl[291] vdd gnd cell_6t
Xbit_r292_c53 bl[53] br[53] wl[292] vdd gnd cell_6t
Xbit_r293_c53 bl[53] br[53] wl[293] vdd gnd cell_6t
Xbit_r294_c53 bl[53] br[53] wl[294] vdd gnd cell_6t
Xbit_r295_c53 bl[53] br[53] wl[295] vdd gnd cell_6t
Xbit_r296_c53 bl[53] br[53] wl[296] vdd gnd cell_6t
Xbit_r297_c53 bl[53] br[53] wl[297] vdd gnd cell_6t
Xbit_r298_c53 bl[53] br[53] wl[298] vdd gnd cell_6t
Xbit_r299_c53 bl[53] br[53] wl[299] vdd gnd cell_6t
Xbit_r300_c53 bl[53] br[53] wl[300] vdd gnd cell_6t
Xbit_r301_c53 bl[53] br[53] wl[301] vdd gnd cell_6t
Xbit_r302_c53 bl[53] br[53] wl[302] vdd gnd cell_6t
Xbit_r303_c53 bl[53] br[53] wl[303] vdd gnd cell_6t
Xbit_r304_c53 bl[53] br[53] wl[304] vdd gnd cell_6t
Xbit_r305_c53 bl[53] br[53] wl[305] vdd gnd cell_6t
Xbit_r306_c53 bl[53] br[53] wl[306] vdd gnd cell_6t
Xbit_r307_c53 bl[53] br[53] wl[307] vdd gnd cell_6t
Xbit_r308_c53 bl[53] br[53] wl[308] vdd gnd cell_6t
Xbit_r309_c53 bl[53] br[53] wl[309] vdd gnd cell_6t
Xbit_r310_c53 bl[53] br[53] wl[310] vdd gnd cell_6t
Xbit_r311_c53 bl[53] br[53] wl[311] vdd gnd cell_6t
Xbit_r312_c53 bl[53] br[53] wl[312] vdd gnd cell_6t
Xbit_r313_c53 bl[53] br[53] wl[313] vdd gnd cell_6t
Xbit_r314_c53 bl[53] br[53] wl[314] vdd gnd cell_6t
Xbit_r315_c53 bl[53] br[53] wl[315] vdd gnd cell_6t
Xbit_r316_c53 bl[53] br[53] wl[316] vdd gnd cell_6t
Xbit_r317_c53 bl[53] br[53] wl[317] vdd gnd cell_6t
Xbit_r318_c53 bl[53] br[53] wl[318] vdd gnd cell_6t
Xbit_r319_c53 bl[53] br[53] wl[319] vdd gnd cell_6t
Xbit_r320_c53 bl[53] br[53] wl[320] vdd gnd cell_6t
Xbit_r321_c53 bl[53] br[53] wl[321] vdd gnd cell_6t
Xbit_r322_c53 bl[53] br[53] wl[322] vdd gnd cell_6t
Xbit_r323_c53 bl[53] br[53] wl[323] vdd gnd cell_6t
Xbit_r324_c53 bl[53] br[53] wl[324] vdd gnd cell_6t
Xbit_r325_c53 bl[53] br[53] wl[325] vdd gnd cell_6t
Xbit_r326_c53 bl[53] br[53] wl[326] vdd gnd cell_6t
Xbit_r327_c53 bl[53] br[53] wl[327] vdd gnd cell_6t
Xbit_r328_c53 bl[53] br[53] wl[328] vdd gnd cell_6t
Xbit_r329_c53 bl[53] br[53] wl[329] vdd gnd cell_6t
Xbit_r330_c53 bl[53] br[53] wl[330] vdd gnd cell_6t
Xbit_r331_c53 bl[53] br[53] wl[331] vdd gnd cell_6t
Xbit_r332_c53 bl[53] br[53] wl[332] vdd gnd cell_6t
Xbit_r333_c53 bl[53] br[53] wl[333] vdd gnd cell_6t
Xbit_r334_c53 bl[53] br[53] wl[334] vdd gnd cell_6t
Xbit_r335_c53 bl[53] br[53] wl[335] vdd gnd cell_6t
Xbit_r336_c53 bl[53] br[53] wl[336] vdd gnd cell_6t
Xbit_r337_c53 bl[53] br[53] wl[337] vdd gnd cell_6t
Xbit_r338_c53 bl[53] br[53] wl[338] vdd gnd cell_6t
Xbit_r339_c53 bl[53] br[53] wl[339] vdd gnd cell_6t
Xbit_r340_c53 bl[53] br[53] wl[340] vdd gnd cell_6t
Xbit_r341_c53 bl[53] br[53] wl[341] vdd gnd cell_6t
Xbit_r342_c53 bl[53] br[53] wl[342] vdd gnd cell_6t
Xbit_r343_c53 bl[53] br[53] wl[343] vdd gnd cell_6t
Xbit_r344_c53 bl[53] br[53] wl[344] vdd gnd cell_6t
Xbit_r345_c53 bl[53] br[53] wl[345] vdd gnd cell_6t
Xbit_r346_c53 bl[53] br[53] wl[346] vdd gnd cell_6t
Xbit_r347_c53 bl[53] br[53] wl[347] vdd gnd cell_6t
Xbit_r348_c53 bl[53] br[53] wl[348] vdd gnd cell_6t
Xbit_r349_c53 bl[53] br[53] wl[349] vdd gnd cell_6t
Xbit_r350_c53 bl[53] br[53] wl[350] vdd gnd cell_6t
Xbit_r351_c53 bl[53] br[53] wl[351] vdd gnd cell_6t
Xbit_r352_c53 bl[53] br[53] wl[352] vdd gnd cell_6t
Xbit_r353_c53 bl[53] br[53] wl[353] vdd gnd cell_6t
Xbit_r354_c53 bl[53] br[53] wl[354] vdd gnd cell_6t
Xbit_r355_c53 bl[53] br[53] wl[355] vdd gnd cell_6t
Xbit_r356_c53 bl[53] br[53] wl[356] vdd gnd cell_6t
Xbit_r357_c53 bl[53] br[53] wl[357] vdd gnd cell_6t
Xbit_r358_c53 bl[53] br[53] wl[358] vdd gnd cell_6t
Xbit_r359_c53 bl[53] br[53] wl[359] vdd gnd cell_6t
Xbit_r360_c53 bl[53] br[53] wl[360] vdd gnd cell_6t
Xbit_r361_c53 bl[53] br[53] wl[361] vdd gnd cell_6t
Xbit_r362_c53 bl[53] br[53] wl[362] vdd gnd cell_6t
Xbit_r363_c53 bl[53] br[53] wl[363] vdd gnd cell_6t
Xbit_r364_c53 bl[53] br[53] wl[364] vdd gnd cell_6t
Xbit_r365_c53 bl[53] br[53] wl[365] vdd gnd cell_6t
Xbit_r366_c53 bl[53] br[53] wl[366] vdd gnd cell_6t
Xbit_r367_c53 bl[53] br[53] wl[367] vdd gnd cell_6t
Xbit_r368_c53 bl[53] br[53] wl[368] vdd gnd cell_6t
Xbit_r369_c53 bl[53] br[53] wl[369] vdd gnd cell_6t
Xbit_r370_c53 bl[53] br[53] wl[370] vdd gnd cell_6t
Xbit_r371_c53 bl[53] br[53] wl[371] vdd gnd cell_6t
Xbit_r372_c53 bl[53] br[53] wl[372] vdd gnd cell_6t
Xbit_r373_c53 bl[53] br[53] wl[373] vdd gnd cell_6t
Xbit_r374_c53 bl[53] br[53] wl[374] vdd gnd cell_6t
Xbit_r375_c53 bl[53] br[53] wl[375] vdd gnd cell_6t
Xbit_r376_c53 bl[53] br[53] wl[376] vdd gnd cell_6t
Xbit_r377_c53 bl[53] br[53] wl[377] vdd gnd cell_6t
Xbit_r378_c53 bl[53] br[53] wl[378] vdd gnd cell_6t
Xbit_r379_c53 bl[53] br[53] wl[379] vdd gnd cell_6t
Xbit_r380_c53 bl[53] br[53] wl[380] vdd gnd cell_6t
Xbit_r381_c53 bl[53] br[53] wl[381] vdd gnd cell_6t
Xbit_r382_c53 bl[53] br[53] wl[382] vdd gnd cell_6t
Xbit_r383_c53 bl[53] br[53] wl[383] vdd gnd cell_6t
Xbit_r384_c53 bl[53] br[53] wl[384] vdd gnd cell_6t
Xbit_r385_c53 bl[53] br[53] wl[385] vdd gnd cell_6t
Xbit_r386_c53 bl[53] br[53] wl[386] vdd gnd cell_6t
Xbit_r387_c53 bl[53] br[53] wl[387] vdd gnd cell_6t
Xbit_r388_c53 bl[53] br[53] wl[388] vdd gnd cell_6t
Xbit_r389_c53 bl[53] br[53] wl[389] vdd gnd cell_6t
Xbit_r390_c53 bl[53] br[53] wl[390] vdd gnd cell_6t
Xbit_r391_c53 bl[53] br[53] wl[391] vdd gnd cell_6t
Xbit_r392_c53 bl[53] br[53] wl[392] vdd gnd cell_6t
Xbit_r393_c53 bl[53] br[53] wl[393] vdd gnd cell_6t
Xbit_r394_c53 bl[53] br[53] wl[394] vdd gnd cell_6t
Xbit_r395_c53 bl[53] br[53] wl[395] vdd gnd cell_6t
Xbit_r396_c53 bl[53] br[53] wl[396] vdd gnd cell_6t
Xbit_r397_c53 bl[53] br[53] wl[397] vdd gnd cell_6t
Xbit_r398_c53 bl[53] br[53] wl[398] vdd gnd cell_6t
Xbit_r399_c53 bl[53] br[53] wl[399] vdd gnd cell_6t
Xbit_r400_c53 bl[53] br[53] wl[400] vdd gnd cell_6t
Xbit_r401_c53 bl[53] br[53] wl[401] vdd gnd cell_6t
Xbit_r402_c53 bl[53] br[53] wl[402] vdd gnd cell_6t
Xbit_r403_c53 bl[53] br[53] wl[403] vdd gnd cell_6t
Xbit_r404_c53 bl[53] br[53] wl[404] vdd gnd cell_6t
Xbit_r405_c53 bl[53] br[53] wl[405] vdd gnd cell_6t
Xbit_r406_c53 bl[53] br[53] wl[406] vdd gnd cell_6t
Xbit_r407_c53 bl[53] br[53] wl[407] vdd gnd cell_6t
Xbit_r408_c53 bl[53] br[53] wl[408] vdd gnd cell_6t
Xbit_r409_c53 bl[53] br[53] wl[409] vdd gnd cell_6t
Xbit_r410_c53 bl[53] br[53] wl[410] vdd gnd cell_6t
Xbit_r411_c53 bl[53] br[53] wl[411] vdd gnd cell_6t
Xbit_r412_c53 bl[53] br[53] wl[412] vdd gnd cell_6t
Xbit_r413_c53 bl[53] br[53] wl[413] vdd gnd cell_6t
Xbit_r414_c53 bl[53] br[53] wl[414] vdd gnd cell_6t
Xbit_r415_c53 bl[53] br[53] wl[415] vdd gnd cell_6t
Xbit_r416_c53 bl[53] br[53] wl[416] vdd gnd cell_6t
Xbit_r417_c53 bl[53] br[53] wl[417] vdd gnd cell_6t
Xbit_r418_c53 bl[53] br[53] wl[418] vdd gnd cell_6t
Xbit_r419_c53 bl[53] br[53] wl[419] vdd gnd cell_6t
Xbit_r420_c53 bl[53] br[53] wl[420] vdd gnd cell_6t
Xbit_r421_c53 bl[53] br[53] wl[421] vdd gnd cell_6t
Xbit_r422_c53 bl[53] br[53] wl[422] vdd gnd cell_6t
Xbit_r423_c53 bl[53] br[53] wl[423] vdd gnd cell_6t
Xbit_r424_c53 bl[53] br[53] wl[424] vdd gnd cell_6t
Xbit_r425_c53 bl[53] br[53] wl[425] vdd gnd cell_6t
Xbit_r426_c53 bl[53] br[53] wl[426] vdd gnd cell_6t
Xbit_r427_c53 bl[53] br[53] wl[427] vdd gnd cell_6t
Xbit_r428_c53 bl[53] br[53] wl[428] vdd gnd cell_6t
Xbit_r429_c53 bl[53] br[53] wl[429] vdd gnd cell_6t
Xbit_r430_c53 bl[53] br[53] wl[430] vdd gnd cell_6t
Xbit_r431_c53 bl[53] br[53] wl[431] vdd gnd cell_6t
Xbit_r432_c53 bl[53] br[53] wl[432] vdd gnd cell_6t
Xbit_r433_c53 bl[53] br[53] wl[433] vdd gnd cell_6t
Xbit_r434_c53 bl[53] br[53] wl[434] vdd gnd cell_6t
Xbit_r435_c53 bl[53] br[53] wl[435] vdd gnd cell_6t
Xbit_r436_c53 bl[53] br[53] wl[436] vdd gnd cell_6t
Xbit_r437_c53 bl[53] br[53] wl[437] vdd gnd cell_6t
Xbit_r438_c53 bl[53] br[53] wl[438] vdd gnd cell_6t
Xbit_r439_c53 bl[53] br[53] wl[439] vdd gnd cell_6t
Xbit_r440_c53 bl[53] br[53] wl[440] vdd gnd cell_6t
Xbit_r441_c53 bl[53] br[53] wl[441] vdd gnd cell_6t
Xbit_r442_c53 bl[53] br[53] wl[442] vdd gnd cell_6t
Xbit_r443_c53 bl[53] br[53] wl[443] vdd gnd cell_6t
Xbit_r444_c53 bl[53] br[53] wl[444] vdd gnd cell_6t
Xbit_r445_c53 bl[53] br[53] wl[445] vdd gnd cell_6t
Xbit_r446_c53 bl[53] br[53] wl[446] vdd gnd cell_6t
Xbit_r447_c53 bl[53] br[53] wl[447] vdd gnd cell_6t
Xbit_r448_c53 bl[53] br[53] wl[448] vdd gnd cell_6t
Xbit_r449_c53 bl[53] br[53] wl[449] vdd gnd cell_6t
Xbit_r450_c53 bl[53] br[53] wl[450] vdd gnd cell_6t
Xbit_r451_c53 bl[53] br[53] wl[451] vdd gnd cell_6t
Xbit_r452_c53 bl[53] br[53] wl[452] vdd gnd cell_6t
Xbit_r453_c53 bl[53] br[53] wl[453] vdd gnd cell_6t
Xbit_r454_c53 bl[53] br[53] wl[454] vdd gnd cell_6t
Xbit_r455_c53 bl[53] br[53] wl[455] vdd gnd cell_6t
Xbit_r456_c53 bl[53] br[53] wl[456] vdd gnd cell_6t
Xbit_r457_c53 bl[53] br[53] wl[457] vdd gnd cell_6t
Xbit_r458_c53 bl[53] br[53] wl[458] vdd gnd cell_6t
Xbit_r459_c53 bl[53] br[53] wl[459] vdd gnd cell_6t
Xbit_r460_c53 bl[53] br[53] wl[460] vdd gnd cell_6t
Xbit_r461_c53 bl[53] br[53] wl[461] vdd gnd cell_6t
Xbit_r462_c53 bl[53] br[53] wl[462] vdd gnd cell_6t
Xbit_r463_c53 bl[53] br[53] wl[463] vdd gnd cell_6t
Xbit_r464_c53 bl[53] br[53] wl[464] vdd gnd cell_6t
Xbit_r465_c53 bl[53] br[53] wl[465] vdd gnd cell_6t
Xbit_r466_c53 bl[53] br[53] wl[466] vdd gnd cell_6t
Xbit_r467_c53 bl[53] br[53] wl[467] vdd gnd cell_6t
Xbit_r468_c53 bl[53] br[53] wl[468] vdd gnd cell_6t
Xbit_r469_c53 bl[53] br[53] wl[469] vdd gnd cell_6t
Xbit_r470_c53 bl[53] br[53] wl[470] vdd gnd cell_6t
Xbit_r471_c53 bl[53] br[53] wl[471] vdd gnd cell_6t
Xbit_r472_c53 bl[53] br[53] wl[472] vdd gnd cell_6t
Xbit_r473_c53 bl[53] br[53] wl[473] vdd gnd cell_6t
Xbit_r474_c53 bl[53] br[53] wl[474] vdd gnd cell_6t
Xbit_r475_c53 bl[53] br[53] wl[475] vdd gnd cell_6t
Xbit_r476_c53 bl[53] br[53] wl[476] vdd gnd cell_6t
Xbit_r477_c53 bl[53] br[53] wl[477] vdd gnd cell_6t
Xbit_r478_c53 bl[53] br[53] wl[478] vdd gnd cell_6t
Xbit_r479_c53 bl[53] br[53] wl[479] vdd gnd cell_6t
Xbit_r480_c53 bl[53] br[53] wl[480] vdd gnd cell_6t
Xbit_r481_c53 bl[53] br[53] wl[481] vdd gnd cell_6t
Xbit_r482_c53 bl[53] br[53] wl[482] vdd gnd cell_6t
Xbit_r483_c53 bl[53] br[53] wl[483] vdd gnd cell_6t
Xbit_r484_c53 bl[53] br[53] wl[484] vdd gnd cell_6t
Xbit_r485_c53 bl[53] br[53] wl[485] vdd gnd cell_6t
Xbit_r486_c53 bl[53] br[53] wl[486] vdd gnd cell_6t
Xbit_r487_c53 bl[53] br[53] wl[487] vdd gnd cell_6t
Xbit_r488_c53 bl[53] br[53] wl[488] vdd gnd cell_6t
Xbit_r489_c53 bl[53] br[53] wl[489] vdd gnd cell_6t
Xbit_r490_c53 bl[53] br[53] wl[490] vdd gnd cell_6t
Xbit_r491_c53 bl[53] br[53] wl[491] vdd gnd cell_6t
Xbit_r492_c53 bl[53] br[53] wl[492] vdd gnd cell_6t
Xbit_r493_c53 bl[53] br[53] wl[493] vdd gnd cell_6t
Xbit_r494_c53 bl[53] br[53] wl[494] vdd gnd cell_6t
Xbit_r495_c53 bl[53] br[53] wl[495] vdd gnd cell_6t
Xbit_r496_c53 bl[53] br[53] wl[496] vdd gnd cell_6t
Xbit_r497_c53 bl[53] br[53] wl[497] vdd gnd cell_6t
Xbit_r498_c53 bl[53] br[53] wl[498] vdd gnd cell_6t
Xbit_r499_c53 bl[53] br[53] wl[499] vdd gnd cell_6t
Xbit_r500_c53 bl[53] br[53] wl[500] vdd gnd cell_6t
Xbit_r501_c53 bl[53] br[53] wl[501] vdd gnd cell_6t
Xbit_r502_c53 bl[53] br[53] wl[502] vdd gnd cell_6t
Xbit_r503_c53 bl[53] br[53] wl[503] vdd gnd cell_6t
Xbit_r504_c53 bl[53] br[53] wl[504] vdd gnd cell_6t
Xbit_r505_c53 bl[53] br[53] wl[505] vdd gnd cell_6t
Xbit_r506_c53 bl[53] br[53] wl[506] vdd gnd cell_6t
Xbit_r507_c53 bl[53] br[53] wl[507] vdd gnd cell_6t
Xbit_r508_c53 bl[53] br[53] wl[508] vdd gnd cell_6t
Xbit_r509_c53 bl[53] br[53] wl[509] vdd gnd cell_6t
Xbit_r510_c53 bl[53] br[53] wl[510] vdd gnd cell_6t
Xbit_r511_c53 bl[53] br[53] wl[511] vdd gnd cell_6t
Xbit_r0_c54 bl[54] br[54] wl[0] vdd gnd cell_6t
Xbit_r1_c54 bl[54] br[54] wl[1] vdd gnd cell_6t
Xbit_r2_c54 bl[54] br[54] wl[2] vdd gnd cell_6t
Xbit_r3_c54 bl[54] br[54] wl[3] vdd gnd cell_6t
Xbit_r4_c54 bl[54] br[54] wl[4] vdd gnd cell_6t
Xbit_r5_c54 bl[54] br[54] wl[5] vdd gnd cell_6t
Xbit_r6_c54 bl[54] br[54] wl[6] vdd gnd cell_6t
Xbit_r7_c54 bl[54] br[54] wl[7] vdd gnd cell_6t
Xbit_r8_c54 bl[54] br[54] wl[8] vdd gnd cell_6t
Xbit_r9_c54 bl[54] br[54] wl[9] vdd gnd cell_6t
Xbit_r10_c54 bl[54] br[54] wl[10] vdd gnd cell_6t
Xbit_r11_c54 bl[54] br[54] wl[11] vdd gnd cell_6t
Xbit_r12_c54 bl[54] br[54] wl[12] vdd gnd cell_6t
Xbit_r13_c54 bl[54] br[54] wl[13] vdd gnd cell_6t
Xbit_r14_c54 bl[54] br[54] wl[14] vdd gnd cell_6t
Xbit_r15_c54 bl[54] br[54] wl[15] vdd gnd cell_6t
Xbit_r16_c54 bl[54] br[54] wl[16] vdd gnd cell_6t
Xbit_r17_c54 bl[54] br[54] wl[17] vdd gnd cell_6t
Xbit_r18_c54 bl[54] br[54] wl[18] vdd gnd cell_6t
Xbit_r19_c54 bl[54] br[54] wl[19] vdd gnd cell_6t
Xbit_r20_c54 bl[54] br[54] wl[20] vdd gnd cell_6t
Xbit_r21_c54 bl[54] br[54] wl[21] vdd gnd cell_6t
Xbit_r22_c54 bl[54] br[54] wl[22] vdd gnd cell_6t
Xbit_r23_c54 bl[54] br[54] wl[23] vdd gnd cell_6t
Xbit_r24_c54 bl[54] br[54] wl[24] vdd gnd cell_6t
Xbit_r25_c54 bl[54] br[54] wl[25] vdd gnd cell_6t
Xbit_r26_c54 bl[54] br[54] wl[26] vdd gnd cell_6t
Xbit_r27_c54 bl[54] br[54] wl[27] vdd gnd cell_6t
Xbit_r28_c54 bl[54] br[54] wl[28] vdd gnd cell_6t
Xbit_r29_c54 bl[54] br[54] wl[29] vdd gnd cell_6t
Xbit_r30_c54 bl[54] br[54] wl[30] vdd gnd cell_6t
Xbit_r31_c54 bl[54] br[54] wl[31] vdd gnd cell_6t
Xbit_r32_c54 bl[54] br[54] wl[32] vdd gnd cell_6t
Xbit_r33_c54 bl[54] br[54] wl[33] vdd gnd cell_6t
Xbit_r34_c54 bl[54] br[54] wl[34] vdd gnd cell_6t
Xbit_r35_c54 bl[54] br[54] wl[35] vdd gnd cell_6t
Xbit_r36_c54 bl[54] br[54] wl[36] vdd gnd cell_6t
Xbit_r37_c54 bl[54] br[54] wl[37] vdd gnd cell_6t
Xbit_r38_c54 bl[54] br[54] wl[38] vdd gnd cell_6t
Xbit_r39_c54 bl[54] br[54] wl[39] vdd gnd cell_6t
Xbit_r40_c54 bl[54] br[54] wl[40] vdd gnd cell_6t
Xbit_r41_c54 bl[54] br[54] wl[41] vdd gnd cell_6t
Xbit_r42_c54 bl[54] br[54] wl[42] vdd gnd cell_6t
Xbit_r43_c54 bl[54] br[54] wl[43] vdd gnd cell_6t
Xbit_r44_c54 bl[54] br[54] wl[44] vdd gnd cell_6t
Xbit_r45_c54 bl[54] br[54] wl[45] vdd gnd cell_6t
Xbit_r46_c54 bl[54] br[54] wl[46] vdd gnd cell_6t
Xbit_r47_c54 bl[54] br[54] wl[47] vdd gnd cell_6t
Xbit_r48_c54 bl[54] br[54] wl[48] vdd gnd cell_6t
Xbit_r49_c54 bl[54] br[54] wl[49] vdd gnd cell_6t
Xbit_r50_c54 bl[54] br[54] wl[50] vdd gnd cell_6t
Xbit_r51_c54 bl[54] br[54] wl[51] vdd gnd cell_6t
Xbit_r52_c54 bl[54] br[54] wl[52] vdd gnd cell_6t
Xbit_r53_c54 bl[54] br[54] wl[53] vdd gnd cell_6t
Xbit_r54_c54 bl[54] br[54] wl[54] vdd gnd cell_6t
Xbit_r55_c54 bl[54] br[54] wl[55] vdd gnd cell_6t
Xbit_r56_c54 bl[54] br[54] wl[56] vdd gnd cell_6t
Xbit_r57_c54 bl[54] br[54] wl[57] vdd gnd cell_6t
Xbit_r58_c54 bl[54] br[54] wl[58] vdd gnd cell_6t
Xbit_r59_c54 bl[54] br[54] wl[59] vdd gnd cell_6t
Xbit_r60_c54 bl[54] br[54] wl[60] vdd gnd cell_6t
Xbit_r61_c54 bl[54] br[54] wl[61] vdd gnd cell_6t
Xbit_r62_c54 bl[54] br[54] wl[62] vdd gnd cell_6t
Xbit_r63_c54 bl[54] br[54] wl[63] vdd gnd cell_6t
Xbit_r64_c54 bl[54] br[54] wl[64] vdd gnd cell_6t
Xbit_r65_c54 bl[54] br[54] wl[65] vdd gnd cell_6t
Xbit_r66_c54 bl[54] br[54] wl[66] vdd gnd cell_6t
Xbit_r67_c54 bl[54] br[54] wl[67] vdd gnd cell_6t
Xbit_r68_c54 bl[54] br[54] wl[68] vdd gnd cell_6t
Xbit_r69_c54 bl[54] br[54] wl[69] vdd gnd cell_6t
Xbit_r70_c54 bl[54] br[54] wl[70] vdd gnd cell_6t
Xbit_r71_c54 bl[54] br[54] wl[71] vdd gnd cell_6t
Xbit_r72_c54 bl[54] br[54] wl[72] vdd gnd cell_6t
Xbit_r73_c54 bl[54] br[54] wl[73] vdd gnd cell_6t
Xbit_r74_c54 bl[54] br[54] wl[74] vdd gnd cell_6t
Xbit_r75_c54 bl[54] br[54] wl[75] vdd gnd cell_6t
Xbit_r76_c54 bl[54] br[54] wl[76] vdd gnd cell_6t
Xbit_r77_c54 bl[54] br[54] wl[77] vdd gnd cell_6t
Xbit_r78_c54 bl[54] br[54] wl[78] vdd gnd cell_6t
Xbit_r79_c54 bl[54] br[54] wl[79] vdd gnd cell_6t
Xbit_r80_c54 bl[54] br[54] wl[80] vdd gnd cell_6t
Xbit_r81_c54 bl[54] br[54] wl[81] vdd gnd cell_6t
Xbit_r82_c54 bl[54] br[54] wl[82] vdd gnd cell_6t
Xbit_r83_c54 bl[54] br[54] wl[83] vdd gnd cell_6t
Xbit_r84_c54 bl[54] br[54] wl[84] vdd gnd cell_6t
Xbit_r85_c54 bl[54] br[54] wl[85] vdd gnd cell_6t
Xbit_r86_c54 bl[54] br[54] wl[86] vdd gnd cell_6t
Xbit_r87_c54 bl[54] br[54] wl[87] vdd gnd cell_6t
Xbit_r88_c54 bl[54] br[54] wl[88] vdd gnd cell_6t
Xbit_r89_c54 bl[54] br[54] wl[89] vdd gnd cell_6t
Xbit_r90_c54 bl[54] br[54] wl[90] vdd gnd cell_6t
Xbit_r91_c54 bl[54] br[54] wl[91] vdd gnd cell_6t
Xbit_r92_c54 bl[54] br[54] wl[92] vdd gnd cell_6t
Xbit_r93_c54 bl[54] br[54] wl[93] vdd gnd cell_6t
Xbit_r94_c54 bl[54] br[54] wl[94] vdd gnd cell_6t
Xbit_r95_c54 bl[54] br[54] wl[95] vdd gnd cell_6t
Xbit_r96_c54 bl[54] br[54] wl[96] vdd gnd cell_6t
Xbit_r97_c54 bl[54] br[54] wl[97] vdd gnd cell_6t
Xbit_r98_c54 bl[54] br[54] wl[98] vdd gnd cell_6t
Xbit_r99_c54 bl[54] br[54] wl[99] vdd gnd cell_6t
Xbit_r100_c54 bl[54] br[54] wl[100] vdd gnd cell_6t
Xbit_r101_c54 bl[54] br[54] wl[101] vdd gnd cell_6t
Xbit_r102_c54 bl[54] br[54] wl[102] vdd gnd cell_6t
Xbit_r103_c54 bl[54] br[54] wl[103] vdd gnd cell_6t
Xbit_r104_c54 bl[54] br[54] wl[104] vdd gnd cell_6t
Xbit_r105_c54 bl[54] br[54] wl[105] vdd gnd cell_6t
Xbit_r106_c54 bl[54] br[54] wl[106] vdd gnd cell_6t
Xbit_r107_c54 bl[54] br[54] wl[107] vdd gnd cell_6t
Xbit_r108_c54 bl[54] br[54] wl[108] vdd gnd cell_6t
Xbit_r109_c54 bl[54] br[54] wl[109] vdd gnd cell_6t
Xbit_r110_c54 bl[54] br[54] wl[110] vdd gnd cell_6t
Xbit_r111_c54 bl[54] br[54] wl[111] vdd gnd cell_6t
Xbit_r112_c54 bl[54] br[54] wl[112] vdd gnd cell_6t
Xbit_r113_c54 bl[54] br[54] wl[113] vdd gnd cell_6t
Xbit_r114_c54 bl[54] br[54] wl[114] vdd gnd cell_6t
Xbit_r115_c54 bl[54] br[54] wl[115] vdd gnd cell_6t
Xbit_r116_c54 bl[54] br[54] wl[116] vdd gnd cell_6t
Xbit_r117_c54 bl[54] br[54] wl[117] vdd gnd cell_6t
Xbit_r118_c54 bl[54] br[54] wl[118] vdd gnd cell_6t
Xbit_r119_c54 bl[54] br[54] wl[119] vdd gnd cell_6t
Xbit_r120_c54 bl[54] br[54] wl[120] vdd gnd cell_6t
Xbit_r121_c54 bl[54] br[54] wl[121] vdd gnd cell_6t
Xbit_r122_c54 bl[54] br[54] wl[122] vdd gnd cell_6t
Xbit_r123_c54 bl[54] br[54] wl[123] vdd gnd cell_6t
Xbit_r124_c54 bl[54] br[54] wl[124] vdd gnd cell_6t
Xbit_r125_c54 bl[54] br[54] wl[125] vdd gnd cell_6t
Xbit_r126_c54 bl[54] br[54] wl[126] vdd gnd cell_6t
Xbit_r127_c54 bl[54] br[54] wl[127] vdd gnd cell_6t
Xbit_r128_c54 bl[54] br[54] wl[128] vdd gnd cell_6t
Xbit_r129_c54 bl[54] br[54] wl[129] vdd gnd cell_6t
Xbit_r130_c54 bl[54] br[54] wl[130] vdd gnd cell_6t
Xbit_r131_c54 bl[54] br[54] wl[131] vdd gnd cell_6t
Xbit_r132_c54 bl[54] br[54] wl[132] vdd gnd cell_6t
Xbit_r133_c54 bl[54] br[54] wl[133] vdd gnd cell_6t
Xbit_r134_c54 bl[54] br[54] wl[134] vdd gnd cell_6t
Xbit_r135_c54 bl[54] br[54] wl[135] vdd gnd cell_6t
Xbit_r136_c54 bl[54] br[54] wl[136] vdd gnd cell_6t
Xbit_r137_c54 bl[54] br[54] wl[137] vdd gnd cell_6t
Xbit_r138_c54 bl[54] br[54] wl[138] vdd gnd cell_6t
Xbit_r139_c54 bl[54] br[54] wl[139] vdd gnd cell_6t
Xbit_r140_c54 bl[54] br[54] wl[140] vdd gnd cell_6t
Xbit_r141_c54 bl[54] br[54] wl[141] vdd gnd cell_6t
Xbit_r142_c54 bl[54] br[54] wl[142] vdd gnd cell_6t
Xbit_r143_c54 bl[54] br[54] wl[143] vdd gnd cell_6t
Xbit_r144_c54 bl[54] br[54] wl[144] vdd gnd cell_6t
Xbit_r145_c54 bl[54] br[54] wl[145] vdd gnd cell_6t
Xbit_r146_c54 bl[54] br[54] wl[146] vdd gnd cell_6t
Xbit_r147_c54 bl[54] br[54] wl[147] vdd gnd cell_6t
Xbit_r148_c54 bl[54] br[54] wl[148] vdd gnd cell_6t
Xbit_r149_c54 bl[54] br[54] wl[149] vdd gnd cell_6t
Xbit_r150_c54 bl[54] br[54] wl[150] vdd gnd cell_6t
Xbit_r151_c54 bl[54] br[54] wl[151] vdd gnd cell_6t
Xbit_r152_c54 bl[54] br[54] wl[152] vdd gnd cell_6t
Xbit_r153_c54 bl[54] br[54] wl[153] vdd gnd cell_6t
Xbit_r154_c54 bl[54] br[54] wl[154] vdd gnd cell_6t
Xbit_r155_c54 bl[54] br[54] wl[155] vdd gnd cell_6t
Xbit_r156_c54 bl[54] br[54] wl[156] vdd gnd cell_6t
Xbit_r157_c54 bl[54] br[54] wl[157] vdd gnd cell_6t
Xbit_r158_c54 bl[54] br[54] wl[158] vdd gnd cell_6t
Xbit_r159_c54 bl[54] br[54] wl[159] vdd gnd cell_6t
Xbit_r160_c54 bl[54] br[54] wl[160] vdd gnd cell_6t
Xbit_r161_c54 bl[54] br[54] wl[161] vdd gnd cell_6t
Xbit_r162_c54 bl[54] br[54] wl[162] vdd gnd cell_6t
Xbit_r163_c54 bl[54] br[54] wl[163] vdd gnd cell_6t
Xbit_r164_c54 bl[54] br[54] wl[164] vdd gnd cell_6t
Xbit_r165_c54 bl[54] br[54] wl[165] vdd gnd cell_6t
Xbit_r166_c54 bl[54] br[54] wl[166] vdd gnd cell_6t
Xbit_r167_c54 bl[54] br[54] wl[167] vdd gnd cell_6t
Xbit_r168_c54 bl[54] br[54] wl[168] vdd gnd cell_6t
Xbit_r169_c54 bl[54] br[54] wl[169] vdd gnd cell_6t
Xbit_r170_c54 bl[54] br[54] wl[170] vdd gnd cell_6t
Xbit_r171_c54 bl[54] br[54] wl[171] vdd gnd cell_6t
Xbit_r172_c54 bl[54] br[54] wl[172] vdd gnd cell_6t
Xbit_r173_c54 bl[54] br[54] wl[173] vdd gnd cell_6t
Xbit_r174_c54 bl[54] br[54] wl[174] vdd gnd cell_6t
Xbit_r175_c54 bl[54] br[54] wl[175] vdd gnd cell_6t
Xbit_r176_c54 bl[54] br[54] wl[176] vdd gnd cell_6t
Xbit_r177_c54 bl[54] br[54] wl[177] vdd gnd cell_6t
Xbit_r178_c54 bl[54] br[54] wl[178] vdd gnd cell_6t
Xbit_r179_c54 bl[54] br[54] wl[179] vdd gnd cell_6t
Xbit_r180_c54 bl[54] br[54] wl[180] vdd gnd cell_6t
Xbit_r181_c54 bl[54] br[54] wl[181] vdd gnd cell_6t
Xbit_r182_c54 bl[54] br[54] wl[182] vdd gnd cell_6t
Xbit_r183_c54 bl[54] br[54] wl[183] vdd gnd cell_6t
Xbit_r184_c54 bl[54] br[54] wl[184] vdd gnd cell_6t
Xbit_r185_c54 bl[54] br[54] wl[185] vdd gnd cell_6t
Xbit_r186_c54 bl[54] br[54] wl[186] vdd gnd cell_6t
Xbit_r187_c54 bl[54] br[54] wl[187] vdd gnd cell_6t
Xbit_r188_c54 bl[54] br[54] wl[188] vdd gnd cell_6t
Xbit_r189_c54 bl[54] br[54] wl[189] vdd gnd cell_6t
Xbit_r190_c54 bl[54] br[54] wl[190] vdd gnd cell_6t
Xbit_r191_c54 bl[54] br[54] wl[191] vdd gnd cell_6t
Xbit_r192_c54 bl[54] br[54] wl[192] vdd gnd cell_6t
Xbit_r193_c54 bl[54] br[54] wl[193] vdd gnd cell_6t
Xbit_r194_c54 bl[54] br[54] wl[194] vdd gnd cell_6t
Xbit_r195_c54 bl[54] br[54] wl[195] vdd gnd cell_6t
Xbit_r196_c54 bl[54] br[54] wl[196] vdd gnd cell_6t
Xbit_r197_c54 bl[54] br[54] wl[197] vdd gnd cell_6t
Xbit_r198_c54 bl[54] br[54] wl[198] vdd gnd cell_6t
Xbit_r199_c54 bl[54] br[54] wl[199] vdd gnd cell_6t
Xbit_r200_c54 bl[54] br[54] wl[200] vdd gnd cell_6t
Xbit_r201_c54 bl[54] br[54] wl[201] vdd gnd cell_6t
Xbit_r202_c54 bl[54] br[54] wl[202] vdd gnd cell_6t
Xbit_r203_c54 bl[54] br[54] wl[203] vdd gnd cell_6t
Xbit_r204_c54 bl[54] br[54] wl[204] vdd gnd cell_6t
Xbit_r205_c54 bl[54] br[54] wl[205] vdd gnd cell_6t
Xbit_r206_c54 bl[54] br[54] wl[206] vdd gnd cell_6t
Xbit_r207_c54 bl[54] br[54] wl[207] vdd gnd cell_6t
Xbit_r208_c54 bl[54] br[54] wl[208] vdd gnd cell_6t
Xbit_r209_c54 bl[54] br[54] wl[209] vdd gnd cell_6t
Xbit_r210_c54 bl[54] br[54] wl[210] vdd gnd cell_6t
Xbit_r211_c54 bl[54] br[54] wl[211] vdd gnd cell_6t
Xbit_r212_c54 bl[54] br[54] wl[212] vdd gnd cell_6t
Xbit_r213_c54 bl[54] br[54] wl[213] vdd gnd cell_6t
Xbit_r214_c54 bl[54] br[54] wl[214] vdd gnd cell_6t
Xbit_r215_c54 bl[54] br[54] wl[215] vdd gnd cell_6t
Xbit_r216_c54 bl[54] br[54] wl[216] vdd gnd cell_6t
Xbit_r217_c54 bl[54] br[54] wl[217] vdd gnd cell_6t
Xbit_r218_c54 bl[54] br[54] wl[218] vdd gnd cell_6t
Xbit_r219_c54 bl[54] br[54] wl[219] vdd gnd cell_6t
Xbit_r220_c54 bl[54] br[54] wl[220] vdd gnd cell_6t
Xbit_r221_c54 bl[54] br[54] wl[221] vdd gnd cell_6t
Xbit_r222_c54 bl[54] br[54] wl[222] vdd gnd cell_6t
Xbit_r223_c54 bl[54] br[54] wl[223] vdd gnd cell_6t
Xbit_r224_c54 bl[54] br[54] wl[224] vdd gnd cell_6t
Xbit_r225_c54 bl[54] br[54] wl[225] vdd gnd cell_6t
Xbit_r226_c54 bl[54] br[54] wl[226] vdd gnd cell_6t
Xbit_r227_c54 bl[54] br[54] wl[227] vdd gnd cell_6t
Xbit_r228_c54 bl[54] br[54] wl[228] vdd gnd cell_6t
Xbit_r229_c54 bl[54] br[54] wl[229] vdd gnd cell_6t
Xbit_r230_c54 bl[54] br[54] wl[230] vdd gnd cell_6t
Xbit_r231_c54 bl[54] br[54] wl[231] vdd gnd cell_6t
Xbit_r232_c54 bl[54] br[54] wl[232] vdd gnd cell_6t
Xbit_r233_c54 bl[54] br[54] wl[233] vdd gnd cell_6t
Xbit_r234_c54 bl[54] br[54] wl[234] vdd gnd cell_6t
Xbit_r235_c54 bl[54] br[54] wl[235] vdd gnd cell_6t
Xbit_r236_c54 bl[54] br[54] wl[236] vdd gnd cell_6t
Xbit_r237_c54 bl[54] br[54] wl[237] vdd gnd cell_6t
Xbit_r238_c54 bl[54] br[54] wl[238] vdd gnd cell_6t
Xbit_r239_c54 bl[54] br[54] wl[239] vdd gnd cell_6t
Xbit_r240_c54 bl[54] br[54] wl[240] vdd gnd cell_6t
Xbit_r241_c54 bl[54] br[54] wl[241] vdd gnd cell_6t
Xbit_r242_c54 bl[54] br[54] wl[242] vdd gnd cell_6t
Xbit_r243_c54 bl[54] br[54] wl[243] vdd gnd cell_6t
Xbit_r244_c54 bl[54] br[54] wl[244] vdd gnd cell_6t
Xbit_r245_c54 bl[54] br[54] wl[245] vdd gnd cell_6t
Xbit_r246_c54 bl[54] br[54] wl[246] vdd gnd cell_6t
Xbit_r247_c54 bl[54] br[54] wl[247] vdd gnd cell_6t
Xbit_r248_c54 bl[54] br[54] wl[248] vdd gnd cell_6t
Xbit_r249_c54 bl[54] br[54] wl[249] vdd gnd cell_6t
Xbit_r250_c54 bl[54] br[54] wl[250] vdd gnd cell_6t
Xbit_r251_c54 bl[54] br[54] wl[251] vdd gnd cell_6t
Xbit_r252_c54 bl[54] br[54] wl[252] vdd gnd cell_6t
Xbit_r253_c54 bl[54] br[54] wl[253] vdd gnd cell_6t
Xbit_r254_c54 bl[54] br[54] wl[254] vdd gnd cell_6t
Xbit_r255_c54 bl[54] br[54] wl[255] vdd gnd cell_6t
Xbit_r256_c54 bl[54] br[54] wl[256] vdd gnd cell_6t
Xbit_r257_c54 bl[54] br[54] wl[257] vdd gnd cell_6t
Xbit_r258_c54 bl[54] br[54] wl[258] vdd gnd cell_6t
Xbit_r259_c54 bl[54] br[54] wl[259] vdd gnd cell_6t
Xbit_r260_c54 bl[54] br[54] wl[260] vdd gnd cell_6t
Xbit_r261_c54 bl[54] br[54] wl[261] vdd gnd cell_6t
Xbit_r262_c54 bl[54] br[54] wl[262] vdd gnd cell_6t
Xbit_r263_c54 bl[54] br[54] wl[263] vdd gnd cell_6t
Xbit_r264_c54 bl[54] br[54] wl[264] vdd gnd cell_6t
Xbit_r265_c54 bl[54] br[54] wl[265] vdd gnd cell_6t
Xbit_r266_c54 bl[54] br[54] wl[266] vdd gnd cell_6t
Xbit_r267_c54 bl[54] br[54] wl[267] vdd gnd cell_6t
Xbit_r268_c54 bl[54] br[54] wl[268] vdd gnd cell_6t
Xbit_r269_c54 bl[54] br[54] wl[269] vdd gnd cell_6t
Xbit_r270_c54 bl[54] br[54] wl[270] vdd gnd cell_6t
Xbit_r271_c54 bl[54] br[54] wl[271] vdd gnd cell_6t
Xbit_r272_c54 bl[54] br[54] wl[272] vdd gnd cell_6t
Xbit_r273_c54 bl[54] br[54] wl[273] vdd gnd cell_6t
Xbit_r274_c54 bl[54] br[54] wl[274] vdd gnd cell_6t
Xbit_r275_c54 bl[54] br[54] wl[275] vdd gnd cell_6t
Xbit_r276_c54 bl[54] br[54] wl[276] vdd gnd cell_6t
Xbit_r277_c54 bl[54] br[54] wl[277] vdd gnd cell_6t
Xbit_r278_c54 bl[54] br[54] wl[278] vdd gnd cell_6t
Xbit_r279_c54 bl[54] br[54] wl[279] vdd gnd cell_6t
Xbit_r280_c54 bl[54] br[54] wl[280] vdd gnd cell_6t
Xbit_r281_c54 bl[54] br[54] wl[281] vdd gnd cell_6t
Xbit_r282_c54 bl[54] br[54] wl[282] vdd gnd cell_6t
Xbit_r283_c54 bl[54] br[54] wl[283] vdd gnd cell_6t
Xbit_r284_c54 bl[54] br[54] wl[284] vdd gnd cell_6t
Xbit_r285_c54 bl[54] br[54] wl[285] vdd gnd cell_6t
Xbit_r286_c54 bl[54] br[54] wl[286] vdd gnd cell_6t
Xbit_r287_c54 bl[54] br[54] wl[287] vdd gnd cell_6t
Xbit_r288_c54 bl[54] br[54] wl[288] vdd gnd cell_6t
Xbit_r289_c54 bl[54] br[54] wl[289] vdd gnd cell_6t
Xbit_r290_c54 bl[54] br[54] wl[290] vdd gnd cell_6t
Xbit_r291_c54 bl[54] br[54] wl[291] vdd gnd cell_6t
Xbit_r292_c54 bl[54] br[54] wl[292] vdd gnd cell_6t
Xbit_r293_c54 bl[54] br[54] wl[293] vdd gnd cell_6t
Xbit_r294_c54 bl[54] br[54] wl[294] vdd gnd cell_6t
Xbit_r295_c54 bl[54] br[54] wl[295] vdd gnd cell_6t
Xbit_r296_c54 bl[54] br[54] wl[296] vdd gnd cell_6t
Xbit_r297_c54 bl[54] br[54] wl[297] vdd gnd cell_6t
Xbit_r298_c54 bl[54] br[54] wl[298] vdd gnd cell_6t
Xbit_r299_c54 bl[54] br[54] wl[299] vdd gnd cell_6t
Xbit_r300_c54 bl[54] br[54] wl[300] vdd gnd cell_6t
Xbit_r301_c54 bl[54] br[54] wl[301] vdd gnd cell_6t
Xbit_r302_c54 bl[54] br[54] wl[302] vdd gnd cell_6t
Xbit_r303_c54 bl[54] br[54] wl[303] vdd gnd cell_6t
Xbit_r304_c54 bl[54] br[54] wl[304] vdd gnd cell_6t
Xbit_r305_c54 bl[54] br[54] wl[305] vdd gnd cell_6t
Xbit_r306_c54 bl[54] br[54] wl[306] vdd gnd cell_6t
Xbit_r307_c54 bl[54] br[54] wl[307] vdd gnd cell_6t
Xbit_r308_c54 bl[54] br[54] wl[308] vdd gnd cell_6t
Xbit_r309_c54 bl[54] br[54] wl[309] vdd gnd cell_6t
Xbit_r310_c54 bl[54] br[54] wl[310] vdd gnd cell_6t
Xbit_r311_c54 bl[54] br[54] wl[311] vdd gnd cell_6t
Xbit_r312_c54 bl[54] br[54] wl[312] vdd gnd cell_6t
Xbit_r313_c54 bl[54] br[54] wl[313] vdd gnd cell_6t
Xbit_r314_c54 bl[54] br[54] wl[314] vdd gnd cell_6t
Xbit_r315_c54 bl[54] br[54] wl[315] vdd gnd cell_6t
Xbit_r316_c54 bl[54] br[54] wl[316] vdd gnd cell_6t
Xbit_r317_c54 bl[54] br[54] wl[317] vdd gnd cell_6t
Xbit_r318_c54 bl[54] br[54] wl[318] vdd gnd cell_6t
Xbit_r319_c54 bl[54] br[54] wl[319] vdd gnd cell_6t
Xbit_r320_c54 bl[54] br[54] wl[320] vdd gnd cell_6t
Xbit_r321_c54 bl[54] br[54] wl[321] vdd gnd cell_6t
Xbit_r322_c54 bl[54] br[54] wl[322] vdd gnd cell_6t
Xbit_r323_c54 bl[54] br[54] wl[323] vdd gnd cell_6t
Xbit_r324_c54 bl[54] br[54] wl[324] vdd gnd cell_6t
Xbit_r325_c54 bl[54] br[54] wl[325] vdd gnd cell_6t
Xbit_r326_c54 bl[54] br[54] wl[326] vdd gnd cell_6t
Xbit_r327_c54 bl[54] br[54] wl[327] vdd gnd cell_6t
Xbit_r328_c54 bl[54] br[54] wl[328] vdd gnd cell_6t
Xbit_r329_c54 bl[54] br[54] wl[329] vdd gnd cell_6t
Xbit_r330_c54 bl[54] br[54] wl[330] vdd gnd cell_6t
Xbit_r331_c54 bl[54] br[54] wl[331] vdd gnd cell_6t
Xbit_r332_c54 bl[54] br[54] wl[332] vdd gnd cell_6t
Xbit_r333_c54 bl[54] br[54] wl[333] vdd gnd cell_6t
Xbit_r334_c54 bl[54] br[54] wl[334] vdd gnd cell_6t
Xbit_r335_c54 bl[54] br[54] wl[335] vdd gnd cell_6t
Xbit_r336_c54 bl[54] br[54] wl[336] vdd gnd cell_6t
Xbit_r337_c54 bl[54] br[54] wl[337] vdd gnd cell_6t
Xbit_r338_c54 bl[54] br[54] wl[338] vdd gnd cell_6t
Xbit_r339_c54 bl[54] br[54] wl[339] vdd gnd cell_6t
Xbit_r340_c54 bl[54] br[54] wl[340] vdd gnd cell_6t
Xbit_r341_c54 bl[54] br[54] wl[341] vdd gnd cell_6t
Xbit_r342_c54 bl[54] br[54] wl[342] vdd gnd cell_6t
Xbit_r343_c54 bl[54] br[54] wl[343] vdd gnd cell_6t
Xbit_r344_c54 bl[54] br[54] wl[344] vdd gnd cell_6t
Xbit_r345_c54 bl[54] br[54] wl[345] vdd gnd cell_6t
Xbit_r346_c54 bl[54] br[54] wl[346] vdd gnd cell_6t
Xbit_r347_c54 bl[54] br[54] wl[347] vdd gnd cell_6t
Xbit_r348_c54 bl[54] br[54] wl[348] vdd gnd cell_6t
Xbit_r349_c54 bl[54] br[54] wl[349] vdd gnd cell_6t
Xbit_r350_c54 bl[54] br[54] wl[350] vdd gnd cell_6t
Xbit_r351_c54 bl[54] br[54] wl[351] vdd gnd cell_6t
Xbit_r352_c54 bl[54] br[54] wl[352] vdd gnd cell_6t
Xbit_r353_c54 bl[54] br[54] wl[353] vdd gnd cell_6t
Xbit_r354_c54 bl[54] br[54] wl[354] vdd gnd cell_6t
Xbit_r355_c54 bl[54] br[54] wl[355] vdd gnd cell_6t
Xbit_r356_c54 bl[54] br[54] wl[356] vdd gnd cell_6t
Xbit_r357_c54 bl[54] br[54] wl[357] vdd gnd cell_6t
Xbit_r358_c54 bl[54] br[54] wl[358] vdd gnd cell_6t
Xbit_r359_c54 bl[54] br[54] wl[359] vdd gnd cell_6t
Xbit_r360_c54 bl[54] br[54] wl[360] vdd gnd cell_6t
Xbit_r361_c54 bl[54] br[54] wl[361] vdd gnd cell_6t
Xbit_r362_c54 bl[54] br[54] wl[362] vdd gnd cell_6t
Xbit_r363_c54 bl[54] br[54] wl[363] vdd gnd cell_6t
Xbit_r364_c54 bl[54] br[54] wl[364] vdd gnd cell_6t
Xbit_r365_c54 bl[54] br[54] wl[365] vdd gnd cell_6t
Xbit_r366_c54 bl[54] br[54] wl[366] vdd gnd cell_6t
Xbit_r367_c54 bl[54] br[54] wl[367] vdd gnd cell_6t
Xbit_r368_c54 bl[54] br[54] wl[368] vdd gnd cell_6t
Xbit_r369_c54 bl[54] br[54] wl[369] vdd gnd cell_6t
Xbit_r370_c54 bl[54] br[54] wl[370] vdd gnd cell_6t
Xbit_r371_c54 bl[54] br[54] wl[371] vdd gnd cell_6t
Xbit_r372_c54 bl[54] br[54] wl[372] vdd gnd cell_6t
Xbit_r373_c54 bl[54] br[54] wl[373] vdd gnd cell_6t
Xbit_r374_c54 bl[54] br[54] wl[374] vdd gnd cell_6t
Xbit_r375_c54 bl[54] br[54] wl[375] vdd gnd cell_6t
Xbit_r376_c54 bl[54] br[54] wl[376] vdd gnd cell_6t
Xbit_r377_c54 bl[54] br[54] wl[377] vdd gnd cell_6t
Xbit_r378_c54 bl[54] br[54] wl[378] vdd gnd cell_6t
Xbit_r379_c54 bl[54] br[54] wl[379] vdd gnd cell_6t
Xbit_r380_c54 bl[54] br[54] wl[380] vdd gnd cell_6t
Xbit_r381_c54 bl[54] br[54] wl[381] vdd gnd cell_6t
Xbit_r382_c54 bl[54] br[54] wl[382] vdd gnd cell_6t
Xbit_r383_c54 bl[54] br[54] wl[383] vdd gnd cell_6t
Xbit_r384_c54 bl[54] br[54] wl[384] vdd gnd cell_6t
Xbit_r385_c54 bl[54] br[54] wl[385] vdd gnd cell_6t
Xbit_r386_c54 bl[54] br[54] wl[386] vdd gnd cell_6t
Xbit_r387_c54 bl[54] br[54] wl[387] vdd gnd cell_6t
Xbit_r388_c54 bl[54] br[54] wl[388] vdd gnd cell_6t
Xbit_r389_c54 bl[54] br[54] wl[389] vdd gnd cell_6t
Xbit_r390_c54 bl[54] br[54] wl[390] vdd gnd cell_6t
Xbit_r391_c54 bl[54] br[54] wl[391] vdd gnd cell_6t
Xbit_r392_c54 bl[54] br[54] wl[392] vdd gnd cell_6t
Xbit_r393_c54 bl[54] br[54] wl[393] vdd gnd cell_6t
Xbit_r394_c54 bl[54] br[54] wl[394] vdd gnd cell_6t
Xbit_r395_c54 bl[54] br[54] wl[395] vdd gnd cell_6t
Xbit_r396_c54 bl[54] br[54] wl[396] vdd gnd cell_6t
Xbit_r397_c54 bl[54] br[54] wl[397] vdd gnd cell_6t
Xbit_r398_c54 bl[54] br[54] wl[398] vdd gnd cell_6t
Xbit_r399_c54 bl[54] br[54] wl[399] vdd gnd cell_6t
Xbit_r400_c54 bl[54] br[54] wl[400] vdd gnd cell_6t
Xbit_r401_c54 bl[54] br[54] wl[401] vdd gnd cell_6t
Xbit_r402_c54 bl[54] br[54] wl[402] vdd gnd cell_6t
Xbit_r403_c54 bl[54] br[54] wl[403] vdd gnd cell_6t
Xbit_r404_c54 bl[54] br[54] wl[404] vdd gnd cell_6t
Xbit_r405_c54 bl[54] br[54] wl[405] vdd gnd cell_6t
Xbit_r406_c54 bl[54] br[54] wl[406] vdd gnd cell_6t
Xbit_r407_c54 bl[54] br[54] wl[407] vdd gnd cell_6t
Xbit_r408_c54 bl[54] br[54] wl[408] vdd gnd cell_6t
Xbit_r409_c54 bl[54] br[54] wl[409] vdd gnd cell_6t
Xbit_r410_c54 bl[54] br[54] wl[410] vdd gnd cell_6t
Xbit_r411_c54 bl[54] br[54] wl[411] vdd gnd cell_6t
Xbit_r412_c54 bl[54] br[54] wl[412] vdd gnd cell_6t
Xbit_r413_c54 bl[54] br[54] wl[413] vdd gnd cell_6t
Xbit_r414_c54 bl[54] br[54] wl[414] vdd gnd cell_6t
Xbit_r415_c54 bl[54] br[54] wl[415] vdd gnd cell_6t
Xbit_r416_c54 bl[54] br[54] wl[416] vdd gnd cell_6t
Xbit_r417_c54 bl[54] br[54] wl[417] vdd gnd cell_6t
Xbit_r418_c54 bl[54] br[54] wl[418] vdd gnd cell_6t
Xbit_r419_c54 bl[54] br[54] wl[419] vdd gnd cell_6t
Xbit_r420_c54 bl[54] br[54] wl[420] vdd gnd cell_6t
Xbit_r421_c54 bl[54] br[54] wl[421] vdd gnd cell_6t
Xbit_r422_c54 bl[54] br[54] wl[422] vdd gnd cell_6t
Xbit_r423_c54 bl[54] br[54] wl[423] vdd gnd cell_6t
Xbit_r424_c54 bl[54] br[54] wl[424] vdd gnd cell_6t
Xbit_r425_c54 bl[54] br[54] wl[425] vdd gnd cell_6t
Xbit_r426_c54 bl[54] br[54] wl[426] vdd gnd cell_6t
Xbit_r427_c54 bl[54] br[54] wl[427] vdd gnd cell_6t
Xbit_r428_c54 bl[54] br[54] wl[428] vdd gnd cell_6t
Xbit_r429_c54 bl[54] br[54] wl[429] vdd gnd cell_6t
Xbit_r430_c54 bl[54] br[54] wl[430] vdd gnd cell_6t
Xbit_r431_c54 bl[54] br[54] wl[431] vdd gnd cell_6t
Xbit_r432_c54 bl[54] br[54] wl[432] vdd gnd cell_6t
Xbit_r433_c54 bl[54] br[54] wl[433] vdd gnd cell_6t
Xbit_r434_c54 bl[54] br[54] wl[434] vdd gnd cell_6t
Xbit_r435_c54 bl[54] br[54] wl[435] vdd gnd cell_6t
Xbit_r436_c54 bl[54] br[54] wl[436] vdd gnd cell_6t
Xbit_r437_c54 bl[54] br[54] wl[437] vdd gnd cell_6t
Xbit_r438_c54 bl[54] br[54] wl[438] vdd gnd cell_6t
Xbit_r439_c54 bl[54] br[54] wl[439] vdd gnd cell_6t
Xbit_r440_c54 bl[54] br[54] wl[440] vdd gnd cell_6t
Xbit_r441_c54 bl[54] br[54] wl[441] vdd gnd cell_6t
Xbit_r442_c54 bl[54] br[54] wl[442] vdd gnd cell_6t
Xbit_r443_c54 bl[54] br[54] wl[443] vdd gnd cell_6t
Xbit_r444_c54 bl[54] br[54] wl[444] vdd gnd cell_6t
Xbit_r445_c54 bl[54] br[54] wl[445] vdd gnd cell_6t
Xbit_r446_c54 bl[54] br[54] wl[446] vdd gnd cell_6t
Xbit_r447_c54 bl[54] br[54] wl[447] vdd gnd cell_6t
Xbit_r448_c54 bl[54] br[54] wl[448] vdd gnd cell_6t
Xbit_r449_c54 bl[54] br[54] wl[449] vdd gnd cell_6t
Xbit_r450_c54 bl[54] br[54] wl[450] vdd gnd cell_6t
Xbit_r451_c54 bl[54] br[54] wl[451] vdd gnd cell_6t
Xbit_r452_c54 bl[54] br[54] wl[452] vdd gnd cell_6t
Xbit_r453_c54 bl[54] br[54] wl[453] vdd gnd cell_6t
Xbit_r454_c54 bl[54] br[54] wl[454] vdd gnd cell_6t
Xbit_r455_c54 bl[54] br[54] wl[455] vdd gnd cell_6t
Xbit_r456_c54 bl[54] br[54] wl[456] vdd gnd cell_6t
Xbit_r457_c54 bl[54] br[54] wl[457] vdd gnd cell_6t
Xbit_r458_c54 bl[54] br[54] wl[458] vdd gnd cell_6t
Xbit_r459_c54 bl[54] br[54] wl[459] vdd gnd cell_6t
Xbit_r460_c54 bl[54] br[54] wl[460] vdd gnd cell_6t
Xbit_r461_c54 bl[54] br[54] wl[461] vdd gnd cell_6t
Xbit_r462_c54 bl[54] br[54] wl[462] vdd gnd cell_6t
Xbit_r463_c54 bl[54] br[54] wl[463] vdd gnd cell_6t
Xbit_r464_c54 bl[54] br[54] wl[464] vdd gnd cell_6t
Xbit_r465_c54 bl[54] br[54] wl[465] vdd gnd cell_6t
Xbit_r466_c54 bl[54] br[54] wl[466] vdd gnd cell_6t
Xbit_r467_c54 bl[54] br[54] wl[467] vdd gnd cell_6t
Xbit_r468_c54 bl[54] br[54] wl[468] vdd gnd cell_6t
Xbit_r469_c54 bl[54] br[54] wl[469] vdd gnd cell_6t
Xbit_r470_c54 bl[54] br[54] wl[470] vdd gnd cell_6t
Xbit_r471_c54 bl[54] br[54] wl[471] vdd gnd cell_6t
Xbit_r472_c54 bl[54] br[54] wl[472] vdd gnd cell_6t
Xbit_r473_c54 bl[54] br[54] wl[473] vdd gnd cell_6t
Xbit_r474_c54 bl[54] br[54] wl[474] vdd gnd cell_6t
Xbit_r475_c54 bl[54] br[54] wl[475] vdd gnd cell_6t
Xbit_r476_c54 bl[54] br[54] wl[476] vdd gnd cell_6t
Xbit_r477_c54 bl[54] br[54] wl[477] vdd gnd cell_6t
Xbit_r478_c54 bl[54] br[54] wl[478] vdd gnd cell_6t
Xbit_r479_c54 bl[54] br[54] wl[479] vdd gnd cell_6t
Xbit_r480_c54 bl[54] br[54] wl[480] vdd gnd cell_6t
Xbit_r481_c54 bl[54] br[54] wl[481] vdd gnd cell_6t
Xbit_r482_c54 bl[54] br[54] wl[482] vdd gnd cell_6t
Xbit_r483_c54 bl[54] br[54] wl[483] vdd gnd cell_6t
Xbit_r484_c54 bl[54] br[54] wl[484] vdd gnd cell_6t
Xbit_r485_c54 bl[54] br[54] wl[485] vdd gnd cell_6t
Xbit_r486_c54 bl[54] br[54] wl[486] vdd gnd cell_6t
Xbit_r487_c54 bl[54] br[54] wl[487] vdd gnd cell_6t
Xbit_r488_c54 bl[54] br[54] wl[488] vdd gnd cell_6t
Xbit_r489_c54 bl[54] br[54] wl[489] vdd gnd cell_6t
Xbit_r490_c54 bl[54] br[54] wl[490] vdd gnd cell_6t
Xbit_r491_c54 bl[54] br[54] wl[491] vdd gnd cell_6t
Xbit_r492_c54 bl[54] br[54] wl[492] vdd gnd cell_6t
Xbit_r493_c54 bl[54] br[54] wl[493] vdd gnd cell_6t
Xbit_r494_c54 bl[54] br[54] wl[494] vdd gnd cell_6t
Xbit_r495_c54 bl[54] br[54] wl[495] vdd gnd cell_6t
Xbit_r496_c54 bl[54] br[54] wl[496] vdd gnd cell_6t
Xbit_r497_c54 bl[54] br[54] wl[497] vdd gnd cell_6t
Xbit_r498_c54 bl[54] br[54] wl[498] vdd gnd cell_6t
Xbit_r499_c54 bl[54] br[54] wl[499] vdd gnd cell_6t
Xbit_r500_c54 bl[54] br[54] wl[500] vdd gnd cell_6t
Xbit_r501_c54 bl[54] br[54] wl[501] vdd gnd cell_6t
Xbit_r502_c54 bl[54] br[54] wl[502] vdd gnd cell_6t
Xbit_r503_c54 bl[54] br[54] wl[503] vdd gnd cell_6t
Xbit_r504_c54 bl[54] br[54] wl[504] vdd gnd cell_6t
Xbit_r505_c54 bl[54] br[54] wl[505] vdd gnd cell_6t
Xbit_r506_c54 bl[54] br[54] wl[506] vdd gnd cell_6t
Xbit_r507_c54 bl[54] br[54] wl[507] vdd gnd cell_6t
Xbit_r508_c54 bl[54] br[54] wl[508] vdd gnd cell_6t
Xbit_r509_c54 bl[54] br[54] wl[509] vdd gnd cell_6t
Xbit_r510_c54 bl[54] br[54] wl[510] vdd gnd cell_6t
Xbit_r511_c54 bl[54] br[54] wl[511] vdd gnd cell_6t
Xbit_r0_c55 bl[55] br[55] wl[0] vdd gnd cell_6t
Xbit_r1_c55 bl[55] br[55] wl[1] vdd gnd cell_6t
Xbit_r2_c55 bl[55] br[55] wl[2] vdd gnd cell_6t
Xbit_r3_c55 bl[55] br[55] wl[3] vdd gnd cell_6t
Xbit_r4_c55 bl[55] br[55] wl[4] vdd gnd cell_6t
Xbit_r5_c55 bl[55] br[55] wl[5] vdd gnd cell_6t
Xbit_r6_c55 bl[55] br[55] wl[6] vdd gnd cell_6t
Xbit_r7_c55 bl[55] br[55] wl[7] vdd gnd cell_6t
Xbit_r8_c55 bl[55] br[55] wl[8] vdd gnd cell_6t
Xbit_r9_c55 bl[55] br[55] wl[9] vdd gnd cell_6t
Xbit_r10_c55 bl[55] br[55] wl[10] vdd gnd cell_6t
Xbit_r11_c55 bl[55] br[55] wl[11] vdd gnd cell_6t
Xbit_r12_c55 bl[55] br[55] wl[12] vdd gnd cell_6t
Xbit_r13_c55 bl[55] br[55] wl[13] vdd gnd cell_6t
Xbit_r14_c55 bl[55] br[55] wl[14] vdd gnd cell_6t
Xbit_r15_c55 bl[55] br[55] wl[15] vdd gnd cell_6t
Xbit_r16_c55 bl[55] br[55] wl[16] vdd gnd cell_6t
Xbit_r17_c55 bl[55] br[55] wl[17] vdd gnd cell_6t
Xbit_r18_c55 bl[55] br[55] wl[18] vdd gnd cell_6t
Xbit_r19_c55 bl[55] br[55] wl[19] vdd gnd cell_6t
Xbit_r20_c55 bl[55] br[55] wl[20] vdd gnd cell_6t
Xbit_r21_c55 bl[55] br[55] wl[21] vdd gnd cell_6t
Xbit_r22_c55 bl[55] br[55] wl[22] vdd gnd cell_6t
Xbit_r23_c55 bl[55] br[55] wl[23] vdd gnd cell_6t
Xbit_r24_c55 bl[55] br[55] wl[24] vdd gnd cell_6t
Xbit_r25_c55 bl[55] br[55] wl[25] vdd gnd cell_6t
Xbit_r26_c55 bl[55] br[55] wl[26] vdd gnd cell_6t
Xbit_r27_c55 bl[55] br[55] wl[27] vdd gnd cell_6t
Xbit_r28_c55 bl[55] br[55] wl[28] vdd gnd cell_6t
Xbit_r29_c55 bl[55] br[55] wl[29] vdd gnd cell_6t
Xbit_r30_c55 bl[55] br[55] wl[30] vdd gnd cell_6t
Xbit_r31_c55 bl[55] br[55] wl[31] vdd gnd cell_6t
Xbit_r32_c55 bl[55] br[55] wl[32] vdd gnd cell_6t
Xbit_r33_c55 bl[55] br[55] wl[33] vdd gnd cell_6t
Xbit_r34_c55 bl[55] br[55] wl[34] vdd gnd cell_6t
Xbit_r35_c55 bl[55] br[55] wl[35] vdd gnd cell_6t
Xbit_r36_c55 bl[55] br[55] wl[36] vdd gnd cell_6t
Xbit_r37_c55 bl[55] br[55] wl[37] vdd gnd cell_6t
Xbit_r38_c55 bl[55] br[55] wl[38] vdd gnd cell_6t
Xbit_r39_c55 bl[55] br[55] wl[39] vdd gnd cell_6t
Xbit_r40_c55 bl[55] br[55] wl[40] vdd gnd cell_6t
Xbit_r41_c55 bl[55] br[55] wl[41] vdd gnd cell_6t
Xbit_r42_c55 bl[55] br[55] wl[42] vdd gnd cell_6t
Xbit_r43_c55 bl[55] br[55] wl[43] vdd gnd cell_6t
Xbit_r44_c55 bl[55] br[55] wl[44] vdd gnd cell_6t
Xbit_r45_c55 bl[55] br[55] wl[45] vdd gnd cell_6t
Xbit_r46_c55 bl[55] br[55] wl[46] vdd gnd cell_6t
Xbit_r47_c55 bl[55] br[55] wl[47] vdd gnd cell_6t
Xbit_r48_c55 bl[55] br[55] wl[48] vdd gnd cell_6t
Xbit_r49_c55 bl[55] br[55] wl[49] vdd gnd cell_6t
Xbit_r50_c55 bl[55] br[55] wl[50] vdd gnd cell_6t
Xbit_r51_c55 bl[55] br[55] wl[51] vdd gnd cell_6t
Xbit_r52_c55 bl[55] br[55] wl[52] vdd gnd cell_6t
Xbit_r53_c55 bl[55] br[55] wl[53] vdd gnd cell_6t
Xbit_r54_c55 bl[55] br[55] wl[54] vdd gnd cell_6t
Xbit_r55_c55 bl[55] br[55] wl[55] vdd gnd cell_6t
Xbit_r56_c55 bl[55] br[55] wl[56] vdd gnd cell_6t
Xbit_r57_c55 bl[55] br[55] wl[57] vdd gnd cell_6t
Xbit_r58_c55 bl[55] br[55] wl[58] vdd gnd cell_6t
Xbit_r59_c55 bl[55] br[55] wl[59] vdd gnd cell_6t
Xbit_r60_c55 bl[55] br[55] wl[60] vdd gnd cell_6t
Xbit_r61_c55 bl[55] br[55] wl[61] vdd gnd cell_6t
Xbit_r62_c55 bl[55] br[55] wl[62] vdd gnd cell_6t
Xbit_r63_c55 bl[55] br[55] wl[63] vdd gnd cell_6t
Xbit_r64_c55 bl[55] br[55] wl[64] vdd gnd cell_6t
Xbit_r65_c55 bl[55] br[55] wl[65] vdd gnd cell_6t
Xbit_r66_c55 bl[55] br[55] wl[66] vdd gnd cell_6t
Xbit_r67_c55 bl[55] br[55] wl[67] vdd gnd cell_6t
Xbit_r68_c55 bl[55] br[55] wl[68] vdd gnd cell_6t
Xbit_r69_c55 bl[55] br[55] wl[69] vdd gnd cell_6t
Xbit_r70_c55 bl[55] br[55] wl[70] vdd gnd cell_6t
Xbit_r71_c55 bl[55] br[55] wl[71] vdd gnd cell_6t
Xbit_r72_c55 bl[55] br[55] wl[72] vdd gnd cell_6t
Xbit_r73_c55 bl[55] br[55] wl[73] vdd gnd cell_6t
Xbit_r74_c55 bl[55] br[55] wl[74] vdd gnd cell_6t
Xbit_r75_c55 bl[55] br[55] wl[75] vdd gnd cell_6t
Xbit_r76_c55 bl[55] br[55] wl[76] vdd gnd cell_6t
Xbit_r77_c55 bl[55] br[55] wl[77] vdd gnd cell_6t
Xbit_r78_c55 bl[55] br[55] wl[78] vdd gnd cell_6t
Xbit_r79_c55 bl[55] br[55] wl[79] vdd gnd cell_6t
Xbit_r80_c55 bl[55] br[55] wl[80] vdd gnd cell_6t
Xbit_r81_c55 bl[55] br[55] wl[81] vdd gnd cell_6t
Xbit_r82_c55 bl[55] br[55] wl[82] vdd gnd cell_6t
Xbit_r83_c55 bl[55] br[55] wl[83] vdd gnd cell_6t
Xbit_r84_c55 bl[55] br[55] wl[84] vdd gnd cell_6t
Xbit_r85_c55 bl[55] br[55] wl[85] vdd gnd cell_6t
Xbit_r86_c55 bl[55] br[55] wl[86] vdd gnd cell_6t
Xbit_r87_c55 bl[55] br[55] wl[87] vdd gnd cell_6t
Xbit_r88_c55 bl[55] br[55] wl[88] vdd gnd cell_6t
Xbit_r89_c55 bl[55] br[55] wl[89] vdd gnd cell_6t
Xbit_r90_c55 bl[55] br[55] wl[90] vdd gnd cell_6t
Xbit_r91_c55 bl[55] br[55] wl[91] vdd gnd cell_6t
Xbit_r92_c55 bl[55] br[55] wl[92] vdd gnd cell_6t
Xbit_r93_c55 bl[55] br[55] wl[93] vdd gnd cell_6t
Xbit_r94_c55 bl[55] br[55] wl[94] vdd gnd cell_6t
Xbit_r95_c55 bl[55] br[55] wl[95] vdd gnd cell_6t
Xbit_r96_c55 bl[55] br[55] wl[96] vdd gnd cell_6t
Xbit_r97_c55 bl[55] br[55] wl[97] vdd gnd cell_6t
Xbit_r98_c55 bl[55] br[55] wl[98] vdd gnd cell_6t
Xbit_r99_c55 bl[55] br[55] wl[99] vdd gnd cell_6t
Xbit_r100_c55 bl[55] br[55] wl[100] vdd gnd cell_6t
Xbit_r101_c55 bl[55] br[55] wl[101] vdd gnd cell_6t
Xbit_r102_c55 bl[55] br[55] wl[102] vdd gnd cell_6t
Xbit_r103_c55 bl[55] br[55] wl[103] vdd gnd cell_6t
Xbit_r104_c55 bl[55] br[55] wl[104] vdd gnd cell_6t
Xbit_r105_c55 bl[55] br[55] wl[105] vdd gnd cell_6t
Xbit_r106_c55 bl[55] br[55] wl[106] vdd gnd cell_6t
Xbit_r107_c55 bl[55] br[55] wl[107] vdd gnd cell_6t
Xbit_r108_c55 bl[55] br[55] wl[108] vdd gnd cell_6t
Xbit_r109_c55 bl[55] br[55] wl[109] vdd gnd cell_6t
Xbit_r110_c55 bl[55] br[55] wl[110] vdd gnd cell_6t
Xbit_r111_c55 bl[55] br[55] wl[111] vdd gnd cell_6t
Xbit_r112_c55 bl[55] br[55] wl[112] vdd gnd cell_6t
Xbit_r113_c55 bl[55] br[55] wl[113] vdd gnd cell_6t
Xbit_r114_c55 bl[55] br[55] wl[114] vdd gnd cell_6t
Xbit_r115_c55 bl[55] br[55] wl[115] vdd gnd cell_6t
Xbit_r116_c55 bl[55] br[55] wl[116] vdd gnd cell_6t
Xbit_r117_c55 bl[55] br[55] wl[117] vdd gnd cell_6t
Xbit_r118_c55 bl[55] br[55] wl[118] vdd gnd cell_6t
Xbit_r119_c55 bl[55] br[55] wl[119] vdd gnd cell_6t
Xbit_r120_c55 bl[55] br[55] wl[120] vdd gnd cell_6t
Xbit_r121_c55 bl[55] br[55] wl[121] vdd gnd cell_6t
Xbit_r122_c55 bl[55] br[55] wl[122] vdd gnd cell_6t
Xbit_r123_c55 bl[55] br[55] wl[123] vdd gnd cell_6t
Xbit_r124_c55 bl[55] br[55] wl[124] vdd gnd cell_6t
Xbit_r125_c55 bl[55] br[55] wl[125] vdd gnd cell_6t
Xbit_r126_c55 bl[55] br[55] wl[126] vdd gnd cell_6t
Xbit_r127_c55 bl[55] br[55] wl[127] vdd gnd cell_6t
Xbit_r128_c55 bl[55] br[55] wl[128] vdd gnd cell_6t
Xbit_r129_c55 bl[55] br[55] wl[129] vdd gnd cell_6t
Xbit_r130_c55 bl[55] br[55] wl[130] vdd gnd cell_6t
Xbit_r131_c55 bl[55] br[55] wl[131] vdd gnd cell_6t
Xbit_r132_c55 bl[55] br[55] wl[132] vdd gnd cell_6t
Xbit_r133_c55 bl[55] br[55] wl[133] vdd gnd cell_6t
Xbit_r134_c55 bl[55] br[55] wl[134] vdd gnd cell_6t
Xbit_r135_c55 bl[55] br[55] wl[135] vdd gnd cell_6t
Xbit_r136_c55 bl[55] br[55] wl[136] vdd gnd cell_6t
Xbit_r137_c55 bl[55] br[55] wl[137] vdd gnd cell_6t
Xbit_r138_c55 bl[55] br[55] wl[138] vdd gnd cell_6t
Xbit_r139_c55 bl[55] br[55] wl[139] vdd gnd cell_6t
Xbit_r140_c55 bl[55] br[55] wl[140] vdd gnd cell_6t
Xbit_r141_c55 bl[55] br[55] wl[141] vdd gnd cell_6t
Xbit_r142_c55 bl[55] br[55] wl[142] vdd gnd cell_6t
Xbit_r143_c55 bl[55] br[55] wl[143] vdd gnd cell_6t
Xbit_r144_c55 bl[55] br[55] wl[144] vdd gnd cell_6t
Xbit_r145_c55 bl[55] br[55] wl[145] vdd gnd cell_6t
Xbit_r146_c55 bl[55] br[55] wl[146] vdd gnd cell_6t
Xbit_r147_c55 bl[55] br[55] wl[147] vdd gnd cell_6t
Xbit_r148_c55 bl[55] br[55] wl[148] vdd gnd cell_6t
Xbit_r149_c55 bl[55] br[55] wl[149] vdd gnd cell_6t
Xbit_r150_c55 bl[55] br[55] wl[150] vdd gnd cell_6t
Xbit_r151_c55 bl[55] br[55] wl[151] vdd gnd cell_6t
Xbit_r152_c55 bl[55] br[55] wl[152] vdd gnd cell_6t
Xbit_r153_c55 bl[55] br[55] wl[153] vdd gnd cell_6t
Xbit_r154_c55 bl[55] br[55] wl[154] vdd gnd cell_6t
Xbit_r155_c55 bl[55] br[55] wl[155] vdd gnd cell_6t
Xbit_r156_c55 bl[55] br[55] wl[156] vdd gnd cell_6t
Xbit_r157_c55 bl[55] br[55] wl[157] vdd gnd cell_6t
Xbit_r158_c55 bl[55] br[55] wl[158] vdd gnd cell_6t
Xbit_r159_c55 bl[55] br[55] wl[159] vdd gnd cell_6t
Xbit_r160_c55 bl[55] br[55] wl[160] vdd gnd cell_6t
Xbit_r161_c55 bl[55] br[55] wl[161] vdd gnd cell_6t
Xbit_r162_c55 bl[55] br[55] wl[162] vdd gnd cell_6t
Xbit_r163_c55 bl[55] br[55] wl[163] vdd gnd cell_6t
Xbit_r164_c55 bl[55] br[55] wl[164] vdd gnd cell_6t
Xbit_r165_c55 bl[55] br[55] wl[165] vdd gnd cell_6t
Xbit_r166_c55 bl[55] br[55] wl[166] vdd gnd cell_6t
Xbit_r167_c55 bl[55] br[55] wl[167] vdd gnd cell_6t
Xbit_r168_c55 bl[55] br[55] wl[168] vdd gnd cell_6t
Xbit_r169_c55 bl[55] br[55] wl[169] vdd gnd cell_6t
Xbit_r170_c55 bl[55] br[55] wl[170] vdd gnd cell_6t
Xbit_r171_c55 bl[55] br[55] wl[171] vdd gnd cell_6t
Xbit_r172_c55 bl[55] br[55] wl[172] vdd gnd cell_6t
Xbit_r173_c55 bl[55] br[55] wl[173] vdd gnd cell_6t
Xbit_r174_c55 bl[55] br[55] wl[174] vdd gnd cell_6t
Xbit_r175_c55 bl[55] br[55] wl[175] vdd gnd cell_6t
Xbit_r176_c55 bl[55] br[55] wl[176] vdd gnd cell_6t
Xbit_r177_c55 bl[55] br[55] wl[177] vdd gnd cell_6t
Xbit_r178_c55 bl[55] br[55] wl[178] vdd gnd cell_6t
Xbit_r179_c55 bl[55] br[55] wl[179] vdd gnd cell_6t
Xbit_r180_c55 bl[55] br[55] wl[180] vdd gnd cell_6t
Xbit_r181_c55 bl[55] br[55] wl[181] vdd gnd cell_6t
Xbit_r182_c55 bl[55] br[55] wl[182] vdd gnd cell_6t
Xbit_r183_c55 bl[55] br[55] wl[183] vdd gnd cell_6t
Xbit_r184_c55 bl[55] br[55] wl[184] vdd gnd cell_6t
Xbit_r185_c55 bl[55] br[55] wl[185] vdd gnd cell_6t
Xbit_r186_c55 bl[55] br[55] wl[186] vdd gnd cell_6t
Xbit_r187_c55 bl[55] br[55] wl[187] vdd gnd cell_6t
Xbit_r188_c55 bl[55] br[55] wl[188] vdd gnd cell_6t
Xbit_r189_c55 bl[55] br[55] wl[189] vdd gnd cell_6t
Xbit_r190_c55 bl[55] br[55] wl[190] vdd gnd cell_6t
Xbit_r191_c55 bl[55] br[55] wl[191] vdd gnd cell_6t
Xbit_r192_c55 bl[55] br[55] wl[192] vdd gnd cell_6t
Xbit_r193_c55 bl[55] br[55] wl[193] vdd gnd cell_6t
Xbit_r194_c55 bl[55] br[55] wl[194] vdd gnd cell_6t
Xbit_r195_c55 bl[55] br[55] wl[195] vdd gnd cell_6t
Xbit_r196_c55 bl[55] br[55] wl[196] vdd gnd cell_6t
Xbit_r197_c55 bl[55] br[55] wl[197] vdd gnd cell_6t
Xbit_r198_c55 bl[55] br[55] wl[198] vdd gnd cell_6t
Xbit_r199_c55 bl[55] br[55] wl[199] vdd gnd cell_6t
Xbit_r200_c55 bl[55] br[55] wl[200] vdd gnd cell_6t
Xbit_r201_c55 bl[55] br[55] wl[201] vdd gnd cell_6t
Xbit_r202_c55 bl[55] br[55] wl[202] vdd gnd cell_6t
Xbit_r203_c55 bl[55] br[55] wl[203] vdd gnd cell_6t
Xbit_r204_c55 bl[55] br[55] wl[204] vdd gnd cell_6t
Xbit_r205_c55 bl[55] br[55] wl[205] vdd gnd cell_6t
Xbit_r206_c55 bl[55] br[55] wl[206] vdd gnd cell_6t
Xbit_r207_c55 bl[55] br[55] wl[207] vdd gnd cell_6t
Xbit_r208_c55 bl[55] br[55] wl[208] vdd gnd cell_6t
Xbit_r209_c55 bl[55] br[55] wl[209] vdd gnd cell_6t
Xbit_r210_c55 bl[55] br[55] wl[210] vdd gnd cell_6t
Xbit_r211_c55 bl[55] br[55] wl[211] vdd gnd cell_6t
Xbit_r212_c55 bl[55] br[55] wl[212] vdd gnd cell_6t
Xbit_r213_c55 bl[55] br[55] wl[213] vdd gnd cell_6t
Xbit_r214_c55 bl[55] br[55] wl[214] vdd gnd cell_6t
Xbit_r215_c55 bl[55] br[55] wl[215] vdd gnd cell_6t
Xbit_r216_c55 bl[55] br[55] wl[216] vdd gnd cell_6t
Xbit_r217_c55 bl[55] br[55] wl[217] vdd gnd cell_6t
Xbit_r218_c55 bl[55] br[55] wl[218] vdd gnd cell_6t
Xbit_r219_c55 bl[55] br[55] wl[219] vdd gnd cell_6t
Xbit_r220_c55 bl[55] br[55] wl[220] vdd gnd cell_6t
Xbit_r221_c55 bl[55] br[55] wl[221] vdd gnd cell_6t
Xbit_r222_c55 bl[55] br[55] wl[222] vdd gnd cell_6t
Xbit_r223_c55 bl[55] br[55] wl[223] vdd gnd cell_6t
Xbit_r224_c55 bl[55] br[55] wl[224] vdd gnd cell_6t
Xbit_r225_c55 bl[55] br[55] wl[225] vdd gnd cell_6t
Xbit_r226_c55 bl[55] br[55] wl[226] vdd gnd cell_6t
Xbit_r227_c55 bl[55] br[55] wl[227] vdd gnd cell_6t
Xbit_r228_c55 bl[55] br[55] wl[228] vdd gnd cell_6t
Xbit_r229_c55 bl[55] br[55] wl[229] vdd gnd cell_6t
Xbit_r230_c55 bl[55] br[55] wl[230] vdd gnd cell_6t
Xbit_r231_c55 bl[55] br[55] wl[231] vdd gnd cell_6t
Xbit_r232_c55 bl[55] br[55] wl[232] vdd gnd cell_6t
Xbit_r233_c55 bl[55] br[55] wl[233] vdd gnd cell_6t
Xbit_r234_c55 bl[55] br[55] wl[234] vdd gnd cell_6t
Xbit_r235_c55 bl[55] br[55] wl[235] vdd gnd cell_6t
Xbit_r236_c55 bl[55] br[55] wl[236] vdd gnd cell_6t
Xbit_r237_c55 bl[55] br[55] wl[237] vdd gnd cell_6t
Xbit_r238_c55 bl[55] br[55] wl[238] vdd gnd cell_6t
Xbit_r239_c55 bl[55] br[55] wl[239] vdd gnd cell_6t
Xbit_r240_c55 bl[55] br[55] wl[240] vdd gnd cell_6t
Xbit_r241_c55 bl[55] br[55] wl[241] vdd gnd cell_6t
Xbit_r242_c55 bl[55] br[55] wl[242] vdd gnd cell_6t
Xbit_r243_c55 bl[55] br[55] wl[243] vdd gnd cell_6t
Xbit_r244_c55 bl[55] br[55] wl[244] vdd gnd cell_6t
Xbit_r245_c55 bl[55] br[55] wl[245] vdd gnd cell_6t
Xbit_r246_c55 bl[55] br[55] wl[246] vdd gnd cell_6t
Xbit_r247_c55 bl[55] br[55] wl[247] vdd gnd cell_6t
Xbit_r248_c55 bl[55] br[55] wl[248] vdd gnd cell_6t
Xbit_r249_c55 bl[55] br[55] wl[249] vdd gnd cell_6t
Xbit_r250_c55 bl[55] br[55] wl[250] vdd gnd cell_6t
Xbit_r251_c55 bl[55] br[55] wl[251] vdd gnd cell_6t
Xbit_r252_c55 bl[55] br[55] wl[252] vdd gnd cell_6t
Xbit_r253_c55 bl[55] br[55] wl[253] vdd gnd cell_6t
Xbit_r254_c55 bl[55] br[55] wl[254] vdd gnd cell_6t
Xbit_r255_c55 bl[55] br[55] wl[255] vdd gnd cell_6t
Xbit_r256_c55 bl[55] br[55] wl[256] vdd gnd cell_6t
Xbit_r257_c55 bl[55] br[55] wl[257] vdd gnd cell_6t
Xbit_r258_c55 bl[55] br[55] wl[258] vdd gnd cell_6t
Xbit_r259_c55 bl[55] br[55] wl[259] vdd gnd cell_6t
Xbit_r260_c55 bl[55] br[55] wl[260] vdd gnd cell_6t
Xbit_r261_c55 bl[55] br[55] wl[261] vdd gnd cell_6t
Xbit_r262_c55 bl[55] br[55] wl[262] vdd gnd cell_6t
Xbit_r263_c55 bl[55] br[55] wl[263] vdd gnd cell_6t
Xbit_r264_c55 bl[55] br[55] wl[264] vdd gnd cell_6t
Xbit_r265_c55 bl[55] br[55] wl[265] vdd gnd cell_6t
Xbit_r266_c55 bl[55] br[55] wl[266] vdd gnd cell_6t
Xbit_r267_c55 bl[55] br[55] wl[267] vdd gnd cell_6t
Xbit_r268_c55 bl[55] br[55] wl[268] vdd gnd cell_6t
Xbit_r269_c55 bl[55] br[55] wl[269] vdd gnd cell_6t
Xbit_r270_c55 bl[55] br[55] wl[270] vdd gnd cell_6t
Xbit_r271_c55 bl[55] br[55] wl[271] vdd gnd cell_6t
Xbit_r272_c55 bl[55] br[55] wl[272] vdd gnd cell_6t
Xbit_r273_c55 bl[55] br[55] wl[273] vdd gnd cell_6t
Xbit_r274_c55 bl[55] br[55] wl[274] vdd gnd cell_6t
Xbit_r275_c55 bl[55] br[55] wl[275] vdd gnd cell_6t
Xbit_r276_c55 bl[55] br[55] wl[276] vdd gnd cell_6t
Xbit_r277_c55 bl[55] br[55] wl[277] vdd gnd cell_6t
Xbit_r278_c55 bl[55] br[55] wl[278] vdd gnd cell_6t
Xbit_r279_c55 bl[55] br[55] wl[279] vdd gnd cell_6t
Xbit_r280_c55 bl[55] br[55] wl[280] vdd gnd cell_6t
Xbit_r281_c55 bl[55] br[55] wl[281] vdd gnd cell_6t
Xbit_r282_c55 bl[55] br[55] wl[282] vdd gnd cell_6t
Xbit_r283_c55 bl[55] br[55] wl[283] vdd gnd cell_6t
Xbit_r284_c55 bl[55] br[55] wl[284] vdd gnd cell_6t
Xbit_r285_c55 bl[55] br[55] wl[285] vdd gnd cell_6t
Xbit_r286_c55 bl[55] br[55] wl[286] vdd gnd cell_6t
Xbit_r287_c55 bl[55] br[55] wl[287] vdd gnd cell_6t
Xbit_r288_c55 bl[55] br[55] wl[288] vdd gnd cell_6t
Xbit_r289_c55 bl[55] br[55] wl[289] vdd gnd cell_6t
Xbit_r290_c55 bl[55] br[55] wl[290] vdd gnd cell_6t
Xbit_r291_c55 bl[55] br[55] wl[291] vdd gnd cell_6t
Xbit_r292_c55 bl[55] br[55] wl[292] vdd gnd cell_6t
Xbit_r293_c55 bl[55] br[55] wl[293] vdd gnd cell_6t
Xbit_r294_c55 bl[55] br[55] wl[294] vdd gnd cell_6t
Xbit_r295_c55 bl[55] br[55] wl[295] vdd gnd cell_6t
Xbit_r296_c55 bl[55] br[55] wl[296] vdd gnd cell_6t
Xbit_r297_c55 bl[55] br[55] wl[297] vdd gnd cell_6t
Xbit_r298_c55 bl[55] br[55] wl[298] vdd gnd cell_6t
Xbit_r299_c55 bl[55] br[55] wl[299] vdd gnd cell_6t
Xbit_r300_c55 bl[55] br[55] wl[300] vdd gnd cell_6t
Xbit_r301_c55 bl[55] br[55] wl[301] vdd gnd cell_6t
Xbit_r302_c55 bl[55] br[55] wl[302] vdd gnd cell_6t
Xbit_r303_c55 bl[55] br[55] wl[303] vdd gnd cell_6t
Xbit_r304_c55 bl[55] br[55] wl[304] vdd gnd cell_6t
Xbit_r305_c55 bl[55] br[55] wl[305] vdd gnd cell_6t
Xbit_r306_c55 bl[55] br[55] wl[306] vdd gnd cell_6t
Xbit_r307_c55 bl[55] br[55] wl[307] vdd gnd cell_6t
Xbit_r308_c55 bl[55] br[55] wl[308] vdd gnd cell_6t
Xbit_r309_c55 bl[55] br[55] wl[309] vdd gnd cell_6t
Xbit_r310_c55 bl[55] br[55] wl[310] vdd gnd cell_6t
Xbit_r311_c55 bl[55] br[55] wl[311] vdd gnd cell_6t
Xbit_r312_c55 bl[55] br[55] wl[312] vdd gnd cell_6t
Xbit_r313_c55 bl[55] br[55] wl[313] vdd gnd cell_6t
Xbit_r314_c55 bl[55] br[55] wl[314] vdd gnd cell_6t
Xbit_r315_c55 bl[55] br[55] wl[315] vdd gnd cell_6t
Xbit_r316_c55 bl[55] br[55] wl[316] vdd gnd cell_6t
Xbit_r317_c55 bl[55] br[55] wl[317] vdd gnd cell_6t
Xbit_r318_c55 bl[55] br[55] wl[318] vdd gnd cell_6t
Xbit_r319_c55 bl[55] br[55] wl[319] vdd gnd cell_6t
Xbit_r320_c55 bl[55] br[55] wl[320] vdd gnd cell_6t
Xbit_r321_c55 bl[55] br[55] wl[321] vdd gnd cell_6t
Xbit_r322_c55 bl[55] br[55] wl[322] vdd gnd cell_6t
Xbit_r323_c55 bl[55] br[55] wl[323] vdd gnd cell_6t
Xbit_r324_c55 bl[55] br[55] wl[324] vdd gnd cell_6t
Xbit_r325_c55 bl[55] br[55] wl[325] vdd gnd cell_6t
Xbit_r326_c55 bl[55] br[55] wl[326] vdd gnd cell_6t
Xbit_r327_c55 bl[55] br[55] wl[327] vdd gnd cell_6t
Xbit_r328_c55 bl[55] br[55] wl[328] vdd gnd cell_6t
Xbit_r329_c55 bl[55] br[55] wl[329] vdd gnd cell_6t
Xbit_r330_c55 bl[55] br[55] wl[330] vdd gnd cell_6t
Xbit_r331_c55 bl[55] br[55] wl[331] vdd gnd cell_6t
Xbit_r332_c55 bl[55] br[55] wl[332] vdd gnd cell_6t
Xbit_r333_c55 bl[55] br[55] wl[333] vdd gnd cell_6t
Xbit_r334_c55 bl[55] br[55] wl[334] vdd gnd cell_6t
Xbit_r335_c55 bl[55] br[55] wl[335] vdd gnd cell_6t
Xbit_r336_c55 bl[55] br[55] wl[336] vdd gnd cell_6t
Xbit_r337_c55 bl[55] br[55] wl[337] vdd gnd cell_6t
Xbit_r338_c55 bl[55] br[55] wl[338] vdd gnd cell_6t
Xbit_r339_c55 bl[55] br[55] wl[339] vdd gnd cell_6t
Xbit_r340_c55 bl[55] br[55] wl[340] vdd gnd cell_6t
Xbit_r341_c55 bl[55] br[55] wl[341] vdd gnd cell_6t
Xbit_r342_c55 bl[55] br[55] wl[342] vdd gnd cell_6t
Xbit_r343_c55 bl[55] br[55] wl[343] vdd gnd cell_6t
Xbit_r344_c55 bl[55] br[55] wl[344] vdd gnd cell_6t
Xbit_r345_c55 bl[55] br[55] wl[345] vdd gnd cell_6t
Xbit_r346_c55 bl[55] br[55] wl[346] vdd gnd cell_6t
Xbit_r347_c55 bl[55] br[55] wl[347] vdd gnd cell_6t
Xbit_r348_c55 bl[55] br[55] wl[348] vdd gnd cell_6t
Xbit_r349_c55 bl[55] br[55] wl[349] vdd gnd cell_6t
Xbit_r350_c55 bl[55] br[55] wl[350] vdd gnd cell_6t
Xbit_r351_c55 bl[55] br[55] wl[351] vdd gnd cell_6t
Xbit_r352_c55 bl[55] br[55] wl[352] vdd gnd cell_6t
Xbit_r353_c55 bl[55] br[55] wl[353] vdd gnd cell_6t
Xbit_r354_c55 bl[55] br[55] wl[354] vdd gnd cell_6t
Xbit_r355_c55 bl[55] br[55] wl[355] vdd gnd cell_6t
Xbit_r356_c55 bl[55] br[55] wl[356] vdd gnd cell_6t
Xbit_r357_c55 bl[55] br[55] wl[357] vdd gnd cell_6t
Xbit_r358_c55 bl[55] br[55] wl[358] vdd gnd cell_6t
Xbit_r359_c55 bl[55] br[55] wl[359] vdd gnd cell_6t
Xbit_r360_c55 bl[55] br[55] wl[360] vdd gnd cell_6t
Xbit_r361_c55 bl[55] br[55] wl[361] vdd gnd cell_6t
Xbit_r362_c55 bl[55] br[55] wl[362] vdd gnd cell_6t
Xbit_r363_c55 bl[55] br[55] wl[363] vdd gnd cell_6t
Xbit_r364_c55 bl[55] br[55] wl[364] vdd gnd cell_6t
Xbit_r365_c55 bl[55] br[55] wl[365] vdd gnd cell_6t
Xbit_r366_c55 bl[55] br[55] wl[366] vdd gnd cell_6t
Xbit_r367_c55 bl[55] br[55] wl[367] vdd gnd cell_6t
Xbit_r368_c55 bl[55] br[55] wl[368] vdd gnd cell_6t
Xbit_r369_c55 bl[55] br[55] wl[369] vdd gnd cell_6t
Xbit_r370_c55 bl[55] br[55] wl[370] vdd gnd cell_6t
Xbit_r371_c55 bl[55] br[55] wl[371] vdd gnd cell_6t
Xbit_r372_c55 bl[55] br[55] wl[372] vdd gnd cell_6t
Xbit_r373_c55 bl[55] br[55] wl[373] vdd gnd cell_6t
Xbit_r374_c55 bl[55] br[55] wl[374] vdd gnd cell_6t
Xbit_r375_c55 bl[55] br[55] wl[375] vdd gnd cell_6t
Xbit_r376_c55 bl[55] br[55] wl[376] vdd gnd cell_6t
Xbit_r377_c55 bl[55] br[55] wl[377] vdd gnd cell_6t
Xbit_r378_c55 bl[55] br[55] wl[378] vdd gnd cell_6t
Xbit_r379_c55 bl[55] br[55] wl[379] vdd gnd cell_6t
Xbit_r380_c55 bl[55] br[55] wl[380] vdd gnd cell_6t
Xbit_r381_c55 bl[55] br[55] wl[381] vdd gnd cell_6t
Xbit_r382_c55 bl[55] br[55] wl[382] vdd gnd cell_6t
Xbit_r383_c55 bl[55] br[55] wl[383] vdd gnd cell_6t
Xbit_r384_c55 bl[55] br[55] wl[384] vdd gnd cell_6t
Xbit_r385_c55 bl[55] br[55] wl[385] vdd gnd cell_6t
Xbit_r386_c55 bl[55] br[55] wl[386] vdd gnd cell_6t
Xbit_r387_c55 bl[55] br[55] wl[387] vdd gnd cell_6t
Xbit_r388_c55 bl[55] br[55] wl[388] vdd gnd cell_6t
Xbit_r389_c55 bl[55] br[55] wl[389] vdd gnd cell_6t
Xbit_r390_c55 bl[55] br[55] wl[390] vdd gnd cell_6t
Xbit_r391_c55 bl[55] br[55] wl[391] vdd gnd cell_6t
Xbit_r392_c55 bl[55] br[55] wl[392] vdd gnd cell_6t
Xbit_r393_c55 bl[55] br[55] wl[393] vdd gnd cell_6t
Xbit_r394_c55 bl[55] br[55] wl[394] vdd gnd cell_6t
Xbit_r395_c55 bl[55] br[55] wl[395] vdd gnd cell_6t
Xbit_r396_c55 bl[55] br[55] wl[396] vdd gnd cell_6t
Xbit_r397_c55 bl[55] br[55] wl[397] vdd gnd cell_6t
Xbit_r398_c55 bl[55] br[55] wl[398] vdd gnd cell_6t
Xbit_r399_c55 bl[55] br[55] wl[399] vdd gnd cell_6t
Xbit_r400_c55 bl[55] br[55] wl[400] vdd gnd cell_6t
Xbit_r401_c55 bl[55] br[55] wl[401] vdd gnd cell_6t
Xbit_r402_c55 bl[55] br[55] wl[402] vdd gnd cell_6t
Xbit_r403_c55 bl[55] br[55] wl[403] vdd gnd cell_6t
Xbit_r404_c55 bl[55] br[55] wl[404] vdd gnd cell_6t
Xbit_r405_c55 bl[55] br[55] wl[405] vdd gnd cell_6t
Xbit_r406_c55 bl[55] br[55] wl[406] vdd gnd cell_6t
Xbit_r407_c55 bl[55] br[55] wl[407] vdd gnd cell_6t
Xbit_r408_c55 bl[55] br[55] wl[408] vdd gnd cell_6t
Xbit_r409_c55 bl[55] br[55] wl[409] vdd gnd cell_6t
Xbit_r410_c55 bl[55] br[55] wl[410] vdd gnd cell_6t
Xbit_r411_c55 bl[55] br[55] wl[411] vdd gnd cell_6t
Xbit_r412_c55 bl[55] br[55] wl[412] vdd gnd cell_6t
Xbit_r413_c55 bl[55] br[55] wl[413] vdd gnd cell_6t
Xbit_r414_c55 bl[55] br[55] wl[414] vdd gnd cell_6t
Xbit_r415_c55 bl[55] br[55] wl[415] vdd gnd cell_6t
Xbit_r416_c55 bl[55] br[55] wl[416] vdd gnd cell_6t
Xbit_r417_c55 bl[55] br[55] wl[417] vdd gnd cell_6t
Xbit_r418_c55 bl[55] br[55] wl[418] vdd gnd cell_6t
Xbit_r419_c55 bl[55] br[55] wl[419] vdd gnd cell_6t
Xbit_r420_c55 bl[55] br[55] wl[420] vdd gnd cell_6t
Xbit_r421_c55 bl[55] br[55] wl[421] vdd gnd cell_6t
Xbit_r422_c55 bl[55] br[55] wl[422] vdd gnd cell_6t
Xbit_r423_c55 bl[55] br[55] wl[423] vdd gnd cell_6t
Xbit_r424_c55 bl[55] br[55] wl[424] vdd gnd cell_6t
Xbit_r425_c55 bl[55] br[55] wl[425] vdd gnd cell_6t
Xbit_r426_c55 bl[55] br[55] wl[426] vdd gnd cell_6t
Xbit_r427_c55 bl[55] br[55] wl[427] vdd gnd cell_6t
Xbit_r428_c55 bl[55] br[55] wl[428] vdd gnd cell_6t
Xbit_r429_c55 bl[55] br[55] wl[429] vdd gnd cell_6t
Xbit_r430_c55 bl[55] br[55] wl[430] vdd gnd cell_6t
Xbit_r431_c55 bl[55] br[55] wl[431] vdd gnd cell_6t
Xbit_r432_c55 bl[55] br[55] wl[432] vdd gnd cell_6t
Xbit_r433_c55 bl[55] br[55] wl[433] vdd gnd cell_6t
Xbit_r434_c55 bl[55] br[55] wl[434] vdd gnd cell_6t
Xbit_r435_c55 bl[55] br[55] wl[435] vdd gnd cell_6t
Xbit_r436_c55 bl[55] br[55] wl[436] vdd gnd cell_6t
Xbit_r437_c55 bl[55] br[55] wl[437] vdd gnd cell_6t
Xbit_r438_c55 bl[55] br[55] wl[438] vdd gnd cell_6t
Xbit_r439_c55 bl[55] br[55] wl[439] vdd gnd cell_6t
Xbit_r440_c55 bl[55] br[55] wl[440] vdd gnd cell_6t
Xbit_r441_c55 bl[55] br[55] wl[441] vdd gnd cell_6t
Xbit_r442_c55 bl[55] br[55] wl[442] vdd gnd cell_6t
Xbit_r443_c55 bl[55] br[55] wl[443] vdd gnd cell_6t
Xbit_r444_c55 bl[55] br[55] wl[444] vdd gnd cell_6t
Xbit_r445_c55 bl[55] br[55] wl[445] vdd gnd cell_6t
Xbit_r446_c55 bl[55] br[55] wl[446] vdd gnd cell_6t
Xbit_r447_c55 bl[55] br[55] wl[447] vdd gnd cell_6t
Xbit_r448_c55 bl[55] br[55] wl[448] vdd gnd cell_6t
Xbit_r449_c55 bl[55] br[55] wl[449] vdd gnd cell_6t
Xbit_r450_c55 bl[55] br[55] wl[450] vdd gnd cell_6t
Xbit_r451_c55 bl[55] br[55] wl[451] vdd gnd cell_6t
Xbit_r452_c55 bl[55] br[55] wl[452] vdd gnd cell_6t
Xbit_r453_c55 bl[55] br[55] wl[453] vdd gnd cell_6t
Xbit_r454_c55 bl[55] br[55] wl[454] vdd gnd cell_6t
Xbit_r455_c55 bl[55] br[55] wl[455] vdd gnd cell_6t
Xbit_r456_c55 bl[55] br[55] wl[456] vdd gnd cell_6t
Xbit_r457_c55 bl[55] br[55] wl[457] vdd gnd cell_6t
Xbit_r458_c55 bl[55] br[55] wl[458] vdd gnd cell_6t
Xbit_r459_c55 bl[55] br[55] wl[459] vdd gnd cell_6t
Xbit_r460_c55 bl[55] br[55] wl[460] vdd gnd cell_6t
Xbit_r461_c55 bl[55] br[55] wl[461] vdd gnd cell_6t
Xbit_r462_c55 bl[55] br[55] wl[462] vdd gnd cell_6t
Xbit_r463_c55 bl[55] br[55] wl[463] vdd gnd cell_6t
Xbit_r464_c55 bl[55] br[55] wl[464] vdd gnd cell_6t
Xbit_r465_c55 bl[55] br[55] wl[465] vdd gnd cell_6t
Xbit_r466_c55 bl[55] br[55] wl[466] vdd gnd cell_6t
Xbit_r467_c55 bl[55] br[55] wl[467] vdd gnd cell_6t
Xbit_r468_c55 bl[55] br[55] wl[468] vdd gnd cell_6t
Xbit_r469_c55 bl[55] br[55] wl[469] vdd gnd cell_6t
Xbit_r470_c55 bl[55] br[55] wl[470] vdd gnd cell_6t
Xbit_r471_c55 bl[55] br[55] wl[471] vdd gnd cell_6t
Xbit_r472_c55 bl[55] br[55] wl[472] vdd gnd cell_6t
Xbit_r473_c55 bl[55] br[55] wl[473] vdd gnd cell_6t
Xbit_r474_c55 bl[55] br[55] wl[474] vdd gnd cell_6t
Xbit_r475_c55 bl[55] br[55] wl[475] vdd gnd cell_6t
Xbit_r476_c55 bl[55] br[55] wl[476] vdd gnd cell_6t
Xbit_r477_c55 bl[55] br[55] wl[477] vdd gnd cell_6t
Xbit_r478_c55 bl[55] br[55] wl[478] vdd gnd cell_6t
Xbit_r479_c55 bl[55] br[55] wl[479] vdd gnd cell_6t
Xbit_r480_c55 bl[55] br[55] wl[480] vdd gnd cell_6t
Xbit_r481_c55 bl[55] br[55] wl[481] vdd gnd cell_6t
Xbit_r482_c55 bl[55] br[55] wl[482] vdd gnd cell_6t
Xbit_r483_c55 bl[55] br[55] wl[483] vdd gnd cell_6t
Xbit_r484_c55 bl[55] br[55] wl[484] vdd gnd cell_6t
Xbit_r485_c55 bl[55] br[55] wl[485] vdd gnd cell_6t
Xbit_r486_c55 bl[55] br[55] wl[486] vdd gnd cell_6t
Xbit_r487_c55 bl[55] br[55] wl[487] vdd gnd cell_6t
Xbit_r488_c55 bl[55] br[55] wl[488] vdd gnd cell_6t
Xbit_r489_c55 bl[55] br[55] wl[489] vdd gnd cell_6t
Xbit_r490_c55 bl[55] br[55] wl[490] vdd gnd cell_6t
Xbit_r491_c55 bl[55] br[55] wl[491] vdd gnd cell_6t
Xbit_r492_c55 bl[55] br[55] wl[492] vdd gnd cell_6t
Xbit_r493_c55 bl[55] br[55] wl[493] vdd gnd cell_6t
Xbit_r494_c55 bl[55] br[55] wl[494] vdd gnd cell_6t
Xbit_r495_c55 bl[55] br[55] wl[495] vdd gnd cell_6t
Xbit_r496_c55 bl[55] br[55] wl[496] vdd gnd cell_6t
Xbit_r497_c55 bl[55] br[55] wl[497] vdd gnd cell_6t
Xbit_r498_c55 bl[55] br[55] wl[498] vdd gnd cell_6t
Xbit_r499_c55 bl[55] br[55] wl[499] vdd gnd cell_6t
Xbit_r500_c55 bl[55] br[55] wl[500] vdd gnd cell_6t
Xbit_r501_c55 bl[55] br[55] wl[501] vdd gnd cell_6t
Xbit_r502_c55 bl[55] br[55] wl[502] vdd gnd cell_6t
Xbit_r503_c55 bl[55] br[55] wl[503] vdd gnd cell_6t
Xbit_r504_c55 bl[55] br[55] wl[504] vdd gnd cell_6t
Xbit_r505_c55 bl[55] br[55] wl[505] vdd gnd cell_6t
Xbit_r506_c55 bl[55] br[55] wl[506] vdd gnd cell_6t
Xbit_r507_c55 bl[55] br[55] wl[507] vdd gnd cell_6t
Xbit_r508_c55 bl[55] br[55] wl[508] vdd gnd cell_6t
Xbit_r509_c55 bl[55] br[55] wl[509] vdd gnd cell_6t
Xbit_r510_c55 bl[55] br[55] wl[510] vdd gnd cell_6t
Xbit_r511_c55 bl[55] br[55] wl[511] vdd gnd cell_6t
Xbit_r0_c56 bl[56] br[56] wl[0] vdd gnd cell_6t
Xbit_r1_c56 bl[56] br[56] wl[1] vdd gnd cell_6t
Xbit_r2_c56 bl[56] br[56] wl[2] vdd gnd cell_6t
Xbit_r3_c56 bl[56] br[56] wl[3] vdd gnd cell_6t
Xbit_r4_c56 bl[56] br[56] wl[4] vdd gnd cell_6t
Xbit_r5_c56 bl[56] br[56] wl[5] vdd gnd cell_6t
Xbit_r6_c56 bl[56] br[56] wl[6] vdd gnd cell_6t
Xbit_r7_c56 bl[56] br[56] wl[7] vdd gnd cell_6t
Xbit_r8_c56 bl[56] br[56] wl[8] vdd gnd cell_6t
Xbit_r9_c56 bl[56] br[56] wl[9] vdd gnd cell_6t
Xbit_r10_c56 bl[56] br[56] wl[10] vdd gnd cell_6t
Xbit_r11_c56 bl[56] br[56] wl[11] vdd gnd cell_6t
Xbit_r12_c56 bl[56] br[56] wl[12] vdd gnd cell_6t
Xbit_r13_c56 bl[56] br[56] wl[13] vdd gnd cell_6t
Xbit_r14_c56 bl[56] br[56] wl[14] vdd gnd cell_6t
Xbit_r15_c56 bl[56] br[56] wl[15] vdd gnd cell_6t
Xbit_r16_c56 bl[56] br[56] wl[16] vdd gnd cell_6t
Xbit_r17_c56 bl[56] br[56] wl[17] vdd gnd cell_6t
Xbit_r18_c56 bl[56] br[56] wl[18] vdd gnd cell_6t
Xbit_r19_c56 bl[56] br[56] wl[19] vdd gnd cell_6t
Xbit_r20_c56 bl[56] br[56] wl[20] vdd gnd cell_6t
Xbit_r21_c56 bl[56] br[56] wl[21] vdd gnd cell_6t
Xbit_r22_c56 bl[56] br[56] wl[22] vdd gnd cell_6t
Xbit_r23_c56 bl[56] br[56] wl[23] vdd gnd cell_6t
Xbit_r24_c56 bl[56] br[56] wl[24] vdd gnd cell_6t
Xbit_r25_c56 bl[56] br[56] wl[25] vdd gnd cell_6t
Xbit_r26_c56 bl[56] br[56] wl[26] vdd gnd cell_6t
Xbit_r27_c56 bl[56] br[56] wl[27] vdd gnd cell_6t
Xbit_r28_c56 bl[56] br[56] wl[28] vdd gnd cell_6t
Xbit_r29_c56 bl[56] br[56] wl[29] vdd gnd cell_6t
Xbit_r30_c56 bl[56] br[56] wl[30] vdd gnd cell_6t
Xbit_r31_c56 bl[56] br[56] wl[31] vdd gnd cell_6t
Xbit_r32_c56 bl[56] br[56] wl[32] vdd gnd cell_6t
Xbit_r33_c56 bl[56] br[56] wl[33] vdd gnd cell_6t
Xbit_r34_c56 bl[56] br[56] wl[34] vdd gnd cell_6t
Xbit_r35_c56 bl[56] br[56] wl[35] vdd gnd cell_6t
Xbit_r36_c56 bl[56] br[56] wl[36] vdd gnd cell_6t
Xbit_r37_c56 bl[56] br[56] wl[37] vdd gnd cell_6t
Xbit_r38_c56 bl[56] br[56] wl[38] vdd gnd cell_6t
Xbit_r39_c56 bl[56] br[56] wl[39] vdd gnd cell_6t
Xbit_r40_c56 bl[56] br[56] wl[40] vdd gnd cell_6t
Xbit_r41_c56 bl[56] br[56] wl[41] vdd gnd cell_6t
Xbit_r42_c56 bl[56] br[56] wl[42] vdd gnd cell_6t
Xbit_r43_c56 bl[56] br[56] wl[43] vdd gnd cell_6t
Xbit_r44_c56 bl[56] br[56] wl[44] vdd gnd cell_6t
Xbit_r45_c56 bl[56] br[56] wl[45] vdd gnd cell_6t
Xbit_r46_c56 bl[56] br[56] wl[46] vdd gnd cell_6t
Xbit_r47_c56 bl[56] br[56] wl[47] vdd gnd cell_6t
Xbit_r48_c56 bl[56] br[56] wl[48] vdd gnd cell_6t
Xbit_r49_c56 bl[56] br[56] wl[49] vdd gnd cell_6t
Xbit_r50_c56 bl[56] br[56] wl[50] vdd gnd cell_6t
Xbit_r51_c56 bl[56] br[56] wl[51] vdd gnd cell_6t
Xbit_r52_c56 bl[56] br[56] wl[52] vdd gnd cell_6t
Xbit_r53_c56 bl[56] br[56] wl[53] vdd gnd cell_6t
Xbit_r54_c56 bl[56] br[56] wl[54] vdd gnd cell_6t
Xbit_r55_c56 bl[56] br[56] wl[55] vdd gnd cell_6t
Xbit_r56_c56 bl[56] br[56] wl[56] vdd gnd cell_6t
Xbit_r57_c56 bl[56] br[56] wl[57] vdd gnd cell_6t
Xbit_r58_c56 bl[56] br[56] wl[58] vdd gnd cell_6t
Xbit_r59_c56 bl[56] br[56] wl[59] vdd gnd cell_6t
Xbit_r60_c56 bl[56] br[56] wl[60] vdd gnd cell_6t
Xbit_r61_c56 bl[56] br[56] wl[61] vdd gnd cell_6t
Xbit_r62_c56 bl[56] br[56] wl[62] vdd gnd cell_6t
Xbit_r63_c56 bl[56] br[56] wl[63] vdd gnd cell_6t
Xbit_r64_c56 bl[56] br[56] wl[64] vdd gnd cell_6t
Xbit_r65_c56 bl[56] br[56] wl[65] vdd gnd cell_6t
Xbit_r66_c56 bl[56] br[56] wl[66] vdd gnd cell_6t
Xbit_r67_c56 bl[56] br[56] wl[67] vdd gnd cell_6t
Xbit_r68_c56 bl[56] br[56] wl[68] vdd gnd cell_6t
Xbit_r69_c56 bl[56] br[56] wl[69] vdd gnd cell_6t
Xbit_r70_c56 bl[56] br[56] wl[70] vdd gnd cell_6t
Xbit_r71_c56 bl[56] br[56] wl[71] vdd gnd cell_6t
Xbit_r72_c56 bl[56] br[56] wl[72] vdd gnd cell_6t
Xbit_r73_c56 bl[56] br[56] wl[73] vdd gnd cell_6t
Xbit_r74_c56 bl[56] br[56] wl[74] vdd gnd cell_6t
Xbit_r75_c56 bl[56] br[56] wl[75] vdd gnd cell_6t
Xbit_r76_c56 bl[56] br[56] wl[76] vdd gnd cell_6t
Xbit_r77_c56 bl[56] br[56] wl[77] vdd gnd cell_6t
Xbit_r78_c56 bl[56] br[56] wl[78] vdd gnd cell_6t
Xbit_r79_c56 bl[56] br[56] wl[79] vdd gnd cell_6t
Xbit_r80_c56 bl[56] br[56] wl[80] vdd gnd cell_6t
Xbit_r81_c56 bl[56] br[56] wl[81] vdd gnd cell_6t
Xbit_r82_c56 bl[56] br[56] wl[82] vdd gnd cell_6t
Xbit_r83_c56 bl[56] br[56] wl[83] vdd gnd cell_6t
Xbit_r84_c56 bl[56] br[56] wl[84] vdd gnd cell_6t
Xbit_r85_c56 bl[56] br[56] wl[85] vdd gnd cell_6t
Xbit_r86_c56 bl[56] br[56] wl[86] vdd gnd cell_6t
Xbit_r87_c56 bl[56] br[56] wl[87] vdd gnd cell_6t
Xbit_r88_c56 bl[56] br[56] wl[88] vdd gnd cell_6t
Xbit_r89_c56 bl[56] br[56] wl[89] vdd gnd cell_6t
Xbit_r90_c56 bl[56] br[56] wl[90] vdd gnd cell_6t
Xbit_r91_c56 bl[56] br[56] wl[91] vdd gnd cell_6t
Xbit_r92_c56 bl[56] br[56] wl[92] vdd gnd cell_6t
Xbit_r93_c56 bl[56] br[56] wl[93] vdd gnd cell_6t
Xbit_r94_c56 bl[56] br[56] wl[94] vdd gnd cell_6t
Xbit_r95_c56 bl[56] br[56] wl[95] vdd gnd cell_6t
Xbit_r96_c56 bl[56] br[56] wl[96] vdd gnd cell_6t
Xbit_r97_c56 bl[56] br[56] wl[97] vdd gnd cell_6t
Xbit_r98_c56 bl[56] br[56] wl[98] vdd gnd cell_6t
Xbit_r99_c56 bl[56] br[56] wl[99] vdd gnd cell_6t
Xbit_r100_c56 bl[56] br[56] wl[100] vdd gnd cell_6t
Xbit_r101_c56 bl[56] br[56] wl[101] vdd gnd cell_6t
Xbit_r102_c56 bl[56] br[56] wl[102] vdd gnd cell_6t
Xbit_r103_c56 bl[56] br[56] wl[103] vdd gnd cell_6t
Xbit_r104_c56 bl[56] br[56] wl[104] vdd gnd cell_6t
Xbit_r105_c56 bl[56] br[56] wl[105] vdd gnd cell_6t
Xbit_r106_c56 bl[56] br[56] wl[106] vdd gnd cell_6t
Xbit_r107_c56 bl[56] br[56] wl[107] vdd gnd cell_6t
Xbit_r108_c56 bl[56] br[56] wl[108] vdd gnd cell_6t
Xbit_r109_c56 bl[56] br[56] wl[109] vdd gnd cell_6t
Xbit_r110_c56 bl[56] br[56] wl[110] vdd gnd cell_6t
Xbit_r111_c56 bl[56] br[56] wl[111] vdd gnd cell_6t
Xbit_r112_c56 bl[56] br[56] wl[112] vdd gnd cell_6t
Xbit_r113_c56 bl[56] br[56] wl[113] vdd gnd cell_6t
Xbit_r114_c56 bl[56] br[56] wl[114] vdd gnd cell_6t
Xbit_r115_c56 bl[56] br[56] wl[115] vdd gnd cell_6t
Xbit_r116_c56 bl[56] br[56] wl[116] vdd gnd cell_6t
Xbit_r117_c56 bl[56] br[56] wl[117] vdd gnd cell_6t
Xbit_r118_c56 bl[56] br[56] wl[118] vdd gnd cell_6t
Xbit_r119_c56 bl[56] br[56] wl[119] vdd gnd cell_6t
Xbit_r120_c56 bl[56] br[56] wl[120] vdd gnd cell_6t
Xbit_r121_c56 bl[56] br[56] wl[121] vdd gnd cell_6t
Xbit_r122_c56 bl[56] br[56] wl[122] vdd gnd cell_6t
Xbit_r123_c56 bl[56] br[56] wl[123] vdd gnd cell_6t
Xbit_r124_c56 bl[56] br[56] wl[124] vdd gnd cell_6t
Xbit_r125_c56 bl[56] br[56] wl[125] vdd gnd cell_6t
Xbit_r126_c56 bl[56] br[56] wl[126] vdd gnd cell_6t
Xbit_r127_c56 bl[56] br[56] wl[127] vdd gnd cell_6t
Xbit_r128_c56 bl[56] br[56] wl[128] vdd gnd cell_6t
Xbit_r129_c56 bl[56] br[56] wl[129] vdd gnd cell_6t
Xbit_r130_c56 bl[56] br[56] wl[130] vdd gnd cell_6t
Xbit_r131_c56 bl[56] br[56] wl[131] vdd gnd cell_6t
Xbit_r132_c56 bl[56] br[56] wl[132] vdd gnd cell_6t
Xbit_r133_c56 bl[56] br[56] wl[133] vdd gnd cell_6t
Xbit_r134_c56 bl[56] br[56] wl[134] vdd gnd cell_6t
Xbit_r135_c56 bl[56] br[56] wl[135] vdd gnd cell_6t
Xbit_r136_c56 bl[56] br[56] wl[136] vdd gnd cell_6t
Xbit_r137_c56 bl[56] br[56] wl[137] vdd gnd cell_6t
Xbit_r138_c56 bl[56] br[56] wl[138] vdd gnd cell_6t
Xbit_r139_c56 bl[56] br[56] wl[139] vdd gnd cell_6t
Xbit_r140_c56 bl[56] br[56] wl[140] vdd gnd cell_6t
Xbit_r141_c56 bl[56] br[56] wl[141] vdd gnd cell_6t
Xbit_r142_c56 bl[56] br[56] wl[142] vdd gnd cell_6t
Xbit_r143_c56 bl[56] br[56] wl[143] vdd gnd cell_6t
Xbit_r144_c56 bl[56] br[56] wl[144] vdd gnd cell_6t
Xbit_r145_c56 bl[56] br[56] wl[145] vdd gnd cell_6t
Xbit_r146_c56 bl[56] br[56] wl[146] vdd gnd cell_6t
Xbit_r147_c56 bl[56] br[56] wl[147] vdd gnd cell_6t
Xbit_r148_c56 bl[56] br[56] wl[148] vdd gnd cell_6t
Xbit_r149_c56 bl[56] br[56] wl[149] vdd gnd cell_6t
Xbit_r150_c56 bl[56] br[56] wl[150] vdd gnd cell_6t
Xbit_r151_c56 bl[56] br[56] wl[151] vdd gnd cell_6t
Xbit_r152_c56 bl[56] br[56] wl[152] vdd gnd cell_6t
Xbit_r153_c56 bl[56] br[56] wl[153] vdd gnd cell_6t
Xbit_r154_c56 bl[56] br[56] wl[154] vdd gnd cell_6t
Xbit_r155_c56 bl[56] br[56] wl[155] vdd gnd cell_6t
Xbit_r156_c56 bl[56] br[56] wl[156] vdd gnd cell_6t
Xbit_r157_c56 bl[56] br[56] wl[157] vdd gnd cell_6t
Xbit_r158_c56 bl[56] br[56] wl[158] vdd gnd cell_6t
Xbit_r159_c56 bl[56] br[56] wl[159] vdd gnd cell_6t
Xbit_r160_c56 bl[56] br[56] wl[160] vdd gnd cell_6t
Xbit_r161_c56 bl[56] br[56] wl[161] vdd gnd cell_6t
Xbit_r162_c56 bl[56] br[56] wl[162] vdd gnd cell_6t
Xbit_r163_c56 bl[56] br[56] wl[163] vdd gnd cell_6t
Xbit_r164_c56 bl[56] br[56] wl[164] vdd gnd cell_6t
Xbit_r165_c56 bl[56] br[56] wl[165] vdd gnd cell_6t
Xbit_r166_c56 bl[56] br[56] wl[166] vdd gnd cell_6t
Xbit_r167_c56 bl[56] br[56] wl[167] vdd gnd cell_6t
Xbit_r168_c56 bl[56] br[56] wl[168] vdd gnd cell_6t
Xbit_r169_c56 bl[56] br[56] wl[169] vdd gnd cell_6t
Xbit_r170_c56 bl[56] br[56] wl[170] vdd gnd cell_6t
Xbit_r171_c56 bl[56] br[56] wl[171] vdd gnd cell_6t
Xbit_r172_c56 bl[56] br[56] wl[172] vdd gnd cell_6t
Xbit_r173_c56 bl[56] br[56] wl[173] vdd gnd cell_6t
Xbit_r174_c56 bl[56] br[56] wl[174] vdd gnd cell_6t
Xbit_r175_c56 bl[56] br[56] wl[175] vdd gnd cell_6t
Xbit_r176_c56 bl[56] br[56] wl[176] vdd gnd cell_6t
Xbit_r177_c56 bl[56] br[56] wl[177] vdd gnd cell_6t
Xbit_r178_c56 bl[56] br[56] wl[178] vdd gnd cell_6t
Xbit_r179_c56 bl[56] br[56] wl[179] vdd gnd cell_6t
Xbit_r180_c56 bl[56] br[56] wl[180] vdd gnd cell_6t
Xbit_r181_c56 bl[56] br[56] wl[181] vdd gnd cell_6t
Xbit_r182_c56 bl[56] br[56] wl[182] vdd gnd cell_6t
Xbit_r183_c56 bl[56] br[56] wl[183] vdd gnd cell_6t
Xbit_r184_c56 bl[56] br[56] wl[184] vdd gnd cell_6t
Xbit_r185_c56 bl[56] br[56] wl[185] vdd gnd cell_6t
Xbit_r186_c56 bl[56] br[56] wl[186] vdd gnd cell_6t
Xbit_r187_c56 bl[56] br[56] wl[187] vdd gnd cell_6t
Xbit_r188_c56 bl[56] br[56] wl[188] vdd gnd cell_6t
Xbit_r189_c56 bl[56] br[56] wl[189] vdd gnd cell_6t
Xbit_r190_c56 bl[56] br[56] wl[190] vdd gnd cell_6t
Xbit_r191_c56 bl[56] br[56] wl[191] vdd gnd cell_6t
Xbit_r192_c56 bl[56] br[56] wl[192] vdd gnd cell_6t
Xbit_r193_c56 bl[56] br[56] wl[193] vdd gnd cell_6t
Xbit_r194_c56 bl[56] br[56] wl[194] vdd gnd cell_6t
Xbit_r195_c56 bl[56] br[56] wl[195] vdd gnd cell_6t
Xbit_r196_c56 bl[56] br[56] wl[196] vdd gnd cell_6t
Xbit_r197_c56 bl[56] br[56] wl[197] vdd gnd cell_6t
Xbit_r198_c56 bl[56] br[56] wl[198] vdd gnd cell_6t
Xbit_r199_c56 bl[56] br[56] wl[199] vdd gnd cell_6t
Xbit_r200_c56 bl[56] br[56] wl[200] vdd gnd cell_6t
Xbit_r201_c56 bl[56] br[56] wl[201] vdd gnd cell_6t
Xbit_r202_c56 bl[56] br[56] wl[202] vdd gnd cell_6t
Xbit_r203_c56 bl[56] br[56] wl[203] vdd gnd cell_6t
Xbit_r204_c56 bl[56] br[56] wl[204] vdd gnd cell_6t
Xbit_r205_c56 bl[56] br[56] wl[205] vdd gnd cell_6t
Xbit_r206_c56 bl[56] br[56] wl[206] vdd gnd cell_6t
Xbit_r207_c56 bl[56] br[56] wl[207] vdd gnd cell_6t
Xbit_r208_c56 bl[56] br[56] wl[208] vdd gnd cell_6t
Xbit_r209_c56 bl[56] br[56] wl[209] vdd gnd cell_6t
Xbit_r210_c56 bl[56] br[56] wl[210] vdd gnd cell_6t
Xbit_r211_c56 bl[56] br[56] wl[211] vdd gnd cell_6t
Xbit_r212_c56 bl[56] br[56] wl[212] vdd gnd cell_6t
Xbit_r213_c56 bl[56] br[56] wl[213] vdd gnd cell_6t
Xbit_r214_c56 bl[56] br[56] wl[214] vdd gnd cell_6t
Xbit_r215_c56 bl[56] br[56] wl[215] vdd gnd cell_6t
Xbit_r216_c56 bl[56] br[56] wl[216] vdd gnd cell_6t
Xbit_r217_c56 bl[56] br[56] wl[217] vdd gnd cell_6t
Xbit_r218_c56 bl[56] br[56] wl[218] vdd gnd cell_6t
Xbit_r219_c56 bl[56] br[56] wl[219] vdd gnd cell_6t
Xbit_r220_c56 bl[56] br[56] wl[220] vdd gnd cell_6t
Xbit_r221_c56 bl[56] br[56] wl[221] vdd gnd cell_6t
Xbit_r222_c56 bl[56] br[56] wl[222] vdd gnd cell_6t
Xbit_r223_c56 bl[56] br[56] wl[223] vdd gnd cell_6t
Xbit_r224_c56 bl[56] br[56] wl[224] vdd gnd cell_6t
Xbit_r225_c56 bl[56] br[56] wl[225] vdd gnd cell_6t
Xbit_r226_c56 bl[56] br[56] wl[226] vdd gnd cell_6t
Xbit_r227_c56 bl[56] br[56] wl[227] vdd gnd cell_6t
Xbit_r228_c56 bl[56] br[56] wl[228] vdd gnd cell_6t
Xbit_r229_c56 bl[56] br[56] wl[229] vdd gnd cell_6t
Xbit_r230_c56 bl[56] br[56] wl[230] vdd gnd cell_6t
Xbit_r231_c56 bl[56] br[56] wl[231] vdd gnd cell_6t
Xbit_r232_c56 bl[56] br[56] wl[232] vdd gnd cell_6t
Xbit_r233_c56 bl[56] br[56] wl[233] vdd gnd cell_6t
Xbit_r234_c56 bl[56] br[56] wl[234] vdd gnd cell_6t
Xbit_r235_c56 bl[56] br[56] wl[235] vdd gnd cell_6t
Xbit_r236_c56 bl[56] br[56] wl[236] vdd gnd cell_6t
Xbit_r237_c56 bl[56] br[56] wl[237] vdd gnd cell_6t
Xbit_r238_c56 bl[56] br[56] wl[238] vdd gnd cell_6t
Xbit_r239_c56 bl[56] br[56] wl[239] vdd gnd cell_6t
Xbit_r240_c56 bl[56] br[56] wl[240] vdd gnd cell_6t
Xbit_r241_c56 bl[56] br[56] wl[241] vdd gnd cell_6t
Xbit_r242_c56 bl[56] br[56] wl[242] vdd gnd cell_6t
Xbit_r243_c56 bl[56] br[56] wl[243] vdd gnd cell_6t
Xbit_r244_c56 bl[56] br[56] wl[244] vdd gnd cell_6t
Xbit_r245_c56 bl[56] br[56] wl[245] vdd gnd cell_6t
Xbit_r246_c56 bl[56] br[56] wl[246] vdd gnd cell_6t
Xbit_r247_c56 bl[56] br[56] wl[247] vdd gnd cell_6t
Xbit_r248_c56 bl[56] br[56] wl[248] vdd gnd cell_6t
Xbit_r249_c56 bl[56] br[56] wl[249] vdd gnd cell_6t
Xbit_r250_c56 bl[56] br[56] wl[250] vdd gnd cell_6t
Xbit_r251_c56 bl[56] br[56] wl[251] vdd gnd cell_6t
Xbit_r252_c56 bl[56] br[56] wl[252] vdd gnd cell_6t
Xbit_r253_c56 bl[56] br[56] wl[253] vdd gnd cell_6t
Xbit_r254_c56 bl[56] br[56] wl[254] vdd gnd cell_6t
Xbit_r255_c56 bl[56] br[56] wl[255] vdd gnd cell_6t
Xbit_r256_c56 bl[56] br[56] wl[256] vdd gnd cell_6t
Xbit_r257_c56 bl[56] br[56] wl[257] vdd gnd cell_6t
Xbit_r258_c56 bl[56] br[56] wl[258] vdd gnd cell_6t
Xbit_r259_c56 bl[56] br[56] wl[259] vdd gnd cell_6t
Xbit_r260_c56 bl[56] br[56] wl[260] vdd gnd cell_6t
Xbit_r261_c56 bl[56] br[56] wl[261] vdd gnd cell_6t
Xbit_r262_c56 bl[56] br[56] wl[262] vdd gnd cell_6t
Xbit_r263_c56 bl[56] br[56] wl[263] vdd gnd cell_6t
Xbit_r264_c56 bl[56] br[56] wl[264] vdd gnd cell_6t
Xbit_r265_c56 bl[56] br[56] wl[265] vdd gnd cell_6t
Xbit_r266_c56 bl[56] br[56] wl[266] vdd gnd cell_6t
Xbit_r267_c56 bl[56] br[56] wl[267] vdd gnd cell_6t
Xbit_r268_c56 bl[56] br[56] wl[268] vdd gnd cell_6t
Xbit_r269_c56 bl[56] br[56] wl[269] vdd gnd cell_6t
Xbit_r270_c56 bl[56] br[56] wl[270] vdd gnd cell_6t
Xbit_r271_c56 bl[56] br[56] wl[271] vdd gnd cell_6t
Xbit_r272_c56 bl[56] br[56] wl[272] vdd gnd cell_6t
Xbit_r273_c56 bl[56] br[56] wl[273] vdd gnd cell_6t
Xbit_r274_c56 bl[56] br[56] wl[274] vdd gnd cell_6t
Xbit_r275_c56 bl[56] br[56] wl[275] vdd gnd cell_6t
Xbit_r276_c56 bl[56] br[56] wl[276] vdd gnd cell_6t
Xbit_r277_c56 bl[56] br[56] wl[277] vdd gnd cell_6t
Xbit_r278_c56 bl[56] br[56] wl[278] vdd gnd cell_6t
Xbit_r279_c56 bl[56] br[56] wl[279] vdd gnd cell_6t
Xbit_r280_c56 bl[56] br[56] wl[280] vdd gnd cell_6t
Xbit_r281_c56 bl[56] br[56] wl[281] vdd gnd cell_6t
Xbit_r282_c56 bl[56] br[56] wl[282] vdd gnd cell_6t
Xbit_r283_c56 bl[56] br[56] wl[283] vdd gnd cell_6t
Xbit_r284_c56 bl[56] br[56] wl[284] vdd gnd cell_6t
Xbit_r285_c56 bl[56] br[56] wl[285] vdd gnd cell_6t
Xbit_r286_c56 bl[56] br[56] wl[286] vdd gnd cell_6t
Xbit_r287_c56 bl[56] br[56] wl[287] vdd gnd cell_6t
Xbit_r288_c56 bl[56] br[56] wl[288] vdd gnd cell_6t
Xbit_r289_c56 bl[56] br[56] wl[289] vdd gnd cell_6t
Xbit_r290_c56 bl[56] br[56] wl[290] vdd gnd cell_6t
Xbit_r291_c56 bl[56] br[56] wl[291] vdd gnd cell_6t
Xbit_r292_c56 bl[56] br[56] wl[292] vdd gnd cell_6t
Xbit_r293_c56 bl[56] br[56] wl[293] vdd gnd cell_6t
Xbit_r294_c56 bl[56] br[56] wl[294] vdd gnd cell_6t
Xbit_r295_c56 bl[56] br[56] wl[295] vdd gnd cell_6t
Xbit_r296_c56 bl[56] br[56] wl[296] vdd gnd cell_6t
Xbit_r297_c56 bl[56] br[56] wl[297] vdd gnd cell_6t
Xbit_r298_c56 bl[56] br[56] wl[298] vdd gnd cell_6t
Xbit_r299_c56 bl[56] br[56] wl[299] vdd gnd cell_6t
Xbit_r300_c56 bl[56] br[56] wl[300] vdd gnd cell_6t
Xbit_r301_c56 bl[56] br[56] wl[301] vdd gnd cell_6t
Xbit_r302_c56 bl[56] br[56] wl[302] vdd gnd cell_6t
Xbit_r303_c56 bl[56] br[56] wl[303] vdd gnd cell_6t
Xbit_r304_c56 bl[56] br[56] wl[304] vdd gnd cell_6t
Xbit_r305_c56 bl[56] br[56] wl[305] vdd gnd cell_6t
Xbit_r306_c56 bl[56] br[56] wl[306] vdd gnd cell_6t
Xbit_r307_c56 bl[56] br[56] wl[307] vdd gnd cell_6t
Xbit_r308_c56 bl[56] br[56] wl[308] vdd gnd cell_6t
Xbit_r309_c56 bl[56] br[56] wl[309] vdd gnd cell_6t
Xbit_r310_c56 bl[56] br[56] wl[310] vdd gnd cell_6t
Xbit_r311_c56 bl[56] br[56] wl[311] vdd gnd cell_6t
Xbit_r312_c56 bl[56] br[56] wl[312] vdd gnd cell_6t
Xbit_r313_c56 bl[56] br[56] wl[313] vdd gnd cell_6t
Xbit_r314_c56 bl[56] br[56] wl[314] vdd gnd cell_6t
Xbit_r315_c56 bl[56] br[56] wl[315] vdd gnd cell_6t
Xbit_r316_c56 bl[56] br[56] wl[316] vdd gnd cell_6t
Xbit_r317_c56 bl[56] br[56] wl[317] vdd gnd cell_6t
Xbit_r318_c56 bl[56] br[56] wl[318] vdd gnd cell_6t
Xbit_r319_c56 bl[56] br[56] wl[319] vdd gnd cell_6t
Xbit_r320_c56 bl[56] br[56] wl[320] vdd gnd cell_6t
Xbit_r321_c56 bl[56] br[56] wl[321] vdd gnd cell_6t
Xbit_r322_c56 bl[56] br[56] wl[322] vdd gnd cell_6t
Xbit_r323_c56 bl[56] br[56] wl[323] vdd gnd cell_6t
Xbit_r324_c56 bl[56] br[56] wl[324] vdd gnd cell_6t
Xbit_r325_c56 bl[56] br[56] wl[325] vdd gnd cell_6t
Xbit_r326_c56 bl[56] br[56] wl[326] vdd gnd cell_6t
Xbit_r327_c56 bl[56] br[56] wl[327] vdd gnd cell_6t
Xbit_r328_c56 bl[56] br[56] wl[328] vdd gnd cell_6t
Xbit_r329_c56 bl[56] br[56] wl[329] vdd gnd cell_6t
Xbit_r330_c56 bl[56] br[56] wl[330] vdd gnd cell_6t
Xbit_r331_c56 bl[56] br[56] wl[331] vdd gnd cell_6t
Xbit_r332_c56 bl[56] br[56] wl[332] vdd gnd cell_6t
Xbit_r333_c56 bl[56] br[56] wl[333] vdd gnd cell_6t
Xbit_r334_c56 bl[56] br[56] wl[334] vdd gnd cell_6t
Xbit_r335_c56 bl[56] br[56] wl[335] vdd gnd cell_6t
Xbit_r336_c56 bl[56] br[56] wl[336] vdd gnd cell_6t
Xbit_r337_c56 bl[56] br[56] wl[337] vdd gnd cell_6t
Xbit_r338_c56 bl[56] br[56] wl[338] vdd gnd cell_6t
Xbit_r339_c56 bl[56] br[56] wl[339] vdd gnd cell_6t
Xbit_r340_c56 bl[56] br[56] wl[340] vdd gnd cell_6t
Xbit_r341_c56 bl[56] br[56] wl[341] vdd gnd cell_6t
Xbit_r342_c56 bl[56] br[56] wl[342] vdd gnd cell_6t
Xbit_r343_c56 bl[56] br[56] wl[343] vdd gnd cell_6t
Xbit_r344_c56 bl[56] br[56] wl[344] vdd gnd cell_6t
Xbit_r345_c56 bl[56] br[56] wl[345] vdd gnd cell_6t
Xbit_r346_c56 bl[56] br[56] wl[346] vdd gnd cell_6t
Xbit_r347_c56 bl[56] br[56] wl[347] vdd gnd cell_6t
Xbit_r348_c56 bl[56] br[56] wl[348] vdd gnd cell_6t
Xbit_r349_c56 bl[56] br[56] wl[349] vdd gnd cell_6t
Xbit_r350_c56 bl[56] br[56] wl[350] vdd gnd cell_6t
Xbit_r351_c56 bl[56] br[56] wl[351] vdd gnd cell_6t
Xbit_r352_c56 bl[56] br[56] wl[352] vdd gnd cell_6t
Xbit_r353_c56 bl[56] br[56] wl[353] vdd gnd cell_6t
Xbit_r354_c56 bl[56] br[56] wl[354] vdd gnd cell_6t
Xbit_r355_c56 bl[56] br[56] wl[355] vdd gnd cell_6t
Xbit_r356_c56 bl[56] br[56] wl[356] vdd gnd cell_6t
Xbit_r357_c56 bl[56] br[56] wl[357] vdd gnd cell_6t
Xbit_r358_c56 bl[56] br[56] wl[358] vdd gnd cell_6t
Xbit_r359_c56 bl[56] br[56] wl[359] vdd gnd cell_6t
Xbit_r360_c56 bl[56] br[56] wl[360] vdd gnd cell_6t
Xbit_r361_c56 bl[56] br[56] wl[361] vdd gnd cell_6t
Xbit_r362_c56 bl[56] br[56] wl[362] vdd gnd cell_6t
Xbit_r363_c56 bl[56] br[56] wl[363] vdd gnd cell_6t
Xbit_r364_c56 bl[56] br[56] wl[364] vdd gnd cell_6t
Xbit_r365_c56 bl[56] br[56] wl[365] vdd gnd cell_6t
Xbit_r366_c56 bl[56] br[56] wl[366] vdd gnd cell_6t
Xbit_r367_c56 bl[56] br[56] wl[367] vdd gnd cell_6t
Xbit_r368_c56 bl[56] br[56] wl[368] vdd gnd cell_6t
Xbit_r369_c56 bl[56] br[56] wl[369] vdd gnd cell_6t
Xbit_r370_c56 bl[56] br[56] wl[370] vdd gnd cell_6t
Xbit_r371_c56 bl[56] br[56] wl[371] vdd gnd cell_6t
Xbit_r372_c56 bl[56] br[56] wl[372] vdd gnd cell_6t
Xbit_r373_c56 bl[56] br[56] wl[373] vdd gnd cell_6t
Xbit_r374_c56 bl[56] br[56] wl[374] vdd gnd cell_6t
Xbit_r375_c56 bl[56] br[56] wl[375] vdd gnd cell_6t
Xbit_r376_c56 bl[56] br[56] wl[376] vdd gnd cell_6t
Xbit_r377_c56 bl[56] br[56] wl[377] vdd gnd cell_6t
Xbit_r378_c56 bl[56] br[56] wl[378] vdd gnd cell_6t
Xbit_r379_c56 bl[56] br[56] wl[379] vdd gnd cell_6t
Xbit_r380_c56 bl[56] br[56] wl[380] vdd gnd cell_6t
Xbit_r381_c56 bl[56] br[56] wl[381] vdd gnd cell_6t
Xbit_r382_c56 bl[56] br[56] wl[382] vdd gnd cell_6t
Xbit_r383_c56 bl[56] br[56] wl[383] vdd gnd cell_6t
Xbit_r384_c56 bl[56] br[56] wl[384] vdd gnd cell_6t
Xbit_r385_c56 bl[56] br[56] wl[385] vdd gnd cell_6t
Xbit_r386_c56 bl[56] br[56] wl[386] vdd gnd cell_6t
Xbit_r387_c56 bl[56] br[56] wl[387] vdd gnd cell_6t
Xbit_r388_c56 bl[56] br[56] wl[388] vdd gnd cell_6t
Xbit_r389_c56 bl[56] br[56] wl[389] vdd gnd cell_6t
Xbit_r390_c56 bl[56] br[56] wl[390] vdd gnd cell_6t
Xbit_r391_c56 bl[56] br[56] wl[391] vdd gnd cell_6t
Xbit_r392_c56 bl[56] br[56] wl[392] vdd gnd cell_6t
Xbit_r393_c56 bl[56] br[56] wl[393] vdd gnd cell_6t
Xbit_r394_c56 bl[56] br[56] wl[394] vdd gnd cell_6t
Xbit_r395_c56 bl[56] br[56] wl[395] vdd gnd cell_6t
Xbit_r396_c56 bl[56] br[56] wl[396] vdd gnd cell_6t
Xbit_r397_c56 bl[56] br[56] wl[397] vdd gnd cell_6t
Xbit_r398_c56 bl[56] br[56] wl[398] vdd gnd cell_6t
Xbit_r399_c56 bl[56] br[56] wl[399] vdd gnd cell_6t
Xbit_r400_c56 bl[56] br[56] wl[400] vdd gnd cell_6t
Xbit_r401_c56 bl[56] br[56] wl[401] vdd gnd cell_6t
Xbit_r402_c56 bl[56] br[56] wl[402] vdd gnd cell_6t
Xbit_r403_c56 bl[56] br[56] wl[403] vdd gnd cell_6t
Xbit_r404_c56 bl[56] br[56] wl[404] vdd gnd cell_6t
Xbit_r405_c56 bl[56] br[56] wl[405] vdd gnd cell_6t
Xbit_r406_c56 bl[56] br[56] wl[406] vdd gnd cell_6t
Xbit_r407_c56 bl[56] br[56] wl[407] vdd gnd cell_6t
Xbit_r408_c56 bl[56] br[56] wl[408] vdd gnd cell_6t
Xbit_r409_c56 bl[56] br[56] wl[409] vdd gnd cell_6t
Xbit_r410_c56 bl[56] br[56] wl[410] vdd gnd cell_6t
Xbit_r411_c56 bl[56] br[56] wl[411] vdd gnd cell_6t
Xbit_r412_c56 bl[56] br[56] wl[412] vdd gnd cell_6t
Xbit_r413_c56 bl[56] br[56] wl[413] vdd gnd cell_6t
Xbit_r414_c56 bl[56] br[56] wl[414] vdd gnd cell_6t
Xbit_r415_c56 bl[56] br[56] wl[415] vdd gnd cell_6t
Xbit_r416_c56 bl[56] br[56] wl[416] vdd gnd cell_6t
Xbit_r417_c56 bl[56] br[56] wl[417] vdd gnd cell_6t
Xbit_r418_c56 bl[56] br[56] wl[418] vdd gnd cell_6t
Xbit_r419_c56 bl[56] br[56] wl[419] vdd gnd cell_6t
Xbit_r420_c56 bl[56] br[56] wl[420] vdd gnd cell_6t
Xbit_r421_c56 bl[56] br[56] wl[421] vdd gnd cell_6t
Xbit_r422_c56 bl[56] br[56] wl[422] vdd gnd cell_6t
Xbit_r423_c56 bl[56] br[56] wl[423] vdd gnd cell_6t
Xbit_r424_c56 bl[56] br[56] wl[424] vdd gnd cell_6t
Xbit_r425_c56 bl[56] br[56] wl[425] vdd gnd cell_6t
Xbit_r426_c56 bl[56] br[56] wl[426] vdd gnd cell_6t
Xbit_r427_c56 bl[56] br[56] wl[427] vdd gnd cell_6t
Xbit_r428_c56 bl[56] br[56] wl[428] vdd gnd cell_6t
Xbit_r429_c56 bl[56] br[56] wl[429] vdd gnd cell_6t
Xbit_r430_c56 bl[56] br[56] wl[430] vdd gnd cell_6t
Xbit_r431_c56 bl[56] br[56] wl[431] vdd gnd cell_6t
Xbit_r432_c56 bl[56] br[56] wl[432] vdd gnd cell_6t
Xbit_r433_c56 bl[56] br[56] wl[433] vdd gnd cell_6t
Xbit_r434_c56 bl[56] br[56] wl[434] vdd gnd cell_6t
Xbit_r435_c56 bl[56] br[56] wl[435] vdd gnd cell_6t
Xbit_r436_c56 bl[56] br[56] wl[436] vdd gnd cell_6t
Xbit_r437_c56 bl[56] br[56] wl[437] vdd gnd cell_6t
Xbit_r438_c56 bl[56] br[56] wl[438] vdd gnd cell_6t
Xbit_r439_c56 bl[56] br[56] wl[439] vdd gnd cell_6t
Xbit_r440_c56 bl[56] br[56] wl[440] vdd gnd cell_6t
Xbit_r441_c56 bl[56] br[56] wl[441] vdd gnd cell_6t
Xbit_r442_c56 bl[56] br[56] wl[442] vdd gnd cell_6t
Xbit_r443_c56 bl[56] br[56] wl[443] vdd gnd cell_6t
Xbit_r444_c56 bl[56] br[56] wl[444] vdd gnd cell_6t
Xbit_r445_c56 bl[56] br[56] wl[445] vdd gnd cell_6t
Xbit_r446_c56 bl[56] br[56] wl[446] vdd gnd cell_6t
Xbit_r447_c56 bl[56] br[56] wl[447] vdd gnd cell_6t
Xbit_r448_c56 bl[56] br[56] wl[448] vdd gnd cell_6t
Xbit_r449_c56 bl[56] br[56] wl[449] vdd gnd cell_6t
Xbit_r450_c56 bl[56] br[56] wl[450] vdd gnd cell_6t
Xbit_r451_c56 bl[56] br[56] wl[451] vdd gnd cell_6t
Xbit_r452_c56 bl[56] br[56] wl[452] vdd gnd cell_6t
Xbit_r453_c56 bl[56] br[56] wl[453] vdd gnd cell_6t
Xbit_r454_c56 bl[56] br[56] wl[454] vdd gnd cell_6t
Xbit_r455_c56 bl[56] br[56] wl[455] vdd gnd cell_6t
Xbit_r456_c56 bl[56] br[56] wl[456] vdd gnd cell_6t
Xbit_r457_c56 bl[56] br[56] wl[457] vdd gnd cell_6t
Xbit_r458_c56 bl[56] br[56] wl[458] vdd gnd cell_6t
Xbit_r459_c56 bl[56] br[56] wl[459] vdd gnd cell_6t
Xbit_r460_c56 bl[56] br[56] wl[460] vdd gnd cell_6t
Xbit_r461_c56 bl[56] br[56] wl[461] vdd gnd cell_6t
Xbit_r462_c56 bl[56] br[56] wl[462] vdd gnd cell_6t
Xbit_r463_c56 bl[56] br[56] wl[463] vdd gnd cell_6t
Xbit_r464_c56 bl[56] br[56] wl[464] vdd gnd cell_6t
Xbit_r465_c56 bl[56] br[56] wl[465] vdd gnd cell_6t
Xbit_r466_c56 bl[56] br[56] wl[466] vdd gnd cell_6t
Xbit_r467_c56 bl[56] br[56] wl[467] vdd gnd cell_6t
Xbit_r468_c56 bl[56] br[56] wl[468] vdd gnd cell_6t
Xbit_r469_c56 bl[56] br[56] wl[469] vdd gnd cell_6t
Xbit_r470_c56 bl[56] br[56] wl[470] vdd gnd cell_6t
Xbit_r471_c56 bl[56] br[56] wl[471] vdd gnd cell_6t
Xbit_r472_c56 bl[56] br[56] wl[472] vdd gnd cell_6t
Xbit_r473_c56 bl[56] br[56] wl[473] vdd gnd cell_6t
Xbit_r474_c56 bl[56] br[56] wl[474] vdd gnd cell_6t
Xbit_r475_c56 bl[56] br[56] wl[475] vdd gnd cell_6t
Xbit_r476_c56 bl[56] br[56] wl[476] vdd gnd cell_6t
Xbit_r477_c56 bl[56] br[56] wl[477] vdd gnd cell_6t
Xbit_r478_c56 bl[56] br[56] wl[478] vdd gnd cell_6t
Xbit_r479_c56 bl[56] br[56] wl[479] vdd gnd cell_6t
Xbit_r480_c56 bl[56] br[56] wl[480] vdd gnd cell_6t
Xbit_r481_c56 bl[56] br[56] wl[481] vdd gnd cell_6t
Xbit_r482_c56 bl[56] br[56] wl[482] vdd gnd cell_6t
Xbit_r483_c56 bl[56] br[56] wl[483] vdd gnd cell_6t
Xbit_r484_c56 bl[56] br[56] wl[484] vdd gnd cell_6t
Xbit_r485_c56 bl[56] br[56] wl[485] vdd gnd cell_6t
Xbit_r486_c56 bl[56] br[56] wl[486] vdd gnd cell_6t
Xbit_r487_c56 bl[56] br[56] wl[487] vdd gnd cell_6t
Xbit_r488_c56 bl[56] br[56] wl[488] vdd gnd cell_6t
Xbit_r489_c56 bl[56] br[56] wl[489] vdd gnd cell_6t
Xbit_r490_c56 bl[56] br[56] wl[490] vdd gnd cell_6t
Xbit_r491_c56 bl[56] br[56] wl[491] vdd gnd cell_6t
Xbit_r492_c56 bl[56] br[56] wl[492] vdd gnd cell_6t
Xbit_r493_c56 bl[56] br[56] wl[493] vdd gnd cell_6t
Xbit_r494_c56 bl[56] br[56] wl[494] vdd gnd cell_6t
Xbit_r495_c56 bl[56] br[56] wl[495] vdd gnd cell_6t
Xbit_r496_c56 bl[56] br[56] wl[496] vdd gnd cell_6t
Xbit_r497_c56 bl[56] br[56] wl[497] vdd gnd cell_6t
Xbit_r498_c56 bl[56] br[56] wl[498] vdd gnd cell_6t
Xbit_r499_c56 bl[56] br[56] wl[499] vdd gnd cell_6t
Xbit_r500_c56 bl[56] br[56] wl[500] vdd gnd cell_6t
Xbit_r501_c56 bl[56] br[56] wl[501] vdd gnd cell_6t
Xbit_r502_c56 bl[56] br[56] wl[502] vdd gnd cell_6t
Xbit_r503_c56 bl[56] br[56] wl[503] vdd gnd cell_6t
Xbit_r504_c56 bl[56] br[56] wl[504] vdd gnd cell_6t
Xbit_r505_c56 bl[56] br[56] wl[505] vdd gnd cell_6t
Xbit_r506_c56 bl[56] br[56] wl[506] vdd gnd cell_6t
Xbit_r507_c56 bl[56] br[56] wl[507] vdd gnd cell_6t
Xbit_r508_c56 bl[56] br[56] wl[508] vdd gnd cell_6t
Xbit_r509_c56 bl[56] br[56] wl[509] vdd gnd cell_6t
Xbit_r510_c56 bl[56] br[56] wl[510] vdd gnd cell_6t
Xbit_r511_c56 bl[56] br[56] wl[511] vdd gnd cell_6t
Xbit_r0_c57 bl[57] br[57] wl[0] vdd gnd cell_6t
Xbit_r1_c57 bl[57] br[57] wl[1] vdd gnd cell_6t
Xbit_r2_c57 bl[57] br[57] wl[2] vdd gnd cell_6t
Xbit_r3_c57 bl[57] br[57] wl[3] vdd gnd cell_6t
Xbit_r4_c57 bl[57] br[57] wl[4] vdd gnd cell_6t
Xbit_r5_c57 bl[57] br[57] wl[5] vdd gnd cell_6t
Xbit_r6_c57 bl[57] br[57] wl[6] vdd gnd cell_6t
Xbit_r7_c57 bl[57] br[57] wl[7] vdd gnd cell_6t
Xbit_r8_c57 bl[57] br[57] wl[8] vdd gnd cell_6t
Xbit_r9_c57 bl[57] br[57] wl[9] vdd gnd cell_6t
Xbit_r10_c57 bl[57] br[57] wl[10] vdd gnd cell_6t
Xbit_r11_c57 bl[57] br[57] wl[11] vdd gnd cell_6t
Xbit_r12_c57 bl[57] br[57] wl[12] vdd gnd cell_6t
Xbit_r13_c57 bl[57] br[57] wl[13] vdd gnd cell_6t
Xbit_r14_c57 bl[57] br[57] wl[14] vdd gnd cell_6t
Xbit_r15_c57 bl[57] br[57] wl[15] vdd gnd cell_6t
Xbit_r16_c57 bl[57] br[57] wl[16] vdd gnd cell_6t
Xbit_r17_c57 bl[57] br[57] wl[17] vdd gnd cell_6t
Xbit_r18_c57 bl[57] br[57] wl[18] vdd gnd cell_6t
Xbit_r19_c57 bl[57] br[57] wl[19] vdd gnd cell_6t
Xbit_r20_c57 bl[57] br[57] wl[20] vdd gnd cell_6t
Xbit_r21_c57 bl[57] br[57] wl[21] vdd gnd cell_6t
Xbit_r22_c57 bl[57] br[57] wl[22] vdd gnd cell_6t
Xbit_r23_c57 bl[57] br[57] wl[23] vdd gnd cell_6t
Xbit_r24_c57 bl[57] br[57] wl[24] vdd gnd cell_6t
Xbit_r25_c57 bl[57] br[57] wl[25] vdd gnd cell_6t
Xbit_r26_c57 bl[57] br[57] wl[26] vdd gnd cell_6t
Xbit_r27_c57 bl[57] br[57] wl[27] vdd gnd cell_6t
Xbit_r28_c57 bl[57] br[57] wl[28] vdd gnd cell_6t
Xbit_r29_c57 bl[57] br[57] wl[29] vdd gnd cell_6t
Xbit_r30_c57 bl[57] br[57] wl[30] vdd gnd cell_6t
Xbit_r31_c57 bl[57] br[57] wl[31] vdd gnd cell_6t
Xbit_r32_c57 bl[57] br[57] wl[32] vdd gnd cell_6t
Xbit_r33_c57 bl[57] br[57] wl[33] vdd gnd cell_6t
Xbit_r34_c57 bl[57] br[57] wl[34] vdd gnd cell_6t
Xbit_r35_c57 bl[57] br[57] wl[35] vdd gnd cell_6t
Xbit_r36_c57 bl[57] br[57] wl[36] vdd gnd cell_6t
Xbit_r37_c57 bl[57] br[57] wl[37] vdd gnd cell_6t
Xbit_r38_c57 bl[57] br[57] wl[38] vdd gnd cell_6t
Xbit_r39_c57 bl[57] br[57] wl[39] vdd gnd cell_6t
Xbit_r40_c57 bl[57] br[57] wl[40] vdd gnd cell_6t
Xbit_r41_c57 bl[57] br[57] wl[41] vdd gnd cell_6t
Xbit_r42_c57 bl[57] br[57] wl[42] vdd gnd cell_6t
Xbit_r43_c57 bl[57] br[57] wl[43] vdd gnd cell_6t
Xbit_r44_c57 bl[57] br[57] wl[44] vdd gnd cell_6t
Xbit_r45_c57 bl[57] br[57] wl[45] vdd gnd cell_6t
Xbit_r46_c57 bl[57] br[57] wl[46] vdd gnd cell_6t
Xbit_r47_c57 bl[57] br[57] wl[47] vdd gnd cell_6t
Xbit_r48_c57 bl[57] br[57] wl[48] vdd gnd cell_6t
Xbit_r49_c57 bl[57] br[57] wl[49] vdd gnd cell_6t
Xbit_r50_c57 bl[57] br[57] wl[50] vdd gnd cell_6t
Xbit_r51_c57 bl[57] br[57] wl[51] vdd gnd cell_6t
Xbit_r52_c57 bl[57] br[57] wl[52] vdd gnd cell_6t
Xbit_r53_c57 bl[57] br[57] wl[53] vdd gnd cell_6t
Xbit_r54_c57 bl[57] br[57] wl[54] vdd gnd cell_6t
Xbit_r55_c57 bl[57] br[57] wl[55] vdd gnd cell_6t
Xbit_r56_c57 bl[57] br[57] wl[56] vdd gnd cell_6t
Xbit_r57_c57 bl[57] br[57] wl[57] vdd gnd cell_6t
Xbit_r58_c57 bl[57] br[57] wl[58] vdd gnd cell_6t
Xbit_r59_c57 bl[57] br[57] wl[59] vdd gnd cell_6t
Xbit_r60_c57 bl[57] br[57] wl[60] vdd gnd cell_6t
Xbit_r61_c57 bl[57] br[57] wl[61] vdd gnd cell_6t
Xbit_r62_c57 bl[57] br[57] wl[62] vdd gnd cell_6t
Xbit_r63_c57 bl[57] br[57] wl[63] vdd gnd cell_6t
Xbit_r64_c57 bl[57] br[57] wl[64] vdd gnd cell_6t
Xbit_r65_c57 bl[57] br[57] wl[65] vdd gnd cell_6t
Xbit_r66_c57 bl[57] br[57] wl[66] vdd gnd cell_6t
Xbit_r67_c57 bl[57] br[57] wl[67] vdd gnd cell_6t
Xbit_r68_c57 bl[57] br[57] wl[68] vdd gnd cell_6t
Xbit_r69_c57 bl[57] br[57] wl[69] vdd gnd cell_6t
Xbit_r70_c57 bl[57] br[57] wl[70] vdd gnd cell_6t
Xbit_r71_c57 bl[57] br[57] wl[71] vdd gnd cell_6t
Xbit_r72_c57 bl[57] br[57] wl[72] vdd gnd cell_6t
Xbit_r73_c57 bl[57] br[57] wl[73] vdd gnd cell_6t
Xbit_r74_c57 bl[57] br[57] wl[74] vdd gnd cell_6t
Xbit_r75_c57 bl[57] br[57] wl[75] vdd gnd cell_6t
Xbit_r76_c57 bl[57] br[57] wl[76] vdd gnd cell_6t
Xbit_r77_c57 bl[57] br[57] wl[77] vdd gnd cell_6t
Xbit_r78_c57 bl[57] br[57] wl[78] vdd gnd cell_6t
Xbit_r79_c57 bl[57] br[57] wl[79] vdd gnd cell_6t
Xbit_r80_c57 bl[57] br[57] wl[80] vdd gnd cell_6t
Xbit_r81_c57 bl[57] br[57] wl[81] vdd gnd cell_6t
Xbit_r82_c57 bl[57] br[57] wl[82] vdd gnd cell_6t
Xbit_r83_c57 bl[57] br[57] wl[83] vdd gnd cell_6t
Xbit_r84_c57 bl[57] br[57] wl[84] vdd gnd cell_6t
Xbit_r85_c57 bl[57] br[57] wl[85] vdd gnd cell_6t
Xbit_r86_c57 bl[57] br[57] wl[86] vdd gnd cell_6t
Xbit_r87_c57 bl[57] br[57] wl[87] vdd gnd cell_6t
Xbit_r88_c57 bl[57] br[57] wl[88] vdd gnd cell_6t
Xbit_r89_c57 bl[57] br[57] wl[89] vdd gnd cell_6t
Xbit_r90_c57 bl[57] br[57] wl[90] vdd gnd cell_6t
Xbit_r91_c57 bl[57] br[57] wl[91] vdd gnd cell_6t
Xbit_r92_c57 bl[57] br[57] wl[92] vdd gnd cell_6t
Xbit_r93_c57 bl[57] br[57] wl[93] vdd gnd cell_6t
Xbit_r94_c57 bl[57] br[57] wl[94] vdd gnd cell_6t
Xbit_r95_c57 bl[57] br[57] wl[95] vdd gnd cell_6t
Xbit_r96_c57 bl[57] br[57] wl[96] vdd gnd cell_6t
Xbit_r97_c57 bl[57] br[57] wl[97] vdd gnd cell_6t
Xbit_r98_c57 bl[57] br[57] wl[98] vdd gnd cell_6t
Xbit_r99_c57 bl[57] br[57] wl[99] vdd gnd cell_6t
Xbit_r100_c57 bl[57] br[57] wl[100] vdd gnd cell_6t
Xbit_r101_c57 bl[57] br[57] wl[101] vdd gnd cell_6t
Xbit_r102_c57 bl[57] br[57] wl[102] vdd gnd cell_6t
Xbit_r103_c57 bl[57] br[57] wl[103] vdd gnd cell_6t
Xbit_r104_c57 bl[57] br[57] wl[104] vdd gnd cell_6t
Xbit_r105_c57 bl[57] br[57] wl[105] vdd gnd cell_6t
Xbit_r106_c57 bl[57] br[57] wl[106] vdd gnd cell_6t
Xbit_r107_c57 bl[57] br[57] wl[107] vdd gnd cell_6t
Xbit_r108_c57 bl[57] br[57] wl[108] vdd gnd cell_6t
Xbit_r109_c57 bl[57] br[57] wl[109] vdd gnd cell_6t
Xbit_r110_c57 bl[57] br[57] wl[110] vdd gnd cell_6t
Xbit_r111_c57 bl[57] br[57] wl[111] vdd gnd cell_6t
Xbit_r112_c57 bl[57] br[57] wl[112] vdd gnd cell_6t
Xbit_r113_c57 bl[57] br[57] wl[113] vdd gnd cell_6t
Xbit_r114_c57 bl[57] br[57] wl[114] vdd gnd cell_6t
Xbit_r115_c57 bl[57] br[57] wl[115] vdd gnd cell_6t
Xbit_r116_c57 bl[57] br[57] wl[116] vdd gnd cell_6t
Xbit_r117_c57 bl[57] br[57] wl[117] vdd gnd cell_6t
Xbit_r118_c57 bl[57] br[57] wl[118] vdd gnd cell_6t
Xbit_r119_c57 bl[57] br[57] wl[119] vdd gnd cell_6t
Xbit_r120_c57 bl[57] br[57] wl[120] vdd gnd cell_6t
Xbit_r121_c57 bl[57] br[57] wl[121] vdd gnd cell_6t
Xbit_r122_c57 bl[57] br[57] wl[122] vdd gnd cell_6t
Xbit_r123_c57 bl[57] br[57] wl[123] vdd gnd cell_6t
Xbit_r124_c57 bl[57] br[57] wl[124] vdd gnd cell_6t
Xbit_r125_c57 bl[57] br[57] wl[125] vdd gnd cell_6t
Xbit_r126_c57 bl[57] br[57] wl[126] vdd gnd cell_6t
Xbit_r127_c57 bl[57] br[57] wl[127] vdd gnd cell_6t
Xbit_r128_c57 bl[57] br[57] wl[128] vdd gnd cell_6t
Xbit_r129_c57 bl[57] br[57] wl[129] vdd gnd cell_6t
Xbit_r130_c57 bl[57] br[57] wl[130] vdd gnd cell_6t
Xbit_r131_c57 bl[57] br[57] wl[131] vdd gnd cell_6t
Xbit_r132_c57 bl[57] br[57] wl[132] vdd gnd cell_6t
Xbit_r133_c57 bl[57] br[57] wl[133] vdd gnd cell_6t
Xbit_r134_c57 bl[57] br[57] wl[134] vdd gnd cell_6t
Xbit_r135_c57 bl[57] br[57] wl[135] vdd gnd cell_6t
Xbit_r136_c57 bl[57] br[57] wl[136] vdd gnd cell_6t
Xbit_r137_c57 bl[57] br[57] wl[137] vdd gnd cell_6t
Xbit_r138_c57 bl[57] br[57] wl[138] vdd gnd cell_6t
Xbit_r139_c57 bl[57] br[57] wl[139] vdd gnd cell_6t
Xbit_r140_c57 bl[57] br[57] wl[140] vdd gnd cell_6t
Xbit_r141_c57 bl[57] br[57] wl[141] vdd gnd cell_6t
Xbit_r142_c57 bl[57] br[57] wl[142] vdd gnd cell_6t
Xbit_r143_c57 bl[57] br[57] wl[143] vdd gnd cell_6t
Xbit_r144_c57 bl[57] br[57] wl[144] vdd gnd cell_6t
Xbit_r145_c57 bl[57] br[57] wl[145] vdd gnd cell_6t
Xbit_r146_c57 bl[57] br[57] wl[146] vdd gnd cell_6t
Xbit_r147_c57 bl[57] br[57] wl[147] vdd gnd cell_6t
Xbit_r148_c57 bl[57] br[57] wl[148] vdd gnd cell_6t
Xbit_r149_c57 bl[57] br[57] wl[149] vdd gnd cell_6t
Xbit_r150_c57 bl[57] br[57] wl[150] vdd gnd cell_6t
Xbit_r151_c57 bl[57] br[57] wl[151] vdd gnd cell_6t
Xbit_r152_c57 bl[57] br[57] wl[152] vdd gnd cell_6t
Xbit_r153_c57 bl[57] br[57] wl[153] vdd gnd cell_6t
Xbit_r154_c57 bl[57] br[57] wl[154] vdd gnd cell_6t
Xbit_r155_c57 bl[57] br[57] wl[155] vdd gnd cell_6t
Xbit_r156_c57 bl[57] br[57] wl[156] vdd gnd cell_6t
Xbit_r157_c57 bl[57] br[57] wl[157] vdd gnd cell_6t
Xbit_r158_c57 bl[57] br[57] wl[158] vdd gnd cell_6t
Xbit_r159_c57 bl[57] br[57] wl[159] vdd gnd cell_6t
Xbit_r160_c57 bl[57] br[57] wl[160] vdd gnd cell_6t
Xbit_r161_c57 bl[57] br[57] wl[161] vdd gnd cell_6t
Xbit_r162_c57 bl[57] br[57] wl[162] vdd gnd cell_6t
Xbit_r163_c57 bl[57] br[57] wl[163] vdd gnd cell_6t
Xbit_r164_c57 bl[57] br[57] wl[164] vdd gnd cell_6t
Xbit_r165_c57 bl[57] br[57] wl[165] vdd gnd cell_6t
Xbit_r166_c57 bl[57] br[57] wl[166] vdd gnd cell_6t
Xbit_r167_c57 bl[57] br[57] wl[167] vdd gnd cell_6t
Xbit_r168_c57 bl[57] br[57] wl[168] vdd gnd cell_6t
Xbit_r169_c57 bl[57] br[57] wl[169] vdd gnd cell_6t
Xbit_r170_c57 bl[57] br[57] wl[170] vdd gnd cell_6t
Xbit_r171_c57 bl[57] br[57] wl[171] vdd gnd cell_6t
Xbit_r172_c57 bl[57] br[57] wl[172] vdd gnd cell_6t
Xbit_r173_c57 bl[57] br[57] wl[173] vdd gnd cell_6t
Xbit_r174_c57 bl[57] br[57] wl[174] vdd gnd cell_6t
Xbit_r175_c57 bl[57] br[57] wl[175] vdd gnd cell_6t
Xbit_r176_c57 bl[57] br[57] wl[176] vdd gnd cell_6t
Xbit_r177_c57 bl[57] br[57] wl[177] vdd gnd cell_6t
Xbit_r178_c57 bl[57] br[57] wl[178] vdd gnd cell_6t
Xbit_r179_c57 bl[57] br[57] wl[179] vdd gnd cell_6t
Xbit_r180_c57 bl[57] br[57] wl[180] vdd gnd cell_6t
Xbit_r181_c57 bl[57] br[57] wl[181] vdd gnd cell_6t
Xbit_r182_c57 bl[57] br[57] wl[182] vdd gnd cell_6t
Xbit_r183_c57 bl[57] br[57] wl[183] vdd gnd cell_6t
Xbit_r184_c57 bl[57] br[57] wl[184] vdd gnd cell_6t
Xbit_r185_c57 bl[57] br[57] wl[185] vdd gnd cell_6t
Xbit_r186_c57 bl[57] br[57] wl[186] vdd gnd cell_6t
Xbit_r187_c57 bl[57] br[57] wl[187] vdd gnd cell_6t
Xbit_r188_c57 bl[57] br[57] wl[188] vdd gnd cell_6t
Xbit_r189_c57 bl[57] br[57] wl[189] vdd gnd cell_6t
Xbit_r190_c57 bl[57] br[57] wl[190] vdd gnd cell_6t
Xbit_r191_c57 bl[57] br[57] wl[191] vdd gnd cell_6t
Xbit_r192_c57 bl[57] br[57] wl[192] vdd gnd cell_6t
Xbit_r193_c57 bl[57] br[57] wl[193] vdd gnd cell_6t
Xbit_r194_c57 bl[57] br[57] wl[194] vdd gnd cell_6t
Xbit_r195_c57 bl[57] br[57] wl[195] vdd gnd cell_6t
Xbit_r196_c57 bl[57] br[57] wl[196] vdd gnd cell_6t
Xbit_r197_c57 bl[57] br[57] wl[197] vdd gnd cell_6t
Xbit_r198_c57 bl[57] br[57] wl[198] vdd gnd cell_6t
Xbit_r199_c57 bl[57] br[57] wl[199] vdd gnd cell_6t
Xbit_r200_c57 bl[57] br[57] wl[200] vdd gnd cell_6t
Xbit_r201_c57 bl[57] br[57] wl[201] vdd gnd cell_6t
Xbit_r202_c57 bl[57] br[57] wl[202] vdd gnd cell_6t
Xbit_r203_c57 bl[57] br[57] wl[203] vdd gnd cell_6t
Xbit_r204_c57 bl[57] br[57] wl[204] vdd gnd cell_6t
Xbit_r205_c57 bl[57] br[57] wl[205] vdd gnd cell_6t
Xbit_r206_c57 bl[57] br[57] wl[206] vdd gnd cell_6t
Xbit_r207_c57 bl[57] br[57] wl[207] vdd gnd cell_6t
Xbit_r208_c57 bl[57] br[57] wl[208] vdd gnd cell_6t
Xbit_r209_c57 bl[57] br[57] wl[209] vdd gnd cell_6t
Xbit_r210_c57 bl[57] br[57] wl[210] vdd gnd cell_6t
Xbit_r211_c57 bl[57] br[57] wl[211] vdd gnd cell_6t
Xbit_r212_c57 bl[57] br[57] wl[212] vdd gnd cell_6t
Xbit_r213_c57 bl[57] br[57] wl[213] vdd gnd cell_6t
Xbit_r214_c57 bl[57] br[57] wl[214] vdd gnd cell_6t
Xbit_r215_c57 bl[57] br[57] wl[215] vdd gnd cell_6t
Xbit_r216_c57 bl[57] br[57] wl[216] vdd gnd cell_6t
Xbit_r217_c57 bl[57] br[57] wl[217] vdd gnd cell_6t
Xbit_r218_c57 bl[57] br[57] wl[218] vdd gnd cell_6t
Xbit_r219_c57 bl[57] br[57] wl[219] vdd gnd cell_6t
Xbit_r220_c57 bl[57] br[57] wl[220] vdd gnd cell_6t
Xbit_r221_c57 bl[57] br[57] wl[221] vdd gnd cell_6t
Xbit_r222_c57 bl[57] br[57] wl[222] vdd gnd cell_6t
Xbit_r223_c57 bl[57] br[57] wl[223] vdd gnd cell_6t
Xbit_r224_c57 bl[57] br[57] wl[224] vdd gnd cell_6t
Xbit_r225_c57 bl[57] br[57] wl[225] vdd gnd cell_6t
Xbit_r226_c57 bl[57] br[57] wl[226] vdd gnd cell_6t
Xbit_r227_c57 bl[57] br[57] wl[227] vdd gnd cell_6t
Xbit_r228_c57 bl[57] br[57] wl[228] vdd gnd cell_6t
Xbit_r229_c57 bl[57] br[57] wl[229] vdd gnd cell_6t
Xbit_r230_c57 bl[57] br[57] wl[230] vdd gnd cell_6t
Xbit_r231_c57 bl[57] br[57] wl[231] vdd gnd cell_6t
Xbit_r232_c57 bl[57] br[57] wl[232] vdd gnd cell_6t
Xbit_r233_c57 bl[57] br[57] wl[233] vdd gnd cell_6t
Xbit_r234_c57 bl[57] br[57] wl[234] vdd gnd cell_6t
Xbit_r235_c57 bl[57] br[57] wl[235] vdd gnd cell_6t
Xbit_r236_c57 bl[57] br[57] wl[236] vdd gnd cell_6t
Xbit_r237_c57 bl[57] br[57] wl[237] vdd gnd cell_6t
Xbit_r238_c57 bl[57] br[57] wl[238] vdd gnd cell_6t
Xbit_r239_c57 bl[57] br[57] wl[239] vdd gnd cell_6t
Xbit_r240_c57 bl[57] br[57] wl[240] vdd gnd cell_6t
Xbit_r241_c57 bl[57] br[57] wl[241] vdd gnd cell_6t
Xbit_r242_c57 bl[57] br[57] wl[242] vdd gnd cell_6t
Xbit_r243_c57 bl[57] br[57] wl[243] vdd gnd cell_6t
Xbit_r244_c57 bl[57] br[57] wl[244] vdd gnd cell_6t
Xbit_r245_c57 bl[57] br[57] wl[245] vdd gnd cell_6t
Xbit_r246_c57 bl[57] br[57] wl[246] vdd gnd cell_6t
Xbit_r247_c57 bl[57] br[57] wl[247] vdd gnd cell_6t
Xbit_r248_c57 bl[57] br[57] wl[248] vdd gnd cell_6t
Xbit_r249_c57 bl[57] br[57] wl[249] vdd gnd cell_6t
Xbit_r250_c57 bl[57] br[57] wl[250] vdd gnd cell_6t
Xbit_r251_c57 bl[57] br[57] wl[251] vdd gnd cell_6t
Xbit_r252_c57 bl[57] br[57] wl[252] vdd gnd cell_6t
Xbit_r253_c57 bl[57] br[57] wl[253] vdd gnd cell_6t
Xbit_r254_c57 bl[57] br[57] wl[254] vdd gnd cell_6t
Xbit_r255_c57 bl[57] br[57] wl[255] vdd gnd cell_6t
Xbit_r256_c57 bl[57] br[57] wl[256] vdd gnd cell_6t
Xbit_r257_c57 bl[57] br[57] wl[257] vdd gnd cell_6t
Xbit_r258_c57 bl[57] br[57] wl[258] vdd gnd cell_6t
Xbit_r259_c57 bl[57] br[57] wl[259] vdd gnd cell_6t
Xbit_r260_c57 bl[57] br[57] wl[260] vdd gnd cell_6t
Xbit_r261_c57 bl[57] br[57] wl[261] vdd gnd cell_6t
Xbit_r262_c57 bl[57] br[57] wl[262] vdd gnd cell_6t
Xbit_r263_c57 bl[57] br[57] wl[263] vdd gnd cell_6t
Xbit_r264_c57 bl[57] br[57] wl[264] vdd gnd cell_6t
Xbit_r265_c57 bl[57] br[57] wl[265] vdd gnd cell_6t
Xbit_r266_c57 bl[57] br[57] wl[266] vdd gnd cell_6t
Xbit_r267_c57 bl[57] br[57] wl[267] vdd gnd cell_6t
Xbit_r268_c57 bl[57] br[57] wl[268] vdd gnd cell_6t
Xbit_r269_c57 bl[57] br[57] wl[269] vdd gnd cell_6t
Xbit_r270_c57 bl[57] br[57] wl[270] vdd gnd cell_6t
Xbit_r271_c57 bl[57] br[57] wl[271] vdd gnd cell_6t
Xbit_r272_c57 bl[57] br[57] wl[272] vdd gnd cell_6t
Xbit_r273_c57 bl[57] br[57] wl[273] vdd gnd cell_6t
Xbit_r274_c57 bl[57] br[57] wl[274] vdd gnd cell_6t
Xbit_r275_c57 bl[57] br[57] wl[275] vdd gnd cell_6t
Xbit_r276_c57 bl[57] br[57] wl[276] vdd gnd cell_6t
Xbit_r277_c57 bl[57] br[57] wl[277] vdd gnd cell_6t
Xbit_r278_c57 bl[57] br[57] wl[278] vdd gnd cell_6t
Xbit_r279_c57 bl[57] br[57] wl[279] vdd gnd cell_6t
Xbit_r280_c57 bl[57] br[57] wl[280] vdd gnd cell_6t
Xbit_r281_c57 bl[57] br[57] wl[281] vdd gnd cell_6t
Xbit_r282_c57 bl[57] br[57] wl[282] vdd gnd cell_6t
Xbit_r283_c57 bl[57] br[57] wl[283] vdd gnd cell_6t
Xbit_r284_c57 bl[57] br[57] wl[284] vdd gnd cell_6t
Xbit_r285_c57 bl[57] br[57] wl[285] vdd gnd cell_6t
Xbit_r286_c57 bl[57] br[57] wl[286] vdd gnd cell_6t
Xbit_r287_c57 bl[57] br[57] wl[287] vdd gnd cell_6t
Xbit_r288_c57 bl[57] br[57] wl[288] vdd gnd cell_6t
Xbit_r289_c57 bl[57] br[57] wl[289] vdd gnd cell_6t
Xbit_r290_c57 bl[57] br[57] wl[290] vdd gnd cell_6t
Xbit_r291_c57 bl[57] br[57] wl[291] vdd gnd cell_6t
Xbit_r292_c57 bl[57] br[57] wl[292] vdd gnd cell_6t
Xbit_r293_c57 bl[57] br[57] wl[293] vdd gnd cell_6t
Xbit_r294_c57 bl[57] br[57] wl[294] vdd gnd cell_6t
Xbit_r295_c57 bl[57] br[57] wl[295] vdd gnd cell_6t
Xbit_r296_c57 bl[57] br[57] wl[296] vdd gnd cell_6t
Xbit_r297_c57 bl[57] br[57] wl[297] vdd gnd cell_6t
Xbit_r298_c57 bl[57] br[57] wl[298] vdd gnd cell_6t
Xbit_r299_c57 bl[57] br[57] wl[299] vdd gnd cell_6t
Xbit_r300_c57 bl[57] br[57] wl[300] vdd gnd cell_6t
Xbit_r301_c57 bl[57] br[57] wl[301] vdd gnd cell_6t
Xbit_r302_c57 bl[57] br[57] wl[302] vdd gnd cell_6t
Xbit_r303_c57 bl[57] br[57] wl[303] vdd gnd cell_6t
Xbit_r304_c57 bl[57] br[57] wl[304] vdd gnd cell_6t
Xbit_r305_c57 bl[57] br[57] wl[305] vdd gnd cell_6t
Xbit_r306_c57 bl[57] br[57] wl[306] vdd gnd cell_6t
Xbit_r307_c57 bl[57] br[57] wl[307] vdd gnd cell_6t
Xbit_r308_c57 bl[57] br[57] wl[308] vdd gnd cell_6t
Xbit_r309_c57 bl[57] br[57] wl[309] vdd gnd cell_6t
Xbit_r310_c57 bl[57] br[57] wl[310] vdd gnd cell_6t
Xbit_r311_c57 bl[57] br[57] wl[311] vdd gnd cell_6t
Xbit_r312_c57 bl[57] br[57] wl[312] vdd gnd cell_6t
Xbit_r313_c57 bl[57] br[57] wl[313] vdd gnd cell_6t
Xbit_r314_c57 bl[57] br[57] wl[314] vdd gnd cell_6t
Xbit_r315_c57 bl[57] br[57] wl[315] vdd gnd cell_6t
Xbit_r316_c57 bl[57] br[57] wl[316] vdd gnd cell_6t
Xbit_r317_c57 bl[57] br[57] wl[317] vdd gnd cell_6t
Xbit_r318_c57 bl[57] br[57] wl[318] vdd gnd cell_6t
Xbit_r319_c57 bl[57] br[57] wl[319] vdd gnd cell_6t
Xbit_r320_c57 bl[57] br[57] wl[320] vdd gnd cell_6t
Xbit_r321_c57 bl[57] br[57] wl[321] vdd gnd cell_6t
Xbit_r322_c57 bl[57] br[57] wl[322] vdd gnd cell_6t
Xbit_r323_c57 bl[57] br[57] wl[323] vdd gnd cell_6t
Xbit_r324_c57 bl[57] br[57] wl[324] vdd gnd cell_6t
Xbit_r325_c57 bl[57] br[57] wl[325] vdd gnd cell_6t
Xbit_r326_c57 bl[57] br[57] wl[326] vdd gnd cell_6t
Xbit_r327_c57 bl[57] br[57] wl[327] vdd gnd cell_6t
Xbit_r328_c57 bl[57] br[57] wl[328] vdd gnd cell_6t
Xbit_r329_c57 bl[57] br[57] wl[329] vdd gnd cell_6t
Xbit_r330_c57 bl[57] br[57] wl[330] vdd gnd cell_6t
Xbit_r331_c57 bl[57] br[57] wl[331] vdd gnd cell_6t
Xbit_r332_c57 bl[57] br[57] wl[332] vdd gnd cell_6t
Xbit_r333_c57 bl[57] br[57] wl[333] vdd gnd cell_6t
Xbit_r334_c57 bl[57] br[57] wl[334] vdd gnd cell_6t
Xbit_r335_c57 bl[57] br[57] wl[335] vdd gnd cell_6t
Xbit_r336_c57 bl[57] br[57] wl[336] vdd gnd cell_6t
Xbit_r337_c57 bl[57] br[57] wl[337] vdd gnd cell_6t
Xbit_r338_c57 bl[57] br[57] wl[338] vdd gnd cell_6t
Xbit_r339_c57 bl[57] br[57] wl[339] vdd gnd cell_6t
Xbit_r340_c57 bl[57] br[57] wl[340] vdd gnd cell_6t
Xbit_r341_c57 bl[57] br[57] wl[341] vdd gnd cell_6t
Xbit_r342_c57 bl[57] br[57] wl[342] vdd gnd cell_6t
Xbit_r343_c57 bl[57] br[57] wl[343] vdd gnd cell_6t
Xbit_r344_c57 bl[57] br[57] wl[344] vdd gnd cell_6t
Xbit_r345_c57 bl[57] br[57] wl[345] vdd gnd cell_6t
Xbit_r346_c57 bl[57] br[57] wl[346] vdd gnd cell_6t
Xbit_r347_c57 bl[57] br[57] wl[347] vdd gnd cell_6t
Xbit_r348_c57 bl[57] br[57] wl[348] vdd gnd cell_6t
Xbit_r349_c57 bl[57] br[57] wl[349] vdd gnd cell_6t
Xbit_r350_c57 bl[57] br[57] wl[350] vdd gnd cell_6t
Xbit_r351_c57 bl[57] br[57] wl[351] vdd gnd cell_6t
Xbit_r352_c57 bl[57] br[57] wl[352] vdd gnd cell_6t
Xbit_r353_c57 bl[57] br[57] wl[353] vdd gnd cell_6t
Xbit_r354_c57 bl[57] br[57] wl[354] vdd gnd cell_6t
Xbit_r355_c57 bl[57] br[57] wl[355] vdd gnd cell_6t
Xbit_r356_c57 bl[57] br[57] wl[356] vdd gnd cell_6t
Xbit_r357_c57 bl[57] br[57] wl[357] vdd gnd cell_6t
Xbit_r358_c57 bl[57] br[57] wl[358] vdd gnd cell_6t
Xbit_r359_c57 bl[57] br[57] wl[359] vdd gnd cell_6t
Xbit_r360_c57 bl[57] br[57] wl[360] vdd gnd cell_6t
Xbit_r361_c57 bl[57] br[57] wl[361] vdd gnd cell_6t
Xbit_r362_c57 bl[57] br[57] wl[362] vdd gnd cell_6t
Xbit_r363_c57 bl[57] br[57] wl[363] vdd gnd cell_6t
Xbit_r364_c57 bl[57] br[57] wl[364] vdd gnd cell_6t
Xbit_r365_c57 bl[57] br[57] wl[365] vdd gnd cell_6t
Xbit_r366_c57 bl[57] br[57] wl[366] vdd gnd cell_6t
Xbit_r367_c57 bl[57] br[57] wl[367] vdd gnd cell_6t
Xbit_r368_c57 bl[57] br[57] wl[368] vdd gnd cell_6t
Xbit_r369_c57 bl[57] br[57] wl[369] vdd gnd cell_6t
Xbit_r370_c57 bl[57] br[57] wl[370] vdd gnd cell_6t
Xbit_r371_c57 bl[57] br[57] wl[371] vdd gnd cell_6t
Xbit_r372_c57 bl[57] br[57] wl[372] vdd gnd cell_6t
Xbit_r373_c57 bl[57] br[57] wl[373] vdd gnd cell_6t
Xbit_r374_c57 bl[57] br[57] wl[374] vdd gnd cell_6t
Xbit_r375_c57 bl[57] br[57] wl[375] vdd gnd cell_6t
Xbit_r376_c57 bl[57] br[57] wl[376] vdd gnd cell_6t
Xbit_r377_c57 bl[57] br[57] wl[377] vdd gnd cell_6t
Xbit_r378_c57 bl[57] br[57] wl[378] vdd gnd cell_6t
Xbit_r379_c57 bl[57] br[57] wl[379] vdd gnd cell_6t
Xbit_r380_c57 bl[57] br[57] wl[380] vdd gnd cell_6t
Xbit_r381_c57 bl[57] br[57] wl[381] vdd gnd cell_6t
Xbit_r382_c57 bl[57] br[57] wl[382] vdd gnd cell_6t
Xbit_r383_c57 bl[57] br[57] wl[383] vdd gnd cell_6t
Xbit_r384_c57 bl[57] br[57] wl[384] vdd gnd cell_6t
Xbit_r385_c57 bl[57] br[57] wl[385] vdd gnd cell_6t
Xbit_r386_c57 bl[57] br[57] wl[386] vdd gnd cell_6t
Xbit_r387_c57 bl[57] br[57] wl[387] vdd gnd cell_6t
Xbit_r388_c57 bl[57] br[57] wl[388] vdd gnd cell_6t
Xbit_r389_c57 bl[57] br[57] wl[389] vdd gnd cell_6t
Xbit_r390_c57 bl[57] br[57] wl[390] vdd gnd cell_6t
Xbit_r391_c57 bl[57] br[57] wl[391] vdd gnd cell_6t
Xbit_r392_c57 bl[57] br[57] wl[392] vdd gnd cell_6t
Xbit_r393_c57 bl[57] br[57] wl[393] vdd gnd cell_6t
Xbit_r394_c57 bl[57] br[57] wl[394] vdd gnd cell_6t
Xbit_r395_c57 bl[57] br[57] wl[395] vdd gnd cell_6t
Xbit_r396_c57 bl[57] br[57] wl[396] vdd gnd cell_6t
Xbit_r397_c57 bl[57] br[57] wl[397] vdd gnd cell_6t
Xbit_r398_c57 bl[57] br[57] wl[398] vdd gnd cell_6t
Xbit_r399_c57 bl[57] br[57] wl[399] vdd gnd cell_6t
Xbit_r400_c57 bl[57] br[57] wl[400] vdd gnd cell_6t
Xbit_r401_c57 bl[57] br[57] wl[401] vdd gnd cell_6t
Xbit_r402_c57 bl[57] br[57] wl[402] vdd gnd cell_6t
Xbit_r403_c57 bl[57] br[57] wl[403] vdd gnd cell_6t
Xbit_r404_c57 bl[57] br[57] wl[404] vdd gnd cell_6t
Xbit_r405_c57 bl[57] br[57] wl[405] vdd gnd cell_6t
Xbit_r406_c57 bl[57] br[57] wl[406] vdd gnd cell_6t
Xbit_r407_c57 bl[57] br[57] wl[407] vdd gnd cell_6t
Xbit_r408_c57 bl[57] br[57] wl[408] vdd gnd cell_6t
Xbit_r409_c57 bl[57] br[57] wl[409] vdd gnd cell_6t
Xbit_r410_c57 bl[57] br[57] wl[410] vdd gnd cell_6t
Xbit_r411_c57 bl[57] br[57] wl[411] vdd gnd cell_6t
Xbit_r412_c57 bl[57] br[57] wl[412] vdd gnd cell_6t
Xbit_r413_c57 bl[57] br[57] wl[413] vdd gnd cell_6t
Xbit_r414_c57 bl[57] br[57] wl[414] vdd gnd cell_6t
Xbit_r415_c57 bl[57] br[57] wl[415] vdd gnd cell_6t
Xbit_r416_c57 bl[57] br[57] wl[416] vdd gnd cell_6t
Xbit_r417_c57 bl[57] br[57] wl[417] vdd gnd cell_6t
Xbit_r418_c57 bl[57] br[57] wl[418] vdd gnd cell_6t
Xbit_r419_c57 bl[57] br[57] wl[419] vdd gnd cell_6t
Xbit_r420_c57 bl[57] br[57] wl[420] vdd gnd cell_6t
Xbit_r421_c57 bl[57] br[57] wl[421] vdd gnd cell_6t
Xbit_r422_c57 bl[57] br[57] wl[422] vdd gnd cell_6t
Xbit_r423_c57 bl[57] br[57] wl[423] vdd gnd cell_6t
Xbit_r424_c57 bl[57] br[57] wl[424] vdd gnd cell_6t
Xbit_r425_c57 bl[57] br[57] wl[425] vdd gnd cell_6t
Xbit_r426_c57 bl[57] br[57] wl[426] vdd gnd cell_6t
Xbit_r427_c57 bl[57] br[57] wl[427] vdd gnd cell_6t
Xbit_r428_c57 bl[57] br[57] wl[428] vdd gnd cell_6t
Xbit_r429_c57 bl[57] br[57] wl[429] vdd gnd cell_6t
Xbit_r430_c57 bl[57] br[57] wl[430] vdd gnd cell_6t
Xbit_r431_c57 bl[57] br[57] wl[431] vdd gnd cell_6t
Xbit_r432_c57 bl[57] br[57] wl[432] vdd gnd cell_6t
Xbit_r433_c57 bl[57] br[57] wl[433] vdd gnd cell_6t
Xbit_r434_c57 bl[57] br[57] wl[434] vdd gnd cell_6t
Xbit_r435_c57 bl[57] br[57] wl[435] vdd gnd cell_6t
Xbit_r436_c57 bl[57] br[57] wl[436] vdd gnd cell_6t
Xbit_r437_c57 bl[57] br[57] wl[437] vdd gnd cell_6t
Xbit_r438_c57 bl[57] br[57] wl[438] vdd gnd cell_6t
Xbit_r439_c57 bl[57] br[57] wl[439] vdd gnd cell_6t
Xbit_r440_c57 bl[57] br[57] wl[440] vdd gnd cell_6t
Xbit_r441_c57 bl[57] br[57] wl[441] vdd gnd cell_6t
Xbit_r442_c57 bl[57] br[57] wl[442] vdd gnd cell_6t
Xbit_r443_c57 bl[57] br[57] wl[443] vdd gnd cell_6t
Xbit_r444_c57 bl[57] br[57] wl[444] vdd gnd cell_6t
Xbit_r445_c57 bl[57] br[57] wl[445] vdd gnd cell_6t
Xbit_r446_c57 bl[57] br[57] wl[446] vdd gnd cell_6t
Xbit_r447_c57 bl[57] br[57] wl[447] vdd gnd cell_6t
Xbit_r448_c57 bl[57] br[57] wl[448] vdd gnd cell_6t
Xbit_r449_c57 bl[57] br[57] wl[449] vdd gnd cell_6t
Xbit_r450_c57 bl[57] br[57] wl[450] vdd gnd cell_6t
Xbit_r451_c57 bl[57] br[57] wl[451] vdd gnd cell_6t
Xbit_r452_c57 bl[57] br[57] wl[452] vdd gnd cell_6t
Xbit_r453_c57 bl[57] br[57] wl[453] vdd gnd cell_6t
Xbit_r454_c57 bl[57] br[57] wl[454] vdd gnd cell_6t
Xbit_r455_c57 bl[57] br[57] wl[455] vdd gnd cell_6t
Xbit_r456_c57 bl[57] br[57] wl[456] vdd gnd cell_6t
Xbit_r457_c57 bl[57] br[57] wl[457] vdd gnd cell_6t
Xbit_r458_c57 bl[57] br[57] wl[458] vdd gnd cell_6t
Xbit_r459_c57 bl[57] br[57] wl[459] vdd gnd cell_6t
Xbit_r460_c57 bl[57] br[57] wl[460] vdd gnd cell_6t
Xbit_r461_c57 bl[57] br[57] wl[461] vdd gnd cell_6t
Xbit_r462_c57 bl[57] br[57] wl[462] vdd gnd cell_6t
Xbit_r463_c57 bl[57] br[57] wl[463] vdd gnd cell_6t
Xbit_r464_c57 bl[57] br[57] wl[464] vdd gnd cell_6t
Xbit_r465_c57 bl[57] br[57] wl[465] vdd gnd cell_6t
Xbit_r466_c57 bl[57] br[57] wl[466] vdd gnd cell_6t
Xbit_r467_c57 bl[57] br[57] wl[467] vdd gnd cell_6t
Xbit_r468_c57 bl[57] br[57] wl[468] vdd gnd cell_6t
Xbit_r469_c57 bl[57] br[57] wl[469] vdd gnd cell_6t
Xbit_r470_c57 bl[57] br[57] wl[470] vdd gnd cell_6t
Xbit_r471_c57 bl[57] br[57] wl[471] vdd gnd cell_6t
Xbit_r472_c57 bl[57] br[57] wl[472] vdd gnd cell_6t
Xbit_r473_c57 bl[57] br[57] wl[473] vdd gnd cell_6t
Xbit_r474_c57 bl[57] br[57] wl[474] vdd gnd cell_6t
Xbit_r475_c57 bl[57] br[57] wl[475] vdd gnd cell_6t
Xbit_r476_c57 bl[57] br[57] wl[476] vdd gnd cell_6t
Xbit_r477_c57 bl[57] br[57] wl[477] vdd gnd cell_6t
Xbit_r478_c57 bl[57] br[57] wl[478] vdd gnd cell_6t
Xbit_r479_c57 bl[57] br[57] wl[479] vdd gnd cell_6t
Xbit_r480_c57 bl[57] br[57] wl[480] vdd gnd cell_6t
Xbit_r481_c57 bl[57] br[57] wl[481] vdd gnd cell_6t
Xbit_r482_c57 bl[57] br[57] wl[482] vdd gnd cell_6t
Xbit_r483_c57 bl[57] br[57] wl[483] vdd gnd cell_6t
Xbit_r484_c57 bl[57] br[57] wl[484] vdd gnd cell_6t
Xbit_r485_c57 bl[57] br[57] wl[485] vdd gnd cell_6t
Xbit_r486_c57 bl[57] br[57] wl[486] vdd gnd cell_6t
Xbit_r487_c57 bl[57] br[57] wl[487] vdd gnd cell_6t
Xbit_r488_c57 bl[57] br[57] wl[488] vdd gnd cell_6t
Xbit_r489_c57 bl[57] br[57] wl[489] vdd gnd cell_6t
Xbit_r490_c57 bl[57] br[57] wl[490] vdd gnd cell_6t
Xbit_r491_c57 bl[57] br[57] wl[491] vdd gnd cell_6t
Xbit_r492_c57 bl[57] br[57] wl[492] vdd gnd cell_6t
Xbit_r493_c57 bl[57] br[57] wl[493] vdd gnd cell_6t
Xbit_r494_c57 bl[57] br[57] wl[494] vdd gnd cell_6t
Xbit_r495_c57 bl[57] br[57] wl[495] vdd gnd cell_6t
Xbit_r496_c57 bl[57] br[57] wl[496] vdd gnd cell_6t
Xbit_r497_c57 bl[57] br[57] wl[497] vdd gnd cell_6t
Xbit_r498_c57 bl[57] br[57] wl[498] vdd gnd cell_6t
Xbit_r499_c57 bl[57] br[57] wl[499] vdd gnd cell_6t
Xbit_r500_c57 bl[57] br[57] wl[500] vdd gnd cell_6t
Xbit_r501_c57 bl[57] br[57] wl[501] vdd gnd cell_6t
Xbit_r502_c57 bl[57] br[57] wl[502] vdd gnd cell_6t
Xbit_r503_c57 bl[57] br[57] wl[503] vdd gnd cell_6t
Xbit_r504_c57 bl[57] br[57] wl[504] vdd gnd cell_6t
Xbit_r505_c57 bl[57] br[57] wl[505] vdd gnd cell_6t
Xbit_r506_c57 bl[57] br[57] wl[506] vdd gnd cell_6t
Xbit_r507_c57 bl[57] br[57] wl[507] vdd gnd cell_6t
Xbit_r508_c57 bl[57] br[57] wl[508] vdd gnd cell_6t
Xbit_r509_c57 bl[57] br[57] wl[509] vdd gnd cell_6t
Xbit_r510_c57 bl[57] br[57] wl[510] vdd gnd cell_6t
Xbit_r511_c57 bl[57] br[57] wl[511] vdd gnd cell_6t
Xbit_r0_c58 bl[58] br[58] wl[0] vdd gnd cell_6t
Xbit_r1_c58 bl[58] br[58] wl[1] vdd gnd cell_6t
Xbit_r2_c58 bl[58] br[58] wl[2] vdd gnd cell_6t
Xbit_r3_c58 bl[58] br[58] wl[3] vdd gnd cell_6t
Xbit_r4_c58 bl[58] br[58] wl[4] vdd gnd cell_6t
Xbit_r5_c58 bl[58] br[58] wl[5] vdd gnd cell_6t
Xbit_r6_c58 bl[58] br[58] wl[6] vdd gnd cell_6t
Xbit_r7_c58 bl[58] br[58] wl[7] vdd gnd cell_6t
Xbit_r8_c58 bl[58] br[58] wl[8] vdd gnd cell_6t
Xbit_r9_c58 bl[58] br[58] wl[9] vdd gnd cell_6t
Xbit_r10_c58 bl[58] br[58] wl[10] vdd gnd cell_6t
Xbit_r11_c58 bl[58] br[58] wl[11] vdd gnd cell_6t
Xbit_r12_c58 bl[58] br[58] wl[12] vdd gnd cell_6t
Xbit_r13_c58 bl[58] br[58] wl[13] vdd gnd cell_6t
Xbit_r14_c58 bl[58] br[58] wl[14] vdd gnd cell_6t
Xbit_r15_c58 bl[58] br[58] wl[15] vdd gnd cell_6t
Xbit_r16_c58 bl[58] br[58] wl[16] vdd gnd cell_6t
Xbit_r17_c58 bl[58] br[58] wl[17] vdd gnd cell_6t
Xbit_r18_c58 bl[58] br[58] wl[18] vdd gnd cell_6t
Xbit_r19_c58 bl[58] br[58] wl[19] vdd gnd cell_6t
Xbit_r20_c58 bl[58] br[58] wl[20] vdd gnd cell_6t
Xbit_r21_c58 bl[58] br[58] wl[21] vdd gnd cell_6t
Xbit_r22_c58 bl[58] br[58] wl[22] vdd gnd cell_6t
Xbit_r23_c58 bl[58] br[58] wl[23] vdd gnd cell_6t
Xbit_r24_c58 bl[58] br[58] wl[24] vdd gnd cell_6t
Xbit_r25_c58 bl[58] br[58] wl[25] vdd gnd cell_6t
Xbit_r26_c58 bl[58] br[58] wl[26] vdd gnd cell_6t
Xbit_r27_c58 bl[58] br[58] wl[27] vdd gnd cell_6t
Xbit_r28_c58 bl[58] br[58] wl[28] vdd gnd cell_6t
Xbit_r29_c58 bl[58] br[58] wl[29] vdd gnd cell_6t
Xbit_r30_c58 bl[58] br[58] wl[30] vdd gnd cell_6t
Xbit_r31_c58 bl[58] br[58] wl[31] vdd gnd cell_6t
Xbit_r32_c58 bl[58] br[58] wl[32] vdd gnd cell_6t
Xbit_r33_c58 bl[58] br[58] wl[33] vdd gnd cell_6t
Xbit_r34_c58 bl[58] br[58] wl[34] vdd gnd cell_6t
Xbit_r35_c58 bl[58] br[58] wl[35] vdd gnd cell_6t
Xbit_r36_c58 bl[58] br[58] wl[36] vdd gnd cell_6t
Xbit_r37_c58 bl[58] br[58] wl[37] vdd gnd cell_6t
Xbit_r38_c58 bl[58] br[58] wl[38] vdd gnd cell_6t
Xbit_r39_c58 bl[58] br[58] wl[39] vdd gnd cell_6t
Xbit_r40_c58 bl[58] br[58] wl[40] vdd gnd cell_6t
Xbit_r41_c58 bl[58] br[58] wl[41] vdd gnd cell_6t
Xbit_r42_c58 bl[58] br[58] wl[42] vdd gnd cell_6t
Xbit_r43_c58 bl[58] br[58] wl[43] vdd gnd cell_6t
Xbit_r44_c58 bl[58] br[58] wl[44] vdd gnd cell_6t
Xbit_r45_c58 bl[58] br[58] wl[45] vdd gnd cell_6t
Xbit_r46_c58 bl[58] br[58] wl[46] vdd gnd cell_6t
Xbit_r47_c58 bl[58] br[58] wl[47] vdd gnd cell_6t
Xbit_r48_c58 bl[58] br[58] wl[48] vdd gnd cell_6t
Xbit_r49_c58 bl[58] br[58] wl[49] vdd gnd cell_6t
Xbit_r50_c58 bl[58] br[58] wl[50] vdd gnd cell_6t
Xbit_r51_c58 bl[58] br[58] wl[51] vdd gnd cell_6t
Xbit_r52_c58 bl[58] br[58] wl[52] vdd gnd cell_6t
Xbit_r53_c58 bl[58] br[58] wl[53] vdd gnd cell_6t
Xbit_r54_c58 bl[58] br[58] wl[54] vdd gnd cell_6t
Xbit_r55_c58 bl[58] br[58] wl[55] vdd gnd cell_6t
Xbit_r56_c58 bl[58] br[58] wl[56] vdd gnd cell_6t
Xbit_r57_c58 bl[58] br[58] wl[57] vdd gnd cell_6t
Xbit_r58_c58 bl[58] br[58] wl[58] vdd gnd cell_6t
Xbit_r59_c58 bl[58] br[58] wl[59] vdd gnd cell_6t
Xbit_r60_c58 bl[58] br[58] wl[60] vdd gnd cell_6t
Xbit_r61_c58 bl[58] br[58] wl[61] vdd gnd cell_6t
Xbit_r62_c58 bl[58] br[58] wl[62] vdd gnd cell_6t
Xbit_r63_c58 bl[58] br[58] wl[63] vdd gnd cell_6t
Xbit_r64_c58 bl[58] br[58] wl[64] vdd gnd cell_6t
Xbit_r65_c58 bl[58] br[58] wl[65] vdd gnd cell_6t
Xbit_r66_c58 bl[58] br[58] wl[66] vdd gnd cell_6t
Xbit_r67_c58 bl[58] br[58] wl[67] vdd gnd cell_6t
Xbit_r68_c58 bl[58] br[58] wl[68] vdd gnd cell_6t
Xbit_r69_c58 bl[58] br[58] wl[69] vdd gnd cell_6t
Xbit_r70_c58 bl[58] br[58] wl[70] vdd gnd cell_6t
Xbit_r71_c58 bl[58] br[58] wl[71] vdd gnd cell_6t
Xbit_r72_c58 bl[58] br[58] wl[72] vdd gnd cell_6t
Xbit_r73_c58 bl[58] br[58] wl[73] vdd gnd cell_6t
Xbit_r74_c58 bl[58] br[58] wl[74] vdd gnd cell_6t
Xbit_r75_c58 bl[58] br[58] wl[75] vdd gnd cell_6t
Xbit_r76_c58 bl[58] br[58] wl[76] vdd gnd cell_6t
Xbit_r77_c58 bl[58] br[58] wl[77] vdd gnd cell_6t
Xbit_r78_c58 bl[58] br[58] wl[78] vdd gnd cell_6t
Xbit_r79_c58 bl[58] br[58] wl[79] vdd gnd cell_6t
Xbit_r80_c58 bl[58] br[58] wl[80] vdd gnd cell_6t
Xbit_r81_c58 bl[58] br[58] wl[81] vdd gnd cell_6t
Xbit_r82_c58 bl[58] br[58] wl[82] vdd gnd cell_6t
Xbit_r83_c58 bl[58] br[58] wl[83] vdd gnd cell_6t
Xbit_r84_c58 bl[58] br[58] wl[84] vdd gnd cell_6t
Xbit_r85_c58 bl[58] br[58] wl[85] vdd gnd cell_6t
Xbit_r86_c58 bl[58] br[58] wl[86] vdd gnd cell_6t
Xbit_r87_c58 bl[58] br[58] wl[87] vdd gnd cell_6t
Xbit_r88_c58 bl[58] br[58] wl[88] vdd gnd cell_6t
Xbit_r89_c58 bl[58] br[58] wl[89] vdd gnd cell_6t
Xbit_r90_c58 bl[58] br[58] wl[90] vdd gnd cell_6t
Xbit_r91_c58 bl[58] br[58] wl[91] vdd gnd cell_6t
Xbit_r92_c58 bl[58] br[58] wl[92] vdd gnd cell_6t
Xbit_r93_c58 bl[58] br[58] wl[93] vdd gnd cell_6t
Xbit_r94_c58 bl[58] br[58] wl[94] vdd gnd cell_6t
Xbit_r95_c58 bl[58] br[58] wl[95] vdd gnd cell_6t
Xbit_r96_c58 bl[58] br[58] wl[96] vdd gnd cell_6t
Xbit_r97_c58 bl[58] br[58] wl[97] vdd gnd cell_6t
Xbit_r98_c58 bl[58] br[58] wl[98] vdd gnd cell_6t
Xbit_r99_c58 bl[58] br[58] wl[99] vdd gnd cell_6t
Xbit_r100_c58 bl[58] br[58] wl[100] vdd gnd cell_6t
Xbit_r101_c58 bl[58] br[58] wl[101] vdd gnd cell_6t
Xbit_r102_c58 bl[58] br[58] wl[102] vdd gnd cell_6t
Xbit_r103_c58 bl[58] br[58] wl[103] vdd gnd cell_6t
Xbit_r104_c58 bl[58] br[58] wl[104] vdd gnd cell_6t
Xbit_r105_c58 bl[58] br[58] wl[105] vdd gnd cell_6t
Xbit_r106_c58 bl[58] br[58] wl[106] vdd gnd cell_6t
Xbit_r107_c58 bl[58] br[58] wl[107] vdd gnd cell_6t
Xbit_r108_c58 bl[58] br[58] wl[108] vdd gnd cell_6t
Xbit_r109_c58 bl[58] br[58] wl[109] vdd gnd cell_6t
Xbit_r110_c58 bl[58] br[58] wl[110] vdd gnd cell_6t
Xbit_r111_c58 bl[58] br[58] wl[111] vdd gnd cell_6t
Xbit_r112_c58 bl[58] br[58] wl[112] vdd gnd cell_6t
Xbit_r113_c58 bl[58] br[58] wl[113] vdd gnd cell_6t
Xbit_r114_c58 bl[58] br[58] wl[114] vdd gnd cell_6t
Xbit_r115_c58 bl[58] br[58] wl[115] vdd gnd cell_6t
Xbit_r116_c58 bl[58] br[58] wl[116] vdd gnd cell_6t
Xbit_r117_c58 bl[58] br[58] wl[117] vdd gnd cell_6t
Xbit_r118_c58 bl[58] br[58] wl[118] vdd gnd cell_6t
Xbit_r119_c58 bl[58] br[58] wl[119] vdd gnd cell_6t
Xbit_r120_c58 bl[58] br[58] wl[120] vdd gnd cell_6t
Xbit_r121_c58 bl[58] br[58] wl[121] vdd gnd cell_6t
Xbit_r122_c58 bl[58] br[58] wl[122] vdd gnd cell_6t
Xbit_r123_c58 bl[58] br[58] wl[123] vdd gnd cell_6t
Xbit_r124_c58 bl[58] br[58] wl[124] vdd gnd cell_6t
Xbit_r125_c58 bl[58] br[58] wl[125] vdd gnd cell_6t
Xbit_r126_c58 bl[58] br[58] wl[126] vdd gnd cell_6t
Xbit_r127_c58 bl[58] br[58] wl[127] vdd gnd cell_6t
Xbit_r128_c58 bl[58] br[58] wl[128] vdd gnd cell_6t
Xbit_r129_c58 bl[58] br[58] wl[129] vdd gnd cell_6t
Xbit_r130_c58 bl[58] br[58] wl[130] vdd gnd cell_6t
Xbit_r131_c58 bl[58] br[58] wl[131] vdd gnd cell_6t
Xbit_r132_c58 bl[58] br[58] wl[132] vdd gnd cell_6t
Xbit_r133_c58 bl[58] br[58] wl[133] vdd gnd cell_6t
Xbit_r134_c58 bl[58] br[58] wl[134] vdd gnd cell_6t
Xbit_r135_c58 bl[58] br[58] wl[135] vdd gnd cell_6t
Xbit_r136_c58 bl[58] br[58] wl[136] vdd gnd cell_6t
Xbit_r137_c58 bl[58] br[58] wl[137] vdd gnd cell_6t
Xbit_r138_c58 bl[58] br[58] wl[138] vdd gnd cell_6t
Xbit_r139_c58 bl[58] br[58] wl[139] vdd gnd cell_6t
Xbit_r140_c58 bl[58] br[58] wl[140] vdd gnd cell_6t
Xbit_r141_c58 bl[58] br[58] wl[141] vdd gnd cell_6t
Xbit_r142_c58 bl[58] br[58] wl[142] vdd gnd cell_6t
Xbit_r143_c58 bl[58] br[58] wl[143] vdd gnd cell_6t
Xbit_r144_c58 bl[58] br[58] wl[144] vdd gnd cell_6t
Xbit_r145_c58 bl[58] br[58] wl[145] vdd gnd cell_6t
Xbit_r146_c58 bl[58] br[58] wl[146] vdd gnd cell_6t
Xbit_r147_c58 bl[58] br[58] wl[147] vdd gnd cell_6t
Xbit_r148_c58 bl[58] br[58] wl[148] vdd gnd cell_6t
Xbit_r149_c58 bl[58] br[58] wl[149] vdd gnd cell_6t
Xbit_r150_c58 bl[58] br[58] wl[150] vdd gnd cell_6t
Xbit_r151_c58 bl[58] br[58] wl[151] vdd gnd cell_6t
Xbit_r152_c58 bl[58] br[58] wl[152] vdd gnd cell_6t
Xbit_r153_c58 bl[58] br[58] wl[153] vdd gnd cell_6t
Xbit_r154_c58 bl[58] br[58] wl[154] vdd gnd cell_6t
Xbit_r155_c58 bl[58] br[58] wl[155] vdd gnd cell_6t
Xbit_r156_c58 bl[58] br[58] wl[156] vdd gnd cell_6t
Xbit_r157_c58 bl[58] br[58] wl[157] vdd gnd cell_6t
Xbit_r158_c58 bl[58] br[58] wl[158] vdd gnd cell_6t
Xbit_r159_c58 bl[58] br[58] wl[159] vdd gnd cell_6t
Xbit_r160_c58 bl[58] br[58] wl[160] vdd gnd cell_6t
Xbit_r161_c58 bl[58] br[58] wl[161] vdd gnd cell_6t
Xbit_r162_c58 bl[58] br[58] wl[162] vdd gnd cell_6t
Xbit_r163_c58 bl[58] br[58] wl[163] vdd gnd cell_6t
Xbit_r164_c58 bl[58] br[58] wl[164] vdd gnd cell_6t
Xbit_r165_c58 bl[58] br[58] wl[165] vdd gnd cell_6t
Xbit_r166_c58 bl[58] br[58] wl[166] vdd gnd cell_6t
Xbit_r167_c58 bl[58] br[58] wl[167] vdd gnd cell_6t
Xbit_r168_c58 bl[58] br[58] wl[168] vdd gnd cell_6t
Xbit_r169_c58 bl[58] br[58] wl[169] vdd gnd cell_6t
Xbit_r170_c58 bl[58] br[58] wl[170] vdd gnd cell_6t
Xbit_r171_c58 bl[58] br[58] wl[171] vdd gnd cell_6t
Xbit_r172_c58 bl[58] br[58] wl[172] vdd gnd cell_6t
Xbit_r173_c58 bl[58] br[58] wl[173] vdd gnd cell_6t
Xbit_r174_c58 bl[58] br[58] wl[174] vdd gnd cell_6t
Xbit_r175_c58 bl[58] br[58] wl[175] vdd gnd cell_6t
Xbit_r176_c58 bl[58] br[58] wl[176] vdd gnd cell_6t
Xbit_r177_c58 bl[58] br[58] wl[177] vdd gnd cell_6t
Xbit_r178_c58 bl[58] br[58] wl[178] vdd gnd cell_6t
Xbit_r179_c58 bl[58] br[58] wl[179] vdd gnd cell_6t
Xbit_r180_c58 bl[58] br[58] wl[180] vdd gnd cell_6t
Xbit_r181_c58 bl[58] br[58] wl[181] vdd gnd cell_6t
Xbit_r182_c58 bl[58] br[58] wl[182] vdd gnd cell_6t
Xbit_r183_c58 bl[58] br[58] wl[183] vdd gnd cell_6t
Xbit_r184_c58 bl[58] br[58] wl[184] vdd gnd cell_6t
Xbit_r185_c58 bl[58] br[58] wl[185] vdd gnd cell_6t
Xbit_r186_c58 bl[58] br[58] wl[186] vdd gnd cell_6t
Xbit_r187_c58 bl[58] br[58] wl[187] vdd gnd cell_6t
Xbit_r188_c58 bl[58] br[58] wl[188] vdd gnd cell_6t
Xbit_r189_c58 bl[58] br[58] wl[189] vdd gnd cell_6t
Xbit_r190_c58 bl[58] br[58] wl[190] vdd gnd cell_6t
Xbit_r191_c58 bl[58] br[58] wl[191] vdd gnd cell_6t
Xbit_r192_c58 bl[58] br[58] wl[192] vdd gnd cell_6t
Xbit_r193_c58 bl[58] br[58] wl[193] vdd gnd cell_6t
Xbit_r194_c58 bl[58] br[58] wl[194] vdd gnd cell_6t
Xbit_r195_c58 bl[58] br[58] wl[195] vdd gnd cell_6t
Xbit_r196_c58 bl[58] br[58] wl[196] vdd gnd cell_6t
Xbit_r197_c58 bl[58] br[58] wl[197] vdd gnd cell_6t
Xbit_r198_c58 bl[58] br[58] wl[198] vdd gnd cell_6t
Xbit_r199_c58 bl[58] br[58] wl[199] vdd gnd cell_6t
Xbit_r200_c58 bl[58] br[58] wl[200] vdd gnd cell_6t
Xbit_r201_c58 bl[58] br[58] wl[201] vdd gnd cell_6t
Xbit_r202_c58 bl[58] br[58] wl[202] vdd gnd cell_6t
Xbit_r203_c58 bl[58] br[58] wl[203] vdd gnd cell_6t
Xbit_r204_c58 bl[58] br[58] wl[204] vdd gnd cell_6t
Xbit_r205_c58 bl[58] br[58] wl[205] vdd gnd cell_6t
Xbit_r206_c58 bl[58] br[58] wl[206] vdd gnd cell_6t
Xbit_r207_c58 bl[58] br[58] wl[207] vdd gnd cell_6t
Xbit_r208_c58 bl[58] br[58] wl[208] vdd gnd cell_6t
Xbit_r209_c58 bl[58] br[58] wl[209] vdd gnd cell_6t
Xbit_r210_c58 bl[58] br[58] wl[210] vdd gnd cell_6t
Xbit_r211_c58 bl[58] br[58] wl[211] vdd gnd cell_6t
Xbit_r212_c58 bl[58] br[58] wl[212] vdd gnd cell_6t
Xbit_r213_c58 bl[58] br[58] wl[213] vdd gnd cell_6t
Xbit_r214_c58 bl[58] br[58] wl[214] vdd gnd cell_6t
Xbit_r215_c58 bl[58] br[58] wl[215] vdd gnd cell_6t
Xbit_r216_c58 bl[58] br[58] wl[216] vdd gnd cell_6t
Xbit_r217_c58 bl[58] br[58] wl[217] vdd gnd cell_6t
Xbit_r218_c58 bl[58] br[58] wl[218] vdd gnd cell_6t
Xbit_r219_c58 bl[58] br[58] wl[219] vdd gnd cell_6t
Xbit_r220_c58 bl[58] br[58] wl[220] vdd gnd cell_6t
Xbit_r221_c58 bl[58] br[58] wl[221] vdd gnd cell_6t
Xbit_r222_c58 bl[58] br[58] wl[222] vdd gnd cell_6t
Xbit_r223_c58 bl[58] br[58] wl[223] vdd gnd cell_6t
Xbit_r224_c58 bl[58] br[58] wl[224] vdd gnd cell_6t
Xbit_r225_c58 bl[58] br[58] wl[225] vdd gnd cell_6t
Xbit_r226_c58 bl[58] br[58] wl[226] vdd gnd cell_6t
Xbit_r227_c58 bl[58] br[58] wl[227] vdd gnd cell_6t
Xbit_r228_c58 bl[58] br[58] wl[228] vdd gnd cell_6t
Xbit_r229_c58 bl[58] br[58] wl[229] vdd gnd cell_6t
Xbit_r230_c58 bl[58] br[58] wl[230] vdd gnd cell_6t
Xbit_r231_c58 bl[58] br[58] wl[231] vdd gnd cell_6t
Xbit_r232_c58 bl[58] br[58] wl[232] vdd gnd cell_6t
Xbit_r233_c58 bl[58] br[58] wl[233] vdd gnd cell_6t
Xbit_r234_c58 bl[58] br[58] wl[234] vdd gnd cell_6t
Xbit_r235_c58 bl[58] br[58] wl[235] vdd gnd cell_6t
Xbit_r236_c58 bl[58] br[58] wl[236] vdd gnd cell_6t
Xbit_r237_c58 bl[58] br[58] wl[237] vdd gnd cell_6t
Xbit_r238_c58 bl[58] br[58] wl[238] vdd gnd cell_6t
Xbit_r239_c58 bl[58] br[58] wl[239] vdd gnd cell_6t
Xbit_r240_c58 bl[58] br[58] wl[240] vdd gnd cell_6t
Xbit_r241_c58 bl[58] br[58] wl[241] vdd gnd cell_6t
Xbit_r242_c58 bl[58] br[58] wl[242] vdd gnd cell_6t
Xbit_r243_c58 bl[58] br[58] wl[243] vdd gnd cell_6t
Xbit_r244_c58 bl[58] br[58] wl[244] vdd gnd cell_6t
Xbit_r245_c58 bl[58] br[58] wl[245] vdd gnd cell_6t
Xbit_r246_c58 bl[58] br[58] wl[246] vdd gnd cell_6t
Xbit_r247_c58 bl[58] br[58] wl[247] vdd gnd cell_6t
Xbit_r248_c58 bl[58] br[58] wl[248] vdd gnd cell_6t
Xbit_r249_c58 bl[58] br[58] wl[249] vdd gnd cell_6t
Xbit_r250_c58 bl[58] br[58] wl[250] vdd gnd cell_6t
Xbit_r251_c58 bl[58] br[58] wl[251] vdd gnd cell_6t
Xbit_r252_c58 bl[58] br[58] wl[252] vdd gnd cell_6t
Xbit_r253_c58 bl[58] br[58] wl[253] vdd gnd cell_6t
Xbit_r254_c58 bl[58] br[58] wl[254] vdd gnd cell_6t
Xbit_r255_c58 bl[58] br[58] wl[255] vdd gnd cell_6t
Xbit_r256_c58 bl[58] br[58] wl[256] vdd gnd cell_6t
Xbit_r257_c58 bl[58] br[58] wl[257] vdd gnd cell_6t
Xbit_r258_c58 bl[58] br[58] wl[258] vdd gnd cell_6t
Xbit_r259_c58 bl[58] br[58] wl[259] vdd gnd cell_6t
Xbit_r260_c58 bl[58] br[58] wl[260] vdd gnd cell_6t
Xbit_r261_c58 bl[58] br[58] wl[261] vdd gnd cell_6t
Xbit_r262_c58 bl[58] br[58] wl[262] vdd gnd cell_6t
Xbit_r263_c58 bl[58] br[58] wl[263] vdd gnd cell_6t
Xbit_r264_c58 bl[58] br[58] wl[264] vdd gnd cell_6t
Xbit_r265_c58 bl[58] br[58] wl[265] vdd gnd cell_6t
Xbit_r266_c58 bl[58] br[58] wl[266] vdd gnd cell_6t
Xbit_r267_c58 bl[58] br[58] wl[267] vdd gnd cell_6t
Xbit_r268_c58 bl[58] br[58] wl[268] vdd gnd cell_6t
Xbit_r269_c58 bl[58] br[58] wl[269] vdd gnd cell_6t
Xbit_r270_c58 bl[58] br[58] wl[270] vdd gnd cell_6t
Xbit_r271_c58 bl[58] br[58] wl[271] vdd gnd cell_6t
Xbit_r272_c58 bl[58] br[58] wl[272] vdd gnd cell_6t
Xbit_r273_c58 bl[58] br[58] wl[273] vdd gnd cell_6t
Xbit_r274_c58 bl[58] br[58] wl[274] vdd gnd cell_6t
Xbit_r275_c58 bl[58] br[58] wl[275] vdd gnd cell_6t
Xbit_r276_c58 bl[58] br[58] wl[276] vdd gnd cell_6t
Xbit_r277_c58 bl[58] br[58] wl[277] vdd gnd cell_6t
Xbit_r278_c58 bl[58] br[58] wl[278] vdd gnd cell_6t
Xbit_r279_c58 bl[58] br[58] wl[279] vdd gnd cell_6t
Xbit_r280_c58 bl[58] br[58] wl[280] vdd gnd cell_6t
Xbit_r281_c58 bl[58] br[58] wl[281] vdd gnd cell_6t
Xbit_r282_c58 bl[58] br[58] wl[282] vdd gnd cell_6t
Xbit_r283_c58 bl[58] br[58] wl[283] vdd gnd cell_6t
Xbit_r284_c58 bl[58] br[58] wl[284] vdd gnd cell_6t
Xbit_r285_c58 bl[58] br[58] wl[285] vdd gnd cell_6t
Xbit_r286_c58 bl[58] br[58] wl[286] vdd gnd cell_6t
Xbit_r287_c58 bl[58] br[58] wl[287] vdd gnd cell_6t
Xbit_r288_c58 bl[58] br[58] wl[288] vdd gnd cell_6t
Xbit_r289_c58 bl[58] br[58] wl[289] vdd gnd cell_6t
Xbit_r290_c58 bl[58] br[58] wl[290] vdd gnd cell_6t
Xbit_r291_c58 bl[58] br[58] wl[291] vdd gnd cell_6t
Xbit_r292_c58 bl[58] br[58] wl[292] vdd gnd cell_6t
Xbit_r293_c58 bl[58] br[58] wl[293] vdd gnd cell_6t
Xbit_r294_c58 bl[58] br[58] wl[294] vdd gnd cell_6t
Xbit_r295_c58 bl[58] br[58] wl[295] vdd gnd cell_6t
Xbit_r296_c58 bl[58] br[58] wl[296] vdd gnd cell_6t
Xbit_r297_c58 bl[58] br[58] wl[297] vdd gnd cell_6t
Xbit_r298_c58 bl[58] br[58] wl[298] vdd gnd cell_6t
Xbit_r299_c58 bl[58] br[58] wl[299] vdd gnd cell_6t
Xbit_r300_c58 bl[58] br[58] wl[300] vdd gnd cell_6t
Xbit_r301_c58 bl[58] br[58] wl[301] vdd gnd cell_6t
Xbit_r302_c58 bl[58] br[58] wl[302] vdd gnd cell_6t
Xbit_r303_c58 bl[58] br[58] wl[303] vdd gnd cell_6t
Xbit_r304_c58 bl[58] br[58] wl[304] vdd gnd cell_6t
Xbit_r305_c58 bl[58] br[58] wl[305] vdd gnd cell_6t
Xbit_r306_c58 bl[58] br[58] wl[306] vdd gnd cell_6t
Xbit_r307_c58 bl[58] br[58] wl[307] vdd gnd cell_6t
Xbit_r308_c58 bl[58] br[58] wl[308] vdd gnd cell_6t
Xbit_r309_c58 bl[58] br[58] wl[309] vdd gnd cell_6t
Xbit_r310_c58 bl[58] br[58] wl[310] vdd gnd cell_6t
Xbit_r311_c58 bl[58] br[58] wl[311] vdd gnd cell_6t
Xbit_r312_c58 bl[58] br[58] wl[312] vdd gnd cell_6t
Xbit_r313_c58 bl[58] br[58] wl[313] vdd gnd cell_6t
Xbit_r314_c58 bl[58] br[58] wl[314] vdd gnd cell_6t
Xbit_r315_c58 bl[58] br[58] wl[315] vdd gnd cell_6t
Xbit_r316_c58 bl[58] br[58] wl[316] vdd gnd cell_6t
Xbit_r317_c58 bl[58] br[58] wl[317] vdd gnd cell_6t
Xbit_r318_c58 bl[58] br[58] wl[318] vdd gnd cell_6t
Xbit_r319_c58 bl[58] br[58] wl[319] vdd gnd cell_6t
Xbit_r320_c58 bl[58] br[58] wl[320] vdd gnd cell_6t
Xbit_r321_c58 bl[58] br[58] wl[321] vdd gnd cell_6t
Xbit_r322_c58 bl[58] br[58] wl[322] vdd gnd cell_6t
Xbit_r323_c58 bl[58] br[58] wl[323] vdd gnd cell_6t
Xbit_r324_c58 bl[58] br[58] wl[324] vdd gnd cell_6t
Xbit_r325_c58 bl[58] br[58] wl[325] vdd gnd cell_6t
Xbit_r326_c58 bl[58] br[58] wl[326] vdd gnd cell_6t
Xbit_r327_c58 bl[58] br[58] wl[327] vdd gnd cell_6t
Xbit_r328_c58 bl[58] br[58] wl[328] vdd gnd cell_6t
Xbit_r329_c58 bl[58] br[58] wl[329] vdd gnd cell_6t
Xbit_r330_c58 bl[58] br[58] wl[330] vdd gnd cell_6t
Xbit_r331_c58 bl[58] br[58] wl[331] vdd gnd cell_6t
Xbit_r332_c58 bl[58] br[58] wl[332] vdd gnd cell_6t
Xbit_r333_c58 bl[58] br[58] wl[333] vdd gnd cell_6t
Xbit_r334_c58 bl[58] br[58] wl[334] vdd gnd cell_6t
Xbit_r335_c58 bl[58] br[58] wl[335] vdd gnd cell_6t
Xbit_r336_c58 bl[58] br[58] wl[336] vdd gnd cell_6t
Xbit_r337_c58 bl[58] br[58] wl[337] vdd gnd cell_6t
Xbit_r338_c58 bl[58] br[58] wl[338] vdd gnd cell_6t
Xbit_r339_c58 bl[58] br[58] wl[339] vdd gnd cell_6t
Xbit_r340_c58 bl[58] br[58] wl[340] vdd gnd cell_6t
Xbit_r341_c58 bl[58] br[58] wl[341] vdd gnd cell_6t
Xbit_r342_c58 bl[58] br[58] wl[342] vdd gnd cell_6t
Xbit_r343_c58 bl[58] br[58] wl[343] vdd gnd cell_6t
Xbit_r344_c58 bl[58] br[58] wl[344] vdd gnd cell_6t
Xbit_r345_c58 bl[58] br[58] wl[345] vdd gnd cell_6t
Xbit_r346_c58 bl[58] br[58] wl[346] vdd gnd cell_6t
Xbit_r347_c58 bl[58] br[58] wl[347] vdd gnd cell_6t
Xbit_r348_c58 bl[58] br[58] wl[348] vdd gnd cell_6t
Xbit_r349_c58 bl[58] br[58] wl[349] vdd gnd cell_6t
Xbit_r350_c58 bl[58] br[58] wl[350] vdd gnd cell_6t
Xbit_r351_c58 bl[58] br[58] wl[351] vdd gnd cell_6t
Xbit_r352_c58 bl[58] br[58] wl[352] vdd gnd cell_6t
Xbit_r353_c58 bl[58] br[58] wl[353] vdd gnd cell_6t
Xbit_r354_c58 bl[58] br[58] wl[354] vdd gnd cell_6t
Xbit_r355_c58 bl[58] br[58] wl[355] vdd gnd cell_6t
Xbit_r356_c58 bl[58] br[58] wl[356] vdd gnd cell_6t
Xbit_r357_c58 bl[58] br[58] wl[357] vdd gnd cell_6t
Xbit_r358_c58 bl[58] br[58] wl[358] vdd gnd cell_6t
Xbit_r359_c58 bl[58] br[58] wl[359] vdd gnd cell_6t
Xbit_r360_c58 bl[58] br[58] wl[360] vdd gnd cell_6t
Xbit_r361_c58 bl[58] br[58] wl[361] vdd gnd cell_6t
Xbit_r362_c58 bl[58] br[58] wl[362] vdd gnd cell_6t
Xbit_r363_c58 bl[58] br[58] wl[363] vdd gnd cell_6t
Xbit_r364_c58 bl[58] br[58] wl[364] vdd gnd cell_6t
Xbit_r365_c58 bl[58] br[58] wl[365] vdd gnd cell_6t
Xbit_r366_c58 bl[58] br[58] wl[366] vdd gnd cell_6t
Xbit_r367_c58 bl[58] br[58] wl[367] vdd gnd cell_6t
Xbit_r368_c58 bl[58] br[58] wl[368] vdd gnd cell_6t
Xbit_r369_c58 bl[58] br[58] wl[369] vdd gnd cell_6t
Xbit_r370_c58 bl[58] br[58] wl[370] vdd gnd cell_6t
Xbit_r371_c58 bl[58] br[58] wl[371] vdd gnd cell_6t
Xbit_r372_c58 bl[58] br[58] wl[372] vdd gnd cell_6t
Xbit_r373_c58 bl[58] br[58] wl[373] vdd gnd cell_6t
Xbit_r374_c58 bl[58] br[58] wl[374] vdd gnd cell_6t
Xbit_r375_c58 bl[58] br[58] wl[375] vdd gnd cell_6t
Xbit_r376_c58 bl[58] br[58] wl[376] vdd gnd cell_6t
Xbit_r377_c58 bl[58] br[58] wl[377] vdd gnd cell_6t
Xbit_r378_c58 bl[58] br[58] wl[378] vdd gnd cell_6t
Xbit_r379_c58 bl[58] br[58] wl[379] vdd gnd cell_6t
Xbit_r380_c58 bl[58] br[58] wl[380] vdd gnd cell_6t
Xbit_r381_c58 bl[58] br[58] wl[381] vdd gnd cell_6t
Xbit_r382_c58 bl[58] br[58] wl[382] vdd gnd cell_6t
Xbit_r383_c58 bl[58] br[58] wl[383] vdd gnd cell_6t
Xbit_r384_c58 bl[58] br[58] wl[384] vdd gnd cell_6t
Xbit_r385_c58 bl[58] br[58] wl[385] vdd gnd cell_6t
Xbit_r386_c58 bl[58] br[58] wl[386] vdd gnd cell_6t
Xbit_r387_c58 bl[58] br[58] wl[387] vdd gnd cell_6t
Xbit_r388_c58 bl[58] br[58] wl[388] vdd gnd cell_6t
Xbit_r389_c58 bl[58] br[58] wl[389] vdd gnd cell_6t
Xbit_r390_c58 bl[58] br[58] wl[390] vdd gnd cell_6t
Xbit_r391_c58 bl[58] br[58] wl[391] vdd gnd cell_6t
Xbit_r392_c58 bl[58] br[58] wl[392] vdd gnd cell_6t
Xbit_r393_c58 bl[58] br[58] wl[393] vdd gnd cell_6t
Xbit_r394_c58 bl[58] br[58] wl[394] vdd gnd cell_6t
Xbit_r395_c58 bl[58] br[58] wl[395] vdd gnd cell_6t
Xbit_r396_c58 bl[58] br[58] wl[396] vdd gnd cell_6t
Xbit_r397_c58 bl[58] br[58] wl[397] vdd gnd cell_6t
Xbit_r398_c58 bl[58] br[58] wl[398] vdd gnd cell_6t
Xbit_r399_c58 bl[58] br[58] wl[399] vdd gnd cell_6t
Xbit_r400_c58 bl[58] br[58] wl[400] vdd gnd cell_6t
Xbit_r401_c58 bl[58] br[58] wl[401] vdd gnd cell_6t
Xbit_r402_c58 bl[58] br[58] wl[402] vdd gnd cell_6t
Xbit_r403_c58 bl[58] br[58] wl[403] vdd gnd cell_6t
Xbit_r404_c58 bl[58] br[58] wl[404] vdd gnd cell_6t
Xbit_r405_c58 bl[58] br[58] wl[405] vdd gnd cell_6t
Xbit_r406_c58 bl[58] br[58] wl[406] vdd gnd cell_6t
Xbit_r407_c58 bl[58] br[58] wl[407] vdd gnd cell_6t
Xbit_r408_c58 bl[58] br[58] wl[408] vdd gnd cell_6t
Xbit_r409_c58 bl[58] br[58] wl[409] vdd gnd cell_6t
Xbit_r410_c58 bl[58] br[58] wl[410] vdd gnd cell_6t
Xbit_r411_c58 bl[58] br[58] wl[411] vdd gnd cell_6t
Xbit_r412_c58 bl[58] br[58] wl[412] vdd gnd cell_6t
Xbit_r413_c58 bl[58] br[58] wl[413] vdd gnd cell_6t
Xbit_r414_c58 bl[58] br[58] wl[414] vdd gnd cell_6t
Xbit_r415_c58 bl[58] br[58] wl[415] vdd gnd cell_6t
Xbit_r416_c58 bl[58] br[58] wl[416] vdd gnd cell_6t
Xbit_r417_c58 bl[58] br[58] wl[417] vdd gnd cell_6t
Xbit_r418_c58 bl[58] br[58] wl[418] vdd gnd cell_6t
Xbit_r419_c58 bl[58] br[58] wl[419] vdd gnd cell_6t
Xbit_r420_c58 bl[58] br[58] wl[420] vdd gnd cell_6t
Xbit_r421_c58 bl[58] br[58] wl[421] vdd gnd cell_6t
Xbit_r422_c58 bl[58] br[58] wl[422] vdd gnd cell_6t
Xbit_r423_c58 bl[58] br[58] wl[423] vdd gnd cell_6t
Xbit_r424_c58 bl[58] br[58] wl[424] vdd gnd cell_6t
Xbit_r425_c58 bl[58] br[58] wl[425] vdd gnd cell_6t
Xbit_r426_c58 bl[58] br[58] wl[426] vdd gnd cell_6t
Xbit_r427_c58 bl[58] br[58] wl[427] vdd gnd cell_6t
Xbit_r428_c58 bl[58] br[58] wl[428] vdd gnd cell_6t
Xbit_r429_c58 bl[58] br[58] wl[429] vdd gnd cell_6t
Xbit_r430_c58 bl[58] br[58] wl[430] vdd gnd cell_6t
Xbit_r431_c58 bl[58] br[58] wl[431] vdd gnd cell_6t
Xbit_r432_c58 bl[58] br[58] wl[432] vdd gnd cell_6t
Xbit_r433_c58 bl[58] br[58] wl[433] vdd gnd cell_6t
Xbit_r434_c58 bl[58] br[58] wl[434] vdd gnd cell_6t
Xbit_r435_c58 bl[58] br[58] wl[435] vdd gnd cell_6t
Xbit_r436_c58 bl[58] br[58] wl[436] vdd gnd cell_6t
Xbit_r437_c58 bl[58] br[58] wl[437] vdd gnd cell_6t
Xbit_r438_c58 bl[58] br[58] wl[438] vdd gnd cell_6t
Xbit_r439_c58 bl[58] br[58] wl[439] vdd gnd cell_6t
Xbit_r440_c58 bl[58] br[58] wl[440] vdd gnd cell_6t
Xbit_r441_c58 bl[58] br[58] wl[441] vdd gnd cell_6t
Xbit_r442_c58 bl[58] br[58] wl[442] vdd gnd cell_6t
Xbit_r443_c58 bl[58] br[58] wl[443] vdd gnd cell_6t
Xbit_r444_c58 bl[58] br[58] wl[444] vdd gnd cell_6t
Xbit_r445_c58 bl[58] br[58] wl[445] vdd gnd cell_6t
Xbit_r446_c58 bl[58] br[58] wl[446] vdd gnd cell_6t
Xbit_r447_c58 bl[58] br[58] wl[447] vdd gnd cell_6t
Xbit_r448_c58 bl[58] br[58] wl[448] vdd gnd cell_6t
Xbit_r449_c58 bl[58] br[58] wl[449] vdd gnd cell_6t
Xbit_r450_c58 bl[58] br[58] wl[450] vdd gnd cell_6t
Xbit_r451_c58 bl[58] br[58] wl[451] vdd gnd cell_6t
Xbit_r452_c58 bl[58] br[58] wl[452] vdd gnd cell_6t
Xbit_r453_c58 bl[58] br[58] wl[453] vdd gnd cell_6t
Xbit_r454_c58 bl[58] br[58] wl[454] vdd gnd cell_6t
Xbit_r455_c58 bl[58] br[58] wl[455] vdd gnd cell_6t
Xbit_r456_c58 bl[58] br[58] wl[456] vdd gnd cell_6t
Xbit_r457_c58 bl[58] br[58] wl[457] vdd gnd cell_6t
Xbit_r458_c58 bl[58] br[58] wl[458] vdd gnd cell_6t
Xbit_r459_c58 bl[58] br[58] wl[459] vdd gnd cell_6t
Xbit_r460_c58 bl[58] br[58] wl[460] vdd gnd cell_6t
Xbit_r461_c58 bl[58] br[58] wl[461] vdd gnd cell_6t
Xbit_r462_c58 bl[58] br[58] wl[462] vdd gnd cell_6t
Xbit_r463_c58 bl[58] br[58] wl[463] vdd gnd cell_6t
Xbit_r464_c58 bl[58] br[58] wl[464] vdd gnd cell_6t
Xbit_r465_c58 bl[58] br[58] wl[465] vdd gnd cell_6t
Xbit_r466_c58 bl[58] br[58] wl[466] vdd gnd cell_6t
Xbit_r467_c58 bl[58] br[58] wl[467] vdd gnd cell_6t
Xbit_r468_c58 bl[58] br[58] wl[468] vdd gnd cell_6t
Xbit_r469_c58 bl[58] br[58] wl[469] vdd gnd cell_6t
Xbit_r470_c58 bl[58] br[58] wl[470] vdd gnd cell_6t
Xbit_r471_c58 bl[58] br[58] wl[471] vdd gnd cell_6t
Xbit_r472_c58 bl[58] br[58] wl[472] vdd gnd cell_6t
Xbit_r473_c58 bl[58] br[58] wl[473] vdd gnd cell_6t
Xbit_r474_c58 bl[58] br[58] wl[474] vdd gnd cell_6t
Xbit_r475_c58 bl[58] br[58] wl[475] vdd gnd cell_6t
Xbit_r476_c58 bl[58] br[58] wl[476] vdd gnd cell_6t
Xbit_r477_c58 bl[58] br[58] wl[477] vdd gnd cell_6t
Xbit_r478_c58 bl[58] br[58] wl[478] vdd gnd cell_6t
Xbit_r479_c58 bl[58] br[58] wl[479] vdd gnd cell_6t
Xbit_r480_c58 bl[58] br[58] wl[480] vdd gnd cell_6t
Xbit_r481_c58 bl[58] br[58] wl[481] vdd gnd cell_6t
Xbit_r482_c58 bl[58] br[58] wl[482] vdd gnd cell_6t
Xbit_r483_c58 bl[58] br[58] wl[483] vdd gnd cell_6t
Xbit_r484_c58 bl[58] br[58] wl[484] vdd gnd cell_6t
Xbit_r485_c58 bl[58] br[58] wl[485] vdd gnd cell_6t
Xbit_r486_c58 bl[58] br[58] wl[486] vdd gnd cell_6t
Xbit_r487_c58 bl[58] br[58] wl[487] vdd gnd cell_6t
Xbit_r488_c58 bl[58] br[58] wl[488] vdd gnd cell_6t
Xbit_r489_c58 bl[58] br[58] wl[489] vdd gnd cell_6t
Xbit_r490_c58 bl[58] br[58] wl[490] vdd gnd cell_6t
Xbit_r491_c58 bl[58] br[58] wl[491] vdd gnd cell_6t
Xbit_r492_c58 bl[58] br[58] wl[492] vdd gnd cell_6t
Xbit_r493_c58 bl[58] br[58] wl[493] vdd gnd cell_6t
Xbit_r494_c58 bl[58] br[58] wl[494] vdd gnd cell_6t
Xbit_r495_c58 bl[58] br[58] wl[495] vdd gnd cell_6t
Xbit_r496_c58 bl[58] br[58] wl[496] vdd gnd cell_6t
Xbit_r497_c58 bl[58] br[58] wl[497] vdd gnd cell_6t
Xbit_r498_c58 bl[58] br[58] wl[498] vdd gnd cell_6t
Xbit_r499_c58 bl[58] br[58] wl[499] vdd gnd cell_6t
Xbit_r500_c58 bl[58] br[58] wl[500] vdd gnd cell_6t
Xbit_r501_c58 bl[58] br[58] wl[501] vdd gnd cell_6t
Xbit_r502_c58 bl[58] br[58] wl[502] vdd gnd cell_6t
Xbit_r503_c58 bl[58] br[58] wl[503] vdd gnd cell_6t
Xbit_r504_c58 bl[58] br[58] wl[504] vdd gnd cell_6t
Xbit_r505_c58 bl[58] br[58] wl[505] vdd gnd cell_6t
Xbit_r506_c58 bl[58] br[58] wl[506] vdd gnd cell_6t
Xbit_r507_c58 bl[58] br[58] wl[507] vdd gnd cell_6t
Xbit_r508_c58 bl[58] br[58] wl[508] vdd gnd cell_6t
Xbit_r509_c58 bl[58] br[58] wl[509] vdd gnd cell_6t
Xbit_r510_c58 bl[58] br[58] wl[510] vdd gnd cell_6t
Xbit_r511_c58 bl[58] br[58] wl[511] vdd gnd cell_6t
Xbit_r0_c59 bl[59] br[59] wl[0] vdd gnd cell_6t
Xbit_r1_c59 bl[59] br[59] wl[1] vdd gnd cell_6t
Xbit_r2_c59 bl[59] br[59] wl[2] vdd gnd cell_6t
Xbit_r3_c59 bl[59] br[59] wl[3] vdd gnd cell_6t
Xbit_r4_c59 bl[59] br[59] wl[4] vdd gnd cell_6t
Xbit_r5_c59 bl[59] br[59] wl[5] vdd gnd cell_6t
Xbit_r6_c59 bl[59] br[59] wl[6] vdd gnd cell_6t
Xbit_r7_c59 bl[59] br[59] wl[7] vdd gnd cell_6t
Xbit_r8_c59 bl[59] br[59] wl[8] vdd gnd cell_6t
Xbit_r9_c59 bl[59] br[59] wl[9] vdd gnd cell_6t
Xbit_r10_c59 bl[59] br[59] wl[10] vdd gnd cell_6t
Xbit_r11_c59 bl[59] br[59] wl[11] vdd gnd cell_6t
Xbit_r12_c59 bl[59] br[59] wl[12] vdd gnd cell_6t
Xbit_r13_c59 bl[59] br[59] wl[13] vdd gnd cell_6t
Xbit_r14_c59 bl[59] br[59] wl[14] vdd gnd cell_6t
Xbit_r15_c59 bl[59] br[59] wl[15] vdd gnd cell_6t
Xbit_r16_c59 bl[59] br[59] wl[16] vdd gnd cell_6t
Xbit_r17_c59 bl[59] br[59] wl[17] vdd gnd cell_6t
Xbit_r18_c59 bl[59] br[59] wl[18] vdd gnd cell_6t
Xbit_r19_c59 bl[59] br[59] wl[19] vdd gnd cell_6t
Xbit_r20_c59 bl[59] br[59] wl[20] vdd gnd cell_6t
Xbit_r21_c59 bl[59] br[59] wl[21] vdd gnd cell_6t
Xbit_r22_c59 bl[59] br[59] wl[22] vdd gnd cell_6t
Xbit_r23_c59 bl[59] br[59] wl[23] vdd gnd cell_6t
Xbit_r24_c59 bl[59] br[59] wl[24] vdd gnd cell_6t
Xbit_r25_c59 bl[59] br[59] wl[25] vdd gnd cell_6t
Xbit_r26_c59 bl[59] br[59] wl[26] vdd gnd cell_6t
Xbit_r27_c59 bl[59] br[59] wl[27] vdd gnd cell_6t
Xbit_r28_c59 bl[59] br[59] wl[28] vdd gnd cell_6t
Xbit_r29_c59 bl[59] br[59] wl[29] vdd gnd cell_6t
Xbit_r30_c59 bl[59] br[59] wl[30] vdd gnd cell_6t
Xbit_r31_c59 bl[59] br[59] wl[31] vdd gnd cell_6t
Xbit_r32_c59 bl[59] br[59] wl[32] vdd gnd cell_6t
Xbit_r33_c59 bl[59] br[59] wl[33] vdd gnd cell_6t
Xbit_r34_c59 bl[59] br[59] wl[34] vdd gnd cell_6t
Xbit_r35_c59 bl[59] br[59] wl[35] vdd gnd cell_6t
Xbit_r36_c59 bl[59] br[59] wl[36] vdd gnd cell_6t
Xbit_r37_c59 bl[59] br[59] wl[37] vdd gnd cell_6t
Xbit_r38_c59 bl[59] br[59] wl[38] vdd gnd cell_6t
Xbit_r39_c59 bl[59] br[59] wl[39] vdd gnd cell_6t
Xbit_r40_c59 bl[59] br[59] wl[40] vdd gnd cell_6t
Xbit_r41_c59 bl[59] br[59] wl[41] vdd gnd cell_6t
Xbit_r42_c59 bl[59] br[59] wl[42] vdd gnd cell_6t
Xbit_r43_c59 bl[59] br[59] wl[43] vdd gnd cell_6t
Xbit_r44_c59 bl[59] br[59] wl[44] vdd gnd cell_6t
Xbit_r45_c59 bl[59] br[59] wl[45] vdd gnd cell_6t
Xbit_r46_c59 bl[59] br[59] wl[46] vdd gnd cell_6t
Xbit_r47_c59 bl[59] br[59] wl[47] vdd gnd cell_6t
Xbit_r48_c59 bl[59] br[59] wl[48] vdd gnd cell_6t
Xbit_r49_c59 bl[59] br[59] wl[49] vdd gnd cell_6t
Xbit_r50_c59 bl[59] br[59] wl[50] vdd gnd cell_6t
Xbit_r51_c59 bl[59] br[59] wl[51] vdd gnd cell_6t
Xbit_r52_c59 bl[59] br[59] wl[52] vdd gnd cell_6t
Xbit_r53_c59 bl[59] br[59] wl[53] vdd gnd cell_6t
Xbit_r54_c59 bl[59] br[59] wl[54] vdd gnd cell_6t
Xbit_r55_c59 bl[59] br[59] wl[55] vdd gnd cell_6t
Xbit_r56_c59 bl[59] br[59] wl[56] vdd gnd cell_6t
Xbit_r57_c59 bl[59] br[59] wl[57] vdd gnd cell_6t
Xbit_r58_c59 bl[59] br[59] wl[58] vdd gnd cell_6t
Xbit_r59_c59 bl[59] br[59] wl[59] vdd gnd cell_6t
Xbit_r60_c59 bl[59] br[59] wl[60] vdd gnd cell_6t
Xbit_r61_c59 bl[59] br[59] wl[61] vdd gnd cell_6t
Xbit_r62_c59 bl[59] br[59] wl[62] vdd gnd cell_6t
Xbit_r63_c59 bl[59] br[59] wl[63] vdd gnd cell_6t
Xbit_r64_c59 bl[59] br[59] wl[64] vdd gnd cell_6t
Xbit_r65_c59 bl[59] br[59] wl[65] vdd gnd cell_6t
Xbit_r66_c59 bl[59] br[59] wl[66] vdd gnd cell_6t
Xbit_r67_c59 bl[59] br[59] wl[67] vdd gnd cell_6t
Xbit_r68_c59 bl[59] br[59] wl[68] vdd gnd cell_6t
Xbit_r69_c59 bl[59] br[59] wl[69] vdd gnd cell_6t
Xbit_r70_c59 bl[59] br[59] wl[70] vdd gnd cell_6t
Xbit_r71_c59 bl[59] br[59] wl[71] vdd gnd cell_6t
Xbit_r72_c59 bl[59] br[59] wl[72] vdd gnd cell_6t
Xbit_r73_c59 bl[59] br[59] wl[73] vdd gnd cell_6t
Xbit_r74_c59 bl[59] br[59] wl[74] vdd gnd cell_6t
Xbit_r75_c59 bl[59] br[59] wl[75] vdd gnd cell_6t
Xbit_r76_c59 bl[59] br[59] wl[76] vdd gnd cell_6t
Xbit_r77_c59 bl[59] br[59] wl[77] vdd gnd cell_6t
Xbit_r78_c59 bl[59] br[59] wl[78] vdd gnd cell_6t
Xbit_r79_c59 bl[59] br[59] wl[79] vdd gnd cell_6t
Xbit_r80_c59 bl[59] br[59] wl[80] vdd gnd cell_6t
Xbit_r81_c59 bl[59] br[59] wl[81] vdd gnd cell_6t
Xbit_r82_c59 bl[59] br[59] wl[82] vdd gnd cell_6t
Xbit_r83_c59 bl[59] br[59] wl[83] vdd gnd cell_6t
Xbit_r84_c59 bl[59] br[59] wl[84] vdd gnd cell_6t
Xbit_r85_c59 bl[59] br[59] wl[85] vdd gnd cell_6t
Xbit_r86_c59 bl[59] br[59] wl[86] vdd gnd cell_6t
Xbit_r87_c59 bl[59] br[59] wl[87] vdd gnd cell_6t
Xbit_r88_c59 bl[59] br[59] wl[88] vdd gnd cell_6t
Xbit_r89_c59 bl[59] br[59] wl[89] vdd gnd cell_6t
Xbit_r90_c59 bl[59] br[59] wl[90] vdd gnd cell_6t
Xbit_r91_c59 bl[59] br[59] wl[91] vdd gnd cell_6t
Xbit_r92_c59 bl[59] br[59] wl[92] vdd gnd cell_6t
Xbit_r93_c59 bl[59] br[59] wl[93] vdd gnd cell_6t
Xbit_r94_c59 bl[59] br[59] wl[94] vdd gnd cell_6t
Xbit_r95_c59 bl[59] br[59] wl[95] vdd gnd cell_6t
Xbit_r96_c59 bl[59] br[59] wl[96] vdd gnd cell_6t
Xbit_r97_c59 bl[59] br[59] wl[97] vdd gnd cell_6t
Xbit_r98_c59 bl[59] br[59] wl[98] vdd gnd cell_6t
Xbit_r99_c59 bl[59] br[59] wl[99] vdd gnd cell_6t
Xbit_r100_c59 bl[59] br[59] wl[100] vdd gnd cell_6t
Xbit_r101_c59 bl[59] br[59] wl[101] vdd gnd cell_6t
Xbit_r102_c59 bl[59] br[59] wl[102] vdd gnd cell_6t
Xbit_r103_c59 bl[59] br[59] wl[103] vdd gnd cell_6t
Xbit_r104_c59 bl[59] br[59] wl[104] vdd gnd cell_6t
Xbit_r105_c59 bl[59] br[59] wl[105] vdd gnd cell_6t
Xbit_r106_c59 bl[59] br[59] wl[106] vdd gnd cell_6t
Xbit_r107_c59 bl[59] br[59] wl[107] vdd gnd cell_6t
Xbit_r108_c59 bl[59] br[59] wl[108] vdd gnd cell_6t
Xbit_r109_c59 bl[59] br[59] wl[109] vdd gnd cell_6t
Xbit_r110_c59 bl[59] br[59] wl[110] vdd gnd cell_6t
Xbit_r111_c59 bl[59] br[59] wl[111] vdd gnd cell_6t
Xbit_r112_c59 bl[59] br[59] wl[112] vdd gnd cell_6t
Xbit_r113_c59 bl[59] br[59] wl[113] vdd gnd cell_6t
Xbit_r114_c59 bl[59] br[59] wl[114] vdd gnd cell_6t
Xbit_r115_c59 bl[59] br[59] wl[115] vdd gnd cell_6t
Xbit_r116_c59 bl[59] br[59] wl[116] vdd gnd cell_6t
Xbit_r117_c59 bl[59] br[59] wl[117] vdd gnd cell_6t
Xbit_r118_c59 bl[59] br[59] wl[118] vdd gnd cell_6t
Xbit_r119_c59 bl[59] br[59] wl[119] vdd gnd cell_6t
Xbit_r120_c59 bl[59] br[59] wl[120] vdd gnd cell_6t
Xbit_r121_c59 bl[59] br[59] wl[121] vdd gnd cell_6t
Xbit_r122_c59 bl[59] br[59] wl[122] vdd gnd cell_6t
Xbit_r123_c59 bl[59] br[59] wl[123] vdd gnd cell_6t
Xbit_r124_c59 bl[59] br[59] wl[124] vdd gnd cell_6t
Xbit_r125_c59 bl[59] br[59] wl[125] vdd gnd cell_6t
Xbit_r126_c59 bl[59] br[59] wl[126] vdd gnd cell_6t
Xbit_r127_c59 bl[59] br[59] wl[127] vdd gnd cell_6t
Xbit_r128_c59 bl[59] br[59] wl[128] vdd gnd cell_6t
Xbit_r129_c59 bl[59] br[59] wl[129] vdd gnd cell_6t
Xbit_r130_c59 bl[59] br[59] wl[130] vdd gnd cell_6t
Xbit_r131_c59 bl[59] br[59] wl[131] vdd gnd cell_6t
Xbit_r132_c59 bl[59] br[59] wl[132] vdd gnd cell_6t
Xbit_r133_c59 bl[59] br[59] wl[133] vdd gnd cell_6t
Xbit_r134_c59 bl[59] br[59] wl[134] vdd gnd cell_6t
Xbit_r135_c59 bl[59] br[59] wl[135] vdd gnd cell_6t
Xbit_r136_c59 bl[59] br[59] wl[136] vdd gnd cell_6t
Xbit_r137_c59 bl[59] br[59] wl[137] vdd gnd cell_6t
Xbit_r138_c59 bl[59] br[59] wl[138] vdd gnd cell_6t
Xbit_r139_c59 bl[59] br[59] wl[139] vdd gnd cell_6t
Xbit_r140_c59 bl[59] br[59] wl[140] vdd gnd cell_6t
Xbit_r141_c59 bl[59] br[59] wl[141] vdd gnd cell_6t
Xbit_r142_c59 bl[59] br[59] wl[142] vdd gnd cell_6t
Xbit_r143_c59 bl[59] br[59] wl[143] vdd gnd cell_6t
Xbit_r144_c59 bl[59] br[59] wl[144] vdd gnd cell_6t
Xbit_r145_c59 bl[59] br[59] wl[145] vdd gnd cell_6t
Xbit_r146_c59 bl[59] br[59] wl[146] vdd gnd cell_6t
Xbit_r147_c59 bl[59] br[59] wl[147] vdd gnd cell_6t
Xbit_r148_c59 bl[59] br[59] wl[148] vdd gnd cell_6t
Xbit_r149_c59 bl[59] br[59] wl[149] vdd gnd cell_6t
Xbit_r150_c59 bl[59] br[59] wl[150] vdd gnd cell_6t
Xbit_r151_c59 bl[59] br[59] wl[151] vdd gnd cell_6t
Xbit_r152_c59 bl[59] br[59] wl[152] vdd gnd cell_6t
Xbit_r153_c59 bl[59] br[59] wl[153] vdd gnd cell_6t
Xbit_r154_c59 bl[59] br[59] wl[154] vdd gnd cell_6t
Xbit_r155_c59 bl[59] br[59] wl[155] vdd gnd cell_6t
Xbit_r156_c59 bl[59] br[59] wl[156] vdd gnd cell_6t
Xbit_r157_c59 bl[59] br[59] wl[157] vdd gnd cell_6t
Xbit_r158_c59 bl[59] br[59] wl[158] vdd gnd cell_6t
Xbit_r159_c59 bl[59] br[59] wl[159] vdd gnd cell_6t
Xbit_r160_c59 bl[59] br[59] wl[160] vdd gnd cell_6t
Xbit_r161_c59 bl[59] br[59] wl[161] vdd gnd cell_6t
Xbit_r162_c59 bl[59] br[59] wl[162] vdd gnd cell_6t
Xbit_r163_c59 bl[59] br[59] wl[163] vdd gnd cell_6t
Xbit_r164_c59 bl[59] br[59] wl[164] vdd gnd cell_6t
Xbit_r165_c59 bl[59] br[59] wl[165] vdd gnd cell_6t
Xbit_r166_c59 bl[59] br[59] wl[166] vdd gnd cell_6t
Xbit_r167_c59 bl[59] br[59] wl[167] vdd gnd cell_6t
Xbit_r168_c59 bl[59] br[59] wl[168] vdd gnd cell_6t
Xbit_r169_c59 bl[59] br[59] wl[169] vdd gnd cell_6t
Xbit_r170_c59 bl[59] br[59] wl[170] vdd gnd cell_6t
Xbit_r171_c59 bl[59] br[59] wl[171] vdd gnd cell_6t
Xbit_r172_c59 bl[59] br[59] wl[172] vdd gnd cell_6t
Xbit_r173_c59 bl[59] br[59] wl[173] vdd gnd cell_6t
Xbit_r174_c59 bl[59] br[59] wl[174] vdd gnd cell_6t
Xbit_r175_c59 bl[59] br[59] wl[175] vdd gnd cell_6t
Xbit_r176_c59 bl[59] br[59] wl[176] vdd gnd cell_6t
Xbit_r177_c59 bl[59] br[59] wl[177] vdd gnd cell_6t
Xbit_r178_c59 bl[59] br[59] wl[178] vdd gnd cell_6t
Xbit_r179_c59 bl[59] br[59] wl[179] vdd gnd cell_6t
Xbit_r180_c59 bl[59] br[59] wl[180] vdd gnd cell_6t
Xbit_r181_c59 bl[59] br[59] wl[181] vdd gnd cell_6t
Xbit_r182_c59 bl[59] br[59] wl[182] vdd gnd cell_6t
Xbit_r183_c59 bl[59] br[59] wl[183] vdd gnd cell_6t
Xbit_r184_c59 bl[59] br[59] wl[184] vdd gnd cell_6t
Xbit_r185_c59 bl[59] br[59] wl[185] vdd gnd cell_6t
Xbit_r186_c59 bl[59] br[59] wl[186] vdd gnd cell_6t
Xbit_r187_c59 bl[59] br[59] wl[187] vdd gnd cell_6t
Xbit_r188_c59 bl[59] br[59] wl[188] vdd gnd cell_6t
Xbit_r189_c59 bl[59] br[59] wl[189] vdd gnd cell_6t
Xbit_r190_c59 bl[59] br[59] wl[190] vdd gnd cell_6t
Xbit_r191_c59 bl[59] br[59] wl[191] vdd gnd cell_6t
Xbit_r192_c59 bl[59] br[59] wl[192] vdd gnd cell_6t
Xbit_r193_c59 bl[59] br[59] wl[193] vdd gnd cell_6t
Xbit_r194_c59 bl[59] br[59] wl[194] vdd gnd cell_6t
Xbit_r195_c59 bl[59] br[59] wl[195] vdd gnd cell_6t
Xbit_r196_c59 bl[59] br[59] wl[196] vdd gnd cell_6t
Xbit_r197_c59 bl[59] br[59] wl[197] vdd gnd cell_6t
Xbit_r198_c59 bl[59] br[59] wl[198] vdd gnd cell_6t
Xbit_r199_c59 bl[59] br[59] wl[199] vdd gnd cell_6t
Xbit_r200_c59 bl[59] br[59] wl[200] vdd gnd cell_6t
Xbit_r201_c59 bl[59] br[59] wl[201] vdd gnd cell_6t
Xbit_r202_c59 bl[59] br[59] wl[202] vdd gnd cell_6t
Xbit_r203_c59 bl[59] br[59] wl[203] vdd gnd cell_6t
Xbit_r204_c59 bl[59] br[59] wl[204] vdd gnd cell_6t
Xbit_r205_c59 bl[59] br[59] wl[205] vdd gnd cell_6t
Xbit_r206_c59 bl[59] br[59] wl[206] vdd gnd cell_6t
Xbit_r207_c59 bl[59] br[59] wl[207] vdd gnd cell_6t
Xbit_r208_c59 bl[59] br[59] wl[208] vdd gnd cell_6t
Xbit_r209_c59 bl[59] br[59] wl[209] vdd gnd cell_6t
Xbit_r210_c59 bl[59] br[59] wl[210] vdd gnd cell_6t
Xbit_r211_c59 bl[59] br[59] wl[211] vdd gnd cell_6t
Xbit_r212_c59 bl[59] br[59] wl[212] vdd gnd cell_6t
Xbit_r213_c59 bl[59] br[59] wl[213] vdd gnd cell_6t
Xbit_r214_c59 bl[59] br[59] wl[214] vdd gnd cell_6t
Xbit_r215_c59 bl[59] br[59] wl[215] vdd gnd cell_6t
Xbit_r216_c59 bl[59] br[59] wl[216] vdd gnd cell_6t
Xbit_r217_c59 bl[59] br[59] wl[217] vdd gnd cell_6t
Xbit_r218_c59 bl[59] br[59] wl[218] vdd gnd cell_6t
Xbit_r219_c59 bl[59] br[59] wl[219] vdd gnd cell_6t
Xbit_r220_c59 bl[59] br[59] wl[220] vdd gnd cell_6t
Xbit_r221_c59 bl[59] br[59] wl[221] vdd gnd cell_6t
Xbit_r222_c59 bl[59] br[59] wl[222] vdd gnd cell_6t
Xbit_r223_c59 bl[59] br[59] wl[223] vdd gnd cell_6t
Xbit_r224_c59 bl[59] br[59] wl[224] vdd gnd cell_6t
Xbit_r225_c59 bl[59] br[59] wl[225] vdd gnd cell_6t
Xbit_r226_c59 bl[59] br[59] wl[226] vdd gnd cell_6t
Xbit_r227_c59 bl[59] br[59] wl[227] vdd gnd cell_6t
Xbit_r228_c59 bl[59] br[59] wl[228] vdd gnd cell_6t
Xbit_r229_c59 bl[59] br[59] wl[229] vdd gnd cell_6t
Xbit_r230_c59 bl[59] br[59] wl[230] vdd gnd cell_6t
Xbit_r231_c59 bl[59] br[59] wl[231] vdd gnd cell_6t
Xbit_r232_c59 bl[59] br[59] wl[232] vdd gnd cell_6t
Xbit_r233_c59 bl[59] br[59] wl[233] vdd gnd cell_6t
Xbit_r234_c59 bl[59] br[59] wl[234] vdd gnd cell_6t
Xbit_r235_c59 bl[59] br[59] wl[235] vdd gnd cell_6t
Xbit_r236_c59 bl[59] br[59] wl[236] vdd gnd cell_6t
Xbit_r237_c59 bl[59] br[59] wl[237] vdd gnd cell_6t
Xbit_r238_c59 bl[59] br[59] wl[238] vdd gnd cell_6t
Xbit_r239_c59 bl[59] br[59] wl[239] vdd gnd cell_6t
Xbit_r240_c59 bl[59] br[59] wl[240] vdd gnd cell_6t
Xbit_r241_c59 bl[59] br[59] wl[241] vdd gnd cell_6t
Xbit_r242_c59 bl[59] br[59] wl[242] vdd gnd cell_6t
Xbit_r243_c59 bl[59] br[59] wl[243] vdd gnd cell_6t
Xbit_r244_c59 bl[59] br[59] wl[244] vdd gnd cell_6t
Xbit_r245_c59 bl[59] br[59] wl[245] vdd gnd cell_6t
Xbit_r246_c59 bl[59] br[59] wl[246] vdd gnd cell_6t
Xbit_r247_c59 bl[59] br[59] wl[247] vdd gnd cell_6t
Xbit_r248_c59 bl[59] br[59] wl[248] vdd gnd cell_6t
Xbit_r249_c59 bl[59] br[59] wl[249] vdd gnd cell_6t
Xbit_r250_c59 bl[59] br[59] wl[250] vdd gnd cell_6t
Xbit_r251_c59 bl[59] br[59] wl[251] vdd gnd cell_6t
Xbit_r252_c59 bl[59] br[59] wl[252] vdd gnd cell_6t
Xbit_r253_c59 bl[59] br[59] wl[253] vdd gnd cell_6t
Xbit_r254_c59 bl[59] br[59] wl[254] vdd gnd cell_6t
Xbit_r255_c59 bl[59] br[59] wl[255] vdd gnd cell_6t
Xbit_r256_c59 bl[59] br[59] wl[256] vdd gnd cell_6t
Xbit_r257_c59 bl[59] br[59] wl[257] vdd gnd cell_6t
Xbit_r258_c59 bl[59] br[59] wl[258] vdd gnd cell_6t
Xbit_r259_c59 bl[59] br[59] wl[259] vdd gnd cell_6t
Xbit_r260_c59 bl[59] br[59] wl[260] vdd gnd cell_6t
Xbit_r261_c59 bl[59] br[59] wl[261] vdd gnd cell_6t
Xbit_r262_c59 bl[59] br[59] wl[262] vdd gnd cell_6t
Xbit_r263_c59 bl[59] br[59] wl[263] vdd gnd cell_6t
Xbit_r264_c59 bl[59] br[59] wl[264] vdd gnd cell_6t
Xbit_r265_c59 bl[59] br[59] wl[265] vdd gnd cell_6t
Xbit_r266_c59 bl[59] br[59] wl[266] vdd gnd cell_6t
Xbit_r267_c59 bl[59] br[59] wl[267] vdd gnd cell_6t
Xbit_r268_c59 bl[59] br[59] wl[268] vdd gnd cell_6t
Xbit_r269_c59 bl[59] br[59] wl[269] vdd gnd cell_6t
Xbit_r270_c59 bl[59] br[59] wl[270] vdd gnd cell_6t
Xbit_r271_c59 bl[59] br[59] wl[271] vdd gnd cell_6t
Xbit_r272_c59 bl[59] br[59] wl[272] vdd gnd cell_6t
Xbit_r273_c59 bl[59] br[59] wl[273] vdd gnd cell_6t
Xbit_r274_c59 bl[59] br[59] wl[274] vdd gnd cell_6t
Xbit_r275_c59 bl[59] br[59] wl[275] vdd gnd cell_6t
Xbit_r276_c59 bl[59] br[59] wl[276] vdd gnd cell_6t
Xbit_r277_c59 bl[59] br[59] wl[277] vdd gnd cell_6t
Xbit_r278_c59 bl[59] br[59] wl[278] vdd gnd cell_6t
Xbit_r279_c59 bl[59] br[59] wl[279] vdd gnd cell_6t
Xbit_r280_c59 bl[59] br[59] wl[280] vdd gnd cell_6t
Xbit_r281_c59 bl[59] br[59] wl[281] vdd gnd cell_6t
Xbit_r282_c59 bl[59] br[59] wl[282] vdd gnd cell_6t
Xbit_r283_c59 bl[59] br[59] wl[283] vdd gnd cell_6t
Xbit_r284_c59 bl[59] br[59] wl[284] vdd gnd cell_6t
Xbit_r285_c59 bl[59] br[59] wl[285] vdd gnd cell_6t
Xbit_r286_c59 bl[59] br[59] wl[286] vdd gnd cell_6t
Xbit_r287_c59 bl[59] br[59] wl[287] vdd gnd cell_6t
Xbit_r288_c59 bl[59] br[59] wl[288] vdd gnd cell_6t
Xbit_r289_c59 bl[59] br[59] wl[289] vdd gnd cell_6t
Xbit_r290_c59 bl[59] br[59] wl[290] vdd gnd cell_6t
Xbit_r291_c59 bl[59] br[59] wl[291] vdd gnd cell_6t
Xbit_r292_c59 bl[59] br[59] wl[292] vdd gnd cell_6t
Xbit_r293_c59 bl[59] br[59] wl[293] vdd gnd cell_6t
Xbit_r294_c59 bl[59] br[59] wl[294] vdd gnd cell_6t
Xbit_r295_c59 bl[59] br[59] wl[295] vdd gnd cell_6t
Xbit_r296_c59 bl[59] br[59] wl[296] vdd gnd cell_6t
Xbit_r297_c59 bl[59] br[59] wl[297] vdd gnd cell_6t
Xbit_r298_c59 bl[59] br[59] wl[298] vdd gnd cell_6t
Xbit_r299_c59 bl[59] br[59] wl[299] vdd gnd cell_6t
Xbit_r300_c59 bl[59] br[59] wl[300] vdd gnd cell_6t
Xbit_r301_c59 bl[59] br[59] wl[301] vdd gnd cell_6t
Xbit_r302_c59 bl[59] br[59] wl[302] vdd gnd cell_6t
Xbit_r303_c59 bl[59] br[59] wl[303] vdd gnd cell_6t
Xbit_r304_c59 bl[59] br[59] wl[304] vdd gnd cell_6t
Xbit_r305_c59 bl[59] br[59] wl[305] vdd gnd cell_6t
Xbit_r306_c59 bl[59] br[59] wl[306] vdd gnd cell_6t
Xbit_r307_c59 bl[59] br[59] wl[307] vdd gnd cell_6t
Xbit_r308_c59 bl[59] br[59] wl[308] vdd gnd cell_6t
Xbit_r309_c59 bl[59] br[59] wl[309] vdd gnd cell_6t
Xbit_r310_c59 bl[59] br[59] wl[310] vdd gnd cell_6t
Xbit_r311_c59 bl[59] br[59] wl[311] vdd gnd cell_6t
Xbit_r312_c59 bl[59] br[59] wl[312] vdd gnd cell_6t
Xbit_r313_c59 bl[59] br[59] wl[313] vdd gnd cell_6t
Xbit_r314_c59 bl[59] br[59] wl[314] vdd gnd cell_6t
Xbit_r315_c59 bl[59] br[59] wl[315] vdd gnd cell_6t
Xbit_r316_c59 bl[59] br[59] wl[316] vdd gnd cell_6t
Xbit_r317_c59 bl[59] br[59] wl[317] vdd gnd cell_6t
Xbit_r318_c59 bl[59] br[59] wl[318] vdd gnd cell_6t
Xbit_r319_c59 bl[59] br[59] wl[319] vdd gnd cell_6t
Xbit_r320_c59 bl[59] br[59] wl[320] vdd gnd cell_6t
Xbit_r321_c59 bl[59] br[59] wl[321] vdd gnd cell_6t
Xbit_r322_c59 bl[59] br[59] wl[322] vdd gnd cell_6t
Xbit_r323_c59 bl[59] br[59] wl[323] vdd gnd cell_6t
Xbit_r324_c59 bl[59] br[59] wl[324] vdd gnd cell_6t
Xbit_r325_c59 bl[59] br[59] wl[325] vdd gnd cell_6t
Xbit_r326_c59 bl[59] br[59] wl[326] vdd gnd cell_6t
Xbit_r327_c59 bl[59] br[59] wl[327] vdd gnd cell_6t
Xbit_r328_c59 bl[59] br[59] wl[328] vdd gnd cell_6t
Xbit_r329_c59 bl[59] br[59] wl[329] vdd gnd cell_6t
Xbit_r330_c59 bl[59] br[59] wl[330] vdd gnd cell_6t
Xbit_r331_c59 bl[59] br[59] wl[331] vdd gnd cell_6t
Xbit_r332_c59 bl[59] br[59] wl[332] vdd gnd cell_6t
Xbit_r333_c59 bl[59] br[59] wl[333] vdd gnd cell_6t
Xbit_r334_c59 bl[59] br[59] wl[334] vdd gnd cell_6t
Xbit_r335_c59 bl[59] br[59] wl[335] vdd gnd cell_6t
Xbit_r336_c59 bl[59] br[59] wl[336] vdd gnd cell_6t
Xbit_r337_c59 bl[59] br[59] wl[337] vdd gnd cell_6t
Xbit_r338_c59 bl[59] br[59] wl[338] vdd gnd cell_6t
Xbit_r339_c59 bl[59] br[59] wl[339] vdd gnd cell_6t
Xbit_r340_c59 bl[59] br[59] wl[340] vdd gnd cell_6t
Xbit_r341_c59 bl[59] br[59] wl[341] vdd gnd cell_6t
Xbit_r342_c59 bl[59] br[59] wl[342] vdd gnd cell_6t
Xbit_r343_c59 bl[59] br[59] wl[343] vdd gnd cell_6t
Xbit_r344_c59 bl[59] br[59] wl[344] vdd gnd cell_6t
Xbit_r345_c59 bl[59] br[59] wl[345] vdd gnd cell_6t
Xbit_r346_c59 bl[59] br[59] wl[346] vdd gnd cell_6t
Xbit_r347_c59 bl[59] br[59] wl[347] vdd gnd cell_6t
Xbit_r348_c59 bl[59] br[59] wl[348] vdd gnd cell_6t
Xbit_r349_c59 bl[59] br[59] wl[349] vdd gnd cell_6t
Xbit_r350_c59 bl[59] br[59] wl[350] vdd gnd cell_6t
Xbit_r351_c59 bl[59] br[59] wl[351] vdd gnd cell_6t
Xbit_r352_c59 bl[59] br[59] wl[352] vdd gnd cell_6t
Xbit_r353_c59 bl[59] br[59] wl[353] vdd gnd cell_6t
Xbit_r354_c59 bl[59] br[59] wl[354] vdd gnd cell_6t
Xbit_r355_c59 bl[59] br[59] wl[355] vdd gnd cell_6t
Xbit_r356_c59 bl[59] br[59] wl[356] vdd gnd cell_6t
Xbit_r357_c59 bl[59] br[59] wl[357] vdd gnd cell_6t
Xbit_r358_c59 bl[59] br[59] wl[358] vdd gnd cell_6t
Xbit_r359_c59 bl[59] br[59] wl[359] vdd gnd cell_6t
Xbit_r360_c59 bl[59] br[59] wl[360] vdd gnd cell_6t
Xbit_r361_c59 bl[59] br[59] wl[361] vdd gnd cell_6t
Xbit_r362_c59 bl[59] br[59] wl[362] vdd gnd cell_6t
Xbit_r363_c59 bl[59] br[59] wl[363] vdd gnd cell_6t
Xbit_r364_c59 bl[59] br[59] wl[364] vdd gnd cell_6t
Xbit_r365_c59 bl[59] br[59] wl[365] vdd gnd cell_6t
Xbit_r366_c59 bl[59] br[59] wl[366] vdd gnd cell_6t
Xbit_r367_c59 bl[59] br[59] wl[367] vdd gnd cell_6t
Xbit_r368_c59 bl[59] br[59] wl[368] vdd gnd cell_6t
Xbit_r369_c59 bl[59] br[59] wl[369] vdd gnd cell_6t
Xbit_r370_c59 bl[59] br[59] wl[370] vdd gnd cell_6t
Xbit_r371_c59 bl[59] br[59] wl[371] vdd gnd cell_6t
Xbit_r372_c59 bl[59] br[59] wl[372] vdd gnd cell_6t
Xbit_r373_c59 bl[59] br[59] wl[373] vdd gnd cell_6t
Xbit_r374_c59 bl[59] br[59] wl[374] vdd gnd cell_6t
Xbit_r375_c59 bl[59] br[59] wl[375] vdd gnd cell_6t
Xbit_r376_c59 bl[59] br[59] wl[376] vdd gnd cell_6t
Xbit_r377_c59 bl[59] br[59] wl[377] vdd gnd cell_6t
Xbit_r378_c59 bl[59] br[59] wl[378] vdd gnd cell_6t
Xbit_r379_c59 bl[59] br[59] wl[379] vdd gnd cell_6t
Xbit_r380_c59 bl[59] br[59] wl[380] vdd gnd cell_6t
Xbit_r381_c59 bl[59] br[59] wl[381] vdd gnd cell_6t
Xbit_r382_c59 bl[59] br[59] wl[382] vdd gnd cell_6t
Xbit_r383_c59 bl[59] br[59] wl[383] vdd gnd cell_6t
Xbit_r384_c59 bl[59] br[59] wl[384] vdd gnd cell_6t
Xbit_r385_c59 bl[59] br[59] wl[385] vdd gnd cell_6t
Xbit_r386_c59 bl[59] br[59] wl[386] vdd gnd cell_6t
Xbit_r387_c59 bl[59] br[59] wl[387] vdd gnd cell_6t
Xbit_r388_c59 bl[59] br[59] wl[388] vdd gnd cell_6t
Xbit_r389_c59 bl[59] br[59] wl[389] vdd gnd cell_6t
Xbit_r390_c59 bl[59] br[59] wl[390] vdd gnd cell_6t
Xbit_r391_c59 bl[59] br[59] wl[391] vdd gnd cell_6t
Xbit_r392_c59 bl[59] br[59] wl[392] vdd gnd cell_6t
Xbit_r393_c59 bl[59] br[59] wl[393] vdd gnd cell_6t
Xbit_r394_c59 bl[59] br[59] wl[394] vdd gnd cell_6t
Xbit_r395_c59 bl[59] br[59] wl[395] vdd gnd cell_6t
Xbit_r396_c59 bl[59] br[59] wl[396] vdd gnd cell_6t
Xbit_r397_c59 bl[59] br[59] wl[397] vdd gnd cell_6t
Xbit_r398_c59 bl[59] br[59] wl[398] vdd gnd cell_6t
Xbit_r399_c59 bl[59] br[59] wl[399] vdd gnd cell_6t
Xbit_r400_c59 bl[59] br[59] wl[400] vdd gnd cell_6t
Xbit_r401_c59 bl[59] br[59] wl[401] vdd gnd cell_6t
Xbit_r402_c59 bl[59] br[59] wl[402] vdd gnd cell_6t
Xbit_r403_c59 bl[59] br[59] wl[403] vdd gnd cell_6t
Xbit_r404_c59 bl[59] br[59] wl[404] vdd gnd cell_6t
Xbit_r405_c59 bl[59] br[59] wl[405] vdd gnd cell_6t
Xbit_r406_c59 bl[59] br[59] wl[406] vdd gnd cell_6t
Xbit_r407_c59 bl[59] br[59] wl[407] vdd gnd cell_6t
Xbit_r408_c59 bl[59] br[59] wl[408] vdd gnd cell_6t
Xbit_r409_c59 bl[59] br[59] wl[409] vdd gnd cell_6t
Xbit_r410_c59 bl[59] br[59] wl[410] vdd gnd cell_6t
Xbit_r411_c59 bl[59] br[59] wl[411] vdd gnd cell_6t
Xbit_r412_c59 bl[59] br[59] wl[412] vdd gnd cell_6t
Xbit_r413_c59 bl[59] br[59] wl[413] vdd gnd cell_6t
Xbit_r414_c59 bl[59] br[59] wl[414] vdd gnd cell_6t
Xbit_r415_c59 bl[59] br[59] wl[415] vdd gnd cell_6t
Xbit_r416_c59 bl[59] br[59] wl[416] vdd gnd cell_6t
Xbit_r417_c59 bl[59] br[59] wl[417] vdd gnd cell_6t
Xbit_r418_c59 bl[59] br[59] wl[418] vdd gnd cell_6t
Xbit_r419_c59 bl[59] br[59] wl[419] vdd gnd cell_6t
Xbit_r420_c59 bl[59] br[59] wl[420] vdd gnd cell_6t
Xbit_r421_c59 bl[59] br[59] wl[421] vdd gnd cell_6t
Xbit_r422_c59 bl[59] br[59] wl[422] vdd gnd cell_6t
Xbit_r423_c59 bl[59] br[59] wl[423] vdd gnd cell_6t
Xbit_r424_c59 bl[59] br[59] wl[424] vdd gnd cell_6t
Xbit_r425_c59 bl[59] br[59] wl[425] vdd gnd cell_6t
Xbit_r426_c59 bl[59] br[59] wl[426] vdd gnd cell_6t
Xbit_r427_c59 bl[59] br[59] wl[427] vdd gnd cell_6t
Xbit_r428_c59 bl[59] br[59] wl[428] vdd gnd cell_6t
Xbit_r429_c59 bl[59] br[59] wl[429] vdd gnd cell_6t
Xbit_r430_c59 bl[59] br[59] wl[430] vdd gnd cell_6t
Xbit_r431_c59 bl[59] br[59] wl[431] vdd gnd cell_6t
Xbit_r432_c59 bl[59] br[59] wl[432] vdd gnd cell_6t
Xbit_r433_c59 bl[59] br[59] wl[433] vdd gnd cell_6t
Xbit_r434_c59 bl[59] br[59] wl[434] vdd gnd cell_6t
Xbit_r435_c59 bl[59] br[59] wl[435] vdd gnd cell_6t
Xbit_r436_c59 bl[59] br[59] wl[436] vdd gnd cell_6t
Xbit_r437_c59 bl[59] br[59] wl[437] vdd gnd cell_6t
Xbit_r438_c59 bl[59] br[59] wl[438] vdd gnd cell_6t
Xbit_r439_c59 bl[59] br[59] wl[439] vdd gnd cell_6t
Xbit_r440_c59 bl[59] br[59] wl[440] vdd gnd cell_6t
Xbit_r441_c59 bl[59] br[59] wl[441] vdd gnd cell_6t
Xbit_r442_c59 bl[59] br[59] wl[442] vdd gnd cell_6t
Xbit_r443_c59 bl[59] br[59] wl[443] vdd gnd cell_6t
Xbit_r444_c59 bl[59] br[59] wl[444] vdd gnd cell_6t
Xbit_r445_c59 bl[59] br[59] wl[445] vdd gnd cell_6t
Xbit_r446_c59 bl[59] br[59] wl[446] vdd gnd cell_6t
Xbit_r447_c59 bl[59] br[59] wl[447] vdd gnd cell_6t
Xbit_r448_c59 bl[59] br[59] wl[448] vdd gnd cell_6t
Xbit_r449_c59 bl[59] br[59] wl[449] vdd gnd cell_6t
Xbit_r450_c59 bl[59] br[59] wl[450] vdd gnd cell_6t
Xbit_r451_c59 bl[59] br[59] wl[451] vdd gnd cell_6t
Xbit_r452_c59 bl[59] br[59] wl[452] vdd gnd cell_6t
Xbit_r453_c59 bl[59] br[59] wl[453] vdd gnd cell_6t
Xbit_r454_c59 bl[59] br[59] wl[454] vdd gnd cell_6t
Xbit_r455_c59 bl[59] br[59] wl[455] vdd gnd cell_6t
Xbit_r456_c59 bl[59] br[59] wl[456] vdd gnd cell_6t
Xbit_r457_c59 bl[59] br[59] wl[457] vdd gnd cell_6t
Xbit_r458_c59 bl[59] br[59] wl[458] vdd gnd cell_6t
Xbit_r459_c59 bl[59] br[59] wl[459] vdd gnd cell_6t
Xbit_r460_c59 bl[59] br[59] wl[460] vdd gnd cell_6t
Xbit_r461_c59 bl[59] br[59] wl[461] vdd gnd cell_6t
Xbit_r462_c59 bl[59] br[59] wl[462] vdd gnd cell_6t
Xbit_r463_c59 bl[59] br[59] wl[463] vdd gnd cell_6t
Xbit_r464_c59 bl[59] br[59] wl[464] vdd gnd cell_6t
Xbit_r465_c59 bl[59] br[59] wl[465] vdd gnd cell_6t
Xbit_r466_c59 bl[59] br[59] wl[466] vdd gnd cell_6t
Xbit_r467_c59 bl[59] br[59] wl[467] vdd gnd cell_6t
Xbit_r468_c59 bl[59] br[59] wl[468] vdd gnd cell_6t
Xbit_r469_c59 bl[59] br[59] wl[469] vdd gnd cell_6t
Xbit_r470_c59 bl[59] br[59] wl[470] vdd gnd cell_6t
Xbit_r471_c59 bl[59] br[59] wl[471] vdd gnd cell_6t
Xbit_r472_c59 bl[59] br[59] wl[472] vdd gnd cell_6t
Xbit_r473_c59 bl[59] br[59] wl[473] vdd gnd cell_6t
Xbit_r474_c59 bl[59] br[59] wl[474] vdd gnd cell_6t
Xbit_r475_c59 bl[59] br[59] wl[475] vdd gnd cell_6t
Xbit_r476_c59 bl[59] br[59] wl[476] vdd gnd cell_6t
Xbit_r477_c59 bl[59] br[59] wl[477] vdd gnd cell_6t
Xbit_r478_c59 bl[59] br[59] wl[478] vdd gnd cell_6t
Xbit_r479_c59 bl[59] br[59] wl[479] vdd gnd cell_6t
Xbit_r480_c59 bl[59] br[59] wl[480] vdd gnd cell_6t
Xbit_r481_c59 bl[59] br[59] wl[481] vdd gnd cell_6t
Xbit_r482_c59 bl[59] br[59] wl[482] vdd gnd cell_6t
Xbit_r483_c59 bl[59] br[59] wl[483] vdd gnd cell_6t
Xbit_r484_c59 bl[59] br[59] wl[484] vdd gnd cell_6t
Xbit_r485_c59 bl[59] br[59] wl[485] vdd gnd cell_6t
Xbit_r486_c59 bl[59] br[59] wl[486] vdd gnd cell_6t
Xbit_r487_c59 bl[59] br[59] wl[487] vdd gnd cell_6t
Xbit_r488_c59 bl[59] br[59] wl[488] vdd gnd cell_6t
Xbit_r489_c59 bl[59] br[59] wl[489] vdd gnd cell_6t
Xbit_r490_c59 bl[59] br[59] wl[490] vdd gnd cell_6t
Xbit_r491_c59 bl[59] br[59] wl[491] vdd gnd cell_6t
Xbit_r492_c59 bl[59] br[59] wl[492] vdd gnd cell_6t
Xbit_r493_c59 bl[59] br[59] wl[493] vdd gnd cell_6t
Xbit_r494_c59 bl[59] br[59] wl[494] vdd gnd cell_6t
Xbit_r495_c59 bl[59] br[59] wl[495] vdd gnd cell_6t
Xbit_r496_c59 bl[59] br[59] wl[496] vdd gnd cell_6t
Xbit_r497_c59 bl[59] br[59] wl[497] vdd gnd cell_6t
Xbit_r498_c59 bl[59] br[59] wl[498] vdd gnd cell_6t
Xbit_r499_c59 bl[59] br[59] wl[499] vdd gnd cell_6t
Xbit_r500_c59 bl[59] br[59] wl[500] vdd gnd cell_6t
Xbit_r501_c59 bl[59] br[59] wl[501] vdd gnd cell_6t
Xbit_r502_c59 bl[59] br[59] wl[502] vdd gnd cell_6t
Xbit_r503_c59 bl[59] br[59] wl[503] vdd gnd cell_6t
Xbit_r504_c59 bl[59] br[59] wl[504] vdd gnd cell_6t
Xbit_r505_c59 bl[59] br[59] wl[505] vdd gnd cell_6t
Xbit_r506_c59 bl[59] br[59] wl[506] vdd gnd cell_6t
Xbit_r507_c59 bl[59] br[59] wl[507] vdd gnd cell_6t
Xbit_r508_c59 bl[59] br[59] wl[508] vdd gnd cell_6t
Xbit_r509_c59 bl[59] br[59] wl[509] vdd gnd cell_6t
Xbit_r510_c59 bl[59] br[59] wl[510] vdd gnd cell_6t
Xbit_r511_c59 bl[59] br[59] wl[511] vdd gnd cell_6t
Xbit_r0_c60 bl[60] br[60] wl[0] vdd gnd cell_6t
Xbit_r1_c60 bl[60] br[60] wl[1] vdd gnd cell_6t
Xbit_r2_c60 bl[60] br[60] wl[2] vdd gnd cell_6t
Xbit_r3_c60 bl[60] br[60] wl[3] vdd gnd cell_6t
Xbit_r4_c60 bl[60] br[60] wl[4] vdd gnd cell_6t
Xbit_r5_c60 bl[60] br[60] wl[5] vdd gnd cell_6t
Xbit_r6_c60 bl[60] br[60] wl[6] vdd gnd cell_6t
Xbit_r7_c60 bl[60] br[60] wl[7] vdd gnd cell_6t
Xbit_r8_c60 bl[60] br[60] wl[8] vdd gnd cell_6t
Xbit_r9_c60 bl[60] br[60] wl[9] vdd gnd cell_6t
Xbit_r10_c60 bl[60] br[60] wl[10] vdd gnd cell_6t
Xbit_r11_c60 bl[60] br[60] wl[11] vdd gnd cell_6t
Xbit_r12_c60 bl[60] br[60] wl[12] vdd gnd cell_6t
Xbit_r13_c60 bl[60] br[60] wl[13] vdd gnd cell_6t
Xbit_r14_c60 bl[60] br[60] wl[14] vdd gnd cell_6t
Xbit_r15_c60 bl[60] br[60] wl[15] vdd gnd cell_6t
Xbit_r16_c60 bl[60] br[60] wl[16] vdd gnd cell_6t
Xbit_r17_c60 bl[60] br[60] wl[17] vdd gnd cell_6t
Xbit_r18_c60 bl[60] br[60] wl[18] vdd gnd cell_6t
Xbit_r19_c60 bl[60] br[60] wl[19] vdd gnd cell_6t
Xbit_r20_c60 bl[60] br[60] wl[20] vdd gnd cell_6t
Xbit_r21_c60 bl[60] br[60] wl[21] vdd gnd cell_6t
Xbit_r22_c60 bl[60] br[60] wl[22] vdd gnd cell_6t
Xbit_r23_c60 bl[60] br[60] wl[23] vdd gnd cell_6t
Xbit_r24_c60 bl[60] br[60] wl[24] vdd gnd cell_6t
Xbit_r25_c60 bl[60] br[60] wl[25] vdd gnd cell_6t
Xbit_r26_c60 bl[60] br[60] wl[26] vdd gnd cell_6t
Xbit_r27_c60 bl[60] br[60] wl[27] vdd gnd cell_6t
Xbit_r28_c60 bl[60] br[60] wl[28] vdd gnd cell_6t
Xbit_r29_c60 bl[60] br[60] wl[29] vdd gnd cell_6t
Xbit_r30_c60 bl[60] br[60] wl[30] vdd gnd cell_6t
Xbit_r31_c60 bl[60] br[60] wl[31] vdd gnd cell_6t
Xbit_r32_c60 bl[60] br[60] wl[32] vdd gnd cell_6t
Xbit_r33_c60 bl[60] br[60] wl[33] vdd gnd cell_6t
Xbit_r34_c60 bl[60] br[60] wl[34] vdd gnd cell_6t
Xbit_r35_c60 bl[60] br[60] wl[35] vdd gnd cell_6t
Xbit_r36_c60 bl[60] br[60] wl[36] vdd gnd cell_6t
Xbit_r37_c60 bl[60] br[60] wl[37] vdd gnd cell_6t
Xbit_r38_c60 bl[60] br[60] wl[38] vdd gnd cell_6t
Xbit_r39_c60 bl[60] br[60] wl[39] vdd gnd cell_6t
Xbit_r40_c60 bl[60] br[60] wl[40] vdd gnd cell_6t
Xbit_r41_c60 bl[60] br[60] wl[41] vdd gnd cell_6t
Xbit_r42_c60 bl[60] br[60] wl[42] vdd gnd cell_6t
Xbit_r43_c60 bl[60] br[60] wl[43] vdd gnd cell_6t
Xbit_r44_c60 bl[60] br[60] wl[44] vdd gnd cell_6t
Xbit_r45_c60 bl[60] br[60] wl[45] vdd gnd cell_6t
Xbit_r46_c60 bl[60] br[60] wl[46] vdd gnd cell_6t
Xbit_r47_c60 bl[60] br[60] wl[47] vdd gnd cell_6t
Xbit_r48_c60 bl[60] br[60] wl[48] vdd gnd cell_6t
Xbit_r49_c60 bl[60] br[60] wl[49] vdd gnd cell_6t
Xbit_r50_c60 bl[60] br[60] wl[50] vdd gnd cell_6t
Xbit_r51_c60 bl[60] br[60] wl[51] vdd gnd cell_6t
Xbit_r52_c60 bl[60] br[60] wl[52] vdd gnd cell_6t
Xbit_r53_c60 bl[60] br[60] wl[53] vdd gnd cell_6t
Xbit_r54_c60 bl[60] br[60] wl[54] vdd gnd cell_6t
Xbit_r55_c60 bl[60] br[60] wl[55] vdd gnd cell_6t
Xbit_r56_c60 bl[60] br[60] wl[56] vdd gnd cell_6t
Xbit_r57_c60 bl[60] br[60] wl[57] vdd gnd cell_6t
Xbit_r58_c60 bl[60] br[60] wl[58] vdd gnd cell_6t
Xbit_r59_c60 bl[60] br[60] wl[59] vdd gnd cell_6t
Xbit_r60_c60 bl[60] br[60] wl[60] vdd gnd cell_6t
Xbit_r61_c60 bl[60] br[60] wl[61] vdd gnd cell_6t
Xbit_r62_c60 bl[60] br[60] wl[62] vdd gnd cell_6t
Xbit_r63_c60 bl[60] br[60] wl[63] vdd gnd cell_6t
Xbit_r64_c60 bl[60] br[60] wl[64] vdd gnd cell_6t
Xbit_r65_c60 bl[60] br[60] wl[65] vdd gnd cell_6t
Xbit_r66_c60 bl[60] br[60] wl[66] vdd gnd cell_6t
Xbit_r67_c60 bl[60] br[60] wl[67] vdd gnd cell_6t
Xbit_r68_c60 bl[60] br[60] wl[68] vdd gnd cell_6t
Xbit_r69_c60 bl[60] br[60] wl[69] vdd gnd cell_6t
Xbit_r70_c60 bl[60] br[60] wl[70] vdd gnd cell_6t
Xbit_r71_c60 bl[60] br[60] wl[71] vdd gnd cell_6t
Xbit_r72_c60 bl[60] br[60] wl[72] vdd gnd cell_6t
Xbit_r73_c60 bl[60] br[60] wl[73] vdd gnd cell_6t
Xbit_r74_c60 bl[60] br[60] wl[74] vdd gnd cell_6t
Xbit_r75_c60 bl[60] br[60] wl[75] vdd gnd cell_6t
Xbit_r76_c60 bl[60] br[60] wl[76] vdd gnd cell_6t
Xbit_r77_c60 bl[60] br[60] wl[77] vdd gnd cell_6t
Xbit_r78_c60 bl[60] br[60] wl[78] vdd gnd cell_6t
Xbit_r79_c60 bl[60] br[60] wl[79] vdd gnd cell_6t
Xbit_r80_c60 bl[60] br[60] wl[80] vdd gnd cell_6t
Xbit_r81_c60 bl[60] br[60] wl[81] vdd gnd cell_6t
Xbit_r82_c60 bl[60] br[60] wl[82] vdd gnd cell_6t
Xbit_r83_c60 bl[60] br[60] wl[83] vdd gnd cell_6t
Xbit_r84_c60 bl[60] br[60] wl[84] vdd gnd cell_6t
Xbit_r85_c60 bl[60] br[60] wl[85] vdd gnd cell_6t
Xbit_r86_c60 bl[60] br[60] wl[86] vdd gnd cell_6t
Xbit_r87_c60 bl[60] br[60] wl[87] vdd gnd cell_6t
Xbit_r88_c60 bl[60] br[60] wl[88] vdd gnd cell_6t
Xbit_r89_c60 bl[60] br[60] wl[89] vdd gnd cell_6t
Xbit_r90_c60 bl[60] br[60] wl[90] vdd gnd cell_6t
Xbit_r91_c60 bl[60] br[60] wl[91] vdd gnd cell_6t
Xbit_r92_c60 bl[60] br[60] wl[92] vdd gnd cell_6t
Xbit_r93_c60 bl[60] br[60] wl[93] vdd gnd cell_6t
Xbit_r94_c60 bl[60] br[60] wl[94] vdd gnd cell_6t
Xbit_r95_c60 bl[60] br[60] wl[95] vdd gnd cell_6t
Xbit_r96_c60 bl[60] br[60] wl[96] vdd gnd cell_6t
Xbit_r97_c60 bl[60] br[60] wl[97] vdd gnd cell_6t
Xbit_r98_c60 bl[60] br[60] wl[98] vdd gnd cell_6t
Xbit_r99_c60 bl[60] br[60] wl[99] vdd gnd cell_6t
Xbit_r100_c60 bl[60] br[60] wl[100] vdd gnd cell_6t
Xbit_r101_c60 bl[60] br[60] wl[101] vdd gnd cell_6t
Xbit_r102_c60 bl[60] br[60] wl[102] vdd gnd cell_6t
Xbit_r103_c60 bl[60] br[60] wl[103] vdd gnd cell_6t
Xbit_r104_c60 bl[60] br[60] wl[104] vdd gnd cell_6t
Xbit_r105_c60 bl[60] br[60] wl[105] vdd gnd cell_6t
Xbit_r106_c60 bl[60] br[60] wl[106] vdd gnd cell_6t
Xbit_r107_c60 bl[60] br[60] wl[107] vdd gnd cell_6t
Xbit_r108_c60 bl[60] br[60] wl[108] vdd gnd cell_6t
Xbit_r109_c60 bl[60] br[60] wl[109] vdd gnd cell_6t
Xbit_r110_c60 bl[60] br[60] wl[110] vdd gnd cell_6t
Xbit_r111_c60 bl[60] br[60] wl[111] vdd gnd cell_6t
Xbit_r112_c60 bl[60] br[60] wl[112] vdd gnd cell_6t
Xbit_r113_c60 bl[60] br[60] wl[113] vdd gnd cell_6t
Xbit_r114_c60 bl[60] br[60] wl[114] vdd gnd cell_6t
Xbit_r115_c60 bl[60] br[60] wl[115] vdd gnd cell_6t
Xbit_r116_c60 bl[60] br[60] wl[116] vdd gnd cell_6t
Xbit_r117_c60 bl[60] br[60] wl[117] vdd gnd cell_6t
Xbit_r118_c60 bl[60] br[60] wl[118] vdd gnd cell_6t
Xbit_r119_c60 bl[60] br[60] wl[119] vdd gnd cell_6t
Xbit_r120_c60 bl[60] br[60] wl[120] vdd gnd cell_6t
Xbit_r121_c60 bl[60] br[60] wl[121] vdd gnd cell_6t
Xbit_r122_c60 bl[60] br[60] wl[122] vdd gnd cell_6t
Xbit_r123_c60 bl[60] br[60] wl[123] vdd gnd cell_6t
Xbit_r124_c60 bl[60] br[60] wl[124] vdd gnd cell_6t
Xbit_r125_c60 bl[60] br[60] wl[125] vdd gnd cell_6t
Xbit_r126_c60 bl[60] br[60] wl[126] vdd gnd cell_6t
Xbit_r127_c60 bl[60] br[60] wl[127] vdd gnd cell_6t
Xbit_r128_c60 bl[60] br[60] wl[128] vdd gnd cell_6t
Xbit_r129_c60 bl[60] br[60] wl[129] vdd gnd cell_6t
Xbit_r130_c60 bl[60] br[60] wl[130] vdd gnd cell_6t
Xbit_r131_c60 bl[60] br[60] wl[131] vdd gnd cell_6t
Xbit_r132_c60 bl[60] br[60] wl[132] vdd gnd cell_6t
Xbit_r133_c60 bl[60] br[60] wl[133] vdd gnd cell_6t
Xbit_r134_c60 bl[60] br[60] wl[134] vdd gnd cell_6t
Xbit_r135_c60 bl[60] br[60] wl[135] vdd gnd cell_6t
Xbit_r136_c60 bl[60] br[60] wl[136] vdd gnd cell_6t
Xbit_r137_c60 bl[60] br[60] wl[137] vdd gnd cell_6t
Xbit_r138_c60 bl[60] br[60] wl[138] vdd gnd cell_6t
Xbit_r139_c60 bl[60] br[60] wl[139] vdd gnd cell_6t
Xbit_r140_c60 bl[60] br[60] wl[140] vdd gnd cell_6t
Xbit_r141_c60 bl[60] br[60] wl[141] vdd gnd cell_6t
Xbit_r142_c60 bl[60] br[60] wl[142] vdd gnd cell_6t
Xbit_r143_c60 bl[60] br[60] wl[143] vdd gnd cell_6t
Xbit_r144_c60 bl[60] br[60] wl[144] vdd gnd cell_6t
Xbit_r145_c60 bl[60] br[60] wl[145] vdd gnd cell_6t
Xbit_r146_c60 bl[60] br[60] wl[146] vdd gnd cell_6t
Xbit_r147_c60 bl[60] br[60] wl[147] vdd gnd cell_6t
Xbit_r148_c60 bl[60] br[60] wl[148] vdd gnd cell_6t
Xbit_r149_c60 bl[60] br[60] wl[149] vdd gnd cell_6t
Xbit_r150_c60 bl[60] br[60] wl[150] vdd gnd cell_6t
Xbit_r151_c60 bl[60] br[60] wl[151] vdd gnd cell_6t
Xbit_r152_c60 bl[60] br[60] wl[152] vdd gnd cell_6t
Xbit_r153_c60 bl[60] br[60] wl[153] vdd gnd cell_6t
Xbit_r154_c60 bl[60] br[60] wl[154] vdd gnd cell_6t
Xbit_r155_c60 bl[60] br[60] wl[155] vdd gnd cell_6t
Xbit_r156_c60 bl[60] br[60] wl[156] vdd gnd cell_6t
Xbit_r157_c60 bl[60] br[60] wl[157] vdd gnd cell_6t
Xbit_r158_c60 bl[60] br[60] wl[158] vdd gnd cell_6t
Xbit_r159_c60 bl[60] br[60] wl[159] vdd gnd cell_6t
Xbit_r160_c60 bl[60] br[60] wl[160] vdd gnd cell_6t
Xbit_r161_c60 bl[60] br[60] wl[161] vdd gnd cell_6t
Xbit_r162_c60 bl[60] br[60] wl[162] vdd gnd cell_6t
Xbit_r163_c60 bl[60] br[60] wl[163] vdd gnd cell_6t
Xbit_r164_c60 bl[60] br[60] wl[164] vdd gnd cell_6t
Xbit_r165_c60 bl[60] br[60] wl[165] vdd gnd cell_6t
Xbit_r166_c60 bl[60] br[60] wl[166] vdd gnd cell_6t
Xbit_r167_c60 bl[60] br[60] wl[167] vdd gnd cell_6t
Xbit_r168_c60 bl[60] br[60] wl[168] vdd gnd cell_6t
Xbit_r169_c60 bl[60] br[60] wl[169] vdd gnd cell_6t
Xbit_r170_c60 bl[60] br[60] wl[170] vdd gnd cell_6t
Xbit_r171_c60 bl[60] br[60] wl[171] vdd gnd cell_6t
Xbit_r172_c60 bl[60] br[60] wl[172] vdd gnd cell_6t
Xbit_r173_c60 bl[60] br[60] wl[173] vdd gnd cell_6t
Xbit_r174_c60 bl[60] br[60] wl[174] vdd gnd cell_6t
Xbit_r175_c60 bl[60] br[60] wl[175] vdd gnd cell_6t
Xbit_r176_c60 bl[60] br[60] wl[176] vdd gnd cell_6t
Xbit_r177_c60 bl[60] br[60] wl[177] vdd gnd cell_6t
Xbit_r178_c60 bl[60] br[60] wl[178] vdd gnd cell_6t
Xbit_r179_c60 bl[60] br[60] wl[179] vdd gnd cell_6t
Xbit_r180_c60 bl[60] br[60] wl[180] vdd gnd cell_6t
Xbit_r181_c60 bl[60] br[60] wl[181] vdd gnd cell_6t
Xbit_r182_c60 bl[60] br[60] wl[182] vdd gnd cell_6t
Xbit_r183_c60 bl[60] br[60] wl[183] vdd gnd cell_6t
Xbit_r184_c60 bl[60] br[60] wl[184] vdd gnd cell_6t
Xbit_r185_c60 bl[60] br[60] wl[185] vdd gnd cell_6t
Xbit_r186_c60 bl[60] br[60] wl[186] vdd gnd cell_6t
Xbit_r187_c60 bl[60] br[60] wl[187] vdd gnd cell_6t
Xbit_r188_c60 bl[60] br[60] wl[188] vdd gnd cell_6t
Xbit_r189_c60 bl[60] br[60] wl[189] vdd gnd cell_6t
Xbit_r190_c60 bl[60] br[60] wl[190] vdd gnd cell_6t
Xbit_r191_c60 bl[60] br[60] wl[191] vdd gnd cell_6t
Xbit_r192_c60 bl[60] br[60] wl[192] vdd gnd cell_6t
Xbit_r193_c60 bl[60] br[60] wl[193] vdd gnd cell_6t
Xbit_r194_c60 bl[60] br[60] wl[194] vdd gnd cell_6t
Xbit_r195_c60 bl[60] br[60] wl[195] vdd gnd cell_6t
Xbit_r196_c60 bl[60] br[60] wl[196] vdd gnd cell_6t
Xbit_r197_c60 bl[60] br[60] wl[197] vdd gnd cell_6t
Xbit_r198_c60 bl[60] br[60] wl[198] vdd gnd cell_6t
Xbit_r199_c60 bl[60] br[60] wl[199] vdd gnd cell_6t
Xbit_r200_c60 bl[60] br[60] wl[200] vdd gnd cell_6t
Xbit_r201_c60 bl[60] br[60] wl[201] vdd gnd cell_6t
Xbit_r202_c60 bl[60] br[60] wl[202] vdd gnd cell_6t
Xbit_r203_c60 bl[60] br[60] wl[203] vdd gnd cell_6t
Xbit_r204_c60 bl[60] br[60] wl[204] vdd gnd cell_6t
Xbit_r205_c60 bl[60] br[60] wl[205] vdd gnd cell_6t
Xbit_r206_c60 bl[60] br[60] wl[206] vdd gnd cell_6t
Xbit_r207_c60 bl[60] br[60] wl[207] vdd gnd cell_6t
Xbit_r208_c60 bl[60] br[60] wl[208] vdd gnd cell_6t
Xbit_r209_c60 bl[60] br[60] wl[209] vdd gnd cell_6t
Xbit_r210_c60 bl[60] br[60] wl[210] vdd gnd cell_6t
Xbit_r211_c60 bl[60] br[60] wl[211] vdd gnd cell_6t
Xbit_r212_c60 bl[60] br[60] wl[212] vdd gnd cell_6t
Xbit_r213_c60 bl[60] br[60] wl[213] vdd gnd cell_6t
Xbit_r214_c60 bl[60] br[60] wl[214] vdd gnd cell_6t
Xbit_r215_c60 bl[60] br[60] wl[215] vdd gnd cell_6t
Xbit_r216_c60 bl[60] br[60] wl[216] vdd gnd cell_6t
Xbit_r217_c60 bl[60] br[60] wl[217] vdd gnd cell_6t
Xbit_r218_c60 bl[60] br[60] wl[218] vdd gnd cell_6t
Xbit_r219_c60 bl[60] br[60] wl[219] vdd gnd cell_6t
Xbit_r220_c60 bl[60] br[60] wl[220] vdd gnd cell_6t
Xbit_r221_c60 bl[60] br[60] wl[221] vdd gnd cell_6t
Xbit_r222_c60 bl[60] br[60] wl[222] vdd gnd cell_6t
Xbit_r223_c60 bl[60] br[60] wl[223] vdd gnd cell_6t
Xbit_r224_c60 bl[60] br[60] wl[224] vdd gnd cell_6t
Xbit_r225_c60 bl[60] br[60] wl[225] vdd gnd cell_6t
Xbit_r226_c60 bl[60] br[60] wl[226] vdd gnd cell_6t
Xbit_r227_c60 bl[60] br[60] wl[227] vdd gnd cell_6t
Xbit_r228_c60 bl[60] br[60] wl[228] vdd gnd cell_6t
Xbit_r229_c60 bl[60] br[60] wl[229] vdd gnd cell_6t
Xbit_r230_c60 bl[60] br[60] wl[230] vdd gnd cell_6t
Xbit_r231_c60 bl[60] br[60] wl[231] vdd gnd cell_6t
Xbit_r232_c60 bl[60] br[60] wl[232] vdd gnd cell_6t
Xbit_r233_c60 bl[60] br[60] wl[233] vdd gnd cell_6t
Xbit_r234_c60 bl[60] br[60] wl[234] vdd gnd cell_6t
Xbit_r235_c60 bl[60] br[60] wl[235] vdd gnd cell_6t
Xbit_r236_c60 bl[60] br[60] wl[236] vdd gnd cell_6t
Xbit_r237_c60 bl[60] br[60] wl[237] vdd gnd cell_6t
Xbit_r238_c60 bl[60] br[60] wl[238] vdd gnd cell_6t
Xbit_r239_c60 bl[60] br[60] wl[239] vdd gnd cell_6t
Xbit_r240_c60 bl[60] br[60] wl[240] vdd gnd cell_6t
Xbit_r241_c60 bl[60] br[60] wl[241] vdd gnd cell_6t
Xbit_r242_c60 bl[60] br[60] wl[242] vdd gnd cell_6t
Xbit_r243_c60 bl[60] br[60] wl[243] vdd gnd cell_6t
Xbit_r244_c60 bl[60] br[60] wl[244] vdd gnd cell_6t
Xbit_r245_c60 bl[60] br[60] wl[245] vdd gnd cell_6t
Xbit_r246_c60 bl[60] br[60] wl[246] vdd gnd cell_6t
Xbit_r247_c60 bl[60] br[60] wl[247] vdd gnd cell_6t
Xbit_r248_c60 bl[60] br[60] wl[248] vdd gnd cell_6t
Xbit_r249_c60 bl[60] br[60] wl[249] vdd gnd cell_6t
Xbit_r250_c60 bl[60] br[60] wl[250] vdd gnd cell_6t
Xbit_r251_c60 bl[60] br[60] wl[251] vdd gnd cell_6t
Xbit_r252_c60 bl[60] br[60] wl[252] vdd gnd cell_6t
Xbit_r253_c60 bl[60] br[60] wl[253] vdd gnd cell_6t
Xbit_r254_c60 bl[60] br[60] wl[254] vdd gnd cell_6t
Xbit_r255_c60 bl[60] br[60] wl[255] vdd gnd cell_6t
Xbit_r256_c60 bl[60] br[60] wl[256] vdd gnd cell_6t
Xbit_r257_c60 bl[60] br[60] wl[257] vdd gnd cell_6t
Xbit_r258_c60 bl[60] br[60] wl[258] vdd gnd cell_6t
Xbit_r259_c60 bl[60] br[60] wl[259] vdd gnd cell_6t
Xbit_r260_c60 bl[60] br[60] wl[260] vdd gnd cell_6t
Xbit_r261_c60 bl[60] br[60] wl[261] vdd gnd cell_6t
Xbit_r262_c60 bl[60] br[60] wl[262] vdd gnd cell_6t
Xbit_r263_c60 bl[60] br[60] wl[263] vdd gnd cell_6t
Xbit_r264_c60 bl[60] br[60] wl[264] vdd gnd cell_6t
Xbit_r265_c60 bl[60] br[60] wl[265] vdd gnd cell_6t
Xbit_r266_c60 bl[60] br[60] wl[266] vdd gnd cell_6t
Xbit_r267_c60 bl[60] br[60] wl[267] vdd gnd cell_6t
Xbit_r268_c60 bl[60] br[60] wl[268] vdd gnd cell_6t
Xbit_r269_c60 bl[60] br[60] wl[269] vdd gnd cell_6t
Xbit_r270_c60 bl[60] br[60] wl[270] vdd gnd cell_6t
Xbit_r271_c60 bl[60] br[60] wl[271] vdd gnd cell_6t
Xbit_r272_c60 bl[60] br[60] wl[272] vdd gnd cell_6t
Xbit_r273_c60 bl[60] br[60] wl[273] vdd gnd cell_6t
Xbit_r274_c60 bl[60] br[60] wl[274] vdd gnd cell_6t
Xbit_r275_c60 bl[60] br[60] wl[275] vdd gnd cell_6t
Xbit_r276_c60 bl[60] br[60] wl[276] vdd gnd cell_6t
Xbit_r277_c60 bl[60] br[60] wl[277] vdd gnd cell_6t
Xbit_r278_c60 bl[60] br[60] wl[278] vdd gnd cell_6t
Xbit_r279_c60 bl[60] br[60] wl[279] vdd gnd cell_6t
Xbit_r280_c60 bl[60] br[60] wl[280] vdd gnd cell_6t
Xbit_r281_c60 bl[60] br[60] wl[281] vdd gnd cell_6t
Xbit_r282_c60 bl[60] br[60] wl[282] vdd gnd cell_6t
Xbit_r283_c60 bl[60] br[60] wl[283] vdd gnd cell_6t
Xbit_r284_c60 bl[60] br[60] wl[284] vdd gnd cell_6t
Xbit_r285_c60 bl[60] br[60] wl[285] vdd gnd cell_6t
Xbit_r286_c60 bl[60] br[60] wl[286] vdd gnd cell_6t
Xbit_r287_c60 bl[60] br[60] wl[287] vdd gnd cell_6t
Xbit_r288_c60 bl[60] br[60] wl[288] vdd gnd cell_6t
Xbit_r289_c60 bl[60] br[60] wl[289] vdd gnd cell_6t
Xbit_r290_c60 bl[60] br[60] wl[290] vdd gnd cell_6t
Xbit_r291_c60 bl[60] br[60] wl[291] vdd gnd cell_6t
Xbit_r292_c60 bl[60] br[60] wl[292] vdd gnd cell_6t
Xbit_r293_c60 bl[60] br[60] wl[293] vdd gnd cell_6t
Xbit_r294_c60 bl[60] br[60] wl[294] vdd gnd cell_6t
Xbit_r295_c60 bl[60] br[60] wl[295] vdd gnd cell_6t
Xbit_r296_c60 bl[60] br[60] wl[296] vdd gnd cell_6t
Xbit_r297_c60 bl[60] br[60] wl[297] vdd gnd cell_6t
Xbit_r298_c60 bl[60] br[60] wl[298] vdd gnd cell_6t
Xbit_r299_c60 bl[60] br[60] wl[299] vdd gnd cell_6t
Xbit_r300_c60 bl[60] br[60] wl[300] vdd gnd cell_6t
Xbit_r301_c60 bl[60] br[60] wl[301] vdd gnd cell_6t
Xbit_r302_c60 bl[60] br[60] wl[302] vdd gnd cell_6t
Xbit_r303_c60 bl[60] br[60] wl[303] vdd gnd cell_6t
Xbit_r304_c60 bl[60] br[60] wl[304] vdd gnd cell_6t
Xbit_r305_c60 bl[60] br[60] wl[305] vdd gnd cell_6t
Xbit_r306_c60 bl[60] br[60] wl[306] vdd gnd cell_6t
Xbit_r307_c60 bl[60] br[60] wl[307] vdd gnd cell_6t
Xbit_r308_c60 bl[60] br[60] wl[308] vdd gnd cell_6t
Xbit_r309_c60 bl[60] br[60] wl[309] vdd gnd cell_6t
Xbit_r310_c60 bl[60] br[60] wl[310] vdd gnd cell_6t
Xbit_r311_c60 bl[60] br[60] wl[311] vdd gnd cell_6t
Xbit_r312_c60 bl[60] br[60] wl[312] vdd gnd cell_6t
Xbit_r313_c60 bl[60] br[60] wl[313] vdd gnd cell_6t
Xbit_r314_c60 bl[60] br[60] wl[314] vdd gnd cell_6t
Xbit_r315_c60 bl[60] br[60] wl[315] vdd gnd cell_6t
Xbit_r316_c60 bl[60] br[60] wl[316] vdd gnd cell_6t
Xbit_r317_c60 bl[60] br[60] wl[317] vdd gnd cell_6t
Xbit_r318_c60 bl[60] br[60] wl[318] vdd gnd cell_6t
Xbit_r319_c60 bl[60] br[60] wl[319] vdd gnd cell_6t
Xbit_r320_c60 bl[60] br[60] wl[320] vdd gnd cell_6t
Xbit_r321_c60 bl[60] br[60] wl[321] vdd gnd cell_6t
Xbit_r322_c60 bl[60] br[60] wl[322] vdd gnd cell_6t
Xbit_r323_c60 bl[60] br[60] wl[323] vdd gnd cell_6t
Xbit_r324_c60 bl[60] br[60] wl[324] vdd gnd cell_6t
Xbit_r325_c60 bl[60] br[60] wl[325] vdd gnd cell_6t
Xbit_r326_c60 bl[60] br[60] wl[326] vdd gnd cell_6t
Xbit_r327_c60 bl[60] br[60] wl[327] vdd gnd cell_6t
Xbit_r328_c60 bl[60] br[60] wl[328] vdd gnd cell_6t
Xbit_r329_c60 bl[60] br[60] wl[329] vdd gnd cell_6t
Xbit_r330_c60 bl[60] br[60] wl[330] vdd gnd cell_6t
Xbit_r331_c60 bl[60] br[60] wl[331] vdd gnd cell_6t
Xbit_r332_c60 bl[60] br[60] wl[332] vdd gnd cell_6t
Xbit_r333_c60 bl[60] br[60] wl[333] vdd gnd cell_6t
Xbit_r334_c60 bl[60] br[60] wl[334] vdd gnd cell_6t
Xbit_r335_c60 bl[60] br[60] wl[335] vdd gnd cell_6t
Xbit_r336_c60 bl[60] br[60] wl[336] vdd gnd cell_6t
Xbit_r337_c60 bl[60] br[60] wl[337] vdd gnd cell_6t
Xbit_r338_c60 bl[60] br[60] wl[338] vdd gnd cell_6t
Xbit_r339_c60 bl[60] br[60] wl[339] vdd gnd cell_6t
Xbit_r340_c60 bl[60] br[60] wl[340] vdd gnd cell_6t
Xbit_r341_c60 bl[60] br[60] wl[341] vdd gnd cell_6t
Xbit_r342_c60 bl[60] br[60] wl[342] vdd gnd cell_6t
Xbit_r343_c60 bl[60] br[60] wl[343] vdd gnd cell_6t
Xbit_r344_c60 bl[60] br[60] wl[344] vdd gnd cell_6t
Xbit_r345_c60 bl[60] br[60] wl[345] vdd gnd cell_6t
Xbit_r346_c60 bl[60] br[60] wl[346] vdd gnd cell_6t
Xbit_r347_c60 bl[60] br[60] wl[347] vdd gnd cell_6t
Xbit_r348_c60 bl[60] br[60] wl[348] vdd gnd cell_6t
Xbit_r349_c60 bl[60] br[60] wl[349] vdd gnd cell_6t
Xbit_r350_c60 bl[60] br[60] wl[350] vdd gnd cell_6t
Xbit_r351_c60 bl[60] br[60] wl[351] vdd gnd cell_6t
Xbit_r352_c60 bl[60] br[60] wl[352] vdd gnd cell_6t
Xbit_r353_c60 bl[60] br[60] wl[353] vdd gnd cell_6t
Xbit_r354_c60 bl[60] br[60] wl[354] vdd gnd cell_6t
Xbit_r355_c60 bl[60] br[60] wl[355] vdd gnd cell_6t
Xbit_r356_c60 bl[60] br[60] wl[356] vdd gnd cell_6t
Xbit_r357_c60 bl[60] br[60] wl[357] vdd gnd cell_6t
Xbit_r358_c60 bl[60] br[60] wl[358] vdd gnd cell_6t
Xbit_r359_c60 bl[60] br[60] wl[359] vdd gnd cell_6t
Xbit_r360_c60 bl[60] br[60] wl[360] vdd gnd cell_6t
Xbit_r361_c60 bl[60] br[60] wl[361] vdd gnd cell_6t
Xbit_r362_c60 bl[60] br[60] wl[362] vdd gnd cell_6t
Xbit_r363_c60 bl[60] br[60] wl[363] vdd gnd cell_6t
Xbit_r364_c60 bl[60] br[60] wl[364] vdd gnd cell_6t
Xbit_r365_c60 bl[60] br[60] wl[365] vdd gnd cell_6t
Xbit_r366_c60 bl[60] br[60] wl[366] vdd gnd cell_6t
Xbit_r367_c60 bl[60] br[60] wl[367] vdd gnd cell_6t
Xbit_r368_c60 bl[60] br[60] wl[368] vdd gnd cell_6t
Xbit_r369_c60 bl[60] br[60] wl[369] vdd gnd cell_6t
Xbit_r370_c60 bl[60] br[60] wl[370] vdd gnd cell_6t
Xbit_r371_c60 bl[60] br[60] wl[371] vdd gnd cell_6t
Xbit_r372_c60 bl[60] br[60] wl[372] vdd gnd cell_6t
Xbit_r373_c60 bl[60] br[60] wl[373] vdd gnd cell_6t
Xbit_r374_c60 bl[60] br[60] wl[374] vdd gnd cell_6t
Xbit_r375_c60 bl[60] br[60] wl[375] vdd gnd cell_6t
Xbit_r376_c60 bl[60] br[60] wl[376] vdd gnd cell_6t
Xbit_r377_c60 bl[60] br[60] wl[377] vdd gnd cell_6t
Xbit_r378_c60 bl[60] br[60] wl[378] vdd gnd cell_6t
Xbit_r379_c60 bl[60] br[60] wl[379] vdd gnd cell_6t
Xbit_r380_c60 bl[60] br[60] wl[380] vdd gnd cell_6t
Xbit_r381_c60 bl[60] br[60] wl[381] vdd gnd cell_6t
Xbit_r382_c60 bl[60] br[60] wl[382] vdd gnd cell_6t
Xbit_r383_c60 bl[60] br[60] wl[383] vdd gnd cell_6t
Xbit_r384_c60 bl[60] br[60] wl[384] vdd gnd cell_6t
Xbit_r385_c60 bl[60] br[60] wl[385] vdd gnd cell_6t
Xbit_r386_c60 bl[60] br[60] wl[386] vdd gnd cell_6t
Xbit_r387_c60 bl[60] br[60] wl[387] vdd gnd cell_6t
Xbit_r388_c60 bl[60] br[60] wl[388] vdd gnd cell_6t
Xbit_r389_c60 bl[60] br[60] wl[389] vdd gnd cell_6t
Xbit_r390_c60 bl[60] br[60] wl[390] vdd gnd cell_6t
Xbit_r391_c60 bl[60] br[60] wl[391] vdd gnd cell_6t
Xbit_r392_c60 bl[60] br[60] wl[392] vdd gnd cell_6t
Xbit_r393_c60 bl[60] br[60] wl[393] vdd gnd cell_6t
Xbit_r394_c60 bl[60] br[60] wl[394] vdd gnd cell_6t
Xbit_r395_c60 bl[60] br[60] wl[395] vdd gnd cell_6t
Xbit_r396_c60 bl[60] br[60] wl[396] vdd gnd cell_6t
Xbit_r397_c60 bl[60] br[60] wl[397] vdd gnd cell_6t
Xbit_r398_c60 bl[60] br[60] wl[398] vdd gnd cell_6t
Xbit_r399_c60 bl[60] br[60] wl[399] vdd gnd cell_6t
Xbit_r400_c60 bl[60] br[60] wl[400] vdd gnd cell_6t
Xbit_r401_c60 bl[60] br[60] wl[401] vdd gnd cell_6t
Xbit_r402_c60 bl[60] br[60] wl[402] vdd gnd cell_6t
Xbit_r403_c60 bl[60] br[60] wl[403] vdd gnd cell_6t
Xbit_r404_c60 bl[60] br[60] wl[404] vdd gnd cell_6t
Xbit_r405_c60 bl[60] br[60] wl[405] vdd gnd cell_6t
Xbit_r406_c60 bl[60] br[60] wl[406] vdd gnd cell_6t
Xbit_r407_c60 bl[60] br[60] wl[407] vdd gnd cell_6t
Xbit_r408_c60 bl[60] br[60] wl[408] vdd gnd cell_6t
Xbit_r409_c60 bl[60] br[60] wl[409] vdd gnd cell_6t
Xbit_r410_c60 bl[60] br[60] wl[410] vdd gnd cell_6t
Xbit_r411_c60 bl[60] br[60] wl[411] vdd gnd cell_6t
Xbit_r412_c60 bl[60] br[60] wl[412] vdd gnd cell_6t
Xbit_r413_c60 bl[60] br[60] wl[413] vdd gnd cell_6t
Xbit_r414_c60 bl[60] br[60] wl[414] vdd gnd cell_6t
Xbit_r415_c60 bl[60] br[60] wl[415] vdd gnd cell_6t
Xbit_r416_c60 bl[60] br[60] wl[416] vdd gnd cell_6t
Xbit_r417_c60 bl[60] br[60] wl[417] vdd gnd cell_6t
Xbit_r418_c60 bl[60] br[60] wl[418] vdd gnd cell_6t
Xbit_r419_c60 bl[60] br[60] wl[419] vdd gnd cell_6t
Xbit_r420_c60 bl[60] br[60] wl[420] vdd gnd cell_6t
Xbit_r421_c60 bl[60] br[60] wl[421] vdd gnd cell_6t
Xbit_r422_c60 bl[60] br[60] wl[422] vdd gnd cell_6t
Xbit_r423_c60 bl[60] br[60] wl[423] vdd gnd cell_6t
Xbit_r424_c60 bl[60] br[60] wl[424] vdd gnd cell_6t
Xbit_r425_c60 bl[60] br[60] wl[425] vdd gnd cell_6t
Xbit_r426_c60 bl[60] br[60] wl[426] vdd gnd cell_6t
Xbit_r427_c60 bl[60] br[60] wl[427] vdd gnd cell_6t
Xbit_r428_c60 bl[60] br[60] wl[428] vdd gnd cell_6t
Xbit_r429_c60 bl[60] br[60] wl[429] vdd gnd cell_6t
Xbit_r430_c60 bl[60] br[60] wl[430] vdd gnd cell_6t
Xbit_r431_c60 bl[60] br[60] wl[431] vdd gnd cell_6t
Xbit_r432_c60 bl[60] br[60] wl[432] vdd gnd cell_6t
Xbit_r433_c60 bl[60] br[60] wl[433] vdd gnd cell_6t
Xbit_r434_c60 bl[60] br[60] wl[434] vdd gnd cell_6t
Xbit_r435_c60 bl[60] br[60] wl[435] vdd gnd cell_6t
Xbit_r436_c60 bl[60] br[60] wl[436] vdd gnd cell_6t
Xbit_r437_c60 bl[60] br[60] wl[437] vdd gnd cell_6t
Xbit_r438_c60 bl[60] br[60] wl[438] vdd gnd cell_6t
Xbit_r439_c60 bl[60] br[60] wl[439] vdd gnd cell_6t
Xbit_r440_c60 bl[60] br[60] wl[440] vdd gnd cell_6t
Xbit_r441_c60 bl[60] br[60] wl[441] vdd gnd cell_6t
Xbit_r442_c60 bl[60] br[60] wl[442] vdd gnd cell_6t
Xbit_r443_c60 bl[60] br[60] wl[443] vdd gnd cell_6t
Xbit_r444_c60 bl[60] br[60] wl[444] vdd gnd cell_6t
Xbit_r445_c60 bl[60] br[60] wl[445] vdd gnd cell_6t
Xbit_r446_c60 bl[60] br[60] wl[446] vdd gnd cell_6t
Xbit_r447_c60 bl[60] br[60] wl[447] vdd gnd cell_6t
Xbit_r448_c60 bl[60] br[60] wl[448] vdd gnd cell_6t
Xbit_r449_c60 bl[60] br[60] wl[449] vdd gnd cell_6t
Xbit_r450_c60 bl[60] br[60] wl[450] vdd gnd cell_6t
Xbit_r451_c60 bl[60] br[60] wl[451] vdd gnd cell_6t
Xbit_r452_c60 bl[60] br[60] wl[452] vdd gnd cell_6t
Xbit_r453_c60 bl[60] br[60] wl[453] vdd gnd cell_6t
Xbit_r454_c60 bl[60] br[60] wl[454] vdd gnd cell_6t
Xbit_r455_c60 bl[60] br[60] wl[455] vdd gnd cell_6t
Xbit_r456_c60 bl[60] br[60] wl[456] vdd gnd cell_6t
Xbit_r457_c60 bl[60] br[60] wl[457] vdd gnd cell_6t
Xbit_r458_c60 bl[60] br[60] wl[458] vdd gnd cell_6t
Xbit_r459_c60 bl[60] br[60] wl[459] vdd gnd cell_6t
Xbit_r460_c60 bl[60] br[60] wl[460] vdd gnd cell_6t
Xbit_r461_c60 bl[60] br[60] wl[461] vdd gnd cell_6t
Xbit_r462_c60 bl[60] br[60] wl[462] vdd gnd cell_6t
Xbit_r463_c60 bl[60] br[60] wl[463] vdd gnd cell_6t
Xbit_r464_c60 bl[60] br[60] wl[464] vdd gnd cell_6t
Xbit_r465_c60 bl[60] br[60] wl[465] vdd gnd cell_6t
Xbit_r466_c60 bl[60] br[60] wl[466] vdd gnd cell_6t
Xbit_r467_c60 bl[60] br[60] wl[467] vdd gnd cell_6t
Xbit_r468_c60 bl[60] br[60] wl[468] vdd gnd cell_6t
Xbit_r469_c60 bl[60] br[60] wl[469] vdd gnd cell_6t
Xbit_r470_c60 bl[60] br[60] wl[470] vdd gnd cell_6t
Xbit_r471_c60 bl[60] br[60] wl[471] vdd gnd cell_6t
Xbit_r472_c60 bl[60] br[60] wl[472] vdd gnd cell_6t
Xbit_r473_c60 bl[60] br[60] wl[473] vdd gnd cell_6t
Xbit_r474_c60 bl[60] br[60] wl[474] vdd gnd cell_6t
Xbit_r475_c60 bl[60] br[60] wl[475] vdd gnd cell_6t
Xbit_r476_c60 bl[60] br[60] wl[476] vdd gnd cell_6t
Xbit_r477_c60 bl[60] br[60] wl[477] vdd gnd cell_6t
Xbit_r478_c60 bl[60] br[60] wl[478] vdd gnd cell_6t
Xbit_r479_c60 bl[60] br[60] wl[479] vdd gnd cell_6t
Xbit_r480_c60 bl[60] br[60] wl[480] vdd gnd cell_6t
Xbit_r481_c60 bl[60] br[60] wl[481] vdd gnd cell_6t
Xbit_r482_c60 bl[60] br[60] wl[482] vdd gnd cell_6t
Xbit_r483_c60 bl[60] br[60] wl[483] vdd gnd cell_6t
Xbit_r484_c60 bl[60] br[60] wl[484] vdd gnd cell_6t
Xbit_r485_c60 bl[60] br[60] wl[485] vdd gnd cell_6t
Xbit_r486_c60 bl[60] br[60] wl[486] vdd gnd cell_6t
Xbit_r487_c60 bl[60] br[60] wl[487] vdd gnd cell_6t
Xbit_r488_c60 bl[60] br[60] wl[488] vdd gnd cell_6t
Xbit_r489_c60 bl[60] br[60] wl[489] vdd gnd cell_6t
Xbit_r490_c60 bl[60] br[60] wl[490] vdd gnd cell_6t
Xbit_r491_c60 bl[60] br[60] wl[491] vdd gnd cell_6t
Xbit_r492_c60 bl[60] br[60] wl[492] vdd gnd cell_6t
Xbit_r493_c60 bl[60] br[60] wl[493] vdd gnd cell_6t
Xbit_r494_c60 bl[60] br[60] wl[494] vdd gnd cell_6t
Xbit_r495_c60 bl[60] br[60] wl[495] vdd gnd cell_6t
Xbit_r496_c60 bl[60] br[60] wl[496] vdd gnd cell_6t
Xbit_r497_c60 bl[60] br[60] wl[497] vdd gnd cell_6t
Xbit_r498_c60 bl[60] br[60] wl[498] vdd gnd cell_6t
Xbit_r499_c60 bl[60] br[60] wl[499] vdd gnd cell_6t
Xbit_r500_c60 bl[60] br[60] wl[500] vdd gnd cell_6t
Xbit_r501_c60 bl[60] br[60] wl[501] vdd gnd cell_6t
Xbit_r502_c60 bl[60] br[60] wl[502] vdd gnd cell_6t
Xbit_r503_c60 bl[60] br[60] wl[503] vdd gnd cell_6t
Xbit_r504_c60 bl[60] br[60] wl[504] vdd gnd cell_6t
Xbit_r505_c60 bl[60] br[60] wl[505] vdd gnd cell_6t
Xbit_r506_c60 bl[60] br[60] wl[506] vdd gnd cell_6t
Xbit_r507_c60 bl[60] br[60] wl[507] vdd gnd cell_6t
Xbit_r508_c60 bl[60] br[60] wl[508] vdd gnd cell_6t
Xbit_r509_c60 bl[60] br[60] wl[509] vdd gnd cell_6t
Xbit_r510_c60 bl[60] br[60] wl[510] vdd gnd cell_6t
Xbit_r511_c60 bl[60] br[60] wl[511] vdd gnd cell_6t
Xbit_r0_c61 bl[61] br[61] wl[0] vdd gnd cell_6t
Xbit_r1_c61 bl[61] br[61] wl[1] vdd gnd cell_6t
Xbit_r2_c61 bl[61] br[61] wl[2] vdd gnd cell_6t
Xbit_r3_c61 bl[61] br[61] wl[3] vdd gnd cell_6t
Xbit_r4_c61 bl[61] br[61] wl[4] vdd gnd cell_6t
Xbit_r5_c61 bl[61] br[61] wl[5] vdd gnd cell_6t
Xbit_r6_c61 bl[61] br[61] wl[6] vdd gnd cell_6t
Xbit_r7_c61 bl[61] br[61] wl[7] vdd gnd cell_6t
Xbit_r8_c61 bl[61] br[61] wl[8] vdd gnd cell_6t
Xbit_r9_c61 bl[61] br[61] wl[9] vdd gnd cell_6t
Xbit_r10_c61 bl[61] br[61] wl[10] vdd gnd cell_6t
Xbit_r11_c61 bl[61] br[61] wl[11] vdd gnd cell_6t
Xbit_r12_c61 bl[61] br[61] wl[12] vdd gnd cell_6t
Xbit_r13_c61 bl[61] br[61] wl[13] vdd gnd cell_6t
Xbit_r14_c61 bl[61] br[61] wl[14] vdd gnd cell_6t
Xbit_r15_c61 bl[61] br[61] wl[15] vdd gnd cell_6t
Xbit_r16_c61 bl[61] br[61] wl[16] vdd gnd cell_6t
Xbit_r17_c61 bl[61] br[61] wl[17] vdd gnd cell_6t
Xbit_r18_c61 bl[61] br[61] wl[18] vdd gnd cell_6t
Xbit_r19_c61 bl[61] br[61] wl[19] vdd gnd cell_6t
Xbit_r20_c61 bl[61] br[61] wl[20] vdd gnd cell_6t
Xbit_r21_c61 bl[61] br[61] wl[21] vdd gnd cell_6t
Xbit_r22_c61 bl[61] br[61] wl[22] vdd gnd cell_6t
Xbit_r23_c61 bl[61] br[61] wl[23] vdd gnd cell_6t
Xbit_r24_c61 bl[61] br[61] wl[24] vdd gnd cell_6t
Xbit_r25_c61 bl[61] br[61] wl[25] vdd gnd cell_6t
Xbit_r26_c61 bl[61] br[61] wl[26] vdd gnd cell_6t
Xbit_r27_c61 bl[61] br[61] wl[27] vdd gnd cell_6t
Xbit_r28_c61 bl[61] br[61] wl[28] vdd gnd cell_6t
Xbit_r29_c61 bl[61] br[61] wl[29] vdd gnd cell_6t
Xbit_r30_c61 bl[61] br[61] wl[30] vdd gnd cell_6t
Xbit_r31_c61 bl[61] br[61] wl[31] vdd gnd cell_6t
Xbit_r32_c61 bl[61] br[61] wl[32] vdd gnd cell_6t
Xbit_r33_c61 bl[61] br[61] wl[33] vdd gnd cell_6t
Xbit_r34_c61 bl[61] br[61] wl[34] vdd gnd cell_6t
Xbit_r35_c61 bl[61] br[61] wl[35] vdd gnd cell_6t
Xbit_r36_c61 bl[61] br[61] wl[36] vdd gnd cell_6t
Xbit_r37_c61 bl[61] br[61] wl[37] vdd gnd cell_6t
Xbit_r38_c61 bl[61] br[61] wl[38] vdd gnd cell_6t
Xbit_r39_c61 bl[61] br[61] wl[39] vdd gnd cell_6t
Xbit_r40_c61 bl[61] br[61] wl[40] vdd gnd cell_6t
Xbit_r41_c61 bl[61] br[61] wl[41] vdd gnd cell_6t
Xbit_r42_c61 bl[61] br[61] wl[42] vdd gnd cell_6t
Xbit_r43_c61 bl[61] br[61] wl[43] vdd gnd cell_6t
Xbit_r44_c61 bl[61] br[61] wl[44] vdd gnd cell_6t
Xbit_r45_c61 bl[61] br[61] wl[45] vdd gnd cell_6t
Xbit_r46_c61 bl[61] br[61] wl[46] vdd gnd cell_6t
Xbit_r47_c61 bl[61] br[61] wl[47] vdd gnd cell_6t
Xbit_r48_c61 bl[61] br[61] wl[48] vdd gnd cell_6t
Xbit_r49_c61 bl[61] br[61] wl[49] vdd gnd cell_6t
Xbit_r50_c61 bl[61] br[61] wl[50] vdd gnd cell_6t
Xbit_r51_c61 bl[61] br[61] wl[51] vdd gnd cell_6t
Xbit_r52_c61 bl[61] br[61] wl[52] vdd gnd cell_6t
Xbit_r53_c61 bl[61] br[61] wl[53] vdd gnd cell_6t
Xbit_r54_c61 bl[61] br[61] wl[54] vdd gnd cell_6t
Xbit_r55_c61 bl[61] br[61] wl[55] vdd gnd cell_6t
Xbit_r56_c61 bl[61] br[61] wl[56] vdd gnd cell_6t
Xbit_r57_c61 bl[61] br[61] wl[57] vdd gnd cell_6t
Xbit_r58_c61 bl[61] br[61] wl[58] vdd gnd cell_6t
Xbit_r59_c61 bl[61] br[61] wl[59] vdd gnd cell_6t
Xbit_r60_c61 bl[61] br[61] wl[60] vdd gnd cell_6t
Xbit_r61_c61 bl[61] br[61] wl[61] vdd gnd cell_6t
Xbit_r62_c61 bl[61] br[61] wl[62] vdd gnd cell_6t
Xbit_r63_c61 bl[61] br[61] wl[63] vdd gnd cell_6t
Xbit_r64_c61 bl[61] br[61] wl[64] vdd gnd cell_6t
Xbit_r65_c61 bl[61] br[61] wl[65] vdd gnd cell_6t
Xbit_r66_c61 bl[61] br[61] wl[66] vdd gnd cell_6t
Xbit_r67_c61 bl[61] br[61] wl[67] vdd gnd cell_6t
Xbit_r68_c61 bl[61] br[61] wl[68] vdd gnd cell_6t
Xbit_r69_c61 bl[61] br[61] wl[69] vdd gnd cell_6t
Xbit_r70_c61 bl[61] br[61] wl[70] vdd gnd cell_6t
Xbit_r71_c61 bl[61] br[61] wl[71] vdd gnd cell_6t
Xbit_r72_c61 bl[61] br[61] wl[72] vdd gnd cell_6t
Xbit_r73_c61 bl[61] br[61] wl[73] vdd gnd cell_6t
Xbit_r74_c61 bl[61] br[61] wl[74] vdd gnd cell_6t
Xbit_r75_c61 bl[61] br[61] wl[75] vdd gnd cell_6t
Xbit_r76_c61 bl[61] br[61] wl[76] vdd gnd cell_6t
Xbit_r77_c61 bl[61] br[61] wl[77] vdd gnd cell_6t
Xbit_r78_c61 bl[61] br[61] wl[78] vdd gnd cell_6t
Xbit_r79_c61 bl[61] br[61] wl[79] vdd gnd cell_6t
Xbit_r80_c61 bl[61] br[61] wl[80] vdd gnd cell_6t
Xbit_r81_c61 bl[61] br[61] wl[81] vdd gnd cell_6t
Xbit_r82_c61 bl[61] br[61] wl[82] vdd gnd cell_6t
Xbit_r83_c61 bl[61] br[61] wl[83] vdd gnd cell_6t
Xbit_r84_c61 bl[61] br[61] wl[84] vdd gnd cell_6t
Xbit_r85_c61 bl[61] br[61] wl[85] vdd gnd cell_6t
Xbit_r86_c61 bl[61] br[61] wl[86] vdd gnd cell_6t
Xbit_r87_c61 bl[61] br[61] wl[87] vdd gnd cell_6t
Xbit_r88_c61 bl[61] br[61] wl[88] vdd gnd cell_6t
Xbit_r89_c61 bl[61] br[61] wl[89] vdd gnd cell_6t
Xbit_r90_c61 bl[61] br[61] wl[90] vdd gnd cell_6t
Xbit_r91_c61 bl[61] br[61] wl[91] vdd gnd cell_6t
Xbit_r92_c61 bl[61] br[61] wl[92] vdd gnd cell_6t
Xbit_r93_c61 bl[61] br[61] wl[93] vdd gnd cell_6t
Xbit_r94_c61 bl[61] br[61] wl[94] vdd gnd cell_6t
Xbit_r95_c61 bl[61] br[61] wl[95] vdd gnd cell_6t
Xbit_r96_c61 bl[61] br[61] wl[96] vdd gnd cell_6t
Xbit_r97_c61 bl[61] br[61] wl[97] vdd gnd cell_6t
Xbit_r98_c61 bl[61] br[61] wl[98] vdd gnd cell_6t
Xbit_r99_c61 bl[61] br[61] wl[99] vdd gnd cell_6t
Xbit_r100_c61 bl[61] br[61] wl[100] vdd gnd cell_6t
Xbit_r101_c61 bl[61] br[61] wl[101] vdd gnd cell_6t
Xbit_r102_c61 bl[61] br[61] wl[102] vdd gnd cell_6t
Xbit_r103_c61 bl[61] br[61] wl[103] vdd gnd cell_6t
Xbit_r104_c61 bl[61] br[61] wl[104] vdd gnd cell_6t
Xbit_r105_c61 bl[61] br[61] wl[105] vdd gnd cell_6t
Xbit_r106_c61 bl[61] br[61] wl[106] vdd gnd cell_6t
Xbit_r107_c61 bl[61] br[61] wl[107] vdd gnd cell_6t
Xbit_r108_c61 bl[61] br[61] wl[108] vdd gnd cell_6t
Xbit_r109_c61 bl[61] br[61] wl[109] vdd gnd cell_6t
Xbit_r110_c61 bl[61] br[61] wl[110] vdd gnd cell_6t
Xbit_r111_c61 bl[61] br[61] wl[111] vdd gnd cell_6t
Xbit_r112_c61 bl[61] br[61] wl[112] vdd gnd cell_6t
Xbit_r113_c61 bl[61] br[61] wl[113] vdd gnd cell_6t
Xbit_r114_c61 bl[61] br[61] wl[114] vdd gnd cell_6t
Xbit_r115_c61 bl[61] br[61] wl[115] vdd gnd cell_6t
Xbit_r116_c61 bl[61] br[61] wl[116] vdd gnd cell_6t
Xbit_r117_c61 bl[61] br[61] wl[117] vdd gnd cell_6t
Xbit_r118_c61 bl[61] br[61] wl[118] vdd gnd cell_6t
Xbit_r119_c61 bl[61] br[61] wl[119] vdd gnd cell_6t
Xbit_r120_c61 bl[61] br[61] wl[120] vdd gnd cell_6t
Xbit_r121_c61 bl[61] br[61] wl[121] vdd gnd cell_6t
Xbit_r122_c61 bl[61] br[61] wl[122] vdd gnd cell_6t
Xbit_r123_c61 bl[61] br[61] wl[123] vdd gnd cell_6t
Xbit_r124_c61 bl[61] br[61] wl[124] vdd gnd cell_6t
Xbit_r125_c61 bl[61] br[61] wl[125] vdd gnd cell_6t
Xbit_r126_c61 bl[61] br[61] wl[126] vdd gnd cell_6t
Xbit_r127_c61 bl[61] br[61] wl[127] vdd gnd cell_6t
Xbit_r128_c61 bl[61] br[61] wl[128] vdd gnd cell_6t
Xbit_r129_c61 bl[61] br[61] wl[129] vdd gnd cell_6t
Xbit_r130_c61 bl[61] br[61] wl[130] vdd gnd cell_6t
Xbit_r131_c61 bl[61] br[61] wl[131] vdd gnd cell_6t
Xbit_r132_c61 bl[61] br[61] wl[132] vdd gnd cell_6t
Xbit_r133_c61 bl[61] br[61] wl[133] vdd gnd cell_6t
Xbit_r134_c61 bl[61] br[61] wl[134] vdd gnd cell_6t
Xbit_r135_c61 bl[61] br[61] wl[135] vdd gnd cell_6t
Xbit_r136_c61 bl[61] br[61] wl[136] vdd gnd cell_6t
Xbit_r137_c61 bl[61] br[61] wl[137] vdd gnd cell_6t
Xbit_r138_c61 bl[61] br[61] wl[138] vdd gnd cell_6t
Xbit_r139_c61 bl[61] br[61] wl[139] vdd gnd cell_6t
Xbit_r140_c61 bl[61] br[61] wl[140] vdd gnd cell_6t
Xbit_r141_c61 bl[61] br[61] wl[141] vdd gnd cell_6t
Xbit_r142_c61 bl[61] br[61] wl[142] vdd gnd cell_6t
Xbit_r143_c61 bl[61] br[61] wl[143] vdd gnd cell_6t
Xbit_r144_c61 bl[61] br[61] wl[144] vdd gnd cell_6t
Xbit_r145_c61 bl[61] br[61] wl[145] vdd gnd cell_6t
Xbit_r146_c61 bl[61] br[61] wl[146] vdd gnd cell_6t
Xbit_r147_c61 bl[61] br[61] wl[147] vdd gnd cell_6t
Xbit_r148_c61 bl[61] br[61] wl[148] vdd gnd cell_6t
Xbit_r149_c61 bl[61] br[61] wl[149] vdd gnd cell_6t
Xbit_r150_c61 bl[61] br[61] wl[150] vdd gnd cell_6t
Xbit_r151_c61 bl[61] br[61] wl[151] vdd gnd cell_6t
Xbit_r152_c61 bl[61] br[61] wl[152] vdd gnd cell_6t
Xbit_r153_c61 bl[61] br[61] wl[153] vdd gnd cell_6t
Xbit_r154_c61 bl[61] br[61] wl[154] vdd gnd cell_6t
Xbit_r155_c61 bl[61] br[61] wl[155] vdd gnd cell_6t
Xbit_r156_c61 bl[61] br[61] wl[156] vdd gnd cell_6t
Xbit_r157_c61 bl[61] br[61] wl[157] vdd gnd cell_6t
Xbit_r158_c61 bl[61] br[61] wl[158] vdd gnd cell_6t
Xbit_r159_c61 bl[61] br[61] wl[159] vdd gnd cell_6t
Xbit_r160_c61 bl[61] br[61] wl[160] vdd gnd cell_6t
Xbit_r161_c61 bl[61] br[61] wl[161] vdd gnd cell_6t
Xbit_r162_c61 bl[61] br[61] wl[162] vdd gnd cell_6t
Xbit_r163_c61 bl[61] br[61] wl[163] vdd gnd cell_6t
Xbit_r164_c61 bl[61] br[61] wl[164] vdd gnd cell_6t
Xbit_r165_c61 bl[61] br[61] wl[165] vdd gnd cell_6t
Xbit_r166_c61 bl[61] br[61] wl[166] vdd gnd cell_6t
Xbit_r167_c61 bl[61] br[61] wl[167] vdd gnd cell_6t
Xbit_r168_c61 bl[61] br[61] wl[168] vdd gnd cell_6t
Xbit_r169_c61 bl[61] br[61] wl[169] vdd gnd cell_6t
Xbit_r170_c61 bl[61] br[61] wl[170] vdd gnd cell_6t
Xbit_r171_c61 bl[61] br[61] wl[171] vdd gnd cell_6t
Xbit_r172_c61 bl[61] br[61] wl[172] vdd gnd cell_6t
Xbit_r173_c61 bl[61] br[61] wl[173] vdd gnd cell_6t
Xbit_r174_c61 bl[61] br[61] wl[174] vdd gnd cell_6t
Xbit_r175_c61 bl[61] br[61] wl[175] vdd gnd cell_6t
Xbit_r176_c61 bl[61] br[61] wl[176] vdd gnd cell_6t
Xbit_r177_c61 bl[61] br[61] wl[177] vdd gnd cell_6t
Xbit_r178_c61 bl[61] br[61] wl[178] vdd gnd cell_6t
Xbit_r179_c61 bl[61] br[61] wl[179] vdd gnd cell_6t
Xbit_r180_c61 bl[61] br[61] wl[180] vdd gnd cell_6t
Xbit_r181_c61 bl[61] br[61] wl[181] vdd gnd cell_6t
Xbit_r182_c61 bl[61] br[61] wl[182] vdd gnd cell_6t
Xbit_r183_c61 bl[61] br[61] wl[183] vdd gnd cell_6t
Xbit_r184_c61 bl[61] br[61] wl[184] vdd gnd cell_6t
Xbit_r185_c61 bl[61] br[61] wl[185] vdd gnd cell_6t
Xbit_r186_c61 bl[61] br[61] wl[186] vdd gnd cell_6t
Xbit_r187_c61 bl[61] br[61] wl[187] vdd gnd cell_6t
Xbit_r188_c61 bl[61] br[61] wl[188] vdd gnd cell_6t
Xbit_r189_c61 bl[61] br[61] wl[189] vdd gnd cell_6t
Xbit_r190_c61 bl[61] br[61] wl[190] vdd gnd cell_6t
Xbit_r191_c61 bl[61] br[61] wl[191] vdd gnd cell_6t
Xbit_r192_c61 bl[61] br[61] wl[192] vdd gnd cell_6t
Xbit_r193_c61 bl[61] br[61] wl[193] vdd gnd cell_6t
Xbit_r194_c61 bl[61] br[61] wl[194] vdd gnd cell_6t
Xbit_r195_c61 bl[61] br[61] wl[195] vdd gnd cell_6t
Xbit_r196_c61 bl[61] br[61] wl[196] vdd gnd cell_6t
Xbit_r197_c61 bl[61] br[61] wl[197] vdd gnd cell_6t
Xbit_r198_c61 bl[61] br[61] wl[198] vdd gnd cell_6t
Xbit_r199_c61 bl[61] br[61] wl[199] vdd gnd cell_6t
Xbit_r200_c61 bl[61] br[61] wl[200] vdd gnd cell_6t
Xbit_r201_c61 bl[61] br[61] wl[201] vdd gnd cell_6t
Xbit_r202_c61 bl[61] br[61] wl[202] vdd gnd cell_6t
Xbit_r203_c61 bl[61] br[61] wl[203] vdd gnd cell_6t
Xbit_r204_c61 bl[61] br[61] wl[204] vdd gnd cell_6t
Xbit_r205_c61 bl[61] br[61] wl[205] vdd gnd cell_6t
Xbit_r206_c61 bl[61] br[61] wl[206] vdd gnd cell_6t
Xbit_r207_c61 bl[61] br[61] wl[207] vdd gnd cell_6t
Xbit_r208_c61 bl[61] br[61] wl[208] vdd gnd cell_6t
Xbit_r209_c61 bl[61] br[61] wl[209] vdd gnd cell_6t
Xbit_r210_c61 bl[61] br[61] wl[210] vdd gnd cell_6t
Xbit_r211_c61 bl[61] br[61] wl[211] vdd gnd cell_6t
Xbit_r212_c61 bl[61] br[61] wl[212] vdd gnd cell_6t
Xbit_r213_c61 bl[61] br[61] wl[213] vdd gnd cell_6t
Xbit_r214_c61 bl[61] br[61] wl[214] vdd gnd cell_6t
Xbit_r215_c61 bl[61] br[61] wl[215] vdd gnd cell_6t
Xbit_r216_c61 bl[61] br[61] wl[216] vdd gnd cell_6t
Xbit_r217_c61 bl[61] br[61] wl[217] vdd gnd cell_6t
Xbit_r218_c61 bl[61] br[61] wl[218] vdd gnd cell_6t
Xbit_r219_c61 bl[61] br[61] wl[219] vdd gnd cell_6t
Xbit_r220_c61 bl[61] br[61] wl[220] vdd gnd cell_6t
Xbit_r221_c61 bl[61] br[61] wl[221] vdd gnd cell_6t
Xbit_r222_c61 bl[61] br[61] wl[222] vdd gnd cell_6t
Xbit_r223_c61 bl[61] br[61] wl[223] vdd gnd cell_6t
Xbit_r224_c61 bl[61] br[61] wl[224] vdd gnd cell_6t
Xbit_r225_c61 bl[61] br[61] wl[225] vdd gnd cell_6t
Xbit_r226_c61 bl[61] br[61] wl[226] vdd gnd cell_6t
Xbit_r227_c61 bl[61] br[61] wl[227] vdd gnd cell_6t
Xbit_r228_c61 bl[61] br[61] wl[228] vdd gnd cell_6t
Xbit_r229_c61 bl[61] br[61] wl[229] vdd gnd cell_6t
Xbit_r230_c61 bl[61] br[61] wl[230] vdd gnd cell_6t
Xbit_r231_c61 bl[61] br[61] wl[231] vdd gnd cell_6t
Xbit_r232_c61 bl[61] br[61] wl[232] vdd gnd cell_6t
Xbit_r233_c61 bl[61] br[61] wl[233] vdd gnd cell_6t
Xbit_r234_c61 bl[61] br[61] wl[234] vdd gnd cell_6t
Xbit_r235_c61 bl[61] br[61] wl[235] vdd gnd cell_6t
Xbit_r236_c61 bl[61] br[61] wl[236] vdd gnd cell_6t
Xbit_r237_c61 bl[61] br[61] wl[237] vdd gnd cell_6t
Xbit_r238_c61 bl[61] br[61] wl[238] vdd gnd cell_6t
Xbit_r239_c61 bl[61] br[61] wl[239] vdd gnd cell_6t
Xbit_r240_c61 bl[61] br[61] wl[240] vdd gnd cell_6t
Xbit_r241_c61 bl[61] br[61] wl[241] vdd gnd cell_6t
Xbit_r242_c61 bl[61] br[61] wl[242] vdd gnd cell_6t
Xbit_r243_c61 bl[61] br[61] wl[243] vdd gnd cell_6t
Xbit_r244_c61 bl[61] br[61] wl[244] vdd gnd cell_6t
Xbit_r245_c61 bl[61] br[61] wl[245] vdd gnd cell_6t
Xbit_r246_c61 bl[61] br[61] wl[246] vdd gnd cell_6t
Xbit_r247_c61 bl[61] br[61] wl[247] vdd gnd cell_6t
Xbit_r248_c61 bl[61] br[61] wl[248] vdd gnd cell_6t
Xbit_r249_c61 bl[61] br[61] wl[249] vdd gnd cell_6t
Xbit_r250_c61 bl[61] br[61] wl[250] vdd gnd cell_6t
Xbit_r251_c61 bl[61] br[61] wl[251] vdd gnd cell_6t
Xbit_r252_c61 bl[61] br[61] wl[252] vdd gnd cell_6t
Xbit_r253_c61 bl[61] br[61] wl[253] vdd gnd cell_6t
Xbit_r254_c61 bl[61] br[61] wl[254] vdd gnd cell_6t
Xbit_r255_c61 bl[61] br[61] wl[255] vdd gnd cell_6t
Xbit_r256_c61 bl[61] br[61] wl[256] vdd gnd cell_6t
Xbit_r257_c61 bl[61] br[61] wl[257] vdd gnd cell_6t
Xbit_r258_c61 bl[61] br[61] wl[258] vdd gnd cell_6t
Xbit_r259_c61 bl[61] br[61] wl[259] vdd gnd cell_6t
Xbit_r260_c61 bl[61] br[61] wl[260] vdd gnd cell_6t
Xbit_r261_c61 bl[61] br[61] wl[261] vdd gnd cell_6t
Xbit_r262_c61 bl[61] br[61] wl[262] vdd gnd cell_6t
Xbit_r263_c61 bl[61] br[61] wl[263] vdd gnd cell_6t
Xbit_r264_c61 bl[61] br[61] wl[264] vdd gnd cell_6t
Xbit_r265_c61 bl[61] br[61] wl[265] vdd gnd cell_6t
Xbit_r266_c61 bl[61] br[61] wl[266] vdd gnd cell_6t
Xbit_r267_c61 bl[61] br[61] wl[267] vdd gnd cell_6t
Xbit_r268_c61 bl[61] br[61] wl[268] vdd gnd cell_6t
Xbit_r269_c61 bl[61] br[61] wl[269] vdd gnd cell_6t
Xbit_r270_c61 bl[61] br[61] wl[270] vdd gnd cell_6t
Xbit_r271_c61 bl[61] br[61] wl[271] vdd gnd cell_6t
Xbit_r272_c61 bl[61] br[61] wl[272] vdd gnd cell_6t
Xbit_r273_c61 bl[61] br[61] wl[273] vdd gnd cell_6t
Xbit_r274_c61 bl[61] br[61] wl[274] vdd gnd cell_6t
Xbit_r275_c61 bl[61] br[61] wl[275] vdd gnd cell_6t
Xbit_r276_c61 bl[61] br[61] wl[276] vdd gnd cell_6t
Xbit_r277_c61 bl[61] br[61] wl[277] vdd gnd cell_6t
Xbit_r278_c61 bl[61] br[61] wl[278] vdd gnd cell_6t
Xbit_r279_c61 bl[61] br[61] wl[279] vdd gnd cell_6t
Xbit_r280_c61 bl[61] br[61] wl[280] vdd gnd cell_6t
Xbit_r281_c61 bl[61] br[61] wl[281] vdd gnd cell_6t
Xbit_r282_c61 bl[61] br[61] wl[282] vdd gnd cell_6t
Xbit_r283_c61 bl[61] br[61] wl[283] vdd gnd cell_6t
Xbit_r284_c61 bl[61] br[61] wl[284] vdd gnd cell_6t
Xbit_r285_c61 bl[61] br[61] wl[285] vdd gnd cell_6t
Xbit_r286_c61 bl[61] br[61] wl[286] vdd gnd cell_6t
Xbit_r287_c61 bl[61] br[61] wl[287] vdd gnd cell_6t
Xbit_r288_c61 bl[61] br[61] wl[288] vdd gnd cell_6t
Xbit_r289_c61 bl[61] br[61] wl[289] vdd gnd cell_6t
Xbit_r290_c61 bl[61] br[61] wl[290] vdd gnd cell_6t
Xbit_r291_c61 bl[61] br[61] wl[291] vdd gnd cell_6t
Xbit_r292_c61 bl[61] br[61] wl[292] vdd gnd cell_6t
Xbit_r293_c61 bl[61] br[61] wl[293] vdd gnd cell_6t
Xbit_r294_c61 bl[61] br[61] wl[294] vdd gnd cell_6t
Xbit_r295_c61 bl[61] br[61] wl[295] vdd gnd cell_6t
Xbit_r296_c61 bl[61] br[61] wl[296] vdd gnd cell_6t
Xbit_r297_c61 bl[61] br[61] wl[297] vdd gnd cell_6t
Xbit_r298_c61 bl[61] br[61] wl[298] vdd gnd cell_6t
Xbit_r299_c61 bl[61] br[61] wl[299] vdd gnd cell_6t
Xbit_r300_c61 bl[61] br[61] wl[300] vdd gnd cell_6t
Xbit_r301_c61 bl[61] br[61] wl[301] vdd gnd cell_6t
Xbit_r302_c61 bl[61] br[61] wl[302] vdd gnd cell_6t
Xbit_r303_c61 bl[61] br[61] wl[303] vdd gnd cell_6t
Xbit_r304_c61 bl[61] br[61] wl[304] vdd gnd cell_6t
Xbit_r305_c61 bl[61] br[61] wl[305] vdd gnd cell_6t
Xbit_r306_c61 bl[61] br[61] wl[306] vdd gnd cell_6t
Xbit_r307_c61 bl[61] br[61] wl[307] vdd gnd cell_6t
Xbit_r308_c61 bl[61] br[61] wl[308] vdd gnd cell_6t
Xbit_r309_c61 bl[61] br[61] wl[309] vdd gnd cell_6t
Xbit_r310_c61 bl[61] br[61] wl[310] vdd gnd cell_6t
Xbit_r311_c61 bl[61] br[61] wl[311] vdd gnd cell_6t
Xbit_r312_c61 bl[61] br[61] wl[312] vdd gnd cell_6t
Xbit_r313_c61 bl[61] br[61] wl[313] vdd gnd cell_6t
Xbit_r314_c61 bl[61] br[61] wl[314] vdd gnd cell_6t
Xbit_r315_c61 bl[61] br[61] wl[315] vdd gnd cell_6t
Xbit_r316_c61 bl[61] br[61] wl[316] vdd gnd cell_6t
Xbit_r317_c61 bl[61] br[61] wl[317] vdd gnd cell_6t
Xbit_r318_c61 bl[61] br[61] wl[318] vdd gnd cell_6t
Xbit_r319_c61 bl[61] br[61] wl[319] vdd gnd cell_6t
Xbit_r320_c61 bl[61] br[61] wl[320] vdd gnd cell_6t
Xbit_r321_c61 bl[61] br[61] wl[321] vdd gnd cell_6t
Xbit_r322_c61 bl[61] br[61] wl[322] vdd gnd cell_6t
Xbit_r323_c61 bl[61] br[61] wl[323] vdd gnd cell_6t
Xbit_r324_c61 bl[61] br[61] wl[324] vdd gnd cell_6t
Xbit_r325_c61 bl[61] br[61] wl[325] vdd gnd cell_6t
Xbit_r326_c61 bl[61] br[61] wl[326] vdd gnd cell_6t
Xbit_r327_c61 bl[61] br[61] wl[327] vdd gnd cell_6t
Xbit_r328_c61 bl[61] br[61] wl[328] vdd gnd cell_6t
Xbit_r329_c61 bl[61] br[61] wl[329] vdd gnd cell_6t
Xbit_r330_c61 bl[61] br[61] wl[330] vdd gnd cell_6t
Xbit_r331_c61 bl[61] br[61] wl[331] vdd gnd cell_6t
Xbit_r332_c61 bl[61] br[61] wl[332] vdd gnd cell_6t
Xbit_r333_c61 bl[61] br[61] wl[333] vdd gnd cell_6t
Xbit_r334_c61 bl[61] br[61] wl[334] vdd gnd cell_6t
Xbit_r335_c61 bl[61] br[61] wl[335] vdd gnd cell_6t
Xbit_r336_c61 bl[61] br[61] wl[336] vdd gnd cell_6t
Xbit_r337_c61 bl[61] br[61] wl[337] vdd gnd cell_6t
Xbit_r338_c61 bl[61] br[61] wl[338] vdd gnd cell_6t
Xbit_r339_c61 bl[61] br[61] wl[339] vdd gnd cell_6t
Xbit_r340_c61 bl[61] br[61] wl[340] vdd gnd cell_6t
Xbit_r341_c61 bl[61] br[61] wl[341] vdd gnd cell_6t
Xbit_r342_c61 bl[61] br[61] wl[342] vdd gnd cell_6t
Xbit_r343_c61 bl[61] br[61] wl[343] vdd gnd cell_6t
Xbit_r344_c61 bl[61] br[61] wl[344] vdd gnd cell_6t
Xbit_r345_c61 bl[61] br[61] wl[345] vdd gnd cell_6t
Xbit_r346_c61 bl[61] br[61] wl[346] vdd gnd cell_6t
Xbit_r347_c61 bl[61] br[61] wl[347] vdd gnd cell_6t
Xbit_r348_c61 bl[61] br[61] wl[348] vdd gnd cell_6t
Xbit_r349_c61 bl[61] br[61] wl[349] vdd gnd cell_6t
Xbit_r350_c61 bl[61] br[61] wl[350] vdd gnd cell_6t
Xbit_r351_c61 bl[61] br[61] wl[351] vdd gnd cell_6t
Xbit_r352_c61 bl[61] br[61] wl[352] vdd gnd cell_6t
Xbit_r353_c61 bl[61] br[61] wl[353] vdd gnd cell_6t
Xbit_r354_c61 bl[61] br[61] wl[354] vdd gnd cell_6t
Xbit_r355_c61 bl[61] br[61] wl[355] vdd gnd cell_6t
Xbit_r356_c61 bl[61] br[61] wl[356] vdd gnd cell_6t
Xbit_r357_c61 bl[61] br[61] wl[357] vdd gnd cell_6t
Xbit_r358_c61 bl[61] br[61] wl[358] vdd gnd cell_6t
Xbit_r359_c61 bl[61] br[61] wl[359] vdd gnd cell_6t
Xbit_r360_c61 bl[61] br[61] wl[360] vdd gnd cell_6t
Xbit_r361_c61 bl[61] br[61] wl[361] vdd gnd cell_6t
Xbit_r362_c61 bl[61] br[61] wl[362] vdd gnd cell_6t
Xbit_r363_c61 bl[61] br[61] wl[363] vdd gnd cell_6t
Xbit_r364_c61 bl[61] br[61] wl[364] vdd gnd cell_6t
Xbit_r365_c61 bl[61] br[61] wl[365] vdd gnd cell_6t
Xbit_r366_c61 bl[61] br[61] wl[366] vdd gnd cell_6t
Xbit_r367_c61 bl[61] br[61] wl[367] vdd gnd cell_6t
Xbit_r368_c61 bl[61] br[61] wl[368] vdd gnd cell_6t
Xbit_r369_c61 bl[61] br[61] wl[369] vdd gnd cell_6t
Xbit_r370_c61 bl[61] br[61] wl[370] vdd gnd cell_6t
Xbit_r371_c61 bl[61] br[61] wl[371] vdd gnd cell_6t
Xbit_r372_c61 bl[61] br[61] wl[372] vdd gnd cell_6t
Xbit_r373_c61 bl[61] br[61] wl[373] vdd gnd cell_6t
Xbit_r374_c61 bl[61] br[61] wl[374] vdd gnd cell_6t
Xbit_r375_c61 bl[61] br[61] wl[375] vdd gnd cell_6t
Xbit_r376_c61 bl[61] br[61] wl[376] vdd gnd cell_6t
Xbit_r377_c61 bl[61] br[61] wl[377] vdd gnd cell_6t
Xbit_r378_c61 bl[61] br[61] wl[378] vdd gnd cell_6t
Xbit_r379_c61 bl[61] br[61] wl[379] vdd gnd cell_6t
Xbit_r380_c61 bl[61] br[61] wl[380] vdd gnd cell_6t
Xbit_r381_c61 bl[61] br[61] wl[381] vdd gnd cell_6t
Xbit_r382_c61 bl[61] br[61] wl[382] vdd gnd cell_6t
Xbit_r383_c61 bl[61] br[61] wl[383] vdd gnd cell_6t
Xbit_r384_c61 bl[61] br[61] wl[384] vdd gnd cell_6t
Xbit_r385_c61 bl[61] br[61] wl[385] vdd gnd cell_6t
Xbit_r386_c61 bl[61] br[61] wl[386] vdd gnd cell_6t
Xbit_r387_c61 bl[61] br[61] wl[387] vdd gnd cell_6t
Xbit_r388_c61 bl[61] br[61] wl[388] vdd gnd cell_6t
Xbit_r389_c61 bl[61] br[61] wl[389] vdd gnd cell_6t
Xbit_r390_c61 bl[61] br[61] wl[390] vdd gnd cell_6t
Xbit_r391_c61 bl[61] br[61] wl[391] vdd gnd cell_6t
Xbit_r392_c61 bl[61] br[61] wl[392] vdd gnd cell_6t
Xbit_r393_c61 bl[61] br[61] wl[393] vdd gnd cell_6t
Xbit_r394_c61 bl[61] br[61] wl[394] vdd gnd cell_6t
Xbit_r395_c61 bl[61] br[61] wl[395] vdd gnd cell_6t
Xbit_r396_c61 bl[61] br[61] wl[396] vdd gnd cell_6t
Xbit_r397_c61 bl[61] br[61] wl[397] vdd gnd cell_6t
Xbit_r398_c61 bl[61] br[61] wl[398] vdd gnd cell_6t
Xbit_r399_c61 bl[61] br[61] wl[399] vdd gnd cell_6t
Xbit_r400_c61 bl[61] br[61] wl[400] vdd gnd cell_6t
Xbit_r401_c61 bl[61] br[61] wl[401] vdd gnd cell_6t
Xbit_r402_c61 bl[61] br[61] wl[402] vdd gnd cell_6t
Xbit_r403_c61 bl[61] br[61] wl[403] vdd gnd cell_6t
Xbit_r404_c61 bl[61] br[61] wl[404] vdd gnd cell_6t
Xbit_r405_c61 bl[61] br[61] wl[405] vdd gnd cell_6t
Xbit_r406_c61 bl[61] br[61] wl[406] vdd gnd cell_6t
Xbit_r407_c61 bl[61] br[61] wl[407] vdd gnd cell_6t
Xbit_r408_c61 bl[61] br[61] wl[408] vdd gnd cell_6t
Xbit_r409_c61 bl[61] br[61] wl[409] vdd gnd cell_6t
Xbit_r410_c61 bl[61] br[61] wl[410] vdd gnd cell_6t
Xbit_r411_c61 bl[61] br[61] wl[411] vdd gnd cell_6t
Xbit_r412_c61 bl[61] br[61] wl[412] vdd gnd cell_6t
Xbit_r413_c61 bl[61] br[61] wl[413] vdd gnd cell_6t
Xbit_r414_c61 bl[61] br[61] wl[414] vdd gnd cell_6t
Xbit_r415_c61 bl[61] br[61] wl[415] vdd gnd cell_6t
Xbit_r416_c61 bl[61] br[61] wl[416] vdd gnd cell_6t
Xbit_r417_c61 bl[61] br[61] wl[417] vdd gnd cell_6t
Xbit_r418_c61 bl[61] br[61] wl[418] vdd gnd cell_6t
Xbit_r419_c61 bl[61] br[61] wl[419] vdd gnd cell_6t
Xbit_r420_c61 bl[61] br[61] wl[420] vdd gnd cell_6t
Xbit_r421_c61 bl[61] br[61] wl[421] vdd gnd cell_6t
Xbit_r422_c61 bl[61] br[61] wl[422] vdd gnd cell_6t
Xbit_r423_c61 bl[61] br[61] wl[423] vdd gnd cell_6t
Xbit_r424_c61 bl[61] br[61] wl[424] vdd gnd cell_6t
Xbit_r425_c61 bl[61] br[61] wl[425] vdd gnd cell_6t
Xbit_r426_c61 bl[61] br[61] wl[426] vdd gnd cell_6t
Xbit_r427_c61 bl[61] br[61] wl[427] vdd gnd cell_6t
Xbit_r428_c61 bl[61] br[61] wl[428] vdd gnd cell_6t
Xbit_r429_c61 bl[61] br[61] wl[429] vdd gnd cell_6t
Xbit_r430_c61 bl[61] br[61] wl[430] vdd gnd cell_6t
Xbit_r431_c61 bl[61] br[61] wl[431] vdd gnd cell_6t
Xbit_r432_c61 bl[61] br[61] wl[432] vdd gnd cell_6t
Xbit_r433_c61 bl[61] br[61] wl[433] vdd gnd cell_6t
Xbit_r434_c61 bl[61] br[61] wl[434] vdd gnd cell_6t
Xbit_r435_c61 bl[61] br[61] wl[435] vdd gnd cell_6t
Xbit_r436_c61 bl[61] br[61] wl[436] vdd gnd cell_6t
Xbit_r437_c61 bl[61] br[61] wl[437] vdd gnd cell_6t
Xbit_r438_c61 bl[61] br[61] wl[438] vdd gnd cell_6t
Xbit_r439_c61 bl[61] br[61] wl[439] vdd gnd cell_6t
Xbit_r440_c61 bl[61] br[61] wl[440] vdd gnd cell_6t
Xbit_r441_c61 bl[61] br[61] wl[441] vdd gnd cell_6t
Xbit_r442_c61 bl[61] br[61] wl[442] vdd gnd cell_6t
Xbit_r443_c61 bl[61] br[61] wl[443] vdd gnd cell_6t
Xbit_r444_c61 bl[61] br[61] wl[444] vdd gnd cell_6t
Xbit_r445_c61 bl[61] br[61] wl[445] vdd gnd cell_6t
Xbit_r446_c61 bl[61] br[61] wl[446] vdd gnd cell_6t
Xbit_r447_c61 bl[61] br[61] wl[447] vdd gnd cell_6t
Xbit_r448_c61 bl[61] br[61] wl[448] vdd gnd cell_6t
Xbit_r449_c61 bl[61] br[61] wl[449] vdd gnd cell_6t
Xbit_r450_c61 bl[61] br[61] wl[450] vdd gnd cell_6t
Xbit_r451_c61 bl[61] br[61] wl[451] vdd gnd cell_6t
Xbit_r452_c61 bl[61] br[61] wl[452] vdd gnd cell_6t
Xbit_r453_c61 bl[61] br[61] wl[453] vdd gnd cell_6t
Xbit_r454_c61 bl[61] br[61] wl[454] vdd gnd cell_6t
Xbit_r455_c61 bl[61] br[61] wl[455] vdd gnd cell_6t
Xbit_r456_c61 bl[61] br[61] wl[456] vdd gnd cell_6t
Xbit_r457_c61 bl[61] br[61] wl[457] vdd gnd cell_6t
Xbit_r458_c61 bl[61] br[61] wl[458] vdd gnd cell_6t
Xbit_r459_c61 bl[61] br[61] wl[459] vdd gnd cell_6t
Xbit_r460_c61 bl[61] br[61] wl[460] vdd gnd cell_6t
Xbit_r461_c61 bl[61] br[61] wl[461] vdd gnd cell_6t
Xbit_r462_c61 bl[61] br[61] wl[462] vdd gnd cell_6t
Xbit_r463_c61 bl[61] br[61] wl[463] vdd gnd cell_6t
Xbit_r464_c61 bl[61] br[61] wl[464] vdd gnd cell_6t
Xbit_r465_c61 bl[61] br[61] wl[465] vdd gnd cell_6t
Xbit_r466_c61 bl[61] br[61] wl[466] vdd gnd cell_6t
Xbit_r467_c61 bl[61] br[61] wl[467] vdd gnd cell_6t
Xbit_r468_c61 bl[61] br[61] wl[468] vdd gnd cell_6t
Xbit_r469_c61 bl[61] br[61] wl[469] vdd gnd cell_6t
Xbit_r470_c61 bl[61] br[61] wl[470] vdd gnd cell_6t
Xbit_r471_c61 bl[61] br[61] wl[471] vdd gnd cell_6t
Xbit_r472_c61 bl[61] br[61] wl[472] vdd gnd cell_6t
Xbit_r473_c61 bl[61] br[61] wl[473] vdd gnd cell_6t
Xbit_r474_c61 bl[61] br[61] wl[474] vdd gnd cell_6t
Xbit_r475_c61 bl[61] br[61] wl[475] vdd gnd cell_6t
Xbit_r476_c61 bl[61] br[61] wl[476] vdd gnd cell_6t
Xbit_r477_c61 bl[61] br[61] wl[477] vdd gnd cell_6t
Xbit_r478_c61 bl[61] br[61] wl[478] vdd gnd cell_6t
Xbit_r479_c61 bl[61] br[61] wl[479] vdd gnd cell_6t
Xbit_r480_c61 bl[61] br[61] wl[480] vdd gnd cell_6t
Xbit_r481_c61 bl[61] br[61] wl[481] vdd gnd cell_6t
Xbit_r482_c61 bl[61] br[61] wl[482] vdd gnd cell_6t
Xbit_r483_c61 bl[61] br[61] wl[483] vdd gnd cell_6t
Xbit_r484_c61 bl[61] br[61] wl[484] vdd gnd cell_6t
Xbit_r485_c61 bl[61] br[61] wl[485] vdd gnd cell_6t
Xbit_r486_c61 bl[61] br[61] wl[486] vdd gnd cell_6t
Xbit_r487_c61 bl[61] br[61] wl[487] vdd gnd cell_6t
Xbit_r488_c61 bl[61] br[61] wl[488] vdd gnd cell_6t
Xbit_r489_c61 bl[61] br[61] wl[489] vdd gnd cell_6t
Xbit_r490_c61 bl[61] br[61] wl[490] vdd gnd cell_6t
Xbit_r491_c61 bl[61] br[61] wl[491] vdd gnd cell_6t
Xbit_r492_c61 bl[61] br[61] wl[492] vdd gnd cell_6t
Xbit_r493_c61 bl[61] br[61] wl[493] vdd gnd cell_6t
Xbit_r494_c61 bl[61] br[61] wl[494] vdd gnd cell_6t
Xbit_r495_c61 bl[61] br[61] wl[495] vdd gnd cell_6t
Xbit_r496_c61 bl[61] br[61] wl[496] vdd gnd cell_6t
Xbit_r497_c61 bl[61] br[61] wl[497] vdd gnd cell_6t
Xbit_r498_c61 bl[61] br[61] wl[498] vdd gnd cell_6t
Xbit_r499_c61 bl[61] br[61] wl[499] vdd gnd cell_6t
Xbit_r500_c61 bl[61] br[61] wl[500] vdd gnd cell_6t
Xbit_r501_c61 bl[61] br[61] wl[501] vdd gnd cell_6t
Xbit_r502_c61 bl[61] br[61] wl[502] vdd gnd cell_6t
Xbit_r503_c61 bl[61] br[61] wl[503] vdd gnd cell_6t
Xbit_r504_c61 bl[61] br[61] wl[504] vdd gnd cell_6t
Xbit_r505_c61 bl[61] br[61] wl[505] vdd gnd cell_6t
Xbit_r506_c61 bl[61] br[61] wl[506] vdd gnd cell_6t
Xbit_r507_c61 bl[61] br[61] wl[507] vdd gnd cell_6t
Xbit_r508_c61 bl[61] br[61] wl[508] vdd gnd cell_6t
Xbit_r509_c61 bl[61] br[61] wl[509] vdd gnd cell_6t
Xbit_r510_c61 bl[61] br[61] wl[510] vdd gnd cell_6t
Xbit_r511_c61 bl[61] br[61] wl[511] vdd gnd cell_6t
Xbit_r0_c62 bl[62] br[62] wl[0] vdd gnd cell_6t
Xbit_r1_c62 bl[62] br[62] wl[1] vdd gnd cell_6t
Xbit_r2_c62 bl[62] br[62] wl[2] vdd gnd cell_6t
Xbit_r3_c62 bl[62] br[62] wl[3] vdd gnd cell_6t
Xbit_r4_c62 bl[62] br[62] wl[4] vdd gnd cell_6t
Xbit_r5_c62 bl[62] br[62] wl[5] vdd gnd cell_6t
Xbit_r6_c62 bl[62] br[62] wl[6] vdd gnd cell_6t
Xbit_r7_c62 bl[62] br[62] wl[7] vdd gnd cell_6t
Xbit_r8_c62 bl[62] br[62] wl[8] vdd gnd cell_6t
Xbit_r9_c62 bl[62] br[62] wl[9] vdd gnd cell_6t
Xbit_r10_c62 bl[62] br[62] wl[10] vdd gnd cell_6t
Xbit_r11_c62 bl[62] br[62] wl[11] vdd gnd cell_6t
Xbit_r12_c62 bl[62] br[62] wl[12] vdd gnd cell_6t
Xbit_r13_c62 bl[62] br[62] wl[13] vdd gnd cell_6t
Xbit_r14_c62 bl[62] br[62] wl[14] vdd gnd cell_6t
Xbit_r15_c62 bl[62] br[62] wl[15] vdd gnd cell_6t
Xbit_r16_c62 bl[62] br[62] wl[16] vdd gnd cell_6t
Xbit_r17_c62 bl[62] br[62] wl[17] vdd gnd cell_6t
Xbit_r18_c62 bl[62] br[62] wl[18] vdd gnd cell_6t
Xbit_r19_c62 bl[62] br[62] wl[19] vdd gnd cell_6t
Xbit_r20_c62 bl[62] br[62] wl[20] vdd gnd cell_6t
Xbit_r21_c62 bl[62] br[62] wl[21] vdd gnd cell_6t
Xbit_r22_c62 bl[62] br[62] wl[22] vdd gnd cell_6t
Xbit_r23_c62 bl[62] br[62] wl[23] vdd gnd cell_6t
Xbit_r24_c62 bl[62] br[62] wl[24] vdd gnd cell_6t
Xbit_r25_c62 bl[62] br[62] wl[25] vdd gnd cell_6t
Xbit_r26_c62 bl[62] br[62] wl[26] vdd gnd cell_6t
Xbit_r27_c62 bl[62] br[62] wl[27] vdd gnd cell_6t
Xbit_r28_c62 bl[62] br[62] wl[28] vdd gnd cell_6t
Xbit_r29_c62 bl[62] br[62] wl[29] vdd gnd cell_6t
Xbit_r30_c62 bl[62] br[62] wl[30] vdd gnd cell_6t
Xbit_r31_c62 bl[62] br[62] wl[31] vdd gnd cell_6t
Xbit_r32_c62 bl[62] br[62] wl[32] vdd gnd cell_6t
Xbit_r33_c62 bl[62] br[62] wl[33] vdd gnd cell_6t
Xbit_r34_c62 bl[62] br[62] wl[34] vdd gnd cell_6t
Xbit_r35_c62 bl[62] br[62] wl[35] vdd gnd cell_6t
Xbit_r36_c62 bl[62] br[62] wl[36] vdd gnd cell_6t
Xbit_r37_c62 bl[62] br[62] wl[37] vdd gnd cell_6t
Xbit_r38_c62 bl[62] br[62] wl[38] vdd gnd cell_6t
Xbit_r39_c62 bl[62] br[62] wl[39] vdd gnd cell_6t
Xbit_r40_c62 bl[62] br[62] wl[40] vdd gnd cell_6t
Xbit_r41_c62 bl[62] br[62] wl[41] vdd gnd cell_6t
Xbit_r42_c62 bl[62] br[62] wl[42] vdd gnd cell_6t
Xbit_r43_c62 bl[62] br[62] wl[43] vdd gnd cell_6t
Xbit_r44_c62 bl[62] br[62] wl[44] vdd gnd cell_6t
Xbit_r45_c62 bl[62] br[62] wl[45] vdd gnd cell_6t
Xbit_r46_c62 bl[62] br[62] wl[46] vdd gnd cell_6t
Xbit_r47_c62 bl[62] br[62] wl[47] vdd gnd cell_6t
Xbit_r48_c62 bl[62] br[62] wl[48] vdd gnd cell_6t
Xbit_r49_c62 bl[62] br[62] wl[49] vdd gnd cell_6t
Xbit_r50_c62 bl[62] br[62] wl[50] vdd gnd cell_6t
Xbit_r51_c62 bl[62] br[62] wl[51] vdd gnd cell_6t
Xbit_r52_c62 bl[62] br[62] wl[52] vdd gnd cell_6t
Xbit_r53_c62 bl[62] br[62] wl[53] vdd gnd cell_6t
Xbit_r54_c62 bl[62] br[62] wl[54] vdd gnd cell_6t
Xbit_r55_c62 bl[62] br[62] wl[55] vdd gnd cell_6t
Xbit_r56_c62 bl[62] br[62] wl[56] vdd gnd cell_6t
Xbit_r57_c62 bl[62] br[62] wl[57] vdd gnd cell_6t
Xbit_r58_c62 bl[62] br[62] wl[58] vdd gnd cell_6t
Xbit_r59_c62 bl[62] br[62] wl[59] vdd gnd cell_6t
Xbit_r60_c62 bl[62] br[62] wl[60] vdd gnd cell_6t
Xbit_r61_c62 bl[62] br[62] wl[61] vdd gnd cell_6t
Xbit_r62_c62 bl[62] br[62] wl[62] vdd gnd cell_6t
Xbit_r63_c62 bl[62] br[62] wl[63] vdd gnd cell_6t
Xbit_r64_c62 bl[62] br[62] wl[64] vdd gnd cell_6t
Xbit_r65_c62 bl[62] br[62] wl[65] vdd gnd cell_6t
Xbit_r66_c62 bl[62] br[62] wl[66] vdd gnd cell_6t
Xbit_r67_c62 bl[62] br[62] wl[67] vdd gnd cell_6t
Xbit_r68_c62 bl[62] br[62] wl[68] vdd gnd cell_6t
Xbit_r69_c62 bl[62] br[62] wl[69] vdd gnd cell_6t
Xbit_r70_c62 bl[62] br[62] wl[70] vdd gnd cell_6t
Xbit_r71_c62 bl[62] br[62] wl[71] vdd gnd cell_6t
Xbit_r72_c62 bl[62] br[62] wl[72] vdd gnd cell_6t
Xbit_r73_c62 bl[62] br[62] wl[73] vdd gnd cell_6t
Xbit_r74_c62 bl[62] br[62] wl[74] vdd gnd cell_6t
Xbit_r75_c62 bl[62] br[62] wl[75] vdd gnd cell_6t
Xbit_r76_c62 bl[62] br[62] wl[76] vdd gnd cell_6t
Xbit_r77_c62 bl[62] br[62] wl[77] vdd gnd cell_6t
Xbit_r78_c62 bl[62] br[62] wl[78] vdd gnd cell_6t
Xbit_r79_c62 bl[62] br[62] wl[79] vdd gnd cell_6t
Xbit_r80_c62 bl[62] br[62] wl[80] vdd gnd cell_6t
Xbit_r81_c62 bl[62] br[62] wl[81] vdd gnd cell_6t
Xbit_r82_c62 bl[62] br[62] wl[82] vdd gnd cell_6t
Xbit_r83_c62 bl[62] br[62] wl[83] vdd gnd cell_6t
Xbit_r84_c62 bl[62] br[62] wl[84] vdd gnd cell_6t
Xbit_r85_c62 bl[62] br[62] wl[85] vdd gnd cell_6t
Xbit_r86_c62 bl[62] br[62] wl[86] vdd gnd cell_6t
Xbit_r87_c62 bl[62] br[62] wl[87] vdd gnd cell_6t
Xbit_r88_c62 bl[62] br[62] wl[88] vdd gnd cell_6t
Xbit_r89_c62 bl[62] br[62] wl[89] vdd gnd cell_6t
Xbit_r90_c62 bl[62] br[62] wl[90] vdd gnd cell_6t
Xbit_r91_c62 bl[62] br[62] wl[91] vdd gnd cell_6t
Xbit_r92_c62 bl[62] br[62] wl[92] vdd gnd cell_6t
Xbit_r93_c62 bl[62] br[62] wl[93] vdd gnd cell_6t
Xbit_r94_c62 bl[62] br[62] wl[94] vdd gnd cell_6t
Xbit_r95_c62 bl[62] br[62] wl[95] vdd gnd cell_6t
Xbit_r96_c62 bl[62] br[62] wl[96] vdd gnd cell_6t
Xbit_r97_c62 bl[62] br[62] wl[97] vdd gnd cell_6t
Xbit_r98_c62 bl[62] br[62] wl[98] vdd gnd cell_6t
Xbit_r99_c62 bl[62] br[62] wl[99] vdd gnd cell_6t
Xbit_r100_c62 bl[62] br[62] wl[100] vdd gnd cell_6t
Xbit_r101_c62 bl[62] br[62] wl[101] vdd gnd cell_6t
Xbit_r102_c62 bl[62] br[62] wl[102] vdd gnd cell_6t
Xbit_r103_c62 bl[62] br[62] wl[103] vdd gnd cell_6t
Xbit_r104_c62 bl[62] br[62] wl[104] vdd gnd cell_6t
Xbit_r105_c62 bl[62] br[62] wl[105] vdd gnd cell_6t
Xbit_r106_c62 bl[62] br[62] wl[106] vdd gnd cell_6t
Xbit_r107_c62 bl[62] br[62] wl[107] vdd gnd cell_6t
Xbit_r108_c62 bl[62] br[62] wl[108] vdd gnd cell_6t
Xbit_r109_c62 bl[62] br[62] wl[109] vdd gnd cell_6t
Xbit_r110_c62 bl[62] br[62] wl[110] vdd gnd cell_6t
Xbit_r111_c62 bl[62] br[62] wl[111] vdd gnd cell_6t
Xbit_r112_c62 bl[62] br[62] wl[112] vdd gnd cell_6t
Xbit_r113_c62 bl[62] br[62] wl[113] vdd gnd cell_6t
Xbit_r114_c62 bl[62] br[62] wl[114] vdd gnd cell_6t
Xbit_r115_c62 bl[62] br[62] wl[115] vdd gnd cell_6t
Xbit_r116_c62 bl[62] br[62] wl[116] vdd gnd cell_6t
Xbit_r117_c62 bl[62] br[62] wl[117] vdd gnd cell_6t
Xbit_r118_c62 bl[62] br[62] wl[118] vdd gnd cell_6t
Xbit_r119_c62 bl[62] br[62] wl[119] vdd gnd cell_6t
Xbit_r120_c62 bl[62] br[62] wl[120] vdd gnd cell_6t
Xbit_r121_c62 bl[62] br[62] wl[121] vdd gnd cell_6t
Xbit_r122_c62 bl[62] br[62] wl[122] vdd gnd cell_6t
Xbit_r123_c62 bl[62] br[62] wl[123] vdd gnd cell_6t
Xbit_r124_c62 bl[62] br[62] wl[124] vdd gnd cell_6t
Xbit_r125_c62 bl[62] br[62] wl[125] vdd gnd cell_6t
Xbit_r126_c62 bl[62] br[62] wl[126] vdd gnd cell_6t
Xbit_r127_c62 bl[62] br[62] wl[127] vdd gnd cell_6t
Xbit_r128_c62 bl[62] br[62] wl[128] vdd gnd cell_6t
Xbit_r129_c62 bl[62] br[62] wl[129] vdd gnd cell_6t
Xbit_r130_c62 bl[62] br[62] wl[130] vdd gnd cell_6t
Xbit_r131_c62 bl[62] br[62] wl[131] vdd gnd cell_6t
Xbit_r132_c62 bl[62] br[62] wl[132] vdd gnd cell_6t
Xbit_r133_c62 bl[62] br[62] wl[133] vdd gnd cell_6t
Xbit_r134_c62 bl[62] br[62] wl[134] vdd gnd cell_6t
Xbit_r135_c62 bl[62] br[62] wl[135] vdd gnd cell_6t
Xbit_r136_c62 bl[62] br[62] wl[136] vdd gnd cell_6t
Xbit_r137_c62 bl[62] br[62] wl[137] vdd gnd cell_6t
Xbit_r138_c62 bl[62] br[62] wl[138] vdd gnd cell_6t
Xbit_r139_c62 bl[62] br[62] wl[139] vdd gnd cell_6t
Xbit_r140_c62 bl[62] br[62] wl[140] vdd gnd cell_6t
Xbit_r141_c62 bl[62] br[62] wl[141] vdd gnd cell_6t
Xbit_r142_c62 bl[62] br[62] wl[142] vdd gnd cell_6t
Xbit_r143_c62 bl[62] br[62] wl[143] vdd gnd cell_6t
Xbit_r144_c62 bl[62] br[62] wl[144] vdd gnd cell_6t
Xbit_r145_c62 bl[62] br[62] wl[145] vdd gnd cell_6t
Xbit_r146_c62 bl[62] br[62] wl[146] vdd gnd cell_6t
Xbit_r147_c62 bl[62] br[62] wl[147] vdd gnd cell_6t
Xbit_r148_c62 bl[62] br[62] wl[148] vdd gnd cell_6t
Xbit_r149_c62 bl[62] br[62] wl[149] vdd gnd cell_6t
Xbit_r150_c62 bl[62] br[62] wl[150] vdd gnd cell_6t
Xbit_r151_c62 bl[62] br[62] wl[151] vdd gnd cell_6t
Xbit_r152_c62 bl[62] br[62] wl[152] vdd gnd cell_6t
Xbit_r153_c62 bl[62] br[62] wl[153] vdd gnd cell_6t
Xbit_r154_c62 bl[62] br[62] wl[154] vdd gnd cell_6t
Xbit_r155_c62 bl[62] br[62] wl[155] vdd gnd cell_6t
Xbit_r156_c62 bl[62] br[62] wl[156] vdd gnd cell_6t
Xbit_r157_c62 bl[62] br[62] wl[157] vdd gnd cell_6t
Xbit_r158_c62 bl[62] br[62] wl[158] vdd gnd cell_6t
Xbit_r159_c62 bl[62] br[62] wl[159] vdd gnd cell_6t
Xbit_r160_c62 bl[62] br[62] wl[160] vdd gnd cell_6t
Xbit_r161_c62 bl[62] br[62] wl[161] vdd gnd cell_6t
Xbit_r162_c62 bl[62] br[62] wl[162] vdd gnd cell_6t
Xbit_r163_c62 bl[62] br[62] wl[163] vdd gnd cell_6t
Xbit_r164_c62 bl[62] br[62] wl[164] vdd gnd cell_6t
Xbit_r165_c62 bl[62] br[62] wl[165] vdd gnd cell_6t
Xbit_r166_c62 bl[62] br[62] wl[166] vdd gnd cell_6t
Xbit_r167_c62 bl[62] br[62] wl[167] vdd gnd cell_6t
Xbit_r168_c62 bl[62] br[62] wl[168] vdd gnd cell_6t
Xbit_r169_c62 bl[62] br[62] wl[169] vdd gnd cell_6t
Xbit_r170_c62 bl[62] br[62] wl[170] vdd gnd cell_6t
Xbit_r171_c62 bl[62] br[62] wl[171] vdd gnd cell_6t
Xbit_r172_c62 bl[62] br[62] wl[172] vdd gnd cell_6t
Xbit_r173_c62 bl[62] br[62] wl[173] vdd gnd cell_6t
Xbit_r174_c62 bl[62] br[62] wl[174] vdd gnd cell_6t
Xbit_r175_c62 bl[62] br[62] wl[175] vdd gnd cell_6t
Xbit_r176_c62 bl[62] br[62] wl[176] vdd gnd cell_6t
Xbit_r177_c62 bl[62] br[62] wl[177] vdd gnd cell_6t
Xbit_r178_c62 bl[62] br[62] wl[178] vdd gnd cell_6t
Xbit_r179_c62 bl[62] br[62] wl[179] vdd gnd cell_6t
Xbit_r180_c62 bl[62] br[62] wl[180] vdd gnd cell_6t
Xbit_r181_c62 bl[62] br[62] wl[181] vdd gnd cell_6t
Xbit_r182_c62 bl[62] br[62] wl[182] vdd gnd cell_6t
Xbit_r183_c62 bl[62] br[62] wl[183] vdd gnd cell_6t
Xbit_r184_c62 bl[62] br[62] wl[184] vdd gnd cell_6t
Xbit_r185_c62 bl[62] br[62] wl[185] vdd gnd cell_6t
Xbit_r186_c62 bl[62] br[62] wl[186] vdd gnd cell_6t
Xbit_r187_c62 bl[62] br[62] wl[187] vdd gnd cell_6t
Xbit_r188_c62 bl[62] br[62] wl[188] vdd gnd cell_6t
Xbit_r189_c62 bl[62] br[62] wl[189] vdd gnd cell_6t
Xbit_r190_c62 bl[62] br[62] wl[190] vdd gnd cell_6t
Xbit_r191_c62 bl[62] br[62] wl[191] vdd gnd cell_6t
Xbit_r192_c62 bl[62] br[62] wl[192] vdd gnd cell_6t
Xbit_r193_c62 bl[62] br[62] wl[193] vdd gnd cell_6t
Xbit_r194_c62 bl[62] br[62] wl[194] vdd gnd cell_6t
Xbit_r195_c62 bl[62] br[62] wl[195] vdd gnd cell_6t
Xbit_r196_c62 bl[62] br[62] wl[196] vdd gnd cell_6t
Xbit_r197_c62 bl[62] br[62] wl[197] vdd gnd cell_6t
Xbit_r198_c62 bl[62] br[62] wl[198] vdd gnd cell_6t
Xbit_r199_c62 bl[62] br[62] wl[199] vdd gnd cell_6t
Xbit_r200_c62 bl[62] br[62] wl[200] vdd gnd cell_6t
Xbit_r201_c62 bl[62] br[62] wl[201] vdd gnd cell_6t
Xbit_r202_c62 bl[62] br[62] wl[202] vdd gnd cell_6t
Xbit_r203_c62 bl[62] br[62] wl[203] vdd gnd cell_6t
Xbit_r204_c62 bl[62] br[62] wl[204] vdd gnd cell_6t
Xbit_r205_c62 bl[62] br[62] wl[205] vdd gnd cell_6t
Xbit_r206_c62 bl[62] br[62] wl[206] vdd gnd cell_6t
Xbit_r207_c62 bl[62] br[62] wl[207] vdd gnd cell_6t
Xbit_r208_c62 bl[62] br[62] wl[208] vdd gnd cell_6t
Xbit_r209_c62 bl[62] br[62] wl[209] vdd gnd cell_6t
Xbit_r210_c62 bl[62] br[62] wl[210] vdd gnd cell_6t
Xbit_r211_c62 bl[62] br[62] wl[211] vdd gnd cell_6t
Xbit_r212_c62 bl[62] br[62] wl[212] vdd gnd cell_6t
Xbit_r213_c62 bl[62] br[62] wl[213] vdd gnd cell_6t
Xbit_r214_c62 bl[62] br[62] wl[214] vdd gnd cell_6t
Xbit_r215_c62 bl[62] br[62] wl[215] vdd gnd cell_6t
Xbit_r216_c62 bl[62] br[62] wl[216] vdd gnd cell_6t
Xbit_r217_c62 bl[62] br[62] wl[217] vdd gnd cell_6t
Xbit_r218_c62 bl[62] br[62] wl[218] vdd gnd cell_6t
Xbit_r219_c62 bl[62] br[62] wl[219] vdd gnd cell_6t
Xbit_r220_c62 bl[62] br[62] wl[220] vdd gnd cell_6t
Xbit_r221_c62 bl[62] br[62] wl[221] vdd gnd cell_6t
Xbit_r222_c62 bl[62] br[62] wl[222] vdd gnd cell_6t
Xbit_r223_c62 bl[62] br[62] wl[223] vdd gnd cell_6t
Xbit_r224_c62 bl[62] br[62] wl[224] vdd gnd cell_6t
Xbit_r225_c62 bl[62] br[62] wl[225] vdd gnd cell_6t
Xbit_r226_c62 bl[62] br[62] wl[226] vdd gnd cell_6t
Xbit_r227_c62 bl[62] br[62] wl[227] vdd gnd cell_6t
Xbit_r228_c62 bl[62] br[62] wl[228] vdd gnd cell_6t
Xbit_r229_c62 bl[62] br[62] wl[229] vdd gnd cell_6t
Xbit_r230_c62 bl[62] br[62] wl[230] vdd gnd cell_6t
Xbit_r231_c62 bl[62] br[62] wl[231] vdd gnd cell_6t
Xbit_r232_c62 bl[62] br[62] wl[232] vdd gnd cell_6t
Xbit_r233_c62 bl[62] br[62] wl[233] vdd gnd cell_6t
Xbit_r234_c62 bl[62] br[62] wl[234] vdd gnd cell_6t
Xbit_r235_c62 bl[62] br[62] wl[235] vdd gnd cell_6t
Xbit_r236_c62 bl[62] br[62] wl[236] vdd gnd cell_6t
Xbit_r237_c62 bl[62] br[62] wl[237] vdd gnd cell_6t
Xbit_r238_c62 bl[62] br[62] wl[238] vdd gnd cell_6t
Xbit_r239_c62 bl[62] br[62] wl[239] vdd gnd cell_6t
Xbit_r240_c62 bl[62] br[62] wl[240] vdd gnd cell_6t
Xbit_r241_c62 bl[62] br[62] wl[241] vdd gnd cell_6t
Xbit_r242_c62 bl[62] br[62] wl[242] vdd gnd cell_6t
Xbit_r243_c62 bl[62] br[62] wl[243] vdd gnd cell_6t
Xbit_r244_c62 bl[62] br[62] wl[244] vdd gnd cell_6t
Xbit_r245_c62 bl[62] br[62] wl[245] vdd gnd cell_6t
Xbit_r246_c62 bl[62] br[62] wl[246] vdd gnd cell_6t
Xbit_r247_c62 bl[62] br[62] wl[247] vdd gnd cell_6t
Xbit_r248_c62 bl[62] br[62] wl[248] vdd gnd cell_6t
Xbit_r249_c62 bl[62] br[62] wl[249] vdd gnd cell_6t
Xbit_r250_c62 bl[62] br[62] wl[250] vdd gnd cell_6t
Xbit_r251_c62 bl[62] br[62] wl[251] vdd gnd cell_6t
Xbit_r252_c62 bl[62] br[62] wl[252] vdd gnd cell_6t
Xbit_r253_c62 bl[62] br[62] wl[253] vdd gnd cell_6t
Xbit_r254_c62 bl[62] br[62] wl[254] vdd gnd cell_6t
Xbit_r255_c62 bl[62] br[62] wl[255] vdd gnd cell_6t
Xbit_r256_c62 bl[62] br[62] wl[256] vdd gnd cell_6t
Xbit_r257_c62 bl[62] br[62] wl[257] vdd gnd cell_6t
Xbit_r258_c62 bl[62] br[62] wl[258] vdd gnd cell_6t
Xbit_r259_c62 bl[62] br[62] wl[259] vdd gnd cell_6t
Xbit_r260_c62 bl[62] br[62] wl[260] vdd gnd cell_6t
Xbit_r261_c62 bl[62] br[62] wl[261] vdd gnd cell_6t
Xbit_r262_c62 bl[62] br[62] wl[262] vdd gnd cell_6t
Xbit_r263_c62 bl[62] br[62] wl[263] vdd gnd cell_6t
Xbit_r264_c62 bl[62] br[62] wl[264] vdd gnd cell_6t
Xbit_r265_c62 bl[62] br[62] wl[265] vdd gnd cell_6t
Xbit_r266_c62 bl[62] br[62] wl[266] vdd gnd cell_6t
Xbit_r267_c62 bl[62] br[62] wl[267] vdd gnd cell_6t
Xbit_r268_c62 bl[62] br[62] wl[268] vdd gnd cell_6t
Xbit_r269_c62 bl[62] br[62] wl[269] vdd gnd cell_6t
Xbit_r270_c62 bl[62] br[62] wl[270] vdd gnd cell_6t
Xbit_r271_c62 bl[62] br[62] wl[271] vdd gnd cell_6t
Xbit_r272_c62 bl[62] br[62] wl[272] vdd gnd cell_6t
Xbit_r273_c62 bl[62] br[62] wl[273] vdd gnd cell_6t
Xbit_r274_c62 bl[62] br[62] wl[274] vdd gnd cell_6t
Xbit_r275_c62 bl[62] br[62] wl[275] vdd gnd cell_6t
Xbit_r276_c62 bl[62] br[62] wl[276] vdd gnd cell_6t
Xbit_r277_c62 bl[62] br[62] wl[277] vdd gnd cell_6t
Xbit_r278_c62 bl[62] br[62] wl[278] vdd gnd cell_6t
Xbit_r279_c62 bl[62] br[62] wl[279] vdd gnd cell_6t
Xbit_r280_c62 bl[62] br[62] wl[280] vdd gnd cell_6t
Xbit_r281_c62 bl[62] br[62] wl[281] vdd gnd cell_6t
Xbit_r282_c62 bl[62] br[62] wl[282] vdd gnd cell_6t
Xbit_r283_c62 bl[62] br[62] wl[283] vdd gnd cell_6t
Xbit_r284_c62 bl[62] br[62] wl[284] vdd gnd cell_6t
Xbit_r285_c62 bl[62] br[62] wl[285] vdd gnd cell_6t
Xbit_r286_c62 bl[62] br[62] wl[286] vdd gnd cell_6t
Xbit_r287_c62 bl[62] br[62] wl[287] vdd gnd cell_6t
Xbit_r288_c62 bl[62] br[62] wl[288] vdd gnd cell_6t
Xbit_r289_c62 bl[62] br[62] wl[289] vdd gnd cell_6t
Xbit_r290_c62 bl[62] br[62] wl[290] vdd gnd cell_6t
Xbit_r291_c62 bl[62] br[62] wl[291] vdd gnd cell_6t
Xbit_r292_c62 bl[62] br[62] wl[292] vdd gnd cell_6t
Xbit_r293_c62 bl[62] br[62] wl[293] vdd gnd cell_6t
Xbit_r294_c62 bl[62] br[62] wl[294] vdd gnd cell_6t
Xbit_r295_c62 bl[62] br[62] wl[295] vdd gnd cell_6t
Xbit_r296_c62 bl[62] br[62] wl[296] vdd gnd cell_6t
Xbit_r297_c62 bl[62] br[62] wl[297] vdd gnd cell_6t
Xbit_r298_c62 bl[62] br[62] wl[298] vdd gnd cell_6t
Xbit_r299_c62 bl[62] br[62] wl[299] vdd gnd cell_6t
Xbit_r300_c62 bl[62] br[62] wl[300] vdd gnd cell_6t
Xbit_r301_c62 bl[62] br[62] wl[301] vdd gnd cell_6t
Xbit_r302_c62 bl[62] br[62] wl[302] vdd gnd cell_6t
Xbit_r303_c62 bl[62] br[62] wl[303] vdd gnd cell_6t
Xbit_r304_c62 bl[62] br[62] wl[304] vdd gnd cell_6t
Xbit_r305_c62 bl[62] br[62] wl[305] vdd gnd cell_6t
Xbit_r306_c62 bl[62] br[62] wl[306] vdd gnd cell_6t
Xbit_r307_c62 bl[62] br[62] wl[307] vdd gnd cell_6t
Xbit_r308_c62 bl[62] br[62] wl[308] vdd gnd cell_6t
Xbit_r309_c62 bl[62] br[62] wl[309] vdd gnd cell_6t
Xbit_r310_c62 bl[62] br[62] wl[310] vdd gnd cell_6t
Xbit_r311_c62 bl[62] br[62] wl[311] vdd gnd cell_6t
Xbit_r312_c62 bl[62] br[62] wl[312] vdd gnd cell_6t
Xbit_r313_c62 bl[62] br[62] wl[313] vdd gnd cell_6t
Xbit_r314_c62 bl[62] br[62] wl[314] vdd gnd cell_6t
Xbit_r315_c62 bl[62] br[62] wl[315] vdd gnd cell_6t
Xbit_r316_c62 bl[62] br[62] wl[316] vdd gnd cell_6t
Xbit_r317_c62 bl[62] br[62] wl[317] vdd gnd cell_6t
Xbit_r318_c62 bl[62] br[62] wl[318] vdd gnd cell_6t
Xbit_r319_c62 bl[62] br[62] wl[319] vdd gnd cell_6t
Xbit_r320_c62 bl[62] br[62] wl[320] vdd gnd cell_6t
Xbit_r321_c62 bl[62] br[62] wl[321] vdd gnd cell_6t
Xbit_r322_c62 bl[62] br[62] wl[322] vdd gnd cell_6t
Xbit_r323_c62 bl[62] br[62] wl[323] vdd gnd cell_6t
Xbit_r324_c62 bl[62] br[62] wl[324] vdd gnd cell_6t
Xbit_r325_c62 bl[62] br[62] wl[325] vdd gnd cell_6t
Xbit_r326_c62 bl[62] br[62] wl[326] vdd gnd cell_6t
Xbit_r327_c62 bl[62] br[62] wl[327] vdd gnd cell_6t
Xbit_r328_c62 bl[62] br[62] wl[328] vdd gnd cell_6t
Xbit_r329_c62 bl[62] br[62] wl[329] vdd gnd cell_6t
Xbit_r330_c62 bl[62] br[62] wl[330] vdd gnd cell_6t
Xbit_r331_c62 bl[62] br[62] wl[331] vdd gnd cell_6t
Xbit_r332_c62 bl[62] br[62] wl[332] vdd gnd cell_6t
Xbit_r333_c62 bl[62] br[62] wl[333] vdd gnd cell_6t
Xbit_r334_c62 bl[62] br[62] wl[334] vdd gnd cell_6t
Xbit_r335_c62 bl[62] br[62] wl[335] vdd gnd cell_6t
Xbit_r336_c62 bl[62] br[62] wl[336] vdd gnd cell_6t
Xbit_r337_c62 bl[62] br[62] wl[337] vdd gnd cell_6t
Xbit_r338_c62 bl[62] br[62] wl[338] vdd gnd cell_6t
Xbit_r339_c62 bl[62] br[62] wl[339] vdd gnd cell_6t
Xbit_r340_c62 bl[62] br[62] wl[340] vdd gnd cell_6t
Xbit_r341_c62 bl[62] br[62] wl[341] vdd gnd cell_6t
Xbit_r342_c62 bl[62] br[62] wl[342] vdd gnd cell_6t
Xbit_r343_c62 bl[62] br[62] wl[343] vdd gnd cell_6t
Xbit_r344_c62 bl[62] br[62] wl[344] vdd gnd cell_6t
Xbit_r345_c62 bl[62] br[62] wl[345] vdd gnd cell_6t
Xbit_r346_c62 bl[62] br[62] wl[346] vdd gnd cell_6t
Xbit_r347_c62 bl[62] br[62] wl[347] vdd gnd cell_6t
Xbit_r348_c62 bl[62] br[62] wl[348] vdd gnd cell_6t
Xbit_r349_c62 bl[62] br[62] wl[349] vdd gnd cell_6t
Xbit_r350_c62 bl[62] br[62] wl[350] vdd gnd cell_6t
Xbit_r351_c62 bl[62] br[62] wl[351] vdd gnd cell_6t
Xbit_r352_c62 bl[62] br[62] wl[352] vdd gnd cell_6t
Xbit_r353_c62 bl[62] br[62] wl[353] vdd gnd cell_6t
Xbit_r354_c62 bl[62] br[62] wl[354] vdd gnd cell_6t
Xbit_r355_c62 bl[62] br[62] wl[355] vdd gnd cell_6t
Xbit_r356_c62 bl[62] br[62] wl[356] vdd gnd cell_6t
Xbit_r357_c62 bl[62] br[62] wl[357] vdd gnd cell_6t
Xbit_r358_c62 bl[62] br[62] wl[358] vdd gnd cell_6t
Xbit_r359_c62 bl[62] br[62] wl[359] vdd gnd cell_6t
Xbit_r360_c62 bl[62] br[62] wl[360] vdd gnd cell_6t
Xbit_r361_c62 bl[62] br[62] wl[361] vdd gnd cell_6t
Xbit_r362_c62 bl[62] br[62] wl[362] vdd gnd cell_6t
Xbit_r363_c62 bl[62] br[62] wl[363] vdd gnd cell_6t
Xbit_r364_c62 bl[62] br[62] wl[364] vdd gnd cell_6t
Xbit_r365_c62 bl[62] br[62] wl[365] vdd gnd cell_6t
Xbit_r366_c62 bl[62] br[62] wl[366] vdd gnd cell_6t
Xbit_r367_c62 bl[62] br[62] wl[367] vdd gnd cell_6t
Xbit_r368_c62 bl[62] br[62] wl[368] vdd gnd cell_6t
Xbit_r369_c62 bl[62] br[62] wl[369] vdd gnd cell_6t
Xbit_r370_c62 bl[62] br[62] wl[370] vdd gnd cell_6t
Xbit_r371_c62 bl[62] br[62] wl[371] vdd gnd cell_6t
Xbit_r372_c62 bl[62] br[62] wl[372] vdd gnd cell_6t
Xbit_r373_c62 bl[62] br[62] wl[373] vdd gnd cell_6t
Xbit_r374_c62 bl[62] br[62] wl[374] vdd gnd cell_6t
Xbit_r375_c62 bl[62] br[62] wl[375] vdd gnd cell_6t
Xbit_r376_c62 bl[62] br[62] wl[376] vdd gnd cell_6t
Xbit_r377_c62 bl[62] br[62] wl[377] vdd gnd cell_6t
Xbit_r378_c62 bl[62] br[62] wl[378] vdd gnd cell_6t
Xbit_r379_c62 bl[62] br[62] wl[379] vdd gnd cell_6t
Xbit_r380_c62 bl[62] br[62] wl[380] vdd gnd cell_6t
Xbit_r381_c62 bl[62] br[62] wl[381] vdd gnd cell_6t
Xbit_r382_c62 bl[62] br[62] wl[382] vdd gnd cell_6t
Xbit_r383_c62 bl[62] br[62] wl[383] vdd gnd cell_6t
Xbit_r384_c62 bl[62] br[62] wl[384] vdd gnd cell_6t
Xbit_r385_c62 bl[62] br[62] wl[385] vdd gnd cell_6t
Xbit_r386_c62 bl[62] br[62] wl[386] vdd gnd cell_6t
Xbit_r387_c62 bl[62] br[62] wl[387] vdd gnd cell_6t
Xbit_r388_c62 bl[62] br[62] wl[388] vdd gnd cell_6t
Xbit_r389_c62 bl[62] br[62] wl[389] vdd gnd cell_6t
Xbit_r390_c62 bl[62] br[62] wl[390] vdd gnd cell_6t
Xbit_r391_c62 bl[62] br[62] wl[391] vdd gnd cell_6t
Xbit_r392_c62 bl[62] br[62] wl[392] vdd gnd cell_6t
Xbit_r393_c62 bl[62] br[62] wl[393] vdd gnd cell_6t
Xbit_r394_c62 bl[62] br[62] wl[394] vdd gnd cell_6t
Xbit_r395_c62 bl[62] br[62] wl[395] vdd gnd cell_6t
Xbit_r396_c62 bl[62] br[62] wl[396] vdd gnd cell_6t
Xbit_r397_c62 bl[62] br[62] wl[397] vdd gnd cell_6t
Xbit_r398_c62 bl[62] br[62] wl[398] vdd gnd cell_6t
Xbit_r399_c62 bl[62] br[62] wl[399] vdd gnd cell_6t
Xbit_r400_c62 bl[62] br[62] wl[400] vdd gnd cell_6t
Xbit_r401_c62 bl[62] br[62] wl[401] vdd gnd cell_6t
Xbit_r402_c62 bl[62] br[62] wl[402] vdd gnd cell_6t
Xbit_r403_c62 bl[62] br[62] wl[403] vdd gnd cell_6t
Xbit_r404_c62 bl[62] br[62] wl[404] vdd gnd cell_6t
Xbit_r405_c62 bl[62] br[62] wl[405] vdd gnd cell_6t
Xbit_r406_c62 bl[62] br[62] wl[406] vdd gnd cell_6t
Xbit_r407_c62 bl[62] br[62] wl[407] vdd gnd cell_6t
Xbit_r408_c62 bl[62] br[62] wl[408] vdd gnd cell_6t
Xbit_r409_c62 bl[62] br[62] wl[409] vdd gnd cell_6t
Xbit_r410_c62 bl[62] br[62] wl[410] vdd gnd cell_6t
Xbit_r411_c62 bl[62] br[62] wl[411] vdd gnd cell_6t
Xbit_r412_c62 bl[62] br[62] wl[412] vdd gnd cell_6t
Xbit_r413_c62 bl[62] br[62] wl[413] vdd gnd cell_6t
Xbit_r414_c62 bl[62] br[62] wl[414] vdd gnd cell_6t
Xbit_r415_c62 bl[62] br[62] wl[415] vdd gnd cell_6t
Xbit_r416_c62 bl[62] br[62] wl[416] vdd gnd cell_6t
Xbit_r417_c62 bl[62] br[62] wl[417] vdd gnd cell_6t
Xbit_r418_c62 bl[62] br[62] wl[418] vdd gnd cell_6t
Xbit_r419_c62 bl[62] br[62] wl[419] vdd gnd cell_6t
Xbit_r420_c62 bl[62] br[62] wl[420] vdd gnd cell_6t
Xbit_r421_c62 bl[62] br[62] wl[421] vdd gnd cell_6t
Xbit_r422_c62 bl[62] br[62] wl[422] vdd gnd cell_6t
Xbit_r423_c62 bl[62] br[62] wl[423] vdd gnd cell_6t
Xbit_r424_c62 bl[62] br[62] wl[424] vdd gnd cell_6t
Xbit_r425_c62 bl[62] br[62] wl[425] vdd gnd cell_6t
Xbit_r426_c62 bl[62] br[62] wl[426] vdd gnd cell_6t
Xbit_r427_c62 bl[62] br[62] wl[427] vdd gnd cell_6t
Xbit_r428_c62 bl[62] br[62] wl[428] vdd gnd cell_6t
Xbit_r429_c62 bl[62] br[62] wl[429] vdd gnd cell_6t
Xbit_r430_c62 bl[62] br[62] wl[430] vdd gnd cell_6t
Xbit_r431_c62 bl[62] br[62] wl[431] vdd gnd cell_6t
Xbit_r432_c62 bl[62] br[62] wl[432] vdd gnd cell_6t
Xbit_r433_c62 bl[62] br[62] wl[433] vdd gnd cell_6t
Xbit_r434_c62 bl[62] br[62] wl[434] vdd gnd cell_6t
Xbit_r435_c62 bl[62] br[62] wl[435] vdd gnd cell_6t
Xbit_r436_c62 bl[62] br[62] wl[436] vdd gnd cell_6t
Xbit_r437_c62 bl[62] br[62] wl[437] vdd gnd cell_6t
Xbit_r438_c62 bl[62] br[62] wl[438] vdd gnd cell_6t
Xbit_r439_c62 bl[62] br[62] wl[439] vdd gnd cell_6t
Xbit_r440_c62 bl[62] br[62] wl[440] vdd gnd cell_6t
Xbit_r441_c62 bl[62] br[62] wl[441] vdd gnd cell_6t
Xbit_r442_c62 bl[62] br[62] wl[442] vdd gnd cell_6t
Xbit_r443_c62 bl[62] br[62] wl[443] vdd gnd cell_6t
Xbit_r444_c62 bl[62] br[62] wl[444] vdd gnd cell_6t
Xbit_r445_c62 bl[62] br[62] wl[445] vdd gnd cell_6t
Xbit_r446_c62 bl[62] br[62] wl[446] vdd gnd cell_6t
Xbit_r447_c62 bl[62] br[62] wl[447] vdd gnd cell_6t
Xbit_r448_c62 bl[62] br[62] wl[448] vdd gnd cell_6t
Xbit_r449_c62 bl[62] br[62] wl[449] vdd gnd cell_6t
Xbit_r450_c62 bl[62] br[62] wl[450] vdd gnd cell_6t
Xbit_r451_c62 bl[62] br[62] wl[451] vdd gnd cell_6t
Xbit_r452_c62 bl[62] br[62] wl[452] vdd gnd cell_6t
Xbit_r453_c62 bl[62] br[62] wl[453] vdd gnd cell_6t
Xbit_r454_c62 bl[62] br[62] wl[454] vdd gnd cell_6t
Xbit_r455_c62 bl[62] br[62] wl[455] vdd gnd cell_6t
Xbit_r456_c62 bl[62] br[62] wl[456] vdd gnd cell_6t
Xbit_r457_c62 bl[62] br[62] wl[457] vdd gnd cell_6t
Xbit_r458_c62 bl[62] br[62] wl[458] vdd gnd cell_6t
Xbit_r459_c62 bl[62] br[62] wl[459] vdd gnd cell_6t
Xbit_r460_c62 bl[62] br[62] wl[460] vdd gnd cell_6t
Xbit_r461_c62 bl[62] br[62] wl[461] vdd gnd cell_6t
Xbit_r462_c62 bl[62] br[62] wl[462] vdd gnd cell_6t
Xbit_r463_c62 bl[62] br[62] wl[463] vdd gnd cell_6t
Xbit_r464_c62 bl[62] br[62] wl[464] vdd gnd cell_6t
Xbit_r465_c62 bl[62] br[62] wl[465] vdd gnd cell_6t
Xbit_r466_c62 bl[62] br[62] wl[466] vdd gnd cell_6t
Xbit_r467_c62 bl[62] br[62] wl[467] vdd gnd cell_6t
Xbit_r468_c62 bl[62] br[62] wl[468] vdd gnd cell_6t
Xbit_r469_c62 bl[62] br[62] wl[469] vdd gnd cell_6t
Xbit_r470_c62 bl[62] br[62] wl[470] vdd gnd cell_6t
Xbit_r471_c62 bl[62] br[62] wl[471] vdd gnd cell_6t
Xbit_r472_c62 bl[62] br[62] wl[472] vdd gnd cell_6t
Xbit_r473_c62 bl[62] br[62] wl[473] vdd gnd cell_6t
Xbit_r474_c62 bl[62] br[62] wl[474] vdd gnd cell_6t
Xbit_r475_c62 bl[62] br[62] wl[475] vdd gnd cell_6t
Xbit_r476_c62 bl[62] br[62] wl[476] vdd gnd cell_6t
Xbit_r477_c62 bl[62] br[62] wl[477] vdd gnd cell_6t
Xbit_r478_c62 bl[62] br[62] wl[478] vdd gnd cell_6t
Xbit_r479_c62 bl[62] br[62] wl[479] vdd gnd cell_6t
Xbit_r480_c62 bl[62] br[62] wl[480] vdd gnd cell_6t
Xbit_r481_c62 bl[62] br[62] wl[481] vdd gnd cell_6t
Xbit_r482_c62 bl[62] br[62] wl[482] vdd gnd cell_6t
Xbit_r483_c62 bl[62] br[62] wl[483] vdd gnd cell_6t
Xbit_r484_c62 bl[62] br[62] wl[484] vdd gnd cell_6t
Xbit_r485_c62 bl[62] br[62] wl[485] vdd gnd cell_6t
Xbit_r486_c62 bl[62] br[62] wl[486] vdd gnd cell_6t
Xbit_r487_c62 bl[62] br[62] wl[487] vdd gnd cell_6t
Xbit_r488_c62 bl[62] br[62] wl[488] vdd gnd cell_6t
Xbit_r489_c62 bl[62] br[62] wl[489] vdd gnd cell_6t
Xbit_r490_c62 bl[62] br[62] wl[490] vdd gnd cell_6t
Xbit_r491_c62 bl[62] br[62] wl[491] vdd gnd cell_6t
Xbit_r492_c62 bl[62] br[62] wl[492] vdd gnd cell_6t
Xbit_r493_c62 bl[62] br[62] wl[493] vdd gnd cell_6t
Xbit_r494_c62 bl[62] br[62] wl[494] vdd gnd cell_6t
Xbit_r495_c62 bl[62] br[62] wl[495] vdd gnd cell_6t
Xbit_r496_c62 bl[62] br[62] wl[496] vdd gnd cell_6t
Xbit_r497_c62 bl[62] br[62] wl[497] vdd gnd cell_6t
Xbit_r498_c62 bl[62] br[62] wl[498] vdd gnd cell_6t
Xbit_r499_c62 bl[62] br[62] wl[499] vdd gnd cell_6t
Xbit_r500_c62 bl[62] br[62] wl[500] vdd gnd cell_6t
Xbit_r501_c62 bl[62] br[62] wl[501] vdd gnd cell_6t
Xbit_r502_c62 bl[62] br[62] wl[502] vdd gnd cell_6t
Xbit_r503_c62 bl[62] br[62] wl[503] vdd gnd cell_6t
Xbit_r504_c62 bl[62] br[62] wl[504] vdd gnd cell_6t
Xbit_r505_c62 bl[62] br[62] wl[505] vdd gnd cell_6t
Xbit_r506_c62 bl[62] br[62] wl[506] vdd gnd cell_6t
Xbit_r507_c62 bl[62] br[62] wl[507] vdd gnd cell_6t
Xbit_r508_c62 bl[62] br[62] wl[508] vdd gnd cell_6t
Xbit_r509_c62 bl[62] br[62] wl[509] vdd gnd cell_6t
Xbit_r510_c62 bl[62] br[62] wl[510] vdd gnd cell_6t
Xbit_r511_c62 bl[62] br[62] wl[511] vdd gnd cell_6t
Xbit_r0_c63 bl[63] br[63] wl[0] vdd gnd cell_6t
Xbit_r1_c63 bl[63] br[63] wl[1] vdd gnd cell_6t
Xbit_r2_c63 bl[63] br[63] wl[2] vdd gnd cell_6t
Xbit_r3_c63 bl[63] br[63] wl[3] vdd gnd cell_6t
Xbit_r4_c63 bl[63] br[63] wl[4] vdd gnd cell_6t
Xbit_r5_c63 bl[63] br[63] wl[5] vdd gnd cell_6t
Xbit_r6_c63 bl[63] br[63] wl[6] vdd gnd cell_6t
Xbit_r7_c63 bl[63] br[63] wl[7] vdd gnd cell_6t
Xbit_r8_c63 bl[63] br[63] wl[8] vdd gnd cell_6t
Xbit_r9_c63 bl[63] br[63] wl[9] vdd gnd cell_6t
Xbit_r10_c63 bl[63] br[63] wl[10] vdd gnd cell_6t
Xbit_r11_c63 bl[63] br[63] wl[11] vdd gnd cell_6t
Xbit_r12_c63 bl[63] br[63] wl[12] vdd gnd cell_6t
Xbit_r13_c63 bl[63] br[63] wl[13] vdd gnd cell_6t
Xbit_r14_c63 bl[63] br[63] wl[14] vdd gnd cell_6t
Xbit_r15_c63 bl[63] br[63] wl[15] vdd gnd cell_6t
Xbit_r16_c63 bl[63] br[63] wl[16] vdd gnd cell_6t
Xbit_r17_c63 bl[63] br[63] wl[17] vdd gnd cell_6t
Xbit_r18_c63 bl[63] br[63] wl[18] vdd gnd cell_6t
Xbit_r19_c63 bl[63] br[63] wl[19] vdd gnd cell_6t
Xbit_r20_c63 bl[63] br[63] wl[20] vdd gnd cell_6t
Xbit_r21_c63 bl[63] br[63] wl[21] vdd gnd cell_6t
Xbit_r22_c63 bl[63] br[63] wl[22] vdd gnd cell_6t
Xbit_r23_c63 bl[63] br[63] wl[23] vdd gnd cell_6t
Xbit_r24_c63 bl[63] br[63] wl[24] vdd gnd cell_6t
Xbit_r25_c63 bl[63] br[63] wl[25] vdd gnd cell_6t
Xbit_r26_c63 bl[63] br[63] wl[26] vdd gnd cell_6t
Xbit_r27_c63 bl[63] br[63] wl[27] vdd gnd cell_6t
Xbit_r28_c63 bl[63] br[63] wl[28] vdd gnd cell_6t
Xbit_r29_c63 bl[63] br[63] wl[29] vdd gnd cell_6t
Xbit_r30_c63 bl[63] br[63] wl[30] vdd gnd cell_6t
Xbit_r31_c63 bl[63] br[63] wl[31] vdd gnd cell_6t
Xbit_r32_c63 bl[63] br[63] wl[32] vdd gnd cell_6t
Xbit_r33_c63 bl[63] br[63] wl[33] vdd gnd cell_6t
Xbit_r34_c63 bl[63] br[63] wl[34] vdd gnd cell_6t
Xbit_r35_c63 bl[63] br[63] wl[35] vdd gnd cell_6t
Xbit_r36_c63 bl[63] br[63] wl[36] vdd gnd cell_6t
Xbit_r37_c63 bl[63] br[63] wl[37] vdd gnd cell_6t
Xbit_r38_c63 bl[63] br[63] wl[38] vdd gnd cell_6t
Xbit_r39_c63 bl[63] br[63] wl[39] vdd gnd cell_6t
Xbit_r40_c63 bl[63] br[63] wl[40] vdd gnd cell_6t
Xbit_r41_c63 bl[63] br[63] wl[41] vdd gnd cell_6t
Xbit_r42_c63 bl[63] br[63] wl[42] vdd gnd cell_6t
Xbit_r43_c63 bl[63] br[63] wl[43] vdd gnd cell_6t
Xbit_r44_c63 bl[63] br[63] wl[44] vdd gnd cell_6t
Xbit_r45_c63 bl[63] br[63] wl[45] vdd gnd cell_6t
Xbit_r46_c63 bl[63] br[63] wl[46] vdd gnd cell_6t
Xbit_r47_c63 bl[63] br[63] wl[47] vdd gnd cell_6t
Xbit_r48_c63 bl[63] br[63] wl[48] vdd gnd cell_6t
Xbit_r49_c63 bl[63] br[63] wl[49] vdd gnd cell_6t
Xbit_r50_c63 bl[63] br[63] wl[50] vdd gnd cell_6t
Xbit_r51_c63 bl[63] br[63] wl[51] vdd gnd cell_6t
Xbit_r52_c63 bl[63] br[63] wl[52] vdd gnd cell_6t
Xbit_r53_c63 bl[63] br[63] wl[53] vdd gnd cell_6t
Xbit_r54_c63 bl[63] br[63] wl[54] vdd gnd cell_6t
Xbit_r55_c63 bl[63] br[63] wl[55] vdd gnd cell_6t
Xbit_r56_c63 bl[63] br[63] wl[56] vdd gnd cell_6t
Xbit_r57_c63 bl[63] br[63] wl[57] vdd gnd cell_6t
Xbit_r58_c63 bl[63] br[63] wl[58] vdd gnd cell_6t
Xbit_r59_c63 bl[63] br[63] wl[59] vdd gnd cell_6t
Xbit_r60_c63 bl[63] br[63] wl[60] vdd gnd cell_6t
Xbit_r61_c63 bl[63] br[63] wl[61] vdd gnd cell_6t
Xbit_r62_c63 bl[63] br[63] wl[62] vdd gnd cell_6t
Xbit_r63_c63 bl[63] br[63] wl[63] vdd gnd cell_6t
Xbit_r64_c63 bl[63] br[63] wl[64] vdd gnd cell_6t
Xbit_r65_c63 bl[63] br[63] wl[65] vdd gnd cell_6t
Xbit_r66_c63 bl[63] br[63] wl[66] vdd gnd cell_6t
Xbit_r67_c63 bl[63] br[63] wl[67] vdd gnd cell_6t
Xbit_r68_c63 bl[63] br[63] wl[68] vdd gnd cell_6t
Xbit_r69_c63 bl[63] br[63] wl[69] vdd gnd cell_6t
Xbit_r70_c63 bl[63] br[63] wl[70] vdd gnd cell_6t
Xbit_r71_c63 bl[63] br[63] wl[71] vdd gnd cell_6t
Xbit_r72_c63 bl[63] br[63] wl[72] vdd gnd cell_6t
Xbit_r73_c63 bl[63] br[63] wl[73] vdd gnd cell_6t
Xbit_r74_c63 bl[63] br[63] wl[74] vdd gnd cell_6t
Xbit_r75_c63 bl[63] br[63] wl[75] vdd gnd cell_6t
Xbit_r76_c63 bl[63] br[63] wl[76] vdd gnd cell_6t
Xbit_r77_c63 bl[63] br[63] wl[77] vdd gnd cell_6t
Xbit_r78_c63 bl[63] br[63] wl[78] vdd gnd cell_6t
Xbit_r79_c63 bl[63] br[63] wl[79] vdd gnd cell_6t
Xbit_r80_c63 bl[63] br[63] wl[80] vdd gnd cell_6t
Xbit_r81_c63 bl[63] br[63] wl[81] vdd gnd cell_6t
Xbit_r82_c63 bl[63] br[63] wl[82] vdd gnd cell_6t
Xbit_r83_c63 bl[63] br[63] wl[83] vdd gnd cell_6t
Xbit_r84_c63 bl[63] br[63] wl[84] vdd gnd cell_6t
Xbit_r85_c63 bl[63] br[63] wl[85] vdd gnd cell_6t
Xbit_r86_c63 bl[63] br[63] wl[86] vdd gnd cell_6t
Xbit_r87_c63 bl[63] br[63] wl[87] vdd gnd cell_6t
Xbit_r88_c63 bl[63] br[63] wl[88] vdd gnd cell_6t
Xbit_r89_c63 bl[63] br[63] wl[89] vdd gnd cell_6t
Xbit_r90_c63 bl[63] br[63] wl[90] vdd gnd cell_6t
Xbit_r91_c63 bl[63] br[63] wl[91] vdd gnd cell_6t
Xbit_r92_c63 bl[63] br[63] wl[92] vdd gnd cell_6t
Xbit_r93_c63 bl[63] br[63] wl[93] vdd gnd cell_6t
Xbit_r94_c63 bl[63] br[63] wl[94] vdd gnd cell_6t
Xbit_r95_c63 bl[63] br[63] wl[95] vdd gnd cell_6t
Xbit_r96_c63 bl[63] br[63] wl[96] vdd gnd cell_6t
Xbit_r97_c63 bl[63] br[63] wl[97] vdd gnd cell_6t
Xbit_r98_c63 bl[63] br[63] wl[98] vdd gnd cell_6t
Xbit_r99_c63 bl[63] br[63] wl[99] vdd gnd cell_6t
Xbit_r100_c63 bl[63] br[63] wl[100] vdd gnd cell_6t
Xbit_r101_c63 bl[63] br[63] wl[101] vdd gnd cell_6t
Xbit_r102_c63 bl[63] br[63] wl[102] vdd gnd cell_6t
Xbit_r103_c63 bl[63] br[63] wl[103] vdd gnd cell_6t
Xbit_r104_c63 bl[63] br[63] wl[104] vdd gnd cell_6t
Xbit_r105_c63 bl[63] br[63] wl[105] vdd gnd cell_6t
Xbit_r106_c63 bl[63] br[63] wl[106] vdd gnd cell_6t
Xbit_r107_c63 bl[63] br[63] wl[107] vdd gnd cell_6t
Xbit_r108_c63 bl[63] br[63] wl[108] vdd gnd cell_6t
Xbit_r109_c63 bl[63] br[63] wl[109] vdd gnd cell_6t
Xbit_r110_c63 bl[63] br[63] wl[110] vdd gnd cell_6t
Xbit_r111_c63 bl[63] br[63] wl[111] vdd gnd cell_6t
Xbit_r112_c63 bl[63] br[63] wl[112] vdd gnd cell_6t
Xbit_r113_c63 bl[63] br[63] wl[113] vdd gnd cell_6t
Xbit_r114_c63 bl[63] br[63] wl[114] vdd gnd cell_6t
Xbit_r115_c63 bl[63] br[63] wl[115] vdd gnd cell_6t
Xbit_r116_c63 bl[63] br[63] wl[116] vdd gnd cell_6t
Xbit_r117_c63 bl[63] br[63] wl[117] vdd gnd cell_6t
Xbit_r118_c63 bl[63] br[63] wl[118] vdd gnd cell_6t
Xbit_r119_c63 bl[63] br[63] wl[119] vdd gnd cell_6t
Xbit_r120_c63 bl[63] br[63] wl[120] vdd gnd cell_6t
Xbit_r121_c63 bl[63] br[63] wl[121] vdd gnd cell_6t
Xbit_r122_c63 bl[63] br[63] wl[122] vdd gnd cell_6t
Xbit_r123_c63 bl[63] br[63] wl[123] vdd gnd cell_6t
Xbit_r124_c63 bl[63] br[63] wl[124] vdd gnd cell_6t
Xbit_r125_c63 bl[63] br[63] wl[125] vdd gnd cell_6t
Xbit_r126_c63 bl[63] br[63] wl[126] vdd gnd cell_6t
Xbit_r127_c63 bl[63] br[63] wl[127] vdd gnd cell_6t
Xbit_r128_c63 bl[63] br[63] wl[128] vdd gnd cell_6t
Xbit_r129_c63 bl[63] br[63] wl[129] vdd gnd cell_6t
Xbit_r130_c63 bl[63] br[63] wl[130] vdd gnd cell_6t
Xbit_r131_c63 bl[63] br[63] wl[131] vdd gnd cell_6t
Xbit_r132_c63 bl[63] br[63] wl[132] vdd gnd cell_6t
Xbit_r133_c63 bl[63] br[63] wl[133] vdd gnd cell_6t
Xbit_r134_c63 bl[63] br[63] wl[134] vdd gnd cell_6t
Xbit_r135_c63 bl[63] br[63] wl[135] vdd gnd cell_6t
Xbit_r136_c63 bl[63] br[63] wl[136] vdd gnd cell_6t
Xbit_r137_c63 bl[63] br[63] wl[137] vdd gnd cell_6t
Xbit_r138_c63 bl[63] br[63] wl[138] vdd gnd cell_6t
Xbit_r139_c63 bl[63] br[63] wl[139] vdd gnd cell_6t
Xbit_r140_c63 bl[63] br[63] wl[140] vdd gnd cell_6t
Xbit_r141_c63 bl[63] br[63] wl[141] vdd gnd cell_6t
Xbit_r142_c63 bl[63] br[63] wl[142] vdd gnd cell_6t
Xbit_r143_c63 bl[63] br[63] wl[143] vdd gnd cell_6t
Xbit_r144_c63 bl[63] br[63] wl[144] vdd gnd cell_6t
Xbit_r145_c63 bl[63] br[63] wl[145] vdd gnd cell_6t
Xbit_r146_c63 bl[63] br[63] wl[146] vdd gnd cell_6t
Xbit_r147_c63 bl[63] br[63] wl[147] vdd gnd cell_6t
Xbit_r148_c63 bl[63] br[63] wl[148] vdd gnd cell_6t
Xbit_r149_c63 bl[63] br[63] wl[149] vdd gnd cell_6t
Xbit_r150_c63 bl[63] br[63] wl[150] vdd gnd cell_6t
Xbit_r151_c63 bl[63] br[63] wl[151] vdd gnd cell_6t
Xbit_r152_c63 bl[63] br[63] wl[152] vdd gnd cell_6t
Xbit_r153_c63 bl[63] br[63] wl[153] vdd gnd cell_6t
Xbit_r154_c63 bl[63] br[63] wl[154] vdd gnd cell_6t
Xbit_r155_c63 bl[63] br[63] wl[155] vdd gnd cell_6t
Xbit_r156_c63 bl[63] br[63] wl[156] vdd gnd cell_6t
Xbit_r157_c63 bl[63] br[63] wl[157] vdd gnd cell_6t
Xbit_r158_c63 bl[63] br[63] wl[158] vdd gnd cell_6t
Xbit_r159_c63 bl[63] br[63] wl[159] vdd gnd cell_6t
Xbit_r160_c63 bl[63] br[63] wl[160] vdd gnd cell_6t
Xbit_r161_c63 bl[63] br[63] wl[161] vdd gnd cell_6t
Xbit_r162_c63 bl[63] br[63] wl[162] vdd gnd cell_6t
Xbit_r163_c63 bl[63] br[63] wl[163] vdd gnd cell_6t
Xbit_r164_c63 bl[63] br[63] wl[164] vdd gnd cell_6t
Xbit_r165_c63 bl[63] br[63] wl[165] vdd gnd cell_6t
Xbit_r166_c63 bl[63] br[63] wl[166] vdd gnd cell_6t
Xbit_r167_c63 bl[63] br[63] wl[167] vdd gnd cell_6t
Xbit_r168_c63 bl[63] br[63] wl[168] vdd gnd cell_6t
Xbit_r169_c63 bl[63] br[63] wl[169] vdd gnd cell_6t
Xbit_r170_c63 bl[63] br[63] wl[170] vdd gnd cell_6t
Xbit_r171_c63 bl[63] br[63] wl[171] vdd gnd cell_6t
Xbit_r172_c63 bl[63] br[63] wl[172] vdd gnd cell_6t
Xbit_r173_c63 bl[63] br[63] wl[173] vdd gnd cell_6t
Xbit_r174_c63 bl[63] br[63] wl[174] vdd gnd cell_6t
Xbit_r175_c63 bl[63] br[63] wl[175] vdd gnd cell_6t
Xbit_r176_c63 bl[63] br[63] wl[176] vdd gnd cell_6t
Xbit_r177_c63 bl[63] br[63] wl[177] vdd gnd cell_6t
Xbit_r178_c63 bl[63] br[63] wl[178] vdd gnd cell_6t
Xbit_r179_c63 bl[63] br[63] wl[179] vdd gnd cell_6t
Xbit_r180_c63 bl[63] br[63] wl[180] vdd gnd cell_6t
Xbit_r181_c63 bl[63] br[63] wl[181] vdd gnd cell_6t
Xbit_r182_c63 bl[63] br[63] wl[182] vdd gnd cell_6t
Xbit_r183_c63 bl[63] br[63] wl[183] vdd gnd cell_6t
Xbit_r184_c63 bl[63] br[63] wl[184] vdd gnd cell_6t
Xbit_r185_c63 bl[63] br[63] wl[185] vdd gnd cell_6t
Xbit_r186_c63 bl[63] br[63] wl[186] vdd gnd cell_6t
Xbit_r187_c63 bl[63] br[63] wl[187] vdd gnd cell_6t
Xbit_r188_c63 bl[63] br[63] wl[188] vdd gnd cell_6t
Xbit_r189_c63 bl[63] br[63] wl[189] vdd gnd cell_6t
Xbit_r190_c63 bl[63] br[63] wl[190] vdd gnd cell_6t
Xbit_r191_c63 bl[63] br[63] wl[191] vdd gnd cell_6t
Xbit_r192_c63 bl[63] br[63] wl[192] vdd gnd cell_6t
Xbit_r193_c63 bl[63] br[63] wl[193] vdd gnd cell_6t
Xbit_r194_c63 bl[63] br[63] wl[194] vdd gnd cell_6t
Xbit_r195_c63 bl[63] br[63] wl[195] vdd gnd cell_6t
Xbit_r196_c63 bl[63] br[63] wl[196] vdd gnd cell_6t
Xbit_r197_c63 bl[63] br[63] wl[197] vdd gnd cell_6t
Xbit_r198_c63 bl[63] br[63] wl[198] vdd gnd cell_6t
Xbit_r199_c63 bl[63] br[63] wl[199] vdd gnd cell_6t
Xbit_r200_c63 bl[63] br[63] wl[200] vdd gnd cell_6t
Xbit_r201_c63 bl[63] br[63] wl[201] vdd gnd cell_6t
Xbit_r202_c63 bl[63] br[63] wl[202] vdd gnd cell_6t
Xbit_r203_c63 bl[63] br[63] wl[203] vdd gnd cell_6t
Xbit_r204_c63 bl[63] br[63] wl[204] vdd gnd cell_6t
Xbit_r205_c63 bl[63] br[63] wl[205] vdd gnd cell_6t
Xbit_r206_c63 bl[63] br[63] wl[206] vdd gnd cell_6t
Xbit_r207_c63 bl[63] br[63] wl[207] vdd gnd cell_6t
Xbit_r208_c63 bl[63] br[63] wl[208] vdd gnd cell_6t
Xbit_r209_c63 bl[63] br[63] wl[209] vdd gnd cell_6t
Xbit_r210_c63 bl[63] br[63] wl[210] vdd gnd cell_6t
Xbit_r211_c63 bl[63] br[63] wl[211] vdd gnd cell_6t
Xbit_r212_c63 bl[63] br[63] wl[212] vdd gnd cell_6t
Xbit_r213_c63 bl[63] br[63] wl[213] vdd gnd cell_6t
Xbit_r214_c63 bl[63] br[63] wl[214] vdd gnd cell_6t
Xbit_r215_c63 bl[63] br[63] wl[215] vdd gnd cell_6t
Xbit_r216_c63 bl[63] br[63] wl[216] vdd gnd cell_6t
Xbit_r217_c63 bl[63] br[63] wl[217] vdd gnd cell_6t
Xbit_r218_c63 bl[63] br[63] wl[218] vdd gnd cell_6t
Xbit_r219_c63 bl[63] br[63] wl[219] vdd gnd cell_6t
Xbit_r220_c63 bl[63] br[63] wl[220] vdd gnd cell_6t
Xbit_r221_c63 bl[63] br[63] wl[221] vdd gnd cell_6t
Xbit_r222_c63 bl[63] br[63] wl[222] vdd gnd cell_6t
Xbit_r223_c63 bl[63] br[63] wl[223] vdd gnd cell_6t
Xbit_r224_c63 bl[63] br[63] wl[224] vdd gnd cell_6t
Xbit_r225_c63 bl[63] br[63] wl[225] vdd gnd cell_6t
Xbit_r226_c63 bl[63] br[63] wl[226] vdd gnd cell_6t
Xbit_r227_c63 bl[63] br[63] wl[227] vdd gnd cell_6t
Xbit_r228_c63 bl[63] br[63] wl[228] vdd gnd cell_6t
Xbit_r229_c63 bl[63] br[63] wl[229] vdd gnd cell_6t
Xbit_r230_c63 bl[63] br[63] wl[230] vdd gnd cell_6t
Xbit_r231_c63 bl[63] br[63] wl[231] vdd gnd cell_6t
Xbit_r232_c63 bl[63] br[63] wl[232] vdd gnd cell_6t
Xbit_r233_c63 bl[63] br[63] wl[233] vdd gnd cell_6t
Xbit_r234_c63 bl[63] br[63] wl[234] vdd gnd cell_6t
Xbit_r235_c63 bl[63] br[63] wl[235] vdd gnd cell_6t
Xbit_r236_c63 bl[63] br[63] wl[236] vdd gnd cell_6t
Xbit_r237_c63 bl[63] br[63] wl[237] vdd gnd cell_6t
Xbit_r238_c63 bl[63] br[63] wl[238] vdd gnd cell_6t
Xbit_r239_c63 bl[63] br[63] wl[239] vdd gnd cell_6t
Xbit_r240_c63 bl[63] br[63] wl[240] vdd gnd cell_6t
Xbit_r241_c63 bl[63] br[63] wl[241] vdd gnd cell_6t
Xbit_r242_c63 bl[63] br[63] wl[242] vdd gnd cell_6t
Xbit_r243_c63 bl[63] br[63] wl[243] vdd gnd cell_6t
Xbit_r244_c63 bl[63] br[63] wl[244] vdd gnd cell_6t
Xbit_r245_c63 bl[63] br[63] wl[245] vdd gnd cell_6t
Xbit_r246_c63 bl[63] br[63] wl[246] vdd gnd cell_6t
Xbit_r247_c63 bl[63] br[63] wl[247] vdd gnd cell_6t
Xbit_r248_c63 bl[63] br[63] wl[248] vdd gnd cell_6t
Xbit_r249_c63 bl[63] br[63] wl[249] vdd gnd cell_6t
Xbit_r250_c63 bl[63] br[63] wl[250] vdd gnd cell_6t
Xbit_r251_c63 bl[63] br[63] wl[251] vdd gnd cell_6t
Xbit_r252_c63 bl[63] br[63] wl[252] vdd gnd cell_6t
Xbit_r253_c63 bl[63] br[63] wl[253] vdd gnd cell_6t
Xbit_r254_c63 bl[63] br[63] wl[254] vdd gnd cell_6t
Xbit_r255_c63 bl[63] br[63] wl[255] vdd gnd cell_6t
Xbit_r256_c63 bl[63] br[63] wl[256] vdd gnd cell_6t
Xbit_r257_c63 bl[63] br[63] wl[257] vdd gnd cell_6t
Xbit_r258_c63 bl[63] br[63] wl[258] vdd gnd cell_6t
Xbit_r259_c63 bl[63] br[63] wl[259] vdd gnd cell_6t
Xbit_r260_c63 bl[63] br[63] wl[260] vdd gnd cell_6t
Xbit_r261_c63 bl[63] br[63] wl[261] vdd gnd cell_6t
Xbit_r262_c63 bl[63] br[63] wl[262] vdd gnd cell_6t
Xbit_r263_c63 bl[63] br[63] wl[263] vdd gnd cell_6t
Xbit_r264_c63 bl[63] br[63] wl[264] vdd gnd cell_6t
Xbit_r265_c63 bl[63] br[63] wl[265] vdd gnd cell_6t
Xbit_r266_c63 bl[63] br[63] wl[266] vdd gnd cell_6t
Xbit_r267_c63 bl[63] br[63] wl[267] vdd gnd cell_6t
Xbit_r268_c63 bl[63] br[63] wl[268] vdd gnd cell_6t
Xbit_r269_c63 bl[63] br[63] wl[269] vdd gnd cell_6t
Xbit_r270_c63 bl[63] br[63] wl[270] vdd gnd cell_6t
Xbit_r271_c63 bl[63] br[63] wl[271] vdd gnd cell_6t
Xbit_r272_c63 bl[63] br[63] wl[272] vdd gnd cell_6t
Xbit_r273_c63 bl[63] br[63] wl[273] vdd gnd cell_6t
Xbit_r274_c63 bl[63] br[63] wl[274] vdd gnd cell_6t
Xbit_r275_c63 bl[63] br[63] wl[275] vdd gnd cell_6t
Xbit_r276_c63 bl[63] br[63] wl[276] vdd gnd cell_6t
Xbit_r277_c63 bl[63] br[63] wl[277] vdd gnd cell_6t
Xbit_r278_c63 bl[63] br[63] wl[278] vdd gnd cell_6t
Xbit_r279_c63 bl[63] br[63] wl[279] vdd gnd cell_6t
Xbit_r280_c63 bl[63] br[63] wl[280] vdd gnd cell_6t
Xbit_r281_c63 bl[63] br[63] wl[281] vdd gnd cell_6t
Xbit_r282_c63 bl[63] br[63] wl[282] vdd gnd cell_6t
Xbit_r283_c63 bl[63] br[63] wl[283] vdd gnd cell_6t
Xbit_r284_c63 bl[63] br[63] wl[284] vdd gnd cell_6t
Xbit_r285_c63 bl[63] br[63] wl[285] vdd gnd cell_6t
Xbit_r286_c63 bl[63] br[63] wl[286] vdd gnd cell_6t
Xbit_r287_c63 bl[63] br[63] wl[287] vdd gnd cell_6t
Xbit_r288_c63 bl[63] br[63] wl[288] vdd gnd cell_6t
Xbit_r289_c63 bl[63] br[63] wl[289] vdd gnd cell_6t
Xbit_r290_c63 bl[63] br[63] wl[290] vdd gnd cell_6t
Xbit_r291_c63 bl[63] br[63] wl[291] vdd gnd cell_6t
Xbit_r292_c63 bl[63] br[63] wl[292] vdd gnd cell_6t
Xbit_r293_c63 bl[63] br[63] wl[293] vdd gnd cell_6t
Xbit_r294_c63 bl[63] br[63] wl[294] vdd gnd cell_6t
Xbit_r295_c63 bl[63] br[63] wl[295] vdd gnd cell_6t
Xbit_r296_c63 bl[63] br[63] wl[296] vdd gnd cell_6t
Xbit_r297_c63 bl[63] br[63] wl[297] vdd gnd cell_6t
Xbit_r298_c63 bl[63] br[63] wl[298] vdd gnd cell_6t
Xbit_r299_c63 bl[63] br[63] wl[299] vdd gnd cell_6t
Xbit_r300_c63 bl[63] br[63] wl[300] vdd gnd cell_6t
Xbit_r301_c63 bl[63] br[63] wl[301] vdd gnd cell_6t
Xbit_r302_c63 bl[63] br[63] wl[302] vdd gnd cell_6t
Xbit_r303_c63 bl[63] br[63] wl[303] vdd gnd cell_6t
Xbit_r304_c63 bl[63] br[63] wl[304] vdd gnd cell_6t
Xbit_r305_c63 bl[63] br[63] wl[305] vdd gnd cell_6t
Xbit_r306_c63 bl[63] br[63] wl[306] vdd gnd cell_6t
Xbit_r307_c63 bl[63] br[63] wl[307] vdd gnd cell_6t
Xbit_r308_c63 bl[63] br[63] wl[308] vdd gnd cell_6t
Xbit_r309_c63 bl[63] br[63] wl[309] vdd gnd cell_6t
Xbit_r310_c63 bl[63] br[63] wl[310] vdd gnd cell_6t
Xbit_r311_c63 bl[63] br[63] wl[311] vdd gnd cell_6t
Xbit_r312_c63 bl[63] br[63] wl[312] vdd gnd cell_6t
Xbit_r313_c63 bl[63] br[63] wl[313] vdd gnd cell_6t
Xbit_r314_c63 bl[63] br[63] wl[314] vdd gnd cell_6t
Xbit_r315_c63 bl[63] br[63] wl[315] vdd gnd cell_6t
Xbit_r316_c63 bl[63] br[63] wl[316] vdd gnd cell_6t
Xbit_r317_c63 bl[63] br[63] wl[317] vdd gnd cell_6t
Xbit_r318_c63 bl[63] br[63] wl[318] vdd gnd cell_6t
Xbit_r319_c63 bl[63] br[63] wl[319] vdd gnd cell_6t
Xbit_r320_c63 bl[63] br[63] wl[320] vdd gnd cell_6t
Xbit_r321_c63 bl[63] br[63] wl[321] vdd gnd cell_6t
Xbit_r322_c63 bl[63] br[63] wl[322] vdd gnd cell_6t
Xbit_r323_c63 bl[63] br[63] wl[323] vdd gnd cell_6t
Xbit_r324_c63 bl[63] br[63] wl[324] vdd gnd cell_6t
Xbit_r325_c63 bl[63] br[63] wl[325] vdd gnd cell_6t
Xbit_r326_c63 bl[63] br[63] wl[326] vdd gnd cell_6t
Xbit_r327_c63 bl[63] br[63] wl[327] vdd gnd cell_6t
Xbit_r328_c63 bl[63] br[63] wl[328] vdd gnd cell_6t
Xbit_r329_c63 bl[63] br[63] wl[329] vdd gnd cell_6t
Xbit_r330_c63 bl[63] br[63] wl[330] vdd gnd cell_6t
Xbit_r331_c63 bl[63] br[63] wl[331] vdd gnd cell_6t
Xbit_r332_c63 bl[63] br[63] wl[332] vdd gnd cell_6t
Xbit_r333_c63 bl[63] br[63] wl[333] vdd gnd cell_6t
Xbit_r334_c63 bl[63] br[63] wl[334] vdd gnd cell_6t
Xbit_r335_c63 bl[63] br[63] wl[335] vdd gnd cell_6t
Xbit_r336_c63 bl[63] br[63] wl[336] vdd gnd cell_6t
Xbit_r337_c63 bl[63] br[63] wl[337] vdd gnd cell_6t
Xbit_r338_c63 bl[63] br[63] wl[338] vdd gnd cell_6t
Xbit_r339_c63 bl[63] br[63] wl[339] vdd gnd cell_6t
Xbit_r340_c63 bl[63] br[63] wl[340] vdd gnd cell_6t
Xbit_r341_c63 bl[63] br[63] wl[341] vdd gnd cell_6t
Xbit_r342_c63 bl[63] br[63] wl[342] vdd gnd cell_6t
Xbit_r343_c63 bl[63] br[63] wl[343] vdd gnd cell_6t
Xbit_r344_c63 bl[63] br[63] wl[344] vdd gnd cell_6t
Xbit_r345_c63 bl[63] br[63] wl[345] vdd gnd cell_6t
Xbit_r346_c63 bl[63] br[63] wl[346] vdd gnd cell_6t
Xbit_r347_c63 bl[63] br[63] wl[347] vdd gnd cell_6t
Xbit_r348_c63 bl[63] br[63] wl[348] vdd gnd cell_6t
Xbit_r349_c63 bl[63] br[63] wl[349] vdd gnd cell_6t
Xbit_r350_c63 bl[63] br[63] wl[350] vdd gnd cell_6t
Xbit_r351_c63 bl[63] br[63] wl[351] vdd gnd cell_6t
Xbit_r352_c63 bl[63] br[63] wl[352] vdd gnd cell_6t
Xbit_r353_c63 bl[63] br[63] wl[353] vdd gnd cell_6t
Xbit_r354_c63 bl[63] br[63] wl[354] vdd gnd cell_6t
Xbit_r355_c63 bl[63] br[63] wl[355] vdd gnd cell_6t
Xbit_r356_c63 bl[63] br[63] wl[356] vdd gnd cell_6t
Xbit_r357_c63 bl[63] br[63] wl[357] vdd gnd cell_6t
Xbit_r358_c63 bl[63] br[63] wl[358] vdd gnd cell_6t
Xbit_r359_c63 bl[63] br[63] wl[359] vdd gnd cell_6t
Xbit_r360_c63 bl[63] br[63] wl[360] vdd gnd cell_6t
Xbit_r361_c63 bl[63] br[63] wl[361] vdd gnd cell_6t
Xbit_r362_c63 bl[63] br[63] wl[362] vdd gnd cell_6t
Xbit_r363_c63 bl[63] br[63] wl[363] vdd gnd cell_6t
Xbit_r364_c63 bl[63] br[63] wl[364] vdd gnd cell_6t
Xbit_r365_c63 bl[63] br[63] wl[365] vdd gnd cell_6t
Xbit_r366_c63 bl[63] br[63] wl[366] vdd gnd cell_6t
Xbit_r367_c63 bl[63] br[63] wl[367] vdd gnd cell_6t
Xbit_r368_c63 bl[63] br[63] wl[368] vdd gnd cell_6t
Xbit_r369_c63 bl[63] br[63] wl[369] vdd gnd cell_6t
Xbit_r370_c63 bl[63] br[63] wl[370] vdd gnd cell_6t
Xbit_r371_c63 bl[63] br[63] wl[371] vdd gnd cell_6t
Xbit_r372_c63 bl[63] br[63] wl[372] vdd gnd cell_6t
Xbit_r373_c63 bl[63] br[63] wl[373] vdd gnd cell_6t
Xbit_r374_c63 bl[63] br[63] wl[374] vdd gnd cell_6t
Xbit_r375_c63 bl[63] br[63] wl[375] vdd gnd cell_6t
Xbit_r376_c63 bl[63] br[63] wl[376] vdd gnd cell_6t
Xbit_r377_c63 bl[63] br[63] wl[377] vdd gnd cell_6t
Xbit_r378_c63 bl[63] br[63] wl[378] vdd gnd cell_6t
Xbit_r379_c63 bl[63] br[63] wl[379] vdd gnd cell_6t
Xbit_r380_c63 bl[63] br[63] wl[380] vdd gnd cell_6t
Xbit_r381_c63 bl[63] br[63] wl[381] vdd gnd cell_6t
Xbit_r382_c63 bl[63] br[63] wl[382] vdd gnd cell_6t
Xbit_r383_c63 bl[63] br[63] wl[383] vdd gnd cell_6t
Xbit_r384_c63 bl[63] br[63] wl[384] vdd gnd cell_6t
Xbit_r385_c63 bl[63] br[63] wl[385] vdd gnd cell_6t
Xbit_r386_c63 bl[63] br[63] wl[386] vdd gnd cell_6t
Xbit_r387_c63 bl[63] br[63] wl[387] vdd gnd cell_6t
Xbit_r388_c63 bl[63] br[63] wl[388] vdd gnd cell_6t
Xbit_r389_c63 bl[63] br[63] wl[389] vdd gnd cell_6t
Xbit_r390_c63 bl[63] br[63] wl[390] vdd gnd cell_6t
Xbit_r391_c63 bl[63] br[63] wl[391] vdd gnd cell_6t
Xbit_r392_c63 bl[63] br[63] wl[392] vdd gnd cell_6t
Xbit_r393_c63 bl[63] br[63] wl[393] vdd gnd cell_6t
Xbit_r394_c63 bl[63] br[63] wl[394] vdd gnd cell_6t
Xbit_r395_c63 bl[63] br[63] wl[395] vdd gnd cell_6t
Xbit_r396_c63 bl[63] br[63] wl[396] vdd gnd cell_6t
Xbit_r397_c63 bl[63] br[63] wl[397] vdd gnd cell_6t
Xbit_r398_c63 bl[63] br[63] wl[398] vdd gnd cell_6t
Xbit_r399_c63 bl[63] br[63] wl[399] vdd gnd cell_6t
Xbit_r400_c63 bl[63] br[63] wl[400] vdd gnd cell_6t
Xbit_r401_c63 bl[63] br[63] wl[401] vdd gnd cell_6t
Xbit_r402_c63 bl[63] br[63] wl[402] vdd gnd cell_6t
Xbit_r403_c63 bl[63] br[63] wl[403] vdd gnd cell_6t
Xbit_r404_c63 bl[63] br[63] wl[404] vdd gnd cell_6t
Xbit_r405_c63 bl[63] br[63] wl[405] vdd gnd cell_6t
Xbit_r406_c63 bl[63] br[63] wl[406] vdd gnd cell_6t
Xbit_r407_c63 bl[63] br[63] wl[407] vdd gnd cell_6t
Xbit_r408_c63 bl[63] br[63] wl[408] vdd gnd cell_6t
Xbit_r409_c63 bl[63] br[63] wl[409] vdd gnd cell_6t
Xbit_r410_c63 bl[63] br[63] wl[410] vdd gnd cell_6t
Xbit_r411_c63 bl[63] br[63] wl[411] vdd gnd cell_6t
Xbit_r412_c63 bl[63] br[63] wl[412] vdd gnd cell_6t
Xbit_r413_c63 bl[63] br[63] wl[413] vdd gnd cell_6t
Xbit_r414_c63 bl[63] br[63] wl[414] vdd gnd cell_6t
Xbit_r415_c63 bl[63] br[63] wl[415] vdd gnd cell_6t
Xbit_r416_c63 bl[63] br[63] wl[416] vdd gnd cell_6t
Xbit_r417_c63 bl[63] br[63] wl[417] vdd gnd cell_6t
Xbit_r418_c63 bl[63] br[63] wl[418] vdd gnd cell_6t
Xbit_r419_c63 bl[63] br[63] wl[419] vdd gnd cell_6t
Xbit_r420_c63 bl[63] br[63] wl[420] vdd gnd cell_6t
Xbit_r421_c63 bl[63] br[63] wl[421] vdd gnd cell_6t
Xbit_r422_c63 bl[63] br[63] wl[422] vdd gnd cell_6t
Xbit_r423_c63 bl[63] br[63] wl[423] vdd gnd cell_6t
Xbit_r424_c63 bl[63] br[63] wl[424] vdd gnd cell_6t
Xbit_r425_c63 bl[63] br[63] wl[425] vdd gnd cell_6t
Xbit_r426_c63 bl[63] br[63] wl[426] vdd gnd cell_6t
Xbit_r427_c63 bl[63] br[63] wl[427] vdd gnd cell_6t
Xbit_r428_c63 bl[63] br[63] wl[428] vdd gnd cell_6t
Xbit_r429_c63 bl[63] br[63] wl[429] vdd gnd cell_6t
Xbit_r430_c63 bl[63] br[63] wl[430] vdd gnd cell_6t
Xbit_r431_c63 bl[63] br[63] wl[431] vdd gnd cell_6t
Xbit_r432_c63 bl[63] br[63] wl[432] vdd gnd cell_6t
Xbit_r433_c63 bl[63] br[63] wl[433] vdd gnd cell_6t
Xbit_r434_c63 bl[63] br[63] wl[434] vdd gnd cell_6t
Xbit_r435_c63 bl[63] br[63] wl[435] vdd gnd cell_6t
Xbit_r436_c63 bl[63] br[63] wl[436] vdd gnd cell_6t
Xbit_r437_c63 bl[63] br[63] wl[437] vdd gnd cell_6t
Xbit_r438_c63 bl[63] br[63] wl[438] vdd gnd cell_6t
Xbit_r439_c63 bl[63] br[63] wl[439] vdd gnd cell_6t
Xbit_r440_c63 bl[63] br[63] wl[440] vdd gnd cell_6t
Xbit_r441_c63 bl[63] br[63] wl[441] vdd gnd cell_6t
Xbit_r442_c63 bl[63] br[63] wl[442] vdd gnd cell_6t
Xbit_r443_c63 bl[63] br[63] wl[443] vdd gnd cell_6t
Xbit_r444_c63 bl[63] br[63] wl[444] vdd gnd cell_6t
Xbit_r445_c63 bl[63] br[63] wl[445] vdd gnd cell_6t
Xbit_r446_c63 bl[63] br[63] wl[446] vdd gnd cell_6t
Xbit_r447_c63 bl[63] br[63] wl[447] vdd gnd cell_6t
Xbit_r448_c63 bl[63] br[63] wl[448] vdd gnd cell_6t
Xbit_r449_c63 bl[63] br[63] wl[449] vdd gnd cell_6t
Xbit_r450_c63 bl[63] br[63] wl[450] vdd gnd cell_6t
Xbit_r451_c63 bl[63] br[63] wl[451] vdd gnd cell_6t
Xbit_r452_c63 bl[63] br[63] wl[452] vdd gnd cell_6t
Xbit_r453_c63 bl[63] br[63] wl[453] vdd gnd cell_6t
Xbit_r454_c63 bl[63] br[63] wl[454] vdd gnd cell_6t
Xbit_r455_c63 bl[63] br[63] wl[455] vdd gnd cell_6t
Xbit_r456_c63 bl[63] br[63] wl[456] vdd gnd cell_6t
Xbit_r457_c63 bl[63] br[63] wl[457] vdd gnd cell_6t
Xbit_r458_c63 bl[63] br[63] wl[458] vdd gnd cell_6t
Xbit_r459_c63 bl[63] br[63] wl[459] vdd gnd cell_6t
Xbit_r460_c63 bl[63] br[63] wl[460] vdd gnd cell_6t
Xbit_r461_c63 bl[63] br[63] wl[461] vdd gnd cell_6t
Xbit_r462_c63 bl[63] br[63] wl[462] vdd gnd cell_6t
Xbit_r463_c63 bl[63] br[63] wl[463] vdd gnd cell_6t
Xbit_r464_c63 bl[63] br[63] wl[464] vdd gnd cell_6t
Xbit_r465_c63 bl[63] br[63] wl[465] vdd gnd cell_6t
Xbit_r466_c63 bl[63] br[63] wl[466] vdd gnd cell_6t
Xbit_r467_c63 bl[63] br[63] wl[467] vdd gnd cell_6t
Xbit_r468_c63 bl[63] br[63] wl[468] vdd gnd cell_6t
Xbit_r469_c63 bl[63] br[63] wl[469] vdd gnd cell_6t
Xbit_r470_c63 bl[63] br[63] wl[470] vdd gnd cell_6t
Xbit_r471_c63 bl[63] br[63] wl[471] vdd gnd cell_6t
Xbit_r472_c63 bl[63] br[63] wl[472] vdd gnd cell_6t
Xbit_r473_c63 bl[63] br[63] wl[473] vdd gnd cell_6t
Xbit_r474_c63 bl[63] br[63] wl[474] vdd gnd cell_6t
Xbit_r475_c63 bl[63] br[63] wl[475] vdd gnd cell_6t
Xbit_r476_c63 bl[63] br[63] wl[476] vdd gnd cell_6t
Xbit_r477_c63 bl[63] br[63] wl[477] vdd gnd cell_6t
Xbit_r478_c63 bl[63] br[63] wl[478] vdd gnd cell_6t
Xbit_r479_c63 bl[63] br[63] wl[479] vdd gnd cell_6t
Xbit_r480_c63 bl[63] br[63] wl[480] vdd gnd cell_6t
Xbit_r481_c63 bl[63] br[63] wl[481] vdd gnd cell_6t
Xbit_r482_c63 bl[63] br[63] wl[482] vdd gnd cell_6t
Xbit_r483_c63 bl[63] br[63] wl[483] vdd gnd cell_6t
Xbit_r484_c63 bl[63] br[63] wl[484] vdd gnd cell_6t
Xbit_r485_c63 bl[63] br[63] wl[485] vdd gnd cell_6t
Xbit_r486_c63 bl[63] br[63] wl[486] vdd gnd cell_6t
Xbit_r487_c63 bl[63] br[63] wl[487] vdd gnd cell_6t
Xbit_r488_c63 bl[63] br[63] wl[488] vdd gnd cell_6t
Xbit_r489_c63 bl[63] br[63] wl[489] vdd gnd cell_6t
Xbit_r490_c63 bl[63] br[63] wl[490] vdd gnd cell_6t
Xbit_r491_c63 bl[63] br[63] wl[491] vdd gnd cell_6t
Xbit_r492_c63 bl[63] br[63] wl[492] vdd gnd cell_6t
Xbit_r493_c63 bl[63] br[63] wl[493] vdd gnd cell_6t
Xbit_r494_c63 bl[63] br[63] wl[494] vdd gnd cell_6t
Xbit_r495_c63 bl[63] br[63] wl[495] vdd gnd cell_6t
Xbit_r496_c63 bl[63] br[63] wl[496] vdd gnd cell_6t
Xbit_r497_c63 bl[63] br[63] wl[497] vdd gnd cell_6t
Xbit_r498_c63 bl[63] br[63] wl[498] vdd gnd cell_6t
Xbit_r499_c63 bl[63] br[63] wl[499] vdd gnd cell_6t
Xbit_r500_c63 bl[63] br[63] wl[500] vdd gnd cell_6t
Xbit_r501_c63 bl[63] br[63] wl[501] vdd gnd cell_6t
Xbit_r502_c63 bl[63] br[63] wl[502] vdd gnd cell_6t
Xbit_r503_c63 bl[63] br[63] wl[503] vdd gnd cell_6t
Xbit_r504_c63 bl[63] br[63] wl[504] vdd gnd cell_6t
Xbit_r505_c63 bl[63] br[63] wl[505] vdd gnd cell_6t
Xbit_r506_c63 bl[63] br[63] wl[506] vdd gnd cell_6t
Xbit_r507_c63 bl[63] br[63] wl[507] vdd gnd cell_6t
Xbit_r508_c63 bl[63] br[63] wl[508] vdd gnd cell_6t
Xbit_r509_c63 bl[63] br[63] wl[509] vdd gnd cell_6t
Xbit_r510_c63 bl[63] br[63] wl[510] vdd gnd cell_6t
Xbit_r511_c63 bl[63] br[63] wl[511] vdd gnd cell_6t
Xbit_r0_c64 bl[64] br[64] wl[0] vdd gnd cell_6t
Xbit_r1_c64 bl[64] br[64] wl[1] vdd gnd cell_6t
Xbit_r2_c64 bl[64] br[64] wl[2] vdd gnd cell_6t
Xbit_r3_c64 bl[64] br[64] wl[3] vdd gnd cell_6t
Xbit_r4_c64 bl[64] br[64] wl[4] vdd gnd cell_6t
Xbit_r5_c64 bl[64] br[64] wl[5] vdd gnd cell_6t
Xbit_r6_c64 bl[64] br[64] wl[6] vdd gnd cell_6t
Xbit_r7_c64 bl[64] br[64] wl[7] vdd gnd cell_6t
Xbit_r8_c64 bl[64] br[64] wl[8] vdd gnd cell_6t
Xbit_r9_c64 bl[64] br[64] wl[9] vdd gnd cell_6t
Xbit_r10_c64 bl[64] br[64] wl[10] vdd gnd cell_6t
Xbit_r11_c64 bl[64] br[64] wl[11] vdd gnd cell_6t
Xbit_r12_c64 bl[64] br[64] wl[12] vdd gnd cell_6t
Xbit_r13_c64 bl[64] br[64] wl[13] vdd gnd cell_6t
Xbit_r14_c64 bl[64] br[64] wl[14] vdd gnd cell_6t
Xbit_r15_c64 bl[64] br[64] wl[15] vdd gnd cell_6t
Xbit_r16_c64 bl[64] br[64] wl[16] vdd gnd cell_6t
Xbit_r17_c64 bl[64] br[64] wl[17] vdd gnd cell_6t
Xbit_r18_c64 bl[64] br[64] wl[18] vdd gnd cell_6t
Xbit_r19_c64 bl[64] br[64] wl[19] vdd gnd cell_6t
Xbit_r20_c64 bl[64] br[64] wl[20] vdd gnd cell_6t
Xbit_r21_c64 bl[64] br[64] wl[21] vdd gnd cell_6t
Xbit_r22_c64 bl[64] br[64] wl[22] vdd gnd cell_6t
Xbit_r23_c64 bl[64] br[64] wl[23] vdd gnd cell_6t
Xbit_r24_c64 bl[64] br[64] wl[24] vdd gnd cell_6t
Xbit_r25_c64 bl[64] br[64] wl[25] vdd gnd cell_6t
Xbit_r26_c64 bl[64] br[64] wl[26] vdd gnd cell_6t
Xbit_r27_c64 bl[64] br[64] wl[27] vdd gnd cell_6t
Xbit_r28_c64 bl[64] br[64] wl[28] vdd gnd cell_6t
Xbit_r29_c64 bl[64] br[64] wl[29] vdd gnd cell_6t
Xbit_r30_c64 bl[64] br[64] wl[30] vdd gnd cell_6t
Xbit_r31_c64 bl[64] br[64] wl[31] vdd gnd cell_6t
Xbit_r32_c64 bl[64] br[64] wl[32] vdd gnd cell_6t
Xbit_r33_c64 bl[64] br[64] wl[33] vdd gnd cell_6t
Xbit_r34_c64 bl[64] br[64] wl[34] vdd gnd cell_6t
Xbit_r35_c64 bl[64] br[64] wl[35] vdd gnd cell_6t
Xbit_r36_c64 bl[64] br[64] wl[36] vdd gnd cell_6t
Xbit_r37_c64 bl[64] br[64] wl[37] vdd gnd cell_6t
Xbit_r38_c64 bl[64] br[64] wl[38] vdd gnd cell_6t
Xbit_r39_c64 bl[64] br[64] wl[39] vdd gnd cell_6t
Xbit_r40_c64 bl[64] br[64] wl[40] vdd gnd cell_6t
Xbit_r41_c64 bl[64] br[64] wl[41] vdd gnd cell_6t
Xbit_r42_c64 bl[64] br[64] wl[42] vdd gnd cell_6t
Xbit_r43_c64 bl[64] br[64] wl[43] vdd gnd cell_6t
Xbit_r44_c64 bl[64] br[64] wl[44] vdd gnd cell_6t
Xbit_r45_c64 bl[64] br[64] wl[45] vdd gnd cell_6t
Xbit_r46_c64 bl[64] br[64] wl[46] vdd gnd cell_6t
Xbit_r47_c64 bl[64] br[64] wl[47] vdd gnd cell_6t
Xbit_r48_c64 bl[64] br[64] wl[48] vdd gnd cell_6t
Xbit_r49_c64 bl[64] br[64] wl[49] vdd gnd cell_6t
Xbit_r50_c64 bl[64] br[64] wl[50] vdd gnd cell_6t
Xbit_r51_c64 bl[64] br[64] wl[51] vdd gnd cell_6t
Xbit_r52_c64 bl[64] br[64] wl[52] vdd gnd cell_6t
Xbit_r53_c64 bl[64] br[64] wl[53] vdd gnd cell_6t
Xbit_r54_c64 bl[64] br[64] wl[54] vdd gnd cell_6t
Xbit_r55_c64 bl[64] br[64] wl[55] vdd gnd cell_6t
Xbit_r56_c64 bl[64] br[64] wl[56] vdd gnd cell_6t
Xbit_r57_c64 bl[64] br[64] wl[57] vdd gnd cell_6t
Xbit_r58_c64 bl[64] br[64] wl[58] vdd gnd cell_6t
Xbit_r59_c64 bl[64] br[64] wl[59] vdd gnd cell_6t
Xbit_r60_c64 bl[64] br[64] wl[60] vdd gnd cell_6t
Xbit_r61_c64 bl[64] br[64] wl[61] vdd gnd cell_6t
Xbit_r62_c64 bl[64] br[64] wl[62] vdd gnd cell_6t
Xbit_r63_c64 bl[64] br[64] wl[63] vdd gnd cell_6t
Xbit_r64_c64 bl[64] br[64] wl[64] vdd gnd cell_6t
Xbit_r65_c64 bl[64] br[64] wl[65] vdd gnd cell_6t
Xbit_r66_c64 bl[64] br[64] wl[66] vdd gnd cell_6t
Xbit_r67_c64 bl[64] br[64] wl[67] vdd gnd cell_6t
Xbit_r68_c64 bl[64] br[64] wl[68] vdd gnd cell_6t
Xbit_r69_c64 bl[64] br[64] wl[69] vdd gnd cell_6t
Xbit_r70_c64 bl[64] br[64] wl[70] vdd gnd cell_6t
Xbit_r71_c64 bl[64] br[64] wl[71] vdd gnd cell_6t
Xbit_r72_c64 bl[64] br[64] wl[72] vdd gnd cell_6t
Xbit_r73_c64 bl[64] br[64] wl[73] vdd gnd cell_6t
Xbit_r74_c64 bl[64] br[64] wl[74] vdd gnd cell_6t
Xbit_r75_c64 bl[64] br[64] wl[75] vdd gnd cell_6t
Xbit_r76_c64 bl[64] br[64] wl[76] vdd gnd cell_6t
Xbit_r77_c64 bl[64] br[64] wl[77] vdd gnd cell_6t
Xbit_r78_c64 bl[64] br[64] wl[78] vdd gnd cell_6t
Xbit_r79_c64 bl[64] br[64] wl[79] vdd gnd cell_6t
Xbit_r80_c64 bl[64] br[64] wl[80] vdd gnd cell_6t
Xbit_r81_c64 bl[64] br[64] wl[81] vdd gnd cell_6t
Xbit_r82_c64 bl[64] br[64] wl[82] vdd gnd cell_6t
Xbit_r83_c64 bl[64] br[64] wl[83] vdd gnd cell_6t
Xbit_r84_c64 bl[64] br[64] wl[84] vdd gnd cell_6t
Xbit_r85_c64 bl[64] br[64] wl[85] vdd gnd cell_6t
Xbit_r86_c64 bl[64] br[64] wl[86] vdd gnd cell_6t
Xbit_r87_c64 bl[64] br[64] wl[87] vdd gnd cell_6t
Xbit_r88_c64 bl[64] br[64] wl[88] vdd gnd cell_6t
Xbit_r89_c64 bl[64] br[64] wl[89] vdd gnd cell_6t
Xbit_r90_c64 bl[64] br[64] wl[90] vdd gnd cell_6t
Xbit_r91_c64 bl[64] br[64] wl[91] vdd gnd cell_6t
Xbit_r92_c64 bl[64] br[64] wl[92] vdd gnd cell_6t
Xbit_r93_c64 bl[64] br[64] wl[93] vdd gnd cell_6t
Xbit_r94_c64 bl[64] br[64] wl[94] vdd gnd cell_6t
Xbit_r95_c64 bl[64] br[64] wl[95] vdd gnd cell_6t
Xbit_r96_c64 bl[64] br[64] wl[96] vdd gnd cell_6t
Xbit_r97_c64 bl[64] br[64] wl[97] vdd gnd cell_6t
Xbit_r98_c64 bl[64] br[64] wl[98] vdd gnd cell_6t
Xbit_r99_c64 bl[64] br[64] wl[99] vdd gnd cell_6t
Xbit_r100_c64 bl[64] br[64] wl[100] vdd gnd cell_6t
Xbit_r101_c64 bl[64] br[64] wl[101] vdd gnd cell_6t
Xbit_r102_c64 bl[64] br[64] wl[102] vdd gnd cell_6t
Xbit_r103_c64 bl[64] br[64] wl[103] vdd gnd cell_6t
Xbit_r104_c64 bl[64] br[64] wl[104] vdd gnd cell_6t
Xbit_r105_c64 bl[64] br[64] wl[105] vdd gnd cell_6t
Xbit_r106_c64 bl[64] br[64] wl[106] vdd gnd cell_6t
Xbit_r107_c64 bl[64] br[64] wl[107] vdd gnd cell_6t
Xbit_r108_c64 bl[64] br[64] wl[108] vdd gnd cell_6t
Xbit_r109_c64 bl[64] br[64] wl[109] vdd gnd cell_6t
Xbit_r110_c64 bl[64] br[64] wl[110] vdd gnd cell_6t
Xbit_r111_c64 bl[64] br[64] wl[111] vdd gnd cell_6t
Xbit_r112_c64 bl[64] br[64] wl[112] vdd gnd cell_6t
Xbit_r113_c64 bl[64] br[64] wl[113] vdd gnd cell_6t
Xbit_r114_c64 bl[64] br[64] wl[114] vdd gnd cell_6t
Xbit_r115_c64 bl[64] br[64] wl[115] vdd gnd cell_6t
Xbit_r116_c64 bl[64] br[64] wl[116] vdd gnd cell_6t
Xbit_r117_c64 bl[64] br[64] wl[117] vdd gnd cell_6t
Xbit_r118_c64 bl[64] br[64] wl[118] vdd gnd cell_6t
Xbit_r119_c64 bl[64] br[64] wl[119] vdd gnd cell_6t
Xbit_r120_c64 bl[64] br[64] wl[120] vdd gnd cell_6t
Xbit_r121_c64 bl[64] br[64] wl[121] vdd gnd cell_6t
Xbit_r122_c64 bl[64] br[64] wl[122] vdd gnd cell_6t
Xbit_r123_c64 bl[64] br[64] wl[123] vdd gnd cell_6t
Xbit_r124_c64 bl[64] br[64] wl[124] vdd gnd cell_6t
Xbit_r125_c64 bl[64] br[64] wl[125] vdd gnd cell_6t
Xbit_r126_c64 bl[64] br[64] wl[126] vdd gnd cell_6t
Xbit_r127_c64 bl[64] br[64] wl[127] vdd gnd cell_6t
Xbit_r128_c64 bl[64] br[64] wl[128] vdd gnd cell_6t
Xbit_r129_c64 bl[64] br[64] wl[129] vdd gnd cell_6t
Xbit_r130_c64 bl[64] br[64] wl[130] vdd gnd cell_6t
Xbit_r131_c64 bl[64] br[64] wl[131] vdd gnd cell_6t
Xbit_r132_c64 bl[64] br[64] wl[132] vdd gnd cell_6t
Xbit_r133_c64 bl[64] br[64] wl[133] vdd gnd cell_6t
Xbit_r134_c64 bl[64] br[64] wl[134] vdd gnd cell_6t
Xbit_r135_c64 bl[64] br[64] wl[135] vdd gnd cell_6t
Xbit_r136_c64 bl[64] br[64] wl[136] vdd gnd cell_6t
Xbit_r137_c64 bl[64] br[64] wl[137] vdd gnd cell_6t
Xbit_r138_c64 bl[64] br[64] wl[138] vdd gnd cell_6t
Xbit_r139_c64 bl[64] br[64] wl[139] vdd gnd cell_6t
Xbit_r140_c64 bl[64] br[64] wl[140] vdd gnd cell_6t
Xbit_r141_c64 bl[64] br[64] wl[141] vdd gnd cell_6t
Xbit_r142_c64 bl[64] br[64] wl[142] vdd gnd cell_6t
Xbit_r143_c64 bl[64] br[64] wl[143] vdd gnd cell_6t
Xbit_r144_c64 bl[64] br[64] wl[144] vdd gnd cell_6t
Xbit_r145_c64 bl[64] br[64] wl[145] vdd gnd cell_6t
Xbit_r146_c64 bl[64] br[64] wl[146] vdd gnd cell_6t
Xbit_r147_c64 bl[64] br[64] wl[147] vdd gnd cell_6t
Xbit_r148_c64 bl[64] br[64] wl[148] vdd gnd cell_6t
Xbit_r149_c64 bl[64] br[64] wl[149] vdd gnd cell_6t
Xbit_r150_c64 bl[64] br[64] wl[150] vdd gnd cell_6t
Xbit_r151_c64 bl[64] br[64] wl[151] vdd gnd cell_6t
Xbit_r152_c64 bl[64] br[64] wl[152] vdd gnd cell_6t
Xbit_r153_c64 bl[64] br[64] wl[153] vdd gnd cell_6t
Xbit_r154_c64 bl[64] br[64] wl[154] vdd gnd cell_6t
Xbit_r155_c64 bl[64] br[64] wl[155] vdd gnd cell_6t
Xbit_r156_c64 bl[64] br[64] wl[156] vdd gnd cell_6t
Xbit_r157_c64 bl[64] br[64] wl[157] vdd gnd cell_6t
Xbit_r158_c64 bl[64] br[64] wl[158] vdd gnd cell_6t
Xbit_r159_c64 bl[64] br[64] wl[159] vdd gnd cell_6t
Xbit_r160_c64 bl[64] br[64] wl[160] vdd gnd cell_6t
Xbit_r161_c64 bl[64] br[64] wl[161] vdd gnd cell_6t
Xbit_r162_c64 bl[64] br[64] wl[162] vdd gnd cell_6t
Xbit_r163_c64 bl[64] br[64] wl[163] vdd gnd cell_6t
Xbit_r164_c64 bl[64] br[64] wl[164] vdd gnd cell_6t
Xbit_r165_c64 bl[64] br[64] wl[165] vdd gnd cell_6t
Xbit_r166_c64 bl[64] br[64] wl[166] vdd gnd cell_6t
Xbit_r167_c64 bl[64] br[64] wl[167] vdd gnd cell_6t
Xbit_r168_c64 bl[64] br[64] wl[168] vdd gnd cell_6t
Xbit_r169_c64 bl[64] br[64] wl[169] vdd gnd cell_6t
Xbit_r170_c64 bl[64] br[64] wl[170] vdd gnd cell_6t
Xbit_r171_c64 bl[64] br[64] wl[171] vdd gnd cell_6t
Xbit_r172_c64 bl[64] br[64] wl[172] vdd gnd cell_6t
Xbit_r173_c64 bl[64] br[64] wl[173] vdd gnd cell_6t
Xbit_r174_c64 bl[64] br[64] wl[174] vdd gnd cell_6t
Xbit_r175_c64 bl[64] br[64] wl[175] vdd gnd cell_6t
Xbit_r176_c64 bl[64] br[64] wl[176] vdd gnd cell_6t
Xbit_r177_c64 bl[64] br[64] wl[177] vdd gnd cell_6t
Xbit_r178_c64 bl[64] br[64] wl[178] vdd gnd cell_6t
Xbit_r179_c64 bl[64] br[64] wl[179] vdd gnd cell_6t
Xbit_r180_c64 bl[64] br[64] wl[180] vdd gnd cell_6t
Xbit_r181_c64 bl[64] br[64] wl[181] vdd gnd cell_6t
Xbit_r182_c64 bl[64] br[64] wl[182] vdd gnd cell_6t
Xbit_r183_c64 bl[64] br[64] wl[183] vdd gnd cell_6t
Xbit_r184_c64 bl[64] br[64] wl[184] vdd gnd cell_6t
Xbit_r185_c64 bl[64] br[64] wl[185] vdd gnd cell_6t
Xbit_r186_c64 bl[64] br[64] wl[186] vdd gnd cell_6t
Xbit_r187_c64 bl[64] br[64] wl[187] vdd gnd cell_6t
Xbit_r188_c64 bl[64] br[64] wl[188] vdd gnd cell_6t
Xbit_r189_c64 bl[64] br[64] wl[189] vdd gnd cell_6t
Xbit_r190_c64 bl[64] br[64] wl[190] vdd gnd cell_6t
Xbit_r191_c64 bl[64] br[64] wl[191] vdd gnd cell_6t
Xbit_r192_c64 bl[64] br[64] wl[192] vdd gnd cell_6t
Xbit_r193_c64 bl[64] br[64] wl[193] vdd gnd cell_6t
Xbit_r194_c64 bl[64] br[64] wl[194] vdd gnd cell_6t
Xbit_r195_c64 bl[64] br[64] wl[195] vdd gnd cell_6t
Xbit_r196_c64 bl[64] br[64] wl[196] vdd gnd cell_6t
Xbit_r197_c64 bl[64] br[64] wl[197] vdd gnd cell_6t
Xbit_r198_c64 bl[64] br[64] wl[198] vdd gnd cell_6t
Xbit_r199_c64 bl[64] br[64] wl[199] vdd gnd cell_6t
Xbit_r200_c64 bl[64] br[64] wl[200] vdd gnd cell_6t
Xbit_r201_c64 bl[64] br[64] wl[201] vdd gnd cell_6t
Xbit_r202_c64 bl[64] br[64] wl[202] vdd gnd cell_6t
Xbit_r203_c64 bl[64] br[64] wl[203] vdd gnd cell_6t
Xbit_r204_c64 bl[64] br[64] wl[204] vdd gnd cell_6t
Xbit_r205_c64 bl[64] br[64] wl[205] vdd gnd cell_6t
Xbit_r206_c64 bl[64] br[64] wl[206] vdd gnd cell_6t
Xbit_r207_c64 bl[64] br[64] wl[207] vdd gnd cell_6t
Xbit_r208_c64 bl[64] br[64] wl[208] vdd gnd cell_6t
Xbit_r209_c64 bl[64] br[64] wl[209] vdd gnd cell_6t
Xbit_r210_c64 bl[64] br[64] wl[210] vdd gnd cell_6t
Xbit_r211_c64 bl[64] br[64] wl[211] vdd gnd cell_6t
Xbit_r212_c64 bl[64] br[64] wl[212] vdd gnd cell_6t
Xbit_r213_c64 bl[64] br[64] wl[213] vdd gnd cell_6t
Xbit_r214_c64 bl[64] br[64] wl[214] vdd gnd cell_6t
Xbit_r215_c64 bl[64] br[64] wl[215] vdd gnd cell_6t
Xbit_r216_c64 bl[64] br[64] wl[216] vdd gnd cell_6t
Xbit_r217_c64 bl[64] br[64] wl[217] vdd gnd cell_6t
Xbit_r218_c64 bl[64] br[64] wl[218] vdd gnd cell_6t
Xbit_r219_c64 bl[64] br[64] wl[219] vdd gnd cell_6t
Xbit_r220_c64 bl[64] br[64] wl[220] vdd gnd cell_6t
Xbit_r221_c64 bl[64] br[64] wl[221] vdd gnd cell_6t
Xbit_r222_c64 bl[64] br[64] wl[222] vdd gnd cell_6t
Xbit_r223_c64 bl[64] br[64] wl[223] vdd gnd cell_6t
Xbit_r224_c64 bl[64] br[64] wl[224] vdd gnd cell_6t
Xbit_r225_c64 bl[64] br[64] wl[225] vdd gnd cell_6t
Xbit_r226_c64 bl[64] br[64] wl[226] vdd gnd cell_6t
Xbit_r227_c64 bl[64] br[64] wl[227] vdd gnd cell_6t
Xbit_r228_c64 bl[64] br[64] wl[228] vdd gnd cell_6t
Xbit_r229_c64 bl[64] br[64] wl[229] vdd gnd cell_6t
Xbit_r230_c64 bl[64] br[64] wl[230] vdd gnd cell_6t
Xbit_r231_c64 bl[64] br[64] wl[231] vdd gnd cell_6t
Xbit_r232_c64 bl[64] br[64] wl[232] vdd gnd cell_6t
Xbit_r233_c64 bl[64] br[64] wl[233] vdd gnd cell_6t
Xbit_r234_c64 bl[64] br[64] wl[234] vdd gnd cell_6t
Xbit_r235_c64 bl[64] br[64] wl[235] vdd gnd cell_6t
Xbit_r236_c64 bl[64] br[64] wl[236] vdd gnd cell_6t
Xbit_r237_c64 bl[64] br[64] wl[237] vdd gnd cell_6t
Xbit_r238_c64 bl[64] br[64] wl[238] vdd gnd cell_6t
Xbit_r239_c64 bl[64] br[64] wl[239] vdd gnd cell_6t
Xbit_r240_c64 bl[64] br[64] wl[240] vdd gnd cell_6t
Xbit_r241_c64 bl[64] br[64] wl[241] vdd gnd cell_6t
Xbit_r242_c64 bl[64] br[64] wl[242] vdd gnd cell_6t
Xbit_r243_c64 bl[64] br[64] wl[243] vdd gnd cell_6t
Xbit_r244_c64 bl[64] br[64] wl[244] vdd gnd cell_6t
Xbit_r245_c64 bl[64] br[64] wl[245] vdd gnd cell_6t
Xbit_r246_c64 bl[64] br[64] wl[246] vdd gnd cell_6t
Xbit_r247_c64 bl[64] br[64] wl[247] vdd gnd cell_6t
Xbit_r248_c64 bl[64] br[64] wl[248] vdd gnd cell_6t
Xbit_r249_c64 bl[64] br[64] wl[249] vdd gnd cell_6t
Xbit_r250_c64 bl[64] br[64] wl[250] vdd gnd cell_6t
Xbit_r251_c64 bl[64] br[64] wl[251] vdd gnd cell_6t
Xbit_r252_c64 bl[64] br[64] wl[252] vdd gnd cell_6t
Xbit_r253_c64 bl[64] br[64] wl[253] vdd gnd cell_6t
Xbit_r254_c64 bl[64] br[64] wl[254] vdd gnd cell_6t
Xbit_r255_c64 bl[64] br[64] wl[255] vdd gnd cell_6t
Xbit_r256_c64 bl[64] br[64] wl[256] vdd gnd cell_6t
Xbit_r257_c64 bl[64] br[64] wl[257] vdd gnd cell_6t
Xbit_r258_c64 bl[64] br[64] wl[258] vdd gnd cell_6t
Xbit_r259_c64 bl[64] br[64] wl[259] vdd gnd cell_6t
Xbit_r260_c64 bl[64] br[64] wl[260] vdd gnd cell_6t
Xbit_r261_c64 bl[64] br[64] wl[261] vdd gnd cell_6t
Xbit_r262_c64 bl[64] br[64] wl[262] vdd gnd cell_6t
Xbit_r263_c64 bl[64] br[64] wl[263] vdd gnd cell_6t
Xbit_r264_c64 bl[64] br[64] wl[264] vdd gnd cell_6t
Xbit_r265_c64 bl[64] br[64] wl[265] vdd gnd cell_6t
Xbit_r266_c64 bl[64] br[64] wl[266] vdd gnd cell_6t
Xbit_r267_c64 bl[64] br[64] wl[267] vdd gnd cell_6t
Xbit_r268_c64 bl[64] br[64] wl[268] vdd gnd cell_6t
Xbit_r269_c64 bl[64] br[64] wl[269] vdd gnd cell_6t
Xbit_r270_c64 bl[64] br[64] wl[270] vdd gnd cell_6t
Xbit_r271_c64 bl[64] br[64] wl[271] vdd gnd cell_6t
Xbit_r272_c64 bl[64] br[64] wl[272] vdd gnd cell_6t
Xbit_r273_c64 bl[64] br[64] wl[273] vdd gnd cell_6t
Xbit_r274_c64 bl[64] br[64] wl[274] vdd gnd cell_6t
Xbit_r275_c64 bl[64] br[64] wl[275] vdd gnd cell_6t
Xbit_r276_c64 bl[64] br[64] wl[276] vdd gnd cell_6t
Xbit_r277_c64 bl[64] br[64] wl[277] vdd gnd cell_6t
Xbit_r278_c64 bl[64] br[64] wl[278] vdd gnd cell_6t
Xbit_r279_c64 bl[64] br[64] wl[279] vdd gnd cell_6t
Xbit_r280_c64 bl[64] br[64] wl[280] vdd gnd cell_6t
Xbit_r281_c64 bl[64] br[64] wl[281] vdd gnd cell_6t
Xbit_r282_c64 bl[64] br[64] wl[282] vdd gnd cell_6t
Xbit_r283_c64 bl[64] br[64] wl[283] vdd gnd cell_6t
Xbit_r284_c64 bl[64] br[64] wl[284] vdd gnd cell_6t
Xbit_r285_c64 bl[64] br[64] wl[285] vdd gnd cell_6t
Xbit_r286_c64 bl[64] br[64] wl[286] vdd gnd cell_6t
Xbit_r287_c64 bl[64] br[64] wl[287] vdd gnd cell_6t
Xbit_r288_c64 bl[64] br[64] wl[288] vdd gnd cell_6t
Xbit_r289_c64 bl[64] br[64] wl[289] vdd gnd cell_6t
Xbit_r290_c64 bl[64] br[64] wl[290] vdd gnd cell_6t
Xbit_r291_c64 bl[64] br[64] wl[291] vdd gnd cell_6t
Xbit_r292_c64 bl[64] br[64] wl[292] vdd gnd cell_6t
Xbit_r293_c64 bl[64] br[64] wl[293] vdd gnd cell_6t
Xbit_r294_c64 bl[64] br[64] wl[294] vdd gnd cell_6t
Xbit_r295_c64 bl[64] br[64] wl[295] vdd gnd cell_6t
Xbit_r296_c64 bl[64] br[64] wl[296] vdd gnd cell_6t
Xbit_r297_c64 bl[64] br[64] wl[297] vdd gnd cell_6t
Xbit_r298_c64 bl[64] br[64] wl[298] vdd gnd cell_6t
Xbit_r299_c64 bl[64] br[64] wl[299] vdd gnd cell_6t
Xbit_r300_c64 bl[64] br[64] wl[300] vdd gnd cell_6t
Xbit_r301_c64 bl[64] br[64] wl[301] vdd gnd cell_6t
Xbit_r302_c64 bl[64] br[64] wl[302] vdd gnd cell_6t
Xbit_r303_c64 bl[64] br[64] wl[303] vdd gnd cell_6t
Xbit_r304_c64 bl[64] br[64] wl[304] vdd gnd cell_6t
Xbit_r305_c64 bl[64] br[64] wl[305] vdd gnd cell_6t
Xbit_r306_c64 bl[64] br[64] wl[306] vdd gnd cell_6t
Xbit_r307_c64 bl[64] br[64] wl[307] vdd gnd cell_6t
Xbit_r308_c64 bl[64] br[64] wl[308] vdd gnd cell_6t
Xbit_r309_c64 bl[64] br[64] wl[309] vdd gnd cell_6t
Xbit_r310_c64 bl[64] br[64] wl[310] vdd gnd cell_6t
Xbit_r311_c64 bl[64] br[64] wl[311] vdd gnd cell_6t
Xbit_r312_c64 bl[64] br[64] wl[312] vdd gnd cell_6t
Xbit_r313_c64 bl[64] br[64] wl[313] vdd gnd cell_6t
Xbit_r314_c64 bl[64] br[64] wl[314] vdd gnd cell_6t
Xbit_r315_c64 bl[64] br[64] wl[315] vdd gnd cell_6t
Xbit_r316_c64 bl[64] br[64] wl[316] vdd gnd cell_6t
Xbit_r317_c64 bl[64] br[64] wl[317] vdd gnd cell_6t
Xbit_r318_c64 bl[64] br[64] wl[318] vdd gnd cell_6t
Xbit_r319_c64 bl[64] br[64] wl[319] vdd gnd cell_6t
Xbit_r320_c64 bl[64] br[64] wl[320] vdd gnd cell_6t
Xbit_r321_c64 bl[64] br[64] wl[321] vdd gnd cell_6t
Xbit_r322_c64 bl[64] br[64] wl[322] vdd gnd cell_6t
Xbit_r323_c64 bl[64] br[64] wl[323] vdd gnd cell_6t
Xbit_r324_c64 bl[64] br[64] wl[324] vdd gnd cell_6t
Xbit_r325_c64 bl[64] br[64] wl[325] vdd gnd cell_6t
Xbit_r326_c64 bl[64] br[64] wl[326] vdd gnd cell_6t
Xbit_r327_c64 bl[64] br[64] wl[327] vdd gnd cell_6t
Xbit_r328_c64 bl[64] br[64] wl[328] vdd gnd cell_6t
Xbit_r329_c64 bl[64] br[64] wl[329] vdd gnd cell_6t
Xbit_r330_c64 bl[64] br[64] wl[330] vdd gnd cell_6t
Xbit_r331_c64 bl[64] br[64] wl[331] vdd gnd cell_6t
Xbit_r332_c64 bl[64] br[64] wl[332] vdd gnd cell_6t
Xbit_r333_c64 bl[64] br[64] wl[333] vdd gnd cell_6t
Xbit_r334_c64 bl[64] br[64] wl[334] vdd gnd cell_6t
Xbit_r335_c64 bl[64] br[64] wl[335] vdd gnd cell_6t
Xbit_r336_c64 bl[64] br[64] wl[336] vdd gnd cell_6t
Xbit_r337_c64 bl[64] br[64] wl[337] vdd gnd cell_6t
Xbit_r338_c64 bl[64] br[64] wl[338] vdd gnd cell_6t
Xbit_r339_c64 bl[64] br[64] wl[339] vdd gnd cell_6t
Xbit_r340_c64 bl[64] br[64] wl[340] vdd gnd cell_6t
Xbit_r341_c64 bl[64] br[64] wl[341] vdd gnd cell_6t
Xbit_r342_c64 bl[64] br[64] wl[342] vdd gnd cell_6t
Xbit_r343_c64 bl[64] br[64] wl[343] vdd gnd cell_6t
Xbit_r344_c64 bl[64] br[64] wl[344] vdd gnd cell_6t
Xbit_r345_c64 bl[64] br[64] wl[345] vdd gnd cell_6t
Xbit_r346_c64 bl[64] br[64] wl[346] vdd gnd cell_6t
Xbit_r347_c64 bl[64] br[64] wl[347] vdd gnd cell_6t
Xbit_r348_c64 bl[64] br[64] wl[348] vdd gnd cell_6t
Xbit_r349_c64 bl[64] br[64] wl[349] vdd gnd cell_6t
Xbit_r350_c64 bl[64] br[64] wl[350] vdd gnd cell_6t
Xbit_r351_c64 bl[64] br[64] wl[351] vdd gnd cell_6t
Xbit_r352_c64 bl[64] br[64] wl[352] vdd gnd cell_6t
Xbit_r353_c64 bl[64] br[64] wl[353] vdd gnd cell_6t
Xbit_r354_c64 bl[64] br[64] wl[354] vdd gnd cell_6t
Xbit_r355_c64 bl[64] br[64] wl[355] vdd gnd cell_6t
Xbit_r356_c64 bl[64] br[64] wl[356] vdd gnd cell_6t
Xbit_r357_c64 bl[64] br[64] wl[357] vdd gnd cell_6t
Xbit_r358_c64 bl[64] br[64] wl[358] vdd gnd cell_6t
Xbit_r359_c64 bl[64] br[64] wl[359] vdd gnd cell_6t
Xbit_r360_c64 bl[64] br[64] wl[360] vdd gnd cell_6t
Xbit_r361_c64 bl[64] br[64] wl[361] vdd gnd cell_6t
Xbit_r362_c64 bl[64] br[64] wl[362] vdd gnd cell_6t
Xbit_r363_c64 bl[64] br[64] wl[363] vdd gnd cell_6t
Xbit_r364_c64 bl[64] br[64] wl[364] vdd gnd cell_6t
Xbit_r365_c64 bl[64] br[64] wl[365] vdd gnd cell_6t
Xbit_r366_c64 bl[64] br[64] wl[366] vdd gnd cell_6t
Xbit_r367_c64 bl[64] br[64] wl[367] vdd gnd cell_6t
Xbit_r368_c64 bl[64] br[64] wl[368] vdd gnd cell_6t
Xbit_r369_c64 bl[64] br[64] wl[369] vdd gnd cell_6t
Xbit_r370_c64 bl[64] br[64] wl[370] vdd gnd cell_6t
Xbit_r371_c64 bl[64] br[64] wl[371] vdd gnd cell_6t
Xbit_r372_c64 bl[64] br[64] wl[372] vdd gnd cell_6t
Xbit_r373_c64 bl[64] br[64] wl[373] vdd gnd cell_6t
Xbit_r374_c64 bl[64] br[64] wl[374] vdd gnd cell_6t
Xbit_r375_c64 bl[64] br[64] wl[375] vdd gnd cell_6t
Xbit_r376_c64 bl[64] br[64] wl[376] vdd gnd cell_6t
Xbit_r377_c64 bl[64] br[64] wl[377] vdd gnd cell_6t
Xbit_r378_c64 bl[64] br[64] wl[378] vdd gnd cell_6t
Xbit_r379_c64 bl[64] br[64] wl[379] vdd gnd cell_6t
Xbit_r380_c64 bl[64] br[64] wl[380] vdd gnd cell_6t
Xbit_r381_c64 bl[64] br[64] wl[381] vdd gnd cell_6t
Xbit_r382_c64 bl[64] br[64] wl[382] vdd gnd cell_6t
Xbit_r383_c64 bl[64] br[64] wl[383] vdd gnd cell_6t
Xbit_r384_c64 bl[64] br[64] wl[384] vdd gnd cell_6t
Xbit_r385_c64 bl[64] br[64] wl[385] vdd gnd cell_6t
Xbit_r386_c64 bl[64] br[64] wl[386] vdd gnd cell_6t
Xbit_r387_c64 bl[64] br[64] wl[387] vdd gnd cell_6t
Xbit_r388_c64 bl[64] br[64] wl[388] vdd gnd cell_6t
Xbit_r389_c64 bl[64] br[64] wl[389] vdd gnd cell_6t
Xbit_r390_c64 bl[64] br[64] wl[390] vdd gnd cell_6t
Xbit_r391_c64 bl[64] br[64] wl[391] vdd gnd cell_6t
Xbit_r392_c64 bl[64] br[64] wl[392] vdd gnd cell_6t
Xbit_r393_c64 bl[64] br[64] wl[393] vdd gnd cell_6t
Xbit_r394_c64 bl[64] br[64] wl[394] vdd gnd cell_6t
Xbit_r395_c64 bl[64] br[64] wl[395] vdd gnd cell_6t
Xbit_r396_c64 bl[64] br[64] wl[396] vdd gnd cell_6t
Xbit_r397_c64 bl[64] br[64] wl[397] vdd gnd cell_6t
Xbit_r398_c64 bl[64] br[64] wl[398] vdd gnd cell_6t
Xbit_r399_c64 bl[64] br[64] wl[399] vdd gnd cell_6t
Xbit_r400_c64 bl[64] br[64] wl[400] vdd gnd cell_6t
Xbit_r401_c64 bl[64] br[64] wl[401] vdd gnd cell_6t
Xbit_r402_c64 bl[64] br[64] wl[402] vdd gnd cell_6t
Xbit_r403_c64 bl[64] br[64] wl[403] vdd gnd cell_6t
Xbit_r404_c64 bl[64] br[64] wl[404] vdd gnd cell_6t
Xbit_r405_c64 bl[64] br[64] wl[405] vdd gnd cell_6t
Xbit_r406_c64 bl[64] br[64] wl[406] vdd gnd cell_6t
Xbit_r407_c64 bl[64] br[64] wl[407] vdd gnd cell_6t
Xbit_r408_c64 bl[64] br[64] wl[408] vdd gnd cell_6t
Xbit_r409_c64 bl[64] br[64] wl[409] vdd gnd cell_6t
Xbit_r410_c64 bl[64] br[64] wl[410] vdd gnd cell_6t
Xbit_r411_c64 bl[64] br[64] wl[411] vdd gnd cell_6t
Xbit_r412_c64 bl[64] br[64] wl[412] vdd gnd cell_6t
Xbit_r413_c64 bl[64] br[64] wl[413] vdd gnd cell_6t
Xbit_r414_c64 bl[64] br[64] wl[414] vdd gnd cell_6t
Xbit_r415_c64 bl[64] br[64] wl[415] vdd gnd cell_6t
Xbit_r416_c64 bl[64] br[64] wl[416] vdd gnd cell_6t
Xbit_r417_c64 bl[64] br[64] wl[417] vdd gnd cell_6t
Xbit_r418_c64 bl[64] br[64] wl[418] vdd gnd cell_6t
Xbit_r419_c64 bl[64] br[64] wl[419] vdd gnd cell_6t
Xbit_r420_c64 bl[64] br[64] wl[420] vdd gnd cell_6t
Xbit_r421_c64 bl[64] br[64] wl[421] vdd gnd cell_6t
Xbit_r422_c64 bl[64] br[64] wl[422] vdd gnd cell_6t
Xbit_r423_c64 bl[64] br[64] wl[423] vdd gnd cell_6t
Xbit_r424_c64 bl[64] br[64] wl[424] vdd gnd cell_6t
Xbit_r425_c64 bl[64] br[64] wl[425] vdd gnd cell_6t
Xbit_r426_c64 bl[64] br[64] wl[426] vdd gnd cell_6t
Xbit_r427_c64 bl[64] br[64] wl[427] vdd gnd cell_6t
Xbit_r428_c64 bl[64] br[64] wl[428] vdd gnd cell_6t
Xbit_r429_c64 bl[64] br[64] wl[429] vdd gnd cell_6t
Xbit_r430_c64 bl[64] br[64] wl[430] vdd gnd cell_6t
Xbit_r431_c64 bl[64] br[64] wl[431] vdd gnd cell_6t
Xbit_r432_c64 bl[64] br[64] wl[432] vdd gnd cell_6t
Xbit_r433_c64 bl[64] br[64] wl[433] vdd gnd cell_6t
Xbit_r434_c64 bl[64] br[64] wl[434] vdd gnd cell_6t
Xbit_r435_c64 bl[64] br[64] wl[435] vdd gnd cell_6t
Xbit_r436_c64 bl[64] br[64] wl[436] vdd gnd cell_6t
Xbit_r437_c64 bl[64] br[64] wl[437] vdd gnd cell_6t
Xbit_r438_c64 bl[64] br[64] wl[438] vdd gnd cell_6t
Xbit_r439_c64 bl[64] br[64] wl[439] vdd gnd cell_6t
Xbit_r440_c64 bl[64] br[64] wl[440] vdd gnd cell_6t
Xbit_r441_c64 bl[64] br[64] wl[441] vdd gnd cell_6t
Xbit_r442_c64 bl[64] br[64] wl[442] vdd gnd cell_6t
Xbit_r443_c64 bl[64] br[64] wl[443] vdd gnd cell_6t
Xbit_r444_c64 bl[64] br[64] wl[444] vdd gnd cell_6t
Xbit_r445_c64 bl[64] br[64] wl[445] vdd gnd cell_6t
Xbit_r446_c64 bl[64] br[64] wl[446] vdd gnd cell_6t
Xbit_r447_c64 bl[64] br[64] wl[447] vdd gnd cell_6t
Xbit_r448_c64 bl[64] br[64] wl[448] vdd gnd cell_6t
Xbit_r449_c64 bl[64] br[64] wl[449] vdd gnd cell_6t
Xbit_r450_c64 bl[64] br[64] wl[450] vdd gnd cell_6t
Xbit_r451_c64 bl[64] br[64] wl[451] vdd gnd cell_6t
Xbit_r452_c64 bl[64] br[64] wl[452] vdd gnd cell_6t
Xbit_r453_c64 bl[64] br[64] wl[453] vdd gnd cell_6t
Xbit_r454_c64 bl[64] br[64] wl[454] vdd gnd cell_6t
Xbit_r455_c64 bl[64] br[64] wl[455] vdd gnd cell_6t
Xbit_r456_c64 bl[64] br[64] wl[456] vdd gnd cell_6t
Xbit_r457_c64 bl[64] br[64] wl[457] vdd gnd cell_6t
Xbit_r458_c64 bl[64] br[64] wl[458] vdd gnd cell_6t
Xbit_r459_c64 bl[64] br[64] wl[459] vdd gnd cell_6t
Xbit_r460_c64 bl[64] br[64] wl[460] vdd gnd cell_6t
Xbit_r461_c64 bl[64] br[64] wl[461] vdd gnd cell_6t
Xbit_r462_c64 bl[64] br[64] wl[462] vdd gnd cell_6t
Xbit_r463_c64 bl[64] br[64] wl[463] vdd gnd cell_6t
Xbit_r464_c64 bl[64] br[64] wl[464] vdd gnd cell_6t
Xbit_r465_c64 bl[64] br[64] wl[465] vdd gnd cell_6t
Xbit_r466_c64 bl[64] br[64] wl[466] vdd gnd cell_6t
Xbit_r467_c64 bl[64] br[64] wl[467] vdd gnd cell_6t
Xbit_r468_c64 bl[64] br[64] wl[468] vdd gnd cell_6t
Xbit_r469_c64 bl[64] br[64] wl[469] vdd gnd cell_6t
Xbit_r470_c64 bl[64] br[64] wl[470] vdd gnd cell_6t
Xbit_r471_c64 bl[64] br[64] wl[471] vdd gnd cell_6t
Xbit_r472_c64 bl[64] br[64] wl[472] vdd gnd cell_6t
Xbit_r473_c64 bl[64] br[64] wl[473] vdd gnd cell_6t
Xbit_r474_c64 bl[64] br[64] wl[474] vdd gnd cell_6t
Xbit_r475_c64 bl[64] br[64] wl[475] vdd gnd cell_6t
Xbit_r476_c64 bl[64] br[64] wl[476] vdd gnd cell_6t
Xbit_r477_c64 bl[64] br[64] wl[477] vdd gnd cell_6t
Xbit_r478_c64 bl[64] br[64] wl[478] vdd gnd cell_6t
Xbit_r479_c64 bl[64] br[64] wl[479] vdd gnd cell_6t
Xbit_r480_c64 bl[64] br[64] wl[480] vdd gnd cell_6t
Xbit_r481_c64 bl[64] br[64] wl[481] vdd gnd cell_6t
Xbit_r482_c64 bl[64] br[64] wl[482] vdd gnd cell_6t
Xbit_r483_c64 bl[64] br[64] wl[483] vdd gnd cell_6t
Xbit_r484_c64 bl[64] br[64] wl[484] vdd gnd cell_6t
Xbit_r485_c64 bl[64] br[64] wl[485] vdd gnd cell_6t
Xbit_r486_c64 bl[64] br[64] wl[486] vdd gnd cell_6t
Xbit_r487_c64 bl[64] br[64] wl[487] vdd gnd cell_6t
Xbit_r488_c64 bl[64] br[64] wl[488] vdd gnd cell_6t
Xbit_r489_c64 bl[64] br[64] wl[489] vdd gnd cell_6t
Xbit_r490_c64 bl[64] br[64] wl[490] vdd gnd cell_6t
Xbit_r491_c64 bl[64] br[64] wl[491] vdd gnd cell_6t
Xbit_r492_c64 bl[64] br[64] wl[492] vdd gnd cell_6t
Xbit_r493_c64 bl[64] br[64] wl[493] vdd gnd cell_6t
Xbit_r494_c64 bl[64] br[64] wl[494] vdd gnd cell_6t
Xbit_r495_c64 bl[64] br[64] wl[495] vdd gnd cell_6t
Xbit_r496_c64 bl[64] br[64] wl[496] vdd gnd cell_6t
Xbit_r497_c64 bl[64] br[64] wl[497] vdd gnd cell_6t
Xbit_r498_c64 bl[64] br[64] wl[498] vdd gnd cell_6t
Xbit_r499_c64 bl[64] br[64] wl[499] vdd gnd cell_6t
Xbit_r500_c64 bl[64] br[64] wl[500] vdd gnd cell_6t
Xbit_r501_c64 bl[64] br[64] wl[501] vdd gnd cell_6t
Xbit_r502_c64 bl[64] br[64] wl[502] vdd gnd cell_6t
Xbit_r503_c64 bl[64] br[64] wl[503] vdd gnd cell_6t
Xbit_r504_c64 bl[64] br[64] wl[504] vdd gnd cell_6t
Xbit_r505_c64 bl[64] br[64] wl[505] vdd gnd cell_6t
Xbit_r506_c64 bl[64] br[64] wl[506] vdd gnd cell_6t
Xbit_r507_c64 bl[64] br[64] wl[507] vdd gnd cell_6t
Xbit_r508_c64 bl[64] br[64] wl[508] vdd gnd cell_6t
Xbit_r509_c64 bl[64] br[64] wl[509] vdd gnd cell_6t
Xbit_r510_c64 bl[64] br[64] wl[510] vdd gnd cell_6t
Xbit_r511_c64 bl[64] br[64] wl[511] vdd gnd cell_6t
Xbit_r0_c65 bl[65] br[65] wl[0] vdd gnd cell_6t
Xbit_r1_c65 bl[65] br[65] wl[1] vdd gnd cell_6t
Xbit_r2_c65 bl[65] br[65] wl[2] vdd gnd cell_6t
Xbit_r3_c65 bl[65] br[65] wl[3] vdd gnd cell_6t
Xbit_r4_c65 bl[65] br[65] wl[4] vdd gnd cell_6t
Xbit_r5_c65 bl[65] br[65] wl[5] vdd gnd cell_6t
Xbit_r6_c65 bl[65] br[65] wl[6] vdd gnd cell_6t
Xbit_r7_c65 bl[65] br[65] wl[7] vdd gnd cell_6t
Xbit_r8_c65 bl[65] br[65] wl[8] vdd gnd cell_6t
Xbit_r9_c65 bl[65] br[65] wl[9] vdd gnd cell_6t
Xbit_r10_c65 bl[65] br[65] wl[10] vdd gnd cell_6t
Xbit_r11_c65 bl[65] br[65] wl[11] vdd gnd cell_6t
Xbit_r12_c65 bl[65] br[65] wl[12] vdd gnd cell_6t
Xbit_r13_c65 bl[65] br[65] wl[13] vdd gnd cell_6t
Xbit_r14_c65 bl[65] br[65] wl[14] vdd gnd cell_6t
Xbit_r15_c65 bl[65] br[65] wl[15] vdd gnd cell_6t
Xbit_r16_c65 bl[65] br[65] wl[16] vdd gnd cell_6t
Xbit_r17_c65 bl[65] br[65] wl[17] vdd gnd cell_6t
Xbit_r18_c65 bl[65] br[65] wl[18] vdd gnd cell_6t
Xbit_r19_c65 bl[65] br[65] wl[19] vdd gnd cell_6t
Xbit_r20_c65 bl[65] br[65] wl[20] vdd gnd cell_6t
Xbit_r21_c65 bl[65] br[65] wl[21] vdd gnd cell_6t
Xbit_r22_c65 bl[65] br[65] wl[22] vdd gnd cell_6t
Xbit_r23_c65 bl[65] br[65] wl[23] vdd gnd cell_6t
Xbit_r24_c65 bl[65] br[65] wl[24] vdd gnd cell_6t
Xbit_r25_c65 bl[65] br[65] wl[25] vdd gnd cell_6t
Xbit_r26_c65 bl[65] br[65] wl[26] vdd gnd cell_6t
Xbit_r27_c65 bl[65] br[65] wl[27] vdd gnd cell_6t
Xbit_r28_c65 bl[65] br[65] wl[28] vdd gnd cell_6t
Xbit_r29_c65 bl[65] br[65] wl[29] vdd gnd cell_6t
Xbit_r30_c65 bl[65] br[65] wl[30] vdd gnd cell_6t
Xbit_r31_c65 bl[65] br[65] wl[31] vdd gnd cell_6t
Xbit_r32_c65 bl[65] br[65] wl[32] vdd gnd cell_6t
Xbit_r33_c65 bl[65] br[65] wl[33] vdd gnd cell_6t
Xbit_r34_c65 bl[65] br[65] wl[34] vdd gnd cell_6t
Xbit_r35_c65 bl[65] br[65] wl[35] vdd gnd cell_6t
Xbit_r36_c65 bl[65] br[65] wl[36] vdd gnd cell_6t
Xbit_r37_c65 bl[65] br[65] wl[37] vdd gnd cell_6t
Xbit_r38_c65 bl[65] br[65] wl[38] vdd gnd cell_6t
Xbit_r39_c65 bl[65] br[65] wl[39] vdd gnd cell_6t
Xbit_r40_c65 bl[65] br[65] wl[40] vdd gnd cell_6t
Xbit_r41_c65 bl[65] br[65] wl[41] vdd gnd cell_6t
Xbit_r42_c65 bl[65] br[65] wl[42] vdd gnd cell_6t
Xbit_r43_c65 bl[65] br[65] wl[43] vdd gnd cell_6t
Xbit_r44_c65 bl[65] br[65] wl[44] vdd gnd cell_6t
Xbit_r45_c65 bl[65] br[65] wl[45] vdd gnd cell_6t
Xbit_r46_c65 bl[65] br[65] wl[46] vdd gnd cell_6t
Xbit_r47_c65 bl[65] br[65] wl[47] vdd gnd cell_6t
Xbit_r48_c65 bl[65] br[65] wl[48] vdd gnd cell_6t
Xbit_r49_c65 bl[65] br[65] wl[49] vdd gnd cell_6t
Xbit_r50_c65 bl[65] br[65] wl[50] vdd gnd cell_6t
Xbit_r51_c65 bl[65] br[65] wl[51] vdd gnd cell_6t
Xbit_r52_c65 bl[65] br[65] wl[52] vdd gnd cell_6t
Xbit_r53_c65 bl[65] br[65] wl[53] vdd gnd cell_6t
Xbit_r54_c65 bl[65] br[65] wl[54] vdd gnd cell_6t
Xbit_r55_c65 bl[65] br[65] wl[55] vdd gnd cell_6t
Xbit_r56_c65 bl[65] br[65] wl[56] vdd gnd cell_6t
Xbit_r57_c65 bl[65] br[65] wl[57] vdd gnd cell_6t
Xbit_r58_c65 bl[65] br[65] wl[58] vdd gnd cell_6t
Xbit_r59_c65 bl[65] br[65] wl[59] vdd gnd cell_6t
Xbit_r60_c65 bl[65] br[65] wl[60] vdd gnd cell_6t
Xbit_r61_c65 bl[65] br[65] wl[61] vdd gnd cell_6t
Xbit_r62_c65 bl[65] br[65] wl[62] vdd gnd cell_6t
Xbit_r63_c65 bl[65] br[65] wl[63] vdd gnd cell_6t
Xbit_r64_c65 bl[65] br[65] wl[64] vdd gnd cell_6t
Xbit_r65_c65 bl[65] br[65] wl[65] vdd gnd cell_6t
Xbit_r66_c65 bl[65] br[65] wl[66] vdd gnd cell_6t
Xbit_r67_c65 bl[65] br[65] wl[67] vdd gnd cell_6t
Xbit_r68_c65 bl[65] br[65] wl[68] vdd gnd cell_6t
Xbit_r69_c65 bl[65] br[65] wl[69] vdd gnd cell_6t
Xbit_r70_c65 bl[65] br[65] wl[70] vdd gnd cell_6t
Xbit_r71_c65 bl[65] br[65] wl[71] vdd gnd cell_6t
Xbit_r72_c65 bl[65] br[65] wl[72] vdd gnd cell_6t
Xbit_r73_c65 bl[65] br[65] wl[73] vdd gnd cell_6t
Xbit_r74_c65 bl[65] br[65] wl[74] vdd gnd cell_6t
Xbit_r75_c65 bl[65] br[65] wl[75] vdd gnd cell_6t
Xbit_r76_c65 bl[65] br[65] wl[76] vdd gnd cell_6t
Xbit_r77_c65 bl[65] br[65] wl[77] vdd gnd cell_6t
Xbit_r78_c65 bl[65] br[65] wl[78] vdd gnd cell_6t
Xbit_r79_c65 bl[65] br[65] wl[79] vdd gnd cell_6t
Xbit_r80_c65 bl[65] br[65] wl[80] vdd gnd cell_6t
Xbit_r81_c65 bl[65] br[65] wl[81] vdd gnd cell_6t
Xbit_r82_c65 bl[65] br[65] wl[82] vdd gnd cell_6t
Xbit_r83_c65 bl[65] br[65] wl[83] vdd gnd cell_6t
Xbit_r84_c65 bl[65] br[65] wl[84] vdd gnd cell_6t
Xbit_r85_c65 bl[65] br[65] wl[85] vdd gnd cell_6t
Xbit_r86_c65 bl[65] br[65] wl[86] vdd gnd cell_6t
Xbit_r87_c65 bl[65] br[65] wl[87] vdd gnd cell_6t
Xbit_r88_c65 bl[65] br[65] wl[88] vdd gnd cell_6t
Xbit_r89_c65 bl[65] br[65] wl[89] vdd gnd cell_6t
Xbit_r90_c65 bl[65] br[65] wl[90] vdd gnd cell_6t
Xbit_r91_c65 bl[65] br[65] wl[91] vdd gnd cell_6t
Xbit_r92_c65 bl[65] br[65] wl[92] vdd gnd cell_6t
Xbit_r93_c65 bl[65] br[65] wl[93] vdd gnd cell_6t
Xbit_r94_c65 bl[65] br[65] wl[94] vdd gnd cell_6t
Xbit_r95_c65 bl[65] br[65] wl[95] vdd gnd cell_6t
Xbit_r96_c65 bl[65] br[65] wl[96] vdd gnd cell_6t
Xbit_r97_c65 bl[65] br[65] wl[97] vdd gnd cell_6t
Xbit_r98_c65 bl[65] br[65] wl[98] vdd gnd cell_6t
Xbit_r99_c65 bl[65] br[65] wl[99] vdd gnd cell_6t
Xbit_r100_c65 bl[65] br[65] wl[100] vdd gnd cell_6t
Xbit_r101_c65 bl[65] br[65] wl[101] vdd gnd cell_6t
Xbit_r102_c65 bl[65] br[65] wl[102] vdd gnd cell_6t
Xbit_r103_c65 bl[65] br[65] wl[103] vdd gnd cell_6t
Xbit_r104_c65 bl[65] br[65] wl[104] vdd gnd cell_6t
Xbit_r105_c65 bl[65] br[65] wl[105] vdd gnd cell_6t
Xbit_r106_c65 bl[65] br[65] wl[106] vdd gnd cell_6t
Xbit_r107_c65 bl[65] br[65] wl[107] vdd gnd cell_6t
Xbit_r108_c65 bl[65] br[65] wl[108] vdd gnd cell_6t
Xbit_r109_c65 bl[65] br[65] wl[109] vdd gnd cell_6t
Xbit_r110_c65 bl[65] br[65] wl[110] vdd gnd cell_6t
Xbit_r111_c65 bl[65] br[65] wl[111] vdd gnd cell_6t
Xbit_r112_c65 bl[65] br[65] wl[112] vdd gnd cell_6t
Xbit_r113_c65 bl[65] br[65] wl[113] vdd gnd cell_6t
Xbit_r114_c65 bl[65] br[65] wl[114] vdd gnd cell_6t
Xbit_r115_c65 bl[65] br[65] wl[115] vdd gnd cell_6t
Xbit_r116_c65 bl[65] br[65] wl[116] vdd gnd cell_6t
Xbit_r117_c65 bl[65] br[65] wl[117] vdd gnd cell_6t
Xbit_r118_c65 bl[65] br[65] wl[118] vdd gnd cell_6t
Xbit_r119_c65 bl[65] br[65] wl[119] vdd gnd cell_6t
Xbit_r120_c65 bl[65] br[65] wl[120] vdd gnd cell_6t
Xbit_r121_c65 bl[65] br[65] wl[121] vdd gnd cell_6t
Xbit_r122_c65 bl[65] br[65] wl[122] vdd gnd cell_6t
Xbit_r123_c65 bl[65] br[65] wl[123] vdd gnd cell_6t
Xbit_r124_c65 bl[65] br[65] wl[124] vdd gnd cell_6t
Xbit_r125_c65 bl[65] br[65] wl[125] vdd gnd cell_6t
Xbit_r126_c65 bl[65] br[65] wl[126] vdd gnd cell_6t
Xbit_r127_c65 bl[65] br[65] wl[127] vdd gnd cell_6t
Xbit_r128_c65 bl[65] br[65] wl[128] vdd gnd cell_6t
Xbit_r129_c65 bl[65] br[65] wl[129] vdd gnd cell_6t
Xbit_r130_c65 bl[65] br[65] wl[130] vdd gnd cell_6t
Xbit_r131_c65 bl[65] br[65] wl[131] vdd gnd cell_6t
Xbit_r132_c65 bl[65] br[65] wl[132] vdd gnd cell_6t
Xbit_r133_c65 bl[65] br[65] wl[133] vdd gnd cell_6t
Xbit_r134_c65 bl[65] br[65] wl[134] vdd gnd cell_6t
Xbit_r135_c65 bl[65] br[65] wl[135] vdd gnd cell_6t
Xbit_r136_c65 bl[65] br[65] wl[136] vdd gnd cell_6t
Xbit_r137_c65 bl[65] br[65] wl[137] vdd gnd cell_6t
Xbit_r138_c65 bl[65] br[65] wl[138] vdd gnd cell_6t
Xbit_r139_c65 bl[65] br[65] wl[139] vdd gnd cell_6t
Xbit_r140_c65 bl[65] br[65] wl[140] vdd gnd cell_6t
Xbit_r141_c65 bl[65] br[65] wl[141] vdd gnd cell_6t
Xbit_r142_c65 bl[65] br[65] wl[142] vdd gnd cell_6t
Xbit_r143_c65 bl[65] br[65] wl[143] vdd gnd cell_6t
Xbit_r144_c65 bl[65] br[65] wl[144] vdd gnd cell_6t
Xbit_r145_c65 bl[65] br[65] wl[145] vdd gnd cell_6t
Xbit_r146_c65 bl[65] br[65] wl[146] vdd gnd cell_6t
Xbit_r147_c65 bl[65] br[65] wl[147] vdd gnd cell_6t
Xbit_r148_c65 bl[65] br[65] wl[148] vdd gnd cell_6t
Xbit_r149_c65 bl[65] br[65] wl[149] vdd gnd cell_6t
Xbit_r150_c65 bl[65] br[65] wl[150] vdd gnd cell_6t
Xbit_r151_c65 bl[65] br[65] wl[151] vdd gnd cell_6t
Xbit_r152_c65 bl[65] br[65] wl[152] vdd gnd cell_6t
Xbit_r153_c65 bl[65] br[65] wl[153] vdd gnd cell_6t
Xbit_r154_c65 bl[65] br[65] wl[154] vdd gnd cell_6t
Xbit_r155_c65 bl[65] br[65] wl[155] vdd gnd cell_6t
Xbit_r156_c65 bl[65] br[65] wl[156] vdd gnd cell_6t
Xbit_r157_c65 bl[65] br[65] wl[157] vdd gnd cell_6t
Xbit_r158_c65 bl[65] br[65] wl[158] vdd gnd cell_6t
Xbit_r159_c65 bl[65] br[65] wl[159] vdd gnd cell_6t
Xbit_r160_c65 bl[65] br[65] wl[160] vdd gnd cell_6t
Xbit_r161_c65 bl[65] br[65] wl[161] vdd gnd cell_6t
Xbit_r162_c65 bl[65] br[65] wl[162] vdd gnd cell_6t
Xbit_r163_c65 bl[65] br[65] wl[163] vdd gnd cell_6t
Xbit_r164_c65 bl[65] br[65] wl[164] vdd gnd cell_6t
Xbit_r165_c65 bl[65] br[65] wl[165] vdd gnd cell_6t
Xbit_r166_c65 bl[65] br[65] wl[166] vdd gnd cell_6t
Xbit_r167_c65 bl[65] br[65] wl[167] vdd gnd cell_6t
Xbit_r168_c65 bl[65] br[65] wl[168] vdd gnd cell_6t
Xbit_r169_c65 bl[65] br[65] wl[169] vdd gnd cell_6t
Xbit_r170_c65 bl[65] br[65] wl[170] vdd gnd cell_6t
Xbit_r171_c65 bl[65] br[65] wl[171] vdd gnd cell_6t
Xbit_r172_c65 bl[65] br[65] wl[172] vdd gnd cell_6t
Xbit_r173_c65 bl[65] br[65] wl[173] vdd gnd cell_6t
Xbit_r174_c65 bl[65] br[65] wl[174] vdd gnd cell_6t
Xbit_r175_c65 bl[65] br[65] wl[175] vdd gnd cell_6t
Xbit_r176_c65 bl[65] br[65] wl[176] vdd gnd cell_6t
Xbit_r177_c65 bl[65] br[65] wl[177] vdd gnd cell_6t
Xbit_r178_c65 bl[65] br[65] wl[178] vdd gnd cell_6t
Xbit_r179_c65 bl[65] br[65] wl[179] vdd gnd cell_6t
Xbit_r180_c65 bl[65] br[65] wl[180] vdd gnd cell_6t
Xbit_r181_c65 bl[65] br[65] wl[181] vdd gnd cell_6t
Xbit_r182_c65 bl[65] br[65] wl[182] vdd gnd cell_6t
Xbit_r183_c65 bl[65] br[65] wl[183] vdd gnd cell_6t
Xbit_r184_c65 bl[65] br[65] wl[184] vdd gnd cell_6t
Xbit_r185_c65 bl[65] br[65] wl[185] vdd gnd cell_6t
Xbit_r186_c65 bl[65] br[65] wl[186] vdd gnd cell_6t
Xbit_r187_c65 bl[65] br[65] wl[187] vdd gnd cell_6t
Xbit_r188_c65 bl[65] br[65] wl[188] vdd gnd cell_6t
Xbit_r189_c65 bl[65] br[65] wl[189] vdd gnd cell_6t
Xbit_r190_c65 bl[65] br[65] wl[190] vdd gnd cell_6t
Xbit_r191_c65 bl[65] br[65] wl[191] vdd gnd cell_6t
Xbit_r192_c65 bl[65] br[65] wl[192] vdd gnd cell_6t
Xbit_r193_c65 bl[65] br[65] wl[193] vdd gnd cell_6t
Xbit_r194_c65 bl[65] br[65] wl[194] vdd gnd cell_6t
Xbit_r195_c65 bl[65] br[65] wl[195] vdd gnd cell_6t
Xbit_r196_c65 bl[65] br[65] wl[196] vdd gnd cell_6t
Xbit_r197_c65 bl[65] br[65] wl[197] vdd gnd cell_6t
Xbit_r198_c65 bl[65] br[65] wl[198] vdd gnd cell_6t
Xbit_r199_c65 bl[65] br[65] wl[199] vdd gnd cell_6t
Xbit_r200_c65 bl[65] br[65] wl[200] vdd gnd cell_6t
Xbit_r201_c65 bl[65] br[65] wl[201] vdd gnd cell_6t
Xbit_r202_c65 bl[65] br[65] wl[202] vdd gnd cell_6t
Xbit_r203_c65 bl[65] br[65] wl[203] vdd gnd cell_6t
Xbit_r204_c65 bl[65] br[65] wl[204] vdd gnd cell_6t
Xbit_r205_c65 bl[65] br[65] wl[205] vdd gnd cell_6t
Xbit_r206_c65 bl[65] br[65] wl[206] vdd gnd cell_6t
Xbit_r207_c65 bl[65] br[65] wl[207] vdd gnd cell_6t
Xbit_r208_c65 bl[65] br[65] wl[208] vdd gnd cell_6t
Xbit_r209_c65 bl[65] br[65] wl[209] vdd gnd cell_6t
Xbit_r210_c65 bl[65] br[65] wl[210] vdd gnd cell_6t
Xbit_r211_c65 bl[65] br[65] wl[211] vdd gnd cell_6t
Xbit_r212_c65 bl[65] br[65] wl[212] vdd gnd cell_6t
Xbit_r213_c65 bl[65] br[65] wl[213] vdd gnd cell_6t
Xbit_r214_c65 bl[65] br[65] wl[214] vdd gnd cell_6t
Xbit_r215_c65 bl[65] br[65] wl[215] vdd gnd cell_6t
Xbit_r216_c65 bl[65] br[65] wl[216] vdd gnd cell_6t
Xbit_r217_c65 bl[65] br[65] wl[217] vdd gnd cell_6t
Xbit_r218_c65 bl[65] br[65] wl[218] vdd gnd cell_6t
Xbit_r219_c65 bl[65] br[65] wl[219] vdd gnd cell_6t
Xbit_r220_c65 bl[65] br[65] wl[220] vdd gnd cell_6t
Xbit_r221_c65 bl[65] br[65] wl[221] vdd gnd cell_6t
Xbit_r222_c65 bl[65] br[65] wl[222] vdd gnd cell_6t
Xbit_r223_c65 bl[65] br[65] wl[223] vdd gnd cell_6t
Xbit_r224_c65 bl[65] br[65] wl[224] vdd gnd cell_6t
Xbit_r225_c65 bl[65] br[65] wl[225] vdd gnd cell_6t
Xbit_r226_c65 bl[65] br[65] wl[226] vdd gnd cell_6t
Xbit_r227_c65 bl[65] br[65] wl[227] vdd gnd cell_6t
Xbit_r228_c65 bl[65] br[65] wl[228] vdd gnd cell_6t
Xbit_r229_c65 bl[65] br[65] wl[229] vdd gnd cell_6t
Xbit_r230_c65 bl[65] br[65] wl[230] vdd gnd cell_6t
Xbit_r231_c65 bl[65] br[65] wl[231] vdd gnd cell_6t
Xbit_r232_c65 bl[65] br[65] wl[232] vdd gnd cell_6t
Xbit_r233_c65 bl[65] br[65] wl[233] vdd gnd cell_6t
Xbit_r234_c65 bl[65] br[65] wl[234] vdd gnd cell_6t
Xbit_r235_c65 bl[65] br[65] wl[235] vdd gnd cell_6t
Xbit_r236_c65 bl[65] br[65] wl[236] vdd gnd cell_6t
Xbit_r237_c65 bl[65] br[65] wl[237] vdd gnd cell_6t
Xbit_r238_c65 bl[65] br[65] wl[238] vdd gnd cell_6t
Xbit_r239_c65 bl[65] br[65] wl[239] vdd gnd cell_6t
Xbit_r240_c65 bl[65] br[65] wl[240] vdd gnd cell_6t
Xbit_r241_c65 bl[65] br[65] wl[241] vdd gnd cell_6t
Xbit_r242_c65 bl[65] br[65] wl[242] vdd gnd cell_6t
Xbit_r243_c65 bl[65] br[65] wl[243] vdd gnd cell_6t
Xbit_r244_c65 bl[65] br[65] wl[244] vdd gnd cell_6t
Xbit_r245_c65 bl[65] br[65] wl[245] vdd gnd cell_6t
Xbit_r246_c65 bl[65] br[65] wl[246] vdd gnd cell_6t
Xbit_r247_c65 bl[65] br[65] wl[247] vdd gnd cell_6t
Xbit_r248_c65 bl[65] br[65] wl[248] vdd gnd cell_6t
Xbit_r249_c65 bl[65] br[65] wl[249] vdd gnd cell_6t
Xbit_r250_c65 bl[65] br[65] wl[250] vdd gnd cell_6t
Xbit_r251_c65 bl[65] br[65] wl[251] vdd gnd cell_6t
Xbit_r252_c65 bl[65] br[65] wl[252] vdd gnd cell_6t
Xbit_r253_c65 bl[65] br[65] wl[253] vdd gnd cell_6t
Xbit_r254_c65 bl[65] br[65] wl[254] vdd gnd cell_6t
Xbit_r255_c65 bl[65] br[65] wl[255] vdd gnd cell_6t
Xbit_r256_c65 bl[65] br[65] wl[256] vdd gnd cell_6t
Xbit_r257_c65 bl[65] br[65] wl[257] vdd gnd cell_6t
Xbit_r258_c65 bl[65] br[65] wl[258] vdd gnd cell_6t
Xbit_r259_c65 bl[65] br[65] wl[259] vdd gnd cell_6t
Xbit_r260_c65 bl[65] br[65] wl[260] vdd gnd cell_6t
Xbit_r261_c65 bl[65] br[65] wl[261] vdd gnd cell_6t
Xbit_r262_c65 bl[65] br[65] wl[262] vdd gnd cell_6t
Xbit_r263_c65 bl[65] br[65] wl[263] vdd gnd cell_6t
Xbit_r264_c65 bl[65] br[65] wl[264] vdd gnd cell_6t
Xbit_r265_c65 bl[65] br[65] wl[265] vdd gnd cell_6t
Xbit_r266_c65 bl[65] br[65] wl[266] vdd gnd cell_6t
Xbit_r267_c65 bl[65] br[65] wl[267] vdd gnd cell_6t
Xbit_r268_c65 bl[65] br[65] wl[268] vdd gnd cell_6t
Xbit_r269_c65 bl[65] br[65] wl[269] vdd gnd cell_6t
Xbit_r270_c65 bl[65] br[65] wl[270] vdd gnd cell_6t
Xbit_r271_c65 bl[65] br[65] wl[271] vdd gnd cell_6t
Xbit_r272_c65 bl[65] br[65] wl[272] vdd gnd cell_6t
Xbit_r273_c65 bl[65] br[65] wl[273] vdd gnd cell_6t
Xbit_r274_c65 bl[65] br[65] wl[274] vdd gnd cell_6t
Xbit_r275_c65 bl[65] br[65] wl[275] vdd gnd cell_6t
Xbit_r276_c65 bl[65] br[65] wl[276] vdd gnd cell_6t
Xbit_r277_c65 bl[65] br[65] wl[277] vdd gnd cell_6t
Xbit_r278_c65 bl[65] br[65] wl[278] vdd gnd cell_6t
Xbit_r279_c65 bl[65] br[65] wl[279] vdd gnd cell_6t
Xbit_r280_c65 bl[65] br[65] wl[280] vdd gnd cell_6t
Xbit_r281_c65 bl[65] br[65] wl[281] vdd gnd cell_6t
Xbit_r282_c65 bl[65] br[65] wl[282] vdd gnd cell_6t
Xbit_r283_c65 bl[65] br[65] wl[283] vdd gnd cell_6t
Xbit_r284_c65 bl[65] br[65] wl[284] vdd gnd cell_6t
Xbit_r285_c65 bl[65] br[65] wl[285] vdd gnd cell_6t
Xbit_r286_c65 bl[65] br[65] wl[286] vdd gnd cell_6t
Xbit_r287_c65 bl[65] br[65] wl[287] vdd gnd cell_6t
Xbit_r288_c65 bl[65] br[65] wl[288] vdd gnd cell_6t
Xbit_r289_c65 bl[65] br[65] wl[289] vdd gnd cell_6t
Xbit_r290_c65 bl[65] br[65] wl[290] vdd gnd cell_6t
Xbit_r291_c65 bl[65] br[65] wl[291] vdd gnd cell_6t
Xbit_r292_c65 bl[65] br[65] wl[292] vdd gnd cell_6t
Xbit_r293_c65 bl[65] br[65] wl[293] vdd gnd cell_6t
Xbit_r294_c65 bl[65] br[65] wl[294] vdd gnd cell_6t
Xbit_r295_c65 bl[65] br[65] wl[295] vdd gnd cell_6t
Xbit_r296_c65 bl[65] br[65] wl[296] vdd gnd cell_6t
Xbit_r297_c65 bl[65] br[65] wl[297] vdd gnd cell_6t
Xbit_r298_c65 bl[65] br[65] wl[298] vdd gnd cell_6t
Xbit_r299_c65 bl[65] br[65] wl[299] vdd gnd cell_6t
Xbit_r300_c65 bl[65] br[65] wl[300] vdd gnd cell_6t
Xbit_r301_c65 bl[65] br[65] wl[301] vdd gnd cell_6t
Xbit_r302_c65 bl[65] br[65] wl[302] vdd gnd cell_6t
Xbit_r303_c65 bl[65] br[65] wl[303] vdd gnd cell_6t
Xbit_r304_c65 bl[65] br[65] wl[304] vdd gnd cell_6t
Xbit_r305_c65 bl[65] br[65] wl[305] vdd gnd cell_6t
Xbit_r306_c65 bl[65] br[65] wl[306] vdd gnd cell_6t
Xbit_r307_c65 bl[65] br[65] wl[307] vdd gnd cell_6t
Xbit_r308_c65 bl[65] br[65] wl[308] vdd gnd cell_6t
Xbit_r309_c65 bl[65] br[65] wl[309] vdd gnd cell_6t
Xbit_r310_c65 bl[65] br[65] wl[310] vdd gnd cell_6t
Xbit_r311_c65 bl[65] br[65] wl[311] vdd gnd cell_6t
Xbit_r312_c65 bl[65] br[65] wl[312] vdd gnd cell_6t
Xbit_r313_c65 bl[65] br[65] wl[313] vdd gnd cell_6t
Xbit_r314_c65 bl[65] br[65] wl[314] vdd gnd cell_6t
Xbit_r315_c65 bl[65] br[65] wl[315] vdd gnd cell_6t
Xbit_r316_c65 bl[65] br[65] wl[316] vdd gnd cell_6t
Xbit_r317_c65 bl[65] br[65] wl[317] vdd gnd cell_6t
Xbit_r318_c65 bl[65] br[65] wl[318] vdd gnd cell_6t
Xbit_r319_c65 bl[65] br[65] wl[319] vdd gnd cell_6t
Xbit_r320_c65 bl[65] br[65] wl[320] vdd gnd cell_6t
Xbit_r321_c65 bl[65] br[65] wl[321] vdd gnd cell_6t
Xbit_r322_c65 bl[65] br[65] wl[322] vdd gnd cell_6t
Xbit_r323_c65 bl[65] br[65] wl[323] vdd gnd cell_6t
Xbit_r324_c65 bl[65] br[65] wl[324] vdd gnd cell_6t
Xbit_r325_c65 bl[65] br[65] wl[325] vdd gnd cell_6t
Xbit_r326_c65 bl[65] br[65] wl[326] vdd gnd cell_6t
Xbit_r327_c65 bl[65] br[65] wl[327] vdd gnd cell_6t
Xbit_r328_c65 bl[65] br[65] wl[328] vdd gnd cell_6t
Xbit_r329_c65 bl[65] br[65] wl[329] vdd gnd cell_6t
Xbit_r330_c65 bl[65] br[65] wl[330] vdd gnd cell_6t
Xbit_r331_c65 bl[65] br[65] wl[331] vdd gnd cell_6t
Xbit_r332_c65 bl[65] br[65] wl[332] vdd gnd cell_6t
Xbit_r333_c65 bl[65] br[65] wl[333] vdd gnd cell_6t
Xbit_r334_c65 bl[65] br[65] wl[334] vdd gnd cell_6t
Xbit_r335_c65 bl[65] br[65] wl[335] vdd gnd cell_6t
Xbit_r336_c65 bl[65] br[65] wl[336] vdd gnd cell_6t
Xbit_r337_c65 bl[65] br[65] wl[337] vdd gnd cell_6t
Xbit_r338_c65 bl[65] br[65] wl[338] vdd gnd cell_6t
Xbit_r339_c65 bl[65] br[65] wl[339] vdd gnd cell_6t
Xbit_r340_c65 bl[65] br[65] wl[340] vdd gnd cell_6t
Xbit_r341_c65 bl[65] br[65] wl[341] vdd gnd cell_6t
Xbit_r342_c65 bl[65] br[65] wl[342] vdd gnd cell_6t
Xbit_r343_c65 bl[65] br[65] wl[343] vdd gnd cell_6t
Xbit_r344_c65 bl[65] br[65] wl[344] vdd gnd cell_6t
Xbit_r345_c65 bl[65] br[65] wl[345] vdd gnd cell_6t
Xbit_r346_c65 bl[65] br[65] wl[346] vdd gnd cell_6t
Xbit_r347_c65 bl[65] br[65] wl[347] vdd gnd cell_6t
Xbit_r348_c65 bl[65] br[65] wl[348] vdd gnd cell_6t
Xbit_r349_c65 bl[65] br[65] wl[349] vdd gnd cell_6t
Xbit_r350_c65 bl[65] br[65] wl[350] vdd gnd cell_6t
Xbit_r351_c65 bl[65] br[65] wl[351] vdd gnd cell_6t
Xbit_r352_c65 bl[65] br[65] wl[352] vdd gnd cell_6t
Xbit_r353_c65 bl[65] br[65] wl[353] vdd gnd cell_6t
Xbit_r354_c65 bl[65] br[65] wl[354] vdd gnd cell_6t
Xbit_r355_c65 bl[65] br[65] wl[355] vdd gnd cell_6t
Xbit_r356_c65 bl[65] br[65] wl[356] vdd gnd cell_6t
Xbit_r357_c65 bl[65] br[65] wl[357] vdd gnd cell_6t
Xbit_r358_c65 bl[65] br[65] wl[358] vdd gnd cell_6t
Xbit_r359_c65 bl[65] br[65] wl[359] vdd gnd cell_6t
Xbit_r360_c65 bl[65] br[65] wl[360] vdd gnd cell_6t
Xbit_r361_c65 bl[65] br[65] wl[361] vdd gnd cell_6t
Xbit_r362_c65 bl[65] br[65] wl[362] vdd gnd cell_6t
Xbit_r363_c65 bl[65] br[65] wl[363] vdd gnd cell_6t
Xbit_r364_c65 bl[65] br[65] wl[364] vdd gnd cell_6t
Xbit_r365_c65 bl[65] br[65] wl[365] vdd gnd cell_6t
Xbit_r366_c65 bl[65] br[65] wl[366] vdd gnd cell_6t
Xbit_r367_c65 bl[65] br[65] wl[367] vdd gnd cell_6t
Xbit_r368_c65 bl[65] br[65] wl[368] vdd gnd cell_6t
Xbit_r369_c65 bl[65] br[65] wl[369] vdd gnd cell_6t
Xbit_r370_c65 bl[65] br[65] wl[370] vdd gnd cell_6t
Xbit_r371_c65 bl[65] br[65] wl[371] vdd gnd cell_6t
Xbit_r372_c65 bl[65] br[65] wl[372] vdd gnd cell_6t
Xbit_r373_c65 bl[65] br[65] wl[373] vdd gnd cell_6t
Xbit_r374_c65 bl[65] br[65] wl[374] vdd gnd cell_6t
Xbit_r375_c65 bl[65] br[65] wl[375] vdd gnd cell_6t
Xbit_r376_c65 bl[65] br[65] wl[376] vdd gnd cell_6t
Xbit_r377_c65 bl[65] br[65] wl[377] vdd gnd cell_6t
Xbit_r378_c65 bl[65] br[65] wl[378] vdd gnd cell_6t
Xbit_r379_c65 bl[65] br[65] wl[379] vdd gnd cell_6t
Xbit_r380_c65 bl[65] br[65] wl[380] vdd gnd cell_6t
Xbit_r381_c65 bl[65] br[65] wl[381] vdd gnd cell_6t
Xbit_r382_c65 bl[65] br[65] wl[382] vdd gnd cell_6t
Xbit_r383_c65 bl[65] br[65] wl[383] vdd gnd cell_6t
Xbit_r384_c65 bl[65] br[65] wl[384] vdd gnd cell_6t
Xbit_r385_c65 bl[65] br[65] wl[385] vdd gnd cell_6t
Xbit_r386_c65 bl[65] br[65] wl[386] vdd gnd cell_6t
Xbit_r387_c65 bl[65] br[65] wl[387] vdd gnd cell_6t
Xbit_r388_c65 bl[65] br[65] wl[388] vdd gnd cell_6t
Xbit_r389_c65 bl[65] br[65] wl[389] vdd gnd cell_6t
Xbit_r390_c65 bl[65] br[65] wl[390] vdd gnd cell_6t
Xbit_r391_c65 bl[65] br[65] wl[391] vdd gnd cell_6t
Xbit_r392_c65 bl[65] br[65] wl[392] vdd gnd cell_6t
Xbit_r393_c65 bl[65] br[65] wl[393] vdd gnd cell_6t
Xbit_r394_c65 bl[65] br[65] wl[394] vdd gnd cell_6t
Xbit_r395_c65 bl[65] br[65] wl[395] vdd gnd cell_6t
Xbit_r396_c65 bl[65] br[65] wl[396] vdd gnd cell_6t
Xbit_r397_c65 bl[65] br[65] wl[397] vdd gnd cell_6t
Xbit_r398_c65 bl[65] br[65] wl[398] vdd gnd cell_6t
Xbit_r399_c65 bl[65] br[65] wl[399] vdd gnd cell_6t
Xbit_r400_c65 bl[65] br[65] wl[400] vdd gnd cell_6t
Xbit_r401_c65 bl[65] br[65] wl[401] vdd gnd cell_6t
Xbit_r402_c65 bl[65] br[65] wl[402] vdd gnd cell_6t
Xbit_r403_c65 bl[65] br[65] wl[403] vdd gnd cell_6t
Xbit_r404_c65 bl[65] br[65] wl[404] vdd gnd cell_6t
Xbit_r405_c65 bl[65] br[65] wl[405] vdd gnd cell_6t
Xbit_r406_c65 bl[65] br[65] wl[406] vdd gnd cell_6t
Xbit_r407_c65 bl[65] br[65] wl[407] vdd gnd cell_6t
Xbit_r408_c65 bl[65] br[65] wl[408] vdd gnd cell_6t
Xbit_r409_c65 bl[65] br[65] wl[409] vdd gnd cell_6t
Xbit_r410_c65 bl[65] br[65] wl[410] vdd gnd cell_6t
Xbit_r411_c65 bl[65] br[65] wl[411] vdd gnd cell_6t
Xbit_r412_c65 bl[65] br[65] wl[412] vdd gnd cell_6t
Xbit_r413_c65 bl[65] br[65] wl[413] vdd gnd cell_6t
Xbit_r414_c65 bl[65] br[65] wl[414] vdd gnd cell_6t
Xbit_r415_c65 bl[65] br[65] wl[415] vdd gnd cell_6t
Xbit_r416_c65 bl[65] br[65] wl[416] vdd gnd cell_6t
Xbit_r417_c65 bl[65] br[65] wl[417] vdd gnd cell_6t
Xbit_r418_c65 bl[65] br[65] wl[418] vdd gnd cell_6t
Xbit_r419_c65 bl[65] br[65] wl[419] vdd gnd cell_6t
Xbit_r420_c65 bl[65] br[65] wl[420] vdd gnd cell_6t
Xbit_r421_c65 bl[65] br[65] wl[421] vdd gnd cell_6t
Xbit_r422_c65 bl[65] br[65] wl[422] vdd gnd cell_6t
Xbit_r423_c65 bl[65] br[65] wl[423] vdd gnd cell_6t
Xbit_r424_c65 bl[65] br[65] wl[424] vdd gnd cell_6t
Xbit_r425_c65 bl[65] br[65] wl[425] vdd gnd cell_6t
Xbit_r426_c65 bl[65] br[65] wl[426] vdd gnd cell_6t
Xbit_r427_c65 bl[65] br[65] wl[427] vdd gnd cell_6t
Xbit_r428_c65 bl[65] br[65] wl[428] vdd gnd cell_6t
Xbit_r429_c65 bl[65] br[65] wl[429] vdd gnd cell_6t
Xbit_r430_c65 bl[65] br[65] wl[430] vdd gnd cell_6t
Xbit_r431_c65 bl[65] br[65] wl[431] vdd gnd cell_6t
Xbit_r432_c65 bl[65] br[65] wl[432] vdd gnd cell_6t
Xbit_r433_c65 bl[65] br[65] wl[433] vdd gnd cell_6t
Xbit_r434_c65 bl[65] br[65] wl[434] vdd gnd cell_6t
Xbit_r435_c65 bl[65] br[65] wl[435] vdd gnd cell_6t
Xbit_r436_c65 bl[65] br[65] wl[436] vdd gnd cell_6t
Xbit_r437_c65 bl[65] br[65] wl[437] vdd gnd cell_6t
Xbit_r438_c65 bl[65] br[65] wl[438] vdd gnd cell_6t
Xbit_r439_c65 bl[65] br[65] wl[439] vdd gnd cell_6t
Xbit_r440_c65 bl[65] br[65] wl[440] vdd gnd cell_6t
Xbit_r441_c65 bl[65] br[65] wl[441] vdd gnd cell_6t
Xbit_r442_c65 bl[65] br[65] wl[442] vdd gnd cell_6t
Xbit_r443_c65 bl[65] br[65] wl[443] vdd gnd cell_6t
Xbit_r444_c65 bl[65] br[65] wl[444] vdd gnd cell_6t
Xbit_r445_c65 bl[65] br[65] wl[445] vdd gnd cell_6t
Xbit_r446_c65 bl[65] br[65] wl[446] vdd gnd cell_6t
Xbit_r447_c65 bl[65] br[65] wl[447] vdd gnd cell_6t
Xbit_r448_c65 bl[65] br[65] wl[448] vdd gnd cell_6t
Xbit_r449_c65 bl[65] br[65] wl[449] vdd gnd cell_6t
Xbit_r450_c65 bl[65] br[65] wl[450] vdd gnd cell_6t
Xbit_r451_c65 bl[65] br[65] wl[451] vdd gnd cell_6t
Xbit_r452_c65 bl[65] br[65] wl[452] vdd gnd cell_6t
Xbit_r453_c65 bl[65] br[65] wl[453] vdd gnd cell_6t
Xbit_r454_c65 bl[65] br[65] wl[454] vdd gnd cell_6t
Xbit_r455_c65 bl[65] br[65] wl[455] vdd gnd cell_6t
Xbit_r456_c65 bl[65] br[65] wl[456] vdd gnd cell_6t
Xbit_r457_c65 bl[65] br[65] wl[457] vdd gnd cell_6t
Xbit_r458_c65 bl[65] br[65] wl[458] vdd gnd cell_6t
Xbit_r459_c65 bl[65] br[65] wl[459] vdd gnd cell_6t
Xbit_r460_c65 bl[65] br[65] wl[460] vdd gnd cell_6t
Xbit_r461_c65 bl[65] br[65] wl[461] vdd gnd cell_6t
Xbit_r462_c65 bl[65] br[65] wl[462] vdd gnd cell_6t
Xbit_r463_c65 bl[65] br[65] wl[463] vdd gnd cell_6t
Xbit_r464_c65 bl[65] br[65] wl[464] vdd gnd cell_6t
Xbit_r465_c65 bl[65] br[65] wl[465] vdd gnd cell_6t
Xbit_r466_c65 bl[65] br[65] wl[466] vdd gnd cell_6t
Xbit_r467_c65 bl[65] br[65] wl[467] vdd gnd cell_6t
Xbit_r468_c65 bl[65] br[65] wl[468] vdd gnd cell_6t
Xbit_r469_c65 bl[65] br[65] wl[469] vdd gnd cell_6t
Xbit_r470_c65 bl[65] br[65] wl[470] vdd gnd cell_6t
Xbit_r471_c65 bl[65] br[65] wl[471] vdd gnd cell_6t
Xbit_r472_c65 bl[65] br[65] wl[472] vdd gnd cell_6t
Xbit_r473_c65 bl[65] br[65] wl[473] vdd gnd cell_6t
Xbit_r474_c65 bl[65] br[65] wl[474] vdd gnd cell_6t
Xbit_r475_c65 bl[65] br[65] wl[475] vdd gnd cell_6t
Xbit_r476_c65 bl[65] br[65] wl[476] vdd gnd cell_6t
Xbit_r477_c65 bl[65] br[65] wl[477] vdd gnd cell_6t
Xbit_r478_c65 bl[65] br[65] wl[478] vdd gnd cell_6t
Xbit_r479_c65 bl[65] br[65] wl[479] vdd gnd cell_6t
Xbit_r480_c65 bl[65] br[65] wl[480] vdd gnd cell_6t
Xbit_r481_c65 bl[65] br[65] wl[481] vdd gnd cell_6t
Xbit_r482_c65 bl[65] br[65] wl[482] vdd gnd cell_6t
Xbit_r483_c65 bl[65] br[65] wl[483] vdd gnd cell_6t
Xbit_r484_c65 bl[65] br[65] wl[484] vdd gnd cell_6t
Xbit_r485_c65 bl[65] br[65] wl[485] vdd gnd cell_6t
Xbit_r486_c65 bl[65] br[65] wl[486] vdd gnd cell_6t
Xbit_r487_c65 bl[65] br[65] wl[487] vdd gnd cell_6t
Xbit_r488_c65 bl[65] br[65] wl[488] vdd gnd cell_6t
Xbit_r489_c65 bl[65] br[65] wl[489] vdd gnd cell_6t
Xbit_r490_c65 bl[65] br[65] wl[490] vdd gnd cell_6t
Xbit_r491_c65 bl[65] br[65] wl[491] vdd gnd cell_6t
Xbit_r492_c65 bl[65] br[65] wl[492] vdd gnd cell_6t
Xbit_r493_c65 bl[65] br[65] wl[493] vdd gnd cell_6t
Xbit_r494_c65 bl[65] br[65] wl[494] vdd gnd cell_6t
Xbit_r495_c65 bl[65] br[65] wl[495] vdd gnd cell_6t
Xbit_r496_c65 bl[65] br[65] wl[496] vdd gnd cell_6t
Xbit_r497_c65 bl[65] br[65] wl[497] vdd gnd cell_6t
Xbit_r498_c65 bl[65] br[65] wl[498] vdd gnd cell_6t
Xbit_r499_c65 bl[65] br[65] wl[499] vdd gnd cell_6t
Xbit_r500_c65 bl[65] br[65] wl[500] vdd gnd cell_6t
Xbit_r501_c65 bl[65] br[65] wl[501] vdd gnd cell_6t
Xbit_r502_c65 bl[65] br[65] wl[502] vdd gnd cell_6t
Xbit_r503_c65 bl[65] br[65] wl[503] vdd gnd cell_6t
Xbit_r504_c65 bl[65] br[65] wl[504] vdd gnd cell_6t
Xbit_r505_c65 bl[65] br[65] wl[505] vdd gnd cell_6t
Xbit_r506_c65 bl[65] br[65] wl[506] vdd gnd cell_6t
Xbit_r507_c65 bl[65] br[65] wl[507] vdd gnd cell_6t
Xbit_r508_c65 bl[65] br[65] wl[508] vdd gnd cell_6t
Xbit_r509_c65 bl[65] br[65] wl[509] vdd gnd cell_6t
Xbit_r510_c65 bl[65] br[65] wl[510] vdd gnd cell_6t
Xbit_r511_c65 bl[65] br[65] wl[511] vdd gnd cell_6t
Xbit_r0_c66 bl[66] br[66] wl[0] vdd gnd cell_6t
Xbit_r1_c66 bl[66] br[66] wl[1] vdd gnd cell_6t
Xbit_r2_c66 bl[66] br[66] wl[2] vdd gnd cell_6t
Xbit_r3_c66 bl[66] br[66] wl[3] vdd gnd cell_6t
Xbit_r4_c66 bl[66] br[66] wl[4] vdd gnd cell_6t
Xbit_r5_c66 bl[66] br[66] wl[5] vdd gnd cell_6t
Xbit_r6_c66 bl[66] br[66] wl[6] vdd gnd cell_6t
Xbit_r7_c66 bl[66] br[66] wl[7] vdd gnd cell_6t
Xbit_r8_c66 bl[66] br[66] wl[8] vdd gnd cell_6t
Xbit_r9_c66 bl[66] br[66] wl[9] vdd gnd cell_6t
Xbit_r10_c66 bl[66] br[66] wl[10] vdd gnd cell_6t
Xbit_r11_c66 bl[66] br[66] wl[11] vdd gnd cell_6t
Xbit_r12_c66 bl[66] br[66] wl[12] vdd gnd cell_6t
Xbit_r13_c66 bl[66] br[66] wl[13] vdd gnd cell_6t
Xbit_r14_c66 bl[66] br[66] wl[14] vdd gnd cell_6t
Xbit_r15_c66 bl[66] br[66] wl[15] vdd gnd cell_6t
Xbit_r16_c66 bl[66] br[66] wl[16] vdd gnd cell_6t
Xbit_r17_c66 bl[66] br[66] wl[17] vdd gnd cell_6t
Xbit_r18_c66 bl[66] br[66] wl[18] vdd gnd cell_6t
Xbit_r19_c66 bl[66] br[66] wl[19] vdd gnd cell_6t
Xbit_r20_c66 bl[66] br[66] wl[20] vdd gnd cell_6t
Xbit_r21_c66 bl[66] br[66] wl[21] vdd gnd cell_6t
Xbit_r22_c66 bl[66] br[66] wl[22] vdd gnd cell_6t
Xbit_r23_c66 bl[66] br[66] wl[23] vdd gnd cell_6t
Xbit_r24_c66 bl[66] br[66] wl[24] vdd gnd cell_6t
Xbit_r25_c66 bl[66] br[66] wl[25] vdd gnd cell_6t
Xbit_r26_c66 bl[66] br[66] wl[26] vdd gnd cell_6t
Xbit_r27_c66 bl[66] br[66] wl[27] vdd gnd cell_6t
Xbit_r28_c66 bl[66] br[66] wl[28] vdd gnd cell_6t
Xbit_r29_c66 bl[66] br[66] wl[29] vdd gnd cell_6t
Xbit_r30_c66 bl[66] br[66] wl[30] vdd gnd cell_6t
Xbit_r31_c66 bl[66] br[66] wl[31] vdd gnd cell_6t
Xbit_r32_c66 bl[66] br[66] wl[32] vdd gnd cell_6t
Xbit_r33_c66 bl[66] br[66] wl[33] vdd gnd cell_6t
Xbit_r34_c66 bl[66] br[66] wl[34] vdd gnd cell_6t
Xbit_r35_c66 bl[66] br[66] wl[35] vdd gnd cell_6t
Xbit_r36_c66 bl[66] br[66] wl[36] vdd gnd cell_6t
Xbit_r37_c66 bl[66] br[66] wl[37] vdd gnd cell_6t
Xbit_r38_c66 bl[66] br[66] wl[38] vdd gnd cell_6t
Xbit_r39_c66 bl[66] br[66] wl[39] vdd gnd cell_6t
Xbit_r40_c66 bl[66] br[66] wl[40] vdd gnd cell_6t
Xbit_r41_c66 bl[66] br[66] wl[41] vdd gnd cell_6t
Xbit_r42_c66 bl[66] br[66] wl[42] vdd gnd cell_6t
Xbit_r43_c66 bl[66] br[66] wl[43] vdd gnd cell_6t
Xbit_r44_c66 bl[66] br[66] wl[44] vdd gnd cell_6t
Xbit_r45_c66 bl[66] br[66] wl[45] vdd gnd cell_6t
Xbit_r46_c66 bl[66] br[66] wl[46] vdd gnd cell_6t
Xbit_r47_c66 bl[66] br[66] wl[47] vdd gnd cell_6t
Xbit_r48_c66 bl[66] br[66] wl[48] vdd gnd cell_6t
Xbit_r49_c66 bl[66] br[66] wl[49] vdd gnd cell_6t
Xbit_r50_c66 bl[66] br[66] wl[50] vdd gnd cell_6t
Xbit_r51_c66 bl[66] br[66] wl[51] vdd gnd cell_6t
Xbit_r52_c66 bl[66] br[66] wl[52] vdd gnd cell_6t
Xbit_r53_c66 bl[66] br[66] wl[53] vdd gnd cell_6t
Xbit_r54_c66 bl[66] br[66] wl[54] vdd gnd cell_6t
Xbit_r55_c66 bl[66] br[66] wl[55] vdd gnd cell_6t
Xbit_r56_c66 bl[66] br[66] wl[56] vdd gnd cell_6t
Xbit_r57_c66 bl[66] br[66] wl[57] vdd gnd cell_6t
Xbit_r58_c66 bl[66] br[66] wl[58] vdd gnd cell_6t
Xbit_r59_c66 bl[66] br[66] wl[59] vdd gnd cell_6t
Xbit_r60_c66 bl[66] br[66] wl[60] vdd gnd cell_6t
Xbit_r61_c66 bl[66] br[66] wl[61] vdd gnd cell_6t
Xbit_r62_c66 bl[66] br[66] wl[62] vdd gnd cell_6t
Xbit_r63_c66 bl[66] br[66] wl[63] vdd gnd cell_6t
Xbit_r64_c66 bl[66] br[66] wl[64] vdd gnd cell_6t
Xbit_r65_c66 bl[66] br[66] wl[65] vdd gnd cell_6t
Xbit_r66_c66 bl[66] br[66] wl[66] vdd gnd cell_6t
Xbit_r67_c66 bl[66] br[66] wl[67] vdd gnd cell_6t
Xbit_r68_c66 bl[66] br[66] wl[68] vdd gnd cell_6t
Xbit_r69_c66 bl[66] br[66] wl[69] vdd gnd cell_6t
Xbit_r70_c66 bl[66] br[66] wl[70] vdd gnd cell_6t
Xbit_r71_c66 bl[66] br[66] wl[71] vdd gnd cell_6t
Xbit_r72_c66 bl[66] br[66] wl[72] vdd gnd cell_6t
Xbit_r73_c66 bl[66] br[66] wl[73] vdd gnd cell_6t
Xbit_r74_c66 bl[66] br[66] wl[74] vdd gnd cell_6t
Xbit_r75_c66 bl[66] br[66] wl[75] vdd gnd cell_6t
Xbit_r76_c66 bl[66] br[66] wl[76] vdd gnd cell_6t
Xbit_r77_c66 bl[66] br[66] wl[77] vdd gnd cell_6t
Xbit_r78_c66 bl[66] br[66] wl[78] vdd gnd cell_6t
Xbit_r79_c66 bl[66] br[66] wl[79] vdd gnd cell_6t
Xbit_r80_c66 bl[66] br[66] wl[80] vdd gnd cell_6t
Xbit_r81_c66 bl[66] br[66] wl[81] vdd gnd cell_6t
Xbit_r82_c66 bl[66] br[66] wl[82] vdd gnd cell_6t
Xbit_r83_c66 bl[66] br[66] wl[83] vdd gnd cell_6t
Xbit_r84_c66 bl[66] br[66] wl[84] vdd gnd cell_6t
Xbit_r85_c66 bl[66] br[66] wl[85] vdd gnd cell_6t
Xbit_r86_c66 bl[66] br[66] wl[86] vdd gnd cell_6t
Xbit_r87_c66 bl[66] br[66] wl[87] vdd gnd cell_6t
Xbit_r88_c66 bl[66] br[66] wl[88] vdd gnd cell_6t
Xbit_r89_c66 bl[66] br[66] wl[89] vdd gnd cell_6t
Xbit_r90_c66 bl[66] br[66] wl[90] vdd gnd cell_6t
Xbit_r91_c66 bl[66] br[66] wl[91] vdd gnd cell_6t
Xbit_r92_c66 bl[66] br[66] wl[92] vdd gnd cell_6t
Xbit_r93_c66 bl[66] br[66] wl[93] vdd gnd cell_6t
Xbit_r94_c66 bl[66] br[66] wl[94] vdd gnd cell_6t
Xbit_r95_c66 bl[66] br[66] wl[95] vdd gnd cell_6t
Xbit_r96_c66 bl[66] br[66] wl[96] vdd gnd cell_6t
Xbit_r97_c66 bl[66] br[66] wl[97] vdd gnd cell_6t
Xbit_r98_c66 bl[66] br[66] wl[98] vdd gnd cell_6t
Xbit_r99_c66 bl[66] br[66] wl[99] vdd gnd cell_6t
Xbit_r100_c66 bl[66] br[66] wl[100] vdd gnd cell_6t
Xbit_r101_c66 bl[66] br[66] wl[101] vdd gnd cell_6t
Xbit_r102_c66 bl[66] br[66] wl[102] vdd gnd cell_6t
Xbit_r103_c66 bl[66] br[66] wl[103] vdd gnd cell_6t
Xbit_r104_c66 bl[66] br[66] wl[104] vdd gnd cell_6t
Xbit_r105_c66 bl[66] br[66] wl[105] vdd gnd cell_6t
Xbit_r106_c66 bl[66] br[66] wl[106] vdd gnd cell_6t
Xbit_r107_c66 bl[66] br[66] wl[107] vdd gnd cell_6t
Xbit_r108_c66 bl[66] br[66] wl[108] vdd gnd cell_6t
Xbit_r109_c66 bl[66] br[66] wl[109] vdd gnd cell_6t
Xbit_r110_c66 bl[66] br[66] wl[110] vdd gnd cell_6t
Xbit_r111_c66 bl[66] br[66] wl[111] vdd gnd cell_6t
Xbit_r112_c66 bl[66] br[66] wl[112] vdd gnd cell_6t
Xbit_r113_c66 bl[66] br[66] wl[113] vdd gnd cell_6t
Xbit_r114_c66 bl[66] br[66] wl[114] vdd gnd cell_6t
Xbit_r115_c66 bl[66] br[66] wl[115] vdd gnd cell_6t
Xbit_r116_c66 bl[66] br[66] wl[116] vdd gnd cell_6t
Xbit_r117_c66 bl[66] br[66] wl[117] vdd gnd cell_6t
Xbit_r118_c66 bl[66] br[66] wl[118] vdd gnd cell_6t
Xbit_r119_c66 bl[66] br[66] wl[119] vdd gnd cell_6t
Xbit_r120_c66 bl[66] br[66] wl[120] vdd gnd cell_6t
Xbit_r121_c66 bl[66] br[66] wl[121] vdd gnd cell_6t
Xbit_r122_c66 bl[66] br[66] wl[122] vdd gnd cell_6t
Xbit_r123_c66 bl[66] br[66] wl[123] vdd gnd cell_6t
Xbit_r124_c66 bl[66] br[66] wl[124] vdd gnd cell_6t
Xbit_r125_c66 bl[66] br[66] wl[125] vdd gnd cell_6t
Xbit_r126_c66 bl[66] br[66] wl[126] vdd gnd cell_6t
Xbit_r127_c66 bl[66] br[66] wl[127] vdd gnd cell_6t
Xbit_r128_c66 bl[66] br[66] wl[128] vdd gnd cell_6t
Xbit_r129_c66 bl[66] br[66] wl[129] vdd gnd cell_6t
Xbit_r130_c66 bl[66] br[66] wl[130] vdd gnd cell_6t
Xbit_r131_c66 bl[66] br[66] wl[131] vdd gnd cell_6t
Xbit_r132_c66 bl[66] br[66] wl[132] vdd gnd cell_6t
Xbit_r133_c66 bl[66] br[66] wl[133] vdd gnd cell_6t
Xbit_r134_c66 bl[66] br[66] wl[134] vdd gnd cell_6t
Xbit_r135_c66 bl[66] br[66] wl[135] vdd gnd cell_6t
Xbit_r136_c66 bl[66] br[66] wl[136] vdd gnd cell_6t
Xbit_r137_c66 bl[66] br[66] wl[137] vdd gnd cell_6t
Xbit_r138_c66 bl[66] br[66] wl[138] vdd gnd cell_6t
Xbit_r139_c66 bl[66] br[66] wl[139] vdd gnd cell_6t
Xbit_r140_c66 bl[66] br[66] wl[140] vdd gnd cell_6t
Xbit_r141_c66 bl[66] br[66] wl[141] vdd gnd cell_6t
Xbit_r142_c66 bl[66] br[66] wl[142] vdd gnd cell_6t
Xbit_r143_c66 bl[66] br[66] wl[143] vdd gnd cell_6t
Xbit_r144_c66 bl[66] br[66] wl[144] vdd gnd cell_6t
Xbit_r145_c66 bl[66] br[66] wl[145] vdd gnd cell_6t
Xbit_r146_c66 bl[66] br[66] wl[146] vdd gnd cell_6t
Xbit_r147_c66 bl[66] br[66] wl[147] vdd gnd cell_6t
Xbit_r148_c66 bl[66] br[66] wl[148] vdd gnd cell_6t
Xbit_r149_c66 bl[66] br[66] wl[149] vdd gnd cell_6t
Xbit_r150_c66 bl[66] br[66] wl[150] vdd gnd cell_6t
Xbit_r151_c66 bl[66] br[66] wl[151] vdd gnd cell_6t
Xbit_r152_c66 bl[66] br[66] wl[152] vdd gnd cell_6t
Xbit_r153_c66 bl[66] br[66] wl[153] vdd gnd cell_6t
Xbit_r154_c66 bl[66] br[66] wl[154] vdd gnd cell_6t
Xbit_r155_c66 bl[66] br[66] wl[155] vdd gnd cell_6t
Xbit_r156_c66 bl[66] br[66] wl[156] vdd gnd cell_6t
Xbit_r157_c66 bl[66] br[66] wl[157] vdd gnd cell_6t
Xbit_r158_c66 bl[66] br[66] wl[158] vdd gnd cell_6t
Xbit_r159_c66 bl[66] br[66] wl[159] vdd gnd cell_6t
Xbit_r160_c66 bl[66] br[66] wl[160] vdd gnd cell_6t
Xbit_r161_c66 bl[66] br[66] wl[161] vdd gnd cell_6t
Xbit_r162_c66 bl[66] br[66] wl[162] vdd gnd cell_6t
Xbit_r163_c66 bl[66] br[66] wl[163] vdd gnd cell_6t
Xbit_r164_c66 bl[66] br[66] wl[164] vdd gnd cell_6t
Xbit_r165_c66 bl[66] br[66] wl[165] vdd gnd cell_6t
Xbit_r166_c66 bl[66] br[66] wl[166] vdd gnd cell_6t
Xbit_r167_c66 bl[66] br[66] wl[167] vdd gnd cell_6t
Xbit_r168_c66 bl[66] br[66] wl[168] vdd gnd cell_6t
Xbit_r169_c66 bl[66] br[66] wl[169] vdd gnd cell_6t
Xbit_r170_c66 bl[66] br[66] wl[170] vdd gnd cell_6t
Xbit_r171_c66 bl[66] br[66] wl[171] vdd gnd cell_6t
Xbit_r172_c66 bl[66] br[66] wl[172] vdd gnd cell_6t
Xbit_r173_c66 bl[66] br[66] wl[173] vdd gnd cell_6t
Xbit_r174_c66 bl[66] br[66] wl[174] vdd gnd cell_6t
Xbit_r175_c66 bl[66] br[66] wl[175] vdd gnd cell_6t
Xbit_r176_c66 bl[66] br[66] wl[176] vdd gnd cell_6t
Xbit_r177_c66 bl[66] br[66] wl[177] vdd gnd cell_6t
Xbit_r178_c66 bl[66] br[66] wl[178] vdd gnd cell_6t
Xbit_r179_c66 bl[66] br[66] wl[179] vdd gnd cell_6t
Xbit_r180_c66 bl[66] br[66] wl[180] vdd gnd cell_6t
Xbit_r181_c66 bl[66] br[66] wl[181] vdd gnd cell_6t
Xbit_r182_c66 bl[66] br[66] wl[182] vdd gnd cell_6t
Xbit_r183_c66 bl[66] br[66] wl[183] vdd gnd cell_6t
Xbit_r184_c66 bl[66] br[66] wl[184] vdd gnd cell_6t
Xbit_r185_c66 bl[66] br[66] wl[185] vdd gnd cell_6t
Xbit_r186_c66 bl[66] br[66] wl[186] vdd gnd cell_6t
Xbit_r187_c66 bl[66] br[66] wl[187] vdd gnd cell_6t
Xbit_r188_c66 bl[66] br[66] wl[188] vdd gnd cell_6t
Xbit_r189_c66 bl[66] br[66] wl[189] vdd gnd cell_6t
Xbit_r190_c66 bl[66] br[66] wl[190] vdd gnd cell_6t
Xbit_r191_c66 bl[66] br[66] wl[191] vdd gnd cell_6t
Xbit_r192_c66 bl[66] br[66] wl[192] vdd gnd cell_6t
Xbit_r193_c66 bl[66] br[66] wl[193] vdd gnd cell_6t
Xbit_r194_c66 bl[66] br[66] wl[194] vdd gnd cell_6t
Xbit_r195_c66 bl[66] br[66] wl[195] vdd gnd cell_6t
Xbit_r196_c66 bl[66] br[66] wl[196] vdd gnd cell_6t
Xbit_r197_c66 bl[66] br[66] wl[197] vdd gnd cell_6t
Xbit_r198_c66 bl[66] br[66] wl[198] vdd gnd cell_6t
Xbit_r199_c66 bl[66] br[66] wl[199] vdd gnd cell_6t
Xbit_r200_c66 bl[66] br[66] wl[200] vdd gnd cell_6t
Xbit_r201_c66 bl[66] br[66] wl[201] vdd gnd cell_6t
Xbit_r202_c66 bl[66] br[66] wl[202] vdd gnd cell_6t
Xbit_r203_c66 bl[66] br[66] wl[203] vdd gnd cell_6t
Xbit_r204_c66 bl[66] br[66] wl[204] vdd gnd cell_6t
Xbit_r205_c66 bl[66] br[66] wl[205] vdd gnd cell_6t
Xbit_r206_c66 bl[66] br[66] wl[206] vdd gnd cell_6t
Xbit_r207_c66 bl[66] br[66] wl[207] vdd gnd cell_6t
Xbit_r208_c66 bl[66] br[66] wl[208] vdd gnd cell_6t
Xbit_r209_c66 bl[66] br[66] wl[209] vdd gnd cell_6t
Xbit_r210_c66 bl[66] br[66] wl[210] vdd gnd cell_6t
Xbit_r211_c66 bl[66] br[66] wl[211] vdd gnd cell_6t
Xbit_r212_c66 bl[66] br[66] wl[212] vdd gnd cell_6t
Xbit_r213_c66 bl[66] br[66] wl[213] vdd gnd cell_6t
Xbit_r214_c66 bl[66] br[66] wl[214] vdd gnd cell_6t
Xbit_r215_c66 bl[66] br[66] wl[215] vdd gnd cell_6t
Xbit_r216_c66 bl[66] br[66] wl[216] vdd gnd cell_6t
Xbit_r217_c66 bl[66] br[66] wl[217] vdd gnd cell_6t
Xbit_r218_c66 bl[66] br[66] wl[218] vdd gnd cell_6t
Xbit_r219_c66 bl[66] br[66] wl[219] vdd gnd cell_6t
Xbit_r220_c66 bl[66] br[66] wl[220] vdd gnd cell_6t
Xbit_r221_c66 bl[66] br[66] wl[221] vdd gnd cell_6t
Xbit_r222_c66 bl[66] br[66] wl[222] vdd gnd cell_6t
Xbit_r223_c66 bl[66] br[66] wl[223] vdd gnd cell_6t
Xbit_r224_c66 bl[66] br[66] wl[224] vdd gnd cell_6t
Xbit_r225_c66 bl[66] br[66] wl[225] vdd gnd cell_6t
Xbit_r226_c66 bl[66] br[66] wl[226] vdd gnd cell_6t
Xbit_r227_c66 bl[66] br[66] wl[227] vdd gnd cell_6t
Xbit_r228_c66 bl[66] br[66] wl[228] vdd gnd cell_6t
Xbit_r229_c66 bl[66] br[66] wl[229] vdd gnd cell_6t
Xbit_r230_c66 bl[66] br[66] wl[230] vdd gnd cell_6t
Xbit_r231_c66 bl[66] br[66] wl[231] vdd gnd cell_6t
Xbit_r232_c66 bl[66] br[66] wl[232] vdd gnd cell_6t
Xbit_r233_c66 bl[66] br[66] wl[233] vdd gnd cell_6t
Xbit_r234_c66 bl[66] br[66] wl[234] vdd gnd cell_6t
Xbit_r235_c66 bl[66] br[66] wl[235] vdd gnd cell_6t
Xbit_r236_c66 bl[66] br[66] wl[236] vdd gnd cell_6t
Xbit_r237_c66 bl[66] br[66] wl[237] vdd gnd cell_6t
Xbit_r238_c66 bl[66] br[66] wl[238] vdd gnd cell_6t
Xbit_r239_c66 bl[66] br[66] wl[239] vdd gnd cell_6t
Xbit_r240_c66 bl[66] br[66] wl[240] vdd gnd cell_6t
Xbit_r241_c66 bl[66] br[66] wl[241] vdd gnd cell_6t
Xbit_r242_c66 bl[66] br[66] wl[242] vdd gnd cell_6t
Xbit_r243_c66 bl[66] br[66] wl[243] vdd gnd cell_6t
Xbit_r244_c66 bl[66] br[66] wl[244] vdd gnd cell_6t
Xbit_r245_c66 bl[66] br[66] wl[245] vdd gnd cell_6t
Xbit_r246_c66 bl[66] br[66] wl[246] vdd gnd cell_6t
Xbit_r247_c66 bl[66] br[66] wl[247] vdd gnd cell_6t
Xbit_r248_c66 bl[66] br[66] wl[248] vdd gnd cell_6t
Xbit_r249_c66 bl[66] br[66] wl[249] vdd gnd cell_6t
Xbit_r250_c66 bl[66] br[66] wl[250] vdd gnd cell_6t
Xbit_r251_c66 bl[66] br[66] wl[251] vdd gnd cell_6t
Xbit_r252_c66 bl[66] br[66] wl[252] vdd gnd cell_6t
Xbit_r253_c66 bl[66] br[66] wl[253] vdd gnd cell_6t
Xbit_r254_c66 bl[66] br[66] wl[254] vdd gnd cell_6t
Xbit_r255_c66 bl[66] br[66] wl[255] vdd gnd cell_6t
Xbit_r256_c66 bl[66] br[66] wl[256] vdd gnd cell_6t
Xbit_r257_c66 bl[66] br[66] wl[257] vdd gnd cell_6t
Xbit_r258_c66 bl[66] br[66] wl[258] vdd gnd cell_6t
Xbit_r259_c66 bl[66] br[66] wl[259] vdd gnd cell_6t
Xbit_r260_c66 bl[66] br[66] wl[260] vdd gnd cell_6t
Xbit_r261_c66 bl[66] br[66] wl[261] vdd gnd cell_6t
Xbit_r262_c66 bl[66] br[66] wl[262] vdd gnd cell_6t
Xbit_r263_c66 bl[66] br[66] wl[263] vdd gnd cell_6t
Xbit_r264_c66 bl[66] br[66] wl[264] vdd gnd cell_6t
Xbit_r265_c66 bl[66] br[66] wl[265] vdd gnd cell_6t
Xbit_r266_c66 bl[66] br[66] wl[266] vdd gnd cell_6t
Xbit_r267_c66 bl[66] br[66] wl[267] vdd gnd cell_6t
Xbit_r268_c66 bl[66] br[66] wl[268] vdd gnd cell_6t
Xbit_r269_c66 bl[66] br[66] wl[269] vdd gnd cell_6t
Xbit_r270_c66 bl[66] br[66] wl[270] vdd gnd cell_6t
Xbit_r271_c66 bl[66] br[66] wl[271] vdd gnd cell_6t
Xbit_r272_c66 bl[66] br[66] wl[272] vdd gnd cell_6t
Xbit_r273_c66 bl[66] br[66] wl[273] vdd gnd cell_6t
Xbit_r274_c66 bl[66] br[66] wl[274] vdd gnd cell_6t
Xbit_r275_c66 bl[66] br[66] wl[275] vdd gnd cell_6t
Xbit_r276_c66 bl[66] br[66] wl[276] vdd gnd cell_6t
Xbit_r277_c66 bl[66] br[66] wl[277] vdd gnd cell_6t
Xbit_r278_c66 bl[66] br[66] wl[278] vdd gnd cell_6t
Xbit_r279_c66 bl[66] br[66] wl[279] vdd gnd cell_6t
Xbit_r280_c66 bl[66] br[66] wl[280] vdd gnd cell_6t
Xbit_r281_c66 bl[66] br[66] wl[281] vdd gnd cell_6t
Xbit_r282_c66 bl[66] br[66] wl[282] vdd gnd cell_6t
Xbit_r283_c66 bl[66] br[66] wl[283] vdd gnd cell_6t
Xbit_r284_c66 bl[66] br[66] wl[284] vdd gnd cell_6t
Xbit_r285_c66 bl[66] br[66] wl[285] vdd gnd cell_6t
Xbit_r286_c66 bl[66] br[66] wl[286] vdd gnd cell_6t
Xbit_r287_c66 bl[66] br[66] wl[287] vdd gnd cell_6t
Xbit_r288_c66 bl[66] br[66] wl[288] vdd gnd cell_6t
Xbit_r289_c66 bl[66] br[66] wl[289] vdd gnd cell_6t
Xbit_r290_c66 bl[66] br[66] wl[290] vdd gnd cell_6t
Xbit_r291_c66 bl[66] br[66] wl[291] vdd gnd cell_6t
Xbit_r292_c66 bl[66] br[66] wl[292] vdd gnd cell_6t
Xbit_r293_c66 bl[66] br[66] wl[293] vdd gnd cell_6t
Xbit_r294_c66 bl[66] br[66] wl[294] vdd gnd cell_6t
Xbit_r295_c66 bl[66] br[66] wl[295] vdd gnd cell_6t
Xbit_r296_c66 bl[66] br[66] wl[296] vdd gnd cell_6t
Xbit_r297_c66 bl[66] br[66] wl[297] vdd gnd cell_6t
Xbit_r298_c66 bl[66] br[66] wl[298] vdd gnd cell_6t
Xbit_r299_c66 bl[66] br[66] wl[299] vdd gnd cell_6t
Xbit_r300_c66 bl[66] br[66] wl[300] vdd gnd cell_6t
Xbit_r301_c66 bl[66] br[66] wl[301] vdd gnd cell_6t
Xbit_r302_c66 bl[66] br[66] wl[302] vdd gnd cell_6t
Xbit_r303_c66 bl[66] br[66] wl[303] vdd gnd cell_6t
Xbit_r304_c66 bl[66] br[66] wl[304] vdd gnd cell_6t
Xbit_r305_c66 bl[66] br[66] wl[305] vdd gnd cell_6t
Xbit_r306_c66 bl[66] br[66] wl[306] vdd gnd cell_6t
Xbit_r307_c66 bl[66] br[66] wl[307] vdd gnd cell_6t
Xbit_r308_c66 bl[66] br[66] wl[308] vdd gnd cell_6t
Xbit_r309_c66 bl[66] br[66] wl[309] vdd gnd cell_6t
Xbit_r310_c66 bl[66] br[66] wl[310] vdd gnd cell_6t
Xbit_r311_c66 bl[66] br[66] wl[311] vdd gnd cell_6t
Xbit_r312_c66 bl[66] br[66] wl[312] vdd gnd cell_6t
Xbit_r313_c66 bl[66] br[66] wl[313] vdd gnd cell_6t
Xbit_r314_c66 bl[66] br[66] wl[314] vdd gnd cell_6t
Xbit_r315_c66 bl[66] br[66] wl[315] vdd gnd cell_6t
Xbit_r316_c66 bl[66] br[66] wl[316] vdd gnd cell_6t
Xbit_r317_c66 bl[66] br[66] wl[317] vdd gnd cell_6t
Xbit_r318_c66 bl[66] br[66] wl[318] vdd gnd cell_6t
Xbit_r319_c66 bl[66] br[66] wl[319] vdd gnd cell_6t
Xbit_r320_c66 bl[66] br[66] wl[320] vdd gnd cell_6t
Xbit_r321_c66 bl[66] br[66] wl[321] vdd gnd cell_6t
Xbit_r322_c66 bl[66] br[66] wl[322] vdd gnd cell_6t
Xbit_r323_c66 bl[66] br[66] wl[323] vdd gnd cell_6t
Xbit_r324_c66 bl[66] br[66] wl[324] vdd gnd cell_6t
Xbit_r325_c66 bl[66] br[66] wl[325] vdd gnd cell_6t
Xbit_r326_c66 bl[66] br[66] wl[326] vdd gnd cell_6t
Xbit_r327_c66 bl[66] br[66] wl[327] vdd gnd cell_6t
Xbit_r328_c66 bl[66] br[66] wl[328] vdd gnd cell_6t
Xbit_r329_c66 bl[66] br[66] wl[329] vdd gnd cell_6t
Xbit_r330_c66 bl[66] br[66] wl[330] vdd gnd cell_6t
Xbit_r331_c66 bl[66] br[66] wl[331] vdd gnd cell_6t
Xbit_r332_c66 bl[66] br[66] wl[332] vdd gnd cell_6t
Xbit_r333_c66 bl[66] br[66] wl[333] vdd gnd cell_6t
Xbit_r334_c66 bl[66] br[66] wl[334] vdd gnd cell_6t
Xbit_r335_c66 bl[66] br[66] wl[335] vdd gnd cell_6t
Xbit_r336_c66 bl[66] br[66] wl[336] vdd gnd cell_6t
Xbit_r337_c66 bl[66] br[66] wl[337] vdd gnd cell_6t
Xbit_r338_c66 bl[66] br[66] wl[338] vdd gnd cell_6t
Xbit_r339_c66 bl[66] br[66] wl[339] vdd gnd cell_6t
Xbit_r340_c66 bl[66] br[66] wl[340] vdd gnd cell_6t
Xbit_r341_c66 bl[66] br[66] wl[341] vdd gnd cell_6t
Xbit_r342_c66 bl[66] br[66] wl[342] vdd gnd cell_6t
Xbit_r343_c66 bl[66] br[66] wl[343] vdd gnd cell_6t
Xbit_r344_c66 bl[66] br[66] wl[344] vdd gnd cell_6t
Xbit_r345_c66 bl[66] br[66] wl[345] vdd gnd cell_6t
Xbit_r346_c66 bl[66] br[66] wl[346] vdd gnd cell_6t
Xbit_r347_c66 bl[66] br[66] wl[347] vdd gnd cell_6t
Xbit_r348_c66 bl[66] br[66] wl[348] vdd gnd cell_6t
Xbit_r349_c66 bl[66] br[66] wl[349] vdd gnd cell_6t
Xbit_r350_c66 bl[66] br[66] wl[350] vdd gnd cell_6t
Xbit_r351_c66 bl[66] br[66] wl[351] vdd gnd cell_6t
Xbit_r352_c66 bl[66] br[66] wl[352] vdd gnd cell_6t
Xbit_r353_c66 bl[66] br[66] wl[353] vdd gnd cell_6t
Xbit_r354_c66 bl[66] br[66] wl[354] vdd gnd cell_6t
Xbit_r355_c66 bl[66] br[66] wl[355] vdd gnd cell_6t
Xbit_r356_c66 bl[66] br[66] wl[356] vdd gnd cell_6t
Xbit_r357_c66 bl[66] br[66] wl[357] vdd gnd cell_6t
Xbit_r358_c66 bl[66] br[66] wl[358] vdd gnd cell_6t
Xbit_r359_c66 bl[66] br[66] wl[359] vdd gnd cell_6t
Xbit_r360_c66 bl[66] br[66] wl[360] vdd gnd cell_6t
Xbit_r361_c66 bl[66] br[66] wl[361] vdd gnd cell_6t
Xbit_r362_c66 bl[66] br[66] wl[362] vdd gnd cell_6t
Xbit_r363_c66 bl[66] br[66] wl[363] vdd gnd cell_6t
Xbit_r364_c66 bl[66] br[66] wl[364] vdd gnd cell_6t
Xbit_r365_c66 bl[66] br[66] wl[365] vdd gnd cell_6t
Xbit_r366_c66 bl[66] br[66] wl[366] vdd gnd cell_6t
Xbit_r367_c66 bl[66] br[66] wl[367] vdd gnd cell_6t
Xbit_r368_c66 bl[66] br[66] wl[368] vdd gnd cell_6t
Xbit_r369_c66 bl[66] br[66] wl[369] vdd gnd cell_6t
Xbit_r370_c66 bl[66] br[66] wl[370] vdd gnd cell_6t
Xbit_r371_c66 bl[66] br[66] wl[371] vdd gnd cell_6t
Xbit_r372_c66 bl[66] br[66] wl[372] vdd gnd cell_6t
Xbit_r373_c66 bl[66] br[66] wl[373] vdd gnd cell_6t
Xbit_r374_c66 bl[66] br[66] wl[374] vdd gnd cell_6t
Xbit_r375_c66 bl[66] br[66] wl[375] vdd gnd cell_6t
Xbit_r376_c66 bl[66] br[66] wl[376] vdd gnd cell_6t
Xbit_r377_c66 bl[66] br[66] wl[377] vdd gnd cell_6t
Xbit_r378_c66 bl[66] br[66] wl[378] vdd gnd cell_6t
Xbit_r379_c66 bl[66] br[66] wl[379] vdd gnd cell_6t
Xbit_r380_c66 bl[66] br[66] wl[380] vdd gnd cell_6t
Xbit_r381_c66 bl[66] br[66] wl[381] vdd gnd cell_6t
Xbit_r382_c66 bl[66] br[66] wl[382] vdd gnd cell_6t
Xbit_r383_c66 bl[66] br[66] wl[383] vdd gnd cell_6t
Xbit_r384_c66 bl[66] br[66] wl[384] vdd gnd cell_6t
Xbit_r385_c66 bl[66] br[66] wl[385] vdd gnd cell_6t
Xbit_r386_c66 bl[66] br[66] wl[386] vdd gnd cell_6t
Xbit_r387_c66 bl[66] br[66] wl[387] vdd gnd cell_6t
Xbit_r388_c66 bl[66] br[66] wl[388] vdd gnd cell_6t
Xbit_r389_c66 bl[66] br[66] wl[389] vdd gnd cell_6t
Xbit_r390_c66 bl[66] br[66] wl[390] vdd gnd cell_6t
Xbit_r391_c66 bl[66] br[66] wl[391] vdd gnd cell_6t
Xbit_r392_c66 bl[66] br[66] wl[392] vdd gnd cell_6t
Xbit_r393_c66 bl[66] br[66] wl[393] vdd gnd cell_6t
Xbit_r394_c66 bl[66] br[66] wl[394] vdd gnd cell_6t
Xbit_r395_c66 bl[66] br[66] wl[395] vdd gnd cell_6t
Xbit_r396_c66 bl[66] br[66] wl[396] vdd gnd cell_6t
Xbit_r397_c66 bl[66] br[66] wl[397] vdd gnd cell_6t
Xbit_r398_c66 bl[66] br[66] wl[398] vdd gnd cell_6t
Xbit_r399_c66 bl[66] br[66] wl[399] vdd gnd cell_6t
Xbit_r400_c66 bl[66] br[66] wl[400] vdd gnd cell_6t
Xbit_r401_c66 bl[66] br[66] wl[401] vdd gnd cell_6t
Xbit_r402_c66 bl[66] br[66] wl[402] vdd gnd cell_6t
Xbit_r403_c66 bl[66] br[66] wl[403] vdd gnd cell_6t
Xbit_r404_c66 bl[66] br[66] wl[404] vdd gnd cell_6t
Xbit_r405_c66 bl[66] br[66] wl[405] vdd gnd cell_6t
Xbit_r406_c66 bl[66] br[66] wl[406] vdd gnd cell_6t
Xbit_r407_c66 bl[66] br[66] wl[407] vdd gnd cell_6t
Xbit_r408_c66 bl[66] br[66] wl[408] vdd gnd cell_6t
Xbit_r409_c66 bl[66] br[66] wl[409] vdd gnd cell_6t
Xbit_r410_c66 bl[66] br[66] wl[410] vdd gnd cell_6t
Xbit_r411_c66 bl[66] br[66] wl[411] vdd gnd cell_6t
Xbit_r412_c66 bl[66] br[66] wl[412] vdd gnd cell_6t
Xbit_r413_c66 bl[66] br[66] wl[413] vdd gnd cell_6t
Xbit_r414_c66 bl[66] br[66] wl[414] vdd gnd cell_6t
Xbit_r415_c66 bl[66] br[66] wl[415] vdd gnd cell_6t
Xbit_r416_c66 bl[66] br[66] wl[416] vdd gnd cell_6t
Xbit_r417_c66 bl[66] br[66] wl[417] vdd gnd cell_6t
Xbit_r418_c66 bl[66] br[66] wl[418] vdd gnd cell_6t
Xbit_r419_c66 bl[66] br[66] wl[419] vdd gnd cell_6t
Xbit_r420_c66 bl[66] br[66] wl[420] vdd gnd cell_6t
Xbit_r421_c66 bl[66] br[66] wl[421] vdd gnd cell_6t
Xbit_r422_c66 bl[66] br[66] wl[422] vdd gnd cell_6t
Xbit_r423_c66 bl[66] br[66] wl[423] vdd gnd cell_6t
Xbit_r424_c66 bl[66] br[66] wl[424] vdd gnd cell_6t
Xbit_r425_c66 bl[66] br[66] wl[425] vdd gnd cell_6t
Xbit_r426_c66 bl[66] br[66] wl[426] vdd gnd cell_6t
Xbit_r427_c66 bl[66] br[66] wl[427] vdd gnd cell_6t
Xbit_r428_c66 bl[66] br[66] wl[428] vdd gnd cell_6t
Xbit_r429_c66 bl[66] br[66] wl[429] vdd gnd cell_6t
Xbit_r430_c66 bl[66] br[66] wl[430] vdd gnd cell_6t
Xbit_r431_c66 bl[66] br[66] wl[431] vdd gnd cell_6t
Xbit_r432_c66 bl[66] br[66] wl[432] vdd gnd cell_6t
Xbit_r433_c66 bl[66] br[66] wl[433] vdd gnd cell_6t
Xbit_r434_c66 bl[66] br[66] wl[434] vdd gnd cell_6t
Xbit_r435_c66 bl[66] br[66] wl[435] vdd gnd cell_6t
Xbit_r436_c66 bl[66] br[66] wl[436] vdd gnd cell_6t
Xbit_r437_c66 bl[66] br[66] wl[437] vdd gnd cell_6t
Xbit_r438_c66 bl[66] br[66] wl[438] vdd gnd cell_6t
Xbit_r439_c66 bl[66] br[66] wl[439] vdd gnd cell_6t
Xbit_r440_c66 bl[66] br[66] wl[440] vdd gnd cell_6t
Xbit_r441_c66 bl[66] br[66] wl[441] vdd gnd cell_6t
Xbit_r442_c66 bl[66] br[66] wl[442] vdd gnd cell_6t
Xbit_r443_c66 bl[66] br[66] wl[443] vdd gnd cell_6t
Xbit_r444_c66 bl[66] br[66] wl[444] vdd gnd cell_6t
Xbit_r445_c66 bl[66] br[66] wl[445] vdd gnd cell_6t
Xbit_r446_c66 bl[66] br[66] wl[446] vdd gnd cell_6t
Xbit_r447_c66 bl[66] br[66] wl[447] vdd gnd cell_6t
Xbit_r448_c66 bl[66] br[66] wl[448] vdd gnd cell_6t
Xbit_r449_c66 bl[66] br[66] wl[449] vdd gnd cell_6t
Xbit_r450_c66 bl[66] br[66] wl[450] vdd gnd cell_6t
Xbit_r451_c66 bl[66] br[66] wl[451] vdd gnd cell_6t
Xbit_r452_c66 bl[66] br[66] wl[452] vdd gnd cell_6t
Xbit_r453_c66 bl[66] br[66] wl[453] vdd gnd cell_6t
Xbit_r454_c66 bl[66] br[66] wl[454] vdd gnd cell_6t
Xbit_r455_c66 bl[66] br[66] wl[455] vdd gnd cell_6t
Xbit_r456_c66 bl[66] br[66] wl[456] vdd gnd cell_6t
Xbit_r457_c66 bl[66] br[66] wl[457] vdd gnd cell_6t
Xbit_r458_c66 bl[66] br[66] wl[458] vdd gnd cell_6t
Xbit_r459_c66 bl[66] br[66] wl[459] vdd gnd cell_6t
Xbit_r460_c66 bl[66] br[66] wl[460] vdd gnd cell_6t
Xbit_r461_c66 bl[66] br[66] wl[461] vdd gnd cell_6t
Xbit_r462_c66 bl[66] br[66] wl[462] vdd gnd cell_6t
Xbit_r463_c66 bl[66] br[66] wl[463] vdd gnd cell_6t
Xbit_r464_c66 bl[66] br[66] wl[464] vdd gnd cell_6t
Xbit_r465_c66 bl[66] br[66] wl[465] vdd gnd cell_6t
Xbit_r466_c66 bl[66] br[66] wl[466] vdd gnd cell_6t
Xbit_r467_c66 bl[66] br[66] wl[467] vdd gnd cell_6t
Xbit_r468_c66 bl[66] br[66] wl[468] vdd gnd cell_6t
Xbit_r469_c66 bl[66] br[66] wl[469] vdd gnd cell_6t
Xbit_r470_c66 bl[66] br[66] wl[470] vdd gnd cell_6t
Xbit_r471_c66 bl[66] br[66] wl[471] vdd gnd cell_6t
Xbit_r472_c66 bl[66] br[66] wl[472] vdd gnd cell_6t
Xbit_r473_c66 bl[66] br[66] wl[473] vdd gnd cell_6t
Xbit_r474_c66 bl[66] br[66] wl[474] vdd gnd cell_6t
Xbit_r475_c66 bl[66] br[66] wl[475] vdd gnd cell_6t
Xbit_r476_c66 bl[66] br[66] wl[476] vdd gnd cell_6t
Xbit_r477_c66 bl[66] br[66] wl[477] vdd gnd cell_6t
Xbit_r478_c66 bl[66] br[66] wl[478] vdd gnd cell_6t
Xbit_r479_c66 bl[66] br[66] wl[479] vdd gnd cell_6t
Xbit_r480_c66 bl[66] br[66] wl[480] vdd gnd cell_6t
Xbit_r481_c66 bl[66] br[66] wl[481] vdd gnd cell_6t
Xbit_r482_c66 bl[66] br[66] wl[482] vdd gnd cell_6t
Xbit_r483_c66 bl[66] br[66] wl[483] vdd gnd cell_6t
Xbit_r484_c66 bl[66] br[66] wl[484] vdd gnd cell_6t
Xbit_r485_c66 bl[66] br[66] wl[485] vdd gnd cell_6t
Xbit_r486_c66 bl[66] br[66] wl[486] vdd gnd cell_6t
Xbit_r487_c66 bl[66] br[66] wl[487] vdd gnd cell_6t
Xbit_r488_c66 bl[66] br[66] wl[488] vdd gnd cell_6t
Xbit_r489_c66 bl[66] br[66] wl[489] vdd gnd cell_6t
Xbit_r490_c66 bl[66] br[66] wl[490] vdd gnd cell_6t
Xbit_r491_c66 bl[66] br[66] wl[491] vdd gnd cell_6t
Xbit_r492_c66 bl[66] br[66] wl[492] vdd gnd cell_6t
Xbit_r493_c66 bl[66] br[66] wl[493] vdd gnd cell_6t
Xbit_r494_c66 bl[66] br[66] wl[494] vdd gnd cell_6t
Xbit_r495_c66 bl[66] br[66] wl[495] vdd gnd cell_6t
Xbit_r496_c66 bl[66] br[66] wl[496] vdd gnd cell_6t
Xbit_r497_c66 bl[66] br[66] wl[497] vdd gnd cell_6t
Xbit_r498_c66 bl[66] br[66] wl[498] vdd gnd cell_6t
Xbit_r499_c66 bl[66] br[66] wl[499] vdd gnd cell_6t
Xbit_r500_c66 bl[66] br[66] wl[500] vdd gnd cell_6t
Xbit_r501_c66 bl[66] br[66] wl[501] vdd gnd cell_6t
Xbit_r502_c66 bl[66] br[66] wl[502] vdd gnd cell_6t
Xbit_r503_c66 bl[66] br[66] wl[503] vdd gnd cell_6t
Xbit_r504_c66 bl[66] br[66] wl[504] vdd gnd cell_6t
Xbit_r505_c66 bl[66] br[66] wl[505] vdd gnd cell_6t
Xbit_r506_c66 bl[66] br[66] wl[506] vdd gnd cell_6t
Xbit_r507_c66 bl[66] br[66] wl[507] vdd gnd cell_6t
Xbit_r508_c66 bl[66] br[66] wl[508] vdd gnd cell_6t
Xbit_r509_c66 bl[66] br[66] wl[509] vdd gnd cell_6t
Xbit_r510_c66 bl[66] br[66] wl[510] vdd gnd cell_6t
Xbit_r511_c66 bl[66] br[66] wl[511] vdd gnd cell_6t
Xbit_r0_c67 bl[67] br[67] wl[0] vdd gnd cell_6t
Xbit_r1_c67 bl[67] br[67] wl[1] vdd gnd cell_6t
Xbit_r2_c67 bl[67] br[67] wl[2] vdd gnd cell_6t
Xbit_r3_c67 bl[67] br[67] wl[3] vdd gnd cell_6t
Xbit_r4_c67 bl[67] br[67] wl[4] vdd gnd cell_6t
Xbit_r5_c67 bl[67] br[67] wl[5] vdd gnd cell_6t
Xbit_r6_c67 bl[67] br[67] wl[6] vdd gnd cell_6t
Xbit_r7_c67 bl[67] br[67] wl[7] vdd gnd cell_6t
Xbit_r8_c67 bl[67] br[67] wl[8] vdd gnd cell_6t
Xbit_r9_c67 bl[67] br[67] wl[9] vdd gnd cell_6t
Xbit_r10_c67 bl[67] br[67] wl[10] vdd gnd cell_6t
Xbit_r11_c67 bl[67] br[67] wl[11] vdd gnd cell_6t
Xbit_r12_c67 bl[67] br[67] wl[12] vdd gnd cell_6t
Xbit_r13_c67 bl[67] br[67] wl[13] vdd gnd cell_6t
Xbit_r14_c67 bl[67] br[67] wl[14] vdd gnd cell_6t
Xbit_r15_c67 bl[67] br[67] wl[15] vdd gnd cell_6t
Xbit_r16_c67 bl[67] br[67] wl[16] vdd gnd cell_6t
Xbit_r17_c67 bl[67] br[67] wl[17] vdd gnd cell_6t
Xbit_r18_c67 bl[67] br[67] wl[18] vdd gnd cell_6t
Xbit_r19_c67 bl[67] br[67] wl[19] vdd gnd cell_6t
Xbit_r20_c67 bl[67] br[67] wl[20] vdd gnd cell_6t
Xbit_r21_c67 bl[67] br[67] wl[21] vdd gnd cell_6t
Xbit_r22_c67 bl[67] br[67] wl[22] vdd gnd cell_6t
Xbit_r23_c67 bl[67] br[67] wl[23] vdd gnd cell_6t
Xbit_r24_c67 bl[67] br[67] wl[24] vdd gnd cell_6t
Xbit_r25_c67 bl[67] br[67] wl[25] vdd gnd cell_6t
Xbit_r26_c67 bl[67] br[67] wl[26] vdd gnd cell_6t
Xbit_r27_c67 bl[67] br[67] wl[27] vdd gnd cell_6t
Xbit_r28_c67 bl[67] br[67] wl[28] vdd gnd cell_6t
Xbit_r29_c67 bl[67] br[67] wl[29] vdd gnd cell_6t
Xbit_r30_c67 bl[67] br[67] wl[30] vdd gnd cell_6t
Xbit_r31_c67 bl[67] br[67] wl[31] vdd gnd cell_6t
Xbit_r32_c67 bl[67] br[67] wl[32] vdd gnd cell_6t
Xbit_r33_c67 bl[67] br[67] wl[33] vdd gnd cell_6t
Xbit_r34_c67 bl[67] br[67] wl[34] vdd gnd cell_6t
Xbit_r35_c67 bl[67] br[67] wl[35] vdd gnd cell_6t
Xbit_r36_c67 bl[67] br[67] wl[36] vdd gnd cell_6t
Xbit_r37_c67 bl[67] br[67] wl[37] vdd gnd cell_6t
Xbit_r38_c67 bl[67] br[67] wl[38] vdd gnd cell_6t
Xbit_r39_c67 bl[67] br[67] wl[39] vdd gnd cell_6t
Xbit_r40_c67 bl[67] br[67] wl[40] vdd gnd cell_6t
Xbit_r41_c67 bl[67] br[67] wl[41] vdd gnd cell_6t
Xbit_r42_c67 bl[67] br[67] wl[42] vdd gnd cell_6t
Xbit_r43_c67 bl[67] br[67] wl[43] vdd gnd cell_6t
Xbit_r44_c67 bl[67] br[67] wl[44] vdd gnd cell_6t
Xbit_r45_c67 bl[67] br[67] wl[45] vdd gnd cell_6t
Xbit_r46_c67 bl[67] br[67] wl[46] vdd gnd cell_6t
Xbit_r47_c67 bl[67] br[67] wl[47] vdd gnd cell_6t
Xbit_r48_c67 bl[67] br[67] wl[48] vdd gnd cell_6t
Xbit_r49_c67 bl[67] br[67] wl[49] vdd gnd cell_6t
Xbit_r50_c67 bl[67] br[67] wl[50] vdd gnd cell_6t
Xbit_r51_c67 bl[67] br[67] wl[51] vdd gnd cell_6t
Xbit_r52_c67 bl[67] br[67] wl[52] vdd gnd cell_6t
Xbit_r53_c67 bl[67] br[67] wl[53] vdd gnd cell_6t
Xbit_r54_c67 bl[67] br[67] wl[54] vdd gnd cell_6t
Xbit_r55_c67 bl[67] br[67] wl[55] vdd gnd cell_6t
Xbit_r56_c67 bl[67] br[67] wl[56] vdd gnd cell_6t
Xbit_r57_c67 bl[67] br[67] wl[57] vdd gnd cell_6t
Xbit_r58_c67 bl[67] br[67] wl[58] vdd gnd cell_6t
Xbit_r59_c67 bl[67] br[67] wl[59] vdd gnd cell_6t
Xbit_r60_c67 bl[67] br[67] wl[60] vdd gnd cell_6t
Xbit_r61_c67 bl[67] br[67] wl[61] vdd gnd cell_6t
Xbit_r62_c67 bl[67] br[67] wl[62] vdd gnd cell_6t
Xbit_r63_c67 bl[67] br[67] wl[63] vdd gnd cell_6t
Xbit_r64_c67 bl[67] br[67] wl[64] vdd gnd cell_6t
Xbit_r65_c67 bl[67] br[67] wl[65] vdd gnd cell_6t
Xbit_r66_c67 bl[67] br[67] wl[66] vdd gnd cell_6t
Xbit_r67_c67 bl[67] br[67] wl[67] vdd gnd cell_6t
Xbit_r68_c67 bl[67] br[67] wl[68] vdd gnd cell_6t
Xbit_r69_c67 bl[67] br[67] wl[69] vdd gnd cell_6t
Xbit_r70_c67 bl[67] br[67] wl[70] vdd gnd cell_6t
Xbit_r71_c67 bl[67] br[67] wl[71] vdd gnd cell_6t
Xbit_r72_c67 bl[67] br[67] wl[72] vdd gnd cell_6t
Xbit_r73_c67 bl[67] br[67] wl[73] vdd gnd cell_6t
Xbit_r74_c67 bl[67] br[67] wl[74] vdd gnd cell_6t
Xbit_r75_c67 bl[67] br[67] wl[75] vdd gnd cell_6t
Xbit_r76_c67 bl[67] br[67] wl[76] vdd gnd cell_6t
Xbit_r77_c67 bl[67] br[67] wl[77] vdd gnd cell_6t
Xbit_r78_c67 bl[67] br[67] wl[78] vdd gnd cell_6t
Xbit_r79_c67 bl[67] br[67] wl[79] vdd gnd cell_6t
Xbit_r80_c67 bl[67] br[67] wl[80] vdd gnd cell_6t
Xbit_r81_c67 bl[67] br[67] wl[81] vdd gnd cell_6t
Xbit_r82_c67 bl[67] br[67] wl[82] vdd gnd cell_6t
Xbit_r83_c67 bl[67] br[67] wl[83] vdd gnd cell_6t
Xbit_r84_c67 bl[67] br[67] wl[84] vdd gnd cell_6t
Xbit_r85_c67 bl[67] br[67] wl[85] vdd gnd cell_6t
Xbit_r86_c67 bl[67] br[67] wl[86] vdd gnd cell_6t
Xbit_r87_c67 bl[67] br[67] wl[87] vdd gnd cell_6t
Xbit_r88_c67 bl[67] br[67] wl[88] vdd gnd cell_6t
Xbit_r89_c67 bl[67] br[67] wl[89] vdd gnd cell_6t
Xbit_r90_c67 bl[67] br[67] wl[90] vdd gnd cell_6t
Xbit_r91_c67 bl[67] br[67] wl[91] vdd gnd cell_6t
Xbit_r92_c67 bl[67] br[67] wl[92] vdd gnd cell_6t
Xbit_r93_c67 bl[67] br[67] wl[93] vdd gnd cell_6t
Xbit_r94_c67 bl[67] br[67] wl[94] vdd gnd cell_6t
Xbit_r95_c67 bl[67] br[67] wl[95] vdd gnd cell_6t
Xbit_r96_c67 bl[67] br[67] wl[96] vdd gnd cell_6t
Xbit_r97_c67 bl[67] br[67] wl[97] vdd gnd cell_6t
Xbit_r98_c67 bl[67] br[67] wl[98] vdd gnd cell_6t
Xbit_r99_c67 bl[67] br[67] wl[99] vdd gnd cell_6t
Xbit_r100_c67 bl[67] br[67] wl[100] vdd gnd cell_6t
Xbit_r101_c67 bl[67] br[67] wl[101] vdd gnd cell_6t
Xbit_r102_c67 bl[67] br[67] wl[102] vdd gnd cell_6t
Xbit_r103_c67 bl[67] br[67] wl[103] vdd gnd cell_6t
Xbit_r104_c67 bl[67] br[67] wl[104] vdd gnd cell_6t
Xbit_r105_c67 bl[67] br[67] wl[105] vdd gnd cell_6t
Xbit_r106_c67 bl[67] br[67] wl[106] vdd gnd cell_6t
Xbit_r107_c67 bl[67] br[67] wl[107] vdd gnd cell_6t
Xbit_r108_c67 bl[67] br[67] wl[108] vdd gnd cell_6t
Xbit_r109_c67 bl[67] br[67] wl[109] vdd gnd cell_6t
Xbit_r110_c67 bl[67] br[67] wl[110] vdd gnd cell_6t
Xbit_r111_c67 bl[67] br[67] wl[111] vdd gnd cell_6t
Xbit_r112_c67 bl[67] br[67] wl[112] vdd gnd cell_6t
Xbit_r113_c67 bl[67] br[67] wl[113] vdd gnd cell_6t
Xbit_r114_c67 bl[67] br[67] wl[114] vdd gnd cell_6t
Xbit_r115_c67 bl[67] br[67] wl[115] vdd gnd cell_6t
Xbit_r116_c67 bl[67] br[67] wl[116] vdd gnd cell_6t
Xbit_r117_c67 bl[67] br[67] wl[117] vdd gnd cell_6t
Xbit_r118_c67 bl[67] br[67] wl[118] vdd gnd cell_6t
Xbit_r119_c67 bl[67] br[67] wl[119] vdd gnd cell_6t
Xbit_r120_c67 bl[67] br[67] wl[120] vdd gnd cell_6t
Xbit_r121_c67 bl[67] br[67] wl[121] vdd gnd cell_6t
Xbit_r122_c67 bl[67] br[67] wl[122] vdd gnd cell_6t
Xbit_r123_c67 bl[67] br[67] wl[123] vdd gnd cell_6t
Xbit_r124_c67 bl[67] br[67] wl[124] vdd gnd cell_6t
Xbit_r125_c67 bl[67] br[67] wl[125] vdd gnd cell_6t
Xbit_r126_c67 bl[67] br[67] wl[126] vdd gnd cell_6t
Xbit_r127_c67 bl[67] br[67] wl[127] vdd gnd cell_6t
Xbit_r128_c67 bl[67] br[67] wl[128] vdd gnd cell_6t
Xbit_r129_c67 bl[67] br[67] wl[129] vdd gnd cell_6t
Xbit_r130_c67 bl[67] br[67] wl[130] vdd gnd cell_6t
Xbit_r131_c67 bl[67] br[67] wl[131] vdd gnd cell_6t
Xbit_r132_c67 bl[67] br[67] wl[132] vdd gnd cell_6t
Xbit_r133_c67 bl[67] br[67] wl[133] vdd gnd cell_6t
Xbit_r134_c67 bl[67] br[67] wl[134] vdd gnd cell_6t
Xbit_r135_c67 bl[67] br[67] wl[135] vdd gnd cell_6t
Xbit_r136_c67 bl[67] br[67] wl[136] vdd gnd cell_6t
Xbit_r137_c67 bl[67] br[67] wl[137] vdd gnd cell_6t
Xbit_r138_c67 bl[67] br[67] wl[138] vdd gnd cell_6t
Xbit_r139_c67 bl[67] br[67] wl[139] vdd gnd cell_6t
Xbit_r140_c67 bl[67] br[67] wl[140] vdd gnd cell_6t
Xbit_r141_c67 bl[67] br[67] wl[141] vdd gnd cell_6t
Xbit_r142_c67 bl[67] br[67] wl[142] vdd gnd cell_6t
Xbit_r143_c67 bl[67] br[67] wl[143] vdd gnd cell_6t
Xbit_r144_c67 bl[67] br[67] wl[144] vdd gnd cell_6t
Xbit_r145_c67 bl[67] br[67] wl[145] vdd gnd cell_6t
Xbit_r146_c67 bl[67] br[67] wl[146] vdd gnd cell_6t
Xbit_r147_c67 bl[67] br[67] wl[147] vdd gnd cell_6t
Xbit_r148_c67 bl[67] br[67] wl[148] vdd gnd cell_6t
Xbit_r149_c67 bl[67] br[67] wl[149] vdd gnd cell_6t
Xbit_r150_c67 bl[67] br[67] wl[150] vdd gnd cell_6t
Xbit_r151_c67 bl[67] br[67] wl[151] vdd gnd cell_6t
Xbit_r152_c67 bl[67] br[67] wl[152] vdd gnd cell_6t
Xbit_r153_c67 bl[67] br[67] wl[153] vdd gnd cell_6t
Xbit_r154_c67 bl[67] br[67] wl[154] vdd gnd cell_6t
Xbit_r155_c67 bl[67] br[67] wl[155] vdd gnd cell_6t
Xbit_r156_c67 bl[67] br[67] wl[156] vdd gnd cell_6t
Xbit_r157_c67 bl[67] br[67] wl[157] vdd gnd cell_6t
Xbit_r158_c67 bl[67] br[67] wl[158] vdd gnd cell_6t
Xbit_r159_c67 bl[67] br[67] wl[159] vdd gnd cell_6t
Xbit_r160_c67 bl[67] br[67] wl[160] vdd gnd cell_6t
Xbit_r161_c67 bl[67] br[67] wl[161] vdd gnd cell_6t
Xbit_r162_c67 bl[67] br[67] wl[162] vdd gnd cell_6t
Xbit_r163_c67 bl[67] br[67] wl[163] vdd gnd cell_6t
Xbit_r164_c67 bl[67] br[67] wl[164] vdd gnd cell_6t
Xbit_r165_c67 bl[67] br[67] wl[165] vdd gnd cell_6t
Xbit_r166_c67 bl[67] br[67] wl[166] vdd gnd cell_6t
Xbit_r167_c67 bl[67] br[67] wl[167] vdd gnd cell_6t
Xbit_r168_c67 bl[67] br[67] wl[168] vdd gnd cell_6t
Xbit_r169_c67 bl[67] br[67] wl[169] vdd gnd cell_6t
Xbit_r170_c67 bl[67] br[67] wl[170] vdd gnd cell_6t
Xbit_r171_c67 bl[67] br[67] wl[171] vdd gnd cell_6t
Xbit_r172_c67 bl[67] br[67] wl[172] vdd gnd cell_6t
Xbit_r173_c67 bl[67] br[67] wl[173] vdd gnd cell_6t
Xbit_r174_c67 bl[67] br[67] wl[174] vdd gnd cell_6t
Xbit_r175_c67 bl[67] br[67] wl[175] vdd gnd cell_6t
Xbit_r176_c67 bl[67] br[67] wl[176] vdd gnd cell_6t
Xbit_r177_c67 bl[67] br[67] wl[177] vdd gnd cell_6t
Xbit_r178_c67 bl[67] br[67] wl[178] vdd gnd cell_6t
Xbit_r179_c67 bl[67] br[67] wl[179] vdd gnd cell_6t
Xbit_r180_c67 bl[67] br[67] wl[180] vdd gnd cell_6t
Xbit_r181_c67 bl[67] br[67] wl[181] vdd gnd cell_6t
Xbit_r182_c67 bl[67] br[67] wl[182] vdd gnd cell_6t
Xbit_r183_c67 bl[67] br[67] wl[183] vdd gnd cell_6t
Xbit_r184_c67 bl[67] br[67] wl[184] vdd gnd cell_6t
Xbit_r185_c67 bl[67] br[67] wl[185] vdd gnd cell_6t
Xbit_r186_c67 bl[67] br[67] wl[186] vdd gnd cell_6t
Xbit_r187_c67 bl[67] br[67] wl[187] vdd gnd cell_6t
Xbit_r188_c67 bl[67] br[67] wl[188] vdd gnd cell_6t
Xbit_r189_c67 bl[67] br[67] wl[189] vdd gnd cell_6t
Xbit_r190_c67 bl[67] br[67] wl[190] vdd gnd cell_6t
Xbit_r191_c67 bl[67] br[67] wl[191] vdd gnd cell_6t
Xbit_r192_c67 bl[67] br[67] wl[192] vdd gnd cell_6t
Xbit_r193_c67 bl[67] br[67] wl[193] vdd gnd cell_6t
Xbit_r194_c67 bl[67] br[67] wl[194] vdd gnd cell_6t
Xbit_r195_c67 bl[67] br[67] wl[195] vdd gnd cell_6t
Xbit_r196_c67 bl[67] br[67] wl[196] vdd gnd cell_6t
Xbit_r197_c67 bl[67] br[67] wl[197] vdd gnd cell_6t
Xbit_r198_c67 bl[67] br[67] wl[198] vdd gnd cell_6t
Xbit_r199_c67 bl[67] br[67] wl[199] vdd gnd cell_6t
Xbit_r200_c67 bl[67] br[67] wl[200] vdd gnd cell_6t
Xbit_r201_c67 bl[67] br[67] wl[201] vdd gnd cell_6t
Xbit_r202_c67 bl[67] br[67] wl[202] vdd gnd cell_6t
Xbit_r203_c67 bl[67] br[67] wl[203] vdd gnd cell_6t
Xbit_r204_c67 bl[67] br[67] wl[204] vdd gnd cell_6t
Xbit_r205_c67 bl[67] br[67] wl[205] vdd gnd cell_6t
Xbit_r206_c67 bl[67] br[67] wl[206] vdd gnd cell_6t
Xbit_r207_c67 bl[67] br[67] wl[207] vdd gnd cell_6t
Xbit_r208_c67 bl[67] br[67] wl[208] vdd gnd cell_6t
Xbit_r209_c67 bl[67] br[67] wl[209] vdd gnd cell_6t
Xbit_r210_c67 bl[67] br[67] wl[210] vdd gnd cell_6t
Xbit_r211_c67 bl[67] br[67] wl[211] vdd gnd cell_6t
Xbit_r212_c67 bl[67] br[67] wl[212] vdd gnd cell_6t
Xbit_r213_c67 bl[67] br[67] wl[213] vdd gnd cell_6t
Xbit_r214_c67 bl[67] br[67] wl[214] vdd gnd cell_6t
Xbit_r215_c67 bl[67] br[67] wl[215] vdd gnd cell_6t
Xbit_r216_c67 bl[67] br[67] wl[216] vdd gnd cell_6t
Xbit_r217_c67 bl[67] br[67] wl[217] vdd gnd cell_6t
Xbit_r218_c67 bl[67] br[67] wl[218] vdd gnd cell_6t
Xbit_r219_c67 bl[67] br[67] wl[219] vdd gnd cell_6t
Xbit_r220_c67 bl[67] br[67] wl[220] vdd gnd cell_6t
Xbit_r221_c67 bl[67] br[67] wl[221] vdd gnd cell_6t
Xbit_r222_c67 bl[67] br[67] wl[222] vdd gnd cell_6t
Xbit_r223_c67 bl[67] br[67] wl[223] vdd gnd cell_6t
Xbit_r224_c67 bl[67] br[67] wl[224] vdd gnd cell_6t
Xbit_r225_c67 bl[67] br[67] wl[225] vdd gnd cell_6t
Xbit_r226_c67 bl[67] br[67] wl[226] vdd gnd cell_6t
Xbit_r227_c67 bl[67] br[67] wl[227] vdd gnd cell_6t
Xbit_r228_c67 bl[67] br[67] wl[228] vdd gnd cell_6t
Xbit_r229_c67 bl[67] br[67] wl[229] vdd gnd cell_6t
Xbit_r230_c67 bl[67] br[67] wl[230] vdd gnd cell_6t
Xbit_r231_c67 bl[67] br[67] wl[231] vdd gnd cell_6t
Xbit_r232_c67 bl[67] br[67] wl[232] vdd gnd cell_6t
Xbit_r233_c67 bl[67] br[67] wl[233] vdd gnd cell_6t
Xbit_r234_c67 bl[67] br[67] wl[234] vdd gnd cell_6t
Xbit_r235_c67 bl[67] br[67] wl[235] vdd gnd cell_6t
Xbit_r236_c67 bl[67] br[67] wl[236] vdd gnd cell_6t
Xbit_r237_c67 bl[67] br[67] wl[237] vdd gnd cell_6t
Xbit_r238_c67 bl[67] br[67] wl[238] vdd gnd cell_6t
Xbit_r239_c67 bl[67] br[67] wl[239] vdd gnd cell_6t
Xbit_r240_c67 bl[67] br[67] wl[240] vdd gnd cell_6t
Xbit_r241_c67 bl[67] br[67] wl[241] vdd gnd cell_6t
Xbit_r242_c67 bl[67] br[67] wl[242] vdd gnd cell_6t
Xbit_r243_c67 bl[67] br[67] wl[243] vdd gnd cell_6t
Xbit_r244_c67 bl[67] br[67] wl[244] vdd gnd cell_6t
Xbit_r245_c67 bl[67] br[67] wl[245] vdd gnd cell_6t
Xbit_r246_c67 bl[67] br[67] wl[246] vdd gnd cell_6t
Xbit_r247_c67 bl[67] br[67] wl[247] vdd gnd cell_6t
Xbit_r248_c67 bl[67] br[67] wl[248] vdd gnd cell_6t
Xbit_r249_c67 bl[67] br[67] wl[249] vdd gnd cell_6t
Xbit_r250_c67 bl[67] br[67] wl[250] vdd gnd cell_6t
Xbit_r251_c67 bl[67] br[67] wl[251] vdd gnd cell_6t
Xbit_r252_c67 bl[67] br[67] wl[252] vdd gnd cell_6t
Xbit_r253_c67 bl[67] br[67] wl[253] vdd gnd cell_6t
Xbit_r254_c67 bl[67] br[67] wl[254] vdd gnd cell_6t
Xbit_r255_c67 bl[67] br[67] wl[255] vdd gnd cell_6t
Xbit_r256_c67 bl[67] br[67] wl[256] vdd gnd cell_6t
Xbit_r257_c67 bl[67] br[67] wl[257] vdd gnd cell_6t
Xbit_r258_c67 bl[67] br[67] wl[258] vdd gnd cell_6t
Xbit_r259_c67 bl[67] br[67] wl[259] vdd gnd cell_6t
Xbit_r260_c67 bl[67] br[67] wl[260] vdd gnd cell_6t
Xbit_r261_c67 bl[67] br[67] wl[261] vdd gnd cell_6t
Xbit_r262_c67 bl[67] br[67] wl[262] vdd gnd cell_6t
Xbit_r263_c67 bl[67] br[67] wl[263] vdd gnd cell_6t
Xbit_r264_c67 bl[67] br[67] wl[264] vdd gnd cell_6t
Xbit_r265_c67 bl[67] br[67] wl[265] vdd gnd cell_6t
Xbit_r266_c67 bl[67] br[67] wl[266] vdd gnd cell_6t
Xbit_r267_c67 bl[67] br[67] wl[267] vdd gnd cell_6t
Xbit_r268_c67 bl[67] br[67] wl[268] vdd gnd cell_6t
Xbit_r269_c67 bl[67] br[67] wl[269] vdd gnd cell_6t
Xbit_r270_c67 bl[67] br[67] wl[270] vdd gnd cell_6t
Xbit_r271_c67 bl[67] br[67] wl[271] vdd gnd cell_6t
Xbit_r272_c67 bl[67] br[67] wl[272] vdd gnd cell_6t
Xbit_r273_c67 bl[67] br[67] wl[273] vdd gnd cell_6t
Xbit_r274_c67 bl[67] br[67] wl[274] vdd gnd cell_6t
Xbit_r275_c67 bl[67] br[67] wl[275] vdd gnd cell_6t
Xbit_r276_c67 bl[67] br[67] wl[276] vdd gnd cell_6t
Xbit_r277_c67 bl[67] br[67] wl[277] vdd gnd cell_6t
Xbit_r278_c67 bl[67] br[67] wl[278] vdd gnd cell_6t
Xbit_r279_c67 bl[67] br[67] wl[279] vdd gnd cell_6t
Xbit_r280_c67 bl[67] br[67] wl[280] vdd gnd cell_6t
Xbit_r281_c67 bl[67] br[67] wl[281] vdd gnd cell_6t
Xbit_r282_c67 bl[67] br[67] wl[282] vdd gnd cell_6t
Xbit_r283_c67 bl[67] br[67] wl[283] vdd gnd cell_6t
Xbit_r284_c67 bl[67] br[67] wl[284] vdd gnd cell_6t
Xbit_r285_c67 bl[67] br[67] wl[285] vdd gnd cell_6t
Xbit_r286_c67 bl[67] br[67] wl[286] vdd gnd cell_6t
Xbit_r287_c67 bl[67] br[67] wl[287] vdd gnd cell_6t
Xbit_r288_c67 bl[67] br[67] wl[288] vdd gnd cell_6t
Xbit_r289_c67 bl[67] br[67] wl[289] vdd gnd cell_6t
Xbit_r290_c67 bl[67] br[67] wl[290] vdd gnd cell_6t
Xbit_r291_c67 bl[67] br[67] wl[291] vdd gnd cell_6t
Xbit_r292_c67 bl[67] br[67] wl[292] vdd gnd cell_6t
Xbit_r293_c67 bl[67] br[67] wl[293] vdd gnd cell_6t
Xbit_r294_c67 bl[67] br[67] wl[294] vdd gnd cell_6t
Xbit_r295_c67 bl[67] br[67] wl[295] vdd gnd cell_6t
Xbit_r296_c67 bl[67] br[67] wl[296] vdd gnd cell_6t
Xbit_r297_c67 bl[67] br[67] wl[297] vdd gnd cell_6t
Xbit_r298_c67 bl[67] br[67] wl[298] vdd gnd cell_6t
Xbit_r299_c67 bl[67] br[67] wl[299] vdd gnd cell_6t
Xbit_r300_c67 bl[67] br[67] wl[300] vdd gnd cell_6t
Xbit_r301_c67 bl[67] br[67] wl[301] vdd gnd cell_6t
Xbit_r302_c67 bl[67] br[67] wl[302] vdd gnd cell_6t
Xbit_r303_c67 bl[67] br[67] wl[303] vdd gnd cell_6t
Xbit_r304_c67 bl[67] br[67] wl[304] vdd gnd cell_6t
Xbit_r305_c67 bl[67] br[67] wl[305] vdd gnd cell_6t
Xbit_r306_c67 bl[67] br[67] wl[306] vdd gnd cell_6t
Xbit_r307_c67 bl[67] br[67] wl[307] vdd gnd cell_6t
Xbit_r308_c67 bl[67] br[67] wl[308] vdd gnd cell_6t
Xbit_r309_c67 bl[67] br[67] wl[309] vdd gnd cell_6t
Xbit_r310_c67 bl[67] br[67] wl[310] vdd gnd cell_6t
Xbit_r311_c67 bl[67] br[67] wl[311] vdd gnd cell_6t
Xbit_r312_c67 bl[67] br[67] wl[312] vdd gnd cell_6t
Xbit_r313_c67 bl[67] br[67] wl[313] vdd gnd cell_6t
Xbit_r314_c67 bl[67] br[67] wl[314] vdd gnd cell_6t
Xbit_r315_c67 bl[67] br[67] wl[315] vdd gnd cell_6t
Xbit_r316_c67 bl[67] br[67] wl[316] vdd gnd cell_6t
Xbit_r317_c67 bl[67] br[67] wl[317] vdd gnd cell_6t
Xbit_r318_c67 bl[67] br[67] wl[318] vdd gnd cell_6t
Xbit_r319_c67 bl[67] br[67] wl[319] vdd gnd cell_6t
Xbit_r320_c67 bl[67] br[67] wl[320] vdd gnd cell_6t
Xbit_r321_c67 bl[67] br[67] wl[321] vdd gnd cell_6t
Xbit_r322_c67 bl[67] br[67] wl[322] vdd gnd cell_6t
Xbit_r323_c67 bl[67] br[67] wl[323] vdd gnd cell_6t
Xbit_r324_c67 bl[67] br[67] wl[324] vdd gnd cell_6t
Xbit_r325_c67 bl[67] br[67] wl[325] vdd gnd cell_6t
Xbit_r326_c67 bl[67] br[67] wl[326] vdd gnd cell_6t
Xbit_r327_c67 bl[67] br[67] wl[327] vdd gnd cell_6t
Xbit_r328_c67 bl[67] br[67] wl[328] vdd gnd cell_6t
Xbit_r329_c67 bl[67] br[67] wl[329] vdd gnd cell_6t
Xbit_r330_c67 bl[67] br[67] wl[330] vdd gnd cell_6t
Xbit_r331_c67 bl[67] br[67] wl[331] vdd gnd cell_6t
Xbit_r332_c67 bl[67] br[67] wl[332] vdd gnd cell_6t
Xbit_r333_c67 bl[67] br[67] wl[333] vdd gnd cell_6t
Xbit_r334_c67 bl[67] br[67] wl[334] vdd gnd cell_6t
Xbit_r335_c67 bl[67] br[67] wl[335] vdd gnd cell_6t
Xbit_r336_c67 bl[67] br[67] wl[336] vdd gnd cell_6t
Xbit_r337_c67 bl[67] br[67] wl[337] vdd gnd cell_6t
Xbit_r338_c67 bl[67] br[67] wl[338] vdd gnd cell_6t
Xbit_r339_c67 bl[67] br[67] wl[339] vdd gnd cell_6t
Xbit_r340_c67 bl[67] br[67] wl[340] vdd gnd cell_6t
Xbit_r341_c67 bl[67] br[67] wl[341] vdd gnd cell_6t
Xbit_r342_c67 bl[67] br[67] wl[342] vdd gnd cell_6t
Xbit_r343_c67 bl[67] br[67] wl[343] vdd gnd cell_6t
Xbit_r344_c67 bl[67] br[67] wl[344] vdd gnd cell_6t
Xbit_r345_c67 bl[67] br[67] wl[345] vdd gnd cell_6t
Xbit_r346_c67 bl[67] br[67] wl[346] vdd gnd cell_6t
Xbit_r347_c67 bl[67] br[67] wl[347] vdd gnd cell_6t
Xbit_r348_c67 bl[67] br[67] wl[348] vdd gnd cell_6t
Xbit_r349_c67 bl[67] br[67] wl[349] vdd gnd cell_6t
Xbit_r350_c67 bl[67] br[67] wl[350] vdd gnd cell_6t
Xbit_r351_c67 bl[67] br[67] wl[351] vdd gnd cell_6t
Xbit_r352_c67 bl[67] br[67] wl[352] vdd gnd cell_6t
Xbit_r353_c67 bl[67] br[67] wl[353] vdd gnd cell_6t
Xbit_r354_c67 bl[67] br[67] wl[354] vdd gnd cell_6t
Xbit_r355_c67 bl[67] br[67] wl[355] vdd gnd cell_6t
Xbit_r356_c67 bl[67] br[67] wl[356] vdd gnd cell_6t
Xbit_r357_c67 bl[67] br[67] wl[357] vdd gnd cell_6t
Xbit_r358_c67 bl[67] br[67] wl[358] vdd gnd cell_6t
Xbit_r359_c67 bl[67] br[67] wl[359] vdd gnd cell_6t
Xbit_r360_c67 bl[67] br[67] wl[360] vdd gnd cell_6t
Xbit_r361_c67 bl[67] br[67] wl[361] vdd gnd cell_6t
Xbit_r362_c67 bl[67] br[67] wl[362] vdd gnd cell_6t
Xbit_r363_c67 bl[67] br[67] wl[363] vdd gnd cell_6t
Xbit_r364_c67 bl[67] br[67] wl[364] vdd gnd cell_6t
Xbit_r365_c67 bl[67] br[67] wl[365] vdd gnd cell_6t
Xbit_r366_c67 bl[67] br[67] wl[366] vdd gnd cell_6t
Xbit_r367_c67 bl[67] br[67] wl[367] vdd gnd cell_6t
Xbit_r368_c67 bl[67] br[67] wl[368] vdd gnd cell_6t
Xbit_r369_c67 bl[67] br[67] wl[369] vdd gnd cell_6t
Xbit_r370_c67 bl[67] br[67] wl[370] vdd gnd cell_6t
Xbit_r371_c67 bl[67] br[67] wl[371] vdd gnd cell_6t
Xbit_r372_c67 bl[67] br[67] wl[372] vdd gnd cell_6t
Xbit_r373_c67 bl[67] br[67] wl[373] vdd gnd cell_6t
Xbit_r374_c67 bl[67] br[67] wl[374] vdd gnd cell_6t
Xbit_r375_c67 bl[67] br[67] wl[375] vdd gnd cell_6t
Xbit_r376_c67 bl[67] br[67] wl[376] vdd gnd cell_6t
Xbit_r377_c67 bl[67] br[67] wl[377] vdd gnd cell_6t
Xbit_r378_c67 bl[67] br[67] wl[378] vdd gnd cell_6t
Xbit_r379_c67 bl[67] br[67] wl[379] vdd gnd cell_6t
Xbit_r380_c67 bl[67] br[67] wl[380] vdd gnd cell_6t
Xbit_r381_c67 bl[67] br[67] wl[381] vdd gnd cell_6t
Xbit_r382_c67 bl[67] br[67] wl[382] vdd gnd cell_6t
Xbit_r383_c67 bl[67] br[67] wl[383] vdd gnd cell_6t
Xbit_r384_c67 bl[67] br[67] wl[384] vdd gnd cell_6t
Xbit_r385_c67 bl[67] br[67] wl[385] vdd gnd cell_6t
Xbit_r386_c67 bl[67] br[67] wl[386] vdd gnd cell_6t
Xbit_r387_c67 bl[67] br[67] wl[387] vdd gnd cell_6t
Xbit_r388_c67 bl[67] br[67] wl[388] vdd gnd cell_6t
Xbit_r389_c67 bl[67] br[67] wl[389] vdd gnd cell_6t
Xbit_r390_c67 bl[67] br[67] wl[390] vdd gnd cell_6t
Xbit_r391_c67 bl[67] br[67] wl[391] vdd gnd cell_6t
Xbit_r392_c67 bl[67] br[67] wl[392] vdd gnd cell_6t
Xbit_r393_c67 bl[67] br[67] wl[393] vdd gnd cell_6t
Xbit_r394_c67 bl[67] br[67] wl[394] vdd gnd cell_6t
Xbit_r395_c67 bl[67] br[67] wl[395] vdd gnd cell_6t
Xbit_r396_c67 bl[67] br[67] wl[396] vdd gnd cell_6t
Xbit_r397_c67 bl[67] br[67] wl[397] vdd gnd cell_6t
Xbit_r398_c67 bl[67] br[67] wl[398] vdd gnd cell_6t
Xbit_r399_c67 bl[67] br[67] wl[399] vdd gnd cell_6t
Xbit_r400_c67 bl[67] br[67] wl[400] vdd gnd cell_6t
Xbit_r401_c67 bl[67] br[67] wl[401] vdd gnd cell_6t
Xbit_r402_c67 bl[67] br[67] wl[402] vdd gnd cell_6t
Xbit_r403_c67 bl[67] br[67] wl[403] vdd gnd cell_6t
Xbit_r404_c67 bl[67] br[67] wl[404] vdd gnd cell_6t
Xbit_r405_c67 bl[67] br[67] wl[405] vdd gnd cell_6t
Xbit_r406_c67 bl[67] br[67] wl[406] vdd gnd cell_6t
Xbit_r407_c67 bl[67] br[67] wl[407] vdd gnd cell_6t
Xbit_r408_c67 bl[67] br[67] wl[408] vdd gnd cell_6t
Xbit_r409_c67 bl[67] br[67] wl[409] vdd gnd cell_6t
Xbit_r410_c67 bl[67] br[67] wl[410] vdd gnd cell_6t
Xbit_r411_c67 bl[67] br[67] wl[411] vdd gnd cell_6t
Xbit_r412_c67 bl[67] br[67] wl[412] vdd gnd cell_6t
Xbit_r413_c67 bl[67] br[67] wl[413] vdd gnd cell_6t
Xbit_r414_c67 bl[67] br[67] wl[414] vdd gnd cell_6t
Xbit_r415_c67 bl[67] br[67] wl[415] vdd gnd cell_6t
Xbit_r416_c67 bl[67] br[67] wl[416] vdd gnd cell_6t
Xbit_r417_c67 bl[67] br[67] wl[417] vdd gnd cell_6t
Xbit_r418_c67 bl[67] br[67] wl[418] vdd gnd cell_6t
Xbit_r419_c67 bl[67] br[67] wl[419] vdd gnd cell_6t
Xbit_r420_c67 bl[67] br[67] wl[420] vdd gnd cell_6t
Xbit_r421_c67 bl[67] br[67] wl[421] vdd gnd cell_6t
Xbit_r422_c67 bl[67] br[67] wl[422] vdd gnd cell_6t
Xbit_r423_c67 bl[67] br[67] wl[423] vdd gnd cell_6t
Xbit_r424_c67 bl[67] br[67] wl[424] vdd gnd cell_6t
Xbit_r425_c67 bl[67] br[67] wl[425] vdd gnd cell_6t
Xbit_r426_c67 bl[67] br[67] wl[426] vdd gnd cell_6t
Xbit_r427_c67 bl[67] br[67] wl[427] vdd gnd cell_6t
Xbit_r428_c67 bl[67] br[67] wl[428] vdd gnd cell_6t
Xbit_r429_c67 bl[67] br[67] wl[429] vdd gnd cell_6t
Xbit_r430_c67 bl[67] br[67] wl[430] vdd gnd cell_6t
Xbit_r431_c67 bl[67] br[67] wl[431] vdd gnd cell_6t
Xbit_r432_c67 bl[67] br[67] wl[432] vdd gnd cell_6t
Xbit_r433_c67 bl[67] br[67] wl[433] vdd gnd cell_6t
Xbit_r434_c67 bl[67] br[67] wl[434] vdd gnd cell_6t
Xbit_r435_c67 bl[67] br[67] wl[435] vdd gnd cell_6t
Xbit_r436_c67 bl[67] br[67] wl[436] vdd gnd cell_6t
Xbit_r437_c67 bl[67] br[67] wl[437] vdd gnd cell_6t
Xbit_r438_c67 bl[67] br[67] wl[438] vdd gnd cell_6t
Xbit_r439_c67 bl[67] br[67] wl[439] vdd gnd cell_6t
Xbit_r440_c67 bl[67] br[67] wl[440] vdd gnd cell_6t
Xbit_r441_c67 bl[67] br[67] wl[441] vdd gnd cell_6t
Xbit_r442_c67 bl[67] br[67] wl[442] vdd gnd cell_6t
Xbit_r443_c67 bl[67] br[67] wl[443] vdd gnd cell_6t
Xbit_r444_c67 bl[67] br[67] wl[444] vdd gnd cell_6t
Xbit_r445_c67 bl[67] br[67] wl[445] vdd gnd cell_6t
Xbit_r446_c67 bl[67] br[67] wl[446] vdd gnd cell_6t
Xbit_r447_c67 bl[67] br[67] wl[447] vdd gnd cell_6t
Xbit_r448_c67 bl[67] br[67] wl[448] vdd gnd cell_6t
Xbit_r449_c67 bl[67] br[67] wl[449] vdd gnd cell_6t
Xbit_r450_c67 bl[67] br[67] wl[450] vdd gnd cell_6t
Xbit_r451_c67 bl[67] br[67] wl[451] vdd gnd cell_6t
Xbit_r452_c67 bl[67] br[67] wl[452] vdd gnd cell_6t
Xbit_r453_c67 bl[67] br[67] wl[453] vdd gnd cell_6t
Xbit_r454_c67 bl[67] br[67] wl[454] vdd gnd cell_6t
Xbit_r455_c67 bl[67] br[67] wl[455] vdd gnd cell_6t
Xbit_r456_c67 bl[67] br[67] wl[456] vdd gnd cell_6t
Xbit_r457_c67 bl[67] br[67] wl[457] vdd gnd cell_6t
Xbit_r458_c67 bl[67] br[67] wl[458] vdd gnd cell_6t
Xbit_r459_c67 bl[67] br[67] wl[459] vdd gnd cell_6t
Xbit_r460_c67 bl[67] br[67] wl[460] vdd gnd cell_6t
Xbit_r461_c67 bl[67] br[67] wl[461] vdd gnd cell_6t
Xbit_r462_c67 bl[67] br[67] wl[462] vdd gnd cell_6t
Xbit_r463_c67 bl[67] br[67] wl[463] vdd gnd cell_6t
Xbit_r464_c67 bl[67] br[67] wl[464] vdd gnd cell_6t
Xbit_r465_c67 bl[67] br[67] wl[465] vdd gnd cell_6t
Xbit_r466_c67 bl[67] br[67] wl[466] vdd gnd cell_6t
Xbit_r467_c67 bl[67] br[67] wl[467] vdd gnd cell_6t
Xbit_r468_c67 bl[67] br[67] wl[468] vdd gnd cell_6t
Xbit_r469_c67 bl[67] br[67] wl[469] vdd gnd cell_6t
Xbit_r470_c67 bl[67] br[67] wl[470] vdd gnd cell_6t
Xbit_r471_c67 bl[67] br[67] wl[471] vdd gnd cell_6t
Xbit_r472_c67 bl[67] br[67] wl[472] vdd gnd cell_6t
Xbit_r473_c67 bl[67] br[67] wl[473] vdd gnd cell_6t
Xbit_r474_c67 bl[67] br[67] wl[474] vdd gnd cell_6t
Xbit_r475_c67 bl[67] br[67] wl[475] vdd gnd cell_6t
Xbit_r476_c67 bl[67] br[67] wl[476] vdd gnd cell_6t
Xbit_r477_c67 bl[67] br[67] wl[477] vdd gnd cell_6t
Xbit_r478_c67 bl[67] br[67] wl[478] vdd gnd cell_6t
Xbit_r479_c67 bl[67] br[67] wl[479] vdd gnd cell_6t
Xbit_r480_c67 bl[67] br[67] wl[480] vdd gnd cell_6t
Xbit_r481_c67 bl[67] br[67] wl[481] vdd gnd cell_6t
Xbit_r482_c67 bl[67] br[67] wl[482] vdd gnd cell_6t
Xbit_r483_c67 bl[67] br[67] wl[483] vdd gnd cell_6t
Xbit_r484_c67 bl[67] br[67] wl[484] vdd gnd cell_6t
Xbit_r485_c67 bl[67] br[67] wl[485] vdd gnd cell_6t
Xbit_r486_c67 bl[67] br[67] wl[486] vdd gnd cell_6t
Xbit_r487_c67 bl[67] br[67] wl[487] vdd gnd cell_6t
Xbit_r488_c67 bl[67] br[67] wl[488] vdd gnd cell_6t
Xbit_r489_c67 bl[67] br[67] wl[489] vdd gnd cell_6t
Xbit_r490_c67 bl[67] br[67] wl[490] vdd gnd cell_6t
Xbit_r491_c67 bl[67] br[67] wl[491] vdd gnd cell_6t
Xbit_r492_c67 bl[67] br[67] wl[492] vdd gnd cell_6t
Xbit_r493_c67 bl[67] br[67] wl[493] vdd gnd cell_6t
Xbit_r494_c67 bl[67] br[67] wl[494] vdd gnd cell_6t
Xbit_r495_c67 bl[67] br[67] wl[495] vdd gnd cell_6t
Xbit_r496_c67 bl[67] br[67] wl[496] vdd gnd cell_6t
Xbit_r497_c67 bl[67] br[67] wl[497] vdd gnd cell_6t
Xbit_r498_c67 bl[67] br[67] wl[498] vdd gnd cell_6t
Xbit_r499_c67 bl[67] br[67] wl[499] vdd gnd cell_6t
Xbit_r500_c67 bl[67] br[67] wl[500] vdd gnd cell_6t
Xbit_r501_c67 bl[67] br[67] wl[501] vdd gnd cell_6t
Xbit_r502_c67 bl[67] br[67] wl[502] vdd gnd cell_6t
Xbit_r503_c67 bl[67] br[67] wl[503] vdd gnd cell_6t
Xbit_r504_c67 bl[67] br[67] wl[504] vdd gnd cell_6t
Xbit_r505_c67 bl[67] br[67] wl[505] vdd gnd cell_6t
Xbit_r506_c67 bl[67] br[67] wl[506] vdd gnd cell_6t
Xbit_r507_c67 bl[67] br[67] wl[507] vdd gnd cell_6t
Xbit_r508_c67 bl[67] br[67] wl[508] vdd gnd cell_6t
Xbit_r509_c67 bl[67] br[67] wl[509] vdd gnd cell_6t
Xbit_r510_c67 bl[67] br[67] wl[510] vdd gnd cell_6t
Xbit_r511_c67 bl[67] br[67] wl[511] vdd gnd cell_6t
Xbit_r0_c68 bl[68] br[68] wl[0] vdd gnd cell_6t
Xbit_r1_c68 bl[68] br[68] wl[1] vdd gnd cell_6t
Xbit_r2_c68 bl[68] br[68] wl[2] vdd gnd cell_6t
Xbit_r3_c68 bl[68] br[68] wl[3] vdd gnd cell_6t
Xbit_r4_c68 bl[68] br[68] wl[4] vdd gnd cell_6t
Xbit_r5_c68 bl[68] br[68] wl[5] vdd gnd cell_6t
Xbit_r6_c68 bl[68] br[68] wl[6] vdd gnd cell_6t
Xbit_r7_c68 bl[68] br[68] wl[7] vdd gnd cell_6t
Xbit_r8_c68 bl[68] br[68] wl[8] vdd gnd cell_6t
Xbit_r9_c68 bl[68] br[68] wl[9] vdd gnd cell_6t
Xbit_r10_c68 bl[68] br[68] wl[10] vdd gnd cell_6t
Xbit_r11_c68 bl[68] br[68] wl[11] vdd gnd cell_6t
Xbit_r12_c68 bl[68] br[68] wl[12] vdd gnd cell_6t
Xbit_r13_c68 bl[68] br[68] wl[13] vdd gnd cell_6t
Xbit_r14_c68 bl[68] br[68] wl[14] vdd gnd cell_6t
Xbit_r15_c68 bl[68] br[68] wl[15] vdd gnd cell_6t
Xbit_r16_c68 bl[68] br[68] wl[16] vdd gnd cell_6t
Xbit_r17_c68 bl[68] br[68] wl[17] vdd gnd cell_6t
Xbit_r18_c68 bl[68] br[68] wl[18] vdd gnd cell_6t
Xbit_r19_c68 bl[68] br[68] wl[19] vdd gnd cell_6t
Xbit_r20_c68 bl[68] br[68] wl[20] vdd gnd cell_6t
Xbit_r21_c68 bl[68] br[68] wl[21] vdd gnd cell_6t
Xbit_r22_c68 bl[68] br[68] wl[22] vdd gnd cell_6t
Xbit_r23_c68 bl[68] br[68] wl[23] vdd gnd cell_6t
Xbit_r24_c68 bl[68] br[68] wl[24] vdd gnd cell_6t
Xbit_r25_c68 bl[68] br[68] wl[25] vdd gnd cell_6t
Xbit_r26_c68 bl[68] br[68] wl[26] vdd gnd cell_6t
Xbit_r27_c68 bl[68] br[68] wl[27] vdd gnd cell_6t
Xbit_r28_c68 bl[68] br[68] wl[28] vdd gnd cell_6t
Xbit_r29_c68 bl[68] br[68] wl[29] vdd gnd cell_6t
Xbit_r30_c68 bl[68] br[68] wl[30] vdd gnd cell_6t
Xbit_r31_c68 bl[68] br[68] wl[31] vdd gnd cell_6t
Xbit_r32_c68 bl[68] br[68] wl[32] vdd gnd cell_6t
Xbit_r33_c68 bl[68] br[68] wl[33] vdd gnd cell_6t
Xbit_r34_c68 bl[68] br[68] wl[34] vdd gnd cell_6t
Xbit_r35_c68 bl[68] br[68] wl[35] vdd gnd cell_6t
Xbit_r36_c68 bl[68] br[68] wl[36] vdd gnd cell_6t
Xbit_r37_c68 bl[68] br[68] wl[37] vdd gnd cell_6t
Xbit_r38_c68 bl[68] br[68] wl[38] vdd gnd cell_6t
Xbit_r39_c68 bl[68] br[68] wl[39] vdd gnd cell_6t
Xbit_r40_c68 bl[68] br[68] wl[40] vdd gnd cell_6t
Xbit_r41_c68 bl[68] br[68] wl[41] vdd gnd cell_6t
Xbit_r42_c68 bl[68] br[68] wl[42] vdd gnd cell_6t
Xbit_r43_c68 bl[68] br[68] wl[43] vdd gnd cell_6t
Xbit_r44_c68 bl[68] br[68] wl[44] vdd gnd cell_6t
Xbit_r45_c68 bl[68] br[68] wl[45] vdd gnd cell_6t
Xbit_r46_c68 bl[68] br[68] wl[46] vdd gnd cell_6t
Xbit_r47_c68 bl[68] br[68] wl[47] vdd gnd cell_6t
Xbit_r48_c68 bl[68] br[68] wl[48] vdd gnd cell_6t
Xbit_r49_c68 bl[68] br[68] wl[49] vdd gnd cell_6t
Xbit_r50_c68 bl[68] br[68] wl[50] vdd gnd cell_6t
Xbit_r51_c68 bl[68] br[68] wl[51] vdd gnd cell_6t
Xbit_r52_c68 bl[68] br[68] wl[52] vdd gnd cell_6t
Xbit_r53_c68 bl[68] br[68] wl[53] vdd gnd cell_6t
Xbit_r54_c68 bl[68] br[68] wl[54] vdd gnd cell_6t
Xbit_r55_c68 bl[68] br[68] wl[55] vdd gnd cell_6t
Xbit_r56_c68 bl[68] br[68] wl[56] vdd gnd cell_6t
Xbit_r57_c68 bl[68] br[68] wl[57] vdd gnd cell_6t
Xbit_r58_c68 bl[68] br[68] wl[58] vdd gnd cell_6t
Xbit_r59_c68 bl[68] br[68] wl[59] vdd gnd cell_6t
Xbit_r60_c68 bl[68] br[68] wl[60] vdd gnd cell_6t
Xbit_r61_c68 bl[68] br[68] wl[61] vdd gnd cell_6t
Xbit_r62_c68 bl[68] br[68] wl[62] vdd gnd cell_6t
Xbit_r63_c68 bl[68] br[68] wl[63] vdd gnd cell_6t
Xbit_r64_c68 bl[68] br[68] wl[64] vdd gnd cell_6t
Xbit_r65_c68 bl[68] br[68] wl[65] vdd gnd cell_6t
Xbit_r66_c68 bl[68] br[68] wl[66] vdd gnd cell_6t
Xbit_r67_c68 bl[68] br[68] wl[67] vdd gnd cell_6t
Xbit_r68_c68 bl[68] br[68] wl[68] vdd gnd cell_6t
Xbit_r69_c68 bl[68] br[68] wl[69] vdd gnd cell_6t
Xbit_r70_c68 bl[68] br[68] wl[70] vdd gnd cell_6t
Xbit_r71_c68 bl[68] br[68] wl[71] vdd gnd cell_6t
Xbit_r72_c68 bl[68] br[68] wl[72] vdd gnd cell_6t
Xbit_r73_c68 bl[68] br[68] wl[73] vdd gnd cell_6t
Xbit_r74_c68 bl[68] br[68] wl[74] vdd gnd cell_6t
Xbit_r75_c68 bl[68] br[68] wl[75] vdd gnd cell_6t
Xbit_r76_c68 bl[68] br[68] wl[76] vdd gnd cell_6t
Xbit_r77_c68 bl[68] br[68] wl[77] vdd gnd cell_6t
Xbit_r78_c68 bl[68] br[68] wl[78] vdd gnd cell_6t
Xbit_r79_c68 bl[68] br[68] wl[79] vdd gnd cell_6t
Xbit_r80_c68 bl[68] br[68] wl[80] vdd gnd cell_6t
Xbit_r81_c68 bl[68] br[68] wl[81] vdd gnd cell_6t
Xbit_r82_c68 bl[68] br[68] wl[82] vdd gnd cell_6t
Xbit_r83_c68 bl[68] br[68] wl[83] vdd gnd cell_6t
Xbit_r84_c68 bl[68] br[68] wl[84] vdd gnd cell_6t
Xbit_r85_c68 bl[68] br[68] wl[85] vdd gnd cell_6t
Xbit_r86_c68 bl[68] br[68] wl[86] vdd gnd cell_6t
Xbit_r87_c68 bl[68] br[68] wl[87] vdd gnd cell_6t
Xbit_r88_c68 bl[68] br[68] wl[88] vdd gnd cell_6t
Xbit_r89_c68 bl[68] br[68] wl[89] vdd gnd cell_6t
Xbit_r90_c68 bl[68] br[68] wl[90] vdd gnd cell_6t
Xbit_r91_c68 bl[68] br[68] wl[91] vdd gnd cell_6t
Xbit_r92_c68 bl[68] br[68] wl[92] vdd gnd cell_6t
Xbit_r93_c68 bl[68] br[68] wl[93] vdd gnd cell_6t
Xbit_r94_c68 bl[68] br[68] wl[94] vdd gnd cell_6t
Xbit_r95_c68 bl[68] br[68] wl[95] vdd gnd cell_6t
Xbit_r96_c68 bl[68] br[68] wl[96] vdd gnd cell_6t
Xbit_r97_c68 bl[68] br[68] wl[97] vdd gnd cell_6t
Xbit_r98_c68 bl[68] br[68] wl[98] vdd gnd cell_6t
Xbit_r99_c68 bl[68] br[68] wl[99] vdd gnd cell_6t
Xbit_r100_c68 bl[68] br[68] wl[100] vdd gnd cell_6t
Xbit_r101_c68 bl[68] br[68] wl[101] vdd gnd cell_6t
Xbit_r102_c68 bl[68] br[68] wl[102] vdd gnd cell_6t
Xbit_r103_c68 bl[68] br[68] wl[103] vdd gnd cell_6t
Xbit_r104_c68 bl[68] br[68] wl[104] vdd gnd cell_6t
Xbit_r105_c68 bl[68] br[68] wl[105] vdd gnd cell_6t
Xbit_r106_c68 bl[68] br[68] wl[106] vdd gnd cell_6t
Xbit_r107_c68 bl[68] br[68] wl[107] vdd gnd cell_6t
Xbit_r108_c68 bl[68] br[68] wl[108] vdd gnd cell_6t
Xbit_r109_c68 bl[68] br[68] wl[109] vdd gnd cell_6t
Xbit_r110_c68 bl[68] br[68] wl[110] vdd gnd cell_6t
Xbit_r111_c68 bl[68] br[68] wl[111] vdd gnd cell_6t
Xbit_r112_c68 bl[68] br[68] wl[112] vdd gnd cell_6t
Xbit_r113_c68 bl[68] br[68] wl[113] vdd gnd cell_6t
Xbit_r114_c68 bl[68] br[68] wl[114] vdd gnd cell_6t
Xbit_r115_c68 bl[68] br[68] wl[115] vdd gnd cell_6t
Xbit_r116_c68 bl[68] br[68] wl[116] vdd gnd cell_6t
Xbit_r117_c68 bl[68] br[68] wl[117] vdd gnd cell_6t
Xbit_r118_c68 bl[68] br[68] wl[118] vdd gnd cell_6t
Xbit_r119_c68 bl[68] br[68] wl[119] vdd gnd cell_6t
Xbit_r120_c68 bl[68] br[68] wl[120] vdd gnd cell_6t
Xbit_r121_c68 bl[68] br[68] wl[121] vdd gnd cell_6t
Xbit_r122_c68 bl[68] br[68] wl[122] vdd gnd cell_6t
Xbit_r123_c68 bl[68] br[68] wl[123] vdd gnd cell_6t
Xbit_r124_c68 bl[68] br[68] wl[124] vdd gnd cell_6t
Xbit_r125_c68 bl[68] br[68] wl[125] vdd gnd cell_6t
Xbit_r126_c68 bl[68] br[68] wl[126] vdd gnd cell_6t
Xbit_r127_c68 bl[68] br[68] wl[127] vdd gnd cell_6t
Xbit_r128_c68 bl[68] br[68] wl[128] vdd gnd cell_6t
Xbit_r129_c68 bl[68] br[68] wl[129] vdd gnd cell_6t
Xbit_r130_c68 bl[68] br[68] wl[130] vdd gnd cell_6t
Xbit_r131_c68 bl[68] br[68] wl[131] vdd gnd cell_6t
Xbit_r132_c68 bl[68] br[68] wl[132] vdd gnd cell_6t
Xbit_r133_c68 bl[68] br[68] wl[133] vdd gnd cell_6t
Xbit_r134_c68 bl[68] br[68] wl[134] vdd gnd cell_6t
Xbit_r135_c68 bl[68] br[68] wl[135] vdd gnd cell_6t
Xbit_r136_c68 bl[68] br[68] wl[136] vdd gnd cell_6t
Xbit_r137_c68 bl[68] br[68] wl[137] vdd gnd cell_6t
Xbit_r138_c68 bl[68] br[68] wl[138] vdd gnd cell_6t
Xbit_r139_c68 bl[68] br[68] wl[139] vdd gnd cell_6t
Xbit_r140_c68 bl[68] br[68] wl[140] vdd gnd cell_6t
Xbit_r141_c68 bl[68] br[68] wl[141] vdd gnd cell_6t
Xbit_r142_c68 bl[68] br[68] wl[142] vdd gnd cell_6t
Xbit_r143_c68 bl[68] br[68] wl[143] vdd gnd cell_6t
Xbit_r144_c68 bl[68] br[68] wl[144] vdd gnd cell_6t
Xbit_r145_c68 bl[68] br[68] wl[145] vdd gnd cell_6t
Xbit_r146_c68 bl[68] br[68] wl[146] vdd gnd cell_6t
Xbit_r147_c68 bl[68] br[68] wl[147] vdd gnd cell_6t
Xbit_r148_c68 bl[68] br[68] wl[148] vdd gnd cell_6t
Xbit_r149_c68 bl[68] br[68] wl[149] vdd gnd cell_6t
Xbit_r150_c68 bl[68] br[68] wl[150] vdd gnd cell_6t
Xbit_r151_c68 bl[68] br[68] wl[151] vdd gnd cell_6t
Xbit_r152_c68 bl[68] br[68] wl[152] vdd gnd cell_6t
Xbit_r153_c68 bl[68] br[68] wl[153] vdd gnd cell_6t
Xbit_r154_c68 bl[68] br[68] wl[154] vdd gnd cell_6t
Xbit_r155_c68 bl[68] br[68] wl[155] vdd gnd cell_6t
Xbit_r156_c68 bl[68] br[68] wl[156] vdd gnd cell_6t
Xbit_r157_c68 bl[68] br[68] wl[157] vdd gnd cell_6t
Xbit_r158_c68 bl[68] br[68] wl[158] vdd gnd cell_6t
Xbit_r159_c68 bl[68] br[68] wl[159] vdd gnd cell_6t
Xbit_r160_c68 bl[68] br[68] wl[160] vdd gnd cell_6t
Xbit_r161_c68 bl[68] br[68] wl[161] vdd gnd cell_6t
Xbit_r162_c68 bl[68] br[68] wl[162] vdd gnd cell_6t
Xbit_r163_c68 bl[68] br[68] wl[163] vdd gnd cell_6t
Xbit_r164_c68 bl[68] br[68] wl[164] vdd gnd cell_6t
Xbit_r165_c68 bl[68] br[68] wl[165] vdd gnd cell_6t
Xbit_r166_c68 bl[68] br[68] wl[166] vdd gnd cell_6t
Xbit_r167_c68 bl[68] br[68] wl[167] vdd gnd cell_6t
Xbit_r168_c68 bl[68] br[68] wl[168] vdd gnd cell_6t
Xbit_r169_c68 bl[68] br[68] wl[169] vdd gnd cell_6t
Xbit_r170_c68 bl[68] br[68] wl[170] vdd gnd cell_6t
Xbit_r171_c68 bl[68] br[68] wl[171] vdd gnd cell_6t
Xbit_r172_c68 bl[68] br[68] wl[172] vdd gnd cell_6t
Xbit_r173_c68 bl[68] br[68] wl[173] vdd gnd cell_6t
Xbit_r174_c68 bl[68] br[68] wl[174] vdd gnd cell_6t
Xbit_r175_c68 bl[68] br[68] wl[175] vdd gnd cell_6t
Xbit_r176_c68 bl[68] br[68] wl[176] vdd gnd cell_6t
Xbit_r177_c68 bl[68] br[68] wl[177] vdd gnd cell_6t
Xbit_r178_c68 bl[68] br[68] wl[178] vdd gnd cell_6t
Xbit_r179_c68 bl[68] br[68] wl[179] vdd gnd cell_6t
Xbit_r180_c68 bl[68] br[68] wl[180] vdd gnd cell_6t
Xbit_r181_c68 bl[68] br[68] wl[181] vdd gnd cell_6t
Xbit_r182_c68 bl[68] br[68] wl[182] vdd gnd cell_6t
Xbit_r183_c68 bl[68] br[68] wl[183] vdd gnd cell_6t
Xbit_r184_c68 bl[68] br[68] wl[184] vdd gnd cell_6t
Xbit_r185_c68 bl[68] br[68] wl[185] vdd gnd cell_6t
Xbit_r186_c68 bl[68] br[68] wl[186] vdd gnd cell_6t
Xbit_r187_c68 bl[68] br[68] wl[187] vdd gnd cell_6t
Xbit_r188_c68 bl[68] br[68] wl[188] vdd gnd cell_6t
Xbit_r189_c68 bl[68] br[68] wl[189] vdd gnd cell_6t
Xbit_r190_c68 bl[68] br[68] wl[190] vdd gnd cell_6t
Xbit_r191_c68 bl[68] br[68] wl[191] vdd gnd cell_6t
Xbit_r192_c68 bl[68] br[68] wl[192] vdd gnd cell_6t
Xbit_r193_c68 bl[68] br[68] wl[193] vdd gnd cell_6t
Xbit_r194_c68 bl[68] br[68] wl[194] vdd gnd cell_6t
Xbit_r195_c68 bl[68] br[68] wl[195] vdd gnd cell_6t
Xbit_r196_c68 bl[68] br[68] wl[196] vdd gnd cell_6t
Xbit_r197_c68 bl[68] br[68] wl[197] vdd gnd cell_6t
Xbit_r198_c68 bl[68] br[68] wl[198] vdd gnd cell_6t
Xbit_r199_c68 bl[68] br[68] wl[199] vdd gnd cell_6t
Xbit_r200_c68 bl[68] br[68] wl[200] vdd gnd cell_6t
Xbit_r201_c68 bl[68] br[68] wl[201] vdd gnd cell_6t
Xbit_r202_c68 bl[68] br[68] wl[202] vdd gnd cell_6t
Xbit_r203_c68 bl[68] br[68] wl[203] vdd gnd cell_6t
Xbit_r204_c68 bl[68] br[68] wl[204] vdd gnd cell_6t
Xbit_r205_c68 bl[68] br[68] wl[205] vdd gnd cell_6t
Xbit_r206_c68 bl[68] br[68] wl[206] vdd gnd cell_6t
Xbit_r207_c68 bl[68] br[68] wl[207] vdd gnd cell_6t
Xbit_r208_c68 bl[68] br[68] wl[208] vdd gnd cell_6t
Xbit_r209_c68 bl[68] br[68] wl[209] vdd gnd cell_6t
Xbit_r210_c68 bl[68] br[68] wl[210] vdd gnd cell_6t
Xbit_r211_c68 bl[68] br[68] wl[211] vdd gnd cell_6t
Xbit_r212_c68 bl[68] br[68] wl[212] vdd gnd cell_6t
Xbit_r213_c68 bl[68] br[68] wl[213] vdd gnd cell_6t
Xbit_r214_c68 bl[68] br[68] wl[214] vdd gnd cell_6t
Xbit_r215_c68 bl[68] br[68] wl[215] vdd gnd cell_6t
Xbit_r216_c68 bl[68] br[68] wl[216] vdd gnd cell_6t
Xbit_r217_c68 bl[68] br[68] wl[217] vdd gnd cell_6t
Xbit_r218_c68 bl[68] br[68] wl[218] vdd gnd cell_6t
Xbit_r219_c68 bl[68] br[68] wl[219] vdd gnd cell_6t
Xbit_r220_c68 bl[68] br[68] wl[220] vdd gnd cell_6t
Xbit_r221_c68 bl[68] br[68] wl[221] vdd gnd cell_6t
Xbit_r222_c68 bl[68] br[68] wl[222] vdd gnd cell_6t
Xbit_r223_c68 bl[68] br[68] wl[223] vdd gnd cell_6t
Xbit_r224_c68 bl[68] br[68] wl[224] vdd gnd cell_6t
Xbit_r225_c68 bl[68] br[68] wl[225] vdd gnd cell_6t
Xbit_r226_c68 bl[68] br[68] wl[226] vdd gnd cell_6t
Xbit_r227_c68 bl[68] br[68] wl[227] vdd gnd cell_6t
Xbit_r228_c68 bl[68] br[68] wl[228] vdd gnd cell_6t
Xbit_r229_c68 bl[68] br[68] wl[229] vdd gnd cell_6t
Xbit_r230_c68 bl[68] br[68] wl[230] vdd gnd cell_6t
Xbit_r231_c68 bl[68] br[68] wl[231] vdd gnd cell_6t
Xbit_r232_c68 bl[68] br[68] wl[232] vdd gnd cell_6t
Xbit_r233_c68 bl[68] br[68] wl[233] vdd gnd cell_6t
Xbit_r234_c68 bl[68] br[68] wl[234] vdd gnd cell_6t
Xbit_r235_c68 bl[68] br[68] wl[235] vdd gnd cell_6t
Xbit_r236_c68 bl[68] br[68] wl[236] vdd gnd cell_6t
Xbit_r237_c68 bl[68] br[68] wl[237] vdd gnd cell_6t
Xbit_r238_c68 bl[68] br[68] wl[238] vdd gnd cell_6t
Xbit_r239_c68 bl[68] br[68] wl[239] vdd gnd cell_6t
Xbit_r240_c68 bl[68] br[68] wl[240] vdd gnd cell_6t
Xbit_r241_c68 bl[68] br[68] wl[241] vdd gnd cell_6t
Xbit_r242_c68 bl[68] br[68] wl[242] vdd gnd cell_6t
Xbit_r243_c68 bl[68] br[68] wl[243] vdd gnd cell_6t
Xbit_r244_c68 bl[68] br[68] wl[244] vdd gnd cell_6t
Xbit_r245_c68 bl[68] br[68] wl[245] vdd gnd cell_6t
Xbit_r246_c68 bl[68] br[68] wl[246] vdd gnd cell_6t
Xbit_r247_c68 bl[68] br[68] wl[247] vdd gnd cell_6t
Xbit_r248_c68 bl[68] br[68] wl[248] vdd gnd cell_6t
Xbit_r249_c68 bl[68] br[68] wl[249] vdd gnd cell_6t
Xbit_r250_c68 bl[68] br[68] wl[250] vdd gnd cell_6t
Xbit_r251_c68 bl[68] br[68] wl[251] vdd gnd cell_6t
Xbit_r252_c68 bl[68] br[68] wl[252] vdd gnd cell_6t
Xbit_r253_c68 bl[68] br[68] wl[253] vdd gnd cell_6t
Xbit_r254_c68 bl[68] br[68] wl[254] vdd gnd cell_6t
Xbit_r255_c68 bl[68] br[68] wl[255] vdd gnd cell_6t
Xbit_r256_c68 bl[68] br[68] wl[256] vdd gnd cell_6t
Xbit_r257_c68 bl[68] br[68] wl[257] vdd gnd cell_6t
Xbit_r258_c68 bl[68] br[68] wl[258] vdd gnd cell_6t
Xbit_r259_c68 bl[68] br[68] wl[259] vdd gnd cell_6t
Xbit_r260_c68 bl[68] br[68] wl[260] vdd gnd cell_6t
Xbit_r261_c68 bl[68] br[68] wl[261] vdd gnd cell_6t
Xbit_r262_c68 bl[68] br[68] wl[262] vdd gnd cell_6t
Xbit_r263_c68 bl[68] br[68] wl[263] vdd gnd cell_6t
Xbit_r264_c68 bl[68] br[68] wl[264] vdd gnd cell_6t
Xbit_r265_c68 bl[68] br[68] wl[265] vdd gnd cell_6t
Xbit_r266_c68 bl[68] br[68] wl[266] vdd gnd cell_6t
Xbit_r267_c68 bl[68] br[68] wl[267] vdd gnd cell_6t
Xbit_r268_c68 bl[68] br[68] wl[268] vdd gnd cell_6t
Xbit_r269_c68 bl[68] br[68] wl[269] vdd gnd cell_6t
Xbit_r270_c68 bl[68] br[68] wl[270] vdd gnd cell_6t
Xbit_r271_c68 bl[68] br[68] wl[271] vdd gnd cell_6t
Xbit_r272_c68 bl[68] br[68] wl[272] vdd gnd cell_6t
Xbit_r273_c68 bl[68] br[68] wl[273] vdd gnd cell_6t
Xbit_r274_c68 bl[68] br[68] wl[274] vdd gnd cell_6t
Xbit_r275_c68 bl[68] br[68] wl[275] vdd gnd cell_6t
Xbit_r276_c68 bl[68] br[68] wl[276] vdd gnd cell_6t
Xbit_r277_c68 bl[68] br[68] wl[277] vdd gnd cell_6t
Xbit_r278_c68 bl[68] br[68] wl[278] vdd gnd cell_6t
Xbit_r279_c68 bl[68] br[68] wl[279] vdd gnd cell_6t
Xbit_r280_c68 bl[68] br[68] wl[280] vdd gnd cell_6t
Xbit_r281_c68 bl[68] br[68] wl[281] vdd gnd cell_6t
Xbit_r282_c68 bl[68] br[68] wl[282] vdd gnd cell_6t
Xbit_r283_c68 bl[68] br[68] wl[283] vdd gnd cell_6t
Xbit_r284_c68 bl[68] br[68] wl[284] vdd gnd cell_6t
Xbit_r285_c68 bl[68] br[68] wl[285] vdd gnd cell_6t
Xbit_r286_c68 bl[68] br[68] wl[286] vdd gnd cell_6t
Xbit_r287_c68 bl[68] br[68] wl[287] vdd gnd cell_6t
Xbit_r288_c68 bl[68] br[68] wl[288] vdd gnd cell_6t
Xbit_r289_c68 bl[68] br[68] wl[289] vdd gnd cell_6t
Xbit_r290_c68 bl[68] br[68] wl[290] vdd gnd cell_6t
Xbit_r291_c68 bl[68] br[68] wl[291] vdd gnd cell_6t
Xbit_r292_c68 bl[68] br[68] wl[292] vdd gnd cell_6t
Xbit_r293_c68 bl[68] br[68] wl[293] vdd gnd cell_6t
Xbit_r294_c68 bl[68] br[68] wl[294] vdd gnd cell_6t
Xbit_r295_c68 bl[68] br[68] wl[295] vdd gnd cell_6t
Xbit_r296_c68 bl[68] br[68] wl[296] vdd gnd cell_6t
Xbit_r297_c68 bl[68] br[68] wl[297] vdd gnd cell_6t
Xbit_r298_c68 bl[68] br[68] wl[298] vdd gnd cell_6t
Xbit_r299_c68 bl[68] br[68] wl[299] vdd gnd cell_6t
Xbit_r300_c68 bl[68] br[68] wl[300] vdd gnd cell_6t
Xbit_r301_c68 bl[68] br[68] wl[301] vdd gnd cell_6t
Xbit_r302_c68 bl[68] br[68] wl[302] vdd gnd cell_6t
Xbit_r303_c68 bl[68] br[68] wl[303] vdd gnd cell_6t
Xbit_r304_c68 bl[68] br[68] wl[304] vdd gnd cell_6t
Xbit_r305_c68 bl[68] br[68] wl[305] vdd gnd cell_6t
Xbit_r306_c68 bl[68] br[68] wl[306] vdd gnd cell_6t
Xbit_r307_c68 bl[68] br[68] wl[307] vdd gnd cell_6t
Xbit_r308_c68 bl[68] br[68] wl[308] vdd gnd cell_6t
Xbit_r309_c68 bl[68] br[68] wl[309] vdd gnd cell_6t
Xbit_r310_c68 bl[68] br[68] wl[310] vdd gnd cell_6t
Xbit_r311_c68 bl[68] br[68] wl[311] vdd gnd cell_6t
Xbit_r312_c68 bl[68] br[68] wl[312] vdd gnd cell_6t
Xbit_r313_c68 bl[68] br[68] wl[313] vdd gnd cell_6t
Xbit_r314_c68 bl[68] br[68] wl[314] vdd gnd cell_6t
Xbit_r315_c68 bl[68] br[68] wl[315] vdd gnd cell_6t
Xbit_r316_c68 bl[68] br[68] wl[316] vdd gnd cell_6t
Xbit_r317_c68 bl[68] br[68] wl[317] vdd gnd cell_6t
Xbit_r318_c68 bl[68] br[68] wl[318] vdd gnd cell_6t
Xbit_r319_c68 bl[68] br[68] wl[319] vdd gnd cell_6t
Xbit_r320_c68 bl[68] br[68] wl[320] vdd gnd cell_6t
Xbit_r321_c68 bl[68] br[68] wl[321] vdd gnd cell_6t
Xbit_r322_c68 bl[68] br[68] wl[322] vdd gnd cell_6t
Xbit_r323_c68 bl[68] br[68] wl[323] vdd gnd cell_6t
Xbit_r324_c68 bl[68] br[68] wl[324] vdd gnd cell_6t
Xbit_r325_c68 bl[68] br[68] wl[325] vdd gnd cell_6t
Xbit_r326_c68 bl[68] br[68] wl[326] vdd gnd cell_6t
Xbit_r327_c68 bl[68] br[68] wl[327] vdd gnd cell_6t
Xbit_r328_c68 bl[68] br[68] wl[328] vdd gnd cell_6t
Xbit_r329_c68 bl[68] br[68] wl[329] vdd gnd cell_6t
Xbit_r330_c68 bl[68] br[68] wl[330] vdd gnd cell_6t
Xbit_r331_c68 bl[68] br[68] wl[331] vdd gnd cell_6t
Xbit_r332_c68 bl[68] br[68] wl[332] vdd gnd cell_6t
Xbit_r333_c68 bl[68] br[68] wl[333] vdd gnd cell_6t
Xbit_r334_c68 bl[68] br[68] wl[334] vdd gnd cell_6t
Xbit_r335_c68 bl[68] br[68] wl[335] vdd gnd cell_6t
Xbit_r336_c68 bl[68] br[68] wl[336] vdd gnd cell_6t
Xbit_r337_c68 bl[68] br[68] wl[337] vdd gnd cell_6t
Xbit_r338_c68 bl[68] br[68] wl[338] vdd gnd cell_6t
Xbit_r339_c68 bl[68] br[68] wl[339] vdd gnd cell_6t
Xbit_r340_c68 bl[68] br[68] wl[340] vdd gnd cell_6t
Xbit_r341_c68 bl[68] br[68] wl[341] vdd gnd cell_6t
Xbit_r342_c68 bl[68] br[68] wl[342] vdd gnd cell_6t
Xbit_r343_c68 bl[68] br[68] wl[343] vdd gnd cell_6t
Xbit_r344_c68 bl[68] br[68] wl[344] vdd gnd cell_6t
Xbit_r345_c68 bl[68] br[68] wl[345] vdd gnd cell_6t
Xbit_r346_c68 bl[68] br[68] wl[346] vdd gnd cell_6t
Xbit_r347_c68 bl[68] br[68] wl[347] vdd gnd cell_6t
Xbit_r348_c68 bl[68] br[68] wl[348] vdd gnd cell_6t
Xbit_r349_c68 bl[68] br[68] wl[349] vdd gnd cell_6t
Xbit_r350_c68 bl[68] br[68] wl[350] vdd gnd cell_6t
Xbit_r351_c68 bl[68] br[68] wl[351] vdd gnd cell_6t
Xbit_r352_c68 bl[68] br[68] wl[352] vdd gnd cell_6t
Xbit_r353_c68 bl[68] br[68] wl[353] vdd gnd cell_6t
Xbit_r354_c68 bl[68] br[68] wl[354] vdd gnd cell_6t
Xbit_r355_c68 bl[68] br[68] wl[355] vdd gnd cell_6t
Xbit_r356_c68 bl[68] br[68] wl[356] vdd gnd cell_6t
Xbit_r357_c68 bl[68] br[68] wl[357] vdd gnd cell_6t
Xbit_r358_c68 bl[68] br[68] wl[358] vdd gnd cell_6t
Xbit_r359_c68 bl[68] br[68] wl[359] vdd gnd cell_6t
Xbit_r360_c68 bl[68] br[68] wl[360] vdd gnd cell_6t
Xbit_r361_c68 bl[68] br[68] wl[361] vdd gnd cell_6t
Xbit_r362_c68 bl[68] br[68] wl[362] vdd gnd cell_6t
Xbit_r363_c68 bl[68] br[68] wl[363] vdd gnd cell_6t
Xbit_r364_c68 bl[68] br[68] wl[364] vdd gnd cell_6t
Xbit_r365_c68 bl[68] br[68] wl[365] vdd gnd cell_6t
Xbit_r366_c68 bl[68] br[68] wl[366] vdd gnd cell_6t
Xbit_r367_c68 bl[68] br[68] wl[367] vdd gnd cell_6t
Xbit_r368_c68 bl[68] br[68] wl[368] vdd gnd cell_6t
Xbit_r369_c68 bl[68] br[68] wl[369] vdd gnd cell_6t
Xbit_r370_c68 bl[68] br[68] wl[370] vdd gnd cell_6t
Xbit_r371_c68 bl[68] br[68] wl[371] vdd gnd cell_6t
Xbit_r372_c68 bl[68] br[68] wl[372] vdd gnd cell_6t
Xbit_r373_c68 bl[68] br[68] wl[373] vdd gnd cell_6t
Xbit_r374_c68 bl[68] br[68] wl[374] vdd gnd cell_6t
Xbit_r375_c68 bl[68] br[68] wl[375] vdd gnd cell_6t
Xbit_r376_c68 bl[68] br[68] wl[376] vdd gnd cell_6t
Xbit_r377_c68 bl[68] br[68] wl[377] vdd gnd cell_6t
Xbit_r378_c68 bl[68] br[68] wl[378] vdd gnd cell_6t
Xbit_r379_c68 bl[68] br[68] wl[379] vdd gnd cell_6t
Xbit_r380_c68 bl[68] br[68] wl[380] vdd gnd cell_6t
Xbit_r381_c68 bl[68] br[68] wl[381] vdd gnd cell_6t
Xbit_r382_c68 bl[68] br[68] wl[382] vdd gnd cell_6t
Xbit_r383_c68 bl[68] br[68] wl[383] vdd gnd cell_6t
Xbit_r384_c68 bl[68] br[68] wl[384] vdd gnd cell_6t
Xbit_r385_c68 bl[68] br[68] wl[385] vdd gnd cell_6t
Xbit_r386_c68 bl[68] br[68] wl[386] vdd gnd cell_6t
Xbit_r387_c68 bl[68] br[68] wl[387] vdd gnd cell_6t
Xbit_r388_c68 bl[68] br[68] wl[388] vdd gnd cell_6t
Xbit_r389_c68 bl[68] br[68] wl[389] vdd gnd cell_6t
Xbit_r390_c68 bl[68] br[68] wl[390] vdd gnd cell_6t
Xbit_r391_c68 bl[68] br[68] wl[391] vdd gnd cell_6t
Xbit_r392_c68 bl[68] br[68] wl[392] vdd gnd cell_6t
Xbit_r393_c68 bl[68] br[68] wl[393] vdd gnd cell_6t
Xbit_r394_c68 bl[68] br[68] wl[394] vdd gnd cell_6t
Xbit_r395_c68 bl[68] br[68] wl[395] vdd gnd cell_6t
Xbit_r396_c68 bl[68] br[68] wl[396] vdd gnd cell_6t
Xbit_r397_c68 bl[68] br[68] wl[397] vdd gnd cell_6t
Xbit_r398_c68 bl[68] br[68] wl[398] vdd gnd cell_6t
Xbit_r399_c68 bl[68] br[68] wl[399] vdd gnd cell_6t
Xbit_r400_c68 bl[68] br[68] wl[400] vdd gnd cell_6t
Xbit_r401_c68 bl[68] br[68] wl[401] vdd gnd cell_6t
Xbit_r402_c68 bl[68] br[68] wl[402] vdd gnd cell_6t
Xbit_r403_c68 bl[68] br[68] wl[403] vdd gnd cell_6t
Xbit_r404_c68 bl[68] br[68] wl[404] vdd gnd cell_6t
Xbit_r405_c68 bl[68] br[68] wl[405] vdd gnd cell_6t
Xbit_r406_c68 bl[68] br[68] wl[406] vdd gnd cell_6t
Xbit_r407_c68 bl[68] br[68] wl[407] vdd gnd cell_6t
Xbit_r408_c68 bl[68] br[68] wl[408] vdd gnd cell_6t
Xbit_r409_c68 bl[68] br[68] wl[409] vdd gnd cell_6t
Xbit_r410_c68 bl[68] br[68] wl[410] vdd gnd cell_6t
Xbit_r411_c68 bl[68] br[68] wl[411] vdd gnd cell_6t
Xbit_r412_c68 bl[68] br[68] wl[412] vdd gnd cell_6t
Xbit_r413_c68 bl[68] br[68] wl[413] vdd gnd cell_6t
Xbit_r414_c68 bl[68] br[68] wl[414] vdd gnd cell_6t
Xbit_r415_c68 bl[68] br[68] wl[415] vdd gnd cell_6t
Xbit_r416_c68 bl[68] br[68] wl[416] vdd gnd cell_6t
Xbit_r417_c68 bl[68] br[68] wl[417] vdd gnd cell_6t
Xbit_r418_c68 bl[68] br[68] wl[418] vdd gnd cell_6t
Xbit_r419_c68 bl[68] br[68] wl[419] vdd gnd cell_6t
Xbit_r420_c68 bl[68] br[68] wl[420] vdd gnd cell_6t
Xbit_r421_c68 bl[68] br[68] wl[421] vdd gnd cell_6t
Xbit_r422_c68 bl[68] br[68] wl[422] vdd gnd cell_6t
Xbit_r423_c68 bl[68] br[68] wl[423] vdd gnd cell_6t
Xbit_r424_c68 bl[68] br[68] wl[424] vdd gnd cell_6t
Xbit_r425_c68 bl[68] br[68] wl[425] vdd gnd cell_6t
Xbit_r426_c68 bl[68] br[68] wl[426] vdd gnd cell_6t
Xbit_r427_c68 bl[68] br[68] wl[427] vdd gnd cell_6t
Xbit_r428_c68 bl[68] br[68] wl[428] vdd gnd cell_6t
Xbit_r429_c68 bl[68] br[68] wl[429] vdd gnd cell_6t
Xbit_r430_c68 bl[68] br[68] wl[430] vdd gnd cell_6t
Xbit_r431_c68 bl[68] br[68] wl[431] vdd gnd cell_6t
Xbit_r432_c68 bl[68] br[68] wl[432] vdd gnd cell_6t
Xbit_r433_c68 bl[68] br[68] wl[433] vdd gnd cell_6t
Xbit_r434_c68 bl[68] br[68] wl[434] vdd gnd cell_6t
Xbit_r435_c68 bl[68] br[68] wl[435] vdd gnd cell_6t
Xbit_r436_c68 bl[68] br[68] wl[436] vdd gnd cell_6t
Xbit_r437_c68 bl[68] br[68] wl[437] vdd gnd cell_6t
Xbit_r438_c68 bl[68] br[68] wl[438] vdd gnd cell_6t
Xbit_r439_c68 bl[68] br[68] wl[439] vdd gnd cell_6t
Xbit_r440_c68 bl[68] br[68] wl[440] vdd gnd cell_6t
Xbit_r441_c68 bl[68] br[68] wl[441] vdd gnd cell_6t
Xbit_r442_c68 bl[68] br[68] wl[442] vdd gnd cell_6t
Xbit_r443_c68 bl[68] br[68] wl[443] vdd gnd cell_6t
Xbit_r444_c68 bl[68] br[68] wl[444] vdd gnd cell_6t
Xbit_r445_c68 bl[68] br[68] wl[445] vdd gnd cell_6t
Xbit_r446_c68 bl[68] br[68] wl[446] vdd gnd cell_6t
Xbit_r447_c68 bl[68] br[68] wl[447] vdd gnd cell_6t
Xbit_r448_c68 bl[68] br[68] wl[448] vdd gnd cell_6t
Xbit_r449_c68 bl[68] br[68] wl[449] vdd gnd cell_6t
Xbit_r450_c68 bl[68] br[68] wl[450] vdd gnd cell_6t
Xbit_r451_c68 bl[68] br[68] wl[451] vdd gnd cell_6t
Xbit_r452_c68 bl[68] br[68] wl[452] vdd gnd cell_6t
Xbit_r453_c68 bl[68] br[68] wl[453] vdd gnd cell_6t
Xbit_r454_c68 bl[68] br[68] wl[454] vdd gnd cell_6t
Xbit_r455_c68 bl[68] br[68] wl[455] vdd gnd cell_6t
Xbit_r456_c68 bl[68] br[68] wl[456] vdd gnd cell_6t
Xbit_r457_c68 bl[68] br[68] wl[457] vdd gnd cell_6t
Xbit_r458_c68 bl[68] br[68] wl[458] vdd gnd cell_6t
Xbit_r459_c68 bl[68] br[68] wl[459] vdd gnd cell_6t
Xbit_r460_c68 bl[68] br[68] wl[460] vdd gnd cell_6t
Xbit_r461_c68 bl[68] br[68] wl[461] vdd gnd cell_6t
Xbit_r462_c68 bl[68] br[68] wl[462] vdd gnd cell_6t
Xbit_r463_c68 bl[68] br[68] wl[463] vdd gnd cell_6t
Xbit_r464_c68 bl[68] br[68] wl[464] vdd gnd cell_6t
Xbit_r465_c68 bl[68] br[68] wl[465] vdd gnd cell_6t
Xbit_r466_c68 bl[68] br[68] wl[466] vdd gnd cell_6t
Xbit_r467_c68 bl[68] br[68] wl[467] vdd gnd cell_6t
Xbit_r468_c68 bl[68] br[68] wl[468] vdd gnd cell_6t
Xbit_r469_c68 bl[68] br[68] wl[469] vdd gnd cell_6t
Xbit_r470_c68 bl[68] br[68] wl[470] vdd gnd cell_6t
Xbit_r471_c68 bl[68] br[68] wl[471] vdd gnd cell_6t
Xbit_r472_c68 bl[68] br[68] wl[472] vdd gnd cell_6t
Xbit_r473_c68 bl[68] br[68] wl[473] vdd gnd cell_6t
Xbit_r474_c68 bl[68] br[68] wl[474] vdd gnd cell_6t
Xbit_r475_c68 bl[68] br[68] wl[475] vdd gnd cell_6t
Xbit_r476_c68 bl[68] br[68] wl[476] vdd gnd cell_6t
Xbit_r477_c68 bl[68] br[68] wl[477] vdd gnd cell_6t
Xbit_r478_c68 bl[68] br[68] wl[478] vdd gnd cell_6t
Xbit_r479_c68 bl[68] br[68] wl[479] vdd gnd cell_6t
Xbit_r480_c68 bl[68] br[68] wl[480] vdd gnd cell_6t
Xbit_r481_c68 bl[68] br[68] wl[481] vdd gnd cell_6t
Xbit_r482_c68 bl[68] br[68] wl[482] vdd gnd cell_6t
Xbit_r483_c68 bl[68] br[68] wl[483] vdd gnd cell_6t
Xbit_r484_c68 bl[68] br[68] wl[484] vdd gnd cell_6t
Xbit_r485_c68 bl[68] br[68] wl[485] vdd gnd cell_6t
Xbit_r486_c68 bl[68] br[68] wl[486] vdd gnd cell_6t
Xbit_r487_c68 bl[68] br[68] wl[487] vdd gnd cell_6t
Xbit_r488_c68 bl[68] br[68] wl[488] vdd gnd cell_6t
Xbit_r489_c68 bl[68] br[68] wl[489] vdd gnd cell_6t
Xbit_r490_c68 bl[68] br[68] wl[490] vdd gnd cell_6t
Xbit_r491_c68 bl[68] br[68] wl[491] vdd gnd cell_6t
Xbit_r492_c68 bl[68] br[68] wl[492] vdd gnd cell_6t
Xbit_r493_c68 bl[68] br[68] wl[493] vdd gnd cell_6t
Xbit_r494_c68 bl[68] br[68] wl[494] vdd gnd cell_6t
Xbit_r495_c68 bl[68] br[68] wl[495] vdd gnd cell_6t
Xbit_r496_c68 bl[68] br[68] wl[496] vdd gnd cell_6t
Xbit_r497_c68 bl[68] br[68] wl[497] vdd gnd cell_6t
Xbit_r498_c68 bl[68] br[68] wl[498] vdd gnd cell_6t
Xbit_r499_c68 bl[68] br[68] wl[499] vdd gnd cell_6t
Xbit_r500_c68 bl[68] br[68] wl[500] vdd gnd cell_6t
Xbit_r501_c68 bl[68] br[68] wl[501] vdd gnd cell_6t
Xbit_r502_c68 bl[68] br[68] wl[502] vdd gnd cell_6t
Xbit_r503_c68 bl[68] br[68] wl[503] vdd gnd cell_6t
Xbit_r504_c68 bl[68] br[68] wl[504] vdd gnd cell_6t
Xbit_r505_c68 bl[68] br[68] wl[505] vdd gnd cell_6t
Xbit_r506_c68 bl[68] br[68] wl[506] vdd gnd cell_6t
Xbit_r507_c68 bl[68] br[68] wl[507] vdd gnd cell_6t
Xbit_r508_c68 bl[68] br[68] wl[508] vdd gnd cell_6t
Xbit_r509_c68 bl[68] br[68] wl[509] vdd gnd cell_6t
Xbit_r510_c68 bl[68] br[68] wl[510] vdd gnd cell_6t
Xbit_r511_c68 bl[68] br[68] wl[511] vdd gnd cell_6t
Xbit_r0_c69 bl[69] br[69] wl[0] vdd gnd cell_6t
Xbit_r1_c69 bl[69] br[69] wl[1] vdd gnd cell_6t
Xbit_r2_c69 bl[69] br[69] wl[2] vdd gnd cell_6t
Xbit_r3_c69 bl[69] br[69] wl[3] vdd gnd cell_6t
Xbit_r4_c69 bl[69] br[69] wl[4] vdd gnd cell_6t
Xbit_r5_c69 bl[69] br[69] wl[5] vdd gnd cell_6t
Xbit_r6_c69 bl[69] br[69] wl[6] vdd gnd cell_6t
Xbit_r7_c69 bl[69] br[69] wl[7] vdd gnd cell_6t
Xbit_r8_c69 bl[69] br[69] wl[8] vdd gnd cell_6t
Xbit_r9_c69 bl[69] br[69] wl[9] vdd gnd cell_6t
Xbit_r10_c69 bl[69] br[69] wl[10] vdd gnd cell_6t
Xbit_r11_c69 bl[69] br[69] wl[11] vdd gnd cell_6t
Xbit_r12_c69 bl[69] br[69] wl[12] vdd gnd cell_6t
Xbit_r13_c69 bl[69] br[69] wl[13] vdd gnd cell_6t
Xbit_r14_c69 bl[69] br[69] wl[14] vdd gnd cell_6t
Xbit_r15_c69 bl[69] br[69] wl[15] vdd gnd cell_6t
Xbit_r16_c69 bl[69] br[69] wl[16] vdd gnd cell_6t
Xbit_r17_c69 bl[69] br[69] wl[17] vdd gnd cell_6t
Xbit_r18_c69 bl[69] br[69] wl[18] vdd gnd cell_6t
Xbit_r19_c69 bl[69] br[69] wl[19] vdd gnd cell_6t
Xbit_r20_c69 bl[69] br[69] wl[20] vdd gnd cell_6t
Xbit_r21_c69 bl[69] br[69] wl[21] vdd gnd cell_6t
Xbit_r22_c69 bl[69] br[69] wl[22] vdd gnd cell_6t
Xbit_r23_c69 bl[69] br[69] wl[23] vdd gnd cell_6t
Xbit_r24_c69 bl[69] br[69] wl[24] vdd gnd cell_6t
Xbit_r25_c69 bl[69] br[69] wl[25] vdd gnd cell_6t
Xbit_r26_c69 bl[69] br[69] wl[26] vdd gnd cell_6t
Xbit_r27_c69 bl[69] br[69] wl[27] vdd gnd cell_6t
Xbit_r28_c69 bl[69] br[69] wl[28] vdd gnd cell_6t
Xbit_r29_c69 bl[69] br[69] wl[29] vdd gnd cell_6t
Xbit_r30_c69 bl[69] br[69] wl[30] vdd gnd cell_6t
Xbit_r31_c69 bl[69] br[69] wl[31] vdd gnd cell_6t
Xbit_r32_c69 bl[69] br[69] wl[32] vdd gnd cell_6t
Xbit_r33_c69 bl[69] br[69] wl[33] vdd gnd cell_6t
Xbit_r34_c69 bl[69] br[69] wl[34] vdd gnd cell_6t
Xbit_r35_c69 bl[69] br[69] wl[35] vdd gnd cell_6t
Xbit_r36_c69 bl[69] br[69] wl[36] vdd gnd cell_6t
Xbit_r37_c69 bl[69] br[69] wl[37] vdd gnd cell_6t
Xbit_r38_c69 bl[69] br[69] wl[38] vdd gnd cell_6t
Xbit_r39_c69 bl[69] br[69] wl[39] vdd gnd cell_6t
Xbit_r40_c69 bl[69] br[69] wl[40] vdd gnd cell_6t
Xbit_r41_c69 bl[69] br[69] wl[41] vdd gnd cell_6t
Xbit_r42_c69 bl[69] br[69] wl[42] vdd gnd cell_6t
Xbit_r43_c69 bl[69] br[69] wl[43] vdd gnd cell_6t
Xbit_r44_c69 bl[69] br[69] wl[44] vdd gnd cell_6t
Xbit_r45_c69 bl[69] br[69] wl[45] vdd gnd cell_6t
Xbit_r46_c69 bl[69] br[69] wl[46] vdd gnd cell_6t
Xbit_r47_c69 bl[69] br[69] wl[47] vdd gnd cell_6t
Xbit_r48_c69 bl[69] br[69] wl[48] vdd gnd cell_6t
Xbit_r49_c69 bl[69] br[69] wl[49] vdd gnd cell_6t
Xbit_r50_c69 bl[69] br[69] wl[50] vdd gnd cell_6t
Xbit_r51_c69 bl[69] br[69] wl[51] vdd gnd cell_6t
Xbit_r52_c69 bl[69] br[69] wl[52] vdd gnd cell_6t
Xbit_r53_c69 bl[69] br[69] wl[53] vdd gnd cell_6t
Xbit_r54_c69 bl[69] br[69] wl[54] vdd gnd cell_6t
Xbit_r55_c69 bl[69] br[69] wl[55] vdd gnd cell_6t
Xbit_r56_c69 bl[69] br[69] wl[56] vdd gnd cell_6t
Xbit_r57_c69 bl[69] br[69] wl[57] vdd gnd cell_6t
Xbit_r58_c69 bl[69] br[69] wl[58] vdd gnd cell_6t
Xbit_r59_c69 bl[69] br[69] wl[59] vdd gnd cell_6t
Xbit_r60_c69 bl[69] br[69] wl[60] vdd gnd cell_6t
Xbit_r61_c69 bl[69] br[69] wl[61] vdd gnd cell_6t
Xbit_r62_c69 bl[69] br[69] wl[62] vdd gnd cell_6t
Xbit_r63_c69 bl[69] br[69] wl[63] vdd gnd cell_6t
Xbit_r64_c69 bl[69] br[69] wl[64] vdd gnd cell_6t
Xbit_r65_c69 bl[69] br[69] wl[65] vdd gnd cell_6t
Xbit_r66_c69 bl[69] br[69] wl[66] vdd gnd cell_6t
Xbit_r67_c69 bl[69] br[69] wl[67] vdd gnd cell_6t
Xbit_r68_c69 bl[69] br[69] wl[68] vdd gnd cell_6t
Xbit_r69_c69 bl[69] br[69] wl[69] vdd gnd cell_6t
Xbit_r70_c69 bl[69] br[69] wl[70] vdd gnd cell_6t
Xbit_r71_c69 bl[69] br[69] wl[71] vdd gnd cell_6t
Xbit_r72_c69 bl[69] br[69] wl[72] vdd gnd cell_6t
Xbit_r73_c69 bl[69] br[69] wl[73] vdd gnd cell_6t
Xbit_r74_c69 bl[69] br[69] wl[74] vdd gnd cell_6t
Xbit_r75_c69 bl[69] br[69] wl[75] vdd gnd cell_6t
Xbit_r76_c69 bl[69] br[69] wl[76] vdd gnd cell_6t
Xbit_r77_c69 bl[69] br[69] wl[77] vdd gnd cell_6t
Xbit_r78_c69 bl[69] br[69] wl[78] vdd gnd cell_6t
Xbit_r79_c69 bl[69] br[69] wl[79] vdd gnd cell_6t
Xbit_r80_c69 bl[69] br[69] wl[80] vdd gnd cell_6t
Xbit_r81_c69 bl[69] br[69] wl[81] vdd gnd cell_6t
Xbit_r82_c69 bl[69] br[69] wl[82] vdd gnd cell_6t
Xbit_r83_c69 bl[69] br[69] wl[83] vdd gnd cell_6t
Xbit_r84_c69 bl[69] br[69] wl[84] vdd gnd cell_6t
Xbit_r85_c69 bl[69] br[69] wl[85] vdd gnd cell_6t
Xbit_r86_c69 bl[69] br[69] wl[86] vdd gnd cell_6t
Xbit_r87_c69 bl[69] br[69] wl[87] vdd gnd cell_6t
Xbit_r88_c69 bl[69] br[69] wl[88] vdd gnd cell_6t
Xbit_r89_c69 bl[69] br[69] wl[89] vdd gnd cell_6t
Xbit_r90_c69 bl[69] br[69] wl[90] vdd gnd cell_6t
Xbit_r91_c69 bl[69] br[69] wl[91] vdd gnd cell_6t
Xbit_r92_c69 bl[69] br[69] wl[92] vdd gnd cell_6t
Xbit_r93_c69 bl[69] br[69] wl[93] vdd gnd cell_6t
Xbit_r94_c69 bl[69] br[69] wl[94] vdd gnd cell_6t
Xbit_r95_c69 bl[69] br[69] wl[95] vdd gnd cell_6t
Xbit_r96_c69 bl[69] br[69] wl[96] vdd gnd cell_6t
Xbit_r97_c69 bl[69] br[69] wl[97] vdd gnd cell_6t
Xbit_r98_c69 bl[69] br[69] wl[98] vdd gnd cell_6t
Xbit_r99_c69 bl[69] br[69] wl[99] vdd gnd cell_6t
Xbit_r100_c69 bl[69] br[69] wl[100] vdd gnd cell_6t
Xbit_r101_c69 bl[69] br[69] wl[101] vdd gnd cell_6t
Xbit_r102_c69 bl[69] br[69] wl[102] vdd gnd cell_6t
Xbit_r103_c69 bl[69] br[69] wl[103] vdd gnd cell_6t
Xbit_r104_c69 bl[69] br[69] wl[104] vdd gnd cell_6t
Xbit_r105_c69 bl[69] br[69] wl[105] vdd gnd cell_6t
Xbit_r106_c69 bl[69] br[69] wl[106] vdd gnd cell_6t
Xbit_r107_c69 bl[69] br[69] wl[107] vdd gnd cell_6t
Xbit_r108_c69 bl[69] br[69] wl[108] vdd gnd cell_6t
Xbit_r109_c69 bl[69] br[69] wl[109] vdd gnd cell_6t
Xbit_r110_c69 bl[69] br[69] wl[110] vdd gnd cell_6t
Xbit_r111_c69 bl[69] br[69] wl[111] vdd gnd cell_6t
Xbit_r112_c69 bl[69] br[69] wl[112] vdd gnd cell_6t
Xbit_r113_c69 bl[69] br[69] wl[113] vdd gnd cell_6t
Xbit_r114_c69 bl[69] br[69] wl[114] vdd gnd cell_6t
Xbit_r115_c69 bl[69] br[69] wl[115] vdd gnd cell_6t
Xbit_r116_c69 bl[69] br[69] wl[116] vdd gnd cell_6t
Xbit_r117_c69 bl[69] br[69] wl[117] vdd gnd cell_6t
Xbit_r118_c69 bl[69] br[69] wl[118] vdd gnd cell_6t
Xbit_r119_c69 bl[69] br[69] wl[119] vdd gnd cell_6t
Xbit_r120_c69 bl[69] br[69] wl[120] vdd gnd cell_6t
Xbit_r121_c69 bl[69] br[69] wl[121] vdd gnd cell_6t
Xbit_r122_c69 bl[69] br[69] wl[122] vdd gnd cell_6t
Xbit_r123_c69 bl[69] br[69] wl[123] vdd gnd cell_6t
Xbit_r124_c69 bl[69] br[69] wl[124] vdd gnd cell_6t
Xbit_r125_c69 bl[69] br[69] wl[125] vdd gnd cell_6t
Xbit_r126_c69 bl[69] br[69] wl[126] vdd gnd cell_6t
Xbit_r127_c69 bl[69] br[69] wl[127] vdd gnd cell_6t
Xbit_r128_c69 bl[69] br[69] wl[128] vdd gnd cell_6t
Xbit_r129_c69 bl[69] br[69] wl[129] vdd gnd cell_6t
Xbit_r130_c69 bl[69] br[69] wl[130] vdd gnd cell_6t
Xbit_r131_c69 bl[69] br[69] wl[131] vdd gnd cell_6t
Xbit_r132_c69 bl[69] br[69] wl[132] vdd gnd cell_6t
Xbit_r133_c69 bl[69] br[69] wl[133] vdd gnd cell_6t
Xbit_r134_c69 bl[69] br[69] wl[134] vdd gnd cell_6t
Xbit_r135_c69 bl[69] br[69] wl[135] vdd gnd cell_6t
Xbit_r136_c69 bl[69] br[69] wl[136] vdd gnd cell_6t
Xbit_r137_c69 bl[69] br[69] wl[137] vdd gnd cell_6t
Xbit_r138_c69 bl[69] br[69] wl[138] vdd gnd cell_6t
Xbit_r139_c69 bl[69] br[69] wl[139] vdd gnd cell_6t
Xbit_r140_c69 bl[69] br[69] wl[140] vdd gnd cell_6t
Xbit_r141_c69 bl[69] br[69] wl[141] vdd gnd cell_6t
Xbit_r142_c69 bl[69] br[69] wl[142] vdd gnd cell_6t
Xbit_r143_c69 bl[69] br[69] wl[143] vdd gnd cell_6t
Xbit_r144_c69 bl[69] br[69] wl[144] vdd gnd cell_6t
Xbit_r145_c69 bl[69] br[69] wl[145] vdd gnd cell_6t
Xbit_r146_c69 bl[69] br[69] wl[146] vdd gnd cell_6t
Xbit_r147_c69 bl[69] br[69] wl[147] vdd gnd cell_6t
Xbit_r148_c69 bl[69] br[69] wl[148] vdd gnd cell_6t
Xbit_r149_c69 bl[69] br[69] wl[149] vdd gnd cell_6t
Xbit_r150_c69 bl[69] br[69] wl[150] vdd gnd cell_6t
Xbit_r151_c69 bl[69] br[69] wl[151] vdd gnd cell_6t
Xbit_r152_c69 bl[69] br[69] wl[152] vdd gnd cell_6t
Xbit_r153_c69 bl[69] br[69] wl[153] vdd gnd cell_6t
Xbit_r154_c69 bl[69] br[69] wl[154] vdd gnd cell_6t
Xbit_r155_c69 bl[69] br[69] wl[155] vdd gnd cell_6t
Xbit_r156_c69 bl[69] br[69] wl[156] vdd gnd cell_6t
Xbit_r157_c69 bl[69] br[69] wl[157] vdd gnd cell_6t
Xbit_r158_c69 bl[69] br[69] wl[158] vdd gnd cell_6t
Xbit_r159_c69 bl[69] br[69] wl[159] vdd gnd cell_6t
Xbit_r160_c69 bl[69] br[69] wl[160] vdd gnd cell_6t
Xbit_r161_c69 bl[69] br[69] wl[161] vdd gnd cell_6t
Xbit_r162_c69 bl[69] br[69] wl[162] vdd gnd cell_6t
Xbit_r163_c69 bl[69] br[69] wl[163] vdd gnd cell_6t
Xbit_r164_c69 bl[69] br[69] wl[164] vdd gnd cell_6t
Xbit_r165_c69 bl[69] br[69] wl[165] vdd gnd cell_6t
Xbit_r166_c69 bl[69] br[69] wl[166] vdd gnd cell_6t
Xbit_r167_c69 bl[69] br[69] wl[167] vdd gnd cell_6t
Xbit_r168_c69 bl[69] br[69] wl[168] vdd gnd cell_6t
Xbit_r169_c69 bl[69] br[69] wl[169] vdd gnd cell_6t
Xbit_r170_c69 bl[69] br[69] wl[170] vdd gnd cell_6t
Xbit_r171_c69 bl[69] br[69] wl[171] vdd gnd cell_6t
Xbit_r172_c69 bl[69] br[69] wl[172] vdd gnd cell_6t
Xbit_r173_c69 bl[69] br[69] wl[173] vdd gnd cell_6t
Xbit_r174_c69 bl[69] br[69] wl[174] vdd gnd cell_6t
Xbit_r175_c69 bl[69] br[69] wl[175] vdd gnd cell_6t
Xbit_r176_c69 bl[69] br[69] wl[176] vdd gnd cell_6t
Xbit_r177_c69 bl[69] br[69] wl[177] vdd gnd cell_6t
Xbit_r178_c69 bl[69] br[69] wl[178] vdd gnd cell_6t
Xbit_r179_c69 bl[69] br[69] wl[179] vdd gnd cell_6t
Xbit_r180_c69 bl[69] br[69] wl[180] vdd gnd cell_6t
Xbit_r181_c69 bl[69] br[69] wl[181] vdd gnd cell_6t
Xbit_r182_c69 bl[69] br[69] wl[182] vdd gnd cell_6t
Xbit_r183_c69 bl[69] br[69] wl[183] vdd gnd cell_6t
Xbit_r184_c69 bl[69] br[69] wl[184] vdd gnd cell_6t
Xbit_r185_c69 bl[69] br[69] wl[185] vdd gnd cell_6t
Xbit_r186_c69 bl[69] br[69] wl[186] vdd gnd cell_6t
Xbit_r187_c69 bl[69] br[69] wl[187] vdd gnd cell_6t
Xbit_r188_c69 bl[69] br[69] wl[188] vdd gnd cell_6t
Xbit_r189_c69 bl[69] br[69] wl[189] vdd gnd cell_6t
Xbit_r190_c69 bl[69] br[69] wl[190] vdd gnd cell_6t
Xbit_r191_c69 bl[69] br[69] wl[191] vdd gnd cell_6t
Xbit_r192_c69 bl[69] br[69] wl[192] vdd gnd cell_6t
Xbit_r193_c69 bl[69] br[69] wl[193] vdd gnd cell_6t
Xbit_r194_c69 bl[69] br[69] wl[194] vdd gnd cell_6t
Xbit_r195_c69 bl[69] br[69] wl[195] vdd gnd cell_6t
Xbit_r196_c69 bl[69] br[69] wl[196] vdd gnd cell_6t
Xbit_r197_c69 bl[69] br[69] wl[197] vdd gnd cell_6t
Xbit_r198_c69 bl[69] br[69] wl[198] vdd gnd cell_6t
Xbit_r199_c69 bl[69] br[69] wl[199] vdd gnd cell_6t
Xbit_r200_c69 bl[69] br[69] wl[200] vdd gnd cell_6t
Xbit_r201_c69 bl[69] br[69] wl[201] vdd gnd cell_6t
Xbit_r202_c69 bl[69] br[69] wl[202] vdd gnd cell_6t
Xbit_r203_c69 bl[69] br[69] wl[203] vdd gnd cell_6t
Xbit_r204_c69 bl[69] br[69] wl[204] vdd gnd cell_6t
Xbit_r205_c69 bl[69] br[69] wl[205] vdd gnd cell_6t
Xbit_r206_c69 bl[69] br[69] wl[206] vdd gnd cell_6t
Xbit_r207_c69 bl[69] br[69] wl[207] vdd gnd cell_6t
Xbit_r208_c69 bl[69] br[69] wl[208] vdd gnd cell_6t
Xbit_r209_c69 bl[69] br[69] wl[209] vdd gnd cell_6t
Xbit_r210_c69 bl[69] br[69] wl[210] vdd gnd cell_6t
Xbit_r211_c69 bl[69] br[69] wl[211] vdd gnd cell_6t
Xbit_r212_c69 bl[69] br[69] wl[212] vdd gnd cell_6t
Xbit_r213_c69 bl[69] br[69] wl[213] vdd gnd cell_6t
Xbit_r214_c69 bl[69] br[69] wl[214] vdd gnd cell_6t
Xbit_r215_c69 bl[69] br[69] wl[215] vdd gnd cell_6t
Xbit_r216_c69 bl[69] br[69] wl[216] vdd gnd cell_6t
Xbit_r217_c69 bl[69] br[69] wl[217] vdd gnd cell_6t
Xbit_r218_c69 bl[69] br[69] wl[218] vdd gnd cell_6t
Xbit_r219_c69 bl[69] br[69] wl[219] vdd gnd cell_6t
Xbit_r220_c69 bl[69] br[69] wl[220] vdd gnd cell_6t
Xbit_r221_c69 bl[69] br[69] wl[221] vdd gnd cell_6t
Xbit_r222_c69 bl[69] br[69] wl[222] vdd gnd cell_6t
Xbit_r223_c69 bl[69] br[69] wl[223] vdd gnd cell_6t
Xbit_r224_c69 bl[69] br[69] wl[224] vdd gnd cell_6t
Xbit_r225_c69 bl[69] br[69] wl[225] vdd gnd cell_6t
Xbit_r226_c69 bl[69] br[69] wl[226] vdd gnd cell_6t
Xbit_r227_c69 bl[69] br[69] wl[227] vdd gnd cell_6t
Xbit_r228_c69 bl[69] br[69] wl[228] vdd gnd cell_6t
Xbit_r229_c69 bl[69] br[69] wl[229] vdd gnd cell_6t
Xbit_r230_c69 bl[69] br[69] wl[230] vdd gnd cell_6t
Xbit_r231_c69 bl[69] br[69] wl[231] vdd gnd cell_6t
Xbit_r232_c69 bl[69] br[69] wl[232] vdd gnd cell_6t
Xbit_r233_c69 bl[69] br[69] wl[233] vdd gnd cell_6t
Xbit_r234_c69 bl[69] br[69] wl[234] vdd gnd cell_6t
Xbit_r235_c69 bl[69] br[69] wl[235] vdd gnd cell_6t
Xbit_r236_c69 bl[69] br[69] wl[236] vdd gnd cell_6t
Xbit_r237_c69 bl[69] br[69] wl[237] vdd gnd cell_6t
Xbit_r238_c69 bl[69] br[69] wl[238] vdd gnd cell_6t
Xbit_r239_c69 bl[69] br[69] wl[239] vdd gnd cell_6t
Xbit_r240_c69 bl[69] br[69] wl[240] vdd gnd cell_6t
Xbit_r241_c69 bl[69] br[69] wl[241] vdd gnd cell_6t
Xbit_r242_c69 bl[69] br[69] wl[242] vdd gnd cell_6t
Xbit_r243_c69 bl[69] br[69] wl[243] vdd gnd cell_6t
Xbit_r244_c69 bl[69] br[69] wl[244] vdd gnd cell_6t
Xbit_r245_c69 bl[69] br[69] wl[245] vdd gnd cell_6t
Xbit_r246_c69 bl[69] br[69] wl[246] vdd gnd cell_6t
Xbit_r247_c69 bl[69] br[69] wl[247] vdd gnd cell_6t
Xbit_r248_c69 bl[69] br[69] wl[248] vdd gnd cell_6t
Xbit_r249_c69 bl[69] br[69] wl[249] vdd gnd cell_6t
Xbit_r250_c69 bl[69] br[69] wl[250] vdd gnd cell_6t
Xbit_r251_c69 bl[69] br[69] wl[251] vdd gnd cell_6t
Xbit_r252_c69 bl[69] br[69] wl[252] vdd gnd cell_6t
Xbit_r253_c69 bl[69] br[69] wl[253] vdd gnd cell_6t
Xbit_r254_c69 bl[69] br[69] wl[254] vdd gnd cell_6t
Xbit_r255_c69 bl[69] br[69] wl[255] vdd gnd cell_6t
Xbit_r256_c69 bl[69] br[69] wl[256] vdd gnd cell_6t
Xbit_r257_c69 bl[69] br[69] wl[257] vdd gnd cell_6t
Xbit_r258_c69 bl[69] br[69] wl[258] vdd gnd cell_6t
Xbit_r259_c69 bl[69] br[69] wl[259] vdd gnd cell_6t
Xbit_r260_c69 bl[69] br[69] wl[260] vdd gnd cell_6t
Xbit_r261_c69 bl[69] br[69] wl[261] vdd gnd cell_6t
Xbit_r262_c69 bl[69] br[69] wl[262] vdd gnd cell_6t
Xbit_r263_c69 bl[69] br[69] wl[263] vdd gnd cell_6t
Xbit_r264_c69 bl[69] br[69] wl[264] vdd gnd cell_6t
Xbit_r265_c69 bl[69] br[69] wl[265] vdd gnd cell_6t
Xbit_r266_c69 bl[69] br[69] wl[266] vdd gnd cell_6t
Xbit_r267_c69 bl[69] br[69] wl[267] vdd gnd cell_6t
Xbit_r268_c69 bl[69] br[69] wl[268] vdd gnd cell_6t
Xbit_r269_c69 bl[69] br[69] wl[269] vdd gnd cell_6t
Xbit_r270_c69 bl[69] br[69] wl[270] vdd gnd cell_6t
Xbit_r271_c69 bl[69] br[69] wl[271] vdd gnd cell_6t
Xbit_r272_c69 bl[69] br[69] wl[272] vdd gnd cell_6t
Xbit_r273_c69 bl[69] br[69] wl[273] vdd gnd cell_6t
Xbit_r274_c69 bl[69] br[69] wl[274] vdd gnd cell_6t
Xbit_r275_c69 bl[69] br[69] wl[275] vdd gnd cell_6t
Xbit_r276_c69 bl[69] br[69] wl[276] vdd gnd cell_6t
Xbit_r277_c69 bl[69] br[69] wl[277] vdd gnd cell_6t
Xbit_r278_c69 bl[69] br[69] wl[278] vdd gnd cell_6t
Xbit_r279_c69 bl[69] br[69] wl[279] vdd gnd cell_6t
Xbit_r280_c69 bl[69] br[69] wl[280] vdd gnd cell_6t
Xbit_r281_c69 bl[69] br[69] wl[281] vdd gnd cell_6t
Xbit_r282_c69 bl[69] br[69] wl[282] vdd gnd cell_6t
Xbit_r283_c69 bl[69] br[69] wl[283] vdd gnd cell_6t
Xbit_r284_c69 bl[69] br[69] wl[284] vdd gnd cell_6t
Xbit_r285_c69 bl[69] br[69] wl[285] vdd gnd cell_6t
Xbit_r286_c69 bl[69] br[69] wl[286] vdd gnd cell_6t
Xbit_r287_c69 bl[69] br[69] wl[287] vdd gnd cell_6t
Xbit_r288_c69 bl[69] br[69] wl[288] vdd gnd cell_6t
Xbit_r289_c69 bl[69] br[69] wl[289] vdd gnd cell_6t
Xbit_r290_c69 bl[69] br[69] wl[290] vdd gnd cell_6t
Xbit_r291_c69 bl[69] br[69] wl[291] vdd gnd cell_6t
Xbit_r292_c69 bl[69] br[69] wl[292] vdd gnd cell_6t
Xbit_r293_c69 bl[69] br[69] wl[293] vdd gnd cell_6t
Xbit_r294_c69 bl[69] br[69] wl[294] vdd gnd cell_6t
Xbit_r295_c69 bl[69] br[69] wl[295] vdd gnd cell_6t
Xbit_r296_c69 bl[69] br[69] wl[296] vdd gnd cell_6t
Xbit_r297_c69 bl[69] br[69] wl[297] vdd gnd cell_6t
Xbit_r298_c69 bl[69] br[69] wl[298] vdd gnd cell_6t
Xbit_r299_c69 bl[69] br[69] wl[299] vdd gnd cell_6t
Xbit_r300_c69 bl[69] br[69] wl[300] vdd gnd cell_6t
Xbit_r301_c69 bl[69] br[69] wl[301] vdd gnd cell_6t
Xbit_r302_c69 bl[69] br[69] wl[302] vdd gnd cell_6t
Xbit_r303_c69 bl[69] br[69] wl[303] vdd gnd cell_6t
Xbit_r304_c69 bl[69] br[69] wl[304] vdd gnd cell_6t
Xbit_r305_c69 bl[69] br[69] wl[305] vdd gnd cell_6t
Xbit_r306_c69 bl[69] br[69] wl[306] vdd gnd cell_6t
Xbit_r307_c69 bl[69] br[69] wl[307] vdd gnd cell_6t
Xbit_r308_c69 bl[69] br[69] wl[308] vdd gnd cell_6t
Xbit_r309_c69 bl[69] br[69] wl[309] vdd gnd cell_6t
Xbit_r310_c69 bl[69] br[69] wl[310] vdd gnd cell_6t
Xbit_r311_c69 bl[69] br[69] wl[311] vdd gnd cell_6t
Xbit_r312_c69 bl[69] br[69] wl[312] vdd gnd cell_6t
Xbit_r313_c69 bl[69] br[69] wl[313] vdd gnd cell_6t
Xbit_r314_c69 bl[69] br[69] wl[314] vdd gnd cell_6t
Xbit_r315_c69 bl[69] br[69] wl[315] vdd gnd cell_6t
Xbit_r316_c69 bl[69] br[69] wl[316] vdd gnd cell_6t
Xbit_r317_c69 bl[69] br[69] wl[317] vdd gnd cell_6t
Xbit_r318_c69 bl[69] br[69] wl[318] vdd gnd cell_6t
Xbit_r319_c69 bl[69] br[69] wl[319] vdd gnd cell_6t
Xbit_r320_c69 bl[69] br[69] wl[320] vdd gnd cell_6t
Xbit_r321_c69 bl[69] br[69] wl[321] vdd gnd cell_6t
Xbit_r322_c69 bl[69] br[69] wl[322] vdd gnd cell_6t
Xbit_r323_c69 bl[69] br[69] wl[323] vdd gnd cell_6t
Xbit_r324_c69 bl[69] br[69] wl[324] vdd gnd cell_6t
Xbit_r325_c69 bl[69] br[69] wl[325] vdd gnd cell_6t
Xbit_r326_c69 bl[69] br[69] wl[326] vdd gnd cell_6t
Xbit_r327_c69 bl[69] br[69] wl[327] vdd gnd cell_6t
Xbit_r328_c69 bl[69] br[69] wl[328] vdd gnd cell_6t
Xbit_r329_c69 bl[69] br[69] wl[329] vdd gnd cell_6t
Xbit_r330_c69 bl[69] br[69] wl[330] vdd gnd cell_6t
Xbit_r331_c69 bl[69] br[69] wl[331] vdd gnd cell_6t
Xbit_r332_c69 bl[69] br[69] wl[332] vdd gnd cell_6t
Xbit_r333_c69 bl[69] br[69] wl[333] vdd gnd cell_6t
Xbit_r334_c69 bl[69] br[69] wl[334] vdd gnd cell_6t
Xbit_r335_c69 bl[69] br[69] wl[335] vdd gnd cell_6t
Xbit_r336_c69 bl[69] br[69] wl[336] vdd gnd cell_6t
Xbit_r337_c69 bl[69] br[69] wl[337] vdd gnd cell_6t
Xbit_r338_c69 bl[69] br[69] wl[338] vdd gnd cell_6t
Xbit_r339_c69 bl[69] br[69] wl[339] vdd gnd cell_6t
Xbit_r340_c69 bl[69] br[69] wl[340] vdd gnd cell_6t
Xbit_r341_c69 bl[69] br[69] wl[341] vdd gnd cell_6t
Xbit_r342_c69 bl[69] br[69] wl[342] vdd gnd cell_6t
Xbit_r343_c69 bl[69] br[69] wl[343] vdd gnd cell_6t
Xbit_r344_c69 bl[69] br[69] wl[344] vdd gnd cell_6t
Xbit_r345_c69 bl[69] br[69] wl[345] vdd gnd cell_6t
Xbit_r346_c69 bl[69] br[69] wl[346] vdd gnd cell_6t
Xbit_r347_c69 bl[69] br[69] wl[347] vdd gnd cell_6t
Xbit_r348_c69 bl[69] br[69] wl[348] vdd gnd cell_6t
Xbit_r349_c69 bl[69] br[69] wl[349] vdd gnd cell_6t
Xbit_r350_c69 bl[69] br[69] wl[350] vdd gnd cell_6t
Xbit_r351_c69 bl[69] br[69] wl[351] vdd gnd cell_6t
Xbit_r352_c69 bl[69] br[69] wl[352] vdd gnd cell_6t
Xbit_r353_c69 bl[69] br[69] wl[353] vdd gnd cell_6t
Xbit_r354_c69 bl[69] br[69] wl[354] vdd gnd cell_6t
Xbit_r355_c69 bl[69] br[69] wl[355] vdd gnd cell_6t
Xbit_r356_c69 bl[69] br[69] wl[356] vdd gnd cell_6t
Xbit_r357_c69 bl[69] br[69] wl[357] vdd gnd cell_6t
Xbit_r358_c69 bl[69] br[69] wl[358] vdd gnd cell_6t
Xbit_r359_c69 bl[69] br[69] wl[359] vdd gnd cell_6t
Xbit_r360_c69 bl[69] br[69] wl[360] vdd gnd cell_6t
Xbit_r361_c69 bl[69] br[69] wl[361] vdd gnd cell_6t
Xbit_r362_c69 bl[69] br[69] wl[362] vdd gnd cell_6t
Xbit_r363_c69 bl[69] br[69] wl[363] vdd gnd cell_6t
Xbit_r364_c69 bl[69] br[69] wl[364] vdd gnd cell_6t
Xbit_r365_c69 bl[69] br[69] wl[365] vdd gnd cell_6t
Xbit_r366_c69 bl[69] br[69] wl[366] vdd gnd cell_6t
Xbit_r367_c69 bl[69] br[69] wl[367] vdd gnd cell_6t
Xbit_r368_c69 bl[69] br[69] wl[368] vdd gnd cell_6t
Xbit_r369_c69 bl[69] br[69] wl[369] vdd gnd cell_6t
Xbit_r370_c69 bl[69] br[69] wl[370] vdd gnd cell_6t
Xbit_r371_c69 bl[69] br[69] wl[371] vdd gnd cell_6t
Xbit_r372_c69 bl[69] br[69] wl[372] vdd gnd cell_6t
Xbit_r373_c69 bl[69] br[69] wl[373] vdd gnd cell_6t
Xbit_r374_c69 bl[69] br[69] wl[374] vdd gnd cell_6t
Xbit_r375_c69 bl[69] br[69] wl[375] vdd gnd cell_6t
Xbit_r376_c69 bl[69] br[69] wl[376] vdd gnd cell_6t
Xbit_r377_c69 bl[69] br[69] wl[377] vdd gnd cell_6t
Xbit_r378_c69 bl[69] br[69] wl[378] vdd gnd cell_6t
Xbit_r379_c69 bl[69] br[69] wl[379] vdd gnd cell_6t
Xbit_r380_c69 bl[69] br[69] wl[380] vdd gnd cell_6t
Xbit_r381_c69 bl[69] br[69] wl[381] vdd gnd cell_6t
Xbit_r382_c69 bl[69] br[69] wl[382] vdd gnd cell_6t
Xbit_r383_c69 bl[69] br[69] wl[383] vdd gnd cell_6t
Xbit_r384_c69 bl[69] br[69] wl[384] vdd gnd cell_6t
Xbit_r385_c69 bl[69] br[69] wl[385] vdd gnd cell_6t
Xbit_r386_c69 bl[69] br[69] wl[386] vdd gnd cell_6t
Xbit_r387_c69 bl[69] br[69] wl[387] vdd gnd cell_6t
Xbit_r388_c69 bl[69] br[69] wl[388] vdd gnd cell_6t
Xbit_r389_c69 bl[69] br[69] wl[389] vdd gnd cell_6t
Xbit_r390_c69 bl[69] br[69] wl[390] vdd gnd cell_6t
Xbit_r391_c69 bl[69] br[69] wl[391] vdd gnd cell_6t
Xbit_r392_c69 bl[69] br[69] wl[392] vdd gnd cell_6t
Xbit_r393_c69 bl[69] br[69] wl[393] vdd gnd cell_6t
Xbit_r394_c69 bl[69] br[69] wl[394] vdd gnd cell_6t
Xbit_r395_c69 bl[69] br[69] wl[395] vdd gnd cell_6t
Xbit_r396_c69 bl[69] br[69] wl[396] vdd gnd cell_6t
Xbit_r397_c69 bl[69] br[69] wl[397] vdd gnd cell_6t
Xbit_r398_c69 bl[69] br[69] wl[398] vdd gnd cell_6t
Xbit_r399_c69 bl[69] br[69] wl[399] vdd gnd cell_6t
Xbit_r400_c69 bl[69] br[69] wl[400] vdd gnd cell_6t
Xbit_r401_c69 bl[69] br[69] wl[401] vdd gnd cell_6t
Xbit_r402_c69 bl[69] br[69] wl[402] vdd gnd cell_6t
Xbit_r403_c69 bl[69] br[69] wl[403] vdd gnd cell_6t
Xbit_r404_c69 bl[69] br[69] wl[404] vdd gnd cell_6t
Xbit_r405_c69 bl[69] br[69] wl[405] vdd gnd cell_6t
Xbit_r406_c69 bl[69] br[69] wl[406] vdd gnd cell_6t
Xbit_r407_c69 bl[69] br[69] wl[407] vdd gnd cell_6t
Xbit_r408_c69 bl[69] br[69] wl[408] vdd gnd cell_6t
Xbit_r409_c69 bl[69] br[69] wl[409] vdd gnd cell_6t
Xbit_r410_c69 bl[69] br[69] wl[410] vdd gnd cell_6t
Xbit_r411_c69 bl[69] br[69] wl[411] vdd gnd cell_6t
Xbit_r412_c69 bl[69] br[69] wl[412] vdd gnd cell_6t
Xbit_r413_c69 bl[69] br[69] wl[413] vdd gnd cell_6t
Xbit_r414_c69 bl[69] br[69] wl[414] vdd gnd cell_6t
Xbit_r415_c69 bl[69] br[69] wl[415] vdd gnd cell_6t
Xbit_r416_c69 bl[69] br[69] wl[416] vdd gnd cell_6t
Xbit_r417_c69 bl[69] br[69] wl[417] vdd gnd cell_6t
Xbit_r418_c69 bl[69] br[69] wl[418] vdd gnd cell_6t
Xbit_r419_c69 bl[69] br[69] wl[419] vdd gnd cell_6t
Xbit_r420_c69 bl[69] br[69] wl[420] vdd gnd cell_6t
Xbit_r421_c69 bl[69] br[69] wl[421] vdd gnd cell_6t
Xbit_r422_c69 bl[69] br[69] wl[422] vdd gnd cell_6t
Xbit_r423_c69 bl[69] br[69] wl[423] vdd gnd cell_6t
Xbit_r424_c69 bl[69] br[69] wl[424] vdd gnd cell_6t
Xbit_r425_c69 bl[69] br[69] wl[425] vdd gnd cell_6t
Xbit_r426_c69 bl[69] br[69] wl[426] vdd gnd cell_6t
Xbit_r427_c69 bl[69] br[69] wl[427] vdd gnd cell_6t
Xbit_r428_c69 bl[69] br[69] wl[428] vdd gnd cell_6t
Xbit_r429_c69 bl[69] br[69] wl[429] vdd gnd cell_6t
Xbit_r430_c69 bl[69] br[69] wl[430] vdd gnd cell_6t
Xbit_r431_c69 bl[69] br[69] wl[431] vdd gnd cell_6t
Xbit_r432_c69 bl[69] br[69] wl[432] vdd gnd cell_6t
Xbit_r433_c69 bl[69] br[69] wl[433] vdd gnd cell_6t
Xbit_r434_c69 bl[69] br[69] wl[434] vdd gnd cell_6t
Xbit_r435_c69 bl[69] br[69] wl[435] vdd gnd cell_6t
Xbit_r436_c69 bl[69] br[69] wl[436] vdd gnd cell_6t
Xbit_r437_c69 bl[69] br[69] wl[437] vdd gnd cell_6t
Xbit_r438_c69 bl[69] br[69] wl[438] vdd gnd cell_6t
Xbit_r439_c69 bl[69] br[69] wl[439] vdd gnd cell_6t
Xbit_r440_c69 bl[69] br[69] wl[440] vdd gnd cell_6t
Xbit_r441_c69 bl[69] br[69] wl[441] vdd gnd cell_6t
Xbit_r442_c69 bl[69] br[69] wl[442] vdd gnd cell_6t
Xbit_r443_c69 bl[69] br[69] wl[443] vdd gnd cell_6t
Xbit_r444_c69 bl[69] br[69] wl[444] vdd gnd cell_6t
Xbit_r445_c69 bl[69] br[69] wl[445] vdd gnd cell_6t
Xbit_r446_c69 bl[69] br[69] wl[446] vdd gnd cell_6t
Xbit_r447_c69 bl[69] br[69] wl[447] vdd gnd cell_6t
Xbit_r448_c69 bl[69] br[69] wl[448] vdd gnd cell_6t
Xbit_r449_c69 bl[69] br[69] wl[449] vdd gnd cell_6t
Xbit_r450_c69 bl[69] br[69] wl[450] vdd gnd cell_6t
Xbit_r451_c69 bl[69] br[69] wl[451] vdd gnd cell_6t
Xbit_r452_c69 bl[69] br[69] wl[452] vdd gnd cell_6t
Xbit_r453_c69 bl[69] br[69] wl[453] vdd gnd cell_6t
Xbit_r454_c69 bl[69] br[69] wl[454] vdd gnd cell_6t
Xbit_r455_c69 bl[69] br[69] wl[455] vdd gnd cell_6t
Xbit_r456_c69 bl[69] br[69] wl[456] vdd gnd cell_6t
Xbit_r457_c69 bl[69] br[69] wl[457] vdd gnd cell_6t
Xbit_r458_c69 bl[69] br[69] wl[458] vdd gnd cell_6t
Xbit_r459_c69 bl[69] br[69] wl[459] vdd gnd cell_6t
Xbit_r460_c69 bl[69] br[69] wl[460] vdd gnd cell_6t
Xbit_r461_c69 bl[69] br[69] wl[461] vdd gnd cell_6t
Xbit_r462_c69 bl[69] br[69] wl[462] vdd gnd cell_6t
Xbit_r463_c69 bl[69] br[69] wl[463] vdd gnd cell_6t
Xbit_r464_c69 bl[69] br[69] wl[464] vdd gnd cell_6t
Xbit_r465_c69 bl[69] br[69] wl[465] vdd gnd cell_6t
Xbit_r466_c69 bl[69] br[69] wl[466] vdd gnd cell_6t
Xbit_r467_c69 bl[69] br[69] wl[467] vdd gnd cell_6t
Xbit_r468_c69 bl[69] br[69] wl[468] vdd gnd cell_6t
Xbit_r469_c69 bl[69] br[69] wl[469] vdd gnd cell_6t
Xbit_r470_c69 bl[69] br[69] wl[470] vdd gnd cell_6t
Xbit_r471_c69 bl[69] br[69] wl[471] vdd gnd cell_6t
Xbit_r472_c69 bl[69] br[69] wl[472] vdd gnd cell_6t
Xbit_r473_c69 bl[69] br[69] wl[473] vdd gnd cell_6t
Xbit_r474_c69 bl[69] br[69] wl[474] vdd gnd cell_6t
Xbit_r475_c69 bl[69] br[69] wl[475] vdd gnd cell_6t
Xbit_r476_c69 bl[69] br[69] wl[476] vdd gnd cell_6t
Xbit_r477_c69 bl[69] br[69] wl[477] vdd gnd cell_6t
Xbit_r478_c69 bl[69] br[69] wl[478] vdd gnd cell_6t
Xbit_r479_c69 bl[69] br[69] wl[479] vdd gnd cell_6t
Xbit_r480_c69 bl[69] br[69] wl[480] vdd gnd cell_6t
Xbit_r481_c69 bl[69] br[69] wl[481] vdd gnd cell_6t
Xbit_r482_c69 bl[69] br[69] wl[482] vdd gnd cell_6t
Xbit_r483_c69 bl[69] br[69] wl[483] vdd gnd cell_6t
Xbit_r484_c69 bl[69] br[69] wl[484] vdd gnd cell_6t
Xbit_r485_c69 bl[69] br[69] wl[485] vdd gnd cell_6t
Xbit_r486_c69 bl[69] br[69] wl[486] vdd gnd cell_6t
Xbit_r487_c69 bl[69] br[69] wl[487] vdd gnd cell_6t
Xbit_r488_c69 bl[69] br[69] wl[488] vdd gnd cell_6t
Xbit_r489_c69 bl[69] br[69] wl[489] vdd gnd cell_6t
Xbit_r490_c69 bl[69] br[69] wl[490] vdd gnd cell_6t
Xbit_r491_c69 bl[69] br[69] wl[491] vdd gnd cell_6t
Xbit_r492_c69 bl[69] br[69] wl[492] vdd gnd cell_6t
Xbit_r493_c69 bl[69] br[69] wl[493] vdd gnd cell_6t
Xbit_r494_c69 bl[69] br[69] wl[494] vdd gnd cell_6t
Xbit_r495_c69 bl[69] br[69] wl[495] vdd gnd cell_6t
Xbit_r496_c69 bl[69] br[69] wl[496] vdd gnd cell_6t
Xbit_r497_c69 bl[69] br[69] wl[497] vdd gnd cell_6t
Xbit_r498_c69 bl[69] br[69] wl[498] vdd gnd cell_6t
Xbit_r499_c69 bl[69] br[69] wl[499] vdd gnd cell_6t
Xbit_r500_c69 bl[69] br[69] wl[500] vdd gnd cell_6t
Xbit_r501_c69 bl[69] br[69] wl[501] vdd gnd cell_6t
Xbit_r502_c69 bl[69] br[69] wl[502] vdd gnd cell_6t
Xbit_r503_c69 bl[69] br[69] wl[503] vdd gnd cell_6t
Xbit_r504_c69 bl[69] br[69] wl[504] vdd gnd cell_6t
Xbit_r505_c69 bl[69] br[69] wl[505] vdd gnd cell_6t
Xbit_r506_c69 bl[69] br[69] wl[506] vdd gnd cell_6t
Xbit_r507_c69 bl[69] br[69] wl[507] vdd gnd cell_6t
Xbit_r508_c69 bl[69] br[69] wl[508] vdd gnd cell_6t
Xbit_r509_c69 bl[69] br[69] wl[509] vdd gnd cell_6t
Xbit_r510_c69 bl[69] br[69] wl[510] vdd gnd cell_6t
Xbit_r511_c69 bl[69] br[69] wl[511] vdd gnd cell_6t
Xbit_r0_c70 bl[70] br[70] wl[0] vdd gnd cell_6t
Xbit_r1_c70 bl[70] br[70] wl[1] vdd gnd cell_6t
Xbit_r2_c70 bl[70] br[70] wl[2] vdd gnd cell_6t
Xbit_r3_c70 bl[70] br[70] wl[3] vdd gnd cell_6t
Xbit_r4_c70 bl[70] br[70] wl[4] vdd gnd cell_6t
Xbit_r5_c70 bl[70] br[70] wl[5] vdd gnd cell_6t
Xbit_r6_c70 bl[70] br[70] wl[6] vdd gnd cell_6t
Xbit_r7_c70 bl[70] br[70] wl[7] vdd gnd cell_6t
Xbit_r8_c70 bl[70] br[70] wl[8] vdd gnd cell_6t
Xbit_r9_c70 bl[70] br[70] wl[9] vdd gnd cell_6t
Xbit_r10_c70 bl[70] br[70] wl[10] vdd gnd cell_6t
Xbit_r11_c70 bl[70] br[70] wl[11] vdd gnd cell_6t
Xbit_r12_c70 bl[70] br[70] wl[12] vdd gnd cell_6t
Xbit_r13_c70 bl[70] br[70] wl[13] vdd gnd cell_6t
Xbit_r14_c70 bl[70] br[70] wl[14] vdd gnd cell_6t
Xbit_r15_c70 bl[70] br[70] wl[15] vdd gnd cell_6t
Xbit_r16_c70 bl[70] br[70] wl[16] vdd gnd cell_6t
Xbit_r17_c70 bl[70] br[70] wl[17] vdd gnd cell_6t
Xbit_r18_c70 bl[70] br[70] wl[18] vdd gnd cell_6t
Xbit_r19_c70 bl[70] br[70] wl[19] vdd gnd cell_6t
Xbit_r20_c70 bl[70] br[70] wl[20] vdd gnd cell_6t
Xbit_r21_c70 bl[70] br[70] wl[21] vdd gnd cell_6t
Xbit_r22_c70 bl[70] br[70] wl[22] vdd gnd cell_6t
Xbit_r23_c70 bl[70] br[70] wl[23] vdd gnd cell_6t
Xbit_r24_c70 bl[70] br[70] wl[24] vdd gnd cell_6t
Xbit_r25_c70 bl[70] br[70] wl[25] vdd gnd cell_6t
Xbit_r26_c70 bl[70] br[70] wl[26] vdd gnd cell_6t
Xbit_r27_c70 bl[70] br[70] wl[27] vdd gnd cell_6t
Xbit_r28_c70 bl[70] br[70] wl[28] vdd gnd cell_6t
Xbit_r29_c70 bl[70] br[70] wl[29] vdd gnd cell_6t
Xbit_r30_c70 bl[70] br[70] wl[30] vdd gnd cell_6t
Xbit_r31_c70 bl[70] br[70] wl[31] vdd gnd cell_6t
Xbit_r32_c70 bl[70] br[70] wl[32] vdd gnd cell_6t
Xbit_r33_c70 bl[70] br[70] wl[33] vdd gnd cell_6t
Xbit_r34_c70 bl[70] br[70] wl[34] vdd gnd cell_6t
Xbit_r35_c70 bl[70] br[70] wl[35] vdd gnd cell_6t
Xbit_r36_c70 bl[70] br[70] wl[36] vdd gnd cell_6t
Xbit_r37_c70 bl[70] br[70] wl[37] vdd gnd cell_6t
Xbit_r38_c70 bl[70] br[70] wl[38] vdd gnd cell_6t
Xbit_r39_c70 bl[70] br[70] wl[39] vdd gnd cell_6t
Xbit_r40_c70 bl[70] br[70] wl[40] vdd gnd cell_6t
Xbit_r41_c70 bl[70] br[70] wl[41] vdd gnd cell_6t
Xbit_r42_c70 bl[70] br[70] wl[42] vdd gnd cell_6t
Xbit_r43_c70 bl[70] br[70] wl[43] vdd gnd cell_6t
Xbit_r44_c70 bl[70] br[70] wl[44] vdd gnd cell_6t
Xbit_r45_c70 bl[70] br[70] wl[45] vdd gnd cell_6t
Xbit_r46_c70 bl[70] br[70] wl[46] vdd gnd cell_6t
Xbit_r47_c70 bl[70] br[70] wl[47] vdd gnd cell_6t
Xbit_r48_c70 bl[70] br[70] wl[48] vdd gnd cell_6t
Xbit_r49_c70 bl[70] br[70] wl[49] vdd gnd cell_6t
Xbit_r50_c70 bl[70] br[70] wl[50] vdd gnd cell_6t
Xbit_r51_c70 bl[70] br[70] wl[51] vdd gnd cell_6t
Xbit_r52_c70 bl[70] br[70] wl[52] vdd gnd cell_6t
Xbit_r53_c70 bl[70] br[70] wl[53] vdd gnd cell_6t
Xbit_r54_c70 bl[70] br[70] wl[54] vdd gnd cell_6t
Xbit_r55_c70 bl[70] br[70] wl[55] vdd gnd cell_6t
Xbit_r56_c70 bl[70] br[70] wl[56] vdd gnd cell_6t
Xbit_r57_c70 bl[70] br[70] wl[57] vdd gnd cell_6t
Xbit_r58_c70 bl[70] br[70] wl[58] vdd gnd cell_6t
Xbit_r59_c70 bl[70] br[70] wl[59] vdd gnd cell_6t
Xbit_r60_c70 bl[70] br[70] wl[60] vdd gnd cell_6t
Xbit_r61_c70 bl[70] br[70] wl[61] vdd gnd cell_6t
Xbit_r62_c70 bl[70] br[70] wl[62] vdd gnd cell_6t
Xbit_r63_c70 bl[70] br[70] wl[63] vdd gnd cell_6t
Xbit_r64_c70 bl[70] br[70] wl[64] vdd gnd cell_6t
Xbit_r65_c70 bl[70] br[70] wl[65] vdd gnd cell_6t
Xbit_r66_c70 bl[70] br[70] wl[66] vdd gnd cell_6t
Xbit_r67_c70 bl[70] br[70] wl[67] vdd gnd cell_6t
Xbit_r68_c70 bl[70] br[70] wl[68] vdd gnd cell_6t
Xbit_r69_c70 bl[70] br[70] wl[69] vdd gnd cell_6t
Xbit_r70_c70 bl[70] br[70] wl[70] vdd gnd cell_6t
Xbit_r71_c70 bl[70] br[70] wl[71] vdd gnd cell_6t
Xbit_r72_c70 bl[70] br[70] wl[72] vdd gnd cell_6t
Xbit_r73_c70 bl[70] br[70] wl[73] vdd gnd cell_6t
Xbit_r74_c70 bl[70] br[70] wl[74] vdd gnd cell_6t
Xbit_r75_c70 bl[70] br[70] wl[75] vdd gnd cell_6t
Xbit_r76_c70 bl[70] br[70] wl[76] vdd gnd cell_6t
Xbit_r77_c70 bl[70] br[70] wl[77] vdd gnd cell_6t
Xbit_r78_c70 bl[70] br[70] wl[78] vdd gnd cell_6t
Xbit_r79_c70 bl[70] br[70] wl[79] vdd gnd cell_6t
Xbit_r80_c70 bl[70] br[70] wl[80] vdd gnd cell_6t
Xbit_r81_c70 bl[70] br[70] wl[81] vdd gnd cell_6t
Xbit_r82_c70 bl[70] br[70] wl[82] vdd gnd cell_6t
Xbit_r83_c70 bl[70] br[70] wl[83] vdd gnd cell_6t
Xbit_r84_c70 bl[70] br[70] wl[84] vdd gnd cell_6t
Xbit_r85_c70 bl[70] br[70] wl[85] vdd gnd cell_6t
Xbit_r86_c70 bl[70] br[70] wl[86] vdd gnd cell_6t
Xbit_r87_c70 bl[70] br[70] wl[87] vdd gnd cell_6t
Xbit_r88_c70 bl[70] br[70] wl[88] vdd gnd cell_6t
Xbit_r89_c70 bl[70] br[70] wl[89] vdd gnd cell_6t
Xbit_r90_c70 bl[70] br[70] wl[90] vdd gnd cell_6t
Xbit_r91_c70 bl[70] br[70] wl[91] vdd gnd cell_6t
Xbit_r92_c70 bl[70] br[70] wl[92] vdd gnd cell_6t
Xbit_r93_c70 bl[70] br[70] wl[93] vdd gnd cell_6t
Xbit_r94_c70 bl[70] br[70] wl[94] vdd gnd cell_6t
Xbit_r95_c70 bl[70] br[70] wl[95] vdd gnd cell_6t
Xbit_r96_c70 bl[70] br[70] wl[96] vdd gnd cell_6t
Xbit_r97_c70 bl[70] br[70] wl[97] vdd gnd cell_6t
Xbit_r98_c70 bl[70] br[70] wl[98] vdd gnd cell_6t
Xbit_r99_c70 bl[70] br[70] wl[99] vdd gnd cell_6t
Xbit_r100_c70 bl[70] br[70] wl[100] vdd gnd cell_6t
Xbit_r101_c70 bl[70] br[70] wl[101] vdd gnd cell_6t
Xbit_r102_c70 bl[70] br[70] wl[102] vdd gnd cell_6t
Xbit_r103_c70 bl[70] br[70] wl[103] vdd gnd cell_6t
Xbit_r104_c70 bl[70] br[70] wl[104] vdd gnd cell_6t
Xbit_r105_c70 bl[70] br[70] wl[105] vdd gnd cell_6t
Xbit_r106_c70 bl[70] br[70] wl[106] vdd gnd cell_6t
Xbit_r107_c70 bl[70] br[70] wl[107] vdd gnd cell_6t
Xbit_r108_c70 bl[70] br[70] wl[108] vdd gnd cell_6t
Xbit_r109_c70 bl[70] br[70] wl[109] vdd gnd cell_6t
Xbit_r110_c70 bl[70] br[70] wl[110] vdd gnd cell_6t
Xbit_r111_c70 bl[70] br[70] wl[111] vdd gnd cell_6t
Xbit_r112_c70 bl[70] br[70] wl[112] vdd gnd cell_6t
Xbit_r113_c70 bl[70] br[70] wl[113] vdd gnd cell_6t
Xbit_r114_c70 bl[70] br[70] wl[114] vdd gnd cell_6t
Xbit_r115_c70 bl[70] br[70] wl[115] vdd gnd cell_6t
Xbit_r116_c70 bl[70] br[70] wl[116] vdd gnd cell_6t
Xbit_r117_c70 bl[70] br[70] wl[117] vdd gnd cell_6t
Xbit_r118_c70 bl[70] br[70] wl[118] vdd gnd cell_6t
Xbit_r119_c70 bl[70] br[70] wl[119] vdd gnd cell_6t
Xbit_r120_c70 bl[70] br[70] wl[120] vdd gnd cell_6t
Xbit_r121_c70 bl[70] br[70] wl[121] vdd gnd cell_6t
Xbit_r122_c70 bl[70] br[70] wl[122] vdd gnd cell_6t
Xbit_r123_c70 bl[70] br[70] wl[123] vdd gnd cell_6t
Xbit_r124_c70 bl[70] br[70] wl[124] vdd gnd cell_6t
Xbit_r125_c70 bl[70] br[70] wl[125] vdd gnd cell_6t
Xbit_r126_c70 bl[70] br[70] wl[126] vdd gnd cell_6t
Xbit_r127_c70 bl[70] br[70] wl[127] vdd gnd cell_6t
Xbit_r128_c70 bl[70] br[70] wl[128] vdd gnd cell_6t
Xbit_r129_c70 bl[70] br[70] wl[129] vdd gnd cell_6t
Xbit_r130_c70 bl[70] br[70] wl[130] vdd gnd cell_6t
Xbit_r131_c70 bl[70] br[70] wl[131] vdd gnd cell_6t
Xbit_r132_c70 bl[70] br[70] wl[132] vdd gnd cell_6t
Xbit_r133_c70 bl[70] br[70] wl[133] vdd gnd cell_6t
Xbit_r134_c70 bl[70] br[70] wl[134] vdd gnd cell_6t
Xbit_r135_c70 bl[70] br[70] wl[135] vdd gnd cell_6t
Xbit_r136_c70 bl[70] br[70] wl[136] vdd gnd cell_6t
Xbit_r137_c70 bl[70] br[70] wl[137] vdd gnd cell_6t
Xbit_r138_c70 bl[70] br[70] wl[138] vdd gnd cell_6t
Xbit_r139_c70 bl[70] br[70] wl[139] vdd gnd cell_6t
Xbit_r140_c70 bl[70] br[70] wl[140] vdd gnd cell_6t
Xbit_r141_c70 bl[70] br[70] wl[141] vdd gnd cell_6t
Xbit_r142_c70 bl[70] br[70] wl[142] vdd gnd cell_6t
Xbit_r143_c70 bl[70] br[70] wl[143] vdd gnd cell_6t
Xbit_r144_c70 bl[70] br[70] wl[144] vdd gnd cell_6t
Xbit_r145_c70 bl[70] br[70] wl[145] vdd gnd cell_6t
Xbit_r146_c70 bl[70] br[70] wl[146] vdd gnd cell_6t
Xbit_r147_c70 bl[70] br[70] wl[147] vdd gnd cell_6t
Xbit_r148_c70 bl[70] br[70] wl[148] vdd gnd cell_6t
Xbit_r149_c70 bl[70] br[70] wl[149] vdd gnd cell_6t
Xbit_r150_c70 bl[70] br[70] wl[150] vdd gnd cell_6t
Xbit_r151_c70 bl[70] br[70] wl[151] vdd gnd cell_6t
Xbit_r152_c70 bl[70] br[70] wl[152] vdd gnd cell_6t
Xbit_r153_c70 bl[70] br[70] wl[153] vdd gnd cell_6t
Xbit_r154_c70 bl[70] br[70] wl[154] vdd gnd cell_6t
Xbit_r155_c70 bl[70] br[70] wl[155] vdd gnd cell_6t
Xbit_r156_c70 bl[70] br[70] wl[156] vdd gnd cell_6t
Xbit_r157_c70 bl[70] br[70] wl[157] vdd gnd cell_6t
Xbit_r158_c70 bl[70] br[70] wl[158] vdd gnd cell_6t
Xbit_r159_c70 bl[70] br[70] wl[159] vdd gnd cell_6t
Xbit_r160_c70 bl[70] br[70] wl[160] vdd gnd cell_6t
Xbit_r161_c70 bl[70] br[70] wl[161] vdd gnd cell_6t
Xbit_r162_c70 bl[70] br[70] wl[162] vdd gnd cell_6t
Xbit_r163_c70 bl[70] br[70] wl[163] vdd gnd cell_6t
Xbit_r164_c70 bl[70] br[70] wl[164] vdd gnd cell_6t
Xbit_r165_c70 bl[70] br[70] wl[165] vdd gnd cell_6t
Xbit_r166_c70 bl[70] br[70] wl[166] vdd gnd cell_6t
Xbit_r167_c70 bl[70] br[70] wl[167] vdd gnd cell_6t
Xbit_r168_c70 bl[70] br[70] wl[168] vdd gnd cell_6t
Xbit_r169_c70 bl[70] br[70] wl[169] vdd gnd cell_6t
Xbit_r170_c70 bl[70] br[70] wl[170] vdd gnd cell_6t
Xbit_r171_c70 bl[70] br[70] wl[171] vdd gnd cell_6t
Xbit_r172_c70 bl[70] br[70] wl[172] vdd gnd cell_6t
Xbit_r173_c70 bl[70] br[70] wl[173] vdd gnd cell_6t
Xbit_r174_c70 bl[70] br[70] wl[174] vdd gnd cell_6t
Xbit_r175_c70 bl[70] br[70] wl[175] vdd gnd cell_6t
Xbit_r176_c70 bl[70] br[70] wl[176] vdd gnd cell_6t
Xbit_r177_c70 bl[70] br[70] wl[177] vdd gnd cell_6t
Xbit_r178_c70 bl[70] br[70] wl[178] vdd gnd cell_6t
Xbit_r179_c70 bl[70] br[70] wl[179] vdd gnd cell_6t
Xbit_r180_c70 bl[70] br[70] wl[180] vdd gnd cell_6t
Xbit_r181_c70 bl[70] br[70] wl[181] vdd gnd cell_6t
Xbit_r182_c70 bl[70] br[70] wl[182] vdd gnd cell_6t
Xbit_r183_c70 bl[70] br[70] wl[183] vdd gnd cell_6t
Xbit_r184_c70 bl[70] br[70] wl[184] vdd gnd cell_6t
Xbit_r185_c70 bl[70] br[70] wl[185] vdd gnd cell_6t
Xbit_r186_c70 bl[70] br[70] wl[186] vdd gnd cell_6t
Xbit_r187_c70 bl[70] br[70] wl[187] vdd gnd cell_6t
Xbit_r188_c70 bl[70] br[70] wl[188] vdd gnd cell_6t
Xbit_r189_c70 bl[70] br[70] wl[189] vdd gnd cell_6t
Xbit_r190_c70 bl[70] br[70] wl[190] vdd gnd cell_6t
Xbit_r191_c70 bl[70] br[70] wl[191] vdd gnd cell_6t
Xbit_r192_c70 bl[70] br[70] wl[192] vdd gnd cell_6t
Xbit_r193_c70 bl[70] br[70] wl[193] vdd gnd cell_6t
Xbit_r194_c70 bl[70] br[70] wl[194] vdd gnd cell_6t
Xbit_r195_c70 bl[70] br[70] wl[195] vdd gnd cell_6t
Xbit_r196_c70 bl[70] br[70] wl[196] vdd gnd cell_6t
Xbit_r197_c70 bl[70] br[70] wl[197] vdd gnd cell_6t
Xbit_r198_c70 bl[70] br[70] wl[198] vdd gnd cell_6t
Xbit_r199_c70 bl[70] br[70] wl[199] vdd gnd cell_6t
Xbit_r200_c70 bl[70] br[70] wl[200] vdd gnd cell_6t
Xbit_r201_c70 bl[70] br[70] wl[201] vdd gnd cell_6t
Xbit_r202_c70 bl[70] br[70] wl[202] vdd gnd cell_6t
Xbit_r203_c70 bl[70] br[70] wl[203] vdd gnd cell_6t
Xbit_r204_c70 bl[70] br[70] wl[204] vdd gnd cell_6t
Xbit_r205_c70 bl[70] br[70] wl[205] vdd gnd cell_6t
Xbit_r206_c70 bl[70] br[70] wl[206] vdd gnd cell_6t
Xbit_r207_c70 bl[70] br[70] wl[207] vdd gnd cell_6t
Xbit_r208_c70 bl[70] br[70] wl[208] vdd gnd cell_6t
Xbit_r209_c70 bl[70] br[70] wl[209] vdd gnd cell_6t
Xbit_r210_c70 bl[70] br[70] wl[210] vdd gnd cell_6t
Xbit_r211_c70 bl[70] br[70] wl[211] vdd gnd cell_6t
Xbit_r212_c70 bl[70] br[70] wl[212] vdd gnd cell_6t
Xbit_r213_c70 bl[70] br[70] wl[213] vdd gnd cell_6t
Xbit_r214_c70 bl[70] br[70] wl[214] vdd gnd cell_6t
Xbit_r215_c70 bl[70] br[70] wl[215] vdd gnd cell_6t
Xbit_r216_c70 bl[70] br[70] wl[216] vdd gnd cell_6t
Xbit_r217_c70 bl[70] br[70] wl[217] vdd gnd cell_6t
Xbit_r218_c70 bl[70] br[70] wl[218] vdd gnd cell_6t
Xbit_r219_c70 bl[70] br[70] wl[219] vdd gnd cell_6t
Xbit_r220_c70 bl[70] br[70] wl[220] vdd gnd cell_6t
Xbit_r221_c70 bl[70] br[70] wl[221] vdd gnd cell_6t
Xbit_r222_c70 bl[70] br[70] wl[222] vdd gnd cell_6t
Xbit_r223_c70 bl[70] br[70] wl[223] vdd gnd cell_6t
Xbit_r224_c70 bl[70] br[70] wl[224] vdd gnd cell_6t
Xbit_r225_c70 bl[70] br[70] wl[225] vdd gnd cell_6t
Xbit_r226_c70 bl[70] br[70] wl[226] vdd gnd cell_6t
Xbit_r227_c70 bl[70] br[70] wl[227] vdd gnd cell_6t
Xbit_r228_c70 bl[70] br[70] wl[228] vdd gnd cell_6t
Xbit_r229_c70 bl[70] br[70] wl[229] vdd gnd cell_6t
Xbit_r230_c70 bl[70] br[70] wl[230] vdd gnd cell_6t
Xbit_r231_c70 bl[70] br[70] wl[231] vdd gnd cell_6t
Xbit_r232_c70 bl[70] br[70] wl[232] vdd gnd cell_6t
Xbit_r233_c70 bl[70] br[70] wl[233] vdd gnd cell_6t
Xbit_r234_c70 bl[70] br[70] wl[234] vdd gnd cell_6t
Xbit_r235_c70 bl[70] br[70] wl[235] vdd gnd cell_6t
Xbit_r236_c70 bl[70] br[70] wl[236] vdd gnd cell_6t
Xbit_r237_c70 bl[70] br[70] wl[237] vdd gnd cell_6t
Xbit_r238_c70 bl[70] br[70] wl[238] vdd gnd cell_6t
Xbit_r239_c70 bl[70] br[70] wl[239] vdd gnd cell_6t
Xbit_r240_c70 bl[70] br[70] wl[240] vdd gnd cell_6t
Xbit_r241_c70 bl[70] br[70] wl[241] vdd gnd cell_6t
Xbit_r242_c70 bl[70] br[70] wl[242] vdd gnd cell_6t
Xbit_r243_c70 bl[70] br[70] wl[243] vdd gnd cell_6t
Xbit_r244_c70 bl[70] br[70] wl[244] vdd gnd cell_6t
Xbit_r245_c70 bl[70] br[70] wl[245] vdd gnd cell_6t
Xbit_r246_c70 bl[70] br[70] wl[246] vdd gnd cell_6t
Xbit_r247_c70 bl[70] br[70] wl[247] vdd gnd cell_6t
Xbit_r248_c70 bl[70] br[70] wl[248] vdd gnd cell_6t
Xbit_r249_c70 bl[70] br[70] wl[249] vdd gnd cell_6t
Xbit_r250_c70 bl[70] br[70] wl[250] vdd gnd cell_6t
Xbit_r251_c70 bl[70] br[70] wl[251] vdd gnd cell_6t
Xbit_r252_c70 bl[70] br[70] wl[252] vdd gnd cell_6t
Xbit_r253_c70 bl[70] br[70] wl[253] vdd gnd cell_6t
Xbit_r254_c70 bl[70] br[70] wl[254] vdd gnd cell_6t
Xbit_r255_c70 bl[70] br[70] wl[255] vdd gnd cell_6t
Xbit_r256_c70 bl[70] br[70] wl[256] vdd gnd cell_6t
Xbit_r257_c70 bl[70] br[70] wl[257] vdd gnd cell_6t
Xbit_r258_c70 bl[70] br[70] wl[258] vdd gnd cell_6t
Xbit_r259_c70 bl[70] br[70] wl[259] vdd gnd cell_6t
Xbit_r260_c70 bl[70] br[70] wl[260] vdd gnd cell_6t
Xbit_r261_c70 bl[70] br[70] wl[261] vdd gnd cell_6t
Xbit_r262_c70 bl[70] br[70] wl[262] vdd gnd cell_6t
Xbit_r263_c70 bl[70] br[70] wl[263] vdd gnd cell_6t
Xbit_r264_c70 bl[70] br[70] wl[264] vdd gnd cell_6t
Xbit_r265_c70 bl[70] br[70] wl[265] vdd gnd cell_6t
Xbit_r266_c70 bl[70] br[70] wl[266] vdd gnd cell_6t
Xbit_r267_c70 bl[70] br[70] wl[267] vdd gnd cell_6t
Xbit_r268_c70 bl[70] br[70] wl[268] vdd gnd cell_6t
Xbit_r269_c70 bl[70] br[70] wl[269] vdd gnd cell_6t
Xbit_r270_c70 bl[70] br[70] wl[270] vdd gnd cell_6t
Xbit_r271_c70 bl[70] br[70] wl[271] vdd gnd cell_6t
Xbit_r272_c70 bl[70] br[70] wl[272] vdd gnd cell_6t
Xbit_r273_c70 bl[70] br[70] wl[273] vdd gnd cell_6t
Xbit_r274_c70 bl[70] br[70] wl[274] vdd gnd cell_6t
Xbit_r275_c70 bl[70] br[70] wl[275] vdd gnd cell_6t
Xbit_r276_c70 bl[70] br[70] wl[276] vdd gnd cell_6t
Xbit_r277_c70 bl[70] br[70] wl[277] vdd gnd cell_6t
Xbit_r278_c70 bl[70] br[70] wl[278] vdd gnd cell_6t
Xbit_r279_c70 bl[70] br[70] wl[279] vdd gnd cell_6t
Xbit_r280_c70 bl[70] br[70] wl[280] vdd gnd cell_6t
Xbit_r281_c70 bl[70] br[70] wl[281] vdd gnd cell_6t
Xbit_r282_c70 bl[70] br[70] wl[282] vdd gnd cell_6t
Xbit_r283_c70 bl[70] br[70] wl[283] vdd gnd cell_6t
Xbit_r284_c70 bl[70] br[70] wl[284] vdd gnd cell_6t
Xbit_r285_c70 bl[70] br[70] wl[285] vdd gnd cell_6t
Xbit_r286_c70 bl[70] br[70] wl[286] vdd gnd cell_6t
Xbit_r287_c70 bl[70] br[70] wl[287] vdd gnd cell_6t
Xbit_r288_c70 bl[70] br[70] wl[288] vdd gnd cell_6t
Xbit_r289_c70 bl[70] br[70] wl[289] vdd gnd cell_6t
Xbit_r290_c70 bl[70] br[70] wl[290] vdd gnd cell_6t
Xbit_r291_c70 bl[70] br[70] wl[291] vdd gnd cell_6t
Xbit_r292_c70 bl[70] br[70] wl[292] vdd gnd cell_6t
Xbit_r293_c70 bl[70] br[70] wl[293] vdd gnd cell_6t
Xbit_r294_c70 bl[70] br[70] wl[294] vdd gnd cell_6t
Xbit_r295_c70 bl[70] br[70] wl[295] vdd gnd cell_6t
Xbit_r296_c70 bl[70] br[70] wl[296] vdd gnd cell_6t
Xbit_r297_c70 bl[70] br[70] wl[297] vdd gnd cell_6t
Xbit_r298_c70 bl[70] br[70] wl[298] vdd gnd cell_6t
Xbit_r299_c70 bl[70] br[70] wl[299] vdd gnd cell_6t
Xbit_r300_c70 bl[70] br[70] wl[300] vdd gnd cell_6t
Xbit_r301_c70 bl[70] br[70] wl[301] vdd gnd cell_6t
Xbit_r302_c70 bl[70] br[70] wl[302] vdd gnd cell_6t
Xbit_r303_c70 bl[70] br[70] wl[303] vdd gnd cell_6t
Xbit_r304_c70 bl[70] br[70] wl[304] vdd gnd cell_6t
Xbit_r305_c70 bl[70] br[70] wl[305] vdd gnd cell_6t
Xbit_r306_c70 bl[70] br[70] wl[306] vdd gnd cell_6t
Xbit_r307_c70 bl[70] br[70] wl[307] vdd gnd cell_6t
Xbit_r308_c70 bl[70] br[70] wl[308] vdd gnd cell_6t
Xbit_r309_c70 bl[70] br[70] wl[309] vdd gnd cell_6t
Xbit_r310_c70 bl[70] br[70] wl[310] vdd gnd cell_6t
Xbit_r311_c70 bl[70] br[70] wl[311] vdd gnd cell_6t
Xbit_r312_c70 bl[70] br[70] wl[312] vdd gnd cell_6t
Xbit_r313_c70 bl[70] br[70] wl[313] vdd gnd cell_6t
Xbit_r314_c70 bl[70] br[70] wl[314] vdd gnd cell_6t
Xbit_r315_c70 bl[70] br[70] wl[315] vdd gnd cell_6t
Xbit_r316_c70 bl[70] br[70] wl[316] vdd gnd cell_6t
Xbit_r317_c70 bl[70] br[70] wl[317] vdd gnd cell_6t
Xbit_r318_c70 bl[70] br[70] wl[318] vdd gnd cell_6t
Xbit_r319_c70 bl[70] br[70] wl[319] vdd gnd cell_6t
Xbit_r320_c70 bl[70] br[70] wl[320] vdd gnd cell_6t
Xbit_r321_c70 bl[70] br[70] wl[321] vdd gnd cell_6t
Xbit_r322_c70 bl[70] br[70] wl[322] vdd gnd cell_6t
Xbit_r323_c70 bl[70] br[70] wl[323] vdd gnd cell_6t
Xbit_r324_c70 bl[70] br[70] wl[324] vdd gnd cell_6t
Xbit_r325_c70 bl[70] br[70] wl[325] vdd gnd cell_6t
Xbit_r326_c70 bl[70] br[70] wl[326] vdd gnd cell_6t
Xbit_r327_c70 bl[70] br[70] wl[327] vdd gnd cell_6t
Xbit_r328_c70 bl[70] br[70] wl[328] vdd gnd cell_6t
Xbit_r329_c70 bl[70] br[70] wl[329] vdd gnd cell_6t
Xbit_r330_c70 bl[70] br[70] wl[330] vdd gnd cell_6t
Xbit_r331_c70 bl[70] br[70] wl[331] vdd gnd cell_6t
Xbit_r332_c70 bl[70] br[70] wl[332] vdd gnd cell_6t
Xbit_r333_c70 bl[70] br[70] wl[333] vdd gnd cell_6t
Xbit_r334_c70 bl[70] br[70] wl[334] vdd gnd cell_6t
Xbit_r335_c70 bl[70] br[70] wl[335] vdd gnd cell_6t
Xbit_r336_c70 bl[70] br[70] wl[336] vdd gnd cell_6t
Xbit_r337_c70 bl[70] br[70] wl[337] vdd gnd cell_6t
Xbit_r338_c70 bl[70] br[70] wl[338] vdd gnd cell_6t
Xbit_r339_c70 bl[70] br[70] wl[339] vdd gnd cell_6t
Xbit_r340_c70 bl[70] br[70] wl[340] vdd gnd cell_6t
Xbit_r341_c70 bl[70] br[70] wl[341] vdd gnd cell_6t
Xbit_r342_c70 bl[70] br[70] wl[342] vdd gnd cell_6t
Xbit_r343_c70 bl[70] br[70] wl[343] vdd gnd cell_6t
Xbit_r344_c70 bl[70] br[70] wl[344] vdd gnd cell_6t
Xbit_r345_c70 bl[70] br[70] wl[345] vdd gnd cell_6t
Xbit_r346_c70 bl[70] br[70] wl[346] vdd gnd cell_6t
Xbit_r347_c70 bl[70] br[70] wl[347] vdd gnd cell_6t
Xbit_r348_c70 bl[70] br[70] wl[348] vdd gnd cell_6t
Xbit_r349_c70 bl[70] br[70] wl[349] vdd gnd cell_6t
Xbit_r350_c70 bl[70] br[70] wl[350] vdd gnd cell_6t
Xbit_r351_c70 bl[70] br[70] wl[351] vdd gnd cell_6t
Xbit_r352_c70 bl[70] br[70] wl[352] vdd gnd cell_6t
Xbit_r353_c70 bl[70] br[70] wl[353] vdd gnd cell_6t
Xbit_r354_c70 bl[70] br[70] wl[354] vdd gnd cell_6t
Xbit_r355_c70 bl[70] br[70] wl[355] vdd gnd cell_6t
Xbit_r356_c70 bl[70] br[70] wl[356] vdd gnd cell_6t
Xbit_r357_c70 bl[70] br[70] wl[357] vdd gnd cell_6t
Xbit_r358_c70 bl[70] br[70] wl[358] vdd gnd cell_6t
Xbit_r359_c70 bl[70] br[70] wl[359] vdd gnd cell_6t
Xbit_r360_c70 bl[70] br[70] wl[360] vdd gnd cell_6t
Xbit_r361_c70 bl[70] br[70] wl[361] vdd gnd cell_6t
Xbit_r362_c70 bl[70] br[70] wl[362] vdd gnd cell_6t
Xbit_r363_c70 bl[70] br[70] wl[363] vdd gnd cell_6t
Xbit_r364_c70 bl[70] br[70] wl[364] vdd gnd cell_6t
Xbit_r365_c70 bl[70] br[70] wl[365] vdd gnd cell_6t
Xbit_r366_c70 bl[70] br[70] wl[366] vdd gnd cell_6t
Xbit_r367_c70 bl[70] br[70] wl[367] vdd gnd cell_6t
Xbit_r368_c70 bl[70] br[70] wl[368] vdd gnd cell_6t
Xbit_r369_c70 bl[70] br[70] wl[369] vdd gnd cell_6t
Xbit_r370_c70 bl[70] br[70] wl[370] vdd gnd cell_6t
Xbit_r371_c70 bl[70] br[70] wl[371] vdd gnd cell_6t
Xbit_r372_c70 bl[70] br[70] wl[372] vdd gnd cell_6t
Xbit_r373_c70 bl[70] br[70] wl[373] vdd gnd cell_6t
Xbit_r374_c70 bl[70] br[70] wl[374] vdd gnd cell_6t
Xbit_r375_c70 bl[70] br[70] wl[375] vdd gnd cell_6t
Xbit_r376_c70 bl[70] br[70] wl[376] vdd gnd cell_6t
Xbit_r377_c70 bl[70] br[70] wl[377] vdd gnd cell_6t
Xbit_r378_c70 bl[70] br[70] wl[378] vdd gnd cell_6t
Xbit_r379_c70 bl[70] br[70] wl[379] vdd gnd cell_6t
Xbit_r380_c70 bl[70] br[70] wl[380] vdd gnd cell_6t
Xbit_r381_c70 bl[70] br[70] wl[381] vdd gnd cell_6t
Xbit_r382_c70 bl[70] br[70] wl[382] vdd gnd cell_6t
Xbit_r383_c70 bl[70] br[70] wl[383] vdd gnd cell_6t
Xbit_r384_c70 bl[70] br[70] wl[384] vdd gnd cell_6t
Xbit_r385_c70 bl[70] br[70] wl[385] vdd gnd cell_6t
Xbit_r386_c70 bl[70] br[70] wl[386] vdd gnd cell_6t
Xbit_r387_c70 bl[70] br[70] wl[387] vdd gnd cell_6t
Xbit_r388_c70 bl[70] br[70] wl[388] vdd gnd cell_6t
Xbit_r389_c70 bl[70] br[70] wl[389] vdd gnd cell_6t
Xbit_r390_c70 bl[70] br[70] wl[390] vdd gnd cell_6t
Xbit_r391_c70 bl[70] br[70] wl[391] vdd gnd cell_6t
Xbit_r392_c70 bl[70] br[70] wl[392] vdd gnd cell_6t
Xbit_r393_c70 bl[70] br[70] wl[393] vdd gnd cell_6t
Xbit_r394_c70 bl[70] br[70] wl[394] vdd gnd cell_6t
Xbit_r395_c70 bl[70] br[70] wl[395] vdd gnd cell_6t
Xbit_r396_c70 bl[70] br[70] wl[396] vdd gnd cell_6t
Xbit_r397_c70 bl[70] br[70] wl[397] vdd gnd cell_6t
Xbit_r398_c70 bl[70] br[70] wl[398] vdd gnd cell_6t
Xbit_r399_c70 bl[70] br[70] wl[399] vdd gnd cell_6t
Xbit_r400_c70 bl[70] br[70] wl[400] vdd gnd cell_6t
Xbit_r401_c70 bl[70] br[70] wl[401] vdd gnd cell_6t
Xbit_r402_c70 bl[70] br[70] wl[402] vdd gnd cell_6t
Xbit_r403_c70 bl[70] br[70] wl[403] vdd gnd cell_6t
Xbit_r404_c70 bl[70] br[70] wl[404] vdd gnd cell_6t
Xbit_r405_c70 bl[70] br[70] wl[405] vdd gnd cell_6t
Xbit_r406_c70 bl[70] br[70] wl[406] vdd gnd cell_6t
Xbit_r407_c70 bl[70] br[70] wl[407] vdd gnd cell_6t
Xbit_r408_c70 bl[70] br[70] wl[408] vdd gnd cell_6t
Xbit_r409_c70 bl[70] br[70] wl[409] vdd gnd cell_6t
Xbit_r410_c70 bl[70] br[70] wl[410] vdd gnd cell_6t
Xbit_r411_c70 bl[70] br[70] wl[411] vdd gnd cell_6t
Xbit_r412_c70 bl[70] br[70] wl[412] vdd gnd cell_6t
Xbit_r413_c70 bl[70] br[70] wl[413] vdd gnd cell_6t
Xbit_r414_c70 bl[70] br[70] wl[414] vdd gnd cell_6t
Xbit_r415_c70 bl[70] br[70] wl[415] vdd gnd cell_6t
Xbit_r416_c70 bl[70] br[70] wl[416] vdd gnd cell_6t
Xbit_r417_c70 bl[70] br[70] wl[417] vdd gnd cell_6t
Xbit_r418_c70 bl[70] br[70] wl[418] vdd gnd cell_6t
Xbit_r419_c70 bl[70] br[70] wl[419] vdd gnd cell_6t
Xbit_r420_c70 bl[70] br[70] wl[420] vdd gnd cell_6t
Xbit_r421_c70 bl[70] br[70] wl[421] vdd gnd cell_6t
Xbit_r422_c70 bl[70] br[70] wl[422] vdd gnd cell_6t
Xbit_r423_c70 bl[70] br[70] wl[423] vdd gnd cell_6t
Xbit_r424_c70 bl[70] br[70] wl[424] vdd gnd cell_6t
Xbit_r425_c70 bl[70] br[70] wl[425] vdd gnd cell_6t
Xbit_r426_c70 bl[70] br[70] wl[426] vdd gnd cell_6t
Xbit_r427_c70 bl[70] br[70] wl[427] vdd gnd cell_6t
Xbit_r428_c70 bl[70] br[70] wl[428] vdd gnd cell_6t
Xbit_r429_c70 bl[70] br[70] wl[429] vdd gnd cell_6t
Xbit_r430_c70 bl[70] br[70] wl[430] vdd gnd cell_6t
Xbit_r431_c70 bl[70] br[70] wl[431] vdd gnd cell_6t
Xbit_r432_c70 bl[70] br[70] wl[432] vdd gnd cell_6t
Xbit_r433_c70 bl[70] br[70] wl[433] vdd gnd cell_6t
Xbit_r434_c70 bl[70] br[70] wl[434] vdd gnd cell_6t
Xbit_r435_c70 bl[70] br[70] wl[435] vdd gnd cell_6t
Xbit_r436_c70 bl[70] br[70] wl[436] vdd gnd cell_6t
Xbit_r437_c70 bl[70] br[70] wl[437] vdd gnd cell_6t
Xbit_r438_c70 bl[70] br[70] wl[438] vdd gnd cell_6t
Xbit_r439_c70 bl[70] br[70] wl[439] vdd gnd cell_6t
Xbit_r440_c70 bl[70] br[70] wl[440] vdd gnd cell_6t
Xbit_r441_c70 bl[70] br[70] wl[441] vdd gnd cell_6t
Xbit_r442_c70 bl[70] br[70] wl[442] vdd gnd cell_6t
Xbit_r443_c70 bl[70] br[70] wl[443] vdd gnd cell_6t
Xbit_r444_c70 bl[70] br[70] wl[444] vdd gnd cell_6t
Xbit_r445_c70 bl[70] br[70] wl[445] vdd gnd cell_6t
Xbit_r446_c70 bl[70] br[70] wl[446] vdd gnd cell_6t
Xbit_r447_c70 bl[70] br[70] wl[447] vdd gnd cell_6t
Xbit_r448_c70 bl[70] br[70] wl[448] vdd gnd cell_6t
Xbit_r449_c70 bl[70] br[70] wl[449] vdd gnd cell_6t
Xbit_r450_c70 bl[70] br[70] wl[450] vdd gnd cell_6t
Xbit_r451_c70 bl[70] br[70] wl[451] vdd gnd cell_6t
Xbit_r452_c70 bl[70] br[70] wl[452] vdd gnd cell_6t
Xbit_r453_c70 bl[70] br[70] wl[453] vdd gnd cell_6t
Xbit_r454_c70 bl[70] br[70] wl[454] vdd gnd cell_6t
Xbit_r455_c70 bl[70] br[70] wl[455] vdd gnd cell_6t
Xbit_r456_c70 bl[70] br[70] wl[456] vdd gnd cell_6t
Xbit_r457_c70 bl[70] br[70] wl[457] vdd gnd cell_6t
Xbit_r458_c70 bl[70] br[70] wl[458] vdd gnd cell_6t
Xbit_r459_c70 bl[70] br[70] wl[459] vdd gnd cell_6t
Xbit_r460_c70 bl[70] br[70] wl[460] vdd gnd cell_6t
Xbit_r461_c70 bl[70] br[70] wl[461] vdd gnd cell_6t
Xbit_r462_c70 bl[70] br[70] wl[462] vdd gnd cell_6t
Xbit_r463_c70 bl[70] br[70] wl[463] vdd gnd cell_6t
Xbit_r464_c70 bl[70] br[70] wl[464] vdd gnd cell_6t
Xbit_r465_c70 bl[70] br[70] wl[465] vdd gnd cell_6t
Xbit_r466_c70 bl[70] br[70] wl[466] vdd gnd cell_6t
Xbit_r467_c70 bl[70] br[70] wl[467] vdd gnd cell_6t
Xbit_r468_c70 bl[70] br[70] wl[468] vdd gnd cell_6t
Xbit_r469_c70 bl[70] br[70] wl[469] vdd gnd cell_6t
Xbit_r470_c70 bl[70] br[70] wl[470] vdd gnd cell_6t
Xbit_r471_c70 bl[70] br[70] wl[471] vdd gnd cell_6t
Xbit_r472_c70 bl[70] br[70] wl[472] vdd gnd cell_6t
Xbit_r473_c70 bl[70] br[70] wl[473] vdd gnd cell_6t
Xbit_r474_c70 bl[70] br[70] wl[474] vdd gnd cell_6t
Xbit_r475_c70 bl[70] br[70] wl[475] vdd gnd cell_6t
Xbit_r476_c70 bl[70] br[70] wl[476] vdd gnd cell_6t
Xbit_r477_c70 bl[70] br[70] wl[477] vdd gnd cell_6t
Xbit_r478_c70 bl[70] br[70] wl[478] vdd gnd cell_6t
Xbit_r479_c70 bl[70] br[70] wl[479] vdd gnd cell_6t
Xbit_r480_c70 bl[70] br[70] wl[480] vdd gnd cell_6t
Xbit_r481_c70 bl[70] br[70] wl[481] vdd gnd cell_6t
Xbit_r482_c70 bl[70] br[70] wl[482] vdd gnd cell_6t
Xbit_r483_c70 bl[70] br[70] wl[483] vdd gnd cell_6t
Xbit_r484_c70 bl[70] br[70] wl[484] vdd gnd cell_6t
Xbit_r485_c70 bl[70] br[70] wl[485] vdd gnd cell_6t
Xbit_r486_c70 bl[70] br[70] wl[486] vdd gnd cell_6t
Xbit_r487_c70 bl[70] br[70] wl[487] vdd gnd cell_6t
Xbit_r488_c70 bl[70] br[70] wl[488] vdd gnd cell_6t
Xbit_r489_c70 bl[70] br[70] wl[489] vdd gnd cell_6t
Xbit_r490_c70 bl[70] br[70] wl[490] vdd gnd cell_6t
Xbit_r491_c70 bl[70] br[70] wl[491] vdd gnd cell_6t
Xbit_r492_c70 bl[70] br[70] wl[492] vdd gnd cell_6t
Xbit_r493_c70 bl[70] br[70] wl[493] vdd gnd cell_6t
Xbit_r494_c70 bl[70] br[70] wl[494] vdd gnd cell_6t
Xbit_r495_c70 bl[70] br[70] wl[495] vdd gnd cell_6t
Xbit_r496_c70 bl[70] br[70] wl[496] vdd gnd cell_6t
Xbit_r497_c70 bl[70] br[70] wl[497] vdd gnd cell_6t
Xbit_r498_c70 bl[70] br[70] wl[498] vdd gnd cell_6t
Xbit_r499_c70 bl[70] br[70] wl[499] vdd gnd cell_6t
Xbit_r500_c70 bl[70] br[70] wl[500] vdd gnd cell_6t
Xbit_r501_c70 bl[70] br[70] wl[501] vdd gnd cell_6t
Xbit_r502_c70 bl[70] br[70] wl[502] vdd gnd cell_6t
Xbit_r503_c70 bl[70] br[70] wl[503] vdd gnd cell_6t
Xbit_r504_c70 bl[70] br[70] wl[504] vdd gnd cell_6t
Xbit_r505_c70 bl[70] br[70] wl[505] vdd gnd cell_6t
Xbit_r506_c70 bl[70] br[70] wl[506] vdd gnd cell_6t
Xbit_r507_c70 bl[70] br[70] wl[507] vdd gnd cell_6t
Xbit_r508_c70 bl[70] br[70] wl[508] vdd gnd cell_6t
Xbit_r509_c70 bl[70] br[70] wl[509] vdd gnd cell_6t
Xbit_r510_c70 bl[70] br[70] wl[510] vdd gnd cell_6t
Xbit_r511_c70 bl[70] br[70] wl[511] vdd gnd cell_6t
Xbit_r0_c71 bl[71] br[71] wl[0] vdd gnd cell_6t
Xbit_r1_c71 bl[71] br[71] wl[1] vdd gnd cell_6t
Xbit_r2_c71 bl[71] br[71] wl[2] vdd gnd cell_6t
Xbit_r3_c71 bl[71] br[71] wl[3] vdd gnd cell_6t
Xbit_r4_c71 bl[71] br[71] wl[4] vdd gnd cell_6t
Xbit_r5_c71 bl[71] br[71] wl[5] vdd gnd cell_6t
Xbit_r6_c71 bl[71] br[71] wl[6] vdd gnd cell_6t
Xbit_r7_c71 bl[71] br[71] wl[7] vdd gnd cell_6t
Xbit_r8_c71 bl[71] br[71] wl[8] vdd gnd cell_6t
Xbit_r9_c71 bl[71] br[71] wl[9] vdd gnd cell_6t
Xbit_r10_c71 bl[71] br[71] wl[10] vdd gnd cell_6t
Xbit_r11_c71 bl[71] br[71] wl[11] vdd gnd cell_6t
Xbit_r12_c71 bl[71] br[71] wl[12] vdd gnd cell_6t
Xbit_r13_c71 bl[71] br[71] wl[13] vdd gnd cell_6t
Xbit_r14_c71 bl[71] br[71] wl[14] vdd gnd cell_6t
Xbit_r15_c71 bl[71] br[71] wl[15] vdd gnd cell_6t
Xbit_r16_c71 bl[71] br[71] wl[16] vdd gnd cell_6t
Xbit_r17_c71 bl[71] br[71] wl[17] vdd gnd cell_6t
Xbit_r18_c71 bl[71] br[71] wl[18] vdd gnd cell_6t
Xbit_r19_c71 bl[71] br[71] wl[19] vdd gnd cell_6t
Xbit_r20_c71 bl[71] br[71] wl[20] vdd gnd cell_6t
Xbit_r21_c71 bl[71] br[71] wl[21] vdd gnd cell_6t
Xbit_r22_c71 bl[71] br[71] wl[22] vdd gnd cell_6t
Xbit_r23_c71 bl[71] br[71] wl[23] vdd gnd cell_6t
Xbit_r24_c71 bl[71] br[71] wl[24] vdd gnd cell_6t
Xbit_r25_c71 bl[71] br[71] wl[25] vdd gnd cell_6t
Xbit_r26_c71 bl[71] br[71] wl[26] vdd gnd cell_6t
Xbit_r27_c71 bl[71] br[71] wl[27] vdd gnd cell_6t
Xbit_r28_c71 bl[71] br[71] wl[28] vdd gnd cell_6t
Xbit_r29_c71 bl[71] br[71] wl[29] vdd gnd cell_6t
Xbit_r30_c71 bl[71] br[71] wl[30] vdd gnd cell_6t
Xbit_r31_c71 bl[71] br[71] wl[31] vdd gnd cell_6t
Xbit_r32_c71 bl[71] br[71] wl[32] vdd gnd cell_6t
Xbit_r33_c71 bl[71] br[71] wl[33] vdd gnd cell_6t
Xbit_r34_c71 bl[71] br[71] wl[34] vdd gnd cell_6t
Xbit_r35_c71 bl[71] br[71] wl[35] vdd gnd cell_6t
Xbit_r36_c71 bl[71] br[71] wl[36] vdd gnd cell_6t
Xbit_r37_c71 bl[71] br[71] wl[37] vdd gnd cell_6t
Xbit_r38_c71 bl[71] br[71] wl[38] vdd gnd cell_6t
Xbit_r39_c71 bl[71] br[71] wl[39] vdd gnd cell_6t
Xbit_r40_c71 bl[71] br[71] wl[40] vdd gnd cell_6t
Xbit_r41_c71 bl[71] br[71] wl[41] vdd gnd cell_6t
Xbit_r42_c71 bl[71] br[71] wl[42] vdd gnd cell_6t
Xbit_r43_c71 bl[71] br[71] wl[43] vdd gnd cell_6t
Xbit_r44_c71 bl[71] br[71] wl[44] vdd gnd cell_6t
Xbit_r45_c71 bl[71] br[71] wl[45] vdd gnd cell_6t
Xbit_r46_c71 bl[71] br[71] wl[46] vdd gnd cell_6t
Xbit_r47_c71 bl[71] br[71] wl[47] vdd gnd cell_6t
Xbit_r48_c71 bl[71] br[71] wl[48] vdd gnd cell_6t
Xbit_r49_c71 bl[71] br[71] wl[49] vdd gnd cell_6t
Xbit_r50_c71 bl[71] br[71] wl[50] vdd gnd cell_6t
Xbit_r51_c71 bl[71] br[71] wl[51] vdd gnd cell_6t
Xbit_r52_c71 bl[71] br[71] wl[52] vdd gnd cell_6t
Xbit_r53_c71 bl[71] br[71] wl[53] vdd gnd cell_6t
Xbit_r54_c71 bl[71] br[71] wl[54] vdd gnd cell_6t
Xbit_r55_c71 bl[71] br[71] wl[55] vdd gnd cell_6t
Xbit_r56_c71 bl[71] br[71] wl[56] vdd gnd cell_6t
Xbit_r57_c71 bl[71] br[71] wl[57] vdd gnd cell_6t
Xbit_r58_c71 bl[71] br[71] wl[58] vdd gnd cell_6t
Xbit_r59_c71 bl[71] br[71] wl[59] vdd gnd cell_6t
Xbit_r60_c71 bl[71] br[71] wl[60] vdd gnd cell_6t
Xbit_r61_c71 bl[71] br[71] wl[61] vdd gnd cell_6t
Xbit_r62_c71 bl[71] br[71] wl[62] vdd gnd cell_6t
Xbit_r63_c71 bl[71] br[71] wl[63] vdd gnd cell_6t
Xbit_r64_c71 bl[71] br[71] wl[64] vdd gnd cell_6t
Xbit_r65_c71 bl[71] br[71] wl[65] vdd gnd cell_6t
Xbit_r66_c71 bl[71] br[71] wl[66] vdd gnd cell_6t
Xbit_r67_c71 bl[71] br[71] wl[67] vdd gnd cell_6t
Xbit_r68_c71 bl[71] br[71] wl[68] vdd gnd cell_6t
Xbit_r69_c71 bl[71] br[71] wl[69] vdd gnd cell_6t
Xbit_r70_c71 bl[71] br[71] wl[70] vdd gnd cell_6t
Xbit_r71_c71 bl[71] br[71] wl[71] vdd gnd cell_6t
Xbit_r72_c71 bl[71] br[71] wl[72] vdd gnd cell_6t
Xbit_r73_c71 bl[71] br[71] wl[73] vdd gnd cell_6t
Xbit_r74_c71 bl[71] br[71] wl[74] vdd gnd cell_6t
Xbit_r75_c71 bl[71] br[71] wl[75] vdd gnd cell_6t
Xbit_r76_c71 bl[71] br[71] wl[76] vdd gnd cell_6t
Xbit_r77_c71 bl[71] br[71] wl[77] vdd gnd cell_6t
Xbit_r78_c71 bl[71] br[71] wl[78] vdd gnd cell_6t
Xbit_r79_c71 bl[71] br[71] wl[79] vdd gnd cell_6t
Xbit_r80_c71 bl[71] br[71] wl[80] vdd gnd cell_6t
Xbit_r81_c71 bl[71] br[71] wl[81] vdd gnd cell_6t
Xbit_r82_c71 bl[71] br[71] wl[82] vdd gnd cell_6t
Xbit_r83_c71 bl[71] br[71] wl[83] vdd gnd cell_6t
Xbit_r84_c71 bl[71] br[71] wl[84] vdd gnd cell_6t
Xbit_r85_c71 bl[71] br[71] wl[85] vdd gnd cell_6t
Xbit_r86_c71 bl[71] br[71] wl[86] vdd gnd cell_6t
Xbit_r87_c71 bl[71] br[71] wl[87] vdd gnd cell_6t
Xbit_r88_c71 bl[71] br[71] wl[88] vdd gnd cell_6t
Xbit_r89_c71 bl[71] br[71] wl[89] vdd gnd cell_6t
Xbit_r90_c71 bl[71] br[71] wl[90] vdd gnd cell_6t
Xbit_r91_c71 bl[71] br[71] wl[91] vdd gnd cell_6t
Xbit_r92_c71 bl[71] br[71] wl[92] vdd gnd cell_6t
Xbit_r93_c71 bl[71] br[71] wl[93] vdd gnd cell_6t
Xbit_r94_c71 bl[71] br[71] wl[94] vdd gnd cell_6t
Xbit_r95_c71 bl[71] br[71] wl[95] vdd gnd cell_6t
Xbit_r96_c71 bl[71] br[71] wl[96] vdd gnd cell_6t
Xbit_r97_c71 bl[71] br[71] wl[97] vdd gnd cell_6t
Xbit_r98_c71 bl[71] br[71] wl[98] vdd gnd cell_6t
Xbit_r99_c71 bl[71] br[71] wl[99] vdd gnd cell_6t
Xbit_r100_c71 bl[71] br[71] wl[100] vdd gnd cell_6t
Xbit_r101_c71 bl[71] br[71] wl[101] vdd gnd cell_6t
Xbit_r102_c71 bl[71] br[71] wl[102] vdd gnd cell_6t
Xbit_r103_c71 bl[71] br[71] wl[103] vdd gnd cell_6t
Xbit_r104_c71 bl[71] br[71] wl[104] vdd gnd cell_6t
Xbit_r105_c71 bl[71] br[71] wl[105] vdd gnd cell_6t
Xbit_r106_c71 bl[71] br[71] wl[106] vdd gnd cell_6t
Xbit_r107_c71 bl[71] br[71] wl[107] vdd gnd cell_6t
Xbit_r108_c71 bl[71] br[71] wl[108] vdd gnd cell_6t
Xbit_r109_c71 bl[71] br[71] wl[109] vdd gnd cell_6t
Xbit_r110_c71 bl[71] br[71] wl[110] vdd gnd cell_6t
Xbit_r111_c71 bl[71] br[71] wl[111] vdd gnd cell_6t
Xbit_r112_c71 bl[71] br[71] wl[112] vdd gnd cell_6t
Xbit_r113_c71 bl[71] br[71] wl[113] vdd gnd cell_6t
Xbit_r114_c71 bl[71] br[71] wl[114] vdd gnd cell_6t
Xbit_r115_c71 bl[71] br[71] wl[115] vdd gnd cell_6t
Xbit_r116_c71 bl[71] br[71] wl[116] vdd gnd cell_6t
Xbit_r117_c71 bl[71] br[71] wl[117] vdd gnd cell_6t
Xbit_r118_c71 bl[71] br[71] wl[118] vdd gnd cell_6t
Xbit_r119_c71 bl[71] br[71] wl[119] vdd gnd cell_6t
Xbit_r120_c71 bl[71] br[71] wl[120] vdd gnd cell_6t
Xbit_r121_c71 bl[71] br[71] wl[121] vdd gnd cell_6t
Xbit_r122_c71 bl[71] br[71] wl[122] vdd gnd cell_6t
Xbit_r123_c71 bl[71] br[71] wl[123] vdd gnd cell_6t
Xbit_r124_c71 bl[71] br[71] wl[124] vdd gnd cell_6t
Xbit_r125_c71 bl[71] br[71] wl[125] vdd gnd cell_6t
Xbit_r126_c71 bl[71] br[71] wl[126] vdd gnd cell_6t
Xbit_r127_c71 bl[71] br[71] wl[127] vdd gnd cell_6t
Xbit_r128_c71 bl[71] br[71] wl[128] vdd gnd cell_6t
Xbit_r129_c71 bl[71] br[71] wl[129] vdd gnd cell_6t
Xbit_r130_c71 bl[71] br[71] wl[130] vdd gnd cell_6t
Xbit_r131_c71 bl[71] br[71] wl[131] vdd gnd cell_6t
Xbit_r132_c71 bl[71] br[71] wl[132] vdd gnd cell_6t
Xbit_r133_c71 bl[71] br[71] wl[133] vdd gnd cell_6t
Xbit_r134_c71 bl[71] br[71] wl[134] vdd gnd cell_6t
Xbit_r135_c71 bl[71] br[71] wl[135] vdd gnd cell_6t
Xbit_r136_c71 bl[71] br[71] wl[136] vdd gnd cell_6t
Xbit_r137_c71 bl[71] br[71] wl[137] vdd gnd cell_6t
Xbit_r138_c71 bl[71] br[71] wl[138] vdd gnd cell_6t
Xbit_r139_c71 bl[71] br[71] wl[139] vdd gnd cell_6t
Xbit_r140_c71 bl[71] br[71] wl[140] vdd gnd cell_6t
Xbit_r141_c71 bl[71] br[71] wl[141] vdd gnd cell_6t
Xbit_r142_c71 bl[71] br[71] wl[142] vdd gnd cell_6t
Xbit_r143_c71 bl[71] br[71] wl[143] vdd gnd cell_6t
Xbit_r144_c71 bl[71] br[71] wl[144] vdd gnd cell_6t
Xbit_r145_c71 bl[71] br[71] wl[145] vdd gnd cell_6t
Xbit_r146_c71 bl[71] br[71] wl[146] vdd gnd cell_6t
Xbit_r147_c71 bl[71] br[71] wl[147] vdd gnd cell_6t
Xbit_r148_c71 bl[71] br[71] wl[148] vdd gnd cell_6t
Xbit_r149_c71 bl[71] br[71] wl[149] vdd gnd cell_6t
Xbit_r150_c71 bl[71] br[71] wl[150] vdd gnd cell_6t
Xbit_r151_c71 bl[71] br[71] wl[151] vdd gnd cell_6t
Xbit_r152_c71 bl[71] br[71] wl[152] vdd gnd cell_6t
Xbit_r153_c71 bl[71] br[71] wl[153] vdd gnd cell_6t
Xbit_r154_c71 bl[71] br[71] wl[154] vdd gnd cell_6t
Xbit_r155_c71 bl[71] br[71] wl[155] vdd gnd cell_6t
Xbit_r156_c71 bl[71] br[71] wl[156] vdd gnd cell_6t
Xbit_r157_c71 bl[71] br[71] wl[157] vdd gnd cell_6t
Xbit_r158_c71 bl[71] br[71] wl[158] vdd gnd cell_6t
Xbit_r159_c71 bl[71] br[71] wl[159] vdd gnd cell_6t
Xbit_r160_c71 bl[71] br[71] wl[160] vdd gnd cell_6t
Xbit_r161_c71 bl[71] br[71] wl[161] vdd gnd cell_6t
Xbit_r162_c71 bl[71] br[71] wl[162] vdd gnd cell_6t
Xbit_r163_c71 bl[71] br[71] wl[163] vdd gnd cell_6t
Xbit_r164_c71 bl[71] br[71] wl[164] vdd gnd cell_6t
Xbit_r165_c71 bl[71] br[71] wl[165] vdd gnd cell_6t
Xbit_r166_c71 bl[71] br[71] wl[166] vdd gnd cell_6t
Xbit_r167_c71 bl[71] br[71] wl[167] vdd gnd cell_6t
Xbit_r168_c71 bl[71] br[71] wl[168] vdd gnd cell_6t
Xbit_r169_c71 bl[71] br[71] wl[169] vdd gnd cell_6t
Xbit_r170_c71 bl[71] br[71] wl[170] vdd gnd cell_6t
Xbit_r171_c71 bl[71] br[71] wl[171] vdd gnd cell_6t
Xbit_r172_c71 bl[71] br[71] wl[172] vdd gnd cell_6t
Xbit_r173_c71 bl[71] br[71] wl[173] vdd gnd cell_6t
Xbit_r174_c71 bl[71] br[71] wl[174] vdd gnd cell_6t
Xbit_r175_c71 bl[71] br[71] wl[175] vdd gnd cell_6t
Xbit_r176_c71 bl[71] br[71] wl[176] vdd gnd cell_6t
Xbit_r177_c71 bl[71] br[71] wl[177] vdd gnd cell_6t
Xbit_r178_c71 bl[71] br[71] wl[178] vdd gnd cell_6t
Xbit_r179_c71 bl[71] br[71] wl[179] vdd gnd cell_6t
Xbit_r180_c71 bl[71] br[71] wl[180] vdd gnd cell_6t
Xbit_r181_c71 bl[71] br[71] wl[181] vdd gnd cell_6t
Xbit_r182_c71 bl[71] br[71] wl[182] vdd gnd cell_6t
Xbit_r183_c71 bl[71] br[71] wl[183] vdd gnd cell_6t
Xbit_r184_c71 bl[71] br[71] wl[184] vdd gnd cell_6t
Xbit_r185_c71 bl[71] br[71] wl[185] vdd gnd cell_6t
Xbit_r186_c71 bl[71] br[71] wl[186] vdd gnd cell_6t
Xbit_r187_c71 bl[71] br[71] wl[187] vdd gnd cell_6t
Xbit_r188_c71 bl[71] br[71] wl[188] vdd gnd cell_6t
Xbit_r189_c71 bl[71] br[71] wl[189] vdd gnd cell_6t
Xbit_r190_c71 bl[71] br[71] wl[190] vdd gnd cell_6t
Xbit_r191_c71 bl[71] br[71] wl[191] vdd gnd cell_6t
Xbit_r192_c71 bl[71] br[71] wl[192] vdd gnd cell_6t
Xbit_r193_c71 bl[71] br[71] wl[193] vdd gnd cell_6t
Xbit_r194_c71 bl[71] br[71] wl[194] vdd gnd cell_6t
Xbit_r195_c71 bl[71] br[71] wl[195] vdd gnd cell_6t
Xbit_r196_c71 bl[71] br[71] wl[196] vdd gnd cell_6t
Xbit_r197_c71 bl[71] br[71] wl[197] vdd gnd cell_6t
Xbit_r198_c71 bl[71] br[71] wl[198] vdd gnd cell_6t
Xbit_r199_c71 bl[71] br[71] wl[199] vdd gnd cell_6t
Xbit_r200_c71 bl[71] br[71] wl[200] vdd gnd cell_6t
Xbit_r201_c71 bl[71] br[71] wl[201] vdd gnd cell_6t
Xbit_r202_c71 bl[71] br[71] wl[202] vdd gnd cell_6t
Xbit_r203_c71 bl[71] br[71] wl[203] vdd gnd cell_6t
Xbit_r204_c71 bl[71] br[71] wl[204] vdd gnd cell_6t
Xbit_r205_c71 bl[71] br[71] wl[205] vdd gnd cell_6t
Xbit_r206_c71 bl[71] br[71] wl[206] vdd gnd cell_6t
Xbit_r207_c71 bl[71] br[71] wl[207] vdd gnd cell_6t
Xbit_r208_c71 bl[71] br[71] wl[208] vdd gnd cell_6t
Xbit_r209_c71 bl[71] br[71] wl[209] vdd gnd cell_6t
Xbit_r210_c71 bl[71] br[71] wl[210] vdd gnd cell_6t
Xbit_r211_c71 bl[71] br[71] wl[211] vdd gnd cell_6t
Xbit_r212_c71 bl[71] br[71] wl[212] vdd gnd cell_6t
Xbit_r213_c71 bl[71] br[71] wl[213] vdd gnd cell_6t
Xbit_r214_c71 bl[71] br[71] wl[214] vdd gnd cell_6t
Xbit_r215_c71 bl[71] br[71] wl[215] vdd gnd cell_6t
Xbit_r216_c71 bl[71] br[71] wl[216] vdd gnd cell_6t
Xbit_r217_c71 bl[71] br[71] wl[217] vdd gnd cell_6t
Xbit_r218_c71 bl[71] br[71] wl[218] vdd gnd cell_6t
Xbit_r219_c71 bl[71] br[71] wl[219] vdd gnd cell_6t
Xbit_r220_c71 bl[71] br[71] wl[220] vdd gnd cell_6t
Xbit_r221_c71 bl[71] br[71] wl[221] vdd gnd cell_6t
Xbit_r222_c71 bl[71] br[71] wl[222] vdd gnd cell_6t
Xbit_r223_c71 bl[71] br[71] wl[223] vdd gnd cell_6t
Xbit_r224_c71 bl[71] br[71] wl[224] vdd gnd cell_6t
Xbit_r225_c71 bl[71] br[71] wl[225] vdd gnd cell_6t
Xbit_r226_c71 bl[71] br[71] wl[226] vdd gnd cell_6t
Xbit_r227_c71 bl[71] br[71] wl[227] vdd gnd cell_6t
Xbit_r228_c71 bl[71] br[71] wl[228] vdd gnd cell_6t
Xbit_r229_c71 bl[71] br[71] wl[229] vdd gnd cell_6t
Xbit_r230_c71 bl[71] br[71] wl[230] vdd gnd cell_6t
Xbit_r231_c71 bl[71] br[71] wl[231] vdd gnd cell_6t
Xbit_r232_c71 bl[71] br[71] wl[232] vdd gnd cell_6t
Xbit_r233_c71 bl[71] br[71] wl[233] vdd gnd cell_6t
Xbit_r234_c71 bl[71] br[71] wl[234] vdd gnd cell_6t
Xbit_r235_c71 bl[71] br[71] wl[235] vdd gnd cell_6t
Xbit_r236_c71 bl[71] br[71] wl[236] vdd gnd cell_6t
Xbit_r237_c71 bl[71] br[71] wl[237] vdd gnd cell_6t
Xbit_r238_c71 bl[71] br[71] wl[238] vdd gnd cell_6t
Xbit_r239_c71 bl[71] br[71] wl[239] vdd gnd cell_6t
Xbit_r240_c71 bl[71] br[71] wl[240] vdd gnd cell_6t
Xbit_r241_c71 bl[71] br[71] wl[241] vdd gnd cell_6t
Xbit_r242_c71 bl[71] br[71] wl[242] vdd gnd cell_6t
Xbit_r243_c71 bl[71] br[71] wl[243] vdd gnd cell_6t
Xbit_r244_c71 bl[71] br[71] wl[244] vdd gnd cell_6t
Xbit_r245_c71 bl[71] br[71] wl[245] vdd gnd cell_6t
Xbit_r246_c71 bl[71] br[71] wl[246] vdd gnd cell_6t
Xbit_r247_c71 bl[71] br[71] wl[247] vdd gnd cell_6t
Xbit_r248_c71 bl[71] br[71] wl[248] vdd gnd cell_6t
Xbit_r249_c71 bl[71] br[71] wl[249] vdd gnd cell_6t
Xbit_r250_c71 bl[71] br[71] wl[250] vdd gnd cell_6t
Xbit_r251_c71 bl[71] br[71] wl[251] vdd gnd cell_6t
Xbit_r252_c71 bl[71] br[71] wl[252] vdd gnd cell_6t
Xbit_r253_c71 bl[71] br[71] wl[253] vdd gnd cell_6t
Xbit_r254_c71 bl[71] br[71] wl[254] vdd gnd cell_6t
Xbit_r255_c71 bl[71] br[71] wl[255] vdd gnd cell_6t
Xbit_r256_c71 bl[71] br[71] wl[256] vdd gnd cell_6t
Xbit_r257_c71 bl[71] br[71] wl[257] vdd gnd cell_6t
Xbit_r258_c71 bl[71] br[71] wl[258] vdd gnd cell_6t
Xbit_r259_c71 bl[71] br[71] wl[259] vdd gnd cell_6t
Xbit_r260_c71 bl[71] br[71] wl[260] vdd gnd cell_6t
Xbit_r261_c71 bl[71] br[71] wl[261] vdd gnd cell_6t
Xbit_r262_c71 bl[71] br[71] wl[262] vdd gnd cell_6t
Xbit_r263_c71 bl[71] br[71] wl[263] vdd gnd cell_6t
Xbit_r264_c71 bl[71] br[71] wl[264] vdd gnd cell_6t
Xbit_r265_c71 bl[71] br[71] wl[265] vdd gnd cell_6t
Xbit_r266_c71 bl[71] br[71] wl[266] vdd gnd cell_6t
Xbit_r267_c71 bl[71] br[71] wl[267] vdd gnd cell_6t
Xbit_r268_c71 bl[71] br[71] wl[268] vdd gnd cell_6t
Xbit_r269_c71 bl[71] br[71] wl[269] vdd gnd cell_6t
Xbit_r270_c71 bl[71] br[71] wl[270] vdd gnd cell_6t
Xbit_r271_c71 bl[71] br[71] wl[271] vdd gnd cell_6t
Xbit_r272_c71 bl[71] br[71] wl[272] vdd gnd cell_6t
Xbit_r273_c71 bl[71] br[71] wl[273] vdd gnd cell_6t
Xbit_r274_c71 bl[71] br[71] wl[274] vdd gnd cell_6t
Xbit_r275_c71 bl[71] br[71] wl[275] vdd gnd cell_6t
Xbit_r276_c71 bl[71] br[71] wl[276] vdd gnd cell_6t
Xbit_r277_c71 bl[71] br[71] wl[277] vdd gnd cell_6t
Xbit_r278_c71 bl[71] br[71] wl[278] vdd gnd cell_6t
Xbit_r279_c71 bl[71] br[71] wl[279] vdd gnd cell_6t
Xbit_r280_c71 bl[71] br[71] wl[280] vdd gnd cell_6t
Xbit_r281_c71 bl[71] br[71] wl[281] vdd gnd cell_6t
Xbit_r282_c71 bl[71] br[71] wl[282] vdd gnd cell_6t
Xbit_r283_c71 bl[71] br[71] wl[283] vdd gnd cell_6t
Xbit_r284_c71 bl[71] br[71] wl[284] vdd gnd cell_6t
Xbit_r285_c71 bl[71] br[71] wl[285] vdd gnd cell_6t
Xbit_r286_c71 bl[71] br[71] wl[286] vdd gnd cell_6t
Xbit_r287_c71 bl[71] br[71] wl[287] vdd gnd cell_6t
Xbit_r288_c71 bl[71] br[71] wl[288] vdd gnd cell_6t
Xbit_r289_c71 bl[71] br[71] wl[289] vdd gnd cell_6t
Xbit_r290_c71 bl[71] br[71] wl[290] vdd gnd cell_6t
Xbit_r291_c71 bl[71] br[71] wl[291] vdd gnd cell_6t
Xbit_r292_c71 bl[71] br[71] wl[292] vdd gnd cell_6t
Xbit_r293_c71 bl[71] br[71] wl[293] vdd gnd cell_6t
Xbit_r294_c71 bl[71] br[71] wl[294] vdd gnd cell_6t
Xbit_r295_c71 bl[71] br[71] wl[295] vdd gnd cell_6t
Xbit_r296_c71 bl[71] br[71] wl[296] vdd gnd cell_6t
Xbit_r297_c71 bl[71] br[71] wl[297] vdd gnd cell_6t
Xbit_r298_c71 bl[71] br[71] wl[298] vdd gnd cell_6t
Xbit_r299_c71 bl[71] br[71] wl[299] vdd gnd cell_6t
Xbit_r300_c71 bl[71] br[71] wl[300] vdd gnd cell_6t
Xbit_r301_c71 bl[71] br[71] wl[301] vdd gnd cell_6t
Xbit_r302_c71 bl[71] br[71] wl[302] vdd gnd cell_6t
Xbit_r303_c71 bl[71] br[71] wl[303] vdd gnd cell_6t
Xbit_r304_c71 bl[71] br[71] wl[304] vdd gnd cell_6t
Xbit_r305_c71 bl[71] br[71] wl[305] vdd gnd cell_6t
Xbit_r306_c71 bl[71] br[71] wl[306] vdd gnd cell_6t
Xbit_r307_c71 bl[71] br[71] wl[307] vdd gnd cell_6t
Xbit_r308_c71 bl[71] br[71] wl[308] vdd gnd cell_6t
Xbit_r309_c71 bl[71] br[71] wl[309] vdd gnd cell_6t
Xbit_r310_c71 bl[71] br[71] wl[310] vdd gnd cell_6t
Xbit_r311_c71 bl[71] br[71] wl[311] vdd gnd cell_6t
Xbit_r312_c71 bl[71] br[71] wl[312] vdd gnd cell_6t
Xbit_r313_c71 bl[71] br[71] wl[313] vdd gnd cell_6t
Xbit_r314_c71 bl[71] br[71] wl[314] vdd gnd cell_6t
Xbit_r315_c71 bl[71] br[71] wl[315] vdd gnd cell_6t
Xbit_r316_c71 bl[71] br[71] wl[316] vdd gnd cell_6t
Xbit_r317_c71 bl[71] br[71] wl[317] vdd gnd cell_6t
Xbit_r318_c71 bl[71] br[71] wl[318] vdd gnd cell_6t
Xbit_r319_c71 bl[71] br[71] wl[319] vdd gnd cell_6t
Xbit_r320_c71 bl[71] br[71] wl[320] vdd gnd cell_6t
Xbit_r321_c71 bl[71] br[71] wl[321] vdd gnd cell_6t
Xbit_r322_c71 bl[71] br[71] wl[322] vdd gnd cell_6t
Xbit_r323_c71 bl[71] br[71] wl[323] vdd gnd cell_6t
Xbit_r324_c71 bl[71] br[71] wl[324] vdd gnd cell_6t
Xbit_r325_c71 bl[71] br[71] wl[325] vdd gnd cell_6t
Xbit_r326_c71 bl[71] br[71] wl[326] vdd gnd cell_6t
Xbit_r327_c71 bl[71] br[71] wl[327] vdd gnd cell_6t
Xbit_r328_c71 bl[71] br[71] wl[328] vdd gnd cell_6t
Xbit_r329_c71 bl[71] br[71] wl[329] vdd gnd cell_6t
Xbit_r330_c71 bl[71] br[71] wl[330] vdd gnd cell_6t
Xbit_r331_c71 bl[71] br[71] wl[331] vdd gnd cell_6t
Xbit_r332_c71 bl[71] br[71] wl[332] vdd gnd cell_6t
Xbit_r333_c71 bl[71] br[71] wl[333] vdd gnd cell_6t
Xbit_r334_c71 bl[71] br[71] wl[334] vdd gnd cell_6t
Xbit_r335_c71 bl[71] br[71] wl[335] vdd gnd cell_6t
Xbit_r336_c71 bl[71] br[71] wl[336] vdd gnd cell_6t
Xbit_r337_c71 bl[71] br[71] wl[337] vdd gnd cell_6t
Xbit_r338_c71 bl[71] br[71] wl[338] vdd gnd cell_6t
Xbit_r339_c71 bl[71] br[71] wl[339] vdd gnd cell_6t
Xbit_r340_c71 bl[71] br[71] wl[340] vdd gnd cell_6t
Xbit_r341_c71 bl[71] br[71] wl[341] vdd gnd cell_6t
Xbit_r342_c71 bl[71] br[71] wl[342] vdd gnd cell_6t
Xbit_r343_c71 bl[71] br[71] wl[343] vdd gnd cell_6t
Xbit_r344_c71 bl[71] br[71] wl[344] vdd gnd cell_6t
Xbit_r345_c71 bl[71] br[71] wl[345] vdd gnd cell_6t
Xbit_r346_c71 bl[71] br[71] wl[346] vdd gnd cell_6t
Xbit_r347_c71 bl[71] br[71] wl[347] vdd gnd cell_6t
Xbit_r348_c71 bl[71] br[71] wl[348] vdd gnd cell_6t
Xbit_r349_c71 bl[71] br[71] wl[349] vdd gnd cell_6t
Xbit_r350_c71 bl[71] br[71] wl[350] vdd gnd cell_6t
Xbit_r351_c71 bl[71] br[71] wl[351] vdd gnd cell_6t
Xbit_r352_c71 bl[71] br[71] wl[352] vdd gnd cell_6t
Xbit_r353_c71 bl[71] br[71] wl[353] vdd gnd cell_6t
Xbit_r354_c71 bl[71] br[71] wl[354] vdd gnd cell_6t
Xbit_r355_c71 bl[71] br[71] wl[355] vdd gnd cell_6t
Xbit_r356_c71 bl[71] br[71] wl[356] vdd gnd cell_6t
Xbit_r357_c71 bl[71] br[71] wl[357] vdd gnd cell_6t
Xbit_r358_c71 bl[71] br[71] wl[358] vdd gnd cell_6t
Xbit_r359_c71 bl[71] br[71] wl[359] vdd gnd cell_6t
Xbit_r360_c71 bl[71] br[71] wl[360] vdd gnd cell_6t
Xbit_r361_c71 bl[71] br[71] wl[361] vdd gnd cell_6t
Xbit_r362_c71 bl[71] br[71] wl[362] vdd gnd cell_6t
Xbit_r363_c71 bl[71] br[71] wl[363] vdd gnd cell_6t
Xbit_r364_c71 bl[71] br[71] wl[364] vdd gnd cell_6t
Xbit_r365_c71 bl[71] br[71] wl[365] vdd gnd cell_6t
Xbit_r366_c71 bl[71] br[71] wl[366] vdd gnd cell_6t
Xbit_r367_c71 bl[71] br[71] wl[367] vdd gnd cell_6t
Xbit_r368_c71 bl[71] br[71] wl[368] vdd gnd cell_6t
Xbit_r369_c71 bl[71] br[71] wl[369] vdd gnd cell_6t
Xbit_r370_c71 bl[71] br[71] wl[370] vdd gnd cell_6t
Xbit_r371_c71 bl[71] br[71] wl[371] vdd gnd cell_6t
Xbit_r372_c71 bl[71] br[71] wl[372] vdd gnd cell_6t
Xbit_r373_c71 bl[71] br[71] wl[373] vdd gnd cell_6t
Xbit_r374_c71 bl[71] br[71] wl[374] vdd gnd cell_6t
Xbit_r375_c71 bl[71] br[71] wl[375] vdd gnd cell_6t
Xbit_r376_c71 bl[71] br[71] wl[376] vdd gnd cell_6t
Xbit_r377_c71 bl[71] br[71] wl[377] vdd gnd cell_6t
Xbit_r378_c71 bl[71] br[71] wl[378] vdd gnd cell_6t
Xbit_r379_c71 bl[71] br[71] wl[379] vdd gnd cell_6t
Xbit_r380_c71 bl[71] br[71] wl[380] vdd gnd cell_6t
Xbit_r381_c71 bl[71] br[71] wl[381] vdd gnd cell_6t
Xbit_r382_c71 bl[71] br[71] wl[382] vdd gnd cell_6t
Xbit_r383_c71 bl[71] br[71] wl[383] vdd gnd cell_6t
Xbit_r384_c71 bl[71] br[71] wl[384] vdd gnd cell_6t
Xbit_r385_c71 bl[71] br[71] wl[385] vdd gnd cell_6t
Xbit_r386_c71 bl[71] br[71] wl[386] vdd gnd cell_6t
Xbit_r387_c71 bl[71] br[71] wl[387] vdd gnd cell_6t
Xbit_r388_c71 bl[71] br[71] wl[388] vdd gnd cell_6t
Xbit_r389_c71 bl[71] br[71] wl[389] vdd gnd cell_6t
Xbit_r390_c71 bl[71] br[71] wl[390] vdd gnd cell_6t
Xbit_r391_c71 bl[71] br[71] wl[391] vdd gnd cell_6t
Xbit_r392_c71 bl[71] br[71] wl[392] vdd gnd cell_6t
Xbit_r393_c71 bl[71] br[71] wl[393] vdd gnd cell_6t
Xbit_r394_c71 bl[71] br[71] wl[394] vdd gnd cell_6t
Xbit_r395_c71 bl[71] br[71] wl[395] vdd gnd cell_6t
Xbit_r396_c71 bl[71] br[71] wl[396] vdd gnd cell_6t
Xbit_r397_c71 bl[71] br[71] wl[397] vdd gnd cell_6t
Xbit_r398_c71 bl[71] br[71] wl[398] vdd gnd cell_6t
Xbit_r399_c71 bl[71] br[71] wl[399] vdd gnd cell_6t
Xbit_r400_c71 bl[71] br[71] wl[400] vdd gnd cell_6t
Xbit_r401_c71 bl[71] br[71] wl[401] vdd gnd cell_6t
Xbit_r402_c71 bl[71] br[71] wl[402] vdd gnd cell_6t
Xbit_r403_c71 bl[71] br[71] wl[403] vdd gnd cell_6t
Xbit_r404_c71 bl[71] br[71] wl[404] vdd gnd cell_6t
Xbit_r405_c71 bl[71] br[71] wl[405] vdd gnd cell_6t
Xbit_r406_c71 bl[71] br[71] wl[406] vdd gnd cell_6t
Xbit_r407_c71 bl[71] br[71] wl[407] vdd gnd cell_6t
Xbit_r408_c71 bl[71] br[71] wl[408] vdd gnd cell_6t
Xbit_r409_c71 bl[71] br[71] wl[409] vdd gnd cell_6t
Xbit_r410_c71 bl[71] br[71] wl[410] vdd gnd cell_6t
Xbit_r411_c71 bl[71] br[71] wl[411] vdd gnd cell_6t
Xbit_r412_c71 bl[71] br[71] wl[412] vdd gnd cell_6t
Xbit_r413_c71 bl[71] br[71] wl[413] vdd gnd cell_6t
Xbit_r414_c71 bl[71] br[71] wl[414] vdd gnd cell_6t
Xbit_r415_c71 bl[71] br[71] wl[415] vdd gnd cell_6t
Xbit_r416_c71 bl[71] br[71] wl[416] vdd gnd cell_6t
Xbit_r417_c71 bl[71] br[71] wl[417] vdd gnd cell_6t
Xbit_r418_c71 bl[71] br[71] wl[418] vdd gnd cell_6t
Xbit_r419_c71 bl[71] br[71] wl[419] vdd gnd cell_6t
Xbit_r420_c71 bl[71] br[71] wl[420] vdd gnd cell_6t
Xbit_r421_c71 bl[71] br[71] wl[421] vdd gnd cell_6t
Xbit_r422_c71 bl[71] br[71] wl[422] vdd gnd cell_6t
Xbit_r423_c71 bl[71] br[71] wl[423] vdd gnd cell_6t
Xbit_r424_c71 bl[71] br[71] wl[424] vdd gnd cell_6t
Xbit_r425_c71 bl[71] br[71] wl[425] vdd gnd cell_6t
Xbit_r426_c71 bl[71] br[71] wl[426] vdd gnd cell_6t
Xbit_r427_c71 bl[71] br[71] wl[427] vdd gnd cell_6t
Xbit_r428_c71 bl[71] br[71] wl[428] vdd gnd cell_6t
Xbit_r429_c71 bl[71] br[71] wl[429] vdd gnd cell_6t
Xbit_r430_c71 bl[71] br[71] wl[430] vdd gnd cell_6t
Xbit_r431_c71 bl[71] br[71] wl[431] vdd gnd cell_6t
Xbit_r432_c71 bl[71] br[71] wl[432] vdd gnd cell_6t
Xbit_r433_c71 bl[71] br[71] wl[433] vdd gnd cell_6t
Xbit_r434_c71 bl[71] br[71] wl[434] vdd gnd cell_6t
Xbit_r435_c71 bl[71] br[71] wl[435] vdd gnd cell_6t
Xbit_r436_c71 bl[71] br[71] wl[436] vdd gnd cell_6t
Xbit_r437_c71 bl[71] br[71] wl[437] vdd gnd cell_6t
Xbit_r438_c71 bl[71] br[71] wl[438] vdd gnd cell_6t
Xbit_r439_c71 bl[71] br[71] wl[439] vdd gnd cell_6t
Xbit_r440_c71 bl[71] br[71] wl[440] vdd gnd cell_6t
Xbit_r441_c71 bl[71] br[71] wl[441] vdd gnd cell_6t
Xbit_r442_c71 bl[71] br[71] wl[442] vdd gnd cell_6t
Xbit_r443_c71 bl[71] br[71] wl[443] vdd gnd cell_6t
Xbit_r444_c71 bl[71] br[71] wl[444] vdd gnd cell_6t
Xbit_r445_c71 bl[71] br[71] wl[445] vdd gnd cell_6t
Xbit_r446_c71 bl[71] br[71] wl[446] vdd gnd cell_6t
Xbit_r447_c71 bl[71] br[71] wl[447] vdd gnd cell_6t
Xbit_r448_c71 bl[71] br[71] wl[448] vdd gnd cell_6t
Xbit_r449_c71 bl[71] br[71] wl[449] vdd gnd cell_6t
Xbit_r450_c71 bl[71] br[71] wl[450] vdd gnd cell_6t
Xbit_r451_c71 bl[71] br[71] wl[451] vdd gnd cell_6t
Xbit_r452_c71 bl[71] br[71] wl[452] vdd gnd cell_6t
Xbit_r453_c71 bl[71] br[71] wl[453] vdd gnd cell_6t
Xbit_r454_c71 bl[71] br[71] wl[454] vdd gnd cell_6t
Xbit_r455_c71 bl[71] br[71] wl[455] vdd gnd cell_6t
Xbit_r456_c71 bl[71] br[71] wl[456] vdd gnd cell_6t
Xbit_r457_c71 bl[71] br[71] wl[457] vdd gnd cell_6t
Xbit_r458_c71 bl[71] br[71] wl[458] vdd gnd cell_6t
Xbit_r459_c71 bl[71] br[71] wl[459] vdd gnd cell_6t
Xbit_r460_c71 bl[71] br[71] wl[460] vdd gnd cell_6t
Xbit_r461_c71 bl[71] br[71] wl[461] vdd gnd cell_6t
Xbit_r462_c71 bl[71] br[71] wl[462] vdd gnd cell_6t
Xbit_r463_c71 bl[71] br[71] wl[463] vdd gnd cell_6t
Xbit_r464_c71 bl[71] br[71] wl[464] vdd gnd cell_6t
Xbit_r465_c71 bl[71] br[71] wl[465] vdd gnd cell_6t
Xbit_r466_c71 bl[71] br[71] wl[466] vdd gnd cell_6t
Xbit_r467_c71 bl[71] br[71] wl[467] vdd gnd cell_6t
Xbit_r468_c71 bl[71] br[71] wl[468] vdd gnd cell_6t
Xbit_r469_c71 bl[71] br[71] wl[469] vdd gnd cell_6t
Xbit_r470_c71 bl[71] br[71] wl[470] vdd gnd cell_6t
Xbit_r471_c71 bl[71] br[71] wl[471] vdd gnd cell_6t
Xbit_r472_c71 bl[71] br[71] wl[472] vdd gnd cell_6t
Xbit_r473_c71 bl[71] br[71] wl[473] vdd gnd cell_6t
Xbit_r474_c71 bl[71] br[71] wl[474] vdd gnd cell_6t
Xbit_r475_c71 bl[71] br[71] wl[475] vdd gnd cell_6t
Xbit_r476_c71 bl[71] br[71] wl[476] vdd gnd cell_6t
Xbit_r477_c71 bl[71] br[71] wl[477] vdd gnd cell_6t
Xbit_r478_c71 bl[71] br[71] wl[478] vdd gnd cell_6t
Xbit_r479_c71 bl[71] br[71] wl[479] vdd gnd cell_6t
Xbit_r480_c71 bl[71] br[71] wl[480] vdd gnd cell_6t
Xbit_r481_c71 bl[71] br[71] wl[481] vdd gnd cell_6t
Xbit_r482_c71 bl[71] br[71] wl[482] vdd gnd cell_6t
Xbit_r483_c71 bl[71] br[71] wl[483] vdd gnd cell_6t
Xbit_r484_c71 bl[71] br[71] wl[484] vdd gnd cell_6t
Xbit_r485_c71 bl[71] br[71] wl[485] vdd gnd cell_6t
Xbit_r486_c71 bl[71] br[71] wl[486] vdd gnd cell_6t
Xbit_r487_c71 bl[71] br[71] wl[487] vdd gnd cell_6t
Xbit_r488_c71 bl[71] br[71] wl[488] vdd gnd cell_6t
Xbit_r489_c71 bl[71] br[71] wl[489] vdd gnd cell_6t
Xbit_r490_c71 bl[71] br[71] wl[490] vdd gnd cell_6t
Xbit_r491_c71 bl[71] br[71] wl[491] vdd gnd cell_6t
Xbit_r492_c71 bl[71] br[71] wl[492] vdd gnd cell_6t
Xbit_r493_c71 bl[71] br[71] wl[493] vdd gnd cell_6t
Xbit_r494_c71 bl[71] br[71] wl[494] vdd gnd cell_6t
Xbit_r495_c71 bl[71] br[71] wl[495] vdd gnd cell_6t
Xbit_r496_c71 bl[71] br[71] wl[496] vdd gnd cell_6t
Xbit_r497_c71 bl[71] br[71] wl[497] vdd gnd cell_6t
Xbit_r498_c71 bl[71] br[71] wl[498] vdd gnd cell_6t
Xbit_r499_c71 bl[71] br[71] wl[499] vdd gnd cell_6t
Xbit_r500_c71 bl[71] br[71] wl[500] vdd gnd cell_6t
Xbit_r501_c71 bl[71] br[71] wl[501] vdd gnd cell_6t
Xbit_r502_c71 bl[71] br[71] wl[502] vdd gnd cell_6t
Xbit_r503_c71 bl[71] br[71] wl[503] vdd gnd cell_6t
Xbit_r504_c71 bl[71] br[71] wl[504] vdd gnd cell_6t
Xbit_r505_c71 bl[71] br[71] wl[505] vdd gnd cell_6t
Xbit_r506_c71 bl[71] br[71] wl[506] vdd gnd cell_6t
Xbit_r507_c71 bl[71] br[71] wl[507] vdd gnd cell_6t
Xbit_r508_c71 bl[71] br[71] wl[508] vdd gnd cell_6t
Xbit_r509_c71 bl[71] br[71] wl[509] vdd gnd cell_6t
Xbit_r510_c71 bl[71] br[71] wl[510] vdd gnd cell_6t
Xbit_r511_c71 bl[71] br[71] wl[511] vdd gnd cell_6t
Xbit_r0_c72 bl[72] br[72] wl[0] vdd gnd cell_6t
Xbit_r1_c72 bl[72] br[72] wl[1] vdd gnd cell_6t
Xbit_r2_c72 bl[72] br[72] wl[2] vdd gnd cell_6t
Xbit_r3_c72 bl[72] br[72] wl[3] vdd gnd cell_6t
Xbit_r4_c72 bl[72] br[72] wl[4] vdd gnd cell_6t
Xbit_r5_c72 bl[72] br[72] wl[5] vdd gnd cell_6t
Xbit_r6_c72 bl[72] br[72] wl[6] vdd gnd cell_6t
Xbit_r7_c72 bl[72] br[72] wl[7] vdd gnd cell_6t
Xbit_r8_c72 bl[72] br[72] wl[8] vdd gnd cell_6t
Xbit_r9_c72 bl[72] br[72] wl[9] vdd gnd cell_6t
Xbit_r10_c72 bl[72] br[72] wl[10] vdd gnd cell_6t
Xbit_r11_c72 bl[72] br[72] wl[11] vdd gnd cell_6t
Xbit_r12_c72 bl[72] br[72] wl[12] vdd gnd cell_6t
Xbit_r13_c72 bl[72] br[72] wl[13] vdd gnd cell_6t
Xbit_r14_c72 bl[72] br[72] wl[14] vdd gnd cell_6t
Xbit_r15_c72 bl[72] br[72] wl[15] vdd gnd cell_6t
Xbit_r16_c72 bl[72] br[72] wl[16] vdd gnd cell_6t
Xbit_r17_c72 bl[72] br[72] wl[17] vdd gnd cell_6t
Xbit_r18_c72 bl[72] br[72] wl[18] vdd gnd cell_6t
Xbit_r19_c72 bl[72] br[72] wl[19] vdd gnd cell_6t
Xbit_r20_c72 bl[72] br[72] wl[20] vdd gnd cell_6t
Xbit_r21_c72 bl[72] br[72] wl[21] vdd gnd cell_6t
Xbit_r22_c72 bl[72] br[72] wl[22] vdd gnd cell_6t
Xbit_r23_c72 bl[72] br[72] wl[23] vdd gnd cell_6t
Xbit_r24_c72 bl[72] br[72] wl[24] vdd gnd cell_6t
Xbit_r25_c72 bl[72] br[72] wl[25] vdd gnd cell_6t
Xbit_r26_c72 bl[72] br[72] wl[26] vdd gnd cell_6t
Xbit_r27_c72 bl[72] br[72] wl[27] vdd gnd cell_6t
Xbit_r28_c72 bl[72] br[72] wl[28] vdd gnd cell_6t
Xbit_r29_c72 bl[72] br[72] wl[29] vdd gnd cell_6t
Xbit_r30_c72 bl[72] br[72] wl[30] vdd gnd cell_6t
Xbit_r31_c72 bl[72] br[72] wl[31] vdd gnd cell_6t
Xbit_r32_c72 bl[72] br[72] wl[32] vdd gnd cell_6t
Xbit_r33_c72 bl[72] br[72] wl[33] vdd gnd cell_6t
Xbit_r34_c72 bl[72] br[72] wl[34] vdd gnd cell_6t
Xbit_r35_c72 bl[72] br[72] wl[35] vdd gnd cell_6t
Xbit_r36_c72 bl[72] br[72] wl[36] vdd gnd cell_6t
Xbit_r37_c72 bl[72] br[72] wl[37] vdd gnd cell_6t
Xbit_r38_c72 bl[72] br[72] wl[38] vdd gnd cell_6t
Xbit_r39_c72 bl[72] br[72] wl[39] vdd gnd cell_6t
Xbit_r40_c72 bl[72] br[72] wl[40] vdd gnd cell_6t
Xbit_r41_c72 bl[72] br[72] wl[41] vdd gnd cell_6t
Xbit_r42_c72 bl[72] br[72] wl[42] vdd gnd cell_6t
Xbit_r43_c72 bl[72] br[72] wl[43] vdd gnd cell_6t
Xbit_r44_c72 bl[72] br[72] wl[44] vdd gnd cell_6t
Xbit_r45_c72 bl[72] br[72] wl[45] vdd gnd cell_6t
Xbit_r46_c72 bl[72] br[72] wl[46] vdd gnd cell_6t
Xbit_r47_c72 bl[72] br[72] wl[47] vdd gnd cell_6t
Xbit_r48_c72 bl[72] br[72] wl[48] vdd gnd cell_6t
Xbit_r49_c72 bl[72] br[72] wl[49] vdd gnd cell_6t
Xbit_r50_c72 bl[72] br[72] wl[50] vdd gnd cell_6t
Xbit_r51_c72 bl[72] br[72] wl[51] vdd gnd cell_6t
Xbit_r52_c72 bl[72] br[72] wl[52] vdd gnd cell_6t
Xbit_r53_c72 bl[72] br[72] wl[53] vdd gnd cell_6t
Xbit_r54_c72 bl[72] br[72] wl[54] vdd gnd cell_6t
Xbit_r55_c72 bl[72] br[72] wl[55] vdd gnd cell_6t
Xbit_r56_c72 bl[72] br[72] wl[56] vdd gnd cell_6t
Xbit_r57_c72 bl[72] br[72] wl[57] vdd gnd cell_6t
Xbit_r58_c72 bl[72] br[72] wl[58] vdd gnd cell_6t
Xbit_r59_c72 bl[72] br[72] wl[59] vdd gnd cell_6t
Xbit_r60_c72 bl[72] br[72] wl[60] vdd gnd cell_6t
Xbit_r61_c72 bl[72] br[72] wl[61] vdd gnd cell_6t
Xbit_r62_c72 bl[72] br[72] wl[62] vdd gnd cell_6t
Xbit_r63_c72 bl[72] br[72] wl[63] vdd gnd cell_6t
Xbit_r64_c72 bl[72] br[72] wl[64] vdd gnd cell_6t
Xbit_r65_c72 bl[72] br[72] wl[65] vdd gnd cell_6t
Xbit_r66_c72 bl[72] br[72] wl[66] vdd gnd cell_6t
Xbit_r67_c72 bl[72] br[72] wl[67] vdd gnd cell_6t
Xbit_r68_c72 bl[72] br[72] wl[68] vdd gnd cell_6t
Xbit_r69_c72 bl[72] br[72] wl[69] vdd gnd cell_6t
Xbit_r70_c72 bl[72] br[72] wl[70] vdd gnd cell_6t
Xbit_r71_c72 bl[72] br[72] wl[71] vdd gnd cell_6t
Xbit_r72_c72 bl[72] br[72] wl[72] vdd gnd cell_6t
Xbit_r73_c72 bl[72] br[72] wl[73] vdd gnd cell_6t
Xbit_r74_c72 bl[72] br[72] wl[74] vdd gnd cell_6t
Xbit_r75_c72 bl[72] br[72] wl[75] vdd gnd cell_6t
Xbit_r76_c72 bl[72] br[72] wl[76] vdd gnd cell_6t
Xbit_r77_c72 bl[72] br[72] wl[77] vdd gnd cell_6t
Xbit_r78_c72 bl[72] br[72] wl[78] vdd gnd cell_6t
Xbit_r79_c72 bl[72] br[72] wl[79] vdd gnd cell_6t
Xbit_r80_c72 bl[72] br[72] wl[80] vdd gnd cell_6t
Xbit_r81_c72 bl[72] br[72] wl[81] vdd gnd cell_6t
Xbit_r82_c72 bl[72] br[72] wl[82] vdd gnd cell_6t
Xbit_r83_c72 bl[72] br[72] wl[83] vdd gnd cell_6t
Xbit_r84_c72 bl[72] br[72] wl[84] vdd gnd cell_6t
Xbit_r85_c72 bl[72] br[72] wl[85] vdd gnd cell_6t
Xbit_r86_c72 bl[72] br[72] wl[86] vdd gnd cell_6t
Xbit_r87_c72 bl[72] br[72] wl[87] vdd gnd cell_6t
Xbit_r88_c72 bl[72] br[72] wl[88] vdd gnd cell_6t
Xbit_r89_c72 bl[72] br[72] wl[89] vdd gnd cell_6t
Xbit_r90_c72 bl[72] br[72] wl[90] vdd gnd cell_6t
Xbit_r91_c72 bl[72] br[72] wl[91] vdd gnd cell_6t
Xbit_r92_c72 bl[72] br[72] wl[92] vdd gnd cell_6t
Xbit_r93_c72 bl[72] br[72] wl[93] vdd gnd cell_6t
Xbit_r94_c72 bl[72] br[72] wl[94] vdd gnd cell_6t
Xbit_r95_c72 bl[72] br[72] wl[95] vdd gnd cell_6t
Xbit_r96_c72 bl[72] br[72] wl[96] vdd gnd cell_6t
Xbit_r97_c72 bl[72] br[72] wl[97] vdd gnd cell_6t
Xbit_r98_c72 bl[72] br[72] wl[98] vdd gnd cell_6t
Xbit_r99_c72 bl[72] br[72] wl[99] vdd gnd cell_6t
Xbit_r100_c72 bl[72] br[72] wl[100] vdd gnd cell_6t
Xbit_r101_c72 bl[72] br[72] wl[101] vdd gnd cell_6t
Xbit_r102_c72 bl[72] br[72] wl[102] vdd gnd cell_6t
Xbit_r103_c72 bl[72] br[72] wl[103] vdd gnd cell_6t
Xbit_r104_c72 bl[72] br[72] wl[104] vdd gnd cell_6t
Xbit_r105_c72 bl[72] br[72] wl[105] vdd gnd cell_6t
Xbit_r106_c72 bl[72] br[72] wl[106] vdd gnd cell_6t
Xbit_r107_c72 bl[72] br[72] wl[107] vdd gnd cell_6t
Xbit_r108_c72 bl[72] br[72] wl[108] vdd gnd cell_6t
Xbit_r109_c72 bl[72] br[72] wl[109] vdd gnd cell_6t
Xbit_r110_c72 bl[72] br[72] wl[110] vdd gnd cell_6t
Xbit_r111_c72 bl[72] br[72] wl[111] vdd gnd cell_6t
Xbit_r112_c72 bl[72] br[72] wl[112] vdd gnd cell_6t
Xbit_r113_c72 bl[72] br[72] wl[113] vdd gnd cell_6t
Xbit_r114_c72 bl[72] br[72] wl[114] vdd gnd cell_6t
Xbit_r115_c72 bl[72] br[72] wl[115] vdd gnd cell_6t
Xbit_r116_c72 bl[72] br[72] wl[116] vdd gnd cell_6t
Xbit_r117_c72 bl[72] br[72] wl[117] vdd gnd cell_6t
Xbit_r118_c72 bl[72] br[72] wl[118] vdd gnd cell_6t
Xbit_r119_c72 bl[72] br[72] wl[119] vdd gnd cell_6t
Xbit_r120_c72 bl[72] br[72] wl[120] vdd gnd cell_6t
Xbit_r121_c72 bl[72] br[72] wl[121] vdd gnd cell_6t
Xbit_r122_c72 bl[72] br[72] wl[122] vdd gnd cell_6t
Xbit_r123_c72 bl[72] br[72] wl[123] vdd gnd cell_6t
Xbit_r124_c72 bl[72] br[72] wl[124] vdd gnd cell_6t
Xbit_r125_c72 bl[72] br[72] wl[125] vdd gnd cell_6t
Xbit_r126_c72 bl[72] br[72] wl[126] vdd gnd cell_6t
Xbit_r127_c72 bl[72] br[72] wl[127] vdd gnd cell_6t
Xbit_r128_c72 bl[72] br[72] wl[128] vdd gnd cell_6t
Xbit_r129_c72 bl[72] br[72] wl[129] vdd gnd cell_6t
Xbit_r130_c72 bl[72] br[72] wl[130] vdd gnd cell_6t
Xbit_r131_c72 bl[72] br[72] wl[131] vdd gnd cell_6t
Xbit_r132_c72 bl[72] br[72] wl[132] vdd gnd cell_6t
Xbit_r133_c72 bl[72] br[72] wl[133] vdd gnd cell_6t
Xbit_r134_c72 bl[72] br[72] wl[134] vdd gnd cell_6t
Xbit_r135_c72 bl[72] br[72] wl[135] vdd gnd cell_6t
Xbit_r136_c72 bl[72] br[72] wl[136] vdd gnd cell_6t
Xbit_r137_c72 bl[72] br[72] wl[137] vdd gnd cell_6t
Xbit_r138_c72 bl[72] br[72] wl[138] vdd gnd cell_6t
Xbit_r139_c72 bl[72] br[72] wl[139] vdd gnd cell_6t
Xbit_r140_c72 bl[72] br[72] wl[140] vdd gnd cell_6t
Xbit_r141_c72 bl[72] br[72] wl[141] vdd gnd cell_6t
Xbit_r142_c72 bl[72] br[72] wl[142] vdd gnd cell_6t
Xbit_r143_c72 bl[72] br[72] wl[143] vdd gnd cell_6t
Xbit_r144_c72 bl[72] br[72] wl[144] vdd gnd cell_6t
Xbit_r145_c72 bl[72] br[72] wl[145] vdd gnd cell_6t
Xbit_r146_c72 bl[72] br[72] wl[146] vdd gnd cell_6t
Xbit_r147_c72 bl[72] br[72] wl[147] vdd gnd cell_6t
Xbit_r148_c72 bl[72] br[72] wl[148] vdd gnd cell_6t
Xbit_r149_c72 bl[72] br[72] wl[149] vdd gnd cell_6t
Xbit_r150_c72 bl[72] br[72] wl[150] vdd gnd cell_6t
Xbit_r151_c72 bl[72] br[72] wl[151] vdd gnd cell_6t
Xbit_r152_c72 bl[72] br[72] wl[152] vdd gnd cell_6t
Xbit_r153_c72 bl[72] br[72] wl[153] vdd gnd cell_6t
Xbit_r154_c72 bl[72] br[72] wl[154] vdd gnd cell_6t
Xbit_r155_c72 bl[72] br[72] wl[155] vdd gnd cell_6t
Xbit_r156_c72 bl[72] br[72] wl[156] vdd gnd cell_6t
Xbit_r157_c72 bl[72] br[72] wl[157] vdd gnd cell_6t
Xbit_r158_c72 bl[72] br[72] wl[158] vdd gnd cell_6t
Xbit_r159_c72 bl[72] br[72] wl[159] vdd gnd cell_6t
Xbit_r160_c72 bl[72] br[72] wl[160] vdd gnd cell_6t
Xbit_r161_c72 bl[72] br[72] wl[161] vdd gnd cell_6t
Xbit_r162_c72 bl[72] br[72] wl[162] vdd gnd cell_6t
Xbit_r163_c72 bl[72] br[72] wl[163] vdd gnd cell_6t
Xbit_r164_c72 bl[72] br[72] wl[164] vdd gnd cell_6t
Xbit_r165_c72 bl[72] br[72] wl[165] vdd gnd cell_6t
Xbit_r166_c72 bl[72] br[72] wl[166] vdd gnd cell_6t
Xbit_r167_c72 bl[72] br[72] wl[167] vdd gnd cell_6t
Xbit_r168_c72 bl[72] br[72] wl[168] vdd gnd cell_6t
Xbit_r169_c72 bl[72] br[72] wl[169] vdd gnd cell_6t
Xbit_r170_c72 bl[72] br[72] wl[170] vdd gnd cell_6t
Xbit_r171_c72 bl[72] br[72] wl[171] vdd gnd cell_6t
Xbit_r172_c72 bl[72] br[72] wl[172] vdd gnd cell_6t
Xbit_r173_c72 bl[72] br[72] wl[173] vdd gnd cell_6t
Xbit_r174_c72 bl[72] br[72] wl[174] vdd gnd cell_6t
Xbit_r175_c72 bl[72] br[72] wl[175] vdd gnd cell_6t
Xbit_r176_c72 bl[72] br[72] wl[176] vdd gnd cell_6t
Xbit_r177_c72 bl[72] br[72] wl[177] vdd gnd cell_6t
Xbit_r178_c72 bl[72] br[72] wl[178] vdd gnd cell_6t
Xbit_r179_c72 bl[72] br[72] wl[179] vdd gnd cell_6t
Xbit_r180_c72 bl[72] br[72] wl[180] vdd gnd cell_6t
Xbit_r181_c72 bl[72] br[72] wl[181] vdd gnd cell_6t
Xbit_r182_c72 bl[72] br[72] wl[182] vdd gnd cell_6t
Xbit_r183_c72 bl[72] br[72] wl[183] vdd gnd cell_6t
Xbit_r184_c72 bl[72] br[72] wl[184] vdd gnd cell_6t
Xbit_r185_c72 bl[72] br[72] wl[185] vdd gnd cell_6t
Xbit_r186_c72 bl[72] br[72] wl[186] vdd gnd cell_6t
Xbit_r187_c72 bl[72] br[72] wl[187] vdd gnd cell_6t
Xbit_r188_c72 bl[72] br[72] wl[188] vdd gnd cell_6t
Xbit_r189_c72 bl[72] br[72] wl[189] vdd gnd cell_6t
Xbit_r190_c72 bl[72] br[72] wl[190] vdd gnd cell_6t
Xbit_r191_c72 bl[72] br[72] wl[191] vdd gnd cell_6t
Xbit_r192_c72 bl[72] br[72] wl[192] vdd gnd cell_6t
Xbit_r193_c72 bl[72] br[72] wl[193] vdd gnd cell_6t
Xbit_r194_c72 bl[72] br[72] wl[194] vdd gnd cell_6t
Xbit_r195_c72 bl[72] br[72] wl[195] vdd gnd cell_6t
Xbit_r196_c72 bl[72] br[72] wl[196] vdd gnd cell_6t
Xbit_r197_c72 bl[72] br[72] wl[197] vdd gnd cell_6t
Xbit_r198_c72 bl[72] br[72] wl[198] vdd gnd cell_6t
Xbit_r199_c72 bl[72] br[72] wl[199] vdd gnd cell_6t
Xbit_r200_c72 bl[72] br[72] wl[200] vdd gnd cell_6t
Xbit_r201_c72 bl[72] br[72] wl[201] vdd gnd cell_6t
Xbit_r202_c72 bl[72] br[72] wl[202] vdd gnd cell_6t
Xbit_r203_c72 bl[72] br[72] wl[203] vdd gnd cell_6t
Xbit_r204_c72 bl[72] br[72] wl[204] vdd gnd cell_6t
Xbit_r205_c72 bl[72] br[72] wl[205] vdd gnd cell_6t
Xbit_r206_c72 bl[72] br[72] wl[206] vdd gnd cell_6t
Xbit_r207_c72 bl[72] br[72] wl[207] vdd gnd cell_6t
Xbit_r208_c72 bl[72] br[72] wl[208] vdd gnd cell_6t
Xbit_r209_c72 bl[72] br[72] wl[209] vdd gnd cell_6t
Xbit_r210_c72 bl[72] br[72] wl[210] vdd gnd cell_6t
Xbit_r211_c72 bl[72] br[72] wl[211] vdd gnd cell_6t
Xbit_r212_c72 bl[72] br[72] wl[212] vdd gnd cell_6t
Xbit_r213_c72 bl[72] br[72] wl[213] vdd gnd cell_6t
Xbit_r214_c72 bl[72] br[72] wl[214] vdd gnd cell_6t
Xbit_r215_c72 bl[72] br[72] wl[215] vdd gnd cell_6t
Xbit_r216_c72 bl[72] br[72] wl[216] vdd gnd cell_6t
Xbit_r217_c72 bl[72] br[72] wl[217] vdd gnd cell_6t
Xbit_r218_c72 bl[72] br[72] wl[218] vdd gnd cell_6t
Xbit_r219_c72 bl[72] br[72] wl[219] vdd gnd cell_6t
Xbit_r220_c72 bl[72] br[72] wl[220] vdd gnd cell_6t
Xbit_r221_c72 bl[72] br[72] wl[221] vdd gnd cell_6t
Xbit_r222_c72 bl[72] br[72] wl[222] vdd gnd cell_6t
Xbit_r223_c72 bl[72] br[72] wl[223] vdd gnd cell_6t
Xbit_r224_c72 bl[72] br[72] wl[224] vdd gnd cell_6t
Xbit_r225_c72 bl[72] br[72] wl[225] vdd gnd cell_6t
Xbit_r226_c72 bl[72] br[72] wl[226] vdd gnd cell_6t
Xbit_r227_c72 bl[72] br[72] wl[227] vdd gnd cell_6t
Xbit_r228_c72 bl[72] br[72] wl[228] vdd gnd cell_6t
Xbit_r229_c72 bl[72] br[72] wl[229] vdd gnd cell_6t
Xbit_r230_c72 bl[72] br[72] wl[230] vdd gnd cell_6t
Xbit_r231_c72 bl[72] br[72] wl[231] vdd gnd cell_6t
Xbit_r232_c72 bl[72] br[72] wl[232] vdd gnd cell_6t
Xbit_r233_c72 bl[72] br[72] wl[233] vdd gnd cell_6t
Xbit_r234_c72 bl[72] br[72] wl[234] vdd gnd cell_6t
Xbit_r235_c72 bl[72] br[72] wl[235] vdd gnd cell_6t
Xbit_r236_c72 bl[72] br[72] wl[236] vdd gnd cell_6t
Xbit_r237_c72 bl[72] br[72] wl[237] vdd gnd cell_6t
Xbit_r238_c72 bl[72] br[72] wl[238] vdd gnd cell_6t
Xbit_r239_c72 bl[72] br[72] wl[239] vdd gnd cell_6t
Xbit_r240_c72 bl[72] br[72] wl[240] vdd gnd cell_6t
Xbit_r241_c72 bl[72] br[72] wl[241] vdd gnd cell_6t
Xbit_r242_c72 bl[72] br[72] wl[242] vdd gnd cell_6t
Xbit_r243_c72 bl[72] br[72] wl[243] vdd gnd cell_6t
Xbit_r244_c72 bl[72] br[72] wl[244] vdd gnd cell_6t
Xbit_r245_c72 bl[72] br[72] wl[245] vdd gnd cell_6t
Xbit_r246_c72 bl[72] br[72] wl[246] vdd gnd cell_6t
Xbit_r247_c72 bl[72] br[72] wl[247] vdd gnd cell_6t
Xbit_r248_c72 bl[72] br[72] wl[248] vdd gnd cell_6t
Xbit_r249_c72 bl[72] br[72] wl[249] vdd gnd cell_6t
Xbit_r250_c72 bl[72] br[72] wl[250] vdd gnd cell_6t
Xbit_r251_c72 bl[72] br[72] wl[251] vdd gnd cell_6t
Xbit_r252_c72 bl[72] br[72] wl[252] vdd gnd cell_6t
Xbit_r253_c72 bl[72] br[72] wl[253] vdd gnd cell_6t
Xbit_r254_c72 bl[72] br[72] wl[254] vdd gnd cell_6t
Xbit_r255_c72 bl[72] br[72] wl[255] vdd gnd cell_6t
Xbit_r256_c72 bl[72] br[72] wl[256] vdd gnd cell_6t
Xbit_r257_c72 bl[72] br[72] wl[257] vdd gnd cell_6t
Xbit_r258_c72 bl[72] br[72] wl[258] vdd gnd cell_6t
Xbit_r259_c72 bl[72] br[72] wl[259] vdd gnd cell_6t
Xbit_r260_c72 bl[72] br[72] wl[260] vdd gnd cell_6t
Xbit_r261_c72 bl[72] br[72] wl[261] vdd gnd cell_6t
Xbit_r262_c72 bl[72] br[72] wl[262] vdd gnd cell_6t
Xbit_r263_c72 bl[72] br[72] wl[263] vdd gnd cell_6t
Xbit_r264_c72 bl[72] br[72] wl[264] vdd gnd cell_6t
Xbit_r265_c72 bl[72] br[72] wl[265] vdd gnd cell_6t
Xbit_r266_c72 bl[72] br[72] wl[266] vdd gnd cell_6t
Xbit_r267_c72 bl[72] br[72] wl[267] vdd gnd cell_6t
Xbit_r268_c72 bl[72] br[72] wl[268] vdd gnd cell_6t
Xbit_r269_c72 bl[72] br[72] wl[269] vdd gnd cell_6t
Xbit_r270_c72 bl[72] br[72] wl[270] vdd gnd cell_6t
Xbit_r271_c72 bl[72] br[72] wl[271] vdd gnd cell_6t
Xbit_r272_c72 bl[72] br[72] wl[272] vdd gnd cell_6t
Xbit_r273_c72 bl[72] br[72] wl[273] vdd gnd cell_6t
Xbit_r274_c72 bl[72] br[72] wl[274] vdd gnd cell_6t
Xbit_r275_c72 bl[72] br[72] wl[275] vdd gnd cell_6t
Xbit_r276_c72 bl[72] br[72] wl[276] vdd gnd cell_6t
Xbit_r277_c72 bl[72] br[72] wl[277] vdd gnd cell_6t
Xbit_r278_c72 bl[72] br[72] wl[278] vdd gnd cell_6t
Xbit_r279_c72 bl[72] br[72] wl[279] vdd gnd cell_6t
Xbit_r280_c72 bl[72] br[72] wl[280] vdd gnd cell_6t
Xbit_r281_c72 bl[72] br[72] wl[281] vdd gnd cell_6t
Xbit_r282_c72 bl[72] br[72] wl[282] vdd gnd cell_6t
Xbit_r283_c72 bl[72] br[72] wl[283] vdd gnd cell_6t
Xbit_r284_c72 bl[72] br[72] wl[284] vdd gnd cell_6t
Xbit_r285_c72 bl[72] br[72] wl[285] vdd gnd cell_6t
Xbit_r286_c72 bl[72] br[72] wl[286] vdd gnd cell_6t
Xbit_r287_c72 bl[72] br[72] wl[287] vdd gnd cell_6t
Xbit_r288_c72 bl[72] br[72] wl[288] vdd gnd cell_6t
Xbit_r289_c72 bl[72] br[72] wl[289] vdd gnd cell_6t
Xbit_r290_c72 bl[72] br[72] wl[290] vdd gnd cell_6t
Xbit_r291_c72 bl[72] br[72] wl[291] vdd gnd cell_6t
Xbit_r292_c72 bl[72] br[72] wl[292] vdd gnd cell_6t
Xbit_r293_c72 bl[72] br[72] wl[293] vdd gnd cell_6t
Xbit_r294_c72 bl[72] br[72] wl[294] vdd gnd cell_6t
Xbit_r295_c72 bl[72] br[72] wl[295] vdd gnd cell_6t
Xbit_r296_c72 bl[72] br[72] wl[296] vdd gnd cell_6t
Xbit_r297_c72 bl[72] br[72] wl[297] vdd gnd cell_6t
Xbit_r298_c72 bl[72] br[72] wl[298] vdd gnd cell_6t
Xbit_r299_c72 bl[72] br[72] wl[299] vdd gnd cell_6t
Xbit_r300_c72 bl[72] br[72] wl[300] vdd gnd cell_6t
Xbit_r301_c72 bl[72] br[72] wl[301] vdd gnd cell_6t
Xbit_r302_c72 bl[72] br[72] wl[302] vdd gnd cell_6t
Xbit_r303_c72 bl[72] br[72] wl[303] vdd gnd cell_6t
Xbit_r304_c72 bl[72] br[72] wl[304] vdd gnd cell_6t
Xbit_r305_c72 bl[72] br[72] wl[305] vdd gnd cell_6t
Xbit_r306_c72 bl[72] br[72] wl[306] vdd gnd cell_6t
Xbit_r307_c72 bl[72] br[72] wl[307] vdd gnd cell_6t
Xbit_r308_c72 bl[72] br[72] wl[308] vdd gnd cell_6t
Xbit_r309_c72 bl[72] br[72] wl[309] vdd gnd cell_6t
Xbit_r310_c72 bl[72] br[72] wl[310] vdd gnd cell_6t
Xbit_r311_c72 bl[72] br[72] wl[311] vdd gnd cell_6t
Xbit_r312_c72 bl[72] br[72] wl[312] vdd gnd cell_6t
Xbit_r313_c72 bl[72] br[72] wl[313] vdd gnd cell_6t
Xbit_r314_c72 bl[72] br[72] wl[314] vdd gnd cell_6t
Xbit_r315_c72 bl[72] br[72] wl[315] vdd gnd cell_6t
Xbit_r316_c72 bl[72] br[72] wl[316] vdd gnd cell_6t
Xbit_r317_c72 bl[72] br[72] wl[317] vdd gnd cell_6t
Xbit_r318_c72 bl[72] br[72] wl[318] vdd gnd cell_6t
Xbit_r319_c72 bl[72] br[72] wl[319] vdd gnd cell_6t
Xbit_r320_c72 bl[72] br[72] wl[320] vdd gnd cell_6t
Xbit_r321_c72 bl[72] br[72] wl[321] vdd gnd cell_6t
Xbit_r322_c72 bl[72] br[72] wl[322] vdd gnd cell_6t
Xbit_r323_c72 bl[72] br[72] wl[323] vdd gnd cell_6t
Xbit_r324_c72 bl[72] br[72] wl[324] vdd gnd cell_6t
Xbit_r325_c72 bl[72] br[72] wl[325] vdd gnd cell_6t
Xbit_r326_c72 bl[72] br[72] wl[326] vdd gnd cell_6t
Xbit_r327_c72 bl[72] br[72] wl[327] vdd gnd cell_6t
Xbit_r328_c72 bl[72] br[72] wl[328] vdd gnd cell_6t
Xbit_r329_c72 bl[72] br[72] wl[329] vdd gnd cell_6t
Xbit_r330_c72 bl[72] br[72] wl[330] vdd gnd cell_6t
Xbit_r331_c72 bl[72] br[72] wl[331] vdd gnd cell_6t
Xbit_r332_c72 bl[72] br[72] wl[332] vdd gnd cell_6t
Xbit_r333_c72 bl[72] br[72] wl[333] vdd gnd cell_6t
Xbit_r334_c72 bl[72] br[72] wl[334] vdd gnd cell_6t
Xbit_r335_c72 bl[72] br[72] wl[335] vdd gnd cell_6t
Xbit_r336_c72 bl[72] br[72] wl[336] vdd gnd cell_6t
Xbit_r337_c72 bl[72] br[72] wl[337] vdd gnd cell_6t
Xbit_r338_c72 bl[72] br[72] wl[338] vdd gnd cell_6t
Xbit_r339_c72 bl[72] br[72] wl[339] vdd gnd cell_6t
Xbit_r340_c72 bl[72] br[72] wl[340] vdd gnd cell_6t
Xbit_r341_c72 bl[72] br[72] wl[341] vdd gnd cell_6t
Xbit_r342_c72 bl[72] br[72] wl[342] vdd gnd cell_6t
Xbit_r343_c72 bl[72] br[72] wl[343] vdd gnd cell_6t
Xbit_r344_c72 bl[72] br[72] wl[344] vdd gnd cell_6t
Xbit_r345_c72 bl[72] br[72] wl[345] vdd gnd cell_6t
Xbit_r346_c72 bl[72] br[72] wl[346] vdd gnd cell_6t
Xbit_r347_c72 bl[72] br[72] wl[347] vdd gnd cell_6t
Xbit_r348_c72 bl[72] br[72] wl[348] vdd gnd cell_6t
Xbit_r349_c72 bl[72] br[72] wl[349] vdd gnd cell_6t
Xbit_r350_c72 bl[72] br[72] wl[350] vdd gnd cell_6t
Xbit_r351_c72 bl[72] br[72] wl[351] vdd gnd cell_6t
Xbit_r352_c72 bl[72] br[72] wl[352] vdd gnd cell_6t
Xbit_r353_c72 bl[72] br[72] wl[353] vdd gnd cell_6t
Xbit_r354_c72 bl[72] br[72] wl[354] vdd gnd cell_6t
Xbit_r355_c72 bl[72] br[72] wl[355] vdd gnd cell_6t
Xbit_r356_c72 bl[72] br[72] wl[356] vdd gnd cell_6t
Xbit_r357_c72 bl[72] br[72] wl[357] vdd gnd cell_6t
Xbit_r358_c72 bl[72] br[72] wl[358] vdd gnd cell_6t
Xbit_r359_c72 bl[72] br[72] wl[359] vdd gnd cell_6t
Xbit_r360_c72 bl[72] br[72] wl[360] vdd gnd cell_6t
Xbit_r361_c72 bl[72] br[72] wl[361] vdd gnd cell_6t
Xbit_r362_c72 bl[72] br[72] wl[362] vdd gnd cell_6t
Xbit_r363_c72 bl[72] br[72] wl[363] vdd gnd cell_6t
Xbit_r364_c72 bl[72] br[72] wl[364] vdd gnd cell_6t
Xbit_r365_c72 bl[72] br[72] wl[365] vdd gnd cell_6t
Xbit_r366_c72 bl[72] br[72] wl[366] vdd gnd cell_6t
Xbit_r367_c72 bl[72] br[72] wl[367] vdd gnd cell_6t
Xbit_r368_c72 bl[72] br[72] wl[368] vdd gnd cell_6t
Xbit_r369_c72 bl[72] br[72] wl[369] vdd gnd cell_6t
Xbit_r370_c72 bl[72] br[72] wl[370] vdd gnd cell_6t
Xbit_r371_c72 bl[72] br[72] wl[371] vdd gnd cell_6t
Xbit_r372_c72 bl[72] br[72] wl[372] vdd gnd cell_6t
Xbit_r373_c72 bl[72] br[72] wl[373] vdd gnd cell_6t
Xbit_r374_c72 bl[72] br[72] wl[374] vdd gnd cell_6t
Xbit_r375_c72 bl[72] br[72] wl[375] vdd gnd cell_6t
Xbit_r376_c72 bl[72] br[72] wl[376] vdd gnd cell_6t
Xbit_r377_c72 bl[72] br[72] wl[377] vdd gnd cell_6t
Xbit_r378_c72 bl[72] br[72] wl[378] vdd gnd cell_6t
Xbit_r379_c72 bl[72] br[72] wl[379] vdd gnd cell_6t
Xbit_r380_c72 bl[72] br[72] wl[380] vdd gnd cell_6t
Xbit_r381_c72 bl[72] br[72] wl[381] vdd gnd cell_6t
Xbit_r382_c72 bl[72] br[72] wl[382] vdd gnd cell_6t
Xbit_r383_c72 bl[72] br[72] wl[383] vdd gnd cell_6t
Xbit_r384_c72 bl[72] br[72] wl[384] vdd gnd cell_6t
Xbit_r385_c72 bl[72] br[72] wl[385] vdd gnd cell_6t
Xbit_r386_c72 bl[72] br[72] wl[386] vdd gnd cell_6t
Xbit_r387_c72 bl[72] br[72] wl[387] vdd gnd cell_6t
Xbit_r388_c72 bl[72] br[72] wl[388] vdd gnd cell_6t
Xbit_r389_c72 bl[72] br[72] wl[389] vdd gnd cell_6t
Xbit_r390_c72 bl[72] br[72] wl[390] vdd gnd cell_6t
Xbit_r391_c72 bl[72] br[72] wl[391] vdd gnd cell_6t
Xbit_r392_c72 bl[72] br[72] wl[392] vdd gnd cell_6t
Xbit_r393_c72 bl[72] br[72] wl[393] vdd gnd cell_6t
Xbit_r394_c72 bl[72] br[72] wl[394] vdd gnd cell_6t
Xbit_r395_c72 bl[72] br[72] wl[395] vdd gnd cell_6t
Xbit_r396_c72 bl[72] br[72] wl[396] vdd gnd cell_6t
Xbit_r397_c72 bl[72] br[72] wl[397] vdd gnd cell_6t
Xbit_r398_c72 bl[72] br[72] wl[398] vdd gnd cell_6t
Xbit_r399_c72 bl[72] br[72] wl[399] vdd gnd cell_6t
Xbit_r400_c72 bl[72] br[72] wl[400] vdd gnd cell_6t
Xbit_r401_c72 bl[72] br[72] wl[401] vdd gnd cell_6t
Xbit_r402_c72 bl[72] br[72] wl[402] vdd gnd cell_6t
Xbit_r403_c72 bl[72] br[72] wl[403] vdd gnd cell_6t
Xbit_r404_c72 bl[72] br[72] wl[404] vdd gnd cell_6t
Xbit_r405_c72 bl[72] br[72] wl[405] vdd gnd cell_6t
Xbit_r406_c72 bl[72] br[72] wl[406] vdd gnd cell_6t
Xbit_r407_c72 bl[72] br[72] wl[407] vdd gnd cell_6t
Xbit_r408_c72 bl[72] br[72] wl[408] vdd gnd cell_6t
Xbit_r409_c72 bl[72] br[72] wl[409] vdd gnd cell_6t
Xbit_r410_c72 bl[72] br[72] wl[410] vdd gnd cell_6t
Xbit_r411_c72 bl[72] br[72] wl[411] vdd gnd cell_6t
Xbit_r412_c72 bl[72] br[72] wl[412] vdd gnd cell_6t
Xbit_r413_c72 bl[72] br[72] wl[413] vdd gnd cell_6t
Xbit_r414_c72 bl[72] br[72] wl[414] vdd gnd cell_6t
Xbit_r415_c72 bl[72] br[72] wl[415] vdd gnd cell_6t
Xbit_r416_c72 bl[72] br[72] wl[416] vdd gnd cell_6t
Xbit_r417_c72 bl[72] br[72] wl[417] vdd gnd cell_6t
Xbit_r418_c72 bl[72] br[72] wl[418] vdd gnd cell_6t
Xbit_r419_c72 bl[72] br[72] wl[419] vdd gnd cell_6t
Xbit_r420_c72 bl[72] br[72] wl[420] vdd gnd cell_6t
Xbit_r421_c72 bl[72] br[72] wl[421] vdd gnd cell_6t
Xbit_r422_c72 bl[72] br[72] wl[422] vdd gnd cell_6t
Xbit_r423_c72 bl[72] br[72] wl[423] vdd gnd cell_6t
Xbit_r424_c72 bl[72] br[72] wl[424] vdd gnd cell_6t
Xbit_r425_c72 bl[72] br[72] wl[425] vdd gnd cell_6t
Xbit_r426_c72 bl[72] br[72] wl[426] vdd gnd cell_6t
Xbit_r427_c72 bl[72] br[72] wl[427] vdd gnd cell_6t
Xbit_r428_c72 bl[72] br[72] wl[428] vdd gnd cell_6t
Xbit_r429_c72 bl[72] br[72] wl[429] vdd gnd cell_6t
Xbit_r430_c72 bl[72] br[72] wl[430] vdd gnd cell_6t
Xbit_r431_c72 bl[72] br[72] wl[431] vdd gnd cell_6t
Xbit_r432_c72 bl[72] br[72] wl[432] vdd gnd cell_6t
Xbit_r433_c72 bl[72] br[72] wl[433] vdd gnd cell_6t
Xbit_r434_c72 bl[72] br[72] wl[434] vdd gnd cell_6t
Xbit_r435_c72 bl[72] br[72] wl[435] vdd gnd cell_6t
Xbit_r436_c72 bl[72] br[72] wl[436] vdd gnd cell_6t
Xbit_r437_c72 bl[72] br[72] wl[437] vdd gnd cell_6t
Xbit_r438_c72 bl[72] br[72] wl[438] vdd gnd cell_6t
Xbit_r439_c72 bl[72] br[72] wl[439] vdd gnd cell_6t
Xbit_r440_c72 bl[72] br[72] wl[440] vdd gnd cell_6t
Xbit_r441_c72 bl[72] br[72] wl[441] vdd gnd cell_6t
Xbit_r442_c72 bl[72] br[72] wl[442] vdd gnd cell_6t
Xbit_r443_c72 bl[72] br[72] wl[443] vdd gnd cell_6t
Xbit_r444_c72 bl[72] br[72] wl[444] vdd gnd cell_6t
Xbit_r445_c72 bl[72] br[72] wl[445] vdd gnd cell_6t
Xbit_r446_c72 bl[72] br[72] wl[446] vdd gnd cell_6t
Xbit_r447_c72 bl[72] br[72] wl[447] vdd gnd cell_6t
Xbit_r448_c72 bl[72] br[72] wl[448] vdd gnd cell_6t
Xbit_r449_c72 bl[72] br[72] wl[449] vdd gnd cell_6t
Xbit_r450_c72 bl[72] br[72] wl[450] vdd gnd cell_6t
Xbit_r451_c72 bl[72] br[72] wl[451] vdd gnd cell_6t
Xbit_r452_c72 bl[72] br[72] wl[452] vdd gnd cell_6t
Xbit_r453_c72 bl[72] br[72] wl[453] vdd gnd cell_6t
Xbit_r454_c72 bl[72] br[72] wl[454] vdd gnd cell_6t
Xbit_r455_c72 bl[72] br[72] wl[455] vdd gnd cell_6t
Xbit_r456_c72 bl[72] br[72] wl[456] vdd gnd cell_6t
Xbit_r457_c72 bl[72] br[72] wl[457] vdd gnd cell_6t
Xbit_r458_c72 bl[72] br[72] wl[458] vdd gnd cell_6t
Xbit_r459_c72 bl[72] br[72] wl[459] vdd gnd cell_6t
Xbit_r460_c72 bl[72] br[72] wl[460] vdd gnd cell_6t
Xbit_r461_c72 bl[72] br[72] wl[461] vdd gnd cell_6t
Xbit_r462_c72 bl[72] br[72] wl[462] vdd gnd cell_6t
Xbit_r463_c72 bl[72] br[72] wl[463] vdd gnd cell_6t
Xbit_r464_c72 bl[72] br[72] wl[464] vdd gnd cell_6t
Xbit_r465_c72 bl[72] br[72] wl[465] vdd gnd cell_6t
Xbit_r466_c72 bl[72] br[72] wl[466] vdd gnd cell_6t
Xbit_r467_c72 bl[72] br[72] wl[467] vdd gnd cell_6t
Xbit_r468_c72 bl[72] br[72] wl[468] vdd gnd cell_6t
Xbit_r469_c72 bl[72] br[72] wl[469] vdd gnd cell_6t
Xbit_r470_c72 bl[72] br[72] wl[470] vdd gnd cell_6t
Xbit_r471_c72 bl[72] br[72] wl[471] vdd gnd cell_6t
Xbit_r472_c72 bl[72] br[72] wl[472] vdd gnd cell_6t
Xbit_r473_c72 bl[72] br[72] wl[473] vdd gnd cell_6t
Xbit_r474_c72 bl[72] br[72] wl[474] vdd gnd cell_6t
Xbit_r475_c72 bl[72] br[72] wl[475] vdd gnd cell_6t
Xbit_r476_c72 bl[72] br[72] wl[476] vdd gnd cell_6t
Xbit_r477_c72 bl[72] br[72] wl[477] vdd gnd cell_6t
Xbit_r478_c72 bl[72] br[72] wl[478] vdd gnd cell_6t
Xbit_r479_c72 bl[72] br[72] wl[479] vdd gnd cell_6t
Xbit_r480_c72 bl[72] br[72] wl[480] vdd gnd cell_6t
Xbit_r481_c72 bl[72] br[72] wl[481] vdd gnd cell_6t
Xbit_r482_c72 bl[72] br[72] wl[482] vdd gnd cell_6t
Xbit_r483_c72 bl[72] br[72] wl[483] vdd gnd cell_6t
Xbit_r484_c72 bl[72] br[72] wl[484] vdd gnd cell_6t
Xbit_r485_c72 bl[72] br[72] wl[485] vdd gnd cell_6t
Xbit_r486_c72 bl[72] br[72] wl[486] vdd gnd cell_6t
Xbit_r487_c72 bl[72] br[72] wl[487] vdd gnd cell_6t
Xbit_r488_c72 bl[72] br[72] wl[488] vdd gnd cell_6t
Xbit_r489_c72 bl[72] br[72] wl[489] vdd gnd cell_6t
Xbit_r490_c72 bl[72] br[72] wl[490] vdd gnd cell_6t
Xbit_r491_c72 bl[72] br[72] wl[491] vdd gnd cell_6t
Xbit_r492_c72 bl[72] br[72] wl[492] vdd gnd cell_6t
Xbit_r493_c72 bl[72] br[72] wl[493] vdd gnd cell_6t
Xbit_r494_c72 bl[72] br[72] wl[494] vdd gnd cell_6t
Xbit_r495_c72 bl[72] br[72] wl[495] vdd gnd cell_6t
Xbit_r496_c72 bl[72] br[72] wl[496] vdd gnd cell_6t
Xbit_r497_c72 bl[72] br[72] wl[497] vdd gnd cell_6t
Xbit_r498_c72 bl[72] br[72] wl[498] vdd gnd cell_6t
Xbit_r499_c72 bl[72] br[72] wl[499] vdd gnd cell_6t
Xbit_r500_c72 bl[72] br[72] wl[500] vdd gnd cell_6t
Xbit_r501_c72 bl[72] br[72] wl[501] vdd gnd cell_6t
Xbit_r502_c72 bl[72] br[72] wl[502] vdd gnd cell_6t
Xbit_r503_c72 bl[72] br[72] wl[503] vdd gnd cell_6t
Xbit_r504_c72 bl[72] br[72] wl[504] vdd gnd cell_6t
Xbit_r505_c72 bl[72] br[72] wl[505] vdd gnd cell_6t
Xbit_r506_c72 bl[72] br[72] wl[506] vdd gnd cell_6t
Xbit_r507_c72 bl[72] br[72] wl[507] vdd gnd cell_6t
Xbit_r508_c72 bl[72] br[72] wl[508] vdd gnd cell_6t
Xbit_r509_c72 bl[72] br[72] wl[509] vdd gnd cell_6t
Xbit_r510_c72 bl[72] br[72] wl[510] vdd gnd cell_6t
Xbit_r511_c72 bl[72] br[72] wl[511] vdd gnd cell_6t
Xbit_r0_c73 bl[73] br[73] wl[0] vdd gnd cell_6t
Xbit_r1_c73 bl[73] br[73] wl[1] vdd gnd cell_6t
Xbit_r2_c73 bl[73] br[73] wl[2] vdd gnd cell_6t
Xbit_r3_c73 bl[73] br[73] wl[3] vdd gnd cell_6t
Xbit_r4_c73 bl[73] br[73] wl[4] vdd gnd cell_6t
Xbit_r5_c73 bl[73] br[73] wl[5] vdd gnd cell_6t
Xbit_r6_c73 bl[73] br[73] wl[6] vdd gnd cell_6t
Xbit_r7_c73 bl[73] br[73] wl[7] vdd gnd cell_6t
Xbit_r8_c73 bl[73] br[73] wl[8] vdd gnd cell_6t
Xbit_r9_c73 bl[73] br[73] wl[9] vdd gnd cell_6t
Xbit_r10_c73 bl[73] br[73] wl[10] vdd gnd cell_6t
Xbit_r11_c73 bl[73] br[73] wl[11] vdd gnd cell_6t
Xbit_r12_c73 bl[73] br[73] wl[12] vdd gnd cell_6t
Xbit_r13_c73 bl[73] br[73] wl[13] vdd gnd cell_6t
Xbit_r14_c73 bl[73] br[73] wl[14] vdd gnd cell_6t
Xbit_r15_c73 bl[73] br[73] wl[15] vdd gnd cell_6t
Xbit_r16_c73 bl[73] br[73] wl[16] vdd gnd cell_6t
Xbit_r17_c73 bl[73] br[73] wl[17] vdd gnd cell_6t
Xbit_r18_c73 bl[73] br[73] wl[18] vdd gnd cell_6t
Xbit_r19_c73 bl[73] br[73] wl[19] vdd gnd cell_6t
Xbit_r20_c73 bl[73] br[73] wl[20] vdd gnd cell_6t
Xbit_r21_c73 bl[73] br[73] wl[21] vdd gnd cell_6t
Xbit_r22_c73 bl[73] br[73] wl[22] vdd gnd cell_6t
Xbit_r23_c73 bl[73] br[73] wl[23] vdd gnd cell_6t
Xbit_r24_c73 bl[73] br[73] wl[24] vdd gnd cell_6t
Xbit_r25_c73 bl[73] br[73] wl[25] vdd gnd cell_6t
Xbit_r26_c73 bl[73] br[73] wl[26] vdd gnd cell_6t
Xbit_r27_c73 bl[73] br[73] wl[27] vdd gnd cell_6t
Xbit_r28_c73 bl[73] br[73] wl[28] vdd gnd cell_6t
Xbit_r29_c73 bl[73] br[73] wl[29] vdd gnd cell_6t
Xbit_r30_c73 bl[73] br[73] wl[30] vdd gnd cell_6t
Xbit_r31_c73 bl[73] br[73] wl[31] vdd gnd cell_6t
Xbit_r32_c73 bl[73] br[73] wl[32] vdd gnd cell_6t
Xbit_r33_c73 bl[73] br[73] wl[33] vdd gnd cell_6t
Xbit_r34_c73 bl[73] br[73] wl[34] vdd gnd cell_6t
Xbit_r35_c73 bl[73] br[73] wl[35] vdd gnd cell_6t
Xbit_r36_c73 bl[73] br[73] wl[36] vdd gnd cell_6t
Xbit_r37_c73 bl[73] br[73] wl[37] vdd gnd cell_6t
Xbit_r38_c73 bl[73] br[73] wl[38] vdd gnd cell_6t
Xbit_r39_c73 bl[73] br[73] wl[39] vdd gnd cell_6t
Xbit_r40_c73 bl[73] br[73] wl[40] vdd gnd cell_6t
Xbit_r41_c73 bl[73] br[73] wl[41] vdd gnd cell_6t
Xbit_r42_c73 bl[73] br[73] wl[42] vdd gnd cell_6t
Xbit_r43_c73 bl[73] br[73] wl[43] vdd gnd cell_6t
Xbit_r44_c73 bl[73] br[73] wl[44] vdd gnd cell_6t
Xbit_r45_c73 bl[73] br[73] wl[45] vdd gnd cell_6t
Xbit_r46_c73 bl[73] br[73] wl[46] vdd gnd cell_6t
Xbit_r47_c73 bl[73] br[73] wl[47] vdd gnd cell_6t
Xbit_r48_c73 bl[73] br[73] wl[48] vdd gnd cell_6t
Xbit_r49_c73 bl[73] br[73] wl[49] vdd gnd cell_6t
Xbit_r50_c73 bl[73] br[73] wl[50] vdd gnd cell_6t
Xbit_r51_c73 bl[73] br[73] wl[51] vdd gnd cell_6t
Xbit_r52_c73 bl[73] br[73] wl[52] vdd gnd cell_6t
Xbit_r53_c73 bl[73] br[73] wl[53] vdd gnd cell_6t
Xbit_r54_c73 bl[73] br[73] wl[54] vdd gnd cell_6t
Xbit_r55_c73 bl[73] br[73] wl[55] vdd gnd cell_6t
Xbit_r56_c73 bl[73] br[73] wl[56] vdd gnd cell_6t
Xbit_r57_c73 bl[73] br[73] wl[57] vdd gnd cell_6t
Xbit_r58_c73 bl[73] br[73] wl[58] vdd gnd cell_6t
Xbit_r59_c73 bl[73] br[73] wl[59] vdd gnd cell_6t
Xbit_r60_c73 bl[73] br[73] wl[60] vdd gnd cell_6t
Xbit_r61_c73 bl[73] br[73] wl[61] vdd gnd cell_6t
Xbit_r62_c73 bl[73] br[73] wl[62] vdd gnd cell_6t
Xbit_r63_c73 bl[73] br[73] wl[63] vdd gnd cell_6t
Xbit_r64_c73 bl[73] br[73] wl[64] vdd gnd cell_6t
Xbit_r65_c73 bl[73] br[73] wl[65] vdd gnd cell_6t
Xbit_r66_c73 bl[73] br[73] wl[66] vdd gnd cell_6t
Xbit_r67_c73 bl[73] br[73] wl[67] vdd gnd cell_6t
Xbit_r68_c73 bl[73] br[73] wl[68] vdd gnd cell_6t
Xbit_r69_c73 bl[73] br[73] wl[69] vdd gnd cell_6t
Xbit_r70_c73 bl[73] br[73] wl[70] vdd gnd cell_6t
Xbit_r71_c73 bl[73] br[73] wl[71] vdd gnd cell_6t
Xbit_r72_c73 bl[73] br[73] wl[72] vdd gnd cell_6t
Xbit_r73_c73 bl[73] br[73] wl[73] vdd gnd cell_6t
Xbit_r74_c73 bl[73] br[73] wl[74] vdd gnd cell_6t
Xbit_r75_c73 bl[73] br[73] wl[75] vdd gnd cell_6t
Xbit_r76_c73 bl[73] br[73] wl[76] vdd gnd cell_6t
Xbit_r77_c73 bl[73] br[73] wl[77] vdd gnd cell_6t
Xbit_r78_c73 bl[73] br[73] wl[78] vdd gnd cell_6t
Xbit_r79_c73 bl[73] br[73] wl[79] vdd gnd cell_6t
Xbit_r80_c73 bl[73] br[73] wl[80] vdd gnd cell_6t
Xbit_r81_c73 bl[73] br[73] wl[81] vdd gnd cell_6t
Xbit_r82_c73 bl[73] br[73] wl[82] vdd gnd cell_6t
Xbit_r83_c73 bl[73] br[73] wl[83] vdd gnd cell_6t
Xbit_r84_c73 bl[73] br[73] wl[84] vdd gnd cell_6t
Xbit_r85_c73 bl[73] br[73] wl[85] vdd gnd cell_6t
Xbit_r86_c73 bl[73] br[73] wl[86] vdd gnd cell_6t
Xbit_r87_c73 bl[73] br[73] wl[87] vdd gnd cell_6t
Xbit_r88_c73 bl[73] br[73] wl[88] vdd gnd cell_6t
Xbit_r89_c73 bl[73] br[73] wl[89] vdd gnd cell_6t
Xbit_r90_c73 bl[73] br[73] wl[90] vdd gnd cell_6t
Xbit_r91_c73 bl[73] br[73] wl[91] vdd gnd cell_6t
Xbit_r92_c73 bl[73] br[73] wl[92] vdd gnd cell_6t
Xbit_r93_c73 bl[73] br[73] wl[93] vdd gnd cell_6t
Xbit_r94_c73 bl[73] br[73] wl[94] vdd gnd cell_6t
Xbit_r95_c73 bl[73] br[73] wl[95] vdd gnd cell_6t
Xbit_r96_c73 bl[73] br[73] wl[96] vdd gnd cell_6t
Xbit_r97_c73 bl[73] br[73] wl[97] vdd gnd cell_6t
Xbit_r98_c73 bl[73] br[73] wl[98] vdd gnd cell_6t
Xbit_r99_c73 bl[73] br[73] wl[99] vdd gnd cell_6t
Xbit_r100_c73 bl[73] br[73] wl[100] vdd gnd cell_6t
Xbit_r101_c73 bl[73] br[73] wl[101] vdd gnd cell_6t
Xbit_r102_c73 bl[73] br[73] wl[102] vdd gnd cell_6t
Xbit_r103_c73 bl[73] br[73] wl[103] vdd gnd cell_6t
Xbit_r104_c73 bl[73] br[73] wl[104] vdd gnd cell_6t
Xbit_r105_c73 bl[73] br[73] wl[105] vdd gnd cell_6t
Xbit_r106_c73 bl[73] br[73] wl[106] vdd gnd cell_6t
Xbit_r107_c73 bl[73] br[73] wl[107] vdd gnd cell_6t
Xbit_r108_c73 bl[73] br[73] wl[108] vdd gnd cell_6t
Xbit_r109_c73 bl[73] br[73] wl[109] vdd gnd cell_6t
Xbit_r110_c73 bl[73] br[73] wl[110] vdd gnd cell_6t
Xbit_r111_c73 bl[73] br[73] wl[111] vdd gnd cell_6t
Xbit_r112_c73 bl[73] br[73] wl[112] vdd gnd cell_6t
Xbit_r113_c73 bl[73] br[73] wl[113] vdd gnd cell_6t
Xbit_r114_c73 bl[73] br[73] wl[114] vdd gnd cell_6t
Xbit_r115_c73 bl[73] br[73] wl[115] vdd gnd cell_6t
Xbit_r116_c73 bl[73] br[73] wl[116] vdd gnd cell_6t
Xbit_r117_c73 bl[73] br[73] wl[117] vdd gnd cell_6t
Xbit_r118_c73 bl[73] br[73] wl[118] vdd gnd cell_6t
Xbit_r119_c73 bl[73] br[73] wl[119] vdd gnd cell_6t
Xbit_r120_c73 bl[73] br[73] wl[120] vdd gnd cell_6t
Xbit_r121_c73 bl[73] br[73] wl[121] vdd gnd cell_6t
Xbit_r122_c73 bl[73] br[73] wl[122] vdd gnd cell_6t
Xbit_r123_c73 bl[73] br[73] wl[123] vdd gnd cell_6t
Xbit_r124_c73 bl[73] br[73] wl[124] vdd gnd cell_6t
Xbit_r125_c73 bl[73] br[73] wl[125] vdd gnd cell_6t
Xbit_r126_c73 bl[73] br[73] wl[126] vdd gnd cell_6t
Xbit_r127_c73 bl[73] br[73] wl[127] vdd gnd cell_6t
Xbit_r128_c73 bl[73] br[73] wl[128] vdd gnd cell_6t
Xbit_r129_c73 bl[73] br[73] wl[129] vdd gnd cell_6t
Xbit_r130_c73 bl[73] br[73] wl[130] vdd gnd cell_6t
Xbit_r131_c73 bl[73] br[73] wl[131] vdd gnd cell_6t
Xbit_r132_c73 bl[73] br[73] wl[132] vdd gnd cell_6t
Xbit_r133_c73 bl[73] br[73] wl[133] vdd gnd cell_6t
Xbit_r134_c73 bl[73] br[73] wl[134] vdd gnd cell_6t
Xbit_r135_c73 bl[73] br[73] wl[135] vdd gnd cell_6t
Xbit_r136_c73 bl[73] br[73] wl[136] vdd gnd cell_6t
Xbit_r137_c73 bl[73] br[73] wl[137] vdd gnd cell_6t
Xbit_r138_c73 bl[73] br[73] wl[138] vdd gnd cell_6t
Xbit_r139_c73 bl[73] br[73] wl[139] vdd gnd cell_6t
Xbit_r140_c73 bl[73] br[73] wl[140] vdd gnd cell_6t
Xbit_r141_c73 bl[73] br[73] wl[141] vdd gnd cell_6t
Xbit_r142_c73 bl[73] br[73] wl[142] vdd gnd cell_6t
Xbit_r143_c73 bl[73] br[73] wl[143] vdd gnd cell_6t
Xbit_r144_c73 bl[73] br[73] wl[144] vdd gnd cell_6t
Xbit_r145_c73 bl[73] br[73] wl[145] vdd gnd cell_6t
Xbit_r146_c73 bl[73] br[73] wl[146] vdd gnd cell_6t
Xbit_r147_c73 bl[73] br[73] wl[147] vdd gnd cell_6t
Xbit_r148_c73 bl[73] br[73] wl[148] vdd gnd cell_6t
Xbit_r149_c73 bl[73] br[73] wl[149] vdd gnd cell_6t
Xbit_r150_c73 bl[73] br[73] wl[150] vdd gnd cell_6t
Xbit_r151_c73 bl[73] br[73] wl[151] vdd gnd cell_6t
Xbit_r152_c73 bl[73] br[73] wl[152] vdd gnd cell_6t
Xbit_r153_c73 bl[73] br[73] wl[153] vdd gnd cell_6t
Xbit_r154_c73 bl[73] br[73] wl[154] vdd gnd cell_6t
Xbit_r155_c73 bl[73] br[73] wl[155] vdd gnd cell_6t
Xbit_r156_c73 bl[73] br[73] wl[156] vdd gnd cell_6t
Xbit_r157_c73 bl[73] br[73] wl[157] vdd gnd cell_6t
Xbit_r158_c73 bl[73] br[73] wl[158] vdd gnd cell_6t
Xbit_r159_c73 bl[73] br[73] wl[159] vdd gnd cell_6t
Xbit_r160_c73 bl[73] br[73] wl[160] vdd gnd cell_6t
Xbit_r161_c73 bl[73] br[73] wl[161] vdd gnd cell_6t
Xbit_r162_c73 bl[73] br[73] wl[162] vdd gnd cell_6t
Xbit_r163_c73 bl[73] br[73] wl[163] vdd gnd cell_6t
Xbit_r164_c73 bl[73] br[73] wl[164] vdd gnd cell_6t
Xbit_r165_c73 bl[73] br[73] wl[165] vdd gnd cell_6t
Xbit_r166_c73 bl[73] br[73] wl[166] vdd gnd cell_6t
Xbit_r167_c73 bl[73] br[73] wl[167] vdd gnd cell_6t
Xbit_r168_c73 bl[73] br[73] wl[168] vdd gnd cell_6t
Xbit_r169_c73 bl[73] br[73] wl[169] vdd gnd cell_6t
Xbit_r170_c73 bl[73] br[73] wl[170] vdd gnd cell_6t
Xbit_r171_c73 bl[73] br[73] wl[171] vdd gnd cell_6t
Xbit_r172_c73 bl[73] br[73] wl[172] vdd gnd cell_6t
Xbit_r173_c73 bl[73] br[73] wl[173] vdd gnd cell_6t
Xbit_r174_c73 bl[73] br[73] wl[174] vdd gnd cell_6t
Xbit_r175_c73 bl[73] br[73] wl[175] vdd gnd cell_6t
Xbit_r176_c73 bl[73] br[73] wl[176] vdd gnd cell_6t
Xbit_r177_c73 bl[73] br[73] wl[177] vdd gnd cell_6t
Xbit_r178_c73 bl[73] br[73] wl[178] vdd gnd cell_6t
Xbit_r179_c73 bl[73] br[73] wl[179] vdd gnd cell_6t
Xbit_r180_c73 bl[73] br[73] wl[180] vdd gnd cell_6t
Xbit_r181_c73 bl[73] br[73] wl[181] vdd gnd cell_6t
Xbit_r182_c73 bl[73] br[73] wl[182] vdd gnd cell_6t
Xbit_r183_c73 bl[73] br[73] wl[183] vdd gnd cell_6t
Xbit_r184_c73 bl[73] br[73] wl[184] vdd gnd cell_6t
Xbit_r185_c73 bl[73] br[73] wl[185] vdd gnd cell_6t
Xbit_r186_c73 bl[73] br[73] wl[186] vdd gnd cell_6t
Xbit_r187_c73 bl[73] br[73] wl[187] vdd gnd cell_6t
Xbit_r188_c73 bl[73] br[73] wl[188] vdd gnd cell_6t
Xbit_r189_c73 bl[73] br[73] wl[189] vdd gnd cell_6t
Xbit_r190_c73 bl[73] br[73] wl[190] vdd gnd cell_6t
Xbit_r191_c73 bl[73] br[73] wl[191] vdd gnd cell_6t
Xbit_r192_c73 bl[73] br[73] wl[192] vdd gnd cell_6t
Xbit_r193_c73 bl[73] br[73] wl[193] vdd gnd cell_6t
Xbit_r194_c73 bl[73] br[73] wl[194] vdd gnd cell_6t
Xbit_r195_c73 bl[73] br[73] wl[195] vdd gnd cell_6t
Xbit_r196_c73 bl[73] br[73] wl[196] vdd gnd cell_6t
Xbit_r197_c73 bl[73] br[73] wl[197] vdd gnd cell_6t
Xbit_r198_c73 bl[73] br[73] wl[198] vdd gnd cell_6t
Xbit_r199_c73 bl[73] br[73] wl[199] vdd gnd cell_6t
Xbit_r200_c73 bl[73] br[73] wl[200] vdd gnd cell_6t
Xbit_r201_c73 bl[73] br[73] wl[201] vdd gnd cell_6t
Xbit_r202_c73 bl[73] br[73] wl[202] vdd gnd cell_6t
Xbit_r203_c73 bl[73] br[73] wl[203] vdd gnd cell_6t
Xbit_r204_c73 bl[73] br[73] wl[204] vdd gnd cell_6t
Xbit_r205_c73 bl[73] br[73] wl[205] vdd gnd cell_6t
Xbit_r206_c73 bl[73] br[73] wl[206] vdd gnd cell_6t
Xbit_r207_c73 bl[73] br[73] wl[207] vdd gnd cell_6t
Xbit_r208_c73 bl[73] br[73] wl[208] vdd gnd cell_6t
Xbit_r209_c73 bl[73] br[73] wl[209] vdd gnd cell_6t
Xbit_r210_c73 bl[73] br[73] wl[210] vdd gnd cell_6t
Xbit_r211_c73 bl[73] br[73] wl[211] vdd gnd cell_6t
Xbit_r212_c73 bl[73] br[73] wl[212] vdd gnd cell_6t
Xbit_r213_c73 bl[73] br[73] wl[213] vdd gnd cell_6t
Xbit_r214_c73 bl[73] br[73] wl[214] vdd gnd cell_6t
Xbit_r215_c73 bl[73] br[73] wl[215] vdd gnd cell_6t
Xbit_r216_c73 bl[73] br[73] wl[216] vdd gnd cell_6t
Xbit_r217_c73 bl[73] br[73] wl[217] vdd gnd cell_6t
Xbit_r218_c73 bl[73] br[73] wl[218] vdd gnd cell_6t
Xbit_r219_c73 bl[73] br[73] wl[219] vdd gnd cell_6t
Xbit_r220_c73 bl[73] br[73] wl[220] vdd gnd cell_6t
Xbit_r221_c73 bl[73] br[73] wl[221] vdd gnd cell_6t
Xbit_r222_c73 bl[73] br[73] wl[222] vdd gnd cell_6t
Xbit_r223_c73 bl[73] br[73] wl[223] vdd gnd cell_6t
Xbit_r224_c73 bl[73] br[73] wl[224] vdd gnd cell_6t
Xbit_r225_c73 bl[73] br[73] wl[225] vdd gnd cell_6t
Xbit_r226_c73 bl[73] br[73] wl[226] vdd gnd cell_6t
Xbit_r227_c73 bl[73] br[73] wl[227] vdd gnd cell_6t
Xbit_r228_c73 bl[73] br[73] wl[228] vdd gnd cell_6t
Xbit_r229_c73 bl[73] br[73] wl[229] vdd gnd cell_6t
Xbit_r230_c73 bl[73] br[73] wl[230] vdd gnd cell_6t
Xbit_r231_c73 bl[73] br[73] wl[231] vdd gnd cell_6t
Xbit_r232_c73 bl[73] br[73] wl[232] vdd gnd cell_6t
Xbit_r233_c73 bl[73] br[73] wl[233] vdd gnd cell_6t
Xbit_r234_c73 bl[73] br[73] wl[234] vdd gnd cell_6t
Xbit_r235_c73 bl[73] br[73] wl[235] vdd gnd cell_6t
Xbit_r236_c73 bl[73] br[73] wl[236] vdd gnd cell_6t
Xbit_r237_c73 bl[73] br[73] wl[237] vdd gnd cell_6t
Xbit_r238_c73 bl[73] br[73] wl[238] vdd gnd cell_6t
Xbit_r239_c73 bl[73] br[73] wl[239] vdd gnd cell_6t
Xbit_r240_c73 bl[73] br[73] wl[240] vdd gnd cell_6t
Xbit_r241_c73 bl[73] br[73] wl[241] vdd gnd cell_6t
Xbit_r242_c73 bl[73] br[73] wl[242] vdd gnd cell_6t
Xbit_r243_c73 bl[73] br[73] wl[243] vdd gnd cell_6t
Xbit_r244_c73 bl[73] br[73] wl[244] vdd gnd cell_6t
Xbit_r245_c73 bl[73] br[73] wl[245] vdd gnd cell_6t
Xbit_r246_c73 bl[73] br[73] wl[246] vdd gnd cell_6t
Xbit_r247_c73 bl[73] br[73] wl[247] vdd gnd cell_6t
Xbit_r248_c73 bl[73] br[73] wl[248] vdd gnd cell_6t
Xbit_r249_c73 bl[73] br[73] wl[249] vdd gnd cell_6t
Xbit_r250_c73 bl[73] br[73] wl[250] vdd gnd cell_6t
Xbit_r251_c73 bl[73] br[73] wl[251] vdd gnd cell_6t
Xbit_r252_c73 bl[73] br[73] wl[252] vdd gnd cell_6t
Xbit_r253_c73 bl[73] br[73] wl[253] vdd gnd cell_6t
Xbit_r254_c73 bl[73] br[73] wl[254] vdd gnd cell_6t
Xbit_r255_c73 bl[73] br[73] wl[255] vdd gnd cell_6t
Xbit_r256_c73 bl[73] br[73] wl[256] vdd gnd cell_6t
Xbit_r257_c73 bl[73] br[73] wl[257] vdd gnd cell_6t
Xbit_r258_c73 bl[73] br[73] wl[258] vdd gnd cell_6t
Xbit_r259_c73 bl[73] br[73] wl[259] vdd gnd cell_6t
Xbit_r260_c73 bl[73] br[73] wl[260] vdd gnd cell_6t
Xbit_r261_c73 bl[73] br[73] wl[261] vdd gnd cell_6t
Xbit_r262_c73 bl[73] br[73] wl[262] vdd gnd cell_6t
Xbit_r263_c73 bl[73] br[73] wl[263] vdd gnd cell_6t
Xbit_r264_c73 bl[73] br[73] wl[264] vdd gnd cell_6t
Xbit_r265_c73 bl[73] br[73] wl[265] vdd gnd cell_6t
Xbit_r266_c73 bl[73] br[73] wl[266] vdd gnd cell_6t
Xbit_r267_c73 bl[73] br[73] wl[267] vdd gnd cell_6t
Xbit_r268_c73 bl[73] br[73] wl[268] vdd gnd cell_6t
Xbit_r269_c73 bl[73] br[73] wl[269] vdd gnd cell_6t
Xbit_r270_c73 bl[73] br[73] wl[270] vdd gnd cell_6t
Xbit_r271_c73 bl[73] br[73] wl[271] vdd gnd cell_6t
Xbit_r272_c73 bl[73] br[73] wl[272] vdd gnd cell_6t
Xbit_r273_c73 bl[73] br[73] wl[273] vdd gnd cell_6t
Xbit_r274_c73 bl[73] br[73] wl[274] vdd gnd cell_6t
Xbit_r275_c73 bl[73] br[73] wl[275] vdd gnd cell_6t
Xbit_r276_c73 bl[73] br[73] wl[276] vdd gnd cell_6t
Xbit_r277_c73 bl[73] br[73] wl[277] vdd gnd cell_6t
Xbit_r278_c73 bl[73] br[73] wl[278] vdd gnd cell_6t
Xbit_r279_c73 bl[73] br[73] wl[279] vdd gnd cell_6t
Xbit_r280_c73 bl[73] br[73] wl[280] vdd gnd cell_6t
Xbit_r281_c73 bl[73] br[73] wl[281] vdd gnd cell_6t
Xbit_r282_c73 bl[73] br[73] wl[282] vdd gnd cell_6t
Xbit_r283_c73 bl[73] br[73] wl[283] vdd gnd cell_6t
Xbit_r284_c73 bl[73] br[73] wl[284] vdd gnd cell_6t
Xbit_r285_c73 bl[73] br[73] wl[285] vdd gnd cell_6t
Xbit_r286_c73 bl[73] br[73] wl[286] vdd gnd cell_6t
Xbit_r287_c73 bl[73] br[73] wl[287] vdd gnd cell_6t
Xbit_r288_c73 bl[73] br[73] wl[288] vdd gnd cell_6t
Xbit_r289_c73 bl[73] br[73] wl[289] vdd gnd cell_6t
Xbit_r290_c73 bl[73] br[73] wl[290] vdd gnd cell_6t
Xbit_r291_c73 bl[73] br[73] wl[291] vdd gnd cell_6t
Xbit_r292_c73 bl[73] br[73] wl[292] vdd gnd cell_6t
Xbit_r293_c73 bl[73] br[73] wl[293] vdd gnd cell_6t
Xbit_r294_c73 bl[73] br[73] wl[294] vdd gnd cell_6t
Xbit_r295_c73 bl[73] br[73] wl[295] vdd gnd cell_6t
Xbit_r296_c73 bl[73] br[73] wl[296] vdd gnd cell_6t
Xbit_r297_c73 bl[73] br[73] wl[297] vdd gnd cell_6t
Xbit_r298_c73 bl[73] br[73] wl[298] vdd gnd cell_6t
Xbit_r299_c73 bl[73] br[73] wl[299] vdd gnd cell_6t
Xbit_r300_c73 bl[73] br[73] wl[300] vdd gnd cell_6t
Xbit_r301_c73 bl[73] br[73] wl[301] vdd gnd cell_6t
Xbit_r302_c73 bl[73] br[73] wl[302] vdd gnd cell_6t
Xbit_r303_c73 bl[73] br[73] wl[303] vdd gnd cell_6t
Xbit_r304_c73 bl[73] br[73] wl[304] vdd gnd cell_6t
Xbit_r305_c73 bl[73] br[73] wl[305] vdd gnd cell_6t
Xbit_r306_c73 bl[73] br[73] wl[306] vdd gnd cell_6t
Xbit_r307_c73 bl[73] br[73] wl[307] vdd gnd cell_6t
Xbit_r308_c73 bl[73] br[73] wl[308] vdd gnd cell_6t
Xbit_r309_c73 bl[73] br[73] wl[309] vdd gnd cell_6t
Xbit_r310_c73 bl[73] br[73] wl[310] vdd gnd cell_6t
Xbit_r311_c73 bl[73] br[73] wl[311] vdd gnd cell_6t
Xbit_r312_c73 bl[73] br[73] wl[312] vdd gnd cell_6t
Xbit_r313_c73 bl[73] br[73] wl[313] vdd gnd cell_6t
Xbit_r314_c73 bl[73] br[73] wl[314] vdd gnd cell_6t
Xbit_r315_c73 bl[73] br[73] wl[315] vdd gnd cell_6t
Xbit_r316_c73 bl[73] br[73] wl[316] vdd gnd cell_6t
Xbit_r317_c73 bl[73] br[73] wl[317] vdd gnd cell_6t
Xbit_r318_c73 bl[73] br[73] wl[318] vdd gnd cell_6t
Xbit_r319_c73 bl[73] br[73] wl[319] vdd gnd cell_6t
Xbit_r320_c73 bl[73] br[73] wl[320] vdd gnd cell_6t
Xbit_r321_c73 bl[73] br[73] wl[321] vdd gnd cell_6t
Xbit_r322_c73 bl[73] br[73] wl[322] vdd gnd cell_6t
Xbit_r323_c73 bl[73] br[73] wl[323] vdd gnd cell_6t
Xbit_r324_c73 bl[73] br[73] wl[324] vdd gnd cell_6t
Xbit_r325_c73 bl[73] br[73] wl[325] vdd gnd cell_6t
Xbit_r326_c73 bl[73] br[73] wl[326] vdd gnd cell_6t
Xbit_r327_c73 bl[73] br[73] wl[327] vdd gnd cell_6t
Xbit_r328_c73 bl[73] br[73] wl[328] vdd gnd cell_6t
Xbit_r329_c73 bl[73] br[73] wl[329] vdd gnd cell_6t
Xbit_r330_c73 bl[73] br[73] wl[330] vdd gnd cell_6t
Xbit_r331_c73 bl[73] br[73] wl[331] vdd gnd cell_6t
Xbit_r332_c73 bl[73] br[73] wl[332] vdd gnd cell_6t
Xbit_r333_c73 bl[73] br[73] wl[333] vdd gnd cell_6t
Xbit_r334_c73 bl[73] br[73] wl[334] vdd gnd cell_6t
Xbit_r335_c73 bl[73] br[73] wl[335] vdd gnd cell_6t
Xbit_r336_c73 bl[73] br[73] wl[336] vdd gnd cell_6t
Xbit_r337_c73 bl[73] br[73] wl[337] vdd gnd cell_6t
Xbit_r338_c73 bl[73] br[73] wl[338] vdd gnd cell_6t
Xbit_r339_c73 bl[73] br[73] wl[339] vdd gnd cell_6t
Xbit_r340_c73 bl[73] br[73] wl[340] vdd gnd cell_6t
Xbit_r341_c73 bl[73] br[73] wl[341] vdd gnd cell_6t
Xbit_r342_c73 bl[73] br[73] wl[342] vdd gnd cell_6t
Xbit_r343_c73 bl[73] br[73] wl[343] vdd gnd cell_6t
Xbit_r344_c73 bl[73] br[73] wl[344] vdd gnd cell_6t
Xbit_r345_c73 bl[73] br[73] wl[345] vdd gnd cell_6t
Xbit_r346_c73 bl[73] br[73] wl[346] vdd gnd cell_6t
Xbit_r347_c73 bl[73] br[73] wl[347] vdd gnd cell_6t
Xbit_r348_c73 bl[73] br[73] wl[348] vdd gnd cell_6t
Xbit_r349_c73 bl[73] br[73] wl[349] vdd gnd cell_6t
Xbit_r350_c73 bl[73] br[73] wl[350] vdd gnd cell_6t
Xbit_r351_c73 bl[73] br[73] wl[351] vdd gnd cell_6t
Xbit_r352_c73 bl[73] br[73] wl[352] vdd gnd cell_6t
Xbit_r353_c73 bl[73] br[73] wl[353] vdd gnd cell_6t
Xbit_r354_c73 bl[73] br[73] wl[354] vdd gnd cell_6t
Xbit_r355_c73 bl[73] br[73] wl[355] vdd gnd cell_6t
Xbit_r356_c73 bl[73] br[73] wl[356] vdd gnd cell_6t
Xbit_r357_c73 bl[73] br[73] wl[357] vdd gnd cell_6t
Xbit_r358_c73 bl[73] br[73] wl[358] vdd gnd cell_6t
Xbit_r359_c73 bl[73] br[73] wl[359] vdd gnd cell_6t
Xbit_r360_c73 bl[73] br[73] wl[360] vdd gnd cell_6t
Xbit_r361_c73 bl[73] br[73] wl[361] vdd gnd cell_6t
Xbit_r362_c73 bl[73] br[73] wl[362] vdd gnd cell_6t
Xbit_r363_c73 bl[73] br[73] wl[363] vdd gnd cell_6t
Xbit_r364_c73 bl[73] br[73] wl[364] vdd gnd cell_6t
Xbit_r365_c73 bl[73] br[73] wl[365] vdd gnd cell_6t
Xbit_r366_c73 bl[73] br[73] wl[366] vdd gnd cell_6t
Xbit_r367_c73 bl[73] br[73] wl[367] vdd gnd cell_6t
Xbit_r368_c73 bl[73] br[73] wl[368] vdd gnd cell_6t
Xbit_r369_c73 bl[73] br[73] wl[369] vdd gnd cell_6t
Xbit_r370_c73 bl[73] br[73] wl[370] vdd gnd cell_6t
Xbit_r371_c73 bl[73] br[73] wl[371] vdd gnd cell_6t
Xbit_r372_c73 bl[73] br[73] wl[372] vdd gnd cell_6t
Xbit_r373_c73 bl[73] br[73] wl[373] vdd gnd cell_6t
Xbit_r374_c73 bl[73] br[73] wl[374] vdd gnd cell_6t
Xbit_r375_c73 bl[73] br[73] wl[375] vdd gnd cell_6t
Xbit_r376_c73 bl[73] br[73] wl[376] vdd gnd cell_6t
Xbit_r377_c73 bl[73] br[73] wl[377] vdd gnd cell_6t
Xbit_r378_c73 bl[73] br[73] wl[378] vdd gnd cell_6t
Xbit_r379_c73 bl[73] br[73] wl[379] vdd gnd cell_6t
Xbit_r380_c73 bl[73] br[73] wl[380] vdd gnd cell_6t
Xbit_r381_c73 bl[73] br[73] wl[381] vdd gnd cell_6t
Xbit_r382_c73 bl[73] br[73] wl[382] vdd gnd cell_6t
Xbit_r383_c73 bl[73] br[73] wl[383] vdd gnd cell_6t
Xbit_r384_c73 bl[73] br[73] wl[384] vdd gnd cell_6t
Xbit_r385_c73 bl[73] br[73] wl[385] vdd gnd cell_6t
Xbit_r386_c73 bl[73] br[73] wl[386] vdd gnd cell_6t
Xbit_r387_c73 bl[73] br[73] wl[387] vdd gnd cell_6t
Xbit_r388_c73 bl[73] br[73] wl[388] vdd gnd cell_6t
Xbit_r389_c73 bl[73] br[73] wl[389] vdd gnd cell_6t
Xbit_r390_c73 bl[73] br[73] wl[390] vdd gnd cell_6t
Xbit_r391_c73 bl[73] br[73] wl[391] vdd gnd cell_6t
Xbit_r392_c73 bl[73] br[73] wl[392] vdd gnd cell_6t
Xbit_r393_c73 bl[73] br[73] wl[393] vdd gnd cell_6t
Xbit_r394_c73 bl[73] br[73] wl[394] vdd gnd cell_6t
Xbit_r395_c73 bl[73] br[73] wl[395] vdd gnd cell_6t
Xbit_r396_c73 bl[73] br[73] wl[396] vdd gnd cell_6t
Xbit_r397_c73 bl[73] br[73] wl[397] vdd gnd cell_6t
Xbit_r398_c73 bl[73] br[73] wl[398] vdd gnd cell_6t
Xbit_r399_c73 bl[73] br[73] wl[399] vdd gnd cell_6t
Xbit_r400_c73 bl[73] br[73] wl[400] vdd gnd cell_6t
Xbit_r401_c73 bl[73] br[73] wl[401] vdd gnd cell_6t
Xbit_r402_c73 bl[73] br[73] wl[402] vdd gnd cell_6t
Xbit_r403_c73 bl[73] br[73] wl[403] vdd gnd cell_6t
Xbit_r404_c73 bl[73] br[73] wl[404] vdd gnd cell_6t
Xbit_r405_c73 bl[73] br[73] wl[405] vdd gnd cell_6t
Xbit_r406_c73 bl[73] br[73] wl[406] vdd gnd cell_6t
Xbit_r407_c73 bl[73] br[73] wl[407] vdd gnd cell_6t
Xbit_r408_c73 bl[73] br[73] wl[408] vdd gnd cell_6t
Xbit_r409_c73 bl[73] br[73] wl[409] vdd gnd cell_6t
Xbit_r410_c73 bl[73] br[73] wl[410] vdd gnd cell_6t
Xbit_r411_c73 bl[73] br[73] wl[411] vdd gnd cell_6t
Xbit_r412_c73 bl[73] br[73] wl[412] vdd gnd cell_6t
Xbit_r413_c73 bl[73] br[73] wl[413] vdd gnd cell_6t
Xbit_r414_c73 bl[73] br[73] wl[414] vdd gnd cell_6t
Xbit_r415_c73 bl[73] br[73] wl[415] vdd gnd cell_6t
Xbit_r416_c73 bl[73] br[73] wl[416] vdd gnd cell_6t
Xbit_r417_c73 bl[73] br[73] wl[417] vdd gnd cell_6t
Xbit_r418_c73 bl[73] br[73] wl[418] vdd gnd cell_6t
Xbit_r419_c73 bl[73] br[73] wl[419] vdd gnd cell_6t
Xbit_r420_c73 bl[73] br[73] wl[420] vdd gnd cell_6t
Xbit_r421_c73 bl[73] br[73] wl[421] vdd gnd cell_6t
Xbit_r422_c73 bl[73] br[73] wl[422] vdd gnd cell_6t
Xbit_r423_c73 bl[73] br[73] wl[423] vdd gnd cell_6t
Xbit_r424_c73 bl[73] br[73] wl[424] vdd gnd cell_6t
Xbit_r425_c73 bl[73] br[73] wl[425] vdd gnd cell_6t
Xbit_r426_c73 bl[73] br[73] wl[426] vdd gnd cell_6t
Xbit_r427_c73 bl[73] br[73] wl[427] vdd gnd cell_6t
Xbit_r428_c73 bl[73] br[73] wl[428] vdd gnd cell_6t
Xbit_r429_c73 bl[73] br[73] wl[429] vdd gnd cell_6t
Xbit_r430_c73 bl[73] br[73] wl[430] vdd gnd cell_6t
Xbit_r431_c73 bl[73] br[73] wl[431] vdd gnd cell_6t
Xbit_r432_c73 bl[73] br[73] wl[432] vdd gnd cell_6t
Xbit_r433_c73 bl[73] br[73] wl[433] vdd gnd cell_6t
Xbit_r434_c73 bl[73] br[73] wl[434] vdd gnd cell_6t
Xbit_r435_c73 bl[73] br[73] wl[435] vdd gnd cell_6t
Xbit_r436_c73 bl[73] br[73] wl[436] vdd gnd cell_6t
Xbit_r437_c73 bl[73] br[73] wl[437] vdd gnd cell_6t
Xbit_r438_c73 bl[73] br[73] wl[438] vdd gnd cell_6t
Xbit_r439_c73 bl[73] br[73] wl[439] vdd gnd cell_6t
Xbit_r440_c73 bl[73] br[73] wl[440] vdd gnd cell_6t
Xbit_r441_c73 bl[73] br[73] wl[441] vdd gnd cell_6t
Xbit_r442_c73 bl[73] br[73] wl[442] vdd gnd cell_6t
Xbit_r443_c73 bl[73] br[73] wl[443] vdd gnd cell_6t
Xbit_r444_c73 bl[73] br[73] wl[444] vdd gnd cell_6t
Xbit_r445_c73 bl[73] br[73] wl[445] vdd gnd cell_6t
Xbit_r446_c73 bl[73] br[73] wl[446] vdd gnd cell_6t
Xbit_r447_c73 bl[73] br[73] wl[447] vdd gnd cell_6t
Xbit_r448_c73 bl[73] br[73] wl[448] vdd gnd cell_6t
Xbit_r449_c73 bl[73] br[73] wl[449] vdd gnd cell_6t
Xbit_r450_c73 bl[73] br[73] wl[450] vdd gnd cell_6t
Xbit_r451_c73 bl[73] br[73] wl[451] vdd gnd cell_6t
Xbit_r452_c73 bl[73] br[73] wl[452] vdd gnd cell_6t
Xbit_r453_c73 bl[73] br[73] wl[453] vdd gnd cell_6t
Xbit_r454_c73 bl[73] br[73] wl[454] vdd gnd cell_6t
Xbit_r455_c73 bl[73] br[73] wl[455] vdd gnd cell_6t
Xbit_r456_c73 bl[73] br[73] wl[456] vdd gnd cell_6t
Xbit_r457_c73 bl[73] br[73] wl[457] vdd gnd cell_6t
Xbit_r458_c73 bl[73] br[73] wl[458] vdd gnd cell_6t
Xbit_r459_c73 bl[73] br[73] wl[459] vdd gnd cell_6t
Xbit_r460_c73 bl[73] br[73] wl[460] vdd gnd cell_6t
Xbit_r461_c73 bl[73] br[73] wl[461] vdd gnd cell_6t
Xbit_r462_c73 bl[73] br[73] wl[462] vdd gnd cell_6t
Xbit_r463_c73 bl[73] br[73] wl[463] vdd gnd cell_6t
Xbit_r464_c73 bl[73] br[73] wl[464] vdd gnd cell_6t
Xbit_r465_c73 bl[73] br[73] wl[465] vdd gnd cell_6t
Xbit_r466_c73 bl[73] br[73] wl[466] vdd gnd cell_6t
Xbit_r467_c73 bl[73] br[73] wl[467] vdd gnd cell_6t
Xbit_r468_c73 bl[73] br[73] wl[468] vdd gnd cell_6t
Xbit_r469_c73 bl[73] br[73] wl[469] vdd gnd cell_6t
Xbit_r470_c73 bl[73] br[73] wl[470] vdd gnd cell_6t
Xbit_r471_c73 bl[73] br[73] wl[471] vdd gnd cell_6t
Xbit_r472_c73 bl[73] br[73] wl[472] vdd gnd cell_6t
Xbit_r473_c73 bl[73] br[73] wl[473] vdd gnd cell_6t
Xbit_r474_c73 bl[73] br[73] wl[474] vdd gnd cell_6t
Xbit_r475_c73 bl[73] br[73] wl[475] vdd gnd cell_6t
Xbit_r476_c73 bl[73] br[73] wl[476] vdd gnd cell_6t
Xbit_r477_c73 bl[73] br[73] wl[477] vdd gnd cell_6t
Xbit_r478_c73 bl[73] br[73] wl[478] vdd gnd cell_6t
Xbit_r479_c73 bl[73] br[73] wl[479] vdd gnd cell_6t
Xbit_r480_c73 bl[73] br[73] wl[480] vdd gnd cell_6t
Xbit_r481_c73 bl[73] br[73] wl[481] vdd gnd cell_6t
Xbit_r482_c73 bl[73] br[73] wl[482] vdd gnd cell_6t
Xbit_r483_c73 bl[73] br[73] wl[483] vdd gnd cell_6t
Xbit_r484_c73 bl[73] br[73] wl[484] vdd gnd cell_6t
Xbit_r485_c73 bl[73] br[73] wl[485] vdd gnd cell_6t
Xbit_r486_c73 bl[73] br[73] wl[486] vdd gnd cell_6t
Xbit_r487_c73 bl[73] br[73] wl[487] vdd gnd cell_6t
Xbit_r488_c73 bl[73] br[73] wl[488] vdd gnd cell_6t
Xbit_r489_c73 bl[73] br[73] wl[489] vdd gnd cell_6t
Xbit_r490_c73 bl[73] br[73] wl[490] vdd gnd cell_6t
Xbit_r491_c73 bl[73] br[73] wl[491] vdd gnd cell_6t
Xbit_r492_c73 bl[73] br[73] wl[492] vdd gnd cell_6t
Xbit_r493_c73 bl[73] br[73] wl[493] vdd gnd cell_6t
Xbit_r494_c73 bl[73] br[73] wl[494] vdd gnd cell_6t
Xbit_r495_c73 bl[73] br[73] wl[495] vdd gnd cell_6t
Xbit_r496_c73 bl[73] br[73] wl[496] vdd gnd cell_6t
Xbit_r497_c73 bl[73] br[73] wl[497] vdd gnd cell_6t
Xbit_r498_c73 bl[73] br[73] wl[498] vdd gnd cell_6t
Xbit_r499_c73 bl[73] br[73] wl[499] vdd gnd cell_6t
Xbit_r500_c73 bl[73] br[73] wl[500] vdd gnd cell_6t
Xbit_r501_c73 bl[73] br[73] wl[501] vdd gnd cell_6t
Xbit_r502_c73 bl[73] br[73] wl[502] vdd gnd cell_6t
Xbit_r503_c73 bl[73] br[73] wl[503] vdd gnd cell_6t
Xbit_r504_c73 bl[73] br[73] wl[504] vdd gnd cell_6t
Xbit_r505_c73 bl[73] br[73] wl[505] vdd gnd cell_6t
Xbit_r506_c73 bl[73] br[73] wl[506] vdd gnd cell_6t
Xbit_r507_c73 bl[73] br[73] wl[507] vdd gnd cell_6t
Xbit_r508_c73 bl[73] br[73] wl[508] vdd gnd cell_6t
Xbit_r509_c73 bl[73] br[73] wl[509] vdd gnd cell_6t
Xbit_r510_c73 bl[73] br[73] wl[510] vdd gnd cell_6t
Xbit_r511_c73 bl[73] br[73] wl[511] vdd gnd cell_6t
Xbit_r0_c74 bl[74] br[74] wl[0] vdd gnd cell_6t
Xbit_r1_c74 bl[74] br[74] wl[1] vdd gnd cell_6t
Xbit_r2_c74 bl[74] br[74] wl[2] vdd gnd cell_6t
Xbit_r3_c74 bl[74] br[74] wl[3] vdd gnd cell_6t
Xbit_r4_c74 bl[74] br[74] wl[4] vdd gnd cell_6t
Xbit_r5_c74 bl[74] br[74] wl[5] vdd gnd cell_6t
Xbit_r6_c74 bl[74] br[74] wl[6] vdd gnd cell_6t
Xbit_r7_c74 bl[74] br[74] wl[7] vdd gnd cell_6t
Xbit_r8_c74 bl[74] br[74] wl[8] vdd gnd cell_6t
Xbit_r9_c74 bl[74] br[74] wl[9] vdd gnd cell_6t
Xbit_r10_c74 bl[74] br[74] wl[10] vdd gnd cell_6t
Xbit_r11_c74 bl[74] br[74] wl[11] vdd gnd cell_6t
Xbit_r12_c74 bl[74] br[74] wl[12] vdd gnd cell_6t
Xbit_r13_c74 bl[74] br[74] wl[13] vdd gnd cell_6t
Xbit_r14_c74 bl[74] br[74] wl[14] vdd gnd cell_6t
Xbit_r15_c74 bl[74] br[74] wl[15] vdd gnd cell_6t
Xbit_r16_c74 bl[74] br[74] wl[16] vdd gnd cell_6t
Xbit_r17_c74 bl[74] br[74] wl[17] vdd gnd cell_6t
Xbit_r18_c74 bl[74] br[74] wl[18] vdd gnd cell_6t
Xbit_r19_c74 bl[74] br[74] wl[19] vdd gnd cell_6t
Xbit_r20_c74 bl[74] br[74] wl[20] vdd gnd cell_6t
Xbit_r21_c74 bl[74] br[74] wl[21] vdd gnd cell_6t
Xbit_r22_c74 bl[74] br[74] wl[22] vdd gnd cell_6t
Xbit_r23_c74 bl[74] br[74] wl[23] vdd gnd cell_6t
Xbit_r24_c74 bl[74] br[74] wl[24] vdd gnd cell_6t
Xbit_r25_c74 bl[74] br[74] wl[25] vdd gnd cell_6t
Xbit_r26_c74 bl[74] br[74] wl[26] vdd gnd cell_6t
Xbit_r27_c74 bl[74] br[74] wl[27] vdd gnd cell_6t
Xbit_r28_c74 bl[74] br[74] wl[28] vdd gnd cell_6t
Xbit_r29_c74 bl[74] br[74] wl[29] vdd gnd cell_6t
Xbit_r30_c74 bl[74] br[74] wl[30] vdd gnd cell_6t
Xbit_r31_c74 bl[74] br[74] wl[31] vdd gnd cell_6t
Xbit_r32_c74 bl[74] br[74] wl[32] vdd gnd cell_6t
Xbit_r33_c74 bl[74] br[74] wl[33] vdd gnd cell_6t
Xbit_r34_c74 bl[74] br[74] wl[34] vdd gnd cell_6t
Xbit_r35_c74 bl[74] br[74] wl[35] vdd gnd cell_6t
Xbit_r36_c74 bl[74] br[74] wl[36] vdd gnd cell_6t
Xbit_r37_c74 bl[74] br[74] wl[37] vdd gnd cell_6t
Xbit_r38_c74 bl[74] br[74] wl[38] vdd gnd cell_6t
Xbit_r39_c74 bl[74] br[74] wl[39] vdd gnd cell_6t
Xbit_r40_c74 bl[74] br[74] wl[40] vdd gnd cell_6t
Xbit_r41_c74 bl[74] br[74] wl[41] vdd gnd cell_6t
Xbit_r42_c74 bl[74] br[74] wl[42] vdd gnd cell_6t
Xbit_r43_c74 bl[74] br[74] wl[43] vdd gnd cell_6t
Xbit_r44_c74 bl[74] br[74] wl[44] vdd gnd cell_6t
Xbit_r45_c74 bl[74] br[74] wl[45] vdd gnd cell_6t
Xbit_r46_c74 bl[74] br[74] wl[46] vdd gnd cell_6t
Xbit_r47_c74 bl[74] br[74] wl[47] vdd gnd cell_6t
Xbit_r48_c74 bl[74] br[74] wl[48] vdd gnd cell_6t
Xbit_r49_c74 bl[74] br[74] wl[49] vdd gnd cell_6t
Xbit_r50_c74 bl[74] br[74] wl[50] vdd gnd cell_6t
Xbit_r51_c74 bl[74] br[74] wl[51] vdd gnd cell_6t
Xbit_r52_c74 bl[74] br[74] wl[52] vdd gnd cell_6t
Xbit_r53_c74 bl[74] br[74] wl[53] vdd gnd cell_6t
Xbit_r54_c74 bl[74] br[74] wl[54] vdd gnd cell_6t
Xbit_r55_c74 bl[74] br[74] wl[55] vdd gnd cell_6t
Xbit_r56_c74 bl[74] br[74] wl[56] vdd gnd cell_6t
Xbit_r57_c74 bl[74] br[74] wl[57] vdd gnd cell_6t
Xbit_r58_c74 bl[74] br[74] wl[58] vdd gnd cell_6t
Xbit_r59_c74 bl[74] br[74] wl[59] vdd gnd cell_6t
Xbit_r60_c74 bl[74] br[74] wl[60] vdd gnd cell_6t
Xbit_r61_c74 bl[74] br[74] wl[61] vdd gnd cell_6t
Xbit_r62_c74 bl[74] br[74] wl[62] vdd gnd cell_6t
Xbit_r63_c74 bl[74] br[74] wl[63] vdd gnd cell_6t
Xbit_r64_c74 bl[74] br[74] wl[64] vdd gnd cell_6t
Xbit_r65_c74 bl[74] br[74] wl[65] vdd gnd cell_6t
Xbit_r66_c74 bl[74] br[74] wl[66] vdd gnd cell_6t
Xbit_r67_c74 bl[74] br[74] wl[67] vdd gnd cell_6t
Xbit_r68_c74 bl[74] br[74] wl[68] vdd gnd cell_6t
Xbit_r69_c74 bl[74] br[74] wl[69] vdd gnd cell_6t
Xbit_r70_c74 bl[74] br[74] wl[70] vdd gnd cell_6t
Xbit_r71_c74 bl[74] br[74] wl[71] vdd gnd cell_6t
Xbit_r72_c74 bl[74] br[74] wl[72] vdd gnd cell_6t
Xbit_r73_c74 bl[74] br[74] wl[73] vdd gnd cell_6t
Xbit_r74_c74 bl[74] br[74] wl[74] vdd gnd cell_6t
Xbit_r75_c74 bl[74] br[74] wl[75] vdd gnd cell_6t
Xbit_r76_c74 bl[74] br[74] wl[76] vdd gnd cell_6t
Xbit_r77_c74 bl[74] br[74] wl[77] vdd gnd cell_6t
Xbit_r78_c74 bl[74] br[74] wl[78] vdd gnd cell_6t
Xbit_r79_c74 bl[74] br[74] wl[79] vdd gnd cell_6t
Xbit_r80_c74 bl[74] br[74] wl[80] vdd gnd cell_6t
Xbit_r81_c74 bl[74] br[74] wl[81] vdd gnd cell_6t
Xbit_r82_c74 bl[74] br[74] wl[82] vdd gnd cell_6t
Xbit_r83_c74 bl[74] br[74] wl[83] vdd gnd cell_6t
Xbit_r84_c74 bl[74] br[74] wl[84] vdd gnd cell_6t
Xbit_r85_c74 bl[74] br[74] wl[85] vdd gnd cell_6t
Xbit_r86_c74 bl[74] br[74] wl[86] vdd gnd cell_6t
Xbit_r87_c74 bl[74] br[74] wl[87] vdd gnd cell_6t
Xbit_r88_c74 bl[74] br[74] wl[88] vdd gnd cell_6t
Xbit_r89_c74 bl[74] br[74] wl[89] vdd gnd cell_6t
Xbit_r90_c74 bl[74] br[74] wl[90] vdd gnd cell_6t
Xbit_r91_c74 bl[74] br[74] wl[91] vdd gnd cell_6t
Xbit_r92_c74 bl[74] br[74] wl[92] vdd gnd cell_6t
Xbit_r93_c74 bl[74] br[74] wl[93] vdd gnd cell_6t
Xbit_r94_c74 bl[74] br[74] wl[94] vdd gnd cell_6t
Xbit_r95_c74 bl[74] br[74] wl[95] vdd gnd cell_6t
Xbit_r96_c74 bl[74] br[74] wl[96] vdd gnd cell_6t
Xbit_r97_c74 bl[74] br[74] wl[97] vdd gnd cell_6t
Xbit_r98_c74 bl[74] br[74] wl[98] vdd gnd cell_6t
Xbit_r99_c74 bl[74] br[74] wl[99] vdd gnd cell_6t
Xbit_r100_c74 bl[74] br[74] wl[100] vdd gnd cell_6t
Xbit_r101_c74 bl[74] br[74] wl[101] vdd gnd cell_6t
Xbit_r102_c74 bl[74] br[74] wl[102] vdd gnd cell_6t
Xbit_r103_c74 bl[74] br[74] wl[103] vdd gnd cell_6t
Xbit_r104_c74 bl[74] br[74] wl[104] vdd gnd cell_6t
Xbit_r105_c74 bl[74] br[74] wl[105] vdd gnd cell_6t
Xbit_r106_c74 bl[74] br[74] wl[106] vdd gnd cell_6t
Xbit_r107_c74 bl[74] br[74] wl[107] vdd gnd cell_6t
Xbit_r108_c74 bl[74] br[74] wl[108] vdd gnd cell_6t
Xbit_r109_c74 bl[74] br[74] wl[109] vdd gnd cell_6t
Xbit_r110_c74 bl[74] br[74] wl[110] vdd gnd cell_6t
Xbit_r111_c74 bl[74] br[74] wl[111] vdd gnd cell_6t
Xbit_r112_c74 bl[74] br[74] wl[112] vdd gnd cell_6t
Xbit_r113_c74 bl[74] br[74] wl[113] vdd gnd cell_6t
Xbit_r114_c74 bl[74] br[74] wl[114] vdd gnd cell_6t
Xbit_r115_c74 bl[74] br[74] wl[115] vdd gnd cell_6t
Xbit_r116_c74 bl[74] br[74] wl[116] vdd gnd cell_6t
Xbit_r117_c74 bl[74] br[74] wl[117] vdd gnd cell_6t
Xbit_r118_c74 bl[74] br[74] wl[118] vdd gnd cell_6t
Xbit_r119_c74 bl[74] br[74] wl[119] vdd gnd cell_6t
Xbit_r120_c74 bl[74] br[74] wl[120] vdd gnd cell_6t
Xbit_r121_c74 bl[74] br[74] wl[121] vdd gnd cell_6t
Xbit_r122_c74 bl[74] br[74] wl[122] vdd gnd cell_6t
Xbit_r123_c74 bl[74] br[74] wl[123] vdd gnd cell_6t
Xbit_r124_c74 bl[74] br[74] wl[124] vdd gnd cell_6t
Xbit_r125_c74 bl[74] br[74] wl[125] vdd gnd cell_6t
Xbit_r126_c74 bl[74] br[74] wl[126] vdd gnd cell_6t
Xbit_r127_c74 bl[74] br[74] wl[127] vdd gnd cell_6t
Xbit_r128_c74 bl[74] br[74] wl[128] vdd gnd cell_6t
Xbit_r129_c74 bl[74] br[74] wl[129] vdd gnd cell_6t
Xbit_r130_c74 bl[74] br[74] wl[130] vdd gnd cell_6t
Xbit_r131_c74 bl[74] br[74] wl[131] vdd gnd cell_6t
Xbit_r132_c74 bl[74] br[74] wl[132] vdd gnd cell_6t
Xbit_r133_c74 bl[74] br[74] wl[133] vdd gnd cell_6t
Xbit_r134_c74 bl[74] br[74] wl[134] vdd gnd cell_6t
Xbit_r135_c74 bl[74] br[74] wl[135] vdd gnd cell_6t
Xbit_r136_c74 bl[74] br[74] wl[136] vdd gnd cell_6t
Xbit_r137_c74 bl[74] br[74] wl[137] vdd gnd cell_6t
Xbit_r138_c74 bl[74] br[74] wl[138] vdd gnd cell_6t
Xbit_r139_c74 bl[74] br[74] wl[139] vdd gnd cell_6t
Xbit_r140_c74 bl[74] br[74] wl[140] vdd gnd cell_6t
Xbit_r141_c74 bl[74] br[74] wl[141] vdd gnd cell_6t
Xbit_r142_c74 bl[74] br[74] wl[142] vdd gnd cell_6t
Xbit_r143_c74 bl[74] br[74] wl[143] vdd gnd cell_6t
Xbit_r144_c74 bl[74] br[74] wl[144] vdd gnd cell_6t
Xbit_r145_c74 bl[74] br[74] wl[145] vdd gnd cell_6t
Xbit_r146_c74 bl[74] br[74] wl[146] vdd gnd cell_6t
Xbit_r147_c74 bl[74] br[74] wl[147] vdd gnd cell_6t
Xbit_r148_c74 bl[74] br[74] wl[148] vdd gnd cell_6t
Xbit_r149_c74 bl[74] br[74] wl[149] vdd gnd cell_6t
Xbit_r150_c74 bl[74] br[74] wl[150] vdd gnd cell_6t
Xbit_r151_c74 bl[74] br[74] wl[151] vdd gnd cell_6t
Xbit_r152_c74 bl[74] br[74] wl[152] vdd gnd cell_6t
Xbit_r153_c74 bl[74] br[74] wl[153] vdd gnd cell_6t
Xbit_r154_c74 bl[74] br[74] wl[154] vdd gnd cell_6t
Xbit_r155_c74 bl[74] br[74] wl[155] vdd gnd cell_6t
Xbit_r156_c74 bl[74] br[74] wl[156] vdd gnd cell_6t
Xbit_r157_c74 bl[74] br[74] wl[157] vdd gnd cell_6t
Xbit_r158_c74 bl[74] br[74] wl[158] vdd gnd cell_6t
Xbit_r159_c74 bl[74] br[74] wl[159] vdd gnd cell_6t
Xbit_r160_c74 bl[74] br[74] wl[160] vdd gnd cell_6t
Xbit_r161_c74 bl[74] br[74] wl[161] vdd gnd cell_6t
Xbit_r162_c74 bl[74] br[74] wl[162] vdd gnd cell_6t
Xbit_r163_c74 bl[74] br[74] wl[163] vdd gnd cell_6t
Xbit_r164_c74 bl[74] br[74] wl[164] vdd gnd cell_6t
Xbit_r165_c74 bl[74] br[74] wl[165] vdd gnd cell_6t
Xbit_r166_c74 bl[74] br[74] wl[166] vdd gnd cell_6t
Xbit_r167_c74 bl[74] br[74] wl[167] vdd gnd cell_6t
Xbit_r168_c74 bl[74] br[74] wl[168] vdd gnd cell_6t
Xbit_r169_c74 bl[74] br[74] wl[169] vdd gnd cell_6t
Xbit_r170_c74 bl[74] br[74] wl[170] vdd gnd cell_6t
Xbit_r171_c74 bl[74] br[74] wl[171] vdd gnd cell_6t
Xbit_r172_c74 bl[74] br[74] wl[172] vdd gnd cell_6t
Xbit_r173_c74 bl[74] br[74] wl[173] vdd gnd cell_6t
Xbit_r174_c74 bl[74] br[74] wl[174] vdd gnd cell_6t
Xbit_r175_c74 bl[74] br[74] wl[175] vdd gnd cell_6t
Xbit_r176_c74 bl[74] br[74] wl[176] vdd gnd cell_6t
Xbit_r177_c74 bl[74] br[74] wl[177] vdd gnd cell_6t
Xbit_r178_c74 bl[74] br[74] wl[178] vdd gnd cell_6t
Xbit_r179_c74 bl[74] br[74] wl[179] vdd gnd cell_6t
Xbit_r180_c74 bl[74] br[74] wl[180] vdd gnd cell_6t
Xbit_r181_c74 bl[74] br[74] wl[181] vdd gnd cell_6t
Xbit_r182_c74 bl[74] br[74] wl[182] vdd gnd cell_6t
Xbit_r183_c74 bl[74] br[74] wl[183] vdd gnd cell_6t
Xbit_r184_c74 bl[74] br[74] wl[184] vdd gnd cell_6t
Xbit_r185_c74 bl[74] br[74] wl[185] vdd gnd cell_6t
Xbit_r186_c74 bl[74] br[74] wl[186] vdd gnd cell_6t
Xbit_r187_c74 bl[74] br[74] wl[187] vdd gnd cell_6t
Xbit_r188_c74 bl[74] br[74] wl[188] vdd gnd cell_6t
Xbit_r189_c74 bl[74] br[74] wl[189] vdd gnd cell_6t
Xbit_r190_c74 bl[74] br[74] wl[190] vdd gnd cell_6t
Xbit_r191_c74 bl[74] br[74] wl[191] vdd gnd cell_6t
Xbit_r192_c74 bl[74] br[74] wl[192] vdd gnd cell_6t
Xbit_r193_c74 bl[74] br[74] wl[193] vdd gnd cell_6t
Xbit_r194_c74 bl[74] br[74] wl[194] vdd gnd cell_6t
Xbit_r195_c74 bl[74] br[74] wl[195] vdd gnd cell_6t
Xbit_r196_c74 bl[74] br[74] wl[196] vdd gnd cell_6t
Xbit_r197_c74 bl[74] br[74] wl[197] vdd gnd cell_6t
Xbit_r198_c74 bl[74] br[74] wl[198] vdd gnd cell_6t
Xbit_r199_c74 bl[74] br[74] wl[199] vdd gnd cell_6t
Xbit_r200_c74 bl[74] br[74] wl[200] vdd gnd cell_6t
Xbit_r201_c74 bl[74] br[74] wl[201] vdd gnd cell_6t
Xbit_r202_c74 bl[74] br[74] wl[202] vdd gnd cell_6t
Xbit_r203_c74 bl[74] br[74] wl[203] vdd gnd cell_6t
Xbit_r204_c74 bl[74] br[74] wl[204] vdd gnd cell_6t
Xbit_r205_c74 bl[74] br[74] wl[205] vdd gnd cell_6t
Xbit_r206_c74 bl[74] br[74] wl[206] vdd gnd cell_6t
Xbit_r207_c74 bl[74] br[74] wl[207] vdd gnd cell_6t
Xbit_r208_c74 bl[74] br[74] wl[208] vdd gnd cell_6t
Xbit_r209_c74 bl[74] br[74] wl[209] vdd gnd cell_6t
Xbit_r210_c74 bl[74] br[74] wl[210] vdd gnd cell_6t
Xbit_r211_c74 bl[74] br[74] wl[211] vdd gnd cell_6t
Xbit_r212_c74 bl[74] br[74] wl[212] vdd gnd cell_6t
Xbit_r213_c74 bl[74] br[74] wl[213] vdd gnd cell_6t
Xbit_r214_c74 bl[74] br[74] wl[214] vdd gnd cell_6t
Xbit_r215_c74 bl[74] br[74] wl[215] vdd gnd cell_6t
Xbit_r216_c74 bl[74] br[74] wl[216] vdd gnd cell_6t
Xbit_r217_c74 bl[74] br[74] wl[217] vdd gnd cell_6t
Xbit_r218_c74 bl[74] br[74] wl[218] vdd gnd cell_6t
Xbit_r219_c74 bl[74] br[74] wl[219] vdd gnd cell_6t
Xbit_r220_c74 bl[74] br[74] wl[220] vdd gnd cell_6t
Xbit_r221_c74 bl[74] br[74] wl[221] vdd gnd cell_6t
Xbit_r222_c74 bl[74] br[74] wl[222] vdd gnd cell_6t
Xbit_r223_c74 bl[74] br[74] wl[223] vdd gnd cell_6t
Xbit_r224_c74 bl[74] br[74] wl[224] vdd gnd cell_6t
Xbit_r225_c74 bl[74] br[74] wl[225] vdd gnd cell_6t
Xbit_r226_c74 bl[74] br[74] wl[226] vdd gnd cell_6t
Xbit_r227_c74 bl[74] br[74] wl[227] vdd gnd cell_6t
Xbit_r228_c74 bl[74] br[74] wl[228] vdd gnd cell_6t
Xbit_r229_c74 bl[74] br[74] wl[229] vdd gnd cell_6t
Xbit_r230_c74 bl[74] br[74] wl[230] vdd gnd cell_6t
Xbit_r231_c74 bl[74] br[74] wl[231] vdd gnd cell_6t
Xbit_r232_c74 bl[74] br[74] wl[232] vdd gnd cell_6t
Xbit_r233_c74 bl[74] br[74] wl[233] vdd gnd cell_6t
Xbit_r234_c74 bl[74] br[74] wl[234] vdd gnd cell_6t
Xbit_r235_c74 bl[74] br[74] wl[235] vdd gnd cell_6t
Xbit_r236_c74 bl[74] br[74] wl[236] vdd gnd cell_6t
Xbit_r237_c74 bl[74] br[74] wl[237] vdd gnd cell_6t
Xbit_r238_c74 bl[74] br[74] wl[238] vdd gnd cell_6t
Xbit_r239_c74 bl[74] br[74] wl[239] vdd gnd cell_6t
Xbit_r240_c74 bl[74] br[74] wl[240] vdd gnd cell_6t
Xbit_r241_c74 bl[74] br[74] wl[241] vdd gnd cell_6t
Xbit_r242_c74 bl[74] br[74] wl[242] vdd gnd cell_6t
Xbit_r243_c74 bl[74] br[74] wl[243] vdd gnd cell_6t
Xbit_r244_c74 bl[74] br[74] wl[244] vdd gnd cell_6t
Xbit_r245_c74 bl[74] br[74] wl[245] vdd gnd cell_6t
Xbit_r246_c74 bl[74] br[74] wl[246] vdd gnd cell_6t
Xbit_r247_c74 bl[74] br[74] wl[247] vdd gnd cell_6t
Xbit_r248_c74 bl[74] br[74] wl[248] vdd gnd cell_6t
Xbit_r249_c74 bl[74] br[74] wl[249] vdd gnd cell_6t
Xbit_r250_c74 bl[74] br[74] wl[250] vdd gnd cell_6t
Xbit_r251_c74 bl[74] br[74] wl[251] vdd gnd cell_6t
Xbit_r252_c74 bl[74] br[74] wl[252] vdd gnd cell_6t
Xbit_r253_c74 bl[74] br[74] wl[253] vdd gnd cell_6t
Xbit_r254_c74 bl[74] br[74] wl[254] vdd gnd cell_6t
Xbit_r255_c74 bl[74] br[74] wl[255] vdd gnd cell_6t
Xbit_r256_c74 bl[74] br[74] wl[256] vdd gnd cell_6t
Xbit_r257_c74 bl[74] br[74] wl[257] vdd gnd cell_6t
Xbit_r258_c74 bl[74] br[74] wl[258] vdd gnd cell_6t
Xbit_r259_c74 bl[74] br[74] wl[259] vdd gnd cell_6t
Xbit_r260_c74 bl[74] br[74] wl[260] vdd gnd cell_6t
Xbit_r261_c74 bl[74] br[74] wl[261] vdd gnd cell_6t
Xbit_r262_c74 bl[74] br[74] wl[262] vdd gnd cell_6t
Xbit_r263_c74 bl[74] br[74] wl[263] vdd gnd cell_6t
Xbit_r264_c74 bl[74] br[74] wl[264] vdd gnd cell_6t
Xbit_r265_c74 bl[74] br[74] wl[265] vdd gnd cell_6t
Xbit_r266_c74 bl[74] br[74] wl[266] vdd gnd cell_6t
Xbit_r267_c74 bl[74] br[74] wl[267] vdd gnd cell_6t
Xbit_r268_c74 bl[74] br[74] wl[268] vdd gnd cell_6t
Xbit_r269_c74 bl[74] br[74] wl[269] vdd gnd cell_6t
Xbit_r270_c74 bl[74] br[74] wl[270] vdd gnd cell_6t
Xbit_r271_c74 bl[74] br[74] wl[271] vdd gnd cell_6t
Xbit_r272_c74 bl[74] br[74] wl[272] vdd gnd cell_6t
Xbit_r273_c74 bl[74] br[74] wl[273] vdd gnd cell_6t
Xbit_r274_c74 bl[74] br[74] wl[274] vdd gnd cell_6t
Xbit_r275_c74 bl[74] br[74] wl[275] vdd gnd cell_6t
Xbit_r276_c74 bl[74] br[74] wl[276] vdd gnd cell_6t
Xbit_r277_c74 bl[74] br[74] wl[277] vdd gnd cell_6t
Xbit_r278_c74 bl[74] br[74] wl[278] vdd gnd cell_6t
Xbit_r279_c74 bl[74] br[74] wl[279] vdd gnd cell_6t
Xbit_r280_c74 bl[74] br[74] wl[280] vdd gnd cell_6t
Xbit_r281_c74 bl[74] br[74] wl[281] vdd gnd cell_6t
Xbit_r282_c74 bl[74] br[74] wl[282] vdd gnd cell_6t
Xbit_r283_c74 bl[74] br[74] wl[283] vdd gnd cell_6t
Xbit_r284_c74 bl[74] br[74] wl[284] vdd gnd cell_6t
Xbit_r285_c74 bl[74] br[74] wl[285] vdd gnd cell_6t
Xbit_r286_c74 bl[74] br[74] wl[286] vdd gnd cell_6t
Xbit_r287_c74 bl[74] br[74] wl[287] vdd gnd cell_6t
Xbit_r288_c74 bl[74] br[74] wl[288] vdd gnd cell_6t
Xbit_r289_c74 bl[74] br[74] wl[289] vdd gnd cell_6t
Xbit_r290_c74 bl[74] br[74] wl[290] vdd gnd cell_6t
Xbit_r291_c74 bl[74] br[74] wl[291] vdd gnd cell_6t
Xbit_r292_c74 bl[74] br[74] wl[292] vdd gnd cell_6t
Xbit_r293_c74 bl[74] br[74] wl[293] vdd gnd cell_6t
Xbit_r294_c74 bl[74] br[74] wl[294] vdd gnd cell_6t
Xbit_r295_c74 bl[74] br[74] wl[295] vdd gnd cell_6t
Xbit_r296_c74 bl[74] br[74] wl[296] vdd gnd cell_6t
Xbit_r297_c74 bl[74] br[74] wl[297] vdd gnd cell_6t
Xbit_r298_c74 bl[74] br[74] wl[298] vdd gnd cell_6t
Xbit_r299_c74 bl[74] br[74] wl[299] vdd gnd cell_6t
Xbit_r300_c74 bl[74] br[74] wl[300] vdd gnd cell_6t
Xbit_r301_c74 bl[74] br[74] wl[301] vdd gnd cell_6t
Xbit_r302_c74 bl[74] br[74] wl[302] vdd gnd cell_6t
Xbit_r303_c74 bl[74] br[74] wl[303] vdd gnd cell_6t
Xbit_r304_c74 bl[74] br[74] wl[304] vdd gnd cell_6t
Xbit_r305_c74 bl[74] br[74] wl[305] vdd gnd cell_6t
Xbit_r306_c74 bl[74] br[74] wl[306] vdd gnd cell_6t
Xbit_r307_c74 bl[74] br[74] wl[307] vdd gnd cell_6t
Xbit_r308_c74 bl[74] br[74] wl[308] vdd gnd cell_6t
Xbit_r309_c74 bl[74] br[74] wl[309] vdd gnd cell_6t
Xbit_r310_c74 bl[74] br[74] wl[310] vdd gnd cell_6t
Xbit_r311_c74 bl[74] br[74] wl[311] vdd gnd cell_6t
Xbit_r312_c74 bl[74] br[74] wl[312] vdd gnd cell_6t
Xbit_r313_c74 bl[74] br[74] wl[313] vdd gnd cell_6t
Xbit_r314_c74 bl[74] br[74] wl[314] vdd gnd cell_6t
Xbit_r315_c74 bl[74] br[74] wl[315] vdd gnd cell_6t
Xbit_r316_c74 bl[74] br[74] wl[316] vdd gnd cell_6t
Xbit_r317_c74 bl[74] br[74] wl[317] vdd gnd cell_6t
Xbit_r318_c74 bl[74] br[74] wl[318] vdd gnd cell_6t
Xbit_r319_c74 bl[74] br[74] wl[319] vdd gnd cell_6t
Xbit_r320_c74 bl[74] br[74] wl[320] vdd gnd cell_6t
Xbit_r321_c74 bl[74] br[74] wl[321] vdd gnd cell_6t
Xbit_r322_c74 bl[74] br[74] wl[322] vdd gnd cell_6t
Xbit_r323_c74 bl[74] br[74] wl[323] vdd gnd cell_6t
Xbit_r324_c74 bl[74] br[74] wl[324] vdd gnd cell_6t
Xbit_r325_c74 bl[74] br[74] wl[325] vdd gnd cell_6t
Xbit_r326_c74 bl[74] br[74] wl[326] vdd gnd cell_6t
Xbit_r327_c74 bl[74] br[74] wl[327] vdd gnd cell_6t
Xbit_r328_c74 bl[74] br[74] wl[328] vdd gnd cell_6t
Xbit_r329_c74 bl[74] br[74] wl[329] vdd gnd cell_6t
Xbit_r330_c74 bl[74] br[74] wl[330] vdd gnd cell_6t
Xbit_r331_c74 bl[74] br[74] wl[331] vdd gnd cell_6t
Xbit_r332_c74 bl[74] br[74] wl[332] vdd gnd cell_6t
Xbit_r333_c74 bl[74] br[74] wl[333] vdd gnd cell_6t
Xbit_r334_c74 bl[74] br[74] wl[334] vdd gnd cell_6t
Xbit_r335_c74 bl[74] br[74] wl[335] vdd gnd cell_6t
Xbit_r336_c74 bl[74] br[74] wl[336] vdd gnd cell_6t
Xbit_r337_c74 bl[74] br[74] wl[337] vdd gnd cell_6t
Xbit_r338_c74 bl[74] br[74] wl[338] vdd gnd cell_6t
Xbit_r339_c74 bl[74] br[74] wl[339] vdd gnd cell_6t
Xbit_r340_c74 bl[74] br[74] wl[340] vdd gnd cell_6t
Xbit_r341_c74 bl[74] br[74] wl[341] vdd gnd cell_6t
Xbit_r342_c74 bl[74] br[74] wl[342] vdd gnd cell_6t
Xbit_r343_c74 bl[74] br[74] wl[343] vdd gnd cell_6t
Xbit_r344_c74 bl[74] br[74] wl[344] vdd gnd cell_6t
Xbit_r345_c74 bl[74] br[74] wl[345] vdd gnd cell_6t
Xbit_r346_c74 bl[74] br[74] wl[346] vdd gnd cell_6t
Xbit_r347_c74 bl[74] br[74] wl[347] vdd gnd cell_6t
Xbit_r348_c74 bl[74] br[74] wl[348] vdd gnd cell_6t
Xbit_r349_c74 bl[74] br[74] wl[349] vdd gnd cell_6t
Xbit_r350_c74 bl[74] br[74] wl[350] vdd gnd cell_6t
Xbit_r351_c74 bl[74] br[74] wl[351] vdd gnd cell_6t
Xbit_r352_c74 bl[74] br[74] wl[352] vdd gnd cell_6t
Xbit_r353_c74 bl[74] br[74] wl[353] vdd gnd cell_6t
Xbit_r354_c74 bl[74] br[74] wl[354] vdd gnd cell_6t
Xbit_r355_c74 bl[74] br[74] wl[355] vdd gnd cell_6t
Xbit_r356_c74 bl[74] br[74] wl[356] vdd gnd cell_6t
Xbit_r357_c74 bl[74] br[74] wl[357] vdd gnd cell_6t
Xbit_r358_c74 bl[74] br[74] wl[358] vdd gnd cell_6t
Xbit_r359_c74 bl[74] br[74] wl[359] vdd gnd cell_6t
Xbit_r360_c74 bl[74] br[74] wl[360] vdd gnd cell_6t
Xbit_r361_c74 bl[74] br[74] wl[361] vdd gnd cell_6t
Xbit_r362_c74 bl[74] br[74] wl[362] vdd gnd cell_6t
Xbit_r363_c74 bl[74] br[74] wl[363] vdd gnd cell_6t
Xbit_r364_c74 bl[74] br[74] wl[364] vdd gnd cell_6t
Xbit_r365_c74 bl[74] br[74] wl[365] vdd gnd cell_6t
Xbit_r366_c74 bl[74] br[74] wl[366] vdd gnd cell_6t
Xbit_r367_c74 bl[74] br[74] wl[367] vdd gnd cell_6t
Xbit_r368_c74 bl[74] br[74] wl[368] vdd gnd cell_6t
Xbit_r369_c74 bl[74] br[74] wl[369] vdd gnd cell_6t
Xbit_r370_c74 bl[74] br[74] wl[370] vdd gnd cell_6t
Xbit_r371_c74 bl[74] br[74] wl[371] vdd gnd cell_6t
Xbit_r372_c74 bl[74] br[74] wl[372] vdd gnd cell_6t
Xbit_r373_c74 bl[74] br[74] wl[373] vdd gnd cell_6t
Xbit_r374_c74 bl[74] br[74] wl[374] vdd gnd cell_6t
Xbit_r375_c74 bl[74] br[74] wl[375] vdd gnd cell_6t
Xbit_r376_c74 bl[74] br[74] wl[376] vdd gnd cell_6t
Xbit_r377_c74 bl[74] br[74] wl[377] vdd gnd cell_6t
Xbit_r378_c74 bl[74] br[74] wl[378] vdd gnd cell_6t
Xbit_r379_c74 bl[74] br[74] wl[379] vdd gnd cell_6t
Xbit_r380_c74 bl[74] br[74] wl[380] vdd gnd cell_6t
Xbit_r381_c74 bl[74] br[74] wl[381] vdd gnd cell_6t
Xbit_r382_c74 bl[74] br[74] wl[382] vdd gnd cell_6t
Xbit_r383_c74 bl[74] br[74] wl[383] vdd gnd cell_6t
Xbit_r384_c74 bl[74] br[74] wl[384] vdd gnd cell_6t
Xbit_r385_c74 bl[74] br[74] wl[385] vdd gnd cell_6t
Xbit_r386_c74 bl[74] br[74] wl[386] vdd gnd cell_6t
Xbit_r387_c74 bl[74] br[74] wl[387] vdd gnd cell_6t
Xbit_r388_c74 bl[74] br[74] wl[388] vdd gnd cell_6t
Xbit_r389_c74 bl[74] br[74] wl[389] vdd gnd cell_6t
Xbit_r390_c74 bl[74] br[74] wl[390] vdd gnd cell_6t
Xbit_r391_c74 bl[74] br[74] wl[391] vdd gnd cell_6t
Xbit_r392_c74 bl[74] br[74] wl[392] vdd gnd cell_6t
Xbit_r393_c74 bl[74] br[74] wl[393] vdd gnd cell_6t
Xbit_r394_c74 bl[74] br[74] wl[394] vdd gnd cell_6t
Xbit_r395_c74 bl[74] br[74] wl[395] vdd gnd cell_6t
Xbit_r396_c74 bl[74] br[74] wl[396] vdd gnd cell_6t
Xbit_r397_c74 bl[74] br[74] wl[397] vdd gnd cell_6t
Xbit_r398_c74 bl[74] br[74] wl[398] vdd gnd cell_6t
Xbit_r399_c74 bl[74] br[74] wl[399] vdd gnd cell_6t
Xbit_r400_c74 bl[74] br[74] wl[400] vdd gnd cell_6t
Xbit_r401_c74 bl[74] br[74] wl[401] vdd gnd cell_6t
Xbit_r402_c74 bl[74] br[74] wl[402] vdd gnd cell_6t
Xbit_r403_c74 bl[74] br[74] wl[403] vdd gnd cell_6t
Xbit_r404_c74 bl[74] br[74] wl[404] vdd gnd cell_6t
Xbit_r405_c74 bl[74] br[74] wl[405] vdd gnd cell_6t
Xbit_r406_c74 bl[74] br[74] wl[406] vdd gnd cell_6t
Xbit_r407_c74 bl[74] br[74] wl[407] vdd gnd cell_6t
Xbit_r408_c74 bl[74] br[74] wl[408] vdd gnd cell_6t
Xbit_r409_c74 bl[74] br[74] wl[409] vdd gnd cell_6t
Xbit_r410_c74 bl[74] br[74] wl[410] vdd gnd cell_6t
Xbit_r411_c74 bl[74] br[74] wl[411] vdd gnd cell_6t
Xbit_r412_c74 bl[74] br[74] wl[412] vdd gnd cell_6t
Xbit_r413_c74 bl[74] br[74] wl[413] vdd gnd cell_6t
Xbit_r414_c74 bl[74] br[74] wl[414] vdd gnd cell_6t
Xbit_r415_c74 bl[74] br[74] wl[415] vdd gnd cell_6t
Xbit_r416_c74 bl[74] br[74] wl[416] vdd gnd cell_6t
Xbit_r417_c74 bl[74] br[74] wl[417] vdd gnd cell_6t
Xbit_r418_c74 bl[74] br[74] wl[418] vdd gnd cell_6t
Xbit_r419_c74 bl[74] br[74] wl[419] vdd gnd cell_6t
Xbit_r420_c74 bl[74] br[74] wl[420] vdd gnd cell_6t
Xbit_r421_c74 bl[74] br[74] wl[421] vdd gnd cell_6t
Xbit_r422_c74 bl[74] br[74] wl[422] vdd gnd cell_6t
Xbit_r423_c74 bl[74] br[74] wl[423] vdd gnd cell_6t
Xbit_r424_c74 bl[74] br[74] wl[424] vdd gnd cell_6t
Xbit_r425_c74 bl[74] br[74] wl[425] vdd gnd cell_6t
Xbit_r426_c74 bl[74] br[74] wl[426] vdd gnd cell_6t
Xbit_r427_c74 bl[74] br[74] wl[427] vdd gnd cell_6t
Xbit_r428_c74 bl[74] br[74] wl[428] vdd gnd cell_6t
Xbit_r429_c74 bl[74] br[74] wl[429] vdd gnd cell_6t
Xbit_r430_c74 bl[74] br[74] wl[430] vdd gnd cell_6t
Xbit_r431_c74 bl[74] br[74] wl[431] vdd gnd cell_6t
Xbit_r432_c74 bl[74] br[74] wl[432] vdd gnd cell_6t
Xbit_r433_c74 bl[74] br[74] wl[433] vdd gnd cell_6t
Xbit_r434_c74 bl[74] br[74] wl[434] vdd gnd cell_6t
Xbit_r435_c74 bl[74] br[74] wl[435] vdd gnd cell_6t
Xbit_r436_c74 bl[74] br[74] wl[436] vdd gnd cell_6t
Xbit_r437_c74 bl[74] br[74] wl[437] vdd gnd cell_6t
Xbit_r438_c74 bl[74] br[74] wl[438] vdd gnd cell_6t
Xbit_r439_c74 bl[74] br[74] wl[439] vdd gnd cell_6t
Xbit_r440_c74 bl[74] br[74] wl[440] vdd gnd cell_6t
Xbit_r441_c74 bl[74] br[74] wl[441] vdd gnd cell_6t
Xbit_r442_c74 bl[74] br[74] wl[442] vdd gnd cell_6t
Xbit_r443_c74 bl[74] br[74] wl[443] vdd gnd cell_6t
Xbit_r444_c74 bl[74] br[74] wl[444] vdd gnd cell_6t
Xbit_r445_c74 bl[74] br[74] wl[445] vdd gnd cell_6t
Xbit_r446_c74 bl[74] br[74] wl[446] vdd gnd cell_6t
Xbit_r447_c74 bl[74] br[74] wl[447] vdd gnd cell_6t
Xbit_r448_c74 bl[74] br[74] wl[448] vdd gnd cell_6t
Xbit_r449_c74 bl[74] br[74] wl[449] vdd gnd cell_6t
Xbit_r450_c74 bl[74] br[74] wl[450] vdd gnd cell_6t
Xbit_r451_c74 bl[74] br[74] wl[451] vdd gnd cell_6t
Xbit_r452_c74 bl[74] br[74] wl[452] vdd gnd cell_6t
Xbit_r453_c74 bl[74] br[74] wl[453] vdd gnd cell_6t
Xbit_r454_c74 bl[74] br[74] wl[454] vdd gnd cell_6t
Xbit_r455_c74 bl[74] br[74] wl[455] vdd gnd cell_6t
Xbit_r456_c74 bl[74] br[74] wl[456] vdd gnd cell_6t
Xbit_r457_c74 bl[74] br[74] wl[457] vdd gnd cell_6t
Xbit_r458_c74 bl[74] br[74] wl[458] vdd gnd cell_6t
Xbit_r459_c74 bl[74] br[74] wl[459] vdd gnd cell_6t
Xbit_r460_c74 bl[74] br[74] wl[460] vdd gnd cell_6t
Xbit_r461_c74 bl[74] br[74] wl[461] vdd gnd cell_6t
Xbit_r462_c74 bl[74] br[74] wl[462] vdd gnd cell_6t
Xbit_r463_c74 bl[74] br[74] wl[463] vdd gnd cell_6t
Xbit_r464_c74 bl[74] br[74] wl[464] vdd gnd cell_6t
Xbit_r465_c74 bl[74] br[74] wl[465] vdd gnd cell_6t
Xbit_r466_c74 bl[74] br[74] wl[466] vdd gnd cell_6t
Xbit_r467_c74 bl[74] br[74] wl[467] vdd gnd cell_6t
Xbit_r468_c74 bl[74] br[74] wl[468] vdd gnd cell_6t
Xbit_r469_c74 bl[74] br[74] wl[469] vdd gnd cell_6t
Xbit_r470_c74 bl[74] br[74] wl[470] vdd gnd cell_6t
Xbit_r471_c74 bl[74] br[74] wl[471] vdd gnd cell_6t
Xbit_r472_c74 bl[74] br[74] wl[472] vdd gnd cell_6t
Xbit_r473_c74 bl[74] br[74] wl[473] vdd gnd cell_6t
Xbit_r474_c74 bl[74] br[74] wl[474] vdd gnd cell_6t
Xbit_r475_c74 bl[74] br[74] wl[475] vdd gnd cell_6t
Xbit_r476_c74 bl[74] br[74] wl[476] vdd gnd cell_6t
Xbit_r477_c74 bl[74] br[74] wl[477] vdd gnd cell_6t
Xbit_r478_c74 bl[74] br[74] wl[478] vdd gnd cell_6t
Xbit_r479_c74 bl[74] br[74] wl[479] vdd gnd cell_6t
Xbit_r480_c74 bl[74] br[74] wl[480] vdd gnd cell_6t
Xbit_r481_c74 bl[74] br[74] wl[481] vdd gnd cell_6t
Xbit_r482_c74 bl[74] br[74] wl[482] vdd gnd cell_6t
Xbit_r483_c74 bl[74] br[74] wl[483] vdd gnd cell_6t
Xbit_r484_c74 bl[74] br[74] wl[484] vdd gnd cell_6t
Xbit_r485_c74 bl[74] br[74] wl[485] vdd gnd cell_6t
Xbit_r486_c74 bl[74] br[74] wl[486] vdd gnd cell_6t
Xbit_r487_c74 bl[74] br[74] wl[487] vdd gnd cell_6t
Xbit_r488_c74 bl[74] br[74] wl[488] vdd gnd cell_6t
Xbit_r489_c74 bl[74] br[74] wl[489] vdd gnd cell_6t
Xbit_r490_c74 bl[74] br[74] wl[490] vdd gnd cell_6t
Xbit_r491_c74 bl[74] br[74] wl[491] vdd gnd cell_6t
Xbit_r492_c74 bl[74] br[74] wl[492] vdd gnd cell_6t
Xbit_r493_c74 bl[74] br[74] wl[493] vdd gnd cell_6t
Xbit_r494_c74 bl[74] br[74] wl[494] vdd gnd cell_6t
Xbit_r495_c74 bl[74] br[74] wl[495] vdd gnd cell_6t
Xbit_r496_c74 bl[74] br[74] wl[496] vdd gnd cell_6t
Xbit_r497_c74 bl[74] br[74] wl[497] vdd gnd cell_6t
Xbit_r498_c74 bl[74] br[74] wl[498] vdd gnd cell_6t
Xbit_r499_c74 bl[74] br[74] wl[499] vdd gnd cell_6t
Xbit_r500_c74 bl[74] br[74] wl[500] vdd gnd cell_6t
Xbit_r501_c74 bl[74] br[74] wl[501] vdd gnd cell_6t
Xbit_r502_c74 bl[74] br[74] wl[502] vdd gnd cell_6t
Xbit_r503_c74 bl[74] br[74] wl[503] vdd gnd cell_6t
Xbit_r504_c74 bl[74] br[74] wl[504] vdd gnd cell_6t
Xbit_r505_c74 bl[74] br[74] wl[505] vdd gnd cell_6t
Xbit_r506_c74 bl[74] br[74] wl[506] vdd gnd cell_6t
Xbit_r507_c74 bl[74] br[74] wl[507] vdd gnd cell_6t
Xbit_r508_c74 bl[74] br[74] wl[508] vdd gnd cell_6t
Xbit_r509_c74 bl[74] br[74] wl[509] vdd gnd cell_6t
Xbit_r510_c74 bl[74] br[74] wl[510] vdd gnd cell_6t
Xbit_r511_c74 bl[74] br[74] wl[511] vdd gnd cell_6t
Xbit_r0_c75 bl[75] br[75] wl[0] vdd gnd cell_6t
Xbit_r1_c75 bl[75] br[75] wl[1] vdd gnd cell_6t
Xbit_r2_c75 bl[75] br[75] wl[2] vdd gnd cell_6t
Xbit_r3_c75 bl[75] br[75] wl[3] vdd gnd cell_6t
Xbit_r4_c75 bl[75] br[75] wl[4] vdd gnd cell_6t
Xbit_r5_c75 bl[75] br[75] wl[5] vdd gnd cell_6t
Xbit_r6_c75 bl[75] br[75] wl[6] vdd gnd cell_6t
Xbit_r7_c75 bl[75] br[75] wl[7] vdd gnd cell_6t
Xbit_r8_c75 bl[75] br[75] wl[8] vdd gnd cell_6t
Xbit_r9_c75 bl[75] br[75] wl[9] vdd gnd cell_6t
Xbit_r10_c75 bl[75] br[75] wl[10] vdd gnd cell_6t
Xbit_r11_c75 bl[75] br[75] wl[11] vdd gnd cell_6t
Xbit_r12_c75 bl[75] br[75] wl[12] vdd gnd cell_6t
Xbit_r13_c75 bl[75] br[75] wl[13] vdd gnd cell_6t
Xbit_r14_c75 bl[75] br[75] wl[14] vdd gnd cell_6t
Xbit_r15_c75 bl[75] br[75] wl[15] vdd gnd cell_6t
Xbit_r16_c75 bl[75] br[75] wl[16] vdd gnd cell_6t
Xbit_r17_c75 bl[75] br[75] wl[17] vdd gnd cell_6t
Xbit_r18_c75 bl[75] br[75] wl[18] vdd gnd cell_6t
Xbit_r19_c75 bl[75] br[75] wl[19] vdd gnd cell_6t
Xbit_r20_c75 bl[75] br[75] wl[20] vdd gnd cell_6t
Xbit_r21_c75 bl[75] br[75] wl[21] vdd gnd cell_6t
Xbit_r22_c75 bl[75] br[75] wl[22] vdd gnd cell_6t
Xbit_r23_c75 bl[75] br[75] wl[23] vdd gnd cell_6t
Xbit_r24_c75 bl[75] br[75] wl[24] vdd gnd cell_6t
Xbit_r25_c75 bl[75] br[75] wl[25] vdd gnd cell_6t
Xbit_r26_c75 bl[75] br[75] wl[26] vdd gnd cell_6t
Xbit_r27_c75 bl[75] br[75] wl[27] vdd gnd cell_6t
Xbit_r28_c75 bl[75] br[75] wl[28] vdd gnd cell_6t
Xbit_r29_c75 bl[75] br[75] wl[29] vdd gnd cell_6t
Xbit_r30_c75 bl[75] br[75] wl[30] vdd gnd cell_6t
Xbit_r31_c75 bl[75] br[75] wl[31] vdd gnd cell_6t
Xbit_r32_c75 bl[75] br[75] wl[32] vdd gnd cell_6t
Xbit_r33_c75 bl[75] br[75] wl[33] vdd gnd cell_6t
Xbit_r34_c75 bl[75] br[75] wl[34] vdd gnd cell_6t
Xbit_r35_c75 bl[75] br[75] wl[35] vdd gnd cell_6t
Xbit_r36_c75 bl[75] br[75] wl[36] vdd gnd cell_6t
Xbit_r37_c75 bl[75] br[75] wl[37] vdd gnd cell_6t
Xbit_r38_c75 bl[75] br[75] wl[38] vdd gnd cell_6t
Xbit_r39_c75 bl[75] br[75] wl[39] vdd gnd cell_6t
Xbit_r40_c75 bl[75] br[75] wl[40] vdd gnd cell_6t
Xbit_r41_c75 bl[75] br[75] wl[41] vdd gnd cell_6t
Xbit_r42_c75 bl[75] br[75] wl[42] vdd gnd cell_6t
Xbit_r43_c75 bl[75] br[75] wl[43] vdd gnd cell_6t
Xbit_r44_c75 bl[75] br[75] wl[44] vdd gnd cell_6t
Xbit_r45_c75 bl[75] br[75] wl[45] vdd gnd cell_6t
Xbit_r46_c75 bl[75] br[75] wl[46] vdd gnd cell_6t
Xbit_r47_c75 bl[75] br[75] wl[47] vdd gnd cell_6t
Xbit_r48_c75 bl[75] br[75] wl[48] vdd gnd cell_6t
Xbit_r49_c75 bl[75] br[75] wl[49] vdd gnd cell_6t
Xbit_r50_c75 bl[75] br[75] wl[50] vdd gnd cell_6t
Xbit_r51_c75 bl[75] br[75] wl[51] vdd gnd cell_6t
Xbit_r52_c75 bl[75] br[75] wl[52] vdd gnd cell_6t
Xbit_r53_c75 bl[75] br[75] wl[53] vdd gnd cell_6t
Xbit_r54_c75 bl[75] br[75] wl[54] vdd gnd cell_6t
Xbit_r55_c75 bl[75] br[75] wl[55] vdd gnd cell_6t
Xbit_r56_c75 bl[75] br[75] wl[56] vdd gnd cell_6t
Xbit_r57_c75 bl[75] br[75] wl[57] vdd gnd cell_6t
Xbit_r58_c75 bl[75] br[75] wl[58] vdd gnd cell_6t
Xbit_r59_c75 bl[75] br[75] wl[59] vdd gnd cell_6t
Xbit_r60_c75 bl[75] br[75] wl[60] vdd gnd cell_6t
Xbit_r61_c75 bl[75] br[75] wl[61] vdd gnd cell_6t
Xbit_r62_c75 bl[75] br[75] wl[62] vdd gnd cell_6t
Xbit_r63_c75 bl[75] br[75] wl[63] vdd gnd cell_6t
Xbit_r64_c75 bl[75] br[75] wl[64] vdd gnd cell_6t
Xbit_r65_c75 bl[75] br[75] wl[65] vdd gnd cell_6t
Xbit_r66_c75 bl[75] br[75] wl[66] vdd gnd cell_6t
Xbit_r67_c75 bl[75] br[75] wl[67] vdd gnd cell_6t
Xbit_r68_c75 bl[75] br[75] wl[68] vdd gnd cell_6t
Xbit_r69_c75 bl[75] br[75] wl[69] vdd gnd cell_6t
Xbit_r70_c75 bl[75] br[75] wl[70] vdd gnd cell_6t
Xbit_r71_c75 bl[75] br[75] wl[71] vdd gnd cell_6t
Xbit_r72_c75 bl[75] br[75] wl[72] vdd gnd cell_6t
Xbit_r73_c75 bl[75] br[75] wl[73] vdd gnd cell_6t
Xbit_r74_c75 bl[75] br[75] wl[74] vdd gnd cell_6t
Xbit_r75_c75 bl[75] br[75] wl[75] vdd gnd cell_6t
Xbit_r76_c75 bl[75] br[75] wl[76] vdd gnd cell_6t
Xbit_r77_c75 bl[75] br[75] wl[77] vdd gnd cell_6t
Xbit_r78_c75 bl[75] br[75] wl[78] vdd gnd cell_6t
Xbit_r79_c75 bl[75] br[75] wl[79] vdd gnd cell_6t
Xbit_r80_c75 bl[75] br[75] wl[80] vdd gnd cell_6t
Xbit_r81_c75 bl[75] br[75] wl[81] vdd gnd cell_6t
Xbit_r82_c75 bl[75] br[75] wl[82] vdd gnd cell_6t
Xbit_r83_c75 bl[75] br[75] wl[83] vdd gnd cell_6t
Xbit_r84_c75 bl[75] br[75] wl[84] vdd gnd cell_6t
Xbit_r85_c75 bl[75] br[75] wl[85] vdd gnd cell_6t
Xbit_r86_c75 bl[75] br[75] wl[86] vdd gnd cell_6t
Xbit_r87_c75 bl[75] br[75] wl[87] vdd gnd cell_6t
Xbit_r88_c75 bl[75] br[75] wl[88] vdd gnd cell_6t
Xbit_r89_c75 bl[75] br[75] wl[89] vdd gnd cell_6t
Xbit_r90_c75 bl[75] br[75] wl[90] vdd gnd cell_6t
Xbit_r91_c75 bl[75] br[75] wl[91] vdd gnd cell_6t
Xbit_r92_c75 bl[75] br[75] wl[92] vdd gnd cell_6t
Xbit_r93_c75 bl[75] br[75] wl[93] vdd gnd cell_6t
Xbit_r94_c75 bl[75] br[75] wl[94] vdd gnd cell_6t
Xbit_r95_c75 bl[75] br[75] wl[95] vdd gnd cell_6t
Xbit_r96_c75 bl[75] br[75] wl[96] vdd gnd cell_6t
Xbit_r97_c75 bl[75] br[75] wl[97] vdd gnd cell_6t
Xbit_r98_c75 bl[75] br[75] wl[98] vdd gnd cell_6t
Xbit_r99_c75 bl[75] br[75] wl[99] vdd gnd cell_6t
Xbit_r100_c75 bl[75] br[75] wl[100] vdd gnd cell_6t
Xbit_r101_c75 bl[75] br[75] wl[101] vdd gnd cell_6t
Xbit_r102_c75 bl[75] br[75] wl[102] vdd gnd cell_6t
Xbit_r103_c75 bl[75] br[75] wl[103] vdd gnd cell_6t
Xbit_r104_c75 bl[75] br[75] wl[104] vdd gnd cell_6t
Xbit_r105_c75 bl[75] br[75] wl[105] vdd gnd cell_6t
Xbit_r106_c75 bl[75] br[75] wl[106] vdd gnd cell_6t
Xbit_r107_c75 bl[75] br[75] wl[107] vdd gnd cell_6t
Xbit_r108_c75 bl[75] br[75] wl[108] vdd gnd cell_6t
Xbit_r109_c75 bl[75] br[75] wl[109] vdd gnd cell_6t
Xbit_r110_c75 bl[75] br[75] wl[110] vdd gnd cell_6t
Xbit_r111_c75 bl[75] br[75] wl[111] vdd gnd cell_6t
Xbit_r112_c75 bl[75] br[75] wl[112] vdd gnd cell_6t
Xbit_r113_c75 bl[75] br[75] wl[113] vdd gnd cell_6t
Xbit_r114_c75 bl[75] br[75] wl[114] vdd gnd cell_6t
Xbit_r115_c75 bl[75] br[75] wl[115] vdd gnd cell_6t
Xbit_r116_c75 bl[75] br[75] wl[116] vdd gnd cell_6t
Xbit_r117_c75 bl[75] br[75] wl[117] vdd gnd cell_6t
Xbit_r118_c75 bl[75] br[75] wl[118] vdd gnd cell_6t
Xbit_r119_c75 bl[75] br[75] wl[119] vdd gnd cell_6t
Xbit_r120_c75 bl[75] br[75] wl[120] vdd gnd cell_6t
Xbit_r121_c75 bl[75] br[75] wl[121] vdd gnd cell_6t
Xbit_r122_c75 bl[75] br[75] wl[122] vdd gnd cell_6t
Xbit_r123_c75 bl[75] br[75] wl[123] vdd gnd cell_6t
Xbit_r124_c75 bl[75] br[75] wl[124] vdd gnd cell_6t
Xbit_r125_c75 bl[75] br[75] wl[125] vdd gnd cell_6t
Xbit_r126_c75 bl[75] br[75] wl[126] vdd gnd cell_6t
Xbit_r127_c75 bl[75] br[75] wl[127] vdd gnd cell_6t
Xbit_r128_c75 bl[75] br[75] wl[128] vdd gnd cell_6t
Xbit_r129_c75 bl[75] br[75] wl[129] vdd gnd cell_6t
Xbit_r130_c75 bl[75] br[75] wl[130] vdd gnd cell_6t
Xbit_r131_c75 bl[75] br[75] wl[131] vdd gnd cell_6t
Xbit_r132_c75 bl[75] br[75] wl[132] vdd gnd cell_6t
Xbit_r133_c75 bl[75] br[75] wl[133] vdd gnd cell_6t
Xbit_r134_c75 bl[75] br[75] wl[134] vdd gnd cell_6t
Xbit_r135_c75 bl[75] br[75] wl[135] vdd gnd cell_6t
Xbit_r136_c75 bl[75] br[75] wl[136] vdd gnd cell_6t
Xbit_r137_c75 bl[75] br[75] wl[137] vdd gnd cell_6t
Xbit_r138_c75 bl[75] br[75] wl[138] vdd gnd cell_6t
Xbit_r139_c75 bl[75] br[75] wl[139] vdd gnd cell_6t
Xbit_r140_c75 bl[75] br[75] wl[140] vdd gnd cell_6t
Xbit_r141_c75 bl[75] br[75] wl[141] vdd gnd cell_6t
Xbit_r142_c75 bl[75] br[75] wl[142] vdd gnd cell_6t
Xbit_r143_c75 bl[75] br[75] wl[143] vdd gnd cell_6t
Xbit_r144_c75 bl[75] br[75] wl[144] vdd gnd cell_6t
Xbit_r145_c75 bl[75] br[75] wl[145] vdd gnd cell_6t
Xbit_r146_c75 bl[75] br[75] wl[146] vdd gnd cell_6t
Xbit_r147_c75 bl[75] br[75] wl[147] vdd gnd cell_6t
Xbit_r148_c75 bl[75] br[75] wl[148] vdd gnd cell_6t
Xbit_r149_c75 bl[75] br[75] wl[149] vdd gnd cell_6t
Xbit_r150_c75 bl[75] br[75] wl[150] vdd gnd cell_6t
Xbit_r151_c75 bl[75] br[75] wl[151] vdd gnd cell_6t
Xbit_r152_c75 bl[75] br[75] wl[152] vdd gnd cell_6t
Xbit_r153_c75 bl[75] br[75] wl[153] vdd gnd cell_6t
Xbit_r154_c75 bl[75] br[75] wl[154] vdd gnd cell_6t
Xbit_r155_c75 bl[75] br[75] wl[155] vdd gnd cell_6t
Xbit_r156_c75 bl[75] br[75] wl[156] vdd gnd cell_6t
Xbit_r157_c75 bl[75] br[75] wl[157] vdd gnd cell_6t
Xbit_r158_c75 bl[75] br[75] wl[158] vdd gnd cell_6t
Xbit_r159_c75 bl[75] br[75] wl[159] vdd gnd cell_6t
Xbit_r160_c75 bl[75] br[75] wl[160] vdd gnd cell_6t
Xbit_r161_c75 bl[75] br[75] wl[161] vdd gnd cell_6t
Xbit_r162_c75 bl[75] br[75] wl[162] vdd gnd cell_6t
Xbit_r163_c75 bl[75] br[75] wl[163] vdd gnd cell_6t
Xbit_r164_c75 bl[75] br[75] wl[164] vdd gnd cell_6t
Xbit_r165_c75 bl[75] br[75] wl[165] vdd gnd cell_6t
Xbit_r166_c75 bl[75] br[75] wl[166] vdd gnd cell_6t
Xbit_r167_c75 bl[75] br[75] wl[167] vdd gnd cell_6t
Xbit_r168_c75 bl[75] br[75] wl[168] vdd gnd cell_6t
Xbit_r169_c75 bl[75] br[75] wl[169] vdd gnd cell_6t
Xbit_r170_c75 bl[75] br[75] wl[170] vdd gnd cell_6t
Xbit_r171_c75 bl[75] br[75] wl[171] vdd gnd cell_6t
Xbit_r172_c75 bl[75] br[75] wl[172] vdd gnd cell_6t
Xbit_r173_c75 bl[75] br[75] wl[173] vdd gnd cell_6t
Xbit_r174_c75 bl[75] br[75] wl[174] vdd gnd cell_6t
Xbit_r175_c75 bl[75] br[75] wl[175] vdd gnd cell_6t
Xbit_r176_c75 bl[75] br[75] wl[176] vdd gnd cell_6t
Xbit_r177_c75 bl[75] br[75] wl[177] vdd gnd cell_6t
Xbit_r178_c75 bl[75] br[75] wl[178] vdd gnd cell_6t
Xbit_r179_c75 bl[75] br[75] wl[179] vdd gnd cell_6t
Xbit_r180_c75 bl[75] br[75] wl[180] vdd gnd cell_6t
Xbit_r181_c75 bl[75] br[75] wl[181] vdd gnd cell_6t
Xbit_r182_c75 bl[75] br[75] wl[182] vdd gnd cell_6t
Xbit_r183_c75 bl[75] br[75] wl[183] vdd gnd cell_6t
Xbit_r184_c75 bl[75] br[75] wl[184] vdd gnd cell_6t
Xbit_r185_c75 bl[75] br[75] wl[185] vdd gnd cell_6t
Xbit_r186_c75 bl[75] br[75] wl[186] vdd gnd cell_6t
Xbit_r187_c75 bl[75] br[75] wl[187] vdd gnd cell_6t
Xbit_r188_c75 bl[75] br[75] wl[188] vdd gnd cell_6t
Xbit_r189_c75 bl[75] br[75] wl[189] vdd gnd cell_6t
Xbit_r190_c75 bl[75] br[75] wl[190] vdd gnd cell_6t
Xbit_r191_c75 bl[75] br[75] wl[191] vdd gnd cell_6t
Xbit_r192_c75 bl[75] br[75] wl[192] vdd gnd cell_6t
Xbit_r193_c75 bl[75] br[75] wl[193] vdd gnd cell_6t
Xbit_r194_c75 bl[75] br[75] wl[194] vdd gnd cell_6t
Xbit_r195_c75 bl[75] br[75] wl[195] vdd gnd cell_6t
Xbit_r196_c75 bl[75] br[75] wl[196] vdd gnd cell_6t
Xbit_r197_c75 bl[75] br[75] wl[197] vdd gnd cell_6t
Xbit_r198_c75 bl[75] br[75] wl[198] vdd gnd cell_6t
Xbit_r199_c75 bl[75] br[75] wl[199] vdd gnd cell_6t
Xbit_r200_c75 bl[75] br[75] wl[200] vdd gnd cell_6t
Xbit_r201_c75 bl[75] br[75] wl[201] vdd gnd cell_6t
Xbit_r202_c75 bl[75] br[75] wl[202] vdd gnd cell_6t
Xbit_r203_c75 bl[75] br[75] wl[203] vdd gnd cell_6t
Xbit_r204_c75 bl[75] br[75] wl[204] vdd gnd cell_6t
Xbit_r205_c75 bl[75] br[75] wl[205] vdd gnd cell_6t
Xbit_r206_c75 bl[75] br[75] wl[206] vdd gnd cell_6t
Xbit_r207_c75 bl[75] br[75] wl[207] vdd gnd cell_6t
Xbit_r208_c75 bl[75] br[75] wl[208] vdd gnd cell_6t
Xbit_r209_c75 bl[75] br[75] wl[209] vdd gnd cell_6t
Xbit_r210_c75 bl[75] br[75] wl[210] vdd gnd cell_6t
Xbit_r211_c75 bl[75] br[75] wl[211] vdd gnd cell_6t
Xbit_r212_c75 bl[75] br[75] wl[212] vdd gnd cell_6t
Xbit_r213_c75 bl[75] br[75] wl[213] vdd gnd cell_6t
Xbit_r214_c75 bl[75] br[75] wl[214] vdd gnd cell_6t
Xbit_r215_c75 bl[75] br[75] wl[215] vdd gnd cell_6t
Xbit_r216_c75 bl[75] br[75] wl[216] vdd gnd cell_6t
Xbit_r217_c75 bl[75] br[75] wl[217] vdd gnd cell_6t
Xbit_r218_c75 bl[75] br[75] wl[218] vdd gnd cell_6t
Xbit_r219_c75 bl[75] br[75] wl[219] vdd gnd cell_6t
Xbit_r220_c75 bl[75] br[75] wl[220] vdd gnd cell_6t
Xbit_r221_c75 bl[75] br[75] wl[221] vdd gnd cell_6t
Xbit_r222_c75 bl[75] br[75] wl[222] vdd gnd cell_6t
Xbit_r223_c75 bl[75] br[75] wl[223] vdd gnd cell_6t
Xbit_r224_c75 bl[75] br[75] wl[224] vdd gnd cell_6t
Xbit_r225_c75 bl[75] br[75] wl[225] vdd gnd cell_6t
Xbit_r226_c75 bl[75] br[75] wl[226] vdd gnd cell_6t
Xbit_r227_c75 bl[75] br[75] wl[227] vdd gnd cell_6t
Xbit_r228_c75 bl[75] br[75] wl[228] vdd gnd cell_6t
Xbit_r229_c75 bl[75] br[75] wl[229] vdd gnd cell_6t
Xbit_r230_c75 bl[75] br[75] wl[230] vdd gnd cell_6t
Xbit_r231_c75 bl[75] br[75] wl[231] vdd gnd cell_6t
Xbit_r232_c75 bl[75] br[75] wl[232] vdd gnd cell_6t
Xbit_r233_c75 bl[75] br[75] wl[233] vdd gnd cell_6t
Xbit_r234_c75 bl[75] br[75] wl[234] vdd gnd cell_6t
Xbit_r235_c75 bl[75] br[75] wl[235] vdd gnd cell_6t
Xbit_r236_c75 bl[75] br[75] wl[236] vdd gnd cell_6t
Xbit_r237_c75 bl[75] br[75] wl[237] vdd gnd cell_6t
Xbit_r238_c75 bl[75] br[75] wl[238] vdd gnd cell_6t
Xbit_r239_c75 bl[75] br[75] wl[239] vdd gnd cell_6t
Xbit_r240_c75 bl[75] br[75] wl[240] vdd gnd cell_6t
Xbit_r241_c75 bl[75] br[75] wl[241] vdd gnd cell_6t
Xbit_r242_c75 bl[75] br[75] wl[242] vdd gnd cell_6t
Xbit_r243_c75 bl[75] br[75] wl[243] vdd gnd cell_6t
Xbit_r244_c75 bl[75] br[75] wl[244] vdd gnd cell_6t
Xbit_r245_c75 bl[75] br[75] wl[245] vdd gnd cell_6t
Xbit_r246_c75 bl[75] br[75] wl[246] vdd gnd cell_6t
Xbit_r247_c75 bl[75] br[75] wl[247] vdd gnd cell_6t
Xbit_r248_c75 bl[75] br[75] wl[248] vdd gnd cell_6t
Xbit_r249_c75 bl[75] br[75] wl[249] vdd gnd cell_6t
Xbit_r250_c75 bl[75] br[75] wl[250] vdd gnd cell_6t
Xbit_r251_c75 bl[75] br[75] wl[251] vdd gnd cell_6t
Xbit_r252_c75 bl[75] br[75] wl[252] vdd gnd cell_6t
Xbit_r253_c75 bl[75] br[75] wl[253] vdd gnd cell_6t
Xbit_r254_c75 bl[75] br[75] wl[254] vdd gnd cell_6t
Xbit_r255_c75 bl[75] br[75] wl[255] vdd gnd cell_6t
Xbit_r256_c75 bl[75] br[75] wl[256] vdd gnd cell_6t
Xbit_r257_c75 bl[75] br[75] wl[257] vdd gnd cell_6t
Xbit_r258_c75 bl[75] br[75] wl[258] vdd gnd cell_6t
Xbit_r259_c75 bl[75] br[75] wl[259] vdd gnd cell_6t
Xbit_r260_c75 bl[75] br[75] wl[260] vdd gnd cell_6t
Xbit_r261_c75 bl[75] br[75] wl[261] vdd gnd cell_6t
Xbit_r262_c75 bl[75] br[75] wl[262] vdd gnd cell_6t
Xbit_r263_c75 bl[75] br[75] wl[263] vdd gnd cell_6t
Xbit_r264_c75 bl[75] br[75] wl[264] vdd gnd cell_6t
Xbit_r265_c75 bl[75] br[75] wl[265] vdd gnd cell_6t
Xbit_r266_c75 bl[75] br[75] wl[266] vdd gnd cell_6t
Xbit_r267_c75 bl[75] br[75] wl[267] vdd gnd cell_6t
Xbit_r268_c75 bl[75] br[75] wl[268] vdd gnd cell_6t
Xbit_r269_c75 bl[75] br[75] wl[269] vdd gnd cell_6t
Xbit_r270_c75 bl[75] br[75] wl[270] vdd gnd cell_6t
Xbit_r271_c75 bl[75] br[75] wl[271] vdd gnd cell_6t
Xbit_r272_c75 bl[75] br[75] wl[272] vdd gnd cell_6t
Xbit_r273_c75 bl[75] br[75] wl[273] vdd gnd cell_6t
Xbit_r274_c75 bl[75] br[75] wl[274] vdd gnd cell_6t
Xbit_r275_c75 bl[75] br[75] wl[275] vdd gnd cell_6t
Xbit_r276_c75 bl[75] br[75] wl[276] vdd gnd cell_6t
Xbit_r277_c75 bl[75] br[75] wl[277] vdd gnd cell_6t
Xbit_r278_c75 bl[75] br[75] wl[278] vdd gnd cell_6t
Xbit_r279_c75 bl[75] br[75] wl[279] vdd gnd cell_6t
Xbit_r280_c75 bl[75] br[75] wl[280] vdd gnd cell_6t
Xbit_r281_c75 bl[75] br[75] wl[281] vdd gnd cell_6t
Xbit_r282_c75 bl[75] br[75] wl[282] vdd gnd cell_6t
Xbit_r283_c75 bl[75] br[75] wl[283] vdd gnd cell_6t
Xbit_r284_c75 bl[75] br[75] wl[284] vdd gnd cell_6t
Xbit_r285_c75 bl[75] br[75] wl[285] vdd gnd cell_6t
Xbit_r286_c75 bl[75] br[75] wl[286] vdd gnd cell_6t
Xbit_r287_c75 bl[75] br[75] wl[287] vdd gnd cell_6t
Xbit_r288_c75 bl[75] br[75] wl[288] vdd gnd cell_6t
Xbit_r289_c75 bl[75] br[75] wl[289] vdd gnd cell_6t
Xbit_r290_c75 bl[75] br[75] wl[290] vdd gnd cell_6t
Xbit_r291_c75 bl[75] br[75] wl[291] vdd gnd cell_6t
Xbit_r292_c75 bl[75] br[75] wl[292] vdd gnd cell_6t
Xbit_r293_c75 bl[75] br[75] wl[293] vdd gnd cell_6t
Xbit_r294_c75 bl[75] br[75] wl[294] vdd gnd cell_6t
Xbit_r295_c75 bl[75] br[75] wl[295] vdd gnd cell_6t
Xbit_r296_c75 bl[75] br[75] wl[296] vdd gnd cell_6t
Xbit_r297_c75 bl[75] br[75] wl[297] vdd gnd cell_6t
Xbit_r298_c75 bl[75] br[75] wl[298] vdd gnd cell_6t
Xbit_r299_c75 bl[75] br[75] wl[299] vdd gnd cell_6t
Xbit_r300_c75 bl[75] br[75] wl[300] vdd gnd cell_6t
Xbit_r301_c75 bl[75] br[75] wl[301] vdd gnd cell_6t
Xbit_r302_c75 bl[75] br[75] wl[302] vdd gnd cell_6t
Xbit_r303_c75 bl[75] br[75] wl[303] vdd gnd cell_6t
Xbit_r304_c75 bl[75] br[75] wl[304] vdd gnd cell_6t
Xbit_r305_c75 bl[75] br[75] wl[305] vdd gnd cell_6t
Xbit_r306_c75 bl[75] br[75] wl[306] vdd gnd cell_6t
Xbit_r307_c75 bl[75] br[75] wl[307] vdd gnd cell_6t
Xbit_r308_c75 bl[75] br[75] wl[308] vdd gnd cell_6t
Xbit_r309_c75 bl[75] br[75] wl[309] vdd gnd cell_6t
Xbit_r310_c75 bl[75] br[75] wl[310] vdd gnd cell_6t
Xbit_r311_c75 bl[75] br[75] wl[311] vdd gnd cell_6t
Xbit_r312_c75 bl[75] br[75] wl[312] vdd gnd cell_6t
Xbit_r313_c75 bl[75] br[75] wl[313] vdd gnd cell_6t
Xbit_r314_c75 bl[75] br[75] wl[314] vdd gnd cell_6t
Xbit_r315_c75 bl[75] br[75] wl[315] vdd gnd cell_6t
Xbit_r316_c75 bl[75] br[75] wl[316] vdd gnd cell_6t
Xbit_r317_c75 bl[75] br[75] wl[317] vdd gnd cell_6t
Xbit_r318_c75 bl[75] br[75] wl[318] vdd gnd cell_6t
Xbit_r319_c75 bl[75] br[75] wl[319] vdd gnd cell_6t
Xbit_r320_c75 bl[75] br[75] wl[320] vdd gnd cell_6t
Xbit_r321_c75 bl[75] br[75] wl[321] vdd gnd cell_6t
Xbit_r322_c75 bl[75] br[75] wl[322] vdd gnd cell_6t
Xbit_r323_c75 bl[75] br[75] wl[323] vdd gnd cell_6t
Xbit_r324_c75 bl[75] br[75] wl[324] vdd gnd cell_6t
Xbit_r325_c75 bl[75] br[75] wl[325] vdd gnd cell_6t
Xbit_r326_c75 bl[75] br[75] wl[326] vdd gnd cell_6t
Xbit_r327_c75 bl[75] br[75] wl[327] vdd gnd cell_6t
Xbit_r328_c75 bl[75] br[75] wl[328] vdd gnd cell_6t
Xbit_r329_c75 bl[75] br[75] wl[329] vdd gnd cell_6t
Xbit_r330_c75 bl[75] br[75] wl[330] vdd gnd cell_6t
Xbit_r331_c75 bl[75] br[75] wl[331] vdd gnd cell_6t
Xbit_r332_c75 bl[75] br[75] wl[332] vdd gnd cell_6t
Xbit_r333_c75 bl[75] br[75] wl[333] vdd gnd cell_6t
Xbit_r334_c75 bl[75] br[75] wl[334] vdd gnd cell_6t
Xbit_r335_c75 bl[75] br[75] wl[335] vdd gnd cell_6t
Xbit_r336_c75 bl[75] br[75] wl[336] vdd gnd cell_6t
Xbit_r337_c75 bl[75] br[75] wl[337] vdd gnd cell_6t
Xbit_r338_c75 bl[75] br[75] wl[338] vdd gnd cell_6t
Xbit_r339_c75 bl[75] br[75] wl[339] vdd gnd cell_6t
Xbit_r340_c75 bl[75] br[75] wl[340] vdd gnd cell_6t
Xbit_r341_c75 bl[75] br[75] wl[341] vdd gnd cell_6t
Xbit_r342_c75 bl[75] br[75] wl[342] vdd gnd cell_6t
Xbit_r343_c75 bl[75] br[75] wl[343] vdd gnd cell_6t
Xbit_r344_c75 bl[75] br[75] wl[344] vdd gnd cell_6t
Xbit_r345_c75 bl[75] br[75] wl[345] vdd gnd cell_6t
Xbit_r346_c75 bl[75] br[75] wl[346] vdd gnd cell_6t
Xbit_r347_c75 bl[75] br[75] wl[347] vdd gnd cell_6t
Xbit_r348_c75 bl[75] br[75] wl[348] vdd gnd cell_6t
Xbit_r349_c75 bl[75] br[75] wl[349] vdd gnd cell_6t
Xbit_r350_c75 bl[75] br[75] wl[350] vdd gnd cell_6t
Xbit_r351_c75 bl[75] br[75] wl[351] vdd gnd cell_6t
Xbit_r352_c75 bl[75] br[75] wl[352] vdd gnd cell_6t
Xbit_r353_c75 bl[75] br[75] wl[353] vdd gnd cell_6t
Xbit_r354_c75 bl[75] br[75] wl[354] vdd gnd cell_6t
Xbit_r355_c75 bl[75] br[75] wl[355] vdd gnd cell_6t
Xbit_r356_c75 bl[75] br[75] wl[356] vdd gnd cell_6t
Xbit_r357_c75 bl[75] br[75] wl[357] vdd gnd cell_6t
Xbit_r358_c75 bl[75] br[75] wl[358] vdd gnd cell_6t
Xbit_r359_c75 bl[75] br[75] wl[359] vdd gnd cell_6t
Xbit_r360_c75 bl[75] br[75] wl[360] vdd gnd cell_6t
Xbit_r361_c75 bl[75] br[75] wl[361] vdd gnd cell_6t
Xbit_r362_c75 bl[75] br[75] wl[362] vdd gnd cell_6t
Xbit_r363_c75 bl[75] br[75] wl[363] vdd gnd cell_6t
Xbit_r364_c75 bl[75] br[75] wl[364] vdd gnd cell_6t
Xbit_r365_c75 bl[75] br[75] wl[365] vdd gnd cell_6t
Xbit_r366_c75 bl[75] br[75] wl[366] vdd gnd cell_6t
Xbit_r367_c75 bl[75] br[75] wl[367] vdd gnd cell_6t
Xbit_r368_c75 bl[75] br[75] wl[368] vdd gnd cell_6t
Xbit_r369_c75 bl[75] br[75] wl[369] vdd gnd cell_6t
Xbit_r370_c75 bl[75] br[75] wl[370] vdd gnd cell_6t
Xbit_r371_c75 bl[75] br[75] wl[371] vdd gnd cell_6t
Xbit_r372_c75 bl[75] br[75] wl[372] vdd gnd cell_6t
Xbit_r373_c75 bl[75] br[75] wl[373] vdd gnd cell_6t
Xbit_r374_c75 bl[75] br[75] wl[374] vdd gnd cell_6t
Xbit_r375_c75 bl[75] br[75] wl[375] vdd gnd cell_6t
Xbit_r376_c75 bl[75] br[75] wl[376] vdd gnd cell_6t
Xbit_r377_c75 bl[75] br[75] wl[377] vdd gnd cell_6t
Xbit_r378_c75 bl[75] br[75] wl[378] vdd gnd cell_6t
Xbit_r379_c75 bl[75] br[75] wl[379] vdd gnd cell_6t
Xbit_r380_c75 bl[75] br[75] wl[380] vdd gnd cell_6t
Xbit_r381_c75 bl[75] br[75] wl[381] vdd gnd cell_6t
Xbit_r382_c75 bl[75] br[75] wl[382] vdd gnd cell_6t
Xbit_r383_c75 bl[75] br[75] wl[383] vdd gnd cell_6t
Xbit_r384_c75 bl[75] br[75] wl[384] vdd gnd cell_6t
Xbit_r385_c75 bl[75] br[75] wl[385] vdd gnd cell_6t
Xbit_r386_c75 bl[75] br[75] wl[386] vdd gnd cell_6t
Xbit_r387_c75 bl[75] br[75] wl[387] vdd gnd cell_6t
Xbit_r388_c75 bl[75] br[75] wl[388] vdd gnd cell_6t
Xbit_r389_c75 bl[75] br[75] wl[389] vdd gnd cell_6t
Xbit_r390_c75 bl[75] br[75] wl[390] vdd gnd cell_6t
Xbit_r391_c75 bl[75] br[75] wl[391] vdd gnd cell_6t
Xbit_r392_c75 bl[75] br[75] wl[392] vdd gnd cell_6t
Xbit_r393_c75 bl[75] br[75] wl[393] vdd gnd cell_6t
Xbit_r394_c75 bl[75] br[75] wl[394] vdd gnd cell_6t
Xbit_r395_c75 bl[75] br[75] wl[395] vdd gnd cell_6t
Xbit_r396_c75 bl[75] br[75] wl[396] vdd gnd cell_6t
Xbit_r397_c75 bl[75] br[75] wl[397] vdd gnd cell_6t
Xbit_r398_c75 bl[75] br[75] wl[398] vdd gnd cell_6t
Xbit_r399_c75 bl[75] br[75] wl[399] vdd gnd cell_6t
Xbit_r400_c75 bl[75] br[75] wl[400] vdd gnd cell_6t
Xbit_r401_c75 bl[75] br[75] wl[401] vdd gnd cell_6t
Xbit_r402_c75 bl[75] br[75] wl[402] vdd gnd cell_6t
Xbit_r403_c75 bl[75] br[75] wl[403] vdd gnd cell_6t
Xbit_r404_c75 bl[75] br[75] wl[404] vdd gnd cell_6t
Xbit_r405_c75 bl[75] br[75] wl[405] vdd gnd cell_6t
Xbit_r406_c75 bl[75] br[75] wl[406] vdd gnd cell_6t
Xbit_r407_c75 bl[75] br[75] wl[407] vdd gnd cell_6t
Xbit_r408_c75 bl[75] br[75] wl[408] vdd gnd cell_6t
Xbit_r409_c75 bl[75] br[75] wl[409] vdd gnd cell_6t
Xbit_r410_c75 bl[75] br[75] wl[410] vdd gnd cell_6t
Xbit_r411_c75 bl[75] br[75] wl[411] vdd gnd cell_6t
Xbit_r412_c75 bl[75] br[75] wl[412] vdd gnd cell_6t
Xbit_r413_c75 bl[75] br[75] wl[413] vdd gnd cell_6t
Xbit_r414_c75 bl[75] br[75] wl[414] vdd gnd cell_6t
Xbit_r415_c75 bl[75] br[75] wl[415] vdd gnd cell_6t
Xbit_r416_c75 bl[75] br[75] wl[416] vdd gnd cell_6t
Xbit_r417_c75 bl[75] br[75] wl[417] vdd gnd cell_6t
Xbit_r418_c75 bl[75] br[75] wl[418] vdd gnd cell_6t
Xbit_r419_c75 bl[75] br[75] wl[419] vdd gnd cell_6t
Xbit_r420_c75 bl[75] br[75] wl[420] vdd gnd cell_6t
Xbit_r421_c75 bl[75] br[75] wl[421] vdd gnd cell_6t
Xbit_r422_c75 bl[75] br[75] wl[422] vdd gnd cell_6t
Xbit_r423_c75 bl[75] br[75] wl[423] vdd gnd cell_6t
Xbit_r424_c75 bl[75] br[75] wl[424] vdd gnd cell_6t
Xbit_r425_c75 bl[75] br[75] wl[425] vdd gnd cell_6t
Xbit_r426_c75 bl[75] br[75] wl[426] vdd gnd cell_6t
Xbit_r427_c75 bl[75] br[75] wl[427] vdd gnd cell_6t
Xbit_r428_c75 bl[75] br[75] wl[428] vdd gnd cell_6t
Xbit_r429_c75 bl[75] br[75] wl[429] vdd gnd cell_6t
Xbit_r430_c75 bl[75] br[75] wl[430] vdd gnd cell_6t
Xbit_r431_c75 bl[75] br[75] wl[431] vdd gnd cell_6t
Xbit_r432_c75 bl[75] br[75] wl[432] vdd gnd cell_6t
Xbit_r433_c75 bl[75] br[75] wl[433] vdd gnd cell_6t
Xbit_r434_c75 bl[75] br[75] wl[434] vdd gnd cell_6t
Xbit_r435_c75 bl[75] br[75] wl[435] vdd gnd cell_6t
Xbit_r436_c75 bl[75] br[75] wl[436] vdd gnd cell_6t
Xbit_r437_c75 bl[75] br[75] wl[437] vdd gnd cell_6t
Xbit_r438_c75 bl[75] br[75] wl[438] vdd gnd cell_6t
Xbit_r439_c75 bl[75] br[75] wl[439] vdd gnd cell_6t
Xbit_r440_c75 bl[75] br[75] wl[440] vdd gnd cell_6t
Xbit_r441_c75 bl[75] br[75] wl[441] vdd gnd cell_6t
Xbit_r442_c75 bl[75] br[75] wl[442] vdd gnd cell_6t
Xbit_r443_c75 bl[75] br[75] wl[443] vdd gnd cell_6t
Xbit_r444_c75 bl[75] br[75] wl[444] vdd gnd cell_6t
Xbit_r445_c75 bl[75] br[75] wl[445] vdd gnd cell_6t
Xbit_r446_c75 bl[75] br[75] wl[446] vdd gnd cell_6t
Xbit_r447_c75 bl[75] br[75] wl[447] vdd gnd cell_6t
Xbit_r448_c75 bl[75] br[75] wl[448] vdd gnd cell_6t
Xbit_r449_c75 bl[75] br[75] wl[449] vdd gnd cell_6t
Xbit_r450_c75 bl[75] br[75] wl[450] vdd gnd cell_6t
Xbit_r451_c75 bl[75] br[75] wl[451] vdd gnd cell_6t
Xbit_r452_c75 bl[75] br[75] wl[452] vdd gnd cell_6t
Xbit_r453_c75 bl[75] br[75] wl[453] vdd gnd cell_6t
Xbit_r454_c75 bl[75] br[75] wl[454] vdd gnd cell_6t
Xbit_r455_c75 bl[75] br[75] wl[455] vdd gnd cell_6t
Xbit_r456_c75 bl[75] br[75] wl[456] vdd gnd cell_6t
Xbit_r457_c75 bl[75] br[75] wl[457] vdd gnd cell_6t
Xbit_r458_c75 bl[75] br[75] wl[458] vdd gnd cell_6t
Xbit_r459_c75 bl[75] br[75] wl[459] vdd gnd cell_6t
Xbit_r460_c75 bl[75] br[75] wl[460] vdd gnd cell_6t
Xbit_r461_c75 bl[75] br[75] wl[461] vdd gnd cell_6t
Xbit_r462_c75 bl[75] br[75] wl[462] vdd gnd cell_6t
Xbit_r463_c75 bl[75] br[75] wl[463] vdd gnd cell_6t
Xbit_r464_c75 bl[75] br[75] wl[464] vdd gnd cell_6t
Xbit_r465_c75 bl[75] br[75] wl[465] vdd gnd cell_6t
Xbit_r466_c75 bl[75] br[75] wl[466] vdd gnd cell_6t
Xbit_r467_c75 bl[75] br[75] wl[467] vdd gnd cell_6t
Xbit_r468_c75 bl[75] br[75] wl[468] vdd gnd cell_6t
Xbit_r469_c75 bl[75] br[75] wl[469] vdd gnd cell_6t
Xbit_r470_c75 bl[75] br[75] wl[470] vdd gnd cell_6t
Xbit_r471_c75 bl[75] br[75] wl[471] vdd gnd cell_6t
Xbit_r472_c75 bl[75] br[75] wl[472] vdd gnd cell_6t
Xbit_r473_c75 bl[75] br[75] wl[473] vdd gnd cell_6t
Xbit_r474_c75 bl[75] br[75] wl[474] vdd gnd cell_6t
Xbit_r475_c75 bl[75] br[75] wl[475] vdd gnd cell_6t
Xbit_r476_c75 bl[75] br[75] wl[476] vdd gnd cell_6t
Xbit_r477_c75 bl[75] br[75] wl[477] vdd gnd cell_6t
Xbit_r478_c75 bl[75] br[75] wl[478] vdd gnd cell_6t
Xbit_r479_c75 bl[75] br[75] wl[479] vdd gnd cell_6t
Xbit_r480_c75 bl[75] br[75] wl[480] vdd gnd cell_6t
Xbit_r481_c75 bl[75] br[75] wl[481] vdd gnd cell_6t
Xbit_r482_c75 bl[75] br[75] wl[482] vdd gnd cell_6t
Xbit_r483_c75 bl[75] br[75] wl[483] vdd gnd cell_6t
Xbit_r484_c75 bl[75] br[75] wl[484] vdd gnd cell_6t
Xbit_r485_c75 bl[75] br[75] wl[485] vdd gnd cell_6t
Xbit_r486_c75 bl[75] br[75] wl[486] vdd gnd cell_6t
Xbit_r487_c75 bl[75] br[75] wl[487] vdd gnd cell_6t
Xbit_r488_c75 bl[75] br[75] wl[488] vdd gnd cell_6t
Xbit_r489_c75 bl[75] br[75] wl[489] vdd gnd cell_6t
Xbit_r490_c75 bl[75] br[75] wl[490] vdd gnd cell_6t
Xbit_r491_c75 bl[75] br[75] wl[491] vdd gnd cell_6t
Xbit_r492_c75 bl[75] br[75] wl[492] vdd gnd cell_6t
Xbit_r493_c75 bl[75] br[75] wl[493] vdd gnd cell_6t
Xbit_r494_c75 bl[75] br[75] wl[494] vdd gnd cell_6t
Xbit_r495_c75 bl[75] br[75] wl[495] vdd gnd cell_6t
Xbit_r496_c75 bl[75] br[75] wl[496] vdd gnd cell_6t
Xbit_r497_c75 bl[75] br[75] wl[497] vdd gnd cell_6t
Xbit_r498_c75 bl[75] br[75] wl[498] vdd gnd cell_6t
Xbit_r499_c75 bl[75] br[75] wl[499] vdd gnd cell_6t
Xbit_r500_c75 bl[75] br[75] wl[500] vdd gnd cell_6t
Xbit_r501_c75 bl[75] br[75] wl[501] vdd gnd cell_6t
Xbit_r502_c75 bl[75] br[75] wl[502] vdd gnd cell_6t
Xbit_r503_c75 bl[75] br[75] wl[503] vdd gnd cell_6t
Xbit_r504_c75 bl[75] br[75] wl[504] vdd gnd cell_6t
Xbit_r505_c75 bl[75] br[75] wl[505] vdd gnd cell_6t
Xbit_r506_c75 bl[75] br[75] wl[506] vdd gnd cell_6t
Xbit_r507_c75 bl[75] br[75] wl[507] vdd gnd cell_6t
Xbit_r508_c75 bl[75] br[75] wl[508] vdd gnd cell_6t
Xbit_r509_c75 bl[75] br[75] wl[509] vdd gnd cell_6t
Xbit_r510_c75 bl[75] br[75] wl[510] vdd gnd cell_6t
Xbit_r511_c75 bl[75] br[75] wl[511] vdd gnd cell_6t
Xbit_r0_c76 bl[76] br[76] wl[0] vdd gnd cell_6t
Xbit_r1_c76 bl[76] br[76] wl[1] vdd gnd cell_6t
Xbit_r2_c76 bl[76] br[76] wl[2] vdd gnd cell_6t
Xbit_r3_c76 bl[76] br[76] wl[3] vdd gnd cell_6t
Xbit_r4_c76 bl[76] br[76] wl[4] vdd gnd cell_6t
Xbit_r5_c76 bl[76] br[76] wl[5] vdd gnd cell_6t
Xbit_r6_c76 bl[76] br[76] wl[6] vdd gnd cell_6t
Xbit_r7_c76 bl[76] br[76] wl[7] vdd gnd cell_6t
Xbit_r8_c76 bl[76] br[76] wl[8] vdd gnd cell_6t
Xbit_r9_c76 bl[76] br[76] wl[9] vdd gnd cell_6t
Xbit_r10_c76 bl[76] br[76] wl[10] vdd gnd cell_6t
Xbit_r11_c76 bl[76] br[76] wl[11] vdd gnd cell_6t
Xbit_r12_c76 bl[76] br[76] wl[12] vdd gnd cell_6t
Xbit_r13_c76 bl[76] br[76] wl[13] vdd gnd cell_6t
Xbit_r14_c76 bl[76] br[76] wl[14] vdd gnd cell_6t
Xbit_r15_c76 bl[76] br[76] wl[15] vdd gnd cell_6t
Xbit_r16_c76 bl[76] br[76] wl[16] vdd gnd cell_6t
Xbit_r17_c76 bl[76] br[76] wl[17] vdd gnd cell_6t
Xbit_r18_c76 bl[76] br[76] wl[18] vdd gnd cell_6t
Xbit_r19_c76 bl[76] br[76] wl[19] vdd gnd cell_6t
Xbit_r20_c76 bl[76] br[76] wl[20] vdd gnd cell_6t
Xbit_r21_c76 bl[76] br[76] wl[21] vdd gnd cell_6t
Xbit_r22_c76 bl[76] br[76] wl[22] vdd gnd cell_6t
Xbit_r23_c76 bl[76] br[76] wl[23] vdd gnd cell_6t
Xbit_r24_c76 bl[76] br[76] wl[24] vdd gnd cell_6t
Xbit_r25_c76 bl[76] br[76] wl[25] vdd gnd cell_6t
Xbit_r26_c76 bl[76] br[76] wl[26] vdd gnd cell_6t
Xbit_r27_c76 bl[76] br[76] wl[27] vdd gnd cell_6t
Xbit_r28_c76 bl[76] br[76] wl[28] vdd gnd cell_6t
Xbit_r29_c76 bl[76] br[76] wl[29] vdd gnd cell_6t
Xbit_r30_c76 bl[76] br[76] wl[30] vdd gnd cell_6t
Xbit_r31_c76 bl[76] br[76] wl[31] vdd gnd cell_6t
Xbit_r32_c76 bl[76] br[76] wl[32] vdd gnd cell_6t
Xbit_r33_c76 bl[76] br[76] wl[33] vdd gnd cell_6t
Xbit_r34_c76 bl[76] br[76] wl[34] vdd gnd cell_6t
Xbit_r35_c76 bl[76] br[76] wl[35] vdd gnd cell_6t
Xbit_r36_c76 bl[76] br[76] wl[36] vdd gnd cell_6t
Xbit_r37_c76 bl[76] br[76] wl[37] vdd gnd cell_6t
Xbit_r38_c76 bl[76] br[76] wl[38] vdd gnd cell_6t
Xbit_r39_c76 bl[76] br[76] wl[39] vdd gnd cell_6t
Xbit_r40_c76 bl[76] br[76] wl[40] vdd gnd cell_6t
Xbit_r41_c76 bl[76] br[76] wl[41] vdd gnd cell_6t
Xbit_r42_c76 bl[76] br[76] wl[42] vdd gnd cell_6t
Xbit_r43_c76 bl[76] br[76] wl[43] vdd gnd cell_6t
Xbit_r44_c76 bl[76] br[76] wl[44] vdd gnd cell_6t
Xbit_r45_c76 bl[76] br[76] wl[45] vdd gnd cell_6t
Xbit_r46_c76 bl[76] br[76] wl[46] vdd gnd cell_6t
Xbit_r47_c76 bl[76] br[76] wl[47] vdd gnd cell_6t
Xbit_r48_c76 bl[76] br[76] wl[48] vdd gnd cell_6t
Xbit_r49_c76 bl[76] br[76] wl[49] vdd gnd cell_6t
Xbit_r50_c76 bl[76] br[76] wl[50] vdd gnd cell_6t
Xbit_r51_c76 bl[76] br[76] wl[51] vdd gnd cell_6t
Xbit_r52_c76 bl[76] br[76] wl[52] vdd gnd cell_6t
Xbit_r53_c76 bl[76] br[76] wl[53] vdd gnd cell_6t
Xbit_r54_c76 bl[76] br[76] wl[54] vdd gnd cell_6t
Xbit_r55_c76 bl[76] br[76] wl[55] vdd gnd cell_6t
Xbit_r56_c76 bl[76] br[76] wl[56] vdd gnd cell_6t
Xbit_r57_c76 bl[76] br[76] wl[57] vdd gnd cell_6t
Xbit_r58_c76 bl[76] br[76] wl[58] vdd gnd cell_6t
Xbit_r59_c76 bl[76] br[76] wl[59] vdd gnd cell_6t
Xbit_r60_c76 bl[76] br[76] wl[60] vdd gnd cell_6t
Xbit_r61_c76 bl[76] br[76] wl[61] vdd gnd cell_6t
Xbit_r62_c76 bl[76] br[76] wl[62] vdd gnd cell_6t
Xbit_r63_c76 bl[76] br[76] wl[63] vdd gnd cell_6t
Xbit_r64_c76 bl[76] br[76] wl[64] vdd gnd cell_6t
Xbit_r65_c76 bl[76] br[76] wl[65] vdd gnd cell_6t
Xbit_r66_c76 bl[76] br[76] wl[66] vdd gnd cell_6t
Xbit_r67_c76 bl[76] br[76] wl[67] vdd gnd cell_6t
Xbit_r68_c76 bl[76] br[76] wl[68] vdd gnd cell_6t
Xbit_r69_c76 bl[76] br[76] wl[69] vdd gnd cell_6t
Xbit_r70_c76 bl[76] br[76] wl[70] vdd gnd cell_6t
Xbit_r71_c76 bl[76] br[76] wl[71] vdd gnd cell_6t
Xbit_r72_c76 bl[76] br[76] wl[72] vdd gnd cell_6t
Xbit_r73_c76 bl[76] br[76] wl[73] vdd gnd cell_6t
Xbit_r74_c76 bl[76] br[76] wl[74] vdd gnd cell_6t
Xbit_r75_c76 bl[76] br[76] wl[75] vdd gnd cell_6t
Xbit_r76_c76 bl[76] br[76] wl[76] vdd gnd cell_6t
Xbit_r77_c76 bl[76] br[76] wl[77] vdd gnd cell_6t
Xbit_r78_c76 bl[76] br[76] wl[78] vdd gnd cell_6t
Xbit_r79_c76 bl[76] br[76] wl[79] vdd gnd cell_6t
Xbit_r80_c76 bl[76] br[76] wl[80] vdd gnd cell_6t
Xbit_r81_c76 bl[76] br[76] wl[81] vdd gnd cell_6t
Xbit_r82_c76 bl[76] br[76] wl[82] vdd gnd cell_6t
Xbit_r83_c76 bl[76] br[76] wl[83] vdd gnd cell_6t
Xbit_r84_c76 bl[76] br[76] wl[84] vdd gnd cell_6t
Xbit_r85_c76 bl[76] br[76] wl[85] vdd gnd cell_6t
Xbit_r86_c76 bl[76] br[76] wl[86] vdd gnd cell_6t
Xbit_r87_c76 bl[76] br[76] wl[87] vdd gnd cell_6t
Xbit_r88_c76 bl[76] br[76] wl[88] vdd gnd cell_6t
Xbit_r89_c76 bl[76] br[76] wl[89] vdd gnd cell_6t
Xbit_r90_c76 bl[76] br[76] wl[90] vdd gnd cell_6t
Xbit_r91_c76 bl[76] br[76] wl[91] vdd gnd cell_6t
Xbit_r92_c76 bl[76] br[76] wl[92] vdd gnd cell_6t
Xbit_r93_c76 bl[76] br[76] wl[93] vdd gnd cell_6t
Xbit_r94_c76 bl[76] br[76] wl[94] vdd gnd cell_6t
Xbit_r95_c76 bl[76] br[76] wl[95] vdd gnd cell_6t
Xbit_r96_c76 bl[76] br[76] wl[96] vdd gnd cell_6t
Xbit_r97_c76 bl[76] br[76] wl[97] vdd gnd cell_6t
Xbit_r98_c76 bl[76] br[76] wl[98] vdd gnd cell_6t
Xbit_r99_c76 bl[76] br[76] wl[99] vdd gnd cell_6t
Xbit_r100_c76 bl[76] br[76] wl[100] vdd gnd cell_6t
Xbit_r101_c76 bl[76] br[76] wl[101] vdd gnd cell_6t
Xbit_r102_c76 bl[76] br[76] wl[102] vdd gnd cell_6t
Xbit_r103_c76 bl[76] br[76] wl[103] vdd gnd cell_6t
Xbit_r104_c76 bl[76] br[76] wl[104] vdd gnd cell_6t
Xbit_r105_c76 bl[76] br[76] wl[105] vdd gnd cell_6t
Xbit_r106_c76 bl[76] br[76] wl[106] vdd gnd cell_6t
Xbit_r107_c76 bl[76] br[76] wl[107] vdd gnd cell_6t
Xbit_r108_c76 bl[76] br[76] wl[108] vdd gnd cell_6t
Xbit_r109_c76 bl[76] br[76] wl[109] vdd gnd cell_6t
Xbit_r110_c76 bl[76] br[76] wl[110] vdd gnd cell_6t
Xbit_r111_c76 bl[76] br[76] wl[111] vdd gnd cell_6t
Xbit_r112_c76 bl[76] br[76] wl[112] vdd gnd cell_6t
Xbit_r113_c76 bl[76] br[76] wl[113] vdd gnd cell_6t
Xbit_r114_c76 bl[76] br[76] wl[114] vdd gnd cell_6t
Xbit_r115_c76 bl[76] br[76] wl[115] vdd gnd cell_6t
Xbit_r116_c76 bl[76] br[76] wl[116] vdd gnd cell_6t
Xbit_r117_c76 bl[76] br[76] wl[117] vdd gnd cell_6t
Xbit_r118_c76 bl[76] br[76] wl[118] vdd gnd cell_6t
Xbit_r119_c76 bl[76] br[76] wl[119] vdd gnd cell_6t
Xbit_r120_c76 bl[76] br[76] wl[120] vdd gnd cell_6t
Xbit_r121_c76 bl[76] br[76] wl[121] vdd gnd cell_6t
Xbit_r122_c76 bl[76] br[76] wl[122] vdd gnd cell_6t
Xbit_r123_c76 bl[76] br[76] wl[123] vdd gnd cell_6t
Xbit_r124_c76 bl[76] br[76] wl[124] vdd gnd cell_6t
Xbit_r125_c76 bl[76] br[76] wl[125] vdd gnd cell_6t
Xbit_r126_c76 bl[76] br[76] wl[126] vdd gnd cell_6t
Xbit_r127_c76 bl[76] br[76] wl[127] vdd gnd cell_6t
Xbit_r128_c76 bl[76] br[76] wl[128] vdd gnd cell_6t
Xbit_r129_c76 bl[76] br[76] wl[129] vdd gnd cell_6t
Xbit_r130_c76 bl[76] br[76] wl[130] vdd gnd cell_6t
Xbit_r131_c76 bl[76] br[76] wl[131] vdd gnd cell_6t
Xbit_r132_c76 bl[76] br[76] wl[132] vdd gnd cell_6t
Xbit_r133_c76 bl[76] br[76] wl[133] vdd gnd cell_6t
Xbit_r134_c76 bl[76] br[76] wl[134] vdd gnd cell_6t
Xbit_r135_c76 bl[76] br[76] wl[135] vdd gnd cell_6t
Xbit_r136_c76 bl[76] br[76] wl[136] vdd gnd cell_6t
Xbit_r137_c76 bl[76] br[76] wl[137] vdd gnd cell_6t
Xbit_r138_c76 bl[76] br[76] wl[138] vdd gnd cell_6t
Xbit_r139_c76 bl[76] br[76] wl[139] vdd gnd cell_6t
Xbit_r140_c76 bl[76] br[76] wl[140] vdd gnd cell_6t
Xbit_r141_c76 bl[76] br[76] wl[141] vdd gnd cell_6t
Xbit_r142_c76 bl[76] br[76] wl[142] vdd gnd cell_6t
Xbit_r143_c76 bl[76] br[76] wl[143] vdd gnd cell_6t
Xbit_r144_c76 bl[76] br[76] wl[144] vdd gnd cell_6t
Xbit_r145_c76 bl[76] br[76] wl[145] vdd gnd cell_6t
Xbit_r146_c76 bl[76] br[76] wl[146] vdd gnd cell_6t
Xbit_r147_c76 bl[76] br[76] wl[147] vdd gnd cell_6t
Xbit_r148_c76 bl[76] br[76] wl[148] vdd gnd cell_6t
Xbit_r149_c76 bl[76] br[76] wl[149] vdd gnd cell_6t
Xbit_r150_c76 bl[76] br[76] wl[150] vdd gnd cell_6t
Xbit_r151_c76 bl[76] br[76] wl[151] vdd gnd cell_6t
Xbit_r152_c76 bl[76] br[76] wl[152] vdd gnd cell_6t
Xbit_r153_c76 bl[76] br[76] wl[153] vdd gnd cell_6t
Xbit_r154_c76 bl[76] br[76] wl[154] vdd gnd cell_6t
Xbit_r155_c76 bl[76] br[76] wl[155] vdd gnd cell_6t
Xbit_r156_c76 bl[76] br[76] wl[156] vdd gnd cell_6t
Xbit_r157_c76 bl[76] br[76] wl[157] vdd gnd cell_6t
Xbit_r158_c76 bl[76] br[76] wl[158] vdd gnd cell_6t
Xbit_r159_c76 bl[76] br[76] wl[159] vdd gnd cell_6t
Xbit_r160_c76 bl[76] br[76] wl[160] vdd gnd cell_6t
Xbit_r161_c76 bl[76] br[76] wl[161] vdd gnd cell_6t
Xbit_r162_c76 bl[76] br[76] wl[162] vdd gnd cell_6t
Xbit_r163_c76 bl[76] br[76] wl[163] vdd gnd cell_6t
Xbit_r164_c76 bl[76] br[76] wl[164] vdd gnd cell_6t
Xbit_r165_c76 bl[76] br[76] wl[165] vdd gnd cell_6t
Xbit_r166_c76 bl[76] br[76] wl[166] vdd gnd cell_6t
Xbit_r167_c76 bl[76] br[76] wl[167] vdd gnd cell_6t
Xbit_r168_c76 bl[76] br[76] wl[168] vdd gnd cell_6t
Xbit_r169_c76 bl[76] br[76] wl[169] vdd gnd cell_6t
Xbit_r170_c76 bl[76] br[76] wl[170] vdd gnd cell_6t
Xbit_r171_c76 bl[76] br[76] wl[171] vdd gnd cell_6t
Xbit_r172_c76 bl[76] br[76] wl[172] vdd gnd cell_6t
Xbit_r173_c76 bl[76] br[76] wl[173] vdd gnd cell_6t
Xbit_r174_c76 bl[76] br[76] wl[174] vdd gnd cell_6t
Xbit_r175_c76 bl[76] br[76] wl[175] vdd gnd cell_6t
Xbit_r176_c76 bl[76] br[76] wl[176] vdd gnd cell_6t
Xbit_r177_c76 bl[76] br[76] wl[177] vdd gnd cell_6t
Xbit_r178_c76 bl[76] br[76] wl[178] vdd gnd cell_6t
Xbit_r179_c76 bl[76] br[76] wl[179] vdd gnd cell_6t
Xbit_r180_c76 bl[76] br[76] wl[180] vdd gnd cell_6t
Xbit_r181_c76 bl[76] br[76] wl[181] vdd gnd cell_6t
Xbit_r182_c76 bl[76] br[76] wl[182] vdd gnd cell_6t
Xbit_r183_c76 bl[76] br[76] wl[183] vdd gnd cell_6t
Xbit_r184_c76 bl[76] br[76] wl[184] vdd gnd cell_6t
Xbit_r185_c76 bl[76] br[76] wl[185] vdd gnd cell_6t
Xbit_r186_c76 bl[76] br[76] wl[186] vdd gnd cell_6t
Xbit_r187_c76 bl[76] br[76] wl[187] vdd gnd cell_6t
Xbit_r188_c76 bl[76] br[76] wl[188] vdd gnd cell_6t
Xbit_r189_c76 bl[76] br[76] wl[189] vdd gnd cell_6t
Xbit_r190_c76 bl[76] br[76] wl[190] vdd gnd cell_6t
Xbit_r191_c76 bl[76] br[76] wl[191] vdd gnd cell_6t
Xbit_r192_c76 bl[76] br[76] wl[192] vdd gnd cell_6t
Xbit_r193_c76 bl[76] br[76] wl[193] vdd gnd cell_6t
Xbit_r194_c76 bl[76] br[76] wl[194] vdd gnd cell_6t
Xbit_r195_c76 bl[76] br[76] wl[195] vdd gnd cell_6t
Xbit_r196_c76 bl[76] br[76] wl[196] vdd gnd cell_6t
Xbit_r197_c76 bl[76] br[76] wl[197] vdd gnd cell_6t
Xbit_r198_c76 bl[76] br[76] wl[198] vdd gnd cell_6t
Xbit_r199_c76 bl[76] br[76] wl[199] vdd gnd cell_6t
Xbit_r200_c76 bl[76] br[76] wl[200] vdd gnd cell_6t
Xbit_r201_c76 bl[76] br[76] wl[201] vdd gnd cell_6t
Xbit_r202_c76 bl[76] br[76] wl[202] vdd gnd cell_6t
Xbit_r203_c76 bl[76] br[76] wl[203] vdd gnd cell_6t
Xbit_r204_c76 bl[76] br[76] wl[204] vdd gnd cell_6t
Xbit_r205_c76 bl[76] br[76] wl[205] vdd gnd cell_6t
Xbit_r206_c76 bl[76] br[76] wl[206] vdd gnd cell_6t
Xbit_r207_c76 bl[76] br[76] wl[207] vdd gnd cell_6t
Xbit_r208_c76 bl[76] br[76] wl[208] vdd gnd cell_6t
Xbit_r209_c76 bl[76] br[76] wl[209] vdd gnd cell_6t
Xbit_r210_c76 bl[76] br[76] wl[210] vdd gnd cell_6t
Xbit_r211_c76 bl[76] br[76] wl[211] vdd gnd cell_6t
Xbit_r212_c76 bl[76] br[76] wl[212] vdd gnd cell_6t
Xbit_r213_c76 bl[76] br[76] wl[213] vdd gnd cell_6t
Xbit_r214_c76 bl[76] br[76] wl[214] vdd gnd cell_6t
Xbit_r215_c76 bl[76] br[76] wl[215] vdd gnd cell_6t
Xbit_r216_c76 bl[76] br[76] wl[216] vdd gnd cell_6t
Xbit_r217_c76 bl[76] br[76] wl[217] vdd gnd cell_6t
Xbit_r218_c76 bl[76] br[76] wl[218] vdd gnd cell_6t
Xbit_r219_c76 bl[76] br[76] wl[219] vdd gnd cell_6t
Xbit_r220_c76 bl[76] br[76] wl[220] vdd gnd cell_6t
Xbit_r221_c76 bl[76] br[76] wl[221] vdd gnd cell_6t
Xbit_r222_c76 bl[76] br[76] wl[222] vdd gnd cell_6t
Xbit_r223_c76 bl[76] br[76] wl[223] vdd gnd cell_6t
Xbit_r224_c76 bl[76] br[76] wl[224] vdd gnd cell_6t
Xbit_r225_c76 bl[76] br[76] wl[225] vdd gnd cell_6t
Xbit_r226_c76 bl[76] br[76] wl[226] vdd gnd cell_6t
Xbit_r227_c76 bl[76] br[76] wl[227] vdd gnd cell_6t
Xbit_r228_c76 bl[76] br[76] wl[228] vdd gnd cell_6t
Xbit_r229_c76 bl[76] br[76] wl[229] vdd gnd cell_6t
Xbit_r230_c76 bl[76] br[76] wl[230] vdd gnd cell_6t
Xbit_r231_c76 bl[76] br[76] wl[231] vdd gnd cell_6t
Xbit_r232_c76 bl[76] br[76] wl[232] vdd gnd cell_6t
Xbit_r233_c76 bl[76] br[76] wl[233] vdd gnd cell_6t
Xbit_r234_c76 bl[76] br[76] wl[234] vdd gnd cell_6t
Xbit_r235_c76 bl[76] br[76] wl[235] vdd gnd cell_6t
Xbit_r236_c76 bl[76] br[76] wl[236] vdd gnd cell_6t
Xbit_r237_c76 bl[76] br[76] wl[237] vdd gnd cell_6t
Xbit_r238_c76 bl[76] br[76] wl[238] vdd gnd cell_6t
Xbit_r239_c76 bl[76] br[76] wl[239] vdd gnd cell_6t
Xbit_r240_c76 bl[76] br[76] wl[240] vdd gnd cell_6t
Xbit_r241_c76 bl[76] br[76] wl[241] vdd gnd cell_6t
Xbit_r242_c76 bl[76] br[76] wl[242] vdd gnd cell_6t
Xbit_r243_c76 bl[76] br[76] wl[243] vdd gnd cell_6t
Xbit_r244_c76 bl[76] br[76] wl[244] vdd gnd cell_6t
Xbit_r245_c76 bl[76] br[76] wl[245] vdd gnd cell_6t
Xbit_r246_c76 bl[76] br[76] wl[246] vdd gnd cell_6t
Xbit_r247_c76 bl[76] br[76] wl[247] vdd gnd cell_6t
Xbit_r248_c76 bl[76] br[76] wl[248] vdd gnd cell_6t
Xbit_r249_c76 bl[76] br[76] wl[249] vdd gnd cell_6t
Xbit_r250_c76 bl[76] br[76] wl[250] vdd gnd cell_6t
Xbit_r251_c76 bl[76] br[76] wl[251] vdd gnd cell_6t
Xbit_r252_c76 bl[76] br[76] wl[252] vdd gnd cell_6t
Xbit_r253_c76 bl[76] br[76] wl[253] vdd gnd cell_6t
Xbit_r254_c76 bl[76] br[76] wl[254] vdd gnd cell_6t
Xbit_r255_c76 bl[76] br[76] wl[255] vdd gnd cell_6t
Xbit_r256_c76 bl[76] br[76] wl[256] vdd gnd cell_6t
Xbit_r257_c76 bl[76] br[76] wl[257] vdd gnd cell_6t
Xbit_r258_c76 bl[76] br[76] wl[258] vdd gnd cell_6t
Xbit_r259_c76 bl[76] br[76] wl[259] vdd gnd cell_6t
Xbit_r260_c76 bl[76] br[76] wl[260] vdd gnd cell_6t
Xbit_r261_c76 bl[76] br[76] wl[261] vdd gnd cell_6t
Xbit_r262_c76 bl[76] br[76] wl[262] vdd gnd cell_6t
Xbit_r263_c76 bl[76] br[76] wl[263] vdd gnd cell_6t
Xbit_r264_c76 bl[76] br[76] wl[264] vdd gnd cell_6t
Xbit_r265_c76 bl[76] br[76] wl[265] vdd gnd cell_6t
Xbit_r266_c76 bl[76] br[76] wl[266] vdd gnd cell_6t
Xbit_r267_c76 bl[76] br[76] wl[267] vdd gnd cell_6t
Xbit_r268_c76 bl[76] br[76] wl[268] vdd gnd cell_6t
Xbit_r269_c76 bl[76] br[76] wl[269] vdd gnd cell_6t
Xbit_r270_c76 bl[76] br[76] wl[270] vdd gnd cell_6t
Xbit_r271_c76 bl[76] br[76] wl[271] vdd gnd cell_6t
Xbit_r272_c76 bl[76] br[76] wl[272] vdd gnd cell_6t
Xbit_r273_c76 bl[76] br[76] wl[273] vdd gnd cell_6t
Xbit_r274_c76 bl[76] br[76] wl[274] vdd gnd cell_6t
Xbit_r275_c76 bl[76] br[76] wl[275] vdd gnd cell_6t
Xbit_r276_c76 bl[76] br[76] wl[276] vdd gnd cell_6t
Xbit_r277_c76 bl[76] br[76] wl[277] vdd gnd cell_6t
Xbit_r278_c76 bl[76] br[76] wl[278] vdd gnd cell_6t
Xbit_r279_c76 bl[76] br[76] wl[279] vdd gnd cell_6t
Xbit_r280_c76 bl[76] br[76] wl[280] vdd gnd cell_6t
Xbit_r281_c76 bl[76] br[76] wl[281] vdd gnd cell_6t
Xbit_r282_c76 bl[76] br[76] wl[282] vdd gnd cell_6t
Xbit_r283_c76 bl[76] br[76] wl[283] vdd gnd cell_6t
Xbit_r284_c76 bl[76] br[76] wl[284] vdd gnd cell_6t
Xbit_r285_c76 bl[76] br[76] wl[285] vdd gnd cell_6t
Xbit_r286_c76 bl[76] br[76] wl[286] vdd gnd cell_6t
Xbit_r287_c76 bl[76] br[76] wl[287] vdd gnd cell_6t
Xbit_r288_c76 bl[76] br[76] wl[288] vdd gnd cell_6t
Xbit_r289_c76 bl[76] br[76] wl[289] vdd gnd cell_6t
Xbit_r290_c76 bl[76] br[76] wl[290] vdd gnd cell_6t
Xbit_r291_c76 bl[76] br[76] wl[291] vdd gnd cell_6t
Xbit_r292_c76 bl[76] br[76] wl[292] vdd gnd cell_6t
Xbit_r293_c76 bl[76] br[76] wl[293] vdd gnd cell_6t
Xbit_r294_c76 bl[76] br[76] wl[294] vdd gnd cell_6t
Xbit_r295_c76 bl[76] br[76] wl[295] vdd gnd cell_6t
Xbit_r296_c76 bl[76] br[76] wl[296] vdd gnd cell_6t
Xbit_r297_c76 bl[76] br[76] wl[297] vdd gnd cell_6t
Xbit_r298_c76 bl[76] br[76] wl[298] vdd gnd cell_6t
Xbit_r299_c76 bl[76] br[76] wl[299] vdd gnd cell_6t
Xbit_r300_c76 bl[76] br[76] wl[300] vdd gnd cell_6t
Xbit_r301_c76 bl[76] br[76] wl[301] vdd gnd cell_6t
Xbit_r302_c76 bl[76] br[76] wl[302] vdd gnd cell_6t
Xbit_r303_c76 bl[76] br[76] wl[303] vdd gnd cell_6t
Xbit_r304_c76 bl[76] br[76] wl[304] vdd gnd cell_6t
Xbit_r305_c76 bl[76] br[76] wl[305] vdd gnd cell_6t
Xbit_r306_c76 bl[76] br[76] wl[306] vdd gnd cell_6t
Xbit_r307_c76 bl[76] br[76] wl[307] vdd gnd cell_6t
Xbit_r308_c76 bl[76] br[76] wl[308] vdd gnd cell_6t
Xbit_r309_c76 bl[76] br[76] wl[309] vdd gnd cell_6t
Xbit_r310_c76 bl[76] br[76] wl[310] vdd gnd cell_6t
Xbit_r311_c76 bl[76] br[76] wl[311] vdd gnd cell_6t
Xbit_r312_c76 bl[76] br[76] wl[312] vdd gnd cell_6t
Xbit_r313_c76 bl[76] br[76] wl[313] vdd gnd cell_6t
Xbit_r314_c76 bl[76] br[76] wl[314] vdd gnd cell_6t
Xbit_r315_c76 bl[76] br[76] wl[315] vdd gnd cell_6t
Xbit_r316_c76 bl[76] br[76] wl[316] vdd gnd cell_6t
Xbit_r317_c76 bl[76] br[76] wl[317] vdd gnd cell_6t
Xbit_r318_c76 bl[76] br[76] wl[318] vdd gnd cell_6t
Xbit_r319_c76 bl[76] br[76] wl[319] vdd gnd cell_6t
Xbit_r320_c76 bl[76] br[76] wl[320] vdd gnd cell_6t
Xbit_r321_c76 bl[76] br[76] wl[321] vdd gnd cell_6t
Xbit_r322_c76 bl[76] br[76] wl[322] vdd gnd cell_6t
Xbit_r323_c76 bl[76] br[76] wl[323] vdd gnd cell_6t
Xbit_r324_c76 bl[76] br[76] wl[324] vdd gnd cell_6t
Xbit_r325_c76 bl[76] br[76] wl[325] vdd gnd cell_6t
Xbit_r326_c76 bl[76] br[76] wl[326] vdd gnd cell_6t
Xbit_r327_c76 bl[76] br[76] wl[327] vdd gnd cell_6t
Xbit_r328_c76 bl[76] br[76] wl[328] vdd gnd cell_6t
Xbit_r329_c76 bl[76] br[76] wl[329] vdd gnd cell_6t
Xbit_r330_c76 bl[76] br[76] wl[330] vdd gnd cell_6t
Xbit_r331_c76 bl[76] br[76] wl[331] vdd gnd cell_6t
Xbit_r332_c76 bl[76] br[76] wl[332] vdd gnd cell_6t
Xbit_r333_c76 bl[76] br[76] wl[333] vdd gnd cell_6t
Xbit_r334_c76 bl[76] br[76] wl[334] vdd gnd cell_6t
Xbit_r335_c76 bl[76] br[76] wl[335] vdd gnd cell_6t
Xbit_r336_c76 bl[76] br[76] wl[336] vdd gnd cell_6t
Xbit_r337_c76 bl[76] br[76] wl[337] vdd gnd cell_6t
Xbit_r338_c76 bl[76] br[76] wl[338] vdd gnd cell_6t
Xbit_r339_c76 bl[76] br[76] wl[339] vdd gnd cell_6t
Xbit_r340_c76 bl[76] br[76] wl[340] vdd gnd cell_6t
Xbit_r341_c76 bl[76] br[76] wl[341] vdd gnd cell_6t
Xbit_r342_c76 bl[76] br[76] wl[342] vdd gnd cell_6t
Xbit_r343_c76 bl[76] br[76] wl[343] vdd gnd cell_6t
Xbit_r344_c76 bl[76] br[76] wl[344] vdd gnd cell_6t
Xbit_r345_c76 bl[76] br[76] wl[345] vdd gnd cell_6t
Xbit_r346_c76 bl[76] br[76] wl[346] vdd gnd cell_6t
Xbit_r347_c76 bl[76] br[76] wl[347] vdd gnd cell_6t
Xbit_r348_c76 bl[76] br[76] wl[348] vdd gnd cell_6t
Xbit_r349_c76 bl[76] br[76] wl[349] vdd gnd cell_6t
Xbit_r350_c76 bl[76] br[76] wl[350] vdd gnd cell_6t
Xbit_r351_c76 bl[76] br[76] wl[351] vdd gnd cell_6t
Xbit_r352_c76 bl[76] br[76] wl[352] vdd gnd cell_6t
Xbit_r353_c76 bl[76] br[76] wl[353] vdd gnd cell_6t
Xbit_r354_c76 bl[76] br[76] wl[354] vdd gnd cell_6t
Xbit_r355_c76 bl[76] br[76] wl[355] vdd gnd cell_6t
Xbit_r356_c76 bl[76] br[76] wl[356] vdd gnd cell_6t
Xbit_r357_c76 bl[76] br[76] wl[357] vdd gnd cell_6t
Xbit_r358_c76 bl[76] br[76] wl[358] vdd gnd cell_6t
Xbit_r359_c76 bl[76] br[76] wl[359] vdd gnd cell_6t
Xbit_r360_c76 bl[76] br[76] wl[360] vdd gnd cell_6t
Xbit_r361_c76 bl[76] br[76] wl[361] vdd gnd cell_6t
Xbit_r362_c76 bl[76] br[76] wl[362] vdd gnd cell_6t
Xbit_r363_c76 bl[76] br[76] wl[363] vdd gnd cell_6t
Xbit_r364_c76 bl[76] br[76] wl[364] vdd gnd cell_6t
Xbit_r365_c76 bl[76] br[76] wl[365] vdd gnd cell_6t
Xbit_r366_c76 bl[76] br[76] wl[366] vdd gnd cell_6t
Xbit_r367_c76 bl[76] br[76] wl[367] vdd gnd cell_6t
Xbit_r368_c76 bl[76] br[76] wl[368] vdd gnd cell_6t
Xbit_r369_c76 bl[76] br[76] wl[369] vdd gnd cell_6t
Xbit_r370_c76 bl[76] br[76] wl[370] vdd gnd cell_6t
Xbit_r371_c76 bl[76] br[76] wl[371] vdd gnd cell_6t
Xbit_r372_c76 bl[76] br[76] wl[372] vdd gnd cell_6t
Xbit_r373_c76 bl[76] br[76] wl[373] vdd gnd cell_6t
Xbit_r374_c76 bl[76] br[76] wl[374] vdd gnd cell_6t
Xbit_r375_c76 bl[76] br[76] wl[375] vdd gnd cell_6t
Xbit_r376_c76 bl[76] br[76] wl[376] vdd gnd cell_6t
Xbit_r377_c76 bl[76] br[76] wl[377] vdd gnd cell_6t
Xbit_r378_c76 bl[76] br[76] wl[378] vdd gnd cell_6t
Xbit_r379_c76 bl[76] br[76] wl[379] vdd gnd cell_6t
Xbit_r380_c76 bl[76] br[76] wl[380] vdd gnd cell_6t
Xbit_r381_c76 bl[76] br[76] wl[381] vdd gnd cell_6t
Xbit_r382_c76 bl[76] br[76] wl[382] vdd gnd cell_6t
Xbit_r383_c76 bl[76] br[76] wl[383] vdd gnd cell_6t
Xbit_r384_c76 bl[76] br[76] wl[384] vdd gnd cell_6t
Xbit_r385_c76 bl[76] br[76] wl[385] vdd gnd cell_6t
Xbit_r386_c76 bl[76] br[76] wl[386] vdd gnd cell_6t
Xbit_r387_c76 bl[76] br[76] wl[387] vdd gnd cell_6t
Xbit_r388_c76 bl[76] br[76] wl[388] vdd gnd cell_6t
Xbit_r389_c76 bl[76] br[76] wl[389] vdd gnd cell_6t
Xbit_r390_c76 bl[76] br[76] wl[390] vdd gnd cell_6t
Xbit_r391_c76 bl[76] br[76] wl[391] vdd gnd cell_6t
Xbit_r392_c76 bl[76] br[76] wl[392] vdd gnd cell_6t
Xbit_r393_c76 bl[76] br[76] wl[393] vdd gnd cell_6t
Xbit_r394_c76 bl[76] br[76] wl[394] vdd gnd cell_6t
Xbit_r395_c76 bl[76] br[76] wl[395] vdd gnd cell_6t
Xbit_r396_c76 bl[76] br[76] wl[396] vdd gnd cell_6t
Xbit_r397_c76 bl[76] br[76] wl[397] vdd gnd cell_6t
Xbit_r398_c76 bl[76] br[76] wl[398] vdd gnd cell_6t
Xbit_r399_c76 bl[76] br[76] wl[399] vdd gnd cell_6t
Xbit_r400_c76 bl[76] br[76] wl[400] vdd gnd cell_6t
Xbit_r401_c76 bl[76] br[76] wl[401] vdd gnd cell_6t
Xbit_r402_c76 bl[76] br[76] wl[402] vdd gnd cell_6t
Xbit_r403_c76 bl[76] br[76] wl[403] vdd gnd cell_6t
Xbit_r404_c76 bl[76] br[76] wl[404] vdd gnd cell_6t
Xbit_r405_c76 bl[76] br[76] wl[405] vdd gnd cell_6t
Xbit_r406_c76 bl[76] br[76] wl[406] vdd gnd cell_6t
Xbit_r407_c76 bl[76] br[76] wl[407] vdd gnd cell_6t
Xbit_r408_c76 bl[76] br[76] wl[408] vdd gnd cell_6t
Xbit_r409_c76 bl[76] br[76] wl[409] vdd gnd cell_6t
Xbit_r410_c76 bl[76] br[76] wl[410] vdd gnd cell_6t
Xbit_r411_c76 bl[76] br[76] wl[411] vdd gnd cell_6t
Xbit_r412_c76 bl[76] br[76] wl[412] vdd gnd cell_6t
Xbit_r413_c76 bl[76] br[76] wl[413] vdd gnd cell_6t
Xbit_r414_c76 bl[76] br[76] wl[414] vdd gnd cell_6t
Xbit_r415_c76 bl[76] br[76] wl[415] vdd gnd cell_6t
Xbit_r416_c76 bl[76] br[76] wl[416] vdd gnd cell_6t
Xbit_r417_c76 bl[76] br[76] wl[417] vdd gnd cell_6t
Xbit_r418_c76 bl[76] br[76] wl[418] vdd gnd cell_6t
Xbit_r419_c76 bl[76] br[76] wl[419] vdd gnd cell_6t
Xbit_r420_c76 bl[76] br[76] wl[420] vdd gnd cell_6t
Xbit_r421_c76 bl[76] br[76] wl[421] vdd gnd cell_6t
Xbit_r422_c76 bl[76] br[76] wl[422] vdd gnd cell_6t
Xbit_r423_c76 bl[76] br[76] wl[423] vdd gnd cell_6t
Xbit_r424_c76 bl[76] br[76] wl[424] vdd gnd cell_6t
Xbit_r425_c76 bl[76] br[76] wl[425] vdd gnd cell_6t
Xbit_r426_c76 bl[76] br[76] wl[426] vdd gnd cell_6t
Xbit_r427_c76 bl[76] br[76] wl[427] vdd gnd cell_6t
Xbit_r428_c76 bl[76] br[76] wl[428] vdd gnd cell_6t
Xbit_r429_c76 bl[76] br[76] wl[429] vdd gnd cell_6t
Xbit_r430_c76 bl[76] br[76] wl[430] vdd gnd cell_6t
Xbit_r431_c76 bl[76] br[76] wl[431] vdd gnd cell_6t
Xbit_r432_c76 bl[76] br[76] wl[432] vdd gnd cell_6t
Xbit_r433_c76 bl[76] br[76] wl[433] vdd gnd cell_6t
Xbit_r434_c76 bl[76] br[76] wl[434] vdd gnd cell_6t
Xbit_r435_c76 bl[76] br[76] wl[435] vdd gnd cell_6t
Xbit_r436_c76 bl[76] br[76] wl[436] vdd gnd cell_6t
Xbit_r437_c76 bl[76] br[76] wl[437] vdd gnd cell_6t
Xbit_r438_c76 bl[76] br[76] wl[438] vdd gnd cell_6t
Xbit_r439_c76 bl[76] br[76] wl[439] vdd gnd cell_6t
Xbit_r440_c76 bl[76] br[76] wl[440] vdd gnd cell_6t
Xbit_r441_c76 bl[76] br[76] wl[441] vdd gnd cell_6t
Xbit_r442_c76 bl[76] br[76] wl[442] vdd gnd cell_6t
Xbit_r443_c76 bl[76] br[76] wl[443] vdd gnd cell_6t
Xbit_r444_c76 bl[76] br[76] wl[444] vdd gnd cell_6t
Xbit_r445_c76 bl[76] br[76] wl[445] vdd gnd cell_6t
Xbit_r446_c76 bl[76] br[76] wl[446] vdd gnd cell_6t
Xbit_r447_c76 bl[76] br[76] wl[447] vdd gnd cell_6t
Xbit_r448_c76 bl[76] br[76] wl[448] vdd gnd cell_6t
Xbit_r449_c76 bl[76] br[76] wl[449] vdd gnd cell_6t
Xbit_r450_c76 bl[76] br[76] wl[450] vdd gnd cell_6t
Xbit_r451_c76 bl[76] br[76] wl[451] vdd gnd cell_6t
Xbit_r452_c76 bl[76] br[76] wl[452] vdd gnd cell_6t
Xbit_r453_c76 bl[76] br[76] wl[453] vdd gnd cell_6t
Xbit_r454_c76 bl[76] br[76] wl[454] vdd gnd cell_6t
Xbit_r455_c76 bl[76] br[76] wl[455] vdd gnd cell_6t
Xbit_r456_c76 bl[76] br[76] wl[456] vdd gnd cell_6t
Xbit_r457_c76 bl[76] br[76] wl[457] vdd gnd cell_6t
Xbit_r458_c76 bl[76] br[76] wl[458] vdd gnd cell_6t
Xbit_r459_c76 bl[76] br[76] wl[459] vdd gnd cell_6t
Xbit_r460_c76 bl[76] br[76] wl[460] vdd gnd cell_6t
Xbit_r461_c76 bl[76] br[76] wl[461] vdd gnd cell_6t
Xbit_r462_c76 bl[76] br[76] wl[462] vdd gnd cell_6t
Xbit_r463_c76 bl[76] br[76] wl[463] vdd gnd cell_6t
Xbit_r464_c76 bl[76] br[76] wl[464] vdd gnd cell_6t
Xbit_r465_c76 bl[76] br[76] wl[465] vdd gnd cell_6t
Xbit_r466_c76 bl[76] br[76] wl[466] vdd gnd cell_6t
Xbit_r467_c76 bl[76] br[76] wl[467] vdd gnd cell_6t
Xbit_r468_c76 bl[76] br[76] wl[468] vdd gnd cell_6t
Xbit_r469_c76 bl[76] br[76] wl[469] vdd gnd cell_6t
Xbit_r470_c76 bl[76] br[76] wl[470] vdd gnd cell_6t
Xbit_r471_c76 bl[76] br[76] wl[471] vdd gnd cell_6t
Xbit_r472_c76 bl[76] br[76] wl[472] vdd gnd cell_6t
Xbit_r473_c76 bl[76] br[76] wl[473] vdd gnd cell_6t
Xbit_r474_c76 bl[76] br[76] wl[474] vdd gnd cell_6t
Xbit_r475_c76 bl[76] br[76] wl[475] vdd gnd cell_6t
Xbit_r476_c76 bl[76] br[76] wl[476] vdd gnd cell_6t
Xbit_r477_c76 bl[76] br[76] wl[477] vdd gnd cell_6t
Xbit_r478_c76 bl[76] br[76] wl[478] vdd gnd cell_6t
Xbit_r479_c76 bl[76] br[76] wl[479] vdd gnd cell_6t
Xbit_r480_c76 bl[76] br[76] wl[480] vdd gnd cell_6t
Xbit_r481_c76 bl[76] br[76] wl[481] vdd gnd cell_6t
Xbit_r482_c76 bl[76] br[76] wl[482] vdd gnd cell_6t
Xbit_r483_c76 bl[76] br[76] wl[483] vdd gnd cell_6t
Xbit_r484_c76 bl[76] br[76] wl[484] vdd gnd cell_6t
Xbit_r485_c76 bl[76] br[76] wl[485] vdd gnd cell_6t
Xbit_r486_c76 bl[76] br[76] wl[486] vdd gnd cell_6t
Xbit_r487_c76 bl[76] br[76] wl[487] vdd gnd cell_6t
Xbit_r488_c76 bl[76] br[76] wl[488] vdd gnd cell_6t
Xbit_r489_c76 bl[76] br[76] wl[489] vdd gnd cell_6t
Xbit_r490_c76 bl[76] br[76] wl[490] vdd gnd cell_6t
Xbit_r491_c76 bl[76] br[76] wl[491] vdd gnd cell_6t
Xbit_r492_c76 bl[76] br[76] wl[492] vdd gnd cell_6t
Xbit_r493_c76 bl[76] br[76] wl[493] vdd gnd cell_6t
Xbit_r494_c76 bl[76] br[76] wl[494] vdd gnd cell_6t
Xbit_r495_c76 bl[76] br[76] wl[495] vdd gnd cell_6t
Xbit_r496_c76 bl[76] br[76] wl[496] vdd gnd cell_6t
Xbit_r497_c76 bl[76] br[76] wl[497] vdd gnd cell_6t
Xbit_r498_c76 bl[76] br[76] wl[498] vdd gnd cell_6t
Xbit_r499_c76 bl[76] br[76] wl[499] vdd gnd cell_6t
Xbit_r500_c76 bl[76] br[76] wl[500] vdd gnd cell_6t
Xbit_r501_c76 bl[76] br[76] wl[501] vdd gnd cell_6t
Xbit_r502_c76 bl[76] br[76] wl[502] vdd gnd cell_6t
Xbit_r503_c76 bl[76] br[76] wl[503] vdd gnd cell_6t
Xbit_r504_c76 bl[76] br[76] wl[504] vdd gnd cell_6t
Xbit_r505_c76 bl[76] br[76] wl[505] vdd gnd cell_6t
Xbit_r506_c76 bl[76] br[76] wl[506] vdd gnd cell_6t
Xbit_r507_c76 bl[76] br[76] wl[507] vdd gnd cell_6t
Xbit_r508_c76 bl[76] br[76] wl[508] vdd gnd cell_6t
Xbit_r509_c76 bl[76] br[76] wl[509] vdd gnd cell_6t
Xbit_r510_c76 bl[76] br[76] wl[510] vdd gnd cell_6t
Xbit_r511_c76 bl[76] br[76] wl[511] vdd gnd cell_6t
Xbit_r0_c77 bl[77] br[77] wl[0] vdd gnd cell_6t
Xbit_r1_c77 bl[77] br[77] wl[1] vdd gnd cell_6t
Xbit_r2_c77 bl[77] br[77] wl[2] vdd gnd cell_6t
Xbit_r3_c77 bl[77] br[77] wl[3] vdd gnd cell_6t
Xbit_r4_c77 bl[77] br[77] wl[4] vdd gnd cell_6t
Xbit_r5_c77 bl[77] br[77] wl[5] vdd gnd cell_6t
Xbit_r6_c77 bl[77] br[77] wl[6] vdd gnd cell_6t
Xbit_r7_c77 bl[77] br[77] wl[7] vdd gnd cell_6t
Xbit_r8_c77 bl[77] br[77] wl[8] vdd gnd cell_6t
Xbit_r9_c77 bl[77] br[77] wl[9] vdd gnd cell_6t
Xbit_r10_c77 bl[77] br[77] wl[10] vdd gnd cell_6t
Xbit_r11_c77 bl[77] br[77] wl[11] vdd gnd cell_6t
Xbit_r12_c77 bl[77] br[77] wl[12] vdd gnd cell_6t
Xbit_r13_c77 bl[77] br[77] wl[13] vdd gnd cell_6t
Xbit_r14_c77 bl[77] br[77] wl[14] vdd gnd cell_6t
Xbit_r15_c77 bl[77] br[77] wl[15] vdd gnd cell_6t
Xbit_r16_c77 bl[77] br[77] wl[16] vdd gnd cell_6t
Xbit_r17_c77 bl[77] br[77] wl[17] vdd gnd cell_6t
Xbit_r18_c77 bl[77] br[77] wl[18] vdd gnd cell_6t
Xbit_r19_c77 bl[77] br[77] wl[19] vdd gnd cell_6t
Xbit_r20_c77 bl[77] br[77] wl[20] vdd gnd cell_6t
Xbit_r21_c77 bl[77] br[77] wl[21] vdd gnd cell_6t
Xbit_r22_c77 bl[77] br[77] wl[22] vdd gnd cell_6t
Xbit_r23_c77 bl[77] br[77] wl[23] vdd gnd cell_6t
Xbit_r24_c77 bl[77] br[77] wl[24] vdd gnd cell_6t
Xbit_r25_c77 bl[77] br[77] wl[25] vdd gnd cell_6t
Xbit_r26_c77 bl[77] br[77] wl[26] vdd gnd cell_6t
Xbit_r27_c77 bl[77] br[77] wl[27] vdd gnd cell_6t
Xbit_r28_c77 bl[77] br[77] wl[28] vdd gnd cell_6t
Xbit_r29_c77 bl[77] br[77] wl[29] vdd gnd cell_6t
Xbit_r30_c77 bl[77] br[77] wl[30] vdd gnd cell_6t
Xbit_r31_c77 bl[77] br[77] wl[31] vdd gnd cell_6t
Xbit_r32_c77 bl[77] br[77] wl[32] vdd gnd cell_6t
Xbit_r33_c77 bl[77] br[77] wl[33] vdd gnd cell_6t
Xbit_r34_c77 bl[77] br[77] wl[34] vdd gnd cell_6t
Xbit_r35_c77 bl[77] br[77] wl[35] vdd gnd cell_6t
Xbit_r36_c77 bl[77] br[77] wl[36] vdd gnd cell_6t
Xbit_r37_c77 bl[77] br[77] wl[37] vdd gnd cell_6t
Xbit_r38_c77 bl[77] br[77] wl[38] vdd gnd cell_6t
Xbit_r39_c77 bl[77] br[77] wl[39] vdd gnd cell_6t
Xbit_r40_c77 bl[77] br[77] wl[40] vdd gnd cell_6t
Xbit_r41_c77 bl[77] br[77] wl[41] vdd gnd cell_6t
Xbit_r42_c77 bl[77] br[77] wl[42] vdd gnd cell_6t
Xbit_r43_c77 bl[77] br[77] wl[43] vdd gnd cell_6t
Xbit_r44_c77 bl[77] br[77] wl[44] vdd gnd cell_6t
Xbit_r45_c77 bl[77] br[77] wl[45] vdd gnd cell_6t
Xbit_r46_c77 bl[77] br[77] wl[46] vdd gnd cell_6t
Xbit_r47_c77 bl[77] br[77] wl[47] vdd gnd cell_6t
Xbit_r48_c77 bl[77] br[77] wl[48] vdd gnd cell_6t
Xbit_r49_c77 bl[77] br[77] wl[49] vdd gnd cell_6t
Xbit_r50_c77 bl[77] br[77] wl[50] vdd gnd cell_6t
Xbit_r51_c77 bl[77] br[77] wl[51] vdd gnd cell_6t
Xbit_r52_c77 bl[77] br[77] wl[52] vdd gnd cell_6t
Xbit_r53_c77 bl[77] br[77] wl[53] vdd gnd cell_6t
Xbit_r54_c77 bl[77] br[77] wl[54] vdd gnd cell_6t
Xbit_r55_c77 bl[77] br[77] wl[55] vdd gnd cell_6t
Xbit_r56_c77 bl[77] br[77] wl[56] vdd gnd cell_6t
Xbit_r57_c77 bl[77] br[77] wl[57] vdd gnd cell_6t
Xbit_r58_c77 bl[77] br[77] wl[58] vdd gnd cell_6t
Xbit_r59_c77 bl[77] br[77] wl[59] vdd gnd cell_6t
Xbit_r60_c77 bl[77] br[77] wl[60] vdd gnd cell_6t
Xbit_r61_c77 bl[77] br[77] wl[61] vdd gnd cell_6t
Xbit_r62_c77 bl[77] br[77] wl[62] vdd gnd cell_6t
Xbit_r63_c77 bl[77] br[77] wl[63] vdd gnd cell_6t
Xbit_r64_c77 bl[77] br[77] wl[64] vdd gnd cell_6t
Xbit_r65_c77 bl[77] br[77] wl[65] vdd gnd cell_6t
Xbit_r66_c77 bl[77] br[77] wl[66] vdd gnd cell_6t
Xbit_r67_c77 bl[77] br[77] wl[67] vdd gnd cell_6t
Xbit_r68_c77 bl[77] br[77] wl[68] vdd gnd cell_6t
Xbit_r69_c77 bl[77] br[77] wl[69] vdd gnd cell_6t
Xbit_r70_c77 bl[77] br[77] wl[70] vdd gnd cell_6t
Xbit_r71_c77 bl[77] br[77] wl[71] vdd gnd cell_6t
Xbit_r72_c77 bl[77] br[77] wl[72] vdd gnd cell_6t
Xbit_r73_c77 bl[77] br[77] wl[73] vdd gnd cell_6t
Xbit_r74_c77 bl[77] br[77] wl[74] vdd gnd cell_6t
Xbit_r75_c77 bl[77] br[77] wl[75] vdd gnd cell_6t
Xbit_r76_c77 bl[77] br[77] wl[76] vdd gnd cell_6t
Xbit_r77_c77 bl[77] br[77] wl[77] vdd gnd cell_6t
Xbit_r78_c77 bl[77] br[77] wl[78] vdd gnd cell_6t
Xbit_r79_c77 bl[77] br[77] wl[79] vdd gnd cell_6t
Xbit_r80_c77 bl[77] br[77] wl[80] vdd gnd cell_6t
Xbit_r81_c77 bl[77] br[77] wl[81] vdd gnd cell_6t
Xbit_r82_c77 bl[77] br[77] wl[82] vdd gnd cell_6t
Xbit_r83_c77 bl[77] br[77] wl[83] vdd gnd cell_6t
Xbit_r84_c77 bl[77] br[77] wl[84] vdd gnd cell_6t
Xbit_r85_c77 bl[77] br[77] wl[85] vdd gnd cell_6t
Xbit_r86_c77 bl[77] br[77] wl[86] vdd gnd cell_6t
Xbit_r87_c77 bl[77] br[77] wl[87] vdd gnd cell_6t
Xbit_r88_c77 bl[77] br[77] wl[88] vdd gnd cell_6t
Xbit_r89_c77 bl[77] br[77] wl[89] vdd gnd cell_6t
Xbit_r90_c77 bl[77] br[77] wl[90] vdd gnd cell_6t
Xbit_r91_c77 bl[77] br[77] wl[91] vdd gnd cell_6t
Xbit_r92_c77 bl[77] br[77] wl[92] vdd gnd cell_6t
Xbit_r93_c77 bl[77] br[77] wl[93] vdd gnd cell_6t
Xbit_r94_c77 bl[77] br[77] wl[94] vdd gnd cell_6t
Xbit_r95_c77 bl[77] br[77] wl[95] vdd gnd cell_6t
Xbit_r96_c77 bl[77] br[77] wl[96] vdd gnd cell_6t
Xbit_r97_c77 bl[77] br[77] wl[97] vdd gnd cell_6t
Xbit_r98_c77 bl[77] br[77] wl[98] vdd gnd cell_6t
Xbit_r99_c77 bl[77] br[77] wl[99] vdd gnd cell_6t
Xbit_r100_c77 bl[77] br[77] wl[100] vdd gnd cell_6t
Xbit_r101_c77 bl[77] br[77] wl[101] vdd gnd cell_6t
Xbit_r102_c77 bl[77] br[77] wl[102] vdd gnd cell_6t
Xbit_r103_c77 bl[77] br[77] wl[103] vdd gnd cell_6t
Xbit_r104_c77 bl[77] br[77] wl[104] vdd gnd cell_6t
Xbit_r105_c77 bl[77] br[77] wl[105] vdd gnd cell_6t
Xbit_r106_c77 bl[77] br[77] wl[106] vdd gnd cell_6t
Xbit_r107_c77 bl[77] br[77] wl[107] vdd gnd cell_6t
Xbit_r108_c77 bl[77] br[77] wl[108] vdd gnd cell_6t
Xbit_r109_c77 bl[77] br[77] wl[109] vdd gnd cell_6t
Xbit_r110_c77 bl[77] br[77] wl[110] vdd gnd cell_6t
Xbit_r111_c77 bl[77] br[77] wl[111] vdd gnd cell_6t
Xbit_r112_c77 bl[77] br[77] wl[112] vdd gnd cell_6t
Xbit_r113_c77 bl[77] br[77] wl[113] vdd gnd cell_6t
Xbit_r114_c77 bl[77] br[77] wl[114] vdd gnd cell_6t
Xbit_r115_c77 bl[77] br[77] wl[115] vdd gnd cell_6t
Xbit_r116_c77 bl[77] br[77] wl[116] vdd gnd cell_6t
Xbit_r117_c77 bl[77] br[77] wl[117] vdd gnd cell_6t
Xbit_r118_c77 bl[77] br[77] wl[118] vdd gnd cell_6t
Xbit_r119_c77 bl[77] br[77] wl[119] vdd gnd cell_6t
Xbit_r120_c77 bl[77] br[77] wl[120] vdd gnd cell_6t
Xbit_r121_c77 bl[77] br[77] wl[121] vdd gnd cell_6t
Xbit_r122_c77 bl[77] br[77] wl[122] vdd gnd cell_6t
Xbit_r123_c77 bl[77] br[77] wl[123] vdd gnd cell_6t
Xbit_r124_c77 bl[77] br[77] wl[124] vdd gnd cell_6t
Xbit_r125_c77 bl[77] br[77] wl[125] vdd gnd cell_6t
Xbit_r126_c77 bl[77] br[77] wl[126] vdd gnd cell_6t
Xbit_r127_c77 bl[77] br[77] wl[127] vdd gnd cell_6t
Xbit_r128_c77 bl[77] br[77] wl[128] vdd gnd cell_6t
Xbit_r129_c77 bl[77] br[77] wl[129] vdd gnd cell_6t
Xbit_r130_c77 bl[77] br[77] wl[130] vdd gnd cell_6t
Xbit_r131_c77 bl[77] br[77] wl[131] vdd gnd cell_6t
Xbit_r132_c77 bl[77] br[77] wl[132] vdd gnd cell_6t
Xbit_r133_c77 bl[77] br[77] wl[133] vdd gnd cell_6t
Xbit_r134_c77 bl[77] br[77] wl[134] vdd gnd cell_6t
Xbit_r135_c77 bl[77] br[77] wl[135] vdd gnd cell_6t
Xbit_r136_c77 bl[77] br[77] wl[136] vdd gnd cell_6t
Xbit_r137_c77 bl[77] br[77] wl[137] vdd gnd cell_6t
Xbit_r138_c77 bl[77] br[77] wl[138] vdd gnd cell_6t
Xbit_r139_c77 bl[77] br[77] wl[139] vdd gnd cell_6t
Xbit_r140_c77 bl[77] br[77] wl[140] vdd gnd cell_6t
Xbit_r141_c77 bl[77] br[77] wl[141] vdd gnd cell_6t
Xbit_r142_c77 bl[77] br[77] wl[142] vdd gnd cell_6t
Xbit_r143_c77 bl[77] br[77] wl[143] vdd gnd cell_6t
Xbit_r144_c77 bl[77] br[77] wl[144] vdd gnd cell_6t
Xbit_r145_c77 bl[77] br[77] wl[145] vdd gnd cell_6t
Xbit_r146_c77 bl[77] br[77] wl[146] vdd gnd cell_6t
Xbit_r147_c77 bl[77] br[77] wl[147] vdd gnd cell_6t
Xbit_r148_c77 bl[77] br[77] wl[148] vdd gnd cell_6t
Xbit_r149_c77 bl[77] br[77] wl[149] vdd gnd cell_6t
Xbit_r150_c77 bl[77] br[77] wl[150] vdd gnd cell_6t
Xbit_r151_c77 bl[77] br[77] wl[151] vdd gnd cell_6t
Xbit_r152_c77 bl[77] br[77] wl[152] vdd gnd cell_6t
Xbit_r153_c77 bl[77] br[77] wl[153] vdd gnd cell_6t
Xbit_r154_c77 bl[77] br[77] wl[154] vdd gnd cell_6t
Xbit_r155_c77 bl[77] br[77] wl[155] vdd gnd cell_6t
Xbit_r156_c77 bl[77] br[77] wl[156] vdd gnd cell_6t
Xbit_r157_c77 bl[77] br[77] wl[157] vdd gnd cell_6t
Xbit_r158_c77 bl[77] br[77] wl[158] vdd gnd cell_6t
Xbit_r159_c77 bl[77] br[77] wl[159] vdd gnd cell_6t
Xbit_r160_c77 bl[77] br[77] wl[160] vdd gnd cell_6t
Xbit_r161_c77 bl[77] br[77] wl[161] vdd gnd cell_6t
Xbit_r162_c77 bl[77] br[77] wl[162] vdd gnd cell_6t
Xbit_r163_c77 bl[77] br[77] wl[163] vdd gnd cell_6t
Xbit_r164_c77 bl[77] br[77] wl[164] vdd gnd cell_6t
Xbit_r165_c77 bl[77] br[77] wl[165] vdd gnd cell_6t
Xbit_r166_c77 bl[77] br[77] wl[166] vdd gnd cell_6t
Xbit_r167_c77 bl[77] br[77] wl[167] vdd gnd cell_6t
Xbit_r168_c77 bl[77] br[77] wl[168] vdd gnd cell_6t
Xbit_r169_c77 bl[77] br[77] wl[169] vdd gnd cell_6t
Xbit_r170_c77 bl[77] br[77] wl[170] vdd gnd cell_6t
Xbit_r171_c77 bl[77] br[77] wl[171] vdd gnd cell_6t
Xbit_r172_c77 bl[77] br[77] wl[172] vdd gnd cell_6t
Xbit_r173_c77 bl[77] br[77] wl[173] vdd gnd cell_6t
Xbit_r174_c77 bl[77] br[77] wl[174] vdd gnd cell_6t
Xbit_r175_c77 bl[77] br[77] wl[175] vdd gnd cell_6t
Xbit_r176_c77 bl[77] br[77] wl[176] vdd gnd cell_6t
Xbit_r177_c77 bl[77] br[77] wl[177] vdd gnd cell_6t
Xbit_r178_c77 bl[77] br[77] wl[178] vdd gnd cell_6t
Xbit_r179_c77 bl[77] br[77] wl[179] vdd gnd cell_6t
Xbit_r180_c77 bl[77] br[77] wl[180] vdd gnd cell_6t
Xbit_r181_c77 bl[77] br[77] wl[181] vdd gnd cell_6t
Xbit_r182_c77 bl[77] br[77] wl[182] vdd gnd cell_6t
Xbit_r183_c77 bl[77] br[77] wl[183] vdd gnd cell_6t
Xbit_r184_c77 bl[77] br[77] wl[184] vdd gnd cell_6t
Xbit_r185_c77 bl[77] br[77] wl[185] vdd gnd cell_6t
Xbit_r186_c77 bl[77] br[77] wl[186] vdd gnd cell_6t
Xbit_r187_c77 bl[77] br[77] wl[187] vdd gnd cell_6t
Xbit_r188_c77 bl[77] br[77] wl[188] vdd gnd cell_6t
Xbit_r189_c77 bl[77] br[77] wl[189] vdd gnd cell_6t
Xbit_r190_c77 bl[77] br[77] wl[190] vdd gnd cell_6t
Xbit_r191_c77 bl[77] br[77] wl[191] vdd gnd cell_6t
Xbit_r192_c77 bl[77] br[77] wl[192] vdd gnd cell_6t
Xbit_r193_c77 bl[77] br[77] wl[193] vdd gnd cell_6t
Xbit_r194_c77 bl[77] br[77] wl[194] vdd gnd cell_6t
Xbit_r195_c77 bl[77] br[77] wl[195] vdd gnd cell_6t
Xbit_r196_c77 bl[77] br[77] wl[196] vdd gnd cell_6t
Xbit_r197_c77 bl[77] br[77] wl[197] vdd gnd cell_6t
Xbit_r198_c77 bl[77] br[77] wl[198] vdd gnd cell_6t
Xbit_r199_c77 bl[77] br[77] wl[199] vdd gnd cell_6t
Xbit_r200_c77 bl[77] br[77] wl[200] vdd gnd cell_6t
Xbit_r201_c77 bl[77] br[77] wl[201] vdd gnd cell_6t
Xbit_r202_c77 bl[77] br[77] wl[202] vdd gnd cell_6t
Xbit_r203_c77 bl[77] br[77] wl[203] vdd gnd cell_6t
Xbit_r204_c77 bl[77] br[77] wl[204] vdd gnd cell_6t
Xbit_r205_c77 bl[77] br[77] wl[205] vdd gnd cell_6t
Xbit_r206_c77 bl[77] br[77] wl[206] vdd gnd cell_6t
Xbit_r207_c77 bl[77] br[77] wl[207] vdd gnd cell_6t
Xbit_r208_c77 bl[77] br[77] wl[208] vdd gnd cell_6t
Xbit_r209_c77 bl[77] br[77] wl[209] vdd gnd cell_6t
Xbit_r210_c77 bl[77] br[77] wl[210] vdd gnd cell_6t
Xbit_r211_c77 bl[77] br[77] wl[211] vdd gnd cell_6t
Xbit_r212_c77 bl[77] br[77] wl[212] vdd gnd cell_6t
Xbit_r213_c77 bl[77] br[77] wl[213] vdd gnd cell_6t
Xbit_r214_c77 bl[77] br[77] wl[214] vdd gnd cell_6t
Xbit_r215_c77 bl[77] br[77] wl[215] vdd gnd cell_6t
Xbit_r216_c77 bl[77] br[77] wl[216] vdd gnd cell_6t
Xbit_r217_c77 bl[77] br[77] wl[217] vdd gnd cell_6t
Xbit_r218_c77 bl[77] br[77] wl[218] vdd gnd cell_6t
Xbit_r219_c77 bl[77] br[77] wl[219] vdd gnd cell_6t
Xbit_r220_c77 bl[77] br[77] wl[220] vdd gnd cell_6t
Xbit_r221_c77 bl[77] br[77] wl[221] vdd gnd cell_6t
Xbit_r222_c77 bl[77] br[77] wl[222] vdd gnd cell_6t
Xbit_r223_c77 bl[77] br[77] wl[223] vdd gnd cell_6t
Xbit_r224_c77 bl[77] br[77] wl[224] vdd gnd cell_6t
Xbit_r225_c77 bl[77] br[77] wl[225] vdd gnd cell_6t
Xbit_r226_c77 bl[77] br[77] wl[226] vdd gnd cell_6t
Xbit_r227_c77 bl[77] br[77] wl[227] vdd gnd cell_6t
Xbit_r228_c77 bl[77] br[77] wl[228] vdd gnd cell_6t
Xbit_r229_c77 bl[77] br[77] wl[229] vdd gnd cell_6t
Xbit_r230_c77 bl[77] br[77] wl[230] vdd gnd cell_6t
Xbit_r231_c77 bl[77] br[77] wl[231] vdd gnd cell_6t
Xbit_r232_c77 bl[77] br[77] wl[232] vdd gnd cell_6t
Xbit_r233_c77 bl[77] br[77] wl[233] vdd gnd cell_6t
Xbit_r234_c77 bl[77] br[77] wl[234] vdd gnd cell_6t
Xbit_r235_c77 bl[77] br[77] wl[235] vdd gnd cell_6t
Xbit_r236_c77 bl[77] br[77] wl[236] vdd gnd cell_6t
Xbit_r237_c77 bl[77] br[77] wl[237] vdd gnd cell_6t
Xbit_r238_c77 bl[77] br[77] wl[238] vdd gnd cell_6t
Xbit_r239_c77 bl[77] br[77] wl[239] vdd gnd cell_6t
Xbit_r240_c77 bl[77] br[77] wl[240] vdd gnd cell_6t
Xbit_r241_c77 bl[77] br[77] wl[241] vdd gnd cell_6t
Xbit_r242_c77 bl[77] br[77] wl[242] vdd gnd cell_6t
Xbit_r243_c77 bl[77] br[77] wl[243] vdd gnd cell_6t
Xbit_r244_c77 bl[77] br[77] wl[244] vdd gnd cell_6t
Xbit_r245_c77 bl[77] br[77] wl[245] vdd gnd cell_6t
Xbit_r246_c77 bl[77] br[77] wl[246] vdd gnd cell_6t
Xbit_r247_c77 bl[77] br[77] wl[247] vdd gnd cell_6t
Xbit_r248_c77 bl[77] br[77] wl[248] vdd gnd cell_6t
Xbit_r249_c77 bl[77] br[77] wl[249] vdd gnd cell_6t
Xbit_r250_c77 bl[77] br[77] wl[250] vdd gnd cell_6t
Xbit_r251_c77 bl[77] br[77] wl[251] vdd gnd cell_6t
Xbit_r252_c77 bl[77] br[77] wl[252] vdd gnd cell_6t
Xbit_r253_c77 bl[77] br[77] wl[253] vdd gnd cell_6t
Xbit_r254_c77 bl[77] br[77] wl[254] vdd gnd cell_6t
Xbit_r255_c77 bl[77] br[77] wl[255] vdd gnd cell_6t
Xbit_r256_c77 bl[77] br[77] wl[256] vdd gnd cell_6t
Xbit_r257_c77 bl[77] br[77] wl[257] vdd gnd cell_6t
Xbit_r258_c77 bl[77] br[77] wl[258] vdd gnd cell_6t
Xbit_r259_c77 bl[77] br[77] wl[259] vdd gnd cell_6t
Xbit_r260_c77 bl[77] br[77] wl[260] vdd gnd cell_6t
Xbit_r261_c77 bl[77] br[77] wl[261] vdd gnd cell_6t
Xbit_r262_c77 bl[77] br[77] wl[262] vdd gnd cell_6t
Xbit_r263_c77 bl[77] br[77] wl[263] vdd gnd cell_6t
Xbit_r264_c77 bl[77] br[77] wl[264] vdd gnd cell_6t
Xbit_r265_c77 bl[77] br[77] wl[265] vdd gnd cell_6t
Xbit_r266_c77 bl[77] br[77] wl[266] vdd gnd cell_6t
Xbit_r267_c77 bl[77] br[77] wl[267] vdd gnd cell_6t
Xbit_r268_c77 bl[77] br[77] wl[268] vdd gnd cell_6t
Xbit_r269_c77 bl[77] br[77] wl[269] vdd gnd cell_6t
Xbit_r270_c77 bl[77] br[77] wl[270] vdd gnd cell_6t
Xbit_r271_c77 bl[77] br[77] wl[271] vdd gnd cell_6t
Xbit_r272_c77 bl[77] br[77] wl[272] vdd gnd cell_6t
Xbit_r273_c77 bl[77] br[77] wl[273] vdd gnd cell_6t
Xbit_r274_c77 bl[77] br[77] wl[274] vdd gnd cell_6t
Xbit_r275_c77 bl[77] br[77] wl[275] vdd gnd cell_6t
Xbit_r276_c77 bl[77] br[77] wl[276] vdd gnd cell_6t
Xbit_r277_c77 bl[77] br[77] wl[277] vdd gnd cell_6t
Xbit_r278_c77 bl[77] br[77] wl[278] vdd gnd cell_6t
Xbit_r279_c77 bl[77] br[77] wl[279] vdd gnd cell_6t
Xbit_r280_c77 bl[77] br[77] wl[280] vdd gnd cell_6t
Xbit_r281_c77 bl[77] br[77] wl[281] vdd gnd cell_6t
Xbit_r282_c77 bl[77] br[77] wl[282] vdd gnd cell_6t
Xbit_r283_c77 bl[77] br[77] wl[283] vdd gnd cell_6t
Xbit_r284_c77 bl[77] br[77] wl[284] vdd gnd cell_6t
Xbit_r285_c77 bl[77] br[77] wl[285] vdd gnd cell_6t
Xbit_r286_c77 bl[77] br[77] wl[286] vdd gnd cell_6t
Xbit_r287_c77 bl[77] br[77] wl[287] vdd gnd cell_6t
Xbit_r288_c77 bl[77] br[77] wl[288] vdd gnd cell_6t
Xbit_r289_c77 bl[77] br[77] wl[289] vdd gnd cell_6t
Xbit_r290_c77 bl[77] br[77] wl[290] vdd gnd cell_6t
Xbit_r291_c77 bl[77] br[77] wl[291] vdd gnd cell_6t
Xbit_r292_c77 bl[77] br[77] wl[292] vdd gnd cell_6t
Xbit_r293_c77 bl[77] br[77] wl[293] vdd gnd cell_6t
Xbit_r294_c77 bl[77] br[77] wl[294] vdd gnd cell_6t
Xbit_r295_c77 bl[77] br[77] wl[295] vdd gnd cell_6t
Xbit_r296_c77 bl[77] br[77] wl[296] vdd gnd cell_6t
Xbit_r297_c77 bl[77] br[77] wl[297] vdd gnd cell_6t
Xbit_r298_c77 bl[77] br[77] wl[298] vdd gnd cell_6t
Xbit_r299_c77 bl[77] br[77] wl[299] vdd gnd cell_6t
Xbit_r300_c77 bl[77] br[77] wl[300] vdd gnd cell_6t
Xbit_r301_c77 bl[77] br[77] wl[301] vdd gnd cell_6t
Xbit_r302_c77 bl[77] br[77] wl[302] vdd gnd cell_6t
Xbit_r303_c77 bl[77] br[77] wl[303] vdd gnd cell_6t
Xbit_r304_c77 bl[77] br[77] wl[304] vdd gnd cell_6t
Xbit_r305_c77 bl[77] br[77] wl[305] vdd gnd cell_6t
Xbit_r306_c77 bl[77] br[77] wl[306] vdd gnd cell_6t
Xbit_r307_c77 bl[77] br[77] wl[307] vdd gnd cell_6t
Xbit_r308_c77 bl[77] br[77] wl[308] vdd gnd cell_6t
Xbit_r309_c77 bl[77] br[77] wl[309] vdd gnd cell_6t
Xbit_r310_c77 bl[77] br[77] wl[310] vdd gnd cell_6t
Xbit_r311_c77 bl[77] br[77] wl[311] vdd gnd cell_6t
Xbit_r312_c77 bl[77] br[77] wl[312] vdd gnd cell_6t
Xbit_r313_c77 bl[77] br[77] wl[313] vdd gnd cell_6t
Xbit_r314_c77 bl[77] br[77] wl[314] vdd gnd cell_6t
Xbit_r315_c77 bl[77] br[77] wl[315] vdd gnd cell_6t
Xbit_r316_c77 bl[77] br[77] wl[316] vdd gnd cell_6t
Xbit_r317_c77 bl[77] br[77] wl[317] vdd gnd cell_6t
Xbit_r318_c77 bl[77] br[77] wl[318] vdd gnd cell_6t
Xbit_r319_c77 bl[77] br[77] wl[319] vdd gnd cell_6t
Xbit_r320_c77 bl[77] br[77] wl[320] vdd gnd cell_6t
Xbit_r321_c77 bl[77] br[77] wl[321] vdd gnd cell_6t
Xbit_r322_c77 bl[77] br[77] wl[322] vdd gnd cell_6t
Xbit_r323_c77 bl[77] br[77] wl[323] vdd gnd cell_6t
Xbit_r324_c77 bl[77] br[77] wl[324] vdd gnd cell_6t
Xbit_r325_c77 bl[77] br[77] wl[325] vdd gnd cell_6t
Xbit_r326_c77 bl[77] br[77] wl[326] vdd gnd cell_6t
Xbit_r327_c77 bl[77] br[77] wl[327] vdd gnd cell_6t
Xbit_r328_c77 bl[77] br[77] wl[328] vdd gnd cell_6t
Xbit_r329_c77 bl[77] br[77] wl[329] vdd gnd cell_6t
Xbit_r330_c77 bl[77] br[77] wl[330] vdd gnd cell_6t
Xbit_r331_c77 bl[77] br[77] wl[331] vdd gnd cell_6t
Xbit_r332_c77 bl[77] br[77] wl[332] vdd gnd cell_6t
Xbit_r333_c77 bl[77] br[77] wl[333] vdd gnd cell_6t
Xbit_r334_c77 bl[77] br[77] wl[334] vdd gnd cell_6t
Xbit_r335_c77 bl[77] br[77] wl[335] vdd gnd cell_6t
Xbit_r336_c77 bl[77] br[77] wl[336] vdd gnd cell_6t
Xbit_r337_c77 bl[77] br[77] wl[337] vdd gnd cell_6t
Xbit_r338_c77 bl[77] br[77] wl[338] vdd gnd cell_6t
Xbit_r339_c77 bl[77] br[77] wl[339] vdd gnd cell_6t
Xbit_r340_c77 bl[77] br[77] wl[340] vdd gnd cell_6t
Xbit_r341_c77 bl[77] br[77] wl[341] vdd gnd cell_6t
Xbit_r342_c77 bl[77] br[77] wl[342] vdd gnd cell_6t
Xbit_r343_c77 bl[77] br[77] wl[343] vdd gnd cell_6t
Xbit_r344_c77 bl[77] br[77] wl[344] vdd gnd cell_6t
Xbit_r345_c77 bl[77] br[77] wl[345] vdd gnd cell_6t
Xbit_r346_c77 bl[77] br[77] wl[346] vdd gnd cell_6t
Xbit_r347_c77 bl[77] br[77] wl[347] vdd gnd cell_6t
Xbit_r348_c77 bl[77] br[77] wl[348] vdd gnd cell_6t
Xbit_r349_c77 bl[77] br[77] wl[349] vdd gnd cell_6t
Xbit_r350_c77 bl[77] br[77] wl[350] vdd gnd cell_6t
Xbit_r351_c77 bl[77] br[77] wl[351] vdd gnd cell_6t
Xbit_r352_c77 bl[77] br[77] wl[352] vdd gnd cell_6t
Xbit_r353_c77 bl[77] br[77] wl[353] vdd gnd cell_6t
Xbit_r354_c77 bl[77] br[77] wl[354] vdd gnd cell_6t
Xbit_r355_c77 bl[77] br[77] wl[355] vdd gnd cell_6t
Xbit_r356_c77 bl[77] br[77] wl[356] vdd gnd cell_6t
Xbit_r357_c77 bl[77] br[77] wl[357] vdd gnd cell_6t
Xbit_r358_c77 bl[77] br[77] wl[358] vdd gnd cell_6t
Xbit_r359_c77 bl[77] br[77] wl[359] vdd gnd cell_6t
Xbit_r360_c77 bl[77] br[77] wl[360] vdd gnd cell_6t
Xbit_r361_c77 bl[77] br[77] wl[361] vdd gnd cell_6t
Xbit_r362_c77 bl[77] br[77] wl[362] vdd gnd cell_6t
Xbit_r363_c77 bl[77] br[77] wl[363] vdd gnd cell_6t
Xbit_r364_c77 bl[77] br[77] wl[364] vdd gnd cell_6t
Xbit_r365_c77 bl[77] br[77] wl[365] vdd gnd cell_6t
Xbit_r366_c77 bl[77] br[77] wl[366] vdd gnd cell_6t
Xbit_r367_c77 bl[77] br[77] wl[367] vdd gnd cell_6t
Xbit_r368_c77 bl[77] br[77] wl[368] vdd gnd cell_6t
Xbit_r369_c77 bl[77] br[77] wl[369] vdd gnd cell_6t
Xbit_r370_c77 bl[77] br[77] wl[370] vdd gnd cell_6t
Xbit_r371_c77 bl[77] br[77] wl[371] vdd gnd cell_6t
Xbit_r372_c77 bl[77] br[77] wl[372] vdd gnd cell_6t
Xbit_r373_c77 bl[77] br[77] wl[373] vdd gnd cell_6t
Xbit_r374_c77 bl[77] br[77] wl[374] vdd gnd cell_6t
Xbit_r375_c77 bl[77] br[77] wl[375] vdd gnd cell_6t
Xbit_r376_c77 bl[77] br[77] wl[376] vdd gnd cell_6t
Xbit_r377_c77 bl[77] br[77] wl[377] vdd gnd cell_6t
Xbit_r378_c77 bl[77] br[77] wl[378] vdd gnd cell_6t
Xbit_r379_c77 bl[77] br[77] wl[379] vdd gnd cell_6t
Xbit_r380_c77 bl[77] br[77] wl[380] vdd gnd cell_6t
Xbit_r381_c77 bl[77] br[77] wl[381] vdd gnd cell_6t
Xbit_r382_c77 bl[77] br[77] wl[382] vdd gnd cell_6t
Xbit_r383_c77 bl[77] br[77] wl[383] vdd gnd cell_6t
Xbit_r384_c77 bl[77] br[77] wl[384] vdd gnd cell_6t
Xbit_r385_c77 bl[77] br[77] wl[385] vdd gnd cell_6t
Xbit_r386_c77 bl[77] br[77] wl[386] vdd gnd cell_6t
Xbit_r387_c77 bl[77] br[77] wl[387] vdd gnd cell_6t
Xbit_r388_c77 bl[77] br[77] wl[388] vdd gnd cell_6t
Xbit_r389_c77 bl[77] br[77] wl[389] vdd gnd cell_6t
Xbit_r390_c77 bl[77] br[77] wl[390] vdd gnd cell_6t
Xbit_r391_c77 bl[77] br[77] wl[391] vdd gnd cell_6t
Xbit_r392_c77 bl[77] br[77] wl[392] vdd gnd cell_6t
Xbit_r393_c77 bl[77] br[77] wl[393] vdd gnd cell_6t
Xbit_r394_c77 bl[77] br[77] wl[394] vdd gnd cell_6t
Xbit_r395_c77 bl[77] br[77] wl[395] vdd gnd cell_6t
Xbit_r396_c77 bl[77] br[77] wl[396] vdd gnd cell_6t
Xbit_r397_c77 bl[77] br[77] wl[397] vdd gnd cell_6t
Xbit_r398_c77 bl[77] br[77] wl[398] vdd gnd cell_6t
Xbit_r399_c77 bl[77] br[77] wl[399] vdd gnd cell_6t
Xbit_r400_c77 bl[77] br[77] wl[400] vdd gnd cell_6t
Xbit_r401_c77 bl[77] br[77] wl[401] vdd gnd cell_6t
Xbit_r402_c77 bl[77] br[77] wl[402] vdd gnd cell_6t
Xbit_r403_c77 bl[77] br[77] wl[403] vdd gnd cell_6t
Xbit_r404_c77 bl[77] br[77] wl[404] vdd gnd cell_6t
Xbit_r405_c77 bl[77] br[77] wl[405] vdd gnd cell_6t
Xbit_r406_c77 bl[77] br[77] wl[406] vdd gnd cell_6t
Xbit_r407_c77 bl[77] br[77] wl[407] vdd gnd cell_6t
Xbit_r408_c77 bl[77] br[77] wl[408] vdd gnd cell_6t
Xbit_r409_c77 bl[77] br[77] wl[409] vdd gnd cell_6t
Xbit_r410_c77 bl[77] br[77] wl[410] vdd gnd cell_6t
Xbit_r411_c77 bl[77] br[77] wl[411] vdd gnd cell_6t
Xbit_r412_c77 bl[77] br[77] wl[412] vdd gnd cell_6t
Xbit_r413_c77 bl[77] br[77] wl[413] vdd gnd cell_6t
Xbit_r414_c77 bl[77] br[77] wl[414] vdd gnd cell_6t
Xbit_r415_c77 bl[77] br[77] wl[415] vdd gnd cell_6t
Xbit_r416_c77 bl[77] br[77] wl[416] vdd gnd cell_6t
Xbit_r417_c77 bl[77] br[77] wl[417] vdd gnd cell_6t
Xbit_r418_c77 bl[77] br[77] wl[418] vdd gnd cell_6t
Xbit_r419_c77 bl[77] br[77] wl[419] vdd gnd cell_6t
Xbit_r420_c77 bl[77] br[77] wl[420] vdd gnd cell_6t
Xbit_r421_c77 bl[77] br[77] wl[421] vdd gnd cell_6t
Xbit_r422_c77 bl[77] br[77] wl[422] vdd gnd cell_6t
Xbit_r423_c77 bl[77] br[77] wl[423] vdd gnd cell_6t
Xbit_r424_c77 bl[77] br[77] wl[424] vdd gnd cell_6t
Xbit_r425_c77 bl[77] br[77] wl[425] vdd gnd cell_6t
Xbit_r426_c77 bl[77] br[77] wl[426] vdd gnd cell_6t
Xbit_r427_c77 bl[77] br[77] wl[427] vdd gnd cell_6t
Xbit_r428_c77 bl[77] br[77] wl[428] vdd gnd cell_6t
Xbit_r429_c77 bl[77] br[77] wl[429] vdd gnd cell_6t
Xbit_r430_c77 bl[77] br[77] wl[430] vdd gnd cell_6t
Xbit_r431_c77 bl[77] br[77] wl[431] vdd gnd cell_6t
Xbit_r432_c77 bl[77] br[77] wl[432] vdd gnd cell_6t
Xbit_r433_c77 bl[77] br[77] wl[433] vdd gnd cell_6t
Xbit_r434_c77 bl[77] br[77] wl[434] vdd gnd cell_6t
Xbit_r435_c77 bl[77] br[77] wl[435] vdd gnd cell_6t
Xbit_r436_c77 bl[77] br[77] wl[436] vdd gnd cell_6t
Xbit_r437_c77 bl[77] br[77] wl[437] vdd gnd cell_6t
Xbit_r438_c77 bl[77] br[77] wl[438] vdd gnd cell_6t
Xbit_r439_c77 bl[77] br[77] wl[439] vdd gnd cell_6t
Xbit_r440_c77 bl[77] br[77] wl[440] vdd gnd cell_6t
Xbit_r441_c77 bl[77] br[77] wl[441] vdd gnd cell_6t
Xbit_r442_c77 bl[77] br[77] wl[442] vdd gnd cell_6t
Xbit_r443_c77 bl[77] br[77] wl[443] vdd gnd cell_6t
Xbit_r444_c77 bl[77] br[77] wl[444] vdd gnd cell_6t
Xbit_r445_c77 bl[77] br[77] wl[445] vdd gnd cell_6t
Xbit_r446_c77 bl[77] br[77] wl[446] vdd gnd cell_6t
Xbit_r447_c77 bl[77] br[77] wl[447] vdd gnd cell_6t
Xbit_r448_c77 bl[77] br[77] wl[448] vdd gnd cell_6t
Xbit_r449_c77 bl[77] br[77] wl[449] vdd gnd cell_6t
Xbit_r450_c77 bl[77] br[77] wl[450] vdd gnd cell_6t
Xbit_r451_c77 bl[77] br[77] wl[451] vdd gnd cell_6t
Xbit_r452_c77 bl[77] br[77] wl[452] vdd gnd cell_6t
Xbit_r453_c77 bl[77] br[77] wl[453] vdd gnd cell_6t
Xbit_r454_c77 bl[77] br[77] wl[454] vdd gnd cell_6t
Xbit_r455_c77 bl[77] br[77] wl[455] vdd gnd cell_6t
Xbit_r456_c77 bl[77] br[77] wl[456] vdd gnd cell_6t
Xbit_r457_c77 bl[77] br[77] wl[457] vdd gnd cell_6t
Xbit_r458_c77 bl[77] br[77] wl[458] vdd gnd cell_6t
Xbit_r459_c77 bl[77] br[77] wl[459] vdd gnd cell_6t
Xbit_r460_c77 bl[77] br[77] wl[460] vdd gnd cell_6t
Xbit_r461_c77 bl[77] br[77] wl[461] vdd gnd cell_6t
Xbit_r462_c77 bl[77] br[77] wl[462] vdd gnd cell_6t
Xbit_r463_c77 bl[77] br[77] wl[463] vdd gnd cell_6t
Xbit_r464_c77 bl[77] br[77] wl[464] vdd gnd cell_6t
Xbit_r465_c77 bl[77] br[77] wl[465] vdd gnd cell_6t
Xbit_r466_c77 bl[77] br[77] wl[466] vdd gnd cell_6t
Xbit_r467_c77 bl[77] br[77] wl[467] vdd gnd cell_6t
Xbit_r468_c77 bl[77] br[77] wl[468] vdd gnd cell_6t
Xbit_r469_c77 bl[77] br[77] wl[469] vdd gnd cell_6t
Xbit_r470_c77 bl[77] br[77] wl[470] vdd gnd cell_6t
Xbit_r471_c77 bl[77] br[77] wl[471] vdd gnd cell_6t
Xbit_r472_c77 bl[77] br[77] wl[472] vdd gnd cell_6t
Xbit_r473_c77 bl[77] br[77] wl[473] vdd gnd cell_6t
Xbit_r474_c77 bl[77] br[77] wl[474] vdd gnd cell_6t
Xbit_r475_c77 bl[77] br[77] wl[475] vdd gnd cell_6t
Xbit_r476_c77 bl[77] br[77] wl[476] vdd gnd cell_6t
Xbit_r477_c77 bl[77] br[77] wl[477] vdd gnd cell_6t
Xbit_r478_c77 bl[77] br[77] wl[478] vdd gnd cell_6t
Xbit_r479_c77 bl[77] br[77] wl[479] vdd gnd cell_6t
Xbit_r480_c77 bl[77] br[77] wl[480] vdd gnd cell_6t
Xbit_r481_c77 bl[77] br[77] wl[481] vdd gnd cell_6t
Xbit_r482_c77 bl[77] br[77] wl[482] vdd gnd cell_6t
Xbit_r483_c77 bl[77] br[77] wl[483] vdd gnd cell_6t
Xbit_r484_c77 bl[77] br[77] wl[484] vdd gnd cell_6t
Xbit_r485_c77 bl[77] br[77] wl[485] vdd gnd cell_6t
Xbit_r486_c77 bl[77] br[77] wl[486] vdd gnd cell_6t
Xbit_r487_c77 bl[77] br[77] wl[487] vdd gnd cell_6t
Xbit_r488_c77 bl[77] br[77] wl[488] vdd gnd cell_6t
Xbit_r489_c77 bl[77] br[77] wl[489] vdd gnd cell_6t
Xbit_r490_c77 bl[77] br[77] wl[490] vdd gnd cell_6t
Xbit_r491_c77 bl[77] br[77] wl[491] vdd gnd cell_6t
Xbit_r492_c77 bl[77] br[77] wl[492] vdd gnd cell_6t
Xbit_r493_c77 bl[77] br[77] wl[493] vdd gnd cell_6t
Xbit_r494_c77 bl[77] br[77] wl[494] vdd gnd cell_6t
Xbit_r495_c77 bl[77] br[77] wl[495] vdd gnd cell_6t
Xbit_r496_c77 bl[77] br[77] wl[496] vdd gnd cell_6t
Xbit_r497_c77 bl[77] br[77] wl[497] vdd gnd cell_6t
Xbit_r498_c77 bl[77] br[77] wl[498] vdd gnd cell_6t
Xbit_r499_c77 bl[77] br[77] wl[499] vdd gnd cell_6t
Xbit_r500_c77 bl[77] br[77] wl[500] vdd gnd cell_6t
Xbit_r501_c77 bl[77] br[77] wl[501] vdd gnd cell_6t
Xbit_r502_c77 bl[77] br[77] wl[502] vdd gnd cell_6t
Xbit_r503_c77 bl[77] br[77] wl[503] vdd gnd cell_6t
Xbit_r504_c77 bl[77] br[77] wl[504] vdd gnd cell_6t
Xbit_r505_c77 bl[77] br[77] wl[505] vdd gnd cell_6t
Xbit_r506_c77 bl[77] br[77] wl[506] vdd gnd cell_6t
Xbit_r507_c77 bl[77] br[77] wl[507] vdd gnd cell_6t
Xbit_r508_c77 bl[77] br[77] wl[508] vdd gnd cell_6t
Xbit_r509_c77 bl[77] br[77] wl[509] vdd gnd cell_6t
Xbit_r510_c77 bl[77] br[77] wl[510] vdd gnd cell_6t
Xbit_r511_c77 bl[77] br[77] wl[511] vdd gnd cell_6t
Xbit_r0_c78 bl[78] br[78] wl[0] vdd gnd cell_6t
Xbit_r1_c78 bl[78] br[78] wl[1] vdd gnd cell_6t
Xbit_r2_c78 bl[78] br[78] wl[2] vdd gnd cell_6t
Xbit_r3_c78 bl[78] br[78] wl[3] vdd gnd cell_6t
Xbit_r4_c78 bl[78] br[78] wl[4] vdd gnd cell_6t
Xbit_r5_c78 bl[78] br[78] wl[5] vdd gnd cell_6t
Xbit_r6_c78 bl[78] br[78] wl[6] vdd gnd cell_6t
Xbit_r7_c78 bl[78] br[78] wl[7] vdd gnd cell_6t
Xbit_r8_c78 bl[78] br[78] wl[8] vdd gnd cell_6t
Xbit_r9_c78 bl[78] br[78] wl[9] vdd gnd cell_6t
Xbit_r10_c78 bl[78] br[78] wl[10] vdd gnd cell_6t
Xbit_r11_c78 bl[78] br[78] wl[11] vdd gnd cell_6t
Xbit_r12_c78 bl[78] br[78] wl[12] vdd gnd cell_6t
Xbit_r13_c78 bl[78] br[78] wl[13] vdd gnd cell_6t
Xbit_r14_c78 bl[78] br[78] wl[14] vdd gnd cell_6t
Xbit_r15_c78 bl[78] br[78] wl[15] vdd gnd cell_6t
Xbit_r16_c78 bl[78] br[78] wl[16] vdd gnd cell_6t
Xbit_r17_c78 bl[78] br[78] wl[17] vdd gnd cell_6t
Xbit_r18_c78 bl[78] br[78] wl[18] vdd gnd cell_6t
Xbit_r19_c78 bl[78] br[78] wl[19] vdd gnd cell_6t
Xbit_r20_c78 bl[78] br[78] wl[20] vdd gnd cell_6t
Xbit_r21_c78 bl[78] br[78] wl[21] vdd gnd cell_6t
Xbit_r22_c78 bl[78] br[78] wl[22] vdd gnd cell_6t
Xbit_r23_c78 bl[78] br[78] wl[23] vdd gnd cell_6t
Xbit_r24_c78 bl[78] br[78] wl[24] vdd gnd cell_6t
Xbit_r25_c78 bl[78] br[78] wl[25] vdd gnd cell_6t
Xbit_r26_c78 bl[78] br[78] wl[26] vdd gnd cell_6t
Xbit_r27_c78 bl[78] br[78] wl[27] vdd gnd cell_6t
Xbit_r28_c78 bl[78] br[78] wl[28] vdd gnd cell_6t
Xbit_r29_c78 bl[78] br[78] wl[29] vdd gnd cell_6t
Xbit_r30_c78 bl[78] br[78] wl[30] vdd gnd cell_6t
Xbit_r31_c78 bl[78] br[78] wl[31] vdd gnd cell_6t
Xbit_r32_c78 bl[78] br[78] wl[32] vdd gnd cell_6t
Xbit_r33_c78 bl[78] br[78] wl[33] vdd gnd cell_6t
Xbit_r34_c78 bl[78] br[78] wl[34] vdd gnd cell_6t
Xbit_r35_c78 bl[78] br[78] wl[35] vdd gnd cell_6t
Xbit_r36_c78 bl[78] br[78] wl[36] vdd gnd cell_6t
Xbit_r37_c78 bl[78] br[78] wl[37] vdd gnd cell_6t
Xbit_r38_c78 bl[78] br[78] wl[38] vdd gnd cell_6t
Xbit_r39_c78 bl[78] br[78] wl[39] vdd gnd cell_6t
Xbit_r40_c78 bl[78] br[78] wl[40] vdd gnd cell_6t
Xbit_r41_c78 bl[78] br[78] wl[41] vdd gnd cell_6t
Xbit_r42_c78 bl[78] br[78] wl[42] vdd gnd cell_6t
Xbit_r43_c78 bl[78] br[78] wl[43] vdd gnd cell_6t
Xbit_r44_c78 bl[78] br[78] wl[44] vdd gnd cell_6t
Xbit_r45_c78 bl[78] br[78] wl[45] vdd gnd cell_6t
Xbit_r46_c78 bl[78] br[78] wl[46] vdd gnd cell_6t
Xbit_r47_c78 bl[78] br[78] wl[47] vdd gnd cell_6t
Xbit_r48_c78 bl[78] br[78] wl[48] vdd gnd cell_6t
Xbit_r49_c78 bl[78] br[78] wl[49] vdd gnd cell_6t
Xbit_r50_c78 bl[78] br[78] wl[50] vdd gnd cell_6t
Xbit_r51_c78 bl[78] br[78] wl[51] vdd gnd cell_6t
Xbit_r52_c78 bl[78] br[78] wl[52] vdd gnd cell_6t
Xbit_r53_c78 bl[78] br[78] wl[53] vdd gnd cell_6t
Xbit_r54_c78 bl[78] br[78] wl[54] vdd gnd cell_6t
Xbit_r55_c78 bl[78] br[78] wl[55] vdd gnd cell_6t
Xbit_r56_c78 bl[78] br[78] wl[56] vdd gnd cell_6t
Xbit_r57_c78 bl[78] br[78] wl[57] vdd gnd cell_6t
Xbit_r58_c78 bl[78] br[78] wl[58] vdd gnd cell_6t
Xbit_r59_c78 bl[78] br[78] wl[59] vdd gnd cell_6t
Xbit_r60_c78 bl[78] br[78] wl[60] vdd gnd cell_6t
Xbit_r61_c78 bl[78] br[78] wl[61] vdd gnd cell_6t
Xbit_r62_c78 bl[78] br[78] wl[62] vdd gnd cell_6t
Xbit_r63_c78 bl[78] br[78] wl[63] vdd gnd cell_6t
Xbit_r64_c78 bl[78] br[78] wl[64] vdd gnd cell_6t
Xbit_r65_c78 bl[78] br[78] wl[65] vdd gnd cell_6t
Xbit_r66_c78 bl[78] br[78] wl[66] vdd gnd cell_6t
Xbit_r67_c78 bl[78] br[78] wl[67] vdd gnd cell_6t
Xbit_r68_c78 bl[78] br[78] wl[68] vdd gnd cell_6t
Xbit_r69_c78 bl[78] br[78] wl[69] vdd gnd cell_6t
Xbit_r70_c78 bl[78] br[78] wl[70] vdd gnd cell_6t
Xbit_r71_c78 bl[78] br[78] wl[71] vdd gnd cell_6t
Xbit_r72_c78 bl[78] br[78] wl[72] vdd gnd cell_6t
Xbit_r73_c78 bl[78] br[78] wl[73] vdd gnd cell_6t
Xbit_r74_c78 bl[78] br[78] wl[74] vdd gnd cell_6t
Xbit_r75_c78 bl[78] br[78] wl[75] vdd gnd cell_6t
Xbit_r76_c78 bl[78] br[78] wl[76] vdd gnd cell_6t
Xbit_r77_c78 bl[78] br[78] wl[77] vdd gnd cell_6t
Xbit_r78_c78 bl[78] br[78] wl[78] vdd gnd cell_6t
Xbit_r79_c78 bl[78] br[78] wl[79] vdd gnd cell_6t
Xbit_r80_c78 bl[78] br[78] wl[80] vdd gnd cell_6t
Xbit_r81_c78 bl[78] br[78] wl[81] vdd gnd cell_6t
Xbit_r82_c78 bl[78] br[78] wl[82] vdd gnd cell_6t
Xbit_r83_c78 bl[78] br[78] wl[83] vdd gnd cell_6t
Xbit_r84_c78 bl[78] br[78] wl[84] vdd gnd cell_6t
Xbit_r85_c78 bl[78] br[78] wl[85] vdd gnd cell_6t
Xbit_r86_c78 bl[78] br[78] wl[86] vdd gnd cell_6t
Xbit_r87_c78 bl[78] br[78] wl[87] vdd gnd cell_6t
Xbit_r88_c78 bl[78] br[78] wl[88] vdd gnd cell_6t
Xbit_r89_c78 bl[78] br[78] wl[89] vdd gnd cell_6t
Xbit_r90_c78 bl[78] br[78] wl[90] vdd gnd cell_6t
Xbit_r91_c78 bl[78] br[78] wl[91] vdd gnd cell_6t
Xbit_r92_c78 bl[78] br[78] wl[92] vdd gnd cell_6t
Xbit_r93_c78 bl[78] br[78] wl[93] vdd gnd cell_6t
Xbit_r94_c78 bl[78] br[78] wl[94] vdd gnd cell_6t
Xbit_r95_c78 bl[78] br[78] wl[95] vdd gnd cell_6t
Xbit_r96_c78 bl[78] br[78] wl[96] vdd gnd cell_6t
Xbit_r97_c78 bl[78] br[78] wl[97] vdd gnd cell_6t
Xbit_r98_c78 bl[78] br[78] wl[98] vdd gnd cell_6t
Xbit_r99_c78 bl[78] br[78] wl[99] vdd gnd cell_6t
Xbit_r100_c78 bl[78] br[78] wl[100] vdd gnd cell_6t
Xbit_r101_c78 bl[78] br[78] wl[101] vdd gnd cell_6t
Xbit_r102_c78 bl[78] br[78] wl[102] vdd gnd cell_6t
Xbit_r103_c78 bl[78] br[78] wl[103] vdd gnd cell_6t
Xbit_r104_c78 bl[78] br[78] wl[104] vdd gnd cell_6t
Xbit_r105_c78 bl[78] br[78] wl[105] vdd gnd cell_6t
Xbit_r106_c78 bl[78] br[78] wl[106] vdd gnd cell_6t
Xbit_r107_c78 bl[78] br[78] wl[107] vdd gnd cell_6t
Xbit_r108_c78 bl[78] br[78] wl[108] vdd gnd cell_6t
Xbit_r109_c78 bl[78] br[78] wl[109] vdd gnd cell_6t
Xbit_r110_c78 bl[78] br[78] wl[110] vdd gnd cell_6t
Xbit_r111_c78 bl[78] br[78] wl[111] vdd gnd cell_6t
Xbit_r112_c78 bl[78] br[78] wl[112] vdd gnd cell_6t
Xbit_r113_c78 bl[78] br[78] wl[113] vdd gnd cell_6t
Xbit_r114_c78 bl[78] br[78] wl[114] vdd gnd cell_6t
Xbit_r115_c78 bl[78] br[78] wl[115] vdd gnd cell_6t
Xbit_r116_c78 bl[78] br[78] wl[116] vdd gnd cell_6t
Xbit_r117_c78 bl[78] br[78] wl[117] vdd gnd cell_6t
Xbit_r118_c78 bl[78] br[78] wl[118] vdd gnd cell_6t
Xbit_r119_c78 bl[78] br[78] wl[119] vdd gnd cell_6t
Xbit_r120_c78 bl[78] br[78] wl[120] vdd gnd cell_6t
Xbit_r121_c78 bl[78] br[78] wl[121] vdd gnd cell_6t
Xbit_r122_c78 bl[78] br[78] wl[122] vdd gnd cell_6t
Xbit_r123_c78 bl[78] br[78] wl[123] vdd gnd cell_6t
Xbit_r124_c78 bl[78] br[78] wl[124] vdd gnd cell_6t
Xbit_r125_c78 bl[78] br[78] wl[125] vdd gnd cell_6t
Xbit_r126_c78 bl[78] br[78] wl[126] vdd gnd cell_6t
Xbit_r127_c78 bl[78] br[78] wl[127] vdd gnd cell_6t
Xbit_r128_c78 bl[78] br[78] wl[128] vdd gnd cell_6t
Xbit_r129_c78 bl[78] br[78] wl[129] vdd gnd cell_6t
Xbit_r130_c78 bl[78] br[78] wl[130] vdd gnd cell_6t
Xbit_r131_c78 bl[78] br[78] wl[131] vdd gnd cell_6t
Xbit_r132_c78 bl[78] br[78] wl[132] vdd gnd cell_6t
Xbit_r133_c78 bl[78] br[78] wl[133] vdd gnd cell_6t
Xbit_r134_c78 bl[78] br[78] wl[134] vdd gnd cell_6t
Xbit_r135_c78 bl[78] br[78] wl[135] vdd gnd cell_6t
Xbit_r136_c78 bl[78] br[78] wl[136] vdd gnd cell_6t
Xbit_r137_c78 bl[78] br[78] wl[137] vdd gnd cell_6t
Xbit_r138_c78 bl[78] br[78] wl[138] vdd gnd cell_6t
Xbit_r139_c78 bl[78] br[78] wl[139] vdd gnd cell_6t
Xbit_r140_c78 bl[78] br[78] wl[140] vdd gnd cell_6t
Xbit_r141_c78 bl[78] br[78] wl[141] vdd gnd cell_6t
Xbit_r142_c78 bl[78] br[78] wl[142] vdd gnd cell_6t
Xbit_r143_c78 bl[78] br[78] wl[143] vdd gnd cell_6t
Xbit_r144_c78 bl[78] br[78] wl[144] vdd gnd cell_6t
Xbit_r145_c78 bl[78] br[78] wl[145] vdd gnd cell_6t
Xbit_r146_c78 bl[78] br[78] wl[146] vdd gnd cell_6t
Xbit_r147_c78 bl[78] br[78] wl[147] vdd gnd cell_6t
Xbit_r148_c78 bl[78] br[78] wl[148] vdd gnd cell_6t
Xbit_r149_c78 bl[78] br[78] wl[149] vdd gnd cell_6t
Xbit_r150_c78 bl[78] br[78] wl[150] vdd gnd cell_6t
Xbit_r151_c78 bl[78] br[78] wl[151] vdd gnd cell_6t
Xbit_r152_c78 bl[78] br[78] wl[152] vdd gnd cell_6t
Xbit_r153_c78 bl[78] br[78] wl[153] vdd gnd cell_6t
Xbit_r154_c78 bl[78] br[78] wl[154] vdd gnd cell_6t
Xbit_r155_c78 bl[78] br[78] wl[155] vdd gnd cell_6t
Xbit_r156_c78 bl[78] br[78] wl[156] vdd gnd cell_6t
Xbit_r157_c78 bl[78] br[78] wl[157] vdd gnd cell_6t
Xbit_r158_c78 bl[78] br[78] wl[158] vdd gnd cell_6t
Xbit_r159_c78 bl[78] br[78] wl[159] vdd gnd cell_6t
Xbit_r160_c78 bl[78] br[78] wl[160] vdd gnd cell_6t
Xbit_r161_c78 bl[78] br[78] wl[161] vdd gnd cell_6t
Xbit_r162_c78 bl[78] br[78] wl[162] vdd gnd cell_6t
Xbit_r163_c78 bl[78] br[78] wl[163] vdd gnd cell_6t
Xbit_r164_c78 bl[78] br[78] wl[164] vdd gnd cell_6t
Xbit_r165_c78 bl[78] br[78] wl[165] vdd gnd cell_6t
Xbit_r166_c78 bl[78] br[78] wl[166] vdd gnd cell_6t
Xbit_r167_c78 bl[78] br[78] wl[167] vdd gnd cell_6t
Xbit_r168_c78 bl[78] br[78] wl[168] vdd gnd cell_6t
Xbit_r169_c78 bl[78] br[78] wl[169] vdd gnd cell_6t
Xbit_r170_c78 bl[78] br[78] wl[170] vdd gnd cell_6t
Xbit_r171_c78 bl[78] br[78] wl[171] vdd gnd cell_6t
Xbit_r172_c78 bl[78] br[78] wl[172] vdd gnd cell_6t
Xbit_r173_c78 bl[78] br[78] wl[173] vdd gnd cell_6t
Xbit_r174_c78 bl[78] br[78] wl[174] vdd gnd cell_6t
Xbit_r175_c78 bl[78] br[78] wl[175] vdd gnd cell_6t
Xbit_r176_c78 bl[78] br[78] wl[176] vdd gnd cell_6t
Xbit_r177_c78 bl[78] br[78] wl[177] vdd gnd cell_6t
Xbit_r178_c78 bl[78] br[78] wl[178] vdd gnd cell_6t
Xbit_r179_c78 bl[78] br[78] wl[179] vdd gnd cell_6t
Xbit_r180_c78 bl[78] br[78] wl[180] vdd gnd cell_6t
Xbit_r181_c78 bl[78] br[78] wl[181] vdd gnd cell_6t
Xbit_r182_c78 bl[78] br[78] wl[182] vdd gnd cell_6t
Xbit_r183_c78 bl[78] br[78] wl[183] vdd gnd cell_6t
Xbit_r184_c78 bl[78] br[78] wl[184] vdd gnd cell_6t
Xbit_r185_c78 bl[78] br[78] wl[185] vdd gnd cell_6t
Xbit_r186_c78 bl[78] br[78] wl[186] vdd gnd cell_6t
Xbit_r187_c78 bl[78] br[78] wl[187] vdd gnd cell_6t
Xbit_r188_c78 bl[78] br[78] wl[188] vdd gnd cell_6t
Xbit_r189_c78 bl[78] br[78] wl[189] vdd gnd cell_6t
Xbit_r190_c78 bl[78] br[78] wl[190] vdd gnd cell_6t
Xbit_r191_c78 bl[78] br[78] wl[191] vdd gnd cell_6t
Xbit_r192_c78 bl[78] br[78] wl[192] vdd gnd cell_6t
Xbit_r193_c78 bl[78] br[78] wl[193] vdd gnd cell_6t
Xbit_r194_c78 bl[78] br[78] wl[194] vdd gnd cell_6t
Xbit_r195_c78 bl[78] br[78] wl[195] vdd gnd cell_6t
Xbit_r196_c78 bl[78] br[78] wl[196] vdd gnd cell_6t
Xbit_r197_c78 bl[78] br[78] wl[197] vdd gnd cell_6t
Xbit_r198_c78 bl[78] br[78] wl[198] vdd gnd cell_6t
Xbit_r199_c78 bl[78] br[78] wl[199] vdd gnd cell_6t
Xbit_r200_c78 bl[78] br[78] wl[200] vdd gnd cell_6t
Xbit_r201_c78 bl[78] br[78] wl[201] vdd gnd cell_6t
Xbit_r202_c78 bl[78] br[78] wl[202] vdd gnd cell_6t
Xbit_r203_c78 bl[78] br[78] wl[203] vdd gnd cell_6t
Xbit_r204_c78 bl[78] br[78] wl[204] vdd gnd cell_6t
Xbit_r205_c78 bl[78] br[78] wl[205] vdd gnd cell_6t
Xbit_r206_c78 bl[78] br[78] wl[206] vdd gnd cell_6t
Xbit_r207_c78 bl[78] br[78] wl[207] vdd gnd cell_6t
Xbit_r208_c78 bl[78] br[78] wl[208] vdd gnd cell_6t
Xbit_r209_c78 bl[78] br[78] wl[209] vdd gnd cell_6t
Xbit_r210_c78 bl[78] br[78] wl[210] vdd gnd cell_6t
Xbit_r211_c78 bl[78] br[78] wl[211] vdd gnd cell_6t
Xbit_r212_c78 bl[78] br[78] wl[212] vdd gnd cell_6t
Xbit_r213_c78 bl[78] br[78] wl[213] vdd gnd cell_6t
Xbit_r214_c78 bl[78] br[78] wl[214] vdd gnd cell_6t
Xbit_r215_c78 bl[78] br[78] wl[215] vdd gnd cell_6t
Xbit_r216_c78 bl[78] br[78] wl[216] vdd gnd cell_6t
Xbit_r217_c78 bl[78] br[78] wl[217] vdd gnd cell_6t
Xbit_r218_c78 bl[78] br[78] wl[218] vdd gnd cell_6t
Xbit_r219_c78 bl[78] br[78] wl[219] vdd gnd cell_6t
Xbit_r220_c78 bl[78] br[78] wl[220] vdd gnd cell_6t
Xbit_r221_c78 bl[78] br[78] wl[221] vdd gnd cell_6t
Xbit_r222_c78 bl[78] br[78] wl[222] vdd gnd cell_6t
Xbit_r223_c78 bl[78] br[78] wl[223] vdd gnd cell_6t
Xbit_r224_c78 bl[78] br[78] wl[224] vdd gnd cell_6t
Xbit_r225_c78 bl[78] br[78] wl[225] vdd gnd cell_6t
Xbit_r226_c78 bl[78] br[78] wl[226] vdd gnd cell_6t
Xbit_r227_c78 bl[78] br[78] wl[227] vdd gnd cell_6t
Xbit_r228_c78 bl[78] br[78] wl[228] vdd gnd cell_6t
Xbit_r229_c78 bl[78] br[78] wl[229] vdd gnd cell_6t
Xbit_r230_c78 bl[78] br[78] wl[230] vdd gnd cell_6t
Xbit_r231_c78 bl[78] br[78] wl[231] vdd gnd cell_6t
Xbit_r232_c78 bl[78] br[78] wl[232] vdd gnd cell_6t
Xbit_r233_c78 bl[78] br[78] wl[233] vdd gnd cell_6t
Xbit_r234_c78 bl[78] br[78] wl[234] vdd gnd cell_6t
Xbit_r235_c78 bl[78] br[78] wl[235] vdd gnd cell_6t
Xbit_r236_c78 bl[78] br[78] wl[236] vdd gnd cell_6t
Xbit_r237_c78 bl[78] br[78] wl[237] vdd gnd cell_6t
Xbit_r238_c78 bl[78] br[78] wl[238] vdd gnd cell_6t
Xbit_r239_c78 bl[78] br[78] wl[239] vdd gnd cell_6t
Xbit_r240_c78 bl[78] br[78] wl[240] vdd gnd cell_6t
Xbit_r241_c78 bl[78] br[78] wl[241] vdd gnd cell_6t
Xbit_r242_c78 bl[78] br[78] wl[242] vdd gnd cell_6t
Xbit_r243_c78 bl[78] br[78] wl[243] vdd gnd cell_6t
Xbit_r244_c78 bl[78] br[78] wl[244] vdd gnd cell_6t
Xbit_r245_c78 bl[78] br[78] wl[245] vdd gnd cell_6t
Xbit_r246_c78 bl[78] br[78] wl[246] vdd gnd cell_6t
Xbit_r247_c78 bl[78] br[78] wl[247] vdd gnd cell_6t
Xbit_r248_c78 bl[78] br[78] wl[248] vdd gnd cell_6t
Xbit_r249_c78 bl[78] br[78] wl[249] vdd gnd cell_6t
Xbit_r250_c78 bl[78] br[78] wl[250] vdd gnd cell_6t
Xbit_r251_c78 bl[78] br[78] wl[251] vdd gnd cell_6t
Xbit_r252_c78 bl[78] br[78] wl[252] vdd gnd cell_6t
Xbit_r253_c78 bl[78] br[78] wl[253] vdd gnd cell_6t
Xbit_r254_c78 bl[78] br[78] wl[254] vdd gnd cell_6t
Xbit_r255_c78 bl[78] br[78] wl[255] vdd gnd cell_6t
Xbit_r256_c78 bl[78] br[78] wl[256] vdd gnd cell_6t
Xbit_r257_c78 bl[78] br[78] wl[257] vdd gnd cell_6t
Xbit_r258_c78 bl[78] br[78] wl[258] vdd gnd cell_6t
Xbit_r259_c78 bl[78] br[78] wl[259] vdd gnd cell_6t
Xbit_r260_c78 bl[78] br[78] wl[260] vdd gnd cell_6t
Xbit_r261_c78 bl[78] br[78] wl[261] vdd gnd cell_6t
Xbit_r262_c78 bl[78] br[78] wl[262] vdd gnd cell_6t
Xbit_r263_c78 bl[78] br[78] wl[263] vdd gnd cell_6t
Xbit_r264_c78 bl[78] br[78] wl[264] vdd gnd cell_6t
Xbit_r265_c78 bl[78] br[78] wl[265] vdd gnd cell_6t
Xbit_r266_c78 bl[78] br[78] wl[266] vdd gnd cell_6t
Xbit_r267_c78 bl[78] br[78] wl[267] vdd gnd cell_6t
Xbit_r268_c78 bl[78] br[78] wl[268] vdd gnd cell_6t
Xbit_r269_c78 bl[78] br[78] wl[269] vdd gnd cell_6t
Xbit_r270_c78 bl[78] br[78] wl[270] vdd gnd cell_6t
Xbit_r271_c78 bl[78] br[78] wl[271] vdd gnd cell_6t
Xbit_r272_c78 bl[78] br[78] wl[272] vdd gnd cell_6t
Xbit_r273_c78 bl[78] br[78] wl[273] vdd gnd cell_6t
Xbit_r274_c78 bl[78] br[78] wl[274] vdd gnd cell_6t
Xbit_r275_c78 bl[78] br[78] wl[275] vdd gnd cell_6t
Xbit_r276_c78 bl[78] br[78] wl[276] vdd gnd cell_6t
Xbit_r277_c78 bl[78] br[78] wl[277] vdd gnd cell_6t
Xbit_r278_c78 bl[78] br[78] wl[278] vdd gnd cell_6t
Xbit_r279_c78 bl[78] br[78] wl[279] vdd gnd cell_6t
Xbit_r280_c78 bl[78] br[78] wl[280] vdd gnd cell_6t
Xbit_r281_c78 bl[78] br[78] wl[281] vdd gnd cell_6t
Xbit_r282_c78 bl[78] br[78] wl[282] vdd gnd cell_6t
Xbit_r283_c78 bl[78] br[78] wl[283] vdd gnd cell_6t
Xbit_r284_c78 bl[78] br[78] wl[284] vdd gnd cell_6t
Xbit_r285_c78 bl[78] br[78] wl[285] vdd gnd cell_6t
Xbit_r286_c78 bl[78] br[78] wl[286] vdd gnd cell_6t
Xbit_r287_c78 bl[78] br[78] wl[287] vdd gnd cell_6t
Xbit_r288_c78 bl[78] br[78] wl[288] vdd gnd cell_6t
Xbit_r289_c78 bl[78] br[78] wl[289] vdd gnd cell_6t
Xbit_r290_c78 bl[78] br[78] wl[290] vdd gnd cell_6t
Xbit_r291_c78 bl[78] br[78] wl[291] vdd gnd cell_6t
Xbit_r292_c78 bl[78] br[78] wl[292] vdd gnd cell_6t
Xbit_r293_c78 bl[78] br[78] wl[293] vdd gnd cell_6t
Xbit_r294_c78 bl[78] br[78] wl[294] vdd gnd cell_6t
Xbit_r295_c78 bl[78] br[78] wl[295] vdd gnd cell_6t
Xbit_r296_c78 bl[78] br[78] wl[296] vdd gnd cell_6t
Xbit_r297_c78 bl[78] br[78] wl[297] vdd gnd cell_6t
Xbit_r298_c78 bl[78] br[78] wl[298] vdd gnd cell_6t
Xbit_r299_c78 bl[78] br[78] wl[299] vdd gnd cell_6t
Xbit_r300_c78 bl[78] br[78] wl[300] vdd gnd cell_6t
Xbit_r301_c78 bl[78] br[78] wl[301] vdd gnd cell_6t
Xbit_r302_c78 bl[78] br[78] wl[302] vdd gnd cell_6t
Xbit_r303_c78 bl[78] br[78] wl[303] vdd gnd cell_6t
Xbit_r304_c78 bl[78] br[78] wl[304] vdd gnd cell_6t
Xbit_r305_c78 bl[78] br[78] wl[305] vdd gnd cell_6t
Xbit_r306_c78 bl[78] br[78] wl[306] vdd gnd cell_6t
Xbit_r307_c78 bl[78] br[78] wl[307] vdd gnd cell_6t
Xbit_r308_c78 bl[78] br[78] wl[308] vdd gnd cell_6t
Xbit_r309_c78 bl[78] br[78] wl[309] vdd gnd cell_6t
Xbit_r310_c78 bl[78] br[78] wl[310] vdd gnd cell_6t
Xbit_r311_c78 bl[78] br[78] wl[311] vdd gnd cell_6t
Xbit_r312_c78 bl[78] br[78] wl[312] vdd gnd cell_6t
Xbit_r313_c78 bl[78] br[78] wl[313] vdd gnd cell_6t
Xbit_r314_c78 bl[78] br[78] wl[314] vdd gnd cell_6t
Xbit_r315_c78 bl[78] br[78] wl[315] vdd gnd cell_6t
Xbit_r316_c78 bl[78] br[78] wl[316] vdd gnd cell_6t
Xbit_r317_c78 bl[78] br[78] wl[317] vdd gnd cell_6t
Xbit_r318_c78 bl[78] br[78] wl[318] vdd gnd cell_6t
Xbit_r319_c78 bl[78] br[78] wl[319] vdd gnd cell_6t
Xbit_r320_c78 bl[78] br[78] wl[320] vdd gnd cell_6t
Xbit_r321_c78 bl[78] br[78] wl[321] vdd gnd cell_6t
Xbit_r322_c78 bl[78] br[78] wl[322] vdd gnd cell_6t
Xbit_r323_c78 bl[78] br[78] wl[323] vdd gnd cell_6t
Xbit_r324_c78 bl[78] br[78] wl[324] vdd gnd cell_6t
Xbit_r325_c78 bl[78] br[78] wl[325] vdd gnd cell_6t
Xbit_r326_c78 bl[78] br[78] wl[326] vdd gnd cell_6t
Xbit_r327_c78 bl[78] br[78] wl[327] vdd gnd cell_6t
Xbit_r328_c78 bl[78] br[78] wl[328] vdd gnd cell_6t
Xbit_r329_c78 bl[78] br[78] wl[329] vdd gnd cell_6t
Xbit_r330_c78 bl[78] br[78] wl[330] vdd gnd cell_6t
Xbit_r331_c78 bl[78] br[78] wl[331] vdd gnd cell_6t
Xbit_r332_c78 bl[78] br[78] wl[332] vdd gnd cell_6t
Xbit_r333_c78 bl[78] br[78] wl[333] vdd gnd cell_6t
Xbit_r334_c78 bl[78] br[78] wl[334] vdd gnd cell_6t
Xbit_r335_c78 bl[78] br[78] wl[335] vdd gnd cell_6t
Xbit_r336_c78 bl[78] br[78] wl[336] vdd gnd cell_6t
Xbit_r337_c78 bl[78] br[78] wl[337] vdd gnd cell_6t
Xbit_r338_c78 bl[78] br[78] wl[338] vdd gnd cell_6t
Xbit_r339_c78 bl[78] br[78] wl[339] vdd gnd cell_6t
Xbit_r340_c78 bl[78] br[78] wl[340] vdd gnd cell_6t
Xbit_r341_c78 bl[78] br[78] wl[341] vdd gnd cell_6t
Xbit_r342_c78 bl[78] br[78] wl[342] vdd gnd cell_6t
Xbit_r343_c78 bl[78] br[78] wl[343] vdd gnd cell_6t
Xbit_r344_c78 bl[78] br[78] wl[344] vdd gnd cell_6t
Xbit_r345_c78 bl[78] br[78] wl[345] vdd gnd cell_6t
Xbit_r346_c78 bl[78] br[78] wl[346] vdd gnd cell_6t
Xbit_r347_c78 bl[78] br[78] wl[347] vdd gnd cell_6t
Xbit_r348_c78 bl[78] br[78] wl[348] vdd gnd cell_6t
Xbit_r349_c78 bl[78] br[78] wl[349] vdd gnd cell_6t
Xbit_r350_c78 bl[78] br[78] wl[350] vdd gnd cell_6t
Xbit_r351_c78 bl[78] br[78] wl[351] vdd gnd cell_6t
Xbit_r352_c78 bl[78] br[78] wl[352] vdd gnd cell_6t
Xbit_r353_c78 bl[78] br[78] wl[353] vdd gnd cell_6t
Xbit_r354_c78 bl[78] br[78] wl[354] vdd gnd cell_6t
Xbit_r355_c78 bl[78] br[78] wl[355] vdd gnd cell_6t
Xbit_r356_c78 bl[78] br[78] wl[356] vdd gnd cell_6t
Xbit_r357_c78 bl[78] br[78] wl[357] vdd gnd cell_6t
Xbit_r358_c78 bl[78] br[78] wl[358] vdd gnd cell_6t
Xbit_r359_c78 bl[78] br[78] wl[359] vdd gnd cell_6t
Xbit_r360_c78 bl[78] br[78] wl[360] vdd gnd cell_6t
Xbit_r361_c78 bl[78] br[78] wl[361] vdd gnd cell_6t
Xbit_r362_c78 bl[78] br[78] wl[362] vdd gnd cell_6t
Xbit_r363_c78 bl[78] br[78] wl[363] vdd gnd cell_6t
Xbit_r364_c78 bl[78] br[78] wl[364] vdd gnd cell_6t
Xbit_r365_c78 bl[78] br[78] wl[365] vdd gnd cell_6t
Xbit_r366_c78 bl[78] br[78] wl[366] vdd gnd cell_6t
Xbit_r367_c78 bl[78] br[78] wl[367] vdd gnd cell_6t
Xbit_r368_c78 bl[78] br[78] wl[368] vdd gnd cell_6t
Xbit_r369_c78 bl[78] br[78] wl[369] vdd gnd cell_6t
Xbit_r370_c78 bl[78] br[78] wl[370] vdd gnd cell_6t
Xbit_r371_c78 bl[78] br[78] wl[371] vdd gnd cell_6t
Xbit_r372_c78 bl[78] br[78] wl[372] vdd gnd cell_6t
Xbit_r373_c78 bl[78] br[78] wl[373] vdd gnd cell_6t
Xbit_r374_c78 bl[78] br[78] wl[374] vdd gnd cell_6t
Xbit_r375_c78 bl[78] br[78] wl[375] vdd gnd cell_6t
Xbit_r376_c78 bl[78] br[78] wl[376] vdd gnd cell_6t
Xbit_r377_c78 bl[78] br[78] wl[377] vdd gnd cell_6t
Xbit_r378_c78 bl[78] br[78] wl[378] vdd gnd cell_6t
Xbit_r379_c78 bl[78] br[78] wl[379] vdd gnd cell_6t
Xbit_r380_c78 bl[78] br[78] wl[380] vdd gnd cell_6t
Xbit_r381_c78 bl[78] br[78] wl[381] vdd gnd cell_6t
Xbit_r382_c78 bl[78] br[78] wl[382] vdd gnd cell_6t
Xbit_r383_c78 bl[78] br[78] wl[383] vdd gnd cell_6t
Xbit_r384_c78 bl[78] br[78] wl[384] vdd gnd cell_6t
Xbit_r385_c78 bl[78] br[78] wl[385] vdd gnd cell_6t
Xbit_r386_c78 bl[78] br[78] wl[386] vdd gnd cell_6t
Xbit_r387_c78 bl[78] br[78] wl[387] vdd gnd cell_6t
Xbit_r388_c78 bl[78] br[78] wl[388] vdd gnd cell_6t
Xbit_r389_c78 bl[78] br[78] wl[389] vdd gnd cell_6t
Xbit_r390_c78 bl[78] br[78] wl[390] vdd gnd cell_6t
Xbit_r391_c78 bl[78] br[78] wl[391] vdd gnd cell_6t
Xbit_r392_c78 bl[78] br[78] wl[392] vdd gnd cell_6t
Xbit_r393_c78 bl[78] br[78] wl[393] vdd gnd cell_6t
Xbit_r394_c78 bl[78] br[78] wl[394] vdd gnd cell_6t
Xbit_r395_c78 bl[78] br[78] wl[395] vdd gnd cell_6t
Xbit_r396_c78 bl[78] br[78] wl[396] vdd gnd cell_6t
Xbit_r397_c78 bl[78] br[78] wl[397] vdd gnd cell_6t
Xbit_r398_c78 bl[78] br[78] wl[398] vdd gnd cell_6t
Xbit_r399_c78 bl[78] br[78] wl[399] vdd gnd cell_6t
Xbit_r400_c78 bl[78] br[78] wl[400] vdd gnd cell_6t
Xbit_r401_c78 bl[78] br[78] wl[401] vdd gnd cell_6t
Xbit_r402_c78 bl[78] br[78] wl[402] vdd gnd cell_6t
Xbit_r403_c78 bl[78] br[78] wl[403] vdd gnd cell_6t
Xbit_r404_c78 bl[78] br[78] wl[404] vdd gnd cell_6t
Xbit_r405_c78 bl[78] br[78] wl[405] vdd gnd cell_6t
Xbit_r406_c78 bl[78] br[78] wl[406] vdd gnd cell_6t
Xbit_r407_c78 bl[78] br[78] wl[407] vdd gnd cell_6t
Xbit_r408_c78 bl[78] br[78] wl[408] vdd gnd cell_6t
Xbit_r409_c78 bl[78] br[78] wl[409] vdd gnd cell_6t
Xbit_r410_c78 bl[78] br[78] wl[410] vdd gnd cell_6t
Xbit_r411_c78 bl[78] br[78] wl[411] vdd gnd cell_6t
Xbit_r412_c78 bl[78] br[78] wl[412] vdd gnd cell_6t
Xbit_r413_c78 bl[78] br[78] wl[413] vdd gnd cell_6t
Xbit_r414_c78 bl[78] br[78] wl[414] vdd gnd cell_6t
Xbit_r415_c78 bl[78] br[78] wl[415] vdd gnd cell_6t
Xbit_r416_c78 bl[78] br[78] wl[416] vdd gnd cell_6t
Xbit_r417_c78 bl[78] br[78] wl[417] vdd gnd cell_6t
Xbit_r418_c78 bl[78] br[78] wl[418] vdd gnd cell_6t
Xbit_r419_c78 bl[78] br[78] wl[419] vdd gnd cell_6t
Xbit_r420_c78 bl[78] br[78] wl[420] vdd gnd cell_6t
Xbit_r421_c78 bl[78] br[78] wl[421] vdd gnd cell_6t
Xbit_r422_c78 bl[78] br[78] wl[422] vdd gnd cell_6t
Xbit_r423_c78 bl[78] br[78] wl[423] vdd gnd cell_6t
Xbit_r424_c78 bl[78] br[78] wl[424] vdd gnd cell_6t
Xbit_r425_c78 bl[78] br[78] wl[425] vdd gnd cell_6t
Xbit_r426_c78 bl[78] br[78] wl[426] vdd gnd cell_6t
Xbit_r427_c78 bl[78] br[78] wl[427] vdd gnd cell_6t
Xbit_r428_c78 bl[78] br[78] wl[428] vdd gnd cell_6t
Xbit_r429_c78 bl[78] br[78] wl[429] vdd gnd cell_6t
Xbit_r430_c78 bl[78] br[78] wl[430] vdd gnd cell_6t
Xbit_r431_c78 bl[78] br[78] wl[431] vdd gnd cell_6t
Xbit_r432_c78 bl[78] br[78] wl[432] vdd gnd cell_6t
Xbit_r433_c78 bl[78] br[78] wl[433] vdd gnd cell_6t
Xbit_r434_c78 bl[78] br[78] wl[434] vdd gnd cell_6t
Xbit_r435_c78 bl[78] br[78] wl[435] vdd gnd cell_6t
Xbit_r436_c78 bl[78] br[78] wl[436] vdd gnd cell_6t
Xbit_r437_c78 bl[78] br[78] wl[437] vdd gnd cell_6t
Xbit_r438_c78 bl[78] br[78] wl[438] vdd gnd cell_6t
Xbit_r439_c78 bl[78] br[78] wl[439] vdd gnd cell_6t
Xbit_r440_c78 bl[78] br[78] wl[440] vdd gnd cell_6t
Xbit_r441_c78 bl[78] br[78] wl[441] vdd gnd cell_6t
Xbit_r442_c78 bl[78] br[78] wl[442] vdd gnd cell_6t
Xbit_r443_c78 bl[78] br[78] wl[443] vdd gnd cell_6t
Xbit_r444_c78 bl[78] br[78] wl[444] vdd gnd cell_6t
Xbit_r445_c78 bl[78] br[78] wl[445] vdd gnd cell_6t
Xbit_r446_c78 bl[78] br[78] wl[446] vdd gnd cell_6t
Xbit_r447_c78 bl[78] br[78] wl[447] vdd gnd cell_6t
Xbit_r448_c78 bl[78] br[78] wl[448] vdd gnd cell_6t
Xbit_r449_c78 bl[78] br[78] wl[449] vdd gnd cell_6t
Xbit_r450_c78 bl[78] br[78] wl[450] vdd gnd cell_6t
Xbit_r451_c78 bl[78] br[78] wl[451] vdd gnd cell_6t
Xbit_r452_c78 bl[78] br[78] wl[452] vdd gnd cell_6t
Xbit_r453_c78 bl[78] br[78] wl[453] vdd gnd cell_6t
Xbit_r454_c78 bl[78] br[78] wl[454] vdd gnd cell_6t
Xbit_r455_c78 bl[78] br[78] wl[455] vdd gnd cell_6t
Xbit_r456_c78 bl[78] br[78] wl[456] vdd gnd cell_6t
Xbit_r457_c78 bl[78] br[78] wl[457] vdd gnd cell_6t
Xbit_r458_c78 bl[78] br[78] wl[458] vdd gnd cell_6t
Xbit_r459_c78 bl[78] br[78] wl[459] vdd gnd cell_6t
Xbit_r460_c78 bl[78] br[78] wl[460] vdd gnd cell_6t
Xbit_r461_c78 bl[78] br[78] wl[461] vdd gnd cell_6t
Xbit_r462_c78 bl[78] br[78] wl[462] vdd gnd cell_6t
Xbit_r463_c78 bl[78] br[78] wl[463] vdd gnd cell_6t
Xbit_r464_c78 bl[78] br[78] wl[464] vdd gnd cell_6t
Xbit_r465_c78 bl[78] br[78] wl[465] vdd gnd cell_6t
Xbit_r466_c78 bl[78] br[78] wl[466] vdd gnd cell_6t
Xbit_r467_c78 bl[78] br[78] wl[467] vdd gnd cell_6t
Xbit_r468_c78 bl[78] br[78] wl[468] vdd gnd cell_6t
Xbit_r469_c78 bl[78] br[78] wl[469] vdd gnd cell_6t
Xbit_r470_c78 bl[78] br[78] wl[470] vdd gnd cell_6t
Xbit_r471_c78 bl[78] br[78] wl[471] vdd gnd cell_6t
Xbit_r472_c78 bl[78] br[78] wl[472] vdd gnd cell_6t
Xbit_r473_c78 bl[78] br[78] wl[473] vdd gnd cell_6t
Xbit_r474_c78 bl[78] br[78] wl[474] vdd gnd cell_6t
Xbit_r475_c78 bl[78] br[78] wl[475] vdd gnd cell_6t
Xbit_r476_c78 bl[78] br[78] wl[476] vdd gnd cell_6t
Xbit_r477_c78 bl[78] br[78] wl[477] vdd gnd cell_6t
Xbit_r478_c78 bl[78] br[78] wl[478] vdd gnd cell_6t
Xbit_r479_c78 bl[78] br[78] wl[479] vdd gnd cell_6t
Xbit_r480_c78 bl[78] br[78] wl[480] vdd gnd cell_6t
Xbit_r481_c78 bl[78] br[78] wl[481] vdd gnd cell_6t
Xbit_r482_c78 bl[78] br[78] wl[482] vdd gnd cell_6t
Xbit_r483_c78 bl[78] br[78] wl[483] vdd gnd cell_6t
Xbit_r484_c78 bl[78] br[78] wl[484] vdd gnd cell_6t
Xbit_r485_c78 bl[78] br[78] wl[485] vdd gnd cell_6t
Xbit_r486_c78 bl[78] br[78] wl[486] vdd gnd cell_6t
Xbit_r487_c78 bl[78] br[78] wl[487] vdd gnd cell_6t
Xbit_r488_c78 bl[78] br[78] wl[488] vdd gnd cell_6t
Xbit_r489_c78 bl[78] br[78] wl[489] vdd gnd cell_6t
Xbit_r490_c78 bl[78] br[78] wl[490] vdd gnd cell_6t
Xbit_r491_c78 bl[78] br[78] wl[491] vdd gnd cell_6t
Xbit_r492_c78 bl[78] br[78] wl[492] vdd gnd cell_6t
Xbit_r493_c78 bl[78] br[78] wl[493] vdd gnd cell_6t
Xbit_r494_c78 bl[78] br[78] wl[494] vdd gnd cell_6t
Xbit_r495_c78 bl[78] br[78] wl[495] vdd gnd cell_6t
Xbit_r496_c78 bl[78] br[78] wl[496] vdd gnd cell_6t
Xbit_r497_c78 bl[78] br[78] wl[497] vdd gnd cell_6t
Xbit_r498_c78 bl[78] br[78] wl[498] vdd gnd cell_6t
Xbit_r499_c78 bl[78] br[78] wl[499] vdd gnd cell_6t
Xbit_r500_c78 bl[78] br[78] wl[500] vdd gnd cell_6t
Xbit_r501_c78 bl[78] br[78] wl[501] vdd gnd cell_6t
Xbit_r502_c78 bl[78] br[78] wl[502] vdd gnd cell_6t
Xbit_r503_c78 bl[78] br[78] wl[503] vdd gnd cell_6t
Xbit_r504_c78 bl[78] br[78] wl[504] vdd gnd cell_6t
Xbit_r505_c78 bl[78] br[78] wl[505] vdd gnd cell_6t
Xbit_r506_c78 bl[78] br[78] wl[506] vdd gnd cell_6t
Xbit_r507_c78 bl[78] br[78] wl[507] vdd gnd cell_6t
Xbit_r508_c78 bl[78] br[78] wl[508] vdd gnd cell_6t
Xbit_r509_c78 bl[78] br[78] wl[509] vdd gnd cell_6t
Xbit_r510_c78 bl[78] br[78] wl[510] vdd gnd cell_6t
Xbit_r511_c78 bl[78] br[78] wl[511] vdd gnd cell_6t
Xbit_r0_c79 bl[79] br[79] wl[0] vdd gnd cell_6t
Xbit_r1_c79 bl[79] br[79] wl[1] vdd gnd cell_6t
Xbit_r2_c79 bl[79] br[79] wl[2] vdd gnd cell_6t
Xbit_r3_c79 bl[79] br[79] wl[3] vdd gnd cell_6t
Xbit_r4_c79 bl[79] br[79] wl[4] vdd gnd cell_6t
Xbit_r5_c79 bl[79] br[79] wl[5] vdd gnd cell_6t
Xbit_r6_c79 bl[79] br[79] wl[6] vdd gnd cell_6t
Xbit_r7_c79 bl[79] br[79] wl[7] vdd gnd cell_6t
Xbit_r8_c79 bl[79] br[79] wl[8] vdd gnd cell_6t
Xbit_r9_c79 bl[79] br[79] wl[9] vdd gnd cell_6t
Xbit_r10_c79 bl[79] br[79] wl[10] vdd gnd cell_6t
Xbit_r11_c79 bl[79] br[79] wl[11] vdd gnd cell_6t
Xbit_r12_c79 bl[79] br[79] wl[12] vdd gnd cell_6t
Xbit_r13_c79 bl[79] br[79] wl[13] vdd gnd cell_6t
Xbit_r14_c79 bl[79] br[79] wl[14] vdd gnd cell_6t
Xbit_r15_c79 bl[79] br[79] wl[15] vdd gnd cell_6t
Xbit_r16_c79 bl[79] br[79] wl[16] vdd gnd cell_6t
Xbit_r17_c79 bl[79] br[79] wl[17] vdd gnd cell_6t
Xbit_r18_c79 bl[79] br[79] wl[18] vdd gnd cell_6t
Xbit_r19_c79 bl[79] br[79] wl[19] vdd gnd cell_6t
Xbit_r20_c79 bl[79] br[79] wl[20] vdd gnd cell_6t
Xbit_r21_c79 bl[79] br[79] wl[21] vdd gnd cell_6t
Xbit_r22_c79 bl[79] br[79] wl[22] vdd gnd cell_6t
Xbit_r23_c79 bl[79] br[79] wl[23] vdd gnd cell_6t
Xbit_r24_c79 bl[79] br[79] wl[24] vdd gnd cell_6t
Xbit_r25_c79 bl[79] br[79] wl[25] vdd gnd cell_6t
Xbit_r26_c79 bl[79] br[79] wl[26] vdd gnd cell_6t
Xbit_r27_c79 bl[79] br[79] wl[27] vdd gnd cell_6t
Xbit_r28_c79 bl[79] br[79] wl[28] vdd gnd cell_6t
Xbit_r29_c79 bl[79] br[79] wl[29] vdd gnd cell_6t
Xbit_r30_c79 bl[79] br[79] wl[30] vdd gnd cell_6t
Xbit_r31_c79 bl[79] br[79] wl[31] vdd gnd cell_6t
Xbit_r32_c79 bl[79] br[79] wl[32] vdd gnd cell_6t
Xbit_r33_c79 bl[79] br[79] wl[33] vdd gnd cell_6t
Xbit_r34_c79 bl[79] br[79] wl[34] vdd gnd cell_6t
Xbit_r35_c79 bl[79] br[79] wl[35] vdd gnd cell_6t
Xbit_r36_c79 bl[79] br[79] wl[36] vdd gnd cell_6t
Xbit_r37_c79 bl[79] br[79] wl[37] vdd gnd cell_6t
Xbit_r38_c79 bl[79] br[79] wl[38] vdd gnd cell_6t
Xbit_r39_c79 bl[79] br[79] wl[39] vdd gnd cell_6t
Xbit_r40_c79 bl[79] br[79] wl[40] vdd gnd cell_6t
Xbit_r41_c79 bl[79] br[79] wl[41] vdd gnd cell_6t
Xbit_r42_c79 bl[79] br[79] wl[42] vdd gnd cell_6t
Xbit_r43_c79 bl[79] br[79] wl[43] vdd gnd cell_6t
Xbit_r44_c79 bl[79] br[79] wl[44] vdd gnd cell_6t
Xbit_r45_c79 bl[79] br[79] wl[45] vdd gnd cell_6t
Xbit_r46_c79 bl[79] br[79] wl[46] vdd gnd cell_6t
Xbit_r47_c79 bl[79] br[79] wl[47] vdd gnd cell_6t
Xbit_r48_c79 bl[79] br[79] wl[48] vdd gnd cell_6t
Xbit_r49_c79 bl[79] br[79] wl[49] vdd gnd cell_6t
Xbit_r50_c79 bl[79] br[79] wl[50] vdd gnd cell_6t
Xbit_r51_c79 bl[79] br[79] wl[51] vdd gnd cell_6t
Xbit_r52_c79 bl[79] br[79] wl[52] vdd gnd cell_6t
Xbit_r53_c79 bl[79] br[79] wl[53] vdd gnd cell_6t
Xbit_r54_c79 bl[79] br[79] wl[54] vdd gnd cell_6t
Xbit_r55_c79 bl[79] br[79] wl[55] vdd gnd cell_6t
Xbit_r56_c79 bl[79] br[79] wl[56] vdd gnd cell_6t
Xbit_r57_c79 bl[79] br[79] wl[57] vdd gnd cell_6t
Xbit_r58_c79 bl[79] br[79] wl[58] vdd gnd cell_6t
Xbit_r59_c79 bl[79] br[79] wl[59] vdd gnd cell_6t
Xbit_r60_c79 bl[79] br[79] wl[60] vdd gnd cell_6t
Xbit_r61_c79 bl[79] br[79] wl[61] vdd gnd cell_6t
Xbit_r62_c79 bl[79] br[79] wl[62] vdd gnd cell_6t
Xbit_r63_c79 bl[79] br[79] wl[63] vdd gnd cell_6t
Xbit_r64_c79 bl[79] br[79] wl[64] vdd gnd cell_6t
Xbit_r65_c79 bl[79] br[79] wl[65] vdd gnd cell_6t
Xbit_r66_c79 bl[79] br[79] wl[66] vdd gnd cell_6t
Xbit_r67_c79 bl[79] br[79] wl[67] vdd gnd cell_6t
Xbit_r68_c79 bl[79] br[79] wl[68] vdd gnd cell_6t
Xbit_r69_c79 bl[79] br[79] wl[69] vdd gnd cell_6t
Xbit_r70_c79 bl[79] br[79] wl[70] vdd gnd cell_6t
Xbit_r71_c79 bl[79] br[79] wl[71] vdd gnd cell_6t
Xbit_r72_c79 bl[79] br[79] wl[72] vdd gnd cell_6t
Xbit_r73_c79 bl[79] br[79] wl[73] vdd gnd cell_6t
Xbit_r74_c79 bl[79] br[79] wl[74] vdd gnd cell_6t
Xbit_r75_c79 bl[79] br[79] wl[75] vdd gnd cell_6t
Xbit_r76_c79 bl[79] br[79] wl[76] vdd gnd cell_6t
Xbit_r77_c79 bl[79] br[79] wl[77] vdd gnd cell_6t
Xbit_r78_c79 bl[79] br[79] wl[78] vdd gnd cell_6t
Xbit_r79_c79 bl[79] br[79] wl[79] vdd gnd cell_6t
Xbit_r80_c79 bl[79] br[79] wl[80] vdd gnd cell_6t
Xbit_r81_c79 bl[79] br[79] wl[81] vdd gnd cell_6t
Xbit_r82_c79 bl[79] br[79] wl[82] vdd gnd cell_6t
Xbit_r83_c79 bl[79] br[79] wl[83] vdd gnd cell_6t
Xbit_r84_c79 bl[79] br[79] wl[84] vdd gnd cell_6t
Xbit_r85_c79 bl[79] br[79] wl[85] vdd gnd cell_6t
Xbit_r86_c79 bl[79] br[79] wl[86] vdd gnd cell_6t
Xbit_r87_c79 bl[79] br[79] wl[87] vdd gnd cell_6t
Xbit_r88_c79 bl[79] br[79] wl[88] vdd gnd cell_6t
Xbit_r89_c79 bl[79] br[79] wl[89] vdd gnd cell_6t
Xbit_r90_c79 bl[79] br[79] wl[90] vdd gnd cell_6t
Xbit_r91_c79 bl[79] br[79] wl[91] vdd gnd cell_6t
Xbit_r92_c79 bl[79] br[79] wl[92] vdd gnd cell_6t
Xbit_r93_c79 bl[79] br[79] wl[93] vdd gnd cell_6t
Xbit_r94_c79 bl[79] br[79] wl[94] vdd gnd cell_6t
Xbit_r95_c79 bl[79] br[79] wl[95] vdd gnd cell_6t
Xbit_r96_c79 bl[79] br[79] wl[96] vdd gnd cell_6t
Xbit_r97_c79 bl[79] br[79] wl[97] vdd gnd cell_6t
Xbit_r98_c79 bl[79] br[79] wl[98] vdd gnd cell_6t
Xbit_r99_c79 bl[79] br[79] wl[99] vdd gnd cell_6t
Xbit_r100_c79 bl[79] br[79] wl[100] vdd gnd cell_6t
Xbit_r101_c79 bl[79] br[79] wl[101] vdd gnd cell_6t
Xbit_r102_c79 bl[79] br[79] wl[102] vdd gnd cell_6t
Xbit_r103_c79 bl[79] br[79] wl[103] vdd gnd cell_6t
Xbit_r104_c79 bl[79] br[79] wl[104] vdd gnd cell_6t
Xbit_r105_c79 bl[79] br[79] wl[105] vdd gnd cell_6t
Xbit_r106_c79 bl[79] br[79] wl[106] vdd gnd cell_6t
Xbit_r107_c79 bl[79] br[79] wl[107] vdd gnd cell_6t
Xbit_r108_c79 bl[79] br[79] wl[108] vdd gnd cell_6t
Xbit_r109_c79 bl[79] br[79] wl[109] vdd gnd cell_6t
Xbit_r110_c79 bl[79] br[79] wl[110] vdd gnd cell_6t
Xbit_r111_c79 bl[79] br[79] wl[111] vdd gnd cell_6t
Xbit_r112_c79 bl[79] br[79] wl[112] vdd gnd cell_6t
Xbit_r113_c79 bl[79] br[79] wl[113] vdd gnd cell_6t
Xbit_r114_c79 bl[79] br[79] wl[114] vdd gnd cell_6t
Xbit_r115_c79 bl[79] br[79] wl[115] vdd gnd cell_6t
Xbit_r116_c79 bl[79] br[79] wl[116] vdd gnd cell_6t
Xbit_r117_c79 bl[79] br[79] wl[117] vdd gnd cell_6t
Xbit_r118_c79 bl[79] br[79] wl[118] vdd gnd cell_6t
Xbit_r119_c79 bl[79] br[79] wl[119] vdd gnd cell_6t
Xbit_r120_c79 bl[79] br[79] wl[120] vdd gnd cell_6t
Xbit_r121_c79 bl[79] br[79] wl[121] vdd gnd cell_6t
Xbit_r122_c79 bl[79] br[79] wl[122] vdd gnd cell_6t
Xbit_r123_c79 bl[79] br[79] wl[123] vdd gnd cell_6t
Xbit_r124_c79 bl[79] br[79] wl[124] vdd gnd cell_6t
Xbit_r125_c79 bl[79] br[79] wl[125] vdd gnd cell_6t
Xbit_r126_c79 bl[79] br[79] wl[126] vdd gnd cell_6t
Xbit_r127_c79 bl[79] br[79] wl[127] vdd gnd cell_6t
Xbit_r128_c79 bl[79] br[79] wl[128] vdd gnd cell_6t
Xbit_r129_c79 bl[79] br[79] wl[129] vdd gnd cell_6t
Xbit_r130_c79 bl[79] br[79] wl[130] vdd gnd cell_6t
Xbit_r131_c79 bl[79] br[79] wl[131] vdd gnd cell_6t
Xbit_r132_c79 bl[79] br[79] wl[132] vdd gnd cell_6t
Xbit_r133_c79 bl[79] br[79] wl[133] vdd gnd cell_6t
Xbit_r134_c79 bl[79] br[79] wl[134] vdd gnd cell_6t
Xbit_r135_c79 bl[79] br[79] wl[135] vdd gnd cell_6t
Xbit_r136_c79 bl[79] br[79] wl[136] vdd gnd cell_6t
Xbit_r137_c79 bl[79] br[79] wl[137] vdd gnd cell_6t
Xbit_r138_c79 bl[79] br[79] wl[138] vdd gnd cell_6t
Xbit_r139_c79 bl[79] br[79] wl[139] vdd gnd cell_6t
Xbit_r140_c79 bl[79] br[79] wl[140] vdd gnd cell_6t
Xbit_r141_c79 bl[79] br[79] wl[141] vdd gnd cell_6t
Xbit_r142_c79 bl[79] br[79] wl[142] vdd gnd cell_6t
Xbit_r143_c79 bl[79] br[79] wl[143] vdd gnd cell_6t
Xbit_r144_c79 bl[79] br[79] wl[144] vdd gnd cell_6t
Xbit_r145_c79 bl[79] br[79] wl[145] vdd gnd cell_6t
Xbit_r146_c79 bl[79] br[79] wl[146] vdd gnd cell_6t
Xbit_r147_c79 bl[79] br[79] wl[147] vdd gnd cell_6t
Xbit_r148_c79 bl[79] br[79] wl[148] vdd gnd cell_6t
Xbit_r149_c79 bl[79] br[79] wl[149] vdd gnd cell_6t
Xbit_r150_c79 bl[79] br[79] wl[150] vdd gnd cell_6t
Xbit_r151_c79 bl[79] br[79] wl[151] vdd gnd cell_6t
Xbit_r152_c79 bl[79] br[79] wl[152] vdd gnd cell_6t
Xbit_r153_c79 bl[79] br[79] wl[153] vdd gnd cell_6t
Xbit_r154_c79 bl[79] br[79] wl[154] vdd gnd cell_6t
Xbit_r155_c79 bl[79] br[79] wl[155] vdd gnd cell_6t
Xbit_r156_c79 bl[79] br[79] wl[156] vdd gnd cell_6t
Xbit_r157_c79 bl[79] br[79] wl[157] vdd gnd cell_6t
Xbit_r158_c79 bl[79] br[79] wl[158] vdd gnd cell_6t
Xbit_r159_c79 bl[79] br[79] wl[159] vdd gnd cell_6t
Xbit_r160_c79 bl[79] br[79] wl[160] vdd gnd cell_6t
Xbit_r161_c79 bl[79] br[79] wl[161] vdd gnd cell_6t
Xbit_r162_c79 bl[79] br[79] wl[162] vdd gnd cell_6t
Xbit_r163_c79 bl[79] br[79] wl[163] vdd gnd cell_6t
Xbit_r164_c79 bl[79] br[79] wl[164] vdd gnd cell_6t
Xbit_r165_c79 bl[79] br[79] wl[165] vdd gnd cell_6t
Xbit_r166_c79 bl[79] br[79] wl[166] vdd gnd cell_6t
Xbit_r167_c79 bl[79] br[79] wl[167] vdd gnd cell_6t
Xbit_r168_c79 bl[79] br[79] wl[168] vdd gnd cell_6t
Xbit_r169_c79 bl[79] br[79] wl[169] vdd gnd cell_6t
Xbit_r170_c79 bl[79] br[79] wl[170] vdd gnd cell_6t
Xbit_r171_c79 bl[79] br[79] wl[171] vdd gnd cell_6t
Xbit_r172_c79 bl[79] br[79] wl[172] vdd gnd cell_6t
Xbit_r173_c79 bl[79] br[79] wl[173] vdd gnd cell_6t
Xbit_r174_c79 bl[79] br[79] wl[174] vdd gnd cell_6t
Xbit_r175_c79 bl[79] br[79] wl[175] vdd gnd cell_6t
Xbit_r176_c79 bl[79] br[79] wl[176] vdd gnd cell_6t
Xbit_r177_c79 bl[79] br[79] wl[177] vdd gnd cell_6t
Xbit_r178_c79 bl[79] br[79] wl[178] vdd gnd cell_6t
Xbit_r179_c79 bl[79] br[79] wl[179] vdd gnd cell_6t
Xbit_r180_c79 bl[79] br[79] wl[180] vdd gnd cell_6t
Xbit_r181_c79 bl[79] br[79] wl[181] vdd gnd cell_6t
Xbit_r182_c79 bl[79] br[79] wl[182] vdd gnd cell_6t
Xbit_r183_c79 bl[79] br[79] wl[183] vdd gnd cell_6t
Xbit_r184_c79 bl[79] br[79] wl[184] vdd gnd cell_6t
Xbit_r185_c79 bl[79] br[79] wl[185] vdd gnd cell_6t
Xbit_r186_c79 bl[79] br[79] wl[186] vdd gnd cell_6t
Xbit_r187_c79 bl[79] br[79] wl[187] vdd gnd cell_6t
Xbit_r188_c79 bl[79] br[79] wl[188] vdd gnd cell_6t
Xbit_r189_c79 bl[79] br[79] wl[189] vdd gnd cell_6t
Xbit_r190_c79 bl[79] br[79] wl[190] vdd gnd cell_6t
Xbit_r191_c79 bl[79] br[79] wl[191] vdd gnd cell_6t
Xbit_r192_c79 bl[79] br[79] wl[192] vdd gnd cell_6t
Xbit_r193_c79 bl[79] br[79] wl[193] vdd gnd cell_6t
Xbit_r194_c79 bl[79] br[79] wl[194] vdd gnd cell_6t
Xbit_r195_c79 bl[79] br[79] wl[195] vdd gnd cell_6t
Xbit_r196_c79 bl[79] br[79] wl[196] vdd gnd cell_6t
Xbit_r197_c79 bl[79] br[79] wl[197] vdd gnd cell_6t
Xbit_r198_c79 bl[79] br[79] wl[198] vdd gnd cell_6t
Xbit_r199_c79 bl[79] br[79] wl[199] vdd gnd cell_6t
Xbit_r200_c79 bl[79] br[79] wl[200] vdd gnd cell_6t
Xbit_r201_c79 bl[79] br[79] wl[201] vdd gnd cell_6t
Xbit_r202_c79 bl[79] br[79] wl[202] vdd gnd cell_6t
Xbit_r203_c79 bl[79] br[79] wl[203] vdd gnd cell_6t
Xbit_r204_c79 bl[79] br[79] wl[204] vdd gnd cell_6t
Xbit_r205_c79 bl[79] br[79] wl[205] vdd gnd cell_6t
Xbit_r206_c79 bl[79] br[79] wl[206] vdd gnd cell_6t
Xbit_r207_c79 bl[79] br[79] wl[207] vdd gnd cell_6t
Xbit_r208_c79 bl[79] br[79] wl[208] vdd gnd cell_6t
Xbit_r209_c79 bl[79] br[79] wl[209] vdd gnd cell_6t
Xbit_r210_c79 bl[79] br[79] wl[210] vdd gnd cell_6t
Xbit_r211_c79 bl[79] br[79] wl[211] vdd gnd cell_6t
Xbit_r212_c79 bl[79] br[79] wl[212] vdd gnd cell_6t
Xbit_r213_c79 bl[79] br[79] wl[213] vdd gnd cell_6t
Xbit_r214_c79 bl[79] br[79] wl[214] vdd gnd cell_6t
Xbit_r215_c79 bl[79] br[79] wl[215] vdd gnd cell_6t
Xbit_r216_c79 bl[79] br[79] wl[216] vdd gnd cell_6t
Xbit_r217_c79 bl[79] br[79] wl[217] vdd gnd cell_6t
Xbit_r218_c79 bl[79] br[79] wl[218] vdd gnd cell_6t
Xbit_r219_c79 bl[79] br[79] wl[219] vdd gnd cell_6t
Xbit_r220_c79 bl[79] br[79] wl[220] vdd gnd cell_6t
Xbit_r221_c79 bl[79] br[79] wl[221] vdd gnd cell_6t
Xbit_r222_c79 bl[79] br[79] wl[222] vdd gnd cell_6t
Xbit_r223_c79 bl[79] br[79] wl[223] vdd gnd cell_6t
Xbit_r224_c79 bl[79] br[79] wl[224] vdd gnd cell_6t
Xbit_r225_c79 bl[79] br[79] wl[225] vdd gnd cell_6t
Xbit_r226_c79 bl[79] br[79] wl[226] vdd gnd cell_6t
Xbit_r227_c79 bl[79] br[79] wl[227] vdd gnd cell_6t
Xbit_r228_c79 bl[79] br[79] wl[228] vdd gnd cell_6t
Xbit_r229_c79 bl[79] br[79] wl[229] vdd gnd cell_6t
Xbit_r230_c79 bl[79] br[79] wl[230] vdd gnd cell_6t
Xbit_r231_c79 bl[79] br[79] wl[231] vdd gnd cell_6t
Xbit_r232_c79 bl[79] br[79] wl[232] vdd gnd cell_6t
Xbit_r233_c79 bl[79] br[79] wl[233] vdd gnd cell_6t
Xbit_r234_c79 bl[79] br[79] wl[234] vdd gnd cell_6t
Xbit_r235_c79 bl[79] br[79] wl[235] vdd gnd cell_6t
Xbit_r236_c79 bl[79] br[79] wl[236] vdd gnd cell_6t
Xbit_r237_c79 bl[79] br[79] wl[237] vdd gnd cell_6t
Xbit_r238_c79 bl[79] br[79] wl[238] vdd gnd cell_6t
Xbit_r239_c79 bl[79] br[79] wl[239] vdd gnd cell_6t
Xbit_r240_c79 bl[79] br[79] wl[240] vdd gnd cell_6t
Xbit_r241_c79 bl[79] br[79] wl[241] vdd gnd cell_6t
Xbit_r242_c79 bl[79] br[79] wl[242] vdd gnd cell_6t
Xbit_r243_c79 bl[79] br[79] wl[243] vdd gnd cell_6t
Xbit_r244_c79 bl[79] br[79] wl[244] vdd gnd cell_6t
Xbit_r245_c79 bl[79] br[79] wl[245] vdd gnd cell_6t
Xbit_r246_c79 bl[79] br[79] wl[246] vdd gnd cell_6t
Xbit_r247_c79 bl[79] br[79] wl[247] vdd gnd cell_6t
Xbit_r248_c79 bl[79] br[79] wl[248] vdd gnd cell_6t
Xbit_r249_c79 bl[79] br[79] wl[249] vdd gnd cell_6t
Xbit_r250_c79 bl[79] br[79] wl[250] vdd gnd cell_6t
Xbit_r251_c79 bl[79] br[79] wl[251] vdd gnd cell_6t
Xbit_r252_c79 bl[79] br[79] wl[252] vdd gnd cell_6t
Xbit_r253_c79 bl[79] br[79] wl[253] vdd gnd cell_6t
Xbit_r254_c79 bl[79] br[79] wl[254] vdd gnd cell_6t
Xbit_r255_c79 bl[79] br[79] wl[255] vdd gnd cell_6t
Xbit_r256_c79 bl[79] br[79] wl[256] vdd gnd cell_6t
Xbit_r257_c79 bl[79] br[79] wl[257] vdd gnd cell_6t
Xbit_r258_c79 bl[79] br[79] wl[258] vdd gnd cell_6t
Xbit_r259_c79 bl[79] br[79] wl[259] vdd gnd cell_6t
Xbit_r260_c79 bl[79] br[79] wl[260] vdd gnd cell_6t
Xbit_r261_c79 bl[79] br[79] wl[261] vdd gnd cell_6t
Xbit_r262_c79 bl[79] br[79] wl[262] vdd gnd cell_6t
Xbit_r263_c79 bl[79] br[79] wl[263] vdd gnd cell_6t
Xbit_r264_c79 bl[79] br[79] wl[264] vdd gnd cell_6t
Xbit_r265_c79 bl[79] br[79] wl[265] vdd gnd cell_6t
Xbit_r266_c79 bl[79] br[79] wl[266] vdd gnd cell_6t
Xbit_r267_c79 bl[79] br[79] wl[267] vdd gnd cell_6t
Xbit_r268_c79 bl[79] br[79] wl[268] vdd gnd cell_6t
Xbit_r269_c79 bl[79] br[79] wl[269] vdd gnd cell_6t
Xbit_r270_c79 bl[79] br[79] wl[270] vdd gnd cell_6t
Xbit_r271_c79 bl[79] br[79] wl[271] vdd gnd cell_6t
Xbit_r272_c79 bl[79] br[79] wl[272] vdd gnd cell_6t
Xbit_r273_c79 bl[79] br[79] wl[273] vdd gnd cell_6t
Xbit_r274_c79 bl[79] br[79] wl[274] vdd gnd cell_6t
Xbit_r275_c79 bl[79] br[79] wl[275] vdd gnd cell_6t
Xbit_r276_c79 bl[79] br[79] wl[276] vdd gnd cell_6t
Xbit_r277_c79 bl[79] br[79] wl[277] vdd gnd cell_6t
Xbit_r278_c79 bl[79] br[79] wl[278] vdd gnd cell_6t
Xbit_r279_c79 bl[79] br[79] wl[279] vdd gnd cell_6t
Xbit_r280_c79 bl[79] br[79] wl[280] vdd gnd cell_6t
Xbit_r281_c79 bl[79] br[79] wl[281] vdd gnd cell_6t
Xbit_r282_c79 bl[79] br[79] wl[282] vdd gnd cell_6t
Xbit_r283_c79 bl[79] br[79] wl[283] vdd gnd cell_6t
Xbit_r284_c79 bl[79] br[79] wl[284] vdd gnd cell_6t
Xbit_r285_c79 bl[79] br[79] wl[285] vdd gnd cell_6t
Xbit_r286_c79 bl[79] br[79] wl[286] vdd gnd cell_6t
Xbit_r287_c79 bl[79] br[79] wl[287] vdd gnd cell_6t
Xbit_r288_c79 bl[79] br[79] wl[288] vdd gnd cell_6t
Xbit_r289_c79 bl[79] br[79] wl[289] vdd gnd cell_6t
Xbit_r290_c79 bl[79] br[79] wl[290] vdd gnd cell_6t
Xbit_r291_c79 bl[79] br[79] wl[291] vdd gnd cell_6t
Xbit_r292_c79 bl[79] br[79] wl[292] vdd gnd cell_6t
Xbit_r293_c79 bl[79] br[79] wl[293] vdd gnd cell_6t
Xbit_r294_c79 bl[79] br[79] wl[294] vdd gnd cell_6t
Xbit_r295_c79 bl[79] br[79] wl[295] vdd gnd cell_6t
Xbit_r296_c79 bl[79] br[79] wl[296] vdd gnd cell_6t
Xbit_r297_c79 bl[79] br[79] wl[297] vdd gnd cell_6t
Xbit_r298_c79 bl[79] br[79] wl[298] vdd gnd cell_6t
Xbit_r299_c79 bl[79] br[79] wl[299] vdd gnd cell_6t
Xbit_r300_c79 bl[79] br[79] wl[300] vdd gnd cell_6t
Xbit_r301_c79 bl[79] br[79] wl[301] vdd gnd cell_6t
Xbit_r302_c79 bl[79] br[79] wl[302] vdd gnd cell_6t
Xbit_r303_c79 bl[79] br[79] wl[303] vdd gnd cell_6t
Xbit_r304_c79 bl[79] br[79] wl[304] vdd gnd cell_6t
Xbit_r305_c79 bl[79] br[79] wl[305] vdd gnd cell_6t
Xbit_r306_c79 bl[79] br[79] wl[306] vdd gnd cell_6t
Xbit_r307_c79 bl[79] br[79] wl[307] vdd gnd cell_6t
Xbit_r308_c79 bl[79] br[79] wl[308] vdd gnd cell_6t
Xbit_r309_c79 bl[79] br[79] wl[309] vdd gnd cell_6t
Xbit_r310_c79 bl[79] br[79] wl[310] vdd gnd cell_6t
Xbit_r311_c79 bl[79] br[79] wl[311] vdd gnd cell_6t
Xbit_r312_c79 bl[79] br[79] wl[312] vdd gnd cell_6t
Xbit_r313_c79 bl[79] br[79] wl[313] vdd gnd cell_6t
Xbit_r314_c79 bl[79] br[79] wl[314] vdd gnd cell_6t
Xbit_r315_c79 bl[79] br[79] wl[315] vdd gnd cell_6t
Xbit_r316_c79 bl[79] br[79] wl[316] vdd gnd cell_6t
Xbit_r317_c79 bl[79] br[79] wl[317] vdd gnd cell_6t
Xbit_r318_c79 bl[79] br[79] wl[318] vdd gnd cell_6t
Xbit_r319_c79 bl[79] br[79] wl[319] vdd gnd cell_6t
Xbit_r320_c79 bl[79] br[79] wl[320] vdd gnd cell_6t
Xbit_r321_c79 bl[79] br[79] wl[321] vdd gnd cell_6t
Xbit_r322_c79 bl[79] br[79] wl[322] vdd gnd cell_6t
Xbit_r323_c79 bl[79] br[79] wl[323] vdd gnd cell_6t
Xbit_r324_c79 bl[79] br[79] wl[324] vdd gnd cell_6t
Xbit_r325_c79 bl[79] br[79] wl[325] vdd gnd cell_6t
Xbit_r326_c79 bl[79] br[79] wl[326] vdd gnd cell_6t
Xbit_r327_c79 bl[79] br[79] wl[327] vdd gnd cell_6t
Xbit_r328_c79 bl[79] br[79] wl[328] vdd gnd cell_6t
Xbit_r329_c79 bl[79] br[79] wl[329] vdd gnd cell_6t
Xbit_r330_c79 bl[79] br[79] wl[330] vdd gnd cell_6t
Xbit_r331_c79 bl[79] br[79] wl[331] vdd gnd cell_6t
Xbit_r332_c79 bl[79] br[79] wl[332] vdd gnd cell_6t
Xbit_r333_c79 bl[79] br[79] wl[333] vdd gnd cell_6t
Xbit_r334_c79 bl[79] br[79] wl[334] vdd gnd cell_6t
Xbit_r335_c79 bl[79] br[79] wl[335] vdd gnd cell_6t
Xbit_r336_c79 bl[79] br[79] wl[336] vdd gnd cell_6t
Xbit_r337_c79 bl[79] br[79] wl[337] vdd gnd cell_6t
Xbit_r338_c79 bl[79] br[79] wl[338] vdd gnd cell_6t
Xbit_r339_c79 bl[79] br[79] wl[339] vdd gnd cell_6t
Xbit_r340_c79 bl[79] br[79] wl[340] vdd gnd cell_6t
Xbit_r341_c79 bl[79] br[79] wl[341] vdd gnd cell_6t
Xbit_r342_c79 bl[79] br[79] wl[342] vdd gnd cell_6t
Xbit_r343_c79 bl[79] br[79] wl[343] vdd gnd cell_6t
Xbit_r344_c79 bl[79] br[79] wl[344] vdd gnd cell_6t
Xbit_r345_c79 bl[79] br[79] wl[345] vdd gnd cell_6t
Xbit_r346_c79 bl[79] br[79] wl[346] vdd gnd cell_6t
Xbit_r347_c79 bl[79] br[79] wl[347] vdd gnd cell_6t
Xbit_r348_c79 bl[79] br[79] wl[348] vdd gnd cell_6t
Xbit_r349_c79 bl[79] br[79] wl[349] vdd gnd cell_6t
Xbit_r350_c79 bl[79] br[79] wl[350] vdd gnd cell_6t
Xbit_r351_c79 bl[79] br[79] wl[351] vdd gnd cell_6t
Xbit_r352_c79 bl[79] br[79] wl[352] vdd gnd cell_6t
Xbit_r353_c79 bl[79] br[79] wl[353] vdd gnd cell_6t
Xbit_r354_c79 bl[79] br[79] wl[354] vdd gnd cell_6t
Xbit_r355_c79 bl[79] br[79] wl[355] vdd gnd cell_6t
Xbit_r356_c79 bl[79] br[79] wl[356] vdd gnd cell_6t
Xbit_r357_c79 bl[79] br[79] wl[357] vdd gnd cell_6t
Xbit_r358_c79 bl[79] br[79] wl[358] vdd gnd cell_6t
Xbit_r359_c79 bl[79] br[79] wl[359] vdd gnd cell_6t
Xbit_r360_c79 bl[79] br[79] wl[360] vdd gnd cell_6t
Xbit_r361_c79 bl[79] br[79] wl[361] vdd gnd cell_6t
Xbit_r362_c79 bl[79] br[79] wl[362] vdd gnd cell_6t
Xbit_r363_c79 bl[79] br[79] wl[363] vdd gnd cell_6t
Xbit_r364_c79 bl[79] br[79] wl[364] vdd gnd cell_6t
Xbit_r365_c79 bl[79] br[79] wl[365] vdd gnd cell_6t
Xbit_r366_c79 bl[79] br[79] wl[366] vdd gnd cell_6t
Xbit_r367_c79 bl[79] br[79] wl[367] vdd gnd cell_6t
Xbit_r368_c79 bl[79] br[79] wl[368] vdd gnd cell_6t
Xbit_r369_c79 bl[79] br[79] wl[369] vdd gnd cell_6t
Xbit_r370_c79 bl[79] br[79] wl[370] vdd gnd cell_6t
Xbit_r371_c79 bl[79] br[79] wl[371] vdd gnd cell_6t
Xbit_r372_c79 bl[79] br[79] wl[372] vdd gnd cell_6t
Xbit_r373_c79 bl[79] br[79] wl[373] vdd gnd cell_6t
Xbit_r374_c79 bl[79] br[79] wl[374] vdd gnd cell_6t
Xbit_r375_c79 bl[79] br[79] wl[375] vdd gnd cell_6t
Xbit_r376_c79 bl[79] br[79] wl[376] vdd gnd cell_6t
Xbit_r377_c79 bl[79] br[79] wl[377] vdd gnd cell_6t
Xbit_r378_c79 bl[79] br[79] wl[378] vdd gnd cell_6t
Xbit_r379_c79 bl[79] br[79] wl[379] vdd gnd cell_6t
Xbit_r380_c79 bl[79] br[79] wl[380] vdd gnd cell_6t
Xbit_r381_c79 bl[79] br[79] wl[381] vdd gnd cell_6t
Xbit_r382_c79 bl[79] br[79] wl[382] vdd gnd cell_6t
Xbit_r383_c79 bl[79] br[79] wl[383] vdd gnd cell_6t
Xbit_r384_c79 bl[79] br[79] wl[384] vdd gnd cell_6t
Xbit_r385_c79 bl[79] br[79] wl[385] vdd gnd cell_6t
Xbit_r386_c79 bl[79] br[79] wl[386] vdd gnd cell_6t
Xbit_r387_c79 bl[79] br[79] wl[387] vdd gnd cell_6t
Xbit_r388_c79 bl[79] br[79] wl[388] vdd gnd cell_6t
Xbit_r389_c79 bl[79] br[79] wl[389] vdd gnd cell_6t
Xbit_r390_c79 bl[79] br[79] wl[390] vdd gnd cell_6t
Xbit_r391_c79 bl[79] br[79] wl[391] vdd gnd cell_6t
Xbit_r392_c79 bl[79] br[79] wl[392] vdd gnd cell_6t
Xbit_r393_c79 bl[79] br[79] wl[393] vdd gnd cell_6t
Xbit_r394_c79 bl[79] br[79] wl[394] vdd gnd cell_6t
Xbit_r395_c79 bl[79] br[79] wl[395] vdd gnd cell_6t
Xbit_r396_c79 bl[79] br[79] wl[396] vdd gnd cell_6t
Xbit_r397_c79 bl[79] br[79] wl[397] vdd gnd cell_6t
Xbit_r398_c79 bl[79] br[79] wl[398] vdd gnd cell_6t
Xbit_r399_c79 bl[79] br[79] wl[399] vdd gnd cell_6t
Xbit_r400_c79 bl[79] br[79] wl[400] vdd gnd cell_6t
Xbit_r401_c79 bl[79] br[79] wl[401] vdd gnd cell_6t
Xbit_r402_c79 bl[79] br[79] wl[402] vdd gnd cell_6t
Xbit_r403_c79 bl[79] br[79] wl[403] vdd gnd cell_6t
Xbit_r404_c79 bl[79] br[79] wl[404] vdd gnd cell_6t
Xbit_r405_c79 bl[79] br[79] wl[405] vdd gnd cell_6t
Xbit_r406_c79 bl[79] br[79] wl[406] vdd gnd cell_6t
Xbit_r407_c79 bl[79] br[79] wl[407] vdd gnd cell_6t
Xbit_r408_c79 bl[79] br[79] wl[408] vdd gnd cell_6t
Xbit_r409_c79 bl[79] br[79] wl[409] vdd gnd cell_6t
Xbit_r410_c79 bl[79] br[79] wl[410] vdd gnd cell_6t
Xbit_r411_c79 bl[79] br[79] wl[411] vdd gnd cell_6t
Xbit_r412_c79 bl[79] br[79] wl[412] vdd gnd cell_6t
Xbit_r413_c79 bl[79] br[79] wl[413] vdd gnd cell_6t
Xbit_r414_c79 bl[79] br[79] wl[414] vdd gnd cell_6t
Xbit_r415_c79 bl[79] br[79] wl[415] vdd gnd cell_6t
Xbit_r416_c79 bl[79] br[79] wl[416] vdd gnd cell_6t
Xbit_r417_c79 bl[79] br[79] wl[417] vdd gnd cell_6t
Xbit_r418_c79 bl[79] br[79] wl[418] vdd gnd cell_6t
Xbit_r419_c79 bl[79] br[79] wl[419] vdd gnd cell_6t
Xbit_r420_c79 bl[79] br[79] wl[420] vdd gnd cell_6t
Xbit_r421_c79 bl[79] br[79] wl[421] vdd gnd cell_6t
Xbit_r422_c79 bl[79] br[79] wl[422] vdd gnd cell_6t
Xbit_r423_c79 bl[79] br[79] wl[423] vdd gnd cell_6t
Xbit_r424_c79 bl[79] br[79] wl[424] vdd gnd cell_6t
Xbit_r425_c79 bl[79] br[79] wl[425] vdd gnd cell_6t
Xbit_r426_c79 bl[79] br[79] wl[426] vdd gnd cell_6t
Xbit_r427_c79 bl[79] br[79] wl[427] vdd gnd cell_6t
Xbit_r428_c79 bl[79] br[79] wl[428] vdd gnd cell_6t
Xbit_r429_c79 bl[79] br[79] wl[429] vdd gnd cell_6t
Xbit_r430_c79 bl[79] br[79] wl[430] vdd gnd cell_6t
Xbit_r431_c79 bl[79] br[79] wl[431] vdd gnd cell_6t
Xbit_r432_c79 bl[79] br[79] wl[432] vdd gnd cell_6t
Xbit_r433_c79 bl[79] br[79] wl[433] vdd gnd cell_6t
Xbit_r434_c79 bl[79] br[79] wl[434] vdd gnd cell_6t
Xbit_r435_c79 bl[79] br[79] wl[435] vdd gnd cell_6t
Xbit_r436_c79 bl[79] br[79] wl[436] vdd gnd cell_6t
Xbit_r437_c79 bl[79] br[79] wl[437] vdd gnd cell_6t
Xbit_r438_c79 bl[79] br[79] wl[438] vdd gnd cell_6t
Xbit_r439_c79 bl[79] br[79] wl[439] vdd gnd cell_6t
Xbit_r440_c79 bl[79] br[79] wl[440] vdd gnd cell_6t
Xbit_r441_c79 bl[79] br[79] wl[441] vdd gnd cell_6t
Xbit_r442_c79 bl[79] br[79] wl[442] vdd gnd cell_6t
Xbit_r443_c79 bl[79] br[79] wl[443] vdd gnd cell_6t
Xbit_r444_c79 bl[79] br[79] wl[444] vdd gnd cell_6t
Xbit_r445_c79 bl[79] br[79] wl[445] vdd gnd cell_6t
Xbit_r446_c79 bl[79] br[79] wl[446] vdd gnd cell_6t
Xbit_r447_c79 bl[79] br[79] wl[447] vdd gnd cell_6t
Xbit_r448_c79 bl[79] br[79] wl[448] vdd gnd cell_6t
Xbit_r449_c79 bl[79] br[79] wl[449] vdd gnd cell_6t
Xbit_r450_c79 bl[79] br[79] wl[450] vdd gnd cell_6t
Xbit_r451_c79 bl[79] br[79] wl[451] vdd gnd cell_6t
Xbit_r452_c79 bl[79] br[79] wl[452] vdd gnd cell_6t
Xbit_r453_c79 bl[79] br[79] wl[453] vdd gnd cell_6t
Xbit_r454_c79 bl[79] br[79] wl[454] vdd gnd cell_6t
Xbit_r455_c79 bl[79] br[79] wl[455] vdd gnd cell_6t
Xbit_r456_c79 bl[79] br[79] wl[456] vdd gnd cell_6t
Xbit_r457_c79 bl[79] br[79] wl[457] vdd gnd cell_6t
Xbit_r458_c79 bl[79] br[79] wl[458] vdd gnd cell_6t
Xbit_r459_c79 bl[79] br[79] wl[459] vdd gnd cell_6t
Xbit_r460_c79 bl[79] br[79] wl[460] vdd gnd cell_6t
Xbit_r461_c79 bl[79] br[79] wl[461] vdd gnd cell_6t
Xbit_r462_c79 bl[79] br[79] wl[462] vdd gnd cell_6t
Xbit_r463_c79 bl[79] br[79] wl[463] vdd gnd cell_6t
Xbit_r464_c79 bl[79] br[79] wl[464] vdd gnd cell_6t
Xbit_r465_c79 bl[79] br[79] wl[465] vdd gnd cell_6t
Xbit_r466_c79 bl[79] br[79] wl[466] vdd gnd cell_6t
Xbit_r467_c79 bl[79] br[79] wl[467] vdd gnd cell_6t
Xbit_r468_c79 bl[79] br[79] wl[468] vdd gnd cell_6t
Xbit_r469_c79 bl[79] br[79] wl[469] vdd gnd cell_6t
Xbit_r470_c79 bl[79] br[79] wl[470] vdd gnd cell_6t
Xbit_r471_c79 bl[79] br[79] wl[471] vdd gnd cell_6t
Xbit_r472_c79 bl[79] br[79] wl[472] vdd gnd cell_6t
Xbit_r473_c79 bl[79] br[79] wl[473] vdd gnd cell_6t
Xbit_r474_c79 bl[79] br[79] wl[474] vdd gnd cell_6t
Xbit_r475_c79 bl[79] br[79] wl[475] vdd gnd cell_6t
Xbit_r476_c79 bl[79] br[79] wl[476] vdd gnd cell_6t
Xbit_r477_c79 bl[79] br[79] wl[477] vdd gnd cell_6t
Xbit_r478_c79 bl[79] br[79] wl[478] vdd gnd cell_6t
Xbit_r479_c79 bl[79] br[79] wl[479] vdd gnd cell_6t
Xbit_r480_c79 bl[79] br[79] wl[480] vdd gnd cell_6t
Xbit_r481_c79 bl[79] br[79] wl[481] vdd gnd cell_6t
Xbit_r482_c79 bl[79] br[79] wl[482] vdd gnd cell_6t
Xbit_r483_c79 bl[79] br[79] wl[483] vdd gnd cell_6t
Xbit_r484_c79 bl[79] br[79] wl[484] vdd gnd cell_6t
Xbit_r485_c79 bl[79] br[79] wl[485] vdd gnd cell_6t
Xbit_r486_c79 bl[79] br[79] wl[486] vdd gnd cell_6t
Xbit_r487_c79 bl[79] br[79] wl[487] vdd gnd cell_6t
Xbit_r488_c79 bl[79] br[79] wl[488] vdd gnd cell_6t
Xbit_r489_c79 bl[79] br[79] wl[489] vdd gnd cell_6t
Xbit_r490_c79 bl[79] br[79] wl[490] vdd gnd cell_6t
Xbit_r491_c79 bl[79] br[79] wl[491] vdd gnd cell_6t
Xbit_r492_c79 bl[79] br[79] wl[492] vdd gnd cell_6t
Xbit_r493_c79 bl[79] br[79] wl[493] vdd gnd cell_6t
Xbit_r494_c79 bl[79] br[79] wl[494] vdd gnd cell_6t
Xbit_r495_c79 bl[79] br[79] wl[495] vdd gnd cell_6t
Xbit_r496_c79 bl[79] br[79] wl[496] vdd gnd cell_6t
Xbit_r497_c79 bl[79] br[79] wl[497] vdd gnd cell_6t
Xbit_r498_c79 bl[79] br[79] wl[498] vdd gnd cell_6t
Xbit_r499_c79 bl[79] br[79] wl[499] vdd gnd cell_6t
Xbit_r500_c79 bl[79] br[79] wl[500] vdd gnd cell_6t
Xbit_r501_c79 bl[79] br[79] wl[501] vdd gnd cell_6t
Xbit_r502_c79 bl[79] br[79] wl[502] vdd gnd cell_6t
Xbit_r503_c79 bl[79] br[79] wl[503] vdd gnd cell_6t
Xbit_r504_c79 bl[79] br[79] wl[504] vdd gnd cell_6t
Xbit_r505_c79 bl[79] br[79] wl[505] vdd gnd cell_6t
Xbit_r506_c79 bl[79] br[79] wl[506] vdd gnd cell_6t
Xbit_r507_c79 bl[79] br[79] wl[507] vdd gnd cell_6t
Xbit_r508_c79 bl[79] br[79] wl[508] vdd gnd cell_6t
Xbit_r509_c79 bl[79] br[79] wl[509] vdd gnd cell_6t
Xbit_r510_c79 bl[79] br[79] wl[510] vdd gnd cell_6t
Xbit_r511_c79 bl[79] br[79] wl[511] vdd gnd cell_6t
Xbit_r0_c80 bl[80] br[80] wl[0] vdd gnd cell_6t
Xbit_r1_c80 bl[80] br[80] wl[1] vdd gnd cell_6t
Xbit_r2_c80 bl[80] br[80] wl[2] vdd gnd cell_6t
Xbit_r3_c80 bl[80] br[80] wl[3] vdd gnd cell_6t
Xbit_r4_c80 bl[80] br[80] wl[4] vdd gnd cell_6t
Xbit_r5_c80 bl[80] br[80] wl[5] vdd gnd cell_6t
Xbit_r6_c80 bl[80] br[80] wl[6] vdd gnd cell_6t
Xbit_r7_c80 bl[80] br[80] wl[7] vdd gnd cell_6t
Xbit_r8_c80 bl[80] br[80] wl[8] vdd gnd cell_6t
Xbit_r9_c80 bl[80] br[80] wl[9] vdd gnd cell_6t
Xbit_r10_c80 bl[80] br[80] wl[10] vdd gnd cell_6t
Xbit_r11_c80 bl[80] br[80] wl[11] vdd gnd cell_6t
Xbit_r12_c80 bl[80] br[80] wl[12] vdd gnd cell_6t
Xbit_r13_c80 bl[80] br[80] wl[13] vdd gnd cell_6t
Xbit_r14_c80 bl[80] br[80] wl[14] vdd gnd cell_6t
Xbit_r15_c80 bl[80] br[80] wl[15] vdd gnd cell_6t
Xbit_r16_c80 bl[80] br[80] wl[16] vdd gnd cell_6t
Xbit_r17_c80 bl[80] br[80] wl[17] vdd gnd cell_6t
Xbit_r18_c80 bl[80] br[80] wl[18] vdd gnd cell_6t
Xbit_r19_c80 bl[80] br[80] wl[19] vdd gnd cell_6t
Xbit_r20_c80 bl[80] br[80] wl[20] vdd gnd cell_6t
Xbit_r21_c80 bl[80] br[80] wl[21] vdd gnd cell_6t
Xbit_r22_c80 bl[80] br[80] wl[22] vdd gnd cell_6t
Xbit_r23_c80 bl[80] br[80] wl[23] vdd gnd cell_6t
Xbit_r24_c80 bl[80] br[80] wl[24] vdd gnd cell_6t
Xbit_r25_c80 bl[80] br[80] wl[25] vdd gnd cell_6t
Xbit_r26_c80 bl[80] br[80] wl[26] vdd gnd cell_6t
Xbit_r27_c80 bl[80] br[80] wl[27] vdd gnd cell_6t
Xbit_r28_c80 bl[80] br[80] wl[28] vdd gnd cell_6t
Xbit_r29_c80 bl[80] br[80] wl[29] vdd gnd cell_6t
Xbit_r30_c80 bl[80] br[80] wl[30] vdd gnd cell_6t
Xbit_r31_c80 bl[80] br[80] wl[31] vdd gnd cell_6t
Xbit_r32_c80 bl[80] br[80] wl[32] vdd gnd cell_6t
Xbit_r33_c80 bl[80] br[80] wl[33] vdd gnd cell_6t
Xbit_r34_c80 bl[80] br[80] wl[34] vdd gnd cell_6t
Xbit_r35_c80 bl[80] br[80] wl[35] vdd gnd cell_6t
Xbit_r36_c80 bl[80] br[80] wl[36] vdd gnd cell_6t
Xbit_r37_c80 bl[80] br[80] wl[37] vdd gnd cell_6t
Xbit_r38_c80 bl[80] br[80] wl[38] vdd gnd cell_6t
Xbit_r39_c80 bl[80] br[80] wl[39] vdd gnd cell_6t
Xbit_r40_c80 bl[80] br[80] wl[40] vdd gnd cell_6t
Xbit_r41_c80 bl[80] br[80] wl[41] vdd gnd cell_6t
Xbit_r42_c80 bl[80] br[80] wl[42] vdd gnd cell_6t
Xbit_r43_c80 bl[80] br[80] wl[43] vdd gnd cell_6t
Xbit_r44_c80 bl[80] br[80] wl[44] vdd gnd cell_6t
Xbit_r45_c80 bl[80] br[80] wl[45] vdd gnd cell_6t
Xbit_r46_c80 bl[80] br[80] wl[46] vdd gnd cell_6t
Xbit_r47_c80 bl[80] br[80] wl[47] vdd gnd cell_6t
Xbit_r48_c80 bl[80] br[80] wl[48] vdd gnd cell_6t
Xbit_r49_c80 bl[80] br[80] wl[49] vdd gnd cell_6t
Xbit_r50_c80 bl[80] br[80] wl[50] vdd gnd cell_6t
Xbit_r51_c80 bl[80] br[80] wl[51] vdd gnd cell_6t
Xbit_r52_c80 bl[80] br[80] wl[52] vdd gnd cell_6t
Xbit_r53_c80 bl[80] br[80] wl[53] vdd gnd cell_6t
Xbit_r54_c80 bl[80] br[80] wl[54] vdd gnd cell_6t
Xbit_r55_c80 bl[80] br[80] wl[55] vdd gnd cell_6t
Xbit_r56_c80 bl[80] br[80] wl[56] vdd gnd cell_6t
Xbit_r57_c80 bl[80] br[80] wl[57] vdd gnd cell_6t
Xbit_r58_c80 bl[80] br[80] wl[58] vdd gnd cell_6t
Xbit_r59_c80 bl[80] br[80] wl[59] vdd gnd cell_6t
Xbit_r60_c80 bl[80] br[80] wl[60] vdd gnd cell_6t
Xbit_r61_c80 bl[80] br[80] wl[61] vdd gnd cell_6t
Xbit_r62_c80 bl[80] br[80] wl[62] vdd gnd cell_6t
Xbit_r63_c80 bl[80] br[80] wl[63] vdd gnd cell_6t
Xbit_r64_c80 bl[80] br[80] wl[64] vdd gnd cell_6t
Xbit_r65_c80 bl[80] br[80] wl[65] vdd gnd cell_6t
Xbit_r66_c80 bl[80] br[80] wl[66] vdd gnd cell_6t
Xbit_r67_c80 bl[80] br[80] wl[67] vdd gnd cell_6t
Xbit_r68_c80 bl[80] br[80] wl[68] vdd gnd cell_6t
Xbit_r69_c80 bl[80] br[80] wl[69] vdd gnd cell_6t
Xbit_r70_c80 bl[80] br[80] wl[70] vdd gnd cell_6t
Xbit_r71_c80 bl[80] br[80] wl[71] vdd gnd cell_6t
Xbit_r72_c80 bl[80] br[80] wl[72] vdd gnd cell_6t
Xbit_r73_c80 bl[80] br[80] wl[73] vdd gnd cell_6t
Xbit_r74_c80 bl[80] br[80] wl[74] vdd gnd cell_6t
Xbit_r75_c80 bl[80] br[80] wl[75] vdd gnd cell_6t
Xbit_r76_c80 bl[80] br[80] wl[76] vdd gnd cell_6t
Xbit_r77_c80 bl[80] br[80] wl[77] vdd gnd cell_6t
Xbit_r78_c80 bl[80] br[80] wl[78] vdd gnd cell_6t
Xbit_r79_c80 bl[80] br[80] wl[79] vdd gnd cell_6t
Xbit_r80_c80 bl[80] br[80] wl[80] vdd gnd cell_6t
Xbit_r81_c80 bl[80] br[80] wl[81] vdd gnd cell_6t
Xbit_r82_c80 bl[80] br[80] wl[82] vdd gnd cell_6t
Xbit_r83_c80 bl[80] br[80] wl[83] vdd gnd cell_6t
Xbit_r84_c80 bl[80] br[80] wl[84] vdd gnd cell_6t
Xbit_r85_c80 bl[80] br[80] wl[85] vdd gnd cell_6t
Xbit_r86_c80 bl[80] br[80] wl[86] vdd gnd cell_6t
Xbit_r87_c80 bl[80] br[80] wl[87] vdd gnd cell_6t
Xbit_r88_c80 bl[80] br[80] wl[88] vdd gnd cell_6t
Xbit_r89_c80 bl[80] br[80] wl[89] vdd gnd cell_6t
Xbit_r90_c80 bl[80] br[80] wl[90] vdd gnd cell_6t
Xbit_r91_c80 bl[80] br[80] wl[91] vdd gnd cell_6t
Xbit_r92_c80 bl[80] br[80] wl[92] vdd gnd cell_6t
Xbit_r93_c80 bl[80] br[80] wl[93] vdd gnd cell_6t
Xbit_r94_c80 bl[80] br[80] wl[94] vdd gnd cell_6t
Xbit_r95_c80 bl[80] br[80] wl[95] vdd gnd cell_6t
Xbit_r96_c80 bl[80] br[80] wl[96] vdd gnd cell_6t
Xbit_r97_c80 bl[80] br[80] wl[97] vdd gnd cell_6t
Xbit_r98_c80 bl[80] br[80] wl[98] vdd gnd cell_6t
Xbit_r99_c80 bl[80] br[80] wl[99] vdd gnd cell_6t
Xbit_r100_c80 bl[80] br[80] wl[100] vdd gnd cell_6t
Xbit_r101_c80 bl[80] br[80] wl[101] vdd gnd cell_6t
Xbit_r102_c80 bl[80] br[80] wl[102] vdd gnd cell_6t
Xbit_r103_c80 bl[80] br[80] wl[103] vdd gnd cell_6t
Xbit_r104_c80 bl[80] br[80] wl[104] vdd gnd cell_6t
Xbit_r105_c80 bl[80] br[80] wl[105] vdd gnd cell_6t
Xbit_r106_c80 bl[80] br[80] wl[106] vdd gnd cell_6t
Xbit_r107_c80 bl[80] br[80] wl[107] vdd gnd cell_6t
Xbit_r108_c80 bl[80] br[80] wl[108] vdd gnd cell_6t
Xbit_r109_c80 bl[80] br[80] wl[109] vdd gnd cell_6t
Xbit_r110_c80 bl[80] br[80] wl[110] vdd gnd cell_6t
Xbit_r111_c80 bl[80] br[80] wl[111] vdd gnd cell_6t
Xbit_r112_c80 bl[80] br[80] wl[112] vdd gnd cell_6t
Xbit_r113_c80 bl[80] br[80] wl[113] vdd gnd cell_6t
Xbit_r114_c80 bl[80] br[80] wl[114] vdd gnd cell_6t
Xbit_r115_c80 bl[80] br[80] wl[115] vdd gnd cell_6t
Xbit_r116_c80 bl[80] br[80] wl[116] vdd gnd cell_6t
Xbit_r117_c80 bl[80] br[80] wl[117] vdd gnd cell_6t
Xbit_r118_c80 bl[80] br[80] wl[118] vdd gnd cell_6t
Xbit_r119_c80 bl[80] br[80] wl[119] vdd gnd cell_6t
Xbit_r120_c80 bl[80] br[80] wl[120] vdd gnd cell_6t
Xbit_r121_c80 bl[80] br[80] wl[121] vdd gnd cell_6t
Xbit_r122_c80 bl[80] br[80] wl[122] vdd gnd cell_6t
Xbit_r123_c80 bl[80] br[80] wl[123] vdd gnd cell_6t
Xbit_r124_c80 bl[80] br[80] wl[124] vdd gnd cell_6t
Xbit_r125_c80 bl[80] br[80] wl[125] vdd gnd cell_6t
Xbit_r126_c80 bl[80] br[80] wl[126] vdd gnd cell_6t
Xbit_r127_c80 bl[80] br[80] wl[127] vdd gnd cell_6t
Xbit_r128_c80 bl[80] br[80] wl[128] vdd gnd cell_6t
Xbit_r129_c80 bl[80] br[80] wl[129] vdd gnd cell_6t
Xbit_r130_c80 bl[80] br[80] wl[130] vdd gnd cell_6t
Xbit_r131_c80 bl[80] br[80] wl[131] vdd gnd cell_6t
Xbit_r132_c80 bl[80] br[80] wl[132] vdd gnd cell_6t
Xbit_r133_c80 bl[80] br[80] wl[133] vdd gnd cell_6t
Xbit_r134_c80 bl[80] br[80] wl[134] vdd gnd cell_6t
Xbit_r135_c80 bl[80] br[80] wl[135] vdd gnd cell_6t
Xbit_r136_c80 bl[80] br[80] wl[136] vdd gnd cell_6t
Xbit_r137_c80 bl[80] br[80] wl[137] vdd gnd cell_6t
Xbit_r138_c80 bl[80] br[80] wl[138] vdd gnd cell_6t
Xbit_r139_c80 bl[80] br[80] wl[139] vdd gnd cell_6t
Xbit_r140_c80 bl[80] br[80] wl[140] vdd gnd cell_6t
Xbit_r141_c80 bl[80] br[80] wl[141] vdd gnd cell_6t
Xbit_r142_c80 bl[80] br[80] wl[142] vdd gnd cell_6t
Xbit_r143_c80 bl[80] br[80] wl[143] vdd gnd cell_6t
Xbit_r144_c80 bl[80] br[80] wl[144] vdd gnd cell_6t
Xbit_r145_c80 bl[80] br[80] wl[145] vdd gnd cell_6t
Xbit_r146_c80 bl[80] br[80] wl[146] vdd gnd cell_6t
Xbit_r147_c80 bl[80] br[80] wl[147] vdd gnd cell_6t
Xbit_r148_c80 bl[80] br[80] wl[148] vdd gnd cell_6t
Xbit_r149_c80 bl[80] br[80] wl[149] vdd gnd cell_6t
Xbit_r150_c80 bl[80] br[80] wl[150] vdd gnd cell_6t
Xbit_r151_c80 bl[80] br[80] wl[151] vdd gnd cell_6t
Xbit_r152_c80 bl[80] br[80] wl[152] vdd gnd cell_6t
Xbit_r153_c80 bl[80] br[80] wl[153] vdd gnd cell_6t
Xbit_r154_c80 bl[80] br[80] wl[154] vdd gnd cell_6t
Xbit_r155_c80 bl[80] br[80] wl[155] vdd gnd cell_6t
Xbit_r156_c80 bl[80] br[80] wl[156] vdd gnd cell_6t
Xbit_r157_c80 bl[80] br[80] wl[157] vdd gnd cell_6t
Xbit_r158_c80 bl[80] br[80] wl[158] vdd gnd cell_6t
Xbit_r159_c80 bl[80] br[80] wl[159] vdd gnd cell_6t
Xbit_r160_c80 bl[80] br[80] wl[160] vdd gnd cell_6t
Xbit_r161_c80 bl[80] br[80] wl[161] vdd gnd cell_6t
Xbit_r162_c80 bl[80] br[80] wl[162] vdd gnd cell_6t
Xbit_r163_c80 bl[80] br[80] wl[163] vdd gnd cell_6t
Xbit_r164_c80 bl[80] br[80] wl[164] vdd gnd cell_6t
Xbit_r165_c80 bl[80] br[80] wl[165] vdd gnd cell_6t
Xbit_r166_c80 bl[80] br[80] wl[166] vdd gnd cell_6t
Xbit_r167_c80 bl[80] br[80] wl[167] vdd gnd cell_6t
Xbit_r168_c80 bl[80] br[80] wl[168] vdd gnd cell_6t
Xbit_r169_c80 bl[80] br[80] wl[169] vdd gnd cell_6t
Xbit_r170_c80 bl[80] br[80] wl[170] vdd gnd cell_6t
Xbit_r171_c80 bl[80] br[80] wl[171] vdd gnd cell_6t
Xbit_r172_c80 bl[80] br[80] wl[172] vdd gnd cell_6t
Xbit_r173_c80 bl[80] br[80] wl[173] vdd gnd cell_6t
Xbit_r174_c80 bl[80] br[80] wl[174] vdd gnd cell_6t
Xbit_r175_c80 bl[80] br[80] wl[175] vdd gnd cell_6t
Xbit_r176_c80 bl[80] br[80] wl[176] vdd gnd cell_6t
Xbit_r177_c80 bl[80] br[80] wl[177] vdd gnd cell_6t
Xbit_r178_c80 bl[80] br[80] wl[178] vdd gnd cell_6t
Xbit_r179_c80 bl[80] br[80] wl[179] vdd gnd cell_6t
Xbit_r180_c80 bl[80] br[80] wl[180] vdd gnd cell_6t
Xbit_r181_c80 bl[80] br[80] wl[181] vdd gnd cell_6t
Xbit_r182_c80 bl[80] br[80] wl[182] vdd gnd cell_6t
Xbit_r183_c80 bl[80] br[80] wl[183] vdd gnd cell_6t
Xbit_r184_c80 bl[80] br[80] wl[184] vdd gnd cell_6t
Xbit_r185_c80 bl[80] br[80] wl[185] vdd gnd cell_6t
Xbit_r186_c80 bl[80] br[80] wl[186] vdd gnd cell_6t
Xbit_r187_c80 bl[80] br[80] wl[187] vdd gnd cell_6t
Xbit_r188_c80 bl[80] br[80] wl[188] vdd gnd cell_6t
Xbit_r189_c80 bl[80] br[80] wl[189] vdd gnd cell_6t
Xbit_r190_c80 bl[80] br[80] wl[190] vdd gnd cell_6t
Xbit_r191_c80 bl[80] br[80] wl[191] vdd gnd cell_6t
Xbit_r192_c80 bl[80] br[80] wl[192] vdd gnd cell_6t
Xbit_r193_c80 bl[80] br[80] wl[193] vdd gnd cell_6t
Xbit_r194_c80 bl[80] br[80] wl[194] vdd gnd cell_6t
Xbit_r195_c80 bl[80] br[80] wl[195] vdd gnd cell_6t
Xbit_r196_c80 bl[80] br[80] wl[196] vdd gnd cell_6t
Xbit_r197_c80 bl[80] br[80] wl[197] vdd gnd cell_6t
Xbit_r198_c80 bl[80] br[80] wl[198] vdd gnd cell_6t
Xbit_r199_c80 bl[80] br[80] wl[199] vdd gnd cell_6t
Xbit_r200_c80 bl[80] br[80] wl[200] vdd gnd cell_6t
Xbit_r201_c80 bl[80] br[80] wl[201] vdd gnd cell_6t
Xbit_r202_c80 bl[80] br[80] wl[202] vdd gnd cell_6t
Xbit_r203_c80 bl[80] br[80] wl[203] vdd gnd cell_6t
Xbit_r204_c80 bl[80] br[80] wl[204] vdd gnd cell_6t
Xbit_r205_c80 bl[80] br[80] wl[205] vdd gnd cell_6t
Xbit_r206_c80 bl[80] br[80] wl[206] vdd gnd cell_6t
Xbit_r207_c80 bl[80] br[80] wl[207] vdd gnd cell_6t
Xbit_r208_c80 bl[80] br[80] wl[208] vdd gnd cell_6t
Xbit_r209_c80 bl[80] br[80] wl[209] vdd gnd cell_6t
Xbit_r210_c80 bl[80] br[80] wl[210] vdd gnd cell_6t
Xbit_r211_c80 bl[80] br[80] wl[211] vdd gnd cell_6t
Xbit_r212_c80 bl[80] br[80] wl[212] vdd gnd cell_6t
Xbit_r213_c80 bl[80] br[80] wl[213] vdd gnd cell_6t
Xbit_r214_c80 bl[80] br[80] wl[214] vdd gnd cell_6t
Xbit_r215_c80 bl[80] br[80] wl[215] vdd gnd cell_6t
Xbit_r216_c80 bl[80] br[80] wl[216] vdd gnd cell_6t
Xbit_r217_c80 bl[80] br[80] wl[217] vdd gnd cell_6t
Xbit_r218_c80 bl[80] br[80] wl[218] vdd gnd cell_6t
Xbit_r219_c80 bl[80] br[80] wl[219] vdd gnd cell_6t
Xbit_r220_c80 bl[80] br[80] wl[220] vdd gnd cell_6t
Xbit_r221_c80 bl[80] br[80] wl[221] vdd gnd cell_6t
Xbit_r222_c80 bl[80] br[80] wl[222] vdd gnd cell_6t
Xbit_r223_c80 bl[80] br[80] wl[223] vdd gnd cell_6t
Xbit_r224_c80 bl[80] br[80] wl[224] vdd gnd cell_6t
Xbit_r225_c80 bl[80] br[80] wl[225] vdd gnd cell_6t
Xbit_r226_c80 bl[80] br[80] wl[226] vdd gnd cell_6t
Xbit_r227_c80 bl[80] br[80] wl[227] vdd gnd cell_6t
Xbit_r228_c80 bl[80] br[80] wl[228] vdd gnd cell_6t
Xbit_r229_c80 bl[80] br[80] wl[229] vdd gnd cell_6t
Xbit_r230_c80 bl[80] br[80] wl[230] vdd gnd cell_6t
Xbit_r231_c80 bl[80] br[80] wl[231] vdd gnd cell_6t
Xbit_r232_c80 bl[80] br[80] wl[232] vdd gnd cell_6t
Xbit_r233_c80 bl[80] br[80] wl[233] vdd gnd cell_6t
Xbit_r234_c80 bl[80] br[80] wl[234] vdd gnd cell_6t
Xbit_r235_c80 bl[80] br[80] wl[235] vdd gnd cell_6t
Xbit_r236_c80 bl[80] br[80] wl[236] vdd gnd cell_6t
Xbit_r237_c80 bl[80] br[80] wl[237] vdd gnd cell_6t
Xbit_r238_c80 bl[80] br[80] wl[238] vdd gnd cell_6t
Xbit_r239_c80 bl[80] br[80] wl[239] vdd gnd cell_6t
Xbit_r240_c80 bl[80] br[80] wl[240] vdd gnd cell_6t
Xbit_r241_c80 bl[80] br[80] wl[241] vdd gnd cell_6t
Xbit_r242_c80 bl[80] br[80] wl[242] vdd gnd cell_6t
Xbit_r243_c80 bl[80] br[80] wl[243] vdd gnd cell_6t
Xbit_r244_c80 bl[80] br[80] wl[244] vdd gnd cell_6t
Xbit_r245_c80 bl[80] br[80] wl[245] vdd gnd cell_6t
Xbit_r246_c80 bl[80] br[80] wl[246] vdd gnd cell_6t
Xbit_r247_c80 bl[80] br[80] wl[247] vdd gnd cell_6t
Xbit_r248_c80 bl[80] br[80] wl[248] vdd gnd cell_6t
Xbit_r249_c80 bl[80] br[80] wl[249] vdd gnd cell_6t
Xbit_r250_c80 bl[80] br[80] wl[250] vdd gnd cell_6t
Xbit_r251_c80 bl[80] br[80] wl[251] vdd gnd cell_6t
Xbit_r252_c80 bl[80] br[80] wl[252] vdd gnd cell_6t
Xbit_r253_c80 bl[80] br[80] wl[253] vdd gnd cell_6t
Xbit_r254_c80 bl[80] br[80] wl[254] vdd gnd cell_6t
Xbit_r255_c80 bl[80] br[80] wl[255] vdd gnd cell_6t
Xbit_r256_c80 bl[80] br[80] wl[256] vdd gnd cell_6t
Xbit_r257_c80 bl[80] br[80] wl[257] vdd gnd cell_6t
Xbit_r258_c80 bl[80] br[80] wl[258] vdd gnd cell_6t
Xbit_r259_c80 bl[80] br[80] wl[259] vdd gnd cell_6t
Xbit_r260_c80 bl[80] br[80] wl[260] vdd gnd cell_6t
Xbit_r261_c80 bl[80] br[80] wl[261] vdd gnd cell_6t
Xbit_r262_c80 bl[80] br[80] wl[262] vdd gnd cell_6t
Xbit_r263_c80 bl[80] br[80] wl[263] vdd gnd cell_6t
Xbit_r264_c80 bl[80] br[80] wl[264] vdd gnd cell_6t
Xbit_r265_c80 bl[80] br[80] wl[265] vdd gnd cell_6t
Xbit_r266_c80 bl[80] br[80] wl[266] vdd gnd cell_6t
Xbit_r267_c80 bl[80] br[80] wl[267] vdd gnd cell_6t
Xbit_r268_c80 bl[80] br[80] wl[268] vdd gnd cell_6t
Xbit_r269_c80 bl[80] br[80] wl[269] vdd gnd cell_6t
Xbit_r270_c80 bl[80] br[80] wl[270] vdd gnd cell_6t
Xbit_r271_c80 bl[80] br[80] wl[271] vdd gnd cell_6t
Xbit_r272_c80 bl[80] br[80] wl[272] vdd gnd cell_6t
Xbit_r273_c80 bl[80] br[80] wl[273] vdd gnd cell_6t
Xbit_r274_c80 bl[80] br[80] wl[274] vdd gnd cell_6t
Xbit_r275_c80 bl[80] br[80] wl[275] vdd gnd cell_6t
Xbit_r276_c80 bl[80] br[80] wl[276] vdd gnd cell_6t
Xbit_r277_c80 bl[80] br[80] wl[277] vdd gnd cell_6t
Xbit_r278_c80 bl[80] br[80] wl[278] vdd gnd cell_6t
Xbit_r279_c80 bl[80] br[80] wl[279] vdd gnd cell_6t
Xbit_r280_c80 bl[80] br[80] wl[280] vdd gnd cell_6t
Xbit_r281_c80 bl[80] br[80] wl[281] vdd gnd cell_6t
Xbit_r282_c80 bl[80] br[80] wl[282] vdd gnd cell_6t
Xbit_r283_c80 bl[80] br[80] wl[283] vdd gnd cell_6t
Xbit_r284_c80 bl[80] br[80] wl[284] vdd gnd cell_6t
Xbit_r285_c80 bl[80] br[80] wl[285] vdd gnd cell_6t
Xbit_r286_c80 bl[80] br[80] wl[286] vdd gnd cell_6t
Xbit_r287_c80 bl[80] br[80] wl[287] vdd gnd cell_6t
Xbit_r288_c80 bl[80] br[80] wl[288] vdd gnd cell_6t
Xbit_r289_c80 bl[80] br[80] wl[289] vdd gnd cell_6t
Xbit_r290_c80 bl[80] br[80] wl[290] vdd gnd cell_6t
Xbit_r291_c80 bl[80] br[80] wl[291] vdd gnd cell_6t
Xbit_r292_c80 bl[80] br[80] wl[292] vdd gnd cell_6t
Xbit_r293_c80 bl[80] br[80] wl[293] vdd gnd cell_6t
Xbit_r294_c80 bl[80] br[80] wl[294] vdd gnd cell_6t
Xbit_r295_c80 bl[80] br[80] wl[295] vdd gnd cell_6t
Xbit_r296_c80 bl[80] br[80] wl[296] vdd gnd cell_6t
Xbit_r297_c80 bl[80] br[80] wl[297] vdd gnd cell_6t
Xbit_r298_c80 bl[80] br[80] wl[298] vdd gnd cell_6t
Xbit_r299_c80 bl[80] br[80] wl[299] vdd gnd cell_6t
Xbit_r300_c80 bl[80] br[80] wl[300] vdd gnd cell_6t
Xbit_r301_c80 bl[80] br[80] wl[301] vdd gnd cell_6t
Xbit_r302_c80 bl[80] br[80] wl[302] vdd gnd cell_6t
Xbit_r303_c80 bl[80] br[80] wl[303] vdd gnd cell_6t
Xbit_r304_c80 bl[80] br[80] wl[304] vdd gnd cell_6t
Xbit_r305_c80 bl[80] br[80] wl[305] vdd gnd cell_6t
Xbit_r306_c80 bl[80] br[80] wl[306] vdd gnd cell_6t
Xbit_r307_c80 bl[80] br[80] wl[307] vdd gnd cell_6t
Xbit_r308_c80 bl[80] br[80] wl[308] vdd gnd cell_6t
Xbit_r309_c80 bl[80] br[80] wl[309] vdd gnd cell_6t
Xbit_r310_c80 bl[80] br[80] wl[310] vdd gnd cell_6t
Xbit_r311_c80 bl[80] br[80] wl[311] vdd gnd cell_6t
Xbit_r312_c80 bl[80] br[80] wl[312] vdd gnd cell_6t
Xbit_r313_c80 bl[80] br[80] wl[313] vdd gnd cell_6t
Xbit_r314_c80 bl[80] br[80] wl[314] vdd gnd cell_6t
Xbit_r315_c80 bl[80] br[80] wl[315] vdd gnd cell_6t
Xbit_r316_c80 bl[80] br[80] wl[316] vdd gnd cell_6t
Xbit_r317_c80 bl[80] br[80] wl[317] vdd gnd cell_6t
Xbit_r318_c80 bl[80] br[80] wl[318] vdd gnd cell_6t
Xbit_r319_c80 bl[80] br[80] wl[319] vdd gnd cell_6t
Xbit_r320_c80 bl[80] br[80] wl[320] vdd gnd cell_6t
Xbit_r321_c80 bl[80] br[80] wl[321] vdd gnd cell_6t
Xbit_r322_c80 bl[80] br[80] wl[322] vdd gnd cell_6t
Xbit_r323_c80 bl[80] br[80] wl[323] vdd gnd cell_6t
Xbit_r324_c80 bl[80] br[80] wl[324] vdd gnd cell_6t
Xbit_r325_c80 bl[80] br[80] wl[325] vdd gnd cell_6t
Xbit_r326_c80 bl[80] br[80] wl[326] vdd gnd cell_6t
Xbit_r327_c80 bl[80] br[80] wl[327] vdd gnd cell_6t
Xbit_r328_c80 bl[80] br[80] wl[328] vdd gnd cell_6t
Xbit_r329_c80 bl[80] br[80] wl[329] vdd gnd cell_6t
Xbit_r330_c80 bl[80] br[80] wl[330] vdd gnd cell_6t
Xbit_r331_c80 bl[80] br[80] wl[331] vdd gnd cell_6t
Xbit_r332_c80 bl[80] br[80] wl[332] vdd gnd cell_6t
Xbit_r333_c80 bl[80] br[80] wl[333] vdd gnd cell_6t
Xbit_r334_c80 bl[80] br[80] wl[334] vdd gnd cell_6t
Xbit_r335_c80 bl[80] br[80] wl[335] vdd gnd cell_6t
Xbit_r336_c80 bl[80] br[80] wl[336] vdd gnd cell_6t
Xbit_r337_c80 bl[80] br[80] wl[337] vdd gnd cell_6t
Xbit_r338_c80 bl[80] br[80] wl[338] vdd gnd cell_6t
Xbit_r339_c80 bl[80] br[80] wl[339] vdd gnd cell_6t
Xbit_r340_c80 bl[80] br[80] wl[340] vdd gnd cell_6t
Xbit_r341_c80 bl[80] br[80] wl[341] vdd gnd cell_6t
Xbit_r342_c80 bl[80] br[80] wl[342] vdd gnd cell_6t
Xbit_r343_c80 bl[80] br[80] wl[343] vdd gnd cell_6t
Xbit_r344_c80 bl[80] br[80] wl[344] vdd gnd cell_6t
Xbit_r345_c80 bl[80] br[80] wl[345] vdd gnd cell_6t
Xbit_r346_c80 bl[80] br[80] wl[346] vdd gnd cell_6t
Xbit_r347_c80 bl[80] br[80] wl[347] vdd gnd cell_6t
Xbit_r348_c80 bl[80] br[80] wl[348] vdd gnd cell_6t
Xbit_r349_c80 bl[80] br[80] wl[349] vdd gnd cell_6t
Xbit_r350_c80 bl[80] br[80] wl[350] vdd gnd cell_6t
Xbit_r351_c80 bl[80] br[80] wl[351] vdd gnd cell_6t
Xbit_r352_c80 bl[80] br[80] wl[352] vdd gnd cell_6t
Xbit_r353_c80 bl[80] br[80] wl[353] vdd gnd cell_6t
Xbit_r354_c80 bl[80] br[80] wl[354] vdd gnd cell_6t
Xbit_r355_c80 bl[80] br[80] wl[355] vdd gnd cell_6t
Xbit_r356_c80 bl[80] br[80] wl[356] vdd gnd cell_6t
Xbit_r357_c80 bl[80] br[80] wl[357] vdd gnd cell_6t
Xbit_r358_c80 bl[80] br[80] wl[358] vdd gnd cell_6t
Xbit_r359_c80 bl[80] br[80] wl[359] vdd gnd cell_6t
Xbit_r360_c80 bl[80] br[80] wl[360] vdd gnd cell_6t
Xbit_r361_c80 bl[80] br[80] wl[361] vdd gnd cell_6t
Xbit_r362_c80 bl[80] br[80] wl[362] vdd gnd cell_6t
Xbit_r363_c80 bl[80] br[80] wl[363] vdd gnd cell_6t
Xbit_r364_c80 bl[80] br[80] wl[364] vdd gnd cell_6t
Xbit_r365_c80 bl[80] br[80] wl[365] vdd gnd cell_6t
Xbit_r366_c80 bl[80] br[80] wl[366] vdd gnd cell_6t
Xbit_r367_c80 bl[80] br[80] wl[367] vdd gnd cell_6t
Xbit_r368_c80 bl[80] br[80] wl[368] vdd gnd cell_6t
Xbit_r369_c80 bl[80] br[80] wl[369] vdd gnd cell_6t
Xbit_r370_c80 bl[80] br[80] wl[370] vdd gnd cell_6t
Xbit_r371_c80 bl[80] br[80] wl[371] vdd gnd cell_6t
Xbit_r372_c80 bl[80] br[80] wl[372] vdd gnd cell_6t
Xbit_r373_c80 bl[80] br[80] wl[373] vdd gnd cell_6t
Xbit_r374_c80 bl[80] br[80] wl[374] vdd gnd cell_6t
Xbit_r375_c80 bl[80] br[80] wl[375] vdd gnd cell_6t
Xbit_r376_c80 bl[80] br[80] wl[376] vdd gnd cell_6t
Xbit_r377_c80 bl[80] br[80] wl[377] vdd gnd cell_6t
Xbit_r378_c80 bl[80] br[80] wl[378] vdd gnd cell_6t
Xbit_r379_c80 bl[80] br[80] wl[379] vdd gnd cell_6t
Xbit_r380_c80 bl[80] br[80] wl[380] vdd gnd cell_6t
Xbit_r381_c80 bl[80] br[80] wl[381] vdd gnd cell_6t
Xbit_r382_c80 bl[80] br[80] wl[382] vdd gnd cell_6t
Xbit_r383_c80 bl[80] br[80] wl[383] vdd gnd cell_6t
Xbit_r384_c80 bl[80] br[80] wl[384] vdd gnd cell_6t
Xbit_r385_c80 bl[80] br[80] wl[385] vdd gnd cell_6t
Xbit_r386_c80 bl[80] br[80] wl[386] vdd gnd cell_6t
Xbit_r387_c80 bl[80] br[80] wl[387] vdd gnd cell_6t
Xbit_r388_c80 bl[80] br[80] wl[388] vdd gnd cell_6t
Xbit_r389_c80 bl[80] br[80] wl[389] vdd gnd cell_6t
Xbit_r390_c80 bl[80] br[80] wl[390] vdd gnd cell_6t
Xbit_r391_c80 bl[80] br[80] wl[391] vdd gnd cell_6t
Xbit_r392_c80 bl[80] br[80] wl[392] vdd gnd cell_6t
Xbit_r393_c80 bl[80] br[80] wl[393] vdd gnd cell_6t
Xbit_r394_c80 bl[80] br[80] wl[394] vdd gnd cell_6t
Xbit_r395_c80 bl[80] br[80] wl[395] vdd gnd cell_6t
Xbit_r396_c80 bl[80] br[80] wl[396] vdd gnd cell_6t
Xbit_r397_c80 bl[80] br[80] wl[397] vdd gnd cell_6t
Xbit_r398_c80 bl[80] br[80] wl[398] vdd gnd cell_6t
Xbit_r399_c80 bl[80] br[80] wl[399] vdd gnd cell_6t
Xbit_r400_c80 bl[80] br[80] wl[400] vdd gnd cell_6t
Xbit_r401_c80 bl[80] br[80] wl[401] vdd gnd cell_6t
Xbit_r402_c80 bl[80] br[80] wl[402] vdd gnd cell_6t
Xbit_r403_c80 bl[80] br[80] wl[403] vdd gnd cell_6t
Xbit_r404_c80 bl[80] br[80] wl[404] vdd gnd cell_6t
Xbit_r405_c80 bl[80] br[80] wl[405] vdd gnd cell_6t
Xbit_r406_c80 bl[80] br[80] wl[406] vdd gnd cell_6t
Xbit_r407_c80 bl[80] br[80] wl[407] vdd gnd cell_6t
Xbit_r408_c80 bl[80] br[80] wl[408] vdd gnd cell_6t
Xbit_r409_c80 bl[80] br[80] wl[409] vdd gnd cell_6t
Xbit_r410_c80 bl[80] br[80] wl[410] vdd gnd cell_6t
Xbit_r411_c80 bl[80] br[80] wl[411] vdd gnd cell_6t
Xbit_r412_c80 bl[80] br[80] wl[412] vdd gnd cell_6t
Xbit_r413_c80 bl[80] br[80] wl[413] vdd gnd cell_6t
Xbit_r414_c80 bl[80] br[80] wl[414] vdd gnd cell_6t
Xbit_r415_c80 bl[80] br[80] wl[415] vdd gnd cell_6t
Xbit_r416_c80 bl[80] br[80] wl[416] vdd gnd cell_6t
Xbit_r417_c80 bl[80] br[80] wl[417] vdd gnd cell_6t
Xbit_r418_c80 bl[80] br[80] wl[418] vdd gnd cell_6t
Xbit_r419_c80 bl[80] br[80] wl[419] vdd gnd cell_6t
Xbit_r420_c80 bl[80] br[80] wl[420] vdd gnd cell_6t
Xbit_r421_c80 bl[80] br[80] wl[421] vdd gnd cell_6t
Xbit_r422_c80 bl[80] br[80] wl[422] vdd gnd cell_6t
Xbit_r423_c80 bl[80] br[80] wl[423] vdd gnd cell_6t
Xbit_r424_c80 bl[80] br[80] wl[424] vdd gnd cell_6t
Xbit_r425_c80 bl[80] br[80] wl[425] vdd gnd cell_6t
Xbit_r426_c80 bl[80] br[80] wl[426] vdd gnd cell_6t
Xbit_r427_c80 bl[80] br[80] wl[427] vdd gnd cell_6t
Xbit_r428_c80 bl[80] br[80] wl[428] vdd gnd cell_6t
Xbit_r429_c80 bl[80] br[80] wl[429] vdd gnd cell_6t
Xbit_r430_c80 bl[80] br[80] wl[430] vdd gnd cell_6t
Xbit_r431_c80 bl[80] br[80] wl[431] vdd gnd cell_6t
Xbit_r432_c80 bl[80] br[80] wl[432] vdd gnd cell_6t
Xbit_r433_c80 bl[80] br[80] wl[433] vdd gnd cell_6t
Xbit_r434_c80 bl[80] br[80] wl[434] vdd gnd cell_6t
Xbit_r435_c80 bl[80] br[80] wl[435] vdd gnd cell_6t
Xbit_r436_c80 bl[80] br[80] wl[436] vdd gnd cell_6t
Xbit_r437_c80 bl[80] br[80] wl[437] vdd gnd cell_6t
Xbit_r438_c80 bl[80] br[80] wl[438] vdd gnd cell_6t
Xbit_r439_c80 bl[80] br[80] wl[439] vdd gnd cell_6t
Xbit_r440_c80 bl[80] br[80] wl[440] vdd gnd cell_6t
Xbit_r441_c80 bl[80] br[80] wl[441] vdd gnd cell_6t
Xbit_r442_c80 bl[80] br[80] wl[442] vdd gnd cell_6t
Xbit_r443_c80 bl[80] br[80] wl[443] vdd gnd cell_6t
Xbit_r444_c80 bl[80] br[80] wl[444] vdd gnd cell_6t
Xbit_r445_c80 bl[80] br[80] wl[445] vdd gnd cell_6t
Xbit_r446_c80 bl[80] br[80] wl[446] vdd gnd cell_6t
Xbit_r447_c80 bl[80] br[80] wl[447] vdd gnd cell_6t
Xbit_r448_c80 bl[80] br[80] wl[448] vdd gnd cell_6t
Xbit_r449_c80 bl[80] br[80] wl[449] vdd gnd cell_6t
Xbit_r450_c80 bl[80] br[80] wl[450] vdd gnd cell_6t
Xbit_r451_c80 bl[80] br[80] wl[451] vdd gnd cell_6t
Xbit_r452_c80 bl[80] br[80] wl[452] vdd gnd cell_6t
Xbit_r453_c80 bl[80] br[80] wl[453] vdd gnd cell_6t
Xbit_r454_c80 bl[80] br[80] wl[454] vdd gnd cell_6t
Xbit_r455_c80 bl[80] br[80] wl[455] vdd gnd cell_6t
Xbit_r456_c80 bl[80] br[80] wl[456] vdd gnd cell_6t
Xbit_r457_c80 bl[80] br[80] wl[457] vdd gnd cell_6t
Xbit_r458_c80 bl[80] br[80] wl[458] vdd gnd cell_6t
Xbit_r459_c80 bl[80] br[80] wl[459] vdd gnd cell_6t
Xbit_r460_c80 bl[80] br[80] wl[460] vdd gnd cell_6t
Xbit_r461_c80 bl[80] br[80] wl[461] vdd gnd cell_6t
Xbit_r462_c80 bl[80] br[80] wl[462] vdd gnd cell_6t
Xbit_r463_c80 bl[80] br[80] wl[463] vdd gnd cell_6t
Xbit_r464_c80 bl[80] br[80] wl[464] vdd gnd cell_6t
Xbit_r465_c80 bl[80] br[80] wl[465] vdd gnd cell_6t
Xbit_r466_c80 bl[80] br[80] wl[466] vdd gnd cell_6t
Xbit_r467_c80 bl[80] br[80] wl[467] vdd gnd cell_6t
Xbit_r468_c80 bl[80] br[80] wl[468] vdd gnd cell_6t
Xbit_r469_c80 bl[80] br[80] wl[469] vdd gnd cell_6t
Xbit_r470_c80 bl[80] br[80] wl[470] vdd gnd cell_6t
Xbit_r471_c80 bl[80] br[80] wl[471] vdd gnd cell_6t
Xbit_r472_c80 bl[80] br[80] wl[472] vdd gnd cell_6t
Xbit_r473_c80 bl[80] br[80] wl[473] vdd gnd cell_6t
Xbit_r474_c80 bl[80] br[80] wl[474] vdd gnd cell_6t
Xbit_r475_c80 bl[80] br[80] wl[475] vdd gnd cell_6t
Xbit_r476_c80 bl[80] br[80] wl[476] vdd gnd cell_6t
Xbit_r477_c80 bl[80] br[80] wl[477] vdd gnd cell_6t
Xbit_r478_c80 bl[80] br[80] wl[478] vdd gnd cell_6t
Xbit_r479_c80 bl[80] br[80] wl[479] vdd gnd cell_6t
Xbit_r480_c80 bl[80] br[80] wl[480] vdd gnd cell_6t
Xbit_r481_c80 bl[80] br[80] wl[481] vdd gnd cell_6t
Xbit_r482_c80 bl[80] br[80] wl[482] vdd gnd cell_6t
Xbit_r483_c80 bl[80] br[80] wl[483] vdd gnd cell_6t
Xbit_r484_c80 bl[80] br[80] wl[484] vdd gnd cell_6t
Xbit_r485_c80 bl[80] br[80] wl[485] vdd gnd cell_6t
Xbit_r486_c80 bl[80] br[80] wl[486] vdd gnd cell_6t
Xbit_r487_c80 bl[80] br[80] wl[487] vdd gnd cell_6t
Xbit_r488_c80 bl[80] br[80] wl[488] vdd gnd cell_6t
Xbit_r489_c80 bl[80] br[80] wl[489] vdd gnd cell_6t
Xbit_r490_c80 bl[80] br[80] wl[490] vdd gnd cell_6t
Xbit_r491_c80 bl[80] br[80] wl[491] vdd gnd cell_6t
Xbit_r492_c80 bl[80] br[80] wl[492] vdd gnd cell_6t
Xbit_r493_c80 bl[80] br[80] wl[493] vdd gnd cell_6t
Xbit_r494_c80 bl[80] br[80] wl[494] vdd gnd cell_6t
Xbit_r495_c80 bl[80] br[80] wl[495] vdd gnd cell_6t
Xbit_r496_c80 bl[80] br[80] wl[496] vdd gnd cell_6t
Xbit_r497_c80 bl[80] br[80] wl[497] vdd gnd cell_6t
Xbit_r498_c80 bl[80] br[80] wl[498] vdd gnd cell_6t
Xbit_r499_c80 bl[80] br[80] wl[499] vdd gnd cell_6t
Xbit_r500_c80 bl[80] br[80] wl[500] vdd gnd cell_6t
Xbit_r501_c80 bl[80] br[80] wl[501] vdd gnd cell_6t
Xbit_r502_c80 bl[80] br[80] wl[502] vdd gnd cell_6t
Xbit_r503_c80 bl[80] br[80] wl[503] vdd gnd cell_6t
Xbit_r504_c80 bl[80] br[80] wl[504] vdd gnd cell_6t
Xbit_r505_c80 bl[80] br[80] wl[505] vdd gnd cell_6t
Xbit_r506_c80 bl[80] br[80] wl[506] vdd gnd cell_6t
Xbit_r507_c80 bl[80] br[80] wl[507] vdd gnd cell_6t
Xbit_r508_c80 bl[80] br[80] wl[508] vdd gnd cell_6t
Xbit_r509_c80 bl[80] br[80] wl[509] vdd gnd cell_6t
Xbit_r510_c80 bl[80] br[80] wl[510] vdd gnd cell_6t
Xbit_r511_c80 bl[80] br[80] wl[511] vdd gnd cell_6t
Xbit_r0_c81 bl[81] br[81] wl[0] vdd gnd cell_6t
Xbit_r1_c81 bl[81] br[81] wl[1] vdd gnd cell_6t
Xbit_r2_c81 bl[81] br[81] wl[2] vdd gnd cell_6t
Xbit_r3_c81 bl[81] br[81] wl[3] vdd gnd cell_6t
Xbit_r4_c81 bl[81] br[81] wl[4] vdd gnd cell_6t
Xbit_r5_c81 bl[81] br[81] wl[5] vdd gnd cell_6t
Xbit_r6_c81 bl[81] br[81] wl[6] vdd gnd cell_6t
Xbit_r7_c81 bl[81] br[81] wl[7] vdd gnd cell_6t
Xbit_r8_c81 bl[81] br[81] wl[8] vdd gnd cell_6t
Xbit_r9_c81 bl[81] br[81] wl[9] vdd gnd cell_6t
Xbit_r10_c81 bl[81] br[81] wl[10] vdd gnd cell_6t
Xbit_r11_c81 bl[81] br[81] wl[11] vdd gnd cell_6t
Xbit_r12_c81 bl[81] br[81] wl[12] vdd gnd cell_6t
Xbit_r13_c81 bl[81] br[81] wl[13] vdd gnd cell_6t
Xbit_r14_c81 bl[81] br[81] wl[14] vdd gnd cell_6t
Xbit_r15_c81 bl[81] br[81] wl[15] vdd gnd cell_6t
Xbit_r16_c81 bl[81] br[81] wl[16] vdd gnd cell_6t
Xbit_r17_c81 bl[81] br[81] wl[17] vdd gnd cell_6t
Xbit_r18_c81 bl[81] br[81] wl[18] vdd gnd cell_6t
Xbit_r19_c81 bl[81] br[81] wl[19] vdd gnd cell_6t
Xbit_r20_c81 bl[81] br[81] wl[20] vdd gnd cell_6t
Xbit_r21_c81 bl[81] br[81] wl[21] vdd gnd cell_6t
Xbit_r22_c81 bl[81] br[81] wl[22] vdd gnd cell_6t
Xbit_r23_c81 bl[81] br[81] wl[23] vdd gnd cell_6t
Xbit_r24_c81 bl[81] br[81] wl[24] vdd gnd cell_6t
Xbit_r25_c81 bl[81] br[81] wl[25] vdd gnd cell_6t
Xbit_r26_c81 bl[81] br[81] wl[26] vdd gnd cell_6t
Xbit_r27_c81 bl[81] br[81] wl[27] vdd gnd cell_6t
Xbit_r28_c81 bl[81] br[81] wl[28] vdd gnd cell_6t
Xbit_r29_c81 bl[81] br[81] wl[29] vdd gnd cell_6t
Xbit_r30_c81 bl[81] br[81] wl[30] vdd gnd cell_6t
Xbit_r31_c81 bl[81] br[81] wl[31] vdd gnd cell_6t
Xbit_r32_c81 bl[81] br[81] wl[32] vdd gnd cell_6t
Xbit_r33_c81 bl[81] br[81] wl[33] vdd gnd cell_6t
Xbit_r34_c81 bl[81] br[81] wl[34] vdd gnd cell_6t
Xbit_r35_c81 bl[81] br[81] wl[35] vdd gnd cell_6t
Xbit_r36_c81 bl[81] br[81] wl[36] vdd gnd cell_6t
Xbit_r37_c81 bl[81] br[81] wl[37] vdd gnd cell_6t
Xbit_r38_c81 bl[81] br[81] wl[38] vdd gnd cell_6t
Xbit_r39_c81 bl[81] br[81] wl[39] vdd gnd cell_6t
Xbit_r40_c81 bl[81] br[81] wl[40] vdd gnd cell_6t
Xbit_r41_c81 bl[81] br[81] wl[41] vdd gnd cell_6t
Xbit_r42_c81 bl[81] br[81] wl[42] vdd gnd cell_6t
Xbit_r43_c81 bl[81] br[81] wl[43] vdd gnd cell_6t
Xbit_r44_c81 bl[81] br[81] wl[44] vdd gnd cell_6t
Xbit_r45_c81 bl[81] br[81] wl[45] vdd gnd cell_6t
Xbit_r46_c81 bl[81] br[81] wl[46] vdd gnd cell_6t
Xbit_r47_c81 bl[81] br[81] wl[47] vdd gnd cell_6t
Xbit_r48_c81 bl[81] br[81] wl[48] vdd gnd cell_6t
Xbit_r49_c81 bl[81] br[81] wl[49] vdd gnd cell_6t
Xbit_r50_c81 bl[81] br[81] wl[50] vdd gnd cell_6t
Xbit_r51_c81 bl[81] br[81] wl[51] vdd gnd cell_6t
Xbit_r52_c81 bl[81] br[81] wl[52] vdd gnd cell_6t
Xbit_r53_c81 bl[81] br[81] wl[53] vdd gnd cell_6t
Xbit_r54_c81 bl[81] br[81] wl[54] vdd gnd cell_6t
Xbit_r55_c81 bl[81] br[81] wl[55] vdd gnd cell_6t
Xbit_r56_c81 bl[81] br[81] wl[56] vdd gnd cell_6t
Xbit_r57_c81 bl[81] br[81] wl[57] vdd gnd cell_6t
Xbit_r58_c81 bl[81] br[81] wl[58] vdd gnd cell_6t
Xbit_r59_c81 bl[81] br[81] wl[59] vdd gnd cell_6t
Xbit_r60_c81 bl[81] br[81] wl[60] vdd gnd cell_6t
Xbit_r61_c81 bl[81] br[81] wl[61] vdd gnd cell_6t
Xbit_r62_c81 bl[81] br[81] wl[62] vdd gnd cell_6t
Xbit_r63_c81 bl[81] br[81] wl[63] vdd gnd cell_6t
Xbit_r64_c81 bl[81] br[81] wl[64] vdd gnd cell_6t
Xbit_r65_c81 bl[81] br[81] wl[65] vdd gnd cell_6t
Xbit_r66_c81 bl[81] br[81] wl[66] vdd gnd cell_6t
Xbit_r67_c81 bl[81] br[81] wl[67] vdd gnd cell_6t
Xbit_r68_c81 bl[81] br[81] wl[68] vdd gnd cell_6t
Xbit_r69_c81 bl[81] br[81] wl[69] vdd gnd cell_6t
Xbit_r70_c81 bl[81] br[81] wl[70] vdd gnd cell_6t
Xbit_r71_c81 bl[81] br[81] wl[71] vdd gnd cell_6t
Xbit_r72_c81 bl[81] br[81] wl[72] vdd gnd cell_6t
Xbit_r73_c81 bl[81] br[81] wl[73] vdd gnd cell_6t
Xbit_r74_c81 bl[81] br[81] wl[74] vdd gnd cell_6t
Xbit_r75_c81 bl[81] br[81] wl[75] vdd gnd cell_6t
Xbit_r76_c81 bl[81] br[81] wl[76] vdd gnd cell_6t
Xbit_r77_c81 bl[81] br[81] wl[77] vdd gnd cell_6t
Xbit_r78_c81 bl[81] br[81] wl[78] vdd gnd cell_6t
Xbit_r79_c81 bl[81] br[81] wl[79] vdd gnd cell_6t
Xbit_r80_c81 bl[81] br[81] wl[80] vdd gnd cell_6t
Xbit_r81_c81 bl[81] br[81] wl[81] vdd gnd cell_6t
Xbit_r82_c81 bl[81] br[81] wl[82] vdd gnd cell_6t
Xbit_r83_c81 bl[81] br[81] wl[83] vdd gnd cell_6t
Xbit_r84_c81 bl[81] br[81] wl[84] vdd gnd cell_6t
Xbit_r85_c81 bl[81] br[81] wl[85] vdd gnd cell_6t
Xbit_r86_c81 bl[81] br[81] wl[86] vdd gnd cell_6t
Xbit_r87_c81 bl[81] br[81] wl[87] vdd gnd cell_6t
Xbit_r88_c81 bl[81] br[81] wl[88] vdd gnd cell_6t
Xbit_r89_c81 bl[81] br[81] wl[89] vdd gnd cell_6t
Xbit_r90_c81 bl[81] br[81] wl[90] vdd gnd cell_6t
Xbit_r91_c81 bl[81] br[81] wl[91] vdd gnd cell_6t
Xbit_r92_c81 bl[81] br[81] wl[92] vdd gnd cell_6t
Xbit_r93_c81 bl[81] br[81] wl[93] vdd gnd cell_6t
Xbit_r94_c81 bl[81] br[81] wl[94] vdd gnd cell_6t
Xbit_r95_c81 bl[81] br[81] wl[95] vdd gnd cell_6t
Xbit_r96_c81 bl[81] br[81] wl[96] vdd gnd cell_6t
Xbit_r97_c81 bl[81] br[81] wl[97] vdd gnd cell_6t
Xbit_r98_c81 bl[81] br[81] wl[98] vdd gnd cell_6t
Xbit_r99_c81 bl[81] br[81] wl[99] vdd gnd cell_6t
Xbit_r100_c81 bl[81] br[81] wl[100] vdd gnd cell_6t
Xbit_r101_c81 bl[81] br[81] wl[101] vdd gnd cell_6t
Xbit_r102_c81 bl[81] br[81] wl[102] vdd gnd cell_6t
Xbit_r103_c81 bl[81] br[81] wl[103] vdd gnd cell_6t
Xbit_r104_c81 bl[81] br[81] wl[104] vdd gnd cell_6t
Xbit_r105_c81 bl[81] br[81] wl[105] vdd gnd cell_6t
Xbit_r106_c81 bl[81] br[81] wl[106] vdd gnd cell_6t
Xbit_r107_c81 bl[81] br[81] wl[107] vdd gnd cell_6t
Xbit_r108_c81 bl[81] br[81] wl[108] vdd gnd cell_6t
Xbit_r109_c81 bl[81] br[81] wl[109] vdd gnd cell_6t
Xbit_r110_c81 bl[81] br[81] wl[110] vdd gnd cell_6t
Xbit_r111_c81 bl[81] br[81] wl[111] vdd gnd cell_6t
Xbit_r112_c81 bl[81] br[81] wl[112] vdd gnd cell_6t
Xbit_r113_c81 bl[81] br[81] wl[113] vdd gnd cell_6t
Xbit_r114_c81 bl[81] br[81] wl[114] vdd gnd cell_6t
Xbit_r115_c81 bl[81] br[81] wl[115] vdd gnd cell_6t
Xbit_r116_c81 bl[81] br[81] wl[116] vdd gnd cell_6t
Xbit_r117_c81 bl[81] br[81] wl[117] vdd gnd cell_6t
Xbit_r118_c81 bl[81] br[81] wl[118] vdd gnd cell_6t
Xbit_r119_c81 bl[81] br[81] wl[119] vdd gnd cell_6t
Xbit_r120_c81 bl[81] br[81] wl[120] vdd gnd cell_6t
Xbit_r121_c81 bl[81] br[81] wl[121] vdd gnd cell_6t
Xbit_r122_c81 bl[81] br[81] wl[122] vdd gnd cell_6t
Xbit_r123_c81 bl[81] br[81] wl[123] vdd gnd cell_6t
Xbit_r124_c81 bl[81] br[81] wl[124] vdd gnd cell_6t
Xbit_r125_c81 bl[81] br[81] wl[125] vdd gnd cell_6t
Xbit_r126_c81 bl[81] br[81] wl[126] vdd gnd cell_6t
Xbit_r127_c81 bl[81] br[81] wl[127] vdd gnd cell_6t
Xbit_r128_c81 bl[81] br[81] wl[128] vdd gnd cell_6t
Xbit_r129_c81 bl[81] br[81] wl[129] vdd gnd cell_6t
Xbit_r130_c81 bl[81] br[81] wl[130] vdd gnd cell_6t
Xbit_r131_c81 bl[81] br[81] wl[131] vdd gnd cell_6t
Xbit_r132_c81 bl[81] br[81] wl[132] vdd gnd cell_6t
Xbit_r133_c81 bl[81] br[81] wl[133] vdd gnd cell_6t
Xbit_r134_c81 bl[81] br[81] wl[134] vdd gnd cell_6t
Xbit_r135_c81 bl[81] br[81] wl[135] vdd gnd cell_6t
Xbit_r136_c81 bl[81] br[81] wl[136] vdd gnd cell_6t
Xbit_r137_c81 bl[81] br[81] wl[137] vdd gnd cell_6t
Xbit_r138_c81 bl[81] br[81] wl[138] vdd gnd cell_6t
Xbit_r139_c81 bl[81] br[81] wl[139] vdd gnd cell_6t
Xbit_r140_c81 bl[81] br[81] wl[140] vdd gnd cell_6t
Xbit_r141_c81 bl[81] br[81] wl[141] vdd gnd cell_6t
Xbit_r142_c81 bl[81] br[81] wl[142] vdd gnd cell_6t
Xbit_r143_c81 bl[81] br[81] wl[143] vdd gnd cell_6t
Xbit_r144_c81 bl[81] br[81] wl[144] vdd gnd cell_6t
Xbit_r145_c81 bl[81] br[81] wl[145] vdd gnd cell_6t
Xbit_r146_c81 bl[81] br[81] wl[146] vdd gnd cell_6t
Xbit_r147_c81 bl[81] br[81] wl[147] vdd gnd cell_6t
Xbit_r148_c81 bl[81] br[81] wl[148] vdd gnd cell_6t
Xbit_r149_c81 bl[81] br[81] wl[149] vdd gnd cell_6t
Xbit_r150_c81 bl[81] br[81] wl[150] vdd gnd cell_6t
Xbit_r151_c81 bl[81] br[81] wl[151] vdd gnd cell_6t
Xbit_r152_c81 bl[81] br[81] wl[152] vdd gnd cell_6t
Xbit_r153_c81 bl[81] br[81] wl[153] vdd gnd cell_6t
Xbit_r154_c81 bl[81] br[81] wl[154] vdd gnd cell_6t
Xbit_r155_c81 bl[81] br[81] wl[155] vdd gnd cell_6t
Xbit_r156_c81 bl[81] br[81] wl[156] vdd gnd cell_6t
Xbit_r157_c81 bl[81] br[81] wl[157] vdd gnd cell_6t
Xbit_r158_c81 bl[81] br[81] wl[158] vdd gnd cell_6t
Xbit_r159_c81 bl[81] br[81] wl[159] vdd gnd cell_6t
Xbit_r160_c81 bl[81] br[81] wl[160] vdd gnd cell_6t
Xbit_r161_c81 bl[81] br[81] wl[161] vdd gnd cell_6t
Xbit_r162_c81 bl[81] br[81] wl[162] vdd gnd cell_6t
Xbit_r163_c81 bl[81] br[81] wl[163] vdd gnd cell_6t
Xbit_r164_c81 bl[81] br[81] wl[164] vdd gnd cell_6t
Xbit_r165_c81 bl[81] br[81] wl[165] vdd gnd cell_6t
Xbit_r166_c81 bl[81] br[81] wl[166] vdd gnd cell_6t
Xbit_r167_c81 bl[81] br[81] wl[167] vdd gnd cell_6t
Xbit_r168_c81 bl[81] br[81] wl[168] vdd gnd cell_6t
Xbit_r169_c81 bl[81] br[81] wl[169] vdd gnd cell_6t
Xbit_r170_c81 bl[81] br[81] wl[170] vdd gnd cell_6t
Xbit_r171_c81 bl[81] br[81] wl[171] vdd gnd cell_6t
Xbit_r172_c81 bl[81] br[81] wl[172] vdd gnd cell_6t
Xbit_r173_c81 bl[81] br[81] wl[173] vdd gnd cell_6t
Xbit_r174_c81 bl[81] br[81] wl[174] vdd gnd cell_6t
Xbit_r175_c81 bl[81] br[81] wl[175] vdd gnd cell_6t
Xbit_r176_c81 bl[81] br[81] wl[176] vdd gnd cell_6t
Xbit_r177_c81 bl[81] br[81] wl[177] vdd gnd cell_6t
Xbit_r178_c81 bl[81] br[81] wl[178] vdd gnd cell_6t
Xbit_r179_c81 bl[81] br[81] wl[179] vdd gnd cell_6t
Xbit_r180_c81 bl[81] br[81] wl[180] vdd gnd cell_6t
Xbit_r181_c81 bl[81] br[81] wl[181] vdd gnd cell_6t
Xbit_r182_c81 bl[81] br[81] wl[182] vdd gnd cell_6t
Xbit_r183_c81 bl[81] br[81] wl[183] vdd gnd cell_6t
Xbit_r184_c81 bl[81] br[81] wl[184] vdd gnd cell_6t
Xbit_r185_c81 bl[81] br[81] wl[185] vdd gnd cell_6t
Xbit_r186_c81 bl[81] br[81] wl[186] vdd gnd cell_6t
Xbit_r187_c81 bl[81] br[81] wl[187] vdd gnd cell_6t
Xbit_r188_c81 bl[81] br[81] wl[188] vdd gnd cell_6t
Xbit_r189_c81 bl[81] br[81] wl[189] vdd gnd cell_6t
Xbit_r190_c81 bl[81] br[81] wl[190] vdd gnd cell_6t
Xbit_r191_c81 bl[81] br[81] wl[191] vdd gnd cell_6t
Xbit_r192_c81 bl[81] br[81] wl[192] vdd gnd cell_6t
Xbit_r193_c81 bl[81] br[81] wl[193] vdd gnd cell_6t
Xbit_r194_c81 bl[81] br[81] wl[194] vdd gnd cell_6t
Xbit_r195_c81 bl[81] br[81] wl[195] vdd gnd cell_6t
Xbit_r196_c81 bl[81] br[81] wl[196] vdd gnd cell_6t
Xbit_r197_c81 bl[81] br[81] wl[197] vdd gnd cell_6t
Xbit_r198_c81 bl[81] br[81] wl[198] vdd gnd cell_6t
Xbit_r199_c81 bl[81] br[81] wl[199] vdd gnd cell_6t
Xbit_r200_c81 bl[81] br[81] wl[200] vdd gnd cell_6t
Xbit_r201_c81 bl[81] br[81] wl[201] vdd gnd cell_6t
Xbit_r202_c81 bl[81] br[81] wl[202] vdd gnd cell_6t
Xbit_r203_c81 bl[81] br[81] wl[203] vdd gnd cell_6t
Xbit_r204_c81 bl[81] br[81] wl[204] vdd gnd cell_6t
Xbit_r205_c81 bl[81] br[81] wl[205] vdd gnd cell_6t
Xbit_r206_c81 bl[81] br[81] wl[206] vdd gnd cell_6t
Xbit_r207_c81 bl[81] br[81] wl[207] vdd gnd cell_6t
Xbit_r208_c81 bl[81] br[81] wl[208] vdd gnd cell_6t
Xbit_r209_c81 bl[81] br[81] wl[209] vdd gnd cell_6t
Xbit_r210_c81 bl[81] br[81] wl[210] vdd gnd cell_6t
Xbit_r211_c81 bl[81] br[81] wl[211] vdd gnd cell_6t
Xbit_r212_c81 bl[81] br[81] wl[212] vdd gnd cell_6t
Xbit_r213_c81 bl[81] br[81] wl[213] vdd gnd cell_6t
Xbit_r214_c81 bl[81] br[81] wl[214] vdd gnd cell_6t
Xbit_r215_c81 bl[81] br[81] wl[215] vdd gnd cell_6t
Xbit_r216_c81 bl[81] br[81] wl[216] vdd gnd cell_6t
Xbit_r217_c81 bl[81] br[81] wl[217] vdd gnd cell_6t
Xbit_r218_c81 bl[81] br[81] wl[218] vdd gnd cell_6t
Xbit_r219_c81 bl[81] br[81] wl[219] vdd gnd cell_6t
Xbit_r220_c81 bl[81] br[81] wl[220] vdd gnd cell_6t
Xbit_r221_c81 bl[81] br[81] wl[221] vdd gnd cell_6t
Xbit_r222_c81 bl[81] br[81] wl[222] vdd gnd cell_6t
Xbit_r223_c81 bl[81] br[81] wl[223] vdd gnd cell_6t
Xbit_r224_c81 bl[81] br[81] wl[224] vdd gnd cell_6t
Xbit_r225_c81 bl[81] br[81] wl[225] vdd gnd cell_6t
Xbit_r226_c81 bl[81] br[81] wl[226] vdd gnd cell_6t
Xbit_r227_c81 bl[81] br[81] wl[227] vdd gnd cell_6t
Xbit_r228_c81 bl[81] br[81] wl[228] vdd gnd cell_6t
Xbit_r229_c81 bl[81] br[81] wl[229] vdd gnd cell_6t
Xbit_r230_c81 bl[81] br[81] wl[230] vdd gnd cell_6t
Xbit_r231_c81 bl[81] br[81] wl[231] vdd gnd cell_6t
Xbit_r232_c81 bl[81] br[81] wl[232] vdd gnd cell_6t
Xbit_r233_c81 bl[81] br[81] wl[233] vdd gnd cell_6t
Xbit_r234_c81 bl[81] br[81] wl[234] vdd gnd cell_6t
Xbit_r235_c81 bl[81] br[81] wl[235] vdd gnd cell_6t
Xbit_r236_c81 bl[81] br[81] wl[236] vdd gnd cell_6t
Xbit_r237_c81 bl[81] br[81] wl[237] vdd gnd cell_6t
Xbit_r238_c81 bl[81] br[81] wl[238] vdd gnd cell_6t
Xbit_r239_c81 bl[81] br[81] wl[239] vdd gnd cell_6t
Xbit_r240_c81 bl[81] br[81] wl[240] vdd gnd cell_6t
Xbit_r241_c81 bl[81] br[81] wl[241] vdd gnd cell_6t
Xbit_r242_c81 bl[81] br[81] wl[242] vdd gnd cell_6t
Xbit_r243_c81 bl[81] br[81] wl[243] vdd gnd cell_6t
Xbit_r244_c81 bl[81] br[81] wl[244] vdd gnd cell_6t
Xbit_r245_c81 bl[81] br[81] wl[245] vdd gnd cell_6t
Xbit_r246_c81 bl[81] br[81] wl[246] vdd gnd cell_6t
Xbit_r247_c81 bl[81] br[81] wl[247] vdd gnd cell_6t
Xbit_r248_c81 bl[81] br[81] wl[248] vdd gnd cell_6t
Xbit_r249_c81 bl[81] br[81] wl[249] vdd gnd cell_6t
Xbit_r250_c81 bl[81] br[81] wl[250] vdd gnd cell_6t
Xbit_r251_c81 bl[81] br[81] wl[251] vdd gnd cell_6t
Xbit_r252_c81 bl[81] br[81] wl[252] vdd gnd cell_6t
Xbit_r253_c81 bl[81] br[81] wl[253] vdd gnd cell_6t
Xbit_r254_c81 bl[81] br[81] wl[254] vdd gnd cell_6t
Xbit_r255_c81 bl[81] br[81] wl[255] vdd gnd cell_6t
Xbit_r256_c81 bl[81] br[81] wl[256] vdd gnd cell_6t
Xbit_r257_c81 bl[81] br[81] wl[257] vdd gnd cell_6t
Xbit_r258_c81 bl[81] br[81] wl[258] vdd gnd cell_6t
Xbit_r259_c81 bl[81] br[81] wl[259] vdd gnd cell_6t
Xbit_r260_c81 bl[81] br[81] wl[260] vdd gnd cell_6t
Xbit_r261_c81 bl[81] br[81] wl[261] vdd gnd cell_6t
Xbit_r262_c81 bl[81] br[81] wl[262] vdd gnd cell_6t
Xbit_r263_c81 bl[81] br[81] wl[263] vdd gnd cell_6t
Xbit_r264_c81 bl[81] br[81] wl[264] vdd gnd cell_6t
Xbit_r265_c81 bl[81] br[81] wl[265] vdd gnd cell_6t
Xbit_r266_c81 bl[81] br[81] wl[266] vdd gnd cell_6t
Xbit_r267_c81 bl[81] br[81] wl[267] vdd gnd cell_6t
Xbit_r268_c81 bl[81] br[81] wl[268] vdd gnd cell_6t
Xbit_r269_c81 bl[81] br[81] wl[269] vdd gnd cell_6t
Xbit_r270_c81 bl[81] br[81] wl[270] vdd gnd cell_6t
Xbit_r271_c81 bl[81] br[81] wl[271] vdd gnd cell_6t
Xbit_r272_c81 bl[81] br[81] wl[272] vdd gnd cell_6t
Xbit_r273_c81 bl[81] br[81] wl[273] vdd gnd cell_6t
Xbit_r274_c81 bl[81] br[81] wl[274] vdd gnd cell_6t
Xbit_r275_c81 bl[81] br[81] wl[275] vdd gnd cell_6t
Xbit_r276_c81 bl[81] br[81] wl[276] vdd gnd cell_6t
Xbit_r277_c81 bl[81] br[81] wl[277] vdd gnd cell_6t
Xbit_r278_c81 bl[81] br[81] wl[278] vdd gnd cell_6t
Xbit_r279_c81 bl[81] br[81] wl[279] vdd gnd cell_6t
Xbit_r280_c81 bl[81] br[81] wl[280] vdd gnd cell_6t
Xbit_r281_c81 bl[81] br[81] wl[281] vdd gnd cell_6t
Xbit_r282_c81 bl[81] br[81] wl[282] vdd gnd cell_6t
Xbit_r283_c81 bl[81] br[81] wl[283] vdd gnd cell_6t
Xbit_r284_c81 bl[81] br[81] wl[284] vdd gnd cell_6t
Xbit_r285_c81 bl[81] br[81] wl[285] vdd gnd cell_6t
Xbit_r286_c81 bl[81] br[81] wl[286] vdd gnd cell_6t
Xbit_r287_c81 bl[81] br[81] wl[287] vdd gnd cell_6t
Xbit_r288_c81 bl[81] br[81] wl[288] vdd gnd cell_6t
Xbit_r289_c81 bl[81] br[81] wl[289] vdd gnd cell_6t
Xbit_r290_c81 bl[81] br[81] wl[290] vdd gnd cell_6t
Xbit_r291_c81 bl[81] br[81] wl[291] vdd gnd cell_6t
Xbit_r292_c81 bl[81] br[81] wl[292] vdd gnd cell_6t
Xbit_r293_c81 bl[81] br[81] wl[293] vdd gnd cell_6t
Xbit_r294_c81 bl[81] br[81] wl[294] vdd gnd cell_6t
Xbit_r295_c81 bl[81] br[81] wl[295] vdd gnd cell_6t
Xbit_r296_c81 bl[81] br[81] wl[296] vdd gnd cell_6t
Xbit_r297_c81 bl[81] br[81] wl[297] vdd gnd cell_6t
Xbit_r298_c81 bl[81] br[81] wl[298] vdd gnd cell_6t
Xbit_r299_c81 bl[81] br[81] wl[299] vdd gnd cell_6t
Xbit_r300_c81 bl[81] br[81] wl[300] vdd gnd cell_6t
Xbit_r301_c81 bl[81] br[81] wl[301] vdd gnd cell_6t
Xbit_r302_c81 bl[81] br[81] wl[302] vdd gnd cell_6t
Xbit_r303_c81 bl[81] br[81] wl[303] vdd gnd cell_6t
Xbit_r304_c81 bl[81] br[81] wl[304] vdd gnd cell_6t
Xbit_r305_c81 bl[81] br[81] wl[305] vdd gnd cell_6t
Xbit_r306_c81 bl[81] br[81] wl[306] vdd gnd cell_6t
Xbit_r307_c81 bl[81] br[81] wl[307] vdd gnd cell_6t
Xbit_r308_c81 bl[81] br[81] wl[308] vdd gnd cell_6t
Xbit_r309_c81 bl[81] br[81] wl[309] vdd gnd cell_6t
Xbit_r310_c81 bl[81] br[81] wl[310] vdd gnd cell_6t
Xbit_r311_c81 bl[81] br[81] wl[311] vdd gnd cell_6t
Xbit_r312_c81 bl[81] br[81] wl[312] vdd gnd cell_6t
Xbit_r313_c81 bl[81] br[81] wl[313] vdd gnd cell_6t
Xbit_r314_c81 bl[81] br[81] wl[314] vdd gnd cell_6t
Xbit_r315_c81 bl[81] br[81] wl[315] vdd gnd cell_6t
Xbit_r316_c81 bl[81] br[81] wl[316] vdd gnd cell_6t
Xbit_r317_c81 bl[81] br[81] wl[317] vdd gnd cell_6t
Xbit_r318_c81 bl[81] br[81] wl[318] vdd gnd cell_6t
Xbit_r319_c81 bl[81] br[81] wl[319] vdd gnd cell_6t
Xbit_r320_c81 bl[81] br[81] wl[320] vdd gnd cell_6t
Xbit_r321_c81 bl[81] br[81] wl[321] vdd gnd cell_6t
Xbit_r322_c81 bl[81] br[81] wl[322] vdd gnd cell_6t
Xbit_r323_c81 bl[81] br[81] wl[323] vdd gnd cell_6t
Xbit_r324_c81 bl[81] br[81] wl[324] vdd gnd cell_6t
Xbit_r325_c81 bl[81] br[81] wl[325] vdd gnd cell_6t
Xbit_r326_c81 bl[81] br[81] wl[326] vdd gnd cell_6t
Xbit_r327_c81 bl[81] br[81] wl[327] vdd gnd cell_6t
Xbit_r328_c81 bl[81] br[81] wl[328] vdd gnd cell_6t
Xbit_r329_c81 bl[81] br[81] wl[329] vdd gnd cell_6t
Xbit_r330_c81 bl[81] br[81] wl[330] vdd gnd cell_6t
Xbit_r331_c81 bl[81] br[81] wl[331] vdd gnd cell_6t
Xbit_r332_c81 bl[81] br[81] wl[332] vdd gnd cell_6t
Xbit_r333_c81 bl[81] br[81] wl[333] vdd gnd cell_6t
Xbit_r334_c81 bl[81] br[81] wl[334] vdd gnd cell_6t
Xbit_r335_c81 bl[81] br[81] wl[335] vdd gnd cell_6t
Xbit_r336_c81 bl[81] br[81] wl[336] vdd gnd cell_6t
Xbit_r337_c81 bl[81] br[81] wl[337] vdd gnd cell_6t
Xbit_r338_c81 bl[81] br[81] wl[338] vdd gnd cell_6t
Xbit_r339_c81 bl[81] br[81] wl[339] vdd gnd cell_6t
Xbit_r340_c81 bl[81] br[81] wl[340] vdd gnd cell_6t
Xbit_r341_c81 bl[81] br[81] wl[341] vdd gnd cell_6t
Xbit_r342_c81 bl[81] br[81] wl[342] vdd gnd cell_6t
Xbit_r343_c81 bl[81] br[81] wl[343] vdd gnd cell_6t
Xbit_r344_c81 bl[81] br[81] wl[344] vdd gnd cell_6t
Xbit_r345_c81 bl[81] br[81] wl[345] vdd gnd cell_6t
Xbit_r346_c81 bl[81] br[81] wl[346] vdd gnd cell_6t
Xbit_r347_c81 bl[81] br[81] wl[347] vdd gnd cell_6t
Xbit_r348_c81 bl[81] br[81] wl[348] vdd gnd cell_6t
Xbit_r349_c81 bl[81] br[81] wl[349] vdd gnd cell_6t
Xbit_r350_c81 bl[81] br[81] wl[350] vdd gnd cell_6t
Xbit_r351_c81 bl[81] br[81] wl[351] vdd gnd cell_6t
Xbit_r352_c81 bl[81] br[81] wl[352] vdd gnd cell_6t
Xbit_r353_c81 bl[81] br[81] wl[353] vdd gnd cell_6t
Xbit_r354_c81 bl[81] br[81] wl[354] vdd gnd cell_6t
Xbit_r355_c81 bl[81] br[81] wl[355] vdd gnd cell_6t
Xbit_r356_c81 bl[81] br[81] wl[356] vdd gnd cell_6t
Xbit_r357_c81 bl[81] br[81] wl[357] vdd gnd cell_6t
Xbit_r358_c81 bl[81] br[81] wl[358] vdd gnd cell_6t
Xbit_r359_c81 bl[81] br[81] wl[359] vdd gnd cell_6t
Xbit_r360_c81 bl[81] br[81] wl[360] vdd gnd cell_6t
Xbit_r361_c81 bl[81] br[81] wl[361] vdd gnd cell_6t
Xbit_r362_c81 bl[81] br[81] wl[362] vdd gnd cell_6t
Xbit_r363_c81 bl[81] br[81] wl[363] vdd gnd cell_6t
Xbit_r364_c81 bl[81] br[81] wl[364] vdd gnd cell_6t
Xbit_r365_c81 bl[81] br[81] wl[365] vdd gnd cell_6t
Xbit_r366_c81 bl[81] br[81] wl[366] vdd gnd cell_6t
Xbit_r367_c81 bl[81] br[81] wl[367] vdd gnd cell_6t
Xbit_r368_c81 bl[81] br[81] wl[368] vdd gnd cell_6t
Xbit_r369_c81 bl[81] br[81] wl[369] vdd gnd cell_6t
Xbit_r370_c81 bl[81] br[81] wl[370] vdd gnd cell_6t
Xbit_r371_c81 bl[81] br[81] wl[371] vdd gnd cell_6t
Xbit_r372_c81 bl[81] br[81] wl[372] vdd gnd cell_6t
Xbit_r373_c81 bl[81] br[81] wl[373] vdd gnd cell_6t
Xbit_r374_c81 bl[81] br[81] wl[374] vdd gnd cell_6t
Xbit_r375_c81 bl[81] br[81] wl[375] vdd gnd cell_6t
Xbit_r376_c81 bl[81] br[81] wl[376] vdd gnd cell_6t
Xbit_r377_c81 bl[81] br[81] wl[377] vdd gnd cell_6t
Xbit_r378_c81 bl[81] br[81] wl[378] vdd gnd cell_6t
Xbit_r379_c81 bl[81] br[81] wl[379] vdd gnd cell_6t
Xbit_r380_c81 bl[81] br[81] wl[380] vdd gnd cell_6t
Xbit_r381_c81 bl[81] br[81] wl[381] vdd gnd cell_6t
Xbit_r382_c81 bl[81] br[81] wl[382] vdd gnd cell_6t
Xbit_r383_c81 bl[81] br[81] wl[383] vdd gnd cell_6t
Xbit_r384_c81 bl[81] br[81] wl[384] vdd gnd cell_6t
Xbit_r385_c81 bl[81] br[81] wl[385] vdd gnd cell_6t
Xbit_r386_c81 bl[81] br[81] wl[386] vdd gnd cell_6t
Xbit_r387_c81 bl[81] br[81] wl[387] vdd gnd cell_6t
Xbit_r388_c81 bl[81] br[81] wl[388] vdd gnd cell_6t
Xbit_r389_c81 bl[81] br[81] wl[389] vdd gnd cell_6t
Xbit_r390_c81 bl[81] br[81] wl[390] vdd gnd cell_6t
Xbit_r391_c81 bl[81] br[81] wl[391] vdd gnd cell_6t
Xbit_r392_c81 bl[81] br[81] wl[392] vdd gnd cell_6t
Xbit_r393_c81 bl[81] br[81] wl[393] vdd gnd cell_6t
Xbit_r394_c81 bl[81] br[81] wl[394] vdd gnd cell_6t
Xbit_r395_c81 bl[81] br[81] wl[395] vdd gnd cell_6t
Xbit_r396_c81 bl[81] br[81] wl[396] vdd gnd cell_6t
Xbit_r397_c81 bl[81] br[81] wl[397] vdd gnd cell_6t
Xbit_r398_c81 bl[81] br[81] wl[398] vdd gnd cell_6t
Xbit_r399_c81 bl[81] br[81] wl[399] vdd gnd cell_6t
Xbit_r400_c81 bl[81] br[81] wl[400] vdd gnd cell_6t
Xbit_r401_c81 bl[81] br[81] wl[401] vdd gnd cell_6t
Xbit_r402_c81 bl[81] br[81] wl[402] vdd gnd cell_6t
Xbit_r403_c81 bl[81] br[81] wl[403] vdd gnd cell_6t
Xbit_r404_c81 bl[81] br[81] wl[404] vdd gnd cell_6t
Xbit_r405_c81 bl[81] br[81] wl[405] vdd gnd cell_6t
Xbit_r406_c81 bl[81] br[81] wl[406] vdd gnd cell_6t
Xbit_r407_c81 bl[81] br[81] wl[407] vdd gnd cell_6t
Xbit_r408_c81 bl[81] br[81] wl[408] vdd gnd cell_6t
Xbit_r409_c81 bl[81] br[81] wl[409] vdd gnd cell_6t
Xbit_r410_c81 bl[81] br[81] wl[410] vdd gnd cell_6t
Xbit_r411_c81 bl[81] br[81] wl[411] vdd gnd cell_6t
Xbit_r412_c81 bl[81] br[81] wl[412] vdd gnd cell_6t
Xbit_r413_c81 bl[81] br[81] wl[413] vdd gnd cell_6t
Xbit_r414_c81 bl[81] br[81] wl[414] vdd gnd cell_6t
Xbit_r415_c81 bl[81] br[81] wl[415] vdd gnd cell_6t
Xbit_r416_c81 bl[81] br[81] wl[416] vdd gnd cell_6t
Xbit_r417_c81 bl[81] br[81] wl[417] vdd gnd cell_6t
Xbit_r418_c81 bl[81] br[81] wl[418] vdd gnd cell_6t
Xbit_r419_c81 bl[81] br[81] wl[419] vdd gnd cell_6t
Xbit_r420_c81 bl[81] br[81] wl[420] vdd gnd cell_6t
Xbit_r421_c81 bl[81] br[81] wl[421] vdd gnd cell_6t
Xbit_r422_c81 bl[81] br[81] wl[422] vdd gnd cell_6t
Xbit_r423_c81 bl[81] br[81] wl[423] vdd gnd cell_6t
Xbit_r424_c81 bl[81] br[81] wl[424] vdd gnd cell_6t
Xbit_r425_c81 bl[81] br[81] wl[425] vdd gnd cell_6t
Xbit_r426_c81 bl[81] br[81] wl[426] vdd gnd cell_6t
Xbit_r427_c81 bl[81] br[81] wl[427] vdd gnd cell_6t
Xbit_r428_c81 bl[81] br[81] wl[428] vdd gnd cell_6t
Xbit_r429_c81 bl[81] br[81] wl[429] vdd gnd cell_6t
Xbit_r430_c81 bl[81] br[81] wl[430] vdd gnd cell_6t
Xbit_r431_c81 bl[81] br[81] wl[431] vdd gnd cell_6t
Xbit_r432_c81 bl[81] br[81] wl[432] vdd gnd cell_6t
Xbit_r433_c81 bl[81] br[81] wl[433] vdd gnd cell_6t
Xbit_r434_c81 bl[81] br[81] wl[434] vdd gnd cell_6t
Xbit_r435_c81 bl[81] br[81] wl[435] vdd gnd cell_6t
Xbit_r436_c81 bl[81] br[81] wl[436] vdd gnd cell_6t
Xbit_r437_c81 bl[81] br[81] wl[437] vdd gnd cell_6t
Xbit_r438_c81 bl[81] br[81] wl[438] vdd gnd cell_6t
Xbit_r439_c81 bl[81] br[81] wl[439] vdd gnd cell_6t
Xbit_r440_c81 bl[81] br[81] wl[440] vdd gnd cell_6t
Xbit_r441_c81 bl[81] br[81] wl[441] vdd gnd cell_6t
Xbit_r442_c81 bl[81] br[81] wl[442] vdd gnd cell_6t
Xbit_r443_c81 bl[81] br[81] wl[443] vdd gnd cell_6t
Xbit_r444_c81 bl[81] br[81] wl[444] vdd gnd cell_6t
Xbit_r445_c81 bl[81] br[81] wl[445] vdd gnd cell_6t
Xbit_r446_c81 bl[81] br[81] wl[446] vdd gnd cell_6t
Xbit_r447_c81 bl[81] br[81] wl[447] vdd gnd cell_6t
Xbit_r448_c81 bl[81] br[81] wl[448] vdd gnd cell_6t
Xbit_r449_c81 bl[81] br[81] wl[449] vdd gnd cell_6t
Xbit_r450_c81 bl[81] br[81] wl[450] vdd gnd cell_6t
Xbit_r451_c81 bl[81] br[81] wl[451] vdd gnd cell_6t
Xbit_r452_c81 bl[81] br[81] wl[452] vdd gnd cell_6t
Xbit_r453_c81 bl[81] br[81] wl[453] vdd gnd cell_6t
Xbit_r454_c81 bl[81] br[81] wl[454] vdd gnd cell_6t
Xbit_r455_c81 bl[81] br[81] wl[455] vdd gnd cell_6t
Xbit_r456_c81 bl[81] br[81] wl[456] vdd gnd cell_6t
Xbit_r457_c81 bl[81] br[81] wl[457] vdd gnd cell_6t
Xbit_r458_c81 bl[81] br[81] wl[458] vdd gnd cell_6t
Xbit_r459_c81 bl[81] br[81] wl[459] vdd gnd cell_6t
Xbit_r460_c81 bl[81] br[81] wl[460] vdd gnd cell_6t
Xbit_r461_c81 bl[81] br[81] wl[461] vdd gnd cell_6t
Xbit_r462_c81 bl[81] br[81] wl[462] vdd gnd cell_6t
Xbit_r463_c81 bl[81] br[81] wl[463] vdd gnd cell_6t
Xbit_r464_c81 bl[81] br[81] wl[464] vdd gnd cell_6t
Xbit_r465_c81 bl[81] br[81] wl[465] vdd gnd cell_6t
Xbit_r466_c81 bl[81] br[81] wl[466] vdd gnd cell_6t
Xbit_r467_c81 bl[81] br[81] wl[467] vdd gnd cell_6t
Xbit_r468_c81 bl[81] br[81] wl[468] vdd gnd cell_6t
Xbit_r469_c81 bl[81] br[81] wl[469] vdd gnd cell_6t
Xbit_r470_c81 bl[81] br[81] wl[470] vdd gnd cell_6t
Xbit_r471_c81 bl[81] br[81] wl[471] vdd gnd cell_6t
Xbit_r472_c81 bl[81] br[81] wl[472] vdd gnd cell_6t
Xbit_r473_c81 bl[81] br[81] wl[473] vdd gnd cell_6t
Xbit_r474_c81 bl[81] br[81] wl[474] vdd gnd cell_6t
Xbit_r475_c81 bl[81] br[81] wl[475] vdd gnd cell_6t
Xbit_r476_c81 bl[81] br[81] wl[476] vdd gnd cell_6t
Xbit_r477_c81 bl[81] br[81] wl[477] vdd gnd cell_6t
Xbit_r478_c81 bl[81] br[81] wl[478] vdd gnd cell_6t
Xbit_r479_c81 bl[81] br[81] wl[479] vdd gnd cell_6t
Xbit_r480_c81 bl[81] br[81] wl[480] vdd gnd cell_6t
Xbit_r481_c81 bl[81] br[81] wl[481] vdd gnd cell_6t
Xbit_r482_c81 bl[81] br[81] wl[482] vdd gnd cell_6t
Xbit_r483_c81 bl[81] br[81] wl[483] vdd gnd cell_6t
Xbit_r484_c81 bl[81] br[81] wl[484] vdd gnd cell_6t
Xbit_r485_c81 bl[81] br[81] wl[485] vdd gnd cell_6t
Xbit_r486_c81 bl[81] br[81] wl[486] vdd gnd cell_6t
Xbit_r487_c81 bl[81] br[81] wl[487] vdd gnd cell_6t
Xbit_r488_c81 bl[81] br[81] wl[488] vdd gnd cell_6t
Xbit_r489_c81 bl[81] br[81] wl[489] vdd gnd cell_6t
Xbit_r490_c81 bl[81] br[81] wl[490] vdd gnd cell_6t
Xbit_r491_c81 bl[81] br[81] wl[491] vdd gnd cell_6t
Xbit_r492_c81 bl[81] br[81] wl[492] vdd gnd cell_6t
Xbit_r493_c81 bl[81] br[81] wl[493] vdd gnd cell_6t
Xbit_r494_c81 bl[81] br[81] wl[494] vdd gnd cell_6t
Xbit_r495_c81 bl[81] br[81] wl[495] vdd gnd cell_6t
Xbit_r496_c81 bl[81] br[81] wl[496] vdd gnd cell_6t
Xbit_r497_c81 bl[81] br[81] wl[497] vdd gnd cell_6t
Xbit_r498_c81 bl[81] br[81] wl[498] vdd gnd cell_6t
Xbit_r499_c81 bl[81] br[81] wl[499] vdd gnd cell_6t
Xbit_r500_c81 bl[81] br[81] wl[500] vdd gnd cell_6t
Xbit_r501_c81 bl[81] br[81] wl[501] vdd gnd cell_6t
Xbit_r502_c81 bl[81] br[81] wl[502] vdd gnd cell_6t
Xbit_r503_c81 bl[81] br[81] wl[503] vdd gnd cell_6t
Xbit_r504_c81 bl[81] br[81] wl[504] vdd gnd cell_6t
Xbit_r505_c81 bl[81] br[81] wl[505] vdd gnd cell_6t
Xbit_r506_c81 bl[81] br[81] wl[506] vdd gnd cell_6t
Xbit_r507_c81 bl[81] br[81] wl[507] vdd gnd cell_6t
Xbit_r508_c81 bl[81] br[81] wl[508] vdd gnd cell_6t
Xbit_r509_c81 bl[81] br[81] wl[509] vdd gnd cell_6t
Xbit_r510_c81 bl[81] br[81] wl[510] vdd gnd cell_6t
Xbit_r511_c81 bl[81] br[81] wl[511] vdd gnd cell_6t
Xbit_r0_c82 bl[82] br[82] wl[0] vdd gnd cell_6t
Xbit_r1_c82 bl[82] br[82] wl[1] vdd gnd cell_6t
Xbit_r2_c82 bl[82] br[82] wl[2] vdd gnd cell_6t
Xbit_r3_c82 bl[82] br[82] wl[3] vdd gnd cell_6t
Xbit_r4_c82 bl[82] br[82] wl[4] vdd gnd cell_6t
Xbit_r5_c82 bl[82] br[82] wl[5] vdd gnd cell_6t
Xbit_r6_c82 bl[82] br[82] wl[6] vdd gnd cell_6t
Xbit_r7_c82 bl[82] br[82] wl[7] vdd gnd cell_6t
Xbit_r8_c82 bl[82] br[82] wl[8] vdd gnd cell_6t
Xbit_r9_c82 bl[82] br[82] wl[9] vdd gnd cell_6t
Xbit_r10_c82 bl[82] br[82] wl[10] vdd gnd cell_6t
Xbit_r11_c82 bl[82] br[82] wl[11] vdd gnd cell_6t
Xbit_r12_c82 bl[82] br[82] wl[12] vdd gnd cell_6t
Xbit_r13_c82 bl[82] br[82] wl[13] vdd gnd cell_6t
Xbit_r14_c82 bl[82] br[82] wl[14] vdd gnd cell_6t
Xbit_r15_c82 bl[82] br[82] wl[15] vdd gnd cell_6t
Xbit_r16_c82 bl[82] br[82] wl[16] vdd gnd cell_6t
Xbit_r17_c82 bl[82] br[82] wl[17] vdd gnd cell_6t
Xbit_r18_c82 bl[82] br[82] wl[18] vdd gnd cell_6t
Xbit_r19_c82 bl[82] br[82] wl[19] vdd gnd cell_6t
Xbit_r20_c82 bl[82] br[82] wl[20] vdd gnd cell_6t
Xbit_r21_c82 bl[82] br[82] wl[21] vdd gnd cell_6t
Xbit_r22_c82 bl[82] br[82] wl[22] vdd gnd cell_6t
Xbit_r23_c82 bl[82] br[82] wl[23] vdd gnd cell_6t
Xbit_r24_c82 bl[82] br[82] wl[24] vdd gnd cell_6t
Xbit_r25_c82 bl[82] br[82] wl[25] vdd gnd cell_6t
Xbit_r26_c82 bl[82] br[82] wl[26] vdd gnd cell_6t
Xbit_r27_c82 bl[82] br[82] wl[27] vdd gnd cell_6t
Xbit_r28_c82 bl[82] br[82] wl[28] vdd gnd cell_6t
Xbit_r29_c82 bl[82] br[82] wl[29] vdd gnd cell_6t
Xbit_r30_c82 bl[82] br[82] wl[30] vdd gnd cell_6t
Xbit_r31_c82 bl[82] br[82] wl[31] vdd gnd cell_6t
Xbit_r32_c82 bl[82] br[82] wl[32] vdd gnd cell_6t
Xbit_r33_c82 bl[82] br[82] wl[33] vdd gnd cell_6t
Xbit_r34_c82 bl[82] br[82] wl[34] vdd gnd cell_6t
Xbit_r35_c82 bl[82] br[82] wl[35] vdd gnd cell_6t
Xbit_r36_c82 bl[82] br[82] wl[36] vdd gnd cell_6t
Xbit_r37_c82 bl[82] br[82] wl[37] vdd gnd cell_6t
Xbit_r38_c82 bl[82] br[82] wl[38] vdd gnd cell_6t
Xbit_r39_c82 bl[82] br[82] wl[39] vdd gnd cell_6t
Xbit_r40_c82 bl[82] br[82] wl[40] vdd gnd cell_6t
Xbit_r41_c82 bl[82] br[82] wl[41] vdd gnd cell_6t
Xbit_r42_c82 bl[82] br[82] wl[42] vdd gnd cell_6t
Xbit_r43_c82 bl[82] br[82] wl[43] vdd gnd cell_6t
Xbit_r44_c82 bl[82] br[82] wl[44] vdd gnd cell_6t
Xbit_r45_c82 bl[82] br[82] wl[45] vdd gnd cell_6t
Xbit_r46_c82 bl[82] br[82] wl[46] vdd gnd cell_6t
Xbit_r47_c82 bl[82] br[82] wl[47] vdd gnd cell_6t
Xbit_r48_c82 bl[82] br[82] wl[48] vdd gnd cell_6t
Xbit_r49_c82 bl[82] br[82] wl[49] vdd gnd cell_6t
Xbit_r50_c82 bl[82] br[82] wl[50] vdd gnd cell_6t
Xbit_r51_c82 bl[82] br[82] wl[51] vdd gnd cell_6t
Xbit_r52_c82 bl[82] br[82] wl[52] vdd gnd cell_6t
Xbit_r53_c82 bl[82] br[82] wl[53] vdd gnd cell_6t
Xbit_r54_c82 bl[82] br[82] wl[54] vdd gnd cell_6t
Xbit_r55_c82 bl[82] br[82] wl[55] vdd gnd cell_6t
Xbit_r56_c82 bl[82] br[82] wl[56] vdd gnd cell_6t
Xbit_r57_c82 bl[82] br[82] wl[57] vdd gnd cell_6t
Xbit_r58_c82 bl[82] br[82] wl[58] vdd gnd cell_6t
Xbit_r59_c82 bl[82] br[82] wl[59] vdd gnd cell_6t
Xbit_r60_c82 bl[82] br[82] wl[60] vdd gnd cell_6t
Xbit_r61_c82 bl[82] br[82] wl[61] vdd gnd cell_6t
Xbit_r62_c82 bl[82] br[82] wl[62] vdd gnd cell_6t
Xbit_r63_c82 bl[82] br[82] wl[63] vdd gnd cell_6t
Xbit_r64_c82 bl[82] br[82] wl[64] vdd gnd cell_6t
Xbit_r65_c82 bl[82] br[82] wl[65] vdd gnd cell_6t
Xbit_r66_c82 bl[82] br[82] wl[66] vdd gnd cell_6t
Xbit_r67_c82 bl[82] br[82] wl[67] vdd gnd cell_6t
Xbit_r68_c82 bl[82] br[82] wl[68] vdd gnd cell_6t
Xbit_r69_c82 bl[82] br[82] wl[69] vdd gnd cell_6t
Xbit_r70_c82 bl[82] br[82] wl[70] vdd gnd cell_6t
Xbit_r71_c82 bl[82] br[82] wl[71] vdd gnd cell_6t
Xbit_r72_c82 bl[82] br[82] wl[72] vdd gnd cell_6t
Xbit_r73_c82 bl[82] br[82] wl[73] vdd gnd cell_6t
Xbit_r74_c82 bl[82] br[82] wl[74] vdd gnd cell_6t
Xbit_r75_c82 bl[82] br[82] wl[75] vdd gnd cell_6t
Xbit_r76_c82 bl[82] br[82] wl[76] vdd gnd cell_6t
Xbit_r77_c82 bl[82] br[82] wl[77] vdd gnd cell_6t
Xbit_r78_c82 bl[82] br[82] wl[78] vdd gnd cell_6t
Xbit_r79_c82 bl[82] br[82] wl[79] vdd gnd cell_6t
Xbit_r80_c82 bl[82] br[82] wl[80] vdd gnd cell_6t
Xbit_r81_c82 bl[82] br[82] wl[81] vdd gnd cell_6t
Xbit_r82_c82 bl[82] br[82] wl[82] vdd gnd cell_6t
Xbit_r83_c82 bl[82] br[82] wl[83] vdd gnd cell_6t
Xbit_r84_c82 bl[82] br[82] wl[84] vdd gnd cell_6t
Xbit_r85_c82 bl[82] br[82] wl[85] vdd gnd cell_6t
Xbit_r86_c82 bl[82] br[82] wl[86] vdd gnd cell_6t
Xbit_r87_c82 bl[82] br[82] wl[87] vdd gnd cell_6t
Xbit_r88_c82 bl[82] br[82] wl[88] vdd gnd cell_6t
Xbit_r89_c82 bl[82] br[82] wl[89] vdd gnd cell_6t
Xbit_r90_c82 bl[82] br[82] wl[90] vdd gnd cell_6t
Xbit_r91_c82 bl[82] br[82] wl[91] vdd gnd cell_6t
Xbit_r92_c82 bl[82] br[82] wl[92] vdd gnd cell_6t
Xbit_r93_c82 bl[82] br[82] wl[93] vdd gnd cell_6t
Xbit_r94_c82 bl[82] br[82] wl[94] vdd gnd cell_6t
Xbit_r95_c82 bl[82] br[82] wl[95] vdd gnd cell_6t
Xbit_r96_c82 bl[82] br[82] wl[96] vdd gnd cell_6t
Xbit_r97_c82 bl[82] br[82] wl[97] vdd gnd cell_6t
Xbit_r98_c82 bl[82] br[82] wl[98] vdd gnd cell_6t
Xbit_r99_c82 bl[82] br[82] wl[99] vdd gnd cell_6t
Xbit_r100_c82 bl[82] br[82] wl[100] vdd gnd cell_6t
Xbit_r101_c82 bl[82] br[82] wl[101] vdd gnd cell_6t
Xbit_r102_c82 bl[82] br[82] wl[102] vdd gnd cell_6t
Xbit_r103_c82 bl[82] br[82] wl[103] vdd gnd cell_6t
Xbit_r104_c82 bl[82] br[82] wl[104] vdd gnd cell_6t
Xbit_r105_c82 bl[82] br[82] wl[105] vdd gnd cell_6t
Xbit_r106_c82 bl[82] br[82] wl[106] vdd gnd cell_6t
Xbit_r107_c82 bl[82] br[82] wl[107] vdd gnd cell_6t
Xbit_r108_c82 bl[82] br[82] wl[108] vdd gnd cell_6t
Xbit_r109_c82 bl[82] br[82] wl[109] vdd gnd cell_6t
Xbit_r110_c82 bl[82] br[82] wl[110] vdd gnd cell_6t
Xbit_r111_c82 bl[82] br[82] wl[111] vdd gnd cell_6t
Xbit_r112_c82 bl[82] br[82] wl[112] vdd gnd cell_6t
Xbit_r113_c82 bl[82] br[82] wl[113] vdd gnd cell_6t
Xbit_r114_c82 bl[82] br[82] wl[114] vdd gnd cell_6t
Xbit_r115_c82 bl[82] br[82] wl[115] vdd gnd cell_6t
Xbit_r116_c82 bl[82] br[82] wl[116] vdd gnd cell_6t
Xbit_r117_c82 bl[82] br[82] wl[117] vdd gnd cell_6t
Xbit_r118_c82 bl[82] br[82] wl[118] vdd gnd cell_6t
Xbit_r119_c82 bl[82] br[82] wl[119] vdd gnd cell_6t
Xbit_r120_c82 bl[82] br[82] wl[120] vdd gnd cell_6t
Xbit_r121_c82 bl[82] br[82] wl[121] vdd gnd cell_6t
Xbit_r122_c82 bl[82] br[82] wl[122] vdd gnd cell_6t
Xbit_r123_c82 bl[82] br[82] wl[123] vdd gnd cell_6t
Xbit_r124_c82 bl[82] br[82] wl[124] vdd gnd cell_6t
Xbit_r125_c82 bl[82] br[82] wl[125] vdd gnd cell_6t
Xbit_r126_c82 bl[82] br[82] wl[126] vdd gnd cell_6t
Xbit_r127_c82 bl[82] br[82] wl[127] vdd gnd cell_6t
Xbit_r128_c82 bl[82] br[82] wl[128] vdd gnd cell_6t
Xbit_r129_c82 bl[82] br[82] wl[129] vdd gnd cell_6t
Xbit_r130_c82 bl[82] br[82] wl[130] vdd gnd cell_6t
Xbit_r131_c82 bl[82] br[82] wl[131] vdd gnd cell_6t
Xbit_r132_c82 bl[82] br[82] wl[132] vdd gnd cell_6t
Xbit_r133_c82 bl[82] br[82] wl[133] vdd gnd cell_6t
Xbit_r134_c82 bl[82] br[82] wl[134] vdd gnd cell_6t
Xbit_r135_c82 bl[82] br[82] wl[135] vdd gnd cell_6t
Xbit_r136_c82 bl[82] br[82] wl[136] vdd gnd cell_6t
Xbit_r137_c82 bl[82] br[82] wl[137] vdd gnd cell_6t
Xbit_r138_c82 bl[82] br[82] wl[138] vdd gnd cell_6t
Xbit_r139_c82 bl[82] br[82] wl[139] vdd gnd cell_6t
Xbit_r140_c82 bl[82] br[82] wl[140] vdd gnd cell_6t
Xbit_r141_c82 bl[82] br[82] wl[141] vdd gnd cell_6t
Xbit_r142_c82 bl[82] br[82] wl[142] vdd gnd cell_6t
Xbit_r143_c82 bl[82] br[82] wl[143] vdd gnd cell_6t
Xbit_r144_c82 bl[82] br[82] wl[144] vdd gnd cell_6t
Xbit_r145_c82 bl[82] br[82] wl[145] vdd gnd cell_6t
Xbit_r146_c82 bl[82] br[82] wl[146] vdd gnd cell_6t
Xbit_r147_c82 bl[82] br[82] wl[147] vdd gnd cell_6t
Xbit_r148_c82 bl[82] br[82] wl[148] vdd gnd cell_6t
Xbit_r149_c82 bl[82] br[82] wl[149] vdd gnd cell_6t
Xbit_r150_c82 bl[82] br[82] wl[150] vdd gnd cell_6t
Xbit_r151_c82 bl[82] br[82] wl[151] vdd gnd cell_6t
Xbit_r152_c82 bl[82] br[82] wl[152] vdd gnd cell_6t
Xbit_r153_c82 bl[82] br[82] wl[153] vdd gnd cell_6t
Xbit_r154_c82 bl[82] br[82] wl[154] vdd gnd cell_6t
Xbit_r155_c82 bl[82] br[82] wl[155] vdd gnd cell_6t
Xbit_r156_c82 bl[82] br[82] wl[156] vdd gnd cell_6t
Xbit_r157_c82 bl[82] br[82] wl[157] vdd gnd cell_6t
Xbit_r158_c82 bl[82] br[82] wl[158] vdd gnd cell_6t
Xbit_r159_c82 bl[82] br[82] wl[159] vdd gnd cell_6t
Xbit_r160_c82 bl[82] br[82] wl[160] vdd gnd cell_6t
Xbit_r161_c82 bl[82] br[82] wl[161] vdd gnd cell_6t
Xbit_r162_c82 bl[82] br[82] wl[162] vdd gnd cell_6t
Xbit_r163_c82 bl[82] br[82] wl[163] vdd gnd cell_6t
Xbit_r164_c82 bl[82] br[82] wl[164] vdd gnd cell_6t
Xbit_r165_c82 bl[82] br[82] wl[165] vdd gnd cell_6t
Xbit_r166_c82 bl[82] br[82] wl[166] vdd gnd cell_6t
Xbit_r167_c82 bl[82] br[82] wl[167] vdd gnd cell_6t
Xbit_r168_c82 bl[82] br[82] wl[168] vdd gnd cell_6t
Xbit_r169_c82 bl[82] br[82] wl[169] vdd gnd cell_6t
Xbit_r170_c82 bl[82] br[82] wl[170] vdd gnd cell_6t
Xbit_r171_c82 bl[82] br[82] wl[171] vdd gnd cell_6t
Xbit_r172_c82 bl[82] br[82] wl[172] vdd gnd cell_6t
Xbit_r173_c82 bl[82] br[82] wl[173] vdd gnd cell_6t
Xbit_r174_c82 bl[82] br[82] wl[174] vdd gnd cell_6t
Xbit_r175_c82 bl[82] br[82] wl[175] vdd gnd cell_6t
Xbit_r176_c82 bl[82] br[82] wl[176] vdd gnd cell_6t
Xbit_r177_c82 bl[82] br[82] wl[177] vdd gnd cell_6t
Xbit_r178_c82 bl[82] br[82] wl[178] vdd gnd cell_6t
Xbit_r179_c82 bl[82] br[82] wl[179] vdd gnd cell_6t
Xbit_r180_c82 bl[82] br[82] wl[180] vdd gnd cell_6t
Xbit_r181_c82 bl[82] br[82] wl[181] vdd gnd cell_6t
Xbit_r182_c82 bl[82] br[82] wl[182] vdd gnd cell_6t
Xbit_r183_c82 bl[82] br[82] wl[183] vdd gnd cell_6t
Xbit_r184_c82 bl[82] br[82] wl[184] vdd gnd cell_6t
Xbit_r185_c82 bl[82] br[82] wl[185] vdd gnd cell_6t
Xbit_r186_c82 bl[82] br[82] wl[186] vdd gnd cell_6t
Xbit_r187_c82 bl[82] br[82] wl[187] vdd gnd cell_6t
Xbit_r188_c82 bl[82] br[82] wl[188] vdd gnd cell_6t
Xbit_r189_c82 bl[82] br[82] wl[189] vdd gnd cell_6t
Xbit_r190_c82 bl[82] br[82] wl[190] vdd gnd cell_6t
Xbit_r191_c82 bl[82] br[82] wl[191] vdd gnd cell_6t
Xbit_r192_c82 bl[82] br[82] wl[192] vdd gnd cell_6t
Xbit_r193_c82 bl[82] br[82] wl[193] vdd gnd cell_6t
Xbit_r194_c82 bl[82] br[82] wl[194] vdd gnd cell_6t
Xbit_r195_c82 bl[82] br[82] wl[195] vdd gnd cell_6t
Xbit_r196_c82 bl[82] br[82] wl[196] vdd gnd cell_6t
Xbit_r197_c82 bl[82] br[82] wl[197] vdd gnd cell_6t
Xbit_r198_c82 bl[82] br[82] wl[198] vdd gnd cell_6t
Xbit_r199_c82 bl[82] br[82] wl[199] vdd gnd cell_6t
Xbit_r200_c82 bl[82] br[82] wl[200] vdd gnd cell_6t
Xbit_r201_c82 bl[82] br[82] wl[201] vdd gnd cell_6t
Xbit_r202_c82 bl[82] br[82] wl[202] vdd gnd cell_6t
Xbit_r203_c82 bl[82] br[82] wl[203] vdd gnd cell_6t
Xbit_r204_c82 bl[82] br[82] wl[204] vdd gnd cell_6t
Xbit_r205_c82 bl[82] br[82] wl[205] vdd gnd cell_6t
Xbit_r206_c82 bl[82] br[82] wl[206] vdd gnd cell_6t
Xbit_r207_c82 bl[82] br[82] wl[207] vdd gnd cell_6t
Xbit_r208_c82 bl[82] br[82] wl[208] vdd gnd cell_6t
Xbit_r209_c82 bl[82] br[82] wl[209] vdd gnd cell_6t
Xbit_r210_c82 bl[82] br[82] wl[210] vdd gnd cell_6t
Xbit_r211_c82 bl[82] br[82] wl[211] vdd gnd cell_6t
Xbit_r212_c82 bl[82] br[82] wl[212] vdd gnd cell_6t
Xbit_r213_c82 bl[82] br[82] wl[213] vdd gnd cell_6t
Xbit_r214_c82 bl[82] br[82] wl[214] vdd gnd cell_6t
Xbit_r215_c82 bl[82] br[82] wl[215] vdd gnd cell_6t
Xbit_r216_c82 bl[82] br[82] wl[216] vdd gnd cell_6t
Xbit_r217_c82 bl[82] br[82] wl[217] vdd gnd cell_6t
Xbit_r218_c82 bl[82] br[82] wl[218] vdd gnd cell_6t
Xbit_r219_c82 bl[82] br[82] wl[219] vdd gnd cell_6t
Xbit_r220_c82 bl[82] br[82] wl[220] vdd gnd cell_6t
Xbit_r221_c82 bl[82] br[82] wl[221] vdd gnd cell_6t
Xbit_r222_c82 bl[82] br[82] wl[222] vdd gnd cell_6t
Xbit_r223_c82 bl[82] br[82] wl[223] vdd gnd cell_6t
Xbit_r224_c82 bl[82] br[82] wl[224] vdd gnd cell_6t
Xbit_r225_c82 bl[82] br[82] wl[225] vdd gnd cell_6t
Xbit_r226_c82 bl[82] br[82] wl[226] vdd gnd cell_6t
Xbit_r227_c82 bl[82] br[82] wl[227] vdd gnd cell_6t
Xbit_r228_c82 bl[82] br[82] wl[228] vdd gnd cell_6t
Xbit_r229_c82 bl[82] br[82] wl[229] vdd gnd cell_6t
Xbit_r230_c82 bl[82] br[82] wl[230] vdd gnd cell_6t
Xbit_r231_c82 bl[82] br[82] wl[231] vdd gnd cell_6t
Xbit_r232_c82 bl[82] br[82] wl[232] vdd gnd cell_6t
Xbit_r233_c82 bl[82] br[82] wl[233] vdd gnd cell_6t
Xbit_r234_c82 bl[82] br[82] wl[234] vdd gnd cell_6t
Xbit_r235_c82 bl[82] br[82] wl[235] vdd gnd cell_6t
Xbit_r236_c82 bl[82] br[82] wl[236] vdd gnd cell_6t
Xbit_r237_c82 bl[82] br[82] wl[237] vdd gnd cell_6t
Xbit_r238_c82 bl[82] br[82] wl[238] vdd gnd cell_6t
Xbit_r239_c82 bl[82] br[82] wl[239] vdd gnd cell_6t
Xbit_r240_c82 bl[82] br[82] wl[240] vdd gnd cell_6t
Xbit_r241_c82 bl[82] br[82] wl[241] vdd gnd cell_6t
Xbit_r242_c82 bl[82] br[82] wl[242] vdd gnd cell_6t
Xbit_r243_c82 bl[82] br[82] wl[243] vdd gnd cell_6t
Xbit_r244_c82 bl[82] br[82] wl[244] vdd gnd cell_6t
Xbit_r245_c82 bl[82] br[82] wl[245] vdd gnd cell_6t
Xbit_r246_c82 bl[82] br[82] wl[246] vdd gnd cell_6t
Xbit_r247_c82 bl[82] br[82] wl[247] vdd gnd cell_6t
Xbit_r248_c82 bl[82] br[82] wl[248] vdd gnd cell_6t
Xbit_r249_c82 bl[82] br[82] wl[249] vdd gnd cell_6t
Xbit_r250_c82 bl[82] br[82] wl[250] vdd gnd cell_6t
Xbit_r251_c82 bl[82] br[82] wl[251] vdd gnd cell_6t
Xbit_r252_c82 bl[82] br[82] wl[252] vdd gnd cell_6t
Xbit_r253_c82 bl[82] br[82] wl[253] vdd gnd cell_6t
Xbit_r254_c82 bl[82] br[82] wl[254] vdd gnd cell_6t
Xbit_r255_c82 bl[82] br[82] wl[255] vdd gnd cell_6t
Xbit_r256_c82 bl[82] br[82] wl[256] vdd gnd cell_6t
Xbit_r257_c82 bl[82] br[82] wl[257] vdd gnd cell_6t
Xbit_r258_c82 bl[82] br[82] wl[258] vdd gnd cell_6t
Xbit_r259_c82 bl[82] br[82] wl[259] vdd gnd cell_6t
Xbit_r260_c82 bl[82] br[82] wl[260] vdd gnd cell_6t
Xbit_r261_c82 bl[82] br[82] wl[261] vdd gnd cell_6t
Xbit_r262_c82 bl[82] br[82] wl[262] vdd gnd cell_6t
Xbit_r263_c82 bl[82] br[82] wl[263] vdd gnd cell_6t
Xbit_r264_c82 bl[82] br[82] wl[264] vdd gnd cell_6t
Xbit_r265_c82 bl[82] br[82] wl[265] vdd gnd cell_6t
Xbit_r266_c82 bl[82] br[82] wl[266] vdd gnd cell_6t
Xbit_r267_c82 bl[82] br[82] wl[267] vdd gnd cell_6t
Xbit_r268_c82 bl[82] br[82] wl[268] vdd gnd cell_6t
Xbit_r269_c82 bl[82] br[82] wl[269] vdd gnd cell_6t
Xbit_r270_c82 bl[82] br[82] wl[270] vdd gnd cell_6t
Xbit_r271_c82 bl[82] br[82] wl[271] vdd gnd cell_6t
Xbit_r272_c82 bl[82] br[82] wl[272] vdd gnd cell_6t
Xbit_r273_c82 bl[82] br[82] wl[273] vdd gnd cell_6t
Xbit_r274_c82 bl[82] br[82] wl[274] vdd gnd cell_6t
Xbit_r275_c82 bl[82] br[82] wl[275] vdd gnd cell_6t
Xbit_r276_c82 bl[82] br[82] wl[276] vdd gnd cell_6t
Xbit_r277_c82 bl[82] br[82] wl[277] vdd gnd cell_6t
Xbit_r278_c82 bl[82] br[82] wl[278] vdd gnd cell_6t
Xbit_r279_c82 bl[82] br[82] wl[279] vdd gnd cell_6t
Xbit_r280_c82 bl[82] br[82] wl[280] vdd gnd cell_6t
Xbit_r281_c82 bl[82] br[82] wl[281] vdd gnd cell_6t
Xbit_r282_c82 bl[82] br[82] wl[282] vdd gnd cell_6t
Xbit_r283_c82 bl[82] br[82] wl[283] vdd gnd cell_6t
Xbit_r284_c82 bl[82] br[82] wl[284] vdd gnd cell_6t
Xbit_r285_c82 bl[82] br[82] wl[285] vdd gnd cell_6t
Xbit_r286_c82 bl[82] br[82] wl[286] vdd gnd cell_6t
Xbit_r287_c82 bl[82] br[82] wl[287] vdd gnd cell_6t
Xbit_r288_c82 bl[82] br[82] wl[288] vdd gnd cell_6t
Xbit_r289_c82 bl[82] br[82] wl[289] vdd gnd cell_6t
Xbit_r290_c82 bl[82] br[82] wl[290] vdd gnd cell_6t
Xbit_r291_c82 bl[82] br[82] wl[291] vdd gnd cell_6t
Xbit_r292_c82 bl[82] br[82] wl[292] vdd gnd cell_6t
Xbit_r293_c82 bl[82] br[82] wl[293] vdd gnd cell_6t
Xbit_r294_c82 bl[82] br[82] wl[294] vdd gnd cell_6t
Xbit_r295_c82 bl[82] br[82] wl[295] vdd gnd cell_6t
Xbit_r296_c82 bl[82] br[82] wl[296] vdd gnd cell_6t
Xbit_r297_c82 bl[82] br[82] wl[297] vdd gnd cell_6t
Xbit_r298_c82 bl[82] br[82] wl[298] vdd gnd cell_6t
Xbit_r299_c82 bl[82] br[82] wl[299] vdd gnd cell_6t
Xbit_r300_c82 bl[82] br[82] wl[300] vdd gnd cell_6t
Xbit_r301_c82 bl[82] br[82] wl[301] vdd gnd cell_6t
Xbit_r302_c82 bl[82] br[82] wl[302] vdd gnd cell_6t
Xbit_r303_c82 bl[82] br[82] wl[303] vdd gnd cell_6t
Xbit_r304_c82 bl[82] br[82] wl[304] vdd gnd cell_6t
Xbit_r305_c82 bl[82] br[82] wl[305] vdd gnd cell_6t
Xbit_r306_c82 bl[82] br[82] wl[306] vdd gnd cell_6t
Xbit_r307_c82 bl[82] br[82] wl[307] vdd gnd cell_6t
Xbit_r308_c82 bl[82] br[82] wl[308] vdd gnd cell_6t
Xbit_r309_c82 bl[82] br[82] wl[309] vdd gnd cell_6t
Xbit_r310_c82 bl[82] br[82] wl[310] vdd gnd cell_6t
Xbit_r311_c82 bl[82] br[82] wl[311] vdd gnd cell_6t
Xbit_r312_c82 bl[82] br[82] wl[312] vdd gnd cell_6t
Xbit_r313_c82 bl[82] br[82] wl[313] vdd gnd cell_6t
Xbit_r314_c82 bl[82] br[82] wl[314] vdd gnd cell_6t
Xbit_r315_c82 bl[82] br[82] wl[315] vdd gnd cell_6t
Xbit_r316_c82 bl[82] br[82] wl[316] vdd gnd cell_6t
Xbit_r317_c82 bl[82] br[82] wl[317] vdd gnd cell_6t
Xbit_r318_c82 bl[82] br[82] wl[318] vdd gnd cell_6t
Xbit_r319_c82 bl[82] br[82] wl[319] vdd gnd cell_6t
Xbit_r320_c82 bl[82] br[82] wl[320] vdd gnd cell_6t
Xbit_r321_c82 bl[82] br[82] wl[321] vdd gnd cell_6t
Xbit_r322_c82 bl[82] br[82] wl[322] vdd gnd cell_6t
Xbit_r323_c82 bl[82] br[82] wl[323] vdd gnd cell_6t
Xbit_r324_c82 bl[82] br[82] wl[324] vdd gnd cell_6t
Xbit_r325_c82 bl[82] br[82] wl[325] vdd gnd cell_6t
Xbit_r326_c82 bl[82] br[82] wl[326] vdd gnd cell_6t
Xbit_r327_c82 bl[82] br[82] wl[327] vdd gnd cell_6t
Xbit_r328_c82 bl[82] br[82] wl[328] vdd gnd cell_6t
Xbit_r329_c82 bl[82] br[82] wl[329] vdd gnd cell_6t
Xbit_r330_c82 bl[82] br[82] wl[330] vdd gnd cell_6t
Xbit_r331_c82 bl[82] br[82] wl[331] vdd gnd cell_6t
Xbit_r332_c82 bl[82] br[82] wl[332] vdd gnd cell_6t
Xbit_r333_c82 bl[82] br[82] wl[333] vdd gnd cell_6t
Xbit_r334_c82 bl[82] br[82] wl[334] vdd gnd cell_6t
Xbit_r335_c82 bl[82] br[82] wl[335] vdd gnd cell_6t
Xbit_r336_c82 bl[82] br[82] wl[336] vdd gnd cell_6t
Xbit_r337_c82 bl[82] br[82] wl[337] vdd gnd cell_6t
Xbit_r338_c82 bl[82] br[82] wl[338] vdd gnd cell_6t
Xbit_r339_c82 bl[82] br[82] wl[339] vdd gnd cell_6t
Xbit_r340_c82 bl[82] br[82] wl[340] vdd gnd cell_6t
Xbit_r341_c82 bl[82] br[82] wl[341] vdd gnd cell_6t
Xbit_r342_c82 bl[82] br[82] wl[342] vdd gnd cell_6t
Xbit_r343_c82 bl[82] br[82] wl[343] vdd gnd cell_6t
Xbit_r344_c82 bl[82] br[82] wl[344] vdd gnd cell_6t
Xbit_r345_c82 bl[82] br[82] wl[345] vdd gnd cell_6t
Xbit_r346_c82 bl[82] br[82] wl[346] vdd gnd cell_6t
Xbit_r347_c82 bl[82] br[82] wl[347] vdd gnd cell_6t
Xbit_r348_c82 bl[82] br[82] wl[348] vdd gnd cell_6t
Xbit_r349_c82 bl[82] br[82] wl[349] vdd gnd cell_6t
Xbit_r350_c82 bl[82] br[82] wl[350] vdd gnd cell_6t
Xbit_r351_c82 bl[82] br[82] wl[351] vdd gnd cell_6t
Xbit_r352_c82 bl[82] br[82] wl[352] vdd gnd cell_6t
Xbit_r353_c82 bl[82] br[82] wl[353] vdd gnd cell_6t
Xbit_r354_c82 bl[82] br[82] wl[354] vdd gnd cell_6t
Xbit_r355_c82 bl[82] br[82] wl[355] vdd gnd cell_6t
Xbit_r356_c82 bl[82] br[82] wl[356] vdd gnd cell_6t
Xbit_r357_c82 bl[82] br[82] wl[357] vdd gnd cell_6t
Xbit_r358_c82 bl[82] br[82] wl[358] vdd gnd cell_6t
Xbit_r359_c82 bl[82] br[82] wl[359] vdd gnd cell_6t
Xbit_r360_c82 bl[82] br[82] wl[360] vdd gnd cell_6t
Xbit_r361_c82 bl[82] br[82] wl[361] vdd gnd cell_6t
Xbit_r362_c82 bl[82] br[82] wl[362] vdd gnd cell_6t
Xbit_r363_c82 bl[82] br[82] wl[363] vdd gnd cell_6t
Xbit_r364_c82 bl[82] br[82] wl[364] vdd gnd cell_6t
Xbit_r365_c82 bl[82] br[82] wl[365] vdd gnd cell_6t
Xbit_r366_c82 bl[82] br[82] wl[366] vdd gnd cell_6t
Xbit_r367_c82 bl[82] br[82] wl[367] vdd gnd cell_6t
Xbit_r368_c82 bl[82] br[82] wl[368] vdd gnd cell_6t
Xbit_r369_c82 bl[82] br[82] wl[369] vdd gnd cell_6t
Xbit_r370_c82 bl[82] br[82] wl[370] vdd gnd cell_6t
Xbit_r371_c82 bl[82] br[82] wl[371] vdd gnd cell_6t
Xbit_r372_c82 bl[82] br[82] wl[372] vdd gnd cell_6t
Xbit_r373_c82 bl[82] br[82] wl[373] vdd gnd cell_6t
Xbit_r374_c82 bl[82] br[82] wl[374] vdd gnd cell_6t
Xbit_r375_c82 bl[82] br[82] wl[375] vdd gnd cell_6t
Xbit_r376_c82 bl[82] br[82] wl[376] vdd gnd cell_6t
Xbit_r377_c82 bl[82] br[82] wl[377] vdd gnd cell_6t
Xbit_r378_c82 bl[82] br[82] wl[378] vdd gnd cell_6t
Xbit_r379_c82 bl[82] br[82] wl[379] vdd gnd cell_6t
Xbit_r380_c82 bl[82] br[82] wl[380] vdd gnd cell_6t
Xbit_r381_c82 bl[82] br[82] wl[381] vdd gnd cell_6t
Xbit_r382_c82 bl[82] br[82] wl[382] vdd gnd cell_6t
Xbit_r383_c82 bl[82] br[82] wl[383] vdd gnd cell_6t
Xbit_r384_c82 bl[82] br[82] wl[384] vdd gnd cell_6t
Xbit_r385_c82 bl[82] br[82] wl[385] vdd gnd cell_6t
Xbit_r386_c82 bl[82] br[82] wl[386] vdd gnd cell_6t
Xbit_r387_c82 bl[82] br[82] wl[387] vdd gnd cell_6t
Xbit_r388_c82 bl[82] br[82] wl[388] vdd gnd cell_6t
Xbit_r389_c82 bl[82] br[82] wl[389] vdd gnd cell_6t
Xbit_r390_c82 bl[82] br[82] wl[390] vdd gnd cell_6t
Xbit_r391_c82 bl[82] br[82] wl[391] vdd gnd cell_6t
Xbit_r392_c82 bl[82] br[82] wl[392] vdd gnd cell_6t
Xbit_r393_c82 bl[82] br[82] wl[393] vdd gnd cell_6t
Xbit_r394_c82 bl[82] br[82] wl[394] vdd gnd cell_6t
Xbit_r395_c82 bl[82] br[82] wl[395] vdd gnd cell_6t
Xbit_r396_c82 bl[82] br[82] wl[396] vdd gnd cell_6t
Xbit_r397_c82 bl[82] br[82] wl[397] vdd gnd cell_6t
Xbit_r398_c82 bl[82] br[82] wl[398] vdd gnd cell_6t
Xbit_r399_c82 bl[82] br[82] wl[399] vdd gnd cell_6t
Xbit_r400_c82 bl[82] br[82] wl[400] vdd gnd cell_6t
Xbit_r401_c82 bl[82] br[82] wl[401] vdd gnd cell_6t
Xbit_r402_c82 bl[82] br[82] wl[402] vdd gnd cell_6t
Xbit_r403_c82 bl[82] br[82] wl[403] vdd gnd cell_6t
Xbit_r404_c82 bl[82] br[82] wl[404] vdd gnd cell_6t
Xbit_r405_c82 bl[82] br[82] wl[405] vdd gnd cell_6t
Xbit_r406_c82 bl[82] br[82] wl[406] vdd gnd cell_6t
Xbit_r407_c82 bl[82] br[82] wl[407] vdd gnd cell_6t
Xbit_r408_c82 bl[82] br[82] wl[408] vdd gnd cell_6t
Xbit_r409_c82 bl[82] br[82] wl[409] vdd gnd cell_6t
Xbit_r410_c82 bl[82] br[82] wl[410] vdd gnd cell_6t
Xbit_r411_c82 bl[82] br[82] wl[411] vdd gnd cell_6t
Xbit_r412_c82 bl[82] br[82] wl[412] vdd gnd cell_6t
Xbit_r413_c82 bl[82] br[82] wl[413] vdd gnd cell_6t
Xbit_r414_c82 bl[82] br[82] wl[414] vdd gnd cell_6t
Xbit_r415_c82 bl[82] br[82] wl[415] vdd gnd cell_6t
Xbit_r416_c82 bl[82] br[82] wl[416] vdd gnd cell_6t
Xbit_r417_c82 bl[82] br[82] wl[417] vdd gnd cell_6t
Xbit_r418_c82 bl[82] br[82] wl[418] vdd gnd cell_6t
Xbit_r419_c82 bl[82] br[82] wl[419] vdd gnd cell_6t
Xbit_r420_c82 bl[82] br[82] wl[420] vdd gnd cell_6t
Xbit_r421_c82 bl[82] br[82] wl[421] vdd gnd cell_6t
Xbit_r422_c82 bl[82] br[82] wl[422] vdd gnd cell_6t
Xbit_r423_c82 bl[82] br[82] wl[423] vdd gnd cell_6t
Xbit_r424_c82 bl[82] br[82] wl[424] vdd gnd cell_6t
Xbit_r425_c82 bl[82] br[82] wl[425] vdd gnd cell_6t
Xbit_r426_c82 bl[82] br[82] wl[426] vdd gnd cell_6t
Xbit_r427_c82 bl[82] br[82] wl[427] vdd gnd cell_6t
Xbit_r428_c82 bl[82] br[82] wl[428] vdd gnd cell_6t
Xbit_r429_c82 bl[82] br[82] wl[429] vdd gnd cell_6t
Xbit_r430_c82 bl[82] br[82] wl[430] vdd gnd cell_6t
Xbit_r431_c82 bl[82] br[82] wl[431] vdd gnd cell_6t
Xbit_r432_c82 bl[82] br[82] wl[432] vdd gnd cell_6t
Xbit_r433_c82 bl[82] br[82] wl[433] vdd gnd cell_6t
Xbit_r434_c82 bl[82] br[82] wl[434] vdd gnd cell_6t
Xbit_r435_c82 bl[82] br[82] wl[435] vdd gnd cell_6t
Xbit_r436_c82 bl[82] br[82] wl[436] vdd gnd cell_6t
Xbit_r437_c82 bl[82] br[82] wl[437] vdd gnd cell_6t
Xbit_r438_c82 bl[82] br[82] wl[438] vdd gnd cell_6t
Xbit_r439_c82 bl[82] br[82] wl[439] vdd gnd cell_6t
Xbit_r440_c82 bl[82] br[82] wl[440] vdd gnd cell_6t
Xbit_r441_c82 bl[82] br[82] wl[441] vdd gnd cell_6t
Xbit_r442_c82 bl[82] br[82] wl[442] vdd gnd cell_6t
Xbit_r443_c82 bl[82] br[82] wl[443] vdd gnd cell_6t
Xbit_r444_c82 bl[82] br[82] wl[444] vdd gnd cell_6t
Xbit_r445_c82 bl[82] br[82] wl[445] vdd gnd cell_6t
Xbit_r446_c82 bl[82] br[82] wl[446] vdd gnd cell_6t
Xbit_r447_c82 bl[82] br[82] wl[447] vdd gnd cell_6t
Xbit_r448_c82 bl[82] br[82] wl[448] vdd gnd cell_6t
Xbit_r449_c82 bl[82] br[82] wl[449] vdd gnd cell_6t
Xbit_r450_c82 bl[82] br[82] wl[450] vdd gnd cell_6t
Xbit_r451_c82 bl[82] br[82] wl[451] vdd gnd cell_6t
Xbit_r452_c82 bl[82] br[82] wl[452] vdd gnd cell_6t
Xbit_r453_c82 bl[82] br[82] wl[453] vdd gnd cell_6t
Xbit_r454_c82 bl[82] br[82] wl[454] vdd gnd cell_6t
Xbit_r455_c82 bl[82] br[82] wl[455] vdd gnd cell_6t
Xbit_r456_c82 bl[82] br[82] wl[456] vdd gnd cell_6t
Xbit_r457_c82 bl[82] br[82] wl[457] vdd gnd cell_6t
Xbit_r458_c82 bl[82] br[82] wl[458] vdd gnd cell_6t
Xbit_r459_c82 bl[82] br[82] wl[459] vdd gnd cell_6t
Xbit_r460_c82 bl[82] br[82] wl[460] vdd gnd cell_6t
Xbit_r461_c82 bl[82] br[82] wl[461] vdd gnd cell_6t
Xbit_r462_c82 bl[82] br[82] wl[462] vdd gnd cell_6t
Xbit_r463_c82 bl[82] br[82] wl[463] vdd gnd cell_6t
Xbit_r464_c82 bl[82] br[82] wl[464] vdd gnd cell_6t
Xbit_r465_c82 bl[82] br[82] wl[465] vdd gnd cell_6t
Xbit_r466_c82 bl[82] br[82] wl[466] vdd gnd cell_6t
Xbit_r467_c82 bl[82] br[82] wl[467] vdd gnd cell_6t
Xbit_r468_c82 bl[82] br[82] wl[468] vdd gnd cell_6t
Xbit_r469_c82 bl[82] br[82] wl[469] vdd gnd cell_6t
Xbit_r470_c82 bl[82] br[82] wl[470] vdd gnd cell_6t
Xbit_r471_c82 bl[82] br[82] wl[471] vdd gnd cell_6t
Xbit_r472_c82 bl[82] br[82] wl[472] vdd gnd cell_6t
Xbit_r473_c82 bl[82] br[82] wl[473] vdd gnd cell_6t
Xbit_r474_c82 bl[82] br[82] wl[474] vdd gnd cell_6t
Xbit_r475_c82 bl[82] br[82] wl[475] vdd gnd cell_6t
Xbit_r476_c82 bl[82] br[82] wl[476] vdd gnd cell_6t
Xbit_r477_c82 bl[82] br[82] wl[477] vdd gnd cell_6t
Xbit_r478_c82 bl[82] br[82] wl[478] vdd gnd cell_6t
Xbit_r479_c82 bl[82] br[82] wl[479] vdd gnd cell_6t
Xbit_r480_c82 bl[82] br[82] wl[480] vdd gnd cell_6t
Xbit_r481_c82 bl[82] br[82] wl[481] vdd gnd cell_6t
Xbit_r482_c82 bl[82] br[82] wl[482] vdd gnd cell_6t
Xbit_r483_c82 bl[82] br[82] wl[483] vdd gnd cell_6t
Xbit_r484_c82 bl[82] br[82] wl[484] vdd gnd cell_6t
Xbit_r485_c82 bl[82] br[82] wl[485] vdd gnd cell_6t
Xbit_r486_c82 bl[82] br[82] wl[486] vdd gnd cell_6t
Xbit_r487_c82 bl[82] br[82] wl[487] vdd gnd cell_6t
Xbit_r488_c82 bl[82] br[82] wl[488] vdd gnd cell_6t
Xbit_r489_c82 bl[82] br[82] wl[489] vdd gnd cell_6t
Xbit_r490_c82 bl[82] br[82] wl[490] vdd gnd cell_6t
Xbit_r491_c82 bl[82] br[82] wl[491] vdd gnd cell_6t
Xbit_r492_c82 bl[82] br[82] wl[492] vdd gnd cell_6t
Xbit_r493_c82 bl[82] br[82] wl[493] vdd gnd cell_6t
Xbit_r494_c82 bl[82] br[82] wl[494] vdd gnd cell_6t
Xbit_r495_c82 bl[82] br[82] wl[495] vdd gnd cell_6t
Xbit_r496_c82 bl[82] br[82] wl[496] vdd gnd cell_6t
Xbit_r497_c82 bl[82] br[82] wl[497] vdd gnd cell_6t
Xbit_r498_c82 bl[82] br[82] wl[498] vdd gnd cell_6t
Xbit_r499_c82 bl[82] br[82] wl[499] vdd gnd cell_6t
Xbit_r500_c82 bl[82] br[82] wl[500] vdd gnd cell_6t
Xbit_r501_c82 bl[82] br[82] wl[501] vdd gnd cell_6t
Xbit_r502_c82 bl[82] br[82] wl[502] vdd gnd cell_6t
Xbit_r503_c82 bl[82] br[82] wl[503] vdd gnd cell_6t
Xbit_r504_c82 bl[82] br[82] wl[504] vdd gnd cell_6t
Xbit_r505_c82 bl[82] br[82] wl[505] vdd gnd cell_6t
Xbit_r506_c82 bl[82] br[82] wl[506] vdd gnd cell_6t
Xbit_r507_c82 bl[82] br[82] wl[507] vdd gnd cell_6t
Xbit_r508_c82 bl[82] br[82] wl[508] vdd gnd cell_6t
Xbit_r509_c82 bl[82] br[82] wl[509] vdd gnd cell_6t
Xbit_r510_c82 bl[82] br[82] wl[510] vdd gnd cell_6t
Xbit_r511_c82 bl[82] br[82] wl[511] vdd gnd cell_6t
Xbit_r0_c83 bl[83] br[83] wl[0] vdd gnd cell_6t
Xbit_r1_c83 bl[83] br[83] wl[1] vdd gnd cell_6t
Xbit_r2_c83 bl[83] br[83] wl[2] vdd gnd cell_6t
Xbit_r3_c83 bl[83] br[83] wl[3] vdd gnd cell_6t
Xbit_r4_c83 bl[83] br[83] wl[4] vdd gnd cell_6t
Xbit_r5_c83 bl[83] br[83] wl[5] vdd gnd cell_6t
Xbit_r6_c83 bl[83] br[83] wl[6] vdd gnd cell_6t
Xbit_r7_c83 bl[83] br[83] wl[7] vdd gnd cell_6t
Xbit_r8_c83 bl[83] br[83] wl[8] vdd gnd cell_6t
Xbit_r9_c83 bl[83] br[83] wl[9] vdd gnd cell_6t
Xbit_r10_c83 bl[83] br[83] wl[10] vdd gnd cell_6t
Xbit_r11_c83 bl[83] br[83] wl[11] vdd gnd cell_6t
Xbit_r12_c83 bl[83] br[83] wl[12] vdd gnd cell_6t
Xbit_r13_c83 bl[83] br[83] wl[13] vdd gnd cell_6t
Xbit_r14_c83 bl[83] br[83] wl[14] vdd gnd cell_6t
Xbit_r15_c83 bl[83] br[83] wl[15] vdd gnd cell_6t
Xbit_r16_c83 bl[83] br[83] wl[16] vdd gnd cell_6t
Xbit_r17_c83 bl[83] br[83] wl[17] vdd gnd cell_6t
Xbit_r18_c83 bl[83] br[83] wl[18] vdd gnd cell_6t
Xbit_r19_c83 bl[83] br[83] wl[19] vdd gnd cell_6t
Xbit_r20_c83 bl[83] br[83] wl[20] vdd gnd cell_6t
Xbit_r21_c83 bl[83] br[83] wl[21] vdd gnd cell_6t
Xbit_r22_c83 bl[83] br[83] wl[22] vdd gnd cell_6t
Xbit_r23_c83 bl[83] br[83] wl[23] vdd gnd cell_6t
Xbit_r24_c83 bl[83] br[83] wl[24] vdd gnd cell_6t
Xbit_r25_c83 bl[83] br[83] wl[25] vdd gnd cell_6t
Xbit_r26_c83 bl[83] br[83] wl[26] vdd gnd cell_6t
Xbit_r27_c83 bl[83] br[83] wl[27] vdd gnd cell_6t
Xbit_r28_c83 bl[83] br[83] wl[28] vdd gnd cell_6t
Xbit_r29_c83 bl[83] br[83] wl[29] vdd gnd cell_6t
Xbit_r30_c83 bl[83] br[83] wl[30] vdd gnd cell_6t
Xbit_r31_c83 bl[83] br[83] wl[31] vdd gnd cell_6t
Xbit_r32_c83 bl[83] br[83] wl[32] vdd gnd cell_6t
Xbit_r33_c83 bl[83] br[83] wl[33] vdd gnd cell_6t
Xbit_r34_c83 bl[83] br[83] wl[34] vdd gnd cell_6t
Xbit_r35_c83 bl[83] br[83] wl[35] vdd gnd cell_6t
Xbit_r36_c83 bl[83] br[83] wl[36] vdd gnd cell_6t
Xbit_r37_c83 bl[83] br[83] wl[37] vdd gnd cell_6t
Xbit_r38_c83 bl[83] br[83] wl[38] vdd gnd cell_6t
Xbit_r39_c83 bl[83] br[83] wl[39] vdd gnd cell_6t
Xbit_r40_c83 bl[83] br[83] wl[40] vdd gnd cell_6t
Xbit_r41_c83 bl[83] br[83] wl[41] vdd gnd cell_6t
Xbit_r42_c83 bl[83] br[83] wl[42] vdd gnd cell_6t
Xbit_r43_c83 bl[83] br[83] wl[43] vdd gnd cell_6t
Xbit_r44_c83 bl[83] br[83] wl[44] vdd gnd cell_6t
Xbit_r45_c83 bl[83] br[83] wl[45] vdd gnd cell_6t
Xbit_r46_c83 bl[83] br[83] wl[46] vdd gnd cell_6t
Xbit_r47_c83 bl[83] br[83] wl[47] vdd gnd cell_6t
Xbit_r48_c83 bl[83] br[83] wl[48] vdd gnd cell_6t
Xbit_r49_c83 bl[83] br[83] wl[49] vdd gnd cell_6t
Xbit_r50_c83 bl[83] br[83] wl[50] vdd gnd cell_6t
Xbit_r51_c83 bl[83] br[83] wl[51] vdd gnd cell_6t
Xbit_r52_c83 bl[83] br[83] wl[52] vdd gnd cell_6t
Xbit_r53_c83 bl[83] br[83] wl[53] vdd gnd cell_6t
Xbit_r54_c83 bl[83] br[83] wl[54] vdd gnd cell_6t
Xbit_r55_c83 bl[83] br[83] wl[55] vdd gnd cell_6t
Xbit_r56_c83 bl[83] br[83] wl[56] vdd gnd cell_6t
Xbit_r57_c83 bl[83] br[83] wl[57] vdd gnd cell_6t
Xbit_r58_c83 bl[83] br[83] wl[58] vdd gnd cell_6t
Xbit_r59_c83 bl[83] br[83] wl[59] vdd gnd cell_6t
Xbit_r60_c83 bl[83] br[83] wl[60] vdd gnd cell_6t
Xbit_r61_c83 bl[83] br[83] wl[61] vdd gnd cell_6t
Xbit_r62_c83 bl[83] br[83] wl[62] vdd gnd cell_6t
Xbit_r63_c83 bl[83] br[83] wl[63] vdd gnd cell_6t
Xbit_r64_c83 bl[83] br[83] wl[64] vdd gnd cell_6t
Xbit_r65_c83 bl[83] br[83] wl[65] vdd gnd cell_6t
Xbit_r66_c83 bl[83] br[83] wl[66] vdd gnd cell_6t
Xbit_r67_c83 bl[83] br[83] wl[67] vdd gnd cell_6t
Xbit_r68_c83 bl[83] br[83] wl[68] vdd gnd cell_6t
Xbit_r69_c83 bl[83] br[83] wl[69] vdd gnd cell_6t
Xbit_r70_c83 bl[83] br[83] wl[70] vdd gnd cell_6t
Xbit_r71_c83 bl[83] br[83] wl[71] vdd gnd cell_6t
Xbit_r72_c83 bl[83] br[83] wl[72] vdd gnd cell_6t
Xbit_r73_c83 bl[83] br[83] wl[73] vdd gnd cell_6t
Xbit_r74_c83 bl[83] br[83] wl[74] vdd gnd cell_6t
Xbit_r75_c83 bl[83] br[83] wl[75] vdd gnd cell_6t
Xbit_r76_c83 bl[83] br[83] wl[76] vdd gnd cell_6t
Xbit_r77_c83 bl[83] br[83] wl[77] vdd gnd cell_6t
Xbit_r78_c83 bl[83] br[83] wl[78] vdd gnd cell_6t
Xbit_r79_c83 bl[83] br[83] wl[79] vdd gnd cell_6t
Xbit_r80_c83 bl[83] br[83] wl[80] vdd gnd cell_6t
Xbit_r81_c83 bl[83] br[83] wl[81] vdd gnd cell_6t
Xbit_r82_c83 bl[83] br[83] wl[82] vdd gnd cell_6t
Xbit_r83_c83 bl[83] br[83] wl[83] vdd gnd cell_6t
Xbit_r84_c83 bl[83] br[83] wl[84] vdd gnd cell_6t
Xbit_r85_c83 bl[83] br[83] wl[85] vdd gnd cell_6t
Xbit_r86_c83 bl[83] br[83] wl[86] vdd gnd cell_6t
Xbit_r87_c83 bl[83] br[83] wl[87] vdd gnd cell_6t
Xbit_r88_c83 bl[83] br[83] wl[88] vdd gnd cell_6t
Xbit_r89_c83 bl[83] br[83] wl[89] vdd gnd cell_6t
Xbit_r90_c83 bl[83] br[83] wl[90] vdd gnd cell_6t
Xbit_r91_c83 bl[83] br[83] wl[91] vdd gnd cell_6t
Xbit_r92_c83 bl[83] br[83] wl[92] vdd gnd cell_6t
Xbit_r93_c83 bl[83] br[83] wl[93] vdd gnd cell_6t
Xbit_r94_c83 bl[83] br[83] wl[94] vdd gnd cell_6t
Xbit_r95_c83 bl[83] br[83] wl[95] vdd gnd cell_6t
Xbit_r96_c83 bl[83] br[83] wl[96] vdd gnd cell_6t
Xbit_r97_c83 bl[83] br[83] wl[97] vdd gnd cell_6t
Xbit_r98_c83 bl[83] br[83] wl[98] vdd gnd cell_6t
Xbit_r99_c83 bl[83] br[83] wl[99] vdd gnd cell_6t
Xbit_r100_c83 bl[83] br[83] wl[100] vdd gnd cell_6t
Xbit_r101_c83 bl[83] br[83] wl[101] vdd gnd cell_6t
Xbit_r102_c83 bl[83] br[83] wl[102] vdd gnd cell_6t
Xbit_r103_c83 bl[83] br[83] wl[103] vdd gnd cell_6t
Xbit_r104_c83 bl[83] br[83] wl[104] vdd gnd cell_6t
Xbit_r105_c83 bl[83] br[83] wl[105] vdd gnd cell_6t
Xbit_r106_c83 bl[83] br[83] wl[106] vdd gnd cell_6t
Xbit_r107_c83 bl[83] br[83] wl[107] vdd gnd cell_6t
Xbit_r108_c83 bl[83] br[83] wl[108] vdd gnd cell_6t
Xbit_r109_c83 bl[83] br[83] wl[109] vdd gnd cell_6t
Xbit_r110_c83 bl[83] br[83] wl[110] vdd gnd cell_6t
Xbit_r111_c83 bl[83] br[83] wl[111] vdd gnd cell_6t
Xbit_r112_c83 bl[83] br[83] wl[112] vdd gnd cell_6t
Xbit_r113_c83 bl[83] br[83] wl[113] vdd gnd cell_6t
Xbit_r114_c83 bl[83] br[83] wl[114] vdd gnd cell_6t
Xbit_r115_c83 bl[83] br[83] wl[115] vdd gnd cell_6t
Xbit_r116_c83 bl[83] br[83] wl[116] vdd gnd cell_6t
Xbit_r117_c83 bl[83] br[83] wl[117] vdd gnd cell_6t
Xbit_r118_c83 bl[83] br[83] wl[118] vdd gnd cell_6t
Xbit_r119_c83 bl[83] br[83] wl[119] vdd gnd cell_6t
Xbit_r120_c83 bl[83] br[83] wl[120] vdd gnd cell_6t
Xbit_r121_c83 bl[83] br[83] wl[121] vdd gnd cell_6t
Xbit_r122_c83 bl[83] br[83] wl[122] vdd gnd cell_6t
Xbit_r123_c83 bl[83] br[83] wl[123] vdd gnd cell_6t
Xbit_r124_c83 bl[83] br[83] wl[124] vdd gnd cell_6t
Xbit_r125_c83 bl[83] br[83] wl[125] vdd gnd cell_6t
Xbit_r126_c83 bl[83] br[83] wl[126] vdd gnd cell_6t
Xbit_r127_c83 bl[83] br[83] wl[127] vdd gnd cell_6t
Xbit_r128_c83 bl[83] br[83] wl[128] vdd gnd cell_6t
Xbit_r129_c83 bl[83] br[83] wl[129] vdd gnd cell_6t
Xbit_r130_c83 bl[83] br[83] wl[130] vdd gnd cell_6t
Xbit_r131_c83 bl[83] br[83] wl[131] vdd gnd cell_6t
Xbit_r132_c83 bl[83] br[83] wl[132] vdd gnd cell_6t
Xbit_r133_c83 bl[83] br[83] wl[133] vdd gnd cell_6t
Xbit_r134_c83 bl[83] br[83] wl[134] vdd gnd cell_6t
Xbit_r135_c83 bl[83] br[83] wl[135] vdd gnd cell_6t
Xbit_r136_c83 bl[83] br[83] wl[136] vdd gnd cell_6t
Xbit_r137_c83 bl[83] br[83] wl[137] vdd gnd cell_6t
Xbit_r138_c83 bl[83] br[83] wl[138] vdd gnd cell_6t
Xbit_r139_c83 bl[83] br[83] wl[139] vdd gnd cell_6t
Xbit_r140_c83 bl[83] br[83] wl[140] vdd gnd cell_6t
Xbit_r141_c83 bl[83] br[83] wl[141] vdd gnd cell_6t
Xbit_r142_c83 bl[83] br[83] wl[142] vdd gnd cell_6t
Xbit_r143_c83 bl[83] br[83] wl[143] vdd gnd cell_6t
Xbit_r144_c83 bl[83] br[83] wl[144] vdd gnd cell_6t
Xbit_r145_c83 bl[83] br[83] wl[145] vdd gnd cell_6t
Xbit_r146_c83 bl[83] br[83] wl[146] vdd gnd cell_6t
Xbit_r147_c83 bl[83] br[83] wl[147] vdd gnd cell_6t
Xbit_r148_c83 bl[83] br[83] wl[148] vdd gnd cell_6t
Xbit_r149_c83 bl[83] br[83] wl[149] vdd gnd cell_6t
Xbit_r150_c83 bl[83] br[83] wl[150] vdd gnd cell_6t
Xbit_r151_c83 bl[83] br[83] wl[151] vdd gnd cell_6t
Xbit_r152_c83 bl[83] br[83] wl[152] vdd gnd cell_6t
Xbit_r153_c83 bl[83] br[83] wl[153] vdd gnd cell_6t
Xbit_r154_c83 bl[83] br[83] wl[154] vdd gnd cell_6t
Xbit_r155_c83 bl[83] br[83] wl[155] vdd gnd cell_6t
Xbit_r156_c83 bl[83] br[83] wl[156] vdd gnd cell_6t
Xbit_r157_c83 bl[83] br[83] wl[157] vdd gnd cell_6t
Xbit_r158_c83 bl[83] br[83] wl[158] vdd gnd cell_6t
Xbit_r159_c83 bl[83] br[83] wl[159] vdd gnd cell_6t
Xbit_r160_c83 bl[83] br[83] wl[160] vdd gnd cell_6t
Xbit_r161_c83 bl[83] br[83] wl[161] vdd gnd cell_6t
Xbit_r162_c83 bl[83] br[83] wl[162] vdd gnd cell_6t
Xbit_r163_c83 bl[83] br[83] wl[163] vdd gnd cell_6t
Xbit_r164_c83 bl[83] br[83] wl[164] vdd gnd cell_6t
Xbit_r165_c83 bl[83] br[83] wl[165] vdd gnd cell_6t
Xbit_r166_c83 bl[83] br[83] wl[166] vdd gnd cell_6t
Xbit_r167_c83 bl[83] br[83] wl[167] vdd gnd cell_6t
Xbit_r168_c83 bl[83] br[83] wl[168] vdd gnd cell_6t
Xbit_r169_c83 bl[83] br[83] wl[169] vdd gnd cell_6t
Xbit_r170_c83 bl[83] br[83] wl[170] vdd gnd cell_6t
Xbit_r171_c83 bl[83] br[83] wl[171] vdd gnd cell_6t
Xbit_r172_c83 bl[83] br[83] wl[172] vdd gnd cell_6t
Xbit_r173_c83 bl[83] br[83] wl[173] vdd gnd cell_6t
Xbit_r174_c83 bl[83] br[83] wl[174] vdd gnd cell_6t
Xbit_r175_c83 bl[83] br[83] wl[175] vdd gnd cell_6t
Xbit_r176_c83 bl[83] br[83] wl[176] vdd gnd cell_6t
Xbit_r177_c83 bl[83] br[83] wl[177] vdd gnd cell_6t
Xbit_r178_c83 bl[83] br[83] wl[178] vdd gnd cell_6t
Xbit_r179_c83 bl[83] br[83] wl[179] vdd gnd cell_6t
Xbit_r180_c83 bl[83] br[83] wl[180] vdd gnd cell_6t
Xbit_r181_c83 bl[83] br[83] wl[181] vdd gnd cell_6t
Xbit_r182_c83 bl[83] br[83] wl[182] vdd gnd cell_6t
Xbit_r183_c83 bl[83] br[83] wl[183] vdd gnd cell_6t
Xbit_r184_c83 bl[83] br[83] wl[184] vdd gnd cell_6t
Xbit_r185_c83 bl[83] br[83] wl[185] vdd gnd cell_6t
Xbit_r186_c83 bl[83] br[83] wl[186] vdd gnd cell_6t
Xbit_r187_c83 bl[83] br[83] wl[187] vdd gnd cell_6t
Xbit_r188_c83 bl[83] br[83] wl[188] vdd gnd cell_6t
Xbit_r189_c83 bl[83] br[83] wl[189] vdd gnd cell_6t
Xbit_r190_c83 bl[83] br[83] wl[190] vdd gnd cell_6t
Xbit_r191_c83 bl[83] br[83] wl[191] vdd gnd cell_6t
Xbit_r192_c83 bl[83] br[83] wl[192] vdd gnd cell_6t
Xbit_r193_c83 bl[83] br[83] wl[193] vdd gnd cell_6t
Xbit_r194_c83 bl[83] br[83] wl[194] vdd gnd cell_6t
Xbit_r195_c83 bl[83] br[83] wl[195] vdd gnd cell_6t
Xbit_r196_c83 bl[83] br[83] wl[196] vdd gnd cell_6t
Xbit_r197_c83 bl[83] br[83] wl[197] vdd gnd cell_6t
Xbit_r198_c83 bl[83] br[83] wl[198] vdd gnd cell_6t
Xbit_r199_c83 bl[83] br[83] wl[199] vdd gnd cell_6t
Xbit_r200_c83 bl[83] br[83] wl[200] vdd gnd cell_6t
Xbit_r201_c83 bl[83] br[83] wl[201] vdd gnd cell_6t
Xbit_r202_c83 bl[83] br[83] wl[202] vdd gnd cell_6t
Xbit_r203_c83 bl[83] br[83] wl[203] vdd gnd cell_6t
Xbit_r204_c83 bl[83] br[83] wl[204] vdd gnd cell_6t
Xbit_r205_c83 bl[83] br[83] wl[205] vdd gnd cell_6t
Xbit_r206_c83 bl[83] br[83] wl[206] vdd gnd cell_6t
Xbit_r207_c83 bl[83] br[83] wl[207] vdd gnd cell_6t
Xbit_r208_c83 bl[83] br[83] wl[208] vdd gnd cell_6t
Xbit_r209_c83 bl[83] br[83] wl[209] vdd gnd cell_6t
Xbit_r210_c83 bl[83] br[83] wl[210] vdd gnd cell_6t
Xbit_r211_c83 bl[83] br[83] wl[211] vdd gnd cell_6t
Xbit_r212_c83 bl[83] br[83] wl[212] vdd gnd cell_6t
Xbit_r213_c83 bl[83] br[83] wl[213] vdd gnd cell_6t
Xbit_r214_c83 bl[83] br[83] wl[214] vdd gnd cell_6t
Xbit_r215_c83 bl[83] br[83] wl[215] vdd gnd cell_6t
Xbit_r216_c83 bl[83] br[83] wl[216] vdd gnd cell_6t
Xbit_r217_c83 bl[83] br[83] wl[217] vdd gnd cell_6t
Xbit_r218_c83 bl[83] br[83] wl[218] vdd gnd cell_6t
Xbit_r219_c83 bl[83] br[83] wl[219] vdd gnd cell_6t
Xbit_r220_c83 bl[83] br[83] wl[220] vdd gnd cell_6t
Xbit_r221_c83 bl[83] br[83] wl[221] vdd gnd cell_6t
Xbit_r222_c83 bl[83] br[83] wl[222] vdd gnd cell_6t
Xbit_r223_c83 bl[83] br[83] wl[223] vdd gnd cell_6t
Xbit_r224_c83 bl[83] br[83] wl[224] vdd gnd cell_6t
Xbit_r225_c83 bl[83] br[83] wl[225] vdd gnd cell_6t
Xbit_r226_c83 bl[83] br[83] wl[226] vdd gnd cell_6t
Xbit_r227_c83 bl[83] br[83] wl[227] vdd gnd cell_6t
Xbit_r228_c83 bl[83] br[83] wl[228] vdd gnd cell_6t
Xbit_r229_c83 bl[83] br[83] wl[229] vdd gnd cell_6t
Xbit_r230_c83 bl[83] br[83] wl[230] vdd gnd cell_6t
Xbit_r231_c83 bl[83] br[83] wl[231] vdd gnd cell_6t
Xbit_r232_c83 bl[83] br[83] wl[232] vdd gnd cell_6t
Xbit_r233_c83 bl[83] br[83] wl[233] vdd gnd cell_6t
Xbit_r234_c83 bl[83] br[83] wl[234] vdd gnd cell_6t
Xbit_r235_c83 bl[83] br[83] wl[235] vdd gnd cell_6t
Xbit_r236_c83 bl[83] br[83] wl[236] vdd gnd cell_6t
Xbit_r237_c83 bl[83] br[83] wl[237] vdd gnd cell_6t
Xbit_r238_c83 bl[83] br[83] wl[238] vdd gnd cell_6t
Xbit_r239_c83 bl[83] br[83] wl[239] vdd gnd cell_6t
Xbit_r240_c83 bl[83] br[83] wl[240] vdd gnd cell_6t
Xbit_r241_c83 bl[83] br[83] wl[241] vdd gnd cell_6t
Xbit_r242_c83 bl[83] br[83] wl[242] vdd gnd cell_6t
Xbit_r243_c83 bl[83] br[83] wl[243] vdd gnd cell_6t
Xbit_r244_c83 bl[83] br[83] wl[244] vdd gnd cell_6t
Xbit_r245_c83 bl[83] br[83] wl[245] vdd gnd cell_6t
Xbit_r246_c83 bl[83] br[83] wl[246] vdd gnd cell_6t
Xbit_r247_c83 bl[83] br[83] wl[247] vdd gnd cell_6t
Xbit_r248_c83 bl[83] br[83] wl[248] vdd gnd cell_6t
Xbit_r249_c83 bl[83] br[83] wl[249] vdd gnd cell_6t
Xbit_r250_c83 bl[83] br[83] wl[250] vdd gnd cell_6t
Xbit_r251_c83 bl[83] br[83] wl[251] vdd gnd cell_6t
Xbit_r252_c83 bl[83] br[83] wl[252] vdd gnd cell_6t
Xbit_r253_c83 bl[83] br[83] wl[253] vdd gnd cell_6t
Xbit_r254_c83 bl[83] br[83] wl[254] vdd gnd cell_6t
Xbit_r255_c83 bl[83] br[83] wl[255] vdd gnd cell_6t
Xbit_r256_c83 bl[83] br[83] wl[256] vdd gnd cell_6t
Xbit_r257_c83 bl[83] br[83] wl[257] vdd gnd cell_6t
Xbit_r258_c83 bl[83] br[83] wl[258] vdd gnd cell_6t
Xbit_r259_c83 bl[83] br[83] wl[259] vdd gnd cell_6t
Xbit_r260_c83 bl[83] br[83] wl[260] vdd gnd cell_6t
Xbit_r261_c83 bl[83] br[83] wl[261] vdd gnd cell_6t
Xbit_r262_c83 bl[83] br[83] wl[262] vdd gnd cell_6t
Xbit_r263_c83 bl[83] br[83] wl[263] vdd gnd cell_6t
Xbit_r264_c83 bl[83] br[83] wl[264] vdd gnd cell_6t
Xbit_r265_c83 bl[83] br[83] wl[265] vdd gnd cell_6t
Xbit_r266_c83 bl[83] br[83] wl[266] vdd gnd cell_6t
Xbit_r267_c83 bl[83] br[83] wl[267] vdd gnd cell_6t
Xbit_r268_c83 bl[83] br[83] wl[268] vdd gnd cell_6t
Xbit_r269_c83 bl[83] br[83] wl[269] vdd gnd cell_6t
Xbit_r270_c83 bl[83] br[83] wl[270] vdd gnd cell_6t
Xbit_r271_c83 bl[83] br[83] wl[271] vdd gnd cell_6t
Xbit_r272_c83 bl[83] br[83] wl[272] vdd gnd cell_6t
Xbit_r273_c83 bl[83] br[83] wl[273] vdd gnd cell_6t
Xbit_r274_c83 bl[83] br[83] wl[274] vdd gnd cell_6t
Xbit_r275_c83 bl[83] br[83] wl[275] vdd gnd cell_6t
Xbit_r276_c83 bl[83] br[83] wl[276] vdd gnd cell_6t
Xbit_r277_c83 bl[83] br[83] wl[277] vdd gnd cell_6t
Xbit_r278_c83 bl[83] br[83] wl[278] vdd gnd cell_6t
Xbit_r279_c83 bl[83] br[83] wl[279] vdd gnd cell_6t
Xbit_r280_c83 bl[83] br[83] wl[280] vdd gnd cell_6t
Xbit_r281_c83 bl[83] br[83] wl[281] vdd gnd cell_6t
Xbit_r282_c83 bl[83] br[83] wl[282] vdd gnd cell_6t
Xbit_r283_c83 bl[83] br[83] wl[283] vdd gnd cell_6t
Xbit_r284_c83 bl[83] br[83] wl[284] vdd gnd cell_6t
Xbit_r285_c83 bl[83] br[83] wl[285] vdd gnd cell_6t
Xbit_r286_c83 bl[83] br[83] wl[286] vdd gnd cell_6t
Xbit_r287_c83 bl[83] br[83] wl[287] vdd gnd cell_6t
Xbit_r288_c83 bl[83] br[83] wl[288] vdd gnd cell_6t
Xbit_r289_c83 bl[83] br[83] wl[289] vdd gnd cell_6t
Xbit_r290_c83 bl[83] br[83] wl[290] vdd gnd cell_6t
Xbit_r291_c83 bl[83] br[83] wl[291] vdd gnd cell_6t
Xbit_r292_c83 bl[83] br[83] wl[292] vdd gnd cell_6t
Xbit_r293_c83 bl[83] br[83] wl[293] vdd gnd cell_6t
Xbit_r294_c83 bl[83] br[83] wl[294] vdd gnd cell_6t
Xbit_r295_c83 bl[83] br[83] wl[295] vdd gnd cell_6t
Xbit_r296_c83 bl[83] br[83] wl[296] vdd gnd cell_6t
Xbit_r297_c83 bl[83] br[83] wl[297] vdd gnd cell_6t
Xbit_r298_c83 bl[83] br[83] wl[298] vdd gnd cell_6t
Xbit_r299_c83 bl[83] br[83] wl[299] vdd gnd cell_6t
Xbit_r300_c83 bl[83] br[83] wl[300] vdd gnd cell_6t
Xbit_r301_c83 bl[83] br[83] wl[301] vdd gnd cell_6t
Xbit_r302_c83 bl[83] br[83] wl[302] vdd gnd cell_6t
Xbit_r303_c83 bl[83] br[83] wl[303] vdd gnd cell_6t
Xbit_r304_c83 bl[83] br[83] wl[304] vdd gnd cell_6t
Xbit_r305_c83 bl[83] br[83] wl[305] vdd gnd cell_6t
Xbit_r306_c83 bl[83] br[83] wl[306] vdd gnd cell_6t
Xbit_r307_c83 bl[83] br[83] wl[307] vdd gnd cell_6t
Xbit_r308_c83 bl[83] br[83] wl[308] vdd gnd cell_6t
Xbit_r309_c83 bl[83] br[83] wl[309] vdd gnd cell_6t
Xbit_r310_c83 bl[83] br[83] wl[310] vdd gnd cell_6t
Xbit_r311_c83 bl[83] br[83] wl[311] vdd gnd cell_6t
Xbit_r312_c83 bl[83] br[83] wl[312] vdd gnd cell_6t
Xbit_r313_c83 bl[83] br[83] wl[313] vdd gnd cell_6t
Xbit_r314_c83 bl[83] br[83] wl[314] vdd gnd cell_6t
Xbit_r315_c83 bl[83] br[83] wl[315] vdd gnd cell_6t
Xbit_r316_c83 bl[83] br[83] wl[316] vdd gnd cell_6t
Xbit_r317_c83 bl[83] br[83] wl[317] vdd gnd cell_6t
Xbit_r318_c83 bl[83] br[83] wl[318] vdd gnd cell_6t
Xbit_r319_c83 bl[83] br[83] wl[319] vdd gnd cell_6t
Xbit_r320_c83 bl[83] br[83] wl[320] vdd gnd cell_6t
Xbit_r321_c83 bl[83] br[83] wl[321] vdd gnd cell_6t
Xbit_r322_c83 bl[83] br[83] wl[322] vdd gnd cell_6t
Xbit_r323_c83 bl[83] br[83] wl[323] vdd gnd cell_6t
Xbit_r324_c83 bl[83] br[83] wl[324] vdd gnd cell_6t
Xbit_r325_c83 bl[83] br[83] wl[325] vdd gnd cell_6t
Xbit_r326_c83 bl[83] br[83] wl[326] vdd gnd cell_6t
Xbit_r327_c83 bl[83] br[83] wl[327] vdd gnd cell_6t
Xbit_r328_c83 bl[83] br[83] wl[328] vdd gnd cell_6t
Xbit_r329_c83 bl[83] br[83] wl[329] vdd gnd cell_6t
Xbit_r330_c83 bl[83] br[83] wl[330] vdd gnd cell_6t
Xbit_r331_c83 bl[83] br[83] wl[331] vdd gnd cell_6t
Xbit_r332_c83 bl[83] br[83] wl[332] vdd gnd cell_6t
Xbit_r333_c83 bl[83] br[83] wl[333] vdd gnd cell_6t
Xbit_r334_c83 bl[83] br[83] wl[334] vdd gnd cell_6t
Xbit_r335_c83 bl[83] br[83] wl[335] vdd gnd cell_6t
Xbit_r336_c83 bl[83] br[83] wl[336] vdd gnd cell_6t
Xbit_r337_c83 bl[83] br[83] wl[337] vdd gnd cell_6t
Xbit_r338_c83 bl[83] br[83] wl[338] vdd gnd cell_6t
Xbit_r339_c83 bl[83] br[83] wl[339] vdd gnd cell_6t
Xbit_r340_c83 bl[83] br[83] wl[340] vdd gnd cell_6t
Xbit_r341_c83 bl[83] br[83] wl[341] vdd gnd cell_6t
Xbit_r342_c83 bl[83] br[83] wl[342] vdd gnd cell_6t
Xbit_r343_c83 bl[83] br[83] wl[343] vdd gnd cell_6t
Xbit_r344_c83 bl[83] br[83] wl[344] vdd gnd cell_6t
Xbit_r345_c83 bl[83] br[83] wl[345] vdd gnd cell_6t
Xbit_r346_c83 bl[83] br[83] wl[346] vdd gnd cell_6t
Xbit_r347_c83 bl[83] br[83] wl[347] vdd gnd cell_6t
Xbit_r348_c83 bl[83] br[83] wl[348] vdd gnd cell_6t
Xbit_r349_c83 bl[83] br[83] wl[349] vdd gnd cell_6t
Xbit_r350_c83 bl[83] br[83] wl[350] vdd gnd cell_6t
Xbit_r351_c83 bl[83] br[83] wl[351] vdd gnd cell_6t
Xbit_r352_c83 bl[83] br[83] wl[352] vdd gnd cell_6t
Xbit_r353_c83 bl[83] br[83] wl[353] vdd gnd cell_6t
Xbit_r354_c83 bl[83] br[83] wl[354] vdd gnd cell_6t
Xbit_r355_c83 bl[83] br[83] wl[355] vdd gnd cell_6t
Xbit_r356_c83 bl[83] br[83] wl[356] vdd gnd cell_6t
Xbit_r357_c83 bl[83] br[83] wl[357] vdd gnd cell_6t
Xbit_r358_c83 bl[83] br[83] wl[358] vdd gnd cell_6t
Xbit_r359_c83 bl[83] br[83] wl[359] vdd gnd cell_6t
Xbit_r360_c83 bl[83] br[83] wl[360] vdd gnd cell_6t
Xbit_r361_c83 bl[83] br[83] wl[361] vdd gnd cell_6t
Xbit_r362_c83 bl[83] br[83] wl[362] vdd gnd cell_6t
Xbit_r363_c83 bl[83] br[83] wl[363] vdd gnd cell_6t
Xbit_r364_c83 bl[83] br[83] wl[364] vdd gnd cell_6t
Xbit_r365_c83 bl[83] br[83] wl[365] vdd gnd cell_6t
Xbit_r366_c83 bl[83] br[83] wl[366] vdd gnd cell_6t
Xbit_r367_c83 bl[83] br[83] wl[367] vdd gnd cell_6t
Xbit_r368_c83 bl[83] br[83] wl[368] vdd gnd cell_6t
Xbit_r369_c83 bl[83] br[83] wl[369] vdd gnd cell_6t
Xbit_r370_c83 bl[83] br[83] wl[370] vdd gnd cell_6t
Xbit_r371_c83 bl[83] br[83] wl[371] vdd gnd cell_6t
Xbit_r372_c83 bl[83] br[83] wl[372] vdd gnd cell_6t
Xbit_r373_c83 bl[83] br[83] wl[373] vdd gnd cell_6t
Xbit_r374_c83 bl[83] br[83] wl[374] vdd gnd cell_6t
Xbit_r375_c83 bl[83] br[83] wl[375] vdd gnd cell_6t
Xbit_r376_c83 bl[83] br[83] wl[376] vdd gnd cell_6t
Xbit_r377_c83 bl[83] br[83] wl[377] vdd gnd cell_6t
Xbit_r378_c83 bl[83] br[83] wl[378] vdd gnd cell_6t
Xbit_r379_c83 bl[83] br[83] wl[379] vdd gnd cell_6t
Xbit_r380_c83 bl[83] br[83] wl[380] vdd gnd cell_6t
Xbit_r381_c83 bl[83] br[83] wl[381] vdd gnd cell_6t
Xbit_r382_c83 bl[83] br[83] wl[382] vdd gnd cell_6t
Xbit_r383_c83 bl[83] br[83] wl[383] vdd gnd cell_6t
Xbit_r384_c83 bl[83] br[83] wl[384] vdd gnd cell_6t
Xbit_r385_c83 bl[83] br[83] wl[385] vdd gnd cell_6t
Xbit_r386_c83 bl[83] br[83] wl[386] vdd gnd cell_6t
Xbit_r387_c83 bl[83] br[83] wl[387] vdd gnd cell_6t
Xbit_r388_c83 bl[83] br[83] wl[388] vdd gnd cell_6t
Xbit_r389_c83 bl[83] br[83] wl[389] vdd gnd cell_6t
Xbit_r390_c83 bl[83] br[83] wl[390] vdd gnd cell_6t
Xbit_r391_c83 bl[83] br[83] wl[391] vdd gnd cell_6t
Xbit_r392_c83 bl[83] br[83] wl[392] vdd gnd cell_6t
Xbit_r393_c83 bl[83] br[83] wl[393] vdd gnd cell_6t
Xbit_r394_c83 bl[83] br[83] wl[394] vdd gnd cell_6t
Xbit_r395_c83 bl[83] br[83] wl[395] vdd gnd cell_6t
Xbit_r396_c83 bl[83] br[83] wl[396] vdd gnd cell_6t
Xbit_r397_c83 bl[83] br[83] wl[397] vdd gnd cell_6t
Xbit_r398_c83 bl[83] br[83] wl[398] vdd gnd cell_6t
Xbit_r399_c83 bl[83] br[83] wl[399] vdd gnd cell_6t
Xbit_r400_c83 bl[83] br[83] wl[400] vdd gnd cell_6t
Xbit_r401_c83 bl[83] br[83] wl[401] vdd gnd cell_6t
Xbit_r402_c83 bl[83] br[83] wl[402] vdd gnd cell_6t
Xbit_r403_c83 bl[83] br[83] wl[403] vdd gnd cell_6t
Xbit_r404_c83 bl[83] br[83] wl[404] vdd gnd cell_6t
Xbit_r405_c83 bl[83] br[83] wl[405] vdd gnd cell_6t
Xbit_r406_c83 bl[83] br[83] wl[406] vdd gnd cell_6t
Xbit_r407_c83 bl[83] br[83] wl[407] vdd gnd cell_6t
Xbit_r408_c83 bl[83] br[83] wl[408] vdd gnd cell_6t
Xbit_r409_c83 bl[83] br[83] wl[409] vdd gnd cell_6t
Xbit_r410_c83 bl[83] br[83] wl[410] vdd gnd cell_6t
Xbit_r411_c83 bl[83] br[83] wl[411] vdd gnd cell_6t
Xbit_r412_c83 bl[83] br[83] wl[412] vdd gnd cell_6t
Xbit_r413_c83 bl[83] br[83] wl[413] vdd gnd cell_6t
Xbit_r414_c83 bl[83] br[83] wl[414] vdd gnd cell_6t
Xbit_r415_c83 bl[83] br[83] wl[415] vdd gnd cell_6t
Xbit_r416_c83 bl[83] br[83] wl[416] vdd gnd cell_6t
Xbit_r417_c83 bl[83] br[83] wl[417] vdd gnd cell_6t
Xbit_r418_c83 bl[83] br[83] wl[418] vdd gnd cell_6t
Xbit_r419_c83 bl[83] br[83] wl[419] vdd gnd cell_6t
Xbit_r420_c83 bl[83] br[83] wl[420] vdd gnd cell_6t
Xbit_r421_c83 bl[83] br[83] wl[421] vdd gnd cell_6t
Xbit_r422_c83 bl[83] br[83] wl[422] vdd gnd cell_6t
Xbit_r423_c83 bl[83] br[83] wl[423] vdd gnd cell_6t
Xbit_r424_c83 bl[83] br[83] wl[424] vdd gnd cell_6t
Xbit_r425_c83 bl[83] br[83] wl[425] vdd gnd cell_6t
Xbit_r426_c83 bl[83] br[83] wl[426] vdd gnd cell_6t
Xbit_r427_c83 bl[83] br[83] wl[427] vdd gnd cell_6t
Xbit_r428_c83 bl[83] br[83] wl[428] vdd gnd cell_6t
Xbit_r429_c83 bl[83] br[83] wl[429] vdd gnd cell_6t
Xbit_r430_c83 bl[83] br[83] wl[430] vdd gnd cell_6t
Xbit_r431_c83 bl[83] br[83] wl[431] vdd gnd cell_6t
Xbit_r432_c83 bl[83] br[83] wl[432] vdd gnd cell_6t
Xbit_r433_c83 bl[83] br[83] wl[433] vdd gnd cell_6t
Xbit_r434_c83 bl[83] br[83] wl[434] vdd gnd cell_6t
Xbit_r435_c83 bl[83] br[83] wl[435] vdd gnd cell_6t
Xbit_r436_c83 bl[83] br[83] wl[436] vdd gnd cell_6t
Xbit_r437_c83 bl[83] br[83] wl[437] vdd gnd cell_6t
Xbit_r438_c83 bl[83] br[83] wl[438] vdd gnd cell_6t
Xbit_r439_c83 bl[83] br[83] wl[439] vdd gnd cell_6t
Xbit_r440_c83 bl[83] br[83] wl[440] vdd gnd cell_6t
Xbit_r441_c83 bl[83] br[83] wl[441] vdd gnd cell_6t
Xbit_r442_c83 bl[83] br[83] wl[442] vdd gnd cell_6t
Xbit_r443_c83 bl[83] br[83] wl[443] vdd gnd cell_6t
Xbit_r444_c83 bl[83] br[83] wl[444] vdd gnd cell_6t
Xbit_r445_c83 bl[83] br[83] wl[445] vdd gnd cell_6t
Xbit_r446_c83 bl[83] br[83] wl[446] vdd gnd cell_6t
Xbit_r447_c83 bl[83] br[83] wl[447] vdd gnd cell_6t
Xbit_r448_c83 bl[83] br[83] wl[448] vdd gnd cell_6t
Xbit_r449_c83 bl[83] br[83] wl[449] vdd gnd cell_6t
Xbit_r450_c83 bl[83] br[83] wl[450] vdd gnd cell_6t
Xbit_r451_c83 bl[83] br[83] wl[451] vdd gnd cell_6t
Xbit_r452_c83 bl[83] br[83] wl[452] vdd gnd cell_6t
Xbit_r453_c83 bl[83] br[83] wl[453] vdd gnd cell_6t
Xbit_r454_c83 bl[83] br[83] wl[454] vdd gnd cell_6t
Xbit_r455_c83 bl[83] br[83] wl[455] vdd gnd cell_6t
Xbit_r456_c83 bl[83] br[83] wl[456] vdd gnd cell_6t
Xbit_r457_c83 bl[83] br[83] wl[457] vdd gnd cell_6t
Xbit_r458_c83 bl[83] br[83] wl[458] vdd gnd cell_6t
Xbit_r459_c83 bl[83] br[83] wl[459] vdd gnd cell_6t
Xbit_r460_c83 bl[83] br[83] wl[460] vdd gnd cell_6t
Xbit_r461_c83 bl[83] br[83] wl[461] vdd gnd cell_6t
Xbit_r462_c83 bl[83] br[83] wl[462] vdd gnd cell_6t
Xbit_r463_c83 bl[83] br[83] wl[463] vdd gnd cell_6t
Xbit_r464_c83 bl[83] br[83] wl[464] vdd gnd cell_6t
Xbit_r465_c83 bl[83] br[83] wl[465] vdd gnd cell_6t
Xbit_r466_c83 bl[83] br[83] wl[466] vdd gnd cell_6t
Xbit_r467_c83 bl[83] br[83] wl[467] vdd gnd cell_6t
Xbit_r468_c83 bl[83] br[83] wl[468] vdd gnd cell_6t
Xbit_r469_c83 bl[83] br[83] wl[469] vdd gnd cell_6t
Xbit_r470_c83 bl[83] br[83] wl[470] vdd gnd cell_6t
Xbit_r471_c83 bl[83] br[83] wl[471] vdd gnd cell_6t
Xbit_r472_c83 bl[83] br[83] wl[472] vdd gnd cell_6t
Xbit_r473_c83 bl[83] br[83] wl[473] vdd gnd cell_6t
Xbit_r474_c83 bl[83] br[83] wl[474] vdd gnd cell_6t
Xbit_r475_c83 bl[83] br[83] wl[475] vdd gnd cell_6t
Xbit_r476_c83 bl[83] br[83] wl[476] vdd gnd cell_6t
Xbit_r477_c83 bl[83] br[83] wl[477] vdd gnd cell_6t
Xbit_r478_c83 bl[83] br[83] wl[478] vdd gnd cell_6t
Xbit_r479_c83 bl[83] br[83] wl[479] vdd gnd cell_6t
Xbit_r480_c83 bl[83] br[83] wl[480] vdd gnd cell_6t
Xbit_r481_c83 bl[83] br[83] wl[481] vdd gnd cell_6t
Xbit_r482_c83 bl[83] br[83] wl[482] vdd gnd cell_6t
Xbit_r483_c83 bl[83] br[83] wl[483] vdd gnd cell_6t
Xbit_r484_c83 bl[83] br[83] wl[484] vdd gnd cell_6t
Xbit_r485_c83 bl[83] br[83] wl[485] vdd gnd cell_6t
Xbit_r486_c83 bl[83] br[83] wl[486] vdd gnd cell_6t
Xbit_r487_c83 bl[83] br[83] wl[487] vdd gnd cell_6t
Xbit_r488_c83 bl[83] br[83] wl[488] vdd gnd cell_6t
Xbit_r489_c83 bl[83] br[83] wl[489] vdd gnd cell_6t
Xbit_r490_c83 bl[83] br[83] wl[490] vdd gnd cell_6t
Xbit_r491_c83 bl[83] br[83] wl[491] vdd gnd cell_6t
Xbit_r492_c83 bl[83] br[83] wl[492] vdd gnd cell_6t
Xbit_r493_c83 bl[83] br[83] wl[493] vdd gnd cell_6t
Xbit_r494_c83 bl[83] br[83] wl[494] vdd gnd cell_6t
Xbit_r495_c83 bl[83] br[83] wl[495] vdd gnd cell_6t
Xbit_r496_c83 bl[83] br[83] wl[496] vdd gnd cell_6t
Xbit_r497_c83 bl[83] br[83] wl[497] vdd gnd cell_6t
Xbit_r498_c83 bl[83] br[83] wl[498] vdd gnd cell_6t
Xbit_r499_c83 bl[83] br[83] wl[499] vdd gnd cell_6t
Xbit_r500_c83 bl[83] br[83] wl[500] vdd gnd cell_6t
Xbit_r501_c83 bl[83] br[83] wl[501] vdd gnd cell_6t
Xbit_r502_c83 bl[83] br[83] wl[502] vdd gnd cell_6t
Xbit_r503_c83 bl[83] br[83] wl[503] vdd gnd cell_6t
Xbit_r504_c83 bl[83] br[83] wl[504] vdd gnd cell_6t
Xbit_r505_c83 bl[83] br[83] wl[505] vdd gnd cell_6t
Xbit_r506_c83 bl[83] br[83] wl[506] vdd gnd cell_6t
Xbit_r507_c83 bl[83] br[83] wl[507] vdd gnd cell_6t
Xbit_r508_c83 bl[83] br[83] wl[508] vdd gnd cell_6t
Xbit_r509_c83 bl[83] br[83] wl[509] vdd gnd cell_6t
Xbit_r510_c83 bl[83] br[83] wl[510] vdd gnd cell_6t
Xbit_r511_c83 bl[83] br[83] wl[511] vdd gnd cell_6t
Xbit_r0_c84 bl[84] br[84] wl[0] vdd gnd cell_6t
Xbit_r1_c84 bl[84] br[84] wl[1] vdd gnd cell_6t
Xbit_r2_c84 bl[84] br[84] wl[2] vdd gnd cell_6t
Xbit_r3_c84 bl[84] br[84] wl[3] vdd gnd cell_6t
Xbit_r4_c84 bl[84] br[84] wl[4] vdd gnd cell_6t
Xbit_r5_c84 bl[84] br[84] wl[5] vdd gnd cell_6t
Xbit_r6_c84 bl[84] br[84] wl[6] vdd gnd cell_6t
Xbit_r7_c84 bl[84] br[84] wl[7] vdd gnd cell_6t
Xbit_r8_c84 bl[84] br[84] wl[8] vdd gnd cell_6t
Xbit_r9_c84 bl[84] br[84] wl[9] vdd gnd cell_6t
Xbit_r10_c84 bl[84] br[84] wl[10] vdd gnd cell_6t
Xbit_r11_c84 bl[84] br[84] wl[11] vdd gnd cell_6t
Xbit_r12_c84 bl[84] br[84] wl[12] vdd gnd cell_6t
Xbit_r13_c84 bl[84] br[84] wl[13] vdd gnd cell_6t
Xbit_r14_c84 bl[84] br[84] wl[14] vdd gnd cell_6t
Xbit_r15_c84 bl[84] br[84] wl[15] vdd gnd cell_6t
Xbit_r16_c84 bl[84] br[84] wl[16] vdd gnd cell_6t
Xbit_r17_c84 bl[84] br[84] wl[17] vdd gnd cell_6t
Xbit_r18_c84 bl[84] br[84] wl[18] vdd gnd cell_6t
Xbit_r19_c84 bl[84] br[84] wl[19] vdd gnd cell_6t
Xbit_r20_c84 bl[84] br[84] wl[20] vdd gnd cell_6t
Xbit_r21_c84 bl[84] br[84] wl[21] vdd gnd cell_6t
Xbit_r22_c84 bl[84] br[84] wl[22] vdd gnd cell_6t
Xbit_r23_c84 bl[84] br[84] wl[23] vdd gnd cell_6t
Xbit_r24_c84 bl[84] br[84] wl[24] vdd gnd cell_6t
Xbit_r25_c84 bl[84] br[84] wl[25] vdd gnd cell_6t
Xbit_r26_c84 bl[84] br[84] wl[26] vdd gnd cell_6t
Xbit_r27_c84 bl[84] br[84] wl[27] vdd gnd cell_6t
Xbit_r28_c84 bl[84] br[84] wl[28] vdd gnd cell_6t
Xbit_r29_c84 bl[84] br[84] wl[29] vdd gnd cell_6t
Xbit_r30_c84 bl[84] br[84] wl[30] vdd gnd cell_6t
Xbit_r31_c84 bl[84] br[84] wl[31] vdd gnd cell_6t
Xbit_r32_c84 bl[84] br[84] wl[32] vdd gnd cell_6t
Xbit_r33_c84 bl[84] br[84] wl[33] vdd gnd cell_6t
Xbit_r34_c84 bl[84] br[84] wl[34] vdd gnd cell_6t
Xbit_r35_c84 bl[84] br[84] wl[35] vdd gnd cell_6t
Xbit_r36_c84 bl[84] br[84] wl[36] vdd gnd cell_6t
Xbit_r37_c84 bl[84] br[84] wl[37] vdd gnd cell_6t
Xbit_r38_c84 bl[84] br[84] wl[38] vdd gnd cell_6t
Xbit_r39_c84 bl[84] br[84] wl[39] vdd gnd cell_6t
Xbit_r40_c84 bl[84] br[84] wl[40] vdd gnd cell_6t
Xbit_r41_c84 bl[84] br[84] wl[41] vdd gnd cell_6t
Xbit_r42_c84 bl[84] br[84] wl[42] vdd gnd cell_6t
Xbit_r43_c84 bl[84] br[84] wl[43] vdd gnd cell_6t
Xbit_r44_c84 bl[84] br[84] wl[44] vdd gnd cell_6t
Xbit_r45_c84 bl[84] br[84] wl[45] vdd gnd cell_6t
Xbit_r46_c84 bl[84] br[84] wl[46] vdd gnd cell_6t
Xbit_r47_c84 bl[84] br[84] wl[47] vdd gnd cell_6t
Xbit_r48_c84 bl[84] br[84] wl[48] vdd gnd cell_6t
Xbit_r49_c84 bl[84] br[84] wl[49] vdd gnd cell_6t
Xbit_r50_c84 bl[84] br[84] wl[50] vdd gnd cell_6t
Xbit_r51_c84 bl[84] br[84] wl[51] vdd gnd cell_6t
Xbit_r52_c84 bl[84] br[84] wl[52] vdd gnd cell_6t
Xbit_r53_c84 bl[84] br[84] wl[53] vdd gnd cell_6t
Xbit_r54_c84 bl[84] br[84] wl[54] vdd gnd cell_6t
Xbit_r55_c84 bl[84] br[84] wl[55] vdd gnd cell_6t
Xbit_r56_c84 bl[84] br[84] wl[56] vdd gnd cell_6t
Xbit_r57_c84 bl[84] br[84] wl[57] vdd gnd cell_6t
Xbit_r58_c84 bl[84] br[84] wl[58] vdd gnd cell_6t
Xbit_r59_c84 bl[84] br[84] wl[59] vdd gnd cell_6t
Xbit_r60_c84 bl[84] br[84] wl[60] vdd gnd cell_6t
Xbit_r61_c84 bl[84] br[84] wl[61] vdd gnd cell_6t
Xbit_r62_c84 bl[84] br[84] wl[62] vdd gnd cell_6t
Xbit_r63_c84 bl[84] br[84] wl[63] vdd gnd cell_6t
Xbit_r64_c84 bl[84] br[84] wl[64] vdd gnd cell_6t
Xbit_r65_c84 bl[84] br[84] wl[65] vdd gnd cell_6t
Xbit_r66_c84 bl[84] br[84] wl[66] vdd gnd cell_6t
Xbit_r67_c84 bl[84] br[84] wl[67] vdd gnd cell_6t
Xbit_r68_c84 bl[84] br[84] wl[68] vdd gnd cell_6t
Xbit_r69_c84 bl[84] br[84] wl[69] vdd gnd cell_6t
Xbit_r70_c84 bl[84] br[84] wl[70] vdd gnd cell_6t
Xbit_r71_c84 bl[84] br[84] wl[71] vdd gnd cell_6t
Xbit_r72_c84 bl[84] br[84] wl[72] vdd gnd cell_6t
Xbit_r73_c84 bl[84] br[84] wl[73] vdd gnd cell_6t
Xbit_r74_c84 bl[84] br[84] wl[74] vdd gnd cell_6t
Xbit_r75_c84 bl[84] br[84] wl[75] vdd gnd cell_6t
Xbit_r76_c84 bl[84] br[84] wl[76] vdd gnd cell_6t
Xbit_r77_c84 bl[84] br[84] wl[77] vdd gnd cell_6t
Xbit_r78_c84 bl[84] br[84] wl[78] vdd gnd cell_6t
Xbit_r79_c84 bl[84] br[84] wl[79] vdd gnd cell_6t
Xbit_r80_c84 bl[84] br[84] wl[80] vdd gnd cell_6t
Xbit_r81_c84 bl[84] br[84] wl[81] vdd gnd cell_6t
Xbit_r82_c84 bl[84] br[84] wl[82] vdd gnd cell_6t
Xbit_r83_c84 bl[84] br[84] wl[83] vdd gnd cell_6t
Xbit_r84_c84 bl[84] br[84] wl[84] vdd gnd cell_6t
Xbit_r85_c84 bl[84] br[84] wl[85] vdd gnd cell_6t
Xbit_r86_c84 bl[84] br[84] wl[86] vdd gnd cell_6t
Xbit_r87_c84 bl[84] br[84] wl[87] vdd gnd cell_6t
Xbit_r88_c84 bl[84] br[84] wl[88] vdd gnd cell_6t
Xbit_r89_c84 bl[84] br[84] wl[89] vdd gnd cell_6t
Xbit_r90_c84 bl[84] br[84] wl[90] vdd gnd cell_6t
Xbit_r91_c84 bl[84] br[84] wl[91] vdd gnd cell_6t
Xbit_r92_c84 bl[84] br[84] wl[92] vdd gnd cell_6t
Xbit_r93_c84 bl[84] br[84] wl[93] vdd gnd cell_6t
Xbit_r94_c84 bl[84] br[84] wl[94] vdd gnd cell_6t
Xbit_r95_c84 bl[84] br[84] wl[95] vdd gnd cell_6t
Xbit_r96_c84 bl[84] br[84] wl[96] vdd gnd cell_6t
Xbit_r97_c84 bl[84] br[84] wl[97] vdd gnd cell_6t
Xbit_r98_c84 bl[84] br[84] wl[98] vdd gnd cell_6t
Xbit_r99_c84 bl[84] br[84] wl[99] vdd gnd cell_6t
Xbit_r100_c84 bl[84] br[84] wl[100] vdd gnd cell_6t
Xbit_r101_c84 bl[84] br[84] wl[101] vdd gnd cell_6t
Xbit_r102_c84 bl[84] br[84] wl[102] vdd gnd cell_6t
Xbit_r103_c84 bl[84] br[84] wl[103] vdd gnd cell_6t
Xbit_r104_c84 bl[84] br[84] wl[104] vdd gnd cell_6t
Xbit_r105_c84 bl[84] br[84] wl[105] vdd gnd cell_6t
Xbit_r106_c84 bl[84] br[84] wl[106] vdd gnd cell_6t
Xbit_r107_c84 bl[84] br[84] wl[107] vdd gnd cell_6t
Xbit_r108_c84 bl[84] br[84] wl[108] vdd gnd cell_6t
Xbit_r109_c84 bl[84] br[84] wl[109] vdd gnd cell_6t
Xbit_r110_c84 bl[84] br[84] wl[110] vdd gnd cell_6t
Xbit_r111_c84 bl[84] br[84] wl[111] vdd gnd cell_6t
Xbit_r112_c84 bl[84] br[84] wl[112] vdd gnd cell_6t
Xbit_r113_c84 bl[84] br[84] wl[113] vdd gnd cell_6t
Xbit_r114_c84 bl[84] br[84] wl[114] vdd gnd cell_6t
Xbit_r115_c84 bl[84] br[84] wl[115] vdd gnd cell_6t
Xbit_r116_c84 bl[84] br[84] wl[116] vdd gnd cell_6t
Xbit_r117_c84 bl[84] br[84] wl[117] vdd gnd cell_6t
Xbit_r118_c84 bl[84] br[84] wl[118] vdd gnd cell_6t
Xbit_r119_c84 bl[84] br[84] wl[119] vdd gnd cell_6t
Xbit_r120_c84 bl[84] br[84] wl[120] vdd gnd cell_6t
Xbit_r121_c84 bl[84] br[84] wl[121] vdd gnd cell_6t
Xbit_r122_c84 bl[84] br[84] wl[122] vdd gnd cell_6t
Xbit_r123_c84 bl[84] br[84] wl[123] vdd gnd cell_6t
Xbit_r124_c84 bl[84] br[84] wl[124] vdd gnd cell_6t
Xbit_r125_c84 bl[84] br[84] wl[125] vdd gnd cell_6t
Xbit_r126_c84 bl[84] br[84] wl[126] vdd gnd cell_6t
Xbit_r127_c84 bl[84] br[84] wl[127] vdd gnd cell_6t
Xbit_r128_c84 bl[84] br[84] wl[128] vdd gnd cell_6t
Xbit_r129_c84 bl[84] br[84] wl[129] vdd gnd cell_6t
Xbit_r130_c84 bl[84] br[84] wl[130] vdd gnd cell_6t
Xbit_r131_c84 bl[84] br[84] wl[131] vdd gnd cell_6t
Xbit_r132_c84 bl[84] br[84] wl[132] vdd gnd cell_6t
Xbit_r133_c84 bl[84] br[84] wl[133] vdd gnd cell_6t
Xbit_r134_c84 bl[84] br[84] wl[134] vdd gnd cell_6t
Xbit_r135_c84 bl[84] br[84] wl[135] vdd gnd cell_6t
Xbit_r136_c84 bl[84] br[84] wl[136] vdd gnd cell_6t
Xbit_r137_c84 bl[84] br[84] wl[137] vdd gnd cell_6t
Xbit_r138_c84 bl[84] br[84] wl[138] vdd gnd cell_6t
Xbit_r139_c84 bl[84] br[84] wl[139] vdd gnd cell_6t
Xbit_r140_c84 bl[84] br[84] wl[140] vdd gnd cell_6t
Xbit_r141_c84 bl[84] br[84] wl[141] vdd gnd cell_6t
Xbit_r142_c84 bl[84] br[84] wl[142] vdd gnd cell_6t
Xbit_r143_c84 bl[84] br[84] wl[143] vdd gnd cell_6t
Xbit_r144_c84 bl[84] br[84] wl[144] vdd gnd cell_6t
Xbit_r145_c84 bl[84] br[84] wl[145] vdd gnd cell_6t
Xbit_r146_c84 bl[84] br[84] wl[146] vdd gnd cell_6t
Xbit_r147_c84 bl[84] br[84] wl[147] vdd gnd cell_6t
Xbit_r148_c84 bl[84] br[84] wl[148] vdd gnd cell_6t
Xbit_r149_c84 bl[84] br[84] wl[149] vdd gnd cell_6t
Xbit_r150_c84 bl[84] br[84] wl[150] vdd gnd cell_6t
Xbit_r151_c84 bl[84] br[84] wl[151] vdd gnd cell_6t
Xbit_r152_c84 bl[84] br[84] wl[152] vdd gnd cell_6t
Xbit_r153_c84 bl[84] br[84] wl[153] vdd gnd cell_6t
Xbit_r154_c84 bl[84] br[84] wl[154] vdd gnd cell_6t
Xbit_r155_c84 bl[84] br[84] wl[155] vdd gnd cell_6t
Xbit_r156_c84 bl[84] br[84] wl[156] vdd gnd cell_6t
Xbit_r157_c84 bl[84] br[84] wl[157] vdd gnd cell_6t
Xbit_r158_c84 bl[84] br[84] wl[158] vdd gnd cell_6t
Xbit_r159_c84 bl[84] br[84] wl[159] vdd gnd cell_6t
Xbit_r160_c84 bl[84] br[84] wl[160] vdd gnd cell_6t
Xbit_r161_c84 bl[84] br[84] wl[161] vdd gnd cell_6t
Xbit_r162_c84 bl[84] br[84] wl[162] vdd gnd cell_6t
Xbit_r163_c84 bl[84] br[84] wl[163] vdd gnd cell_6t
Xbit_r164_c84 bl[84] br[84] wl[164] vdd gnd cell_6t
Xbit_r165_c84 bl[84] br[84] wl[165] vdd gnd cell_6t
Xbit_r166_c84 bl[84] br[84] wl[166] vdd gnd cell_6t
Xbit_r167_c84 bl[84] br[84] wl[167] vdd gnd cell_6t
Xbit_r168_c84 bl[84] br[84] wl[168] vdd gnd cell_6t
Xbit_r169_c84 bl[84] br[84] wl[169] vdd gnd cell_6t
Xbit_r170_c84 bl[84] br[84] wl[170] vdd gnd cell_6t
Xbit_r171_c84 bl[84] br[84] wl[171] vdd gnd cell_6t
Xbit_r172_c84 bl[84] br[84] wl[172] vdd gnd cell_6t
Xbit_r173_c84 bl[84] br[84] wl[173] vdd gnd cell_6t
Xbit_r174_c84 bl[84] br[84] wl[174] vdd gnd cell_6t
Xbit_r175_c84 bl[84] br[84] wl[175] vdd gnd cell_6t
Xbit_r176_c84 bl[84] br[84] wl[176] vdd gnd cell_6t
Xbit_r177_c84 bl[84] br[84] wl[177] vdd gnd cell_6t
Xbit_r178_c84 bl[84] br[84] wl[178] vdd gnd cell_6t
Xbit_r179_c84 bl[84] br[84] wl[179] vdd gnd cell_6t
Xbit_r180_c84 bl[84] br[84] wl[180] vdd gnd cell_6t
Xbit_r181_c84 bl[84] br[84] wl[181] vdd gnd cell_6t
Xbit_r182_c84 bl[84] br[84] wl[182] vdd gnd cell_6t
Xbit_r183_c84 bl[84] br[84] wl[183] vdd gnd cell_6t
Xbit_r184_c84 bl[84] br[84] wl[184] vdd gnd cell_6t
Xbit_r185_c84 bl[84] br[84] wl[185] vdd gnd cell_6t
Xbit_r186_c84 bl[84] br[84] wl[186] vdd gnd cell_6t
Xbit_r187_c84 bl[84] br[84] wl[187] vdd gnd cell_6t
Xbit_r188_c84 bl[84] br[84] wl[188] vdd gnd cell_6t
Xbit_r189_c84 bl[84] br[84] wl[189] vdd gnd cell_6t
Xbit_r190_c84 bl[84] br[84] wl[190] vdd gnd cell_6t
Xbit_r191_c84 bl[84] br[84] wl[191] vdd gnd cell_6t
Xbit_r192_c84 bl[84] br[84] wl[192] vdd gnd cell_6t
Xbit_r193_c84 bl[84] br[84] wl[193] vdd gnd cell_6t
Xbit_r194_c84 bl[84] br[84] wl[194] vdd gnd cell_6t
Xbit_r195_c84 bl[84] br[84] wl[195] vdd gnd cell_6t
Xbit_r196_c84 bl[84] br[84] wl[196] vdd gnd cell_6t
Xbit_r197_c84 bl[84] br[84] wl[197] vdd gnd cell_6t
Xbit_r198_c84 bl[84] br[84] wl[198] vdd gnd cell_6t
Xbit_r199_c84 bl[84] br[84] wl[199] vdd gnd cell_6t
Xbit_r200_c84 bl[84] br[84] wl[200] vdd gnd cell_6t
Xbit_r201_c84 bl[84] br[84] wl[201] vdd gnd cell_6t
Xbit_r202_c84 bl[84] br[84] wl[202] vdd gnd cell_6t
Xbit_r203_c84 bl[84] br[84] wl[203] vdd gnd cell_6t
Xbit_r204_c84 bl[84] br[84] wl[204] vdd gnd cell_6t
Xbit_r205_c84 bl[84] br[84] wl[205] vdd gnd cell_6t
Xbit_r206_c84 bl[84] br[84] wl[206] vdd gnd cell_6t
Xbit_r207_c84 bl[84] br[84] wl[207] vdd gnd cell_6t
Xbit_r208_c84 bl[84] br[84] wl[208] vdd gnd cell_6t
Xbit_r209_c84 bl[84] br[84] wl[209] vdd gnd cell_6t
Xbit_r210_c84 bl[84] br[84] wl[210] vdd gnd cell_6t
Xbit_r211_c84 bl[84] br[84] wl[211] vdd gnd cell_6t
Xbit_r212_c84 bl[84] br[84] wl[212] vdd gnd cell_6t
Xbit_r213_c84 bl[84] br[84] wl[213] vdd gnd cell_6t
Xbit_r214_c84 bl[84] br[84] wl[214] vdd gnd cell_6t
Xbit_r215_c84 bl[84] br[84] wl[215] vdd gnd cell_6t
Xbit_r216_c84 bl[84] br[84] wl[216] vdd gnd cell_6t
Xbit_r217_c84 bl[84] br[84] wl[217] vdd gnd cell_6t
Xbit_r218_c84 bl[84] br[84] wl[218] vdd gnd cell_6t
Xbit_r219_c84 bl[84] br[84] wl[219] vdd gnd cell_6t
Xbit_r220_c84 bl[84] br[84] wl[220] vdd gnd cell_6t
Xbit_r221_c84 bl[84] br[84] wl[221] vdd gnd cell_6t
Xbit_r222_c84 bl[84] br[84] wl[222] vdd gnd cell_6t
Xbit_r223_c84 bl[84] br[84] wl[223] vdd gnd cell_6t
Xbit_r224_c84 bl[84] br[84] wl[224] vdd gnd cell_6t
Xbit_r225_c84 bl[84] br[84] wl[225] vdd gnd cell_6t
Xbit_r226_c84 bl[84] br[84] wl[226] vdd gnd cell_6t
Xbit_r227_c84 bl[84] br[84] wl[227] vdd gnd cell_6t
Xbit_r228_c84 bl[84] br[84] wl[228] vdd gnd cell_6t
Xbit_r229_c84 bl[84] br[84] wl[229] vdd gnd cell_6t
Xbit_r230_c84 bl[84] br[84] wl[230] vdd gnd cell_6t
Xbit_r231_c84 bl[84] br[84] wl[231] vdd gnd cell_6t
Xbit_r232_c84 bl[84] br[84] wl[232] vdd gnd cell_6t
Xbit_r233_c84 bl[84] br[84] wl[233] vdd gnd cell_6t
Xbit_r234_c84 bl[84] br[84] wl[234] vdd gnd cell_6t
Xbit_r235_c84 bl[84] br[84] wl[235] vdd gnd cell_6t
Xbit_r236_c84 bl[84] br[84] wl[236] vdd gnd cell_6t
Xbit_r237_c84 bl[84] br[84] wl[237] vdd gnd cell_6t
Xbit_r238_c84 bl[84] br[84] wl[238] vdd gnd cell_6t
Xbit_r239_c84 bl[84] br[84] wl[239] vdd gnd cell_6t
Xbit_r240_c84 bl[84] br[84] wl[240] vdd gnd cell_6t
Xbit_r241_c84 bl[84] br[84] wl[241] vdd gnd cell_6t
Xbit_r242_c84 bl[84] br[84] wl[242] vdd gnd cell_6t
Xbit_r243_c84 bl[84] br[84] wl[243] vdd gnd cell_6t
Xbit_r244_c84 bl[84] br[84] wl[244] vdd gnd cell_6t
Xbit_r245_c84 bl[84] br[84] wl[245] vdd gnd cell_6t
Xbit_r246_c84 bl[84] br[84] wl[246] vdd gnd cell_6t
Xbit_r247_c84 bl[84] br[84] wl[247] vdd gnd cell_6t
Xbit_r248_c84 bl[84] br[84] wl[248] vdd gnd cell_6t
Xbit_r249_c84 bl[84] br[84] wl[249] vdd gnd cell_6t
Xbit_r250_c84 bl[84] br[84] wl[250] vdd gnd cell_6t
Xbit_r251_c84 bl[84] br[84] wl[251] vdd gnd cell_6t
Xbit_r252_c84 bl[84] br[84] wl[252] vdd gnd cell_6t
Xbit_r253_c84 bl[84] br[84] wl[253] vdd gnd cell_6t
Xbit_r254_c84 bl[84] br[84] wl[254] vdd gnd cell_6t
Xbit_r255_c84 bl[84] br[84] wl[255] vdd gnd cell_6t
Xbit_r256_c84 bl[84] br[84] wl[256] vdd gnd cell_6t
Xbit_r257_c84 bl[84] br[84] wl[257] vdd gnd cell_6t
Xbit_r258_c84 bl[84] br[84] wl[258] vdd gnd cell_6t
Xbit_r259_c84 bl[84] br[84] wl[259] vdd gnd cell_6t
Xbit_r260_c84 bl[84] br[84] wl[260] vdd gnd cell_6t
Xbit_r261_c84 bl[84] br[84] wl[261] vdd gnd cell_6t
Xbit_r262_c84 bl[84] br[84] wl[262] vdd gnd cell_6t
Xbit_r263_c84 bl[84] br[84] wl[263] vdd gnd cell_6t
Xbit_r264_c84 bl[84] br[84] wl[264] vdd gnd cell_6t
Xbit_r265_c84 bl[84] br[84] wl[265] vdd gnd cell_6t
Xbit_r266_c84 bl[84] br[84] wl[266] vdd gnd cell_6t
Xbit_r267_c84 bl[84] br[84] wl[267] vdd gnd cell_6t
Xbit_r268_c84 bl[84] br[84] wl[268] vdd gnd cell_6t
Xbit_r269_c84 bl[84] br[84] wl[269] vdd gnd cell_6t
Xbit_r270_c84 bl[84] br[84] wl[270] vdd gnd cell_6t
Xbit_r271_c84 bl[84] br[84] wl[271] vdd gnd cell_6t
Xbit_r272_c84 bl[84] br[84] wl[272] vdd gnd cell_6t
Xbit_r273_c84 bl[84] br[84] wl[273] vdd gnd cell_6t
Xbit_r274_c84 bl[84] br[84] wl[274] vdd gnd cell_6t
Xbit_r275_c84 bl[84] br[84] wl[275] vdd gnd cell_6t
Xbit_r276_c84 bl[84] br[84] wl[276] vdd gnd cell_6t
Xbit_r277_c84 bl[84] br[84] wl[277] vdd gnd cell_6t
Xbit_r278_c84 bl[84] br[84] wl[278] vdd gnd cell_6t
Xbit_r279_c84 bl[84] br[84] wl[279] vdd gnd cell_6t
Xbit_r280_c84 bl[84] br[84] wl[280] vdd gnd cell_6t
Xbit_r281_c84 bl[84] br[84] wl[281] vdd gnd cell_6t
Xbit_r282_c84 bl[84] br[84] wl[282] vdd gnd cell_6t
Xbit_r283_c84 bl[84] br[84] wl[283] vdd gnd cell_6t
Xbit_r284_c84 bl[84] br[84] wl[284] vdd gnd cell_6t
Xbit_r285_c84 bl[84] br[84] wl[285] vdd gnd cell_6t
Xbit_r286_c84 bl[84] br[84] wl[286] vdd gnd cell_6t
Xbit_r287_c84 bl[84] br[84] wl[287] vdd gnd cell_6t
Xbit_r288_c84 bl[84] br[84] wl[288] vdd gnd cell_6t
Xbit_r289_c84 bl[84] br[84] wl[289] vdd gnd cell_6t
Xbit_r290_c84 bl[84] br[84] wl[290] vdd gnd cell_6t
Xbit_r291_c84 bl[84] br[84] wl[291] vdd gnd cell_6t
Xbit_r292_c84 bl[84] br[84] wl[292] vdd gnd cell_6t
Xbit_r293_c84 bl[84] br[84] wl[293] vdd gnd cell_6t
Xbit_r294_c84 bl[84] br[84] wl[294] vdd gnd cell_6t
Xbit_r295_c84 bl[84] br[84] wl[295] vdd gnd cell_6t
Xbit_r296_c84 bl[84] br[84] wl[296] vdd gnd cell_6t
Xbit_r297_c84 bl[84] br[84] wl[297] vdd gnd cell_6t
Xbit_r298_c84 bl[84] br[84] wl[298] vdd gnd cell_6t
Xbit_r299_c84 bl[84] br[84] wl[299] vdd gnd cell_6t
Xbit_r300_c84 bl[84] br[84] wl[300] vdd gnd cell_6t
Xbit_r301_c84 bl[84] br[84] wl[301] vdd gnd cell_6t
Xbit_r302_c84 bl[84] br[84] wl[302] vdd gnd cell_6t
Xbit_r303_c84 bl[84] br[84] wl[303] vdd gnd cell_6t
Xbit_r304_c84 bl[84] br[84] wl[304] vdd gnd cell_6t
Xbit_r305_c84 bl[84] br[84] wl[305] vdd gnd cell_6t
Xbit_r306_c84 bl[84] br[84] wl[306] vdd gnd cell_6t
Xbit_r307_c84 bl[84] br[84] wl[307] vdd gnd cell_6t
Xbit_r308_c84 bl[84] br[84] wl[308] vdd gnd cell_6t
Xbit_r309_c84 bl[84] br[84] wl[309] vdd gnd cell_6t
Xbit_r310_c84 bl[84] br[84] wl[310] vdd gnd cell_6t
Xbit_r311_c84 bl[84] br[84] wl[311] vdd gnd cell_6t
Xbit_r312_c84 bl[84] br[84] wl[312] vdd gnd cell_6t
Xbit_r313_c84 bl[84] br[84] wl[313] vdd gnd cell_6t
Xbit_r314_c84 bl[84] br[84] wl[314] vdd gnd cell_6t
Xbit_r315_c84 bl[84] br[84] wl[315] vdd gnd cell_6t
Xbit_r316_c84 bl[84] br[84] wl[316] vdd gnd cell_6t
Xbit_r317_c84 bl[84] br[84] wl[317] vdd gnd cell_6t
Xbit_r318_c84 bl[84] br[84] wl[318] vdd gnd cell_6t
Xbit_r319_c84 bl[84] br[84] wl[319] vdd gnd cell_6t
Xbit_r320_c84 bl[84] br[84] wl[320] vdd gnd cell_6t
Xbit_r321_c84 bl[84] br[84] wl[321] vdd gnd cell_6t
Xbit_r322_c84 bl[84] br[84] wl[322] vdd gnd cell_6t
Xbit_r323_c84 bl[84] br[84] wl[323] vdd gnd cell_6t
Xbit_r324_c84 bl[84] br[84] wl[324] vdd gnd cell_6t
Xbit_r325_c84 bl[84] br[84] wl[325] vdd gnd cell_6t
Xbit_r326_c84 bl[84] br[84] wl[326] vdd gnd cell_6t
Xbit_r327_c84 bl[84] br[84] wl[327] vdd gnd cell_6t
Xbit_r328_c84 bl[84] br[84] wl[328] vdd gnd cell_6t
Xbit_r329_c84 bl[84] br[84] wl[329] vdd gnd cell_6t
Xbit_r330_c84 bl[84] br[84] wl[330] vdd gnd cell_6t
Xbit_r331_c84 bl[84] br[84] wl[331] vdd gnd cell_6t
Xbit_r332_c84 bl[84] br[84] wl[332] vdd gnd cell_6t
Xbit_r333_c84 bl[84] br[84] wl[333] vdd gnd cell_6t
Xbit_r334_c84 bl[84] br[84] wl[334] vdd gnd cell_6t
Xbit_r335_c84 bl[84] br[84] wl[335] vdd gnd cell_6t
Xbit_r336_c84 bl[84] br[84] wl[336] vdd gnd cell_6t
Xbit_r337_c84 bl[84] br[84] wl[337] vdd gnd cell_6t
Xbit_r338_c84 bl[84] br[84] wl[338] vdd gnd cell_6t
Xbit_r339_c84 bl[84] br[84] wl[339] vdd gnd cell_6t
Xbit_r340_c84 bl[84] br[84] wl[340] vdd gnd cell_6t
Xbit_r341_c84 bl[84] br[84] wl[341] vdd gnd cell_6t
Xbit_r342_c84 bl[84] br[84] wl[342] vdd gnd cell_6t
Xbit_r343_c84 bl[84] br[84] wl[343] vdd gnd cell_6t
Xbit_r344_c84 bl[84] br[84] wl[344] vdd gnd cell_6t
Xbit_r345_c84 bl[84] br[84] wl[345] vdd gnd cell_6t
Xbit_r346_c84 bl[84] br[84] wl[346] vdd gnd cell_6t
Xbit_r347_c84 bl[84] br[84] wl[347] vdd gnd cell_6t
Xbit_r348_c84 bl[84] br[84] wl[348] vdd gnd cell_6t
Xbit_r349_c84 bl[84] br[84] wl[349] vdd gnd cell_6t
Xbit_r350_c84 bl[84] br[84] wl[350] vdd gnd cell_6t
Xbit_r351_c84 bl[84] br[84] wl[351] vdd gnd cell_6t
Xbit_r352_c84 bl[84] br[84] wl[352] vdd gnd cell_6t
Xbit_r353_c84 bl[84] br[84] wl[353] vdd gnd cell_6t
Xbit_r354_c84 bl[84] br[84] wl[354] vdd gnd cell_6t
Xbit_r355_c84 bl[84] br[84] wl[355] vdd gnd cell_6t
Xbit_r356_c84 bl[84] br[84] wl[356] vdd gnd cell_6t
Xbit_r357_c84 bl[84] br[84] wl[357] vdd gnd cell_6t
Xbit_r358_c84 bl[84] br[84] wl[358] vdd gnd cell_6t
Xbit_r359_c84 bl[84] br[84] wl[359] vdd gnd cell_6t
Xbit_r360_c84 bl[84] br[84] wl[360] vdd gnd cell_6t
Xbit_r361_c84 bl[84] br[84] wl[361] vdd gnd cell_6t
Xbit_r362_c84 bl[84] br[84] wl[362] vdd gnd cell_6t
Xbit_r363_c84 bl[84] br[84] wl[363] vdd gnd cell_6t
Xbit_r364_c84 bl[84] br[84] wl[364] vdd gnd cell_6t
Xbit_r365_c84 bl[84] br[84] wl[365] vdd gnd cell_6t
Xbit_r366_c84 bl[84] br[84] wl[366] vdd gnd cell_6t
Xbit_r367_c84 bl[84] br[84] wl[367] vdd gnd cell_6t
Xbit_r368_c84 bl[84] br[84] wl[368] vdd gnd cell_6t
Xbit_r369_c84 bl[84] br[84] wl[369] vdd gnd cell_6t
Xbit_r370_c84 bl[84] br[84] wl[370] vdd gnd cell_6t
Xbit_r371_c84 bl[84] br[84] wl[371] vdd gnd cell_6t
Xbit_r372_c84 bl[84] br[84] wl[372] vdd gnd cell_6t
Xbit_r373_c84 bl[84] br[84] wl[373] vdd gnd cell_6t
Xbit_r374_c84 bl[84] br[84] wl[374] vdd gnd cell_6t
Xbit_r375_c84 bl[84] br[84] wl[375] vdd gnd cell_6t
Xbit_r376_c84 bl[84] br[84] wl[376] vdd gnd cell_6t
Xbit_r377_c84 bl[84] br[84] wl[377] vdd gnd cell_6t
Xbit_r378_c84 bl[84] br[84] wl[378] vdd gnd cell_6t
Xbit_r379_c84 bl[84] br[84] wl[379] vdd gnd cell_6t
Xbit_r380_c84 bl[84] br[84] wl[380] vdd gnd cell_6t
Xbit_r381_c84 bl[84] br[84] wl[381] vdd gnd cell_6t
Xbit_r382_c84 bl[84] br[84] wl[382] vdd gnd cell_6t
Xbit_r383_c84 bl[84] br[84] wl[383] vdd gnd cell_6t
Xbit_r384_c84 bl[84] br[84] wl[384] vdd gnd cell_6t
Xbit_r385_c84 bl[84] br[84] wl[385] vdd gnd cell_6t
Xbit_r386_c84 bl[84] br[84] wl[386] vdd gnd cell_6t
Xbit_r387_c84 bl[84] br[84] wl[387] vdd gnd cell_6t
Xbit_r388_c84 bl[84] br[84] wl[388] vdd gnd cell_6t
Xbit_r389_c84 bl[84] br[84] wl[389] vdd gnd cell_6t
Xbit_r390_c84 bl[84] br[84] wl[390] vdd gnd cell_6t
Xbit_r391_c84 bl[84] br[84] wl[391] vdd gnd cell_6t
Xbit_r392_c84 bl[84] br[84] wl[392] vdd gnd cell_6t
Xbit_r393_c84 bl[84] br[84] wl[393] vdd gnd cell_6t
Xbit_r394_c84 bl[84] br[84] wl[394] vdd gnd cell_6t
Xbit_r395_c84 bl[84] br[84] wl[395] vdd gnd cell_6t
Xbit_r396_c84 bl[84] br[84] wl[396] vdd gnd cell_6t
Xbit_r397_c84 bl[84] br[84] wl[397] vdd gnd cell_6t
Xbit_r398_c84 bl[84] br[84] wl[398] vdd gnd cell_6t
Xbit_r399_c84 bl[84] br[84] wl[399] vdd gnd cell_6t
Xbit_r400_c84 bl[84] br[84] wl[400] vdd gnd cell_6t
Xbit_r401_c84 bl[84] br[84] wl[401] vdd gnd cell_6t
Xbit_r402_c84 bl[84] br[84] wl[402] vdd gnd cell_6t
Xbit_r403_c84 bl[84] br[84] wl[403] vdd gnd cell_6t
Xbit_r404_c84 bl[84] br[84] wl[404] vdd gnd cell_6t
Xbit_r405_c84 bl[84] br[84] wl[405] vdd gnd cell_6t
Xbit_r406_c84 bl[84] br[84] wl[406] vdd gnd cell_6t
Xbit_r407_c84 bl[84] br[84] wl[407] vdd gnd cell_6t
Xbit_r408_c84 bl[84] br[84] wl[408] vdd gnd cell_6t
Xbit_r409_c84 bl[84] br[84] wl[409] vdd gnd cell_6t
Xbit_r410_c84 bl[84] br[84] wl[410] vdd gnd cell_6t
Xbit_r411_c84 bl[84] br[84] wl[411] vdd gnd cell_6t
Xbit_r412_c84 bl[84] br[84] wl[412] vdd gnd cell_6t
Xbit_r413_c84 bl[84] br[84] wl[413] vdd gnd cell_6t
Xbit_r414_c84 bl[84] br[84] wl[414] vdd gnd cell_6t
Xbit_r415_c84 bl[84] br[84] wl[415] vdd gnd cell_6t
Xbit_r416_c84 bl[84] br[84] wl[416] vdd gnd cell_6t
Xbit_r417_c84 bl[84] br[84] wl[417] vdd gnd cell_6t
Xbit_r418_c84 bl[84] br[84] wl[418] vdd gnd cell_6t
Xbit_r419_c84 bl[84] br[84] wl[419] vdd gnd cell_6t
Xbit_r420_c84 bl[84] br[84] wl[420] vdd gnd cell_6t
Xbit_r421_c84 bl[84] br[84] wl[421] vdd gnd cell_6t
Xbit_r422_c84 bl[84] br[84] wl[422] vdd gnd cell_6t
Xbit_r423_c84 bl[84] br[84] wl[423] vdd gnd cell_6t
Xbit_r424_c84 bl[84] br[84] wl[424] vdd gnd cell_6t
Xbit_r425_c84 bl[84] br[84] wl[425] vdd gnd cell_6t
Xbit_r426_c84 bl[84] br[84] wl[426] vdd gnd cell_6t
Xbit_r427_c84 bl[84] br[84] wl[427] vdd gnd cell_6t
Xbit_r428_c84 bl[84] br[84] wl[428] vdd gnd cell_6t
Xbit_r429_c84 bl[84] br[84] wl[429] vdd gnd cell_6t
Xbit_r430_c84 bl[84] br[84] wl[430] vdd gnd cell_6t
Xbit_r431_c84 bl[84] br[84] wl[431] vdd gnd cell_6t
Xbit_r432_c84 bl[84] br[84] wl[432] vdd gnd cell_6t
Xbit_r433_c84 bl[84] br[84] wl[433] vdd gnd cell_6t
Xbit_r434_c84 bl[84] br[84] wl[434] vdd gnd cell_6t
Xbit_r435_c84 bl[84] br[84] wl[435] vdd gnd cell_6t
Xbit_r436_c84 bl[84] br[84] wl[436] vdd gnd cell_6t
Xbit_r437_c84 bl[84] br[84] wl[437] vdd gnd cell_6t
Xbit_r438_c84 bl[84] br[84] wl[438] vdd gnd cell_6t
Xbit_r439_c84 bl[84] br[84] wl[439] vdd gnd cell_6t
Xbit_r440_c84 bl[84] br[84] wl[440] vdd gnd cell_6t
Xbit_r441_c84 bl[84] br[84] wl[441] vdd gnd cell_6t
Xbit_r442_c84 bl[84] br[84] wl[442] vdd gnd cell_6t
Xbit_r443_c84 bl[84] br[84] wl[443] vdd gnd cell_6t
Xbit_r444_c84 bl[84] br[84] wl[444] vdd gnd cell_6t
Xbit_r445_c84 bl[84] br[84] wl[445] vdd gnd cell_6t
Xbit_r446_c84 bl[84] br[84] wl[446] vdd gnd cell_6t
Xbit_r447_c84 bl[84] br[84] wl[447] vdd gnd cell_6t
Xbit_r448_c84 bl[84] br[84] wl[448] vdd gnd cell_6t
Xbit_r449_c84 bl[84] br[84] wl[449] vdd gnd cell_6t
Xbit_r450_c84 bl[84] br[84] wl[450] vdd gnd cell_6t
Xbit_r451_c84 bl[84] br[84] wl[451] vdd gnd cell_6t
Xbit_r452_c84 bl[84] br[84] wl[452] vdd gnd cell_6t
Xbit_r453_c84 bl[84] br[84] wl[453] vdd gnd cell_6t
Xbit_r454_c84 bl[84] br[84] wl[454] vdd gnd cell_6t
Xbit_r455_c84 bl[84] br[84] wl[455] vdd gnd cell_6t
Xbit_r456_c84 bl[84] br[84] wl[456] vdd gnd cell_6t
Xbit_r457_c84 bl[84] br[84] wl[457] vdd gnd cell_6t
Xbit_r458_c84 bl[84] br[84] wl[458] vdd gnd cell_6t
Xbit_r459_c84 bl[84] br[84] wl[459] vdd gnd cell_6t
Xbit_r460_c84 bl[84] br[84] wl[460] vdd gnd cell_6t
Xbit_r461_c84 bl[84] br[84] wl[461] vdd gnd cell_6t
Xbit_r462_c84 bl[84] br[84] wl[462] vdd gnd cell_6t
Xbit_r463_c84 bl[84] br[84] wl[463] vdd gnd cell_6t
Xbit_r464_c84 bl[84] br[84] wl[464] vdd gnd cell_6t
Xbit_r465_c84 bl[84] br[84] wl[465] vdd gnd cell_6t
Xbit_r466_c84 bl[84] br[84] wl[466] vdd gnd cell_6t
Xbit_r467_c84 bl[84] br[84] wl[467] vdd gnd cell_6t
Xbit_r468_c84 bl[84] br[84] wl[468] vdd gnd cell_6t
Xbit_r469_c84 bl[84] br[84] wl[469] vdd gnd cell_6t
Xbit_r470_c84 bl[84] br[84] wl[470] vdd gnd cell_6t
Xbit_r471_c84 bl[84] br[84] wl[471] vdd gnd cell_6t
Xbit_r472_c84 bl[84] br[84] wl[472] vdd gnd cell_6t
Xbit_r473_c84 bl[84] br[84] wl[473] vdd gnd cell_6t
Xbit_r474_c84 bl[84] br[84] wl[474] vdd gnd cell_6t
Xbit_r475_c84 bl[84] br[84] wl[475] vdd gnd cell_6t
Xbit_r476_c84 bl[84] br[84] wl[476] vdd gnd cell_6t
Xbit_r477_c84 bl[84] br[84] wl[477] vdd gnd cell_6t
Xbit_r478_c84 bl[84] br[84] wl[478] vdd gnd cell_6t
Xbit_r479_c84 bl[84] br[84] wl[479] vdd gnd cell_6t
Xbit_r480_c84 bl[84] br[84] wl[480] vdd gnd cell_6t
Xbit_r481_c84 bl[84] br[84] wl[481] vdd gnd cell_6t
Xbit_r482_c84 bl[84] br[84] wl[482] vdd gnd cell_6t
Xbit_r483_c84 bl[84] br[84] wl[483] vdd gnd cell_6t
Xbit_r484_c84 bl[84] br[84] wl[484] vdd gnd cell_6t
Xbit_r485_c84 bl[84] br[84] wl[485] vdd gnd cell_6t
Xbit_r486_c84 bl[84] br[84] wl[486] vdd gnd cell_6t
Xbit_r487_c84 bl[84] br[84] wl[487] vdd gnd cell_6t
Xbit_r488_c84 bl[84] br[84] wl[488] vdd gnd cell_6t
Xbit_r489_c84 bl[84] br[84] wl[489] vdd gnd cell_6t
Xbit_r490_c84 bl[84] br[84] wl[490] vdd gnd cell_6t
Xbit_r491_c84 bl[84] br[84] wl[491] vdd gnd cell_6t
Xbit_r492_c84 bl[84] br[84] wl[492] vdd gnd cell_6t
Xbit_r493_c84 bl[84] br[84] wl[493] vdd gnd cell_6t
Xbit_r494_c84 bl[84] br[84] wl[494] vdd gnd cell_6t
Xbit_r495_c84 bl[84] br[84] wl[495] vdd gnd cell_6t
Xbit_r496_c84 bl[84] br[84] wl[496] vdd gnd cell_6t
Xbit_r497_c84 bl[84] br[84] wl[497] vdd gnd cell_6t
Xbit_r498_c84 bl[84] br[84] wl[498] vdd gnd cell_6t
Xbit_r499_c84 bl[84] br[84] wl[499] vdd gnd cell_6t
Xbit_r500_c84 bl[84] br[84] wl[500] vdd gnd cell_6t
Xbit_r501_c84 bl[84] br[84] wl[501] vdd gnd cell_6t
Xbit_r502_c84 bl[84] br[84] wl[502] vdd gnd cell_6t
Xbit_r503_c84 bl[84] br[84] wl[503] vdd gnd cell_6t
Xbit_r504_c84 bl[84] br[84] wl[504] vdd gnd cell_6t
Xbit_r505_c84 bl[84] br[84] wl[505] vdd gnd cell_6t
Xbit_r506_c84 bl[84] br[84] wl[506] vdd gnd cell_6t
Xbit_r507_c84 bl[84] br[84] wl[507] vdd gnd cell_6t
Xbit_r508_c84 bl[84] br[84] wl[508] vdd gnd cell_6t
Xbit_r509_c84 bl[84] br[84] wl[509] vdd gnd cell_6t
Xbit_r510_c84 bl[84] br[84] wl[510] vdd gnd cell_6t
Xbit_r511_c84 bl[84] br[84] wl[511] vdd gnd cell_6t
Xbit_r0_c85 bl[85] br[85] wl[0] vdd gnd cell_6t
Xbit_r1_c85 bl[85] br[85] wl[1] vdd gnd cell_6t
Xbit_r2_c85 bl[85] br[85] wl[2] vdd gnd cell_6t
Xbit_r3_c85 bl[85] br[85] wl[3] vdd gnd cell_6t
Xbit_r4_c85 bl[85] br[85] wl[4] vdd gnd cell_6t
Xbit_r5_c85 bl[85] br[85] wl[5] vdd gnd cell_6t
Xbit_r6_c85 bl[85] br[85] wl[6] vdd gnd cell_6t
Xbit_r7_c85 bl[85] br[85] wl[7] vdd gnd cell_6t
Xbit_r8_c85 bl[85] br[85] wl[8] vdd gnd cell_6t
Xbit_r9_c85 bl[85] br[85] wl[9] vdd gnd cell_6t
Xbit_r10_c85 bl[85] br[85] wl[10] vdd gnd cell_6t
Xbit_r11_c85 bl[85] br[85] wl[11] vdd gnd cell_6t
Xbit_r12_c85 bl[85] br[85] wl[12] vdd gnd cell_6t
Xbit_r13_c85 bl[85] br[85] wl[13] vdd gnd cell_6t
Xbit_r14_c85 bl[85] br[85] wl[14] vdd gnd cell_6t
Xbit_r15_c85 bl[85] br[85] wl[15] vdd gnd cell_6t
Xbit_r16_c85 bl[85] br[85] wl[16] vdd gnd cell_6t
Xbit_r17_c85 bl[85] br[85] wl[17] vdd gnd cell_6t
Xbit_r18_c85 bl[85] br[85] wl[18] vdd gnd cell_6t
Xbit_r19_c85 bl[85] br[85] wl[19] vdd gnd cell_6t
Xbit_r20_c85 bl[85] br[85] wl[20] vdd gnd cell_6t
Xbit_r21_c85 bl[85] br[85] wl[21] vdd gnd cell_6t
Xbit_r22_c85 bl[85] br[85] wl[22] vdd gnd cell_6t
Xbit_r23_c85 bl[85] br[85] wl[23] vdd gnd cell_6t
Xbit_r24_c85 bl[85] br[85] wl[24] vdd gnd cell_6t
Xbit_r25_c85 bl[85] br[85] wl[25] vdd gnd cell_6t
Xbit_r26_c85 bl[85] br[85] wl[26] vdd gnd cell_6t
Xbit_r27_c85 bl[85] br[85] wl[27] vdd gnd cell_6t
Xbit_r28_c85 bl[85] br[85] wl[28] vdd gnd cell_6t
Xbit_r29_c85 bl[85] br[85] wl[29] vdd gnd cell_6t
Xbit_r30_c85 bl[85] br[85] wl[30] vdd gnd cell_6t
Xbit_r31_c85 bl[85] br[85] wl[31] vdd gnd cell_6t
Xbit_r32_c85 bl[85] br[85] wl[32] vdd gnd cell_6t
Xbit_r33_c85 bl[85] br[85] wl[33] vdd gnd cell_6t
Xbit_r34_c85 bl[85] br[85] wl[34] vdd gnd cell_6t
Xbit_r35_c85 bl[85] br[85] wl[35] vdd gnd cell_6t
Xbit_r36_c85 bl[85] br[85] wl[36] vdd gnd cell_6t
Xbit_r37_c85 bl[85] br[85] wl[37] vdd gnd cell_6t
Xbit_r38_c85 bl[85] br[85] wl[38] vdd gnd cell_6t
Xbit_r39_c85 bl[85] br[85] wl[39] vdd gnd cell_6t
Xbit_r40_c85 bl[85] br[85] wl[40] vdd gnd cell_6t
Xbit_r41_c85 bl[85] br[85] wl[41] vdd gnd cell_6t
Xbit_r42_c85 bl[85] br[85] wl[42] vdd gnd cell_6t
Xbit_r43_c85 bl[85] br[85] wl[43] vdd gnd cell_6t
Xbit_r44_c85 bl[85] br[85] wl[44] vdd gnd cell_6t
Xbit_r45_c85 bl[85] br[85] wl[45] vdd gnd cell_6t
Xbit_r46_c85 bl[85] br[85] wl[46] vdd gnd cell_6t
Xbit_r47_c85 bl[85] br[85] wl[47] vdd gnd cell_6t
Xbit_r48_c85 bl[85] br[85] wl[48] vdd gnd cell_6t
Xbit_r49_c85 bl[85] br[85] wl[49] vdd gnd cell_6t
Xbit_r50_c85 bl[85] br[85] wl[50] vdd gnd cell_6t
Xbit_r51_c85 bl[85] br[85] wl[51] vdd gnd cell_6t
Xbit_r52_c85 bl[85] br[85] wl[52] vdd gnd cell_6t
Xbit_r53_c85 bl[85] br[85] wl[53] vdd gnd cell_6t
Xbit_r54_c85 bl[85] br[85] wl[54] vdd gnd cell_6t
Xbit_r55_c85 bl[85] br[85] wl[55] vdd gnd cell_6t
Xbit_r56_c85 bl[85] br[85] wl[56] vdd gnd cell_6t
Xbit_r57_c85 bl[85] br[85] wl[57] vdd gnd cell_6t
Xbit_r58_c85 bl[85] br[85] wl[58] vdd gnd cell_6t
Xbit_r59_c85 bl[85] br[85] wl[59] vdd gnd cell_6t
Xbit_r60_c85 bl[85] br[85] wl[60] vdd gnd cell_6t
Xbit_r61_c85 bl[85] br[85] wl[61] vdd gnd cell_6t
Xbit_r62_c85 bl[85] br[85] wl[62] vdd gnd cell_6t
Xbit_r63_c85 bl[85] br[85] wl[63] vdd gnd cell_6t
Xbit_r64_c85 bl[85] br[85] wl[64] vdd gnd cell_6t
Xbit_r65_c85 bl[85] br[85] wl[65] vdd gnd cell_6t
Xbit_r66_c85 bl[85] br[85] wl[66] vdd gnd cell_6t
Xbit_r67_c85 bl[85] br[85] wl[67] vdd gnd cell_6t
Xbit_r68_c85 bl[85] br[85] wl[68] vdd gnd cell_6t
Xbit_r69_c85 bl[85] br[85] wl[69] vdd gnd cell_6t
Xbit_r70_c85 bl[85] br[85] wl[70] vdd gnd cell_6t
Xbit_r71_c85 bl[85] br[85] wl[71] vdd gnd cell_6t
Xbit_r72_c85 bl[85] br[85] wl[72] vdd gnd cell_6t
Xbit_r73_c85 bl[85] br[85] wl[73] vdd gnd cell_6t
Xbit_r74_c85 bl[85] br[85] wl[74] vdd gnd cell_6t
Xbit_r75_c85 bl[85] br[85] wl[75] vdd gnd cell_6t
Xbit_r76_c85 bl[85] br[85] wl[76] vdd gnd cell_6t
Xbit_r77_c85 bl[85] br[85] wl[77] vdd gnd cell_6t
Xbit_r78_c85 bl[85] br[85] wl[78] vdd gnd cell_6t
Xbit_r79_c85 bl[85] br[85] wl[79] vdd gnd cell_6t
Xbit_r80_c85 bl[85] br[85] wl[80] vdd gnd cell_6t
Xbit_r81_c85 bl[85] br[85] wl[81] vdd gnd cell_6t
Xbit_r82_c85 bl[85] br[85] wl[82] vdd gnd cell_6t
Xbit_r83_c85 bl[85] br[85] wl[83] vdd gnd cell_6t
Xbit_r84_c85 bl[85] br[85] wl[84] vdd gnd cell_6t
Xbit_r85_c85 bl[85] br[85] wl[85] vdd gnd cell_6t
Xbit_r86_c85 bl[85] br[85] wl[86] vdd gnd cell_6t
Xbit_r87_c85 bl[85] br[85] wl[87] vdd gnd cell_6t
Xbit_r88_c85 bl[85] br[85] wl[88] vdd gnd cell_6t
Xbit_r89_c85 bl[85] br[85] wl[89] vdd gnd cell_6t
Xbit_r90_c85 bl[85] br[85] wl[90] vdd gnd cell_6t
Xbit_r91_c85 bl[85] br[85] wl[91] vdd gnd cell_6t
Xbit_r92_c85 bl[85] br[85] wl[92] vdd gnd cell_6t
Xbit_r93_c85 bl[85] br[85] wl[93] vdd gnd cell_6t
Xbit_r94_c85 bl[85] br[85] wl[94] vdd gnd cell_6t
Xbit_r95_c85 bl[85] br[85] wl[95] vdd gnd cell_6t
Xbit_r96_c85 bl[85] br[85] wl[96] vdd gnd cell_6t
Xbit_r97_c85 bl[85] br[85] wl[97] vdd gnd cell_6t
Xbit_r98_c85 bl[85] br[85] wl[98] vdd gnd cell_6t
Xbit_r99_c85 bl[85] br[85] wl[99] vdd gnd cell_6t
Xbit_r100_c85 bl[85] br[85] wl[100] vdd gnd cell_6t
Xbit_r101_c85 bl[85] br[85] wl[101] vdd gnd cell_6t
Xbit_r102_c85 bl[85] br[85] wl[102] vdd gnd cell_6t
Xbit_r103_c85 bl[85] br[85] wl[103] vdd gnd cell_6t
Xbit_r104_c85 bl[85] br[85] wl[104] vdd gnd cell_6t
Xbit_r105_c85 bl[85] br[85] wl[105] vdd gnd cell_6t
Xbit_r106_c85 bl[85] br[85] wl[106] vdd gnd cell_6t
Xbit_r107_c85 bl[85] br[85] wl[107] vdd gnd cell_6t
Xbit_r108_c85 bl[85] br[85] wl[108] vdd gnd cell_6t
Xbit_r109_c85 bl[85] br[85] wl[109] vdd gnd cell_6t
Xbit_r110_c85 bl[85] br[85] wl[110] vdd gnd cell_6t
Xbit_r111_c85 bl[85] br[85] wl[111] vdd gnd cell_6t
Xbit_r112_c85 bl[85] br[85] wl[112] vdd gnd cell_6t
Xbit_r113_c85 bl[85] br[85] wl[113] vdd gnd cell_6t
Xbit_r114_c85 bl[85] br[85] wl[114] vdd gnd cell_6t
Xbit_r115_c85 bl[85] br[85] wl[115] vdd gnd cell_6t
Xbit_r116_c85 bl[85] br[85] wl[116] vdd gnd cell_6t
Xbit_r117_c85 bl[85] br[85] wl[117] vdd gnd cell_6t
Xbit_r118_c85 bl[85] br[85] wl[118] vdd gnd cell_6t
Xbit_r119_c85 bl[85] br[85] wl[119] vdd gnd cell_6t
Xbit_r120_c85 bl[85] br[85] wl[120] vdd gnd cell_6t
Xbit_r121_c85 bl[85] br[85] wl[121] vdd gnd cell_6t
Xbit_r122_c85 bl[85] br[85] wl[122] vdd gnd cell_6t
Xbit_r123_c85 bl[85] br[85] wl[123] vdd gnd cell_6t
Xbit_r124_c85 bl[85] br[85] wl[124] vdd gnd cell_6t
Xbit_r125_c85 bl[85] br[85] wl[125] vdd gnd cell_6t
Xbit_r126_c85 bl[85] br[85] wl[126] vdd gnd cell_6t
Xbit_r127_c85 bl[85] br[85] wl[127] vdd gnd cell_6t
Xbit_r128_c85 bl[85] br[85] wl[128] vdd gnd cell_6t
Xbit_r129_c85 bl[85] br[85] wl[129] vdd gnd cell_6t
Xbit_r130_c85 bl[85] br[85] wl[130] vdd gnd cell_6t
Xbit_r131_c85 bl[85] br[85] wl[131] vdd gnd cell_6t
Xbit_r132_c85 bl[85] br[85] wl[132] vdd gnd cell_6t
Xbit_r133_c85 bl[85] br[85] wl[133] vdd gnd cell_6t
Xbit_r134_c85 bl[85] br[85] wl[134] vdd gnd cell_6t
Xbit_r135_c85 bl[85] br[85] wl[135] vdd gnd cell_6t
Xbit_r136_c85 bl[85] br[85] wl[136] vdd gnd cell_6t
Xbit_r137_c85 bl[85] br[85] wl[137] vdd gnd cell_6t
Xbit_r138_c85 bl[85] br[85] wl[138] vdd gnd cell_6t
Xbit_r139_c85 bl[85] br[85] wl[139] vdd gnd cell_6t
Xbit_r140_c85 bl[85] br[85] wl[140] vdd gnd cell_6t
Xbit_r141_c85 bl[85] br[85] wl[141] vdd gnd cell_6t
Xbit_r142_c85 bl[85] br[85] wl[142] vdd gnd cell_6t
Xbit_r143_c85 bl[85] br[85] wl[143] vdd gnd cell_6t
Xbit_r144_c85 bl[85] br[85] wl[144] vdd gnd cell_6t
Xbit_r145_c85 bl[85] br[85] wl[145] vdd gnd cell_6t
Xbit_r146_c85 bl[85] br[85] wl[146] vdd gnd cell_6t
Xbit_r147_c85 bl[85] br[85] wl[147] vdd gnd cell_6t
Xbit_r148_c85 bl[85] br[85] wl[148] vdd gnd cell_6t
Xbit_r149_c85 bl[85] br[85] wl[149] vdd gnd cell_6t
Xbit_r150_c85 bl[85] br[85] wl[150] vdd gnd cell_6t
Xbit_r151_c85 bl[85] br[85] wl[151] vdd gnd cell_6t
Xbit_r152_c85 bl[85] br[85] wl[152] vdd gnd cell_6t
Xbit_r153_c85 bl[85] br[85] wl[153] vdd gnd cell_6t
Xbit_r154_c85 bl[85] br[85] wl[154] vdd gnd cell_6t
Xbit_r155_c85 bl[85] br[85] wl[155] vdd gnd cell_6t
Xbit_r156_c85 bl[85] br[85] wl[156] vdd gnd cell_6t
Xbit_r157_c85 bl[85] br[85] wl[157] vdd gnd cell_6t
Xbit_r158_c85 bl[85] br[85] wl[158] vdd gnd cell_6t
Xbit_r159_c85 bl[85] br[85] wl[159] vdd gnd cell_6t
Xbit_r160_c85 bl[85] br[85] wl[160] vdd gnd cell_6t
Xbit_r161_c85 bl[85] br[85] wl[161] vdd gnd cell_6t
Xbit_r162_c85 bl[85] br[85] wl[162] vdd gnd cell_6t
Xbit_r163_c85 bl[85] br[85] wl[163] vdd gnd cell_6t
Xbit_r164_c85 bl[85] br[85] wl[164] vdd gnd cell_6t
Xbit_r165_c85 bl[85] br[85] wl[165] vdd gnd cell_6t
Xbit_r166_c85 bl[85] br[85] wl[166] vdd gnd cell_6t
Xbit_r167_c85 bl[85] br[85] wl[167] vdd gnd cell_6t
Xbit_r168_c85 bl[85] br[85] wl[168] vdd gnd cell_6t
Xbit_r169_c85 bl[85] br[85] wl[169] vdd gnd cell_6t
Xbit_r170_c85 bl[85] br[85] wl[170] vdd gnd cell_6t
Xbit_r171_c85 bl[85] br[85] wl[171] vdd gnd cell_6t
Xbit_r172_c85 bl[85] br[85] wl[172] vdd gnd cell_6t
Xbit_r173_c85 bl[85] br[85] wl[173] vdd gnd cell_6t
Xbit_r174_c85 bl[85] br[85] wl[174] vdd gnd cell_6t
Xbit_r175_c85 bl[85] br[85] wl[175] vdd gnd cell_6t
Xbit_r176_c85 bl[85] br[85] wl[176] vdd gnd cell_6t
Xbit_r177_c85 bl[85] br[85] wl[177] vdd gnd cell_6t
Xbit_r178_c85 bl[85] br[85] wl[178] vdd gnd cell_6t
Xbit_r179_c85 bl[85] br[85] wl[179] vdd gnd cell_6t
Xbit_r180_c85 bl[85] br[85] wl[180] vdd gnd cell_6t
Xbit_r181_c85 bl[85] br[85] wl[181] vdd gnd cell_6t
Xbit_r182_c85 bl[85] br[85] wl[182] vdd gnd cell_6t
Xbit_r183_c85 bl[85] br[85] wl[183] vdd gnd cell_6t
Xbit_r184_c85 bl[85] br[85] wl[184] vdd gnd cell_6t
Xbit_r185_c85 bl[85] br[85] wl[185] vdd gnd cell_6t
Xbit_r186_c85 bl[85] br[85] wl[186] vdd gnd cell_6t
Xbit_r187_c85 bl[85] br[85] wl[187] vdd gnd cell_6t
Xbit_r188_c85 bl[85] br[85] wl[188] vdd gnd cell_6t
Xbit_r189_c85 bl[85] br[85] wl[189] vdd gnd cell_6t
Xbit_r190_c85 bl[85] br[85] wl[190] vdd gnd cell_6t
Xbit_r191_c85 bl[85] br[85] wl[191] vdd gnd cell_6t
Xbit_r192_c85 bl[85] br[85] wl[192] vdd gnd cell_6t
Xbit_r193_c85 bl[85] br[85] wl[193] vdd gnd cell_6t
Xbit_r194_c85 bl[85] br[85] wl[194] vdd gnd cell_6t
Xbit_r195_c85 bl[85] br[85] wl[195] vdd gnd cell_6t
Xbit_r196_c85 bl[85] br[85] wl[196] vdd gnd cell_6t
Xbit_r197_c85 bl[85] br[85] wl[197] vdd gnd cell_6t
Xbit_r198_c85 bl[85] br[85] wl[198] vdd gnd cell_6t
Xbit_r199_c85 bl[85] br[85] wl[199] vdd gnd cell_6t
Xbit_r200_c85 bl[85] br[85] wl[200] vdd gnd cell_6t
Xbit_r201_c85 bl[85] br[85] wl[201] vdd gnd cell_6t
Xbit_r202_c85 bl[85] br[85] wl[202] vdd gnd cell_6t
Xbit_r203_c85 bl[85] br[85] wl[203] vdd gnd cell_6t
Xbit_r204_c85 bl[85] br[85] wl[204] vdd gnd cell_6t
Xbit_r205_c85 bl[85] br[85] wl[205] vdd gnd cell_6t
Xbit_r206_c85 bl[85] br[85] wl[206] vdd gnd cell_6t
Xbit_r207_c85 bl[85] br[85] wl[207] vdd gnd cell_6t
Xbit_r208_c85 bl[85] br[85] wl[208] vdd gnd cell_6t
Xbit_r209_c85 bl[85] br[85] wl[209] vdd gnd cell_6t
Xbit_r210_c85 bl[85] br[85] wl[210] vdd gnd cell_6t
Xbit_r211_c85 bl[85] br[85] wl[211] vdd gnd cell_6t
Xbit_r212_c85 bl[85] br[85] wl[212] vdd gnd cell_6t
Xbit_r213_c85 bl[85] br[85] wl[213] vdd gnd cell_6t
Xbit_r214_c85 bl[85] br[85] wl[214] vdd gnd cell_6t
Xbit_r215_c85 bl[85] br[85] wl[215] vdd gnd cell_6t
Xbit_r216_c85 bl[85] br[85] wl[216] vdd gnd cell_6t
Xbit_r217_c85 bl[85] br[85] wl[217] vdd gnd cell_6t
Xbit_r218_c85 bl[85] br[85] wl[218] vdd gnd cell_6t
Xbit_r219_c85 bl[85] br[85] wl[219] vdd gnd cell_6t
Xbit_r220_c85 bl[85] br[85] wl[220] vdd gnd cell_6t
Xbit_r221_c85 bl[85] br[85] wl[221] vdd gnd cell_6t
Xbit_r222_c85 bl[85] br[85] wl[222] vdd gnd cell_6t
Xbit_r223_c85 bl[85] br[85] wl[223] vdd gnd cell_6t
Xbit_r224_c85 bl[85] br[85] wl[224] vdd gnd cell_6t
Xbit_r225_c85 bl[85] br[85] wl[225] vdd gnd cell_6t
Xbit_r226_c85 bl[85] br[85] wl[226] vdd gnd cell_6t
Xbit_r227_c85 bl[85] br[85] wl[227] vdd gnd cell_6t
Xbit_r228_c85 bl[85] br[85] wl[228] vdd gnd cell_6t
Xbit_r229_c85 bl[85] br[85] wl[229] vdd gnd cell_6t
Xbit_r230_c85 bl[85] br[85] wl[230] vdd gnd cell_6t
Xbit_r231_c85 bl[85] br[85] wl[231] vdd gnd cell_6t
Xbit_r232_c85 bl[85] br[85] wl[232] vdd gnd cell_6t
Xbit_r233_c85 bl[85] br[85] wl[233] vdd gnd cell_6t
Xbit_r234_c85 bl[85] br[85] wl[234] vdd gnd cell_6t
Xbit_r235_c85 bl[85] br[85] wl[235] vdd gnd cell_6t
Xbit_r236_c85 bl[85] br[85] wl[236] vdd gnd cell_6t
Xbit_r237_c85 bl[85] br[85] wl[237] vdd gnd cell_6t
Xbit_r238_c85 bl[85] br[85] wl[238] vdd gnd cell_6t
Xbit_r239_c85 bl[85] br[85] wl[239] vdd gnd cell_6t
Xbit_r240_c85 bl[85] br[85] wl[240] vdd gnd cell_6t
Xbit_r241_c85 bl[85] br[85] wl[241] vdd gnd cell_6t
Xbit_r242_c85 bl[85] br[85] wl[242] vdd gnd cell_6t
Xbit_r243_c85 bl[85] br[85] wl[243] vdd gnd cell_6t
Xbit_r244_c85 bl[85] br[85] wl[244] vdd gnd cell_6t
Xbit_r245_c85 bl[85] br[85] wl[245] vdd gnd cell_6t
Xbit_r246_c85 bl[85] br[85] wl[246] vdd gnd cell_6t
Xbit_r247_c85 bl[85] br[85] wl[247] vdd gnd cell_6t
Xbit_r248_c85 bl[85] br[85] wl[248] vdd gnd cell_6t
Xbit_r249_c85 bl[85] br[85] wl[249] vdd gnd cell_6t
Xbit_r250_c85 bl[85] br[85] wl[250] vdd gnd cell_6t
Xbit_r251_c85 bl[85] br[85] wl[251] vdd gnd cell_6t
Xbit_r252_c85 bl[85] br[85] wl[252] vdd gnd cell_6t
Xbit_r253_c85 bl[85] br[85] wl[253] vdd gnd cell_6t
Xbit_r254_c85 bl[85] br[85] wl[254] vdd gnd cell_6t
Xbit_r255_c85 bl[85] br[85] wl[255] vdd gnd cell_6t
Xbit_r256_c85 bl[85] br[85] wl[256] vdd gnd cell_6t
Xbit_r257_c85 bl[85] br[85] wl[257] vdd gnd cell_6t
Xbit_r258_c85 bl[85] br[85] wl[258] vdd gnd cell_6t
Xbit_r259_c85 bl[85] br[85] wl[259] vdd gnd cell_6t
Xbit_r260_c85 bl[85] br[85] wl[260] vdd gnd cell_6t
Xbit_r261_c85 bl[85] br[85] wl[261] vdd gnd cell_6t
Xbit_r262_c85 bl[85] br[85] wl[262] vdd gnd cell_6t
Xbit_r263_c85 bl[85] br[85] wl[263] vdd gnd cell_6t
Xbit_r264_c85 bl[85] br[85] wl[264] vdd gnd cell_6t
Xbit_r265_c85 bl[85] br[85] wl[265] vdd gnd cell_6t
Xbit_r266_c85 bl[85] br[85] wl[266] vdd gnd cell_6t
Xbit_r267_c85 bl[85] br[85] wl[267] vdd gnd cell_6t
Xbit_r268_c85 bl[85] br[85] wl[268] vdd gnd cell_6t
Xbit_r269_c85 bl[85] br[85] wl[269] vdd gnd cell_6t
Xbit_r270_c85 bl[85] br[85] wl[270] vdd gnd cell_6t
Xbit_r271_c85 bl[85] br[85] wl[271] vdd gnd cell_6t
Xbit_r272_c85 bl[85] br[85] wl[272] vdd gnd cell_6t
Xbit_r273_c85 bl[85] br[85] wl[273] vdd gnd cell_6t
Xbit_r274_c85 bl[85] br[85] wl[274] vdd gnd cell_6t
Xbit_r275_c85 bl[85] br[85] wl[275] vdd gnd cell_6t
Xbit_r276_c85 bl[85] br[85] wl[276] vdd gnd cell_6t
Xbit_r277_c85 bl[85] br[85] wl[277] vdd gnd cell_6t
Xbit_r278_c85 bl[85] br[85] wl[278] vdd gnd cell_6t
Xbit_r279_c85 bl[85] br[85] wl[279] vdd gnd cell_6t
Xbit_r280_c85 bl[85] br[85] wl[280] vdd gnd cell_6t
Xbit_r281_c85 bl[85] br[85] wl[281] vdd gnd cell_6t
Xbit_r282_c85 bl[85] br[85] wl[282] vdd gnd cell_6t
Xbit_r283_c85 bl[85] br[85] wl[283] vdd gnd cell_6t
Xbit_r284_c85 bl[85] br[85] wl[284] vdd gnd cell_6t
Xbit_r285_c85 bl[85] br[85] wl[285] vdd gnd cell_6t
Xbit_r286_c85 bl[85] br[85] wl[286] vdd gnd cell_6t
Xbit_r287_c85 bl[85] br[85] wl[287] vdd gnd cell_6t
Xbit_r288_c85 bl[85] br[85] wl[288] vdd gnd cell_6t
Xbit_r289_c85 bl[85] br[85] wl[289] vdd gnd cell_6t
Xbit_r290_c85 bl[85] br[85] wl[290] vdd gnd cell_6t
Xbit_r291_c85 bl[85] br[85] wl[291] vdd gnd cell_6t
Xbit_r292_c85 bl[85] br[85] wl[292] vdd gnd cell_6t
Xbit_r293_c85 bl[85] br[85] wl[293] vdd gnd cell_6t
Xbit_r294_c85 bl[85] br[85] wl[294] vdd gnd cell_6t
Xbit_r295_c85 bl[85] br[85] wl[295] vdd gnd cell_6t
Xbit_r296_c85 bl[85] br[85] wl[296] vdd gnd cell_6t
Xbit_r297_c85 bl[85] br[85] wl[297] vdd gnd cell_6t
Xbit_r298_c85 bl[85] br[85] wl[298] vdd gnd cell_6t
Xbit_r299_c85 bl[85] br[85] wl[299] vdd gnd cell_6t
Xbit_r300_c85 bl[85] br[85] wl[300] vdd gnd cell_6t
Xbit_r301_c85 bl[85] br[85] wl[301] vdd gnd cell_6t
Xbit_r302_c85 bl[85] br[85] wl[302] vdd gnd cell_6t
Xbit_r303_c85 bl[85] br[85] wl[303] vdd gnd cell_6t
Xbit_r304_c85 bl[85] br[85] wl[304] vdd gnd cell_6t
Xbit_r305_c85 bl[85] br[85] wl[305] vdd gnd cell_6t
Xbit_r306_c85 bl[85] br[85] wl[306] vdd gnd cell_6t
Xbit_r307_c85 bl[85] br[85] wl[307] vdd gnd cell_6t
Xbit_r308_c85 bl[85] br[85] wl[308] vdd gnd cell_6t
Xbit_r309_c85 bl[85] br[85] wl[309] vdd gnd cell_6t
Xbit_r310_c85 bl[85] br[85] wl[310] vdd gnd cell_6t
Xbit_r311_c85 bl[85] br[85] wl[311] vdd gnd cell_6t
Xbit_r312_c85 bl[85] br[85] wl[312] vdd gnd cell_6t
Xbit_r313_c85 bl[85] br[85] wl[313] vdd gnd cell_6t
Xbit_r314_c85 bl[85] br[85] wl[314] vdd gnd cell_6t
Xbit_r315_c85 bl[85] br[85] wl[315] vdd gnd cell_6t
Xbit_r316_c85 bl[85] br[85] wl[316] vdd gnd cell_6t
Xbit_r317_c85 bl[85] br[85] wl[317] vdd gnd cell_6t
Xbit_r318_c85 bl[85] br[85] wl[318] vdd gnd cell_6t
Xbit_r319_c85 bl[85] br[85] wl[319] vdd gnd cell_6t
Xbit_r320_c85 bl[85] br[85] wl[320] vdd gnd cell_6t
Xbit_r321_c85 bl[85] br[85] wl[321] vdd gnd cell_6t
Xbit_r322_c85 bl[85] br[85] wl[322] vdd gnd cell_6t
Xbit_r323_c85 bl[85] br[85] wl[323] vdd gnd cell_6t
Xbit_r324_c85 bl[85] br[85] wl[324] vdd gnd cell_6t
Xbit_r325_c85 bl[85] br[85] wl[325] vdd gnd cell_6t
Xbit_r326_c85 bl[85] br[85] wl[326] vdd gnd cell_6t
Xbit_r327_c85 bl[85] br[85] wl[327] vdd gnd cell_6t
Xbit_r328_c85 bl[85] br[85] wl[328] vdd gnd cell_6t
Xbit_r329_c85 bl[85] br[85] wl[329] vdd gnd cell_6t
Xbit_r330_c85 bl[85] br[85] wl[330] vdd gnd cell_6t
Xbit_r331_c85 bl[85] br[85] wl[331] vdd gnd cell_6t
Xbit_r332_c85 bl[85] br[85] wl[332] vdd gnd cell_6t
Xbit_r333_c85 bl[85] br[85] wl[333] vdd gnd cell_6t
Xbit_r334_c85 bl[85] br[85] wl[334] vdd gnd cell_6t
Xbit_r335_c85 bl[85] br[85] wl[335] vdd gnd cell_6t
Xbit_r336_c85 bl[85] br[85] wl[336] vdd gnd cell_6t
Xbit_r337_c85 bl[85] br[85] wl[337] vdd gnd cell_6t
Xbit_r338_c85 bl[85] br[85] wl[338] vdd gnd cell_6t
Xbit_r339_c85 bl[85] br[85] wl[339] vdd gnd cell_6t
Xbit_r340_c85 bl[85] br[85] wl[340] vdd gnd cell_6t
Xbit_r341_c85 bl[85] br[85] wl[341] vdd gnd cell_6t
Xbit_r342_c85 bl[85] br[85] wl[342] vdd gnd cell_6t
Xbit_r343_c85 bl[85] br[85] wl[343] vdd gnd cell_6t
Xbit_r344_c85 bl[85] br[85] wl[344] vdd gnd cell_6t
Xbit_r345_c85 bl[85] br[85] wl[345] vdd gnd cell_6t
Xbit_r346_c85 bl[85] br[85] wl[346] vdd gnd cell_6t
Xbit_r347_c85 bl[85] br[85] wl[347] vdd gnd cell_6t
Xbit_r348_c85 bl[85] br[85] wl[348] vdd gnd cell_6t
Xbit_r349_c85 bl[85] br[85] wl[349] vdd gnd cell_6t
Xbit_r350_c85 bl[85] br[85] wl[350] vdd gnd cell_6t
Xbit_r351_c85 bl[85] br[85] wl[351] vdd gnd cell_6t
Xbit_r352_c85 bl[85] br[85] wl[352] vdd gnd cell_6t
Xbit_r353_c85 bl[85] br[85] wl[353] vdd gnd cell_6t
Xbit_r354_c85 bl[85] br[85] wl[354] vdd gnd cell_6t
Xbit_r355_c85 bl[85] br[85] wl[355] vdd gnd cell_6t
Xbit_r356_c85 bl[85] br[85] wl[356] vdd gnd cell_6t
Xbit_r357_c85 bl[85] br[85] wl[357] vdd gnd cell_6t
Xbit_r358_c85 bl[85] br[85] wl[358] vdd gnd cell_6t
Xbit_r359_c85 bl[85] br[85] wl[359] vdd gnd cell_6t
Xbit_r360_c85 bl[85] br[85] wl[360] vdd gnd cell_6t
Xbit_r361_c85 bl[85] br[85] wl[361] vdd gnd cell_6t
Xbit_r362_c85 bl[85] br[85] wl[362] vdd gnd cell_6t
Xbit_r363_c85 bl[85] br[85] wl[363] vdd gnd cell_6t
Xbit_r364_c85 bl[85] br[85] wl[364] vdd gnd cell_6t
Xbit_r365_c85 bl[85] br[85] wl[365] vdd gnd cell_6t
Xbit_r366_c85 bl[85] br[85] wl[366] vdd gnd cell_6t
Xbit_r367_c85 bl[85] br[85] wl[367] vdd gnd cell_6t
Xbit_r368_c85 bl[85] br[85] wl[368] vdd gnd cell_6t
Xbit_r369_c85 bl[85] br[85] wl[369] vdd gnd cell_6t
Xbit_r370_c85 bl[85] br[85] wl[370] vdd gnd cell_6t
Xbit_r371_c85 bl[85] br[85] wl[371] vdd gnd cell_6t
Xbit_r372_c85 bl[85] br[85] wl[372] vdd gnd cell_6t
Xbit_r373_c85 bl[85] br[85] wl[373] vdd gnd cell_6t
Xbit_r374_c85 bl[85] br[85] wl[374] vdd gnd cell_6t
Xbit_r375_c85 bl[85] br[85] wl[375] vdd gnd cell_6t
Xbit_r376_c85 bl[85] br[85] wl[376] vdd gnd cell_6t
Xbit_r377_c85 bl[85] br[85] wl[377] vdd gnd cell_6t
Xbit_r378_c85 bl[85] br[85] wl[378] vdd gnd cell_6t
Xbit_r379_c85 bl[85] br[85] wl[379] vdd gnd cell_6t
Xbit_r380_c85 bl[85] br[85] wl[380] vdd gnd cell_6t
Xbit_r381_c85 bl[85] br[85] wl[381] vdd gnd cell_6t
Xbit_r382_c85 bl[85] br[85] wl[382] vdd gnd cell_6t
Xbit_r383_c85 bl[85] br[85] wl[383] vdd gnd cell_6t
Xbit_r384_c85 bl[85] br[85] wl[384] vdd gnd cell_6t
Xbit_r385_c85 bl[85] br[85] wl[385] vdd gnd cell_6t
Xbit_r386_c85 bl[85] br[85] wl[386] vdd gnd cell_6t
Xbit_r387_c85 bl[85] br[85] wl[387] vdd gnd cell_6t
Xbit_r388_c85 bl[85] br[85] wl[388] vdd gnd cell_6t
Xbit_r389_c85 bl[85] br[85] wl[389] vdd gnd cell_6t
Xbit_r390_c85 bl[85] br[85] wl[390] vdd gnd cell_6t
Xbit_r391_c85 bl[85] br[85] wl[391] vdd gnd cell_6t
Xbit_r392_c85 bl[85] br[85] wl[392] vdd gnd cell_6t
Xbit_r393_c85 bl[85] br[85] wl[393] vdd gnd cell_6t
Xbit_r394_c85 bl[85] br[85] wl[394] vdd gnd cell_6t
Xbit_r395_c85 bl[85] br[85] wl[395] vdd gnd cell_6t
Xbit_r396_c85 bl[85] br[85] wl[396] vdd gnd cell_6t
Xbit_r397_c85 bl[85] br[85] wl[397] vdd gnd cell_6t
Xbit_r398_c85 bl[85] br[85] wl[398] vdd gnd cell_6t
Xbit_r399_c85 bl[85] br[85] wl[399] vdd gnd cell_6t
Xbit_r400_c85 bl[85] br[85] wl[400] vdd gnd cell_6t
Xbit_r401_c85 bl[85] br[85] wl[401] vdd gnd cell_6t
Xbit_r402_c85 bl[85] br[85] wl[402] vdd gnd cell_6t
Xbit_r403_c85 bl[85] br[85] wl[403] vdd gnd cell_6t
Xbit_r404_c85 bl[85] br[85] wl[404] vdd gnd cell_6t
Xbit_r405_c85 bl[85] br[85] wl[405] vdd gnd cell_6t
Xbit_r406_c85 bl[85] br[85] wl[406] vdd gnd cell_6t
Xbit_r407_c85 bl[85] br[85] wl[407] vdd gnd cell_6t
Xbit_r408_c85 bl[85] br[85] wl[408] vdd gnd cell_6t
Xbit_r409_c85 bl[85] br[85] wl[409] vdd gnd cell_6t
Xbit_r410_c85 bl[85] br[85] wl[410] vdd gnd cell_6t
Xbit_r411_c85 bl[85] br[85] wl[411] vdd gnd cell_6t
Xbit_r412_c85 bl[85] br[85] wl[412] vdd gnd cell_6t
Xbit_r413_c85 bl[85] br[85] wl[413] vdd gnd cell_6t
Xbit_r414_c85 bl[85] br[85] wl[414] vdd gnd cell_6t
Xbit_r415_c85 bl[85] br[85] wl[415] vdd gnd cell_6t
Xbit_r416_c85 bl[85] br[85] wl[416] vdd gnd cell_6t
Xbit_r417_c85 bl[85] br[85] wl[417] vdd gnd cell_6t
Xbit_r418_c85 bl[85] br[85] wl[418] vdd gnd cell_6t
Xbit_r419_c85 bl[85] br[85] wl[419] vdd gnd cell_6t
Xbit_r420_c85 bl[85] br[85] wl[420] vdd gnd cell_6t
Xbit_r421_c85 bl[85] br[85] wl[421] vdd gnd cell_6t
Xbit_r422_c85 bl[85] br[85] wl[422] vdd gnd cell_6t
Xbit_r423_c85 bl[85] br[85] wl[423] vdd gnd cell_6t
Xbit_r424_c85 bl[85] br[85] wl[424] vdd gnd cell_6t
Xbit_r425_c85 bl[85] br[85] wl[425] vdd gnd cell_6t
Xbit_r426_c85 bl[85] br[85] wl[426] vdd gnd cell_6t
Xbit_r427_c85 bl[85] br[85] wl[427] vdd gnd cell_6t
Xbit_r428_c85 bl[85] br[85] wl[428] vdd gnd cell_6t
Xbit_r429_c85 bl[85] br[85] wl[429] vdd gnd cell_6t
Xbit_r430_c85 bl[85] br[85] wl[430] vdd gnd cell_6t
Xbit_r431_c85 bl[85] br[85] wl[431] vdd gnd cell_6t
Xbit_r432_c85 bl[85] br[85] wl[432] vdd gnd cell_6t
Xbit_r433_c85 bl[85] br[85] wl[433] vdd gnd cell_6t
Xbit_r434_c85 bl[85] br[85] wl[434] vdd gnd cell_6t
Xbit_r435_c85 bl[85] br[85] wl[435] vdd gnd cell_6t
Xbit_r436_c85 bl[85] br[85] wl[436] vdd gnd cell_6t
Xbit_r437_c85 bl[85] br[85] wl[437] vdd gnd cell_6t
Xbit_r438_c85 bl[85] br[85] wl[438] vdd gnd cell_6t
Xbit_r439_c85 bl[85] br[85] wl[439] vdd gnd cell_6t
Xbit_r440_c85 bl[85] br[85] wl[440] vdd gnd cell_6t
Xbit_r441_c85 bl[85] br[85] wl[441] vdd gnd cell_6t
Xbit_r442_c85 bl[85] br[85] wl[442] vdd gnd cell_6t
Xbit_r443_c85 bl[85] br[85] wl[443] vdd gnd cell_6t
Xbit_r444_c85 bl[85] br[85] wl[444] vdd gnd cell_6t
Xbit_r445_c85 bl[85] br[85] wl[445] vdd gnd cell_6t
Xbit_r446_c85 bl[85] br[85] wl[446] vdd gnd cell_6t
Xbit_r447_c85 bl[85] br[85] wl[447] vdd gnd cell_6t
Xbit_r448_c85 bl[85] br[85] wl[448] vdd gnd cell_6t
Xbit_r449_c85 bl[85] br[85] wl[449] vdd gnd cell_6t
Xbit_r450_c85 bl[85] br[85] wl[450] vdd gnd cell_6t
Xbit_r451_c85 bl[85] br[85] wl[451] vdd gnd cell_6t
Xbit_r452_c85 bl[85] br[85] wl[452] vdd gnd cell_6t
Xbit_r453_c85 bl[85] br[85] wl[453] vdd gnd cell_6t
Xbit_r454_c85 bl[85] br[85] wl[454] vdd gnd cell_6t
Xbit_r455_c85 bl[85] br[85] wl[455] vdd gnd cell_6t
Xbit_r456_c85 bl[85] br[85] wl[456] vdd gnd cell_6t
Xbit_r457_c85 bl[85] br[85] wl[457] vdd gnd cell_6t
Xbit_r458_c85 bl[85] br[85] wl[458] vdd gnd cell_6t
Xbit_r459_c85 bl[85] br[85] wl[459] vdd gnd cell_6t
Xbit_r460_c85 bl[85] br[85] wl[460] vdd gnd cell_6t
Xbit_r461_c85 bl[85] br[85] wl[461] vdd gnd cell_6t
Xbit_r462_c85 bl[85] br[85] wl[462] vdd gnd cell_6t
Xbit_r463_c85 bl[85] br[85] wl[463] vdd gnd cell_6t
Xbit_r464_c85 bl[85] br[85] wl[464] vdd gnd cell_6t
Xbit_r465_c85 bl[85] br[85] wl[465] vdd gnd cell_6t
Xbit_r466_c85 bl[85] br[85] wl[466] vdd gnd cell_6t
Xbit_r467_c85 bl[85] br[85] wl[467] vdd gnd cell_6t
Xbit_r468_c85 bl[85] br[85] wl[468] vdd gnd cell_6t
Xbit_r469_c85 bl[85] br[85] wl[469] vdd gnd cell_6t
Xbit_r470_c85 bl[85] br[85] wl[470] vdd gnd cell_6t
Xbit_r471_c85 bl[85] br[85] wl[471] vdd gnd cell_6t
Xbit_r472_c85 bl[85] br[85] wl[472] vdd gnd cell_6t
Xbit_r473_c85 bl[85] br[85] wl[473] vdd gnd cell_6t
Xbit_r474_c85 bl[85] br[85] wl[474] vdd gnd cell_6t
Xbit_r475_c85 bl[85] br[85] wl[475] vdd gnd cell_6t
Xbit_r476_c85 bl[85] br[85] wl[476] vdd gnd cell_6t
Xbit_r477_c85 bl[85] br[85] wl[477] vdd gnd cell_6t
Xbit_r478_c85 bl[85] br[85] wl[478] vdd gnd cell_6t
Xbit_r479_c85 bl[85] br[85] wl[479] vdd gnd cell_6t
Xbit_r480_c85 bl[85] br[85] wl[480] vdd gnd cell_6t
Xbit_r481_c85 bl[85] br[85] wl[481] vdd gnd cell_6t
Xbit_r482_c85 bl[85] br[85] wl[482] vdd gnd cell_6t
Xbit_r483_c85 bl[85] br[85] wl[483] vdd gnd cell_6t
Xbit_r484_c85 bl[85] br[85] wl[484] vdd gnd cell_6t
Xbit_r485_c85 bl[85] br[85] wl[485] vdd gnd cell_6t
Xbit_r486_c85 bl[85] br[85] wl[486] vdd gnd cell_6t
Xbit_r487_c85 bl[85] br[85] wl[487] vdd gnd cell_6t
Xbit_r488_c85 bl[85] br[85] wl[488] vdd gnd cell_6t
Xbit_r489_c85 bl[85] br[85] wl[489] vdd gnd cell_6t
Xbit_r490_c85 bl[85] br[85] wl[490] vdd gnd cell_6t
Xbit_r491_c85 bl[85] br[85] wl[491] vdd gnd cell_6t
Xbit_r492_c85 bl[85] br[85] wl[492] vdd gnd cell_6t
Xbit_r493_c85 bl[85] br[85] wl[493] vdd gnd cell_6t
Xbit_r494_c85 bl[85] br[85] wl[494] vdd gnd cell_6t
Xbit_r495_c85 bl[85] br[85] wl[495] vdd gnd cell_6t
Xbit_r496_c85 bl[85] br[85] wl[496] vdd gnd cell_6t
Xbit_r497_c85 bl[85] br[85] wl[497] vdd gnd cell_6t
Xbit_r498_c85 bl[85] br[85] wl[498] vdd gnd cell_6t
Xbit_r499_c85 bl[85] br[85] wl[499] vdd gnd cell_6t
Xbit_r500_c85 bl[85] br[85] wl[500] vdd gnd cell_6t
Xbit_r501_c85 bl[85] br[85] wl[501] vdd gnd cell_6t
Xbit_r502_c85 bl[85] br[85] wl[502] vdd gnd cell_6t
Xbit_r503_c85 bl[85] br[85] wl[503] vdd gnd cell_6t
Xbit_r504_c85 bl[85] br[85] wl[504] vdd gnd cell_6t
Xbit_r505_c85 bl[85] br[85] wl[505] vdd gnd cell_6t
Xbit_r506_c85 bl[85] br[85] wl[506] vdd gnd cell_6t
Xbit_r507_c85 bl[85] br[85] wl[507] vdd gnd cell_6t
Xbit_r508_c85 bl[85] br[85] wl[508] vdd gnd cell_6t
Xbit_r509_c85 bl[85] br[85] wl[509] vdd gnd cell_6t
Xbit_r510_c85 bl[85] br[85] wl[510] vdd gnd cell_6t
Xbit_r511_c85 bl[85] br[85] wl[511] vdd gnd cell_6t
Xbit_r0_c86 bl[86] br[86] wl[0] vdd gnd cell_6t
Xbit_r1_c86 bl[86] br[86] wl[1] vdd gnd cell_6t
Xbit_r2_c86 bl[86] br[86] wl[2] vdd gnd cell_6t
Xbit_r3_c86 bl[86] br[86] wl[3] vdd gnd cell_6t
Xbit_r4_c86 bl[86] br[86] wl[4] vdd gnd cell_6t
Xbit_r5_c86 bl[86] br[86] wl[5] vdd gnd cell_6t
Xbit_r6_c86 bl[86] br[86] wl[6] vdd gnd cell_6t
Xbit_r7_c86 bl[86] br[86] wl[7] vdd gnd cell_6t
Xbit_r8_c86 bl[86] br[86] wl[8] vdd gnd cell_6t
Xbit_r9_c86 bl[86] br[86] wl[9] vdd gnd cell_6t
Xbit_r10_c86 bl[86] br[86] wl[10] vdd gnd cell_6t
Xbit_r11_c86 bl[86] br[86] wl[11] vdd gnd cell_6t
Xbit_r12_c86 bl[86] br[86] wl[12] vdd gnd cell_6t
Xbit_r13_c86 bl[86] br[86] wl[13] vdd gnd cell_6t
Xbit_r14_c86 bl[86] br[86] wl[14] vdd gnd cell_6t
Xbit_r15_c86 bl[86] br[86] wl[15] vdd gnd cell_6t
Xbit_r16_c86 bl[86] br[86] wl[16] vdd gnd cell_6t
Xbit_r17_c86 bl[86] br[86] wl[17] vdd gnd cell_6t
Xbit_r18_c86 bl[86] br[86] wl[18] vdd gnd cell_6t
Xbit_r19_c86 bl[86] br[86] wl[19] vdd gnd cell_6t
Xbit_r20_c86 bl[86] br[86] wl[20] vdd gnd cell_6t
Xbit_r21_c86 bl[86] br[86] wl[21] vdd gnd cell_6t
Xbit_r22_c86 bl[86] br[86] wl[22] vdd gnd cell_6t
Xbit_r23_c86 bl[86] br[86] wl[23] vdd gnd cell_6t
Xbit_r24_c86 bl[86] br[86] wl[24] vdd gnd cell_6t
Xbit_r25_c86 bl[86] br[86] wl[25] vdd gnd cell_6t
Xbit_r26_c86 bl[86] br[86] wl[26] vdd gnd cell_6t
Xbit_r27_c86 bl[86] br[86] wl[27] vdd gnd cell_6t
Xbit_r28_c86 bl[86] br[86] wl[28] vdd gnd cell_6t
Xbit_r29_c86 bl[86] br[86] wl[29] vdd gnd cell_6t
Xbit_r30_c86 bl[86] br[86] wl[30] vdd gnd cell_6t
Xbit_r31_c86 bl[86] br[86] wl[31] vdd gnd cell_6t
Xbit_r32_c86 bl[86] br[86] wl[32] vdd gnd cell_6t
Xbit_r33_c86 bl[86] br[86] wl[33] vdd gnd cell_6t
Xbit_r34_c86 bl[86] br[86] wl[34] vdd gnd cell_6t
Xbit_r35_c86 bl[86] br[86] wl[35] vdd gnd cell_6t
Xbit_r36_c86 bl[86] br[86] wl[36] vdd gnd cell_6t
Xbit_r37_c86 bl[86] br[86] wl[37] vdd gnd cell_6t
Xbit_r38_c86 bl[86] br[86] wl[38] vdd gnd cell_6t
Xbit_r39_c86 bl[86] br[86] wl[39] vdd gnd cell_6t
Xbit_r40_c86 bl[86] br[86] wl[40] vdd gnd cell_6t
Xbit_r41_c86 bl[86] br[86] wl[41] vdd gnd cell_6t
Xbit_r42_c86 bl[86] br[86] wl[42] vdd gnd cell_6t
Xbit_r43_c86 bl[86] br[86] wl[43] vdd gnd cell_6t
Xbit_r44_c86 bl[86] br[86] wl[44] vdd gnd cell_6t
Xbit_r45_c86 bl[86] br[86] wl[45] vdd gnd cell_6t
Xbit_r46_c86 bl[86] br[86] wl[46] vdd gnd cell_6t
Xbit_r47_c86 bl[86] br[86] wl[47] vdd gnd cell_6t
Xbit_r48_c86 bl[86] br[86] wl[48] vdd gnd cell_6t
Xbit_r49_c86 bl[86] br[86] wl[49] vdd gnd cell_6t
Xbit_r50_c86 bl[86] br[86] wl[50] vdd gnd cell_6t
Xbit_r51_c86 bl[86] br[86] wl[51] vdd gnd cell_6t
Xbit_r52_c86 bl[86] br[86] wl[52] vdd gnd cell_6t
Xbit_r53_c86 bl[86] br[86] wl[53] vdd gnd cell_6t
Xbit_r54_c86 bl[86] br[86] wl[54] vdd gnd cell_6t
Xbit_r55_c86 bl[86] br[86] wl[55] vdd gnd cell_6t
Xbit_r56_c86 bl[86] br[86] wl[56] vdd gnd cell_6t
Xbit_r57_c86 bl[86] br[86] wl[57] vdd gnd cell_6t
Xbit_r58_c86 bl[86] br[86] wl[58] vdd gnd cell_6t
Xbit_r59_c86 bl[86] br[86] wl[59] vdd gnd cell_6t
Xbit_r60_c86 bl[86] br[86] wl[60] vdd gnd cell_6t
Xbit_r61_c86 bl[86] br[86] wl[61] vdd gnd cell_6t
Xbit_r62_c86 bl[86] br[86] wl[62] vdd gnd cell_6t
Xbit_r63_c86 bl[86] br[86] wl[63] vdd gnd cell_6t
Xbit_r64_c86 bl[86] br[86] wl[64] vdd gnd cell_6t
Xbit_r65_c86 bl[86] br[86] wl[65] vdd gnd cell_6t
Xbit_r66_c86 bl[86] br[86] wl[66] vdd gnd cell_6t
Xbit_r67_c86 bl[86] br[86] wl[67] vdd gnd cell_6t
Xbit_r68_c86 bl[86] br[86] wl[68] vdd gnd cell_6t
Xbit_r69_c86 bl[86] br[86] wl[69] vdd gnd cell_6t
Xbit_r70_c86 bl[86] br[86] wl[70] vdd gnd cell_6t
Xbit_r71_c86 bl[86] br[86] wl[71] vdd gnd cell_6t
Xbit_r72_c86 bl[86] br[86] wl[72] vdd gnd cell_6t
Xbit_r73_c86 bl[86] br[86] wl[73] vdd gnd cell_6t
Xbit_r74_c86 bl[86] br[86] wl[74] vdd gnd cell_6t
Xbit_r75_c86 bl[86] br[86] wl[75] vdd gnd cell_6t
Xbit_r76_c86 bl[86] br[86] wl[76] vdd gnd cell_6t
Xbit_r77_c86 bl[86] br[86] wl[77] vdd gnd cell_6t
Xbit_r78_c86 bl[86] br[86] wl[78] vdd gnd cell_6t
Xbit_r79_c86 bl[86] br[86] wl[79] vdd gnd cell_6t
Xbit_r80_c86 bl[86] br[86] wl[80] vdd gnd cell_6t
Xbit_r81_c86 bl[86] br[86] wl[81] vdd gnd cell_6t
Xbit_r82_c86 bl[86] br[86] wl[82] vdd gnd cell_6t
Xbit_r83_c86 bl[86] br[86] wl[83] vdd gnd cell_6t
Xbit_r84_c86 bl[86] br[86] wl[84] vdd gnd cell_6t
Xbit_r85_c86 bl[86] br[86] wl[85] vdd gnd cell_6t
Xbit_r86_c86 bl[86] br[86] wl[86] vdd gnd cell_6t
Xbit_r87_c86 bl[86] br[86] wl[87] vdd gnd cell_6t
Xbit_r88_c86 bl[86] br[86] wl[88] vdd gnd cell_6t
Xbit_r89_c86 bl[86] br[86] wl[89] vdd gnd cell_6t
Xbit_r90_c86 bl[86] br[86] wl[90] vdd gnd cell_6t
Xbit_r91_c86 bl[86] br[86] wl[91] vdd gnd cell_6t
Xbit_r92_c86 bl[86] br[86] wl[92] vdd gnd cell_6t
Xbit_r93_c86 bl[86] br[86] wl[93] vdd gnd cell_6t
Xbit_r94_c86 bl[86] br[86] wl[94] vdd gnd cell_6t
Xbit_r95_c86 bl[86] br[86] wl[95] vdd gnd cell_6t
Xbit_r96_c86 bl[86] br[86] wl[96] vdd gnd cell_6t
Xbit_r97_c86 bl[86] br[86] wl[97] vdd gnd cell_6t
Xbit_r98_c86 bl[86] br[86] wl[98] vdd gnd cell_6t
Xbit_r99_c86 bl[86] br[86] wl[99] vdd gnd cell_6t
Xbit_r100_c86 bl[86] br[86] wl[100] vdd gnd cell_6t
Xbit_r101_c86 bl[86] br[86] wl[101] vdd gnd cell_6t
Xbit_r102_c86 bl[86] br[86] wl[102] vdd gnd cell_6t
Xbit_r103_c86 bl[86] br[86] wl[103] vdd gnd cell_6t
Xbit_r104_c86 bl[86] br[86] wl[104] vdd gnd cell_6t
Xbit_r105_c86 bl[86] br[86] wl[105] vdd gnd cell_6t
Xbit_r106_c86 bl[86] br[86] wl[106] vdd gnd cell_6t
Xbit_r107_c86 bl[86] br[86] wl[107] vdd gnd cell_6t
Xbit_r108_c86 bl[86] br[86] wl[108] vdd gnd cell_6t
Xbit_r109_c86 bl[86] br[86] wl[109] vdd gnd cell_6t
Xbit_r110_c86 bl[86] br[86] wl[110] vdd gnd cell_6t
Xbit_r111_c86 bl[86] br[86] wl[111] vdd gnd cell_6t
Xbit_r112_c86 bl[86] br[86] wl[112] vdd gnd cell_6t
Xbit_r113_c86 bl[86] br[86] wl[113] vdd gnd cell_6t
Xbit_r114_c86 bl[86] br[86] wl[114] vdd gnd cell_6t
Xbit_r115_c86 bl[86] br[86] wl[115] vdd gnd cell_6t
Xbit_r116_c86 bl[86] br[86] wl[116] vdd gnd cell_6t
Xbit_r117_c86 bl[86] br[86] wl[117] vdd gnd cell_6t
Xbit_r118_c86 bl[86] br[86] wl[118] vdd gnd cell_6t
Xbit_r119_c86 bl[86] br[86] wl[119] vdd gnd cell_6t
Xbit_r120_c86 bl[86] br[86] wl[120] vdd gnd cell_6t
Xbit_r121_c86 bl[86] br[86] wl[121] vdd gnd cell_6t
Xbit_r122_c86 bl[86] br[86] wl[122] vdd gnd cell_6t
Xbit_r123_c86 bl[86] br[86] wl[123] vdd gnd cell_6t
Xbit_r124_c86 bl[86] br[86] wl[124] vdd gnd cell_6t
Xbit_r125_c86 bl[86] br[86] wl[125] vdd gnd cell_6t
Xbit_r126_c86 bl[86] br[86] wl[126] vdd gnd cell_6t
Xbit_r127_c86 bl[86] br[86] wl[127] vdd gnd cell_6t
Xbit_r128_c86 bl[86] br[86] wl[128] vdd gnd cell_6t
Xbit_r129_c86 bl[86] br[86] wl[129] vdd gnd cell_6t
Xbit_r130_c86 bl[86] br[86] wl[130] vdd gnd cell_6t
Xbit_r131_c86 bl[86] br[86] wl[131] vdd gnd cell_6t
Xbit_r132_c86 bl[86] br[86] wl[132] vdd gnd cell_6t
Xbit_r133_c86 bl[86] br[86] wl[133] vdd gnd cell_6t
Xbit_r134_c86 bl[86] br[86] wl[134] vdd gnd cell_6t
Xbit_r135_c86 bl[86] br[86] wl[135] vdd gnd cell_6t
Xbit_r136_c86 bl[86] br[86] wl[136] vdd gnd cell_6t
Xbit_r137_c86 bl[86] br[86] wl[137] vdd gnd cell_6t
Xbit_r138_c86 bl[86] br[86] wl[138] vdd gnd cell_6t
Xbit_r139_c86 bl[86] br[86] wl[139] vdd gnd cell_6t
Xbit_r140_c86 bl[86] br[86] wl[140] vdd gnd cell_6t
Xbit_r141_c86 bl[86] br[86] wl[141] vdd gnd cell_6t
Xbit_r142_c86 bl[86] br[86] wl[142] vdd gnd cell_6t
Xbit_r143_c86 bl[86] br[86] wl[143] vdd gnd cell_6t
Xbit_r144_c86 bl[86] br[86] wl[144] vdd gnd cell_6t
Xbit_r145_c86 bl[86] br[86] wl[145] vdd gnd cell_6t
Xbit_r146_c86 bl[86] br[86] wl[146] vdd gnd cell_6t
Xbit_r147_c86 bl[86] br[86] wl[147] vdd gnd cell_6t
Xbit_r148_c86 bl[86] br[86] wl[148] vdd gnd cell_6t
Xbit_r149_c86 bl[86] br[86] wl[149] vdd gnd cell_6t
Xbit_r150_c86 bl[86] br[86] wl[150] vdd gnd cell_6t
Xbit_r151_c86 bl[86] br[86] wl[151] vdd gnd cell_6t
Xbit_r152_c86 bl[86] br[86] wl[152] vdd gnd cell_6t
Xbit_r153_c86 bl[86] br[86] wl[153] vdd gnd cell_6t
Xbit_r154_c86 bl[86] br[86] wl[154] vdd gnd cell_6t
Xbit_r155_c86 bl[86] br[86] wl[155] vdd gnd cell_6t
Xbit_r156_c86 bl[86] br[86] wl[156] vdd gnd cell_6t
Xbit_r157_c86 bl[86] br[86] wl[157] vdd gnd cell_6t
Xbit_r158_c86 bl[86] br[86] wl[158] vdd gnd cell_6t
Xbit_r159_c86 bl[86] br[86] wl[159] vdd gnd cell_6t
Xbit_r160_c86 bl[86] br[86] wl[160] vdd gnd cell_6t
Xbit_r161_c86 bl[86] br[86] wl[161] vdd gnd cell_6t
Xbit_r162_c86 bl[86] br[86] wl[162] vdd gnd cell_6t
Xbit_r163_c86 bl[86] br[86] wl[163] vdd gnd cell_6t
Xbit_r164_c86 bl[86] br[86] wl[164] vdd gnd cell_6t
Xbit_r165_c86 bl[86] br[86] wl[165] vdd gnd cell_6t
Xbit_r166_c86 bl[86] br[86] wl[166] vdd gnd cell_6t
Xbit_r167_c86 bl[86] br[86] wl[167] vdd gnd cell_6t
Xbit_r168_c86 bl[86] br[86] wl[168] vdd gnd cell_6t
Xbit_r169_c86 bl[86] br[86] wl[169] vdd gnd cell_6t
Xbit_r170_c86 bl[86] br[86] wl[170] vdd gnd cell_6t
Xbit_r171_c86 bl[86] br[86] wl[171] vdd gnd cell_6t
Xbit_r172_c86 bl[86] br[86] wl[172] vdd gnd cell_6t
Xbit_r173_c86 bl[86] br[86] wl[173] vdd gnd cell_6t
Xbit_r174_c86 bl[86] br[86] wl[174] vdd gnd cell_6t
Xbit_r175_c86 bl[86] br[86] wl[175] vdd gnd cell_6t
Xbit_r176_c86 bl[86] br[86] wl[176] vdd gnd cell_6t
Xbit_r177_c86 bl[86] br[86] wl[177] vdd gnd cell_6t
Xbit_r178_c86 bl[86] br[86] wl[178] vdd gnd cell_6t
Xbit_r179_c86 bl[86] br[86] wl[179] vdd gnd cell_6t
Xbit_r180_c86 bl[86] br[86] wl[180] vdd gnd cell_6t
Xbit_r181_c86 bl[86] br[86] wl[181] vdd gnd cell_6t
Xbit_r182_c86 bl[86] br[86] wl[182] vdd gnd cell_6t
Xbit_r183_c86 bl[86] br[86] wl[183] vdd gnd cell_6t
Xbit_r184_c86 bl[86] br[86] wl[184] vdd gnd cell_6t
Xbit_r185_c86 bl[86] br[86] wl[185] vdd gnd cell_6t
Xbit_r186_c86 bl[86] br[86] wl[186] vdd gnd cell_6t
Xbit_r187_c86 bl[86] br[86] wl[187] vdd gnd cell_6t
Xbit_r188_c86 bl[86] br[86] wl[188] vdd gnd cell_6t
Xbit_r189_c86 bl[86] br[86] wl[189] vdd gnd cell_6t
Xbit_r190_c86 bl[86] br[86] wl[190] vdd gnd cell_6t
Xbit_r191_c86 bl[86] br[86] wl[191] vdd gnd cell_6t
Xbit_r192_c86 bl[86] br[86] wl[192] vdd gnd cell_6t
Xbit_r193_c86 bl[86] br[86] wl[193] vdd gnd cell_6t
Xbit_r194_c86 bl[86] br[86] wl[194] vdd gnd cell_6t
Xbit_r195_c86 bl[86] br[86] wl[195] vdd gnd cell_6t
Xbit_r196_c86 bl[86] br[86] wl[196] vdd gnd cell_6t
Xbit_r197_c86 bl[86] br[86] wl[197] vdd gnd cell_6t
Xbit_r198_c86 bl[86] br[86] wl[198] vdd gnd cell_6t
Xbit_r199_c86 bl[86] br[86] wl[199] vdd gnd cell_6t
Xbit_r200_c86 bl[86] br[86] wl[200] vdd gnd cell_6t
Xbit_r201_c86 bl[86] br[86] wl[201] vdd gnd cell_6t
Xbit_r202_c86 bl[86] br[86] wl[202] vdd gnd cell_6t
Xbit_r203_c86 bl[86] br[86] wl[203] vdd gnd cell_6t
Xbit_r204_c86 bl[86] br[86] wl[204] vdd gnd cell_6t
Xbit_r205_c86 bl[86] br[86] wl[205] vdd gnd cell_6t
Xbit_r206_c86 bl[86] br[86] wl[206] vdd gnd cell_6t
Xbit_r207_c86 bl[86] br[86] wl[207] vdd gnd cell_6t
Xbit_r208_c86 bl[86] br[86] wl[208] vdd gnd cell_6t
Xbit_r209_c86 bl[86] br[86] wl[209] vdd gnd cell_6t
Xbit_r210_c86 bl[86] br[86] wl[210] vdd gnd cell_6t
Xbit_r211_c86 bl[86] br[86] wl[211] vdd gnd cell_6t
Xbit_r212_c86 bl[86] br[86] wl[212] vdd gnd cell_6t
Xbit_r213_c86 bl[86] br[86] wl[213] vdd gnd cell_6t
Xbit_r214_c86 bl[86] br[86] wl[214] vdd gnd cell_6t
Xbit_r215_c86 bl[86] br[86] wl[215] vdd gnd cell_6t
Xbit_r216_c86 bl[86] br[86] wl[216] vdd gnd cell_6t
Xbit_r217_c86 bl[86] br[86] wl[217] vdd gnd cell_6t
Xbit_r218_c86 bl[86] br[86] wl[218] vdd gnd cell_6t
Xbit_r219_c86 bl[86] br[86] wl[219] vdd gnd cell_6t
Xbit_r220_c86 bl[86] br[86] wl[220] vdd gnd cell_6t
Xbit_r221_c86 bl[86] br[86] wl[221] vdd gnd cell_6t
Xbit_r222_c86 bl[86] br[86] wl[222] vdd gnd cell_6t
Xbit_r223_c86 bl[86] br[86] wl[223] vdd gnd cell_6t
Xbit_r224_c86 bl[86] br[86] wl[224] vdd gnd cell_6t
Xbit_r225_c86 bl[86] br[86] wl[225] vdd gnd cell_6t
Xbit_r226_c86 bl[86] br[86] wl[226] vdd gnd cell_6t
Xbit_r227_c86 bl[86] br[86] wl[227] vdd gnd cell_6t
Xbit_r228_c86 bl[86] br[86] wl[228] vdd gnd cell_6t
Xbit_r229_c86 bl[86] br[86] wl[229] vdd gnd cell_6t
Xbit_r230_c86 bl[86] br[86] wl[230] vdd gnd cell_6t
Xbit_r231_c86 bl[86] br[86] wl[231] vdd gnd cell_6t
Xbit_r232_c86 bl[86] br[86] wl[232] vdd gnd cell_6t
Xbit_r233_c86 bl[86] br[86] wl[233] vdd gnd cell_6t
Xbit_r234_c86 bl[86] br[86] wl[234] vdd gnd cell_6t
Xbit_r235_c86 bl[86] br[86] wl[235] vdd gnd cell_6t
Xbit_r236_c86 bl[86] br[86] wl[236] vdd gnd cell_6t
Xbit_r237_c86 bl[86] br[86] wl[237] vdd gnd cell_6t
Xbit_r238_c86 bl[86] br[86] wl[238] vdd gnd cell_6t
Xbit_r239_c86 bl[86] br[86] wl[239] vdd gnd cell_6t
Xbit_r240_c86 bl[86] br[86] wl[240] vdd gnd cell_6t
Xbit_r241_c86 bl[86] br[86] wl[241] vdd gnd cell_6t
Xbit_r242_c86 bl[86] br[86] wl[242] vdd gnd cell_6t
Xbit_r243_c86 bl[86] br[86] wl[243] vdd gnd cell_6t
Xbit_r244_c86 bl[86] br[86] wl[244] vdd gnd cell_6t
Xbit_r245_c86 bl[86] br[86] wl[245] vdd gnd cell_6t
Xbit_r246_c86 bl[86] br[86] wl[246] vdd gnd cell_6t
Xbit_r247_c86 bl[86] br[86] wl[247] vdd gnd cell_6t
Xbit_r248_c86 bl[86] br[86] wl[248] vdd gnd cell_6t
Xbit_r249_c86 bl[86] br[86] wl[249] vdd gnd cell_6t
Xbit_r250_c86 bl[86] br[86] wl[250] vdd gnd cell_6t
Xbit_r251_c86 bl[86] br[86] wl[251] vdd gnd cell_6t
Xbit_r252_c86 bl[86] br[86] wl[252] vdd gnd cell_6t
Xbit_r253_c86 bl[86] br[86] wl[253] vdd gnd cell_6t
Xbit_r254_c86 bl[86] br[86] wl[254] vdd gnd cell_6t
Xbit_r255_c86 bl[86] br[86] wl[255] vdd gnd cell_6t
Xbit_r256_c86 bl[86] br[86] wl[256] vdd gnd cell_6t
Xbit_r257_c86 bl[86] br[86] wl[257] vdd gnd cell_6t
Xbit_r258_c86 bl[86] br[86] wl[258] vdd gnd cell_6t
Xbit_r259_c86 bl[86] br[86] wl[259] vdd gnd cell_6t
Xbit_r260_c86 bl[86] br[86] wl[260] vdd gnd cell_6t
Xbit_r261_c86 bl[86] br[86] wl[261] vdd gnd cell_6t
Xbit_r262_c86 bl[86] br[86] wl[262] vdd gnd cell_6t
Xbit_r263_c86 bl[86] br[86] wl[263] vdd gnd cell_6t
Xbit_r264_c86 bl[86] br[86] wl[264] vdd gnd cell_6t
Xbit_r265_c86 bl[86] br[86] wl[265] vdd gnd cell_6t
Xbit_r266_c86 bl[86] br[86] wl[266] vdd gnd cell_6t
Xbit_r267_c86 bl[86] br[86] wl[267] vdd gnd cell_6t
Xbit_r268_c86 bl[86] br[86] wl[268] vdd gnd cell_6t
Xbit_r269_c86 bl[86] br[86] wl[269] vdd gnd cell_6t
Xbit_r270_c86 bl[86] br[86] wl[270] vdd gnd cell_6t
Xbit_r271_c86 bl[86] br[86] wl[271] vdd gnd cell_6t
Xbit_r272_c86 bl[86] br[86] wl[272] vdd gnd cell_6t
Xbit_r273_c86 bl[86] br[86] wl[273] vdd gnd cell_6t
Xbit_r274_c86 bl[86] br[86] wl[274] vdd gnd cell_6t
Xbit_r275_c86 bl[86] br[86] wl[275] vdd gnd cell_6t
Xbit_r276_c86 bl[86] br[86] wl[276] vdd gnd cell_6t
Xbit_r277_c86 bl[86] br[86] wl[277] vdd gnd cell_6t
Xbit_r278_c86 bl[86] br[86] wl[278] vdd gnd cell_6t
Xbit_r279_c86 bl[86] br[86] wl[279] vdd gnd cell_6t
Xbit_r280_c86 bl[86] br[86] wl[280] vdd gnd cell_6t
Xbit_r281_c86 bl[86] br[86] wl[281] vdd gnd cell_6t
Xbit_r282_c86 bl[86] br[86] wl[282] vdd gnd cell_6t
Xbit_r283_c86 bl[86] br[86] wl[283] vdd gnd cell_6t
Xbit_r284_c86 bl[86] br[86] wl[284] vdd gnd cell_6t
Xbit_r285_c86 bl[86] br[86] wl[285] vdd gnd cell_6t
Xbit_r286_c86 bl[86] br[86] wl[286] vdd gnd cell_6t
Xbit_r287_c86 bl[86] br[86] wl[287] vdd gnd cell_6t
Xbit_r288_c86 bl[86] br[86] wl[288] vdd gnd cell_6t
Xbit_r289_c86 bl[86] br[86] wl[289] vdd gnd cell_6t
Xbit_r290_c86 bl[86] br[86] wl[290] vdd gnd cell_6t
Xbit_r291_c86 bl[86] br[86] wl[291] vdd gnd cell_6t
Xbit_r292_c86 bl[86] br[86] wl[292] vdd gnd cell_6t
Xbit_r293_c86 bl[86] br[86] wl[293] vdd gnd cell_6t
Xbit_r294_c86 bl[86] br[86] wl[294] vdd gnd cell_6t
Xbit_r295_c86 bl[86] br[86] wl[295] vdd gnd cell_6t
Xbit_r296_c86 bl[86] br[86] wl[296] vdd gnd cell_6t
Xbit_r297_c86 bl[86] br[86] wl[297] vdd gnd cell_6t
Xbit_r298_c86 bl[86] br[86] wl[298] vdd gnd cell_6t
Xbit_r299_c86 bl[86] br[86] wl[299] vdd gnd cell_6t
Xbit_r300_c86 bl[86] br[86] wl[300] vdd gnd cell_6t
Xbit_r301_c86 bl[86] br[86] wl[301] vdd gnd cell_6t
Xbit_r302_c86 bl[86] br[86] wl[302] vdd gnd cell_6t
Xbit_r303_c86 bl[86] br[86] wl[303] vdd gnd cell_6t
Xbit_r304_c86 bl[86] br[86] wl[304] vdd gnd cell_6t
Xbit_r305_c86 bl[86] br[86] wl[305] vdd gnd cell_6t
Xbit_r306_c86 bl[86] br[86] wl[306] vdd gnd cell_6t
Xbit_r307_c86 bl[86] br[86] wl[307] vdd gnd cell_6t
Xbit_r308_c86 bl[86] br[86] wl[308] vdd gnd cell_6t
Xbit_r309_c86 bl[86] br[86] wl[309] vdd gnd cell_6t
Xbit_r310_c86 bl[86] br[86] wl[310] vdd gnd cell_6t
Xbit_r311_c86 bl[86] br[86] wl[311] vdd gnd cell_6t
Xbit_r312_c86 bl[86] br[86] wl[312] vdd gnd cell_6t
Xbit_r313_c86 bl[86] br[86] wl[313] vdd gnd cell_6t
Xbit_r314_c86 bl[86] br[86] wl[314] vdd gnd cell_6t
Xbit_r315_c86 bl[86] br[86] wl[315] vdd gnd cell_6t
Xbit_r316_c86 bl[86] br[86] wl[316] vdd gnd cell_6t
Xbit_r317_c86 bl[86] br[86] wl[317] vdd gnd cell_6t
Xbit_r318_c86 bl[86] br[86] wl[318] vdd gnd cell_6t
Xbit_r319_c86 bl[86] br[86] wl[319] vdd gnd cell_6t
Xbit_r320_c86 bl[86] br[86] wl[320] vdd gnd cell_6t
Xbit_r321_c86 bl[86] br[86] wl[321] vdd gnd cell_6t
Xbit_r322_c86 bl[86] br[86] wl[322] vdd gnd cell_6t
Xbit_r323_c86 bl[86] br[86] wl[323] vdd gnd cell_6t
Xbit_r324_c86 bl[86] br[86] wl[324] vdd gnd cell_6t
Xbit_r325_c86 bl[86] br[86] wl[325] vdd gnd cell_6t
Xbit_r326_c86 bl[86] br[86] wl[326] vdd gnd cell_6t
Xbit_r327_c86 bl[86] br[86] wl[327] vdd gnd cell_6t
Xbit_r328_c86 bl[86] br[86] wl[328] vdd gnd cell_6t
Xbit_r329_c86 bl[86] br[86] wl[329] vdd gnd cell_6t
Xbit_r330_c86 bl[86] br[86] wl[330] vdd gnd cell_6t
Xbit_r331_c86 bl[86] br[86] wl[331] vdd gnd cell_6t
Xbit_r332_c86 bl[86] br[86] wl[332] vdd gnd cell_6t
Xbit_r333_c86 bl[86] br[86] wl[333] vdd gnd cell_6t
Xbit_r334_c86 bl[86] br[86] wl[334] vdd gnd cell_6t
Xbit_r335_c86 bl[86] br[86] wl[335] vdd gnd cell_6t
Xbit_r336_c86 bl[86] br[86] wl[336] vdd gnd cell_6t
Xbit_r337_c86 bl[86] br[86] wl[337] vdd gnd cell_6t
Xbit_r338_c86 bl[86] br[86] wl[338] vdd gnd cell_6t
Xbit_r339_c86 bl[86] br[86] wl[339] vdd gnd cell_6t
Xbit_r340_c86 bl[86] br[86] wl[340] vdd gnd cell_6t
Xbit_r341_c86 bl[86] br[86] wl[341] vdd gnd cell_6t
Xbit_r342_c86 bl[86] br[86] wl[342] vdd gnd cell_6t
Xbit_r343_c86 bl[86] br[86] wl[343] vdd gnd cell_6t
Xbit_r344_c86 bl[86] br[86] wl[344] vdd gnd cell_6t
Xbit_r345_c86 bl[86] br[86] wl[345] vdd gnd cell_6t
Xbit_r346_c86 bl[86] br[86] wl[346] vdd gnd cell_6t
Xbit_r347_c86 bl[86] br[86] wl[347] vdd gnd cell_6t
Xbit_r348_c86 bl[86] br[86] wl[348] vdd gnd cell_6t
Xbit_r349_c86 bl[86] br[86] wl[349] vdd gnd cell_6t
Xbit_r350_c86 bl[86] br[86] wl[350] vdd gnd cell_6t
Xbit_r351_c86 bl[86] br[86] wl[351] vdd gnd cell_6t
Xbit_r352_c86 bl[86] br[86] wl[352] vdd gnd cell_6t
Xbit_r353_c86 bl[86] br[86] wl[353] vdd gnd cell_6t
Xbit_r354_c86 bl[86] br[86] wl[354] vdd gnd cell_6t
Xbit_r355_c86 bl[86] br[86] wl[355] vdd gnd cell_6t
Xbit_r356_c86 bl[86] br[86] wl[356] vdd gnd cell_6t
Xbit_r357_c86 bl[86] br[86] wl[357] vdd gnd cell_6t
Xbit_r358_c86 bl[86] br[86] wl[358] vdd gnd cell_6t
Xbit_r359_c86 bl[86] br[86] wl[359] vdd gnd cell_6t
Xbit_r360_c86 bl[86] br[86] wl[360] vdd gnd cell_6t
Xbit_r361_c86 bl[86] br[86] wl[361] vdd gnd cell_6t
Xbit_r362_c86 bl[86] br[86] wl[362] vdd gnd cell_6t
Xbit_r363_c86 bl[86] br[86] wl[363] vdd gnd cell_6t
Xbit_r364_c86 bl[86] br[86] wl[364] vdd gnd cell_6t
Xbit_r365_c86 bl[86] br[86] wl[365] vdd gnd cell_6t
Xbit_r366_c86 bl[86] br[86] wl[366] vdd gnd cell_6t
Xbit_r367_c86 bl[86] br[86] wl[367] vdd gnd cell_6t
Xbit_r368_c86 bl[86] br[86] wl[368] vdd gnd cell_6t
Xbit_r369_c86 bl[86] br[86] wl[369] vdd gnd cell_6t
Xbit_r370_c86 bl[86] br[86] wl[370] vdd gnd cell_6t
Xbit_r371_c86 bl[86] br[86] wl[371] vdd gnd cell_6t
Xbit_r372_c86 bl[86] br[86] wl[372] vdd gnd cell_6t
Xbit_r373_c86 bl[86] br[86] wl[373] vdd gnd cell_6t
Xbit_r374_c86 bl[86] br[86] wl[374] vdd gnd cell_6t
Xbit_r375_c86 bl[86] br[86] wl[375] vdd gnd cell_6t
Xbit_r376_c86 bl[86] br[86] wl[376] vdd gnd cell_6t
Xbit_r377_c86 bl[86] br[86] wl[377] vdd gnd cell_6t
Xbit_r378_c86 bl[86] br[86] wl[378] vdd gnd cell_6t
Xbit_r379_c86 bl[86] br[86] wl[379] vdd gnd cell_6t
Xbit_r380_c86 bl[86] br[86] wl[380] vdd gnd cell_6t
Xbit_r381_c86 bl[86] br[86] wl[381] vdd gnd cell_6t
Xbit_r382_c86 bl[86] br[86] wl[382] vdd gnd cell_6t
Xbit_r383_c86 bl[86] br[86] wl[383] vdd gnd cell_6t
Xbit_r384_c86 bl[86] br[86] wl[384] vdd gnd cell_6t
Xbit_r385_c86 bl[86] br[86] wl[385] vdd gnd cell_6t
Xbit_r386_c86 bl[86] br[86] wl[386] vdd gnd cell_6t
Xbit_r387_c86 bl[86] br[86] wl[387] vdd gnd cell_6t
Xbit_r388_c86 bl[86] br[86] wl[388] vdd gnd cell_6t
Xbit_r389_c86 bl[86] br[86] wl[389] vdd gnd cell_6t
Xbit_r390_c86 bl[86] br[86] wl[390] vdd gnd cell_6t
Xbit_r391_c86 bl[86] br[86] wl[391] vdd gnd cell_6t
Xbit_r392_c86 bl[86] br[86] wl[392] vdd gnd cell_6t
Xbit_r393_c86 bl[86] br[86] wl[393] vdd gnd cell_6t
Xbit_r394_c86 bl[86] br[86] wl[394] vdd gnd cell_6t
Xbit_r395_c86 bl[86] br[86] wl[395] vdd gnd cell_6t
Xbit_r396_c86 bl[86] br[86] wl[396] vdd gnd cell_6t
Xbit_r397_c86 bl[86] br[86] wl[397] vdd gnd cell_6t
Xbit_r398_c86 bl[86] br[86] wl[398] vdd gnd cell_6t
Xbit_r399_c86 bl[86] br[86] wl[399] vdd gnd cell_6t
Xbit_r400_c86 bl[86] br[86] wl[400] vdd gnd cell_6t
Xbit_r401_c86 bl[86] br[86] wl[401] vdd gnd cell_6t
Xbit_r402_c86 bl[86] br[86] wl[402] vdd gnd cell_6t
Xbit_r403_c86 bl[86] br[86] wl[403] vdd gnd cell_6t
Xbit_r404_c86 bl[86] br[86] wl[404] vdd gnd cell_6t
Xbit_r405_c86 bl[86] br[86] wl[405] vdd gnd cell_6t
Xbit_r406_c86 bl[86] br[86] wl[406] vdd gnd cell_6t
Xbit_r407_c86 bl[86] br[86] wl[407] vdd gnd cell_6t
Xbit_r408_c86 bl[86] br[86] wl[408] vdd gnd cell_6t
Xbit_r409_c86 bl[86] br[86] wl[409] vdd gnd cell_6t
Xbit_r410_c86 bl[86] br[86] wl[410] vdd gnd cell_6t
Xbit_r411_c86 bl[86] br[86] wl[411] vdd gnd cell_6t
Xbit_r412_c86 bl[86] br[86] wl[412] vdd gnd cell_6t
Xbit_r413_c86 bl[86] br[86] wl[413] vdd gnd cell_6t
Xbit_r414_c86 bl[86] br[86] wl[414] vdd gnd cell_6t
Xbit_r415_c86 bl[86] br[86] wl[415] vdd gnd cell_6t
Xbit_r416_c86 bl[86] br[86] wl[416] vdd gnd cell_6t
Xbit_r417_c86 bl[86] br[86] wl[417] vdd gnd cell_6t
Xbit_r418_c86 bl[86] br[86] wl[418] vdd gnd cell_6t
Xbit_r419_c86 bl[86] br[86] wl[419] vdd gnd cell_6t
Xbit_r420_c86 bl[86] br[86] wl[420] vdd gnd cell_6t
Xbit_r421_c86 bl[86] br[86] wl[421] vdd gnd cell_6t
Xbit_r422_c86 bl[86] br[86] wl[422] vdd gnd cell_6t
Xbit_r423_c86 bl[86] br[86] wl[423] vdd gnd cell_6t
Xbit_r424_c86 bl[86] br[86] wl[424] vdd gnd cell_6t
Xbit_r425_c86 bl[86] br[86] wl[425] vdd gnd cell_6t
Xbit_r426_c86 bl[86] br[86] wl[426] vdd gnd cell_6t
Xbit_r427_c86 bl[86] br[86] wl[427] vdd gnd cell_6t
Xbit_r428_c86 bl[86] br[86] wl[428] vdd gnd cell_6t
Xbit_r429_c86 bl[86] br[86] wl[429] vdd gnd cell_6t
Xbit_r430_c86 bl[86] br[86] wl[430] vdd gnd cell_6t
Xbit_r431_c86 bl[86] br[86] wl[431] vdd gnd cell_6t
Xbit_r432_c86 bl[86] br[86] wl[432] vdd gnd cell_6t
Xbit_r433_c86 bl[86] br[86] wl[433] vdd gnd cell_6t
Xbit_r434_c86 bl[86] br[86] wl[434] vdd gnd cell_6t
Xbit_r435_c86 bl[86] br[86] wl[435] vdd gnd cell_6t
Xbit_r436_c86 bl[86] br[86] wl[436] vdd gnd cell_6t
Xbit_r437_c86 bl[86] br[86] wl[437] vdd gnd cell_6t
Xbit_r438_c86 bl[86] br[86] wl[438] vdd gnd cell_6t
Xbit_r439_c86 bl[86] br[86] wl[439] vdd gnd cell_6t
Xbit_r440_c86 bl[86] br[86] wl[440] vdd gnd cell_6t
Xbit_r441_c86 bl[86] br[86] wl[441] vdd gnd cell_6t
Xbit_r442_c86 bl[86] br[86] wl[442] vdd gnd cell_6t
Xbit_r443_c86 bl[86] br[86] wl[443] vdd gnd cell_6t
Xbit_r444_c86 bl[86] br[86] wl[444] vdd gnd cell_6t
Xbit_r445_c86 bl[86] br[86] wl[445] vdd gnd cell_6t
Xbit_r446_c86 bl[86] br[86] wl[446] vdd gnd cell_6t
Xbit_r447_c86 bl[86] br[86] wl[447] vdd gnd cell_6t
Xbit_r448_c86 bl[86] br[86] wl[448] vdd gnd cell_6t
Xbit_r449_c86 bl[86] br[86] wl[449] vdd gnd cell_6t
Xbit_r450_c86 bl[86] br[86] wl[450] vdd gnd cell_6t
Xbit_r451_c86 bl[86] br[86] wl[451] vdd gnd cell_6t
Xbit_r452_c86 bl[86] br[86] wl[452] vdd gnd cell_6t
Xbit_r453_c86 bl[86] br[86] wl[453] vdd gnd cell_6t
Xbit_r454_c86 bl[86] br[86] wl[454] vdd gnd cell_6t
Xbit_r455_c86 bl[86] br[86] wl[455] vdd gnd cell_6t
Xbit_r456_c86 bl[86] br[86] wl[456] vdd gnd cell_6t
Xbit_r457_c86 bl[86] br[86] wl[457] vdd gnd cell_6t
Xbit_r458_c86 bl[86] br[86] wl[458] vdd gnd cell_6t
Xbit_r459_c86 bl[86] br[86] wl[459] vdd gnd cell_6t
Xbit_r460_c86 bl[86] br[86] wl[460] vdd gnd cell_6t
Xbit_r461_c86 bl[86] br[86] wl[461] vdd gnd cell_6t
Xbit_r462_c86 bl[86] br[86] wl[462] vdd gnd cell_6t
Xbit_r463_c86 bl[86] br[86] wl[463] vdd gnd cell_6t
Xbit_r464_c86 bl[86] br[86] wl[464] vdd gnd cell_6t
Xbit_r465_c86 bl[86] br[86] wl[465] vdd gnd cell_6t
Xbit_r466_c86 bl[86] br[86] wl[466] vdd gnd cell_6t
Xbit_r467_c86 bl[86] br[86] wl[467] vdd gnd cell_6t
Xbit_r468_c86 bl[86] br[86] wl[468] vdd gnd cell_6t
Xbit_r469_c86 bl[86] br[86] wl[469] vdd gnd cell_6t
Xbit_r470_c86 bl[86] br[86] wl[470] vdd gnd cell_6t
Xbit_r471_c86 bl[86] br[86] wl[471] vdd gnd cell_6t
Xbit_r472_c86 bl[86] br[86] wl[472] vdd gnd cell_6t
Xbit_r473_c86 bl[86] br[86] wl[473] vdd gnd cell_6t
Xbit_r474_c86 bl[86] br[86] wl[474] vdd gnd cell_6t
Xbit_r475_c86 bl[86] br[86] wl[475] vdd gnd cell_6t
Xbit_r476_c86 bl[86] br[86] wl[476] vdd gnd cell_6t
Xbit_r477_c86 bl[86] br[86] wl[477] vdd gnd cell_6t
Xbit_r478_c86 bl[86] br[86] wl[478] vdd gnd cell_6t
Xbit_r479_c86 bl[86] br[86] wl[479] vdd gnd cell_6t
Xbit_r480_c86 bl[86] br[86] wl[480] vdd gnd cell_6t
Xbit_r481_c86 bl[86] br[86] wl[481] vdd gnd cell_6t
Xbit_r482_c86 bl[86] br[86] wl[482] vdd gnd cell_6t
Xbit_r483_c86 bl[86] br[86] wl[483] vdd gnd cell_6t
Xbit_r484_c86 bl[86] br[86] wl[484] vdd gnd cell_6t
Xbit_r485_c86 bl[86] br[86] wl[485] vdd gnd cell_6t
Xbit_r486_c86 bl[86] br[86] wl[486] vdd gnd cell_6t
Xbit_r487_c86 bl[86] br[86] wl[487] vdd gnd cell_6t
Xbit_r488_c86 bl[86] br[86] wl[488] vdd gnd cell_6t
Xbit_r489_c86 bl[86] br[86] wl[489] vdd gnd cell_6t
Xbit_r490_c86 bl[86] br[86] wl[490] vdd gnd cell_6t
Xbit_r491_c86 bl[86] br[86] wl[491] vdd gnd cell_6t
Xbit_r492_c86 bl[86] br[86] wl[492] vdd gnd cell_6t
Xbit_r493_c86 bl[86] br[86] wl[493] vdd gnd cell_6t
Xbit_r494_c86 bl[86] br[86] wl[494] vdd gnd cell_6t
Xbit_r495_c86 bl[86] br[86] wl[495] vdd gnd cell_6t
Xbit_r496_c86 bl[86] br[86] wl[496] vdd gnd cell_6t
Xbit_r497_c86 bl[86] br[86] wl[497] vdd gnd cell_6t
Xbit_r498_c86 bl[86] br[86] wl[498] vdd gnd cell_6t
Xbit_r499_c86 bl[86] br[86] wl[499] vdd gnd cell_6t
Xbit_r500_c86 bl[86] br[86] wl[500] vdd gnd cell_6t
Xbit_r501_c86 bl[86] br[86] wl[501] vdd gnd cell_6t
Xbit_r502_c86 bl[86] br[86] wl[502] vdd gnd cell_6t
Xbit_r503_c86 bl[86] br[86] wl[503] vdd gnd cell_6t
Xbit_r504_c86 bl[86] br[86] wl[504] vdd gnd cell_6t
Xbit_r505_c86 bl[86] br[86] wl[505] vdd gnd cell_6t
Xbit_r506_c86 bl[86] br[86] wl[506] vdd gnd cell_6t
Xbit_r507_c86 bl[86] br[86] wl[507] vdd gnd cell_6t
Xbit_r508_c86 bl[86] br[86] wl[508] vdd gnd cell_6t
Xbit_r509_c86 bl[86] br[86] wl[509] vdd gnd cell_6t
Xbit_r510_c86 bl[86] br[86] wl[510] vdd gnd cell_6t
Xbit_r511_c86 bl[86] br[86] wl[511] vdd gnd cell_6t
Xbit_r0_c87 bl[87] br[87] wl[0] vdd gnd cell_6t
Xbit_r1_c87 bl[87] br[87] wl[1] vdd gnd cell_6t
Xbit_r2_c87 bl[87] br[87] wl[2] vdd gnd cell_6t
Xbit_r3_c87 bl[87] br[87] wl[3] vdd gnd cell_6t
Xbit_r4_c87 bl[87] br[87] wl[4] vdd gnd cell_6t
Xbit_r5_c87 bl[87] br[87] wl[5] vdd gnd cell_6t
Xbit_r6_c87 bl[87] br[87] wl[6] vdd gnd cell_6t
Xbit_r7_c87 bl[87] br[87] wl[7] vdd gnd cell_6t
Xbit_r8_c87 bl[87] br[87] wl[8] vdd gnd cell_6t
Xbit_r9_c87 bl[87] br[87] wl[9] vdd gnd cell_6t
Xbit_r10_c87 bl[87] br[87] wl[10] vdd gnd cell_6t
Xbit_r11_c87 bl[87] br[87] wl[11] vdd gnd cell_6t
Xbit_r12_c87 bl[87] br[87] wl[12] vdd gnd cell_6t
Xbit_r13_c87 bl[87] br[87] wl[13] vdd gnd cell_6t
Xbit_r14_c87 bl[87] br[87] wl[14] vdd gnd cell_6t
Xbit_r15_c87 bl[87] br[87] wl[15] vdd gnd cell_6t
Xbit_r16_c87 bl[87] br[87] wl[16] vdd gnd cell_6t
Xbit_r17_c87 bl[87] br[87] wl[17] vdd gnd cell_6t
Xbit_r18_c87 bl[87] br[87] wl[18] vdd gnd cell_6t
Xbit_r19_c87 bl[87] br[87] wl[19] vdd gnd cell_6t
Xbit_r20_c87 bl[87] br[87] wl[20] vdd gnd cell_6t
Xbit_r21_c87 bl[87] br[87] wl[21] vdd gnd cell_6t
Xbit_r22_c87 bl[87] br[87] wl[22] vdd gnd cell_6t
Xbit_r23_c87 bl[87] br[87] wl[23] vdd gnd cell_6t
Xbit_r24_c87 bl[87] br[87] wl[24] vdd gnd cell_6t
Xbit_r25_c87 bl[87] br[87] wl[25] vdd gnd cell_6t
Xbit_r26_c87 bl[87] br[87] wl[26] vdd gnd cell_6t
Xbit_r27_c87 bl[87] br[87] wl[27] vdd gnd cell_6t
Xbit_r28_c87 bl[87] br[87] wl[28] vdd gnd cell_6t
Xbit_r29_c87 bl[87] br[87] wl[29] vdd gnd cell_6t
Xbit_r30_c87 bl[87] br[87] wl[30] vdd gnd cell_6t
Xbit_r31_c87 bl[87] br[87] wl[31] vdd gnd cell_6t
Xbit_r32_c87 bl[87] br[87] wl[32] vdd gnd cell_6t
Xbit_r33_c87 bl[87] br[87] wl[33] vdd gnd cell_6t
Xbit_r34_c87 bl[87] br[87] wl[34] vdd gnd cell_6t
Xbit_r35_c87 bl[87] br[87] wl[35] vdd gnd cell_6t
Xbit_r36_c87 bl[87] br[87] wl[36] vdd gnd cell_6t
Xbit_r37_c87 bl[87] br[87] wl[37] vdd gnd cell_6t
Xbit_r38_c87 bl[87] br[87] wl[38] vdd gnd cell_6t
Xbit_r39_c87 bl[87] br[87] wl[39] vdd gnd cell_6t
Xbit_r40_c87 bl[87] br[87] wl[40] vdd gnd cell_6t
Xbit_r41_c87 bl[87] br[87] wl[41] vdd gnd cell_6t
Xbit_r42_c87 bl[87] br[87] wl[42] vdd gnd cell_6t
Xbit_r43_c87 bl[87] br[87] wl[43] vdd gnd cell_6t
Xbit_r44_c87 bl[87] br[87] wl[44] vdd gnd cell_6t
Xbit_r45_c87 bl[87] br[87] wl[45] vdd gnd cell_6t
Xbit_r46_c87 bl[87] br[87] wl[46] vdd gnd cell_6t
Xbit_r47_c87 bl[87] br[87] wl[47] vdd gnd cell_6t
Xbit_r48_c87 bl[87] br[87] wl[48] vdd gnd cell_6t
Xbit_r49_c87 bl[87] br[87] wl[49] vdd gnd cell_6t
Xbit_r50_c87 bl[87] br[87] wl[50] vdd gnd cell_6t
Xbit_r51_c87 bl[87] br[87] wl[51] vdd gnd cell_6t
Xbit_r52_c87 bl[87] br[87] wl[52] vdd gnd cell_6t
Xbit_r53_c87 bl[87] br[87] wl[53] vdd gnd cell_6t
Xbit_r54_c87 bl[87] br[87] wl[54] vdd gnd cell_6t
Xbit_r55_c87 bl[87] br[87] wl[55] vdd gnd cell_6t
Xbit_r56_c87 bl[87] br[87] wl[56] vdd gnd cell_6t
Xbit_r57_c87 bl[87] br[87] wl[57] vdd gnd cell_6t
Xbit_r58_c87 bl[87] br[87] wl[58] vdd gnd cell_6t
Xbit_r59_c87 bl[87] br[87] wl[59] vdd gnd cell_6t
Xbit_r60_c87 bl[87] br[87] wl[60] vdd gnd cell_6t
Xbit_r61_c87 bl[87] br[87] wl[61] vdd gnd cell_6t
Xbit_r62_c87 bl[87] br[87] wl[62] vdd gnd cell_6t
Xbit_r63_c87 bl[87] br[87] wl[63] vdd gnd cell_6t
Xbit_r64_c87 bl[87] br[87] wl[64] vdd gnd cell_6t
Xbit_r65_c87 bl[87] br[87] wl[65] vdd gnd cell_6t
Xbit_r66_c87 bl[87] br[87] wl[66] vdd gnd cell_6t
Xbit_r67_c87 bl[87] br[87] wl[67] vdd gnd cell_6t
Xbit_r68_c87 bl[87] br[87] wl[68] vdd gnd cell_6t
Xbit_r69_c87 bl[87] br[87] wl[69] vdd gnd cell_6t
Xbit_r70_c87 bl[87] br[87] wl[70] vdd gnd cell_6t
Xbit_r71_c87 bl[87] br[87] wl[71] vdd gnd cell_6t
Xbit_r72_c87 bl[87] br[87] wl[72] vdd gnd cell_6t
Xbit_r73_c87 bl[87] br[87] wl[73] vdd gnd cell_6t
Xbit_r74_c87 bl[87] br[87] wl[74] vdd gnd cell_6t
Xbit_r75_c87 bl[87] br[87] wl[75] vdd gnd cell_6t
Xbit_r76_c87 bl[87] br[87] wl[76] vdd gnd cell_6t
Xbit_r77_c87 bl[87] br[87] wl[77] vdd gnd cell_6t
Xbit_r78_c87 bl[87] br[87] wl[78] vdd gnd cell_6t
Xbit_r79_c87 bl[87] br[87] wl[79] vdd gnd cell_6t
Xbit_r80_c87 bl[87] br[87] wl[80] vdd gnd cell_6t
Xbit_r81_c87 bl[87] br[87] wl[81] vdd gnd cell_6t
Xbit_r82_c87 bl[87] br[87] wl[82] vdd gnd cell_6t
Xbit_r83_c87 bl[87] br[87] wl[83] vdd gnd cell_6t
Xbit_r84_c87 bl[87] br[87] wl[84] vdd gnd cell_6t
Xbit_r85_c87 bl[87] br[87] wl[85] vdd gnd cell_6t
Xbit_r86_c87 bl[87] br[87] wl[86] vdd gnd cell_6t
Xbit_r87_c87 bl[87] br[87] wl[87] vdd gnd cell_6t
Xbit_r88_c87 bl[87] br[87] wl[88] vdd gnd cell_6t
Xbit_r89_c87 bl[87] br[87] wl[89] vdd gnd cell_6t
Xbit_r90_c87 bl[87] br[87] wl[90] vdd gnd cell_6t
Xbit_r91_c87 bl[87] br[87] wl[91] vdd gnd cell_6t
Xbit_r92_c87 bl[87] br[87] wl[92] vdd gnd cell_6t
Xbit_r93_c87 bl[87] br[87] wl[93] vdd gnd cell_6t
Xbit_r94_c87 bl[87] br[87] wl[94] vdd gnd cell_6t
Xbit_r95_c87 bl[87] br[87] wl[95] vdd gnd cell_6t
Xbit_r96_c87 bl[87] br[87] wl[96] vdd gnd cell_6t
Xbit_r97_c87 bl[87] br[87] wl[97] vdd gnd cell_6t
Xbit_r98_c87 bl[87] br[87] wl[98] vdd gnd cell_6t
Xbit_r99_c87 bl[87] br[87] wl[99] vdd gnd cell_6t
Xbit_r100_c87 bl[87] br[87] wl[100] vdd gnd cell_6t
Xbit_r101_c87 bl[87] br[87] wl[101] vdd gnd cell_6t
Xbit_r102_c87 bl[87] br[87] wl[102] vdd gnd cell_6t
Xbit_r103_c87 bl[87] br[87] wl[103] vdd gnd cell_6t
Xbit_r104_c87 bl[87] br[87] wl[104] vdd gnd cell_6t
Xbit_r105_c87 bl[87] br[87] wl[105] vdd gnd cell_6t
Xbit_r106_c87 bl[87] br[87] wl[106] vdd gnd cell_6t
Xbit_r107_c87 bl[87] br[87] wl[107] vdd gnd cell_6t
Xbit_r108_c87 bl[87] br[87] wl[108] vdd gnd cell_6t
Xbit_r109_c87 bl[87] br[87] wl[109] vdd gnd cell_6t
Xbit_r110_c87 bl[87] br[87] wl[110] vdd gnd cell_6t
Xbit_r111_c87 bl[87] br[87] wl[111] vdd gnd cell_6t
Xbit_r112_c87 bl[87] br[87] wl[112] vdd gnd cell_6t
Xbit_r113_c87 bl[87] br[87] wl[113] vdd gnd cell_6t
Xbit_r114_c87 bl[87] br[87] wl[114] vdd gnd cell_6t
Xbit_r115_c87 bl[87] br[87] wl[115] vdd gnd cell_6t
Xbit_r116_c87 bl[87] br[87] wl[116] vdd gnd cell_6t
Xbit_r117_c87 bl[87] br[87] wl[117] vdd gnd cell_6t
Xbit_r118_c87 bl[87] br[87] wl[118] vdd gnd cell_6t
Xbit_r119_c87 bl[87] br[87] wl[119] vdd gnd cell_6t
Xbit_r120_c87 bl[87] br[87] wl[120] vdd gnd cell_6t
Xbit_r121_c87 bl[87] br[87] wl[121] vdd gnd cell_6t
Xbit_r122_c87 bl[87] br[87] wl[122] vdd gnd cell_6t
Xbit_r123_c87 bl[87] br[87] wl[123] vdd gnd cell_6t
Xbit_r124_c87 bl[87] br[87] wl[124] vdd gnd cell_6t
Xbit_r125_c87 bl[87] br[87] wl[125] vdd gnd cell_6t
Xbit_r126_c87 bl[87] br[87] wl[126] vdd gnd cell_6t
Xbit_r127_c87 bl[87] br[87] wl[127] vdd gnd cell_6t
Xbit_r128_c87 bl[87] br[87] wl[128] vdd gnd cell_6t
Xbit_r129_c87 bl[87] br[87] wl[129] vdd gnd cell_6t
Xbit_r130_c87 bl[87] br[87] wl[130] vdd gnd cell_6t
Xbit_r131_c87 bl[87] br[87] wl[131] vdd gnd cell_6t
Xbit_r132_c87 bl[87] br[87] wl[132] vdd gnd cell_6t
Xbit_r133_c87 bl[87] br[87] wl[133] vdd gnd cell_6t
Xbit_r134_c87 bl[87] br[87] wl[134] vdd gnd cell_6t
Xbit_r135_c87 bl[87] br[87] wl[135] vdd gnd cell_6t
Xbit_r136_c87 bl[87] br[87] wl[136] vdd gnd cell_6t
Xbit_r137_c87 bl[87] br[87] wl[137] vdd gnd cell_6t
Xbit_r138_c87 bl[87] br[87] wl[138] vdd gnd cell_6t
Xbit_r139_c87 bl[87] br[87] wl[139] vdd gnd cell_6t
Xbit_r140_c87 bl[87] br[87] wl[140] vdd gnd cell_6t
Xbit_r141_c87 bl[87] br[87] wl[141] vdd gnd cell_6t
Xbit_r142_c87 bl[87] br[87] wl[142] vdd gnd cell_6t
Xbit_r143_c87 bl[87] br[87] wl[143] vdd gnd cell_6t
Xbit_r144_c87 bl[87] br[87] wl[144] vdd gnd cell_6t
Xbit_r145_c87 bl[87] br[87] wl[145] vdd gnd cell_6t
Xbit_r146_c87 bl[87] br[87] wl[146] vdd gnd cell_6t
Xbit_r147_c87 bl[87] br[87] wl[147] vdd gnd cell_6t
Xbit_r148_c87 bl[87] br[87] wl[148] vdd gnd cell_6t
Xbit_r149_c87 bl[87] br[87] wl[149] vdd gnd cell_6t
Xbit_r150_c87 bl[87] br[87] wl[150] vdd gnd cell_6t
Xbit_r151_c87 bl[87] br[87] wl[151] vdd gnd cell_6t
Xbit_r152_c87 bl[87] br[87] wl[152] vdd gnd cell_6t
Xbit_r153_c87 bl[87] br[87] wl[153] vdd gnd cell_6t
Xbit_r154_c87 bl[87] br[87] wl[154] vdd gnd cell_6t
Xbit_r155_c87 bl[87] br[87] wl[155] vdd gnd cell_6t
Xbit_r156_c87 bl[87] br[87] wl[156] vdd gnd cell_6t
Xbit_r157_c87 bl[87] br[87] wl[157] vdd gnd cell_6t
Xbit_r158_c87 bl[87] br[87] wl[158] vdd gnd cell_6t
Xbit_r159_c87 bl[87] br[87] wl[159] vdd gnd cell_6t
Xbit_r160_c87 bl[87] br[87] wl[160] vdd gnd cell_6t
Xbit_r161_c87 bl[87] br[87] wl[161] vdd gnd cell_6t
Xbit_r162_c87 bl[87] br[87] wl[162] vdd gnd cell_6t
Xbit_r163_c87 bl[87] br[87] wl[163] vdd gnd cell_6t
Xbit_r164_c87 bl[87] br[87] wl[164] vdd gnd cell_6t
Xbit_r165_c87 bl[87] br[87] wl[165] vdd gnd cell_6t
Xbit_r166_c87 bl[87] br[87] wl[166] vdd gnd cell_6t
Xbit_r167_c87 bl[87] br[87] wl[167] vdd gnd cell_6t
Xbit_r168_c87 bl[87] br[87] wl[168] vdd gnd cell_6t
Xbit_r169_c87 bl[87] br[87] wl[169] vdd gnd cell_6t
Xbit_r170_c87 bl[87] br[87] wl[170] vdd gnd cell_6t
Xbit_r171_c87 bl[87] br[87] wl[171] vdd gnd cell_6t
Xbit_r172_c87 bl[87] br[87] wl[172] vdd gnd cell_6t
Xbit_r173_c87 bl[87] br[87] wl[173] vdd gnd cell_6t
Xbit_r174_c87 bl[87] br[87] wl[174] vdd gnd cell_6t
Xbit_r175_c87 bl[87] br[87] wl[175] vdd gnd cell_6t
Xbit_r176_c87 bl[87] br[87] wl[176] vdd gnd cell_6t
Xbit_r177_c87 bl[87] br[87] wl[177] vdd gnd cell_6t
Xbit_r178_c87 bl[87] br[87] wl[178] vdd gnd cell_6t
Xbit_r179_c87 bl[87] br[87] wl[179] vdd gnd cell_6t
Xbit_r180_c87 bl[87] br[87] wl[180] vdd gnd cell_6t
Xbit_r181_c87 bl[87] br[87] wl[181] vdd gnd cell_6t
Xbit_r182_c87 bl[87] br[87] wl[182] vdd gnd cell_6t
Xbit_r183_c87 bl[87] br[87] wl[183] vdd gnd cell_6t
Xbit_r184_c87 bl[87] br[87] wl[184] vdd gnd cell_6t
Xbit_r185_c87 bl[87] br[87] wl[185] vdd gnd cell_6t
Xbit_r186_c87 bl[87] br[87] wl[186] vdd gnd cell_6t
Xbit_r187_c87 bl[87] br[87] wl[187] vdd gnd cell_6t
Xbit_r188_c87 bl[87] br[87] wl[188] vdd gnd cell_6t
Xbit_r189_c87 bl[87] br[87] wl[189] vdd gnd cell_6t
Xbit_r190_c87 bl[87] br[87] wl[190] vdd gnd cell_6t
Xbit_r191_c87 bl[87] br[87] wl[191] vdd gnd cell_6t
Xbit_r192_c87 bl[87] br[87] wl[192] vdd gnd cell_6t
Xbit_r193_c87 bl[87] br[87] wl[193] vdd gnd cell_6t
Xbit_r194_c87 bl[87] br[87] wl[194] vdd gnd cell_6t
Xbit_r195_c87 bl[87] br[87] wl[195] vdd gnd cell_6t
Xbit_r196_c87 bl[87] br[87] wl[196] vdd gnd cell_6t
Xbit_r197_c87 bl[87] br[87] wl[197] vdd gnd cell_6t
Xbit_r198_c87 bl[87] br[87] wl[198] vdd gnd cell_6t
Xbit_r199_c87 bl[87] br[87] wl[199] vdd gnd cell_6t
Xbit_r200_c87 bl[87] br[87] wl[200] vdd gnd cell_6t
Xbit_r201_c87 bl[87] br[87] wl[201] vdd gnd cell_6t
Xbit_r202_c87 bl[87] br[87] wl[202] vdd gnd cell_6t
Xbit_r203_c87 bl[87] br[87] wl[203] vdd gnd cell_6t
Xbit_r204_c87 bl[87] br[87] wl[204] vdd gnd cell_6t
Xbit_r205_c87 bl[87] br[87] wl[205] vdd gnd cell_6t
Xbit_r206_c87 bl[87] br[87] wl[206] vdd gnd cell_6t
Xbit_r207_c87 bl[87] br[87] wl[207] vdd gnd cell_6t
Xbit_r208_c87 bl[87] br[87] wl[208] vdd gnd cell_6t
Xbit_r209_c87 bl[87] br[87] wl[209] vdd gnd cell_6t
Xbit_r210_c87 bl[87] br[87] wl[210] vdd gnd cell_6t
Xbit_r211_c87 bl[87] br[87] wl[211] vdd gnd cell_6t
Xbit_r212_c87 bl[87] br[87] wl[212] vdd gnd cell_6t
Xbit_r213_c87 bl[87] br[87] wl[213] vdd gnd cell_6t
Xbit_r214_c87 bl[87] br[87] wl[214] vdd gnd cell_6t
Xbit_r215_c87 bl[87] br[87] wl[215] vdd gnd cell_6t
Xbit_r216_c87 bl[87] br[87] wl[216] vdd gnd cell_6t
Xbit_r217_c87 bl[87] br[87] wl[217] vdd gnd cell_6t
Xbit_r218_c87 bl[87] br[87] wl[218] vdd gnd cell_6t
Xbit_r219_c87 bl[87] br[87] wl[219] vdd gnd cell_6t
Xbit_r220_c87 bl[87] br[87] wl[220] vdd gnd cell_6t
Xbit_r221_c87 bl[87] br[87] wl[221] vdd gnd cell_6t
Xbit_r222_c87 bl[87] br[87] wl[222] vdd gnd cell_6t
Xbit_r223_c87 bl[87] br[87] wl[223] vdd gnd cell_6t
Xbit_r224_c87 bl[87] br[87] wl[224] vdd gnd cell_6t
Xbit_r225_c87 bl[87] br[87] wl[225] vdd gnd cell_6t
Xbit_r226_c87 bl[87] br[87] wl[226] vdd gnd cell_6t
Xbit_r227_c87 bl[87] br[87] wl[227] vdd gnd cell_6t
Xbit_r228_c87 bl[87] br[87] wl[228] vdd gnd cell_6t
Xbit_r229_c87 bl[87] br[87] wl[229] vdd gnd cell_6t
Xbit_r230_c87 bl[87] br[87] wl[230] vdd gnd cell_6t
Xbit_r231_c87 bl[87] br[87] wl[231] vdd gnd cell_6t
Xbit_r232_c87 bl[87] br[87] wl[232] vdd gnd cell_6t
Xbit_r233_c87 bl[87] br[87] wl[233] vdd gnd cell_6t
Xbit_r234_c87 bl[87] br[87] wl[234] vdd gnd cell_6t
Xbit_r235_c87 bl[87] br[87] wl[235] vdd gnd cell_6t
Xbit_r236_c87 bl[87] br[87] wl[236] vdd gnd cell_6t
Xbit_r237_c87 bl[87] br[87] wl[237] vdd gnd cell_6t
Xbit_r238_c87 bl[87] br[87] wl[238] vdd gnd cell_6t
Xbit_r239_c87 bl[87] br[87] wl[239] vdd gnd cell_6t
Xbit_r240_c87 bl[87] br[87] wl[240] vdd gnd cell_6t
Xbit_r241_c87 bl[87] br[87] wl[241] vdd gnd cell_6t
Xbit_r242_c87 bl[87] br[87] wl[242] vdd gnd cell_6t
Xbit_r243_c87 bl[87] br[87] wl[243] vdd gnd cell_6t
Xbit_r244_c87 bl[87] br[87] wl[244] vdd gnd cell_6t
Xbit_r245_c87 bl[87] br[87] wl[245] vdd gnd cell_6t
Xbit_r246_c87 bl[87] br[87] wl[246] vdd gnd cell_6t
Xbit_r247_c87 bl[87] br[87] wl[247] vdd gnd cell_6t
Xbit_r248_c87 bl[87] br[87] wl[248] vdd gnd cell_6t
Xbit_r249_c87 bl[87] br[87] wl[249] vdd gnd cell_6t
Xbit_r250_c87 bl[87] br[87] wl[250] vdd gnd cell_6t
Xbit_r251_c87 bl[87] br[87] wl[251] vdd gnd cell_6t
Xbit_r252_c87 bl[87] br[87] wl[252] vdd gnd cell_6t
Xbit_r253_c87 bl[87] br[87] wl[253] vdd gnd cell_6t
Xbit_r254_c87 bl[87] br[87] wl[254] vdd gnd cell_6t
Xbit_r255_c87 bl[87] br[87] wl[255] vdd gnd cell_6t
Xbit_r256_c87 bl[87] br[87] wl[256] vdd gnd cell_6t
Xbit_r257_c87 bl[87] br[87] wl[257] vdd gnd cell_6t
Xbit_r258_c87 bl[87] br[87] wl[258] vdd gnd cell_6t
Xbit_r259_c87 bl[87] br[87] wl[259] vdd gnd cell_6t
Xbit_r260_c87 bl[87] br[87] wl[260] vdd gnd cell_6t
Xbit_r261_c87 bl[87] br[87] wl[261] vdd gnd cell_6t
Xbit_r262_c87 bl[87] br[87] wl[262] vdd gnd cell_6t
Xbit_r263_c87 bl[87] br[87] wl[263] vdd gnd cell_6t
Xbit_r264_c87 bl[87] br[87] wl[264] vdd gnd cell_6t
Xbit_r265_c87 bl[87] br[87] wl[265] vdd gnd cell_6t
Xbit_r266_c87 bl[87] br[87] wl[266] vdd gnd cell_6t
Xbit_r267_c87 bl[87] br[87] wl[267] vdd gnd cell_6t
Xbit_r268_c87 bl[87] br[87] wl[268] vdd gnd cell_6t
Xbit_r269_c87 bl[87] br[87] wl[269] vdd gnd cell_6t
Xbit_r270_c87 bl[87] br[87] wl[270] vdd gnd cell_6t
Xbit_r271_c87 bl[87] br[87] wl[271] vdd gnd cell_6t
Xbit_r272_c87 bl[87] br[87] wl[272] vdd gnd cell_6t
Xbit_r273_c87 bl[87] br[87] wl[273] vdd gnd cell_6t
Xbit_r274_c87 bl[87] br[87] wl[274] vdd gnd cell_6t
Xbit_r275_c87 bl[87] br[87] wl[275] vdd gnd cell_6t
Xbit_r276_c87 bl[87] br[87] wl[276] vdd gnd cell_6t
Xbit_r277_c87 bl[87] br[87] wl[277] vdd gnd cell_6t
Xbit_r278_c87 bl[87] br[87] wl[278] vdd gnd cell_6t
Xbit_r279_c87 bl[87] br[87] wl[279] vdd gnd cell_6t
Xbit_r280_c87 bl[87] br[87] wl[280] vdd gnd cell_6t
Xbit_r281_c87 bl[87] br[87] wl[281] vdd gnd cell_6t
Xbit_r282_c87 bl[87] br[87] wl[282] vdd gnd cell_6t
Xbit_r283_c87 bl[87] br[87] wl[283] vdd gnd cell_6t
Xbit_r284_c87 bl[87] br[87] wl[284] vdd gnd cell_6t
Xbit_r285_c87 bl[87] br[87] wl[285] vdd gnd cell_6t
Xbit_r286_c87 bl[87] br[87] wl[286] vdd gnd cell_6t
Xbit_r287_c87 bl[87] br[87] wl[287] vdd gnd cell_6t
Xbit_r288_c87 bl[87] br[87] wl[288] vdd gnd cell_6t
Xbit_r289_c87 bl[87] br[87] wl[289] vdd gnd cell_6t
Xbit_r290_c87 bl[87] br[87] wl[290] vdd gnd cell_6t
Xbit_r291_c87 bl[87] br[87] wl[291] vdd gnd cell_6t
Xbit_r292_c87 bl[87] br[87] wl[292] vdd gnd cell_6t
Xbit_r293_c87 bl[87] br[87] wl[293] vdd gnd cell_6t
Xbit_r294_c87 bl[87] br[87] wl[294] vdd gnd cell_6t
Xbit_r295_c87 bl[87] br[87] wl[295] vdd gnd cell_6t
Xbit_r296_c87 bl[87] br[87] wl[296] vdd gnd cell_6t
Xbit_r297_c87 bl[87] br[87] wl[297] vdd gnd cell_6t
Xbit_r298_c87 bl[87] br[87] wl[298] vdd gnd cell_6t
Xbit_r299_c87 bl[87] br[87] wl[299] vdd gnd cell_6t
Xbit_r300_c87 bl[87] br[87] wl[300] vdd gnd cell_6t
Xbit_r301_c87 bl[87] br[87] wl[301] vdd gnd cell_6t
Xbit_r302_c87 bl[87] br[87] wl[302] vdd gnd cell_6t
Xbit_r303_c87 bl[87] br[87] wl[303] vdd gnd cell_6t
Xbit_r304_c87 bl[87] br[87] wl[304] vdd gnd cell_6t
Xbit_r305_c87 bl[87] br[87] wl[305] vdd gnd cell_6t
Xbit_r306_c87 bl[87] br[87] wl[306] vdd gnd cell_6t
Xbit_r307_c87 bl[87] br[87] wl[307] vdd gnd cell_6t
Xbit_r308_c87 bl[87] br[87] wl[308] vdd gnd cell_6t
Xbit_r309_c87 bl[87] br[87] wl[309] vdd gnd cell_6t
Xbit_r310_c87 bl[87] br[87] wl[310] vdd gnd cell_6t
Xbit_r311_c87 bl[87] br[87] wl[311] vdd gnd cell_6t
Xbit_r312_c87 bl[87] br[87] wl[312] vdd gnd cell_6t
Xbit_r313_c87 bl[87] br[87] wl[313] vdd gnd cell_6t
Xbit_r314_c87 bl[87] br[87] wl[314] vdd gnd cell_6t
Xbit_r315_c87 bl[87] br[87] wl[315] vdd gnd cell_6t
Xbit_r316_c87 bl[87] br[87] wl[316] vdd gnd cell_6t
Xbit_r317_c87 bl[87] br[87] wl[317] vdd gnd cell_6t
Xbit_r318_c87 bl[87] br[87] wl[318] vdd gnd cell_6t
Xbit_r319_c87 bl[87] br[87] wl[319] vdd gnd cell_6t
Xbit_r320_c87 bl[87] br[87] wl[320] vdd gnd cell_6t
Xbit_r321_c87 bl[87] br[87] wl[321] vdd gnd cell_6t
Xbit_r322_c87 bl[87] br[87] wl[322] vdd gnd cell_6t
Xbit_r323_c87 bl[87] br[87] wl[323] vdd gnd cell_6t
Xbit_r324_c87 bl[87] br[87] wl[324] vdd gnd cell_6t
Xbit_r325_c87 bl[87] br[87] wl[325] vdd gnd cell_6t
Xbit_r326_c87 bl[87] br[87] wl[326] vdd gnd cell_6t
Xbit_r327_c87 bl[87] br[87] wl[327] vdd gnd cell_6t
Xbit_r328_c87 bl[87] br[87] wl[328] vdd gnd cell_6t
Xbit_r329_c87 bl[87] br[87] wl[329] vdd gnd cell_6t
Xbit_r330_c87 bl[87] br[87] wl[330] vdd gnd cell_6t
Xbit_r331_c87 bl[87] br[87] wl[331] vdd gnd cell_6t
Xbit_r332_c87 bl[87] br[87] wl[332] vdd gnd cell_6t
Xbit_r333_c87 bl[87] br[87] wl[333] vdd gnd cell_6t
Xbit_r334_c87 bl[87] br[87] wl[334] vdd gnd cell_6t
Xbit_r335_c87 bl[87] br[87] wl[335] vdd gnd cell_6t
Xbit_r336_c87 bl[87] br[87] wl[336] vdd gnd cell_6t
Xbit_r337_c87 bl[87] br[87] wl[337] vdd gnd cell_6t
Xbit_r338_c87 bl[87] br[87] wl[338] vdd gnd cell_6t
Xbit_r339_c87 bl[87] br[87] wl[339] vdd gnd cell_6t
Xbit_r340_c87 bl[87] br[87] wl[340] vdd gnd cell_6t
Xbit_r341_c87 bl[87] br[87] wl[341] vdd gnd cell_6t
Xbit_r342_c87 bl[87] br[87] wl[342] vdd gnd cell_6t
Xbit_r343_c87 bl[87] br[87] wl[343] vdd gnd cell_6t
Xbit_r344_c87 bl[87] br[87] wl[344] vdd gnd cell_6t
Xbit_r345_c87 bl[87] br[87] wl[345] vdd gnd cell_6t
Xbit_r346_c87 bl[87] br[87] wl[346] vdd gnd cell_6t
Xbit_r347_c87 bl[87] br[87] wl[347] vdd gnd cell_6t
Xbit_r348_c87 bl[87] br[87] wl[348] vdd gnd cell_6t
Xbit_r349_c87 bl[87] br[87] wl[349] vdd gnd cell_6t
Xbit_r350_c87 bl[87] br[87] wl[350] vdd gnd cell_6t
Xbit_r351_c87 bl[87] br[87] wl[351] vdd gnd cell_6t
Xbit_r352_c87 bl[87] br[87] wl[352] vdd gnd cell_6t
Xbit_r353_c87 bl[87] br[87] wl[353] vdd gnd cell_6t
Xbit_r354_c87 bl[87] br[87] wl[354] vdd gnd cell_6t
Xbit_r355_c87 bl[87] br[87] wl[355] vdd gnd cell_6t
Xbit_r356_c87 bl[87] br[87] wl[356] vdd gnd cell_6t
Xbit_r357_c87 bl[87] br[87] wl[357] vdd gnd cell_6t
Xbit_r358_c87 bl[87] br[87] wl[358] vdd gnd cell_6t
Xbit_r359_c87 bl[87] br[87] wl[359] vdd gnd cell_6t
Xbit_r360_c87 bl[87] br[87] wl[360] vdd gnd cell_6t
Xbit_r361_c87 bl[87] br[87] wl[361] vdd gnd cell_6t
Xbit_r362_c87 bl[87] br[87] wl[362] vdd gnd cell_6t
Xbit_r363_c87 bl[87] br[87] wl[363] vdd gnd cell_6t
Xbit_r364_c87 bl[87] br[87] wl[364] vdd gnd cell_6t
Xbit_r365_c87 bl[87] br[87] wl[365] vdd gnd cell_6t
Xbit_r366_c87 bl[87] br[87] wl[366] vdd gnd cell_6t
Xbit_r367_c87 bl[87] br[87] wl[367] vdd gnd cell_6t
Xbit_r368_c87 bl[87] br[87] wl[368] vdd gnd cell_6t
Xbit_r369_c87 bl[87] br[87] wl[369] vdd gnd cell_6t
Xbit_r370_c87 bl[87] br[87] wl[370] vdd gnd cell_6t
Xbit_r371_c87 bl[87] br[87] wl[371] vdd gnd cell_6t
Xbit_r372_c87 bl[87] br[87] wl[372] vdd gnd cell_6t
Xbit_r373_c87 bl[87] br[87] wl[373] vdd gnd cell_6t
Xbit_r374_c87 bl[87] br[87] wl[374] vdd gnd cell_6t
Xbit_r375_c87 bl[87] br[87] wl[375] vdd gnd cell_6t
Xbit_r376_c87 bl[87] br[87] wl[376] vdd gnd cell_6t
Xbit_r377_c87 bl[87] br[87] wl[377] vdd gnd cell_6t
Xbit_r378_c87 bl[87] br[87] wl[378] vdd gnd cell_6t
Xbit_r379_c87 bl[87] br[87] wl[379] vdd gnd cell_6t
Xbit_r380_c87 bl[87] br[87] wl[380] vdd gnd cell_6t
Xbit_r381_c87 bl[87] br[87] wl[381] vdd gnd cell_6t
Xbit_r382_c87 bl[87] br[87] wl[382] vdd gnd cell_6t
Xbit_r383_c87 bl[87] br[87] wl[383] vdd gnd cell_6t
Xbit_r384_c87 bl[87] br[87] wl[384] vdd gnd cell_6t
Xbit_r385_c87 bl[87] br[87] wl[385] vdd gnd cell_6t
Xbit_r386_c87 bl[87] br[87] wl[386] vdd gnd cell_6t
Xbit_r387_c87 bl[87] br[87] wl[387] vdd gnd cell_6t
Xbit_r388_c87 bl[87] br[87] wl[388] vdd gnd cell_6t
Xbit_r389_c87 bl[87] br[87] wl[389] vdd gnd cell_6t
Xbit_r390_c87 bl[87] br[87] wl[390] vdd gnd cell_6t
Xbit_r391_c87 bl[87] br[87] wl[391] vdd gnd cell_6t
Xbit_r392_c87 bl[87] br[87] wl[392] vdd gnd cell_6t
Xbit_r393_c87 bl[87] br[87] wl[393] vdd gnd cell_6t
Xbit_r394_c87 bl[87] br[87] wl[394] vdd gnd cell_6t
Xbit_r395_c87 bl[87] br[87] wl[395] vdd gnd cell_6t
Xbit_r396_c87 bl[87] br[87] wl[396] vdd gnd cell_6t
Xbit_r397_c87 bl[87] br[87] wl[397] vdd gnd cell_6t
Xbit_r398_c87 bl[87] br[87] wl[398] vdd gnd cell_6t
Xbit_r399_c87 bl[87] br[87] wl[399] vdd gnd cell_6t
Xbit_r400_c87 bl[87] br[87] wl[400] vdd gnd cell_6t
Xbit_r401_c87 bl[87] br[87] wl[401] vdd gnd cell_6t
Xbit_r402_c87 bl[87] br[87] wl[402] vdd gnd cell_6t
Xbit_r403_c87 bl[87] br[87] wl[403] vdd gnd cell_6t
Xbit_r404_c87 bl[87] br[87] wl[404] vdd gnd cell_6t
Xbit_r405_c87 bl[87] br[87] wl[405] vdd gnd cell_6t
Xbit_r406_c87 bl[87] br[87] wl[406] vdd gnd cell_6t
Xbit_r407_c87 bl[87] br[87] wl[407] vdd gnd cell_6t
Xbit_r408_c87 bl[87] br[87] wl[408] vdd gnd cell_6t
Xbit_r409_c87 bl[87] br[87] wl[409] vdd gnd cell_6t
Xbit_r410_c87 bl[87] br[87] wl[410] vdd gnd cell_6t
Xbit_r411_c87 bl[87] br[87] wl[411] vdd gnd cell_6t
Xbit_r412_c87 bl[87] br[87] wl[412] vdd gnd cell_6t
Xbit_r413_c87 bl[87] br[87] wl[413] vdd gnd cell_6t
Xbit_r414_c87 bl[87] br[87] wl[414] vdd gnd cell_6t
Xbit_r415_c87 bl[87] br[87] wl[415] vdd gnd cell_6t
Xbit_r416_c87 bl[87] br[87] wl[416] vdd gnd cell_6t
Xbit_r417_c87 bl[87] br[87] wl[417] vdd gnd cell_6t
Xbit_r418_c87 bl[87] br[87] wl[418] vdd gnd cell_6t
Xbit_r419_c87 bl[87] br[87] wl[419] vdd gnd cell_6t
Xbit_r420_c87 bl[87] br[87] wl[420] vdd gnd cell_6t
Xbit_r421_c87 bl[87] br[87] wl[421] vdd gnd cell_6t
Xbit_r422_c87 bl[87] br[87] wl[422] vdd gnd cell_6t
Xbit_r423_c87 bl[87] br[87] wl[423] vdd gnd cell_6t
Xbit_r424_c87 bl[87] br[87] wl[424] vdd gnd cell_6t
Xbit_r425_c87 bl[87] br[87] wl[425] vdd gnd cell_6t
Xbit_r426_c87 bl[87] br[87] wl[426] vdd gnd cell_6t
Xbit_r427_c87 bl[87] br[87] wl[427] vdd gnd cell_6t
Xbit_r428_c87 bl[87] br[87] wl[428] vdd gnd cell_6t
Xbit_r429_c87 bl[87] br[87] wl[429] vdd gnd cell_6t
Xbit_r430_c87 bl[87] br[87] wl[430] vdd gnd cell_6t
Xbit_r431_c87 bl[87] br[87] wl[431] vdd gnd cell_6t
Xbit_r432_c87 bl[87] br[87] wl[432] vdd gnd cell_6t
Xbit_r433_c87 bl[87] br[87] wl[433] vdd gnd cell_6t
Xbit_r434_c87 bl[87] br[87] wl[434] vdd gnd cell_6t
Xbit_r435_c87 bl[87] br[87] wl[435] vdd gnd cell_6t
Xbit_r436_c87 bl[87] br[87] wl[436] vdd gnd cell_6t
Xbit_r437_c87 bl[87] br[87] wl[437] vdd gnd cell_6t
Xbit_r438_c87 bl[87] br[87] wl[438] vdd gnd cell_6t
Xbit_r439_c87 bl[87] br[87] wl[439] vdd gnd cell_6t
Xbit_r440_c87 bl[87] br[87] wl[440] vdd gnd cell_6t
Xbit_r441_c87 bl[87] br[87] wl[441] vdd gnd cell_6t
Xbit_r442_c87 bl[87] br[87] wl[442] vdd gnd cell_6t
Xbit_r443_c87 bl[87] br[87] wl[443] vdd gnd cell_6t
Xbit_r444_c87 bl[87] br[87] wl[444] vdd gnd cell_6t
Xbit_r445_c87 bl[87] br[87] wl[445] vdd gnd cell_6t
Xbit_r446_c87 bl[87] br[87] wl[446] vdd gnd cell_6t
Xbit_r447_c87 bl[87] br[87] wl[447] vdd gnd cell_6t
Xbit_r448_c87 bl[87] br[87] wl[448] vdd gnd cell_6t
Xbit_r449_c87 bl[87] br[87] wl[449] vdd gnd cell_6t
Xbit_r450_c87 bl[87] br[87] wl[450] vdd gnd cell_6t
Xbit_r451_c87 bl[87] br[87] wl[451] vdd gnd cell_6t
Xbit_r452_c87 bl[87] br[87] wl[452] vdd gnd cell_6t
Xbit_r453_c87 bl[87] br[87] wl[453] vdd gnd cell_6t
Xbit_r454_c87 bl[87] br[87] wl[454] vdd gnd cell_6t
Xbit_r455_c87 bl[87] br[87] wl[455] vdd gnd cell_6t
Xbit_r456_c87 bl[87] br[87] wl[456] vdd gnd cell_6t
Xbit_r457_c87 bl[87] br[87] wl[457] vdd gnd cell_6t
Xbit_r458_c87 bl[87] br[87] wl[458] vdd gnd cell_6t
Xbit_r459_c87 bl[87] br[87] wl[459] vdd gnd cell_6t
Xbit_r460_c87 bl[87] br[87] wl[460] vdd gnd cell_6t
Xbit_r461_c87 bl[87] br[87] wl[461] vdd gnd cell_6t
Xbit_r462_c87 bl[87] br[87] wl[462] vdd gnd cell_6t
Xbit_r463_c87 bl[87] br[87] wl[463] vdd gnd cell_6t
Xbit_r464_c87 bl[87] br[87] wl[464] vdd gnd cell_6t
Xbit_r465_c87 bl[87] br[87] wl[465] vdd gnd cell_6t
Xbit_r466_c87 bl[87] br[87] wl[466] vdd gnd cell_6t
Xbit_r467_c87 bl[87] br[87] wl[467] vdd gnd cell_6t
Xbit_r468_c87 bl[87] br[87] wl[468] vdd gnd cell_6t
Xbit_r469_c87 bl[87] br[87] wl[469] vdd gnd cell_6t
Xbit_r470_c87 bl[87] br[87] wl[470] vdd gnd cell_6t
Xbit_r471_c87 bl[87] br[87] wl[471] vdd gnd cell_6t
Xbit_r472_c87 bl[87] br[87] wl[472] vdd gnd cell_6t
Xbit_r473_c87 bl[87] br[87] wl[473] vdd gnd cell_6t
Xbit_r474_c87 bl[87] br[87] wl[474] vdd gnd cell_6t
Xbit_r475_c87 bl[87] br[87] wl[475] vdd gnd cell_6t
Xbit_r476_c87 bl[87] br[87] wl[476] vdd gnd cell_6t
Xbit_r477_c87 bl[87] br[87] wl[477] vdd gnd cell_6t
Xbit_r478_c87 bl[87] br[87] wl[478] vdd gnd cell_6t
Xbit_r479_c87 bl[87] br[87] wl[479] vdd gnd cell_6t
Xbit_r480_c87 bl[87] br[87] wl[480] vdd gnd cell_6t
Xbit_r481_c87 bl[87] br[87] wl[481] vdd gnd cell_6t
Xbit_r482_c87 bl[87] br[87] wl[482] vdd gnd cell_6t
Xbit_r483_c87 bl[87] br[87] wl[483] vdd gnd cell_6t
Xbit_r484_c87 bl[87] br[87] wl[484] vdd gnd cell_6t
Xbit_r485_c87 bl[87] br[87] wl[485] vdd gnd cell_6t
Xbit_r486_c87 bl[87] br[87] wl[486] vdd gnd cell_6t
Xbit_r487_c87 bl[87] br[87] wl[487] vdd gnd cell_6t
Xbit_r488_c87 bl[87] br[87] wl[488] vdd gnd cell_6t
Xbit_r489_c87 bl[87] br[87] wl[489] vdd gnd cell_6t
Xbit_r490_c87 bl[87] br[87] wl[490] vdd gnd cell_6t
Xbit_r491_c87 bl[87] br[87] wl[491] vdd gnd cell_6t
Xbit_r492_c87 bl[87] br[87] wl[492] vdd gnd cell_6t
Xbit_r493_c87 bl[87] br[87] wl[493] vdd gnd cell_6t
Xbit_r494_c87 bl[87] br[87] wl[494] vdd gnd cell_6t
Xbit_r495_c87 bl[87] br[87] wl[495] vdd gnd cell_6t
Xbit_r496_c87 bl[87] br[87] wl[496] vdd gnd cell_6t
Xbit_r497_c87 bl[87] br[87] wl[497] vdd gnd cell_6t
Xbit_r498_c87 bl[87] br[87] wl[498] vdd gnd cell_6t
Xbit_r499_c87 bl[87] br[87] wl[499] vdd gnd cell_6t
Xbit_r500_c87 bl[87] br[87] wl[500] vdd gnd cell_6t
Xbit_r501_c87 bl[87] br[87] wl[501] vdd gnd cell_6t
Xbit_r502_c87 bl[87] br[87] wl[502] vdd gnd cell_6t
Xbit_r503_c87 bl[87] br[87] wl[503] vdd gnd cell_6t
Xbit_r504_c87 bl[87] br[87] wl[504] vdd gnd cell_6t
Xbit_r505_c87 bl[87] br[87] wl[505] vdd gnd cell_6t
Xbit_r506_c87 bl[87] br[87] wl[506] vdd gnd cell_6t
Xbit_r507_c87 bl[87] br[87] wl[507] vdd gnd cell_6t
Xbit_r508_c87 bl[87] br[87] wl[508] vdd gnd cell_6t
Xbit_r509_c87 bl[87] br[87] wl[509] vdd gnd cell_6t
Xbit_r510_c87 bl[87] br[87] wl[510] vdd gnd cell_6t
Xbit_r511_c87 bl[87] br[87] wl[511] vdd gnd cell_6t
Xbit_r0_c88 bl[88] br[88] wl[0] vdd gnd cell_6t
Xbit_r1_c88 bl[88] br[88] wl[1] vdd gnd cell_6t
Xbit_r2_c88 bl[88] br[88] wl[2] vdd gnd cell_6t
Xbit_r3_c88 bl[88] br[88] wl[3] vdd gnd cell_6t
Xbit_r4_c88 bl[88] br[88] wl[4] vdd gnd cell_6t
Xbit_r5_c88 bl[88] br[88] wl[5] vdd gnd cell_6t
Xbit_r6_c88 bl[88] br[88] wl[6] vdd gnd cell_6t
Xbit_r7_c88 bl[88] br[88] wl[7] vdd gnd cell_6t
Xbit_r8_c88 bl[88] br[88] wl[8] vdd gnd cell_6t
Xbit_r9_c88 bl[88] br[88] wl[9] vdd gnd cell_6t
Xbit_r10_c88 bl[88] br[88] wl[10] vdd gnd cell_6t
Xbit_r11_c88 bl[88] br[88] wl[11] vdd gnd cell_6t
Xbit_r12_c88 bl[88] br[88] wl[12] vdd gnd cell_6t
Xbit_r13_c88 bl[88] br[88] wl[13] vdd gnd cell_6t
Xbit_r14_c88 bl[88] br[88] wl[14] vdd gnd cell_6t
Xbit_r15_c88 bl[88] br[88] wl[15] vdd gnd cell_6t
Xbit_r16_c88 bl[88] br[88] wl[16] vdd gnd cell_6t
Xbit_r17_c88 bl[88] br[88] wl[17] vdd gnd cell_6t
Xbit_r18_c88 bl[88] br[88] wl[18] vdd gnd cell_6t
Xbit_r19_c88 bl[88] br[88] wl[19] vdd gnd cell_6t
Xbit_r20_c88 bl[88] br[88] wl[20] vdd gnd cell_6t
Xbit_r21_c88 bl[88] br[88] wl[21] vdd gnd cell_6t
Xbit_r22_c88 bl[88] br[88] wl[22] vdd gnd cell_6t
Xbit_r23_c88 bl[88] br[88] wl[23] vdd gnd cell_6t
Xbit_r24_c88 bl[88] br[88] wl[24] vdd gnd cell_6t
Xbit_r25_c88 bl[88] br[88] wl[25] vdd gnd cell_6t
Xbit_r26_c88 bl[88] br[88] wl[26] vdd gnd cell_6t
Xbit_r27_c88 bl[88] br[88] wl[27] vdd gnd cell_6t
Xbit_r28_c88 bl[88] br[88] wl[28] vdd gnd cell_6t
Xbit_r29_c88 bl[88] br[88] wl[29] vdd gnd cell_6t
Xbit_r30_c88 bl[88] br[88] wl[30] vdd gnd cell_6t
Xbit_r31_c88 bl[88] br[88] wl[31] vdd gnd cell_6t
Xbit_r32_c88 bl[88] br[88] wl[32] vdd gnd cell_6t
Xbit_r33_c88 bl[88] br[88] wl[33] vdd gnd cell_6t
Xbit_r34_c88 bl[88] br[88] wl[34] vdd gnd cell_6t
Xbit_r35_c88 bl[88] br[88] wl[35] vdd gnd cell_6t
Xbit_r36_c88 bl[88] br[88] wl[36] vdd gnd cell_6t
Xbit_r37_c88 bl[88] br[88] wl[37] vdd gnd cell_6t
Xbit_r38_c88 bl[88] br[88] wl[38] vdd gnd cell_6t
Xbit_r39_c88 bl[88] br[88] wl[39] vdd gnd cell_6t
Xbit_r40_c88 bl[88] br[88] wl[40] vdd gnd cell_6t
Xbit_r41_c88 bl[88] br[88] wl[41] vdd gnd cell_6t
Xbit_r42_c88 bl[88] br[88] wl[42] vdd gnd cell_6t
Xbit_r43_c88 bl[88] br[88] wl[43] vdd gnd cell_6t
Xbit_r44_c88 bl[88] br[88] wl[44] vdd gnd cell_6t
Xbit_r45_c88 bl[88] br[88] wl[45] vdd gnd cell_6t
Xbit_r46_c88 bl[88] br[88] wl[46] vdd gnd cell_6t
Xbit_r47_c88 bl[88] br[88] wl[47] vdd gnd cell_6t
Xbit_r48_c88 bl[88] br[88] wl[48] vdd gnd cell_6t
Xbit_r49_c88 bl[88] br[88] wl[49] vdd gnd cell_6t
Xbit_r50_c88 bl[88] br[88] wl[50] vdd gnd cell_6t
Xbit_r51_c88 bl[88] br[88] wl[51] vdd gnd cell_6t
Xbit_r52_c88 bl[88] br[88] wl[52] vdd gnd cell_6t
Xbit_r53_c88 bl[88] br[88] wl[53] vdd gnd cell_6t
Xbit_r54_c88 bl[88] br[88] wl[54] vdd gnd cell_6t
Xbit_r55_c88 bl[88] br[88] wl[55] vdd gnd cell_6t
Xbit_r56_c88 bl[88] br[88] wl[56] vdd gnd cell_6t
Xbit_r57_c88 bl[88] br[88] wl[57] vdd gnd cell_6t
Xbit_r58_c88 bl[88] br[88] wl[58] vdd gnd cell_6t
Xbit_r59_c88 bl[88] br[88] wl[59] vdd gnd cell_6t
Xbit_r60_c88 bl[88] br[88] wl[60] vdd gnd cell_6t
Xbit_r61_c88 bl[88] br[88] wl[61] vdd gnd cell_6t
Xbit_r62_c88 bl[88] br[88] wl[62] vdd gnd cell_6t
Xbit_r63_c88 bl[88] br[88] wl[63] vdd gnd cell_6t
Xbit_r64_c88 bl[88] br[88] wl[64] vdd gnd cell_6t
Xbit_r65_c88 bl[88] br[88] wl[65] vdd gnd cell_6t
Xbit_r66_c88 bl[88] br[88] wl[66] vdd gnd cell_6t
Xbit_r67_c88 bl[88] br[88] wl[67] vdd gnd cell_6t
Xbit_r68_c88 bl[88] br[88] wl[68] vdd gnd cell_6t
Xbit_r69_c88 bl[88] br[88] wl[69] vdd gnd cell_6t
Xbit_r70_c88 bl[88] br[88] wl[70] vdd gnd cell_6t
Xbit_r71_c88 bl[88] br[88] wl[71] vdd gnd cell_6t
Xbit_r72_c88 bl[88] br[88] wl[72] vdd gnd cell_6t
Xbit_r73_c88 bl[88] br[88] wl[73] vdd gnd cell_6t
Xbit_r74_c88 bl[88] br[88] wl[74] vdd gnd cell_6t
Xbit_r75_c88 bl[88] br[88] wl[75] vdd gnd cell_6t
Xbit_r76_c88 bl[88] br[88] wl[76] vdd gnd cell_6t
Xbit_r77_c88 bl[88] br[88] wl[77] vdd gnd cell_6t
Xbit_r78_c88 bl[88] br[88] wl[78] vdd gnd cell_6t
Xbit_r79_c88 bl[88] br[88] wl[79] vdd gnd cell_6t
Xbit_r80_c88 bl[88] br[88] wl[80] vdd gnd cell_6t
Xbit_r81_c88 bl[88] br[88] wl[81] vdd gnd cell_6t
Xbit_r82_c88 bl[88] br[88] wl[82] vdd gnd cell_6t
Xbit_r83_c88 bl[88] br[88] wl[83] vdd gnd cell_6t
Xbit_r84_c88 bl[88] br[88] wl[84] vdd gnd cell_6t
Xbit_r85_c88 bl[88] br[88] wl[85] vdd gnd cell_6t
Xbit_r86_c88 bl[88] br[88] wl[86] vdd gnd cell_6t
Xbit_r87_c88 bl[88] br[88] wl[87] vdd gnd cell_6t
Xbit_r88_c88 bl[88] br[88] wl[88] vdd gnd cell_6t
Xbit_r89_c88 bl[88] br[88] wl[89] vdd gnd cell_6t
Xbit_r90_c88 bl[88] br[88] wl[90] vdd gnd cell_6t
Xbit_r91_c88 bl[88] br[88] wl[91] vdd gnd cell_6t
Xbit_r92_c88 bl[88] br[88] wl[92] vdd gnd cell_6t
Xbit_r93_c88 bl[88] br[88] wl[93] vdd gnd cell_6t
Xbit_r94_c88 bl[88] br[88] wl[94] vdd gnd cell_6t
Xbit_r95_c88 bl[88] br[88] wl[95] vdd gnd cell_6t
Xbit_r96_c88 bl[88] br[88] wl[96] vdd gnd cell_6t
Xbit_r97_c88 bl[88] br[88] wl[97] vdd gnd cell_6t
Xbit_r98_c88 bl[88] br[88] wl[98] vdd gnd cell_6t
Xbit_r99_c88 bl[88] br[88] wl[99] vdd gnd cell_6t
Xbit_r100_c88 bl[88] br[88] wl[100] vdd gnd cell_6t
Xbit_r101_c88 bl[88] br[88] wl[101] vdd gnd cell_6t
Xbit_r102_c88 bl[88] br[88] wl[102] vdd gnd cell_6t
Xbit_r103_c88 bl[88] br[88] wl[103] vdd gnd cell_6t
Xbit_r104_c88 bl[88] br[88] wl[104] vdd gnd cell_6t
Xbit_r105_c88 bl[88] br[88] wl[105] vdd gnd cell_6t
Xbit_r106_c88 bl[88] br[88] wl[106] vdd gnd cell_6t
Xbit_r107_c88 bl[88] br[88] wl[107] vdd gnd cell_6t
Xbit_r108_c88 bl[88] br[88] wl[108] vdd gnd cell_6t
Xbit_r109_c88 bl[88] br[88] wl[109] vdd gnd cell_6t
Xbit_r110_c88 bl[88] br[88] wl[110] vdd gnd cell_6t
Xbit_r111_c88 bl[88] br[88] wl[111] vdd gnd cell_6t
Xbit_r112_c88 bl[88] br[88] wl[112] vdd gnd cell_6t
Xbit_r113_c88 bl[88] br[88] wl[113] vdd gnd cell_6t
Xbit_r114_c88 bl[88] br[88] wl[114] vdd gnd cell_6t
Xbit_r115_c88 bl[88] br[88] wl[115] vdd gnd cell_6t
Xbit_r116_c88 bl[88] br[88] wl[116] vdd gnd cell_6t
Xbit_r117_c88 bl[88] br[88] wl[117] vdd gnd cell_6t
Xbit_r118_c88 bl[88] br[88] wl[118] vdd gnd cell_6t
Xbit_r119_c88 bl[88] br[88] wl[119] vdd gnd cell_6t
Xbit_r120_c88 bl[88] br[88] wl[120] vdd gnd cell_6t
Xbit_r121_c88 bl[88] br[88] wl[121] vdd gnd cell_6t
Xbit_r122_c88 bl[88] br[88] wl[122] vdd gnd cell_6t
Xbit_r123_c88 bl[88] br[88] wl[123] vdd gnd cell_6t
Xbit_r124_c88 bl[88] br[88] wl[124] vdd gnd cell_6t
Xbit_r125_c88 bl[88] br[88] wl[125] vdd gnd cell_6t
Xbit_r126_c88 bl[88] br[88] wl[126] vdd gnd cell_6t
Xbit_r127_c88 bl[88] br[88] wl[127] vdd gnd cell_6t
Xbit_r128_c88 bl[88] br[88] wl[128] vdd gnd cell_6t
Xbit_r129_c88 bl[88] br[88] wl[129] vdd gnd cell_6t
Xbit_r130_c88 bl[88] br[88] wl[130] vdd gnd cell_6t
Xbit_r131_c88 bl[88] br[88] wl[131] vdd gnd cell_6t
Xbit_r132_c88 bl[88] br[88] wl[132] vdd gnd cell_6t
Xbit_r133_c88 bl[88] br[88] wl[133] vdd gnd cell_6t
Xbit_r134_c88 bl[88] br[88] wl[134] vdd gnd cell_6t
Xbit_r135_c88 bl[88] br[88] wl[135] vdd gnd cell_6t
Xbit_r136_c88 bl[88] br[88] wl[136] vdd gnd cell_6t
Xbit_r137_c88 bl[88] br[88] wl[137] vdd gnd cell_6t
Xbit_r138_c88 bl[88] br[88] wl[138] vdd gnd cell_6t
Xbit_r139_c88 bl[88] br[88] wl[139] vdd gnd cell_6t
Xbit_r140_c88 bl[88] br[88] wl[140] vdd gnd cell_6t
Xbit_r141_c88 bl[88] br[88] wl[141] vdd gnd cell_6t
Xbit_r142_c88 bl[88] br[88] wl[142] vdd gnd cell_6t
Xbit_r143_c88 bl[88] br[88] wl[143] vdd gnd cell_6t
Xbit_r144_c88 bl[88] br[88] wl[144] vdd gnd cell_6t
Xbit_r145_c88 bl[88] br[88] wl[145] vdd gnd cell_6t
Xbit_r146_c88 bl[88] br[88] wl[146] vdd gnd cell_6t
Xbit_r147_c88 bl[88] br[88] wl[147] vdd gnd cell_6t
Xbit_r148_c88 bl[88] br[88] wl[148] vdd gnd cell_6t
Xbit_r149_c88 bl[88] br[88] wl[149] vdd gnd cell_6t
Xbit_r150_c88 bl[88] br[88] wl[150] vdd gnd cell_6t
Xbit_r151_c88 bl[88] br[88] wl[151] vdd gnd cell_6t
Xbit_r152_c88 bl[88] br[88] wl[152] vdd gnd cell_6t
Xbit_r153_c88 bl[88] br[88] wl[153] vdd gnd cell_6t
Xbit_r154_c88 bl[88] br[88] wl[154] vdd gnd cell_6t
Xbit_r155_c88 bl[88] br[88] wl[155] vdd gnd cell_6t
Xbit_r156_c88 bl[88] br[88] wl[156] vdd gnd cell_6t
Xbit_r157_c88 bl[88] br[88] wl[157] vdd gnd cell_6t
Xbit_r158_c88 bl[88] br[88] wl[158] vdd gnd cell_6t
Xbit_r159_c88 bl[88] br[88] wl[159] vdd gnd cell_6t
Xbit_r160_c88 bl[88] br[88] wl[160] vdd gnd cell_6t
Xbit_r161_c88 bl[88] br[88] wl[161] vdd gnd cell_6t
Xbit_r162_c88 bl[88] br[88] wl[162] vdd gnd cell_6t
Xbit_r163_c88 bl[88] br[88] wl[163] vdd gnd cell_6t
Xbit_r164_c88 bl[88] br[88] wl[164] vdd gnd cell_6t
Xbit_r165_c88 bl[88] br[88] wl[165] vdd gnd cell_6t
Xbit_r166_c88 bl[88] br[88] wl[166] vdd gnd cell_6t
Xbit_r167_c88 bl[88] br[88] wl[167] vdd gnd cell_6t
Xbit_r168_c88 bl[88] br[88] wl[168] vdd gnd cell_6t
Xbit_r169_c88 bl[88] br[88] wl[169] vdd gnd cell_6t
Xbit_r170_c88 bl[88] br[88] wl[170] vdd gnd cell_6t
Xbit_r171_c88 bl[88] br[88] wl[171] vdd gnd cell_6t
Xbit_r172_c88 bl[88] br[88] wl[172] vdd gnd cell_6t
Xbit_r173_c88 bl[88] br[88] wl[173] vdd gnd cell_6t
Xbit_r174_c88 bl[88] br[88] wl[174] vdd gnd cell_6t
Xbit_r175_c88 bl[88] br[88] wl[175] vdd gnd cell_6t
Xbit_r176_c88 bl[88] br[88] wl[176] vdd gnd cell_6t
Xbit_r177_c88 bl[88] br[88] wl[177] vdd gnd cell_6t
Xbit_r178_c88 bl[88] br[88] wl[178] vdd gnd cell_6t
Xbit_r179_c88 bl[88] br[88] wl[179] vdd gnd cell_6t
Xbit_r180_c88 bl[88] br[88] wl[180] vdd gnd cell_6t
Xbit_r181_c88 bl[88] br[88] wl[181] vdd gnd cell_6t
Xbit_r182_c88 bl[88] br[88] wl[182] vdd gnd cell_6t
Xbit_r183_c88 bl[88] br[88] wl[183] vdd gnd cell_6t
Xbit_r184_c88 bl[88] br[88] wl[184] vdd gnd cell_6t
Xbit_r185_c88 bl[88] br[88] wl[185] vdd gnd cell_6t
Xbit_r186_c88 bl[88] br[88] wl[186] vdd gnd cell_6t
Xbit_r187_c88 bl[88] br[88] wl[187] vdd gnd cell_6t
Xbit_r188_c88 bl[88] br[88] wl[188] vdd gnd cell_6t
Xbit_r189_c88 bl[88] br[88] wl[189] vdd gnd cell_6t
Xbit_r190_c88 bl[88] br[88] wl[190] vdd gnd cell_6t
Xbit_r191_c88 bl[88] br[88] wl[191] vdd gnd cell_6t
Xbit_r192_c88 bl[88] br[88] wl[192] vdd gnd cell_6t
Xbit_r193_c88 bl[88] br[88] wl[193] vdd gnd cell_6t
Xbit_r194_c88 bl[88] br[88] wl[194] vdd gnd cell_6t
Xbit_r195_c88 bl[88] br[88] wl[195] vdd gnd cell_6t
Xbit_r196_c88 bl[88] br[88] wl[196] vdd gnd cell_6t
Xbit_r197_c88 bl[88] br[88] wl[197] vdd gnd cell_6t
Xbit_r198_c88 bl[88] br[88] wl[198] vdd gnd cell_6t
Xbit_r199_c88 bl[88] br[88] wl[199] vdd gnd cell_6t
Xbit_r200_c88 bl[88] br[88] wl[200] vdd gnd cell_6t
Xbit_r201_c88 bl[88] br[88] wl[201] vdd gnd cell_6t
Xbit_r202_c88 bl[88] br[88] wl[202] vdd gnd cell_6t
Xbit_r203_c88 bl[88] br[88] wl[203] vdd gnd cell_6t
Xbit_r204_c88 bl[88] br[88] wl[204] vdd gnd cell_6t
Xbit_r205_c88 bl[88] br[88] wl[205] vdd gnd cell_6t
Xbit_r206_c88 bl[88] br[88] wl[206] vdd gnd cell_6t
Xbit_r207_c88 bl[88] br[88] wl[207] vdd gnd cell_6t
Xbit_r208_c88 bl[88] br[88] wl[208] vdd gnd cell_6t
Xbit_r209_c88 bl[88] br[88] wl[209] vdd gnd cell_6t
Xbit_r210_c88 bl[88] br[88] wl[210] vdd gnd cell_6t
Xbit_r211_c88 bl[88] br[88] wl[211] vdd gnd cell_6t
Xbit_r212_c88 bl[88] br[88] wl[212] vdd gnd cell_6t
Xbit_r213_c88 bl[88] br[88] wl[213] vdd gnd cell_6t
Xbit_r214_c88 bl[88] br[88] wl[214] vdd gnd cell_6t
Xbit_r215_c88 bl[88] br[88] wl[215] vdd gnd cell_6t
Xbit_r216_c88 bl[88] br[88] wl[216] vdd gnd cell_6t
Xbit_r217_c88 bl[88] br[88] wl[217] vdd gnd cell_6t
Xbit_r218_c88 bl[88] br[88] wl[218] vdd gnd cell_6t
Xbit_r219_c88 bl[88] br[88] wl[219] vdd gnd cell_6t
Xbit_r220_c88 bl[88] br[88] wl[220] vdd gnd cell_6t
Xbit_r221_c88 bl[88] br[88] wl[221] vdd gnd cell_6t
Xbit_r222_c88 bl[88] br[88] wl[222] vdd gnd cell_6t
Xbit_r223_c88 bl[88] br[88] wl[223] vdd gnd cell_6t
Xbit_r224_c88 bl[88] br[88] wl[224] vdd gnd cell_6t
Xbit_r225_c88 bl[88] br[88] wl[225] vdd gnd cell_6t
Xbit_r226_c88 bl[88] br[88] wl[226] vdd gnd cell_6t
Xbit_r227_c88 bl[88] br[88] wl[227] vdd gnd cell_6t
Xbit_r228_c88 bl[88] br[88] wl[228] vdd gnd cell_6t
Xbit_r229_c88 bl[88] br[88] wl[229] vdd gnd cell_6t
Xbit_r230_c88 bl[88] br[88] wl[230] vdd gnd cell_6t
Xbit_r231_c88 bl[88] br[88] wl[231] vdd gnd cell_6t
Xbit_r232_c88 bl[88] br[88] wl[232] vdd gnd cell_6t
Xbit_r233_c88 bl[88] br[88] wl[233] vdd gnd cell_6t
Xbit_r234_c88 bl[88] br[88] wl[234] vdd gnd cell_6t
Xbit_r235_c88 bl[88] br[88] wl[235] vdd gnd cell_6t
Xbit_r236_c88 bl[88] br[88] wl[236] vdd gnd cell_6t
Xbit_r237_c88 bl[88] br[88] wl[237] vdd gnd cell_6t
Xbit_r238_c88 bl[88] br[88] wl[238] vdd gnd cell_6t
Xbit_r239_c88 bl[88] br[88] wl[239] vdd gnd cell_6t
Xbit_r240_c88 bl[88] br[88] wl[240] vdd gnd cell_6t
Xbit_r241_c88 bl[88] br[88] wl[241] vdd gnd cell_6t
Xbit_r242_c88 bl[88] br[88] wl[242] vdd gnd cell_6t
Xbit_r243_c88 bl[88] br[88] wl[243] vdd gnd cell_6t
Xbit_r244_c88 bl[88] br[88] wl[244] vdd gnd cell_6t
Xbit_r245_c88 bl[88] br[88] wl[245] vdd gnd cell_6t
Xbit_r246_c88 bl[88] br[88] wl[246] vdd gnd cell_6t
Xbit_r247_c88 bl[88] br[88] wl[247] vdd gnd cell_6t
Xbit_r248_c88 bl[88] br[88] wl[248] vdd gnd cell_6t
Xbit_r249_c88 bl[88] br[88] wl[249] vdd gnd cell_6t
Xbit_r250_c88 bl[88] br[88] wl[250] vdd gnd cell_6t
Xbit_r251_c88 bl[88] br[88] wl[251] vdd gnd cell_6t
Xbit_r252_c88 bl[88] br[88] wl[252] vdd gnd cell_6t
Xbit_r253_c88 bl[88] br[88] wl[253] vdd gnd cell_6t
Xbit_r254_c88 bl[88] br[88] wl[254] vdd gnd cell_6t
Xbit_r255_c88 bl[88] br[88] wl[255] vdd gnd cell_6t
Xbit_r256_c88 bl[88] br[88] wl[256] vdd gnd cell_6t
Xbit_r257_c88 bl[88] br[88] wl[257] vdd gnd cell_6t
Xbit_r258_c88 bl[88] br[88] wl[258] vdd gnd cell_6t
Xbit_r259_c88 bl[88] br[88] wl[259] vdd gnd cell_6t
Xbit_r260_c88 bl[88] br[88] wl[260] vdd gnd cell_6t
Xbit_r261_c88 bl[88] br[88] wl[261] vdd gnd cell_6t
Xbit_r262_c88 bl[88] br[88] wl[262] vdd gnd cell_6t
Xbit_r263_c88 bl[88] br[88] wl[263] vdd gnd cell_6t
Xbit_r264_c88 bl[88] br[88] wl[264] vdd gnd cell_6t
Xbit_r265_c88 bl[88] br[88] wl[265] vdd gnd cell_6t
Xbit_r266_c88 bl[88] br[88] wl[266] vdd gnd cell_6t
Xbit_r267_c88 bl[88] br[88] wl[267] vdd gnd cell_6t
Xbit_r268_c88 bl[88] br[88] wl[268] vdd gnd cell_6t
Xbit_r269_c88 bl[88] br[88] wl[269] vdd gnd cell_6t
Xbit_r270_c88 bl[88] br[88] wl[270] vdd gnd cell_6t
Xbit_r271_c88 bl[88] br[88] wl[271] vdd gnd cell_6t
Xbit_r272_c88 bl[88] br[88] wl[272] vdd gnd cell_6t
Xbit_r273_c88 bl[88] br[88] wl[273] vdd gnd cell_6t
Xbit_r274_c88 bl[88] br[88] wl[274] vdd gnd cell_6t
Xbit_r275_c88 bl[88] br[88] wl[275] vdd gnd cell_6t
Xbit_r276_c88 bl[88] br[88] wl[276] vdd gnd cell_6t
Xbit_r277_c88 bl[88] br[88] wl[277] vdd gnd cell_6t
Xbit_r278_c88 bl[88] br[88] wl[278] vdd gnd cell_6t
Xbit_r279_c88 bl[88] br[88] wl[279] vdd gnd cell_6t
Xbit_r280_c88 bl[88] br[88] wl[280] vdd gnd cell_6t
Xbit_r281_c88 bl[88] br[88] wl[281] vdd gnd cell_6t
Xbit_r282_c88 bl[88] br[88] wl[282] vdd gnd cell_6t
Xbit_r283_c88 bl[88] br[88] wl[283] vdd gnd cell_6t
Xbit_r284_c88 bl[88] br[88] wl[284] vdd gnd cell_6t
Xbit_r285_c88 bl[88] br[88] wl[285] vdd gnd cell_6t
Xbit_r286_c88 bl[88] br[88] wl[286] vdd gnd cell_6t
Xbit_r287_c88 bl[88] br[88] wl[287] vdd gnd cell_6t
Xbit_r288_c88 bl[88] br[88] wl[288] vdd gnd cell_6t
Xbit_r289_c88 bl[88] br[88] wl[289] vdd gnd cell_6t
Xbit_r290_c88 bl[88] br[88] wl[290] vdd gnd cell_6t
Xbit_r291_c88 bl[88] br[88] wl[291] vdd gnd cell_6t
Xbit_r292_c88 bl[88] br[88] wl[292] vdd gnd cell_6t
Xbit_r293_c88 bl[88] br[88] wl[293] vdd gnd cell_6t
Xbit_r294_c88 bl[88] br[88] wl[294] vdd gnd cell_6t
Xbit_r295_c88 bl[88] br[88] wl[295] vdd gnd cell_6t
Xbit_r296_c88 bl[88] br[88] wl[296] vdd gnd cell_6t
Xbit_r297_c88 bl[88] br[88] wl[297] vdd gnd cell_6t
Xbit_r298_c88 bl[88] br[88] wl[298] vdd gnd cell_6t
Xbit_r299_c88 bl[88] br[88] wl[299] vdd gnd cell_6t
Xbit_r300_c88 bl[88] br[88] wl[300] vdd gnd cell_6t
Xbit_r301_c88 bl[88] br[88] wl[301] vdd gnd cell_6t
Xbit_r302_c88 bl[88] br[88] wl[302] vdd gnd cell_6t
Xbit_r303_c88 bl[88] br[88] wl[303] vdd gnd cell_6t
Xbit_r304_c88 bl[88] br[88] wl[304] vdd gnd cell_6t
Xbit_r305_c88 bl[88] br[88] wl[305] vdd gnd cell_6t
Xbit_r306_c88 bl[88] br[88] wl[306] vdd gnd cell_6t
Xbit_r307_c88 bl[88] br[88] wl[307] vdd gnd cell_6t
Xbit_r308_c88 bl[88] br[88] wl[308] vdd gnd cell_6t
Xbit_r309_c88 bl[88] br[88] wl[309] vdd gnd cell_6t
Xbit_r310_c88 bl[88] br[88] wl[310] vdd gnd cell_6t
Xbit_r311_c88 bl[88] br[88] wl[311] vdd gnd cell_6t
Xbit_r312_c88 bl[88] br[88] wl[312] vdd gnd cell_6t
Xbit_r313_c88 bl[88] br[88] wl[313] vdd gnd cell_6t
Xbit_r314_c88 bl[88] br[88] wl[314] vdd gnd cell_6t
Xbit_r315_c88 bl[88] br[88] wl[315] vdd gnd cell_6t
Xbit_r316_c88 bl[88] br[88] wl[316] vdd gnd cell_6t
Xbit_r317_c88 bl[88] br[88] wl[317] vdd gnd cell_6t
Xbit_r318_c88 bl[88] br[88] wl[318] vdd gnd cell_6t
Xbit_r319_c88 bl[88] br[88] wl[319] vdd gnd cell_6t
Xbit_r320_c88 bl[88] br[88] wl[320] vdd gnd cell_6t
Xbit_r321_c88 bl[88] br[88] wl[321] vdd gnd cell_6t
Xbit_r322_c88 bl[88] br[88] wl[322] vdd gnd cell_6t
Xbit_r323_c88 bl[88] br[88] wl[323] vdd gnd cell_6t
Xbit_r324_c88 bl[88] br[88] wl[324] vdd gnd cell_6t
Xbit_r325_c88 bl[88] br[88] wl[325] vdd gnd cell_6t
Xbit_r326_c88 bl[88] br[88] wl[326] vdd gnd cell_6t
Xbit_r327_c88 bl[88] br[88] wl[327] vdd gnd cell_6t
Xbit_r328_c88 bl[88] br[88] wl[328] vdd gnd cell_6t
Xbit_r329_c88 bl[88] br[88] wl[329] vdd gnd cell_6t
Xbit_r330_c88 bl[88] br[88] wl[330] vdd gnd cell_6t
Xbit_r331_c88 bl[88] br[88] wl[331] vdd gnd cell_6t
Xbit_r332_c88 bl[88] br[88] wl[332] vdd gnd cell_6t
Xbit_r333_c88 bl[88] br[88] wl[333] vdd gnd cell_6t
Xbit_r334_c88 bl[88] br[88] wl[334] vdd gnd cell_6t
Xbit_r335_c88 bl[88] br[88] wl[335] vdd gnd cell_6t
Xbit_r336_c88 bl[88] br[88] wl[336] vdd gnd cell_6t
Xbit_r337_c88 bl[88] br[88] wl[337] vdd gnd cell_6t
Xbit_r338_c88 bl[88] br[88] wl[338] vdd gnd cell_6t
Xbit_r339_c88 bl[88] br[88] wl[339] vdd gnd cell_6t
Xbit_r340_c88 bl[88] br[88] wl[340] vdd gnd cell_6t
Xbit_r341_c88 bl[88] br[88] wl[341] vdd gnd cell_6t
Xbit_r342_c88 bl[88] br[88] wl[342] vdd gnd cell_6t
Xbit_r343_c88 bl[88] br[88] wl[343] vdd gnd cell_6t
Xbit_r344_c88 bl[88] br[88] wl[344] vdd gnd cell_6t
Xbit_r345_c88 bl[88] br[88] wl[345] vdd gnd cell_6t
Xbit_r346_c88 bl[88] br[88] wl[346] vdd gnd cell_6t
Xbit_r347_c88 bl[88] br[88] wl[347] vdd gnd cell_6t
Xbit_r348_c88 bl[88] br[88] wl[348] vdd gnd cell_6t
Xbit_r349_c88 bl[88] br[88] wl[349] vdd gnd cell_6t
Xbit_r350_c88 bl[88] br[88] wl[350] vdd gnd cell_6t
Xbit_r351_c88 bl[88] br[88] wl[351] vdd gnd cell_6t
Xbit_r352_c88 bl[88] br[88] wl[352] vdd gnd cell_6t
Xbit_r353_c88 bl[88] br[88] wl[353] vdd gnd cell_6t
Xbit_r354_c88 bl[88] br[88] wl[354] vdd gnd cell_6t
Xbit_r355_c88 bl[88] br[88] wl[355] vdd gnd cell_6t
Xbit_r356_c88 bl[88] br[88] wl[356] vdd gnd cell_6t
Xbit_r357_c88 bl[88] br[88] wl[357] vdd gnd cell_6t
Xbit_r358_c88 bl[88] br[88] wl[358] vdd gnd cell_6t
Xbit_r359_c88 bl[88] br[88] wl[359] vdd gnd cell_6t
Xbit_r360_c88 bl[88] br[88] wl[360] vdd gnd cell_6t
Xbit_r361_c88 bl[88] br[88] wl[361] vdd gnd cell_6t
Xbit_r362_c88 bl[88] br[88] wl[362] vdd gnd cell_6t
Xbit_r363_c88 bl[88] br[88] wl[363] vdd gnd cell_6t
Xbit_r364_c88 bl[88] br[88] wl[364] vdd gnd cell_6t
Xbit_r365_c88 bl[88] br[88] wl[365] vdd gnd cell_6t
Xbit_r366_c88 bl[88] br[88] wl[366] vdd gnd cell_6t
Xbit_r367_c88 bl[88] br[88] wl[367] vdd gnd cell_6t
Xbit_r368_c88 bl[88] br[88] wl[368] vdd gnd cell_6t
Xbit_r369_c88 bl[88] br[88] wl[369] vdd gnd cell_6t
Xbit_r370_c88 bl[88] br[88] wl[370] vdd gnd cell_6t
Xbit_r371_c88 bl[88] br[88] wl[371] vdd gnd cell_6t
Xbit_r372_c88 bl[88] br[88] wl[372] vdd gnd cell_6t
Xbit_r373_c88 bl[88] br[88] wl[373] vdd gnd cell_6t
Xbit_r374_c88 bl[88] br[88] wl[374] vdd gnd cell_6t
Xbit_r375_c88 bl[88] br[88] wl[375] vdd gnd cell_6t
Xbit_r376_c88 bl[88] br[88] wl[376] vdd gnd cell_6t
Xbit_r377_c88 bl[88] br[88] wl[377] vdd gnd cell_6t
Xbit_r378_c88 bl[88] br[88] wl[378] vdd gnd cell_6t
Xbit_r379_c88 bl[88] br[88] wl[379] vdd gnd cell_6t
Xbit_r380_c88 bl[88] br[88] wl[380] vdd gnd cell_6t
Xbit_r381_c88 bl[88] br[88] wl[381] vdd gnd cell_6t
Xbit_r382_c88 bl[88] br[88] wl[382] vdd gnd cell_6t
Xbit_r383_c88 bl[88] br[88] wl[383] vdd gnd cell_6t
Xbit_r384_c88 bl[88] br[88] wl[384] vdd gnd cell_6t
Xbit_r385_c88 bl[88] br[88] wl[385] vdd gnd cell_6t
Xbit_r386_c88 bl[88] br[88] wl[386] vdd gnd cell_6t
Xbit_r387_c88 bl[88] br[88] wl[387] vdd gnd cell_6t
Xbit_r388_c88 bl[88] br[88] wl[388] vdd gnd cell_6t
Xbit_r389_c88 bl[88] br[88] wl[389] vdd gnd cell_6t
Xbit_r390_c88 bl[88] br[88] wl[390] vdd gnd cell_6t
Xbit_r391_c88 bl[88] br[88] wl[391] vdd gnd cell_6t
Xbit_r392_c88 bl[88] br[88] wl[392] vdd gnd cell_6t
Xbit_r393_c88 bl[88] br[88] wl[393] vdd gnd cell_6t
Xbit_r394_c88 bl[88] br[88] wl[394] vdd gnd cell_6t
Xbit_r395_c88 bl[88] br[88] wl[395] vdd gnd cell_6t
Xbit_r396_c88 bl[88] br[88] wl[396] vdd gnd cell_6t
Xbit_r397_c88 bl[88] br[88] wl[397] vdd gnd cell_6t
Xbit_r398_c88 bl[88] br[88] wl[398] vdd gnd cell_6t
Xbit_r399_c88 bl[88] br[88] wl[399] vdd gnd cell_6t
Xbit_r400_c88 bl[88] br[88] wl[400] vdd gnd cell_6t
Xbit_r401_c88 bl[88] br[88] wl[401] vdd gnd cell_6t
Xbit_r402_c88 bl[88] br[88] wl[402] vdd gnd cell_6t
Xbit_r403_c88 bl[88] br[88] wl[403] vdd gnd cell_6t
Xbit_r404_c88 bl[88] br[88] wl[404] vdd gnd cell_6t
Xbit_r405_c88 bl[88] br[88] wl[405] vdd gnd cell_6t
Xbit_r406_c88 bl[88] br[88] wl[406] vdd gnd cell_6t
Xbit_r407_c88 bl[88] br[88] wl[407] vdd gnd cell_6t
Xbit_r408_c88 bl[88] br[88] wl[408] vdd gnd cell_6t
Xbit_r409_c88 bl[88] br[88] wl[409] vdd gnd cell_6t
Xbit_r410_c88 bl[88] br[88] wl[410] vdd gnd cell_6t
Xbit_r411_c88 bl[88] br[88] wl[411] vdd gnd cell_6t
Xbit_r412_c88 bl[88] br[88] wl[412] vdd gnd cell_6t
Xbit_r413_c88 bl[88] br[88] wl[413] vdd gnd cell_6t
Xbit_r414_c88 bl[88] br[88] wl[414] vdd gnd cell_6t
Xbit_r415_c88 bl[88] br[88] wl[415] vdd gnd cell_6t
Xbit_r416_c88 bl[88] br[88] wl[416] vdd gnd cell_6t
Xbit_r417_c88 bl[88] br[88] wl[417] vdd gnd cell_6t
Xbit_r418_c88 bl[88] br[88] wl[418] vdd gnd cell_6t
Xbit_r419_c88 bl[88] br[88] wl[419] vdd gnd cell_6t
Xbit_r420_c88 bl[88] br[88] wl[420] vdd gnd cell_6t
Xbit_r421_c88 bl[88] br[88] wl[421] vdd gnd cell_6t
Xbit_r422_c88 bl[88] br[88] wl[422] vdd gnd cell_6t
Xbit_r423_c88 bl[88] br[88] wl[423] vdd gnd cell_6t
Xbit_r424_c88 bl[88] br[88] wl[424] vdd gnd cell_6t
Xbit_r425_c88 bl[88] br[88] wl[425] vdd gnd cell_6t
Xbit_r426_c88 bl[88] br[88] wl[426] vdd gnd cell_6t
Xbit_r427_c88 bl[88] br[88] wl[427] vdd gnd cell_6t
Xbit_r428_c88 bl[88] br[88] wl[428] vdd gnd cell_6t
Xbit_r429_c88 bl[88] br[88] wl[429] vdd gnd cell_6t
Xbit_r430_c88 bl[88] br[88] wl[430] vdd gnd cell_6t
Xbit_r431_c88 bl[88] br[88] wl[431] vdd gnd cell_6t
Xbit_r432_c88 bl[88] br[88] wl[432] vdd gnd cell_6t
Xbit_r433_c88 bl[88] br[88] wl[433] vdd gnd cell_6t
Xbit_r434_c88 bl[88] br[88] wl[434] vdd gnd cell_6t
Xbit_r435_c88 bl[88] br[88] wl[435] vdd gnd cell_6t
Xbit_r436_c88 bl[88] br[88] wl[436] vdd gnd cell_6t
Xbit_r437_c88 bl[88] br[88] wl[437] vdd gnd cell_6t
Xbit_r438_c88 bl[88] br[88] wl[438] vdd gnd cell_6t
Xbit_r439_c88 bl[88] br[88] wl[439] vdd gnd cell_6t
Xbit_r440_c88 bl[88] br[88] wl[440] vdd gnd cell_6t
Xbit_r441_c88 bl[88] br[88] wl[441] vdd gnd cell_6t
Xbit_r442_c88 bl[88] br[88] wl[442] vdd gnd cell_6t
Xbit_r443_c88 bl[88] br[88] wl[443] vdd gnd cell_6t
Xbit_r444_c88 bl[88] br[88] wl[444] vdd gnd cell_6t
Xbit_r445_c88 bl[88] br[88] wl[445] vdd gnd cell_6t
Xbit_r446_c88 bl[88] br[88] wl[446] vdd gnd cell_6t
Xbit_r447_c88 bl[88] br[88] wl[447] vdd gnd cell_6t
Xbit_r448_c88 bl[88] br[88] wl[448] vdd gnd cell_6t
Xbit_r449_c88 bl[88] br[88] wl[449] vdd gnd cell_6t
Xbit_r450_c88 bl[88] br[88] wl[450] vdd gnd cell_6t
Xbit_r451_c88 bl[88] br[88] wl[451] vdd gnd cell_6t
Xbit_r452_c88 bl[88] br[88] wl[452] vdd gnd cell_6t
Xbit_r453_c88 bl[88] br[88] wl[453] vdd gnd cell_6t
Xbit_r454_c88 bl[88] br[88] wl[454] vdd gnd cell_6t
Xbit_r455_c88 bl[88] br[88] wl[455] vdd gnd cell_6t
Xbit_r456_c88 bl[88] br[88] wl[456] vdd gnd cell_6t
Xbit_r457_c88 bl[88] br[88] wl[457] vdd gnd cell_6t
Xbit_r458_c88 bl[88] br[88] wl[458] vdd gnd cell_6t
Xbit_r459_c88 bl[88] br[88] wl[459] vdd gnd cell_6t
Xbit_r460_c88 bl[88] br[88] wl[460] vdd gnd cell_6t
Xbit_r461_c88 bl[88] br[88] wl[461] vdd gnd cell_6t
Xbit_r462_c88 bl[88] br[88] wl[462] vdd gnd cell_6t
Xbit_r463_c88 bl[88] br[88] wl[463] vdd gnd cell_6t
Xbit_r464_c88 bl[88] br[88] wl[464] vdd gnd cell_6t
Xbit_r465_c88 bl[88] br[88] wl[465] vdd gnd cell_6t
Xbit_r466_c88 bl[88] br[88] wl[466] vdd gnd cell_6t
Xbit_r467_c88 bl[88] br[88] wl[467] vdd gnd cell_6t
Xbit_r468_c88 bl[88] br[88] wl[468] vdd gnd cell_6t
Xbit_r469_c88 bl[88] br[88] wl[469] vdd gnd cell_6t
Xbit_r470_c88 bl[88] br[88] wl[470] vdd gnd cell_6t
Xbit_r471_c88 bl[88] br[88] wl[471] vdd gnd cell_6t
Xbit_r472_c88 bl[88] br[88] wl[472] vdd gnd cell_6t
Xbit_r473_c88 bl[88] br[88] wl[473] vdd gnd cell_6t
Xbit_r474_c88 bl[88] br[88] wl[474] vdd gnd cell_6t
Xbit_r475_c88 bl[88] br[88] wl[475] vdd gnd cell_6t
Xbit_r476_c88 bl[88] br[88] wl[476] vdd gnd cell_6t
Xbit_r477_c88 bl[88] br[88] wl[477] vdd gnd cell_6t
Xbit_r478_c88 bl[88] br[88] wl[478] vdd gnd cell_6t
Xbit_r479_c88 bl[88] br[88] wl[479] vdd gnd cell_6t
Xbit_r480_c88 bl[88] br[88] wl[480] vdd gnd cell_6t
Xbit_r481_c88 bl[88] br[88] wl[481] vdd gnd cell_6t
Xbit_r482_c88 bl[88] br[88] wl[482] vdd gnd cell_6t
Xbit_r483_c88 bl[88] br[88] wl[483] vdd gnd cell_6t
Xbit_r484_c88 bl[88] br[88] wl[484] vdd gnd cell_6t
Xbit_r485_c88 bl[88] br[88] wl[485] vdd gnd cell_6t
Xbit_r486_c88 bl[88] br[88] wl[486] vdd gnd cell_6t
Xbit_r487_c88 bl[88] br[88] wl[487] vdd gnd cell_6t
Xbit_r488_c88 bl[88] br[88] wl[488] vdd gnd cell_6t
Xbit_r489_c88 bl[88] br[88] wl[489] vdd gnd cell_6t
Xbit_r490_c88 bl[88] br[88] wl[490] vdd gnd cell_6t
Xbit_r491_c88 bl[88] br[88] wl[491] vdd gnd cell_6t
Xbit_r492_c88 bl[88] br[88] wl[492] vdd gnd cell_6t
Xbit_r493_c88 bl[88] br[88] wl[493] vdd gnd cell_6t
Xbit_r494_c88 bl[88] br[88] wl[494] vdd gnd cell_6t
Xbit_r495_c88 bl[88] br[88] wl[495] vdd gnd cell_6t
Xbit_r496_c88 bl[88] br[88] wl[496] vdd gnd cell_6t
Xbit_r497_c88 bl[88] br[88] wl[497] vdd gnd cell_6t
Xbit_r498_c88 bl[88] br[88] wl[498] vdd gnd cell_6t
Xbit_r499_c88 bl[88] br[88] wl[499] vdd gnd cell_6t
Xbit_r500_c88 bl[88] br[88] wl[500] vdd gnd cell_6t
Xbit_r501_c88 bl[88] br[88] wl[501] vdd gnd cell_6t
Xbit_r502_c88 bl[88] br[88] wl[502] vdd gnd cell_6t
Xbit_r503_c88 bl[88] br[88] wl[503] vdd gnd cell_6t
Xbit_r504_c88 bl[88] br[88] wl[504] vdd gnd cell_6t
Xbit_r505_c88 bl[88] br[88] wl[505] vdd gnd cell_6t
Xbit_r506_c88 bl[88] br[88] wl[506] vdd gnd cell_6t
Xbit_r507_c88 bl[88] br[88] wl[507] vdd gnd cell_6t
Xbit_r508_c88 bl[88] br[88] wl[508] vdd gnd cell_6t
Xbit_r509_c88 bl[88] br[88] wl[509] vdd gnd cell_6t
Xbit_r510_c88 bl[88] br[88] wl[510] vdd gnd cell_6t
Xbit_r511_c88 bl[88] br[88] wl[511] vdd gnd cell_6t
Xbit_r0_c89 bl[89] br[89] wl[0] vdd gnd cell_6t
Xbit_r1_c89 bl[89] br[89] wl[1] vdd gnd cell_6t
Xbit_r2_c89 bl[89] br[89] wl[2] vdd gnd cell_6t
Xbit_r3_c89 bl[89] br[89] wl[3] vdd gnd cell_6t
Xbit_r4_c89 bl[89] br[89] wl[4] vdd gnd cell_6t
Xbit_r5_c89 bl[89] br[89] wl[5] vdd gnd cell_6t
Xbit_r6_c89 bl[89] br[89] wl[6] vdd gnd cell_6t
Xbit_r7_c89 bl[89] br[89] wl[7] vdd gnd cell_6t
Xbit_r8_c89 bl[89] br[89] wl[8] vdd gnd cell_6t
Xbit_r9_c89 bl[89] br[89] wl[9] vdd gnd cell_6t
Xbit_r10_c89 bl[89] br[89] wl[10] vdd gnd cell_6t
Xbit_r11_c89 bl[89] br[89] wl[11] vdd gnd cell_6t
Xbit_r12_c89 bl[89] br[89] wl[12] vdd gnd cell_6t
Xbit_r13_c89 bl[89] br[89] wl[13] vdd gnd cell_6t
Xbit_r14_c89 bl[89] br[89] wl[14] vdd gnd cell_6t
Xbit_r15_c89 bl[89] br[89] wl[15] vdd gnd cell_6t
Xbit_r16_c89 bl[89] br[89] wl[16] vdd gnd cell_6t
Xbit_r17_c89 bl[89] br[89] wl[17] vdd gnd cell_6t
Xbit_r18_c89 bl[89] br[89] wl[18] vdd gnd cell_6t
Xbit_r19_c89 bl[89] br[89] wl[19] vdd gnd cell_6t
Xbit_r20_c89 bl[89] br[89] wl[20] vdd gnd cell_6t
Xbit_r21_c89 bl[89] br[89] wl[21] vdd gnd cell_6t
Xbit_r22_c89 bl[89] br[89] wl[22] vdd gnd cell_6t
Xbit_r23_c89 bl[89] br[89] wl[23] vdd gnd cell_6t
Xbit_r24_c89 bl[89] br[89] wl[24] vdd gnd cell_6t
Xbit_r25_c89 bl[89] br[89] wl[25] vdd gnd cell_6t
Xbit_r26_c89 bl[89] br[89] wl[26] vdd gnd cell_6t
Xbit_r27_c89 bl[89] br[89] wl[27] vdd gnd cell_6t
Xbit_r28_c89 bl[89] br[89] wl[28] vdd gnd cell_6t
Xbit_r29_c89 bl[89] br[89] wl[29] vdd gnd cell_6t
Xbit_r30_c89 bl[89] br[89] wl[30] vdd gnd cell_6t
Xbit_r31_c89 bl[89] br[89] wl[31] vdd gnd cell_6t
Xbit_r32_c89 bl[89] br[89] wl[32] vdd gnd cell_6t
Xbit_r33_c89 bl[89] br[89] wl[33] vdd gnd cell_6t
Xbit_r34_c89 bl[89] br[89] wl[34] vdd gnd cell_6t
Xbit_r35_c89 bl[89] br[89] wl[35] vdd gnd cell_6t
Xbit_r36_c89 bl[89] br[89] wl[36] vdd gnd cell_6t
Xbit_r37_c89 bl[89] br[89] wl[37] vdd gnd cell_6t
Xbit_r38_c89 bl[89] br[89] wl[38] vdd gnd cell_6t
Xbit_r39_c89 bl[89] br[89] wl[39] vdd gnd cell_6t
Xbit_r40_c89 bl[89] br[89] wl[40] vdd gnd cell_6t
Xbit_r41_c89 bl[89] br[89] wl[41] vdd gnd cell_6t
Xbit_r42_c89 bl[89] br[89] wl[42] vdd gnd cell_6t
Xbit_r43_c89 bl[89] br[89] wl[43] vdd gnd cell_6t
Xbit_r44_c89 bl[89] br[89] wl[44] vdd gnd cell_6t
Xbit_r45_c89 bl[89] br[89] wl[45] vdd gnd cell_6t
Xbit_r46_c89 bl[89] br[89] wl[46] vdd gnd cell_6t
Xbit_r47_c89 bl[89] br[89] wl[47] vdd gnd cell_6t
Xbit_r48_c89 bl[89] br[89] wl[48] vdd gnd cell_6t
Xbit_r49_c89 bl[89] br[89] wl[49] vdd gnd cell_6t
Xbit_r50_c89 bl[89] br[89] wl[50] vdd gnd cell_6t
Xbit_r51_c89 bl[89] br[89] wl[51] vdd gnd cell_6t
Xbit_r52_c89 bl[89] br[89] wl[52] vdd gnd cell_6t
Xbit_r53_c89 bl[89] br[89] wl[53] vdd gnd cell_6t
Xbit_r54_c89 bl[89] br[89] wl[54] vdd gnd cell_6t
Xbit_r55_c89 bl[89] br[89] wl[55] vdd gnd cell_6t
Xbit_r56_c89 bl[89] br[89] wl[56] vdd gnd cell_6t
Xbit_r57_c89 bl[89] br[89] wl[57] vdd gnd cell_6t
Xbit_r58_c89 bl[89] br[89] wl[58] vdd gnd cell_6t
Xbit_r59_c89 bl[89] br[89] wl[59] vdd gnd cell_6t
Xbit_r60_c89 bl[89] br[89] wl[60] vdd gnd cell_6t
Xbit_r61_c89 bl[89] br[89] wl[61] vdd gnd cell_6t
Xbit_r62_c89 bl[89] br[89] wl[62] vdd gnd cell_6t
Xbit_r63_c89 bl[89] br[89] wl[63] vdd gnd cell_6t
Xbit_r64_c89 bl[89] br[89] wl[64] vdd gnd cell_6t
Xbit_r65_c89 bl[89] br[89] wl[65] vdd gnd cell_6t
Xbit_r66_c89 bl[89] br[89] wl[66] vdd gnd cell_6t
Xbit_r67_c89 bl[89] br[89] wl[67] vdd gnd cell_6t
Xbit_r68_c89 bl[89] br[89] wl[68] vdd gnd cell_6t
Xbit_r69_c89 bl[89] br[89] wl[69] vdd gnd cell_6t
Xbit_r70_c89 bl[89] br[89] wl[70] vdd gnd cell_6t
Xbit_r71_c89 bl[89] br[89] wl[71] vdd gnd cell_6t
Xbit_r72_c89 bl[89] br[89] wl[72] vdd gnd cell_6t
Xbit_r73_c89 bl[89] br[89] wl[73] vdd gnd cell_6t
Xbit_r74_c89 bl[89] br[89] wl[74] vdd gnd cell_6t
Xbit_r75_c89 bl[89] br[89] wl[75] vdd gnd cell_6t
Xbit_r76_c89 bl[89] br[89] wl[76] vdd gnd cell_6t
Xbit_r77_c89 bl[89] br[89] wl[77] vdd gnd cell_6t
Xbit_r78_c89 bl[89] br[89] wl[78] vdd gnd cell_6t
Xbit_r79_c89 bl[89] br[89] wl[79] vdd gnd cell_6t
Xbit_r80_c89 bl[89] br[89] wl[80] vdd gnd cell_6t
Xbit_r81_c89 bl[89] br[89] wl[81] vdd gnd cell_6t
Xbit_r82_c89 bl[89] br[89] wl[82] vdd gnd cell_6t
Xbit_r83_c89 bl[89] br[89] wl[83] vdd gnd cell_6t
Xbit_r84_c89 bl[89] br[89] wl[84] vdd gnd cell_6t
Xbit_r85_c89 bl[89] br[89] wl[85] vdd gnd cell_6t
Xbit_r86_c89 bl[89] br[89] wl[86] vdd gnd cell_6t
Xbit_r87_c89 bl[89] br[89] wl[87] vdd gnd cell_6t
Xbit_r88_c89 bl[89] br[89] wl[88] vdd gnd cell_6t
Xbit_r89_c89 bl[89] br[89] wl[89] vdd gnd cell_6t
Xbit_r90_c89 bl[89] br[89] wl[90] vdd gnd cell_6t
Xbit_r91_c89 bl[89] br[89] wl[91] vdd gnd cell_6t
Xbit_r92_c89 bl[89] br[89] wl[92] vdd gnd cell_6t
Xbit_r93_c89 bl[89] br[89] wl[93] vdd gnd cell_6t
Xbit_r94_c89 bl[89] br[89] wl[94] vdd gnd cell_6t
Xbit_r95_c89 bl[89] br[89] wl[95] vdd gnd cell_6t
Xbit_r96_c89 bl[89] br[89] wl[96] vdd gnd cell_6t
Xbit_r97_c89 bl[89] br[89] wl[97] vdd gnd cell_6t
Xbit_r98_c89 bl[89] br[89] wl[98] vdd gnd cell_6t
Xbit_r99_c89 bl[89] br[89] wl[99] vdd gnd cell_6t
Xbit_r100_c89 bl[89] br[89] wl[100] vdd gnd cell_6t
Xbit_r101_c89 bl[89] br[89] wl[101] vdd gnd cell_6t
Xbit_r102_c89 bl[89] br[89] wl[102] vdd gnd cell_6t
Xbit_r103_c89 bl[89] br[89] wl[103] vdd gnd cell_6t
Xbit_r104_c89 bl[89] br[89] wl[104] vdd gnd cell_6t
Xbit_r105_c89 bl[89] br[89] wl[105] vdd gnd cell_6t
Xbit_r106_c89 bl[89] br[89] wl[106] vdd gnd cell_6t
Xbit_r107_c89 bl[89] br[89] wl[107] vdd gnd cell_6t
Xbit_r108_c89 bl[89] br[89] wl[108] vdd gnd cell_6t
Xbit_r109_c89 bl[89] br[89] wl[109] vdd gnd cell_6t
Xbit_r110_c89 bl[89] br[89] wl[110] vdd gnd cell_6t
Xbit_r111_c89 bl[89] br[89] wl[111] vdd gnd cell_6t
Xbit_r112_c89 bl[89] br[89] wl[112] vdd gnd cell_6t
Xbit_r113_c89 bl[89] br[89] wl[113] vdd gnd cell_6t
Xbit_r114_c89 bl[89] br[89] wl[114] vdd gnd cell_6t
Xbit_r115_c89 bl[89] br[89] wl[115] vdd gnd cell_6t
Xbit_r116_c89 bl[89] br[89] wl[116] vdd gnd cell_6t
Xbit_r117_c89 bl[89] br[89] wl[117] vdd gnd cell_6t
Xbit_r118_c89 bl[89] br[89] wl[118] vdd gnd cell_6t
Xbit_r119_c89 bl[89] br[89] wl[119] vdd gnd cell_6t
Xbit_r120_c89 bl[89] br[89] wl[120] vdd gnd cell_6t
Xbit_r121_c89 bl[89] br[89] wl[121] vdd gnd cell_6t
Xbit_r122_c89 bl[89] br[89] wl[122] vdd gnd cell_6t
Xbit_r123_c89 bl[89] br[89] wl[123] vdd gnd cell_6t
Xbit_r124_c89 bl[89] br[89] wl[124] vdd gnd cell_6t
Xbit_r125_c89 bl[89] br[89] wl[125] vdd gnd cell_6t
Xbit_r126_c89 bl[89] br[89] wl[126] vdd gnd cell_6t
Xbit_r127_c89 bl[89] br[89] wl[127] vdd gnd cell_6t
Xbit_r128_c89 bl[89] br[89] wl[128] vdd gnd cell_6t
Xbit_r129_c89 bl[89] br[89] wl[129] vdd gnd cell_6t
Xbit_r130_c89 bl[89] br[89] wl[130] vdd gnd cell_6t
Xbit_r131_c89 bl[89] br[89] wl[131] vdd gnd cell_6t
Xbit_r132_c89 bl[89] br[89] wl[132] vdd gnd cell_6t
Xbit_r133_c89 bl[89] br[89] wl[133] vdd gnd cell_6t
Xbit_r134_c89 bl[89] br[89] wl[134] vdd gnd cell_6t
Xbit_r135_c89 bl[89] br[89] wl[135] vdd gnd cell_6t
Xbit_r136_c89 bl[89] br[89] wl[136] vdd gnd cell_6t
Xbit_r137_c89 bl[89] br[89] wl[137] vdd gnd cell_6t
Xbit_r138_c89 bl[89] br[89] wl[138] vdd gnd cell_6t
Xbit_r139_c89 bl[89] br[89] wl[139] vdd gnd cell_6t
Xbit_r140_c89 bl[89] br[89] wl[140] vdd gnd cell_6t
Xbit_r141_c89 bl[89] br[89] wl[141] vdd gnd cell_6t
Xbit_r142_c89 bl[89] br[89] wl[142] vdd gnd cell_6t
Xbit_r143_c89 bl[89] br[89] wl[143] vdd gnd cell_6t
Xbit_r144_c89 bl[89] br[89] wl[144] vdd gnd cell_6t
Xbit_r145_c89 bl[89] br[89] wl[145] vdd gnd cell_6t
Xbit_r146_c89 bl[89] br[89] wl[146] vdd gnd cell_6t
Xbit_r147_c89 bl[89] br[89] wl[147] vdd gnd cell_6t
Xbit_r148_c89 bl[89] br[89] wl[148] vdd gnd cell_6t
Xbit_r149_c89 bl[89] br[89] wl[149] vdd gnd cell_6t
Xbit_r150_c89 bl[89] br[89] wl[150] vdd gnd cell_6t
Xbit_r151_c89 bl[89] br[89] wl[151] vdd gnd cell_6t
Xbit_r152_c89 bl[89] br[89] wl[152] vdd gnd cell_6t
Xbit_r153_c89 bl[89] br[89] wl[153] vdd gnd cell_6t
Xbit_r154_c89 bl[89] br[89] wl[154] vdd gnd cell_6t
Xbit_r155_c89 bl[89] br[89] wl[155] vdd gnd cell_6t
Xbit_r156_c89 bl[89] br[89] wl[156] vdd gnd cell_6t
Xbit_r157_c89 bl[89] br[89] wl[157] vdd gnd cell_6t
Xbit_r158_c89 bl[89] br[89] wl[158] vdd gnd cell_6t
Xbit_r159_c89 bl[89] br[89] wl[159] vdd gnd cell_6t
Xbit_r160_c89 bl[89] br[89] wl[160] vdd gnd cell_6t
Xbit_r161_c89 bl[89] br[89] wl[161] vdd gnd cell_6t
Xbit_r162_c89 bl[89] br[89] wl[162] vdd gnd cell_6t
Xbit_r163_c89 bl[89] br[89] wl[163] vdd gnd cell_6t
Xbit_r164_c89 bl[89] br[89] wl[164] vdd gnd cell_6t
Xbit_r165_c89 bl[89] br[89] wl[165] vdd gnd cell_6t
Xbit_r166_c89 bl[89] br[89] wl[166] vdd gnd cell_6t
Xbit_r167_c89 bl[89] br[89] wl[167] vdd gnd cell_6t
Xbit_r168_c89 bl[89] br[89] wl[168] vdd gnd cell_6t
Xbit_r169_c89 bl[89] br[89] wl[169] vdd gnd cell_6t
Xbit_r170_c89 bl[89] br[89] wl[170] vdd gnd cell_6t
Xbit_r171_c89 bl[89] br[89] wl[171] vdd gnd cell_6t
Xbit_r172_c89 bl[89] br[89] wl[172] vdd gnd cell_6t
Xbit_r173_c89 bl[89] br[89] wl[173] vdd gnd cell_6t
Xbit_r174_c89 bl[89] br[89] wl[174] vdd gnd cell_6t
Xbit_r175_c89 bl[89] br[89] wl[175] vdd gnd cell_6t
Xbit_r176_c89 bl[89] br[89] wl[176] vdd gnd cell_6t
Xbit_r177_c89 bl[89] br[89] wl[177] vdd gnd cell_6t
Xbit_r178_c89 bl[89] br[89] wl[178] vdd gnd cell_6t
Xbit_r179_c89 bl[89] br[89] wl[179] vdd gnd cell_6t
Xbit_r180_c89 bl[89] br[89] wl[180] vdd gnd cell_6t
Xbit_r181_c89 bl[89] br[89] wl[181] vdd gnd cell_6t
Xbit_r182_c89 bl[89] br[89] wl[182] vdd gnd cell_6t
Xbit_r183_c89 bl[89] br[89] wl[183] vdd gnd cell_6t
Xbit_r184_c89 bl[89] br[89] wl[184] vdd gnd cell_6t
Xbit_r185_c89 bl[89] br[89] wl[185] vdd gnd cell_6t
Xbit_r186_c89 bl[89] br[89] wl[186] vdd gnd cell_6t
Xbit_r187_c89 bl[89] br[89] wl[187] vdd gnd cell_6t
Xbit_r188_c89 bl[89] br[89] wl[188] vdd gnd cell_6t
Xbit_r189_c89 bl[89] br[89] wl[189] vdd gnd cell_6t
Xbit_r190_c89 bl[89] br[89] wl[190] vdd gnd cell_6t
Xbit_r191_c89 bl[89] br[89] wl[191] vdd gnd cell_6t
Xbit_r192_c89 bl[89] br[89] wl[192] vdd gnd cell_6t
Xbit_r193_c89 bl[89] br[89] wl[193] vdd gnd cell_6t
Xbit_r194_c89 bl[89] br[89] wl[194] vdd gnd cell_6t
Xbit_r195_c89 bl[89] br[89] wl[195] vdd gnd cell_6t
Xbit_r196_c89 bl[89] br[89] wl[196] vdd gnd cell_6t
Xbit_r197_c89 bl[89] br[89] wl[197] vdd gnd cell_6t
Xbit_r198_c89 bl[89] br[89] wl[198] vdd gnd cell_6t
Xbit_r199_c89 bl[89] br[89] wl[199] vdd gnd cell_6t
Xbit_r200_c89 bl[89] br[89] wl[200] vdd gnd cell_6t
Xbit_r201_c89 bl[89] br[89] wl[201] vdd gnd cell_6t
Xbit_r202_c89 bl[89] br[89] wl[202] vdd gnd cell_6t
Xbit_r203_c89 bl[89] br[89] wl[203] vdd gnd cell_6t
Xbit_r204_c89 bl[89] br[89] wl[204] vdd gnd cell_6t
Xbit_r205_c89 bl[89] br[89] wl[205] vdd gnd cell_6t
Xbit_r206_c89 bl[89] br[89] wl[206] vdd gnd cell_6t
Xbit_r207_c89 bl[89] br[89] wl[207] vdd gnd cell_6t
Xbit_r208_c89 bl[89] br[89] wl[208] vdd gnd cell_6t
Xbit_r209_c89 bl[89] br[89] wl[209] vdd gnd cell_6t
Xbit_r210_c89 bl[89] br[89] wl[210] vdd gnd cell_6t
Xbit_r211_c89 bl[89] br[89] wl[211] vdd gnd cell_6t
Xbit_r212_c89 bl[89] br[89] wl[212] vdd gnd cell_6t
Xbit_r213_c89 bl[89] br[89] wl[213] vdd gnd cell_6t
Xbit_r214_c89 bl[89] br[89] wl[214] vdd gnd cell_6t
Xbit_r215_c89 bl[89] br[89] wl[215] vdd gnd cell_6t
Xbit_r216_c89 bl[89] br[89] wl[216] vdd gnd cell_6t
Xbit_r217_c89 bl[89] br[89] wl[217] vdd gnd cell_6t
Xbit_r218_c89 bl[89] br[89] wl[218] vdd gnd cell_6t
Xbit_r219_c89 bl[89] br[89] wl[219] vdd gnd cell_6t
Xbit_r220_c89 bl[89] br[89] wl[220] vdd gnd cell_6t
Xbit_r221_c89 bl[89] br[89] wl[221] vdd gnd cell_6t
Xbit_r222_c89 bl[89] br[89] wl[222] vdd gnd cell_6t
Xbit_r223_c89 bl[89] br[89] wl[223] vdd gnd cell_6t
Xbit_r224_c89 bl[89] br[89] wl[224] vdd gnd cell_6t
Xbit_r225_c89 bl[89] br[89] wl[225] vdd gnd cell_6t
Xbit_r226_c89 bl[89] br[89] wl[226] vdd gnd cell_6t
Xbit_r227_c89 bl[89] br[89] wl[227] vdd gnd cell_6t
Xbit_r228_c89 bl[89] br[89] wl[228] vdd gnd cell_6t
Xbit_r229_c89 bl[89] br[89] wl[229] vdd gnd cell_6t
Xbit_r230_c89 bl[89] br[89] wl[230] vdd gnd cell_6t
Xbit_r231_c89 bl[89] br[89] wl[231] vdd gnd cell_6t
Xbit_r232_c89 bl[89] br[89] wl[232] vdd gnd cell_6t
Xbit_r233_c89 bl[89] br[89] wl[233] vdd gnd cell_6t
Xbit_r234_c89 bl[89] br[89] wl[234] vdd gnd cell_6t
Xbit_r235_c89 bl[89] br[89] wl[235] vdd gnd cell_6t
Xbit_r236_c89 bl[89] br[89] wl[236] vdd gnd cell_6t
Xbit_r237_c89 bl[89] br[89] wl[237] vdd gnd cell_6t
Xbit_r238_c89 bl[89] br[89] wl[238] vdd gnd cell_6t
Xbit_r239_c89 bl[89] br[89] wl[239] vdd gnd cell_6t
Xbit_r240_c89 bl[89] br[89] wl[240] vdd gnd cell_6t
Xbit_r241_c89 bl[89] br[89] wl[241] vdd gnd cell_6t
Xbit_r242_c89 bl[89] br[89] wl[242] vdd gnd cell_6t
Xbit_r243_c89 bl[89] br[89] wl[243] vdd gnd cell_6t
Xbit_r244_c89 bl[89] br[89] wl[244] vdd gnd cell_6t
Xbit_r245_c89 bl[89] br[89] wl[245] vdd gnd cell_6t
Xbit_r246_c89 bl[89] br[89] wl[246] vdd gnd cell_6t
Xbit_r247_c89 bl[89] br[89] wl[247] vdd gnd cell_6t
Xbit_r248_c89 bl[89] br[89] wl[248] vdd gnd cell_6t
Xbit_r249_c89 bl[89] br[89] wl[249] vdd gnd cell_6t
Xbit_r250_c89 bl[89] br[89] wl[250] vdd gnd cell_6t
Xbit_r251_c89 bl[89] br[89] wl[251] vdd gnd cell_6t
Xbit_r252_c89 bl[89] br[89] wl[252] vdd gnd cell_6t
Xbit_r253_c89 bl[89] br[89] wl[253] vdd gnd cell_6t
Xbit_r254_c89 bl[89] br[89] wl[254] vdd gnd cell_6t
Xbit_r255_c89 bl[89] br[89] wl[255] vdd gnd cell_6t
Xbit_r256_c89 bl[89] br[89] wl[256] vdd gnd cell_6t
Xbit_r257_c89 bl[89] br[89] wl[257] vdd gnd cell_6t
Xbit_r258_c89 bl[89] br[89] wl[258] vdd gnd cell_6t
Xbit_r259_c89 bl[89] br[89] wl[259] vdd gnd cell_6t
Xbit_r260_c89 bl[89] br[89] wl[260] vdd gnd cell_6t
Xbit_r261_c89 bl[89] br[89] wl[261] vdd gnd cell_6t
Xbit_r262_c89 bl[89] br[89] wl[262] vdd gnd cell_6t
Xbit_r263_c89 bl[89] br[89] wl[263] vdd gnd cell_6t
Xbit_r264_c89 bl[89] br[89] wl[264] vdd gnd cell_6t
Xbit_r265_c89 bl[89] br[89] wl[265] vdd gnd cell_6t
Xbit_r266_c89 bl[89] br[89] wl[266] vdd gnd cell_6t
Xbit_r267_c89 bl[89] br[89] wl[267] vdd gnd cell_6t
Xbit_r268_c89 bl[89] br[89] wl[268] vdd gnd cell_6t
Xbit_r269_c89 bl[89] br[89] wl[269] vdd gnd cell_6t
Xbit_r270_c89 bl[89] br[89] wl[270] vdd gnd cell_6t
Xbit_r271_c89 bl[89] br[89] wl[271] vdd gnd cell_6t
Xbit_r272_c89 bl[89] br[89] wl[272] vdd gnd cell_6t
Xbit_r273_c89 bl[89] br[89] wl[273] vdd gnd cell_6t
Xbit_r274_c89 bl[89] br[89] wl[274] vdd gnd cell_6t
Xbit_r275_c89 bl[89] br[89] wl[275] vdd gnd cell_6t
Xbit_r276_c89 bl[89] br[89] wl[276] vdd gnd cell_6t
Xbit_r277_c89 bl[89] br[89] wl[277] vdd gnd cell_6t
Xbit_r278_c89 bl[89] br[89] wl[278] vdd gnd cell_6t
Xbit_r279_c89 bl[89] br[89] wl[279] vdd gnd cell_6t
Xbit_r280_c89 bl[89] br[89] wl[280] vdd gnd cell_6t
Xbit_r281_c89 bl[89] br[89] wl[281] vdd gnd cell_6t
Xbit_r282_c89 bl[89] br[89] wl[282] vdd gnd cell_6t
Xbit_r283_c89 bl[89] br[89] wl[283] vdd gnd cell_6t
Xbit_r284_c89 bl[89] br[89] wl[284] vdd gnd cell_6t
Xbit_r285_c89 bl[89] br[89] wl[285] vdd gnd cell_6t
Xbit_r286_c89 bl[89] br[89] wl[286] vdd gnd cell_6t
Xbit_r287_c89 bl[89] br[89] wl[287] vdd gnd cell_6t
Xbit_r288_c89 bl[89] br[89] wl[288] vdd gnd cell_6t
Xbit_r289_c89 bl[89] br[89] wl[289] vdd gnd cell_6t
Xbit_r290_c89 bl[89] br[89] wl[290] vdd gnd cell_6t
Xbit_r291_c89 bl[89] br[89] wl[291] vdd gnd cell_6t
Xbit_r292_c89 bl[89] br[89] wl[292] vdd gnd cell_6t
Xbit_r293_c89 bl[89] br[89] wl[293] vdd gnd cell_6t
Xbit_r294_c89 bl[89] br[89] wl[294] vdd gnd cell_6t
Xbit_r295_c89 bl[89] br[89] wl[295] vdd gnd cell_6t
Xbit_r296_c89 bl[89] br[89] wl[296] vdd gnd cell_6t
Xbit_r297_c89 bl[89] br[89] wl[297] vdd gnd cell_6t
Xbit_r298_c89 bl[89] br[89] wl[298] vdd gnd cell_6t
Xbit_r299_c89 bl[89] br[89] wl[299] vdd gnd cell_6t
Xbit_r300_c89 bl[89] br[89] wl[300] vdd gnd cell_6t
Xbit_r301_c89 bl[89] br[89] wl[301] vdd gnd cell_6t
Xbit_r302_c89 bl[89] br[89] wl[302] vdd gnd cell_6t
Xbit_r303_c89 bl[89] br[89] wl[303] vdd gnd cell_6t
Xbit_r304_c89 bl[89] br[89] wl[304] vdd gnd cell_6t
Xbit_r305_c89 bl[89] br[89] wl[305] vdd gnd cell_6t
Xbit_r306_c89 bl[89] br[89] wl[306] vdd gnd cell_6t
Xbit_r307_c89 bl[89] br[89] wl[307] vdd gnd cell_6t
Xbit_r308_c89 bl[89] br[89] wl[308] vdd gnd cell_6t
Xbit_r309_c89 bl[89] br[89] wl[309] vdd gnd cell_6t
Xbit_r310_c89 bl[89] br[89] wl[310] vdd gnd cell_6t
Xbit_r311_c89 bl[89] br[89] wl[311] vdd gnd cell_6t
Xbit_r312_c89 bl[89] br[89] wl[312] vdd gnd cell_6t
Xbit_r313_c89 bl[89] br[89] wl[313] vdd gnd cell_6t
Xbit_r314_c89 bl[89] br[89] wl[314] vdd gnd cell_6t
Xbit_r315_c89 bl[89] br[89] wl[315] vdd gnd cell_6t
Xbit_r316_c89 bl[89] br[89] wl[316] vdd gnd cell_6t
Xbit_r317_c89 bl[89] br[89] wl[317] vdd gnd cell_6t
Xbit_r318_c89 bl[89] br[89] wl[318] vdd gnd cell_6t
Xbit_r319_c89 bl[89] br[89] wl[319] vdd gnd cell_6t
Xbit_r320_c89 bl[89] br[89] wl[320] vdd gnd cell_6t
Xbit_r321_c89 bl[89] br[89] wl[321] vdd gnd cell_6t
Xbit_r322_c89 bl[89] br[89] wl[322] vdd gnd cell_6t
Xbit_r323_c89 bl[89] br[89] wl[323] vdd gnd cell_6t
Xbit_r324_c89 bl[89] br[89] wl[324] vdd gnd cell_6t
Xbit_r325_c89 bl[89] br[89] wl[325] vdd gnd cell_6t
Xbit_r326_c89 bl[89] br[89] wl[326] vdd gnd cell_6t
Xbit_r327_c89 bl[89] br[89] wl[327] vdd gnd cell_6t
Xbit_r328_c89 bl[89] br[89] wl[328] vdd gnd cell_6t
Xbit_r329_c89 bl[89] br[89] wl[329] vdd gnd cell_6t
Xbit_r330_c89 bl[89] br[89] wl[330] vdd gnd cell_6t
Xbit_r331_c89 bl[89] br[89] wl[331] vdd gnd cell_6t
Xbit_r332_c89 bl[89] br[89] wl[332] vdd gnd cell_6t
Xbit_r333_c89 bl[89] br[89] wl[333] vdd gnd cell_6t
Xbit_r334_c89 bl[89] br[89] wl[334] vdd gnd cell_6t
Xbit_r335_c89 bl[89] br[89] wl[335] vdd gnd cell_6t
Xbit_r336_c89 bl[89] br[89] wl[336] vdd gnd cell_6t
Xbit_r337_c89 bl[89] br[89] wl[337] vdd gnd cell_6t
Xbit_r338_c89 bl[89] br[89] wl[338] vdd gnd cell_6t
Xbit_r339_c89 bl[89] br[89] wl[339] vdd gnd cell_6t
Xbit_r340_c89 bl[89] br[89] wl[340] vdd gnd cell_6t
Xbit_r341_c89 bl[89] br[89] wl[341] vdd gnd cell_6t
Xbit_r342_c89 bl[89] br[89] wl[342] vdd gnd cell_6t
Xbit_r343_c89 bl[89] br[89] wl[343] vdd gnd cell_6t
Xbit_r344_c89 bl[89] br[89] wl[344] vdd gnd cell_6t
Xbit_r345_c89 bl[89] br[89] wl[345] vdd gnd cell_6t
Xbit_r346_c89 bl[89] br[89] wl[346] vdd gnd cell_6t
Xbit_r347_c89 bl[89] br[89] wl[347] vdd gnd cell_6t
Xbit_r348_c89 bl[89] br[89] wl[348] vdd gnd cell_6t
Xbit_r349_c89 bl[89] br[89] wl[349] vdd gnd cell_6t
Xbit_r350_c89 bl[89] br[89] wl[350] vdd gnd cell_6t
Xbit_r351_c89 bl[89] br[89] wl[351] vdd gnd cell_6t
Xbit_r352_c89 bl[89] br[89] wl[352] vdd gnd cell_6t
Xbit_r353_c89 bl[89] br[89] wl[353] vdd gnd cell_6t
Xbit_r354_c89 bl[89] br[89] wl[354] vdd gnd cell_6t
Xbit_r355_c89 bl[89] br[89] wl[355] vdd gnd cell_6t
Xbit_r356_c89 bl[89] br[89] wl[356] vdd gnd cell_6t
Xbit_r357_c89 bl[89] br[89] wl[357] vdd gnd cell_6t
Xbit_r358_c89 bl[89] br[89] wl[358] vdd gnd cell_6t
Xbit_r359_c89 bl[89] br[89] wl[359] vdd gnd cell_6t
Xbit_r360_c89 bl[89] br[89] wl[360] vdd gnd cell_6t
Xbit_r361_c89 bl[89] br[89] wl[361] vdd gnd cell_6t
Xbit_r362_c89 bl[89] br[89] wl[362] vdd gnd cell_6t
Xbit_r363_c89 bl[89] br[89] wl[363] vdd gnd cell_6t
Xbit_r364_c89 bl[89] br[89] wl[364] vdd gnd cell_6t
Xbit_r365_c89 bl[89] br[89] wl[365] vdd gnd cell_6t
Xbit_r366_c89 bl[89] br[89] wl[366] vdd gnd cell_6t
Xbit_r367_c89 bl[89] br[89] wl[367] vdd gnd cell_6t
Xbit_r368_c89 bl[89] br[89] wl[368] vdd gnd cell_6t
Xbit_r369_c89 bl[89] br[89] wl[369] vdd gnd cell_6t
Xbit_r370_c89 bl[89] br[89] wl[370] vdd gnd cell_6t
Xbit_r371_c89 bl[89] br[89] wl[371] vdd gnd cell_6t
Xbit_r372_c89 bl[89] br[89] wl[372] vdd gnd cell_6t
Xbit_r373_c89 bl[89] br[89] wl[373] vdd gnd cell_6t
Xbit_r374_c89 bl[89] br[89] wl[374] vdd gnd cell_6t
Xbit_r375_c89 bl[89] br[89] wl[375] vdd gnd cell_6t
Xbit_r376_c89 bl[89] br[89] wl[376] vdd gnd cell_6t
Xbit_r377_c89 bl[89] br[89] wl[377] vdd gnd cell_6t
Xbit_r378_c89 bl[89] br[89] wl[378] vdd gnd cell_6t
Xbit_r379_c89 bl[89] br[89] wl[379] vdd gnd cell_6t
Xbit_r380_c89 bl[89] br[89] wl[380] vdd gnd cell_6t
Xbit_r381_c89 bl[89] br[89] wl[381] vdd gnd cell_6t
Xbit_r382_c89 bl[89] br[89] wl[382] vdd gnd cell_6t
Xbit_r383_c89 bl[89] br[89] wl[383] vdd gnd cell_6t
Xbit_r384_c89 bl[89] br[89] wl[384] vdd gnd cell_6t
Xbit_r385_c89 bl[89] br[89] wl[385] vdd gnd cell_6t
Xbit_r386_c89 bl[89] br[89] wl[386] vdd gnd cell_6t
Xbit_r387_c89 bl[89] br[89] wl[387] vdd gnd cell_6t
Xbit_r388_c89 bl[89] br[89] wl[388] vdd gnd cell_6t
Xbit_r389_c89 bl[89] br[89] wl[389] vdd gnd cell_6t
Xbit_r390_c89 bl[89] br[89] wl[390] vdd gnd cell_6t
Xbit_r391_c89 bl[89] br[89] wl[391] vdd gnd cell_6t
Xbit_r392_c89 bl[89] br[89] wl[392] vdd gnd cell_6t
Xbit_r393_c89 bl[89] br[89] wl[393] vdd gnd cell_6t
Xbit_r394_c89 bl[89] br[89] wl[394] vdd gnd cell_6t
Xbit_r395_c89 bl[89] br[89] wl[395] vdd gnd cell_6t
Xbit_r396_c89 bl[89] br[89] wl[396] vdd gnd cell_6t
Xbit_r397_c89 bl[89] br[89] wl[397] vdd gnd cell_6t
Xbit_r398_c89 bl[89] br[89] wl[398] vdd gnd cell_6t
Xbit_r399_c89 bl[89] br[89] wl[399] vdd gnd cell_6t
Xbit_r400_c89 bl[89] br[89] wl[400] vdd gnd cell_6t
Xbit_r401_c89 bl[89] br[89] wl[401] vdd gnd cell_6t
Xbit_r402_c89 bl[89] br[89] wl[402] vdd gnd cell_6t
Xbit_r403_c89 bl[89] br[89] wl[403] vdd gnd cell_6t
Xbit_r404_c89 bl[89] br[89] wl[404] vdd gnd cell_6t
Xbit_r405_c89 bl[89] br[89] wl[405] vdd gnd cell_6t
Xbit_r406_c89 bl[89] br[89] wl[406] vdd gnd cell_6t
Xbit_r407_c89 bl[89] br[89] wl[407] vdd gnd cell_6t
Xbit_r408_c89 bl[89] br[89] wl[408] vdd gnd cell_6t
Xbit_r409_c89 bl[89] br[89] wl[409] vdd gnd cell_6t
Xbit_r410_c89 bl[89] br[89] wl[410] vdd gnd cell_6t
Xbit_r411_c89 bl[89] br[89] wl[411] vdd gnd cell_6t
Xbit_r412_c89 bl[89] br[89] wl[412] vdd gnd cell_6t
Xbit_r413_c89 bl[89] br[89] wl[413] vdd gnd cell_6t
Xbit_r414_c89 bl[89] br[89] wl[414] vdd gnd cell_6t
Xbit_r415_c89 bl[89] br[89] wl[415] vdd gnd cell_6t
Xbit_r416_c89 bl[89] br[89] wl[416] vdd gnd cell_6t
Xbit_r417_c89 bl[89] br[89] wl[417] vdd gnd cell_6t
Xbit_r418_c89 bl[89] br[89] wl[418] vdd gnd cell_6t
Xbit_r419_c89 bl[89] br[89] wl[419] vdd gnd cell_6t
Xbit_r420_c89 bl[89] br[89] wl[420] vdd gnd cell_6t
Xbit_r421_c89 bl[89] br[89] wl[421] vdd gnd cell_6t
Xbit_r422_c89 bl[89] br[89] wl[422] vdd gnd cell_6t
Xbit_r423_c89 bl[89] br[89] wl[423] vdd gnd cell_6t
Xbit_r424_c89 bl[89] br[89] wl[424] vdd gnd cell_6t
Xbit_r425_c89 bl[89] br[89] wl[425] vdd gnd cell_6t
Xbit_r426_c89 bl[89] br[89] wl[426] vdd gnd cell_6t
Xbit_r427_c89 bl[89] br[89] wl[427] vdd gnd cell_6t
Xbit_r428_c89 bl[89] br[89] wl[428] vdd gnd cell_6t
Xbit_r429_c89 bl[89] br[89] wl[429] vdd gnd cell_6t
Xbit_r430_c89 bl[89] br[89] wl[430] vdd gnd cell_6t
Xbit_r431_c89 bl[89] br[89] wl[431] vdd gnd cell_6t
Xbit_r432_c89 bl[89] br[89] wl[432] vdd gnd cell_6t
Xbit_r433_c89 bl[89] br[89] wl[433] vdd gnd cell_6t
Xbit_r434_c89 bl[89] br[89] wl[434] vdd gnd cell_6t
Xbit_r435_c89 bl[89] br[89] wl[435] vdd gnd cell_6t
Xbit_r436_c89 bl[89] br[89] wl[436] vdd gnd cell_6t
Xbit_r437_c89 bl[89] br[89] wl[437] vdd gnd cell_6t
Xbit_r438_c89 bl[89] br[89] wl[438] vdd gnd cell_6t
Xbit_r439_c89 bl[89] br[89] wl[439] vdd gnd cell_6t
Xbit_r440_c89 bl[89] br[89] wl[440] vdd gnd cell_6t
Xbit_r441_c89 bl[89] br[89] wl[441] vdd gnd cell_6t
Xbit_r442_c89 bl[89] br[89] wl[442] vdd gnd cell_6t
Xbit_r443_c89 bl[89] br[89] wl[443] vdd gnd cell_6t
Xbit_r444_c89 bl[89] br[89] wl[444] vdd gnd cell_6t
Xbit_r445_c89 bl[89] br[89] wl[445] vdd gnd cell_6t
Xbit_r446_c89 bl[89] br[89] wl[446] vdd gnd cell_6t
Xbit_r447_c89 bl[89] br[89] wl[447] vdd gnd cell_6t
Xbit_r448_c89 bl[89] br[89] wl[448] vdd gnd cell_6t
Xbit_r449_c89 bl[89] br[89] wl[449] vdd gnd cell_6t
Xbit_r450_c89 bl[89] br[89] wl[450] vdd gnd cell_6t
Xbit_r451_c89 bl[89] br[89] wl[451] vdd gnd cell_6t
Xbit_r452_c89 bl[89] br[89] wl[452] vdd gnd cell_6t
Xbit_r453_c89 bl[89] br[89] wl[453] vdd gnd cell_6t
Xbit_r454_c89 bl[89] br[89] wl[454] vdd gnd cell_6t
Xbit_r455_c89 bl[89] br[89] wl[455] vdd gnd cell_6t
Xbit_r456_c89 bl[89] br[89] wl[456] vdd gnd cell_6t
Xbit_r457_c89 bl[89] br[89] wl[457] vdd gnd cell_6t
Xbit_r458_c89 bl[89] br[89] wl[458] vdd gnd cell_6t
Xbit_r459_c89 bl[89] br[89] wl[459] vdd gnd cell_6t
Xbit_r460_c89 bl[89] br[89] wl[460] vdd gnd cell_6t
Xbit_r461_c89 bl[89] br[89] wl[461] vdd gnd cell_6t
Xbit_r462_c89 bl[89] br[89] wl[462] vdd gnd cell_6t
Xbit_r463_c89 bl[89] br[89] wl[463] vdd gnd cell_6t
Xbit_r464_c89 bl[89] br[89] wl[464] vdd gnd cell_6t
Xbit_r465_c89 bl[89] br[89] wl[465] vdd gnd cell_6t
Xbit_r466_c89 bl[89] br[89] wl[466] vdd gnd cell_6t
Xbit_r467_c89 bl[89] br[89] wl[467] vdd gnd cell_6t
Xbit_r468_c89 bl[89] br[89] wl[468] vdd gnd cell_6t
Xbit_r469_c89 bl[89] br[89] wl[469] vdd gnd cell_6t
Xbit_r470_c89 bl[89] br[89] wl[470] vdd gnd cell_6t
Xbit_r471_c89 bl[89] br[89] wl[471] vdd gnd cell_6t
Xbit_r472_c89 bl[89] br[89] wl[472] vdd gnd cell_6t
Xbit_r473_c89 bl[89] br[89] wl[473] vdd gnd cell_6t
Xbit_r474_c89 bl[89] br[89] wl[474] vdd gnd cell_6t
Xbit_r475_c89 bl[89] br[89] wl[475] vdd gnd cell_6t
Xbit_r476_c89 bl[89] br[89] wl[476] vdd gnd cell_6t
Xbit_r477_c89 bl[89] br[89] wl[477] vdd gnd cell_6t
Xbit_r478_c89 bl[89] br[89] wl[478] vdd gnd cell_6t
Xbit_r479_c89 bl[89] br[89] wl[479] vdd gnd cell_6t
Xbit_r480_c89 bl[89] br[89] wl[480] vdd gnd cell_6t
Xbit_r481_c89 bl[89] br[89] wl[481] vdd gnd cell_6t
Xbit_r482_c89 bl[89] br[89] wl[482] vdd gnd cell_6t
Xbit_r483_c89 bl[89] br[89] wl[483] vdd gnd cell_6t
Xbit_r484_c89 bl[89] br[89] wl[484] vdd gnd cell_6t
Xbit_r485_c89 bl[89] br[89] wl[485] vdd gnd cell_6t
Xbit_r486_c89 bl[89] br[89] wl[486] vdd gnd cell_6t
Xbit_r487_c89 bl[89] br[89] wl[487] vdd gnd cell_6t
Xbit_r488_c89 bl[89] br[89] wl[488] vdd gnd cell_6t
Xbit_r489_c89 bl[89] br[89] wl[489] vdd gnd cell_6t
Xbit_r490_c89 bl[89] br[89] wl[490] vdd gnd cell_6t
Xbit_r491_c89 bl[89] br[89] wl[491] vdd gnd cell_6t
Xbit_r492_c89 bl[89] br[89] wl[492] vdd gnd cell_6t
Xbit_r493_c89 bl[89] br[89] wl[493] vdd gnd cell_6t
Xbit_r494_c89 bl[89] br[89] wl[494] vdd gnd cell_6t
Xbit_r495_c89 bl[89] br[89] wl[495] vdd gnd cell_6t
Xbit_r496_c89 bl[89] br[89] wl[496] vdd gnd cell_6t
Xbit_r497_c89 bl[89] br[89] wl[497] vdd gnd cell_6t
Xbit_r498_c89 bl[89] br[89] wl[498] vdd gnd cell_6t
Xbit_r499_c89 bl[89] br[89] wl[499] vdd gnd cell_6t
Xbit_r500_c89 bl[89] br[89] wl[500] vdd gnd cell_6t
Xbit_r501_c89 bl[89] br[89] wl[501] vdd gnd cell_6t
Xbit_r502_c89 bl[89] br[89] wl[502] vdd gnd cell_6t
Xbit_r503_c89 bl[89] br[89] wl[503] vdd gnd cell_6t
Xbit_r504_c89 bl[89] br[89] wl[504] vdd gnd cell_6t
Xbit_r505_c89 bl[89] br[89] wl[505] vdd gnd cell_6t
Xbit_r506_c89 bl[89] br[89] wl[506] vdd gnd cell_6t
Xbit_r507_c89 bl[89] br[89] wl[507] vdd gnd cell_6t
Xbit_r508_c89 bl[89] br[89] wl[508] vdd gnd cell_6t
Xbit_r509_c89 bl[89] br[89] wl[509] vdd gnd cell_6t
Xbit_r510_c89 bl[89] br[89] wl[510] vdd gnd cell_6t
Xbit_r511_c89 bl[89] br[89] wl[511] vdd gnd cell_6t
Xbit_r0_c90 bl[90] br[90] wl[0] vdd gnd cell_6t
Xbit_r1_c90 bl[90] br[90] wl[1] vdd gnd cell_6t
Xbit_r2_c90 bl[90] br[90] wl[2] vdd gnd cell_6t
Xbit_r3_c90 bl[90] br[90] wl[3] vdd gnd cell_6t
Xbit_r4_c90 bl[90] br[90] wl[4] vdd gnd cell_6t
Xbit_r5_c90 bl[90] br[90] wl[5] vdd gnd cell_6t
Xbit_r6_c90 bl[90] br[90] wl[6] vdd gnd cell_6t
Xbit_r7_c90 bl[90] br[90] wl[7] vdd gnd cell_6t
Xbit_r8_c90 bl[90] br[90] wl[8] vdd gnd cell_6t
Xbit_r9_c90 bl[90] br[90] wl[9] vdd gnd cell_6t
Xbit_r10_c90 bl[90] br[90] wl[10] vdd gnd cell_6t
Xbit_r11_c90 bl[90] br[90] wl[11] vdd gnd cell_6t
Xbit_r12_c90 bl[90] br[90] wl[12] vdd gnd cell_6t
Xbit_r13_c90 bl[90] br[90] wl[13] vdd gnd cell_6t
Xbit_r14_c90 bl[90] br[90] wl[14] vdd gnd cell_6t
Xbit_r15_c90 bl[90] br[90] wl[15] vdd gnd cell_6t
Xbit_r16_c90 bl[90] br[90] wl[16] vdd gnd cell_6t
Xbit_r17_c90 bl[90] br[90] wl[17] vdd gnd cell_6t
Xbit_r18_c90 bl[90] br[90] wl[18] vdd gnd cell_6t
Xbit_r19_c90 bl[90] br[90] wl[19] vdd gnd cell_6t
Xbit_r20_c90 bl[90] br[90] wl[20] vdd gnd cell_6t
Xbit_r21_c90 bl[90] br[90] wl[21] vdd gnd cell_6t
Xbit_r22_c90 bl[90] br[90] wl[22] vdd gnd cell_6t
Xbit_r23_c90 bl[90] br[90] wl[23] vdd gnd cell_6t
Xbit_r24_c90 bl[90] br[90] wl[24] vdd gnd cell_6t
Xbit_r25_c90 bl[90] br[90] wl[25] vdd gnd cell_6t
Xbit_r26_c90 bl[90] br[90] wl[26] vdd gnd cell_6t
Xbit_r27_c90 bl[90] br[90] wl[27] vdd gnd cell_6t
Xbit_r28_c90 bl[90] br[90] wl[28] vdd gnd cell_6t
Xbit_r29_c90 bl[90] br[90] wl[29] vdd gnd cell_6t
Xbit_r30_c90 bl[90] br[90] wl[30] vdd gnd cell_6t
Xbit_r31_c90 bl[90] br[90] wl[31] vdd gnd cell_6t
Xbit_r32_c90 bl[90] br[90] wl[32] vdd gnd cell_6t
Xbit_r33_c90 bl[90] br[90] wl[33] vdd gnd cell_6t
Xbit_r34_c90 bl[90] br[90] wl[34] vdd gnd cell_6t
Xbit_r35_c90 bl[90] br[90] wl[35] vdd gnd cell_6t
Xbit_r36_c90 bl[90] br[90] wl[36] vdd gnd cell_6t
Xbit_r37_c90 bl[90] br[90] wl[37] vdd gnd cell_6t
Xbit_r38_c90 bl[90] br[90] wl[38] vdd gnd cell_6t
Xbit_r39_c90 bl[90] br[90] wl[39] vdd gnd cell_6t
Xbit_r40_c90 bl[90] br[90] wl[40] vdd gnd cell_6t
Xbit_r41_c90 bl[90] br[90] wl[41] vdd gnd cell_6t
Xbit_r42_c90 bl[90] br[90] wl[42] vdd gnd cell_6t
Xbit_r43_c90 bl[90] br[90] wl[43] vdd gnd cell_6t
Xbit_r44_c90 bl[90] br[90] wl[44] vdd gnd cell_6t
Xbit_r45_c90 bl[90] br[90] wl[45] vdd gnd cell_6t
Xbit_r46_c90 bl[90] br[90] wl[46] vdd gnd cell_6t
Xbit_r47_c90 bl[90] br[90] wl[47] vdd gnd cell_6t
Xbit_r48_c90 bl[90] br[90] wl[48] vdd gnd cell_6t
Xbit_r49_c90 bl[90] br[90] wl[49] vdd gnd cell_6t
Xbit_r50_c90 bl[90] br[90] wl[50] vdd gnd cell_6t
Xbit_r51_c90 bl[90] br[90] wl[51] vdd gnd cell_6t
Xbit_r52_c90 bl[90] br[90] wl[52] vdd gnd cell_6t
Xbit_r53_c90 bl[90] br[90] wl[53] vdd gnd cell_6t
Xbit_r54_c90 bl[90] br[90] wl[54] vdd gnd cell_6t
Xbit_r55_c90 bl[90] br[90] wl[55] vdd gnd cell_6t
Xbit_r56_c90 bl[90] br[90] wl[56] vdd gnd cell_6t
Xbit_r57_c90 bl[90] br[90] wl[57] vdd gnd cell_6t
Xbit_r58_c90 bl[90] br[90] wl[58] vdd gnd cell_6t
Xbit_r59_c90 bl[90] br[90] wl[59] vdd gnd cell_6t
Xbit_r60_c90 bl[90] br[90] wl[60] vdd gnd cell_6t
Xbit_r61_c90 bl[90] br[90] wl[61] vdd gnd cell_6t
Xbit_r62_c90 bl[90] br[90] wl[62] vdd gnd cell_6t
Xbit_r63_c90 bl[90] br[90] wl[63] vdd gnd cell_6t
Xbit_r64_c90 bl[90] br[90] wl[64] vdd gnd cell_6t
Xbit_r65_c90 bl[90] br[90] wl[65] vdd gnd cell_6t
Xbit_r66_c90 bl[90] br[90] wl[66] vdd gnd cell_6t
Xbit_r67_c90 bl[90] br[90] wl[67] vdd gnd cell_6t
Xbit_r68_c90 bl[90] br[90] wl[68] vdd gnd cell_6t
Xbit_r69_c90 bl[90] br[90] wl[69] vdd gnd cell_6t
Xbit_r70_c90 bl[90] br[90] wl[70] vdd gnd cell_6t
Xbit_r71_c90 bl[90] br[90] wl[71] vdd gnd cell_6t
Xbit_r72_c90 bl[90] br[90] wl[72] vdd gnd cell_6t
Xbit_r73_c90 bl[90] br[90] wl[73] vdd gnd cell_6t
Xbit_r74_c90 bl[90] br[90] wl[74] vdd gnd cell_6t
Xbit_r75_c90 bl[90] br[90] wl[75] vdd gnd cell_6t
Xbit_r76_c90 bl[90] br[90] wl[76] vdd gnd cell_6t
Xbit_r77_c90 bl[90] br[90] wl[77] vdd gnd cell_6t
Xbit_r78_c90 bl[90] br[90] wl[78] vdd gnd cell_6t
Xbit_r79_c90 bl[90] br[90] wl[79] vdd gnd cell_6t
Xbit_r80_c90 bl[90] br[90] wl[80] vdd gnd cell_6t
Xbit_r81_c90 bl[90] br[90] wl[81] vdd gnd cell_6t
Xbit_r82_c90 bl[90] br[90] wl[82] vdd gnd cell_6t
Xbit_r83_c90 bl[90] br[90] wl[83] vdd gnd cell_6t
Xbit_r84_c90 bl[90] br[90] wl[84] vdd gnd cell_6t
Xbit_r85_c90 bl[90] br[90] wl[85] vdd gnd cell_6t
Xbit_r86_c90 bl[90] br[90] wl[86] vdd gnd cell_6t
Xbit_r87_c90 bl[90] br[90] wl[87] vdd gnd cell_6t
Xbit_r88_c90 bl[90] br[90] wl[88] vdd gnd cell_6t
Xbit_r89_c90 bl[90] br[90] wl[89] vdd gnd cell_6t
Xbit_r90_c90 bl[90] br[90] wl[90] vdd gnd cell_6t
Xbit_r91_c90 bl[90] br[90] wl[91] vdd gnd cell_6t
Xbit_r92_c90 bl[90] br[90] wl[92] vdd gnd cell_6t
Xbit_r93_c90 bl[90] br[90] wl[93] vdd gnd cell_6t
Xbit_r94_c90 bl[90] br[90] wl[94] vdd gnd cell_6t
Xbit_r95_c90 bl[90] br[90] wl[95] vdd gnd cell_6t
Xbit_r96_c90 bl[90] br[90] wl[96] vdd gnd cell_6t
Xbit_r97_c90 bl[90] br[90] wl[97] vdd gnd cell_6t
Xbit_r98_c90 bl[90] br[90] wl[98] vdd gnd cell_6t
Xbit_r99_c90 bl[90] br[90] wl[99] vdd gnd cell_6t
Xbit_r100_c90 bl[90] br[90] wl[100] vdd gnd cell_6t
Xbit_r101_c90 bl[90] br[90] wl[101] vdd gnd cell_6t
Xbit_r102_c90 bl[90] br[90] wl[102] vdd gnd cell_6t
Xbit_r103_c90 bl[90] br[90] wl[103] vdd gnd cell_6t
Xbit_r104_c90 bl[90] br[90] wl[104] vdd gnd cell_6t
Xbit_r105_c90 bl[90] br[90] wl[105] vdd gnd cell_6t
Xbit_r106_c90 bl[90] br[90] wl[106] vdd gnd cell_6t
Xbit_r107_c90 bl[90] br[90] wl[107] vdd gnd cell_6t
Xbit_r108_c90 bl[90] br[90] wl[108] vdd gnd cell_6t
Xbit_r109_c90 bl[90] br[90] wl[109] vdd gnd cell_6t
Xbit_r110_c90 bl[90] br[90] wl[110] vdd gnd cell_6t
Xbit_r111_c90 bl[90] br[90] wl[111] vdd gnd cell_6t
Xbit_r112_c90 bl[90] br[90] wl[112] vdd gnd cell_6t
Xbit_r113_c90 bl[90] br[90] wl[113] vdd gnd cell_6t
Xbit_r114_c90 bl[90] br[90] wl[114] vdd gnd cell_6t
Xbit_r115_c90 bl[90] br[90] wl[115] vdd gnd cell_6t
Xbit_r116_c90 bl[90] br[90] wl[116] vdd gnd cell_6t
Xbit_r117_c90 bl[90] br[90] wl[117] vdd gnd cell_6t
Xbit_r118_c90 bl[90] br[90] wl[118] vdd gnd cell_6t
Xbit_r119_c90 bl[90] br[90] wl[119] vdd gnd cell_6t
Xbit_r120_c90 bl[90] br[90] wl[120] vdd gnd cell_6t
Xbit_r121_c90 bl[90] br[90] wl[121] vdd gnd cell_6t
Xbit_r122_c90 bl[90] br[90] wl[122] vdd gnd cell_6t
Xbit_r123_c90 bl[90] br[90] wl[123] vdd gnd cell_6t
Xbit_r124_c90 bl[90] br[90] wl[124] vdd gnd cell_6t
Xbit_r125_c90 bl[90] br[90] wl[125] vdd gnd cell_6t
Xbit_r126_c90 bl[90] br[90] wl[126] vdd gnd cell_6t
Xbit_r127_c90 bl[90] br[90] wl[127] vdd gnd cell_6t
Xbit_r128_c90 bl[90] br[90] wl[128] vdd gnd cell_6t
Xbit_r129_c90 bl[90] br[90] wl[129] vdd gnd cell_6t
Xbit_r130_c90 bl[90] br[90] wl[130] vdd gnd cell_6t
Xbit_r131_c90 bl[90] br[90] wl[131] vdd gnd cell_6t
Xbit_r132_c90 bl[90] br[90] wl[132] vdd gnd cell_6t
Xbit_r133_c90 bl[90] br[90] wl[133] vdd gnd cell_6t
Xbit_r134_c90 bl[90] br[90] wl[134] vdd gnd cell_6t
Xbit_r135_c90 bl[90] br[90] wl[135] vdd gnd cell_6t
Xbit_r136_c90 bl[90] br[90] wl[136] vdd gnd cell_6t
Xbit_r137_c90 bl[90] br[90] wl[137] vdd gnd cell_6t
Xbit_r138_c90 bl[90] br[90] wl[138] vdd gnd cell_6t
Xbit_r139_c90 bl[90] br[90] wl[139] vdd gnd cell_6t
Xbit_r140_c90 bl[90] br[90] wl[140] vdd gnd cell_6t
Xbit_r141_c90 bl[90] br[90] wl[141] vdd gnd cell_6t
Xbit_r142_c90 bl[90] br[90] wl[142] vdd gnd cell_6t
Xbit_r143_c90 bl[90] br[90] wl[143] vdd gnd cell_6t
Xbit_r144_c90 bl[90] br[90] wl[144] vdd gnd cell_6t
Xbit_r145_c90 bl[90] br[90] wl[145] vdd gnd cell_6t
Xbit_r146_c90 bl[90] br[90] wl[146] vdd gnd cell_6t
Xbit_r147_c90 bl[90] br[90] wl[147] vdd gnd cell_6t
Xbit_r148_c90 bl[90] br[90] wl[148] vdd gnd cell_6t
Xbit_r149_c90 bl[90] br[90] wl[149] vdd gnd cell_6t
Xbit_r150_c90 bl[90] br[90] wl[150] vdd gnd cell_6t
Xbit_r151_c90 bl[90] br[90] wl[151] vdd gnd cell_6t
Xbit_r152_c90 bl[90] br[90] wl[152] vdd gnd cell_6t
Xbit_r153_c90 bl[90] br[90] wl[153] vdd gnd cell_6t
Xbit_r154_c90 bl[90] br[90] wl[154] vdd gnd cell_6t
Xbit_r155_c90 bl[90] br[90] wl[155] vdd gnd cell_6t
Xbit_r156_c90 bl[90] br[90] wl[156] vdd gnd cell_6t
Xbit_r157_c90 bl[90] br[90] wl[157] vdd gnd cell_6t
Xbit_r158_c90 bl[90] br[90] wl[158] vdd gnd cell_6t
Xbit_r159_c90 bl[90] br[90] wl[159] vdd gnd cell_6t
Xbit_r160_c90 bl[90] br[90] wl[160] vdd gnd cell_6t
Xbit_r161_c90 bl[90] br[90] wl[161] vdd gnd cell_6t
Xbit_r162_c90 bl[90] br[90] wl[162] vdd gnd cell_6t
Xbit_r163_c90 bl[90] br[90] wl[163] vdd gnd cell_6t
Xbit_r164_c90 bl[90] br[90] wl[164] vdd gnd cell_6t
Xbit_r165_c90 bl[90] br[90] wl[165] vdd gnd cell_6t
Xbit_r166_c90 bl[90] br[90] wl[166] vdd gnd cell_6t
Xbit_r167_c90 bl[90] br[90] wl[167] vdd gnd cell_6t
Xbit_r168_c90 bl[90] br[90] wl[168] vdd gnd cell_6t
Xbit_r169_c90 bl[90] br[90] wl[169] vdd gnd cell_6t
Xbit_r170_c90 bl[90] br[90] wl[170] vdd gnd cell_6t
Xbit_r171_c90 bl[90] br[90] wl[171] vdd gnd cell_6t
Xbit_r172_c90 bl[90] br[90] wl[172] vdd gnd cell_6t
Xbit_r173_c90 bl[90] br[90] wl[173] vdd gnd cell_6t
Xbit_r174_c90 bl[90] br[90] wl[174] vdd gnd cell_6t
Xbit_r175_c90 bl[90] br[90] wl[175] vdd gnd cell_6t
Xbit_r176_c90 bl[90] br[90] wl[176] vdd gnd cell_6t
Xbit_r177_c90 bl[90] br[90] wl[177] vdd gnd cell_6t
Xbit_r178_c90 bl[90] br[90] wl[178] vdd gnd cell_6t
Xbit_r179_c90 bl[90] br[90] wl[179] vdd gnd cell_6t
Xbit_r180_c90 bl[90] br[90] wl[180] vdd gnd cell_6t
Xbit_r181_c90 bl[90] br[90] wl[181] vdd gnd cell_6t
Xbit_r182_c90 bl[90] br[90] wl[182] vdd gnd cell_6t
Xbit_r183_c90 bl[90] br[90] wl[183] vdd gnd cell_6t
Xbit_r184_c90 bl[90] br[90] wl[184] vdd gnd cell_6t
Xbit_r185_c90 bl[90] br[90] wl[185] vdd gnd cell_6t
Xbit_r186_c90 bl[90] br[90] wl[186] vdd gnd cell_6t
Xbit_r187_c90 bl[90] br[90] wl[187] vdd gnd cell_6t
Xbit_r188_c90 bl[90] br[90] wl[188] vdd gnd cell_6t
Xbit_r189_c90 bl[90] br[90] wl[189] vdd gnd cell_6t
Xbit_r190_c90 bl[90] br[90] wl[190] vdd gnd cell_6t
Xbit_r191_c90 bl[90] br[90] wl[191] vdd gnd cell_6t
Xbit_r192_c90 bl[90] br[90] wl[192] vdd gnd cell_6t
Xbit_r193_c90 bl[90] br[90] wl[193] vdd gnd cell_6t
Xbit_r194_c90 bl[90] br[90] wl[194] vdd gnd cell_6t
Xbit_r195_c90 bl[90] br[90] wl[195] vdd gnd cell_6t
Xbit_r196_c90 bl[90] br[90] wl[196] vdd gnd cell_6t
Xbit_r197_c90 bl[90] br[90] wl[197] vdd gnd cell_6t
Xbit_r198_c90 bl[90] br[90] wl[198] vdd gnd cell_6t
Xbit_r199_c90 bl[90] br[90] wl[199] vdd gnd cell_6t
Xbit_r200_c90 bl[90] br[90] wl[200] vdd gnd cell_6t
Xbit_r201_c90 bl[90] br[90] wl[201] vdd gnd cell_6t
Xbit_r202_c90 bl[90] br[90] wl[202] vdd gnd cell_6t
Xbit_r203_c90 bl[90] br[90] wl[203] vdd gnd cell_6t
Xbit_r204_c90 bl[90] br[90] wl[204] vdd gnd cell_6t
Xbit_r205_c90 bl[90] br[90] wl[205] vdd gnd cell_6t
Xbit_r206_c90 bl[90] br[90] wl[206] vdd gnd cell_6t
Xbit_r207_c90 bl[90] br[90] wl[207] vdd gnd cell_6t
Xbit_r208_c90 bl[90] br[90] wl[208] vdd gnd cell_6t
Xbit_r209_c90 bl[90] br[90] wl[209] vdd gnd cell_6t
Xbit_r210_c90 bl[90] br[90] wl[210] vdd gnd cell_6t
Xbit_r211_c90 bl[90] br[90] wl[211] vdd gnd cell_6t
Xbit_r212_c90 bl[90] br[90] wl[212] vdd gnd cell_6t
Xbit_r213_c90 bl[90] br[90] wl[213] vdd gnd cell_6t
Xbit_r214_c90 bl[90] br[90] wl[214] vdd gnd cell_6t
Xbit_r215_c90 bl[90] br[90] wl[215] vdd gnd cell_6t
Xbit_r216_c90 bl[90] br[90] wl[216] vdd gnd cell_6t
Xbit_r217_c90 bl[90] br[90] wl[217] vdd gnd cell_6t
Xbit_r218_c90 bl[90] br[90] wl[218] vdd gnd cell_6t
Xbit_r219_c90 bl[90] br[90] wl[219] vdd gnd cell_6t
Xbit_r220_c90 bl[90] br[90] wl[220] vdd gnd cell_6t
Xbit_r221_c90 bl[90] br[90] wl[221] vdd gnd cell_6t
Xbit_r222_c90 bl[90] br[90] wl[222] vdd gnd cell_6t
Xbit_r223_c90 bl[90] br[90] wl[223] vdd gnd cell_6t
Xbit_r224_c90 bl[90] br[90] wl[224] vdd gnd cell_6t
Xbit_r225_c90 bl[90] br[90] wl[225] vdd gnd cell_6t
Xbit_r226_c90 bl[90] br[90] wl[226] vdd gnd cell_6t
Xbit_r227_c90 bl[90] br[90] wl[227] vdd gnd cell_6t
Xbit_r228_c90 bl[90] br[90] wl[228] vdd gnd cell_6t
Xbit_r229_c90 bl[90] br[90] wl[229] vdd gnd cell_6t
Xbit_r230_c90 bl[90] br[90] wl[230] vdd gnd cell_6t
Xbit_r231_c90 bl[90] br[90] wl[231] vdd gnd cell_6t
Xbit_r232_c90 bl[90] br[90] wl[232] vdd gnd cell_6t
Xbit_r233_c90 bl[90] br[90] wl[233] vdd gnd cell_6t
Xbit_r234_c90 bl[90] br[90] wl[234] vdd gnd cell_6t
Xbit_r235_c90 bl[90] br[90] wl[235] vdd gnd cell_6t
Xbit_r236_c90 bl[90] br[90] wl[236] vdd gnd cell_6t
Xbit_r237_c90 bl[90] br[90] wl[237] vdd gnd cell_6t
Xbit_r238_c90 bl[90] br[90] wl[238] vdd gnd cell_6t
Xbit_r239_c90 bl[90] br[90] wl[239] vdd gnd cell_6t
Xbit_r240_c90 bl[90] br[90] wl[240] vdd gnd cell_6t
Xbit_r241_c90 bl[90] br[90] wl[241] vdd gnd cell_6t
Xbit_r242_c90 bl[90] br[90] wl[242] vdd gnd cell_6t
Xbit_r243_c90 bl[90] br[90] wl[243] vdd gnd cell_6t
Xbit_r244_c90 bl[90] br[90] wl[244] vdd gnd cell_6t
Xbit_r245_c90 bl[90] br[90] wl[245] vdd gnd cell_6t
Xbit_r246_c90 bl[90] br[90] wl[246] vdd gnd cell_6t
Xbit_r247_c90 bl[90] br[90] wl[247] vdd gnd cell_6t
Xbit_r248_c90 bl[90] br[90] wl[248] vdd gnd cell_6t
Xbit_r249_c90 bl[90] br[90] wl[249] vdd gnd cell_6t
Xbit_r250_c90 bl[90] br[90] wl[250] vdd gnd cell_6t
Xbit_r251_c90 bl[90] br[90] wl[251] vdd gnd cell_6t
Xbit_r252_c90 bl[90] br[90] wl[252] vdd gnd cell_6t
Xbit_r253_c90 bl[90] br[90] wl[253] vdd gnd cell_6t
Xbit_r254_c90 bl[90] br[90] wl[254] vdd gnd cell_6t
Xbit_r255_c90 bl[90] br[90] wl[255] vdd gnd cell_6t
Xbit_r256_c90 bl[90] br[90] wl[256] vdd gnd cell_6t
Xbit_r257_c90 bl[90] br[90] wl[257] vdd gnd cell_6t
Xbit_r258_c90 bl[90] br[90] wl[258] vdd gnd cell_6t
Xbit_r259_c90 bl[90] br[90] wl[259] vdd gnd cell_6t
Xbit_r260_c90 bl[90] br[90] wl[260] vdd gnd cell_6t
Xbit_r261_c90 bl[90] br[90] wl[261] vdd gnd cell_6t
Xbit_r262_c90 bl[90] br[90] wl[262] vdd gnd cell_6t
Xbit_r263_c90 bl[90] br[90] wl[263] vdd gnd cell_6t
Xbit_r264_c90 bl[90] br[90] wl[264] vdd gnd cell_6t
Xbit_r265_c90 bl[90] br[90] wl[265] vdd gnd cell_6t
Xbit_r266_c90 bl[90] br[90] wl[266] vdd gnd cell_6t
Xbit_r267_c90 bl[90] br[90] wl[267] vdd gnd cell_6t
Xbit_r268_c90 bl[90] br[90] wl[268] vdd gnd cell_6t
Xbit_r269_c90 bl[90] br[90] wl[269] vdd gnd cell_6t
Xbit_r270_c90 bl[90] br[90] wl[270] vdd gnd cell_6t
Xbit_r271_c90 bl[90] br[90] wl[271] vdd gnd cell_6t
Xbit_r272_c90 bl[90] br[90] wl[272] vdd gnd cell_6t
Xbit_r273_c90 bl[90] br[90] wl[273] vdd gnd cell_6t
Xbit_r274_c90 bl[90] br[90] wl[274] vdd gnd cell_6t
Xbit_r275_c90 bl[90] br[90] wl[275] vdd gnd cell_6t
Xbit_r276_c90 bl[90] br[90] wl[276] vdd gnd cell_6t
Xbit_r277_c90 bl[90] br[90] wl[277] vdd gnd cell_6t
Xbit_r278_c90 bl[90] br[90] wl[278] vdd gnd cell_6t
Xbit_r279_c90 bl[90] br[90] wl[279] vdd gnd cell_6t
Xbit_r280_c90 bl[90] br[90] wl[280] vdd gnd cell_6t
Xbit_r281_c90 bl[90] br[90] wl[281] vdd gnd cell_6t
Xbit_r282_c90 bl[90] br[90] wl[282] vdd gnd cell_6t
Xbit_r283_c90 bl[90] br[90] wl[283] vdd gnd cell_6t
Xbit_r284_c90 bl[90] br[90] wl[284] vdd gnd cell_6t
Xbit_r285_c90 bl[90] br[90] wl[285] vdd gnd cell_6t
Xbit_r286_c90 bl[90] br[90] wl[286] vdd gnd cell_6t
Xbit_r287_c90 bl[90] br[90] wl[287] vdd gnd cell_6t
Xbit_r288_c90 bl[90] br[90] wl[288] vdd gnd cell_6t
Xbit_r289_c90 bl[90] br[90] wl[289] vdd gnd cell_6t
Xbit_r290_c90 bl[90] br[90] wl[290] vdd gnd cell_6t
Xbit_r291_c90 bl[90] br[90] wl[291] vdd gnd cell_6t
Xbit_r292_c90 bl[90] br[90] wl[292] vdd gnd cell_6t
Xbit_r293_c90 bl[90] br[90] wl[293] vdd gnd cell_6t
Xbit_r294_c90 bl[90] br[90] wl[294] vdd gnd cell_6t
Xbit_r295_c90 bl[90] br[90] wl[295] vdd gnd cell_6t
Xbit_r296_c90 bl[90] br[90] wl[296] vdd gnd cell_6t
Xbit_r297_c90 bl[90] br[90] wl[297] vdd gnd cell_6t
Xbit_r298_c90 bl[90] br[90] wl[298] vdd gnd cell_6t
Xbit_r299_c90 bl[90] br[90] wl[299] vdd gnd cell_6t
Xbit_r300_c90 bl[90] br[90] wl[300] vdd gnd cell_6t
Xbit_r301_c90 bl[90] br[90] wl[301] vdd gnd cell_6t
Xbit_r302_c90 bl[90] br[90] wl[302] vdd gnd cell_6t
Xbit_r303_c90 bl[90] br[90] wl[303] vdd gnd cell_6t
Xbit_r304_c90 bl[90] br[90] wl[304] vdd gnd cell_6t
Xbit_r305_c90 bl[90] br[90] wl[305] vdd gnd cell_6t
Xbit_r306_c90 bl[90] br[90] wl[306] vdd gnd cell_6t
Xbit_r307_c90 bl[90] br[90] wl[307] vdd gnd cell_6t
Xbit_r308_c90 bl[90] br[90] wl[308] vdd gnd cell_6t
Xbit_r309_c90 bl[90] br[90] wl[309] vdd gnd cell_6t
Xbit_r310_c90 bl[90] br[90] wl[310] vdd gnd cell_6t
Xbit_r311_c90 bl[90] br[90] wl[311] vdd gnd cell_6t
Xbit_r312_c90 bl[90] br[90] wl[312] vdd gnd cell_6t
Xbit_r313_c90 bl[90] br[90] wl[313] vdd gnd cell_6t
Xbit_r314_c90 bl[90] br[90] wl[314] vdd gnd cell_6t
Xbit_r315_c90 bl[90] br[90] wl[315] vdd gnd cell_6t
Xbit_r316_c90 bl[90] br[90] wl[316] vdd gnd cell_6t
Xbit_r317_c90 bl[90] br[90] wl[317] vdd gnd cell_6t
Xbit_r318_c90 bl[90] br[90] wl[318] vdd gnd cell_6t
Xbit_r319_c90 bl[90] br[90] wl[319] vdd gnd cell_6t
Xbit_r320_c90 bl[90] br[90] wl[320] vdd gnd cell_6t
Xbit_r321_c90 bl[90] br[90] wl[321] vdd gnd cell_6t
Xbit_r322_c90 bl[90] br[90] wl[322] vdd gnd cell_6t
Xbit_r323_c90 bl[90] br[90] wl[323] vdd gnd cell_6t
Xbit_r324_c90 bl[90] br[90] wl[324] vdd gnd cell_6t
Xbit_r325_c90 bl[90] br[90] wl[325] vdd gnd cell_6t
Xbit_r326_c90 bl[90] br[90] wl[326] vdd gnd cell_6t
Xbit_r327_c90 bl[90] br[90] wl[327] vdd gnd cell_6t
Xbit_r328_c90 bl[90] br[90] wl[328] vdd gnd cell_6t
Xbit_r329_c90 bl[90] br[90] wl[329] vdd gnd cell_6t
Xbit_r330_c90 bl[90] br[90] wl[330] vdd gnd cell_6t
Xbit_r331_c90 bl[90] br[90] wl[331] vdd gnd cell_6t
Xbit_r332_c90 bl[90] br[90] wl[332] vdd gnd cell_6t
Xbit_r333_c90 bl[90] br[90] wl[333] vdd gnd cell_6t
Xbit_r334_c90 bl[90] br[90] wl[334] vdd gnd cell_6t
Xbit_r335_c90 bl[90] br[90] wl[335] vdd gnd cell_6t
Xbit_r336_c90 bl[90] br[90] wl[336] vdd gnd cell_6t
Xbit_r337_c90 bl[90] br[90] wl[337] vdd gnd cell_6t
Xbit_r338_c90 bl[90] br[90] wl[338] vdd gnd cell_6t
Xbit_r339_c90 bl[90] br[90] wl[339] vdd gnd cell_6t
Xbit_r340_c90 bl[90] br[90] wl[340] vdd gnd cell_6t
Xbit_r341_c90 bl[90] br[90] wl[341] vdd gnd cell_6t
Xbit_r342_c90 bl[90] br[90] wl[342] vdd gnd cell_6t
Xbit_r343_c90 bl[90] br[90] wl[343] vdd gnd cell_6t
Xbit_r344_c90 bl[90] br[90] wl[344] vdd gnd cell_6t
Xbit_r345_c90 bl[90] br[90] wl[345] vdd gnd cell_6t
Xbit_r346_c90 bl[90] br[90] wl[346] vdd gnd cell_6t
Xbit_r347_c90 bl[90] br[90] wl[347] vdd gnd cell_6t
Xbit_r348_c90 bl[90] br[90] wl[348] vdd gnd cell_6t
Xbit_r349_c90 bl[90] br[90] wl[349] vdd gnd cell_6t
Xbit_r350_c90 bl[90] br[90] wl[350] vdd gnd cell_6t
Xbit_r351_c90 bl[90] br[90] wl[351] vdd gnd cell_6t
Xbit_r352_c90 bl[90] br[90] wl[352] vdd gnd cell_6t
Xbit_r353_c90 bl[90] br[90] wl[353] vdd gnd cell_6t
Xbit_r354_c90 bl[90] br[90] wl[354] vdd gnd cell_6t
Xbit_r355_c90 bl[90] br[90] wl[355] vdd gnd cell_6t
Xbit_r356_c90 bl[90] br[90] wl[356] vdd gnd cell_6t
Xbit_r357_c90 bl[90] br[90] wl[357] vdd gnd cell_6t
Xbit_r358_c90 bl[90] br[90] wl[358] vdd gnd cell_6t
Xbit_r359_c90 bl[90] br[90] wl[359] vdd gnd cell_6t
Xbit_r360_c90 bl[90] br[90] wl[360] vdd gnd cell_6t
Xbit_r361_c90 bl[90] br[90] wl[361] vdd gnd cell_6t
Xbit_r362_c90 bl[90] br[90] wl[362] vdd gnd cell_6t
Xbit_r363_c90 bl[90] br[90] wl[363] vdd gnd cell_6t
Xbit_r364_c90 bl[90] br[90] wl[364] vdd gnd cell_6t
Xbit_r365_c90 bl[90] br[90] wl[365] vdd gnd cell_6t
Xbit_r366_c90 bl[90] br[90] wl[366] vdd gnd cell_6t
Xbit_r367_c90 bl[90] br[90] wl[367] vdd gnd cell_6t
Xbit_r368_c90 bl[90] br[90] wl[368] vdd gnd cell_6t
Xbit_r369_c90 bl[90] br[90] wl[369] vdd gnd cell_6t
Xbit_r370_c90 bl[90] br[90] wl[370] vdd gnd cell_6t
Xbit_r371_c90 bl[90] br[90] wl[371] vdd gnd cell_6t
Xbit_r372_c90 bl[90] br[90] wl[372] vdd gnd cell_6t
Xbit_r373_c90 bl[90] br[90] wl[373] vdd gnd cell_6t
Xbit_r374_c90 bl[90] br[90] wl[374] vdd gnd cell_6t
Xbit_r375_c90 bl[90] br[90] wl[375] vdd gnd cell_6t
Xbit_r376_c90 bl[90] br[90] wl[376] vdd gnd cell_6t
Xbit_r377_c90 bl[90] br[90] wl[377] vdd gnd cell_6t
Xbit_r378_c90 bl[90] br[90] wl[378] vdd gnd cell_6t
Xbit_r379_c90 bl[90] br[90] wl[379] vdd gnd cell_6t
Xbit_r380_c90 bl[90] br[90] wl[380] vdd gnd cell_6t
Xbit_r381_c90 bl[90] br[90] wl[381] vdd gnd cell_6t
Xbit_r382_c90 bl[90] br[90] wl[382] vdd gnd cell_6t
Xbit_r383_c90 bl[90] br[90] wl[383] vdd gnd cell_6t
Xbit_r384_c90 bl[90] br[90] wl[384] vdd gnd cell_6t
Xbit_r385_c90 bl[90] br[90] wl[385] vdd gnd cell_6t
Xbit_r386_c90 bl[90] br[90] wl[386] vdd gnd cell_6t
Xbit_r387_c90 bl[90] br[90] wl[387] vdd gnd cell_6t
Xbit_r388_c90 bl[90] br[90] wl[388] vdd gnd cell_6t
Xbit_r389_c90 bl[90] br[90] wl[389] vdd gnd cell_6t
Xbit_r390_c90 bl[90] br[90] wl[390] vdd gnd cell_6t
Xbit_r391_c90 bl[90] br[90] wl[391] vdd gnd cell_6t
Xbit_r392_c90 bl[90] br[90] wl[392] vdd gnd cell_6t
Xbit_r393_c90 bl[90] br[90] wl[393] vdd gnd cell_6t
Xbit_r394_c90 bl[90] br[90] wl[394] vdd gnd cell_6t
Xbit_r395_c90 bl[90] br[90] wl[395] vdd gnd cell_6t
Xbit_r396_c90 bl[90] br[90] wl[396] vdd gnd cell_6t
Xbit_r397_c90 bl[90] br[90] wl[397] vdd gnd cell_6t
Xbit_r398_c90 bl[90] br[90] wl[398] vdd gnd cell_6t
Xbit_r399_c90 bl[90] br[90] wl[399] vdd gnd cell_6t
Xbit_r400_c90 bl[90] br[90] wl[400] vdd gnd cell_6t
Xbit_r401_c90 bl[90] br[90] wl[401] vdd gnd cell_6t
Xbit_r402_c90 bl[90] br[90] wl[402] vdd gnd cell_6t
Xbit_r403_c90 bl[90] br[90] wl[403] vdd gnd cell_6t
Xbit_r404_c90 bl[90] br[90] wl[404] vdd gnd cell_6t
Xbit_r405_c90 bl[90] br[90] wl[405] vdd gnd cell_6t
Xbit_r406_c90 bl[90] br[90] wl[406] vdd gnd cell_6t
Xbit_r407_c90 bl[90] br[90] wl[407] vdd gnd cell_6t
Xbit_r408_c90 bl[90] br[90] wl[408] vdd gnd cell_6t
Xbit_r409_c90 bl[90] br[90] wl[409] vdd gnd cell_6t
Xbit_r410_c90 bl[90] br[90] wl[410] vdd gnd cell_6t
Xbit_r411_c90 bl[90] br[90] wl[411] vdd gnd cell_6t
Xbit_r412_c90 bl[90] br[90] wl[412] vdd gnd cell_6t
Xbit_r413_c90 bl[90] br[90] wl[413] vdd gnd cell_6t
Xbit_r414_c90 bl[90] br[90] wl[414] vdd gnd cell_6t
Xbit_r415_c90 bl[90] br[90] wl[415] vdd gnd cell_6t
Xbit_r416_c90 bl[90] br[90] wl[416] vdd gnd cell_6t
Xbit_r417_c90 bl[90] br[90] wl[417] vdd gnd cell_6t
Xbit_r418_c90 bl[90] br[90] wl[418] vdd gnd cell_6t
Xbit_r419_c90 bl[90] br[90] wl[419] vdd gnd cell_6t
Xbit_r420_c90 bl[90] br[90] wl[420] vdd gnd cell_6t
Xbit_r421_c90 bl[90] br[90] wl[421] vdd gnd cell_6t
Xbit_r422_c90 bl[90] br[90] wl[422] vdd gnd cell_6t
Xbit_r423_c90 bl[90] br[90] wl[423] vdd gnd cell_6t
Xbit_r424_c90 bl[90] br[90] wl[424] vdd gnd cell_6t
Xbit_r425_c90 bl[90] br[90] wl[425] vdd gnd cell_6t
Xbit_r426_c90 bl[90] br[90] wl[426] vdd gnd cell_6t
Xbit_r427_c90 bl[90] br[90] wl[427] vdd gnd cell_6t
Xbit_r428_c90 bl[90] br[90] wl[428] vdd gnd cell_6t
Xbit_r429_c90 bl[90] br[90] wl[429] vdd gnd cell_6t
Xbit_r430_c90 bl[90] br[90] wl[430] vdd gnd cell_6t
Xbit_r431_c90 bl[90] br[90] wl[431] vdd gnd cell_6t
Xbit_r432_c90 bl[90] br[90] wl[432] vdd gnd cell_6t
Xbit_r433_c90 bl[90] br[90] wl[433] vdd gnd cell_6t
Xbit_r434_c90 bl[90] br[90] wl[434] vdd gnd cell_6t
Xbit_r435_c90 bl[90] br[90] wl[435] vdd gnd cell_6t
Xbit_r436_c90 bl[90] br[90] wl[436] vdd gnd cell_6t
Xbit_r437_c90 bl[90] br[90] wl[437] vdd gnd cell_6t
Xbit_r438_c90 bl[90] br[90] wl[438] vdd gnd cell_6t
Xbit_r439_c90 bl[90] br[90] wl[439] vdd gnd cell_6t
Xbit_r440_c90 bl[90] br[90] wl[440] vdd gnd cell_6t
Xbit_r441_c90 bl[90] br[90] wl[441] vdd gnd cell_6t
Xbit_r442_c90 bl[90] br[90] wl[442] vdd gnd cell_6t
Xbit_r443_c90 bl[90] br[90] wl[443] vdd gnd cell_6t
Xbit_r444_c90 bl[90] br[90] wl[444] vdd gnd cell_6t
Xbit_r445_c90 bl[90] br[90] wl[445] vdd gnd cell_6t
Xbit_r446_c90 bl[90] br[90] wl[446] vdd gnd cell_6t
Xbit_r447_c90 bl[90] br[90] wl[447] vdd gnd cell_6t
Xbit_r448_c90 bl[90] br[90] wl[448] vdd gnd cell_6t
Xbit_r449_c90 bl[90] br[90] wl[449] vdd gnd cell_6t
Xbit_r450_c90 bl[90] br[90] wl[450] vdd gnd cell_6t
Xbit_r451_c90 bl[90] br[90] wl[451] vdd gnd cell_6t
Xbit_r452_c90 bl[90] br[90] wl[452] vdd gnd cell_6t
Xbit_r453_c90 bl[90] br[90] wl[453] vdd gnd cell_6t
Xbit_r454_c90 bl[90] br[90] wl[454] vdd gnd cell_6t
Xbit_r455_c90 bl[90] br[90] wl[455] vdd gnd cell_6t
Xbit_r456_c90 bl[90] br[90] wl[456] vdd gnd cell_6t
Xbit_r457_c90 bl[90] br[90] wl[457] vdd gnd cell_6t
Xbit_r458_c90 bl[90] br[90] wl[458] vdd gnd cell_6t
Xbit_r459_c90 bl[90] br[90] wl[459] vdd gnd cell_6t
Xbit_r460_c90 bl[90] br[90] wl[460] vdd gnd cell_6t
Xbit_r461_c90 bl[90] br[90] wl[461] vdd gnd cell_6t
Xbit_r462_c90 bl[90] br[90] wl[462] vdd gnd cell_6t
Xbit_r463_c90 bl[90] br[90] wl[463] vdd gnd cell_6t
Xbit_r464_c90 bl[90] br[90] wl[464] vdd gnd cell_6t
Xbit_r465_c90 bl[90] br[90] wl[465] vdd gnd cell_6t
Xbit_r466_c90 bl[90] br[90] wl[466] vdd gnd cell_6t
Xbit_r467_c90 bl[90] br[90] wl[467] vdd gnd cell_6t
Xbit_r468_c90 bl[90] br[90] wl[468] vdd gnd cell_6t
Xbit_r469_c90 bl[90] br[90] wl[469] vdd gnd cell_6t
Xbit_r470_c90 bl[90] br[90] wl[470] vdd gnd cell_6t
Xbit_r471_c90 bl[90] br[90] wl[471] vdd gnd cell_6t
Xbit_r472_c90 bl[90] br[90] wl[472] vdd gnd cell_6t
Xbit_r473_c90 bl[90] br[90] wl[473] vdd gnd cell_6t
Xbit_r474_c90 bl[90] br[90] wl[474] vdd gnd cell_6t
Xbit_r475_c90 bl[90] br[90] wl[475] vdd gnd cell_6t
Xbit_r476_c90 bl[90] br[90] wl[476] vdd gnd cell_6t
Xbit_r477_c90 bl[90] br[90] wl[477] vdd gnd cell_6t
Xbit_r478_c90 bl[90] br[90] wl[478] vdd gnd cell_6t
Xbit_r479_c90 bl[90] br[90] wl[479] vdd gnd cell_6t
Xbit_r480_c90 bl[90] br[90] wl[480] vdd gnd cell_6t
Xbit_r481_c90 bl[90] br[90] wl[481] vdd gnd cell_6t
Xbit_r482_c90 bl[90] br[90] wl[482] vdd gnd cell_6t
Xbit_r483_c90 bl[90] br[90] wl[483] vdd gnd cell_6t
Xbit_r484_c90 bl[90] br[90] wl[484] vdd gnd cell_6t
Xbit_r485_c90 bl[90] br[90] wl[485] vdd gnd cell_6t
Xbit_r486_c90 bl[90] br[90] wl[486] vdd gnd cell_6t
Xbit_r487_c90 bl[90] br[90] wl[487] vdd gnd cell_6t
Xbit_r488_c90 bl[90] br[90] wl[488] vdd gnd cell_6t
Xbit_r489_c90 bl[90] br[90] wl[489] vdd gnd cell_6t
Xbit_r490_c90 bl[90] br[90] wl[490] vdd gnd cell_6t
Xbit_r491_c90 bl[90] br[90] wl[491] vdd gnd cell_6t
Xbit_r492_c90 bl[90] br[90] wl[492] vdd gnd cell_6t
Xbit_r493_c90 bl[90] br[90] wl[493] vdd gnd cell_6t
Xbit_r494_c90 bl[90] br[90] wl[494] vdd gnd cell_6t
Xbit_r495_c90 bl[90] br[90] wl[495] vdd gnd cell_6t
Xbit_r496_c90 bl[90] br[90] wl[496] vdd gnd cell_6t
Xbit_r497_c90 bl[90] br[90] wl[497] vdd gnd cell_6t
Xbit_r498_c90 bl[90] br[90] wl[498] vdd gnd cell_6t
Xbit_r499_c90 bl[90] br[90] wl[499] vdd gnd cell_6t
Xbit_r500_c90 bl[90] br[90] wl[500] vdd gnd cell_6t
Xbit_r501_c90 bl[90] br[90] wl[501] vdd gnd cell_6t
Xbit_r502_c90 bl[90] br[90] wl[502] vdd gnd cell_6t
Xbit_r503_c90 bl[90] br[90] wl[503] vdd gnd cell_6t
Xbit_r504_c90 bl[90] br[90] wl[504] vdd gnd cell_6t
Xbit_r505_c90 bl[90] br[90] wl[505] vdd gnd cell_6t
Xbit_r506_c90 bl[90] br[90] wl[506] vdd gnd cell_6t
Xbit_r507_c90 bl[90] br[90] wl[507] vdd gnd cell_6t
Xbit_r508_c90 bl[90] br[90] wl[508] vdd gnd cell_6t
Xbit_r509_c90 bl[90] br[90] wl[509] vdd gnd cell_6t
Xbit_r510_c90 bl[90] br[90] wl[510] vdd gnd cell_6t
Xbit_r511_c90 bl[90] br[90] wl[511] vdd gnd cell_6t
Xbit_r0_c91 bl[91] br[91] wl[0] vdd gnd cell_6t
Xbit_r1_c91 bl[91] br[91] wl[1] vdd gnd cell_6t
Xbit_r2_c91 bl[91] br[91] wl[2] vdd gnd cell_6t
Xbit_r3_c91 bl[91] br[91] wl[3] vdd gnd cell_6t
Xbit_r4_c91 bl[91] br[91] wl[4] vdd gnd cell_6t
Xbit_r5_c91 bl[91] br[91] wl[5] vdd gnd cell_6t
Xbit_r6_c91 bl[91] br[91] wl[6] vdd gnd cell_6t
Xbit_r7_c91 bl[91] br[91] wl[7] vdd gnd cell_6t
Xbit_r8_c91 bl[91] br[91] wl[8] vdd gnd cell_6t
Xbit_r9_c91 bl[91] br[91] wl[9] vdd gnd cell_6t
Xbit_r10_c91 bl[91] br[91] wl[10] vdd gnd cell_6t
Xbit_r11_c91 bl[91] br[91] wl[11] vdd gnd cell_6t
Xbit_r12_c91 bl[91] br[91] wl[12] vdd gnd cell_6t
Xbit_r13_c91 bl[91] br[91] wl[13] vdd gnd cell_6t
Xbit_r14_c91 bl[91] br[91] wl[14] vdd gnd cell_6t
Xbit_r15_c91 bl[91] br[91] wl[15] vdd gnd cell_6t
Xbit_r16_c91 bl[91] br[91] wl[16] vdd gnd cell_6t
Xbit_r17_c91 bl[91] br[91] wl[17] vdd gnd cell_6t
Xbit_r18_c91 bl[91] br[91] wl[18] vdd gnd cell_6t
Xbit_r19_c91 bl[91] br[91] wl[19] vdd gnd cell_6t
Xbit_r20_c91 bl[91] br[91] wl[20] vdd gnd cell_6t
Xbit_r21_c91 bl[91] br[91] wl[21] vdd gnd cell_6t
Xbit_r22_c91 bl[91] br[91] wl[22] vdd gnd cell_6t
Xbit_r23_c91 bl[91] br[91] wl[23] vdd gnd cell_6t
Xbit_r24_c91 bl[91] br[91] wl[24] vdd gnd cell_6t
Xbit_r25_c91 bl[91] br[91] wl[25] vdd gnd cell_6t
Xbit_r26_c91 bl[91] br[91] wl[26] vdd gnd cell_6t
Xbit_r27_c91 bl[91] br[91] wl[27] vdd gnd cell_6t
Xbit_r28_c91 bl[91] br[91] wl[28] vdd gnd cell_6t
Xbit_r29_c91 bl[91] br[91] wl[29] vdd gnd cell_6t
Xbit_r30_c91 bl[91] br[91] wl[30] vdd gnd cell_6t
Xbit_r31_c91 bl[91] br[91] wl[31] vdd gnd cell_6t
Xbit_r32_c91 bl[91] br[91] wl[32] vdd gnd cell_6t
Xbit_r33_c91 bl[91] br[91] wl[33] vdd gnd cell_6t
Xbit_r34_c91 bl[91] br[91] wl[34] vdd gnd cell_6t
Xbit_r35_c91 bl[91] br[91] wl[35] vdd gnd cell_6t
Xbit_r36_c91 bl[91] br[91] wl[36] vdd gnd cell_6t
Xbit_r37_c91 bl[91] br[91] wl[37] vdd gnd cell_6t
Xbit_r38_c91 bl[91] br[91] wl[38] vdd gnd cell_6t
Xbit_r39_c91 bl[91] br[91] wl[39] vdd gnd cell_6t
Xbit_r40_c91 bl[91] br[91] wl[40] vdd gnd cell_6t
Xbit_r41_c91 bl[91] br[91] wl[41] vdd gnd cell_6t
Xbit_r42_c91 bl[91] br[91] wl[42] vdd gnd cell_6t
Xbit_r43_c91 bl[91] br[91] wl[43] vdd gnd cell_6t
Xbit_r44_c91 bl[91] br[91] wl[44] vdd gnd cell_6t
Xbit_r45_c91 bl[91] br[91] wl[45] vdd gnd cell_6t
Xbit_r46_c91 bl[91] br[91] wl[46] vdd gnd cell_6t
Xbit_r47_c91 bl[91] br[91] wl[47] vdd gnd cell_6t
Xbit_r48_c91 bl[91] br[91] wl[48] vdd gnd cell_6t
Xbit_r49_c91 bl[91] br[91] wl[49] vdd gnd cell_6t
Xbit_r50_c91 bl[91] br[91] wl[50] vdd gnd cell_6t
Xbit_r51_c91 bl[91] br[91] wl[51] vdd gnd cell_6t
Xbit_r52_c91 bl[91] br[91] wl[52] vdd gnd cell_6t
Xbit_r53_c91 bl[91] br[91] wl[53] vdd gnd cell_6t
Xbit_r54_c91 bl[91] br[91] wl[54] vdd gnd cell_6t
Xbit_r55_c91 bl[91] br[91] wl[55] vdd gnd cell_6t
Xbit_r56_c91 bl[91] br[91] wl[56] vdd gnd cell_6t
Xbit_r57_c91 bl[91] br[91] wl[57] vdd gnd cell_6t
Xbit_r58_c91 bl[91] br[91] wl[58] vdd gnd cell_6t
Xbit_r59_c91 bl[91] br[91] wl[59] vdd gnd cell_6t
Xbit_r60_c91 bl[91] br[91] wl[60] vdd gnd cell_6t
Xbit_r61_c91 bl[91] br[91] wl[61] vdd gnd cell_6t
Xbit_r62_c91 bl[91] br[91] wl[62] vdd gnd cell_6t
Xbit_r63_c91 bl[91] br[91] wl[63] vdd gnd cell_6t
Xbit_r64_c91 bl[91] br[91] wl[64] vdd gnd cell_6t
Xbit_r65_c91 bl[91] br[91] wl[65] vdd gnd cell_6t
Xbit_r66_c91 bl[91] br[91] wl[66] vdd gnd cell_6t
Xbit_r67_c91 bl[91] br[91] wl[67] vdd gnd cell_6t
Xbit_r68_c91 bl[91] br[91] wl[68] vdd gnd cell_6t
Xbit_r69_c91 bl[91] br[91] wl[69] vdd gnd cell_6t
Xbit_r70_c91 bl[91] br[91] wl[70] vdd gnd cell_6t
Xbit_r71_c91 bl[91] br[91] wl[71] vdd gnd cell_6t
Xbit_r72_c91 bl[91] br[91] wl[72] vdd gnd cell_6t
Xbit_r73_c91 bl[91] br[91] wl[73] vdd gnd cell_6t
Xbit_r74_c91 bl[91] br[91] wl[74] vdd gnd cell_6t
Xbit_r75_c91 bl[91] br[91] wl[75] vdd gnd cell_6t
Xbit_r76_c91 bl[91] br[91] wl[76] vdd gnd cell_6t
Xbit_r77_c91 bl[91] br[91] wl[77] vdd gnd cell_6t
Xbit_r78_c91 bl[91] br[91] wl[78] vdd gnd cell_6t
Xbit_r79_c91 bl[91] br[91] wl[79] vdd gnd cell_6t
Xbit_r80_c91 bl[91] br[91] wl[80] vdd gnd cell_6t
Xbit_r81_c91 bl[91] br[91] wl[81] vdd gnd cell_6t
Xbit_r82_c91 bl[91] br[91] wl[82] vdd gnd cell_6t
Xbit_r83_c91 bl[91] br[91] wl[83] vdd gnd cell_6t
Xbit_r84_c91 bl[91] br[91] wl[84] vdd gnd cell_6t
Xbit_r85_c91 bl[91] br[91] wl[85] vdd gnd cell_6t
Xbit_r86_c91 bl[91] br[91] wl[86] vdd gnd cell_6t
Xbit_r87_c91 bl[91] br[91] wl[87] vdd gnd cell_6t
Xbit_r88_c91 bl[91] br[91] wl[88] vdd gnd cell_6t
Xbit_r89_c91 bl[91] br[91] wl[89] vdd gnd cell_6t
Xbit_r90_c91 bl[91] br[91] wl[90] vdd gnd cell_6t
Xbit_r91_c91 bl[91] br[91] wl[91] vdd gnd cell_6t
Xbit_r92_c91 bl[91] br[91] wl[92] vdd gnd cell_6t
Xbit_r93_c91 bl[91] br[91] wl[93] vdd gnd cell_6t
Xbit_r94_c91 bl[91] br[91] wl[94] vdd gnd cell_6t
Xbit_r95_c91 bl[91] br[91] wl[95] vdd gnd cell_6t
Xbit_r96_c91 bl[91] br[91] wl[96] vdd gnd cell_6t
Xbit_r97_c91 bl[91] br[91] wl[97] vdd gnd cell_6t
Xbit_r98_c91 bl[91] br[91] wl[98] vdd gnd cell_6t
Xbit_r99_c91 bl[91] br[91] wl[99] vdd gnd cell_6t
Xbit_r100_c91 bl[91] br[91] wl[100] vdd gnd cell_6t
Xbit_r101_c91 bl[91] br[91] wl[101] vdd gnd cell_6t
Xbit_r102_c91 bl[91] br[91] wl[102] vdd gnd cell_6t
Xbit_r103_c91 bl[91] br[91] wl[103] vdd gnd cell_6t
Xbit_r104_c91 bl[91] br[91] wl[104] vdd gnd cell_6t
Xbit_r105_c91 bl[91] br[91] wl[105] vdd gnd cell_6t
Xbit_r106_c91 bl[91] br[91] wl[106] vdd gnd cell_6t
Xbit_r107_c91 bl[91] br[91] wl[107] vdd gnd cell_6t
Xbit_r108_c91 bl[91] br[91] wl[108] vdd gnd cell_6t
Xbit_r109_c91 bl[91] br[91] wl[109] vdd gnd cell_6t
Xbit_r110_c91 bl[91] br[91] wl[110] vdd gnd cell_6t
Xbit_r111_c91 bl[91] br[91] wl[111] vdd gnd cell_6t
Xbit_r112_c91 bl[91] br[91] wl[112] vdd gnd cell_6t
Xbit_r113_c91 bl[91] br[91] wl[113] vdd gnd cell_6t
Xbit_r114_c91 bl[91] br[91] wl[114] vdd gnd cell_6t
Xbit_r115_c91 bl[91] br[91] wl[115] vdd gnd cell_6t
Xbit_r116_c91 bl[91] br[91] wl[116] vdd gnd cell_6t
Xbit_r117_c91 bl[91] br[91] wl[117] vdd gnd cell_6t
Xbit_r118_c91 bl[91] br[91] wl[118] vdd gnd cell_6t
Xbit_r119_c91 bl[91] br[91] wl[119] vdd gnd cell_6t
Xbit_r120_c91 bl[91] br[91] wl[120] vdd gnd cell_6t
Xbit_r121_c91 bl[91] br[91] wl[121] vdd gnd cell_6t
Xbit_r122_c91 bl[91] br[91] wl[122] vdd gnd cell_6t
Xbit_r123_c91 bl[91] br[91] wl[123] vdd gnd cell_6t
Xbit_r124_c91 bl[91] br[91] wl[124] vdd gnd cell_6t
Xbit_r125_c91 bl[91] br[91] wl[125] vdd gnd cell_6t
Xbit_r126_c91 bl[91] br[91] wl[126] vdd gnd cell_6t
Xbit_r127_c91 bl[91] br[91] wl[127] vdd gnd cell_6t
Xbit_r128_c91 bl[91] br[91] wl[128] vdd gnd cell_6t
Xbit_r129_c91 bl[91] br[91] wl[129] vdd gnd cell_6t
Xbit_r130_c91 bl[91] br[91] wl[130] vdd gnd cell_6t
Xbit_r131_c91 bl[91] br[91] wl[131] vdd gnd cell_6t
Xbit_r132_c91 bl[91] br[91] wl[132] vdd gnd cell_6t
Xbit_r133_c91 bl[91] br[91] wl[133] vdd gnd cell_6t
Xbit_r134_c91 bl[91] br[91] wl[134] vdd gnd cell_6t
Xbit_r135_c91 bl[91] br[91] wl[135] vdd gnd cell_6t
Xbit_r136_c91 bl[91] br[91] wl[136] vdd gnd cell_6t
Xbit_r137_c91 bl[91] br[91] wl[137] vdd gnd cell_6t
Xbit_r138_c91 bl[91] br[91] wl[138] vdd gnd cell_6t
Xbit_r139_c91 bl[91] br[91] wl[139] vdd gnd cell_6t
Xbit_r140_c91 bl[91] br[91] wl[140] vdd gnd cell_6t
Xbit_r141_c91 bl[91] br[91] wl[141] vdd gnd cell_6t
Xbit_r142_c91 bl[91] br[91] wl[142] vdd gnd cell_6t
Xbit_r143_c91 bl[91] br[91] wl[143] vdd gnd cell_6t
Xbit_r144_c91 bl[91] br[91] wl[144] vdd gnd cell_6t
Xbit_r145_c91 bl[91] br[91] wl[145] vdd gnd cell_6t
Xbit_r146_c91 bl[91] br[91] wl[146] vdd gnd cell_6t
Xbit_r147_c91 bl[91] br[91] wl[147] vdd gnd cell_6t
Xbit_r148_c91 bl[91] br[91] wl[148] vdd gnd cell_6t
Xbit_r149_c91 bl[91] br[91] wl[149] vdd gnd cell_6t
Xbit_r150_c91 bl[91] br[91] wl[150] vdd gnd cell_6t
Xbit_r151_c91 bl[91] br[91] wl[151] vdd gnd cell_6t
Xbit_r152_c91 bl[91] br[91] wl[152] vdd gnd cell_6t
Xbit_r153_c91 bl[91] br[91] wl[153] vdd gnd cell_6t
Xbit_r154_c91 bl[91] br[91] wl[154] vdd gnd cell_6t
Xbit_r155_c91 bl[91] br[91] wl[155] vdd gnd cell_6t
Xbit_r156_c91 bl[91] br[91] wl[156] vdd gnd cell_6t
Xbit_r157_c91 bl[91] br[91] wl[157] vdd gnd cell_6t
Xbit_r158_c91 bl[91] br[91] wl[158] vdd gnd cell_6t
Xbit_r159_c91 bl[91] br[91] wl[159] vdd gnd cell_6t
Xbit_r160_c91 bl[91] br[91] wl[160] vdd gnd cell_6t
Xbit_r161_c91 bl[91] br[91] wl[161] vdd gnd cell_6t
Xbit_r162_c91 bl[91] br[91] wl[162] vdd gnd cell_6t
Xbit_r163_c91 bl[91] br[91] wl[163] vdd gnd cell_6t
Xbit_r164_c91 bl[91] br[91] wl[164] vdd gnd cell_6t
Xbit_r165_c91 bl[91] br[91] wl[165] vdd gnd cell_6t
Xbit_r166_c91 bl[91] br[91] wl[166] vdd gnd cell_6t
Xbit_r167_c91 bl[91] br[91] wl[167] vdd gnd cell_6t
Xbit_r168_c91 bl[91] br[91] wl[168] vdd gnd cell_6t
Xbit_r169_c91 bl[91] br[91] wl[169] vdd gnd cell_6t
Xbit_r170_c91 bl[91] br[91] wl[170] vdd gnd cell_6t
Xbit_r171_c91 bl[91] br[91] wl[171] vdd gnd cell_6t
Xbit_r172_c91 bl[91] br[91] wl[172] vdd gnd cell_6t
Xbit_r173_c91 bl[91] br[91] wl[173] vdd gnd cell_6t
Xbit_r174_c91 bl[91] br[91] wl[174] vdd gnd cell_6t
Xbit_r175_c91 bl[91] br[91] wl[175] vdd gnd cell_6t
Xbit_r176_c91 bl[91] br[91] wl[176] vdd gnd cell_6t
Xbit_r177_c91 bl[91] br[91] wl[177] vdd gnd cell_6t
Xbit_r178_c91 bl[91] br[91] wl[178] vdd gnd cell_6t
Xbit_r179_c91 bl[91] br[91] wl[179] vdd gnd cell_6t
Xbit_r180_c91 bl[91] br[91] wl[180] vdd gnd cell_6t
Xbit_r181_c91 bl[91] br[91] wl[181] vdd gnd cell_6t
Xbit_r182_c91 bl[91] br[91] wl[182] vdd gnd cell_6t
Xbit_r183_c91 bl[91] br[91] wl[183] vdd gnd cell_6t
Xbit_r184_c91 bl[91] br[91] wl[184] vdd gnd cell_6t
Xbit_r185_c91 bl[91] br[91] wl[185] vdd gnd cell_6t
Xbit_r186_c91 bl[91] br[91] wl[186] vdd gnd cell_6t
Xbit_r187_c91 bl[91] br[91] wl[187] vdd gnd cell_6t
Xbit_r188_c91 bl[91] br[91] wl[188] vdd gnd cell_6t
Xbit_r189_c91 bl[91] br[91] wl[189] vdd gnd cell_6t
Xbit_r190_c91 bl[91] br[91] wl[190] vdd gnd cell_6t
Xbit_r191_c91 bl[91] br[91] wl[191] vdd gnd cell_6t
Xbit_r192_c91 bl[91] br[91] wl[192] vdd gnd cell_6t
Xbit_r193_c91 bl[91] br[91] wl[193] vdd gnd cell_6t
Xbit_r194_c91 bl[91] br[91] wl[194] vdd gnd cell_6t
Xbit_r195_c91 bl[91] br[91] wl[195] vdd gnd cell_6t
Xbit_r196_c91 bl[91] br[91] wl[196] vdd gnd cell_6t
Xbit_r197_c91 bl[91] br[91] wl[197] vdd gnd cell_6t
Xbit_r198_c91 bl[91] br[91] wl[198] vdd gnd cell_6t
Xbit_r199_c91 bl[91] br[91] wl[199] vdd gnd cell_6t
Xbit_r200_c91 bl[91] br[91] wl[200] vdd gnd cell_6t
Xbit_r201_c91 bl[91] br[91] wl[201] vdd gnd cell_6t
Xbit_r202_c91 bl[91] br[91] wl[202] vdd gnd cell_6t
Xbit_r203_c91 bl[91] br[91] wl[203] vdd gnd cell_6t
Xbit_r204_c91 bl[91] br[91] wl[204] vdd gnd cell_6t
Xbit_r205_c91 bl[91] br[91] wl[205] vdd gnd cell_6t
Xbit_r206_c91 bl[91] br[91] wl[206] vdd gnd cell_6t
Xbit_r207_c91 bl[91] br[91] wl[207] vdd gnd cell_6t
Xbit_r208_c91 bl[91] br[91] wl[208] vdd gnd cell_6t
Xbit_r209_c91 bl[91] br[91] wl[209] vdd gnd cell_6t
Xbit_r210_c91 bl[91] br[91] wl[210] vdd gnd cell_6t
Xbit_r211_c91 bl[91] br[91] wl[211] vdd gnd cell_6t
Xbit_r212_c91 bl[91] br[91] wl[212] vdd gnd cell_6t
Xbit_r213_c91 bl[91] br[91] wl[213] vdd gnd cell_6t
Xbit_r214_c91 bl[91] br[91] wl[214] vdd gnd cell_6t
Xbit_r215_c91 bl[91] br[91] wl[215] vdd gnd cell_6t
Xbit_r216_c91 bl[91] br[91] wl[216] vdd gnd cell_6t
Xbit_r217_c91 bl[91] br[91] wl[217] vdd gnd cell_6t
Xbit_r218_c91 bl[91] br[91] wl[218] vdd gnd cell_6t
Xbit_r219_c91 bl[91] br[91] wl[219] vdd gnd cell_6t
Xbit_r220_c91 bl[91] br[91] wl[220] vdd gnd cell_6t
Xbit_r221_c91 bl[91] br[91] wl[221] vdd gnd cell_6t
Xbit_r222_c91 bl[91] br[91] wl[222] vdd gnd cell_6t
Xbit_r223_c91 bl[91] br[91] wl[223] vdd gnd cell_6t
Xbit_r224_c91 bl[91] br[91] wl[224] vdd gnd cell_6t
Xbit_r225_c91 bl[91] br[91] wl[225] vdd gnd cell_6t
Xbit_r226_c91 bl[91] br[91] wl[226] vdd gnd cell_6t
Xbit_r227_c91 bl[91] br[91] wl[227] vdd gnd cell_6t
Xbit_r228_c91 bl[91] br[91] wl[228] vdd gnd cell_6t
Xbit_r229_c91 bl[91] br[91] wl[229] vdd gnd cell_6t
Xbit_r230_c91 bl[91] br[91] wl[230] vdd gnd cell_6t
Xbit_r231_c91 bl[91] br[91] wl[231] vdd gnd cell_6t
Xbit_r232_c91 bl[91] br[91] wl[232] vdd gnd cell_6t
Xbit_r233_c91 bl[91] br[91] wl[233] vdd gnd cell_6t
Xbit_r234_c91 bl[91] br[91] wl[234] vdd gnd cell_6t
Xbit_r235_c91 bl[91] br[91] wl[235] vdd gnd cell_6t
Xbit_r236_c91 bl[91] br[91] wl[236] vdd gnd cell_6t
Xbit_r237_c91 bl[91] br[91] wl[237] vdd gnd cell_6t
Xbit_r238_c91 bl[91] br[91] wl[238] vdd gnd cell_6t
Xbit_r239_c91 bl[91] br[91] wl[239] vdd gnd cell_6t
Xbit_r240_c91 bl[91] br[91] wl[240] vdd gnd cell_6t
Xbit_r241_c91 bl[91] br[91] wl[241] vdd gnd cell_6t
Xbit_r242_c91 bl[91] br[91] wl[242] vdd gnd cell_6t
Xbit_r243_c91 bl[91] br[91] wl[243] vdd gnd cell_6t
Xbit_r244_c91 bl[91] br[91] wl[244] vdd gnd cell_6t
Xbit_r245_c91 bl[91] br[91] wl[245] vdd gnd cell_6t
Xbit_r246_c91 bl[91] br[91] wl[246] vdd gnd cell_6t
Xbit_r247_c91 bl[91] br[91] wl[247] vdd gnd cell_6t
Xbit_r248_c91 bl[91] br[91] wl[248] vdd gnd cell_6t
Xbit_r249_c91 bl[91] br[91] wl[249] vdd gnd cell_6t
Xbit_r250_c91 bl[91] br[91] wl[250] vdd gnd cell_6t
Xbit_r251_c91 bl[91] br[91] wl[251] vdd gnd cell_6t
Xbit_r252_c91 bl[91] br[91] wl[252] vdd gnd cell_6t
Xbit_r253_c91 bl[91] br[91] wl[253] vdd gnd cell_6t
Xbit_r254_c91 bl[91] br[91] wl[254] vdd gnd cell_6t
Xbit_r255_c91 bl[91] br[91] wl[255] vdd gnd cell_6t
Xbit_r256_c91 bl[91] br[91] wl[256] vdd gnd cell_6t
Xbit_r257_c91 bl[91] br[91] wl[257] vdd gnd cell_6t
Xbit_r258_c91 bl[91] br[91] wl[258] vdd gnd cell_6t
Xbit_r259_c91 bl[91] br[91] wl[259] vdd gnd cell_6t
Xbit_r260_c91 bl[91] br[91] wl[260] vdd gnd cell_6t
Xbit_r261_c91 bl[91] br[91] wl[261] vdd gnd cell_6t
Xbit_r262_c91 bl[91] br[91] wl[262] vdd gnd cell_6t
Xbit_r263_c91 bl[91] br[91] wl[263] vdd gnd cell_6t
Xbit_r264_c91 bl[91] br[91] wl[264] vdd gnd cell_6t
Xbit_r265_c91 bl[91] br[91] wl[265] vdd gnd cell_6t
Xbit_r266_c91 bl[91] br[91] wl[266] vdd gnd cell_6t
Xbit_r267_c91 bl[91] br[91] wl[267] vdd gnd cell_6t
Xbit_r268_c91 bl[91] br[91] wl[268] vdd gnd cell_6t
Xbit_r269_c91 bl[91] br[91] wl[269] vdd gnd cell_6t
Xbit_r270_c91 bl[91] br[91] wl[270] vdd gnd cell_6t
Xbit_r271_c91 bl[91] br[91] wl[271] vdd gnd cell_6t
Xbit_r272_c91 bl[91] br[91] wl[272] vdd gnd cell_6t
Xbit_r273_c91 bl[91] br[91] wl[273] vdd gnd cell_6t
Xbit_r274_c91 bl[91] br[91] wl[274] vdd gnd cell_6t
Xbit_r275_c91 bl[91] br[91] wl[275] vdd gnd cell_6t
Xbit_r276_c91 bl[91] br[91] wl[276] vdd gnd cell_6t
Xbit_r277_c91 bl[91] br[91] wl[277] vdd gnd cell_6t
Xbit_r278_c91 bl[91] br[91] wl[278] vdd gnd cell_6t
Xbit_r279_c91 bl[91] br[91] wl[279] vdd gnd cell_6t
Xbit_r280_c91 bl[91] br[91] wl[280] vdd gnd cell_6t
Xbit_r281_c91 bl[91] br[91] wl[281] vdd gnd cell_6t
Xbit_r282_c91 bl[91] br[91] wl[282] vdd gnd cell_6t
Xbit_r283_c91 bl[91] br[91] wl[283] vdd gnd cell_6t
Xbit_r284_c91 bl[91] br[91] wl[284] vdd gnd cell_6t
Xbit_r285_c91 bl[91] br[91] wl[285] vdd gnd cell_6t
Xbit_r286_c91 bl[91] br[91] wl[286] vdd gnd cell_6t
Xbit_r287_c91 bl[91] br[91] wl[287] vdd gnd cell_6t
Xbit_r288_c91 bl[91] br[91] wl[288] vdd gnd cell_6t
Xbit_r289_c91 bl[91] br[91] wl[289] vdd gnd cell_6t
Xbit_r290_c91 bl[91] br[91] wl[290] vdd gnd cell_6t
Xbit_r291_c91 bl[91] br[91] wl[291] vdd gnd cell_6t
Xbit_r292_c91 bl[91] br[91] wl[292] vdd gnd cell_6t
Xbit_r293_c91 bl[91] br[91] wl[293] vdd gnd cell_6t
Xbit_r294_c91 bl[91] br[91] wl[294] vdd gnd cell_6t
Xbit_r295_c91 bl[91] br[91] wl[295] vdd gnd cell_6t
Xbit_r296_c91 bl[91] br[91] wl[296] vdd gnd cell_6t
Xbit_r297_c91 bl[91] br[91] wl[297] vdd gnd cell_6t
Xbit_r298_c91 bl[91] br[91] wl[298] vdd gnd cell_6t
Xbit_r299_c91 bl[91] br[91] wl[299] vdd gnd cell_6t
Xbit_r300_c91 bl[91] br[91] wl[300] vdd gnd cell_6t
Xbit_r301_c91 bl[91] br[91] wl[301] vdd gnd cell_6t
Xbit_r302_c91 bl[91] br[91] wl[302] vdd gnd cell_6t
Xbit_r303_c91 bl[91] br[91] wl[303] vdd gnd cell_6t
Xbit_r304_c91 bl[91] br[91] wl[304] vdd gnd cell_6t
Xbit_r305_c91 bl[91] br[91] wl[305] vdd gnd cell_6t
Xbit_r306_c91 bl[91] br[91] wl[306] vdd gnd cell_6t
Xbit_r307_c91 bl[91] br[91] wl[307] vdd gnd cell_6t
Xbit_r308_c91 bl[91] br[91] wl[308] vdd gnd cell_6t
Xbit_r309_c91 bl[91] br[91] wl[309] vdd gnd cell_6t
Xbit_r310_c91 bl[91] br[91] wl[310] vdd gnd cell_6t
Xbit_r311_c91 bl[91] br[91] wl[311] vdd gnd cell_6t
Xbit_r312_c91 bl[91] br[91] wl[312] vdd gnd cell_6t
Xbit_r313_c91 bl[91] br[91] wl[313] vdd gnd cell_6t
Xbit_r314_c91 bl[91] br[91] wl[314] vdd gnd cell_6t
Xbit_r315_c91 bl[91] br[91] wl[315] vdd gnd cell_6t
Xbit_r316_c91 bl[91] br[91] wl[316] vdd gnd cell_6t
Xbit_r317_c91 bl[91] br[91] wl[317] vdd gnd cell_6t
Xbit_r318_c91 bl[91] br[91] wl[318] vdd gnd cell_6t
Xbit_r319_c91 bl[91] br[91] wl[319] vdd gnd cell_6t
Xbit_r320_c91 bl[91] br[91] wl[320] vdd gnd cell_6t
Xbit_r321_c91 bl[91] br[91] wl[321] vdd gnd cell_6t
Xbit_r322_c91 bl[91] br[91] wl[322] vdd gnd cell_6t
Xbit_r323_c91 bl[91] br[91] wl[323] vdd gnd cell_6t
Xbit_r324_c91 bl[91] br[91] wl[324] vdd gnd cell_6t
Xbit_r325_c91 bl[91] br[91] wl[325] vdd gnd cell_6t
Xbit_r326_c91 bl[91] br[91] wl[326] vdd gnd cell_6t
Xbit_r327_c91 bl[91] br[91] wl[327] vdd gnd cell_6t
Xbit_r328_c91 bl[91] br[91] wl[328] vdd gnd cell_6t
Xbit_r329_c91 bl[91] br[91] wl[329] vdd gnd cell_6t
Xbit_r330_c91 bl[91] br[91] wl[330] vdd gnd cell_6t
Xbit_r331_c91 bl[91] br[91] wl[331] vdd gnd cell_6t
Xbit_r332_c91 bl[91] br[91] wl[332] vdd gnd cell_6t
Xbit_r333_c91 bl[91] br[91] wl[333] vdd gnd cell_6t
Xbit_r334_c91 bl[91] br[91] wl[334] vdd gnd cell_6t
Xbit_r335_c91 bl[91] br[91] wl[335] vdd gnd cell_6t
Xbit_r336_c91 bl[91] br[91] wl[336] vdd gnd cell_6t
Xbit_r337_c91 bl[91] br[91] wl[337] vdd gnd cell_6t
Xbit_r338_c91 bl[91] br[91] wl[338] vdd gnd cell_6t
Xbit_r339_c91 bl[91] br[91] wl[339] vdd gnd cell_6t
Xbit_r340_c91 bl[91] br[91] wl[340] vdd gnd cell_6t
Xbit_r341_c91 bl[91] br[91] wl[341] vdd gnd cell_6t
Xbit_r342_c91 bl[91] br[91] wl[342] vdd gnd cell_6t
Xbit_r343_c91 bl[91] br[91] wl[343] vdd gnd cell_6t
Xbit_r344_c91 bl[91] br[91] wl[344] vdd gnd cell_6t
Xbit_r345_c91 bl[91] br[91] wl[345] vdd gnd cell_6t
Xbit_r346_c91 bl[91] br[91] wl[346] vdd gnd cell_6t
Xbit_r347_c91 bl[91] br[91] wl[347] vdd gnd cell_6t
Xbit_r348_c91 bl[91] br[91] wl[348] vdd gnd cell_6t
Xbit_r349_c91 bl[91] br[91] wl[349] vdd gnd cell_6t
Xbit_r350_c91 bl[91] br[91] wl[350] vdd gnd cell_6t
Xbit_r351_c91 bl[91] br[91] wl[351] vdd gnd cell_6t
Xbit_r352_c91 bl[91] br[91] wl[352] vdd gnd cell_6t
Xbit_r353_c91 bl[91] br[91] wl[353] vdd gnd cell_6t
Xbit_r354_c91 bl[91] br[91] wl[354] vdd gnd cell_6t
Xbit_r355_c91 bl[91] br[91] wl[355] vdd gnd cell_6t
Xbit_r356_c91 bl[91] br[91] wl[356] vdd gnd cell_6t
Xbit_r357_c91 bl[91] br[91] wl[357] vdd gnd cell_6t
Xbit_r358_c91 bl[91] br[91] wl[358] vdd gnd cell_6t
Xbit_r359_c91 bl[91] br[91] wl[359] vdd gnd cell_6t
Xbit_r360_c91 bl[91] br[91] wl[360] vdd gnd cell_6t
Xbit_r361_c91 bl[91] br[91] wl[361] vdd gnd cell_6t
Xbit_r362_c91 bl[91] br[91] wl[362] vdd gnd cell_6t
Xbit_r363_c91 bl[91] br[91] wl[363] vdd gnd cell_6t
Xbit_r364_c91 bl[91] br[91] wl[364] vdd gnd cell_6t
Xbit_r365_c91 bl[91] br[91] wl[365] vdd gnd cell_6t
Xbit_r366_c91 bl[91] br[91] wl[366] vdd gnd cell_6t
Xbit_r367_c91 bl[91] br[91] wl[367] vdd gnd cell_6t
Xbit_r368_c91 bl[91] br[91] wl[368] vdd gnd cell_6t
Xbit_r369_c91 bl[91] br[91] wl[369] vdd gnd cell_6t
Xbit_r370_c91 bl[91] br[91] wl[370] vdd gnd cell_6t
Xbit_r371_c91 bl[91] br[91] wl[371] vdd gnd cell_6t
Xbit_r372_c91 bl[91] br[91] wl[372] vdd gnd cell_6t
Xbit_r373_c91 bl[91] br[91] wl[373] vdd gnd cell_6t
Xbit_r374_c91 bl[91] br[91] wl[374] vdd gnd cell_6t
Xbit_r375_c91 bl[91] br[91] wl[375] vdd gnd cell_6t
Xbit_r376_c91 bl[91] br[91] wl[376] vdd gnd cell_6t
Xbit_r377_c91 bl[91] br[91] wl[377] vdd gnd cell_6t
Xbit_r378_c91 bl[91] br[91] wl[378] vdd gnd cell_6t
Xbit_r379_c91 bl[91] br[91] wl[379] vdd gnd cell_6t
Xbit_r380_c91 bl[91] br[91] wl[380] vdd gnd cell_6t
Xbit_r381_c91 bl[91] br[91] wl[381] vdd gnd cell_6t
Xbit_r382_c91 bl[91] br[91] wl[382] vdd gnd cell_6t
Xbit_r383_c91 bl[91] br[91] wl[383] vdd gnd cell_6t
Xbit_r384_c91 bl[91] br[91] wl[384] vdd gnd cell_6t
Xbit_r385_c91 bl[91] br[91] wl[385] vdd gnd cell_6t
Xbit_r386_c91 bl[91] br[91] wl[386] vdd gnd cell_6t
Xbit_r387_c91 bl[91] br[91] wl[387] vdd gnd cell_6t
Xbit_r388_c91 bl[91] br[91] wl[388] vdd gnd cell_6t
Xbit_r389_c91 bl[91] br[91] wl[389] vdd gnd cell_6t
Xbit_r390_c91 bl[91] br[91] wl[390] vdd gnd cell_6t
Xbit_r391_c91 bl[91] br[91] wl[391] vdd gnd cell_6t
Xbit_r392_c91 bl[91] br[91] wl[392] vdd gnd cell_6t
Xbit_r393_c91 bl[91] br[91] wl[393] vdd gnd cell_6t
Xbit_r394_c91 bl[91] br[91] wl[394] vdd gnd cell_6t
Xbit_r395_c91 bl[91] br[91] wl[395] vdd gnd cell_6t
Xbit_r396_c91 bl[91] br[91] wl[396] vdd gnd cell_6t
Xbit_r397_c91 bl[91] br[91] wl[397] vdd gnd cell_6t
Xbit_r398_c91 bl[91] br[91] wl[398] vdd gnd cell_6t
Xbit_r399_c91 bl[91] br[91] wl[399] vdd gnd cell_6t
Xbit_r400_c91 bl[91] br[91] wl[400] vdd gnd cell_6t
Xbit_r401_c91 bl[91] br[91] wl[401] vdd gnd cell_6t
Xbit_r402_c91 bl[91] br[91] wl[402] vdd gnd cell_6t
Xbit_r403_c91 bl[91] br[91] wl[403] vdd gnd cell_6t
Xbit_r404_c91 bl[91] br[91] wl[404] vdd gnd cell_6t
Xbit_r405_c91 bl[91] br[91] wl[405] vdd gnd cell_6t
Xbit_r406_c91 bl[91] br[91] wl[406] vdd gnd cell_6t
Xbit_r407_c91 bl[91] br[91] wl[407] vdd gnd cell_6t
Xbit_r408_c91 bl[91] br[91] wl[408] vdd gnd cell_6t
Xbit_r409_c91 bl[91] br[91] wl[409] vdd gnd cell_6t
Xbit_r410_c91 bl[91] br[91] wl[410] vdd gnd cell_6t
Xbit_r411_c91 bl[91] br[91] wl[411] vdd gnd cell_6t
Xbit_r412_c91 bl[91] br[91] wl[412] vdd gnd cell_6t
Xbit_r413_c91 bl[91] br[91] wl[413] vdd gnd cell_6t
Xbit_r414_c91 bl[91] br[91] wl[414] vdd gnd cell_6t
Xbit_r415_c91 bl[91] br[91] wl[415] vdd gnd cell_6t
Xbit_r416_c91 bl[91] br[91] wl[416] vdd gnd cell_6t
Xbit_r417_c91 bl[91] br[91] wl[417] vdd gnd cell_6t
Xbit_r418_c91 bl[91] br[91] wl[418] vdd gnd cell_6t
Xbit_r419_c91 bl[91] br[91] wl[419] vdd gnd cell_6t
Xbit_r420_c91 bl[91] br[91] wl[420] vdd gnd cell_6t
Xbit_r421_c91 bl[91] br[91] wl[421] vdd gnd cell_6t
Xbit_r422_c91 bl[91] br[91] wl[422] vdd gnd cell_6t
Xbit_r423_c91 bl[91] br[91] wl[423] vdd gnd cell_6t
Xbit_r424_c91 bl[91] br[91] wl[424] vdd gnd cell_6t
Xbit_r425_c91 bl[91] br[91] wl[425] vdd gnd cell_6t
Xbit_r426_c91 bl[91] br[91] wl[426] vdd gnd cell_6t
Xbit_r427_c91 bl[91] br[91] wl[427] vdd gnd cell_6t
Xbit_r428_c91 bl[91] br[91] wl[428] vdd gnd cell_6t
Xbit_r429_c91 bl[91] br[91] wl[429] vdd gnd cell_6t
Xbit_r430_c91 bl[91] br[91] wl[430] vdd gnd cell_6t
Xbit_r431_c91 bl[91] br[91] wl[431] vdd gnd cell_6t
Xbit_r432_c91 bl[91] br[91] wl[432] vdd gnd cell_6t
Xbit_r433_c91 bl[91] br[91] wl[433] vdd gnd cell_6t
Xbit_r434_c91 bl[91] br[91] wl[434] vdd gnd cell_6t
Xbit_r435_c91 bl[91] br[91] wl[435] vdd gnd cell_6t
Xbit_r436_c91 bl[91] br[91] wl[436] vdd gnd cell_6t
Xbit_r437_c91 bl[91] br[91] wl[437] vdd gnd cell_6t
Xbit_r438_c91 bl[91] br[91] wl[438] vdd gnd cell_6t
Xbit_r439_c91 bl[91] br[91] wl[439] vdd gnd cell_6t
Xbit_r440_c91 bl[91] br[91] wl[440] vdd gnd cell_6t
Xbit_r441_c91 bl[91] br[91] wl[441] vdd gnd cell_6t
Xbit_r442_c91 bl[91] br[91] wl[442] vdd gnd cell_6t
Xbit_r443_c91 bl[91] br[91] wl[443] vdd gnd cell_6t
Xbit_r444_c91 bl[91] br[91] wl[444] vdd gnd cell_6t
Xbit_r445_c91 bl[91] br[91] wl[445] vdd gnd cell_6t
Xbit_r446_c91 bl[91] br[91] wl[446] vdd gnd cell_6t
Xbit_r447_c91 bl[91] br[91] wl[447] vdd gnd cell_6t
Xbit_r448_c91 bl[91] br[91] wl[448] vdd gnd cell_6t
Xbit_r449_c91 bl[91] br[91] wl[449] vdd gnd cell_6t
Xbit_r450_c91 bl[91] br[91] wl[450] vdd gnd cell_6t
Xbit_r451_c91 bl[91] br[91] wl[451] vdd gnd cell_6t
Xbit_r452_c91 bl[91] br[91] wl[452] vdd gnd cell_6t
Xbit_r453_c91 bl[91] br[91] wl[453] vdd gnd cell_6t
Xbit_r454_c91 bl[91] br[91] wl[454] vdd gnd cell_6t
Xbit_r455_c91 bl[91] br[91] wl[455] vdd gnd cell_6t
Xbit_r456_c91 bl[91] br[91] wl[456] vdd gnd cell_6t
Xbit_r457_c91 bl[91] br[91] wl[457] vdd gnd cell_6t
Xbit_r458_c91 bl[91] br[91] wl[458] vdd gnd cell_6t
Xbit_r459_c91 bl[91] br[91] wl[459] vdd gnd cell_6t
Xbit_r460_c91 bl[91] br[91] wl[460] vdd gnd cell_6t
Xbit_r461_c91 bl[91] br[91] wl[461] vdd gnd cell_6t
Xbit_r462_c91 bl[91] br[91] wl[462] vdd gnd cell_6t
Xbit_r463_c91 bl[91] br[91] wl[463] vdd gnd cell_6t
Xbit_r464_c91 bl[91] br[91] wl[464] vdd gnd cell_6t
Xbit_r465_c91 bl[91] br[91] wl[465] vdd gnd cell_6t
Xbit_r466_c91 bl[91] br[91] wl[466] vdd gnd cell_6t
Xbit_r467_c91 bl[91] br[91] wl[467] vdd gnd cell_6t
Xbit_r468_c91 bl[91] br[91] wl[468] vdd gnd cell_6t
Xbit_r469_c91 bl[91] br[91] wl[469] vdd gnd cell_6t
Xbit_r470_c91 bl[91] br[91] wl[470] vdd gnd cell_6t
Xbit_r471_c91 bl[91] br[91] wl[471] vdd gnd cell_6t
Xbit_r472_c91 bl[91] br[91] wl[472] vdd gnd cell_6t
Xbit_r473_c91 bl[91] br[91] wl[473] vdd gnd cell_6t
Xbit_r474_c91 bl[91] br[91] wl[474] vdd gnd cell_6t
Xbit_r475_c91 bl[91] br[91] wl[475] vdd gnd cell_6t
Xbit_r476_c91 bl[91] br[91] wl[476] vdd gnd cell_6t
Xbit_r477_c91 bl[91] br[91] wl[477] vdd gnd cell_6t
Xbit_r478_c91 bl[91] br[91] wl[478] vdd gnd cell_6t
Xbit_r479_c91 bl[91] br[91] wl[479] vdd gnd cell_6t
Xbit_r480_c91 bl[91] br[91] wl[480] vdd gnd cell_6t
Xbit_r481_c91 bl[91] br[91] wl[481] vdd gnd cell_6t
Xbit_r482_c91 bl[91] br[91] wl[482] vdd gnd cell_6t
Xbit_r483_c91 bl[91] br[91] wl[483] vdd gnd cell_6t
Xbit_r484_c91 bl[91] br[91] wl[484] vdd gnd cell_6t
Xbit_r485_c91 bl[91] br[91] wl[485] vdd gnd cell_6t
Xbit_r486_c91 bl[91] br[91] wl[486] vdd gnd cell_6t
Xbit_r487_c91 bl[91] br[91] wl[487] vdd gnd cell_6t
Xbit_r488_c91 bl[91] br[91] wl[488] vdd gnd cell_6t
Xbit_r489_c91 bl[91] br[91] wl[489] vdd gnd cell_6t
Xbit_r490_c91 bl[91] br[91] wl[490] vdd gnd cell_6t
Xbit_r491_c91 bl[91] br[91] wl[491] vdd gnd cell_6t
Xbit_r492_c91 bl[91] br[91] wl[492] vdd gnd cell_6t
Xbit_r493_c91 bl[91] br[91] wl[493] vdd gnd cell_6t
Xbit_r494_c91 bl[91] br[91] wl[494] vdd gnd cell_6t
Xbit_r495_c91 bl[91] br[91] wl[495] vdd gnd cell_6t
Xbit_r496_c91 bl[91] br[91] wl[496] vdd gnd cell_6t
Xbit_r497_c91 bl[91] br[91] wl[497] vdd gnd cell_6t
Xbit_r498_c91 bl[91] br[91] wl[498] vdd gnd cell_6t
Xbit_r499_c91 bl[91] br[91] wl[499] vdd gnd cell_6t
Xbit_r500_c91 bl[91] br[91] wl[500] vdd gnd cell_6t
Xbit_r501_c91 bl[91] br[91] wl[501] vdd gnd cell_6t
Xbit_r502_c91 bl[91] br[91] wl[502] vdd gnd cell_6t
Xbit_r503_c91 bl[91] br[91] wl[503] vdd gnd cell_6t
Xbit_r504_c91 bl[91] br[91] wl[504] vdd gnd cell_6t
Xbit_r505_c91 bl[91] br[91] wl[505] vdd gnd cell_6t
Xbit_r506_c91 bl[91] br[91] wl[506] vdd gnd cell_6t
Xbit_r507_c91 bl[91] br[91] wl[507] vdd gnd cell_6t
Xbit_r508_c91 bl[91] br[91] wl[508] vdd gnd cell_6t
Xbit_r509_c91 bl[91] br[91] wl[509] vdd gnd cell_6t
Xbit_r510_c91 bl[91] br[91] wl[510] vdd gnd cell_6t
Xbit_r511_c91 bl[91] br[91] wl[511] vdd gnd cell_6t
Xbit_r0_c92 bl[92] br[92] wl[0] vdd gnd cell_6t
Xbit_r1_c92 bl[92] br[92] wl[1] vdd gnd cell_6t
Xbit_r2_c92 bl[92] br[92] wl[2] vdd gnd cell_6t
Xbit_r3_c92 bl[92] br[92] wl[3] vdd gnd cell_6t
Xbit_r4_c92 bl[92] br[92] wl[4] vdd gnd cell_6t
Xbit_r5_c92 bl[92] br[92] wl[5] vdd gnd cell_6t
Xbit_r6_c92 bl[92] br[92] wl[6] vdd gnd cell_6t
Xbit_r7_c92 bl[92] br[92] wl[7] vdd gnd cell_6t
Xbit_r8_c92 bl[92] br[92] wl[8] vdd gnd cell_6t
Xbit_r9_c92 bl[92] br[92] wl[9] vdd gnd cell_6t
Xbit_r10_c92 bl[92] br[92] wl[10] vdd gnd cell_6t
Xbit_r11_c92 bl[92] br[92] wl[11] vdd gnd cell_6t
Xbit_r12_c92 bl[92] br[92] wl[12] vdd gnd cell_6t
Xbit_r13_c92 bl[92] br[92] wl[13] vdd gnd cell_6t
Xbit_r14_c92 bl[92] br[92] wl[14] vdd gnd cell_6t
Xbit_r15_c92 bl[92] br[92] wl[15] vdd gnd cell_6t
Xbit_r16_c92 bl[92] br[92] wl[16] vdd gnd cell_6t
Xbit_r17_c92 bl[92] br[92] wl[17] vdd gnd cell_6t
Xbit_r18_c92 bl[92] br[92] wl[18] vdd gnd cell_6t
Xbit_r19_c92 bl[92] br[92] wl[19] vdd gnd cell_6t
Xbit_r20_c92 bl[92] br[92] wl[20] vdd gnd cell_6t
Xbit_r21_c92 bl[92] br[92] wl[21] vdd gnd cell_6t
Xbit_r22_c92 bl[92] br[92] wl[22] vdd gnd cell_6t
Xbit_r23_c92 bl[92] br[92] wl[23] vdd gnd cell_6t
Xbit_r24_c92 bl[92] br[92] wl[24] vdd gnd cell_6t
Xbit_r25_c92 bl[92] br[92] wl[25] vdd gnd cell_6t
Xbit_r26_c92 bl[92] br[92] wl[26] vdd gnd cell_6t
Xbit_r27_c92 bl[92] br[92] wl[27] vdd gnd cell_6t
Xbit_r28_c92 bl[92] br[92] wl[28] vdd gnd cell_6t
Xbit_r29_c92 bl[92] br[92] wl[29] vdd gnd cell_6t
Xbit_r30_c92 bl[92] br[92] wl[30] vdd gnd cell_6t
Xbit_r31_c92 bl[92] br[92] wl[31] vdd gnd cell_6t
Xbit_r32_c92 bl[92] br[92] wl[32] vdd gnd cell_6t
Xbit_r33_c92 bl[92] br[92] wl[33] vdd gnd cell_6t
Xbit_r34_c92 bl[92] br[92] wl[34] vdd gnd cell_6t
Xbit_r35_c92 bl[92] br[92] wl[35] vdd gnd cell_6t
Xbit_r36_c92 bl[92] br[92] wl[36] vdd gnd cell_6t
Xbit_r37_c92 bl[92] br[92] wl[37] vdd gnd cell_6t
Xbit_r38_c92 bl[92] br[92] wl[38] vdd gnd cell_6t
Xbit_r39_c92 bl[92] br[92] wl[39] vdd gnd cell_6t
Xbit_r40_c92 bl[92] br[92] wl[40] vdd gnd cell_6t
Xbit_r41_c92 bl[92] br[92] wl[41] vdd gnd cell_6t
Xbit_r42_c92 bl[92] br[92] wl[42] vdd gnd cell_6t
Xbit_r43_c92 bl[92] br[92] wl[43] vdd gnd cell_6t
Xbit_r44_c92 bl[92] br[92] wl[44] vdd gnd cell_6t
Xbit_r45_c92 bl[92] br[92] wl[45] vdd gnd cell_6t
Xbit_r46_c92 bl[92] br[92] wl[46] vdd gnd cell_6t
Xbit_r47_c92 bl[92] br[92] wl[47] vdd gnd cell_6t
Xbit_r48_c92 bl[92] br[92] wl[48] vdd gnd cell_6t
Xbit_r49_c92 bl[92] br[92] wl[49] vdd gnd cell_6t
Xbit_r50_c92 bl[92] br[92] wl[50] vdd gnd cell_6t
Xbit_r51_c92 bl[92] br[92] wl[51] vdd gnd cell_6t
Xbit_r52_c92 bl[92] br[92] wl[52] vdd gnd cell_6t
Xbit_r53_c92 bl[92] br[92] wl[53] vdd gnd cell_6t
Xbit_r54_c92 bl[92] br[92] wl[54] vdd gnd cell_6t
Xbit_r55_c92 bl[92] br[92] wl[55] vdd gnd cell_6t
Xbit_r56_c92 bl[92] br[92] wl[56] vdd gnd cell_6t
Xbit_r57_c92 bl[92] br[92] wl[57] vdd gnd cell_6t
Xbit_r58_c92 bl[92] br[92] wl[58] vdd gnd cell_6t
Xbit_r59_c92 bl[92] br[92] wl[59] vdd gnd cell_6t
Xbit_r60_c92 bl[92] br[92] wl[60] vdd gnd cell_6t
Xbit_r61_c92 bl[92] br[92] wl[61] vdd gnd cell_6t
Xbit_r62_c92 bl[92] br[92] wl[62] vdd gnd cell_6t
Xbit_r63_c92 bl[92] br[92] wl[63] vdd gnd cell_6t
Xbit_r64_c92 bl[92] br[92] wl[64] vdd gnd cell_6t
Xbit_r65_c92 bl[92] br[92] wl[65] vdd gnd cell_6t
Xbit_r66_c92 bl[92] br[92] wl[66] vdd gnd cell_6t
Xbit_r67_c92 bl[92] br[92] wl[67] vdd gnd cell_6t
Xbit_r68_c92 bl[92] br[92] wl[68] vdd gnd cell_6t
Xbit_r69_c92 bl[92] br[92] wl[69] vdd gnd cell_6t
Xbit_r70_c92 bl[92] br[92] wl[70] vdd gnd cell_6t
Xbit_r71_c92 bl[92] br[92] wl[71] vdd gnd cell_6t
Xbit_r72_c92 bl[92] br[92] wl[72] vdd gnd cell_6t
Xbit_r73_c92 bl[92] br[92] wl[73] vdd gnd cell_6t
Xbit_r74_c92 bl[92] br[92] wl[74] vdd gnd cell_6t
Xbit_r75_c92 bl[92] br[92] wl[75] vdd gnd cell_6t
Xbit_r76_c92 bl[92] br[92] wl[76] vdd gnd cell_6t
Xbit_r77_c92 bl[92] br[92] wl[77] vdd gnd cell_6t
Xbit_r78_c92 bl[92] br[92] wl[78] vdd gnd cell_6t
Xbit_r79_c92 bl[92] br[92] wl[79] vdd gnd cell_6t
Xbit_r80_c92 bl[92] br[92] wl[80] vdd gnd cell_6t
Xbit_r81_c92 bl[92] br[92] wl[81] vdd gnd cell_6t
Xbit_r82_c92 bl[92] br[92] wl[82] vdd gnd cell_6t
Xbit_r83_c92 bl[92] br[92] wl[83] vdd gnd cell_6t
Xbit_r84_c92 bl[92] br[92] wl[84] vdd gnd cell_6t
Xbit_r85_c92 bl[92] br[92] wl[85] vdd gnd cell_6t
Xbit_r86_c92 bl[92] br[92] wl[86] vdd gnd cell_6t
Xbit_r87_c92 bl[92] br[92] wl[87] vdd gnd cell_6t
Xbit_r88_c92 bl[92] br[92] wl[88] vdd gnd cell_6t
Xbit_r89_c92 bl[92] br[92] wl[89] vdd gnd cell_6t
Xbit_r90_c92 bl[92] br[92] wl[90] vdd gnd cell_6t
Xbit_r91_c92 bl[92] br[92] wl[91] vdd gnd cell_6t
Xbit_r92_c92 bl[92] br[92] wl[92] vdd gnd cell_6t
Xbit_r93_c92 bl[92] br[92] wl[93] vdd gnd cell_6t
Xbit_r94_c92 bl[92] br[92] wl[94] vdd gnd cell_6t
Xbit_r95_c92 bl[92] br[92] wl[95] vdd gnd cell_6t
Xbit_r96_c92 bl[92] br[92] wl[96] vdd gnd cell_6t
Xbit_r97_c92 bl[92] br[92] wl[97] vdd gnd cell_6t
Xbit_r98_c92 bl[92] br[92] wl[98] vdd gnd cell_6t
Xbit_r99_c92 bl[92] br[92] wl[99] vdd gnd cell_6t
Xbit_r100_c92 bl[92] br[92] wl[100] vdd gnd cell_6t
Xbit_r101_c92 bl[92] br[92] wl[101] vdd gnd cell_6t
Xbit_r102_c92 bl[92] br[92] wl[102] vdd gnd cell_6t
Xbit_r103_c92 bl[92] br[92] wl[103] vdd gnd cell_6t
Xbit_r104_c92 bl[92] br[92] wl[104] vdd gnd cell_6t
Xbit_r105_c92 bl[92] br[92] wl[105] vdd gnd cell_6t
Xbit_r106_c92 bl[92] br[92] wl[106] vdd gnd cell_6t
Xbit_r107_c92 bl[92] br[92] wl[107] vdd gnd cell_6t
Xbit_r108_c92 bl[92] br[92] wl[108] vdd gnd cell_6t
Xbit_r109_c92 bl[92] br[92] wl[109] vdd gnd cell_6t
Xbit_r110_c92 bl[92] br[92] wl[110] vdd gnd cell_6t
Xbit_r111_c92 bl[92] br[92] wl[111] vdd gnd cell_6t
Xbit_r112_c92 bl[92] br[92] wl[112] vdd gnd cell_6t
Xbit_r113_c92 bl[92] br[92] wl[113] vdd gnd cell_6t
Xbit_r114_c92 bl[92] br[92] wl[114] vdd gnd cell_6t
Xbit_r115_c92 bl[92] br[92] wl[115] vdd gnd cell_6t
Xbit_r116_c92 bl[92] br[92] wl[116] vdd gnd cell_6t
Xbit_r117_c92 bl[92] br[92] wl[117] vdd gnd cell_6t
Xbit_r118_c92 bl[92] br[92] wl[118] vdd gnd cell_6t
Xbit_r119_c92 bl[92] br[92] wl[119] vdd gnd cell_6t
Xbit_r120_c92 bl[92] br[92] wl[120] vdd gnd cell_6t
Xbit_r121_c92 bl[92] br[92] wl[121] vdd gnd cell_6t
Xbit_r122_c92 bl[92] br[92] wl[122] vdd gnd cell_6t
Xbit_r123_c92 bl[92] br[92] wl[123] vdd gnd cell_6t
Xbit_r124_c92 bl[92] br[92] wl[124] vdd gnd cell_6t
Xbit_r125_c92 bl[92] br[92] wl[125] vdd gnd cell_6t
Xbit_r126_c92 bl[92] br[92] wl[126] vdd gnd cell_6t
Xbit_r127_c92 bl[92] br[92] wl[127] vdd gnd cell_6t
Xbit_r128_c92 bl[92] br[92] wl[128] vdd gnd cell_6t
Xbit_r129_c92 bl[92] br[92] wl[129] vdd gnd cell_6t
Xbit_r130_c92 bl[92] br[92] wl[130] vdd gnd cell_6t
Xbit_r131_c92 bl[92] br[92] wl[131] vdd gnd cell_6t
Xbit_r132_c92 bl[92] br[92] wl[132] vdd gnd cell_6t
Xbit_r133_c92 bl[92] br[92] wl[133] vdd gnd cell_6t
Xbit_r134_c92 bl[92] br[92] wl[134] vdd gnd cell_6t
Xbit_r135_c92 bl[92] br[92] wl[135] vdd gnd cell_6t
Xbit_r136_c92 bl[92] br[92] wl[136] vdd gnd cell_6t
Xbit_r137_c92 bl[92] br[92] wl[137] vdd gnd cell_6t
Xbit_r138_c92 bl[92] br[92] wl[138] vdd gnd cell_6t
Xbit_r139_c92 bl[92] br[92] wl[139] vdd gnd cell_6t
Xbit_r140_c92 bl[92] br[92] wl[140] vdd gnd cell_6t
Xbit_r141_c92 bl[92] br[92] wl[141] vdd gnd cell_6t
Xbit_r142_c92 bl[92] br[92] wl[142] vdd gnd cell_6t
Xbit_r143_c92 bl[92] br[92] wl[143] vdd gnd cell_6t
Xbit_r144_c92 bl[92] br[92] wl[144] vdd gnd cell_6t
Xbit_r145_c92 bl[92] br[92] wl[145] vdd gnd cell_6t
Xbit_r146_c92 bl[92] br[92] wl[146] vdd gnd cell_6t
Xbit_r147_c92 bl[92] br[92] wl[147] vdd gnd cell_6t
Xbit_r148_c92 bl[92] br[92] wl[148] vdd gnd cell_6t
Xbit_r149_c92 bl[92] br[92] wl[149] vdd gnd cell_6t
Xbit_r150_c92 bl[92] br[92] wl[150] vdd gnd cell_6t
Xbit_r151_c92 bl[92] br[92] wl[151] vdd gnd cell_6t
Xbit_r152_c92 bl[92] br[92] wl[152] vdd gnd cell_6t
Xbit_r153_c92 bl[92] br[92] wl[153] vdd gnd cell_6t
Xbit_r154_c92 bl[92] br[92] wl[154] vdd gnd cell_6t
Xbit_r155_c92 bl[92] br[92] wl[155] vdd gnd cell_6t
Xbit_r156_c92 bl[92] br[92] wl[156] vdd gnd cell_6t
Xbit_r157_c92 bl[92] br[92] wl[157] vdd gnd cell_6t
Xbit_r158_c92 bl[92] br[92] wl[158] vdd gnd cell_6t
Xbit_r159_c92 bl[92] br[92] wl[159] vdd gnd cell_6t
Xbit_r160_c92 bl[92] br[92] wl[160] vdd gnd cell_6t
Xbit_r161_c92 bl[92] br[92] wl[161] vdd gnd cell_6t
Xbit_r162_c92 bl[92] br[92] wl[162] vdd gnd cell_6t
Xbit_r163_c92 bl[92] br[92] wl[163] vdd gnd cell_6t
Xbit_r164_c92 bl[92] br[92] wl[164] vdd gnd cell_6t
Xbit_r165_c92 bl[92] br[92] wl[165] vdd gnd cell_6t
Xbit_r166_c92 bl[92] br[92] wl[166] vdd gnd cell_6t
Xbit_r167_c92 bl[92] br[92] wl[167] vdd gnd cell_6t
Xbit_r168_c92 bl[92] br[92] wl[168] vdd gnd cell_6t
Xbit_r169_c92 bl[92] br[92] wl[169] vdd gnd cell_6t
Xbit_r170_c92 bl[92] br[92] wl[170] vdd gnd cell_6t
Xbit_r171_c92 bl[92] br[92] wl[171] vdd gnd cell_6t
Xbit_r172_c92 bl[92] br[92] wl[172] vdd gnd cell_6t
Xbit_r173_c92 bl[92] br[92] wl[173] vdd gnd cell_6t
Xbit_r174_c92 bl[92] br[92] wl[174] vdd gnd cell_6t
Xbit_r175_c92 bl[92] br[92] wl[175] vdd gnd cell_6t
Xbit_r176_c92 bl[92] br[92] wl[176] vdd gnd cell_6t
Xbit_r177_c92 bl[92] br[92] wl[177] vdd gnd cell_6t
Xbit_r178_c92 bl[92] br[92] wl[178] vdd gnd cell_6t
Xbit_r179_c92 bl[92] br[92] wl[179] vdd gnd cell_6t
Xbit_r180_c92 bl[92] br[92] wl[180] vdd gnd cell_6t
Xbit_r181_c92 bl[92] br[92] wl[181] vdd gnd cell_6t
Xbit_r182_c92 bl[92] br[92] wl[182] vdd gnd cell_6t
Xbit_r183_c92 bl[92] br[92] wl[183] vdd gnd cell_6t
Xbit_r184_c92 bl[92] br[92] wl[184] vdd gnd cell_6t
Xbit_r185_c92 bl[92] br[92] wl[185] vdd gnd cell_6t
Xbit_r186_c92 bl[92] br[92] wl[186] vdd gnd cell_6t
Xbit_r187_c92 bl[92] br[92] wl[187] vdd gnd cell_6t
Xbit_r188_c92 bl[92] br[92] wl[188] vdd gnd cell_6t
Xbit_r189_c92 bl[92] br[92] wl[189] vdd gnd cell_6t
Xbit_r190_c92 bl[92] br[92] wl[190] vdd gnd cell_6t
Xbit_r191_c92 bl[92] br[92] wl[191] vdd gnd cell_6t
Xbit_r192_c92 bl[92] br[92] wl[192] vdd gnd cell_6t
Xbit_r193_c92 bl[92] br[92] wl[193] vdd gnd cell_6t
Xbit_r194_c92 bl[92] br[92] wl[194] vdd gnd cell_6t
Xbit_r195_c92 bl[92] br[92] wl[195] vdd gnd cell_6t
Xbit_r196_c92 bl[92] br[92] wl[196] vdd gnd cell_6t
Xbit_r197_c92 bl[92] br[92] wl[197] vdd gnd cell_6t
Xbit_r198_c92 bl[92] br[92] wl[198] vdd gnd cell_6t
Xbit_r199_c92 bl[92] br[92] wl[199] vdd gnd cell_6t
Xbit_r200_c92 bl[92] br[92] wl[200] vdd gnd cell_6t
Xbit_r201_c92 bl[92] br[92] wl[201] vdd gnd cell_6t
Xbit_r202_c92 bl[92] br[92] wl[202] vdd gnd cell_6t
Xbit_r203_c92 bl[92] br[92] wl[203] vdd gnd cell_6t
Xbit_r204_c92 bl[92] br[92] wl[204] vdd gnd cell_6t
Xbit_r205_c92 bl[92] br[92] wl[205] vdd gnd cell_6t
Xbit_r206_c92 bl[92] br[92] wl[206] vdd gnd cell_6t
Xbit_r207_c92 bl[92] br[92] wl[207] vdd gnd cell_6t
Xbit_r208_c92 bl[92] br[92] wl[208] vdd gnd cell_6t
Xbit_r209_c92 bl[92] br[92] wl[209] vdd gnd cell_6t
Xbit_r210_c92 bl[92] br[92] wl[210] vdd gnd cell_6t
Xbit_r211_c92 bl[92] br[92] wl[211] vdd gnd cell_6t
Xbit_r212_c92 bl[92] br[92] wl[212] vdd gnd cell_6t
Xbit_r213_c92 bl[92] br[92] wl[213] vdd gnd cell_6t
Xbit_r214_c92 bl[92] br[92] wl[214] vdd gnd cell_6t
Xbit_r215_c92 bl[92] br[92] wl[215] vdd gnd cell_6t
Xbit_r216_c92 bl[92] br[92] wl[216] vdd gnd cell_6t
Xbit_r217_c92 bl[92] br[92] wl[217] vdd gnd cell_6t
Xbit_r218_c92 bl[92] br[92] wl[218] vdd gnd cell_6t
Xbit_r219_c92 bl[92] br[92] wl[219] vdd gnd cell_6t
Xbit_r220_c92 bl[92] br[92] wl[220] vdd gnd cell_6t
Xbit_r221_c92 bl[92] br[92] wl[221] vdd gnd cell_6t
Xbit_r222_c92 bl[92] br[92] wl[222] vdd gnd cell_6t
Xbit_r223_c92 bl[92] br[92] wl[223] vdd gnd cell_6t
Xbit_r224_c92 bl[92] br[92] wl[224] vdd gnd cell_6t
Xbit_r225_c92 bl[92] br[92] wl[225] vdd gnd cell_6t
Xbit_r226_c92 bl[92] br[92] wl[226] vdd gnd cell_6t
Xbit_r227_c92 bl[92] br[92] wl[227] vdd gnd cell_6t
Xbit_r228_c92 bl[92] br[92] wl[228] vdd gnd cell_6t
Xbit_r229_c92 bl[92] br[92] wl[229] vdd gnd cell_6t
Xbit_r230_c92 bl[92] br[92] wl[230] vdd gnd cell_6t
Xbit_r231_c92 bl[92] br[92] wl[231] vdd gnd cell_6t
Xbit_r232_c92 bl[92] br[92] wl[232] vdd gnd cell_6t
Xbit_r233_c92 bl[92] br[92] wl[233] vdd gnd cell_6t
Xbit_r234_c92 bl[92] br[92] wl[234] vdd gnd cell_6t
Xbit_r235_c92 bl[92] br[92] wl[235] vdd gnd cell_6t
Xbit_r236_c92 bl[92] br[92] wl[236] vdd gnd cell_6t
Xbit_r237_c92 bl[92] br[92] wl[237] vdd gnd cell_6t
Xbit_r238_c92 bl[92] br[92] wl[238] vdd gnd cell_6t
Xbit_r239_c92 bl[92] br[92] wl[239] vdd gnd cell_6t
Xbit_r240_c92 bl[92] br[92] wl[240] vdd gnd cell_6t
Xbit_r241_c92 bl[92] br[92] wl[241] vdd gnd cell_6t
Xbit_r242_c92 bl[92] br[92] wl[242] vdd gnd cell_6t
Xbit_r243_c92 bl[92] br[92] wl[243] vdd gnd cell_6t
Xbit_r244_c92 bl[92] br[92] wl[244] vdd gnd cell_6t
Xbit_r245_c92 bl[92] br[92] wl[245] vdd gnd cell_6t
Xbit_r246_c92 bl[92] br[92] wl[246] vdd gnd cell_6t
Xbit_r247_c92 bl[92] br[92] wl[247] vdd gnd cell_6t
Xbit_r248_c92 bl[92] br[92] wl[248] vdd gnd cell_6t
Xbit_r249_c92 bl[92] br[92] wl[249] vdd gnd cell_6t
Xbit_r250_c92 bl[92] br[92] wl[250] vdd gnd cell_6t
Xbit_r251_c92 bl[92] br[92] wl[251] vdd gnd cell_6t
Xbit_r252_c92 bl[92] br[92] wl[252] vdd gnd cell_6t
Xbit_r253_c92 bl[92] br[92] wl[253] vdd gnd cell_6t
Xbit_r254_c92 bl[92] br[92] wl[254] vdd gnd cell_6t
Xbit_r255_c92 bl[92] br[92] wl[255] vdd gnd cell_6t
Xbit_r256_c92 bl[92] br[92] wl[256] vdd gnd cell_6t
Xbit_r257_c92 bl[92] br[92] wl[257] vdd gnd cell_6t
Xbit_r258_c92 bl[92] br[92] wl[258] vdd gnd cell_6t
Xbit_r259_c92 bl[92] br[92] wl[259] vdd gnd cell_6t
Xbit_r260_c92 bl[92] br[92] wl[260] vdd gnd cell_6t
Xbit_r261_c92 bl[92] br[92] wl[261] vdd gnd cell_6t
Xbit_r262_c92 bl[92] br[92] wl[262] vdd gnd cell_6t
Xbit_r263_c92 bl[92] br[92] wl[263] vdd gnd cell_6t
Xbit_r264_c92 bl[92] br[92] wl[264] vdd gnd cell_6t
Xbit_r265_c92 bl[92] br[92] wl[265] vdd gnd cell_6t
Xbit_r266_c92 bl[92] br[92] wl[266] vdd gnd cell_6t
Xbit_r267_c92 bl[92] br[92] wl[267] vdd gnd cell_6t
Xbit_r268_c92 bl[92] br[92] wl[268] vdd gnd cell_6t
Xbit_r269_c92 bl[92] br[92] wl[269] vdd gnd cell_6t
Xbit_r270_c92 bl[92] br[92] wl[270] vdd gnd cell_6t
Xbit_r271_c92 bl[92] br[92] wl[271] vdd gnd cell_6t
Xbit_r272_c92 bl[92] br[92] wl[272] vdd gnd cell_6t
Xbit_r273_c92 bl[92] br[92] wl[273] vdd gnd cell_6t
Xbit_r274_c92 bl[92] br[92] wl[274] vdd gnd cell_6t
Xbit_r275_c92 bl[92] br[92] wl[275] vdd gnd cell_6t
Xbit_r276_c92 bl[92] br[92] wl[276] vdd gnd cell_6t
Xbit_r277_c92 bl[92] br[92] wl[277] vdd gnd cell_6t
Xbit_r278_c92 bl[92] br[92] wl[278] vdd gnd cell_6t
Xbit_r279_c92 bl[92] br[92] wl[279] vdd gnd cell_6t
Xbit_r280_c92 bl[92] br[92] wl[280] vdd gnd cell_6t
Xbit_r281_c92 bl[92] br[92] wl[281] vdd gnd cell_6t
Xbit_r282_c92 bl[92] br[92] wl[282] vdd gnd cell_6t
Xbit_r283_c92 bl[92] br[92] wl[283] vdd gnd cell_6t
Xbit_r284_c92 bl[92] br[92] wl[284] vdd gnd cell_6t
Xbit_r285_c92 bl[92] br[92] wl[285] vdd gnd cell_6t
Xbit_r286_c92 bl[92] br[92] wl[286] vdd gnd cell_6t
Xbit_r287_c92 bl[92] br[92] wl[287] vdd gnd cell_6t
Xbit_r288_c92 bl[92] br[92] wl[288] vdd gnd cell_6t
Xbit_r289_c92 bl[92] br[92] wl[289] vdd gnd cell_6t
Xbit_r290_c92 bl[92] br[92] wl[290] vdd gnd cell_6t
Xbit_r291_c92 bl[92] br[92] wl[291] vdd gnd cell_6t
Xbit_r292_c92 bl[92] br[92] wl[292] vdd gnd cell_6t
Xbit_r293_c92 bl[92] br[92] wl[293] vdd gnd cell_6t
Xbit_r294_c92 bl[92] br[92] wl[294] vdd gnd cell_6t
Xbit_r295_c92 bl[92] br[92] wl[295] vdd gnd cell_6t
Xbit_r296_c92 bl[92] br[92] wl[296] vdd gnd cell_6t
Xbit_r297_c92 bl[92] br[92] wl[297] vdd gnd cell_6t
Xbit_r298_c92 bl[92] br[92] wl[298] vdd gnd cell_6t
Xbit_r299_c92 bl[92] br[92] wl[299] vdd gnd cell_6t
Xbit_r300_c92 bl[92] br[92] wl[300] vdd gnd cell_6t
Xbit_r301_c92 bl[92] br[92] wl[301] vdd gnd cell_6t
Xbit_r302_c92 bl[92] br[92] wl[302] vdd gnd cell_6t
Xbit_r303_c92 bl[92] br[92] wl[303] vdd gnd cell_6t
Xbit_r304_c92 bl[92] br[92] wl[304] vdd gnd cell_6t
Xbit_r305_c92 bl[92] br[92] wl[305] vdd gnd cell_6t
Xbit_r306_c92 bl[92] br[92] wl[306] vdd gnd cell_6t
Xbit_r307_c92 bl[92] br[92] wl[307] vdd gnd cell_6t
Xbit_r308_c92 bl[92] br[92] wl[308] vdd gnd cell_6t
Xbit_r309_c92 bl[92] br[92] wl[309] vdd gnd cell_6t
Xbit_r310_c92 bl[92] br[92] wl[310] vdd gnd cell_6t
Xbit_r311_c92 bl[92] br[92] wl[311] vdd gnd cell_6t
Xbit_r312_c92 bl[92] br[92] wl[312] vdd gnd cell_6t
Xbit_r313_c92 bl[92] br[92] wl[313] vdd gnd cell_6t
Xbit_r314_c92 bl[92] br[92] wl[314] vdd gnd cell_6t
Xbit_r315_c92 bl[92] br[92] wl[315] vdd gnd cell_6t
Xbit_r316_c92 bl[92] br[92] wl[316] vdd gnd cell_6t
Xbit_r317_c92 bl[92] br[92] wl[317] vdd gnd cell_6t
Xbit_r318_c92 bl[92] br[92] wl[318] vdd gnd cell_6t
Xbit_r319_c92 bl[92] br[92] wl[319] vdd gnd cell_6t
Xbit_r320_c92 bl[92] br[92] wl[320] vdd gnd cell_6t
Xbit_r321_c92 bl[92] br[92] wl[321] vdd gnd cell_6t
Xbit_r322_c92 bl[92] br[92] wl[322] vdd gnd cell_6t
Xbit_r323_c92 bl[92] br[92] wl[323] vdd gnd cell_6t
Xbit_r324_c92 bl[92] br[92] wl[324] vdd gnd cell_6t
Xbit_r325_c92 bl[92] br[92] wl[325] vdd gnd cell_6t
Xbit_r326_c92 bl[92] br[92] wl[326] vdd gnd cell_6t
Xbit_r327_c92 bl[92] br[92] wl[327] vdd gnd cell_6t
Xbit_r328_c92 bl[92] br[92] wl[328] vdd gnd cell_6t
Xbit_r329_c92 bl[92] br[92] wl[329] vdd gnd cell_6t
Xbit_r330_c92 bl[92] br[92] wl[330] vdd gnd cell_6t
Xbit_r331_c92 bl[92] br[92] wl[331] vdd gnd cell_6t
Xbit_r332_c92 bl[92] br[92] wl[332] vdd gnd cell_6t
Xbit_r333_c92 bl[92] br[92] wl[333] vdd gnd cell_6t
Xbit_r334_c92 bl[92] br[92] wl[334] vdd gnd cell_6t
Xbit_r335_c92 bl[92] br[92] wl[335] vdd gnd cell_6t
Xbit_r336_c92 bl[92] br[92] wl[336] vdd gnd cell_6t
Xbit_r337_c92 bl[92] br[92] wl[337] vdd gnd cell_6t
Xbit_r338_c92 bl[92] br[92] wl[338] vdd gnd cell_6t
Xbit_r339_c92 bl[92] br[92] wl[339] vdd gnd cell_6t
Xbit_r340_c92 bl[92] br[92] wl[340] vdd gnd cell_6t
Xbit_r341_c92 bl[92] br[92] wl[341] vdd gnd cell_6t
Xbit_r342_c92 bl[92] br[92] wl[342] vdd gnd cell_6t
Xbit_r343_c92 bl[92] br[92] wl[343] vdd gnd cell_6t
Xbit_r344_c92 bl[92] br[92] wl[344] vdd gnd cell_6t
Xbit_r345_c92 bl[92] br[92] wl[345] vdd gnd cell_6t
Xbit_r346_c92 bl[92] br[92] wl[346] vdd gnd cell_6t
Xbit_r347_c92 bl[92] br[92] wl[347] vdd gnd cell_6t
Xbit_r348_c92 bl[92] br[92] wl[348] vdd gnd cell_6t
Xbit_r349_c92 bl[92] br[92] wl[349] vdd gnd cell_6t
Xbit_r350_c92 bl[92] br[92] wl[350] vdd gnd cell_6t
Xbit_r351_c92 bl[92] br[92] wl[351] vdd gnd cell_6t
Xbit_r352_c92 bl[92] br[92] wl[352] vdd gnd cell_6t
Xbit_r353_c92 bl[92] br[92] wl[353] vdd gnd cell_6t
Xbit_r354_c92 bl[92] br[92] wl[354] vdd gnd cell_6t
Xbit_r355_c92 bl[92] br[92] wl[355] vdd gnd cell_6t
Xbit_r356_c92 bl[92] br[92] wl[356] vdd gnd cell_6t
Xbit_r357_c92 bl[92] br[92] wl[357] vdd gnd cell_6t
Xbit_r358_c92 bl[92] br[92] wl[358] vdd gnd cell_6t
Xbit_r359_c92 bl[92] br[92] wl[359] vdd gnd cell_6t
Xbit_r360_c92 bl[92] br[92] wl[360] vdd gnd cell_6t
Xbit_r361_c92 bl[92] br[92] wl[361] vdd gnd cell_6t
Xbit_r362_c92 bl[92] br[92] wl[362] vdd gnd cell_6t
Xbit_r363_c92 bl[92] br[92] wl[363] vdd gnd cell_6t
Xbit_r364_c92 bl[92] br[92] wl[364] vdd gnd cell_6t
Xbit_r365_c92 bl[92] br[92] wl[365] vdd gnd cell_6t
Xbit_r366_c92 bl[92] br[92] wl[366] vdd gnd cell_6t
Xbit_r367_c92 bl[92] br[92] wl[367] vdd gnd cell_6t
Xbit_r368_c92 bl[92] br[92] wl[368] vdd gnd cell_6t
Xbit_r369_c92 bl[92] br[92] wl[369] vdd gnd cell_6t
Xbit_r370_c92 bl[92] br[92] wl[370] vdd gnd cell_6t
Xbit_r371_c92 bl[92] br[92] wl[371] vdd gnd cell_6t
Xbit_r372_c92 bl[92] br[92] wl[372] vdd gnd cell_6t
Xbit_r373_c92 bl[92] br[92] wl[373] vdd gnd cell_6t
Xbit_r374_c92 bl[92] br[92] wl[374] vdd gnd cell_6t
Xbit_r375_c92 bl[92] br[92] wl[375] vdd gnd cell_6t
Xbit_r376_c92 bl[92] br[92] wl[376] vdd gnd cell_6t
Xbit_r377_c92 bl[92] br[92] wl[377] vdd gnd cell_6t
Xbit_r378_c92 bl[92] br[92] wl[378] vdd gnd cell_6t
Xbit_r379_c92 bl[92] br[92] wl[379] vdd gnd cell_6t
Xbit_r380_c92 bl[92] br[92] wl[380] vdd gnd cell_6t
Xbit_r381_c92 bl[92] br[92] wl[381] vdd gnd cell_6t
Xbit_r382_c92 bl[92] br[92] wl[382] vdd gnd cell_6t
Xbit_r383_c92 bl[92] br[92] wl[383] vdd gnd cell_6t
Xbit_r384_c92 bl[92] br[92] wl[384] vdd gnd cell_6t
Xbit_r385_c92 bl[92] br[92] wl[385] vdd gnd cell_6t
Xbit_r386_c92 bl[92] br[92] wl[386] vdd gnd cell_6t
Xbit_r387_c92 bl[92] br[92] wl[387] vdd gnd cell_6t
Xbit_r388_c92 bl[92] br[92] wl[388] vdd gnd cell_6t
Xbit_r389_c92 bl[92] br[92] wl[389] vdd gnd cell_6t
Xbit_r390_c92 bl[92] br[92] wl[390] vdd gnd cell_6t
Xbit_r391_c92 bl[92] br[92] wl[391] vdd gnd cell_6t
Xbit_r392_c92 bl[92] br[92] wl[392] vdd gnd cell_6t
Xbit_r393_c92 bl[92] br[92] wl[393] vdd gnd cell_6t
Xbit_r394_c92 bl[92] br[92] wl[394] vdd gnd cell_6t
Xbit_r395_c92 bl[92] br[92] wl[395] vdd gnd cell_6t
Xbit_r396_c92 bl[92] br[92] wl[396] vdd gnd cell_6t
Xbit_r397_c92 bl[92] br[92] wl[397] vdd gnd cell_6t
Xbit_r398_c92 bl[92] br[92] wl[398] vdd gnd cell_6t
Xbit_r399_c92 bl[92] br[92] wl[399] vdd gnd cell_6t
Xbit_r400_c92 bl[92] br[92] wl[400] vdd gnd cell_6t
Xbit_r401_c92 bl[92] br[92] wl[401] vdd gnd cell_6t
Xbit_r402_c92 bl[92] br[92] wl[402] vdd gnd cell_6t
Xbit_r403_c92 bl[92] br[92] wl[403] vdd gnd cell_6t
Xbit_r404_c92 bl[92] br[92] wl[404] vdd gnd cell_6t
Xbit_r405_c92 bl[92] br[92] wl[405] vdd gnd cell_6t
Xbit_r406_c92 bl[92] br[92] wl[406] vdd gnd cell_6t
Xbit_r407_c92 bl[92] br[92] wl[407] vdd gnd cell_6t
Xbit_r408_c92 bl[92] br[92] wl[408] vdd gnd cell_6t
Xbit_r409_c92 bl[92] br[92] wl[409] vdd gnd cell_6t
Xbit_r410_c92 bl[92] br[92] wl[410] vdd gnd cell_6t
Xbit_r411_c92 bl[92] br[92] wl[411] vdd gnd cell_6t
Xbit_r412_c92 bl[92] br[92] wl[412] vdd gnd cell_6t
Xbit_r413_c92 bl[92] br[92] wl[413] vdd gnd cell_6t
Xbit_r414_c92 bl[92] br[92] wl[414] vdd gnd cell_6t
Xbit_r415_c92 bl[92] br[92] wl[415] vdd gnd cell_6t
Xbit_r416_c92 bl[92] br[92] wl[416] vdd gnd cell_6t
Xbit_r417_c92 bl[92] br[92] wl[417] vdd gnd cell_6t
Xbit_r418_c92 bl[92] br[92] wl[418] vdd gnd cell_6t
Xbit_r419_c92 bl[92] br[92] wl[419] vdd gnd cell_6t
Xbit_r420_c92 bl[92] br[92] wl[420] vdd gnd cell_6t
Xbit_r421_c92 bl[92] br[92] wl[421] vdd gnd cell_6t
Xbit_r422_c92 bl[92] br[92] wl[422] vdd gnd cell_6t
Xbit_r423_c92 bl[92] br[92] wl[423] vdd gnd cell_6t
Xbit_r424_c92 bl[92] br[92] wl[424] vdd gnd cell_6t
Xbit_r425_c92 bl[92] br[92] wl[425] vdd gnd cell_6t
Xbit_r426_c92 bl[92] br[92] wl[426] vdd gnd cell_6t
Xbit_r427_c92 bl[92] br[92] wl[427] vdd gnd cell_6t
Xbit_r428_c92 bl[92] br[92] wl[428] vdd gnd cell_6t
Xbit_r429_c92 bl[92] br[92] wl[429] vdd gnd cell_6t
Xbit_r430_c92 bl[92] br[92] wl[430] vdd gnd cell_6t
Xbit_r431_c92 bl[92] br[92] wl[431] vdd gnd cell_6t
Xbit_r432_c92 bl[92] br[92] wl[432] vdd gnd cell_6t
Xbit_r433_c92 bl[92] br[92] wl[433] vdd gnd cell_6t
Xbit_r434_c92 bl[92] br[92] wl[434] vdd gnd cell_6t
Xbit_r435_c92 bl[92] br[92] wl[435] vdd gnd cell_6t
Xbit_r436_c92 bl[92] br[92] wl[436] vdd gnd cell_6t
Xbit_r437_c92 bl[92] br[92] wl[437] vdd gnd cell_6t
Xbit_r438_c92 bl[92] br[92] wl[438] vdd gnd cell_6t
Xbit_r439_c92 bl[92] br[92] wl[439] vdd gnd cell_6t
Xbit_r440_c92 bl[92] br[92] wl[440] vdd gnd cell_6t
Xbit_r441_c92 bl[92] br[92] wl[441] vdd gnd cell_6t
Xbit_r442_c92 bl[92] br[92] wl[442] vdd gnd cell_6t
Xbit_r443_c92 bl[92] br[92] wl[443] vdd gnd cell_6t
Xbit_r444_c92 bl[92] br[92] wl[444] vdd gnd cell_6t
Xbit_r445_c92 bl[92] br[92] wl[445] vdd gnd cell_6t
Xbit_r446_c92 bl[92] br[92] wl[446] vdd gnd cell_6t
Xbit_r447_c92 bl[92] br[92] wl[447] vdd gnd cell_6t
Xbit_r448_c92 bl[92] br[92] wl[448] vdd gnd cell_6t
Xbit_r449_c92 bl[92] br[92] wl[449] vdd gnd cell_6t
Xbit_r450_c92 bl[92] br[92] wl[450] vdd gnd cell_6t
Xbit_r451_c92 bl[92] br[92] wl[451] vdd gnd cell_6t
Xbit_r452_c92 bl[92] br[92] wl[452] vdd gnd cell_6t
Xbit_r453_c92 bl[92] br[92] wl[453] vdd gnd cell_6t
Xbit_r454_c92 bl[92] br[92] wl[454] vdd gnd cell_6t
Xbit_r455_c92 bl[92] br[92] wl[455] vdd gnd cell_6t
Xbit_r456_c92 bl[92] br[92] wl[456] vdd gnd cell_6t
Xbit_r457_c92 bl[92] br[92] wl[457] vdd gnd cell_6t
Xbit_r458_c92 bl[92] br[92] wl[458] vdd gnd cell_6t
Xbit_r459_c92 bl[92] br[92] wl[459] vdd gnd cell_6t
Xbit_r460_c92 bl[92] br[92] wl[460] vdd gnd cell_6t
Xbit_r461_c92 bl[92] br[92] wl[461] vdd gnd cell_6t
Xbit_r462_c92 bl[92] br[92] wl[462] vdd gnd cell_6t
Xbit_r463_c92 bl[92] br[92] wl[463] vdd gnd cell_6t
Xbit_r464_c92 bl[92] br[92] wl[464] vdd gnd cell_6t
Xbit_r465_c92 bl[92] br[92] wl[465] vdd gnd cell_6t
Xbit_r466_c92 bl[92] br[92] wl[466] vdd gnd cell_6t
Xbit_r467_c92 bl[92] br[92] wl[467] vdd gnd cell_6t
Xbit_r468_c92 bl[92] br[92] wl[468] vdd gnd cell_6t
Xbit_r469_c92 bl[92] br[92] wl[469] vdd gnd cell_6t
Xbit_r470_c92 bl[92] br[92] wl[470] vdd gnd cell_6t
Xbit_r471_c92 bl[92] br[92] wl[471] vdd gnd cell_6t
Xbit_r472_c92 bl[92] br[92] wl[472] vdd gnd cell_6t
Xbit_r473_c92 bl[92] br[92] wl[473] vdd gnd cell_6t
Xbit_r474_c92 bl[92] br[92] wl[474] vdd gnd cell_6t
Xbit_r475_c92 bl[92] br[92] wl[475] vdd gnd cell_6t
Xbit_r476_c92 bl[92] br[92] wl[476] vdd gnd cell_6t
Xbit_r477_c92 bl[92] br[92] wl[477] vdd gnd cell_6t
Xbit_r478_c92 bl[92] br[92] wl[478] vdd gnd cell_6t
Xbit_r479_c92 bl[92] br[92] wl[479] vdd gnd cell_6t
Xbit_r480_c92 bl[92] br[92] wl[480] vdd gnd cell_6t
Xbit_r481_c92 bl[92] br[92] wl[481] vdd gnd cell_6t
Xbit_r482_c92 bl[92] br[92] wl[482] vdd gnd cell_6t
Xbit_r483_c92 bl[92] br[92] wl[483] vdd gnd cell_6t
Xbit_r484_c92 bl[92] br[92] wl[484] vdd gnd cell_6t
Xbit_r485_c92 bl[92] br[92] wl[485] vdd gnd cell_6t
Xbit_r486_c92 bl[92] br[92] wl[486] vdd gnd cell_6t
Xbit_r487_c92 bl[92] br[92] wl[487] vdd gnd cell_6t
Xbit_r488_c92 bl[92] br[92] wl[488] vdd gnd cell_6t
Xbit_r489_c92 bl[92] br[92] wl[489] vdd gnd cell_6t
Xbit_r490_c92 bl[92] br[92] wl[490] vdd gnd cell_6t
Xbit_r491_c92 bl[92] br[92] wl[491] vdd gnd cell_6t
Xbit_r492_c92 bl[92] br[92] wl[492] vdd gnd cell_6t
Xbit_r493_c92 bl[92] br[92] wl[493] vdd gnd cell_6t
Xbit_r494_c92 bl[92] br[92] wl[494] vdd gnd cell_6t
Xbit_r495_c92 bl[92] br[92] wl[495] vdd gnd cell_6t
Xbit_r496_c92 bl[92] br[92] wl[496] vdd gnd cell_6t
Xbit_r497_c92 bl[92] br[92] wl[497] vdd gnd cell_6t
Xbit_r498_c92 bl[92] br[92] wl[498] vdd gnd cell_6t
Xbit_r499_c92 bl[92] br[92] wl[499] vdd gnd cell_6t
Xbit_r500_c92 bl[92] br[92] wl[500] vdd gnd cell_6t
Xbit_r501_c92 bl[92] br[92] wl[501] vdd gnd cell_6t
Xbit_r502_c92 bl[92] br[92] wl[502] vdd gnd cell_6t
Xbit_r503_c92 bl[92] br[92] wl[503] vdd gnd cell_6t
Xbit_r504_c92 bl[92] br[92] wl[504] vdd gnd cell_6t
Xbit_r505_c92 bl[92] br[92] wl[505] vdd gnd cell_6t
Xbit_r506_c92 bl[92] br[92] wl[506] vdd gnd cell_6t
Xbit_r507_c92 bl[92] br[92] wl[507] vdd gnd cell_6t
Xbit_r508_c92 bl[92] br[92] wl[508] vdd gnd cell_6t
Xbit_r509_c92 bl[92] br[92] wl[509] vdd gnd cell_6t
Xbit_r510_c92 bl[92] br[92] wl[510] vdd gnd cell_6t
Xbit_r511_c92 bl[92] br[92] wl[511] vdd gnd cell_6t
Xbit_r0_c93 bl[93] br[93] wl[0] vdd gnd cell_6t
Xbit_r1_c93 bl[93] br[93] wl[1] vdd gnd cell_6t
Xbit_r2_c93 bl[93] br[93] wl[2] vdd gnd cell_6t
Xbit_r3_c93 bl[93] br[93] wl[3] vdd gnd cell_6t
Xbit_r4_c93 bl[93] br[93] wl[4] vdd gnd cell_6t
Xbit_r5_c93 bl[93] br[93] wl[5] vdd gnd cell_6t
Xbit_r6_c93 bl[93] br[93] wl[6] vdd gnd cell_6t
Xbit_r7_c93 bl[93] br[93] wl[7] vdd gnd cell_6t
Xbit_r8_c93 bl[93] br[93] wl[8] vdd gnd cell_6t
Xbit_r9_c93 bl[93] br[93] wl[9] vdd gnd cell_6t
Xbit_r10_c93 bl[93] br[93] wl[10] vdd gnd cell_6t
Xbit_r11_c93 bl[93] br[93] wl[11] vdd gnd cell_6t
Xbit_r12_c93 bl[93] br[93] wl[12] vdd gnd cell_6t
Xbit_r13_c93 bl[93] br[93] wl[13] vdd gnd cell_6t
Xbit_r14_c93 bl[93] br[93] wl[14] vdd gnd cell_6t
Xbit_r15_c93 bl[93] br[93] wl[15] vdd gnd cell_6t
Xbit_r16_c93 bl[93] br[93] wl[16] vdd gnd cell_6t
Xbit_r17_c93 bl[93] br[93] wl[17] vdd gnd cell_6t
Xbit_r18_c93 bl[93] br[93] wl[18] vdd gnd cell_6t
Xbit_r19_c93 bl[93] br[93] wl[19] vdd gnd cell_6t
Xbit_r20_c93 bl[93] br[93] wl[20] vdd gnd cell_6t
Xbit_r21_c93 bl[93] br[93] wl[21] vdd gnd cell_6t
Xbit_r22_c93 bl[93] br[93] wl[22] vdd gnd cell_6t
Xbit_r23_c93 bl[93] br[93] wl[23] vdd gnd cell_6t
Xbit_r24_c93 bl[93] br[93] wl[24] vdd gnd cell_6t
Xbit_r25_c93 bl[93] br[93] wl[25] vdd gnd cell_6t
Xbit_r26_c93 bl[93] br[93] wl[26] vdd gnd cell_6t
Xbit_r27_c93 bl[93] br[93] wl[27] vdd gnd cell_6t
Xbit_r28_c93 bl[93] br[93] wl[28] vdd gnd cell_6t
Xbit_r29_c93 bl[93] br[93] wl[29] vdd gnd cell_6t
Xbit_r30_c93 bl[93] br[93] wl[30] vdd gnd cell_6t
Xbit_r31_c93 bl[93] br[93] wl[31] vdd gnd cell_6t
Xbit_r32_c93 bl[93] br[93] wl[32] vdd gnd cell_6t
Xbit_r33_c93 bl[93] br[93] wl[33] vdd gnd cell_6t
Xbit_r34_c93 bl[93] br[93] wl[34] vdd gnd cell_6t
Xbit_r35_c93 bl[93] br[93] wl[35] vdd gnd cell_6t
Xbit_r36_c93 bl[93] br[93] wl[36] vdd gnd cell_6t
Xbit_r37_c93 bl[93] br[93] wl[37] vdd gnd cell_6t
Xbit_r38_c93 bl[93] br[93] wl[38] vdd gnd cell_6t
Xbit_r39_c93 bl[93] br[93] wl[39] vdd gnd cell_6t
Xbit_r40_c93 bl[93] br[93] wl[40] vdd gnd cell_6t
Xbit_r41_c93 bl[93] br[93] wl[41] vdd gnd cell_6t
Xbit_r42_c93 bl[93] br[93] wl[42] vdd gnd cell_6t
Xbit_r43_c93 bl[93] br[93] wl[43] vdd gnd cell_6t
Xbit_r44_c93 bl[93] br[93] wl[44] vdd gnd cell_6t
Xbit_r45_c93 bl[93] br[93] wl[45] vdd gnd cell_6t
Xbit_r46_c93 bl[93] br[93] wl[46] vdd gnd cell_6t
Xbit_r47_c93 bl[93] br[93] wl[47] vdd gnd cell_6t
Xbit_r48_c93 bl[93] br[93] wl[48] vdd gnd cell_6t
Xbit_r49_c93 bl[93] br[93] wl[49] vdd gnd cell_6t
Xbit_r50_c93 bl[93] br[93] wl[50] vdd gnd cell_6t
Xbit_r51_c93 bl[93] br[93] wl[51] vdd gnd cell_6t
Xbit_r52_c93 bl[93] br[93] wl[52] vdd gnd cell_6t
Xbit_r53_c93 bl[93] br[93] wl[53] vdd gnd cell_6t
Xbit_r54_c93 bl[93] br[93] wl[54] vdd gnd cell_6t
Xbit_r55_c93 bl[93] br[93] wl[55] vdd gnd cell_6t
Xbit_r56_c93 bl[93] br[93] wl[56] vdd gnd cell_6t
Xbit_r57_c93 bl[93] br[93] wl[57] vdd gnd cell_6t
Xbit_r58_c93 bl[93] br[93] wl[58] vdd gnd cell_6t
Xbit_r59_c93 bl[93] br[93] wl[59] vdd gnd cell_6t
Xbit_r60_c93 bl[93] br[93] wl[60] vdd gnd cell_6t
Xbit_r61_c93 bl[93] br[93] wl[61] vdd gnd cell_6t
Xbit_r62_c93 bl[93] br[93] wl[62] vdd gnd cell_6t
Xbit_r63_c93 bl[93] br[93] wl[63] vdd gnd cell_6t
Xbit_r64_c93 bl[93] br[93] wl[64] vdd gnd cell_6t
Xbit_r65_c93 bl[93] br[93] wl[65] vdd gnd cell_6t
Xbit_r66_c93 bl[93] br[93] wl[66] vdd gnd cell_6t
Xbit_r67_c93 bl[93] br[93] wl[67] vdd gnd cell_6t
Xbit_r68_c93 bl[93] br[93] wl[68] vdd gnd cell_6t
Xbit_r69_c93 bl[93] br[93] wl[69] vdd gnd cell_6t
Xbit_r70_c93 bl[93] br[93] wl[70] vdd gnd cell_6t
Xbit_r71_c93 bl[93] br[93] wl[71] vdd gnd cell_6t
Xbit_r72_c93 bl[93] br[93] wl[72] vdd gnd cell_6t
Xbit_r73_c93 bl[93] br[93] wl[73] vdd gnd cell_6t
Xbit_r74_c93 bl[93] br[93] wl[74] vdd gnd cell_6t
Xbit_r75_c93 bl[93] br[93] wl[75] vdd gnd cell_6t
Xbit_r76_c93 bl[93] br[93] wl[76] vdd gnd cell_6t
Xbit_r77_c93 bl[93] br[93] wl[77] vdd gnd cell_6t
Xbit_r78_c93 bl[93] br[93] wl[78] vdd gnd cell_6t
Xbit_r79_c93 bl[93] br[93] wl[79] vdd gnd cell_6t
Xbit_r80_c93 bl[93] br[93] wl[80] vdd gnd cell_6t
Xbit_r81_c93 bl[93] br[93] wl[81] vdd gnd cell_6t
Xbit_r82_c93 bl[93] br[93] wl[82] vdd gnd cell_6t
Xbit_r83_c93 bl[93] br[93] wl[83] vdd gnd cell_6t
Xbit_r84_c93 bl[93] br[93] wl[84] vdd gnd cell_6t
Xbit_r85_c93 bl[93] br[93] wl[85] vdd gnd cell_6t
Xbit_r86_c93 bl[93] br[93] wl[86] vdd gnd cell_6t
Xbit_r87_c93 bl[93] br[93] wl[87] vdd gnd cell_6t
Xbit_r88_c93 bl[93] br[93] wl[88] vdd gnd cell_6t
Xbit_r89_c93 bl[93] br[93] wl[89] vdd gnd cell_6t
Xbit_r90_c93 bl[93] br[93] wl[90] vdd gnd cell_6t
Xbit_r91_c93 bl[93] br[93] wl[91] vdd gnd cell_6t
Xbit_r92_c93 bl[93] br[93] wl[92] vdd gnd cell_6t
Xbit_r93_c93 bl[93] br[93] wl[93] vdd gnd cell_6t
Xbit_r94_c93 bl[93] br[93] wl[94] vdd gnd cell_6t
Xbit_r95_c93 bl[93] br[93] wl[95] vdd gnd cell_6t
Xbit_r96_c93 bl[93] br[93] wl[96] vdd gnd cell_6t
Xbit_r97_c93 bl[93] br[93] wl[97] vdd gnd cell_6t
Xbit_r98_c93 bl[93] br[93] wl[98] vdd gnd cell_6t
Xbit_r99_c93 bl[93] br[93] wl[99] vdd gnd cell_6t
Xbit_r100_c93 bl[93] br[93] wl[100] vdd gnd cell_6t
Xbit_r101_c93 bl[93] br[93] wl[101] vdd gnd cell_6t
Xbit_r102_c93 bl[93] br[93] wl[102] vdd gnd cell_6t
Xbit_r103_c93 bl[93] br[93] wl[103] vdd gnd cell_6t
Xbit_r104_c93 bl[93] br[93] wl[104] vdd gnd cell_6t
Xbit_r105_c93 bl[93] br[93] wl[105] vdd gnd cell_6t
Xbit_r106_c93 bl[93] br[93] wl[106] vdd gnd cell_6t
Xbit_r107_c93 bl[93] br[93] wl[107] vdd gnd cell_6t
Xbit_r108_c93 bl[93] br[93] wl[108] vdd gnd cell_6t
Xbit_r109_c93 bl[93] br[93] wl[109] vdd gnd cell_6t
Xbit_r110_c93 bl[93] br[93] wl[110] vdd gnd cell_6t
Xbit_r111_c93 bl[93] br[93] wl[111] vdd gnd cell_6t
Xbit_r112_c93 bl[93] br[93] wl[112] vdd gnd cell_6t
Xbit_r113_c93 bl[93] br[93] wl[113] vdd gnd cell_6t
Xbit_r114_c93 bl[93] br[93] wl[114] vdd gnd cell_6t
Xbit_r115_c93 bl[93] br[93] wl[115] vdd gnd cell_6t
Xbit_r116_c93 bl[93] br[93] wl[116] vdd gnd cell_6t
Xbit_r117_c93 bl[93] br[93] wl[117] vdd gnd cell_6t
Xbit_r118_c93 bl[93] br[93] wl[118] vdd gnd cell_6t
Xbit_r119_c93 bl[93] br[93] wl[119] vdd gnd cell_6t
Xbit_r120_c93 bl[93] br[93] wl[120] vdd gnd cell_6t
Xbit_r121_c93 bl[93] br[93] wl[121] vdd gnd cell_6t
Xbit_r122_c93 bl[93] br[93] wl[122] vdd gnd cell_6t
Xbit_r123_c93 bl[93] br[93] wl[123] vdd gnd cell_6t
Xbit_r124_c93 bl[93] br[93] wl[124] vdd gnd cell_6t
Xbit_r125_c93 bl[93] br[93] wl[125] vdd gnd cell_6t
Xbit_r126_c93 bl[93] br[93] wl[126] vdd gnd cell_6t
Xbit_r127_c93 bl[93] br[93] wl[127] vdd gnd cell_6t
Xbit_r128_c93 bl[93] br[93] wl[128] vdd gnd cell_6t
Xbit_r129_c93 bl[93] br[93] wl[129] vdd gnd cell_6t
Xbit_r130_c93 bl[93] br[93] wl[130] vdd gnd cell_6t
Xbit_r131_c93 bl[93] br[93] wl[131] vdd gnd cell_6t
Xbit_r132_c93 bl[93] br[93] wl[132] vdd gnd cell_6t
Xbit_r133_c93 bl[93] br[93] wl[133] vdd gnd cell_6t
Xbit_r134_c93 bl[93] br[93] wl[134] vdd gnd cell_6t
Xbit_r135_c93 bl[93] br[93] wl[135] vdd gnd cell_6t
Xbit_r136_c93 bl[93] br[93] wl[136] vdd gnd cell_6t
Xbit_r137_c93 bl[93] br[93] wl[137] vdd gnd cell_6t
Xbit_r138_c93 bl[93] br[93] wl[138] vdd gnd cell_6t
Xbit_r139_c93 bl[93] br[93] wl[139] vdd gnd cell_6t
Xbit_r140_c93 bl[93] br[93] wl[140] vdd gnd cell_6t
Xbit_r141_c93 bl[93] br[93] wl[141] vdd gnd cell_6t
Xbit_r142_c93 bl[93] br[93] wl[142] vdd gnd cell_6t
Xbit_r143_c93 bl[93] br[93] wl[143] vdd gnd cell_6t
Xbit_r144_c93 bl[93] br[93] wl[144] vdd gnd cell_6t
Xbit_r145_c93 bl[93] br[93] wl[145] vdd gnd cell_6t
Xbit_r146_c93 bl[93] br[93] wl[146] vdd gnd cell_6t
Xbit_r147_c93 bl[93] br[93] wl[147] vdd gnd cell_6t
Xbit_r148_c93 bl[93] br[93] wl[148] vdd gnd cell_6t
Xbit_r149_c93 bl[93] br[93] wl[149] vdd gnd cell_6t
Xbit_r150_c93 bl[93] br[93] wl[150] vdd gnd cell_6t
Xbit_r151_c93 bl[93] br[93] wl[151] vdd gnd cell_6t
Xbit_r152_c93 bl[93] br[93] wl[152] vdd gnd cell_6t
Xbit_r153_c93 bl[93] br[93] wl[153] vdd gnd cell_6t
Xbit_r154_c93 bl[93] br[93] wl[154] vdd gnd cell_6t
Xbit_r155_c93 bl[93] br[93] wl[155] vdd gnd cell_6t
Xbit_r156_c93 bl[93] br[93] wl[156] vdd gnd cell_6t
Xbit_r157_c93 bl[93] br[93] wl[157] vdd gnd cell_6t
Xbit_r158_c93 bl[93] br[93] wl[158] vdd gnd cell_6t
Xbit_r159_c93 bl[93] br[93] wl[159] vdd gnd cell_6t
Xbit_r160_c93 bl[93] br[93] wl[160] vdd gnd cell_6t
Xbit_r161_c93 bl[93] br[93] wl[161] vdd gnd cell_6t
Xbit_r162_c93 bl[93] br[93] wl[162] vdd gnd cell_6t
Xbit_r163_c93 bl[93] br[93] wl[163] vdd gnd cell_6t
Xbit_r164_c93 bl[93] br[93] wl[164] vdd gnd cell_6t
Xbit_r165_c93 bl[93] br[93] wl[165] vdd gnd cell_6t
Xbit_r166_c93 bl[93] br[93] wl[166] vdd gnd cell_6t
Xbit_r167_c93 bl[93] br[93] wl[167] vdd gnd cell_6t
Xbit_r168_c93 bl[93] br[93] wl[168] vdd gnd cell_6t
Xbit_r169_c93 bl[93] br[93] wl[169] vdd gnd cell_6t
Xbit_r170_c93 bl[93] br[93] wl[170] vdd gnd cell_6t
Xbit_r171_c93 bl[93] br[93] wl[171] vdd gnd cell_6t
Xbit_r172_c93 bl[93] br[93] wl[172] vdd gnd cell_6t
Xbit_r173_c93 bl[93] br[93] wl[173] vdd gnd cell_6t
Xbit_r174_c93 bl[93] br[93] wl[174] vdd gnd cell_6t
Xbit_r175_c93 bl[93] br[93] wl[175] vdd gnd cell_6t
Xbit_r176_c93 bl[93] br[93] wl[176] vdd gnd cell_6t
Xbit_r177_c93 bl[93] br[93] wl[177] vdd gnd cell_6t
Xbit_r178_c93 bl[93] br[93] wl[178] vdd gnd cell_6t
Xbit_r179_c93 bl[93] br[93] wl[179] vdd gnd cell_6t
Xbit_r180_c93 bl[93] br[93] wl[180] vdd gnd cell_6t
Xbit_r181_c93 bl[93] br[93] wl[181] vdd gnd cell_6t
Xbit_r182_c93 bl[93] br[93] wl[182] vdd gnd cell_6t
Xbit_r183_c93 bl[93] br[93] wl[183] vdd gnd cell_6t
Xbit_r184_c93 bl[93] br[93] wl[184] vdd gnd cell_6t
Xbit_r185_c93 bl[93] br[93] wl[185] vdd gnd cell_6t
Xbit_r186_c93 bl[93] br[93] wl[186] vdd gnd cell_6t
Xbit_r187_c93 bl[93] br[93] wl[187] vdd gnd cell_6t
Xbit_r188_c93 bl[93] br[93] wl[188] vdd gnd cell_6t
Xbit_r189_c93 bl[93] br[93] wl[189] vdd gnd cell_6t
Xbit_r190_c93 bl[93] br[93] wl[190] vdd gnd cell_6t
Xbit_r191_c93 bl[93] br[93] wl[191] vdd gnd cell_6t
Xbit_r192_c93 bl[93] br[93] wl[192] vdd gnd cell_6t
Xbit_r193_c93 bl[93] br[93] wl[193] vdd gnd cell_6t
Xbit_r194_c93 bl[93] br[93] wl[194] vdd gnd cell_6t
Xbit_r195_c93 bl[93] br[93] wl[195] vdd gnd cell_6t
Xbit_r196_c93 bl[93] br[93] wl[196] vdd gnd cell_6t
Xbit_r197_c93 bl[93] br[93] wl[197] vdd gnd cell_6t
Xbit_r198_c93 bl[93] br[93] wl[198] vdd gnd cell_6t
Xbit_r199_c93 bl[93] br[93] wl[199] vdd gnd cell_6t
Xbit_r200_c93 bl[93] br[93] wl[200] vdd gnd cell_6t
Xbit_r201_c93 bl[93] br[93] wl[201] vdd gnd cell_6t
Xbit_r202_c93 bl[93] br[93] wl[202] vdd gnd cell_6t
Xbit_r203_c93 bl[93] br[93] wl[203] vdd gnd cell_6t
Xbit_r204_c93 bl[93] br[93] wl[204] vdd gnd cell_6t
Xbit_r205_c93 bl[93] br[93] wl[205] vdd gnd cell_6t
Xbit_r206_c93 bl[93] br[93] wl[206] vdd gnd cell_6t
Xbit_r207_c93 bl[93] br[93] wl[207] vdd gnd cell_6t
Xbit_r208_c93 bl[93] br[93] wl[208] vdd gnd cell_6t
Xbit_r209_c93 bl[93] br[93] wl[209] vdd gnd cell_6t
Xbit_r210_c93 bl[93] br[93] wl[210] vdd gnd cell_6t
Xbit_r211_c93 bl[93] br[93] wl[211] vdd gnd cell_6t
Xbit_r212_c93 bl[93] br[93] wl[212] vdd gnd cell_6t
Xbit_r213_c93 bl[93] br[93] wl[213] vdd gnd cell_6t
Xbit_r214_c93 bl[93] br[93] wl[214] vdd gnd cell_6t
Xbit_r215_c93 bl[93] br[93] wl[215] vdd gnd cell_6t
Xbit_r216_c93 bl[93] br[93] wl[216] vdd gnd cell_6t
Xbit_r217_c93 bl[93] br[93] wl[217] vdd gnd cell_6t
Xbit_r218_c93 bl[93] br[93] wl[218] vdd gnd cell_6t
Xbit_r219_c93 bl[93] br[93] wl[219] vdd gnd cell_6t
Xbit_r220_c93 bl[93] br[93] wl[220] vdd gnd cell_6t
Xbit_r221_c93 bl[93] br[93] wl[221] vdd gnd cell_6t
Xbit_r222_c93 bl[93] br[93] wl[222] vdd gnd cell_6t
Xbit_r223_c93 bl[93] br[93] wl[223] vdd gnd cell_6t
Xbit_r224_c93 bl[93] br[93] wl[224] vdd gnd cell_6t
Xbit_r225_c93 bl[93] br[93] wl[225] vdd gnd cell_6t
Xbit_r226_c93 bl[93] br[93] wl[226] vdd gnd cell_6t
Xbit_r227_c93 bl[93] br[93] wl[227] vdd gnd cell_6t
Xbit_r228_c93 bl[93] br[93] wl[228] vdd gnd cell_6t
Xbit_r229_c93 bl[93] br[93] wl[229] vdd gnd cell_6t
Xbit_r230_c93 bl[93] br[93] wl[230] vdd gnd cell_6t
Xbit_r231_c93 bl[93] br[93] wl[231] vdd gnd cell_6t
Xbit_r232_c93 bl[93] br[93] wl[232] vdd gnd cell_6t
Xbit_r233_c93 bl[93] br[93] wl[233] vdd gnd cell_6t
Xbit_r234_c93 bl[93] br[93] wl[234] vdd gnd cell_6t
Xbit_r235_c93 bl[93] br[93] wl[235] vdd gnd cell_6t
Xbit_r236_c93 bl[93] br[93] wl[236] vdd gnd cell_6t
Xbit_r237_c93 bl[93] br[93] wl[237] vdd gnd cell_6t
Xbit_r238_c93 bl[93] br[93] wl[238] vdd gnd cell_6t
Xbit_r239_c93 bl[93] br[93] wl[239] vdd gnd cell_6t
Xbit_r240_c93 bl[93] br[93] wl[240] vdd gnd cell_6t
Xbit_r241_c93 bl[93] br[93] wl[241] vdd gnd cell_6t
Xbit_r242_c93 bl[93] br[93] wl[242] vdd gnd cell_6t
Xbit_r243_c93 bl[93] br[93] wl[243] vdd gnd cell_6t
Xbit_r244_c93 bl[93] br[93] wl[244] vdd gnd cell_6t
Xbit_r245_c93 bl[93] br[93] wl[245] vdd gnd cell_6t
Xbit_r246_c93 bl[93] br[93] wl[246] vdd gnd cell_6t
Xbit_r247_c93 bl[93] br[93] wl[247] vdd gnd cell_6t
Xbit_r248_c93 bl[93] br[93] wl[248] vdd gnd cell_6t
Xbit_r249_c93 bl[93] br[93] wl[249] vdd gnd cell_6t
Xbit_r250_c93 bl[93] br[93] wl[250] vdd gnd cell_6t
Xbit_r251_c93 bl[93] br[93] wl[251] vdd gnd cell_6t
Xbit_r252_c93 bl[93] br[93] wl[252] vdd gnd cell_6t
Xbit_r253_c93 bl[93] br[93] wl[253] vdd gnd cell_6t
Xbit_r254_c93 bl[93] br[93] wl[254] vdd gnd cell_6t
Xbit_r255_c93 bl[93] br[93] wl[255] vdd gnd cell_6t
Xbit_r256_c93 bl[93] br[93] wl[256] vdd gnd cell_6t
Xbit_r257_c93 bl[93] br[93] wl[257] vdd gnd cell_6t
Xbit_r258_c93 bl[93] br[93] wl[258] vdd gnd cell_6t
Xbit_r259_c93 bl[93] br[93] wl[259] vdd gnd cell_6t
Xbit_r260_c93 bl[93] br[93] wl[260] vdd gnd cell_6t
Xbit_r261_c93 bl[93] br[93] wl[261] vdd gnd cell_6t
Xbit_r262_c93 bl[93] br[93] wl[262] vdd gnd cell_6t
Xbit_r263_c93 bl[93] br[93] wl[263] vdd gnd cell_6t
Xbit_r264_c93 bl[93] br[93] wl[264] vdd gnd cell_6t
Xbit_r265_c93 bl[93] br[93] wl[265] vdd gnd cell_6t
Xbit_r266_c93 bl[93] br[93] wl[266] vdd gnd cell_6t
Xbit_r267_c93 bl[93] br[93] wl[267] vdd gnd cell_6t
Xbit_r268_c93 bl[93] br[93] wl[268] vdd gnd cell_6t
Xbit_r269_c93 bl[93] br[93] wl[269] vdd gnd cell_6t
Xbit_r270_c93 bl[93] br[93] wl[270] vdd gnd cell_6t
Xbit_r271_c93 bl[93] br[93] wl[271] vdd gnd cell_6t
Xbit_r272_c93 bl[93] br[93] wl[272] vdd gnd cell_6t
Xbit_r273_c93 bl[93] br[93] wl[273] vdd gnd cell_6t
Xbit_r274_c93 bl[93] br[93] wl[274] vdd gnd cell_6t
Xbit_r275_c93 bl[93] br[93] wl[275] vdd gnd cell_6t
Xbit_r276_c93 bl[93] br[93] wl[276] vdd gnd cell_6t
Xbit_r277_c93 bl[93] br[93] wl[277] vdd gnd cell_6t
Xbit_r278_c93 bl[93] br[93] wl[278] vdd gnd cell_6t
Xbit_r279_c93 bl[93] br[93] wl[279] vdd gnd cell_6t
Xbit_r280_c93 bl[93] br[93] wl[280] vdd gnd cell_6t
Xbit_r281_c93 bl[93] br[93] wl[281] vdd gnd cell_6t
Xbit_r282_c93 bl[93] br[93] wl[282] vdd gnd cell_6t
Xbit_r283_c93 bl[93] br[93] wl[283] vdd gnd cell_6t
Xbit_r284_c93 bl[93] br[93] wl[284] vdd gnd cell_6t
Xbit_r285_c93 bl[93] br[93] wl[285] vdd gnd cell_6t
Xbit_r286_c93 bl[93] br[93] wl[286] vdd gnd cell_6t
Xbit_r287_c93 bl[93] br[93] wl[287] vdd gnd cell_6t
Xbit_r288_c93 bl[93] br[93] wl[288] vdd gnd cell_6t
Xbit_r289_c93 bl[93] br[93] wl[289] vdd gnd cell_6t
Xbit_r290_c93 bl[93] br[93] wl[290] vdd gnd cell_6t
Xbit_r291_c93 bl[93] br[93] wl[291] vdd gnd cell_6t
Xbit_r292_c93 bl[93] br[93] wl[292] vdd gnd cell_6t
Xbit_r293_c93 bl[93] br[93] wl[293] vdd gnd cell_6t
Xbit_r294_c93 bl[93] br[93] wl[294] vdd gnd cell_6t
Xbit_r295_c93 bl[93] br[93] wl[295] vdd gnd cell_6t
Xbit_r296_c93 bl[93] br[93] wl[296] vdd gnd cell_6t
Xbit_r297_c93 bl[93] br[93] wl[297] vdd gnd cell_6t
Xbit_r298_c93 bl[93] br[93] wl[298] vdd gnd cell_6t
Xbit_r299_c93 bl[93] br[93] wl[299] vdd gnd cell_6t
Xbit_r300_c93 bl[93] br[93] wl[300] vdd gnd cell_6t
Xbit_r301_c93 bl[93] br[93] wl[301] vdd gnd cell_6t
Xbit_r302_c93 bl[93] br[93] wl[302] vdd gnd cell_6t
Xbit_r303_c93 bl[93] br[93] wl[303] vdd gnd cell_6t
Xbit_r304_c93 bl[93] br[93] wl[304] vdd gnd cell_6t
Xbit_r305_c93 bl[93] br[93] wl[305] vdd gnd cell_6t
Xbit_r306_c93 bl[93] br[93] wl[306] vdd gnd cell_6t
Xbit_r307_c93 bl[93] br[93] wl[307] vdd gnd cell_6t
Xbit_r308_c93 bl[93] br[93] wl[308] vdd gnd cell_6t
Xbit_r309_c93 bl[93] br[93] wl[309] vdd gnd cell_6t
Xbit_r310_c93 bl[93] br[93] wl[310] vdd gnd cell_6t
Xbit_r311_c93 bl[93] br[93] wl[311] vdd gnd cell_6t
Xbit_r312_c93 bl[93] br[93] wl[312] vdd gnd cell_6t
Xbit_r313_c93 bl[93] br[93] wl[313] vdd gnd cell_6t
Xbit_r314_c93 bl[93] br[93] wl[314] vdd gnd cell_6t
Xbit_r315_c93 bl[93] br[93] wl[315] vdd gnd cell_6t
Xbit_r316_c93 bl[93] br[93] wl[316] vdd gnd cell_6t
Xbit_r317_c93 bl[93] br[93] wl[317] vdd gnd cell_6t
Xbit_r318_c93 bl[93] br[93] wl[318] vdd gnd cell_6t
Xbit_r319_c93 bl[93] br[93] wl[319] vdd gnd cell_6t
Xbit_r320_c93 bl[93] br[93] wl[320] vdd gnd cell_6t
Xbit_r321_c93 bl[93] br[93] wl[321] vdd gnd cell_6t
Xbit_r322_c93 bl[93] br[93] wl[322] vdd gnd cell_6t
Xbit_r323_c93 bl[93] br[93] wl[323] vdd gnd cell_6t
Xbit_r324_c93 bl[93] br[93] wl[324] vdd gnd cell_6t
Xbit_r325_c93 bl[93] br[93] wl[325] vdd gnd cell_6t
Xbit_r326_c93 bl[93] br[93] wl[326] vdd gnd cell_6t
Xbit_r327_c93 bl[93] br[93] wl[327] vdd gnd cell_6t
Xbit_r328_c93 bl[93] br[93] wl[328] vdd gnd cell_6t
Xbit_r329_c93 bl[93] br[93] wl[329] vdd gnd cell_6t
Xbit_r330_c93 bl[93] br[93] wl[330] vdd gnd cell_6t
Xbit_r331_c93 bl[93] br[93] wl[331] vdd gnd cell_6t
Xbit_r332_c93 bl[93] br[93] wl[332] vdd gnd cell_6t
Xbit_r333_c93 bl[93] br[93] wl[333] vdd gnd cell_6t
Xbit_r334_c93 bl[93] br[93] wl[334] vdd gnd cell_6t
Xbit_r335_c93 bl[93] br[93] wl[335] vdd gnd cell_6t
Xbit_r336_c93 bl[93] br[93] wl[336] vdd gnd cell_6t
Xbit_r337_c93 bl[93] br[93] wl[337] vdd gnd cell_6t
Xbit_r338_c93 bl[93] br[93] wl[338] vdd gnd cell_6t
Xbit_r339_c93 bl[93] br[93] wl[339] vdd gnd cell_6t
Xbit_r340_c93 bl[93] br[93] wl[340] vdd gnd cell_6t
Xbit_r341_c93 bl[93] br[93] wl[341] vdd gnd cell_6t
Xbit_r342_c93 bl[93] br[93] wl[342] vdd gnd cell_6t
Xbit_r343_c93 bl[93] br[93] wl[343] vdd gnd cell_6t
Xbit_r344_c93 bl[93] br[93] wl[344] vdd gnd cell_6t
Xbit_r345_c93 bl[93] br[93] wl[345] vdd gnd cell_6t
Xbit_r346_c93 bl[93] br[93] wl[346] vdd gnd cell_6t
Xbit_r347_c93 bl[93] br[93] wl[347] vdd gnd cell_6t
Xbit_r348_c93 bl[93] br[93] wl[348] vdd gnd cell_6t
Xbit_r349_c93 bl[93] br[93] wl[349] vdd gnd cell_6t
Xbit_r350_c93 bl[93] br[93] wl[350] vdd gnd cell_6t
Xbit_r351_c93 bl[93] br[93] wl[351] vdd gnd cell_6t
Xbit_r352_c93 bl[93] br[93] wl[352] vdd gnd cell_6t
Xbit_r353_c93 bl[93] br[93] wl[353] vdd gnd cell_6t
Xbit_r354_c93 bl[93] br[93] wl[354] vdd gnd cell_6t
Xbit_r355_c93 bl[93] br[93] wl[355] vdd gnd cell_6t
Xbit_r356_c93 bl[93] br[93] wl[356] vdd gnd cell_6t
Xbit_r357_c93 bl[93] br[93] wl[357] vdd gnd cell_6t
Xbit_r358_c93 bl[93] br[93] wl[358] vdd gnd cell_6t
Xbit_r359_c93 bl[93] br[93] wl[359] vdd gnd cell_6t
Xbit_r360_c93 bl[93] br[93] wl[360] vdd gnd cell_6t
Xbit_r361_c93 bl[93] br[93] wl[361] vdd gnd cell_6t
Xbit_r362_c93 bl[93] br[93] wl[362] vdd gnd cell_6t
Xbit_r363_c93 bl[93] br[93] wl[363] vdd gnd cell_6t
Xbit_r364_c93 bl[93] br[93] wl[364] vdd gnd cell_6t
Xbit_r365_c93 bl[93] br[93] wl[365] vdd gnd cell_6t
Xbit_r366_c93 bl[93] br[93] wl[366] vdd gnd cell_6t
Xbit_r367_c93 bl[93] br[93] wl[367] vdd gnd cell_6t
Xbit_r368_c93 bl[93] br[93] wl[368] vdd gnd cell_6t
Xbit_r369_c93 bl[93] br[93] wl[369] vdd gnd cell_6t
Xbit_r370_c93 bl[93] br[93] wl[370] vdd gnd cell_6t
Xbit_r371_c93 bl[93] br[93] wl[371] vdd gnd cell_6t
Xbit_r372_c93 bl[93] br[93] wl[372] vdd gnd cell_6t
Xbit_r373_c93 bl[93] br[93] wl[373] vdd gnd cell_6t
Xbit_r374_c93 bl[93] br[93] wl[374] vdd gnd cell_6t
Xbit_r375_c93 bl[93] br[93] wl[375] vdd gnd cell_6t
Xbit_r376_c93 bl[93] br[93] wl[376] vdd gnd cell_6t
Xbit_r377_c93 bl[93] br[93] wl[377] vdd gnd cell_6t
Xbit_r378_c93 bl[93] br[93] wl[378] vdd gnd cell_6t
Xbit_r379_c93 bl[93] br[93] wl[379] vdd gnd cell_6t
Xbit_r380_c93 bl[93] br[93] wl[380] vdd gnd cell_6t
Xbit_r381_c93 bl[93] br[93] wl[381] vdd gnd cell_6t
Xbit_r382_c93 bl[93] br[93] wl[382] vdd gnd cell_6t
Xbit_r383_c93 bl[93] br[93] wl[383] vdd gnd cell_6t
Xbit_r384_c93 bl[93] br[93] wl[384] vdd gnd cell_6t
Xbit_r385_c93 bl[93] br[93] wl[385] vdd gnd cell_6t
Xbit_r386_c93 bl[93] br[93] wl[386] vdd gnd cell_6t
Xbit_r387_c93 bl[93] br[93] wl[387] vdd gnd cell_6t
Xbit_r388_c93 bl[93] br[93] wl[388] vdd gnd cell_6t
Xbit_r389_c93 bl[93] br[93] wl[389] vdd gnd cell_6t
Xbit_r390_c93 bl[93] br[93] wl[390] vdd gnd cell_6t
Xbit_r391_c93 bl[93] br[93] wl[391] vdd gnd cell_6t
Xbit_r392_c93 bl[93] br[93] wl[392] vdd gnd cell_6t
Xbit_r393_c93 bl[93] br[93] wl[393] vdd gnd cell_6t
Xbit_r394_c93 bl[93] br[93] wl[394] vdd gnd cell_6t
Xbit_r395_c93 bl[93] br[93] wl[395] vdd gnd cell_6t
Xbit_r396_c93 bl[93] br[93] wl[396] vdd gnd cell_6t
Xbit_r397_c93 bl[93] br[93] wl[397] vdd gnd cell_6t
Xbit_r398_c93 bl[93] br[93] wl[398] vdd gnd cell_6t
Xbit_r399_c93 bl[93] br[93] wl[399] vdd gnd cell_6t
Xbit_r400_c93 bl[93] br[93] wl[400] vdd gnd cell_6t
Xbit_r401_c93 bl[93] br[93] wl[401] vdd gnd cell_6t
Xbit_r402_c93 bl[93] br[93] wl[402] vdd gnd cell_6t
Xbit_r403_c93 bl[93] br[93] wl[403] vdd gnd cell_6t
Xbit_r404_c93 bl[93] br[93] wl[404] vdd gnd cell_6t
Xbit_r405_c93 bl[93] br[93] wl[405] vdd gnd cell_6t
Xbit_r406_c93 bl[93] br[93] wl[406] vdd gnd cell_6t
Xbit_r407_c93 bl[93] br[93] wl[407] vdd gnd cell_6t
Xbit_r408_c93 bl[93] br[93] wl[408] vdd gnd cell_6t
Xbit_r409_c93 bl[93] br[93] wl[409] vdd gnd cell_6t
Xbit_r410_c93 bl[93] br[93] wl[410] vdd gnd cell_6t
Xbit_r411_c93 bl[93] br[93] wl[411] vdd gnd cell_6t
Xbit_r412_c93 bl[93] br[93] wl[412] vdd gnd cell_6t
Xbit_r413_c93 bl[93] br[93] wl[413] vdd gnd cell_6t
Xbit_r414_c93 bl[93] br[93] wl[414] vdd gnd cell_6t
Xbit_r415_c93 bl[93] br[93] wl[415] vdd gnd cell_6t
Xbit_r416_c93 bl[93] br[93] wl[416] vdd gnd cell_6t
Xbit_r417_c93 bl[93] br[93] wl[417] vdd gnd cell_6t
Xbit_r418_c93 bl[93] br[93] wl[418] vdd gnd cell_6t
Xbit_r419_c93 bl[93] br[93] wl[419] vdd gnd cell_6t
Xbit_r420_c93 bl[93] br[93] wl[420] vdd gnd cell_6t
Xbit_r421_c93 bl[93] br[93] wl[421] vdd gnd cell_6t
Xbit_r422_c93 bl[93] br[93] wl[422] vdd gnd cell_6t
Xbit_r423_c93 bl[93] br[93] wl[423] vdd gnd cell_6t
Xbit_r424_c93 bl[93] br[93] wl[424] vdd gnd cell_6t
Xbit_r425_c93 bl[93] br[93] wl[425] vdd gnd cell_6t
Xbit_r426_c93 bl[93] br[93] wl[426] vdd gnd cell_6t
Xbit_r427_c93 bl[93] br[93] wl[427] vdd gnd cell_6t
Xbit_r428_c93 bl[93] br[93] wl[428] vdd gnd cell_6t
Xbit_r429_c93 bl[93] br[93] wl[429] vdd gnd cell_6t
Xbit_r430_c93 bl[93] br[93] wl[430] vdd gnd cell_6t
Xbit_r431_c93 bl[93] br[93] wl[431] vdd gnd cell_6t
Xbit_r432_c93 bl[93] br[93] wl[432] vdd gnd cell_6t
Xbit_r433_c93 bl[93] br[93] wl[433] vdd gnd cell_6t
Xbit_r434_c93 bl[93] br[93] wl[434] vdd gnd cell_6t
Xbit_r435_c93 bl[93] br[93] wl[435] vdd gnd cell_6t
Xbit_r436_c93 bl[93] br[93] wl[436] vdd gnd cell_6t
Xbit_r437_c93 bl[93] br[93] wl[437] vdd gnd cell_6t
Xbit_r438_c93 bl[93] br[93] wl[438] vdd gnd cell_6t
Xbit_r439_c93 bl[93] br[93] wl[439] vdd gnd cell_6t
Xbit_r440_c93 bl[93] br[93] wl[440] vdd gnd cell_6t
Xbit_r441_c93 bl[93] br[93] wl[441] vdd gnd cell_6t
Xbit_r442_c93 bl[93] br[93] wl[442] vdd gnd cell_6t
Xbit_r443_c93 bl[93] br[93] wl[443] vdd gnd cell_6t
Xbit_r444_c93 bl[93] br[93] wl[444] vdd gnd cell_6t
Xbit_r445_c93 bl[93] br[93] wl[445] vdd gnd cell_6t
Xbit_r446_c93 bl[93] br[93] wl[446] vdd gnd cell_6t
Xbit_r447_c93 bl[93] br[93] wl[447] vdd gnd cell_6t
Xbit_r448_c93 bl[93] br[93] wl[448] vdd gnd cell_6t
Xbit_r449_c93 bl[93] br[93] wl[449] vdd gnd cell_6t
Xbit_r450_c93 bl[93] br[93] wl[450] vdd gnd cell_6t
Xbit_r451_c93 bl[93] br[93] wl[451] vdd gnd cell_6t
Xbit_r452_c93 bl[93] br[93] wl[452] vdd gnd cell_6t
Xbit_r453_c93 bl[93] br[93] wl[453] vdd gnd cell_6t
Xbit_r454_c93 bl[93] br[93] wl[454] vdd gnd cell_6t
Xbit_r455_c93 bl[93] br[93] wl[455] vdd gnd cell_6t
Xbit_r456_c93 bl[93] br[93] wl[456] vdd gnd cell_6t
Xbit_r457_c93 bl[93] br[93] wl[457] vdd gnd cell_6t
Xbit_r458_c93 bl[93] br[93] wl[458] vdd gnd cell_6t
Xbit_r459_c93 bl[93] br[93] wl[459] vdd gnd cell_6t
Xbit_r460_c93 bl[93] br[93] wl[460] vdd gnd cell_6t
Xbit_r461_c93 bl[93] br[93] wl[461] vdd gnd cell_6t
Xbit_r462_c93 bl[93] br[93] wl[462] vdd gnd cell_6t
Xbit_r463_c93 bl[93] br[93] wl[463] vdd gnd cell_6t
Xbit_r464_c93 bl[93] br[93] wl[464] vdd gnd cell_6t
Xbit_r465_c93 bl[93] br[93] wl[465] vdd gnd cell_6t
Xbit_r466_c93 bl[93] br[93] wl[466] vdd gnd cell_6t
Xbit_r467_c93 bl[93] br[93] wl[467] vdd gnd cell_6t
Xbit_r468_c93 bl[93] br[93] wl[468] vdd gnd cell_6t
Xbit_r469_c93 bl[93] br[93] wl[469] vdd gnd cell_6t
Xbit_r470_c93 bl[93] br[93] wl[470] vdd gnd cell_6t
Xbit_r471_c93 bl[93] br[93] wl[471] vdd gnd cell_6t
Xbit_r472_c93 bl[93] br[93] wl[472] vdd gnd cell_6t
Xbit_r473_c93 bl[93] br[93] wl[473] vdd gnd cell_6t
Xbit_r474_c93 bl[93] br[93] wl[474] vdd gnd cell_6t
Xbit_r475_c93 bl[93] br[93] wl[475] vdd gnd cell_6t
Xbit_r476_c93 bl[93] br[93] wl[476] vdd gnd cell_6t
Xbit_r477_c93 bl[93] br[93] wl[477] vdd gnd cell_6t
Xbit_r478_c93 bl[93] br[93] wl[478] vdd gnd cell_6t
Xbit_r479_c93 bl[93] br[93] wl[479] vdd gnd cell_6t
Xbit_r480_c93 bl[93] br[93] wl[480] vdd gnd cell_6t
Xbit_r481_c93 bl[93] br[93] wl[481] vdd gnd cell_6t
Xbit_r482_c93 bl[93] br[93] wl[482] vdd gnd cell_6t
Xbit_r483_c93 bl[93] br[93] wl[483] vdd gnd cell_6t
Xbit_r484_c93 bl[93] br[93] wl[484] vdd gnd cell_6t
Xbit_r485_c93 bl[93] br[93] wl[485] vdd gnd cell_6t
Xbit_r486_c93 bl[93] br[93] wl[486] vdd gnd cell_6t
Xbit_r487_c93 bl[93] br[93] wl[487] vdd gnd cell_6t
Xbit_r488_c93 bl[93] br[93] wl[488] vdd gnd cell_6t
Xbit_r489_c93 bl[93] br[93] wl[489] vdd gnd cell_6t
Xbit_r490_c93 bl[93] br[93] wl[490] vdd gnd cell_6t
Xbit_r491_c93 bl[93] br[93] wl[491] vdd gnd cell_6t
Xbit_r492_c93 bl[93] br[93] wl[492] vdd gnd cell_6t
Xbit_r493_c93 bl[93] br[93] wl[493] vdd gnd cell_6t
Xbit_r494_c93 bl[93] br[93] wl[494] vdd gnd cell_6t
Xbit_r495_c93 bl[93] br[93] wl[495] vdd gnd cell_6t
Xbit_r496_c93 bl[93] br[93] wl[496] vdd gnd cell_6t
Xbit_r497_c93 bl[93] br[93] wl[497] vdd gnd cell_6t
Xbit_r498_c93 bl[93] br[93] wl[498] vdd gnd cell_6t
Xbit_r499_c93 bl[93] br[93] wl[499] vdd gnd cell_6t
Xbit_r500_c93 bl[93] br[93] wl[500] vdd gnd cell_6t
Xbit_r501_c93 bl[93] br[93] wl[501] vdd gnd cell_6t
Xbit_r502_c93 bl[93] br[93] wl[502] vdd gnd cell_6t
Xbit_r503_c93 bl[93] br[93] wl[503] vdd gnd cell_6t
Xbit_r504_c93 bl[93] br[93] wl[504] vdd gnd cell_6t
Xbit_r505_c93 bl[93] br[93] wl[505] vdd gnd cell_6t
Xbit_r506_c93 bl[93] br[93] wl[506] vdd gnd cell_6t
Xbit_r507_c93 bl[93] br[93] wl[507] vdd gnd cell_6t
Xbit_r508_c93 bl[93] br[93] wl[508] vdd gnd cell_6t
Xbit_r509_c93 bl[93] br[93] wl[509] vdd gnd cell_6t
Xbit_r510_c93 bl[93] br[93] wl[510] vdd gnd cell_6t
Xbit_r511_c93 bl[93] br[93] wl[511] vdd gnd cell_6t
Xbit_r0_c94 bl[94] br[94] wl[0] vdd gnd cell_6t
Xbit_r1_c94 bl[94] br[94] wl[1] vdd gnd cell_6t
Xbit_r2_c94 bl[94] br[94] wl[2] vdd gnd cell_6t
Xbit_r3_c94 bl[94] br[94] wl[3] vdd gnd cell_6t
Xbit_r4_c94 bl[94] br[94] wl[4] vdd gnd cell_6t
Xbit_r5_c94 bl[94] br[94] wl[5] vdd gnd cell_6t
Xbit_r6_c94 bl[94] br[94] wl[6] vdd gnd cell_6t
Xbit_r7_c94 bl[94] br[94] wl[7] vdd gnd cell_6t
Xbit_r8_c94 bl[94] br[94] wl[8] vdd gnd cell_6t
Xbit_r9_c94 bl[94] br[94] wl[9] vdd gnd cell_6t
Xbit_r10_c94 bl[94] br[94] wl[10] vdd gnd cell_6t
Xbit_r11_c94 bl[94] br[94] wl[11] vdd gnd cell_6t
Xbit_r12_c94 bl[94] br[94] wl[12] vdd gnd cell_6t
Xbit_r13_c94 bl[94] br[94] wl[13] vdd gnd cell_6t
Xbit_r14_c94 bl[94] br[94] wl[14] vdd gnd cell_6t
Xbit_r15_c94 bl[94] br[94] wl[15] vdd gnd cell_6t
Xbit_r16_c94 bl[94] br[94] wl[16] vdd gnd cell_6t
Xbit_r17_c94 bl[94] br[94] wl[17] vdd gnd cell_6t
Xbit_r18_c94 bl[94] br[94] wl[18] vdd gnd cell_6t
Xbit_r19_c94 bl[94] br[94] wl[19] vdd gnd cell_6t
Xbit_r20_c94 bl[94] br[94] wl[20] vdd gnd cell_6t
Xbit_r21_c94 bl[94] br[94] wl[21] vdd gnd cell_6t
Xbit_r22_c94 bl[94] br[94] wl[22] vdd gnd cell_6t
Xbit_r23_c94 bl[94] br[94] wl[23] vdd gnd cell_6t
Xbit_r24_c94 bl[94] br[94] wl[24] vdd gnd cell_6t
Xbit_r25_c94 bl[94] br[94] wl[25] vdd gnd cell_6t
Xbit_r26_c94 bl[94] br[94] wl[26] vdd gnd cell_6t
Xbit_r27_c94 bl[94] br[94] wl[27] vdd gnd cell_6t
Xbit_r28_c94 bl[94] br[94] wl[28] vdd gnd cell_6t
Xbit_r29_c94 bl[94] br[94] wl[29] vdd gnd cell_6t
Xbit_r30_c94 bl[94] br[94] wl[30] vdd gnd cell_6t
Xbit_r31_c94 bl[94] br[94] wl[31] vdd gnd cell_6t
Xbit_r32_c94 bl[94] br[94] wl[32] vdd gnd cell_6t
Xbit_r33_c94 bl[94] br[94] wl[33] vdd gnd cell_6t
Xbit_r34_c94 bl[94] br[94] wl[34] vdd gnd cell_6t
Xbit_r35_c94 bl[94] br[94] wl[35] vdd gnd cell_6t
Xbit_r36_c94 bl[94] br[94] wl[36] vdd gnd cell_6t
Xbit_r37_c94 bl[94] br[94] wl[37] vdd gnd cell_6t
Xbit_r38_c94 bl[94] br[94] wl[38] vdd gnd cell_6t
Xbit_r39_c94 bl[94] br[94] wl[39] vdd gnd cell_6t
Xbit_r40_c94 bl[94] br[94] wl[40] vdd gnd cell_6t
Xbit_r41_c94 bl[94] br[94] wl[41] vdd gnd cell_6t
Xbit_r42_c94 bl[94] br[94] wl[42] vdd gnd cell_6t
Xbit_r43_c94 bl[94] br[94] wl[43] vdd gnd cell_6t
Xbit_r44_c94 bl[94] br[94] wl[44] vdd gnd cell_6t
Xbit_r45_c94 bl[94] br[94] wl[45] vdd gnd cell_6t
Xbit_r46_c94 bl[94] br[94] wl[46] vdd gnd cell_6t
Xbit_r47_c94 bl[94] br[94] wl[47] vdd gnd cell_6t
Xbit_r48_c94 bl[94] br[94] wl[48] vdd gnd cell_6t
Xbit_r49_c94 bl[94] br[94] wl[49] vdd gnd cell_6t
Xbit_r50_c94 bl[94] br[94] wl[50] vdd gnd cell_6t
Xbit_r51_c94 bl[94] br[94] wl[51] vdd gnd cell_6t
Xbit_r52_c94 bl[94] br[94] wl[52] vdd gnd cell_6t
Xbit_r53_c94 bl[94] br[94] wl[53] vdd gnd cell_6t
Xbit_r54_c94 bl[94] br[94] wl[54] vdd gnd cell_6t
Xbit_r55_c94 bl[94] br[94] wl[55] vdd gnd cell_6t
Xbit_r56_c94 bl[94] br[94] wl[56] vdd gnd cell_6t
Xbit_r57_c94 bl[94] br[94] wl[57] vdd gnd cell_6t
Xbit_r58_c94 bl[94] br[94] wl[58] vdd gnd cell_6t
Xbit_r59_c94 bl[94] br[94] wl[59] vdd gnd cell_6t
Xbit_r60_c94 bl[94] br[94] wl[60] vdd gnd cell_6t
Xbit_r61_c94 bl[94] br[94] wl[61] vdd gnd cell_6t
Xbit_r62_c94 bl[94] br[94] wl[62] vdd gnd cell_6t
Xbit_r63_c94 bl[94] br[94] wl[63] vdd gnd cell_6t
Xbit_r64_c94 bl[94] br[94] wl[64] vdd gnd cell_6t
Xbit_r65_c94 bl[94] br[94] wl[65] vdd gnd cell_6t
Xbit_r66_c94 bl[94] br[94] wl[66] vdd gnd cell_6t
Xbit_r67_c94 bl[94] br[94] wl[67] vdd gnd cell_6t
Xbit_r68_c94 bl[94] br[94] wl[68] vdd gnd cell_6t
Xbit_r69_c94 bl[94] br[94] wl[69] vdd gnd cell_6t
Xbit_r70_c94 bl[94] br[94] wl[70] vdd gnd cell_6t
Xbit_r71_c94 bl[94] br[94] wl[71] vdd gnd cell_6t
Xbit_r72_c94 bl[94] br[94] wl[72] vdd gnd cell_6t
Xbit_r73_c94 bl[94] br[94] wl[73] vdd gnd cell_6t
Xbit_r74_c94 bl[94] br[94] wl[74] vdd gnd cell_6t
Xbit_r75_c94 bl[94] br[94] wl[75] vdd gnd cell_6t
Xbit_r76_c94 bl[94] br[94] wl[76] vdd gnd cell_6t
Xbit_r77_c94 bl[94] br[94] wl[77] vdd gnd cell_6t
Xbit_r78_c94 bl[94] br[94] wl[78] vdd gnd cell_6t
Xbit_r79_c94 bl[94] br[94] wl[79] vdd gnd cell_6t
Xbit_r80_c94 bl[94] br[94] wl[80] vdd gnd cell_6t
Xbit_r81_c94 bl[94] br[94] wl[81] vdd gnd cell_6t
Xbit_r82_c94 bl[94] br[94] wl[82] vdd gnd cell_6t
Xbit_r83_c94 bl[94] br[94] wl[83] vdd gnd cell_6t
Xbit_r84_c94 bl[94] br[94] wl[84] vdd gnd cell_6t
Xbit_r85_c94 bl[94] br[94] wl[85] vdd gnd cell_6t
Xbit_r86_c94 bl[94] br[94] wl[86] vdd gnd cell_6t
Xbit_r87_c94 bl[94] br[94] wl[87] vdd gnd cell_6t
Xbit_r88_c94 bl[94] br[94] wl[88] vdd gnd cell_6t
Xbit_r89_c94 bl[94] br[94] wl[89] vdd gnd cell_6t
Xbit_r90_c94 bl[94] br[94] wl[90] vdd gnd cell_6t
Xbit_r91_c94 bl[94] br[94] wl[91] vdd gnd cell_6t
Xbit_r92_c94 bl[94] br[94] wl[92] vdd gnd cell_6t
Xbit_r93_c94 bl[94] br[94] wl[93] vdd gnd cell_6t
Xbit_r94_c94 bl[94] br[94] wl[94] vdd gnd cell_6t
Xbit_r95_c94 bl[94] br[94] wl[95] vdd gnd cell_6t
Xbit_r96_c94 bl[94] br[94] wl[96] vdd gnd cell_6t
Xbit_r97_c94 bl[94] br[94] wl[97] vdd gnd cell_6t
Xbit_r98_c94 bl[94] br[94] wl[98] vdd gnd cell_6t
Xbit_r99_c94 bl[94] br[94] wl[99] vdd gnd cell_6t
Xbit_r100_c94 bl[94] br[94] wl[100] vdd gnd cell_6t
Xbit_r101_c94 bl[94] br[94] wl[101] vdd gnd cell_6t
Xbit_r102_c94 bl[94] br[94] wl[102] vdd gnd cell_6t
Xbit_r103_c94 bl[94] br[94] wl[103] vdd gnd cell_6t
Xbit_r104_c94 bl[94] br[94] wl[104] vdd gnd cell_6t
Xbit_r105_c94 bl[94] br[94] wl[105] vdd gnd cell_6t
Xbit_r106_c94 bl[94] br[94] wl[106] vdd gnd cell_6t
Xbit_r107_c94 bl[94] br[94] wl[107] vdd gnd cell_6t
Xbit_r108_c94 bl[94] br[94] wl[108] vdd gnd cell_6t
Xbit_r109_c94 bl[94] br[94] wl[109] vdd gnd cell_6t
Xbit_r110_c94 bl[94] br[94] wl[110] vdd gnd cell_6t
Xbit_r111_c94 bl[94] br[94] wl[111] vdd gnd cell_6t
Xbit_r112_c94 bl[94] br[94] wl[112] vdd gnd cell_6t
Xbit_r113_c94 bl[94] br[94] wl[113] vdd gnd cell_6t
Xbit_r114_c94 bl[94] br[94] wl[114] vdd gnd cell_6t
Xbit_r115_c94 bl[94] br[94] wl[115] vdd gnd cell_6t
Xbit_r116_c94 bl[94] br[94] wl[116] vdd gnd cell_6t
Xbit_r117_c94 bl[94] br[94] wl[117] vdd gnd cell_6t
Xbit_r118_c94 bl[94] br[94] wl[118] vdd gnd cell_6t
Xbit_r119_c94 bl[94] br[94] wl[119] vdd gnd cell_6t
Xbit_r120_c94 bl[94] br[94] wl[120] vdd gnd cell_6t
Xbit_r121_c94 bl[94] br[94] wl[121] vdd gnd cell_6t
Xbit_r122_c94 bl[94] br[94] wl[122] vdd gnd cell_6t
Xbit_r123_c94 bl[94] br[94] wl[123] vdd gnd cell_6t
Xbit_r124_c94 bl[94] br[94] wl[124] vdd gnd cell_6t
Xbit_r125_c94 bl[94] br[94] wl[125] vdd gnd cell_6t
Xbit_r126_c94 bl[94] br[94] wl[126] vdd gnd cell_6t
Xbit_r127_c94 bl[94] br[94] wl[127] vdd gnd cell_6t
Xbit_r128_c94 bl[94] br[94] wl[128] vdd gnd cell_6t
Xbit_r129_c94 bl[94] br[94] wl[129] vdd gnd cell_6t
Xbit_r130_c94 bl[94] br[94] wl[130] vdd gnd cell_6t
Xbit_r131_c94 bl[94] br[94] wl[131] vdd gnd cell_6t
Xbit_r132_c94 bl[94] br[94] wl[132] vdd gnd cell_6t
Xbit_r133_c94 bl[94] br[94] wl[133] vdd gnd cell_6t
Xbit_r134_c94 bl[94] br[94] wl[134] vdd gnd cell_6t
Xbit_r135_c94 bl[94] br[94] wl[135] vdd gnd cell_6t
Xbit_r136_c94 bl[94] br[94] wl[136] vdd gnd cell_6t
Xbit_r137_c94 bl[94] br[94] wl[137] vdd gnd cell_6t
Xbit_r138_c94 bl[94] br[94] wl[138] vdd gnd cell_6t
Xbit_r139_c94 bl[94] br[94] wl[139] vdd gnd cell_6t
Xbit_r140_c94 bl[94] br[94] wl[140] vdd gnd cell_6t
Xbit_r141_c94 bl[94] br[94] wl[141] vdd gnd cell_6t
Xbit_r142_c94 bl[94] br[94] wl[142] vdd gnd cell_6t
Xbit_r143_c94 bl[94] br[94] wl[143] vdd gnd cell_6t
Xbit_r144_c94 bl[94] br[94] wl[144] vdd gnd cell_6t
Xbit_r145_c94 bl[94] br[94] wl[145] vdd gnd cell_6t
Xbit_r146_c94 bl[94] br[94] wl[146] vdd gnd cell_6t
Xbit_r147_c94 bl[94] br[94] wl[147] vdd gnd cell_6t
Xbit_r148_c94 bl[94] br[94] wl[148] vdd gnd cell_6t
Xbit_r149_c94 bl[94] br[94] wl[149] vdd gnd cell_6t
Xbit_r150_c94 bl[94] br[94] wl[150] vdd gnd cell_6t
Xbit_r151_c94 bl[94] br[94] wl[151] vdd gnd cell_6t
Xbit_r152_c94 bl[94] br[94] wl[152] vdd gnd cell_6t
Xbit_r153_c94 bl[94] br[94] wl[153] vdd gnd cell_6t
Xbit_r154_c94 bl[94] br[94] wl[154] vdd gnd cell_6t
Xbit_r155_c94 bl[94] br[94] wl[155] vdd gnd cell_6t
Xbit_r156_c94 bl[94] br[94] wl[156] vdd gnd cell_6t
Xbit_r157_c94 bl[94] br[94] wl[157] vdd gnd cell_6t
Xbit_r158_c94 bl[94] br[94] wl[158] vdd gnd cell_6t
Xbit_r159_c94 bl[94] br[94] wl[159] vdd gnd cell_6t
Xbit_r160_c94 bl[94] br[94] wl[160] vdd gnd cell_6t
Xbit_r161_c94 bl[94] br[94] wl[161] vdd gnd cell_6t
Xbit_r162_c94 bl[94] br[94] wl[162] vdd gnd cell_6t
Xbit_r163_c94 bl[94] br[94] wl[163] vdd gnd cell_6t
Xbit_r164_c94 bl[94] br[94] wl[164] vdd gnd cell_6t
Xbit_r165_c94 bl[94] br[94] wl[165] vdd gnd cell_6t
Xbit_r166_c94 bl[94] br[94] wl[166] vdd gnd cell_6t
Xbit_r167_c94 bl[94] br[94] wl[167] vdd gnd cell_6t
Xbit_r168_c94 bl[94] br[94] wl[168] vdd gnd cell_6t
Xbit_r169_c94 bl[94] br[94] wl[169] vdd gnd cell_6t
Xbit_r170_c94 bl[94] br[94] wl[170] vdd gnd cell_6t
Xbit_r171_c94 bl[94] br[94] wl[171] vdd gnd cell_6t
Xbit_r172_c94 bl[94] br[94] wl[172] vdd gnd cell_6t
Xbit_r173_c94 bl[94] br[94] wl[173] vdd gnd cell_6t
Xbit_r174_c94 bl[94] br[94] wl[174] vdd gnd cell_6t
Xbit_r175_c94 bl[94] br[94] wl[175] vdd gnd cell_6t
Xbit_r176_c94 bl[94] br[94] wl[176] vdd gnd cell_6t
Xbit_r177_c94 bl[94] br[94] wl[177] vdd gnd cell_6t
Xbit_r178_c94 bl[94] br[94] wl[178] vdd gnd cell_6t
Xbit_r179_c94 bl[94] br[94] wl[179] vdd gnd cell_6t
Xbit_r180_c94 bl[94] br[94] wl[180] vdd gnd cell_6t
Xbit_r181_c94 bl[94] br[94] wl[181] vdd gnd cell_6t
Xbit_r182_c94 bl[94] br[94] wl[182] vdd gnd cell_6t
Xbit_r183_c94 bl[94] br[94] wl[183] vdd gnd cell_6t
Xbit_r184_c94 bl[94] br[94] wl[184] vdd gnd cell_6t
Xbit_r185_c94 bl[94] br[94] wl[185] vdd gnd cell_6t
Xbit_r186_c94 bl[94] br[94] wl[186] vdd gnd cell_6t
Xbit_r187_c94 bl[94] br[94] wl[187] vdd gnd cell_6t
Xbit_r188_c94 bl[94] br[94] wl[188] vdd gnd cell_6t
Xbit_r189_c94 bl[94] br[94] wl[189] vdd gnd cell_6t
Xbit_r190_c94 bl[94] br[94] wl[190] vdd gnd cell_6t
Xbit_r191_c94 bl[94] br[94] wl[191] vdd gnd cell_6t
Xbit_r192_c94 bl[94] br[94] wl[192] vdd gnd cell_6t
Xbit_r193_c94 bl[94] br[94] wl[193] vdd gnd cell_6t
Xbit_r194_c94 bl[94] br[94] wl[194] vdd gnd cell_6t
Xbit_r195_c94 bl[94] br[94] wl[195] vdd gnd cell_6t
Xbit_r196_c94 bl[94] br[94] wl[196] vdd gnd cell_6t
Xbit_r197_c94 bl[94] br[94] wl[197] vdd gnd cell_6t
Xbit_r198_c94 bl[94] br[94] wl[198] vdd gnd cell_6t
Xbit_r199_c94 bl[94] br[94] wl[199] vdd gnd cell_6t
Xbit_r200_c94 bl[94] br[94] wl[200] vdd gnd cell_6t
Xbit_r201_c94 bl[94] br[94] wl[201] vdd gnd cell_6t
Xbit_r202_c94 bl[94] br[94] wl[202] vdd gnd cell_6t
Xbit_r203_c94 bl[94] br[94] wl[203] vdd gnd cell_6t
Xbit_r204_c94 bl[94] br[94] wl[204] vdd gnd cell_6t
Xbit_r205_c94 bl[94] br[94] wl[205] vdd gnd cell_6t
Xbit_r206_c94 bl[94] br[94] wl[206] vdd gnd cell_6t
Xbit_r207_c94 bl[94] br[94] wl[207] vdd gnd cell_6t
Xbit_r208_c94 bl[94] br[94] wl[208] vdd gnd cell_6t
Xbit_r209_c94 bl[94] br[94] wl[209] vdd gnd cell_6t
Xbit_r210_c94 bl[94] br[94] wl[210] vdd gnd cell_6t
Xbit_r211_c94 bl[94] br[94] wl[211] vdd gnd cell_6t
Xbit_r212_c94 bl[94] br[94] wl[212] vdd gnd cell_6t
Xbit_r213_c94 bl[94] br[94] wl[213] vdd gnd cell_6t
Xbit_r214_c94 bl[94] br[94] wl[214] vdd gnd cell_6t
Xbit_r215_c94 bl[94] br[94] wl[215] vdd gnd cell_6t
Xbit_r216_c94 bl[94] br[94] wl[216] vdd gnd cell_6t
Xbit_r217_c94 bl[94] br[94] wl[217] vdd gnd cell_6t
Xbit_r218_c94 bl[94] br[94] wl[218] vdd gnd cell_6t
Xbit_r219_c94 bl[94] br[94] wl[219] vdd gnd cell_6t
Xbit_r220_c94 bl[94] br[94] wl[220] vdd gnd cell_6t
Xbit_r221_c94 bl[94] br[94] wl[221] vdd gnd cell_6t
Xbit_r222_c94 bl[94] br[94] wl[222] vdd gnd cell_6t
Xbit_r223_c94 bl[94] br[94] wl[223] vdd gnd cell_6t
Xbit_r224_c94 bl[94] br[94] wl[224] vdd gnd cell_6t
Xbit_r225_c94 bl[94] br[94] wl[225] vdd gnd cell_6t
Xbit_r226_c94 bl[94] br[94] wl[226] vdd gnd cell_6t
Xbit_r227_c94 bl[94] br[94] wl[227] vdd gnd cell_6t
Xbit_r228_c94 bl[94] br[94] wl[228] vdd gnd cell_6t
Xbit_r229_c94 bl[94] br[94] wl[229] vdd gnd cell_6t
Xbit_r230_c94 bl[94] br[94] wl[230] vdd gnd cell_6t
Xbit_r231_c94 bl[94] br[94] wl[231] vdd gnd cell_6t
Xbit_r232_c94 bl[94] br[94] wl[232] vdd gnd cell_6t
Xbit_r233_c94 bl[94] br[94] wl[233] vdd gnd cell_6t
Xbit_r234_c94 bl[94] br[94] wl[234] vdd gnd cell_6t
Xbit_r235_c94 bl[94] br[94] wl[235] vdd gnd cell_6t
Xbit_r236_c94 bl[94] br[94] wl[236] vdd gnd cell_6t
Xbit_r237_c94 bl[94] br[94] wl[237] vdd gnd cell_6t
Xbit_r238_c94 bl[94] br[94] wl[238] vdd gnd cell_6t
Xbit_r239_c94 bl[94] br[94] wl[239] vdd gnd cell_6t
Xbit_r240_c94 bl[94] br[94] wl[240] vdd gnd cell_6t
Xbit_r241_c94 bl[94] br[94] wl[241] vdd gnd cell_6t
Xbit_r242_c94 bl[94] br[94] wl[242] vdd gnd cell_6t
Xbit_r243_c94 bl[94] br[94] wl[243] vdd gnd cell_6t
Xbit_r244_c94 bl[94] br[94] wl[244] vdd gnd cell_6t
Xbit_r245_c94 bl[94] br[94] wl[245] vdd gnd cell_6t
Xbit_r246_c94 bl[94] br[94] wl[246] vdd gnd cell_6t
Xbit_r247_c94 bl[94] br[94] wl[247] vdd gnd cell_6t
Xbit_r248_c94 bl[94] br[94] wl[248] vdd gnd cell_6t
Xbit_r249_c94 bl[94] br[94] wl[249] vdd gnd cell_6t
Xbit_r250_c94 bl[94] br[94] wl[250] vdd gnd cell_6t
Xbit_r251_c94 bl[94] br[94] wl[251] vdd gnd cell_6t
Xbit_r252_c94 bl[94] br[94] wl[252] vdd gnd cell_6t
Xbit_r253_c94 bl[94] br[94] wl[253] vdd gnd cell_6t
Xbit_r254_c94 bl[94] br[94] wl[254] vdd gnd cell_6t
Xbit_r255_c94 bl[94] br[94] wl[255] vdd gnd cell_6t
Xbit_r256_c94 bl[94] br[94] wl[256] vdd gnd cell_6t
Xbit_r257_c94 bl[94] br[94] wl[257] vdd gnd cell_6t
Xbit_r258_c94 bl[94] br[94] wl[258] vdd gnd cell_6t
Xbit_r259_c94 bl[94] br[94] wl[259] vdd gnd cell_6t
Xbit_r260_c94 bl[94] br[94] wl[260] vdd gnd cell_6t
Xbit_r261_c94 bl[94] br[94] wl[261] vdd gnd cell_6t
Xbit_r262_c94 bl[94] br[94] wl[262] vdd gnd cell_6t
Xbit_r263_c94 bl[94] br[94] wl[263] vdd gnd cell_6t
Xbit_r264_c94 bl[94] br[94] wl[264] vdd gnd cell_6t
Xbit_r265_c94 bl[94] br[94] wl[265] vdd gnd cell_6t
Xbit_r266_c94 bl[94] br[94] wl[266] vdd gnd cell_6t
Xbit_r267_c94 bl[94] br[94] wl[267] vdd gnd cell_6t
Xbit_r268_c94 bl[94] br[94] wl[268] vdd gnd cell_6t
Xbit_r269_c94 bl[94] br[94] wl[269] vdd gnd cell_6t
Xbit_r270_c94 bl[94] br[94] wl[270] vdd gnd cell_6t
Xbit_r271_c94 bl[94] br[94] wl[271] vdd gnd cell_6t
Xbit_r272_c94 bl[94] br[94] wl[272] vdd gnd cell_6t
Xbit_r273_c94 bl[94] br[94] wl[273] vdd gnd cell_6t
Xbit_r274_c94 bl[94] br[94] wl[274] vdd gnd cell_6t
Xbit_r275_c94 bl[94] br[94] wl[275] vdd gnd cell_6t
Xbit_r276_c94 bl[94] br[94] wl[276] vdd gnd cell_6t
Xbit_r277_c94 bl[94] br[94] wl[277] vdd gnd cell_6t
Xbit_r278_c94 bl[94] br[94] wl[278] vdd gnd cell_6t
Xbit_r279_c94 bl[94] br[94] wl[279] vdd gnd cell_6t
Xbit_r280_c94 bl[94] br[94] wl[280] vdd gnd cell_6t
Xbit_r281_c94 bl[94] br[94] wl[281] vdd gnd cell_6t
Xbit_r282_c94 bl[94] br[94] wl[282] vdd gnd cell_6t
Xbit_r283_c94 bl[94] br[94] wl[283] vdd gnd cell_6t
Xbit_r284_c94 bl[94] br[94] wl[284] vdd gnd cell_6t
Xbit_r285_c94 bl[94] br[94] wl[285] vdd gnd cell_6t
Xbit_r286_c94 bl[94] br[94] wl[286] vdd gnd cell_6t
Xbit_r287_c94 bl[94] br[94] wl[287] vdd gnd cell_6t
Xbit_r288_c94 bl[94] br[94] wl[288] vdd gnd cell_6t
Xbit_r289_c94 bl[94] br[94] wl[289] vdd gnd cell_6t
Xbit_r290_c94 bl[94] br[94] wl[290] vdd gnd cell_6t
Xbit_r291_c94 bl[94] br[94] wl[291] vdd gnd cell_6t
Xbit_r292_c94 bl[94] br[94] wl[292] vdd gnd cell_6t
Xbit_r293_c94 bl[94] br[94] wl[293] vdd gnd cell_6t
Xbit_r294_c94 bl[94] br[94] wl[294] vdd gnd cell_6t
Xbit_r295_c94 bl[94] br[94] wl[295] vdd gnd cell_6t
Xbit_r296_c94 bl[94] br[94] wl[296] vdd gnd cell_6t
Xbit_r297_c94 bl[94] br[94] wl[297] vdd gnd cell_6t
Xbit_r298_c94 bl[94] br[94] wl[298] vdd gnd cell_6t
Xbit_r299_c94 bl[94] br[94] wl[299] vdd gnd cell_6t
Xbit_r300_c94 bl[94] br[94] wl[300] vdd gnd cell_6t
Xbit_r301_c94 bl[94] br[94] wl[301] vdd gnd cell_6t
Xbit_r302_c94 bl[94] br[94] wl[302] vdd gnd cell_6t
Xbit_r303_c94 bl[94] br[94] wl[303] vdd gnd cell_6t
Xbit_r304_c94 bl[94] br[94] wl[304] vdd gnd cell_6t
Xbit_r305_c94 bl[94] br[94] wl[305] vdd gnd cell_6t
Xbit_r306_c94 bl[94] br[94] wl[306] vdd gnd cell_6t
Xbit_r307_c94 bl[94] br[94] wl[307] vdd gnd cell_6t
Xbit_r308_c94 bl[94] br[94] wl[308] vdd gnd cell_6t
Xbit_r309_c94 bl[94] br[94] wl[309] vdd gnd cell_6t
Xbit_r310_c94 bl[94] br[94] wl[310] vdd gnd cell_6t
Xbit_r311_c94 bl[94] br[94] wl[311] vdd gnd cell_6t
Xbit_r312_c94 bl[94] br[94] wl[312] vdd gnd cell_6t
Xbit_r313_c94 bl[94] br[94] wl[313] vdd gnd cell_6t
Xbit_r314_c94 bl[94] br[94] wl[314] vdd gnd cell_6t
Xbit_r315_c94 bl[94] br[94] wl[315] vdd gnd cell_6t
Xbit_r316_c94 bl[94] br[94] wl[316] vdd gnd cell_6t
Xbit_r317_c94 bl[94] br[94] wl[317] vdd gnd cell_6t
Xbit_r318_c94 bl[94] br[94] wl[318] vdd gnd cell_6t
Xbit_r319_c94 bl[94] br[94] wl[319] vdd gnd cell_6t
Xbit_r320_c94 bl[94] br[94] wl[320] vdd gnd cell_6t
Xbit_r321_c94 bl[94] br[94] wl[321] vdd gnd cell_6t
Xbit_r322_c94 bl[94] br[94] wl[322] vdd gnd cell_6t
Xbit_r323_c94 bl[94] br[94] wl[323] vdd gnd cell_6t
Xbit_r324_c94 bl[94] br[94] wl[324] vdd gnd cell_6t
Xbit_r325_c94 bl[94] br[94] wl[325] vdd gnd cell_6t
Xbit_r326_c94 bl[94] br[94] wl[326] vdd gnd cell_6t
Xbit_r327_c94 bl[94] br[94] wl[327] vdd gnd cell_6t
Xbit_r328_c94 bl[94] br[94] wl[328] vdd gnd cell_6t
Xbit_r329_c94 bl[94] br[94] wl[329] vdd gnd cell_6t
Xbit_r330_c94 bl[94] br[94] wl[330] vdd gnd cell_6t
Xbit_r331_c94 bl[94] br[94] wl[331] vdd gnd cell_6t
Xbit_r332_c94 bl[94] br[94] wl[332] vdd gnd cell_6t
Xbit_r333_c94 bl[94] br[94] wl[333] vdd gnd cell_6t
Xbit_r334_c94 bl[94] br[94] wl[334] vdd gnd cell_6t
Xbit_r335_c94 bl[94] br[94] wl[335] vdd gnd cell_6t
Xbit_r336_c94 bl[94] br[94] wl[336] vdd gnd cell_6t
Xbit_r337_c94 bl[94] br[94] wl[337] vdd gnd cell_6t
Xbit_r338_c94 bl[94] br[94] wl[338] vdd gnd cell_6t
Xbit_r339_c94 bl[94] br[94] wl[339] vdd gnd cell_6t
Xbit_r340_c94 bl[94] br[94] wl[340] vdd gnd cell_6t
Xbit_r341_c94 bl[94] br[94] wl[341] vdd gnd cell_6t
Xbit_r342_c94 bl[94] br[94] wl[342] vdd gnd cell_6t
Xbit_r343_c94 bl[94] br[94] wl[343] vdd gnd cell_6t
Xbit_r344_c94 bl[94] br[94] wl[344] vdd gnd cell_6t
Xbit_r345_c94 bl[94] br[94] wl[345] vdd gnd cell_6t
Xbit_r346_c94 bl[94] br[94] wl[346] vdd gnd cell_6t
Xbit_r347_c94 bl[94] br[94] wl[347] vdd gnd cell_6t
Xbit_r348_c94 bl[94] br[94] wl[348] vdd gnd cell_6t
Xbit_r349_c94 bl[94] br[94] wl[349] vdd gnd cell_6t
Xbit_r350_c94 bl[94] br[94] wl[350] vdd gnd cell_6t
Xbit_r351_c94 bl[94] br[94] wl[351] vdd gnd cell_6t
Xbit_r352_c94 bl[94] br[94] wl[352] vdd gnd cell_6t
Xbit_r353_c94 bl[94] br[94] wl[353] vdd gnd cell_6t
Xbit_r354_c94 bl[94] br[94] wl[354] vdd gnd cell_6t
Xbit_r355_c94 bl[94] br[94] wl[355] vdd gnd cell_6t
Xbit_r356_c94 bl[94] br[94] wl[356] vdd gnd cell_6t
Xbit_r357_c94 bl[94] br[94] wl[357] vdd gnd cell_6t
Xbit_r358_c94 bl[94] br[94] wl[358] vdd gnd cell_6t
Xbit_r359_c94 bl[94] br[94] wl[359] vdd gnd cell_6t
Xbit_r360_c94 bl[94] br[94] wl[360] vdd gnd cell_6t
Xbit_r361_c94 bl[94] br[94] wl[361] vdd gnd cell_6t
Xbit_r362_c94 bl[94] br[94] wl[362] vdd gnd cell_6t
Xbit_r363_c94 bl[94] br[94] wl[363] vdd gnd cell_6t
Xbit_r364_c94 bl[94] br[94] wl[364] vdd gnd cell_6t
Xbit_r365_c94 bl[94] br[94] wl[365] vdd gnd cell_6t
Xbit_r366_c94 bl[94] br[94] wl[366] vdd gnd cell_6t
Xbit_r367_c94 bl[94] br[94] wl[367] vdd gnd cell_6t
Xbit_r368_c94 bl[94] br[94] wl[368] vdd gnd cell_6t
Xbit_r369_c94 bl[94] br[94] wl[369] vdd gnd cell_6t
Xbit_r370_c94 bl[94] br[94] wl[370] vdd gnd cell_6t
Xbit_r371_c94 bl[94] br[94] wl[371] vdd gnd cell_6t
Xbit_r372_c94 bl[94] br[94] wl[372] vdd gnd cell_6t
Xbit_r373_c94 bl[94] br[94] wl[373] vdd gnd cell_6t
Xbit_r374_c94 bl[94] br[94] wl[374] vdd gnd cell_6t
Xbit_r375_c94 bl[94] br[94] wl[375] vdd gnd cell_6t
Xbit_r376_c94 bl[94] br[94] wl[376] vdd gnd cell_6t
Xbit_r377_c94 bl[94] br[94] wl[377] vdd gnd cell_6t
Xbit_r378_c94 bl[94] br[94] wl[378] vdd gnd cell_6t
Xbit_r379_c94 bl[94] br[94] wl[379] vdd gnd cell_6t
Xbit_r380_c94 bl[94] br[94] wl[380] vdd gnd cell_6t
Xbit_r381_c94 bl[94] br[94] wl[381] vdd gnd cell_6t
Xbit_r382_c94 bl[94] br[94] wl[382] vdd gnd cell_6t
Xbit_r383_c94 bl[94] br[94] wl[383] vdd gnd cell_6t
Xbit_r384_c94 bl[94] br[94] wl[384] vdd gnd cell_6t
Xbit_r385_c94 bl[94] br[94] wl[385] vdd gnd cell_6t
Xbit_r386_c94 bl[94] br[94] wl[386] vdd gnd cell_6t
Xbit_r387_c94 bl[94] br[94] wl[387] vdd gnd cell_6t
Xbit_r388_c94 bl[94] br[94] wl[388] vdd gnd cell_6t
Xbit_r389_c94 bl[94] br[94] wl[389] vdd gnd cell_6t
Xbit_r390_c94 bl[94] br[94] wl[390] vdd gnd cell_6t
Xbit_r391_c94 bl[94] br[94] wl[391] vdd gnd cell_6t
Xbit_r392_c94 bl[94] br[94] wl[392] vdd gnd cell_6t
Xbit_r393_c94 bl[94] br[94] wl[393] vdd gnd cell_6t
Xbit_r394_c94 bl[94] br[94] wl[394] vdd gnd cell_6t
Xbit_r395_c94 bl[94] br[94] wl[395] vdd gnd cell_6t
Xbit_r396_c94 bl[94] br[94] wl[396] vdd gnd cell_6t
Xbit_r397_c94 bl[94] br[94] wl[397] vdd gnd cell_6t
Xbit_r398_c94 bl[94] br[94] wl[398] vdd gnd cell_6t
Xbit_r399_c94 bl[94] br[94] wl[399] vdd gnd cell_6t
Xbit_r400_c94 bl[94] br[94] wl[400] vdd gnd cell_6t
Xbit_r401_c94 bl[94] br[94] wl[401] vdd gnd cell_6t
Xbit_r402_c94 bl[94] br[94] wl[402] vdd gnd cell_6t
Xbit_r403_c94 bl[94] br[94] wl[403] vdd gnd cell_6t
Xbit_r404_c94 bl[94] br[94] wl[404] vdd gnd cell_6t
Xbit_r405_c94 bl[94] br[94] wl[405] vdd gnd cell_6t
Xbit_r406_c94 bl[94] br[94] wl[406] vdd gnd cell_6t
Xbit_r407_c94 bl[94] br[94] wl[407] vdd gnd cell_6t
Xbit_r408_c94 bl[94] br[94] wl[408] vdd gnd cell_6t
Xbit_r409_c94 bl[94] br[94] wl[409] vdd gnd cell_6t
Xbit_r410_c94 bl[94] br[94] wl[410] vdd gnd cell_6t
Xbit_r411_c94 bl[94] br[94] wl[411] vdd gnd cell_6t
Xbit_r412_c94 bl[94] br[94] wl[412] vdd gnd cell_6t
Xbit_r413_c94 bl[94] br[94] wl[413] vdd gnd cell_6t
Xbit_r414_c94 bl[94] br[94] wl[414] vdd gnd cell_6t
Xbit_r415_c94 bl[94] br[94] wl[415] vdd gnd cell_6t
Xbit_r416_c94 bl[94] br[94] wl[416] vdd gnd cell_6t
Xbit_r417_c94 bl[94] br[94] wl[417] vdd gnd cell_6t
Xbit_r418_c94 bl[94] br[94] wl[418] vdd gnd cell_6t
Xbit_r419_c94 bl[94] br[94] wl[419] vdd gnd cell_6t
Xbit_r420_c94 bl[94] br[94] wl[420] vdd gnd cell_6t
Xbit_r421_c94 bl[94] br[94] wl[421] vdd gnd cell_6t
Xbit_r422_c94 bl[94] br[94] wl[422] vdd gnd cell_6t
Xbit_r423_c94 bl[94] br[94] wl[423] vdd gnd cell_6t
Xbit_r424_c94 bl[94] br[94] wl[424] vdd gnd cell_6t
Xbit_r425_c94 bl[94] br[94] wl[425] vdd gnd cell_6t
Xbit_r426_c94 bl[94] br[94] wl[426] vdd gnd cell_6t
Xbit_r427_c94 bl[94] br[94] wl[427] vdd gnd cell_6t
Xbit_r428_c94 bl[94] br[94] wl[428] vdd gnd cell_6t
Xbit_r429_c94 bl[94] br[94] wl[429] vdd gnd cell_6t
Xbit_r430_c94 bl[94] br[94] wl[430] vdd gnd cell_6t
Xbit_r431_c94 bl[94] br[94] wl[431] vdd gnd cell_6t
Xbit_r432_c94 bl[94] br[94] wl[432] vdd gnd cell_6t
Xbit_r433_c94 bl[94] br[94] wl[433] vdd gnd cell_6t
Xbit_r434_c94 bl[94] br[94] wl[434] vdd gnd cell_6t
Xbit_r435_c94 bl[94] br[94] wl[435] vdd gnd cell_6t
Xbit_r436_c94 bl[94] br[94] wl[436] vdd gnd cell_6t
Xbit_r437_c94 bl[94] br[94] wl[437] vdd gnd cell_6t
Xbit_r438_c94 bl[94] br[94] wl[438] vdd gnd cell_6t
Xbit_r439_c94 bl[94] br[94] wl[439] vdd gnd cell_6t
Xbit_r440_c94 bl[94] br[94] wl[440] vdd gnd cell_6t
Xbit_r441_c94 bl[94] br[94] wl[441] vdd gnd cell_6t
Xbit_r442_c94 bl[94] br[94] wl[442] vdd gnd cell_6t
Xbit_r443_c94 bl[94] br[94] wl[443] vdd gnd cell_6t
Xbit_r444_c94 bl[94] br[94] wl[444] vdd gnd cell_6t
Xbit_r445_c94 bl[94] br[94] wl[445] vdd gnd cell_6t
Xbit_r446_c94 bl[94] br[94] wl[446] vdd gnd cell_6t
Xbit_r447_c94 bl[94] br[94] wl[447] vdd gnd cell_6t
Xbit_r448_c94 bl[94] br[94] wl[448] vdd gnd cell_6t
Xbit_r449_c94 bl[94] br[94] wl[449] vdd gnd cell_6t
Xbit_r450_c94 bl[94] br[94] wl[450] vdd gnd cell_6t
Xbit_r451_c94 bl[94] br[94] wl[451] vdd gnd cell_6t
Xbit_r452_c94 bl[94] br[94] wl[452] vdd gnd cell_6t
Xbit_r453_c94 bl[94] br[94] wl[453] vdd gnd cell_6t
Xbit_r454_c94 bl[94] br[94] wl[454] vdd gnd cell_6t
Xbit_r455_c94 bl[94] br[94] wl[455] vdd gnd cell_6t
Xbit_r456_c94 bl[94] br[94] wl[456] vdd gnd cell_6t
Xbit_r457_c94 bl[94] br[94] wl[457] vdd gnd cell_6t
Xbit_r458_c94 bl[94] br[94] wl[458] vdd gnd cell_6t
Xbit_r459_c94 bl[94] br[94] wl[459] vdd gnd cell_6t
Xbit_r460_c94 bl[94] br[94] wl[460] vdd gnd cell_6t
Xbit_r461_c94 bl[94] br[94] wl[461] vdd gnd cell_6t
Xbit_r462_c94 bl[94] br[94] wl[462] vdd gnd cell_6t
Xbit_r463_c94 bl[94] br[94] wl[463] vdd gnd cell_6t
Xbit_r464_c94 bl[94] br[94] wl[464] vdd gnd cell_6t
Xbit_r465_c94 bl[94] br[94] wl[465] vdd gnd cell_6t
Xbit_r466_c94 bl[94] br[94] wl[466] vdd gnd cell_6t
Xbit_r467_c94 bl[94] br[94] wl[467] vdd gnd cell_6t
Xbit_r468_c94 bl[94] br[94] wl[468] vdd gnd cell_6t
Xbit_r469_c94 bl[94] br[94] wl[469] vdd gnd cell_6t
Xbit_r470_c94 bl[94] br[94] wl[470] vdd gnd cell_6t
Xbit_r471_c94 bl[94] br[94] wl[471] vdd gnd cell_6t
Xbit_r472_c94 bl[94] br[94] wl[472] vdd gnd cell_6t
Xbit_r473_c94 bl[94] br[94] wl[473] vdd gnd cell_6t
Xbit_r474_c94 bl[94] br[94] wl[474] vdd gnd cell_6t
Xbit_r475_c94 bl[94] br[94] wl[475] vdd gnd cell_6t
Xbit_r476_c94 bl[94] br[94] wl[476] vdd gnd cell_6t
Xbit_r477_c94 bl[94] br[94] wl[477] vdd gnd cell_6t
Xbit_r478_c94 bl[94] br[94] wl[478] vdd gnd cell_6t
Xbit_r479_c94 bl[94] br[94] wl[479] vdd gnd cell_6t
Xbit_r480_c94 bl[94] br[94] wl[480] vdd gnd cell_6t
Xbit_r481_c94 bl[94] br[94] wl[481] vdd gnd cell_6t
Xbit_r482_c94 bl[94] br[94] wl[482] vdd gnd cell_6t
Xbit_r483_c94 bl[94] br[94] wl[483] vdd gnd cell_6t
Xbit_r484_c94 bl[94] br[94] wl[484] vdd gnd cell_6t
Xbit_r485_c94 bl[94] br[94] wl[485] vdd gnd cell_6t
Xbit_r486_c94 bl[94] br[94] wl[486] vdd gnd cell_6t
Xbit_r487_c94 bl[94] br[94] wl[487] vdd gnd cell_6t
Xbit_r488_c94 bl[94] br[94] wl[488] vdd gnd cell_6t
Xbit_r489_c94 bl[94] br[94] wl[489] vdd gnd cell_6t
Xbit_r490_c94 bl[94] br[94] wl[490] vdd gnd cell_6t
Xbit_r491_c94 bl[94] br[94] wl[491] vdd gnd cell_6t
Xbit_r492_c94 bl[94] br[94] wl[492] vdd gnd cell_6t
Xbit_r493_c94 bl[94] br[94] wl[493] vdd gnd cell_6t
Xbit_r494_c94 bl[94] br[94] wl[494] vdd gnd cell_6t
Xbit_r495_c94 bl[94] br[94] wl[495] vdd gnd cell_6t
Xbit_r496_c94 bl[94] br[94] wl[496] vdd gnd cell_6t
Xbit_r497_c94 bl[94] br[94] wl[497] vdd gnd cell_6t
Xbit_r498_c94 bl[94] br[94] wl[498] vdd gnd cell_6t
Xbit_r499_c94 bl[94] br[94] wl[499] vdd gnd cell_6t
Xbit_r500_c94 bl[94] br[94] wl[500] vdd gnd cell_6t
Xbit_r501_c94 bl[94] br[94] wl[501] vdd gnd cell_6t
Xbit_r502_c94 bl[94] br[94] wl[502] vdd gnd cell_6t
Xbit_r503_c94 bl[94] br[94] wl[503] vdd gnd cell_6t
Xbit_r504_c94 bl[94] br[94] wl[504] vdd gnd cell_6t
Xbit_r505_c94 bl[94] br[94] wl[505] vdd gnd cell_6t
Xbit_r506_c94 bl[94] br[94] wl[506] vdd gnd cell_6t
Xbit_r507_c94 bl[94] br[94] wl[507] vdd gnd cell_6t
Xbit_r508_c94 bl[94] br[94] wl[508] vdd gnd cell_6t
Xbit_r509_c94 bl[94] br[94] wl[509] vdd gnd cell_6t
Xbit_r510_c94 bl[94] br[94] wl[510] vdd gnd cell_6t
Xbit_r511_c94 bl[94] br[94] wl[511] vdd gnd cell_6t
Xbit_r0_c95 bl[95] br[95] wl[0] vdd gnd cell_6t
Xbit_r1_c95 bl[95] br[95] wl[1] vdd gnd cell_6t
Xbit_r2_c95 bl[95] br[95] wl[2] vdd gnd cell_6t
Xbit_r3_c95 bl[95] br[95] wl[3] vdd gnd cell_6t
Xbit_r4_c95 bl[95] br[95] wl[4] vdd gnd cell_6t
Xbit_r5_c95 bl[95] br[95] wl[5] vdd gnd cell_6t
Xbit_r6_c95 bl[95] br[95] wl[6] vdd gnd cell_6t
Xbit_r7_c95 bl[95] br[95] wl[7] vdd gnd cell_6t
Xbit_r8_c95 bl[95] br[95] wl[8] vdd gnd cell_6t
Xbit_r9_c95 bl[95] br[95] wl[9] vdd gnd cell_6t
Xbit_r10_c95 bl[95] br[95] wl[10] vdd gnd cell_6t
Xbit_r11_c95 bl[95] br[95] wl[11] vdd gnd cell_6t
Xbit_r12_c95 bl[95] br[95] wl[12] vdd gnd cell_6t
Xbit_r13_c95 bl[95] br[95] wl[13] vdd gnd cell_6t
Xbit_r14_c95 bl[95] br[95] wl[14] vdd gnd cell_6t
Xbit_r15_c95 bl[95] br[95] wl[15] vdd gnd cell_6t
Xbit_r16_c95 bl[95] br[95] wl[16] vdd gnd cell_6t
Xbit_r17_c95 bl[95] br[95] wl[17] vdd gnd cell_6t
Xbit_r18_c95 bl[95] br[95] wl[18] vdd gnd cell_6t
Xbit_r19_c95 bl[95] br[95] wl[19] vdd gnd cell_6t
Xbit_r20_c95 bl[95] br[95] wl[20] vdd gnd cell_6t
Xbit_r21_c95 bl[95] br[95] wl[21] vdd gnd cell_6t
Xbit_r22_c95 bl[95] br[95] wl[22] vdd gnd cell_6t
Xbit_r23_c95 bl[95] br[95] wl[23] vdd gnd cell_6t
Xbit_r24_c95 bl[95] br[95] wl[24] vdd gnd cell_6t
Xbit_r25_c95 bl[95] br[95] wl[25] vdd gnd cell_6t
Xbit_r26_c95 bl[95] br[95] wl[26] vdd gnd cell_6t
Xbit_r27_c95 bl[95] br[95] wl[27] vdd gnd cell_6t
Xbit_r28_c95 bl[95] br[95] wl[28] vdd gnd cell_6t
Xbit_r29_c95 bl[95] br[95] wl[29] vdd gnd cell_6t
Xbit_r30_c95 bl[95] br[95] wl[30] vdd gnd cell_6t
Xbit_r31_c95 bl[95] br[95] wl[31] vdd gnd cell_6t
Xbit_r32_c95 bl[95] br[95] wl[32] vdd gnd cell_6t
Xbit_r33_c95 bl[95] br[95] wl[33] vdd gnd cell_6t
Xbit_r34_c95 bl[95] br[95] wl[34] vdd gnd cell_6t
Xbit_r35_c95 bl[95] br[95] wl[35] vdd gnd cell_6t
Xbit_r36_c95 bl[95] br[95] wl[36] vdd gnd cell_6t
Xbit_r37_c95 bl[95] br[95] wl[37] vdd gnd cell_6t
Xbit_r38_c95 bl[95] br[95] wl[38] vdd gnd cell_6t
Xbit_r39_c95 bl[95] br[95] wl[39] vdd gnd cell_6t
Xbit_r40_c95 bl[95] br[95] wl[40] vdd gnd cell_6t
Xbit_r41_c95 bl[95] br[95] wl[41] vdd gnd cell_6t
Xbit_r42_c95 bl[95] br[95] wl[42] vdd gnd cell_6t
Xbit_r43_c95 bl[95] br[95] wl[43] vdd gnd cell_6t
Xbit_r44_c95 bl[95] br[95] wl[44] vdd gnd cell_6t
Xbit_r45_c95 bl[95] br[95] wl[45] vdd gnd cell_6t
Xbit_r46_c95 bl[95] br[95] wl[46] vdd gnd cell_6t
Xbit_r47_c95 bl[95] br[95] wl[47] vdd gnd cell_6t
Xbit_r48_c95 bl[95] br[95] wl[48] vdd gnd cell_6t
Xbit_r49_c95 bl[95] br[95] wl[49] vdd gnd cell_6t
Xbit_r50_c95 bl[95] br[95] wl[50] vdd gnd cell_6t
Xbit_r51_c95 bl[95] br[95] wl[51] vdd gnd cell_6t
Xbit_r52_c95 bl[95] br[95] wl[52] vdd gnd cell_6t
Xbit_r53_c95 bl[95] br[95] wl[53] vdd gnd cell_6t
Xbit_r54_c95 bl[95] br[95] wl[54] vdd gnd cell_6t
Xbit_r55_c95 bl[95] br[95] wl[55] vdd gnd cell_6t
Xbit_r56_c95 bl[95] br[95] wl[56] vdd gnd cell_6t
Xbit_r57_c95 bl[95] br[95] wl[57] vdd gnd cell_6t
Xbit_r58_c95 bl[95] br[95] wl[58] vdd gnd cell_6t
Xbit_r59_c95 bl[95] br[95] wl[59] vdd gnd cell_6t
Xbit_r60_c95 bl[95] br[95] wl[60] vdd gnd cell_6t
Xbit_r61_c95 bl[95] br[95] wl[61] vdd gnd cell_6t
Xbit_r62_c95 bl[95] br[95] wl[62] vdd gnd cell_6t
Xbit_r63_c95 bl[95] br[95] wl[63] vdd gnd cell_6t
Xbit_r64_c95 bl[95] br[95] wl[64] vdd gnd cell_6t
Xbit_r65_c95 bl[95] br[95] wl[65] vdd gnd cell_6t
Xbit_r66_c95 bl[95] br[95] wl[66] vdd gnd cell_6t
Xbit_r67_c95 bl[95] br[95] wl[67] vdd gnd cell_6t
Xbit_r68_c95 bl[95] br[95] wl[68] vdd gnd cell_6t
Xbit_r69_c95 bl[95] br[95] wl[69] vdd gnd cell_6t
Xbit_r70_c95 bl[95] br[95] wl[70] vdd gnd cell_6t
Xbit_r71_c95 bl[95] br[95] wl[71] vdd gnd cell_6t
Xbit_r72_c95 bl[95] br[95] wl[72] vdd gnd cell_6t
Xbit_r73_c95 bl[95] br[95] wl[73] vdd gnd cell_6t
Xbit_r74_c95 bl[95] br[95] wl[74] vdd gnd cell_6t
Xbit_r75_c95 bl[95] br[95] wl[75] vdd gnd cell_6t
Xbit_r76_c95 bl[95] br[95] wl[76] vdd gnd cell_6t
Xbit_r77_c95 bl[95] br[95] wl[77] vdd gnd cell_6t
Xbit_r78_c95 bl[95] br[95] wl[78] vdd gnd cell_6t
Xbit_r79_c95 bl[95] br[95] wl[79] vdd gnd cell_6t
Xbit_r80_c95 bl[95] br[95] wl[80] vdd gnd cell_6t
Xbit_r81_c95 bl[95] br[95] wl[81] vdd gnd cell_6t
Xbit_r82_c95 bl[95] br[95] wl[82] vdd gnd cell_6t
Xbit_r83_c95 bl[95] br[95] wl[83] vdd gnd cell_6t
Xbit_r84_c95 bl[95] br[95] wl[84] vdd gnd cell_6t
Xbit_r85_c95 bl[95] br[95] wl[85] vdd gnd cell_6t
Xbit_r86_c95 bl[95] br[95] wl[86] vdd gnd cell_6t
Xbit_r87_c95 bl[95] br[95] wl[87] vdd gnd cell_6t
Xbit_r88_c95 bl[95] br[95] wl[88] vdd gnd cell_6t
Xbit_r89_c95 bl[95] br[95] wl[89] vdd gnd cell_6t
Xbit_r90_c95 bl[95] br[95] wl[90] vdd gnd cell_6t
Xbit_r91_c95 bl[95] br[95] wl[91] vdd gnd cell_6t
Xbit_r92_c95 bl[95] br[95] wl[92] vdd gnd cell_6t
Xbit_r93_c95 bl[95] br[95] wl[93] vdd gnd cell_6t
Xbit_r94_c95 bl[95] br[95] wl[94] vdd gnd cell_6t
Xbit_r95_c95 bl[95] br[95] wl[95] vdd gnd cell_6t
Xbit_r96_c95 bl[95] br[95] wl[96] vdd gnd cell_6t
Xbit_r97_c95 bl[95] br[95] wl[97] vdd gnd cell_6t
Xbit_r98_c95 bl[95] br[95] wl[98] vdd gnd cell_6t
Xbit_r99_c95 bl[95] br[95] wl[99] vdd gnd cell_6t
Xbit_r100_c95 bl[95] br[95] wl[100] vdd gnd cell_6t
Xbit_r101_c95 bl[95] br[95] wl[101] vdd gnd cell_6t
Xbit_r102_c95 bl[95] br[95] wl[102] vdd gnd cell_6t
Xbit_r103_c95 bl[95] br[95] wl[103] vdd gnd cell_6t
Xbit_r104_c95 bl[95] br[95] wl[104] vdd gnd cell_6t
Xbit_r105_c95 bl[95] br[95] wl[105] vdd gnd cell_6t
Xbit_r106_c95 bl[95] br[95] wl[106] vdd gnd cell_6t
Xbit_r107_c95 bl[95] br[95] wl[107] vdd gnd cell_6t
Xbit_r108_c95 bl[95] br[95] wl[108] vdd gnd cell_6t
Xbit_r109_c95 bl[95] br[95] wl[109] vdd gnd cell_6t
Xbit_r110_c95 bl[95] br[95] wl[110] vdd gnd cell_6t
Xbit_r111_c95 bl[95] br[95] wl[111] vdd gnd cell_6t
Xbit_r112_c95 bl[95] br[95] wl[112] vdd gnd cell_6t
Xbit_r113_c95 bl[95] br[95] wl[113] vdd gnd cell_6t
Xbit_r114_c95 bl[95] br[95] wl[114] vdd gnd cell_6t
Xbit_r115_c95 bl[95] br[95] wl[115] vdd gnd cell_6t
Xbit_r116_c95 bl[95] br[95] wl[116] vdd gnd cell_6t
Xbit_r117_c95 bl[95] br[95] wl[117] vdd gnd cell_6t
Xbit_r118_c95 bl[95] br[95] wl[118] vdd gnd cell_6t
Xbit_r119_c95 bl[95] br[95] wl[119] vdd gnd cell_6t
Xbit_r120_c95 bl[95] br[95] wl[120] vdd gnd cell_6t
Xbit_r121_c95 bl[95] br[95] wl[121] vdd gnd cell_6t
Xbit_r122_c95 bl[95] br[95] wl[122] vdd gnd cell_6t
Xbit_r123_c95 bl[95] br[95] wl[123] vdd gnd cell_6t
Xbit_r124_c95 bl[95] br[95] wl[124] vdd gnd cell_6t
Xbit_r125_c95 bl[95] br[95] wl[125] vdd gnd cell_6t
Xbit_r126_c95 bl[95] br[95] wl[126] vdd gnd cell_6t
Xbit_r127_c95 bl[95] br[95] wl[127] vdd gnd cell_6t
Xbit_r128_c95 bl[95] br[95] wl[128] vdd gnd cell_6t
Xbit_r129_c95 bl[95] br[95] wl[129] vdd gnd cell_6t
Xbit_r130_c95 bl[95] br[95] wl[130] vdd gnd cell_6t
Xbit_r131_c95 bl[95] br[95] wl[131] vdd gnd cell_6t
Xbit_r132_c95 bl[95] br[95] wl[132] vdd gnd cell_6t
Xbit_r133_c95 bl[95] br[95] wl[133] vdd gnd cell_6t
Xbit_r134_c95 bl[95] br[95] wl[134] vdd gnd cell_6t
Xbit_r135_c95 bl[95] br[95] wl[135] vdd gnd cell_6t
Xbit_r136_c95 bl[95] br[95] wl[136] vdd gnd cell_6t
Xbit_r137_c95 bl[95] br[95] wl[137] vdd gnd cell_6t
Xbit_r138_c95 bl[95] br[95] wl[138] vdd gnd cell_6t
Xbit_r139_c95 bl[95] br[95] wl[139] vdd gnd cell_6t
Xbit_r140_c95 bl[95] br[95] wl[140] vdd gnd cell_6t
Xbit_r141_c95 bl[95] br[95] wl[141] vdd gnd cell_6t
Xbit_r142_c95 bl[95] br[95] wl[142] vdd gnd cell_6t
Xbit_r143_c95 bl[95] br[95] wl[143] vdd gnd cell_6t
Xbit_r144_c95 bl[95] br[95] wl[144] vdd gnd cell_6t
Xbit_r145_c95 bl[95] br[95] wl[145] vdd gnd cell_6t
Xbit_r146_c95 bl[95] br[95] wl[146] vdd gnd cell_6t
Xbit_r147_c95 bl[95] br[95] wl[147] vdd gnd cell_6t
Xbit_r148_c95 bl[95] br[95] wl[148] vdd gnd cell_6t
Xbit_r149_c95 bl[95] br[95] wl[149] vdd gnd cell_6t
Xbit_r150_c95 bl[95] br[95] wl[150] vdd gnd cell_6t
Xbit_r151_c95 bl[95] br[95] wl[151] vdd gnd cell_6t
Xbit_r152_c95 bl[95] br[95] wl[152] vdd gnd cell_6t
Xbit_r153_c95 bl[95] br[95] wl[153] vdd gnd cell_6t
Xbit_r154_c95 bl[95] br[95] wl[154] vdd gnd cell_6t
Xbit_r155_c95 bl[95] br[95] wl[155] vdd gnd cell_6t
Xbit_r156_c95 bl[95] br[95] wl[156] vdd gnd cell_6t
Xbit_r157_c95 bl[95] br[95] wl[157] vdd gnd cell_6t
Xbit_r158_c95 bl[95] br[95] wl[158] vdd gnd cell_6t
Xbit_r159_c95 bl[95] br[95] wl[159] vdd gnd cell_6t
Xbit_r160_c95 bl[95] br[95] wl[160] vdd gnd cell_6t
Xbit_r161_c95 bl[95] br[95] wl[161] vdd gnd cell_6t
Xbit_r162_c95 bl[95] br[95] wl[162] vdd gnd cell_6t
Xbit_r163_c95 bl[95] br[95] wl[163] vdd gnd cell_6t
Xbit_r164_c95 bl[95] br[95] wl[164] vdd gnd cell_6t
Xbit_r165_c95 bl[95] br[95] wl[165] vdd gnd cell_6t
Xbit_r166_c95 bl[95] br[95] wl[166] vdd gnd cell_6t
Xbit_r167_c95 bl[95] br[95] wl[167] vdd gnd cell_6t
Xbit_r168_c95 bl[95] br[95] wl[168] vdd gnd cell_6t
Xbit_r169_c95 bl[95] br[95] wl[169] vdd gnd cell_6t
Xbit_r170_c95 bl[95] br[95] wl[170] vdd gnd cell_6t
Xbit_r171_c95 bl[95] br[95] wl[171] vdd gnd cell_6t
Xbit_r172_c95 bl[95] br[95] wl[172] vdd gnd cell_6t
Xbit_r173_c95 bl[95] br[95] wl[173] vdd gnd cell_6t
Xbit_r174_c95 bl[95] br[95] wl[174] vdd gnd cell_6t
Xbit_r175_c95 bl[95] br[95] wl[175] vdd gnd cell_6t
Xbit_r176_c95 bl[95] br[95] wl[176] vdd gnd cell_6t
Xbit_r177_c95 bl[95] br[95] wl[177] vdd gnd cell_6t
Xbit_r178_c95 bl[95] br[95] wl[178] vdd gnd cell_6t
Xbit_r179_c95 bl[95] br[95] wl[179] vdd gnd cell_6t
Xbit_r180_c95 bl[95] br[95] wl[180] vdd gnd cell_6t
Xbit_r181_c95 bl[95] br[95] wl[181] vdd gnd cell_6t
Xbit_r182_c95 bl[95] br[95] wl[182] vdd gnd cell_6t
Xbit_r183_c95 bl[95] br[95] wl[183] vdd gnd cell_6t
Xbit_r184_c95 bl[95] br[95] wl[184] vdd gnd cell_6t
Xbit_r185_c95 bl[95] br[95] wl[185] vdd gnd cell_6t
Xbit_r186_c95 bl[95] br[95] wl[186] vdd gnd cell_6t
Xbit_r187_c95 bl[95] br[95] wl[187] vdd gnd cell_6t
Xbit_r188_c95 bl[95] br[95] wl[188] vdd gnd cell_6t
Xbit_r189_c95 bl[95] br[95] wl[189] vdd gnd cell_6t
Xbit_r190_c95 bl[95] br[95] wl[190] vdd gnd cell_6t
Xbit_r191_c95 bl[95] br[95] wl[191] vdd gnd cell_6t
Xbit_r192_c95 bl[95] br[95] wl[192] vdd gnd cell_6t
Xbit_r193_c95 bl[95] br[95] wl[193] vdd gnd cell_6t
Xbit_r194_c95 bl[95] br[95] wl[194] vdd gnd cell_6t
Xbit_r195_c95 bl[95] br[95] wl[195] vdd gnd cell_6t
Xbit_r196_c95 bl[95] br[95] wl[196] vdd gnd cell_6t
Xbit_r197_c95 bl[95] br[95] wl[197] vdd gnd cell_6t
Xbit_r198_c95 bl[95] br[95] wl[198] vdd gnd cell_6t
Xbit_r199_c95 bl[95] br[95] wl[199] vdd gnd cell_6t
Xbit_r200_c95 bl[95] br[95] wl[200] vdd gnd cell_6t
Xbit_r201_c95 bl[95] br[95] wl[201] vdd gnd cell_6t
Xbit_r202_c95 bl[95] br[95] wl[202] vdd gnd cell_6t
Xbit_r203_c95 bl[95] br[95] wl[203] vdd gnd cell_6t
Xbit_r204_c95 bl[95] br[95] wl[204] vdd gnd cell_6t
Xbit_r205_c95 bl[95] br[95] wl[205] vdd gnd cell_6t
Xbit_r206_c95 bl[95] br[95] wl[206] vdd gnd cell_6t
Xbit_r207_c95 bl[95] br[95] wl[207] vdd gnd cell_6t
Xbit_r208_c95 bl[95] br[95] wl[208] vdd gnd cell_6t
Xbit_r209_c95 bl[95] br[95] wl[209] vdd gnd cell_6t
Xbit_r210_c95 bl[95] br[95] wl[210] vdd gnd cell_6t
Xbit_r211_c95 bl[95] br[95] wl[211] vdd gnd cell_6t
Xbit_r212_c95 bl[95] br[95] wl[212] vdd gnd cell_6t
Xbit_r213_c95 bl[95] br[95] wl[213] vdd gnd cell_6t
Xbit_r214_c95 bl[95] br[95] wl[214] vdd gnd cell_6t
Xbit_r215_c95 bl[95] br[95] wl[215] vdd gnd cell_6t
Xbit_r216_c95 bl[95] br[95] wl[216] vdd gnd cell_6t
Xbit_r217_c95 bl[95] br[95] wl[217] vdd gnd cell_6t
Xbit_r218_c95 bl[95] br[95] wl[218] vdd gnd cell_6t
Xbit_r219_c95 bl[95] br[95] wl[219] vdd gnd cell_6t
Xbit_r220_c95 bl[95] br[95] wl[220] vdd gnd cell_6t
Xbit_r221_c95 bl[95] br[95] wl[221] vdd gnd cell_6t
Xbit_r222_c95 bl[95] br[95] wl[222] vdd gnd cell_6t
Xbit_r223_c95 bl[95] br[95] wl[223] vdd gnd cell_6t
Xbit_r224_c95 bl[95] br[95] wl[224] vdd gnd cell_6t
Xbit_r225_c95 bl[95] br[95] wl[225] vdd gnd cell_6t
Xbit_r226_c95 bl[95] br[95] wl[226] vdd gnd cell_6t
Xbit_r227_c95 bl[95] br[95] wl[227] vdd gnd cell_6t
Xbit_r228_c95 bl[95] br[95] wl[228] vdd gnd cell_6t
Xbit_r229_c95 bl[95] br[95] wl[229] vdd gnd cell_6t
Xbit_r230_c95 bl[95] br[95] wl[230] vdd gnd cell_6t
Xbit_r231_c95 bl[95] br[95] wl[231] vdd gnd cell_6t
Xbit_r232_c95 bl[95] br[95] wl[232] vdd gnd cell_6t
Xbit_r233_c95 bl[95] br[95] wl[233] vdd gnd cell_6t
Xbit_r234_c95 bl[95] br[95] wl[234] vdd gnd cell_6t
Xbit_r235_c95 bl[95] br[95] wl[235] vdd gnd cell_6t
Xbit_r236_c95 bl[95] br[95] wl[236] vdd gnd cell_6t
Xbit_r237_c95 bl[95] br[95] wl[237] vdd gnd cell_6t
Xbit_r238_c95 bl[95] br[95] wl[238] vdd gnd cell_6t
Xbit_r239_c95 bl[95] br[95] wl[239] vdd gnd cell_6t
Xbit_r240_c95 bl[95] br[95] wl[240] vdd gnd cell_6t
Xbit_r241_c95 bl[95] br[95] wl[241] vdd gnd cell_6t
Xbit_r242_c95 bl[95] br[95] wl[242] vdd gnd cell_6t
Xbit_r243_c95 bl[95] br[95] wl[243] vdd gnd cell_6t
Xbit_r244_c95 bl[95] br[95] wl[244] vdd gnd cell_6t
Xbit_r245_c95 bl[95] br[95] wl[245] vdd gnd cell_6t
Xbit_r246_c95 bl[95] br[95] wl[246] vdd gnd cell_6t
Xbit_r247_c95 bl[95] br[95] wl[247] vdd gnd cell_6t
Xbit_r248_c95 bl[95] br[95] wl[248] vdd gnd cell_6t
Xbit_r249_c95 bl[95] br[95] wl[249] vdd gnd cell_6t
Xbit_r250_c95 bl[95] br[95] wl[250] vdd gnd cell_6t
Xbit_r251_c95 bl[95] br[95] wl[251] vdd gnd cell_6t
Xbit_r252_c95 bl[95] br[95] wl[252] vdd gnd cell_6t
Xbit_r253_c95 bl[95] br[95] wl[253] vdd gnd cell_6t
Xbit_r254_c95 bl[95] br[95] wl[254] vdd gnd cell_6t
Xbit_r255_c95 bl[95] br[95] wl[255] vdd gnd cell_6t
Xbit_r256_c95 bl[95] br[95] wl[256] vdd gnd cell_6t
Xbit_r257_c95 bl[95] br[95] wl[257] vdd gnd cell_6t
Xbit_r258_c95 bl[95] br[95] wl[258] vdd gnd cell_6t
Xbit_r259_c95 bl[95] br[95] wl[259] vdd gnd cell_6t
Xbit_r260_c95 bl[95] br[95] wl[260] vdd gnd cell_6t
Xbit_r261_c95 bl[95] br[95] wl[261] vdd gnd cell_6t
Xbit_r262_c95 bl[95] br[95] wl[262] vdd gnd cell_6t
Xbit_r263_c95 bl[95] br[95] wl[263] vdd gnd cell_6t
Xbit_r264_c95 bl[95] br[95] wl[264] vdd gnd cell_6t
Xbit_r265_c95 bl[95] br[95] wl[265] vdd gnd cell_6t
Xbit_r266_c95 bl[95] br[95] wl[266] vdd gnd cell_6t
Xbit_r267_c95 bl[95] br[95] wl[267] vdd gnd cell_6t
Xbit_r268_c95 bl[95] br[95] wl[268] vdd gnd cell_6t
Xbit_r269_c95 bl[95] br[95] wl[269] vdd gnd cell_6t
Xbit_r270_c95 bl[95] br[95] wl[270] vdd gnd cell_6t
Xbit_r271_c95 bl[95] br[95] wl[271] vdd gnd cell_6t
Xbit_r272_c95 bl[95] br[95] wl[272] vdd gnd cell_6t
Xbit_r273_c95 bl[95] br[95] wl[273] vdd gnd cell_6t
Xbit_r274_c95 bl[95] br[95] wl[274] vdd gnd cell_6t
Xbit_r275_c95 bl[95] br[95] wl[275] vdd gnd cell_6t
Xbit_r276_c95 bl[95] br[95] wl[276] vdd gnd cell_6t
Xbit_r277_c95 bl[95] br[95] wl[277] vdd gnd cell_6t
Xbit_r278_c95 bl[95] br[95] wl[278] vdd gnd cell_6t
Xbit_r279_c95 bl[95] br[95] wl[279] vdd gnd cell_6t
Xbit_r280_c95 bl[95] br[95] wl[280] vdd gnd cell_6t
Xbit_r281_c95 bl[95] br[95] wl[281] vdd gnd cell_6t
Xbit_r282_c95 bl[95] br[95] wl[282] vdd gnd cell_6t
Xbit_r283_c95 bl[95] br[95] wl[283] vdd gnd cell_6t
Xbit_r284_c95 bl[95] br[95] wl[284] vdd gnd cell_6t
Xbit_r285_c95 bl[95] br[95] wl[285] vdd gnd cell_6t
Xbit_r286_c95 bl[95] br[95] wl[286] vdd gnd cell_6t
Xbit_r287_c95 bl[95] br[95] wl[287] vdd gnd cell_6t
Xbit_r288_c95 bl[95] br[95] wl[288] vdd gnd cell_6t
Xbit_r289_c95 bl[95] br[95] wl[289] vdd gnd cell_6t
Xbit_r290_c95 bl[95] br[95] wl[290] vdd gnd cell_6t
Xbit_r291_c95 bl[95] br[95] wl[291] vdd gnd cell_6t
Xbit_r292_c95 bl[95] br[95] wl[292] vdd gnd cell_6t
Xbit_r293_c95 bl[95] br[95] wl[293] vdd gnd cell_6t
Xbit_r294_c95 bl[95] br[95] wl[294] vdd gnd cell_6t
Xbit_r295_c95 bl[95] br[95] wl[295] vdd gnd cell_6t
Xbit_r296_c95 bl[95] br[95] wl[296] vdd gnd cell_6t
Xbit_r297_c95 bl[95] br[95] wl[297] vdd gnd cell_6t
Xbit_r298_c95 bl[95] br[95] wl[298] vdd gnd cell_6t
Xbit_r299_c95 bl[95] br[95] wl[299] vdd gnd cell_6t
Xbit_r300_c95 bl[95] br[95] wl[300] vdd gnd cell_6t
Xbit_r301_c95 bl[95] br[95] wl[301] vdd gnd cell_6t
Xbit_r302_c95 bl[95] br[95] wl[302] vdd gnd cell_6t
Xbit_r303_c95 bl[95] br[95] wl[303] vdd gnd cell_6t
Xbit_r304_c95 bl[95] br[95] wl[304] vdd gnd cell_6t
Xbit_r305_c95 bl[95] br[95] wl[305] vdd gnd cell_6t
Xbit_r306_c95 bl[95] br[95] wl[306] vdd gnd cell_6t
Xbit_r307_c95 bl[95] br[95] wl[307] vdd gnd cell_6t
Xbit_r308_c95 bl[95] br[95] wl[308] vdd gnd cell_6t
Xbit_r309_c95 bl[95] br[95] wl[309] vdd gnd cell_6t
Xbit_r310_c95 bl[95] br[95] wl[310] vdd gnd cell_6t
Xbit_r311_c95 bl[95] br[95] wl[311] vdd gnd cell_6t
Xbit_r312_c95 bl[95] br[95] wl[312] vdd gnd cell_6t
Xbit_r313_c95 bl[95] br[95] wl[313] vdd gnd cell_6t
Xbit_r314_c95 bl[95] br[95] wl[314] vdd gnd cell_6t
Xbit_r315_c95 bl[95] br[95] wl[315] vdd gnd cell_6t
Xbit_r316_c95 bl[95] br[95] wl[316] vdd gnd cell_6t
Xbit_r317_c95 bl[95] br[95] wl[317] vdd gnd cell_6t
Xbit_r318_c95 bl[95] br[95] wl[318] vdd gnd cell_6t
Xbit_r319_c95 bl[95] br[95] wl[319] vdd gnd cell_6t
Xbit_r320_c95 bl[95] br[95] wl[320] vdd gnd cell_6t
Xbit_r321_c95 bl[95] br[95] wl[321] vdd gnd cell_6t
Xbit_r322_c95 bl[95] br[95] wl[322] vdd gnd cell_6t
Xbit_r323_c95 bl[95] br[95] wl[323] vdd gnd cell_6t
Xbit_r324_c95 bl[95] br[95] wl[324] vdd gnd cell_6t
Xbit_r325_c95 bl[95] br[95] wl[325] vdd gnd cell_6t
Xbit_r326_c95 bl[95] br[95] wl[326] vdd gnd cell_6t
Xbit_r327_c95 bl[95] br[95] wl[327] vdd gnd cell_6t
Xbit_r328_c95 bl[95] br[95] wl[328] vdd gnd cell_6t
Xbit_r329_c95 bl[95] br[95] wl[329] vdd gnd cell_6t
Xbit_r330_c95 bl[95] br[95] wl[330] vdd gnd cell_6t
Xbit_r331_c95 bl[95] br[95] wl[331] vdd gnd cell_6t
Xbit_r332_c95 bl[95] br[95] wl[332] vdd gnd cell_6t
Xbit_r333_c95 bl[95] br[95] wl[333] vdd gnd cell_6t
Xbit_r334_c95 bl[95] br[95] wl[334] vdd gnd cell_6t
Xbit_r335_c95 bl[95] br[95] wl[335] vdd gnd cell_6t
Xbit_r336_c95 bl[95] br[95] wl[336] vdd gnd cell_6t
Xbit_r337_c95 bl[95] br[95] wl[337] vdd gnd cell_6t
Xbit_r338_c95 bl[95] br[95] wl[338] vdd gnd cell_6t
Xbit_r339_c95 bl[95] br[95] wl[339] vdd gnd cell_6t
Xbit_r340_c95 bl[95] br[95] wl[340] vdd gnd cell_6t
Xbit_r341_c95 bl[95] br[95] wl[341] vdd gnd cell_6t
Xbit_r342_c95 bl[95] br[95] wl[342] vdd gnd cell_6t
Xbit_r343_c95 bl[95] br[95] wl[343] vdd gnd cell_6t
Xbit_r344_c95 bl[95] br[95] wl[344] vdd gnd cell_6t
Xbit_r345_c95 bl[95] br[95] wl[345] vdd gnd cell_6t
Xbit_r346_c95 bl[95] br[95] wl[346] vdd gnd cell_6t
Xbit_r347_c95 bl[95] br[95] wl[347] vdd gnd cell_6t
Xbit_r348_c95 bl[95] br[95] wl[348] vdd gnd cell_6t
Xbit_r349_c95 bl[95] br[95] wl[349] vdd gnd cell_6t
Xbit_r350_c95 bl[95] br[95] wl[350] vdd gnd cell_6t
Xbit_r351_c95 bl[95] br[95] wl[351] vdd gnd cell_6t
Xbit_r352_c95 bl[95] br[95] wl[352] vdd gnd cell_6t
Xbit_r353_c95 bl[95] br[95] wl[353] vdd gnd cell_6t
Xbit_r354_c95 bl[95] br[95] wl[354] vdd gnd cell_6t
Xbit_r355_c95 bl[95] br[95] wl[355] vdd gnd cell_6t
Xbit_r356_c95 bl[95] br[95] wl[356] vdd gnd cell_6t
Xbit_r357_c95 bl[95] br[95] wl[357] vdd gnd cell_6t
Xbit_r358_c95 bl[95] br[95] wl[358] vdd gnd cell_6t
Xbit_r359_c95 bl[95] br[95] wl[359] vdd gnd cell_6t
Xbit_r360_c95 bl[95] br[95] wl[360] vdd gnd cell_6t
Xbit_r361_c95 bl[95] br[95] wl[361] vdd gnd cell_6t
Xbit_r362_c95 bl[95] br[95] wl[362] vdd gnd cell_6t
Xbit_r363_c95 bl[95] br[95] wl[363] vdd gnd cell_6t
Xbit_r364_c95 bl[95] br[95] wl[364] vdd gnd cell_6t
Xbit_r365_c95 bl[95] br[95] wl[365] vdd gnd cell_6t
Xbit_r366_c95 bl[95] br[95] wl[366] vdd gnd cell_6t
Xbit_r367_c95 bl[95] br[95] wl[367] vdd gnd cell_6t
Xbit_r368_c95 bl[95] br[95] wl[368] vdd gnd cell_6t
Xbit_r369_c95 bl[95] br[95] wl[369] vdd gnd cell_6t
Xbit_r370_c95 bl[95] br[95] wl[370] vdd gnd cell_6t
Xbit_r371_c95 bl[95] br[95] wl[371] vdd gnd cell_6t
Xbit_r372_c95 bl[95] br[95] wl[372] vdd gnd cell_6t
Xbit_r373_c95 bl[95] br[95] wl[373] vdd gnd cell_6t
Xbit_r374_c95 bl[95] br[95] wl[374] vdd gnd cell_6t
Xbit_r375_c95 bl[95] br[95] wl[375] vdd gnd cell_6t
Xbit_r376_c95 bl[95] br[95] wl[376] vdd gnd cell_6t
Xbit_r377_c95 bl[95] br[95] wl[377] vdd gnd cell_6t
Xbit_r378_c95 bl[95] br[95] wl[378] vdd gnd cell_6t
Xbit_r379_c95 bl[95] br[95] wl[379] vdd gnd cell_6t
Xbit_r380_c95 bl[95] br[95] wl[380] vdd gnd cell_6t
Xbit_r381_c95 bl[95] br[95] wl[381] vdd gnd cell_6t
Xbit_r382_c95 bl[95] br[95] wl[382] vdd gnd cell_6t
Xbit_r383_c95 bl[95] br[95] wl[383] vdd gnd cell_6t
Xbit_r384_c95 bl[95] br[95] wl[384] vdd gnd cell_6t
Xbit_r385_c95 bl[95] br[95] wl[385] vdd gnd cell_6t
Xbit_r386_c95 bl[95] br[95] wl[386] vdd gnd cell_6t
Xbit_r387_c95 bl[95] br[95] wl[387] vdd gnd cell_6t
Xbit_r388_c95 bl[95] br[95] wl[388] vdd gnd cell_6t
Xbit_r389_c95 bl[95] br[95] wl[389] vdd gnd cell_6t
Xbit_r390_c95 bl[95] br[95] wl[390] vdd gnd cell_6t
Xbit_r391_c95 bl[95] br[95] wl[391] vdd gnd cell_6t
Xbit_r392_c95 bl[95] br[95] wl[392] vdd gnd cell_6t
Xbit_r393_c95 bl[95] br[95] wl[393] vdd gnd cell_6t
Xbit_r394_c95 bl[95] br[95] wl[394] vdd gnd cell_6t
Xbit_r395_c95 bl[95] br[95] wl[395] vdd gnd cell_6t
Xbit_r396_c95 bl[95] br[95] wl[396] vdd gnd cell_6t
Xbit_r397_c95 bl[95] br[95] wl[397] vdd gnd cell_6t
Xbit_r398_c95 bl[95] br[95] wl[398] vdd gnd cell_6t
Xbit_r399_c95 bl[95] br[95] wl[399] vdd gnd cell_6t
Xbit_r400_c95 bl[95] br[95] wl[400] vdd gnd cell_6t
Xbit_r401_c95 bl[95] br[95] wl[401] vdd gnd cell_6t
Xbit_r402_c95 bl[95] br[95] wl[402] vdd gnd cell_6t
Xbit_r403_c95 bl[95] br[95] wl[403] vdd gnd cell_6t
Xbit_r404_c95 bl[95] br[95] wl[404] vdd gnd cell_6t
Xbit_r405_c95 bl[95] br[95] wl[405] vdd gnd cell_6t
Xbit_r406_c95 bl[95] br[95] wl[406] vdd gnd cell_6t
Xbit_r407_c95 bl[95] br[95] wl[407] vdd gnd cell_6t
Xbit_r408_c95 bl[95] br[95] wl[408] vdd gnd cell_6t
Xbit_r409_c95 bl[95] br[95] wl[409] vdd gnd cell_6t
Xbit_r410_c95 bl[95] br[95] wl[410] vdd gnd cell_6t
Xbit_r411_c95 bl[95] br[95] wl[411] vdd gnd cell_6t
Xbit_r412_c95 bl[95] br[95] wl[412] vdd gnd cell_6t
Xbit_r413_c95 bl[95] br[95] wl[413] vdd gnd cell_6t
Xbit_r414_c95 bl[95] br[95] wl[414] vdd gnd cell_6t
Xbit_r415_c95 bl[95] br[95] wl[415] vdd gnd cell_6t
Xbit_r416_c95 bl[95] br[95] wl[416] vdd gnd cell_6t
Xbit_r417_c95 bl[95] br[95] wl[417] vdd gnd cell_6t
Xbit_r418_c95 bl[95] br[95] wl[418] vdd gnd cell_6t
Xbit_r419_c95 bl[95] br[95] wl[419] vdd gnd cell_6t
Xbit_r420_c95 bl[95] br[95] wl[420] vdd gnd cell_6t
Xbit_r421_c95 bl[95] br[95] wl[421] vdd gnd cell_6t
Xbit_r422_c95 bl[95] br[95] wl[422] vdd gnd cell_6t
Xbit_r423_c95 bl[95] br[95] wl[423] vdd gnd cell_6t
Xbit_r424_c95 bl[95] br[95] wl[424] vdd gnd cell_6t
Xbit_r425_c95 bl[95] br[95] wl[425] vdd gnd cell_6t
Xbit_r426_c95 bl[95] br[95] wl[426] vdd gnd cell_6t
Xbit_r427_c95 bl[95] br[95] wl[427] vdd gnd cell_6t
Xbit_r428_c95 bl[95] br[95] wl[428] vdd gnd cell_6t
Xbit_r429_c95 bl[95] br[95] wl[429] vdd gnd cell_6t
Xbit_r430_c95 bl[95] br[95] wl[430] vdd gnd cell_6t
Xbit_r431_c95 bl[95] br[95] wl[431] vdd gnd cell_6t
Xbit_r432_c95 bl[95] br[95] wl[432] vdd gnd cell_6t
Xbit_r433_c95 bl[95] br[95] wl[433] vdd gnd cell_6t
Xbit_r434_c95 bl[95] br[95] wl[434] vdd gnd cell_6t
Xbit_r435_c95 bl[95] br[95] wl[435] vdd gnd cell_6t
Xbit_r436_c95 bl[95] br[95] wl[436] vdd gnd cell_6t
Xbit_r437_c95 bl[95] br[95] wl[437] vdd gnd cell_6t
Xbit_r438_c95 bl[95] br[95] wl[438] vdd gnd cell_6t
Xbit_r439_c95 bl[95] br[95] wl[439] vdd gnd cell_6t
Xbit_r440_c95 bl[95] br[95] wl[440] vdd gnd cell_6t
Xbit_r441_c95 bl[95] br[95] wl[441] vdd gnd cell_6t
Xbit_r442_c95 bl[95] br[95] wl[442] vdd gnd cell_6t
Xbit_r443_c95 bl[95] br[95] wl[443] vdd gnd cell_6t
Xbit_r444_c95 bl[95] br[95] wl[444] vdd gnd cell_6t
Xbit_r445_c95 bl[95] br[95] wl[445] vdd gnd cell_6t
Xbit_r446_c95 bl[95] br[95] wl[446] vdd gnd cell_6t
Xbit_r447_c95 bl[95] br[95] wl[447] vdd gnd cell_6t
Xbit_r448_c95 bl[95] br[95] wl[448] vdd gnd cell_6t
Xbit_r449_c95 bl[95] br[95] wl[449] vdd gnd cell_6t
Xbit_r450_c95 bl[95] br[95] wl[450] vdd gnd cell_6t
Xbit_r451_c95 bl[95] br[95] wl[451] vdd gnd cell_6t
Xbit_r452_c95 bl[95] br[95] wl[452] vdd gnd cell_6t
Xbit_r453_c95 bl[95] br[95] wl[453] vdd gnd cell_6t
Xbit_r454_c95 bl[95] br[95] wl[454] vdd gnd cell_6t
Xbit_r455_c95 bl[95] br[95] wl[455] vdd gnd cell_6t
Xbit_r456_c95 bl[95] br[95] wl[456] vdd gnd cell_6t
Xbit_r457_c95 bl[95] br[95] wl[457] vdd gnd cell_6t
Xbit_r458_c95 bl[95] br[95] wl[458] vdd gnd cell_6t
Xbit_r459_c95 bl[95] br[95] wl[459] vdd gnd cell_6t
Xbit_r460_c95 bl[95] br[95] wl[460] vdd gnd cell_6t
Xbit_r461_c95 bl[95] br[95] wl[461] vdd gnd cell_6t
Xbit_r462_c95 bl[95] br[95] wl[462] vdd gnd cell_6t
Xbit_r463_c95 bl[95] br[95] wl[463] vdd gnd cell_6t
Xbit_r464_c95 bl[95] br[95] wl[464] vdd gnd cell_6t
Xbit_r465_c95 bl[95] br[95] wl[465] vdd gnd cell_6t
Xbit_r466_c95 bl[95] br[95] wl[466] vdd gnd cell_6t
Xbit_r467_c95 bl[95] br[95] wl[467] vdd gnd cell_6t
Xbit_r468_c95 bl[95] br[95] wl[468] vdd gnd cell_6t
Xbit_r469_c95 bl[95] br[95] wl[469] vdd gnd cell_6t
Xbit_r470_c95 bl[95] br[95] wl[470] vdd gnd cell_6t
Xbit_r471_c95 bl[95] br[95] wl[471] vdd gnd cell_6t
Xbit_r472_c95 bl[95] br[95] wl[472] vdd gnd cell_6t
Xbit_r473_c95 bl[95] br[95] wl[473] vdd gnd cell_6t
Xbit_r474_c95 bl[95] br[95] wl[474] vdd gnd cell_6t
Xbit_r475_c95 bl[95] br[95] wl[475] vdd gnd cell_6t
Xbit_r476_c95 bl[95] br[95] wl[476] vdd gnd cell_6t
Xbit_r477_c95 bl[95] br[95] wl[477] vdd gnd cell_6t
Xbit_r478_c95 bl[95] br[95] wl[478] vdd gnd cell_6t
Xbit_r479_c95 bl[95] br[95] wl[479] vdd gnd cell_6t
Xbit_r480_c95 bl[95] br[95] wl[480] vdd gnd cell_6t
Xbit_r481_c95 bl[95] br[95] wl[481] vdd gnd cell_6t
Xbit_r482_c95 bl[95] br[95] wl[482] vdd gnd cell_6t
Xbit_r483_c95 bl[95] br[95] wl[483] vdd gnd cell_6t
Xbit_r484_c95 bl[95] br[95] wl[484] vdd gnd cell_6t
Xbit_r485_c95 bl[95] br[95] wl[485] vdd gnd cell_6t
Xbit_r486_c95 bl[95] br[95] wl[486] vdd gnd cell_6t
Xbit_r487_c95 bl[95] br[95] wl[487] vdd gnd cell_6t
Xbit_r488_c95 bl[95] br[95] wl[488] vdd gnd cell_6t
Xbit_r489_c95 bl[95] br[95] wl[489] vdd gnd cell_6t
Xbit_r490_c95 bl[95] br[95] wl[490] vdd gnd cell_6t
Xbit_r491_c95 bl[95] br[95] wl[491] vdd gnd cell_6t
Xbit_r492_c95 bl[95] br[95] wl[492] vdd gnd cell_6t
Xbit_r493_c95 bl[95] br[95] wl[493] vdd gnd cell_6t
Xbit_r494_c95 bl[95] br[95] wl[494] vdd gnd cell_6t
Xbit_r495_c95 bl[95] br[95] wl[495] vdd gnd cell_6t
Xbit_r496_c95 bl[95] br[95] wl[496] vdd gnd cell_6t
Xbit_r497_c95 bl[95] br[95] wl[497] vdd gnd cell_6t
Xbit_r498_c95 bl[95] br[95] wl[498] vdd gnd cell_6t
Xbit_r499_c95 bl[95] br[95] wl[499] vdd gnd cell_6t
Xbit_r500_c95 bl[95] br[95] wl[500] vdd gnd cell_6t
Xbit_r501_c95 bl[95] br[95] wl[501] vdd gnd cell_6t
Xbit_r502_c95 bl[95] br[95] wl[502] vdd gnd cell_6t
Xbit_r503_c95 bl[95] br[95] wl[503] vdd gnd cell_6t
Xbit_r504_c95 bl[95] br[95] wl[504] vdd gnd cell_6t
Xbit_r505_c95 bl[95] br[95] wl[505] vdd gnd cell_6t
Xbit_r506_c95 bl[95] br[95] wl[506] vdd gnd cell_6t
Xbit_r507_c95 bl[95] br[95] wl[507] vdd gnd cell_6t
Xbit_r508_c95 bl[95] br[95] wl[508] vdd gnd cell_6t
Xbit_r509_c95 bl[95] br[95] wl[509] vdd gnd cell_6t
Xbit_r510_c95 bl[95] br[95] wl[510] vdd gnd cell_6t
Xbit_r511_c95 bl[95] br[95] wl[511] vdd gnd cell_6t
Xbit_r0_c96 bl[96] br[96] wl[0] vdd gnd cell_6t
Xbit_r1_c96 bl[96] br[96] wl[1] vdd gnd cell_6t
Xbit_r2_c96 bl[96] br[96] wl[2] vdd gnd cell_6t
Xbit_r3_c96 bl[96] br[96] wl[3] vdd gnd cell_6t
Xbit_r4_c96 bl[96] br[96] wl[4] vdd gnd cell_6t
Xbit_r5_c96 bl[96] br[96] wl[5] vdd gnd cell_6t
Xbit_r6_c96 bl[96] br[96] wl[6] vdd gnd cell_6t
Xbit_r7_c96 bl[96] br[96] wl[7] vdd gnd cell_6t
Xbit_r8_c96 bl[96] br[96] wl[8] vdd gnd cell_6t
Xbit_r9_c96 bl[96] br[96] wl[9] vdd gnd cell_6t
Xbit_r10_c96 bl[96] br[96] wl[10] vdd gnd cell_6t
Xbit_r11_c96 bl[96] br[96] wl[11] vdd gnd cell_6t
Xbit_r12_c96 bl[96] br[96] wl[12] vdd gnd cell_6t
Xbit_r13_c96 bl[96] br[96] wl[13] vdd gnd cell_6t
Xbit_r14_c96 bl[96] br[96] wl[14] vdd gnd cell_6t
Xbit_r15_c96 bl[96] br[96] wl[15] vdd gnd cell_6t
Xbit_r16_c96 bl[96] br[96] wl[16] vdd gnd cell_6t
Xbit_r17_c96 bl[96] br[96] wl[17] vdd gnd cell_6t
Xbit_r18_c96 bl[96] br[96] wl[18] vdd gnd cell_6t
Xbit_r19_c96 bl[96] br[96] wl[19] vdd gnd cell_6t
Xbit_r20_c96 bl[96] br[96] wl[20] vdd gnd cell_6t
Xbit_r21_c96 bl[96] br[96] wl[21] vdd gnd cell_6t
Xbit_r22_c96 bl[96] br[96] wl[22] vdd gnd cell_6t
Xbit_r23_c96 bl[96] br[96] wl[23] vdd gnd cell_6t
Xbit_r24_c96 bl[96] br[96] wl[24] vdd gnd cell_6t
Xbit_r25_c96 bl[96] br[96] wl[25] vdd gnd cell_6t
Xbit_r26_c96 bl[96] br[96] wl[26] vdd gnd cell_6t
Xbit_r27_c96 bl[96] br[96] wl[27] vdd gnd cell_6t
Xbit_r28_c96 bl[96] br[96] wl[28] vdd gnd cell_6t
Xbit_r29_c96 bl[96] br[96] wl[29] vdd gnd cell_6t
Xbit_r30_c96 bl[96] br[96] wl[30] vdd gnd cell_6t
Xbit_r31_c96 bl[96] br[96] wl[31] vdd gnd cell_6t
Xbit_r32_c96 bl[96] br[96] wl[32] vdd gnd cell_6t
Xbit_r33_c96 bl[96] br[96] wl[33] vdd gnd cell_6t
Xbit_r34_c96 bl[96] br[96] wl[34] vdd gnd cell_6t
Xbit_r35_c96 bl[96] br[96] wl[35] vdd gnd cell_6t
Xbit_r36_c96 bl[96] br[96] wl[36] vdd gnd cell_6t
Xbit_r37_c96 bl[96] br[96] wl[37] vdd gnd cell_6t
Xbit_r38_c96 bl[96] br[96] wl[38] vdd gnd cell_6t
Xbit_r39_c96 bl[96] br[96] wl[39] vdd gnd cell_6t
Xbit_r40_c96 bl[96] br[96] wl[40] vdd gnd cell_6t
Xbit_r41_c96 bl[96] br[96] wl[41] vdd gnd cell_6t
Xbit_r42_c96 bl[96] br[96] wl[42] vdd gnd cell_6t
Xbit_r43_c96 bl[96] br[96] wl[43] vdd gnd cell_6t
Xbit_r44_c96 bl[96] br[96] wl[44] vdd gnd cell_6t
Xbit_r45_c96 bl[96] br[96] wl[45] vdd gnd cell_6t
Xbit_r46_c96 bl[96] br[96] wl[46] vdd gnd cell_6t
Xbit_r47_c96 bl[96] br[96] wl[47] vdd gnd cell_6t
Xbit_r48_c96 bl[96] br[96] wl[48] vdd gnd cell_6t
Xbit_r49_c96 bl[96] br[96] wl[49] vdd gnd cell_6t
Xbit_r50_c96 bl[96] br[96] wl[50] vdd gnd cell_6t
Xbit_r51_c96 bl[96] br[96] wl[51] vdd gnd cell_6t
Xbit_r52_c96 bl[96] br[96] wl[52] vdd gnd cell_6t
Xbit_r53_c96 bl[96] br[96] wl[53] vdd gnd cell_6t
Xbit_r54_c96 bl[96] br[96] wl[54] vdd gnd cell_6t
Xbit_r55_c96 bl[96] br[96] wl[55] vdd gnd cell_6t
Xbit_r56_c96 bl[96] br[96] wl[56] vdd gnd cell_6t
Xbit_r57_c96 bl[96] br[96] wl[57] vdd gnd cell_6t
Xbit_r58_c96 bl[96] br[96] wl[58] vdd gnd cell_6t
Xbit_r59_c96 bl[96] br[96] wl[59] vdd gnd cell_6t
Xbit_r60_c96 bl[96] br[96] wl[60] vdd gnd cell_6t
Xbit_r61_c96 bl[96] br[96] wl[61] vdd gnd cell_6t
Xbit_r62_c96 bl[96] br[96] wl[62] vdd gnd cell_6t
Xbit_r63_c96 bl[96] br[96] wl[63] vdd gnd cell_6t
Xbit_r64_c96 bl[96] br[96] wl[64] vdd gnd cell_6t
Xbit_r65_c96 bl[96] br[96] wl[65] vdd gnd cell_6t
Xbit_r66_c96 bl[96] br[96] wl[66] vdd gnd cell_6t
Xbit_r67_c96 bl[96] br[96] wl[67] vdd gnd cell_6t
Xbit_r68_c96 bl[96] br[96] wl[68] vdd gnd cell_6t
Xbit_r69_c96 bl[96] br[96] wl[69] vdd gnd cell_6t
Xbit_r70_c96 bl[96] br[96] wl[70] vdd gnd cell_6t
Xbit_r71_c96 bl[96] br[96] wl[71] vdd gnd cell_6t
Xbit_r72_c96 bl[96] br[96] wl[72] vdd gnd cell_6t
Xbit_r73_c96 bl[96] br[96] wl[73] vdd gnd cell_6t
Xbit_r74_c96 bl[96] br[96] wl[74] vdd gnd cell_6t
Xbit_r75_c96 bl[96] br[96] wl[75] vdd gnd cell_6t
Xbit_r76_c96 bl[96] br[96] wl[76] vdd gnd cell_6t
Xbit_r77_c96 bl[96] br[96] wl[77] vdd gnd cell_6t
Xbit_r78_c96 bl[96] br[96] wl[78] vdd gnd cell_6t
Xbit_r79_c96 bl[96] br[96] wl[79] vdd gnd cell_6t
Xbit_r80_c96 bl[96] br[96] wl[80] vdd gnd cell_6t
Xbit_r81_c96 bl[96] br[96] wl[81] vdd gnd cell_6t
Xbit_r82_c96 bl[96] br[96] wl[82] vdd gnd cell_6t
Xbit_r83_c96 bl[96] br[96] wl[83] vdd gnd cell_6t
Xbit_r84_c96 bl[96] br[96] wl[84] vdd gnd cell_6t
Xbit_r85_c96 bl[96] br[96] wl[85] vdd gnd cell_6t
Xbit_r86_c96 bl[96] br[96] wl[86] vdd gnd cell_6t
Xbit_r87_c96 bl[96] br[96] wl[87] vdd gnd cell_6t
Xbit_r88_c96 bl[96] br[96] wl[88] vdd gnd cell_6t
Xbit_r89_c96 bl[96] br[96] wl[89] vdd gnd cell_6t
Xbit_r90_c96 bl[96] br[96] wl[90] vdd gnd cell_6t
Xbit_r91_c96 bl[96] br[96] wl[91] vdd gnd cell_6t
Xbit_r92_c96 bl[96] br[96] wl[92] vdd gnd cell_6t
Xbit_r93_c96 bl[96] br[96] wl[93] vdd gnd cell_6t
Xbit_r94_c96 bl[96] br[96] wl[94] vdd gnd cell_6t
Xbit_r95_c96 bl[96] br[96] wl[95] vdd gnd cell_6t
Xbit_r96_c96 bl[96] br[96] wl[96] vdd gnd cell_6t
Xbit_r97_c96 bl[96] br[96] wl[97] vdd gnd cell_6t
Xbit_r98_c96 bl[96] br[96] wl[98] vdd gnd cell_6t
Xbit_r99_c96 bl[96] br[96] wl[99] vdd gnd cell_6t
Xbit_r100_c96 bl[96] br[96] wl[100] vdd gnd cell_6t
Xbit_r101_c96 bl[96] br[96] wl[101] vdd gnd cell_6t
Xbit_r102_c96 bl[96] br[96] wl[102] vdd gnd cell_6t
Xbit_r103_c96 bl[96] br[96] wl[103] vdd gnd cell_6t
Xbit_r104_c96 bl[96] br[96] wl[104] vdd gnd cell_6t
Xbit_r105_c96 bl[96] br[96] wl[105] vdd gnd cell_6t
Xbit_r106_c96 bl[96] br[96] wl[106] vdd gnd cell_6t
Xbit_r107_c96 bl[96] br[96] wl[107] vdd gnd cell_6t
Xbit_r108_c96 bl[96] br[96] wl[108] vdd gnd cell_6t
Xbit_r109_c96 bl[96] br[96] wl[109] vdd gnd cell_6t
Xbit_r110_c96 bl[96] br[96] wl[110] vdd gnd cell_6t
Xbit_r111_c96 bl[96] br[96] wl[111] vdd gnd cell_6t
Xbit_r112_c96 bl[96] br[96] wl[112] vdd gnd cell_6t
Xbit_r113_c96 bl[96] br[96] wl[113] vdd gnd cell_6t
Xbit_r114_c96 bl[96] br[96] wl[114] vdd gnd cell_6t
Xbit_r115_c96 bl[96] br[96] wl[115] vdd gnd cell_6t
Xbit_r116_c96 bl[96] br[96] wl[116] vdd gnd cell_6t
Xbit_r117_c96 bl[96] br[96] wl[117] vdd gnd cell_6t
Xbit_r118_c96 bl[96] br[96] wl[118] vdd gnd cell_6t
Xbit_r119_c96 bl[96] br[96] wl[119] vdd gnd cell_6t
Xbit_r120_c96 bl[96] br[96] wl[120] vdd gnd cell_6t
Xbit_r121_c96 bl[96] br[96] wl[121] vdd gnd cell_6t
Xbit_r122_c96 bl[96] br[96] wl[122] vdd gnd cell_6t
Xbit_r123_c96 bl[96] br[96] wl[123] vdd gnd cell_6t
Xbit_r124_c96 bl[96] br[96] wl[124] vdd gnd cell_6t
Xbit_r125_c96 bl[96] br[96] wl[125] vdd gnd cell_6t
Xbit_r126_c96 bl[96] br[96] wl[126] vdd gnd cell_6t
Xbit_r127_c96 bl[96] br[96] wl[127] vdd gnd cell_6t
Xbit_r128_c96 bl[96] br[96] wl[128] vdd gnd cell_6t
Xbit_r129_c96 bl[96] br[96] wl[129] vdd gnd cell_6t
Xbit_r130_c96 bl[96] br[96] wl[130] vdd gnd cell_6t
Xbit_r131_c96 bl[96] br[96] wl[131] vdd gnd cell_6t
Xbit_r132_c96 bl[96] br[96] wl[132] vdd gnd cell_6t
Xbit_r133_c96 bl[96] br[96] wl[133] vdd gnd cell_6t
Xbit_r134_c96 bl[96] br[96] wl[134] vdd gnd cell_6t
Xbit_r135_c96 bl[96] br[96] wl[135] vdd gnd cell_6t
Xbit_r136_c96 bl[96] br[96] wl[136] vdd gnd cell_6t
Xbit_r137_c96 bl[96] br[96] wl[137] vdd gnd cell_6t
Xbit_r138_c96 bl[96] br[96] wl[138] vdd gnd cell_6t
Xbit_r139_c96 bl[96] br[96] wl[139] vdd gnd cell_6t
Xbit_r140_c96 bl[96] br[96] wl[140] vdd gnd cell_6t
Xbit_r141_c96 bl[96] br[96] wl[141] vdd gnd cell_6t
Xbit_r142_c96 bl[96] br[96] wl[142] vdd gnd cell_6t
Xbit_r143_c96 bl[96] br[96] wl[143] vdd gnd cell_6t
Xbit_r144_c96 bl[96] br[96] wl[144] vdd gnd cell_6t
Xbit_r145_c96 bl[96] br[96] wl[145] vdd gnd cell_6t
Xbit_r146_c96 bl[96] br[96] wl[146] vdd gnd cell_6t
Xbit_r147_c96 bl[96] br[96] wl[147] vdd gnd cell_6t
Xbit_r148_c96 bl[96] br[96] wl[148] vdd gnd cell_6t
Xbit_r149_c96 bl[96] br[96] wl[149] vdd gnd cell_6t
Xbit_r150_c96 bl[96] br[96] wl[150] vdd gnd cell_6t
Xbit_r151_c96 bl[96] br[96] wl[151] vdd gnd cell_6t
Xbit_r152_c96 bl[96] br[96] wl[152] vdd gnd cell_6t
Xbit_r153_c96 bl[96] br[96] wl[153] vdd gnd cell_6t
Xbit_r154_c96 bl[96] br[96] wl[154] vdd gnd cell_6t
Xbit_r155_c96 bl[96] br[96] wl[155] vdd gnd cell_6t
Xbit_r156_c96 bl[96] br[96] wl[156] vdd gnd cell_6t
Xbit_r157_c96 bl[96] br[96] wl[157] vdd gnd cell_6t
Xbit_r158_c96 bl[96] br[96] wl[158] vdd gnd cell_6t
Xbit_r159_c96 bl[96] br[96] wl[159] vdd gnd cell_6t
Xbit_r160_c96 bl[96] br[96] wl[160] vdd gnd cell_6t
Xbit_r161_c96 bl[96] br[96] wl[161] vdd gnd cell_6t
Xbit_r162_c96 bl[96] br[96] wl[162] vdd gnd cell_6t
Xbit_r163_c96 bl[96] br[96] wl[163] vdd gnd cell_6t
Xbit_r164_c96 bl[96] br[96] wl[164] vdd gnd cell_6t
Xbit_r165_c96 bl[96] br[96] wl[165] vdd gnd cell_6t
Xbit_r166_c96 bl[96] br[96] wl[166] vdd gnd cell_6t
Xbit_r167_c96 bl[96] br[96] wl[167] vdd gnd cell_6t
Xbit_r168_c96 bl[96] br[96] wl[168] vdd gnd cell_6t
Xbit_r169_c96 bl[96] br[96] wl[169] vdd gnd cell_6t
Xbit_r170_c96 bl[96] br[96] wl[170] vdd gnd cell_6t
Xbit_r171_c96 bl[96] br[96] wl[171] vdd gnd cell_6t
Xbit_r172_c96 bl[96] br[96] wl[172] vdd gnd cell_6t
Xbit_r173_c96 bl[96] br[96] wl[173] vdd gnd cell_6t
Xbit_r174_c96 bl[96] br[96] wl[174] vdd gnd cell_6t
Xbit_r175_c96 bl[96] br[96] wl[175] vdd gnd cell_6t
Xbit_r176_c96 bl[96] br[96] wl[176] vdd gnd cell_6t
Xbit_r177_c96 bl[96] br[96] wl[177] vdd gnd cell_6t
Xbit_r178_c96 bl[96] br[96] wl[178] vdd gnd cell_6t
Xbit_r179_c96 bl[96] br[96] wl[179] vdd gnd cell_6t
Xbit_r180_c96 bl[96] br[96] wl[180] vdd gnd cell_6t
Xbit_r181_c96 bl[96] br[96] wl[181] vdd gnd cell_6t
Xbit_r182_c96 bl[96] br[96] wl[182] vdd gnd cell_6t
Xbit_r183_c96 bl[96] br[96] wl[183] vdd gnd cell_6t
Xbit_r184_c96 bl[96] br[96] wl[184] vdd gnd cell_6t
Xbit_r185_c96 bl[96] br[96] wl[185] vdd gnd cell_6t
Xbit_r186_c96 bl[96] br[96] wl[186] vdd gnd cell_6t
Xbit_r187_c96 bl[96] br[96] wl[187] vdd gnd cell_6t
Xbit_r188_c96 bl[96] br[96] wl[188] vdd gnd cell_6t
Xbit_r189_c96 bl[96] br[96] wl[189] vdd gnd cell_6t
Xbit_r190_c96 bl[96] br[96] wl[190] vdd gnd cell_6t
Xbit_r191_c96 bl[96] br[96] wl[191] vdd gnd cell_6t
Xbit_r192_c96 bl[96] br[96] wl[192] vdd gnd cell_6t
Xbit_r193_c96 bl[96] br[96] wl[193] vdd gnd cell_6t
Xbit_r194_c96 bl[96] br[96] wl[194] vdd gnd cell_6t
Xbit_r195_c96 bl[96] br[96] wl[195] vdd gnd cell_6t
Xbit_r196_c96 bl[96] br[96] wl[196] vdd gnd cell_6t
Xbit_r197_c96 bl[96] br[96] wl[197] vdd gnd cell_6t
Xbit_r198_c96 bl[96] br[96] wl[198] vdd gnd cell_6t
Xbit_r199_c96 bl[96] br[96] wl[199] vdd gnd cell_6t
Xbit_r200_c96 bl[96] br[96] wl[200] vdd gnd cell_6t
Xbit_r201_c96 bl[96] br[96] wl[201] vdd gnd cell_6t
Xbit_r202_c96 bl[96] br[96] wl[202] vdd gnd cell_6t
Xbit_r203_c96 bl[96] br[96] wl[203] vdd gnd cell_6t
Xbit_r204_c96 bl[96] br[96] wl[204] vdd gnd cell_6t
Xbit_r205_c96 bl[96] br[96] wl[205] vdd gnd cell_6t
Xbit_r206_c96 bl[96] br[96] wl[206] vdd gnd cell_6t
Xbit_r207_c96 bl[96] br[96] wl[207] vdd gnd cell_6t
Xbit_r208_c96 bl[96] br[96] wl[208] vdd gnd cell_6t
Xbit_r209_c96 bl[96] br[96] wl[209] vdd gnd cell_6t
Xbit_r210_c96 bl[96] br[96] wl[210] vdd gnd cell_6t
Xbit_r211_c96 bl[96] br[96] wl[211] vdd gnd cell_6t
Xbit_r212_c96 bl[96] br[96] wl[212] vdd gnd cell_6t
Xbit_r213_c96 bl[96] br[96] wl[213] vdd gnd cell_6t
Xbit_r214_c96 bl[96] br[96] wl[214] vdd gnd cell_6t
Xbit_r215_c96 bl[96] br[96] wl[215] vdd gnd cell_6t
Xbit_r216_c96 bl[96] br[96] wl[216] vdd gnd cell_6t
Xbit_r217_c96 bl[96] br[96] wl[217] vdd gnd cell_6t
Xbit_r218_c96 bl[96] br[96] wl[218] vdd gnd cell_6t
Xbit_r219_c96 bl[96] br[96] wl[219] vdd gnd cell_6t
Xbit_r220_c96 bl[96] br[96] wl[220] vdd gnd cell_6t
Xbit_r221_c96 bl[96] br[96] wl[221] vdd gnd cell_6t
Xbit_r222_c96 bl[96] br[96] wl[222] vdd gnd cell_6t
Xbit_r223_c96 bl[96] br[96] wl[223] vdd gnd cell_6t
Xbit_r224_c96 bl[96] br[96] wl[224] vdd gnd cell_6t
Xbit_r225_c96 bl[96] br[96] wl[225] vdd gnd cell_6t
Xbit_r226_c96 bl[96] br[96] wl[226] vdd gnd cell_6t
Xbit_r227_c96 bl[96] br[96] wl[227] vdd gnd cell_6t
Xbit_r228_c96 bl[96] br[96] wl[228] vdd gnd cell_6t
Xbit_r229_c96 bl[96] br[96] wl[229] vdd gnd cell_6t
Xbit_r230_c96 bl[96] br[96] wl[230] vdd gnd cell_6t
Xbit_r231_c96 bl[96] br[96] wl[231] vdd gnd cell_6t
Xbit_r232_c96 bl[96] br[96] wl[232] vdd gnd cell_6t
Xbit_r233_c96 bl[96] br[96] wl[233] vdd gnd cell_6t
Xbit_r234_c96 bl[96] br[96] wl[234] vdd gnd cell_6t
Xbit_r235_c96 bl[96] br[96] wl[235] vdd gnd cell_6t
Xbit_r236_c96 bl[96] br[96] wl[236] vdd gnd cell_6t
Xbit_r237_c96 bl[96] br[96] wl[237] vdd gnd cell_6t
Xbit_r238_c96 bl[96] br[96] wl[238] vdd gnd cell_6t
Xbit_r239_c96 bl[96] br[96] wl[239] vdd gnd cell_6t
Xbit_r240_c96 bl[96] br[96] wl[240] vdd gnd cell_6t
Xbit_r241_c96 bl[96] br[96] wl[241] vdd gnd cell_6t
Xbit_r242_c96 bl[96] br[96] wl[242] vdd gnd cell_6t
Xbit_r243_c96 bl[96] br[96] wl[243] vdd gnd cell_6t
Xbit_r244_c96 bl[96] br[96] wl[244] vdd gnd cell_6t
Xbit_r245_c96 bl[96] br[96] wl[245] vdd gnd cell_6t
Xbit_r246_c96 bl[96] br[96] wl[246] vdd gnd cell_6t
Xbit_r247_c96 bl[96] br[96] wl[247] vdd gnd cell_6t
Xbit_r248_c96 bl[96] br[96] wl[248] vdd gnd cell_6t
Xbit_r249_c96 bl[96] br[96] wl[249] vdd gnd cell_6t
Xbit_r250_c96 bl[96] br[96] wl[250] vdd gnd cell_6t
Xbit_r251_c96 bl[96] br[96] wl[251] vdd gnd cell_6t
Xbit_r252_c96 bl[96] br[96] wl[252] vdd gnd cell_6t
Xbit_r253_c96 bl[96] br[96] wl[253] vdd gnd cell_6t
Xbit_r254_c96 bl[96] br[96] wl[254] vdd gnd cell_6t
Xbit_r255_c96 bl[96] br[96] wl[255] vdd gnd cell_6t
Xbit_r256_c96 bl[96] br[96] wl[256] vdd gnd cell_6t
Xbit_r257_c96 bl[96] br[96] wl[257] vdd gnd cell_6t
Xbit_r258_c96 bl[96] br[96] wl[258] vdd gnd cell_6t
Xbit_r259_c96 bl[96] br[96] wl[259] vdd gnd cell_6t
Xbit_r260_c96 bl[96] br[96] wl[260] vdd gnd cell_6t
Xbit_r261_c96 bl[96] br[96] wl[261] vdd gnd cell_6t
Xbit_r262_c96 bl[96] br[96] wl[262] vdd gnd cell_6t
Xbit_r263_c96 bl[96] br[96] wl[263] vdd gnd cell_6t
Xbit_r264_c96 bl[96] br[96] wl[264] vdd gnd cell_6t
Xbit_r265_c96 bl[96] br[96] wl[265] vdd gnd cell_6t
Xbit_r266_c96 bl[96] br[96] wl[266] vdd gnd cell_6t
Xbit_r267_c96 bl[96] br[96] wl[267] vdd gnd cell_6t
Xbit_r268_c96 bl[96] br[96] wl[268] vdd gnd cell_6t
Xbit_r269_c96 bl[96] br[96] wl[269] vdd gnd cell_6t
Xbit_r270_c96 bl[96] br[96] wl[270] vdd gnd cell_6t
Xbit_r271_c96 bl[96] br[96] wl[271] vdd gnd cell_6t
Xbit_r272_c96 bl[96] br[96] wl[272] vdd gnd cell_6t
Xbit_r273_c96 bl[96] br[96] wl[273] vdd gnd cell_6t
Xbit_r274_c96 bl[96] br[96] wl[274] vdd gnd cell_6t
Xbit_r275_c96 bl[96] br[96] wl[275] vdd gnd cell_6t
Xbit_r276_c96 bl[96] br[96] wl[276] vdd gnd cell_6t
Xbit_r277_c96 bl[96] br[96] wl[277] vdd gnd cell_6t
Xbit_r278_c96 bl[96] br[96] wl[278] vdd gnd cell_6t
Xbit_r279_c96 bl[96] br[96] wl[279] vdd gnd cell_6t
Xbit_r280_c96 bl[96] br[96] wl[280] vdd gnd cell_6t
Xbit_r281_c96 bl[96] br[96] wl[281] vdd gnd cell_6t
Xbit_r282_c96 bl[96] br[96] wl[282] vdd gnd cell_6t
Xbit_r283_c96 bl[96] br[96] wl[283] vdd gnd cell_6t
Xbit_r284_c96 bl[96] br[96] wl[284] vdd gnd cell_6t
Xbit_r285_c96 bl[96] br[96] wl[285] vdd gnd cell_6t
Xbit_r286_c96 bl[96] br[96] wl[286] vdd gnd cell_6t
Xbit_r287_c96 bl[96] br[96] wl[287] vdd gnd cell_6t
Xbit_r288_c96 bl[96] br[96] wl[288] vdd gnd cell_6t
Xbit_r289_c96 bl[96] br[96] wl[289] vdd gnd cell_6t
Xbit_r290_c96 bl[96] br[96] wl[290] vdd gnd cell_6t
Xbit_r291_c96 bl[96] br[96] wl[291] vdd gnd cell_6t
Xbit_r292_c96 bl[96] br[96] wl[292] vdd gnd cell_6t
Xbit_r293_c96 bl[96] br[96] wl[293] vdd gnd cell_6t
Xbit_r294_c96 bl[96] br[96] wl[294] vdd gnd cell_6t
Xbit_r295_c96 bl[96] br[96] wl[295] vdd gnd cell_6t
Xbit_r296_c96 bl[96] br[96] wl[296] vdd gnd cell_6t
Xbit_r297_c96 bl[96] br[96] wl[297] vdd gnd cell_6t
Xbit_r298_c96 bl[96] br[96] wl[298] vdd gnd cell_6t
Xbit_r299_c96 bl[96] br[96] wl[299] vdd gnd cell_6t
Xbit_r300_c96 bl[96] br[96] wl[300] vdd gnd cell_6t
Xbit_r301_c96 bl[96] br[96] wl[301] vdd gnd cell_6t
Xbit_r302_c96 bl[96] br[96] wl[302] vdd gnd cell_6t
Xbit_r303_c96 bl[96] br[96] wl[303] vdd gnd cell_6t
Xbit_r304_c96 bl[96] br[96] wl[304] vdd gnd cell_6t
Xbit_r305_c96 bl[96] br[96] wl[305] vdd gnd cell_6t
Xbit_r306_c96 bl[96] br[96] wl[306] vdd gnd cell_6t
Xbit_r307_c96 bl[96] br[96] wl[307] vdd gnd cell_6t
Xbit_r308_c96 bl[96] br[96] wl[308] vdd gnd cell_6t
Xbit_r309_c96 bl[96] br[96] wl[309] vdd gnd cell_6t
Xbit_r310_c96 bl[96] br[96] wl[310] vdd gnd cell_6t
Xbit_r311_c96 bl[96] br[96] wl[311] vdd gnd cell_6t
Xbit_r312_c96 bl[96] br[96] wl[312] vdd gnd cell_6t
Xbit_r313_c96 bl[96] br[96] wl[313] vdd gnd cell_6t
Xbit_r314_c96 bl[96] br[96] wl[314] vdd gnd cell_6t
Xbit_r315_c96 bl[96] br[96] wl[315] vdd gnd cell_6t
Xbit_r316_c96 bl[96] br[96] wl[316] vdd gnd cell_6t
Xbit_r317_c96 bl[96] br[96] wl[317] vdd gnd cell_6t
Xbit_r318_c96 bl[96] br[96] wl[318] vdd gnd cell_6t
Xbit_r319_c96 bl[96] br[96] wl[319] vdd gnd cell_6t
Xbit_r320_c96 bl[96] br[96] wl[320] vdd gnd cell_6t
Xbit_r321_c96 bl[96] br[96] wl[321] vdd gnd cell_6t
Xbit_r322_c96 bl[96] br[96] wl[322] vdd gnd cell_6t
Xbit_r323_c96 bl[96] br[96] wl[323] vdd gnd cell_6t
Xbit_r324_c96 bl[96] br[96] wl[324] vdd gnd cell_6t
Xbit_r325_c96 bl[96] br[96] wl[325] vdd gnd cell_6t
Xbit_r326_c96 bl[96] br[96] wl[326] vdd gnd cell_6t
Xbit_r327_c96 bl[96] br[96] wl[327] vdd gnd cell_6t
Xbit_r328_c96 bl[96] br[96] wl[328] vdd gnd cell_6t
Xbit_r329_c96 bl[96] br[96] wl[329] vdd gnd cell_6t
Xbit_r330_c96 bl[96] br[96] wl[330] vdd gnd cell_6t
Xbit_r331_c96 bl[96] br[96] wl[331] vdd gnd cell_6t
Xbit_r332_c96 bl[96] br[96] wl[332] vdd gnd cell_6t
Xbit_r333_c96 bl[96] br[96] wl[333] vdd gnd cell_6t
Xbit_r334_c96 bl[96] br[96] wl[334] vdd gnd cell_6t
Xbit_r335_c96 bl[96] br[96] wl[335] vdd gnd cell_6t
Xbit_r336_c96 bl[96] br[96] wl[336] vdd gnd cell_6t
Xbit_r337_c96 bl[96] br[96] wl[337] vdd gnd cell_6t
Xbit_r338_c96 bl[96] br[96] wl[338] vdd gnd cell_6t
Xbit_r339_c96 bl[96] br[96] wl[339] vdd gnd cell_6t
Xbit_r340_c96 bl[96] br[96] wl[340] vdd gnd cell_6t
Xbit_r341_c96 bl[96] br[96] wl[341] vdd gnd cell_6t
Xbit_r342_c96 bl[96] br[96] wl[342] vdd gnd cell_6t
Xbit_r343_c96 bl[96] br[96] wl[343] vdd gnd cell_6t
Xbit_r344_c96 bl[96] br[96] wl[344] vdd gnd cell_6t
Xbit_r345_c96 bl[96] br[96] wl[345] vdd gnd cell_6t
Xbit_r346_c96 bl[96] br[96] wl[346] vdd gnd cell_6t
Xbit_r347_c96 bl[96] br[96] wl[347] vdd gnd cell_6t
Xbit_r348_c96 bl[96] br[96] wl[348] vdd gnd cell_6t
Xbit_r349_c96 bl[96] br[96] wl[349] vdd gnd cell_6t
Xbit_r350_c96 bl[96] br[96] wl[350] vdd gnd cell_6t
Xbit_r351_c96 bl[96] br[96] wl[351] vdd gnd cell_6t
Xbit_r352_c96 bl[96] br[96] wl[352] vdd gnd cell_6t
Xbit_r353_c96 bl[96] br[96] wl[353] vdd gnd cell_6t
Xbit_r354_c96 bl[96] br[96] wl[354] vdd gnd cell_6t
Xbit_r355_c96 bl[96] br[96] wl[355] vdd gnd cell_6t
Xbit_r356_c96 bl[96] br[96] wl[356] vdd gnd cell_6t
Xbit_r357_c96 bl[96] br[96] wl[357] vdd gnd cell_6t
Xbit_r358_c96 bl[96] br[96] wl[358] vdd gnd cell_6t
Xbit_r359_c96 bl[96] br[96] wl[359] vdd gnd cell_6t
Xbit_r360_c96 bl[96] br[96] wl[360] vdd gnd cell_6t
Xbit_r361_c96 bl[96] br[96] wl[361] vdd gnd cell_6t
Xbit_r362_c96 bl[96] br[96] wl[362] vdd gnd cell_6t
Xbit_r363_c96 bl[96] br[96] wl[363] vdd gnd cell_6t
Xbit_r364_c96 bl[96] br[96] wl[364] vdd gnd cell_6t
Xbit_r365_c96 bl[96] br[96] wl[365] vdd gnd cell_6t
Xbit_r366_c96 bl[96] br[96] wl[366] vdd gnd cell_6t
Xbit_r367_c96 bl[96] br[96] wl[367] vdd gnd cell_6t
Xbit_r368_c96 bl[96] br[96] wl[368] vdd gnd cell_6t
Xbit_r369_c96 bl[96] br[96] wl[369] vdd gnd cell_6t
Xbit_r370_c96 bl[96] br[96] wl[370] vdd gnd cell_6t
Xbit_r371_c96 bl[96] br[96] wl[371] vdd gnd cell_6t
Xbit_r372_c96 bl[96] br[96] wl[372] vdd gnd cell_6t
Xbit_r373_c96 bl[96] br[96] wl[373] vdd gnd cell_6t
Xbit_r374_c96 bl[96] br[96] wl[374] vdd gnd cell_6t
Xbit_r375_c96 bl[96] br[96] wl[375] vdd gnd cell_6t
Xbit_r376_c96 bl[96] br[96] wl[376] vdd gnd cell_6t
Xbit_r377_c96 bl[96] br[96] wl[377] vdd gnd cell_6t
Xbit_r378_c96 bl[96] br[96] wl[378] vdd gnd cell_6t
Xbit_r379_c96 bl[96] br[96] wl[379] vdd gnd cell_6t
Xbit_r380_c96 bl[96] br[96] wl[380] vdd gnd cell_6t
Xbit_r381_c96 bl[96] br[96] wl[381] vdd gnd cell_6t
Xbit_r382_c96 bl[96] br[96] wl[382] vdd gnd cell_6t
Xbit_r383_c96 bl[96] br[96] wl[383] vdd gnd cell_6t
Xbit_r384_c96 bl[96] br[96] wl[384] vdd gnd cell_6t
Xbit_r385_c96 bl[96] br[96] wl[385] vdd gnd cell_6t
Xbit_r386_c96 bl[96] br[96] wl[386] vdd gnd cell_6t
Xbit_r387_c96 bl[96] br[96] wl[387] vdd gnd cell_6t
Xbit_r388_c96 bl[96] br[96] wl[388] vdd gnd cell_6t
Xbit_r389_c96 bl[96] br[96] wl[389] vdd gnd cell_6t
Xbit_r390_c96 bl[96] br[96] wl[390] vdd gnd cell_6t
Xbit_r391_c96 bl[96] br[96] wl[391] vdd gnd cell_6t
Xbit_r392_c96 bl[96] br[96] wl[392] vdd gnd cell_6t
Xbit_r393_c96 bl[96] br[96] wl[393] vdd gnd cell_6t
Xbit_r394_c96 bl[96] br[96] wl[394] vdd gnd cell_6t
Xbit_r395_c96 bl[96] br[96] wl[395] vdd gnd cell_6t
Xbit_r396_c96 bl[96] br[96] wl[396] vdd gnd cell_6t
Xbit_r397_c96 bl[96] br[96] wl[397] vdd gnd cell_6t
Xbit_r398_c96 bl[96] br[96] wl[398] vdd gnd cell_6t
Xbit_r399_c96 bl[96] br[96] wl[399] vdd gnd cell_6t
Xbit_r400_c96 bl[96] br[96] wl[400] vdd gnd cell_6t
Xbit_r401_c96 bl[96] br[96] wl[401] vdd gnd cell_6t
Xbit_r402_c96 bl[96] br[96] wl[402] vdd gnd cell_6t
Xbit_r403_c96 bl[96] br[96] wl[403] vdd gnd cell_6t
Xbit_r404_c96 bl[96] br[96] wl[404] vdd gnd cell_6t
Xbit_r405_c96 bl[96] br[96] wl[405] vdd gnd cell_6t
Xbit_r406_c96 bl[96] br[96] wl[406] vdd gnd cell_6t
Xbit_r407_c96 bl[96] br[96] wl[407] vdd gnd cell_6t
Xbit_r408_c96 bl[96] br[96] wl[408] vdd gnd cell_6t
Xbit_r409_c96 bl[96] br[96] wl[409] vdd gnd cell_6t
Xbit_r410_c96 bl[96] br[96] wl[410] vdd gnd cell_6t
Xbit_r411_c96 bl[96] br[96] wl[411] vdd gnd cell_6t
Xbit_r412_c96 bl[96] br[96] wl[412] vdd gnd cell_6t
Xbit_r413_c96 bl[96] br[96] wl[413] vdd gnd cell_6t
Xbit_r414_c96 bl[96] br[96] wl[414] vdd gnd cell_6t
Xbit_r415_c96 bl[96] br[96] wl[415] vdd gnd cell_6t
Xbit_r416_c96 bl[96] br[96] wl[416] vdd gnd cell_6t
Xbit_r417_c96 bl[96] br[96] wl[417] vdd gnd cell_6t
Xbit_r418_c96 bl[96] br[96] wl[418] vdd gnd cell_6t
Xbit_r419_c96 bl[96] br[96] wl[419] vdd gnd cell_6t
Xbit_r420_c96 bl[96] br[96] wl[420] vdd gnd cell_6t
Xbit_r421_c96 bl[96] br[96] wl[421] vdd gnd cell_6t
Xbit_r422_c96 bl[96] br[96] wl[422] vdd gnd cell_6t
Xbit_r423_c96 bl[96] br[96] wl[423] vdd gnd cell_6t
Xbit_r424_c96 bl[96] br[96] wl[424] vdd gnd cell_6t
Xbit_r425_c96 bl[96] br[96] wl[425] vdd gnd cell_6t
Xbit_r426_c96 bl[96] br[96] wl[426] vdd gnd cell_6t
Xbit_r427_c96 bl[96] br[96] wl[427] vdd gnd cell_6t
Xbit_r428_c96 bl[96] br[96] wl[428] vdd gnd cell_6t
Xbit_r429_c96 bl[96] br[96] wl[429] vdd gnd cell_6t
Xbit_r430_c96 bl[96] br[96] wl[430] vdd gnd cell_6t
Xbit_r431_c96 bl[96] br[96] wl[431] vdd gnd cell_6t
Xbit_r432_c96 bl[96] br[96] wl[432] vdd gnd cell_6t
Xbit_r433_c96 bl[96] br[96] wl[433] vdd gnd cell_6t
Xbit_r434_c96 bl[96] br[96] wl[434] vdd gnd cell_6t
Xbit_r435_c96 bl[96] br[96] wl[435] vdd gnd cell_6t
Xbit_r436_c96 bl[96] br[96] wl[436] vdd gnd cell_6t
Xbit_r437_c96 bl[96] br[96] wl[437] vdd gnd cell_6t
Xbit_r438_c96 bl[96] br[96] wl[438] vdd gnd cell_6t
Xbit_r439_c96 bl[96] br[96] wl[439] vdd gnd cell_6t
Xbit_r440_c96 bl[96] br[96] wl[440] vdd gnd cell_6t
Xbit_r441_c96 bl[96] br[96] wl[441] vdd gnd cell_6t
Xbit_r442_c96 bl[96] br[96] wl[442] vdd gnd cell_6t
Xbit_r443_c96 bl[96] br[96] wl[443] vdd gnd cell_6t
Xbit_r444_c96 bl[96] br[96] wl[444] vdd gnd cell_6t
Xbit_r445_c96 bl[96] br[96] wl[445] vdd gnd cell_6t
Xbit_r446_c96 bl[96] br[96] wl[446] vdd gnd cell_6t
Xbit_r447_c96 bl[96] br[96] wl[447] vdd gnd cell_6t
Xbit_r448_c96 bl[96] br[96] wl[448] vdd gnd cell_6t
Xbit_r449_c96 bl[96] br[96] wl[449] vdd gnd cell_6t
Xbit_r450_c96 bl[96] br[96] wl[450] vdd gnd cell_6t
Xbit_r451_c96 bl[96] br[96] wl[451] vdd gnd cell_6t
Xbit_r452_c96 bl[96] br[96] wl[452] vdd gnd cell_6t
Xbit_r453_c96 bl[96] br[96] wl[453] vdd gnd cell_6t
Xbit_r454_c96 bl[96] br[96] wl[454] vdd gnd cell_6t
Xbit_r455_c96 bl[96] br[96] wl[455] vdd gnd cell_6t
Xbit_r456_c96 bl[96] br[96] wl[456] vdd gnd cell_6t
Xbit_r457_c96 bl[96] br[96] wl[457] vdd gnd cell_6t
Xbit_r458_c96 bl[96] br[96] wl[458] vdd gnd cell_6t
Xbit_r459_c96 bl[96] br[96] wl[459] vdd gnd cell_6t
Xbit_r460_c96 bl[96] br[96] wl[460] vdd gnd cell_6t
Xbit_r461_c96 bl[96] br[96] wl[461] vdd gnd cell_6t
Xbit_r462_c96 bl[96] br[96] wl[462] vdd gnd cell_6t
Xbit_r463_c96 bl[96] br[96] wl[463] vdd gnd cell_6t
Xbit_r464_c96 bl[96] br[96] wl[464] vdd gnd cell_6t
Xbit_r465_c96 bl[96] br[96] wl[465] vdd gnd cell_6t
Xbit_r466_c96 bl[96] br[96] wl[466] vdd gnd cell_6t
Xbit_r467_c96 bl[96] br[96] wl[467] vdd gnd cell_6t
Xbit_r468_c96 bl[96] br[96] wl[468] vdd gnd cell_6t
Xbit_r469_c96 bl[96] br[96] wl[469] vdd gnd cell_6t
Xbit_r470_c96 bl[96] br[96] wl[470] vdd gnd cell_6t
Xbit_r471_c96 bl[96] br[96] wl[471] vdd gnd cell_6t
Xbit_r472_c96 bl[96] br[96] wl[472] vdd gnd cell_6t
Xbit_r473_c96 bl[96] br[96] wl[473] vdd gnd cell_6t
Xbit_r474_c96 bl[96] br[96] wl[474] vdd gnd cell_6t
Xbit_r475_c96 bl[96] br[96] wl[475] vdd gnd cell_6t
Xbit_r476_c96 bl[96] br[96] wl[476] vdd gnd cell_6t
Xbit_r477_c96 bl[96] br[96] wl[477] vdd gnd cell_6t
Xbit_r478_c96 bl[96] br[96] wl[478] vdd gnd cell_6t
Xbit_r479_c96 bl[96] br[96] wl[479] vdd gnd cell_6t
Xbit_r480_c96 bl[96] br[96] wl[480] vdd gnd cell_6t
Xbit_r481_c96 bl[96] br[96] wl[481] vdd gnd cell_6t
Xbit_r482_c96 bl[96] br[96] wl[482] vdd gnd cell_6t
Xbit_r483_c96 bl[96] br[96] wl[483] vdd gnd cell_6t
Xbit_r484_c96 bl[96] br[96] wl[484] vdd gnd cell_6t
Xbit_r485_c96 bl[96] br[96] wl[485] vdd gnd cell_6t
Xbit_r486_c96 bl[96] br[96] wl[486] vdd gnd cell_6t
Xbit_r487_c96 bl[96] br[96] wl[487] vdd gnd cell_6t
Xbit_r488_c96 bl[96] br[96] wl[488] vdd gnd cell_6t
Xbit_r489_c96 bl[96] br[96] wl[489] vdd gnd cell_6t
Xbit_r490_c96 bl[96] br[96] wl[490] vdd gnd cell_6t
Xbit_r491_c96 bl[96] br[96] wl[491] vdd gnd cell_6t
Xbit_r492_c96 bl[96] br[96] wl[492] vdd gnd cell_6t
Xbit_r493_c96 bl[96] br[96] wl[493] vdd gnd cell_6t
Xbit_r494_c96 bl[96] br[96] wl[494] vdd gnd cell_6t
Xbit_r495_c96 bl[96] br[96] wl[495] vdd gnd cell_6t
Xbit_r496_c96 bl[96] br[96] wl[496] vdd gnd cell_6t
Xbit_r497_c96 bl[96] br[96] wl[497] vdd gnd cell_6t
Xbit_r498_c96 bl[96] br[96] wl[498] vdd gnd cell_6t
Xbit_r499_c96 bl[96] br[96] wl[499] vdd gnd cell_6t
Xbit_r500_c96 bl[96] br[96] wl[500] vdd gnd cell_6t
Xbit_r501_c96 bl[96] br[96] wl[501] vdd gnd cell_6t
Xbit_r502_c96 bl[96] br[96] wl[502] vdd gnd cell_6t
Xbit_r503_c96 bl[96] br[96] wl[503] vdd gnd cell_6t
Xbit_r504_c96 bl[96] br[96] wl[504] vdd gnd cell_6t
Xbit_r505_c96 bl[96] br[96] wl[505] vdd gnd cell_6t
Xbit_r506_c96 bl[96] br[96] wl[506] vdd gnd cell_6t
Xbit_r507_c96 bl[96] br[96] wl[507] vdd gnd cell_6t
Xbit_r508_c96 bl[96] br[96] wl[508] vdd gnd cell_6t
Xbit_r509_c96 bl[96] br[96] wl[509] vdd gnd cell_6t
Xbit_r510_c96 bl[96] br[96] wl[510] vdd gnd cell_6t
Xbit_r511_c96 bl[96] br[96] wl[511] vdd gnd cell_6t
Xbit_r0_c97 bl[97] br[97] wl[0] vdd gnd cell_6t
Xbit_r1_c97 bl[97] br[97] wl[1] vdd gnd cell_6t
Xbit_r2_c97 bl[97] br[97] wl[2] vdd gnd cell_6t
Xbit_r3_c97 bl[97] br[97] wl[3] vdd gnd cell_6t
Xbit_r4_c97 bl[97] br[97] wl[4] vdd gnd cell_6t
Xbit_r5_c97 bl[97] br[97] wl[5] vdd gnd cell_6t
Xbit_r6_c97 bl[97] br[97] wl[6] vdd gnd cell_6t
Xbit_r7_c97 bl[97] br[97] wl[7] vdd gnd cell_6t
Xbit_r8_c97 bl[97] br[97] wl[8] vdd gnd cell_6t
Xbit_r9_c97 bl[97] br[97] wl[9] vdd gnd cell_6t
Xbit_r10_c97 bl[97] br[97] wl[10] vdd gnd cell_6t
Xbit_r11_c97 bl[97] br[97] wl[11] vdd gnd cell_6t
Xbit_r12_c97 bl[97] br[97] wl[12] vdd gnd cell_6t
Xbit_r13_c97 bl[97] br[97] wl[13] vdd gnd cell_6t
Xbit_r14_c97 bl[97] br[97] wl[14] vdd gnd cell_6t
Xbit_r15_c97 bl[97] br[97] wl[15] vdd gnd cell_6t
Xbit_r16_c97 bl[97] br[97] wl[16] vdd gnd cell_6t
Xbit_r17_c97 bl[97] br[97] wl[17] vdd gnd cell_6t
Xbit_r18_c97 bl[97] br[97] wl[18] vdd gnd cell_6t
Xbit_r19_c97 bl[97] br[97] wl[19] vdd gnd cell_6t
Xbit_r20_c97 bl[97] br[97] wl[20] vdd gnd cell_6t
Xbit_r21_c97 bl[97] br[97] wl[21] vdd gnd cell_6t
Xbit_r22_c97 bl[97] br[97] wl[22] vdd gnd cell_6t
Xbit_r23_c97 bl[97] br[97] wl[23] vdd gnd cell_6t
Xbit_r24_c97 bl[97] br[97] wl[24] vdd gnd cell_6t
Xbit_r25_c97 bl[97] br[97] wl[25] vdd gnd cell_6t
Xbit_r26_c97 bl[97] br[97] wl[26] vdd gnd cell_6t
Xbit_r27_c97 bl[97] br[97] wl[27] vdd gnd cell_6t
Xbit_r28_c97 bl[97] br[97] wl[28] vdd gnd cell_6t
Xbit_r29_c97 bl[97] br[97] wl[29] vdd gnd cell_6t
Xbit_r30_c97 bl[97] br[97] wl[30] vdd gnd cell_6t
Xbit_r31_c97 bl[97] br[97] wl[31] vdd gnd cell_6t
Xbit_r32_c97 bl[97] br[97] wl[32] vdd gnd cell_6t
Xbit_r33_c97 bl[97] br[97] wl[33] vdd gnd cell_6t
Xbit_r34_c97 bl[97] br[97] wl[34] vdd gnd cell_6t
Xbit_r35_c97 bl[97] br[97] wl[35] vdd gnd cell_6t
Xbit_r36_c97 bl[97] br[97] wl[36] vdd gnd cell_6t
Xbit_r37_c97 bl[97] br[97] wl[37] vdd gnd cell_6t
Xbit_r38_c97 bl[97] br[97] wl[38] vdd gnd cell_6t
Xbit_r39_c97 bl[97] br[97] wl[39] vdd gnd cell_6t
Xbit_r40_c97 bl[97] br[97] wl[40] vdd gnd cell_6t
Xbit_r41_c97 bl[97] br[97] wl[41] vdd gnd cell_6t
Xbit_r42_c97 bl[97] br[97] wl[42] vdd gnd cell_6t
Xbit_r43_c97 bl[97] br[97] wl[43] vdd gnd cell_6t
Xbit_r44_c97 bl[97] br[97] wl[44] vdd gnd cell_6t
Xbit_r45_c97 bl[97] br[97] wl[45] vdd gnd cell_6t
Xbit_r46_c97 bl[97] br[97] wl[46] vdd gnd cell_6t
Xbit_r47_c97 bl[97] br[97] wl[47] vdd gnd cell_6t
Xbit_r48_c97 bl[97] br[97] wl[48] vdd gnd cell_6t
Xbit_r49_c97 bl[97] br[97] wl[49] vdd gnd cell_6t
Xbit_r50_c97 bl[97] br[97] wl[50] vdd gnd cell_6t
Xbit_r51_c97 bl[97] br[97] wl[51] vdd gnd cell_6t
Xbit_r52_c97 bl[97] br[97] wl[52] vdd gnd cell_6t
Xbit_r53_c97 bl[97] br[97] wl[53] vdd gnd cell_6t
Xbit_r54_c97 bl[97] br[97] wl[54] vdd gnd cell_6t
Xbit_r55_c97 bl[97] br[97] wl[55] vdd gnd cell_6t
Xbit_r56_c97 bl[97] br[97] wl[56] vdd gnd cell_6t
Xbit_r57_c97 bl[97] br[97] wl[57] vdd gnd cell_6t
Xbit_r58_c97 bl[97] br[97] wl[58] vdd gnd cell_6t
Xbit_r59_c97 bl[97] br[97] wl[59] vdd gnd cell_6t
Xbit_r60_c97 bl[97] br[97] wl[60] vdd gnd cell_6t
Xbit_r61_c97 bl[97] br[97] wl[61] vdd gnd cell_6t
Xbit_r62_c97 bl[97] br[97] wl[62] vdd gnd cell_6t
Xbit_r63_c97 bl[97] br[97] wl[63] vdd gnd cell_6t
Xbit_r64_c97 bl[97] br[97] wl[64] vdd gnd cell_6t
Xbit_r65_c97 bl[97] br[97] wl[65] vdd gnd cell_6t
Xbit_r66_c97 bl[97] br[97] wl[66] vdd gnd cell_6t
Xbit_r67_c97 bl[97] br[97] wl[67] vdd gnd cell_6t
Xbit_r68_c97 bl[97] br[97] wl[68] vdd gnd cell_6t
Xbit_r69_c97 bl[97] br[97] wl[69] vdd gnd cell_6t
Xbit_r70_c97 bl[97] br[97] wl[70] vdd gnd cell_6t
Xbit_r71_c97 bl[97] br[97] wl[71] vdd gnd cell_6t
Xbit_r72_c97 bl[97] br[97] wl[72] vdd gnd cell_6t
Xbit_r73_c97 bl[97] br[97] wl[73] vdd gnd cell_6t
Xbit_r74_c97 bl[97] br[97] wl[74] vdd gnd cell_6t
Xbit_r75_c97 bl[97] br[97] wl[75] vdd gnd cell_6t
Xbit_r76_c97 bl[97] br[97] wl[76] vdd gnd cell_6t
Xbit_r77_c97 bl[97] br[97] wl[77] vdd gnd cell_6t
Xbit_r78_c97 bl[97] br[97] wl[78] vdd gnd cell_6t
Xbit_r79_c97 bl[97] br[97] wl[79] vdd gnd cell_6t
Xbit_r80_c97 bl[97] br[97] wl[80] vdd gnd cell_6t
Xbit_r81_c97 bl[97] br[97] wl[81] vdd gnd cell_6t
Xbit_r82_c97 bl[97] br[97] wl[82] vdd gnd cell_6t
Xbit_r83_c97 bl[97] br[97] wl[83] vdd gnd cell_6t
Xbit_r84_c97 bl[97] br[97] wl[84] vdd gnd cell_6t
Xbit_r85_c97 bl[97] br[97] wl[85] vdd gnd cell_6t
Xbit_r86_c97 bl[97] br[97] wl[86] vdd gnd cell_6t
Xbit_r87_c97 bl[97] br[97] wl[87] vdd gnd cell_6t
Xbit_r88_c97 bl[97] br[97] wl[88] vdd gnd cell_6t
Xbit_r89_c97 bl[97] br[97] wl[89] vdd gnd cell_6t
Xbit_r90_c97 bl[97] br[97] wl[90] vdd gnd cell_6t
Xbit_r91_c97 bl[97] br[97] wl[91] vdd gnd cell_6t
Xbit_r92_c97 bl[97] br[97] wl[92] vdd gnd cell_6t
Xbit_r93_c97 bl[97] br[97] wl[93] vdd gnd cell_6t
Xbit_r94_c97 bl[97] br[97] wl[94] vdd gnd cell_6t
Xbit_r95_c97 bl[97] br[97] wl[95] vdd gnd cell_6t
Xbit_r96_c97 bl[97] br[97] wl[96] vdd gnd cell_6t
Xbit_r97_c97 bl[97] br[97] wl[97] vdd gnd cell_6t
Xbit_r98_c97 bl[97] br[97] wl[98] vdd gnd cell_6t
Xbit_r99_c97 bl[97] br[97] wl[99] vdd gnd cell_6t
Xbit_r100_c97 bl[97] br[97] wl[100] vdd gnd cell_6t
Xbit_r101_c97 bl[97] br[97] wl[101] vdd gnd cell_6t
Xbit_r102_c97 bl[97] br[97] wl[102] vdd gnd cell_6t
Xbit_r103_c97 bl[97] br[97] wl[103] vdd gnd cell_6t
Xbit_r104_c97 bl[97] br[97] wl[104] vdd gnd cell_6t
Xbit_r105_c97 bl[97] br[97] wl[105] vdd gnd cell_6t
Xbit_r106_c97 bl[97] br[97] wl[106] vdd gnd cell_6t
Xbit_r107_c97 bl[97] br[97] wl[107] vdd gnd cell_6t
Xbit_r108_c97 bl[97] br[97] wl[108] vdd gnd cell_6t
Xbit_r109_c97 bl[97] br[97] wl[109] vdd gnd cell_6t
Xbit_r110_c97 bl[97] br[97] wl[110] vdd gnd cell_6t
Xbit_r111_c97 bl[97] br[97] wl[111] vdd gnd cell_6t
Xbit_r112_c97 bl[97] br[97] wl[112] vdd gnd cell_6t
Xbit_r113_c97 bl[97] br[97] wl[113] vdd gnd cell_6t
Xbit_r114_c97 bl[97] br[97] wl[114] vdd gnd cell_6t
Xbit_r115_c97 bl[97] br[97] wl[115] vdd gnd cell_6t
Xbit_r116_c97 bl[97] br[97] wl[116] vdd gnd cell_6t
Xbit_r117_c97 bl[97] br[97] wl[117] vdd gnd cell_6t
Xbit_r118_c97 bl[97] br[97] wl[118] vdd gnd cell_6t
Xbit_r119_c97 bl[97] br[97] wl[119] vdd gnd cell_6t
Xbit_r120_c97 bl[97] br[97] wl[120] vdd gnd cell_6t
Xbit_r121_c97 bl[97] br[97] wl[121] vdd gnd cell_6t
Xbit_r122_c97 bl[97] br[97] wl[122] vdd gnd cell_6t
Xbit_r123_c97 bl[97] br[97] wl[123] vdd gnd cell_6t
Xbit_r124_c97 bl[97] br[97] wl[124] vdd gnd cell_6t
Xbit_r125_c97 bl[97] br[97] wl[125] vdd gnd cell_6t
Xbit_r126_c97 bl[97] br[97] wl[126] vdd gnd cell_6t
Xbit_r127_c97 bl[97] br[97] wl[127] vdd gnd cell_6t
Xbit_r128_c97 bl[97] br[97] wl[128] vdd gnd cell_6t
Xbit_r129_c97 bl[97] br[97] wl[129] vdd gnd cell_6t
Xbit_r130_c97 bl[97] br[97] wl[130] vdd gnd cell_6t
Xbit_r131_c97 bl[97] br[97] wl[131] vdd gnd cell_6t
Xbit_r132_c97 bl[97] br[97] wl[132] vdd gnd cell_6t
Xbit_r133_c97 bl[97] br[97] wl[133] vdd gnd cell_6t
Xbit_r134_c97 bl[97] br[97] wl[134] vdd gnd cell_6t
Xbit_r135_c97 bl[97] br[97] wl[135] vdd gnd cell_6t
Xbit_r136_c97 bl[97] br[97] wl[136] vdd gnd cell_6t
Xbit_r137_c97 bl[97] br[97] wl[137] vdd gnd cell_6t
Xbit_r138_c97 bl[97] br[97] wl[138] vdd gnd cell_6t
Xbit_r139_c97 bl[97] br[97] wl[139] vdd gnd cell_6t
Xbit_r140_c97 bl[97] br[97] wl[140] vdd gnd cell_6t
Xbit_r141_c97 bl[97] br[97] wl[141] vdd gnd cell_6t
Xbit_r142_c97 bl[97] br[97] wl[142] vdd gnd cell_6t
Xbit_r143_c97 bl[97] br[97] wl[143] vdd gnd cell_6t
Xbit_r144_c97 bl[97] br[97] wl[144] vdd gnd cell_6t
Xbit_r145_c97 bl[97] br[97] wl[145] vdd gnd cell_6t
Xbit_r146_c97 bl[97] br[97] wl[146] vdd gnd cell_6t
Xbit_r147_c97 bl[97] br[97] wl[147] vdd gnd cell_6t
Xbit_r148_c97 bl[97] br[97] wl[148] vdd gnd cell_6t
Xbit_r149_c97 bl[97] br[97] wl[149] vdd gnd cell_6t
Xbit_r150_c97 bl[97] br[97] wl[150] vdd gnd cell_6t
Xbit_r151_c97 bl[97] br[97] wl[151] vdd gnd cell_6t
Xbit_r152_c97 bl[97] br[97] wl[152] vdd gnd cell_6t
Xbit_r153_c97 bl[97] br[97] wl[153] vdd gnd cell_6t
Xbit_r154_c97 bl[97] br[97] wl[154] vdd gnd cell_6t
Xbit_r155_c97 bl[97] br[97] wl[155] vdd gnd cell_6t
Xbit_r156_c97 bl[97] br[97] wl[156] vdd gnd cell_6t
Xbit_r157_c97 bl[97] br[97] wl[157] vdd gnd cell_6t
Xbit_r158_c97 bl[97] br[97] wl[158] vdd gnd cell_6t
Xbit_r159_c97 bl[97] br[97] wl[159] vdd gnd cell_6t
Xbit_r160_c97 bl[97] br[97] wl[160] vdd gnd cell_6t
Xbit_r161_c97 bl[97] br[97] wl[161] vdd gnd cell_6t
Xbit_r162_c97 bl[97] br[97] wl[162] vdd gnd cell_6t
Xbit_r163_c97 bl[97] br[97] wl[163] vdd gnd cell_6t
Xbit_r164_c97 bl[97] br[97] wl[164] vdd gnd cell_6t
Xbit_r165_c97 bl[97] br[97] wl[165] vdd gnd cell_6t
Xbit_r166_c97 bl[97] br[97] wl[166] vdd gnd cell_6t
Xbit_r167_c97 bl[97] br[97] wl[167] vdd gnd cell_6t
Xbit_r168_c97 bl[97] br[97] wl[168] vdd gnd cell_6t
Xbit_r169_c97 bl[97] br[97] wl[169] vdd gnd cell_6t
Xbit_r170_c97 bl[97] br[97] wl[170] vdd gnd cell_6t
Xbit_r171_c97 bl[97] br[97] wl[171] vdd gnd cell_6t
Xbit_r172_c97 bl[97] br[97] wl[172] vdd gnd cell_6t
Xbit_r173_c97 bl[97] br[97] wl[173] vdd gnd cell_6t
Xbit_r174_c97 bl[97] br[97] wl[174] vdd gnd cell_6t
Xbit_r175_c97 bl[97] br[97] wl[175] vdd gnd cell_6t
Xbit_r176_c97 bl[97] br[97] wl[176] vdd gnd cell_6t
Xbit_r177_c97 bl[97] br[97] wl[177] vdd gnd cell_6t
Xbit_r178_c97 bl[97] br[97] wl[178] vdd gnd cell_6t
Xbit_r179_c97 bl[97] br[97] wl[179] vdd gnd cell_6t
Xbit_r180_c97 bl[97] br[97] wl[180] vdd gnd cell_6t
Xbit_r181_c97 bl[97] br[97] wl[181] vdd gnd cell_6t
Xbit_r182_c97 bl[97] br[97] wl[182] vdd gnd cell_6t
Xbit_r183_c97 bl[97] br[97] wl[183] vdd gnd cell_6t
Xbit_r184_c97 bl[97] br[97] wl[184] vdd gnd cell_6t
Xbit_r185_c97 bl[97] br[97] wl[185] vdd gnd cell_6t
Xbit_r186_c97 bl[97] br[97] wl[186] vdd gnd cell_6t
Xbit_r187_c97 bl[97] br[97] wl[187] vdd gnd cell_6t
Xbit_r188_c97 bl[97] br[97] wl[188] vdd gnd cell_6t
Xbit_r189_c97 bl[97] br[97] wl[189] vdd gnd cell_6t
Xbit_r190_c97 bl[97] br[97] wl[190] vdd gnd cell_6t
Xbit_r191_c97 bl[97] br[97] wl[191] vdd gnd cell_6t
Xbit_r192_c97 bl[97] br[97] wl[192] vdd gnd cell_6t
Xbit_r193_c97 bl[97] br[97] wl[193] vdd gnd cell_6t
Xbit_r194_c97 bl[97] br[97] wl[194] vdd gnd cell_6t
Xbit_r195_c97 bl[97] br[97] wl[195] vdd gnd cell_6t
Xbit_r196_c97 bl[97] br[97] wl[196] vdd gnd cell_6t
Xbit_r197_c97 bl[97] br[97] wl[197] vdd gnd cell_6t
Xbit_r198_c97 bl[97] br[97] wl[198] vdd gnd cell_6t
Xbit_r199_c97 bl[97] br[97] wl[199] vdd gnd cell_6t
Xbit_r200_c97 bl[97] br[97] wl[200] vdd gnd cell_6t
Xbit_r201_c97 bl[97] br[97] wl[201] vdd gnd cell_6t
Xbit_r202_c97 bl[97] br[97] wl[202] vdd gnd cell_6t
Xbit_r203_c97 bl[97] br[97] wl[203] vdd gnd cell_6t
Xbit_r204_c97 bl[97] br[97] wl[204] vdd gnd cell_6t
Xbit_r205_c97 bl[97] br[97] wl[205] vdd gnd cell_6t
Xbit_r206_c97 bl[97] br[97] wl[206] vdd gnd cell_6t
Xbit_r207_c97 bl[97] br[97] wl[207] vdd gnd cell_6t
Xbit_r208_c97 bl[97] br[97] wl[208] vdd gnd cell_6t
Xbit_r209_c97 bl[97] br[97] wl[209] vdd gnd cell_6t
Xbit_r210_c97 bl[97] br[97] wl[210] vdd gnd cell_6t
Xbit_r211_c97 bl[97] br[97] wl[211] vdd gnd cell_6t
Xbit_r212_c97 bl[97] br[97] wl[212] vdd gnd cell_6t
Xbit_r213_c97 bl[97] br[97] wl[213] vdd gnd cell_6t
Xbit_r214_c97 bl[97] br[97] wl[214] vdd gnd cell_6t
Xbit_r215_c97 bl[97] br[97] wl[215] vdd gnd cell_6t
Xbit_r216_c97 bl[97] br[97] wl[216] vdd gnd cell_6t
Xbit_r217_c97 bl[97] br[97] wl[217] vdd gnd cell_6t
Xbit_r218_c97 bl[97] br[97] wl[218] vdd gnd cell_6t
Xbit_r219_c97 bl[97] br[97] wl[219] vdd gnd cell_6t
Xbit_r220_c97 bl[97] br[97] wl[220] vdd gnd cell_6t
Xbit_r221_c97 bl[97] br[97] wl[221] vdd gnd cell_6t
Xbit_r222_c97 bl[97] br[97] wl[222] vdd gnd cell_6t
Xbit_r223_c97 bl[97] br[97] wl[223] vdd gnd cell_6t
Xbit_r224_c97 bl[97] br[97] wl[224] vdd gnd cell_6t
Xbit_r225_c97 bl[97] br[97] wl[225] vdd gnd cell_6t
Xbit_r226_c97 bl[97] br[97] wl[226] vdd gnd cell_6t
Xbit_r227_c97 bl[97] br[97] wl[227] vdd gnd cell_6t
Xbit_r228_c97 bl[97] br[97] wl[228] vdd gnd cell_6t
Xbit_r229_c97 bl[97] br[97] wl[229] vdd gnd cell_6t
Xbit_r230_c97 bl[97] br[97] wl[230] vdd gnd cell_6t
Xbit_r231_c97 bl[97] br[97] wl[231] vdd gnd cell_6t
Xbit_r232_c97 bl[97] br[97] wl[232] vdd gnd cell_6t
Xbit_r233_c97 bl[97] br[97] wl[233] vdd gnd cell_6t
Xbit_r234_c97 bl[97] br[97] wl[234] vdd gnd cell_6t
Xbit_r235_c97 bl[97] br[97] wl[235] vdd gnd cell_6t
Xbit_r236_c97 bl[97] br[97] wl[236] vdd gnd cell_6t
Xbit_r237_c97 bl[97] br[97] wl[237] vdd gnd cell_6t
Xbit_r238_c97 bl[97] br[97] wl[238] vdd gnd cell_6t
Xbit_r239_c97 bl[97] br[97] wl[239] vdd gnd cell_6t
Xbit_r240_c97 bl[97] br[97] wl[240] vdd gnd cell_6t
Xbit_r241_c97 bl[97] br[97] wl[241] vdd gnd cell_6t
Xbit_r242_c97 bl[97] br[97] wl[242] vdd gnd cell_6t
Xbit_r243_c97 bl[97] br[97] wl[243] vdd gnd cell_6t
Xbit_r244_c97 bl[97] br[97] wl[244] vdd gnd cell_6t
Xbit_r245_c97 bl[97] br[97] wl[245] vdd gnd cell_6t
Xbit_r246_c97 bl[97] br[97] wl[246] vdd gnd cell_6t
Xbit_r247_c97 bl[97] br[97] wl[247] vdd gnd cell_6t
Xbit_r248_c97 bl[97] br[97] wl[248] vdd gnd cell_6t
Xbit_r249_c97 bl[97] br[97] wl[249] vdd gnd cell_6t
Xbit_r250_c97 bl[97] br[97] wl[250] vdd gnd cell_6t
Xbit_r251_c97 bl[97] br[97] wl[251] vdd gnd cell_6t
Xbit_r252_c97 bl[97] br[97] wl[252] vdd gnd cell_6t
Xbit_r253_c97 bl[97] br[97] wl[253] vdd gnd cell_6t
Xbit_r254_c97 bl[97] br[97] wl[254] vdd gnd cell_6t
Xbit_r255_c97 bl[97] br[97] wl[255] vdd gnd cell_6t
Xbit_r256_c97 bl[97] br[97] wl[256] vdd gnd cell_6t
Xbit_r257_c97 bl[97] br[97] wl[257] vdd gnd cell_6t
Xbit_r258_c97 bl[97] br[97] wl[258] vdd gnd cell_6t
Xbit_r259_c97 bl[97] br[97] wl[259] vdd gnd cell_6t
Xbit_r260_c97 bl[97] br[97] wl[260] vdd gnd cell_6t
Xbit_r261_c97 bl[97] br[97] wl[261] vdd gnd cell_6t
Xbit_r262_c97 bl[97] br[97] wl[262] vdd gnd cell_6t
Xbit_r263_c97 bl[97] br[97] wl[263] vdd gnd cell_6t
Xbit_r264_c97 bl[97] br[97] wl[264] vdd gnd cell_6t
Xbit_r265_c97 bl[97] br[97] wl[265] vdd gnd cell_6t
Xbit_r266_c97 bl[97] br[97] wl[266] vdd gnd cell_6t
Xbit_r267_c97 bl[97] br[97] wl[267] vdd gnd cell_6t
Xbit_r268_c97 bl[97] br[97] wl[268] vdd gnd cell_6t
Xbit_r269_c97 bl[97] br[97] wl[269] vdd gnd cell_6t
Xbit_r270_c97 bl[97] br[97] wl[270] vdd gnd cell_6t
Xbit_r271_c97 bl[97] br[97] wl[271] vdd gnd cell_6t
Xbit_r272_c97 bl[97] br[97] wl[272] vdd gnd cell_6t
Xbit_r273_c97 bl[97] br[97] wl[273] vdd gnd cell_6t
Xbit_r274_c97 bl[97] br[97] wl[274] vdd gnd cell_6t
Xbit_r275_c97 bl[97] br[97] wl[275] vdd gnd cell_6t
Xbit_r276_c97 bl[97] br[97] wl[276] vdd gnd cell_6t
Xbit_r277_c97 bl[97] br[97] wl[277] vdd gnd cell_6t
Xbit_r278_c97 bl[97] br[97] wl[278] vdd gnd cell_6t
Xbit_r279_c97 bl[97] br[97] wl[279] vdd gnd cell_6t
Xbit_r280_c97 bl[97] br[97] wl[280] vdd gnd cell_6t
Xbit_r281_c97 bl[97] br[97] wl[281] vdd gnd cell_6t
Xbit_r282_c97 bl[97] br[97] wl[282] vdd gnd cell_6t
Xbit_r283_c97 bl[97] br[97] wl[283] vdd gnd cell_6t
Xbit_r284_c97 bl[97] br[97] wl[284] vdd gnd cell_6t
Xbit_r285_c97 bl[97] br[97] wl[285] vdd gnd cell_6t
Xbit_r286_c97 bl[97] br[97] wl[286] vdd gnd cell_6t
Xbit_r287_c97 bl[97] br[97] wl[287] vdd gnd cell_6t
Xbit_r288_c97 bl[97] br[97] wl[288] vdd gnd cell_6t
Xbit_r289_c97 bl[97] br[97] wl[289] vdd gnd cell_6t
Xbit_r290_c97 bl[97] br[97] wl[290] vdd gnd cell_6t
Xbit_r291_c97 bl[97] br[97] wl[291] vdd gnd cell_6t
Xbit_r292_c97 bl[97] br[97] wl[292] vdd gnd cell_6t
Xbit_r293_c97 bl[97] br[97] wl[293] vdd gnd cell_6t
Xbit_r294_c97 bl[97] br[97] wl[294] vdd gnd cell_6t
Xbit_r295_c97 bl[97] br[97] wl[295] vdd gnd cell_6t
Xbit_r296_c97 bl[97] br[97] wl[296] vdd gnd cell_6t
Xbit_r297_c97 bl[97] br[97] wl[297] vdd gnd cell_6t
Xbit_r298_c97 bl[97] br[97] wl[298] vdd gnd cell_6t
Xbit_r299_c97 bl[97] br[97] wl[299] vdd gnd cell_6t
Xbit_r300_c97 bl[97] br[97] wl[300] vdd gnd cell_6t
Xbit_r301_c97 bl[97] br[97] wl[301] vdd gnd cell_6t
Xbit_r302_c97 bl[97] br[97] wl[302] vdd gnd cell_6t
Xbit_r303_c97 bl[97] br[97] wl[303] vdd gnd cell_6t
Xbit_r304_c97 bl[97] br[97] wl[304] vdd gnd cell_6t
Xbit_r305_c97 bl[97] br[97] wl[305] vdd gnd cell_6t
Xbit_r306_c97 bl[97] br[97] wl[306] vdd gnd cell_6t
Xbit_r307_c97 bl[97] br[97] wl[307] vdd gnd cell_6t
Xbit_r308_c97 bl[97] br[97] wl[308] vdd gnd cell_6t
Xbit_r309_c97 bl[97] br[97] wl[309] vdd gnd cell_6t
Xbit_r310_c97 bl[97] br[97] wl[310] vdd gnd cell_6t
Xbit_r311_c97 bl[97] br[97] wl[311] vdd gnd cell_6t
Xbit_r312_c97 bl[97] br[97] wl[312] vdd gnd cell_6t
Xbit_r313_c97 bl[97] br[97] wl[313] vdd gnd cell_6t
Xbit_r314_c97 bl[97] br[97] wl[314] vdd gnd cell_6t
Xbit_r315_c97 bl[97] br[97] wl[315] vdd gnd cell_6t
Xbit_r316_c97 bl[97] br[97] wl[316] vdd gnd cell_6t
Xbit_r317_c97 bl[97] br[97] wl[317] vdd gnd cell_6t
Xbit_r318_c97 bl[97] br[97] wl[318] vdd gnd cell_6t
Xbit_r319_c97 bl[97] br[97] wl[319] vdd gnd cell_6t
Xbit_r320_c97 bl[97] br[97] wl[320] vdd gnd cell_6t
Xbit_r321_c97 bl[97] br[97] wl[321] vdd gnd cell_6t
Xbit_r322_c97 bl[97] br[97] wl[322] vdd gnd cell_6t
Xbit_r323_c97 bl[97] br[97] wl[323] vdd gnd cell_6t
Xbit_r324_c97 bl[97] br[97] wl[324] vdd gnd cell_6t
Xbit_r325_c97 bl[97] br[97] wl[325] vdd gnd cell_6t
Xbit_r326_c97 bl[97] br[97] wl[326] vdd gnd cell_6t
Xbit_r327_c97 bl[97] br[97] wl[327] vdd gnd cell_6t
Xbit_r328_c97 bl[97] br[97] wl[328] vdd gnd cell_6t
Xbit_r329_c97 bl[97] br[97] wl[329] vdd gnd cell_6t
Xbit_r330_c97 bl[97] br[97] wl[330] vdd gnd cell_6t
Xbit_r331_c97 bl[97] br[97] wl[331] vdd gnd cell_6t
Xbit_r332_c97 bl[97] br[97] wl[332] vdd gnd cell_6t
Xbit_r333_c97 bl[97] br[97] wl[333] vdd gnd cell_6t
Xbit_r334_c97 bl[97] br[97] wl[334] vdd gnd cell_6t
Xbit_r335_c97 bl[97] br[97] wl[335] vdd gnd cell_6t
Xbit_r336_c97 bl[97] br[97] wl[336] vdd gnd cell_6t
Xbit_r337_c97 bl[97] br[97] wl[337] vdd gnd cell_6t
Xbit_r338_c97 bl[97] br[97] wl[338] vdd gnd cell_6t
Xbit_r339_c97 bl[97] br[97] wl[339] vdd gnd cell_6t
Xbit_r340_c97 bl[97] br[97] wl[340] vdd gnd cell_6t
Xbit_r341_c97 bl[97] br[97] wl[341] vdd gnd cell_6t
Xbit_r342_c97 bl[97] br[97] wl[342] vdd gnd cell_6t
Xbit_r343_c97 bl[97] br[97] wl[343] vdd gnd cell_6t
Xbit_r344_c97 bl[97] br[97] wl[344] vdd gnd cell_6t
Xbit_r345_c97 bl[97] br[97] wl[345] vdd gnd cell_6t
Xbit_r346_c97 bl[97] br[97] wl[346] vdd gnd cell_6t
Xbit_r347_c97 bl[97] br[97] wl[347] vdd gnd cell_6t
Xbit_r348_c97 bl[97] br[97] wl[348] vdd gnd cell_6t
Xbit_r349_c97 bl[97] br[97] wl[349] vdd gnd cell_6t
Xbit_r350_c97 bl[97] br[97] wl[350] vdd gnd cell_6t
Xbit_r351_c97 bl[97] br[97] wl[351] vdd gnd cell_6t
Xbit_r352_c97 bl[97] br[97] wl[352] vdd gnd cell_6t
Xbit_r353_c97 bl[97] br[97] wl[353] vdd gnd cell_6t
Xbit_r354_c97 bl[97] br[97] wl[354] vdd gnd cell_6t
Xbit_r355_c97 bl[97] br[97] wl[355] vdd gnd cell_6t
Xbit_r356_c97 bl[97] br[97] wl[356] vdd gnd cell_6t
Xbit_r357_c97 bl[97] br[97] wl[357] vdd gnd cell_6t
Xbit_r358_c97 bl[97] br[97] wl[358] vdd gnd cell_6t
Xbit_r359_c97 bl[97] br[97] wl[359] vdd gnd cell_6t
Xbit_r360_c97 bl[97] br[97] wl[360] vdd gnd cell_6t
Xbit_r361_c97 bl[97] br[97] wl[361] vdd gnd cell_6t
Xbit_r362_c97 bl[97] br[97] wl[362] vdd gnd cell_6t
Xbit_r363_c97 bl[97] br[97] wl[363] vdd gnd cell_6t
Xbit_r364_c97 bl[97] br[97] wl[364] vdd gnd cell_6t
Xbit_r365_c97 bl[97] br[97] wl[365] vdd gnd cell_6t
Xbit_r366_c97 bl[97] br[97] wl[366] vdd gnd cell_6t
Xbit_r367_c97 bl[97] br[97] wl[367] vdd gnd cell_6t
Xbit_r368_c97 bl[97] br[97] wl[368] vdd gnd cell_6t
Xbit_r369_c97 bl[97] br[97] wl[369] vdd gnd cell_6t
Xbit_r370_c97 bl[97] br[97] wl[370] vdd gnd cell_6t
Xbit_r371_c97 bl[97] br[97] wl[371] vdd gnd cell_6t
Xbit_r372_c97 bl[97] br[97] wl[372] vdd gnd cell_6t
Xbit_r373_c97 bl[97] br[97] wl[373] vdd gnd cell_6t
Xbit_r374_c97 bl[97] br[97] wl[374] vdd gnd cell_6t
Xbit_r375_c97 bl[97] br[97] wl[375] vdd gnd cell_6t
Xbit_r376_c97 bl[97] br[97] wl[376] vdd gnd cell_6t
Xbit_r377_c97 bl[97] br[97] wl[377] vdd gnd cell_6t
Xbit_r378_c97 bl[97] br[97] wl[378] vdd gnd cell_6t
Xbit_r379_c97 bl[97] br[97] wl[379] vdd gnd cell_6t
Xbit_r380_c97 bl[97] br[97] wl[380] vdd gnd cell_6t
Xbit_r381_c97 bl[97] br[97] wl[381] vdd gnd cell_6t
Xbit_r382_c97 bl[97] br[97] wl[382] vdd gnd cell_6t
Xbit_r383_c97 bl[97] br[97] wl[383] vdd gnd cell_6t
Xbit_r384_c97 bl[97] br[97] wl[384] vdd gnd cell_6t
Xbit_r385_c97 bl[97] br[97] wl[385] vdd gnd cell_6t
Xbit_r386_c97 bl[97] br[97] wl[386] vdd gnd cell_6t
Xbit_r387_c97 bl[97] br[97] wl[387] vdd gnd cell_6t
Xbit_r388_c97 bl[97] br[97] wl[388] vdd gnd cell_6t
Xbit_r389_c97 bl[97] br[97] wl[389] vdd gnd cell_6t
Xbit_r390_c97 bl[97] br[97] wl[390] vdd gnd cell_6t
Xbit_r391_c97 bl[97] br[97] wl[391] vdd gnd cell_6t
Xbit_r392_c97 bl[97] br[97] wl[392] vdd gnd cell_6t
Xbit_r393_c97 bl[97] br[97] wl[393] vdd gnd cell_6t
Xbit_r394_c97 bl[97] br[97] wl[394] vdd gnd cell_6t
Xbit_r395_c97 bl[97] br[97] wl[395] vdd gnd cell_6t
Xbit_r396_c97 bl[97] br[97] wl[396] vdd gnd cell_6t
Xbit_r397_c97 bl[97] br[97] wl[397] vdd gnd cell_6t
Xbit_r398_c97 bl[97] br[97] wl[398] vdd gnd cell_6t
Xbit_r399_c97 bl[97] br[97] wl[399] vdd gnd cell_6t
Xbit_r400_c97 bl[97] br[97] wl[400] vdd gnd cell_6t
Xbit_r401_c97 bl[97] br[97] wl[401] vdd gnd cell_6t
Xbit_r402_c97 bl[97] br[97] wl[402] vdd gnd cell_6t
Xbit_r403_c97 bl[97] br[97] wl[403] vdd gnd cell_6t
Xbit_r404_c97 bl[97] br[97] wl[404] vdd gnd cell_6t
Xbit_r405_c97 bl[97] br[97] wl[405] vdd gnd cell_6t
Xbit_r406_c97 bl[97] br[97] wl[406] vdd gnd cell_6t
Xbit_r407_c97 bl[97] br[97] wl[407] vdd gnd cell_6t
Xbit_r408_c97 bl[97] br[97] wl[408] vdd gnd cell_6t
Xbit_r409_c97 bl[97] br[97] wl[409] vdd gnd cell_6t
Xbit_r410_c97 bl[97] br[97] wl[410] vdd gnd cell_6t
Xbit_r411_c97 bl[97] br[97] wl[411] vdd gnd cell_6t
Xbit_r412_c97 bl[97] br[97] wl[412] vdd gnd cell_6t
Xbit_r413_c97 bl[97] br[97] wl[413] vdd gnd cell_6t
Xbit_r414_c97 bl[97] br[97] wl[414] vdd gnd cell_6t
Xbit_r415_c97 bl[97] br[97] wl[415] vdd gnd cell_6t
Xbit_r416_c97 bl[97] br[97] wl[416] vdd gnd cell_6t
Xbit_r417_c97 bl[97] br[97] wl[417] vdd gnd cell_6t
Xbit_r418_c97 bl[97] br[97] wl[418] vdd gnd cell_6t
Xbit_r419_c97 bl[97] br[97] wl[419] vdd gnd cell_6t
Xbit_r420_c97 bl[97] br[97] wl[420] vdd gnd cell_6t
Xbit_r421_c97 bl[97] br[97] wl[421] vdd gnd cell_6t
Xbit_r422_c97 bl[97] br[97] wl[422] vdd gnd cell_6t
Xbit_r423_c97 bl[97] br[97] wl[423] vdd gnd cell_6t
Xbit_r424_c97 bl[97] br[97] wl[424] vdd gnd cell_6t
Xbit_r425_c97 bl[97] br[97] wl[425] vdd gnd cell_6t
Xbit_r426_c97 bl[97] br[97] wl[426] vdd gnd cell_6t
Xbit_r427_c97 bl[97] br[97] wl[427] vdd gnd cell_6t
Xbit_r428_c97 bl[97] br[97] wl[428] vdd gnd cell_6t
Xbit_r429_c97 bl[97] br[97] wl[429] vdd gnd cell_6t
Xbit_r430_c97 bl[97] br[97] wl[430] vdd gnd cell_6t
Xbit_r431_c97 bl[97] br[97] wl[431] vdd gnd cell_6t
Xbit_r432_c97 bl[97] br[97] wl[432] vdd gnd cell_6t
Xbit_r433_c97 bl[97] br[97] wl[433] vdd gnd cell_6t
Xbit_r434_c97 bl[97] br[97] wl[434] vdd gnd cell_6t
Xbit_r435_c97 bl[97] br[97] wl[435] vdd gnd cell_6t
Xbit_r436_c97 bl[97] br[97] wl[436] vdd gnd cell_6t
Xbit_r437_c97 bl[97] br[97] wl[437] vdd gnd cell_6t
Xbit_r438_c97 bl[97] br[97] wl[438] vdd gnd cell_6t
Xbit_r439_c97 bl[97] br[97] wl[439] vdd gnd cell_6t
Xbit_r440_c97 bl[97] br[97] wl[440] vdd gnd cell_6t
Xbit_r441_c97 bl[97] br[97] wl[441] vdd gnd cell_6t
Xbit_r442_c97 bl[97] br[97] wl[442] vdd gnd cell_6t
Xbit_r443_c97 bl[97] br[97] wl[443] vdd gnd cell_6t
Xbit_r444_c97 bl[97] br[97] wl[444] vdd gnd cell_6t
Xbit_r445_c97 bl[97] br[97] wl[445] vdd gnd cell_6t
Xbit_r446_c97 bl[97] br[97] wl[446] vdd gnd cell_6t
Xbit_r447_c97 bl[97] br[97] wl[447] vdd gnd cell_6t
Xbit_r448_c97 bl[97] br[97] wl[448] vdd gnd cell_6t
Xbit_r449_c97 bl[97] br[97] wl[449] vdd gnd cell_6t
Xbit_r450_c97 bl[97] br[97] wl[450] vdd gnd cell_6t
Xbit_r451_c97 bl[97] br[97] wl[451] vdd gnd cell_6t
Xbit_r452_c97 bl[97] br[97] wl[452] vdd gnd cell_6t
Xbit_r453_c97 bl[97] br[97] wl[453] vdd gnd cell_6t
Xbit_r454_c97 bl[97] br[97] wl[454] vdd gnd cell_6t
Xbit_r455_c97 bl[97] br[97] wl[455] vdd gnd cell_6t
Xbit_r456_c97 bl[97] br[97] wl[456] vdd gnd cell_6t
Xbit_r457_c97 bl[97] br[97] wl[457] vdd gnd cell_6t
Xbit_r458_c97 bl[97] br[97] wl[458] vdd gnd cell_6t
Xbit_r459_c97 bl[97] br[97] wl[459] vdd gnd cell_6t
Xbit_r460_c97 bl[97] br[97] wl[460] vdd gnd cell_6t
Xbit_r461_c97 bl[97] br[97] wl[461] vdd gnd cell_6t
Xbit_r462_c97 bl[97] br[97] wl[462] vdd gnd cell_6t
Xbit_r463_c97 bl[97] br[97] wl[463] vdd gnd cell_6t
Xbit_r464_c97 bl[97] br[97] wl[464] vdd gnd cell_6t
Xbit_r465_c97 bl[97] br[97] wl[465] vdd gnd cell_6t
Xbit_r466_c97 bl[97] br[97] wl[466] vdd gnd cell_6t
Xbit_r467_c97 bl[97] br[97] wl[467] vdd gnd cell_6t
Xbit_r468_c97 bl[97] br[97] wl[468] vdd gnd cell_6t
Xbit_r469_c97 bl[97] br[97] wl[469] vdd gnd cell_6t
Xbit_r470_c97 bl[97] br[97] wl[470] vdd gnd cell_6t
Xbit_r471_c97 bl[97] br[97] wl[471] vdd gnd cell_6t
Xbit_r472_c97 bl[97] br[97] wl[472] vdd gnd cell_6t
Xbit_r473_c97 bl[97] br[97] wl[473] vdd gnd cell_6t
Xbit_r474_c97 bl[97] br[97] wl[474] vdd gnd cell_6t
Xbit_r475_c97 bl[97] br[97] wl[475] vdd gnd cell_6t
Xbit_r476_c97 bl[97] br[97] wl[476] vdd gnd cell_6t
Xbit_r477_c97 bl[97] br[97] wl[477] vdd gnd cell_6t
Xbit_r478_c97 bl[97] br[97] wl[478] vdd gnd cell_6t
Xbit_r479_c97 bl[97] br[97] wl[479] vdd gnd cell_6t
Xbit_r480_c97 bl[97] br[97] wl[480] vdd gnd cell_6t
Xbit_r481_c97 bl[97] br[97] wl[481] vdd gnd cell_6t
Xbit_r482_c97 bl[97] br[97] wl[482] vdd gnd cell_6t
Xbit_r483_c97 bl[97] br[97] wl[483] vdd gnd cell_6t
Xbit_r484_c97 bl[97] br[97] wl[484] vdd gnd cell_6t
Xbit_r485_c97 bl[97] br[97] wl[485] vdd gnd cell_6t
Xbit_r486_c97 bl[97] br[97] wl[486] vdd gnd cell_6t
Xbit_r487_c97 bl[97] br[97] wl[487] vdd gnd cell_6t
Xbit_r488_c97 bl[97] br[97] wl[488] vdd gnd cell_6t
Xbit_r489_c97 bl[97] br[97] wl[489] vdd gnd cell_6t
Xbit_r490_c97 bl[97] br[97] wl[490] vdd gnd cell_6t
Xbit_r491_c97 bl[97] br[97] wl[491] vdd gnd cell_6t
Xbit_r492_c97 bl[97] br[97] wl[492] vdd gnd cell_6t
Xbit_r493_c97 bl[97] br[97] wl[493] vdd gnd cell_6t
Xbit_r494_c97 bl[97] br[97] wl[494] vdd gnd cell_6t
Xbit_r495_c97 bl[97] br[97] wl[495] vdd gnd cell_6t
Xbit_r496_c97 bl[97] br[97] wl[496] vdd gnd cell_6t
Xbit_r497_c97 bl[97] br[97] wl[497] vdd gnd cell_6t
Xbit_r498_c97 bl[97] br[97] wl[498] vdd gnd cell_6t
Xbit_r499_c97 bl[97] br[97] wl[499] vdd gnd cell_6t
Xbit_r500_c97 bl[97] br[97] wl[500] vdd gnd cell_6t
Xbit_r501_c97 bl[97] br[97] wl[501] vdd gnd cell_6t
Xbit_r502_c97 bl[97] br[97] wl[502] vdd gnd cell_6t
Xbit_r503_c97 bl[97] br[97] wl[503] vdd gnd cell_6t
Xbit_r504_c97 bl[97] br[97] wl[504] vdd gnd cell_6t
Xbit_r505_c97 bl[97] br[97] wl[505] vdd gnd cell_6t
Xbit_r506_c97 bl[97] br[97] wl[506] vdd gnd cell_6t
Xbit_r507_c97 bl[97] br[97] wl[507] vdd gnd cell_6t
Xbit_r508_c97 bl[97] br[97] wl[508] vdd gnd cell_6t
Xbit_r509_c97 bl[97] br[97] wl[509] vdd gnd cell_6t
Xbit_r510_c97 bl[97] br[97] wl[510] vdd gnd cell_6t
Xbit_r511_c97 bl[97] br[97] wl[511] vdd gnd cell_6t
Xbit_r0_c98 bl[98] br[98] wl[0] vdd gnd cell_6t
Xbit_r1_c98 bl[98] br[98] wl[1] vdd gnd cell_6t
Xbit_r2_c98 bl[98] br[98] wl[2] vdd gnd cell_6t
Xbit_r3_c98 bl[98] br[98] wl[3] vdd gnd cell_6t
Xbit_r4_c98 bl[98] br[98] wl[4] vdd gnd cell_6t
Xbit_r5_c98 bl[98] br[98] wl[5] vdd gnd cell_6t
Xbit_r6_c98 bl[98] br[98] wl[6] vdd gnd cell_6t
Xbit_r7_c98 bl[98] br[98] wl[7] vdd gnd cell_6t
Xbit_r8_c98 bl[98] br[98] wl[8] vdd gnd cell_6t
Xbit_r9_c98 bl[98] br[98] wl[9] vdd gnd cell_6t
Xbit_r10_c98 bl[98] br[98] wl[10] vdd gnd cell_6t
Xbit_r11_c98 bl[98] br[98] wl[11] vdd gnd cell_6t
Xbit_r12_c98 bl[98] br[98] wl[12] vdd gnd cell_6t
Xbit_r13_c98 bl[98] br[98] wl[13] vdd gnd cell_6t
Xbit_r14_c98 bl[98] br[98] wl[14] vdd gnd cell_6t
Xbit_r15_c98 bl[98] br[98] wl[15] vdd gnd cell_6t
Xbit_r16_c98 bl[98] br[98] wl[16] vdd gnd cell_6t
Xbit_r17_c98 bl[98] br[98] wl[17] vdd gnd cell_6t
Xbit_r18_c98 bl[98] br[98] wl[18] vdd gnd cell_6t
Xbit_r19_c98 bl[98] br[98] wl[19] vdd gnd cell_6t
Xbit_r20_c98 bl[98] br[98] wl[20] vdd gnd cell_6t
Xbit_r21_c98 bl[98] br[98] wl[21] vdd gnd cell_6t
Xbit_r22_c98 bl[98] br[98] wl[22] vdd gnd cell_6t
Xbit_r23_c98 bl[98] br[98] wl[23] vdd gnd cell_6t
Xbit_r24_c98 bl[98] br[98] wl[24] vdd gnd cell_6t
Xbit_r25_c98 bl[98] br[98] wl[25] vdd gnd cell_6t
Xbit_r26_c98 bl[98] br[98] wl[26] vdd gnd cell_6t
Xbit_r27_c98 bl[98] br[98] wl[27] vdd gnd cell_6t
Xbit_r28_c98 bl[98] br[98] wl[28] vdd gnd cell_6t
Xbit_r29_c98 bl[98] br[98] wl[29] vdd gnd cell_6t
Xbit_r30_c98 bl[98] br[98] wl[30] vdd gnd cell_6t
Xbit_r31_c98 bl[98] br[98] wl[31] vdd gnd cell_6t
Xbit_r32_c98 bl[98] br[98] wl[32] vdd gnd cell_6t
Xbit_r33_c98 bl[98] br[98] wl[33] vdd gnd cell_6t
Xbit_r34_c98 bl[98] br[98] wl[34] vdd gnd cell_6t
Xbit_r35_c98 bl[98] br[98] wl[35] vdd gnd cell_6t
Xbit_r36_c98 bl[98] br[98] wl[36] vdd gnd cell_6t
Xbit_r37_c98 bl[98] br[98] wl[37] vdd gnd cell_6t
Xbit_r38_c98 bl[98] br[98] wl[38] vdd gnd cell_6t
Xbit_r39_c98 bl[98] br[98] wl[39] vdd gnd cell_6t
Xbit_r40_c98 bl[98] br[98] wl[40] vdd gnd cell_6t
Xbit_r41_c98 bl[98] br[98] wl[41] vdd gnd cell_6t
Xbit_r42_c98 bl[98] br[98] wl[42] vdd gnd cell_6t
Xbit_r43_c98 bl[98] br[98] wl[43] vdd gnd cell_6t
Xbit_r44_c98 bl[98] br[98] wl[44] vdd gnd cell_6t
Xbit_r45_c98 bl[98] br[98] wl[45] vdd gnd cell_6t
Xbit_r46_c98 bl[98] br[98] wl[46] vdd gnd cell_6t
Xbit_r47_c98 bl[98] br[98] wl[47] vdd gnd cell_6t
Xbit_r48_c98 bl[98] br[98] wl[48] vdd gnd cell_6t
Xbit_r49_c98 bl[98] br[98] wl[49] vdd gnd cell_6t
Xbit_r50_c98 bl[98] br[98] wl[50] vdd gnd cell_6t
Xbit_r51_c98 bl[98] br[98] wl[51] vdd gnd cell_6t
Xbit_r52_c98 bl[98] br[98] wl[52] vdd gnd cell_6t
Xbit_r53_c98 bl[98] br[98] wl[53] vdd gnd cell_6t
Xbit_r54_c98 bl[98] br[98] wl[54] vdd gnd cell_6t
Xbit_r55_c98 bl[98] br[98] wl[55] vdd gnd cell_6t
Xbit_r56_c98 bl[98] br[98] wl[56] vdd gnd cell_6t
Xbit_r57_c98 bl[98] br[98] wl[57] vdd gnd cell_6t
Xbit_r58_c98 bl[98] br[98] wl[58] vdd gnd cell_6t
Xbit_r59_c98 bl[98] br[98] wl[59] vdd gnd cell_6t
Xbit_r60_c98 bl[98] br[98] wl[60] vdd gnd cell_6t
Xbit_r61_c98 bl[98] br[98] wl[61] vdd gnd cell_6t
Xbit_r62_c98 bl[98] br[98] wl[62] vdd gnd cell_6t
Xbit_r63_c98 bl[98] br[98] wl[63] vdd gnd cell_6t
Xbit_r64_c98 bl[98] br[98] wl[64] vdd gnd cell_6t
Xbit_r65_c98 bl[98] br[98] wl[65] vdd gnd cell_6t
Xbit_r66_c98 bl[98] br[98] wl[66] vdd gnd cell_6t
Xbit_r67_c98 bl[98] br[98] wl[67] vdd gnd cell_6t
Xbit_r68_c98 bl[98] br[98] wl[68] vdd gnd cell_6t
Xbit_r69_c98 bl[98] br[98] wl[69] vdd gnd cell_6t
Xbit_r70_c98 bl[98] br[98] wl[70] vdd gnd cell_6t
Xbit_r71_c98 bl[98] br[98] wl[71] vdd gnd cell_6t
Xbit_r72_c98 bl[98] br[98] wl[72] vdd gnd cell_6t
Xbit_r73_c98 bl[98] br[98] wl[73] vdd gnd cell_6t
Xbit_r74_c98 bl[98] br[98] wl[74] vdd gnd cell_6t
Xbit_r75_c98 bl[98] br[98] wl[75] vdd gnd cell_6t
Xbit_r76_c98 bl[98] br[98] wl[76] vdd gnd cell_6t
Xbit_r77_c98 bl[98] br[98] wl[77] vdd gnd cell_6t
Xbit_r78_c98 bl[98] br[98] wl[78] vdd gnd cell_6t
Xbit_r79_c98 bl[98] br[98] wl[79] vdd gnd cell_6t
Xbit_r80_c98 bl[98] br[98] wl[80] vdd gnd cell_6t
Xbit_r81_c98 bl[98] br[98] wl[81] vdd gnd cell_6t
Xbit_r82_c98 bl[98] br[98] wl[82] vdd gnd cell_6t
Xbit_r83_c98 bl[98] br[98] wl[83] vdd gnd cell_6t
Xbit_r84_c98 bl[98] br[98] wl[84] vdd gnd cell_6t
Xbit_r85_c98 bl[98] br[98] wl[85] vdd gnd cell_6t
Xbit_r86_c98 bl[98] br[98] wl[86] vdd gnd cell_6t
Xbit_r87_c98 bl[98] br[98] wl[87] vdd gnd cell_6t
Xbit_r88_c98 bl[98] br[98] wl[88] vdd gnd cell_6t
Xbit_r89_c98 bl[98] br[98] wl[89] vdd gnd cell_6t
Xbit_r90_c98 bl[98] br[98] wl[90] vdd gnd cell_6t
Xbit_r91_c98 bl[98] br[98] wl[91] vdd gnd cell_6t
Xbit_r92_c98 bl[98] br[98] wl[92] vdd gnd cell_6t
Xbit_r93_c98 bl[98] br[98] wl[93] vdd gnd cell_6t
Xbit_r94_c98 bl[98] br[98] wl[94] vdd gnd cell_6t
Xbit_r95_c98 bl[98] br[98] wl[95] vdd gnd cell_6t
Xbit_r96_c98 bl[98] br[98] wl[96] vdd gnd cell_6t
Xbit_r97_c98 bl[98] br[98] wl[97] vdd gnd cell_6t
Xbit_r98_c98 bl[98] br[98] wl[98] vdd gnd cell_6t
Xbit_r99_c98 bl[98] br[98] wl[99] vdd gnd cell_6t
Xbit_r100_c98 bl[98] br[98] wl[100] vdd gnd cell_6t
Xbit_r101_c98 bl[98] br[98] wl[101] vdd gnd cell_6t
Xbit_r102_c98 bl[98] br[98] wl[102] vdd gnd cell_6t
Xbit_r103_c98 bl[98] br[98] wl[103] vdd gnd cell_6t
Xbit_r104_c98 bl[98] br[98] wl[104] vdd gnd cell_6t
Xbit_r105_c98 bl[98] br[98] wl[105] vdd gnd cell_6t
Xbit_r106_c98 bl[98] br[98] wl[106] vdd gnd cell_6t
Xbit_r107_c98 bl[98] br[98] wl[107] vdd gnd cell_6t
Xbit_r108_c98 bl[98] br[98] wl[108] vdd gnd cell_6t
Xbit_r109_c98 bl[98] br[98] wl[109] vdd gnd cell_6t
Xbit_r110_c98 bl[98] br[98] wl[110] vdd gnd cell_6t
Xbit_r111_c98 bl[98] br[98] wl[111] vdd gnd cell_6t
Xbit_r112_c98 bl[98] br[98] wl[112] vdd gnd cell_6t
Xbit_r113_c98 bl[98] br[98] wl[113] vdd gnd cell_6t
Xbit_r114_c98 bl[98] br[98] wl[114] vdd gnd cell_6t
Xbit_r115_c98 bl[98] br[98] wl[115] vdd gnd cell_6t
Xbit_r116_c98 bl[98] br[98] wl[116] vdd gnd cell_6t
Xbit_r117_c98 bl[98] br[98] wl[117] vdd gnd cell_6t
Xbit_r118_c98 bl[98] br[98] wl[118] vdd gnd cell_6t
Xbit_r119_c98 bl[98] br[98] wl[119] vdd gnd cell_6t
Xbit_r120_c98 bl[98] br[98] wl[120] vdd gnd cell_6t
Xbit_r121_c98 bl[98] br[98] wl[121] vdd gnd cell_6t
Xbit_r122_c98 bl[98] br[98] wl[122] vdd gnd cell_6t
Xbit_r123_c98 bl[98] br[98] wl[123] vdd gnd cell_6t
Xbit_r124_c98 bl[98] br[98] wl[124] vdd gnd cell_6t
Xbit_r125_c98 bl[98] br[98] wl[125] vdd gnd cell_6t
Xbit_r126_c98 bl[98] br[98] wl[126] vdd gnd cell_6t
Xbit_r127_c98 bl[98] br[98] wl[127] vdd gnd cell_6t
Xbit_r128_c98 bl[98] br[98] wl[128] vdd gnd cell_6t
Xbit_r129_c98 bl[98] br[98] wl[129] vdd gnd cell_6t
Xbit_r130_c98 bl[98] br[98] wl[130] vdd gnd cell_6t
Xbit_r131_c98 bl[98] br[98] wl[131] vdd gnd cell_6t
Xbit_r132_c98 bl[98] br[98] wl[132] vdd gnd cell_6t
Xbit_r133_c98 bl[98] br[98] wl[133] vdd gnd cell_6t
Xbit_r134_c98 bl[98] br[98] wl[134] vdd gnd cell_6t
Xbit_r135_c98 bl[98] br[98] wl[135] vdd gnd cell_6t
Xbit_r136_c98 bl[98] br[98] wl[136] vdd gnd cell_6t
Xbit_r137_c98 bl[98] br[98] wl[137] vdd gnd cell_6t
Xbit_r138_c98 bl[98] br[98] wl[138] vdd gnd cell_6t
Xbit_r139_c98 bl[98] br[98] wl[139] vdd gnd cell_6t
Xbit_r140_c98 bl[98] br[98] wl[140] vdd gnd cell_6t
Xbit_r141_c98 bl[98] br[98] wl[141] vdd gnd cell_6t
Xbit_r142_c98 bl[98] br[98] wl[142] vdd gnd cell_6t
Xbit_r143_c98 bl[98] br[98] wl[143] vdd gnd cell_6t
Xbit_r144_c98 bl[98] br[98] wl[144] vdd gnd cell_6t
Xbit_r145_c98 bl[98] br[98] wl[145] vdd gnd cell_6t
Xbit_r146_c98 bl[98] br[98] wl[146] vdd gnd cell_6t
Xbit_r147_c98 bl[98] br[98] wl[147] vdd gnd cell_6t
Xbit_r148_c98 bl[98] br[98] wl[148] vdd gnd cell_6t
Xbit_r149_c98 bl[98] br[98] wl[149] vdd gnd cell_6t
Xbit_r150_c98 bl[98] br[98] wl[150] vdd gnd cell_6t
Xbit_r151_c98 bl[98] br[98] wl[151] vdd gnd cell_6t
Xbit_r152_c98 bl[98] br[98] wl[152] vdd gnd cell_6t
Xbit_r153_c98 bl[98] br[98] wl[153] vdd gnd cell_6t
Xbit_r154_c98 bl[98] br[98] wl[154] vdd gnd cell_6t
Xbit_r155_c98 bl[98] br[98] wl[155] vdd gnd cell_6t
Xbit_r156_c98 bl[98] br[98] wl[156] vdd gnd cell_6t
Xbit_r157_c98 bl[98] br[98] wl[157] vdd gnd cell_6t
Xbit_r158_c98 bl[98] br[98] wl[158] vdd gnd cell_6t
Xbit_r159_c98 bl[98] br[98] wl[159] vdd gnd cell_6t
Xbit_r160_c98 bl[98] br[98] wl[160] vdd gnd cell_6t
Xbit_r161_c98 bl[98] br[98] wl[161] vdd gnd cell_6t
Xbit_r162_c98 bl[98] br[98] wl[162] vdd gnd cell_6t
Xbit_r163_c98 bl[98] br[98] wl[163] vdd gnd cell_6t
Xbit_r164_c98 bl[98] br[98] wl[164] vdd gnd cell_6t
Xbit_r165_c98 bl[98] br[98] wl[165] vdd gnd cell_6t
Xbit_r166_c98 bl[98] br[98] wl[166] vdd gnd cell_6t
Xbit_r167_c98 bl[98] br[98] wl[167] vdd gnd cell_6t
Xbit_r168_c98 bl[98] br[98] wl[168] vdd gnd cell_6t
Xbit_r169_c98 bl[98] br[98] wl[169] vdd gnd cell_6t
Xbit_r170_c98 bl[98] br[98] wl[170] vdd gnd cell_6t
Xbit_r171_c98 bl[98] br[98] wl[171] vdd gnd cell_6t
Xbit_r172_c98 bl[98] br[98] wl[172] vdd gnd cell_6t
Xbit_r173_c98 bl[98] br[98] wl[173] vdd gnd cell_6t
Xbit_r174_c98 bl[98] br[98] wl[174] vdd gnd cell_6t
Xbit_r175_c98 bl[98] br[98] wl[175] vdd gnd cell_6t
Xbit_r176_c98 bl[98] br[98] wl[176] vdd gnd cell_6t
Xbit_r177_c98 bl[98] br[98] wl[177] vdd gnd cell_6t
Xbit_r178_c98 bl[98] br[98] wl[178] vdd gnd cell_6t
Xbit_r179_c98 bl[98] br[98] wl[179] vdd gnd cell_6t
Xbit_r180_c98 bl[98] br[98] wl[180] vdd gnd cell_6t
Xbit_r181_c98 bl[98] br[98] wl[181] vdd gnd cell_6t
Xbit_r182_c98 bl[98] br[98] wl[182] vdd gnd cell_6t
Xbit_r183_c98 bl[98] br[98] wl[183] vdd gnd cell_6t
Xbit_r184_c98 bl[98] br[98] wl[184] vdd gnd cell_6t
Xbit_r185_c98 bl[98] br[98] wl[185] vdd gnd cell_6t
Xbit_r186_c98 bl[98] br[98] wl[186] vdd gnd cell_6t
Xbit_r187_c98 bl[98] br[98] wl[187] vdd gnd cell_6t
Xbit_r188_c98 bl[98] br[98] wl[188] vdd gnd cell_6t
Xbit_r189_c98 bl[98] br[98] wl[189] vdd gnd cell_6t
Xbit_r190_c98 bl[98] br[98] wl[190] vdd gnd cell_6t
Xbit_r191_c98 bl[98] br[98] wl[191] vdd gnd cell_6t
Xbit_r192_c98 bl[98] br[98] wl[192] vdd gnd cell_6t
Xbit_r193_c98 bl[98] br[98] wl[193] vdd gnd cell_6t
Xbit_r194_c98 bl[98] br[98] wl[194] vdd gnd cell_6t
Xbit_r195_c98 bl[98] br[98] wl[195] vdd gnd cell_6t
Xbit_r196_c98 bl[98] br[98] wl[196] vdd gnd cell_6t
Xbit_r197_c98 bl[98] br[98] wl[197] vdd gnd cell_6t
Xbit_r198_c98 bl[98] br[98] wl[198] vdd gnd cell_6t
Xbit_r199_c98 bl[98] br[98] wl[199] vdd gnd cell_6t
Xbit_r200_c98 bl[98] br[98] wl[200] vdd gnd cell_6t
Xbit_r201_c98 bl[98] br[98] wl[201] vdd gnd cell_6t
Xbit_r202_c98 bl[98] br[98] wl[202] vdd gnd cell_6t
Xbit_r203_c98 bl[98] br[98] wl[203] vdd gnd cell_6t
Xbit_r204_c98 bl[98] br[98] wl[204] vdd gnd cell_6t
Xbit_r205_c98 bl[98] br[98] wl[205] vdd gnd cell_6t
Xbit_r206_c98 bl[98] br[98] wl[206] vdd gnd cell_6t
Xbit_r207_c98 bl[98] br[98] wl[207] vdd gnd cell_6t
Xbit_r208_c98 bl[98] br[98] wl[208] vdd gnd cell_6t
Xbit_r209_c98 bl[98] br[98] wl[209] vdd gnd cell_6t
Xbit_r210_c98 bl[98] br[98] wl[210] vdd gnd cell_6t
Xbit_r211_c98 bl[98] br[98] wl[211] vdd gnd cell_6t
Xbit_r212_c98 bl[98] br[98] wl[212] vdd gnd cell_6t
Xbit_r213_c98 bl[98] br[98] wl[213] vdd gnd cell_6t
Xbit_r214_c98 bl[98] br[98] wl[214] vdd gnd cell_6t
Xbit_r215_c98 bl[98] br[98] wl[215] vdd gnd cell_6t
Xbit_r216_c98 bl[98] br[98] wl[216] vdd gnd cell_6t
Xbit_r217_c98 bl[98] br[98] wl[217] vdd gnd cell_6t
Xbit_r218_c98 bl[98] br[98] wl[218] vdd gnd cell_6t
Xbit_r219_c98 bl[98] br[98] wl[219] vdd gnd cell_6t
Xbit_r220_c98 bl[98] br[98] wl[220] vdd gnd cell_6t
Xbit_r221_c98 bl[98] br[98] wl[221] vdd gnd cell_6t
Xbit_r222_c98 bl[98] br[98] wl[222] vdd gnd cell_6t
Xbit_r223_c98 bl[98] br[98] wl[223] vdd gnd cell_6t
Xbit_r224_c98 bl[98] br[98] wl[224] vdd gnd cell_6t
Xbit_r225_c98 bl[98] br[98] wl[225] vdd gnd cell_6t
Xbit_r226_c98 bl[98] br[98] wl[226] vdd gnd cell_6t
Xbit_r227_c98 bl[98] br[98] wl[227] vdd gnd cell_6t
Xbit_r228_c98 bl[98] br[98] wl[228] vdd gnd cell_6t
Xbit_r229_c98 bl[98] br[98] wl[229] vdd gnd cell_6t
Xbit_r230_c98 bl[98] br[98] wl[230] vdd gnd cell_6t
Xbit_r231_c98 bl[98] br[98] wl[231] vdd gnd cell_6t
Xbit_r232_c98 bl[98] br[98] wl[232] vdd gnd cell_6t
Xbit_r233_c98 bl[98] br[98] wl[233] vdd gnd cell_6t
Xbit_r234_c98 bl[98] br[98] wl[234] vdd gnd cell_6t
Xbit_r235_c98 bl[98] br[98] wl[235] vdd gnd cell_6t
Xbit_r236_c98 bl[98] br[98] wl[236] vdd gnd cell_6t
Xbit_r237_c98 bl[98] br[98] wl[237] vdd gnd cell_6t
Xbit_r238_c98 bl[98] br[98] wl[238] vdd gnd cell_6t
Xbit_r239_c98 bl[98] br[98] wl[239] vdd gnd cell_6t
Xbit_r240_c98 bl[98] br[98] wl[240] vdd gnd cell_6t
Xbit_r241_c98 bl[98] br[98] wl[241] vdd gnd cell_6t
Xbit_r242_c98 bl[98] br[98] wl[242] vdd gnd cell_6t
Xbit_r243_c98 bl[98] br[98] wl[243] vdd gnd cell_6t
Xbit_r244_c98 bl[98] br[98] wl[244] vdd gnd cell_6t
Xbit_r245_c98 bl[98] br[98] wl[245] vdd gnd cell_6t
Xbit_r246_c98 bl[98] br[98] wl[246] vdd gnd cell_6t
Xbit_r247_c98 bl[98] br[98] wl[247] vdd gnd cell_6t
Xbit_r248_c98 bl[98] br[98] wl[248] vdd gnd cell_6t
Xbit_r249_c98 bl[98] br[98] wl[249] vdd gnd cell_6t
Xbit_r250_c98 bl[98] br[98] wl[250] vdd gnd cell_6t
Xbit_r251_c98 bl[98] br[98] wl[251] vdd gnd cell_6t
Xbit_r252_c98 bl[98] br[98] wl[252] vdd gnd cell_6t
Xbit_r253_c98 bl[98] br[98] wl[253] vdd gnd cell_6t
Xbit_r254_c98 bl[98] br[98] wl[254] vdd gnd cell_6t
Xbit_r255_c98 bl[98] br[98] wl[255] vdd gnd cell_6t
Xbit_r256_c98 bl[98] br[98] wl[256] vdd gnd cell_6t
Xbit_r257_c98 bl[98] br[98] wl[257] vdd gnd cell_6t
Xbit_r258_c98 bl[98] br[98] wl[258] vdd gnd cell_6t
Xbit_r259_c98 bl[98] br[98] wl[259] vdd gnd cell_6t
Xbit_r260_c98 bl[98] br[98] wl[260] vdd gnd cell_6t
Xbit_r261_c98 bl[98] br[98] wl[261] vdd gnd cell_6t
Xbit_r262_c98 bl[98] br[98] wl[262] vdd gnd cell_6t
Xbit_r263_c98 bl[98] br[98] wl[263] vdd gnd cell_6t
Xbit_r264_c98 bl[98] br[98] wl[264] vdd gnd cell_6t
Xbit_r265_c98 bl[98] br[98] wl[265] vdd gnd cell_6t
Xbit_r266_c98 bl[98] br[98] wl[266] vdd gnd cell_6t
Xbit_r267_c98 bl[98] br[98] wl[267] vdd gnd cell_6t
Xbit_r268_c98 bl[98] br[98] wl[268] vdd gnd cell_6t
Xbit_r269_c98 bl[98] br[98] wl[269] vdd gnd cell_6t
Xbit_r270_c98 bl[98] br[98] wl[270] vdd gnd cell_6t
Xbit_r271_c98 bl[98] br[98] wl[271] vdd gnd cell_6t
Xbit_r272_c98 bl[98] br[98] wl[272] vdd gnd cell_6t
Xbit_r273_c98 bl[98] br[98] wl[273] vdd gnd cell_6t
Xbit_r274_c98 bl[98] br[98] wl[274] vdd gnd cell_6t
Xbit_r275_c98 bl[98] br[98] wl[275] vdd gnd cell_6t
Xbit_r276_c98 bl[98] br[98] wl[276] vdd gnd cell_6t
Xbit_r277_c98 bl[98] br[98] wl[277] vdd gnd cell_6t
Xbit_r278_c98 bl[98] br[98] wl[278] vdd gnd cell_6t
Xbit_r279_c98 bl[98] br[98] wl[279] vdd gnd cell_6t
Xbit_r280_c98 bl[98] br[98] wl[280] vdd gnd cell_6t
Xbit_r281_c98 bl[98] br[98] wl[281] vdd gnd cell_6t
Xbit_r282_c98 bl[98] br[98] wl[282] vdd gnd cell_6t
Xbit_r283_c98 bl[98] br[98] wl[283] vdd gnd cell_6t
Xbit_r284_c98 bl[98] br[98] wl[284] vdd gnd cell_6t
Xbit_r285_c98 bl[98] br[98] wl[285] vdd gnd cell_6t
Xbit_r286_c98 bl[98] br[98] wl[286] vdd gnd cell_6t
Xbit_r287_c98 bl[98] br[98] wl[287] vdd gnd cell_6t
Xbit_r288_c98 bl[98] br[98] wl[288] vdd gnd cell_6t
Xbit_r289_c98 bl[98] br[98] wl[289] vdd gnd cell_6t
Xbit_r290_c98 bl[98] br[98] wl[290] vdd gnd cell_6t
Xbit_r291_c98 bl[98] br[98] wl[291] vdd gnd cell_6t
Xbit_r292_c98 bl[98] br[98] wl[292] vdd gnd cell_6t
Xbit_r293_c98 bl[98] br[98] wl[293] vdd gnd cell_6t
Xbit_r294_c98 bl[98] br[98] wl[294] vdd gnd cell_6t
Xbit_r295_c98 bl[98] br[98] wl[295] vdd gnd cell_6t
Xbit_r296_c98 bl[98] br[98] wl[296] vdd gnd cell_6t
Xbit_r297_c98 bl[98] br[98] wl[297] vdd gnd cell_6t
Xbit_r298_c98 bl[98] br[98] wl[298] vdd gnd cell_6t
Xbit_r299_c98 bl[98] br[98] wl[299] vdd gnd cell_6t
Xbit_r300_c98 bl[98] br[98] wl[300] vdd gnd cell_6t
Xbit_r301_c98 bl[98] br[98] wl[301] vdd gnd cell_6t
Xbit_r302_c98 bl[98] br[98] wl[302] vdd gnd cell_6t
Xbit_r303_c98 bl[98] br[98] wl[303] vdd gnd cell_6t
Xbit_r304_c98 bl[98] br[98] wl[304] vdd gnd cell_6t
Xbit_r305_c98 bl[98] br[98] wl[305] vdd gnd cell_6t
Xbit_r306_c98 bl[98] br[98] wl[306] vdd gnd cell_6t
Xbit_r307_c98 bl[98] br[98] wl[307] vdd gnd cell_6t
Xbit_r308_c98 bl[98] br[98] wl[308] vdd gnd cell_6t
Xbit_r309_c98 bl[98] br[98] wl[309] vdd gnd cell_6t
Xbit_r310_c98 bl[98] br[98] wl[310] vdd gnd cell_6t
Xbit_r311_c98 bl[98] br[98] wl[311] vdd gnd cell_6t
Xbit_r312_c98 bl[98] br[98] wl[312] vdd gnd cell_6t
Xbit_r313_c98 bl[98] br[98] wl[313] vdd gnd cell_6t
Xbit_r314_c98 bl[98] br[98] wl[314] vdd gnd cell_6t
Xbit_r315_c98 bl[98] br[98] wl[315] vdd gnd cell_6t
Xbit_r316_c98 bl[98] br[98] wl[316] vdd gnd cell_6t
Xbit_r317_c98 bl[98] br[98] wl[317] vdd gnd cell_6t
Xbit_r318_c98 bl[98] br[98] wl[318] vdd gnd cell_6t
Xbit_r319_c98 bl[98] br[98] wl[319] vdd gnd cell_6t
Xbit_r320_c98 bl[98] br[98] wl[320] vdd gnd cell_6t
Xbit_r321_c98 bl[98] br[98] wl[321] vdd gnd cell_6t
Xbit_r322_c98 bl[98] br[98] wl[322] vdd gnd cell_6t
Xbit_r323_c98 bl[98] br[98] wl[323] vdd gnd cell_6t
Xbit_r324_c98 bl[98] br[98] wl[324] vdd gnd cell_6t
Xbit_r325_c98 bl[98] br[98] wl[325] vdd gnd cell_6t
Xbit_r326_c98 bl[98] br[98] wl[326] vdd gnd cell_6t
Xbit_r327_c98 bl[98] br[98] wl[327] vdd gnd cell_6t
Xbit_r328_c98 bl[98] br[98] wl[328] vdd gnd cell_6t
Xbit_r329_c98 bl[98] br[98] wl[329] vdd gnd cell_6t
Xbit_r330_c98 bl[98] br[98] wl[330] vdd gnd cell_6t
Xbit_r331_c98 bl[98] br[98] wl[331] vdd gnd cell_6t
Xbit_r332_c98 bl[98] br[98] wl[332] vdd gnd cell_6t
Xbit_r333_c98 bl[98] br[98] wl[333] vdd gnd cell_6t
Xbit_r334_c98 bl[98] br[98] wl[334] vdd gnd cell_6t
Xbit_r335_c98 bl[98] br[98] wl[335] vdd gnd cell_6t
Xbit_r336_c98 bl[98] br[98] wl[336] vdd gnd cell_6t
Xbit_r337_c98 bl[98] br[98] wl[337] vdd gnd cell_6t
Xbit_r338_c98 bl[98] br[98] wl[338] vdd gnd cell_6t
Xbit_r339_c98 bl[98] br[98] wl[339] vdd gnd cell_6t
Xbit_r340_c98 bl[98] br[98] wl[340] vdd gnd cell_6t
Xbit_r341_c98 bl[98] br[98] wl[341] vdd gnd cell_6t
Xbit_r342_c98 bl[98] br[98] wl[342] vdd gnd cell_6t
Xbit_r343_c98 bl[98] br[98] wl[343] vdd gnd cell_6t
Xbit_r344_c98 bl[98] br[98] wl[344] vdd gnd cell_6t
Xbit_r345_c98 bl[98] br[98] wl[345] vdd gnd cell_6t
Xbit_r346_c98 bl[98] br[98] wl[346] vdd gnd cell_6t
Xbit_r347_c98 bl[98] br[98] wl[347] vdd gnd cell_6t
Xbit_r348_c98 bl[98] br[98] wl[348] vdd gnd cell_6t
Xbit_r349_c98 bl[98] br[98] wl[349] vdd gnd cell_6t
Xbit_r350_c98 bl[98] br[98] wl[350] vdd gnd cell_6t
Xbit_r351_c98 bl[98] br[98] wl[351] vdd gnd cell_6t
Xbit_r352_c98 bl[98] br[98] wl[352] vdd gnd cell_6t
Xbit_r353_c98 bl[98] br[98] wl[353] vdd gnd cell_6t
Xbit_r354_c98 bl[98] br[98] wl[354] vdd gnd cell_6t
Xbit_r355_c98 bl[98] br[98] wl[355] vdd gnd cell_6t
Xbit_r356_c98 bl[98] br[98] wl[356] vdd gnd cell_6t
Xbit_r357_c98 bl[98] br[98] wl[357] vdd gnd cell_6t
Xbit_r358_c98 bl[98] br[98] wl[358] vdd gnd cell_6t
Xbit_r359_c98 bl[98] br[98] wl[359] vdd gnd cell_6t
Xbit_r360_c98 bl[98] br[98] wl[360] vdd gnd cell_6t
Xbit_r361_c98 bl[98] br[98] wl[361] vdd gnd cell_6t
Xbit_r362_c98 bl[98] br[98] wl[362] vdd gnd cell_6t
Xbit_r363_c98 bl[98] br[98] wl[363] vdd gnd cell_6t
Xbit_r364_c98 bl[98] br[98] wl[364] vdd gnd cell_6t
Xbit_r365_c98 bl[98] br[98] wl[365] vdd gnd cell_6t
Xbit_r366_c98 bl[98] br[98] wl[366] vdd gnd cell_6t
Xbit_r367_c98 bl[98] br[98] wl[367] vdd gnd cell_6t
Xbit_r368_c98 bl[98] br[98] wl[368] vdd gnd cell_6t
Xbit_r369_c98 bl[98] br[98] wl[369] vdd gnd cell_6t
Xbit_r370_c98 bl[98] br[98] wl[370] vdd gnd cell_6t
Xbit_r371_c98 bl[98] br[98] wl[371] vdd gnd cell_6t
Xbit_r372_c98 bl[98] br[98] wl[372] vdd gnd cell_6t
Xbit_r373_c98 bl[98] br[98] wl[373] vdd gnd cell_6t
Xbit_r374_c98 bl[98] br[98] wl[374] vdd gnd cell_6t
Xbit_r375_c98 bl[98] br[98] wl[375] vdd gnd cell_6t
Xbit_r376_c98 bl[98] br[98] wl[376] vdd gnd cell_6t
Xbit_r377_c98 bl[98] br[98] wl[377] vdd gnd cell_6t
Xbit_r378_c98 bl[98] br[98] wl[378] vdd gnd cell_6t
Xbit_r379_c98 bl[98] br[98] wl[379] vdd gnd cell_6t
Xbit_r380_c98 bl[98] br[98] wl[380] vdd gnd cell_6t
Xbit_r381_c98 bl[98] br[98] wl[381] vdd gnd cell_6t
Xbit_r382_c98 bl[98] br[98] wl[382] vdd gnd cell_6t
Xbit_r383_c98 bl[98] br[98] wl[383] vdd gnd cell_6t
Xbit_r384_c98 bl[98] br[98] wl[384] vdd gnd cell_6t
Xbit_r385_c98 bl[98] br[98] wl[385] vdd gnd cell_6t
Xbit_r386_c98 bl[98] br[98] wl[386] vdd gnd cell_6t
Xbit_r387_c98 bl[98] br[98] wl[387] vdd gnd cell_6t
Xbit_r388_c98 bl[98] br[98] wl[388] vdd gnd cell_6t
Xbit_r389_c98 bl[98] br[98] wl[389] vdd gnd cell_6t
Xbit_r390_c98 bl[98] br[98] wl[390] vdd gnd cell_6t
Xbit_r391_c98 bl[98] br[98] wl[391] vdd gnd cell_6t
Xbit_r392_c98 bl[98] br[98] wl[392] vdd gnd cell_6t
Xbit_r393_c98 bl[98] br[98] wl[393] vdd gnd cell_6t
Xbit_r394_c98 bl[98] br[98] wl[394] vdd gnd cell_6t
Xbit_r395_c98 bl[98] br[98] wl[395] vdd gnd cell_6t
Xbit_r396_c98 bl[98] br[98] wl[396] vdd gnd cell_6t
Xbit_r397_c98 bl[98] br[98] wl[397] vdd gnd cell_6t
Xbit_r398_c98 bl[98] br[98] wl[398] vdd gnd cell_6t
Xbit_r399_c98 bl[98] br[98] wl[399] vdd gnd cell_6t
Xbit_r400_c98 bl[98] br[98] wl[400] vdd gnd cell_6t
Xbit_r401_c98 bl[98] br[98] wl[401] vdd gnd cell_6t
Xbit_r402_c98 bl[98] br[98] wl[402] vdd gnd cell_6t
Xbit_r403_c98 bl[98] br[98] wl[403] vdd gnd cell_6t
Xbit_r404_c98 bl[98] br[98] wl[404] vdd gnd cell_6t
Xbit_r405_c98 bl[98] br[98] wl[405] vdd gnd cell_6t
Xbit_r406_c98 bl[98] br[98] wl[406] vdd gnd cell_6t
Xbit_r407_c98 bl[98] br[98] wl[407] vdd gnd cell_6t
Xbit_r408_c98 bl[98] br[98] wl[408] vdd gnd cell_6t
Xbit_r409_c98 bl[98] br[98] wl[409] vdd gnd cell_6t
Xbit_r410_c98 bl[98] br[98] wl[410] vdd gnd cell_6t
Xbit_r411_c98 bl[98] br[98] wl[411] vdd gnd cell_6t
Xbit_r412_c98 bl[98] br[98] wl[412] vdd gnd cell_6t
Xbit_r413_c98 bl[98] br[98] wl[413] vdd gnd cell_6t
Xbit_r414_c98 bl[98] br[98] wl[414] vdd gnd cell_6t
Xbit_r415_c98 bl[98] br[98] wl[415] vdd gnd cell_6t
Xbit_r416_c98 bl[98] br[98] wl[416] vdd gnd cell_6t
Xbit_r417_c98 bl[98] br[98] wl[417] vdd gnd cell_6t
Xbit_r418_c98 bl[98] br[98] wl[418] vdd gnd cell_6t
Xbit_r419_c98 bl[98] br[98] wl[419] vdd gnd cell_6t
Xbit_r420_c98 bl[98] br[98] wl[420] vdd gnd cell_6t
Xbit_r421_c98 bl[98] br[98] wl[421] vdd gnd cell_6t
Xbit_r422_c98 bl[98] br[98] wl[422] vdd gnd cell_6t
Xbit_r423_c98 bl[98] br[98] wl[423] vdd gnd cell_6t
Xbit_r424_c98 bl[98] br[98] wl[424] vdd gnd cell_6t
Xbit_r425_c98 bl[98] br[98] wl[425] vdd gnd cell_6t
Xbit_r426_c98 bl[98] br[98] wl[426] vdd gnd cell_6t
Xbit_r427_c98 bl[98] br[98] wl[427] vdd gnd cell_6t
Xbit_r428_c98 bl[98] br[98] wl[428] vdd gnd cell_6t
Xbit_r429_c98 bl[98] br[98] wl[429] vdd gnd cell_6t
Xbit_r430_c98 bl[98] br[98] wl[430] vdd gnd cell_6t
Xbit_r431_c98 bl[98] br[98] wl[431] vdd gnd cell_6t
Xbit_r432_c98 bl[98] br[98] wl[432] vdd gnd cell_6t
Xbit_r433_c98 bl[98] br[98] wl[433] vdd gnd cell_6t
Xbit_r434_c98 bl[98] br[98] wl[434] vdd gnd cell_6t
Xbit_r435_c98 bl[98] br[98] wl[435] vdd gnd cell_6t
Xbit_r436_c98 bl[98] br[98] wl[436] vdd gnd cell_6t
Xbit_r437_c98 bl[98] br[98] wl[437] vdd gnd cell_6t
Xbit_r438_c98 bl[98] br[98] wl[438] vdd gnd cell_6t
Xbit_r439_c98 bl[98] br[98] wl[439] vdd gnd cell_6t
Xbit_r440_c98 bl[98] br[98] wl[440] vdd gnd cell_6t
Xbit_r441_c98 bl[98] br[98] wl[441] vdd gnd cell_6t
Xbit_r442_c98 bl[98] br[98] wl[442] vdd gnd cell_6t
Xbit_r443_c98 bl[98] br[98] wl[443] vdd gnd cell_6t
Xbit_r444_c98 bl[98] br[98] wl[444] vdd gnd cell_6t
Xbit_r445_c98 bl[98] br[98] wl[445] vdd gnd cell_6t
Xbit_r446_c98 bl[98] br[98] wl[446] vdd gnd cell_6t
Xbit_r447_c98 bl[98] br[98] wl[447] vdd gnd cell_6t
Xbit_r448_c98 bl[98] br[98] wl[448] vdd gnd cell_6t
Xbit_r449_c98 bl[98] br[98] wl[449] vdd gnd cell_6t
Xbit_r450_c98 bl[98] br[98] wl[450] vdd gnd cell_6t
Xbit_r451_c98 bl[98] br[98] wl[451] vdd gnd cell_6t
Xbit_r452_c98 bl[98] br[98] wl[452] vdd gnd cell_6t
Xbit_r453_c98 bl[98] br[98] wl[453] vdd gnd cell_6t
Xbit_r454_c98 bl[98] br[98] wl[454] vdd gnd cell_6t
Xbit_r455_c98 bl[98] br[98] wl[455] vdd gnd cell_6t
Xbit_r456_c98 bl[98] br[98] wl[456] vdd gnd cell_6t
Xbit_r457_c98 bl[98] br[98] wl[457] vdd gnd cell_6t
Xbit_r458_c98 bl[98] br[98] wl[458] vdd gnd cell_6t
Xbit_r459_c98 bl[98] br[98] wl[459] vdd gnd cell_6t
Xbit_r460_c98 bl[98] br[98] wl[460] vdd gnd cell_6t
Xbit_r461_c98 bl[98] br[98] wl[461] vdd gnd cell_6t
Xbit_r462_c98 bl[98] br[98] wl[462] vdd gnd cell_6t
Xbit_r463_c98 bl[98] br[98] wl[463] vdd gnd cell_6t
Xbit_r464_c98 bl[98] br[98] wl[464] vdd gnd cell_6t
Xbit_r465_c98 bl[98] br[98] wl[465] vdd gnd cell_6t
Xbit_r466_c98 bl[98] br[98] wl[466] vdd gnd cell_6t
Xbit_r467_c98 bl[98] br[98] wl[467] vdd gnd cell_6t
Xbit_r468_c98 bl[98] br[98] wl[468] vdd gnd cell_6t
Xbit_r469_c98 bl[98] br[98] wl[469] vdd gnd cell_6t
Xbit_r470_c98 bl[98] br[98] wl[470] vdd gnd cell_6t
Xbit_r471_c98 bl[98] br[98] wl[471] vdd gnd cell_6t
Xbit_r472_c98 bl[98] br[98] wl[472] vdd gnd cell_6t
Xbit_r473_c98 bl[98] br[98] wl[473] vdd gnd cell_6t
Xbit_r474_c98 bl[98] br[98] wl[474] vdd gnd cell_6t
Xbit_r475_c98 bl[98] br[98] wl[475] vdd gnd cell_6t
Xbit_r476_c98 bl[98] br[98] wl[476] vdd gnd cell_6t
Xbit_r477_c98 bl[98] br[98] wl[477] vdd gnd cell_6t
Xbit_r478_c98 bl[98] br[98] wl[478] vdd gnd cell_6t
Xbit_r479_c98 bl[98] br[98] wl[479] vdd gnd cell_6t
Xbit_r480_c98 bl[98] br[98] wl[480] vdd gnd cell_6t
Xbit_r481_c98 bl[98] br[98] wl[481] vdd gnd cell_6t
Xbit_r482_c98 bl[98] br[98] wl[482] vdd gnd cell_6t
Xbit_r483_c98 bl[98] br[98] wl[483] vdd gnd cell_6t
Xbit_r484_c98 bl[98] br[98] wl[484] vdd gnd cell_6t
Xbit_r485_c98 bl[98] br[98] wl[485] vdd gnd cell_6t
Xbit_r486_c98 bl[98] br[98] wl[486] vdd gnd cell_6t
Xbit_r487_c98 bl[98] br[98] wl[487] vdd gnd cell_6t
Xbit_r488_c98 bl[98] br[98] wl[488] vdd gnd cell_6t
Xbit_r489_c98 bl[98] br[98] wl[489] vdd gnd cell_6t
Xbit_r490_c98 bl[98] br[98] wl[490] vdd gnd cell_6t
Xbit_r491_c98 bl[98] br[98] wl[491] vdd gnd cell_6t
Xbit_r492_c98 bl[98] br[98] wl[492] vdd gnd cell_6t
Xbit_r493_c98 bl[98] br[98] wl[493] vdd gnd cell_6t
Xbit_r494_c98 bl[98] br[98] wl[494] vdd gnd cell_6t
Xbit_r495_c98 bl[98] br[98] wl[495] vdd gnd cell_6t
Xbit_r496_c98 bl[98] br[98] wl[496] vdd gnd cell_6t
Xbit_r497_c98 bl[98] br[98] wl[497] vdd gnd cell_6t
Xbit_r498_c98 bl[98] br[98] wl[498] vdd gnd cell_6t
Xbit_r499_c98 bl[98] br[98] wl[499] vdd gnd cell_6t
Xbit_r500_c98 bl[98] br[98] wl[500] vdd gnd cell_6t
Xbit_r501_c98 bl[98] br[98] wl[501] vdd gnd cell_6t
Xbit_r502_c98 bl[98] br[98] wl[502] vdd gnd cell_6t
Xbit_r503_c98 bl[98] br[98] wl[503] vdd gnd cell_6t
Xbit_r504_c98 bl[98] br[98] wl[504] vdd gnd cell_6t
Xbit_r505_c98 bl[98] br[98] wl[505] vdd gnd cell_6t
Xbit_r506_c98 bl[98] br[98] wl[506] vdd gnd cell_6t
Xbit_r507_c98 bl[98] br[98] wl[507] vdd gnd cell_6t
Xbit_r508_c98 bl[98] br[98] wl[508] vdd gnd cell_6t
Xbit_r509_c98 bl[98] br[98] wl[509] vdd gnd cell_6t
Xbit_r510_c98 bl[98] br[98] wl[510] vdd gnd cell_6t
Xbit_r511_c98 bl[98] br[98] wl[511] vdd gnd cell_6t
Xbit_r0_c99 bl[99] br[99] wl[0] vdd gnd cell_6t
Xbit_r1_c99 bl[99] br[99] wl[1] vdd gnd cell_6t
Xbit_r2_c99 bl[99] br[99] wl[2] vdd gnd cell_6t
Xbit_r3_c99 bl[99] br[99] wl[3] vdd gnd cell_6t
Xbit_r4_c99 bl[99] br[99] wl[4] vdd gnd cell_6t
Xbit_r5_c99 bl[99] br[99] wl[5] vdd gnd cell_6t
Xbit_r6_c99 bl[99] br[99] wl[6] vdd gnd cell_6t
Xbit_r7_c99 bl[99] br[99] wl[7] vdd gnd cell_6t
Xbit_r8_c99 bl[99] br[99] wl[8] vdd gnd cell_6t
Xbit_r9_c99 bl[99] br[99] wl[9] vdd gnd cell_6t
Xbit_r10_c99 bl[99] br[99] wl[10] vdd gnd cell_6t
Xbit_r11_c99 bl[99] br[99] wl[11] vdd gnd cell_6t
Xbit_r12_c99 bl[99] br[99] wl[12] vdd gnd cell_6t
Xbit_r13_c99 bl[99] br[99] wl[13] vdd gnd cell_6t
Xbit_r14_c99 bl[99] br[99] wl[14] vdd gnd cell_6t
Xbit_r15_c99 bl[99] br[99] wl[15] vdd gnd cell_6t
Xbit_r16_c99 bl[99] br[99] wl[16] vdd gnd cell_6t
Xbit_r17_c99 bl[99] br[99] wl[17] vdd gnd cell_6t
Xbit_r18_c99 bl[99] br[99] wl[18] vdd gnd cell_6t
Xbit_r19_c99 bl[99] br[99] wl[19] vdd gnd cell_6t
Xbit_r20_c99 bl[99] br[99] wl[20] vdd gnd cell_6t
Xbit_r21_c99 bl[99] br[99] wl[21] vdd gnd cell_6t
Xbit_r22_c99 bl[99] br[99] wl[22] vdd gnd cell_6t
Xbit_r23_c99 bl[99] br[99] wl[23] vdd gnd cell_6t
Xbit_r24_c99 bl[99] br[99] wl[24] vdd gnd cell_6t
Xbit_r25_c99 bl[99] br[99] wl[25] vdd gnd cell_6t
Xbit_r26_c99 bl[99] br[99] wl[26] vdd gnd cell_6t
Xbit_r27_c99 bl[99] br[99] wl[27] vdd gnd cell_6t
Xbit_r28_c99 bl[99] br[99] wl[28] vdd gnd cell_6t
Xbit_r29_c99 bl[99] br[99] wl[29] vdd gnd cell_6t
Xbit_r30_c99 bl[99] br[99] wl[30] vdd gnd cell_6t
Xbit_r31_c99 bl[99] br[99] wl[31] vdd gnd cell_6t
Xbit_r32_c99 bl[99] br[99] wl[32] vdd gnd cell_6t
Xbit_r33_c99 bl[99] br[99] wl[33] vdd gnd cell_6t
Xbit_r34_c99 bl[99] br[99] wl[34] vdd gnd cell_6t
Xbit_r35_c99 bl[99] br[99] wl[35] vdd gnd cell_6t
Xbit_r36_c99 bl[99] br[99] wl[36] vdd gnd cell_6t
Xbit_r37_c99 bl[99] br[99] wl[37] vdd gnd cell_6t
Xbit_r38_c99 bl[99] br[99] wl[38] vdd gnd cell_6t
Xbit_r39_c99 bl[99] br[99] wl[39] vdd gnd cell_6t
Xbit_r40_c99 bl[99] br[99] wl[40] vdd gnd cell_6t
Xbit_r41_c99 bl[99] br[99] wl[41] vdd gnd cell_6t
Xbit_r42_c99 bl[99] br[99] wl[42] vdd gnd cell_6t
Xbit_r43_c99 bl[99] br[99] wl[43] vdd gnd cell_6t
Xbit_r44_c99 bl[99] br[99] wl[44] vdd gnd cell_6t
Xbit_r45_c99 bl[99] br[99] wl[45] vdd gnd cell_6t
Xbit_r46_c99 bl[99] br[99] wl[46] vdd gnd cell_6t
Xbit_r47_c99 bl[99] br[99] wl[47] vdd gnd cell_6t
Xbit_r48_c99 bl[99] br[99] wl[48] vdd gnd cell_6t
Xbit_r49_c99 bl[99] br[99] wl[49] vdd gnd cell_6t
Xbit_r50_c99 bl[99] br[99] wl[50] vdd gnd cell_6t
Xbit_r51_c99 bl[99] br[99] wl[51] vdd gnd cell_6t
Xbit_r52_c99 bl[99] br[99] wl[52] vdd gnd cell_6t
Xbit_r53_c99 bl[99] br[99] wl[53] vdd gnd cell_6t
Xbit_r54_c99 bl[99] br[99] wl[54] vdd gnd cell_6t
Xbit_r55_c99 bl[99] br[99] wl[55] vdd gnd cell_6t
Xbit_r56_c99 bl[99] br[99] wl[56] vdd gnd cell_6t
Xbit_r57_c99 bl[99] br[99] wl[57] vdd gnd cell_6t
Xbit_r58_c99 bl[99] br[99] wl[58] vdd gnd cell_6t
Xbit_r59_c99 bl[99] br[99] wl[59] vdd gnd cell_6t
Xbit_r60_c99 bl[99] br[99] wl[60] vdd gnd cell_6t
Xbit_r61_c99 bl[99] br[99] wl[61] vdd gnd cell_6t
Xbit_r62_c99 bl[99] br[99] wl[62] vdd gnd cell_6t
Xbit_r63_c99 bl[99] br[99] wl[63] vdd gnd cell_6t
Xbit_r64_c99 bl[99] br[99] wl[64] vdd gnd cell_6t
Xbit_r65_c99 bl[99] br[99] wl[65] vdd gnd cell_6t
Xbit_r66_c99 bl[99] br[99] wl[66] vdd gnd cell_6t
Xbit_r67_c99 bl[99] br[99] wl[67] vdd gnd cell_6t
Xbit_r68_c99 bl[99] br[99] wl[68] vdd gnd cell_6t
Xbit_r69_c99 bl[99] br[99] wl[69] vdd gnd cell_6t
Xbit_r70_c99 bl[99] br[99] wl[70] vdd gnd cell_6t
Xbit_r71_c99 bl[99] br[99] wl[71] vdd gnd cell_6t
Xbit_r72_c99 bl[99] br[99] wl[72] vdd gnd cell_6t
Xbit_r73_c99 bl[99] br[99] wl[73] vdd gnd cell_6t
Xbit_r74_c99 bl[99] br[99] wl[74] vdd gnd cell_6t
Xbit_r75_c99 bl[99] br[99] wl[75] vdd gnd cell_6t
Xbit_r76_c99 bl[99] br[99] wl[76] vdd gnd cell_6t
Xbit_r77_c99 bl[99] br[99] wl[77] vdd gnd cell_6t
Xbit_r78_c99 bl[99] br[99] wl[78] vdd gnd cell_6t
Xbit_r79_c99 bl[99] br[99] wl[79] vdd gnd cell_6t
Xbit_r80_c99 bl[99] br[99] wl[80] vdd gnd cell_6t
Xbit_r81_c99 bl[99] br[99] wl[81] vdd gnd cell_6t
Xbit_r82_c99 bl[99] br[99] wl[82] vdd gnd cell_6t
Xbit_r83_c99 bl[99] br[99] wl[83] vdd gnd cell_6t
Xbit_r84_c99 bl[99] br[99] wl[84] vdd gnd cell_6t
Xbit_r85_c99 bl[99] br[99] wl[85] vdd gnd cell_6t
Xbit_r86_c99 bl[99] br[99] wl[86] vdd gnd cell_6t
Xbit_r87_c99 bl[99] br[99] wl[87] vdd gnd cell_6t
Xbit_r88_c99 bl[99] br[99] wl[88] vdd gnd cell_6t
Xbit_r89_c99 bl[99] br[99] wl[89] vdd gnd cell_6t
Xbit_r90_c99 bl[99] br[99] wl[90] vdd gnd cell_6t
Xbit_r91_c99 bl[99] br[99] wl[91] vdd gnd cell_6t
Xbit_r92_c99 bl[99] br[99] wl[92] vdd gnd cell_6t
Xbit_r93_c99 bl[99] br[99] wl[93] vdd gnd cell_6t
Xbit_r94_c99 bl[99] br[99] wl[94] vdd gnd cell_6t
Xbit_r95_c99 bl[99] br[99] wl[95] vdd gnd cell_6t
Xbit_r96_c99 bl[99] br[99] wl[96] vdd gnd cell_6t
Xbit_r97_c99 bl[99] br[99] wl[97] vdd gnd cell_6t
Xbit_r98_c99 bl[99] br[99] wl[98] vdd gnd cell_6t
Xbit_r99_c99 bl[99] br[99] wl[99] vdd gnd cell_6t
Xbit_r100_c99 bl[99] br[99] wl[100] vdd gnd cell_6t
Xbit_r101_c99 bl[99] br[99] wl[101] vdd gnd cell_6t
Xbit_r102_c99 bl[99] br[99] wl[102] vdd gnd cell_6t
Xbit_r103_c99 bl[99] br[99] wl[103] vdd gnd cell_6t
Xbit_r104_c99 bl[99] br[99] wl[104] vdd gnd cell_6t
Xbit_r105_c99 bl[99] br[99] wl[105] vdd gnd cell_6t
Xbit_r106_c99 bl[99] br[99] wl[106] vdd gnd cell_6t
Xbit_r107_c99 bl[99] br[99] wl[107] vdd gnd cell_6t
Xbit_r108_c99 bl[99] br[99] wl[108] vdd gnd cell_6t
Xbit_r109_c99 bl[99] br[99] wl[109] vdd gnd cell_6t
Xbit_r110_c99 bl[99] br[99] wl[110] vdd gnd cell_6t
Xbit_r111_c99 bl[99] br[99] wl[111] vdd gnd cell_6t
Xbit_r112_c99 bl[99] br[99] wl[112] vdd gnd cell_6t
Xbit_r113_c99 bl[99] br[99] wl[113] vdd gnd cell_6t
Xbit_r114_c99 bl[99] br[99] wl[114] vdd gnd cell_6t
Xbit_r115_c99 bl[99] br[99] wl[115] vdd gnd cell_6t
Xbit_r116_c99 bl[99] br[99] wl[116] vdd gnd cell_6t
Xbit_r117_c99 bl[99] br[99] wl[117] vdd gnd cell_6t
Xbit_r118_c99 bl[99] br[99] wl[118] vdd gnd cell_6t
Xbit_r119_c99 bl[99] br[99] wl[119] vdd gnd cell_6t
Xbit_r120_c99 bl[99] br[99] wl[120] vdd gnd cell_6t
Xbit_r121_c99 bl[99] br[99] wl[121] vdd gnd cell_6t
Xbit_r122_c99 bl[99] br[99] wl[122] vdd gnd cell_6t
Xbit_r123_c99 bl[99] br[99] wl[123] vdd gnd cell_6t
Xbit_r124_c99 bl[99] br[99] wl[124] vdd gnd cell_6t
Xbit_r125_c99 bl[99] br[99] wl[125] vdd gnd cell_6t
Xbit_r126_c99 bl[99] br[99] wl[126] vdd gnd cell_6t
Xbit_r127_c99 bl[99] br[99] wl[127] vdd gnd cell_6t
Xbit_r128_c99 bl[99] br[99] wl[128] vdd gnd cell_6t
Xbit_r129_c99 bl[99] br[99] wl[129] vdd gnd cell_6t
Xbit_r130_c99 bl[99] br[99] wl[130] vdd gnd cell_6t
Xbit_r131_c99 bl[99] br[99] wl[131] vdd gnd cell_6t
Xbit_r132_c99 bl[99] br[99] wl[132] vdd gnd cell_6t
Xbit_r133_c99 bl[99] br[99] wl[133] vdd gnd cell_6t
Xbit_r134_c99 bl[99] br[99] wl[134] vdd gnd cell_6t
Xbit_r135_c99 bl[99] br[99] wl[135] vdd gnd cell_6t
Xbit_r136_c99 bl[99] br[99] wl[136] vdd gnd cell_6t
Xbit_r137_c99 bl[99] br[99] wl[137] vdd gnd cell_6t
Xbit_r138_c99 bl[99] br[99] wl[138] vdd gnd cell_6t
Xbit_r139_c99 bl[99] br[99] wl[139] vdd gnd cell_6t
Xbit_r140_c99 bl[99] br[99] wl[140] vdd gnd cell_6t
Xbit_r141_c99 bl[99] br[99] wl[141] vdd gnd cell_6t
Xbit_r142_c99 bl[99] br[99] wl[142] vdd gnd cell_6t
Xbit_r143_c99 bl[99] br[99] wl[143] vdd gnd cell_6t
Xbit_r144_c99 bl[99] br[99] wl[144] vdd gnd cell_6t
Xbit_r145_c99 bl[99] br[99] wl[145] vdd gnd cell_6t
Xbit_r146_c99 bl[99] br[99] wl[146] vdd gnd cell_6t
Xbit_r147_c99 bl[99] br[99] wl[147] vdd gnd cell_6t
Xbit_r148_c99 bl[99] br[99] wl[148] vdd gnd cell_6t
Xbit_r149_c99 bl[99] br[99] wl[149] vdd gnd cell_6t
Xbit_r150_c99 bl[99] br[99] wl[150] vdd gnd cell_6t
Xbit_r151_c99 bl[99] br[99] wl[151] vdd gnd cell_6t
Xbit_r152_c99 bl[99] br[99] wl[152] vdd gnd cell_6t
Xbit_r153_c99 bl[99] br[99] wl[153] vdd gnd cell_6t
Xbit_r154_c99 bl[99] br[99] wl[154] vdd gnd cell_6t
Xbit_r155_c99 bl[99] br[99] wl[155] vdd gnd cell_6t
Xbit_r156_c99 bl[99] br[99] wl[156] vdd gnd cell_6t
Xbit_r157_c99 bl[99] br[99] wl[157] vdd gnd cell_6t
Xbit_r158_c99 bl[99] br[99] wl[158] vdd gnd cell_6t
Xbit_r159_c99 bl[99] br[99] wl[159] vdd gnd cell_6t
Xbit_r160_c99 bl[99] br[99] wl[160] vdd gnd cell_6t
Xbit_r161_c99 bl[99] br[99] wl[161] vdd gnd cell_6t
Xbit_r162_c99 bl[99] br[99] wl[162] vdd gnd cell_6t
Xbit_r163_c99 bl[99] br[99] wl[163] vdd gnd cell_6t
Xbit_r164_c99 bl[99] br[99] wl[164] vdd gnd cell_6t
Xbit_r165_c99 bl[99] br[99] wl[165] vdd gnd cell_6t
Xbit_r166_c99 bl[99] br[99] wl[166] vdd gnd cell_6t
Xbit_r167_c99 bl[99] br[99] wl[167] vdd gnd cell_6t
Xbit_r168_c99 bl[99] br[99] wl[168] vdd gnd cell_6t
Xbit_r169_c99 bl[99] br[99] wl[169] vdd gnd cell_6t
Xbit_r170_c99 bl[99] br[99] wl[170] vdd gnd cell_6t
Xbit_r171_c99 bl[99] br[99] wl[171] vdd gnd cell_6t
Xbit_r172_c99 bl[99] br[99] wl[172] vdd gnd cell_6t
Xbit_r173_c99 bl[99] br[99] wl[173] vdd gnd cell_6t
Xbit_r174_c99 bl[99] br[99] wl[174] vdd gnd cell_6t
Xbit_r175_c99 bl[99] br[99] wl[175] vdd gnd cell_6t
Xbit_r176_c99 bl[99] br[99] wl[176] vdd gnd cell_6t
Xbit_r177_c99 bl[99] br[99] wl[177] vdd gnd cell_6t
Xbit_r178_c99 bl[99] br[99] wl[178] vdd gnd cell_6t
Xbit_r179_c99 bl[99] br[99] wl[179] vdd gnd cell_6t
Xbit_r180_c99 bl[99] br[99] wl[180] vdd gnd cell_6t
Xbit_r181_c99 bl[99] br[99] wl[181] vdd gnd cell_6t
Xbit_r182_c99 bl[99] br[99] wl[182] vdd gnd cell_6t
Xbit_r183_c99 bl[99] br[99] wl[183] vdd gnd cell_6t
Xbit_r184_c99 bl[99] br[99] wl[184] vdd gnd cell_6t
Xbit_r185_c99 bl[99] br[99] wl[185] vdd gnd cell_6t
Xbit_r186_c99 bl[99] br[99] wl[186] vdd gnd cell_6t
Xbit_r187_c99 bl[99] br[99] wl[187] vdd gnd cell_6t
Xbit_r188_c99 bl[99] br[99] wl[188] vdd gnd cell_6t
Xbit_r189_c99 bl[99] br[99] wl[189] vdd gnd cell_6t
Xbit_r190_c99 bl[99] br[99] wl[190] vdd gnd cell_6t
Xbit_r191_c99 bl[99] br[99] wl[191] vdd gnd cell_6t
Xbit_r192_c99 bl[99] br[99] wl[192] vdd gnd cell_6t
Xbit_r193_c99 bl[99] br[99] wl[193] vdd gnd cell_6t
Xbit_r194_c99 bl[99] br[99] wl[194] vdd gnd cell_6t
Xbit_r195_c99 bl[99] br[99] wl[195] vdd gnd cell_6t
Xbit_r196_c99 bl[99] br[99] wl[196] vdd gnd cell_6t
Xbit_r197_c99 bl[99] br[99] wl[197] vdd gnd cell_6t
Xbit_r198_c99 bl[99] br[99] wl[198] vdd gnd cell_6t
Xbit_r199_c99 bl[99] br[99] wl[199] vdd gnd cell_6t
Xbit_r200_c99 bl[99] br[99] wl[200] vdd gnd cell_6t
Xbit_r201_c99 bl[99] br[99] wl[201] vdd gnd cell_6t
Xbit_r202_c99 bl[99] br[99] wl[202] vdd gnd cell_6t
Xbit_r203_c99 bl[99] br[99] wl[203] vdd gnd cell_6t
Xbit_r204_c99 bl[99] br[99] wl[204] vdd gnd cell_6t
Xbit_r205_c99 bl[99] br[99] wl[205] vdd gnd cell_6t
Xbit_r206_c99 bl[99] br[99] wl[206] vdd gnd cell_6t
Xbit_r207_c99 bl[99] br[99] wl[207] vdd gnd cell_6t
Xbit_r208_c99 bl[99] br[99] wl[208] vdd gnd cell_6t
Xbit_r209_c99 bl[99] br[99] wl[209] vdd gnd cell_6t
Xbit_r210_c99 bl[99] br[99] wl[210] vdd gnd cell_6t
Xbit_r211_c99 bl[99] br[99] wl[211] vdd gnd cell_6t
Xbit_r212_c99 bl[99] br[99] wl[212] vdd gnd cell_6t
Xbit_r213_c99 bl[99] br[99] wl[213] vdd gnd cell_6t
Xbit_r214_c99 bl[99] br[99] wl[214] vdd gnd cell_6t
Xbit_r215_c99 bl[99] br[99] wl[215] vdd gnd cell_6t
Xbit_r216_c99 bl[99] br[99] wl[216] vdd gnd cell_6t
Xbit_r217_c99 bl[99] br[99] wl[217] vdd gnd cell_6t
Xbit_r218_c99 bl[99] br[99] wl[218] vdd gnd cell_6t
Xbit_r219_c99 bl[99] br[99] wl[219] vdd gnd cell_6t
Xbit_r220_c99 bl[99] br[99] wl[220] vdd gnd cell_6t
Xbit_r221_c99 bl[99] br[99] wl[221] vdd gnd cell_6t
Xbit_r222_c99 bl[99] br[99] wl[222] vdd gnd cell_6t
Xbit_r223_c99 bl[99] br[99] wl[223] vdd gnd cell_6t
Xbit_r224_c99 bl[99] br[99] wl[224] vdd gnd cell_6t
Xbit_r225_c99 bl[99] br[99] wl[225] vdd gnd cell_6t
Xbit_r226_c99 bl[99] br[99] wl[226] vdd gnd cell_6t
Xbit_r227_c99 bl[99] br[99] wl[227] vdd gnd cell_6t
Xbit_r228_c99 bl[99] br[99] wl[228] vdd gnd cell_6t
Xbit_r229_c99 bl[99] br[99] wl[229] vdd gnd cell_6t
Xbit_r230_c99 bl[99] br[99] wl[230] vdd gnd cell_6t
Xbit_r231_c99 bl[99] br[99] wl[231] vdd gnd cell_6t
Xbit_r232_c99 bl[99] br[99] wl[232] vdd gnd cell_6t
Xbit_r233_c99 bl[99] br[99] wl[233] vdd gnd cell_6t
Xbit_r234_c99 bl[99] br[99] wl[234] vdd gnd cell_6t
Xbit_r235_c99 bl[99] br[99] wl[235] vdd gnd cell_6t
Xbit_r236_c99 bl[99] br[99] wl[236] vdd gnd cell_6t
Xbit_r237_c99 bl[99] br[99] wl[237] vdd gnd cell_6t
Xbit_r238_c99 bl[99] br[99] wl[238] vdd gnd cell_6t
Xbit_r239_c99 bl[99] br[99] wl[239] vdd gnd cell_6t
Xbit_r240_c99 bl[99] br[99] wl[240] vdd gnd cell_6t
Xbit_r241_c99 bl[99] br[99] wl[241] vdd gnd cell_6t
Xbit_r242_c99 bl[99] br[99] wl[242] vdd gnd cell_6t
Xbit_r243_c99 bl[99] br[99] wl[243] vdd gnd cell_6t
Xbit_r244_c99 bl[99] br[99] wl[244] vdd gnd cell_6t
Xbit_r245_c99 bl[99] br[99] wl[245] vdd gnd cell_6t
Xbit_r246_c99 bl[99] br[99] wl[246] vdd gnd cell_6t
Xbit_r247_c99 bl[99] br[99] wl[247] vdd gnd cell_6t
Xbit_r248_c99 bl[99] br[99] wl[248] vdd gnd cell_6t
Xbit_r249_c99 bl[99] br[99] wl[249] vdd gnd cell_6t
Xbit_r250_c99 bl[99] br[99] wl[250] vdd gnd cell_6t
Xbit_r251_c99 bl[99] br[99] wl[251] vdd gnd cell_6t
Xbit_r252_c99 bl[99] br[99] wl[252] vdd gnd cell_6t
Xbit_r253_c99 bl[99] br[99] wl[253] vdd gnd cell_6t
Xbit_r254_c99 bl[99] br[99] wl[254] vdd gnd cell_6t
Xbit_r255_c99 bl[99] br[99] wl[255] vdd gnd cell_6t
Xbit_r256_c99 bl[99] br[99] wl[256] vdd gnd cell_6t
Xbit_r257_c99 bl[99] br[99] wl[257] vdd gnd cell_6t
Xbit_r258_c99 bl[99] br[99] wl[258] vdd gnd cell_6t
Xbit_r259_c99 bl[99] br[99] wl[259] vdd gnd cell_6t
Xbit_r260_c99 bl[99] br[99] wl[260] vdd gnd cell_6t
Xbit_r261_c99 bl[99] br[99] wl[261] vdd gnd cell_6t
Xbit_r262_c99 bl[99] br[99] wl[262] vdd gnd cell_6t
Xbit_r263_c99 bl[99] br[99] wl[263] vdd gnd cell_6t
Xbit_r264_c99 bl[99] br[99] wl[264] vdd gnd cell_6t
Xbit_r265_c99 bl[99] br[99] wl[265] vdd gnd cell_6t
Xbit_r266_c99 bl[99] br[99] wl[266] vdd gnd cell_6t
Xbit_r267_c99 bl[99] br[99] wl[267] vdd gnd cell_6t
Xbit_r268_c99 bl[99] br[99] wl[268] vdd gnd cell_6t
Xbit_r269_c99 bl[99] br[99] wl[269] vdd gnd cell_6t
Xbit_r270_c99 bl[99] br[99] wl[270] vdd gnd cell_6t
Xbit_r271_c99 bl[99] br[99] wl[271] vdd gnd cell_6t
Xbit_r272_c99 bl[99] br[99] wl[272] vdd gnd cell_6t
Xbit_r273_c99 bl[99] br[99] wl[273] vdd gnd cell_6t
Xbit_r274_c99 bl[99] br[99] wl[274] vdd gnd cell_6t
Xbit_r275_c99 bl[99] br[99] wl[275] vdd gnd cell_6t
Xbit_r276_c99 bl[99] br[99] wl[276] vdd gnd cell_6t
Xbit_r277_c99 bl[99] br[99] wl[277] vdd gnd cell_6t
Xbit_r278_c99 bl[99] br[99] wl[278] vdd gnd cell_6t
Xbit_r279_c99 bl[99] br[99] wl[279] vdd gnd cell_6t
Xbit_r280_c99 bl[99] br[99] wl[280] vdd gnd cell_6t
Xbit_r281_c99 bl[99] br[99] wl[281] vdd gnd cell_6t
Xbit_r282_c99 bl[99] br[99] wl[282] vdd gnd cell_6t
Xbit_r283_c99 bl[99] br[99] wl[283] vdd gnd cell_6t
Xbit_r284_c99 bl[99] br[99] wl[284] vdd gnd cell_6t
Xbit_r285_c99 bl[99] br[99] wl[285] vdd gnd cell_6t
Xbit_r286_c99 bl[99] br[99] wl[286] vdd gnd cell_6t
Xbit_r287_c99 bl[99] br[99] wl[287] vdd gnd cell_6t
Xbit_r288_c99 bl[99] br[99] wl[288] vdd gnd cell_6t
Xbit_r289_c99 bl[99] br[99] wl[289] vdd gnd cell_6t
Xbit_r290_c99 bl[99] br[99] wl[290] vdd gnd cell_6t
Xbit_r291_c99 bl[99] br[99] wl[291] vdd gnd cell_6t
Xbit_r292_c99 bl[99] br[99] wl[292] vdd gnd cell_6t
Xbit_r293_c99 bl[99] br[99] wl[293] vdd gnd cell_6t
Xbit_r294_c99 bl[99] br[99] wl[294] vdd gnd cell_6t
Xbit_r295_c99 bl[99] br[99] wl[295] vdd gnd cell_6t
Xbit_r296_c99 bl[99] br[99] wl[296] vdd gnd cell_6t
Xbit_r297_c99 bl[99] br[99] wl[297] vdd gnd cell_6t
Xbit_r298_c99 bl[99] br[99] wl[298] vdd gnd cell_6t
Xbit_r299_c99 bl[99] br[99] wl[299] vdd gnd cell_6t
Xbit_r300_c99 bl[99] br[99] wl[300] vdd gnd cell_6t
Xbit_r301_c99 bl[99] br[99] wl[301] vdd gnd cell_6t
Xbit_r302_c99 bl[99] br[99] wl[302] vdd gnd cell_6t
Xbit_r303_c99 bl[99] br[99] wl[303] vdd gnd cell_6t
Xbit_r304_c99 bl[99] br[99] wl[304] vdd gnd cell_6t
Xbit_r305_c99 bl[99] br[99] wl[305] vdd gnd cell_6t
Xbit_r306_c99 bl[99] br[99] wl[306] vdd gnd cell_6t
Xbit_r307_c99 bl[99] br[99] wl[307] vdd gnd cell_6t
Xbit_r308_c99 bl[99] br[99] wl[308] vdd gnd cell_6t
Xbit_r309_c99 bl[99] br[99] wl[309] vdd gnd cell_6t
Xbit_r310_c99 bl[99] br[99] wl[310] vdd gnd cell_6t
Xbit_r311_c99 bl[99] br[99] wl[311] vdd gnd cell_6t
Xbit_r312_c99 bl[99] br[99] wl[312] vdd gnd cell_6t
Xbit_r313_c99 bl[99] br[99] wl[313] vdd gnd cell_6t
Xbit_r314_c99 bl[99] br[99] wl[314] vdd gnd cell_6t
Xbit_r315_c99 bl[99] br[99] wl[315] vdd gnd cell_6t
Xbit_r316_c99 bl[99] br[99] wl[316] vdd gnd cell_6t
Xbit_r317_c99 bl[99] br[99] wl[317] vdd gnd cell_6t
Xbit_r318_c99 bl[99] br[99] wl[318] vdd gnd cell_6t
Xbit_r319_c99 bl[99] br[99] wl[319] vdd gnd cell_6t
Xbit_r320_c99 bl[99] br[99] wl[320] vdd gnd cell_6t
Xbit_r321_c99 bl[99] br[99] wl[321] vdd gnd cell_6t
Xbit_r322_c99 bl[99] br[99] wl[322] vdd gnd cell_6t
Xbit_r323_c99 bl[99] br[99] wl[323] vdd gnd cell_6t
Xbit_r324_c99 bl[99] br[99] wl[324] vdd gnd cell_6t
Xbit_r325_c99 bl[99] br[99] wl[325] vdd gnd cell_6t
Xbit_r326_c99 bl[99] br[99] wl[326] vdd gnd cell_6t
Xbit_r327_c99 bl[99] br[99] wl[327] vdd gnd cell_6t
Xbit_r328_c99 bl[99] br[99] wl[328] vdd gnd cell_6t
Xbit_r329_c99 bl[99] br[99] wl[329] vdd gnd cell_6t
Xbit_r330_c99 bl[99] br[99] wl[330] vdd gnd cell_6t
Xbit_r331_c99 bl[99] br[99] wl[331] vdd gnd cell_6t
Xbit_r332_c99 bl[99] br[99] wl[332] vdd gnd cell_6t
Xbit_r333_c99 bl[99] br[99] wl[333] vdd gnd cell_6t
Xbit_r334_c99 bl[99] br[99] wl[334] vdd gnd cell_6t
Xbit_r335_c99 bl[99] br[99] wl[335] vdd gnd cell_6t
Xbit_r336_c99 bl[99] br[99] wl[336] vdd gnd cell_6t
Xbit_r337_c99 bl[99] br[99] wl[337] vdd gnd cell_6t
Xbit_r338_c99 bl[99] br[99] wl[338] vdd gnd cell_6t
Xbit_r339_c99 bl[99] br[99] wl[339] vdd gnd cell_6t
Xbit_r340_c99 bl[99] br[99] wl[340] vdd gnd cell_6t
Xbit_r341_c99 bl[99] br[99] wl[341] vdd gnd cell_6t
Xbit_r342_c99 bl[99] br[99] wl[342] vdd gnd cell_6t
Xbit_r343_c99 bl[99] br[99] wl[343] vdd gnd cell_6t
Xbit_r344_c99 bl[99] br[99] wl[344] vdd gnd cell_6t
Xbit_r345_c99 bl[99] br[99] wl[345] vdd gnd cell_6t
Xbit_r346_c99 bl[99] br[99] wl[346] vdd gnd cell_6t
Xbit_r347_c99 bl[99] br[99] wl[347] vdd gnd cell_6t
Xbit_r348_c99 bl[99] br[99] wl[348] vdd gnd cell_6t
Xbit_r349_c99 bl[99] br[99] wl[349] vdd gnd cell_6t
Xbit_r350_c99 bl[99] br[99] wl[350] vdd gnd cell_6t
Xbit_r351_c99 bl[99] br[99] wl[351] vdd gnd cell_6t
Xbit_r352_c99 bl[99] br[99] wl[352] vdd gnd cell_6t
Xbit_r353_c99 bl[99] br[99] wl[353] vdd gnd cell_6t
Xbit_r354_c99 bl[99] br[99] wl[354] vdd gnd cell_6t
Xbit_r355_c99 bl[99] br[99] wl[355] vdd gnd cell_6t
Xbit_r356_c99 bl[99] br[99] wl[356] vdd gnd cell_6t
Xbit_r357_c99 bl[99] br[99] wl[357] vdd gnd cell_6t
Xbit_r358_c99 bl[99] br[99] wl[358] vdd gnd cell_6t
Xbit_r359_c99 bl[99] br[99] wl[359] vdd gnd cell_6t
Xbit_r360_c99 bl[99] br[99] wl[360] vdd gnd cell_6t
Xbit_r361_c99 bl[99] br[99] wl[361] vdd gnd cell_6t
Xbit_r362_c99 bl[99] br[99] wl[362] vdd gnd cell_6t
Xbit_r363_c99 bl[99] br[99] wl[363] vdd gnd cell_6t
Xbit_r364_c99 bl[99] br[99] wl[364] vdd gnd cell_6t
Xbit_r365_c99 bl[99] br[99] wl[365] vdd gnd cell_6t
Xbit_r366_c99 bl[99] br[99] wl[366] vdd gnd cell_6t
Xbit_r367_c99 bl[99] br[99] wl[367] vdd gnd cell_6t
Xbit_r368_c99 bl[99] br[99] wl[368] vdd gnd cell_6t
Xbit_r369_c99 bl[99] br[99] wl[369] vdd gnd cell_6t
Xbit_r370_c99 bl[99] br[99] wl[370] vdd gnd cell_6t
Xbit_r371_c99 bl[99] br[99] wl[371] vdd gnd cell_6t
Xbit_r372_c99 bl[99] br[99] wl[372] vdd gnd cell_6t
Xbit_r373_c99 bl[99] br[99] wl[373] vdd gnd cell_6t
Xbit_r374_c99 bl[99] br[99] wl[374] vdd gnd cell_6t
Xbit_r375_c99 bl[99] br[99] wl[375] vdd gnd cell_6t
Xbit_r376_c99 bl[99] br[99] wl[376] vdd gnd cell_6t
Xbit_r377_c99 bl[99] br[99] wl[377] vdd gnd cell_6t
Xbit_r378_c99 bl[99] br[99] wl[378] vdd gnd cell_6t
Xbit_r379_c99 bl[99] br[99] wl[379] vdd gnd cell_6t
Xbit_r380_c99 bl[99] br[99] wl[380] vdd gnd cell_6t
Xbit_r381_c99 bl[99] br[99] wl[381] vdd gnd cell_6t
Xbit_r382_c99 bl[99] br[99] wl[382] vdd gnd cell_6t
Xbit_r383_c99 bl[99] br[99] wl[383] vdd gnd cell_6t
Xbit_r384_c99 bl[99] br[99] wl[384] vdd gnd cell_6t
Xbit_r385_c99 bl[99] br[99] wl[385] vdd gnd cell_6t
Xbit_r386_c99 bl[99] br[99] wl[386] vdd gnd cell_6t
Xbit_r387_c99 bl[99] br[99] wl[387] vdd gnd cell_6t
Xbit_r388_c99 bl[99] br[99] wl[388] vdd gnd cell_6t
Xbit_r389_c99 bl[99] br[99] wl[389] vdd gnd cell_6t
Xbit_r390_c99 bl[99] br[99] wl[390] vdd gnd cell_6t
Xbit_r391_c99 bl[99] br[99] wl[391] vdd gnd cell_6t
Xbit_r392_c99 bl[99] br[99] wl[392] vdd gnd cell_6t
Xbit_r393_c99 bl[99] br[99] wl[393] vdd gnd cell_6t
Xbit_r394_c99 bl[99] br[99] wl[394] vdd gnd cell_6t
Xbit_r395_c99 bl[99] br[99] wl[395] vdd gnd cell_6t
Xbit_r396_c99 bl[99] br[99] wl[396] vdd gnd cell_6t
Xbit_r397_c99 bl[99] br[99] wl[397] vdd gnd cell_6t
Xbit_r398_c99 bl[99] br[99] wl[398] vdd gnd cell_6t
Xbit_r399_c99 bl[99] br[99] wl[399] vdd gnd cell_6t
Xbit_r400_c99 bl[99] br[99] wl[400] vdd gnd cell_6t
Xbit_r401_c99 bl[99] br[99] wl[401] vdd gnd cell_6t
Xbit_r402_c99 bl[99] br[99] wl[402] vdd gnd cell_6t
Xbit_r403_c99 bl[99] br[99] wl[403] vdd gnd cell_6t
Xbit_r404_c99 bl[99] br[99] wl[404] vdd gnd cell_6t
Xbit_r405_c99 bl[99] br[99] wl[405] vdd gnd cell_6t
Xbit_r406_c99 bl[99] br[99] wl[406] vdd gnd cell_6t
Xbit_r407_c99 bl[99] br[99] wl[407] vdd gnd cell_6t
Xbit_r408_c99 bl[99] br[99] wl[408] vdd gnd cell_6t
Xbit_r409_c99 bl[99] br[99] wl[409] vdd gnd cell_6t
Xbit_r410_c99 bl[99] br[99] wl[410] vdd gnd cell_6t
Xbit_r411_c99 bl[99] br[99] wl[411] vdd gnd cell_6t
Xbit_r412_c99 bl[99] br[99] wl[412] vdd gnd cell_6t
Xbit_r413_c99 bl[99] br[99] wl[413] vdd gnd cell_6t
Xbit_r414_c99 bl[99] br[99] wl[414] vdd gnd cell_6t
Xbit_r415_c99 bl[99] br[99] wl[415] vdd gnd cell_6t
Xbit_r416_c99 bl[99] br[99] wl[416] vdd gnd cell_6t
Xbit_r417_c99 bl[99] br[99] wl[417] vdd gnd cell_6t
Xbit_r418_c99 bl[99] br[99] wl[418] vdd gnd cell_6t
Xbit_r419_c99 bl[99] br[99] wl[419] vdd gnd cell_6t
Xbit_r420_c99 bl[99] br[99] wl[420] vdd gnd cell_6t
Xbit_r421_c99 bl[99] br[99] wl[421] vdd gnd cell_6t
Xbit_r422_c99 bl[99] br[99] wl[422] vdd gnd cell_6t
Xbit_r423_c99 bl[99] br[99] wl[423] vdd gnd cell_6t
Xbit_r424_c99 bl[99] br[99] wl[424] vdd gnd cell_6t
Xbit_r425_c99 bl[99] br[99] wl[425] vdd gnd cell_6t
Xbit_r426_c99 bl[99] br[99] wl[426] vdd gnd cell_6t
Xbit_r427_c99 bl[99] br[99] wl[427] vdd gnd cell_6t
Xbit_r428_c99 bl[99] br[99] wl[428] vdd gnd cell_6t
Xbit_r429_c99 bl[99] br[99] wl[429] vdd gnd cell_6t
Xbit_r430_c99 bl[99] br[99] wl[430] vdd gnd cell_6t
Xbit_r431_c99 bl[99] br[99] wl[431] vdd gnd cell_6t
Xbit_r432_c99 bl[99] br[99] wl[432] vdd gnd cell_6t
Xbit_r433_c99 bl[99] br[99] wl[433] vdd gnd cell_6t
Xbit_r434_c99 bl[99] br[99] wl[434] vdd gnd cell_6t
Xbit_r435_c99 bl[99] br[99] wl[435] vdd gnd cell_6t
Xbit_r436_c99 bl[99] br[99] wl[436] vdd gnd cell_6t
Xbit_r437_c99 bl[99] br[99] wl[437] vdd gnd cell_6t
Xbit_r438_c99 bl[99] br[99] wl[438] vdd gnd cell_6t
Xbit_r439_c99 bl[99] br[99] wl[439] vdd gnd cell_6t
Xbit_r440_c99 bl[99] br[99] wl[440] vdd gnd cell_6t
Xbit_r441_c99 bl[99] br[99] wl[441] vdd gnd cell_6t
Xbit_r442_c99 bl[99] br[99] wl[442] vdd gnd cell_6t
Xbit_r443_c99 bl[99] br[99] wl[443] vdd gnd cell_6t
Xbit_r444_c99 bl[99] br[99] wl[444] vdd gnd cell_6t
Xbit_r445_c99 bl[99] br[99] wl[445] vdd gnd cell_6t
Xbit_r446_c99 bl[99] br[99] wl[446] vdd gnd cell_6t
Xbit_r447_c99 bl[99] br[99] wl[447] vdd gnd cell_6t
Xbit_r448_c99 bl[99] br[99] wl[448] vdd gnd cell_6t
Xbit_r449_c99 bl[99] br[99] wl[449] vdd gnd cell_6t
Xbit_r450_c99 bl[99] br[99] wl[450] vdd gnd cell_6t
Xbit_r451_c99 bl[99] br[99] wl[451] vdd gnd cell_6t
Xbit_r452_c99 bl[99] br[99] wl[452] vdd gnd cell_6t
Xbit_r453_c99 bl[99] br[99] wl[453] vdd gnd cell_6t
Xbit_r454_c99 bl[99] br[99] wl[454] vdd gnd cell_6t
Xbit_r455_c99 bl[99] br[99] wl[455] vdd gnd cell_6t
Xbit_r456_c99 bl[99] br[99] wl[456] vdd gnd cell_6t
Xbit_r457_c99 bl[99] br[99] wl[457] vdd gnd cell_6t
Xbit_r458_c99 bl[99] br[99] wl[458] vdd gnd cell_6t
Xbit_r459_c99 bl[99] br[99] wl[459] vdd gnd cell_6t
Xbit_r460_c99 bl[99] br[99] wl[460] vdd gnd cell_6t
Xbit_r461_c99 bl[99] br[99] wl[461] vdd gnd cell_6t
Xbit_r462_c99 bl[99] br[99] wl[462] vdd gnd cell_6t
Xbit_r463_c99 bl[99] br[99] wl[463] vdd gnd cell_6t
Xbit_r464_c99 bl[99] br[99] wl[464] vdd gnd cell_6t
Xbit_r465_c99 bl[99] br[99] wl[465] vdd gnd cell_6t
Xbit_r466_c99 bl[99] br[99] wl[466] vdd gnd cell_6t
Xbit_r467_c99 bl[99] br[99] wl[467] vdd gnd cell_6t
Xbit_r468_c99 bl[99] br[99] wl[468] vdd gnd cell_6t
Xbit_r469_c99 bl[99] br[99] wl[469] vdd gnd cell_6t
Xbit_r470_c99 bl[99] br[99] wl[470] vdd gnd cell_6t
Xbit_r471_c99 bl[99] br[99] wl[471] vdd gnd cell_6t
Xbit_r472_c99 bl[99] br[99] wl[472] vdd gnd cell_6t
Xbit_r473_c99 bl[99] br[99] wl[473] vdd gnd cell_6t
Xbit_r474_c99 bl[99] br[99] wl[474] vdd gnd cell_6t
Xbit_r475_c99 bl[99] br[99] wl[475] vdd gnd cell_6t
Xbit_r476_c99 bl[99] br[99] wl[476] vdd gnd cell_6t
Xbit_r477_c99 bl[99] br[99] wl[477] vdd gnd cell_6t
Xbit_r478_c99 bl[99] br[99] wl[478] vdd gnd cell_6t
Xbit_r479_c99 bl[99] br[99] wl[479] vdd gnd cell_6t
Xbit_r480_c99 bl[99] br[99] wl[480] vdd gnd cell_6t
Xbit_r481_c99 bl[99] br[99] wl[481] vdd gnd cell_6t
Xbit_r482_c99 bl[99] br[99] wl[482] vdd gnd cell_6t
Xbit_r483_c99 bl[99] br[99] wl[483] vdd gnd cell_6t
Xbit_r484_c99 bl[99] br[99] wl[484] vdd gnd cell_6t
Xbit_r485_c99 bl[99] br[99] wl[485] vdd gnd cell_6t
Xbit_r486_c99 bl[99] br[99] wl[486] vdd gnd cell_6t
Xbit_r487_c99 bl[99] br[99] wl[487] vdd gnd cell_6t
Xbit_r488_c99 bl[99] br[99] wl[488] vdd gnd cell_6t
Xbit_r489_c99 bl[99] br[99] wl[489] vdd gnd cell_6t
Xbit_r490_c99 bl[99] br[99] wl[490] vdd gnd cell_6t
Xbit_r491_c99 bl[99] br[99] wl[491] vdd gnd cell_6t
Xbit_r492_c99 bl[99] br[99] wl[492] vdd gnd cell_6t
Xbit_r493_c99 bl[99] br[99] wl[493] vdd gnd cell_6t
Xbit_r494_c99 bl[99] br[99] wl[494] vdd gnd cell_6t
Xbit_r495_c99 bl[99] br[99] wl[495] vdd gnd cell_6t
Xbit_r496_c99 bl[99] br[99] wl[496] vdd gnd cell_6t
Xbit_r497_c99 bl[99] br[99] wl[497] vdd gnd cell_6t
Xbit_r498_c99 bl[99] br[99] wl[498] vdd gnd cell_6t
Xbit_r499_c99 bl[99] br[99] wl[499] vdd gnd cell_6t
Xbit_r500_c99 bl[99] br[99] wl[500] vdd gnd cell_6t
Xbit_r501_c99 bl[99] br[99] wl[501] vdd gnd cell_6t
Xbit_r502_c99 bl[99] br[99] wl[502] vdd gnd cell_6t
Xbit_r503_c99 bl[99] br[99] wl[503] vdd gnd cell_6t
Xbit_r504_c99 bl[99] br[99] wl[504] vdd gnd cell_6t
Xbit_r505_c99 bl[99] br[99] wl[505] vdd gnd cell_6t
Xbit_r506_c99 bl[99] br[99] wl[506] vdd gnd cell_6t
Xbit_r507_c99 bl[99] br[99] wl[507] vdd gnd cell_6t
Xbit_r508_c99 bl[99] br[99] wl[508] vdd gnd cell_6t
Xbit_r509_c99 bl[99] br[99] wl[509] vdd gnd cell_6t
Xbit_r510_c99 bl[99] br[99] wl[510] vdd gnd cell_6t
Xbit_r511_c99 bl[99] br[99] wl[511] vdd gnd cell_6t
Xbit_r0_c100 bl[100] br[100] wl[0] vdd gnd cell_6t
Xbit_r1_c100 bl[100] br[100] wl[1] vdd gnd cell_6t
Xbit_r2_c100 bl[100] br[100] wl[2] vdd gnd cell_6t
Xbit_r3_c100 bl[100] br[100] wl[3] vdd gnd cell_6t
Xbit_r4_c100 bl[100] br[100] wl[4] vdd gnd cell_6t
Xbit_r5_c100 bl[100] br[100] wl[5] vdd gnd cell_6t
Xbit_r6_c100 bl[100] br[100] wl[6] vdd gnd cell_6t
Xbit_r7_c100 bl[100] br[100] wl[7] vdd gnd cell_6t
Xbit_r8_c100 bl[100] br[100] wl[8] vdd gnd cell_6t
Xbit_r9_c100 bl[100] br[100] wl[9] vdd gnd cell_6t
Xbit_r10_c100 bl[100] br[100] wl[10] vdd gnd cell_6t
Xbit_r11_c100 bl[100] br[100] wl[11] vdd gnd cell_6t
Xbit_r12_c100 bl[100] br[100] wl[12] vdd gnd cell_6t
Xbit_r13_c100 bl[100] br[100] wl[13] vdd gnd cell_6t
Xbit_r14_c100 bl[100] br[100] wl[14] vdd gnd cell_6t
Xbit_r15_c100 bl[100] br[100] wl[15] vdd gnd cell_6t
Xbit_r16_c100 bl[100] br[100] wl[16] vdd gnd cell_6t
Xbit_r17_c100 bl[100] br[100] wl[17] vdd gnd cell_6t
Xbit_r18_c100 bl[100] br[100] wl[18] vdd gnd cell_6t
Xbit_r19_c100 bl[100] br[100] wl[19] vdd gnd cell_6t
Xbit_r20_c100 bl[100] br[100] wl[20] vdd gnd cell_6t
Xbit_r21_c100 bl[100] br[100] wl[21] vdd gnd cell_6t
Xbit_r22_c100 bl[100] br[100] wl[22] vdd gnd cell_6t
Xbit_r23_c100 bl[100] br[100] wl[23] vdd gnd cell_6t
Xbit_r24_c100 bl[100] br[100] wl[24] vdd gnd cell_6t
Xbit_r25_c100 bl[100] br[100] wl[25] vdd gnd cell_6t
Xbit_r26_c100 bl[100] br[100] wl[26] vdd gnd cell_6t
Xbit_r27_c100 bl[100] br[100] wl[27] vdd gnd cell_6t
Xbit_r28_c100 bl[100] br[100] wl[28] vdd gnd cell_6t
Xbit_r29_c100 bl[100] br[100] wl[29] vdd gnd cell_6t
Xbit_r30_c100 bl[100] br[100] wl[30] vdd gnd cell_6t
Xbit_r31_c100 bl[100] br[100] wl[31] vdd gnd cell_6t
Xbit_r32_c100 bl[100] br[100] wl[32] vdd gnd cell_6t
Xbit_r33_c100 bl[100] br[100] wl[33] vdd gnd cell_6t
Xbit_r34_c100 bl[100] br[100] wl[34] vdd gnd cell_6t
Xbit_r35_c100 bl[100] br[100] wl[35] vdd gnd cell_6t
Xbit_r36_c100 bl[100] br[100] wl[36] vdd gnd cell_6t
Xbit_r37_c100 bl[100] br[100] wl[37] vdd gnd cell_6t
Xbit_r38_c100 bl[100] br[100] wl[38] vdd gnd cell_6t
Xbit_r39_c100 bl[100] br[100] wl[39] vdd gnd cell_6t
Xbit_r40_c100 bl[100] br[100] wl[40] vdd gnd cell_6t
Xbit_r41_c100 bl[100] br[100] wl[41] vdd gnd cell_6t
Xbit_r42_c100 bl[100] br[100] wl[42] vdd gnd cell_6t
Xbit_r43_c100 bl[100] br[100] wl[43] vdd gnd cell_6t
Xbit_r44_c100 bl[100] br[100] wl[44] vdd gnd cell_6t
Xbit_r45_c100 bl[100] br[100] wl[45] vdd gnd cell_6t
Xbit_r46_c100 bl[100] br[100] wl[46] vdd gnd cell_6t
Xbit_r47_c100 bl[100] br[100] wl[47] vdd gnd cell_6t
Xbit_r48_c100 bl[100] br[100] wl[48] vdd gnd cell_6t
Xbit_r49_c100 bl[100] br[100] wl[49] vdd gnd cell_6t
Xbit_r50_c100 bl[100] br[100] wl[50] vdd gnd cell_6t
Xbit_r51_c100 bl[100] br[100] wl[51] vdd gnd cell_6t
Xbit_r52_c100 bl[100] br[100] wl[52] vdd gnd cell_6t
Xbit_r53_c100 bl[100] br[100] wl[53] vdd gnd cell_6t
Xbit_r54_c100 bl[100] br[100] wl[54] vdd gnd cell_6t
Xbit_r55_c100 bl[100] br[100] wl[55] vdd gnd cell_6t
Xbit_r56_c100 bl[100] br[100] wl[56] vdd gnd cell_6t
Xbit_r57_c100 bl[100] br[100] wl[57] vdd gnd cell_6t
Xbit_r58_c100 bl[100] br[100] wl[58] vdd gnd cell_6t
Xbit_r59_c100 bl[100] br[100] wl[59] vdd gnd cell_6t
Xbit_r60_c100 bl[100] br[100] wl[60] vdd gnd cell_6t
Xbit_r61_c100 bl[100] br[100] wl[61] vdd gnd cell_6t
Xbit_r62_c100 bl[100] br[100] wl[62] vdd gnd cell_6t
Xbit_r63_c100 bl[100] br[100] wl[63] vdd gnd cell_6t
Xbit_r64_c100 bl[100] br[100] wl[64] vdd gnd cell_6t
Xbit_r65_c100 bl[100] br[100] wl[65] vdd gnd cell_6t
Xbit_r66_c100 bl[100] br[100] wl[66] vdd gnd cell_6t
Xbit_r67_c100 bl[100] br[100] wl[67] vdd gnd cell_6t
Xbit_r68_c100 bl[100] br[100] wl[68] vdd gnd cell_6t
Xbit_r69_c100 bl[100] br[100] wl[69] vdd gnd cell_6t
Xbit_r70_c100 bl[100] br[100] wl[70] vdd gnd cell_6t
Xbit_r71_c100 bl[100] br[100] wl[71] vdd gnd cell_6t
Xbit_r72_c100 bl[100] br[100] wl[72] vdd gnd cell_6t
Xbit_r73_c100 bl[100] br[100] wl[73] vdd gnd cell_6t
Xbit_r74_c100 bl[100] br[100] wl[74] vdd gnd cell_6t
Xbit_r75_c100 bl[100] br[100] wl[75] vdd gnd cell_6t
Xbit_r76_c100 bl[100] br[100] wl[76] vdd gnd cell_6t
Xbit_r77_c100 bl[100] br[100] wl[77] vdd gnd cell_6t
Xbit_r78_c100 bl[100] br[100] wl[78] vdd gnd cell_6t
Xbit_r79_c100 bl[100] br[100] wl[79] vdd gnd cell_6t
Xbit_r80_c100 bl[100] br[100] wl[80] vdd gnd cell_6t
Xbit_r81_c100 bl[100] br[100] wl[81] vdd gnd cell_6t
Xbit_r82_c100 bl[100] br[100] wl[82] vdd gnd cell_6t
Xbit_r83_c100 bl[100] br[100] wl[83] vdd gnd cell_6t
Xbit_r84_c100 bl[100] br[100] wl[84] vdd gnd cell_6t
Xbit_r85_c100 bl[100] br[100] wl[85] vdd gnd cell_6t
Xbit_r86_c100 bl[100] br[100] wl[86] vdd gnd cell_6t
Xbit_r87_c100 bl[100] br[100] wl[87] vdd gnd cell_6t
Xbit_r88_c100 bl[100] br[100] wl[88] vdd gnd cell_6t
Xbit_r89_c100 bl[100] br[100] wl[89] vdd gnd cell_6t
Xbit_r90_c100 bl[100] br[100] wl[90] vdd gnd cell_6t
Xbit_r91_c100 bl[100] br[100] wl[91] vdd gnd cell_6t
Xbit_r92_c100 bl[100] br[100] wl[92] vdd gnd cell_6t
Xbit_r93_c100 bl[100] br[100] wl[93] vdd gnd cell_6t
Xbit_r94_c100 bl[100] br[100] wl[94] vdd gnd cell_6t
Xbit_r95_c100 bl[100] br[100] wl[95] vdd gnd cell_6t
Xbit_r96_c100 bl[100] br[100] wl[96] vdd gnd cell_6t
Xbit_r97_c100 bl[100] br[100] wl[97] vdd gnd cell_6t
Xbit_r98_c100 bl[100] br[100] wl[98] vdd gnd cell_6t
Xbit_r99_c100 bl[100] br[100] wl[99] vdd gnd cell_6t
Xbit_r100_c100 bl[100] br[100] wl[100] vdd gnd cell_6t
Xbit_r101_c100 bl[100] br[100] wl[101] vdd gnd cell_6t
Xbit_r102_c100 bl[100] br[100] wl[102] vdd gnd cell_6t
Xbit_r103_c100 bl[100] br[100] wl[103] vdd gnd cell_6t
Xbit_r104_c100 bl[100] br[100] wl[104] vdd gnd cell_6t
Xbit_r105_c100 bl[100] br[100] wl[105] vdd gnd cell_6t
Xbit_r106_c100 bl[100] br[100] wl[106] vdd gnd cell_6t
Xbit_r107_c100 bl[100] br[100] wl[107] vdd gnd cell_6t
Xbit_r108_c100 bl[100] br[100] wl[108] vdd gnd cell_6t
Xbit_r109_c100 bl[100] br[100] wl[109] vdd gnd cell_6t
Xbit_r110_c100 bl[100] br[100] wl[110] vdd gnd cell_6t
Xbit_r111_c100 bl[100] br[100] wl[111] vdd gnd cell_6t
Xbit_r112_c100 bl[100] br[100] wl[112] vdd gnd cell_6t
Xbit_r113_c100 bl[100] br[100] wl[113] vdd gnd cell_6t
Xbit_r114_c100 bl[100] br[100] wl[114] vdd gnd cell_6t
Xbit_r115_c100 bl[100] br[100] wl[115] vdd gnd cell_6t
Xbit_r116_c100 bl[100] br[100] wl[116] vdd gnd cell_6t
Xbit_r117_c100 bl[100] br[100] wl[117] vdd gnd cell_6t
Xbit_r118_c100 bl[100] br[100] wl[118] vdd gnd cell_6t
Xbit_r119_c100 bl[100] br[100] wl[119] vdd gnd cell_6t
Xbit_r120_c100 bl[100] br[100] wl[120] vdd gnd cell_6t
Xbit_r121_c100 bl[100] br[100] wl[121] vdd gnd cell_6t
Xbit_r122_c100 bl[100] br[100] wl[122] vdd gnd cell_6t
Xbit_r123_c100 bl[100] br[100] wl[123] vdd gnd cell_6t
Xbit_r124_c100 bl[100] br[100] wl[124] vdd gnd cell_6t
Xbit_r125_c100 bl[100] br[100] wl[125] vdd gnd cell_6t
Xbit_r126_c100 bl[100] br[100] wl[126] vdd gnd cell_6t
Xbit_r127_c100 bl[100] br[100] wl[127] vdd gnd cell_6t
Xbit_r128_c100 bl[100] br[100] wl[128] vdd gnd cell_6t
Xbit_r129_c100 bl[100] br[100] wl[129] vdd gnd cell_6t
Xbit_r130_c100 bl[100] br[100] wl[130] vdd gnd cell_6t
Xbit_r131_c100 bl[100] br[100] wl[131] vdd gnd cell_6t
Xbit_r132_c100 bl[100] br[100] wl[132] vdd gnd cell_6t
Xbit_r133_c100 bl[100] br[100] wl[133] vdd gnd cell_6t
Xbit_r134_c100 bl[100] br[100] wl[134] vdd gnd cell_6t
Xbit_r135_c100 bl[100] br[100] wl[135] vdd gnd cell_6t
Xbit_r136_c100 bl[100] br[100] wl[136] vdd gnd cell_6t
Xbit_r137_c100 bl[100] br[100] wl[137] vdd gnd cell_6t
Xbit_r138_c100 bl[100] br[100] wl[138] vdd gnd cell_6t
Xbit_r139_c100 bl[100] br[100] wl[139] vdd gnd cell_6t
Xbit_r140_c100 bl[100] br[100] wl[140] vdd gnd cell_6t
Xbit_r141_c100 bl[100] br[100] wl[141] vdd gnd cell_6t
Xbit_r142_c100 bl[100] br[100] wl[142] vdd gnd cell_6t
Xbit_r143_c100 bl[100] br[100] wl[143] vdd gnd cell_6t
Xbit_r144_c100 bl[100] br[100] wl[144] vdd gnd cell_6t
Xbit_r145_c100 bl[100] br[100] wl[145] vdd gnd cell_6t
Xbit_r146_c100 bl[100] br[100] wl[146] vdd gnd cell_6t
Xbit_r147_c100 bl[100] br[100] wl[147] vdd gnd cell_6t
Xbit_r148_c100 bl[100] br[100] wl[148] vdd gnd cell_6t
Xbit_r149_c100 bl[100] br[100] wl[149] vdd gnd cell_6t
Xbit_r150_c100 bl[100] br[100] wl[150] vdd gnd cell_6t
Xbit_r151_c100 bl[100] br[100] wl[151] vdd gnd cell_6t
Xbit_r152_c100 bl[100] br[100] wl[152] vdd gnd cell_6t
Xbit_r153_c100 bl[100] br[100] wl[153] vdd gnd cell_6t
Xbit_r154_c100 bl[100] br[100] wl[154] vdd gnd cell_6t
Xbit_r155_c100 bl[100] br[100] wl[155] vdd gnd cell_6t
Xbit_r156_c100 bl[100] br[100] wl[156] vdd gnd cell_6t
Xbit_r157_c100 bl[100] br[100] wl[157] vdd gnd cell_6t
Xbit_r158_c100 bl[100] br[100] wl[158] vdd gnd cell_6t
Xbit_r159_c100 bl[100] br[100] wl[159] vdd gnd cell_6t
Xbit_r160_c100 bl[100] br[100] wl[160] vdd gnd cell_6t
Xbit_r161_c100 bl[100] br[100] wl[161] vdd gnd cell_6t
Xbit_r162_c100 bl[100] br[100] wl[162] vdd gnd cell_6t
Xbit_r163_c100 bl[100] br[100] wl[163] vdd gnd cell_6t
Xbit_r164_c100 bl[100] br[100] wl[164] vdd gnd cell_6t
Xbit_r165_c100 bl[100] br[100] wl[165] vdd gnd cell_6t
Xbit_r166_c100 bl[100] br[100] wl[166] vdd gnd cell_6t
Xbit_r167_c100 bl[100] br[100] wl[167] vdd gnd cell_6t
Xbit_r168_c100 bl[100] br[100] wl[168] vdd gnd cell_6t
Xbit_r169_c100 bl[100] br[100] wl[169] vdd gnd cell_6t
Xbit_r170_c100 bl[100] br[100] wl[170] vdd gnd cell_6t
Xbit_r171_c100 bl[100] br[100] wl[171] vdd gnd cell_6t
Xbit_r172_c100 bl[100] br[100] wl[172] vdd gnd cell_6t
Xbit_r173_c100 bl[100] br[100] wl[173] vdd gnd cell_6t
Xbit_r174_c100 bl[100] br[100] wl[174] vdd gnd cell_6t
Xbit_r175_c100 bl[100] br[100] wl[175] vdd gnd cell_6t
Xbit_r176_c100 bl[100] br[100] wl[176] vdd gnd cell_6t
Xbit_r177_c100 bl[100] br[100] wl[177] vdd gnd cell_6t
Xbit_r178_c100 bl[100] br[100] wl[178] vdd gnd cell_6t
Xbit_r179_c100 bl[100] br[100] wl[179] vdd gnd cell_6t
Xbit_r180_c100 bl[100] br[100] wl[180] vdd gnd cell_6t
Xbit_r181_c100 bl[100] br[100] wl[181] vdd gnd cell_6t
Xbit_r182_c100 bl[100] br[100] wl[182] vdd gnd cell_6t
Xbit_r183_c100 bl[100] br[100] wl[183] vdd gnd cell_6t
Xbit_r184_c100 bl[100] br[100] wl[184] vdd gnd cell_6t
Xbit_r185_c100 bl[100] br[100] wl[185] vdd gnd cell_6t
Xbit_r186_c100 bl[100] br[100] wl[186] vdd gnd cell_6t
Xbit_r187_c100 bl[100] br[100] wl[187] vdd gnd cell_6t
Xbit_r188_c100 bl[100] br[100] wl[188] vdd gnd cell_6t
Xbit_r189_c100 bl[100] br[100] wl[189] vdd gnd cell_6t
Xbit_r190_c100 bl[100] br[100] wl[190] vdd gnd cell_6t
Xbit_r191_c100 bl[100] br[100] wl[191] vdd gnd cell_6t
Xbit_r192_c100 bl[100] br[100] wl[192] vdd gnd cell_6t
Xbit_r193_c100 bl[100] br[100] wl[193] vdd gnd cell_6t
Xbit_r194_c100 bl[100] br[100] wl[194] vdd gnd cell_6t
Xbit_r195_c100 bl[100] br[100] wl[195] vdd gnd cell_6t
Xbit_r196_c100 bl[100] br[100] wl[196] vdd gnd cell_6t
Xbit_r197_c100 bl[100] br[100] wl[197] vdd gnd cell_6t
Xbit_r198_c100 bl[100] br[100] wl[198] vdd gnd cell_6t
Xbit_r199_c100 bl[100] br[100] wl[199] vdd gnd cell_6t
Xbit_r200_c100 bl[100] br[100] wl[200] vdd gnd cell_6t
Xbit_r201_c100 bl[100] br[100] wl[201] vdd gnd cell_6t
Xbit_r202_c100 bl[100] br[100] wl[202] vdd gnd cell_6t
Xbit_r203_c100 bl[100] br[100] wl[203] vdd gnd cell_6t
Xbit_r204_c100 bl[100] br[100] wl[204] vdd gnd cell_6t
Xbit_r205_c100 bl[100] br[100] wl[205] vdd gnd cell_6t
Xbit_r206_c100 bl[100] br[100] wl[206] vdd gnd cell_6t
Xbit_r207_c100 bl[100] br[100] wl[207] vdd gnd cell_6t
Xbit_r208_c100 bl[100] br[100] wl[208] vdd gnd cell_6t
Xbit_r209_c100 bl[100] br[100] wl[209] vdd gnd cell_6t
Xbit_r210_c100 bl[100] br[100] wl[210] vdd gnd cell_6t
Xbit_r211_c100 bl[100] br[100] wl[211] vdd gnd cell_6t
Xbit_r212_c100 bl[100] br[100] wl[212] vdd gnd cell_6t
Xbit_r213_c100 bl[100] br[100] wl[213] vdd gnd cell_6t
Xbit_r214_c100 bl[100] br[100] wl[214] vdd gnd cell_6t
Xbit_r215_c100 bl[100] br[100] wl[215] vdd gnd cell_6t
Xbit_r216_c100 bl[100] br[100] wl[216] vdd gnd cell_6t
Xbit_r217_c100 bl[100] br[100] wl[217] vdd gnd cell_6t
Xbit_r218_c100 bl[100] br[100] wl[218] vdd gnd cell_6t
Xbit_r219_c100 bl[100] br[100] wl[219] vdd gnd cell_6t
Xbit_r220_c100 bl[100] br[100] wl[220] vdd gnd cell_6t
Xbit_r221_c100 bl[100] br[100] wl[221] vdd gnd cell_6t
Xbit_r222_c100 bl[100] br[100] wl[222] vdd gnd cell_6t
Xbit_r223_c100 bl[100] br[100] wl[223] vdd gnd cell_6t
Xbit_r224_c100 bl[100] br[100] wl[224] vdd gnd cell_6t
Xbit_r225_c100 bl[100] br[100] wl[225] vdd gnd cell_6t
Xbit_r226_c100 bl[100] br[100] wl[226] vdd gnd cell_6t
Xbit_r227_c100 bl[100] br[100] wl[227] vdd gnd cell_6t
Xbit_r228_c100 bl[100] br[100] wl[228] vdd gnd cell_6t
Xbit_r229_c100 bl[100] br[100] wl[229] vdd gnd cell_6t
Xbit_r230_c100 bl[100] br[100] wl[230] vdd gnd cell_6t
Xbit_r231_c100 bl[100] br[100] wl[231] vdd gnd cell_6t
Xbit_r232_c100 bl[100] br[100] wl[232] vdd gnd cell_6t
Xbit_r233_c100 bl[100] br[100] wl[233] vdd gnd cell_6t
Xbit_r234_c100 bl[100] br[100] wl[234] vdd gnd cell_6t
Xbit_r235_c100 bl[100] br[100] wl[235] vdd gnd cell_6t
Xbit_r236_c100 bl[100] br[100] wl[236] vdd gnd cell_6t
Xbit_r237_c100 bl[100] br[100] wl[237] vdd gnd cell_6t
Xbit_r238_c100 bl[100] br[100] wl[238] vdd gnd cell_6t
Xbit_r239_c100 bl[100] br[100] wl[239] vdd gnd cell_6t
Xbit_r240_c100 bl[100] br[100] wl[240] vdd gnd cell_6t
Xbit_r241_c100 bl[100] br[100] wl[241] vdd gnd cell_6t
Xbit_r242_c100 bl[100] br[100] wl[242] vdd gnd cell_6t
Xbit_r243_c100 bl[100] br[100] wl[243] vdd gnd cell_6t
Xbit_r244_c100 bl[100] br[100] wl[244] vdd gnd cell_6t
Xbit_r245_c100 bl[100] br[100] wl[245] vdd gnd cell_6t
Xbit_r246_c100 bl[100] br[100] wl[246] vdd gnd cell_6t
Xbit_r247_c100 bl[100] br[100] wl[247] vdd gnd cell_6t
Xbit_r248_c100 bl[100] br[100] wl[248] vdd gnd cell_6t
Xbit_r249_c100 bl[100] br[100] wl[249] vdd gnd cell_6t
Xbit_r250_c100 bl[100] br[100] wl[250] vdd gnd cell_6t
Xbit_r251_c100 bl[100] br[100] wl[251] vdd gnd cell_6t
Xbit_r252_c100 bl[100] br[100] wl[252] vdd gnd cell_6t
Xbit_r253_c100 bl[100] br[100] wl[253] vdd gnd cell_6t
Xbit_r254_c100 bl[100] br[100] wl[254] vdd gnd cell_6t
Xbit_r255_c100 bl[100] br[100] wl[255] vdd gnd cell_6t
Xbit_r256_c100 bl[100] br[100] wl[256] vdd gnd cell_6t
Xbit_r257_c100 bl[100] br[100] wl[257] vdd gnd cell_6t
Xbit_r258_c100 bl[100] br[100] wl[258] vdd gnd cell_6t
Xbit_r259_c100 bl[100] br[100] wl[259] vdd gnd cell_6t
Xbit_r260_c100 bl[100] br[100] wl[260] vdd gnd cell_6t
Xbit_r261_c100 bl[100] br[100] wl[261] vdd gnd cell_6t
Xbit_r262_c100 bl[100] br[100] wl[262] vdd gnd cell_6t
Xbit_r263_c100 bl[100] br[100] wl[263] vdd gnd cell_6t
Xbit_r264_c100 bl[100] br[100] wl[264] vdd gnd cell_6t
Xbit_r265_c100 bl[100] br[100] wl[265] vdd gnd cell_6t
Xbit_r266_c100 bl[100] br[100] wl[266] vdd gnd cell_6t
Xbit_r267_c100 bl[100] br[100] wl[267] vdd gnd cell_6t
Xbit_r268_c100 bl[100] br[100] wl[268] vdd gnd cell_6t
Xbit_r269_c100 bl[100] br[100] wl[269] vdd gnd cell_6t
Xbit_r270_c100 bl[100] br[100] wl[270] vdd gnd cell_6t
Xbit_r271_c100 bl[100] br[100] wl[271] vdd gnd cell_6t
Xbit_r272_c100 bl[100] br[100] wl[272] vdd gnd cell_6t
Xbit_r273_c100 bl[100] br[100] wl[273] vdd gnd cell_6t
Xbit_r274_c100 bl[100] br[100] wl[274] vdd gnd cell_6t
Xbit_r275_c100 bl[100] br[100] wl[275] vdd gnd cell_6t
Xbit_r276_c100 bl[100] br[100] wl[276] vdd gnd cell_6t
Xbit_r277_c100 bl[100] br[100] wl[277] vdd gnd cell_6t
Xbit_r278_c100 bl[100] br[100] wl[278] vdd gnd cell_6t
Xbit_r279_c100 bl[100] br[100] wl[279] vdd gnd cell_6t
Xbit_r280_c100 bl[100] br[100] wl[280] vdd gnd cell_6t
Xbit_r281_c100 bl[100] br[100] wl[281] vdd gnd cell_6t
Xbit_r282_c100 bl[100] br[100] wl[282] vdd gnd cell_6t
Xbit_r283_c100 bl[100] br[100] wl[283] vdd gnd cell_6t
Xbit_r284_c100 bl[100] br[100] wl[284] vdd gnd cell_6t
Xbit_r285_c100 bl[100] br[100] wl[285] vdd gnd cell_6t
Xbit_r286_c100 bl[100] br[100] wl[286] vdd gnd cell_6t
Xbit_r287_c100 bl[100] br[100] wl[287] vdd gnd cell_6t
Xbit_r288_c100 bl[100] br[100] wl[288] vdd gnd cell_6t
Xbit_r289_c100 bl[100] br[100] wl[289] vdd gnd cell_6t
Xbit_r290_c100 bl[100] br[100] wl[290] vdd gnd cell_6t
Xbit_r291_c100 bl[100] br[100] wl[291] vdd gnd cell_6t
Xbit_r292_c100 bl[100] br[100] wl[292] vdd gnd cell_6t
Xbit_r293_c100 bl[100] br[100] wl[293] vdd gnd cell_6t
Xbit_r294_c100 bl[100] br[100] wl[294] vdd gnd cell_6t
Xbit_r295_c100 bl[100] br[100] wl[295] vdd gnd cell_6t
Xbit_r296_c100 bl[100] br[100] wl[296] vdd gnd cell_6t
Xbit_r297_c100 bl[100] br[100] wl[297] vdd gnd cell_6t
Xbit_r298_c100 bl[100] br[100] wl[298] vdd gnd cell_6t
Xbit_r299_c100 bl[100] br[100] wl[299] vdd gnd cell_6t
Xbit_r300_c100 bl[100] br[100] wl[300] vdd gnd cell_6t
Xbit_r301_c100 bl[100] br[100] wl[301] vdd gnd cell_6t
Xbit_r302_c100 bl[100] br[100] wl[302] vdd gnd cell_6t
Xbit_r303_c100 bl[100] br[100] wl[303] vdd gnd cell_6t
Xbit_r304_c100 bl[100] br[100] wl[304] vdd gnd cell_6t
Xbit_r305_c100 bl[100] br[100] wl[305] vdd gnd cell_6t
Xbit_r306_c100 bl[100] br[100] wl[306] vdd gnd cell_6t
Xbit_r307_c100 bl[100] br[100] wl[307] vdd gnd cell_6t
Xbit_r308_c100 bl[100] br[100] wl[308] vdd gnd cell_6t
Xbit_r309_c100 bl[100] br[100] wl[309] vdd gnd cell_6t
Xbit_r310_c100 bl[100] br[100] wl[310] vdd gnd cell_6t
Xbit_r311_c100 bl[100] br[100] wl[311] vdd gnd cell_6t
Xbit_r312_c100 bl[100] br[100] wl[312] vdd gnd cell_6t
Xbit_r313_c100 bl[100] br[100] wl[313] vdd gnd cell_6t
Xbit_r314_c100 bl[100] br[100] wl[314] vdd gnd cell_6t
Xbit_r315_c100 bl[100] br[100] wl[315] vdd gnd cell_6t
Xbit_r316_c100 bl[100] br[100] wl[316] vdd gnd cell_6t
Xbit_r317_c100 bl[100] br[100] wl[317] vdd gnd cell_6t
Xbit_r318_c100 bl[100] br[100] wl[318] vdd gnd cell_6t
Xbit_r319_c100 bl[100] br[100] wl[319] vdd gnd cell_6t
Xbit_r320_c100 bl[100] br[100] wl[320] vdd gnd cell_6t
Xbit_r321_c100 bl[100] br[100] wl[321] vdd gnd cell_6t
Xbit_r322_c100 bl[100] br[100] wl[322] vdd gnd cell_6t
Xbit_r323_c100 bl[100] br[100] wl[323] vdd gnd cell_6t
Xbit_r324_c100 bl[100] br[100] wl[324] vdd gnd cell_6t
Xbit_r325_c100 bl[100] br[100] wl[325] vdd gnd cell_6t
Xbit_r326_c100 bl[100] br[100] wl[326] vdd gnd cell_6t
Xbit_r327_c100 bl[100] br[100] wl[327] vdd gnd cell_6t
Xbit_r328_c100 bl[100] br[100] wl[328] vdd gnd cell_6t
Xbit_r329_c100 bl[100] br[100] wl[329] vdd gnd cell_6t
Xbit_r330_c100 bl[100] br[100] wl[330] vdd gnd cell_6t
Xbit_r331_c100 bl[100] br[100] wl[331] vdd gnd cell_6t
Xbit_r332_c100 bl[100] br[100] wl[332] vdd gnd cell_6t
Xbit_r333_c100 bl[100] br[100] wl[333] vdd gnd cell_6t
Xbit_r334_c100 bl[100] br[100] wl[334] vdd gnd cell_6t
Xbit_r335_c100 bl[100] br[100] wl[335] vdd gnd cell_6t
Xbit_r336_c100 bl[100] br[100] wl[336] vdd gnd cell_6t
Xbit_r337_c100 bl[100] br[100] wl[337] vdd gnd cell_6t
Xbit_r338_c100 bl[100] br[100] wl[338] vdd gnd cell_6t
Xbit_r339_c100 bl[100] br[100] wl[339] vdd gnd cell_6t
Xbit_r340_c100 bl[100] br[100] wl[340] vdd gnd cell_6t
Xbit_r341_c100 bl[100] br[100] wl[341] vdd gnd cell_6t
Xbit_r342_c100 bl[100] br[100] wl[342] vdd gnd cell_6t
Xbit_r343_c100 bl[100] br[100] wl[343] vdd gnd cell_6t
Xbit_r344_c100 bl[100] br[100] wl[344] vdd gnd cell_6t
Xbit_r345_c100 bl[100] br[100] wl[345] vdd gnd cell_6t
Xbit_r346_c100 bl[100] br[100] wl[346] vdd gnd cell_6t
Xbit_r347_c100 bl[100] br[100] wl[347] vdd gnd cell_6t
Xbit_r348_c100 bl[100] br[100] wl[348] vdd gnd cell_6t
Xbit_r349_c100 bl[100] br[100] wl[349] vdd gnd cell_6t
Xbit_r350_c100 bl[100] br[100] wl[350] vdd gnd cell_6t
Xbit_r351_c100 bl[100] br[100] wl[351] vdd gnd cell_6t
Xbit_r352_c100 bl[100] br[100] wl[352] vdd gnd cell_6t
Xbit_r353_c100 bl[100] br[100] wl[353] vdd gnd cell_6t
Xbit_r354_c100 bl[100] br[100] wl[354] vdd gnd cell_6t
Xbit_r355_c100 bl[100] br[100] wl[355] vdd gnd cell_6t
Xbit_r356_c100 bl[100] br[100] wl[356] vdd gnd cell_6t
Xbit_r357_c100 bl[100] br[100] wl[357] vdd gnd cell_6t
Xbit_r358_c100 bl[100] br[100] wl[358] vdd gnd cell_6t
Xbit_r359_c100 bl[100] br[100] wl[359] vdd gnd cell_6t
Xbit_r360_c100 bl[100] br[100] wl[360] vdd gnd cell_6t
Xbit_r361_c100 bl[100] br[100] wl[361] vdd gnd cell_6t
Xbit_r362_c100 bl[100] br[100] wl[362] vdd gnd cell_6t
Xbit_r363_c100 bl[100] br[100] wl[363] vdd gnd cell_6t
Xbit_r364_c100 bl[100] br[100] wl[364] vdd gnd cell_6t
Xbit_r365_c100 bl[100] br[100] wl[365] vdd gnd cell_6t
Xbit_r366_c100 bl[100] br[100] wl[366] vdd gnd cell_6t
Xbit_r367_c100 bl[100] br[100] wl[367] vdd gnd cell_6t
Xbit_r368_c100 bl[100] br[100] wl[368] vdd gnd cell_6t
Xbit_r369_c100 bl[100] br[100] wl[369] vdd gnd cell_6t
Xbit_r370_c100 bl[100] br[100] wl[370] vdd gnd cell_6t
Xbit_r371_c100 bl[100] br[100] wl[371] vdd gnd cell_6t
Xbit_r372_c100 bl[100] br[100] wl[372] vdd gnd cell_6t
Xbit_r373_c100 bl[100] br[100] wl[373] vdd gnd cell_6t
Xbit_r374_c100 bl[100] br[100] wl[374] vdd gnd cell_6t
Xbit_r375_c100 bl[100] br[100] wl[375] vdd gnd cell_6t
Xbit_r376_c100 bl[100] br[100] wl[376] vdd gnd cell_6t
Xbit_r377_c100 bl[100] br[100] wl[377] vdd gnd cell_6t
Xbit_r378_c100 bl[100] br[100] wl[378] vdd gnd cell_6t
Xbit_r379_c100 bl[100] br[100] wl[379] vdd gnd cell_6t
Xbit_r380_c100 bl[100] br[100] wl[380] vdd gnd cell_6t
Xbit_r381_c100 bl[100] br[100] wl[381] vdd gnd cell_6t
Xbit_r382_c100 bl[100] br[100] wl[382] vdd gnd cell_6t
Xbit_r383_c100 bl[100] br[100] wl[383] vdd gnd cell_6t
Xbit_r384_c100 bl[100] br[100] wl[384] vdd gnd cell_6t
Xbit_r385_c100 bl[100] br[100] wl[385] vdd gnd cell_6t
Xbit_r386_c100 bl[100] br[100] wl[386] vdd gnd cell_6t
Xbit_r387_c100 bl[100] br[100] wl[387] vdd gnd cell_6t
Xbit_r388_c100 bl[100] br[100] wl[388] vdd gnd cell_6t
Xbit_r389_c100 bl[100] br[100] wl[389] vdd gnd cell_6t
Xbit_r390_c100 bl[100] br[100] wl[390] vdd gnd cell_6t
Xbit_r391_c100 bl[100] br[100] wl[391] vdd gnd cell_6t
Xbit_r392_c100 bl[100] br[100] wl[392] vdd gnd cell_6t
Xbit_r393_c100 bl[100] br[100] wl[393] vdd gnd cell_6t
Xbit_r394_c100 bl[100] br[100] wl[394] vdd gnd cell_6t
Xbit_r395_c100 bl[100] br[100] wl[395] vdd gnd cell_6t
Xbit_r396_c100 bl[100] br[100] wl[396] vdd gnd cell_6t
Xbit_r397_c100 bl[100] br[100] wl[397] vdd gnd cell_6t
Xbit_r398_c100 bl[100] br[100] wl[398] vdd gnd cell_6t
Xbit_r399_c100 bl[100] br[100] wl[399] vdd gnd cell_6t
Xbit_r400_c100 bl[100] br[100] wl[400] vdd gnd cell_6t
Xbit_r401_c100 bl[100] br[100] wl[401] vdd gnd cell_6t
Xbit_r402_c100 bl[100] br[100] wl[402] vdd gnd cell_6t
Xbit_r403_c100 bl[100] br[100] wl[403] vdd gnd cell_6t
Xbit_r404_c100 bl[100] br[100] wl[404] vdd gnd cell_6t
Xbit_r405_c100 bl[100] br[100] wl[405] vdd gnd cell_6t
Xbit_r406_c100 bl[100] br[100] wl[406] vdd gnd cell_6t
Xbit_r407_c100 bl[100] br[100] wl[407] vdd gnd cell_6t
Xbit_r408_c100 bl[100] br[100] wl[408] vdd gnd cell_6t
Xbit_r409_c100 bl[100] br[100] wl[409] vdd gnd cell_6t
Xbit_r410_c100 bl[100] br[100] wl[410] vdd gnd cell_6t
Xbit_r411_c100 bl[100] br[100] wl[411] vdd gnd cell_6t
Xbit_r412_c100 bl[100] br[100] wl[412] vdd gnd cell_6t
Xbit_r413_c100 bl[100] br[100] wl[413] vdd gnd cell_6t
Xbit_r414_c100 bl[100] br[100] wl[414] vdd gnd cell_6t
Xbit_r415_c100 bl[100] br[100] wl[415] vdd gnd cell_6t
Xbit_r416_c100 bl[100] br[100] wl[416] vdd gnd cell_6t
Xbit_r417_c100 bl[100] br[100] wl[417] vdd gnd cell_6t
Xbit_r418_c100 bl[100] br[100] wl[418] vdd gnd cell_6t
Xbit_r419_c100 bl[100] br[100] wl[419] vdd gnd cell_6t
Xbit_r420_c100 bl[100] br[100] wl[420] vdd gnd cell_6t
Xbit_r421_c100 bl[100] br[100] wl[421] vdd gnd cell_6t
Xbit_r422_c100 bl[100] br[100] wl[422] vdd gnd cell_6t
Xbit_r423_c100 bl[100] br[100] wl[423] vdd gnd cell_6t
Xbit_r424_c100 bl[100] br[100] wl[424] vdd gnd cell_6t
Xbit_r425_c100 bl[100] br[100] wl[425] vdd gnd cell_6t
Xbit_r426_c100 bl[100] br[100] wl[426] vdd gnd cell_6t
Xbit_r427_c100 bl[100] br[100] wl[427] vdd gnd cell_6t
Xbit_r428_c100 bl[100] br[100] wl[428] vdd gnd cell_6t
Xbit_r429_c100 bl[100] br[100] wl[429] vdd gnd cell_6t
Xbit_r430_c100 bl[100] br[100] wl[430] vdd gnd cell_6t
Xbit_r431_c100 bl[100] br[100] wl[431] vdd gnd cell_6t
Xbit_r432_c100 bl[100] br[100] wl[432] vdd gnd cell_6t
Xbit_r433_c100 bl[100] br[100] wl[433] vdd gnd cell_6t
Xbit_r434_c100 bl[100] br[100] wl[434] vdd gnd cell_6t
Xbit_r435_c100 bl[100] br[100] wl[435] vdd gnd cell_6t
Xbit_r436_c100 bl[100] br[100] wl[436] vdd gnd cell_6t
Xbit_r437_c100 bl[100] br[100] wl[437] vdd gnd cell_6t
Xbit_r438_c100 bl[100] br[100] wl[438] vdd gnd cell_6t
Xbit_r439_c100 bl[100] br[100] wl[439] vdd gnd cell_6t
Xbit_r440_c100 bl[100] br[100] wl[440] vdd gnd cell_6t
Xbit_r441_c100 bl[100] br[100] wl[441] vdd gnd cell_6t
Xbit_r442_c100 bl[100] br[100] wl[442] vdd gnd cell_6t
Xbit_r443_c100 bl[100] br[100] wl[443] vdd gnd cell_6t
Xbit_r444_c100 bl[100] br[100] wl[444] vdd gnd cell_6t
Xbit_r445_c100 bl[100] br[100] wl[445] vdd gnd cell_6t
Xbit_r446_c100 bl[100] br[100] wl[446] vdd gnd cell_6t
Xbit_r447_c100 bl[100] br[100] wl[447] vdd gnd cell_6t
Xbit_r448_c100 bl[100] br[100] wl[448] vdd gnd cell_6t
Xbit_r449_c100 bl[100] br[100] wl[449] vdd gnd cell_6t
Xbit_r450_c100 bl[100] br[100] wl[450] vdd gnd cell_6t
Xbit_r451_c100 bl[100] br[100] wl[451] vdd gnd cell_6t
Xbit_r452_c100 bl[100] br[100] wl[452] vdd gnd cell_6t
Xbit_r453_c100 bl[100] br[100] wl[453] vdd gnd cell_6t
Xbit_r454_c100 bl[100] br[100] wl[454] vdd gnd cell_6t
Xbit_r455_c100 bl[100] br[100] wl[455] vdd gnd cell_6t
Xbit_r456_c100 bl[100] br[100] wl[456] vdd gnd cell_6t
Xbit_r457_c100 bl[100] br[100] wl[457] vdd gnd cell_6t
Xbit_r458_c100 bl[100] br[100] wl[458] vdd gnd cell_6t
Xbit_r459_c100 bl[100] br[100] wl[459] vdd gnd cell_6t
Xbit_r460_c100 bl[100] br[100] wl[460] vdd gnd cell_6t
Xbit_r461_c100 bl[100] br[100] wl[461] vdd gnd cell_6t
Xbit_r462_c100 bl[100] br[100] wl[462] vdd gnd cell_6t
Xbit_r463_c100 bl[100] br[100] wl[463] vdd gnd cell_6t
Xbit_r464_c100 bl[100] br[100] wl[464] vdd gnd cell_6t
Xbit_r465_c100 bl[100] br[100] wl[465] vdd gnd cell_6t
Xbit_r466_c100 bl[100] br[100] wl[466] vdd gnd cell_6t
Xbit_r467_c100 bl[100] br[100] wl[467] vdd gnd cell_6t
Xbit_r468_c100 bl[100] br[100] wl[468] vdd gnd cell_6t
Xbit_r469_c100 bl[100] br[100] wl[469] vdd gnd cell_6t
Xbit_r470_c100 bl[100] br[100] wl[470] vdd gnd cell_6t
Xbit_r471_c100 bl[100] br[100] wl[471] vdd gnd cell_6t
Xbit_r472_c100 bl[100] br[100] wl[472] vdd gnd cell_6t
Xbit_r473_c100 bl[100] br[100] wl[473] vdd gnd cell_6t
Xbit_r474_c100 bl[100] br[100] wl[474] vdd gnd cell_6t
Xbit_r475_c100 bl[100] br[100] wl[475] vdd gnd cell_6t
Xbit_r476_c100 bl[100] br[100] wl[476] vdd gnd cell_6t
Xbit_r477_c100 bl[100] br[100] wl[477] vdd gnd cell_6t
Xbit_r478_c100 bl[100] br[100] wl[478] vdd gnd cell_6t
Xbit_r479_c100 bl[100] br[100] wl[479] vdd gnd cell_6t
Xbit_r480_c100 bl[100] br[100] wl[480] vdd gnd cell_6t
Xbit_r481_c100 bl[100] br[100] wl[481] vdd gnd cell_6t
Xbit_r482_c100 bl[100] br[100] wl[482] vdd gnd cell_6t
Xbit_r483_c100 bl[100] br[100] wl[483] vdd gnd cell_6t
Xbit_r484_c100 bl[100] br[100] wl[484] vdd gnd cell_6t
Xbit_r485_c100 bl[100] br[100] wl[485] vdd gnd cell_6t
Xbit_r486_c100 bl[100] br[100] wl[486] vdd gnd cell_6t
Xbit_r487_c100 bl[100] br[100] wl[487] vdd gnd cell_6t
Xbit_r488_c100 bl[100] br[100] wl[488] vdd gnd cell_6t
Xbit_r489_c100 bl[100] br[100] wl[489] vdd gnd cell_6t
Xbit_r490_c100 bl[100] br[100] wl[490] vdd gnd cell_6t
Xbit_r491_c100 bl[100] br[100] wl[491] vdd gnd cell_6t
Xbit_r492_c100 bl[100] br[100] wl[492] vdd gnd cell_6t
Xbit_r493_c100 bl[100] br[100] wl[493] vdd gnd cell_6t
Xbit_r494_c100 bl[100] br[100] wl[494] vdd gnd cell_6t
Xbit_r495_c100 bl[100] br[100] wl[495] vdd gnd cell_6t
Xbit_r496_c100 bl[100] br[100] wl[496] vdd gnd cell_6t
Xbit_r497_c100 bl[100] br[100] wl[497] vdd gnd cell_6t
Xbit_r498_c100 bl[100] br[100] wl[498] vdd gnd cell_6t
Xbit_r499_c100 bl[100] br[100] wl[499] vdd gnd cell_6t
Xbit_r500_c100 bl[100] br[100] wl[500] vdd gnd cell_6t
Xbit_r501_c100 bl[100] br[100] wl[501] vdd gnd cell_6t
Xbit_r502_c100 bl[100] br[100] wl[502] vdd gnd cell_6t
Xbit_r503_c100 bl[100] br[100] wl[503] vdd gnd cell_6t
Xbit_r504_c100 bl[100] br[100] wl[504] vdd gnd cell_6t
Xbit_r505_c100 bl[100] br[100] wl[505] vdd gnd cell_6t
Xbit_r506_c100 bl[100] br[100] wl[506] vdd gnd cell_6t
Xbit_r507_c100 bl[100] br[100] wl[507] vdd gnd cell_6t
Xbit_r508_c100 bl[100] br[100] wl[508] vdd gnd cell_6t
Xbit_r509_c100 bl[100] br[100] wl[509] vdd gnd cell_6t
Xbit_r510_c100 bl[100] br[100] wl[510] vdd gnd cell_6t
Xbit_r511_c100 bl[100] br[100] wl[511] vdd gnd cell_6t
Xbit_r0_c101 bl[101] br[101] wl[0] vdd gnd cell_6t
Xbit_r1_c101 bl[101] br[101] wl[1] vdd gnd cell_6t
Xbit_r2_c101 bl[101] br[101] wl[2] vdd gnd cell_6t
Xbit_r3_c101 bl[101] br[101] wl[3] vdd gnd cell_6t
Xbit_r4_c101 bl[101] br[101] wl[4] vdd gnd cell_6t
Xbit_r5_c101 bl[101] br[101] wl[5] vdd gnd cell_6t
Xbit_r6_c101 bl[101] br[101] wl[6] vdd gnd cell_6t
Xbit_r7_c101 bl[101] br[101] wl[7] vdd gnd cell_6t
Xbit_r8_c101 bl[101] br[101] wl[8] vdd gnd cell_6t
Xbit_r9_c101 bl[101] br[101] wl[9] vdd gnd cell_6t
Xbit_r10_c101 bl[101] br[101] wl[10] vdd gnd cell_6t
Xbit_r11_c101 bl[101] br[101] wl[11] vdd gnd cell_6t
Xbit_r12_c101 bl[101] br[101] wl[12] vdd gnd cell_6t
Xbit_r13_c101 bl[101] br[101] wl[13] vdd gnd cell_6t
Xbit_r14_c101 bl[101] br[101] wl[14] vdd gnd cell_6t
Xbit_r15_c101 bl[101] br[101] wl[15] vdd gnd cell_6t
Xbit_r16_c101 bl[101] br[101] wl[16] vdd gnd cell_6t
Xbit_r17_c101 bl[101] br[101] wl[17] vdd gnd cell_6t
Xbit_r18_c101 bl[101] br[101] wl[18] vdd gnd cell_6t
Xbit_r19_c101 bl[101] br[101] wl[19] vdd gnd cell_6t
Xbit_r20_c101 bl[101] br[101] wl[20] vdd gnd cell_6t
Xbit_r21_c101 bl[101] br[101] wl[21] vdd gnd cell_6t
Xbit_r22_c101 bl[101] br[101] wl[22] vdd gnd cell_6t
Xbit_r23_c101 bl[101] br[101] wl[23] vdd gnd cell_6t
Xbit_r24_c101 bl[101] br[101] wl[24] vdd gnd cell_6t
Xbit_r25_c101 bl[101] br[101] wl[25] vdd gnd cell_6t
Xbit_r26_c101 bl[101] br[101] wl[26] vdd gnd cell_6t
Xbit_r27_c101 bl[101] br[101] wl[27] vdd gnd cell_6t
Xbit_r28_c101 bl[101] br[101] wl[28] vdd gnd cell_6t
Xbit_r29_c101 bl[101] br[101] wl[29] vdd gnd cell_6t
Xbit_r30_c101 bl[101] br[101] wl[30] vdd gnd cell_6t
Xbit_r31_c101 bl[101] br[101] wl[31] vdd gnd cell_6t
Xbit_r32_c101 bl[101] br[101] wl[32] vdd gnd cell_6t
Xbit_r33_c101 bl[101] br[101] wl[33] vdd gnd cell_6t
Xbit_r34_c101 bl[101] br[101] wl[34] vdd gnd cell_6t
Xbit_r35_c101 bl[101] br[101] wl[35] vdd gnd cell_6t
Xbit_r36_c101 bl[101] br[101] wl[36] vdd gnd cell_6t
Xbit_r37_c101 bl[101] br[101] wl[37] vdd gnd cell_6t
Xbit_r38_c101 bl[101] br[101] wl[38] vdd gnd cell_6t
Xbit_r39_c101 bl[101] br[101] wl[39] vdd gnd cell_6t
Xbit_r40_c101 bl[101] br[101] wl[40] vdd gnd cell_6t
Xbit_r41_c101 bl[101] br[101] wl[41] vdd gnd cell_6t
Xbit_r42_c101 bl[101] br[101] wl[42] vdd gnd cell_6t
Xbit_r43_c101 bl[101] br[101] wl[43] vdd gnd cell_6t
Xbit_r44_c101 bl[101] br[101] wl[44] vdd gnd cell_6t
Xbit_r45_c101 bl[101] br[101] wl[45] vdd gnd cell_6t
Xbit_r46_c101 bl[101] br[101] wl[46] vdd gnd cell_6t
Xbit_r47_c101 bl[101] br[101] wl[47] vdd gnd cell_6t
Xbit_r48_c101 bl[101] br[101] wl[48] vdd gnd cell_6t
Xbit_r49_c101 bl[101] br[101] wl[49] vdd gnd cell_6t
Xbit_r50_c101 bl[101] br[101] wl[50] vdd gnd cell_6t
Xbit_r51_c101 bl[101] br[101] wl[51] vdd gnd cell_6t
Xbit_r52_c101 bl[101] br[101] wl[52] vdd gnd cell_6t
Xbit_r53_c101 bl[101] br[101] wl[53] vdd gnd cell_6t
Xbit_r54_c101 bl[101] br[101] wl[54] vdd gnd cell_6t
Xbit_r55_c101 bl[101] br[101] wl[55] vdd gnd cell_6t
Xbit_r56_c101 bl[101] br[101] wl[56] vdd gnd cell_6t
Xbit_r57_c101 bl[101] br[101] wl[57] vdd gnd cell_6t
Xbit_r58_c101 bl[101] br[101] wl[58] vdd gnd cell_6t
Xbit_r59_c101 bl[101] br[101] wl[59] vdd gnd cell_6t
Xbit_r60_c101 bl[101] br[101] wl[60] vdd gnd cell_6t
Xbit_r61_c101 bl[101] br[101] wl[61] vdd gnd cell_6t
Xbit_r62_c101 bl[101] br[101] wl[62] vdd gnd cell_6t
Xbit_r63_c101 bl[101] br[101] wl[63] vdd gnd cell_6t
Xbit_r64_c101 bl[101] br[101] wl[64] vdd gnd cell_6t
Xbit_r65_c101 bl[101] br[101] wl[65] vdd gnd cell_6t
Xbit_r66_c101 bl[101] br[101] wl[66] vdd gnd cell_6t
Xbit_r67_c101 bl[101] br[101] wl[67] vdd gnd cell_6t
Xbit_r68_c101 bl[101] br[101] wl[68] vdd gnd cell_6t
Xbit_r69_c101 bl[101] br[101] wl[69] vdd gnd cell_6t
Xbit_r70_c101 bl[101] br[101] wl[70] vdd gnd cell_6t
Xbit_r71_c101 bl[101] br[101] wl[71] vdd gnd cell_6t
Xbit_r72_c101 bl[101] br[101] wl[72] vdd gnd cell_6t
Xbit_r73_c101 bl[101] br[101] wl[73] vdd gnd cell_6t
Xbit_r74_c101 bl[101] br[101] wl[74] vdd gnd cell_6t
Xbit_r75_c101 bl[101] br[101] wl[75] vdd gnd cell_6t
Xbit_r76_c101 bl[101] br[101] wl[76] vdd gnd cell_6t
Xbit_r77_c101 bl[101] br[101] wl[77] vdd gnd cell_6t
Xbit_r78_c101 bl[101] br[101] wl[78] vdd gnd cell_6t
Xbit_r79_c101 bl[101] br[101] wl[79] vdd gnd cell_6t
Xbit_r80_c101 bl[101] br[101] wl[80] vdd gnd cell_6t
Xbit_r81_c101 bl[101] br[101] wl[81] vdd gnd cell_6t
Xbit_r82_c101 bl[101] br[101] wl[82] vdd gnd cell_6t
Xbit_r83_c101 bl[101] br[101] wl[83] vdd gnd cell_6t
Xbit_r84_c101 bl[101] br[101] wl[84] vdd gnd cell_6t
Xbit_r85_c101 bl[101] br[101] wl[85] vdd gnd cell_6t
Xbit_r86_c101 bl[101] br[101] wl[86] vdd gnd cell_6t
Xbit_r87_c101 bl[101] br[101] wl[87] vdd gnd cell_6t
Xbit_r88_c101 bl[101] br[101] wl[88] vdd gnd cell_6t
Xbit_r89_c101 bl[101] br[101] wl[89] vdd gnd cell_6t
Xbit_r90_c101 bl[101] br[101] wl[90] vdd gnd cell_6t
Xbit_r91_c101 bl[101] br[101] wl[91] vdd gnd cell_6t
Xbit_r92_c101 bl[101] br[101] wl[92] vdd gnd cell_6t
Xbit_r93_c101 bl[101] br[101] wl[93] vdd gnd cell_6t
Xbit_r94_c101 bl[101] br[101] wl[94] vdd gnd cell_6t
Xbit_r95_c101 bl[101] br[101] wl[95] vdd gnd cell_6t
Xbit_r96_c101 bl[101] br[101] wl[96] vdd gnd cell_6t
Xbit_r97_c101 bl[101] br[101] wl[97] vdd gnd cell_6t
Xbit_r98_c101 bl[101] br[101] wl[98] vdd gnd cell_6t
Xbit_r99_c101 bl[101] br[101] wl[99] vdd gnd cell_6t
Xbit_r100_c101 bl[101] br[101] wl[100] vdd gnd cell_6t
Xbit_r101_c101 bl[101] br[101] wl[101] vdd gnd cell_6t
Xbit_r102_c101 bl[101] br[101] wl[102] vdd gnd cell_6t
Xbit_r103_c101 bl[101] br[101] wl[103] vdd gnd cell_6t
Xbit_r104_c101 bl[101] br[101] wl[104] vdd gnd cell_6t
Xbit_r105_c101 bl[101] br[101] wl[105] vdd gnd cell_6t
Xbit_r106_c101 bl[101] br[101] wl[106] vdd gnd cell_6t
Xbit_r107_c101 bl[101] br[101] wl[107] vdd gnd cell_6t
Xbit_r108_c101 bl[101] br[101] wl[108] vdd gnd cell_6t
Xbit_r109_c101 bl[101] br[101] wl[109] vdd gnd cell_6t
Xbit_r110_c101 bl[101] br[101] wl[110] vdd gnd cell_6t
Xbit_r111_c101 bl[101] br[101] wl[111] vdd gnd cell_6t
Xbit_r112_c101 bl[101] br[101] wl[112] vdd gnd cell_6t
Xbit_r113_c101 bl[101] br[101] wl[113] vdd gnd cell_6t
Xbit_r114_c101 bl[101] br[101] wl[114] vdd gnd cell_6t
Xbit_r115_c101 bl[101] br[101] wl[115] vdd gnd cell_6t
Xbit_r116_c101 bl[101] br[101] wl[116] vdd gnd cell_6t
Xbit_r117_c101 bl[101] br[101] wl[117] vdd gnd cell_6t
Xbit_r118_c101 bl[101] br[101] wl[118] vdd gnd cell_6t
Xbit_r119_c101 bl[101] br[101] wl[119] vdd gnd cell_6t
Xbit_r120_c101 bl[101] br[101] wl[120] vdd gnd cell_6t
Xbit_r121_c101 bl[101] br[101] wl[121] vdd gnd cell_6t
Xbit_r122_c101 bl[101] br[101] wl[122] vdd gnd cell_6t
Xbit_r123_c101 bl[101] br[101] wl[123] vdd gnd cell_6t
Xbit_r124_c101 bl[101] br[101] wl[124] vdd gnd cell_6t
Xbit_r125_c101 bl[101] br[101] wl[125] vdd gnd cell_6t
Xbit_r126_c101 bl[101] br[101] wl[126] vdd gnd cell_6t
Xbit_r127_c101 bl[101] br[101] wl[127] vdd gnd cell_6t
Xbit_r128_c101 bl[101] br[101] wl[128] vdd gnd cell_6t
Xbit_r129_c101 bl[101] br[101] wl[129] vdd gnd cell_6t
Xbit_r130_c101 bl[101] br[101] wl[130] vdd gnd cell_6t
Xbit_r131_c101 bl[101] br[101] wl[131] vdd gnd cell_6t
Xbit_r132_c101 bl[101] br[101] wl[132] vdd gnd cell_6t
Xbit_r133_c101 bl[101] br[101] wl[133] vdd gnd cell_6t
Xbit_r134_c101 bl[101] br[101] wl[134] vdd gnd cell_6t
Xbit_r135_c101 bl[101] br[101] wl[135] vdd gnd cell_6t
Xbit_r136_c101 bl[101] br[101] wl[136] vdd gnd cell_6t
Xbit_r137_c101 bl[101] br[101] wl[137] vdd gnd cell_6t
Xbit_r138_c101 bl[101] br[101] wl[138] vdd gnd cell_6t
Xbit_r139_c101 bl[101] br[101] wl[139] vdd gnd cell_6t
Xbit_r140_c101 bl[101] br[101] wl[140] vdd gnd cell_6t
Xbit_r141_c101 bl[101] br[101] wl[141] vdd gnd cell_6t
Xbit_r142_c101 bl[101] br[101] wl[142] vdd gnd cell_6t
Xbit_r143_c101 bl[101] br[101] wl[143] vdd gnd cell_6t
Xbit_r144_c101 bl[101] br[101] wl[144] vdd gnd cell_6t
Xbit_r145_c101 bl[101] br[101] wl[145] vdd gnd cell_6t
Xbit_r146_c101 bl[101] br[101] wl[146] vdd gnd cell_6t
Xbit_r147_c101 bl[101] br[101] wl[147] vdd gnd cell_6t
Xbit_r148_c101 bl[101] br[101] wl[148] vdd gnd cell_6t
Xbit_r149_c101 bl[101] br[101] wl[149] vdd gnd cell_6t
Xbit_r150_c101 bl[101] br[101] wl[150] vdd gnd cell_6t
Xbit_r151_c101 bl[101] br[101] wl[151] vdd gnd cell_6t
Xbit_r152_c101 bl[101] br[101] wl[152] vdd gnd cell_6t
Xbit_r153_c101 bl[101] br[101] wl[153] vdd gnd cell_6t
Xbit_r154_c101 bl[101] br[101] wl[154] vdd gnd cell_6t
Xbit_r155_c101 bl[101] br[101] wl[155] vdd gnd cell_6t
Xbit_r156_c101 bl[101] br[101] wl[156] vdd gnd cell_6t
Xbit_r157_c101 bl[101] br[101] wl[157] vdd gnd cell_6t
Xbit_r158_c101 bl[101] br[101] wl[158] vdd gnd cell_6t
Xbit_r159_c101 bl[101] br[101] wl[159] vdd gnd cell_6t
Xbit_r160_c101 bl[101] br[101] wl[160] vdd gnd cell_6t
Xbit_r161_c101 bl[101] br[101] wl[161] vdd gnd cell_6t
Xbit_r162_c101 bl[101] br[101] wl[162] vdd gnd cell_6t
Xbit_r163_c101 bl[101] br[101] wl[163] vdd gnd cell_6t
Xbit_r164_c101 bl[101] br[101] wl[164] vdd gnd cell_6t
Xbit_r165_c101 bl[101] br[101] wl[165] vdd gnd cell_6t
Xbit_r166_c101 bl[101] br[101] wl[166] vdd gnd cell_6t
Xbit_r167_c101 bl[101] br[101] wl[167] vdd gnd cell_6t
Xbit_r168_c101 bl[101] br[101] wl[168] vdd gnd cell_6t
Xbit_r169_c101 bl[101] br[101] wl[169] vdd gnd cell_6t
Xbit_r170_c101 bl[101] br[101] wl[170] vdd gnd cell_6t
Xbit_r171_c101 bl[101] br[101] wl[171] vdd gnd cell_6t
Xbit_r172_c101 bl[101] br[101] wl[172] vdd gnd cell_6t
Xbit_r173_c101 bl[101] br[101] wl[173] vdd gnd cell_6t
Xbit_r174_c101 bl[101] br[101] wl[174] vdd gnd cell_6t
Xbit_r175_c101 bl[101] br[101] wl[175] vdd gnd cell_6t
Xbit_r176_c101 bl[101] br[101] wl[176] vdd gnd cell_6t
Xbit_r177_c101 bl[101] br[101] wl[177] vdd gnd cell_6t
Xbit_r178_c101 bl[101] br[101] wl[178] vdd gnd cell_6t
Xbit_r179_c101 bl[101] br[101] wl[179] vdd gnd cell_6t
Xbit_r180_c101 bl[101] br[101] wl[180] vdd gnd cell_6t
Xbit_r181_c101 bl[101] br[101] wl[181] vdd gnd cell_6t
Xbit_r182_c101 bl[101] br[101] wl[182] vdd gnd cell_6t
Xbit_r183_c101 bl[101] br[101] wl[183] vdd gnd cell_6t
Xbit_r184_c101 bl[101] br[101] wl[184] vdd gnd cell_6t
Xbit_r185_c101 bl[101] br[101] wl[185] vdd gnd cell_6t
Xbit_r186_c101 bl[101] br[101] wl[186] vdd gnd cell_6t
Xbit_r187_c101 bl[101] br[101] wl[187] vdd gnd cell_6t
Xbit_r188_c101 bl[101] br[101] wl[188] vdd gnd cell_6t
Xbit_r189_c101 bl[101] br[101] wl[189] vdd gnd cell_6t
Xbit_r190_c101 bl[101] br[101] wl[190] vdd gnd cell_6t
Xbit_r191_c101 bl[101] br[101] wl[191] vdd gnd cell_6t
Xbit_r192_c101 bl[101] br[101] wl[192] vdd gnd cell_6t
Xbit_r193_c101 bl[101] br[101] wl[193] vdd gnd cell_6t
Xbit_r194_c101 bl[101] br[101] wl[194] vdd gnd cell_6t
Xbit_r195_c101 bl[101] br[101] wl[195] vdd gnd cell_6t
Xbit_r196_c101 bl[101] br[101] wl[196] vdd gnd cell_6t
Xbit_r197_c101 bl[101] br[101] wl[197] vdd gnd cell_6t
Xbit_r198_c101 bl[101] br[101] wl[198] vdd gnd cell_6t
Xbit_r199_c101 bl[101] br[101] wl[199] vdd gnd cell_6t
Xbit_r200_c101 bl[101] br[101] wl[200] vdd gnd cell_6t
Xbit_r201_c101 bl[101] br[101] wl[201] vdd gnd cell_6t
Xbit_r202_c101 bl[101] br[101] wl[202] vdd gnd cell_6t
Xbit_r203_c101 bl[101] br[101] wl[203] vdd gnd cell_6t
Xbit_r204_c101 bl[101] br[101] wl[204] vdd gnd cell_6t
Xbit_r205_c101 bl[101] br[101] wl[205] vdd gnd cell_6t
Xbit_r206_c101 bl[101] br[101] wl[206] vdd gnd cell_6t
Xbit_r207_c101 bl[101] br[101] wl[207] vdd gnd cell_6t
Xbit_r208_c101 bl[101] br[101] wl[208] vdd gnd cell_6t
Xbit_r209_c101 bl[101] br[101] wl[209] vdd gnd cell_6t
Xbit_r210_c101 bl[101] br[101] wl[210] vdd gnd cell_6t
Xbit_r211_c101 bl[101] br[101] wl[211] vdd gnd cell_6t
Xbit_r212_c101 bl[101] br[101] wl[212] vdd gnd cell_6t
Xbit_r213_c101 bl[101] br[101] wl[213] vdd gnd cell_6t
Xbit_r214_c101 bl[101] br[101] wl[214] vdd gnd cell_6t
Xbit_r215_c101 bl[101] br[101] wl[215] vdd gnd cell_6t
Xbit_r216_c101 bl[101] br[101] wl[216] vdd gnd cell_6t
Xbit_r217_c101 bl[101] br[101] wl[217] vdd gnd cell_6t
Xbit_r218_c101 bl[101] br[101] wl[218] vdd gnd cell_6t
Xbit_r219_c101 bl[101] br[101] wl[219] vdd gnd cell_6t
Xbit_r220_c101 bl[101] br[101] wl[220] vdd gnd cell_6t
Xbit_r221_c101 bl[101] br[101] wl[221] vdd gnd cell_6t
Xbit_r222_c101 bl[101] br[101] wl[222] vdd gnd cell_6t
Xbit_r223_c101 bl[101] br[101] wl[223] vdd gnd cell_6t
Xbit_r224_c101 bl[101] br[101] wl[224] vdd gnd cell_6t
Xbit_r225_c101 bl[101] br[101] wl[225] vdd gnd cell_6t
Xbit_r226_c101 bl[101] br[101] wl[226] vdd gnd cell_6t
Xbit_r227_c101 bl[101] br[101] wl[227] vdd gnd cell_6t
Xbit_r228_c101 bl[101] br[101] wl[228] vdd gnd cell_6t
Xbit_r229_c101 bl[101] br[101] wl[229] vdd gnd cell_6t
Xbit_r230_c101 bl[101] br[101] wl[230] vdd gnd cell_6t
Xbit_r231_c101 bl[101] br[101] wl[231] vdd gnd cell_6t
Xbit_r232_c101 bl[101] br[101] wl[232] vdd gnd cell_6t
Xbit_r233_c101 bl[101] br[101] wl[233] vdd gnd cell_6t
Xbit_r234_c101 bl[101] br[101] wl[234] vdd gnd cell_6t
Xbit_r235_c101 bl[101] br[101] wl[235] vdd gnd cell_6t
Xbit_r236_c101 bl[101] br[101] wl[236] vdd gnd cell_6t
Xbit_r237_c101 bl[101] br[101] wl[237] vdd gnd cell_6t
Xbit_r238_c101 bl[101] br[101] wl[238] vdd gnd cell_6t
Xbit_r239_c101 bl[101] br[101] wl[239] vdd gnd cell_6t
Xbit_r240_c101 bl[101] br[101] wl[240] vdd gnd cell_6t
Xbit_r241_c101 bl[101] br[101] wl[241] vdd gnd cell_6t
Xbit_r242_c101 bl[101] br[101] wl[242] vdd gnd cell_6t
Xbit_r243_c101 bl[101] br[101] wl[243] vdd gnd cell_6t
Xbit_r244_c101 bl[101] br[101] wl[244] vdd gnd cell_6t
Xbit_r245_c101 bl[101] br[101] wl[245] vdd gnd cell_6t
Xbit_r246_c101 bl[101] br[101] wl[246] vdd gnd cell_6t
Xbit_r247_c101 bl[101] br[101] wl[247] vdd gnd cell_6t
Xbit_r248_c101 bl[101] br[101] wl[248] vdd gnd cell_6t
Xbit_r249_c101 bl[101] br[101] wl[249] vdd gnd cell_6t
Xbit_r250_c101 bl[101] br[101] wl[250] vdd gnd cell_6t
Xbit_r251_c101 bl[101] br[101] wl[251] vdd gnd cell_6t
Xbit_r252_c101 bl[101] br[101] wl[252] vdd gnd cell_6t
Xbit_r253_c101 bl[101] br[101] wl[253] vdd gnd cell_6t
Xbit_r254_c101 bl[101] br[101] wl[254] vdd gnd cell_6t
Xbit_r255_c101 bl[101] br[101] wl[255] vdd gnd cell_6t
Xbit_r256_c101 bl[101] br[101] wl[256] vdd gnd cell_6t
Xbit_r257_c101 bl[101] br[101] wl[257] vdd gnd cell_6t
Xbit_r258_c101 bl[101] br[101] wl[258] vdd gnd cell_6t
Xbit_r259_c101 bl[101] br[101] wl[259] vdd gnd cell_6t
Xbit_r260_c101 bl[101] br[101] wl[260] vdd gnd cell_6t
Xbit_r261_c101 bl[101] br[101] wl[261] vdd gnd cell_6t
Xbit_r262_c101 bl[101] br[101] wl[262] vdd gnd cell_6t
Xbit_r263_c101 bl[101] br[101] wl[263] vdd gnd cell_6t
Xbit_r264_c101 bl[101] br[101] wl[264] vdd gnd cell_6t
Xbit_r265_c101 bl[101] br[101] wl[265] vdd gnd cell_6t
Xbit_r266_c101 bl[101] br[101] wl[266] vdd gnd cell_6t
Xbit_r267_c101 bl[101] br[101] wl[267] vdd gnd cell_6t
Xbit_r268_c101 bl[101] br[101] wl[268] vdd gnd cell_6t
Xbit_r269_c101 bl[101] br[101] wl[269] vdd gnd cell_6t
Xbit_r270_c101 bl[101] br[101] wl[270] vdd gnd cell_6t
Xbit_r271_c101 bl[101] br[101] wl[271] vdd gnd cell_6t
Xbit_r272_c101 bl[101] br[101] wl[272] vdd gnd cell_6t
Xbit_r273_c101 bl[101] br[101] wl[273] vdd gnd cell_6t
Xbit_r274_c101 bl[101] br[101] wl[274] vdd gnd cell_6t
Xbit_r275_c101 bl[101] br[101] wl[275] vdd gnd cell_6t
Xbit_r276_c101 bl[101] br[101] wl[276] vdd gnd cell_6t
Xbit_r277_c101 bl[101] br[101] wl[277] vdd gnd cell_6t
Xbit_r278_c101 bl[101] br[101] wl[278] vdd gnd cell_6t
Xbit_r279_c101 bl[101] br[101] wl[279] vdd gnd cell_6t
Xbit_r280_c101 bl[101] br[101] wl[280] vdd gnd cell_6t
Xbit_r281_c101 bl[101] br[101] wl[281] vdd gnd cell_6t
Xbit_r282_c101 bl[101] br[101] wl[282] vdd gnd cell_6t
Xbit_r283_c101 bl[101] br[101] wl[283] vdd gnd cell_6t
Xbit_r284_c101 bl[101] br[101] wl[284] vdd gnd cell_6t
Xbit_r285_c101 bl[101] br[101] wl[285] vdd gnd cell_6t
Xbit_r286_c101 bl[101] br[101] wl[286] vdd gnd cell_6t
Xbit_r287_c101 bl[101] br[101] wl[287] vdd gnd cell_6t
Xbit_r288_c101 bl[101] br[101] wl[288] vdd gnd cell_6t
Xbit_r289_c101 bl[101] br[101] wl[289] vdd gnd cell_6t
Xbit_r290_c101 bl[101] br[101] wl[290] vdd gnd cell_6t
Xbit_r291_c101 bl[101] br[101] wl[291] vdd gnd cell_6t
Xbit_r292_c101 bl[101] br[101] wl[292] vdd gnd cell_6t
Xbit_r293_c101 bl[101] br[101] wl[293] vdd gnd cell_6t
Xbit_r294_c101 bl[101] br[101] wl[294] vdd gnd cell_6t
Xbit_r295_c101 bl[101] br[101] wl[295] vdd gnd cell_6t
Xbit_r296_c101 bl[101] br[101] wl[296] vdd gnd cell_6t
Xbit_r297_c101 bl[101] br[101] wl[297] vdd gnd cell_6t
Xbit_r298_c101 bl[101] br[101] wl[298] vdd gnd cell_6t
Xbit_r299_c101 bl[101] br[101] wl[299] vdd gnd cell_6t
Xbit_r300_c101 bl[101] br[101] wl[300] vdd gnd cell_6t
Xbit_r301_c101 bl[101] br[101] wl[301] vdd gnd cell_6t
Xbit_r302_c101 bl[101] br[101] wl[302] vdd gnd cell_6t
Xbit_r303_c101 bl[101] br[101] wl[303] vdd gnd cell_6t
Xbit_r304_c101 bl[101] br[101] wl[304] vdd gnd cell_6t
Xbit_r305_c101 bl[101] br[101] wl[305] vdd gnd cell_6t
Xbit_r306_c101 bl[101] br[101] wl[306] vdd gnd cell_6t
Xbit_r307_c101 bl[101] br[101] wl[307] vdd gnd cell_6t
Xbit_r308_c101 bl[101] br[101] wl[308] vdd gnd cell_6t
Xbit_r309_c101 bl[101] br[101] wl[309] vdd gnd cell_6t
Xbit_r310_c101 bl[101] br[101] wl[310] vdd gnd cell_6t
Xbit_r311_c101 bl[101] br[101] wl[311] vdd gnd cell_6t
Xbit_r312_c101 bl[101] br[101] wl[312] vdd gnd cell_6t
Xbit_r313_c101 bl[101] br[101] wl[313] vdd gnd cell_6t
Xbit_r314_c101 bl[101] br[101] wl[314] vdd gnd cell_6t
Xbit_r315_c101 bl[101] br[101] wl[315] vdd gnd cell_6t
Xbit_r316_c101 bl[101] br[101] wl[316] vdd gnd cell_6t
Xbit_r317_c101 bl[101] br[101] wl[317] vdd gnd cell_6t
Xbit_r318_c101 bl[101] br[101] wl[318] vdd gnd cell_6t
Xbit_r319_c101 bl[101] br[101] wl[319] vdd gnd cell_6t
Xbit_r320_c101 bl[101] br[101] wl[320] vdd gnd cell_6t
Xbit_r321_c101 bl[101] br[101] wl[321] vdd gnd cell_6t
Xbit_r322_c101 bl[101] br[101] wl[322] vdd gnd cell_6t
Xbit_r323_c101 bl[101] br[101] wl[323] vdd gnd cell_6t
Xbit_r324_c101 bl[101] br[101] wl[324] vdd gnd cell_6t
Xbit_r325_c101 bl[101] br[101] wl[325] vdd gnd cell_6t
Xbit_r326_c101 bl[101] br[101] wl[326] vdd gnd cell_6t
Xbit_r327_c101 bl[101] br[101] wl[327] vdd gnd cell_6t
Xbit_r328_c101 bl[101] br[101] wl[328] vdd gnd cell_6t
Xbit_r329_c101 bl[101] br[101] wl[329] vdd gnd cell_6t
Xbit_r330_c101 bl[101] br[101] wl[330] vdd gnd cell_6t
Xbit_r331_c101 bl[101] br[101] wl[331] vdd gnd cell_6t
Xbit_r332_c101 bl[101] br[101] wl[332] vdd gnd cell_6t
Xbit_r333_c101 bl[101] br[101] wl[333] vdd gnd cell_6t
Xbit_r334_c101 bl[101] br[101] wl[334] vdd gnd cell_6t
Xbit_r335_c101 bl[101] br[101] wl[335] vdd gnd cell_6t
Xbit_r336_c101 bl[101] br[101] wl[336] vdd gnd cell_6t
Xbit_r337_c101 bl[101] br[101] wl[337] vdd gnd cell_6t
Xbit_r338_c101 bl[101] br[101] wl[338] vdd gnd cell_6t
Xbit_r339_c101 bl[101] br[101] wl[339] vdd gnd cell_6t
Xbit_r340_c101 bl[101] br[101] wl[340] vdd gnd cell_6t
Xbit_r341_c101 bl[101] br[101] wl[341] vdd gnd cell_6t
Xbit_r342_c101 bl[101] br[101] wl[342] vdd gnd cell_6t
Xbit_r343_c101 bl[101] br[101] wl[343] vdd gnd cell_6t
Xbit_r344_c101 bl[101] br[101] wl[344] vdd gnd cell_6t
Xbit_r345_c101 bl[101] br[101] wl[345] vdd gnd cell_6t
Xbit_r346_c101 bl[101] br[101] wl[346] vdd gnd cell_6t
Xbit_r347_c101 bl[101] br[101] wl[347] vdd gnd cell_6t
Xbit_r348_c101 bl[101] br[101] wl[348] vdd gnd cell_6t
Xbit_r349_c101 bl[101] br[101] wl[349] vdd gnd cell_6t
Xbit_r350_c101 bl[101] br[101] wl[350] vdd gnd cell_6t
Xbit_r351_c101 bl[101] br[101] wl[351] vdd gnd cell_6t
Xbit_r352_c101 bl[101] br[101] wl[352] vdd gnd cell_6t
Xbit_r353_c101 bl[101] br[101] wl[353] vdd gnd cell_6t
Xbit_r354_c101 bl[101] br[101] wl[354] vdd gnd cell_6t
Xbit_r355_c101 bl[101] br[101] wl[355] vdd gnd cell_6t
Xbit_r356_c101 bl[101] br[101] wl[356] vdd gnd cell_6t
Xbit_r357_c101 bl[101] br[101] wl[357] vdd gnd cell_6t
Xbit_r358_c101 bl[101] br[101] wl[358] vdd gnd cell_6t
Xbit_r359_c101 bl[101] br[101] wl[359] vdd gnd cell_6t
Xbit_r360_c101 bl[101] br[101] wl[360] vdd gnd cell_6t
Xbit_r361_c101 bl[101] br[101] wl[361] vdd gnd cell_6t
Xbit_r362_c101 bl[101] br[101] wl[362] vdd gnd cell_6t
Xbit_r363_c101 bl[101] br[101] wl[363] vdd gnd cell_6t
Xbit_r364_c101 bl[101] br[101] wl[364] vdd gnd cell_6t
Xbit_r365_c101 bl[101] br[101] wl[365] vdd gnd cell_6t
Xbit_r366_c101 bl[101] br[101] wl[366] vdd gnd cell_6t
Xbit_r367_c101 bl[101] br[101] wl[367] vdd gnd cell_6t
Xbit_r368_c101 bl[101] br[101] wl[368] vdd gnd cell_6t
Xbit_r369_c101 bl[101] br[101] wl[369] vdd gnd cell_6t
Xbit_r370_c101 bl[101] br[101] wl[370] vdd gnd cell_6t
Xbit_r371_c101 bl[101] br[101] wl[371] vdd gnd cell_6t
Xbit_r372_c101 bl[101] br[101] wl[372] vdd gnd cell_6t
Xbit_r373_c101 bl[101] br[101] wl[373] vdd gnd cell_6t
Xbit_r374_c101 bl[101] br[101] wl[374] vdd gnd cell_6t
Xbit_r375_c101 bl[101] br[101] wl[375] vdd gnd cell_6t
Xbit_r376_c101 bl[101] br[101] wl[376] vdd gnd cell_6t
Xbit_r377_c101 bl[101] br[101] wl[377] vdd gnd cell_6t
Xbit_r378_c101 bl[101] br[101] wl[378] vdd gnd cell_6t
Xbit_r379_c101 bl[101] br[101] wl[379] vdd gnd cell_6t
Xbit_r380_c101 bl[101] br[101] wl[380] vdd gnd cell_6t
Xbit_r381_c101 bl[101] br[101] wl[381] vdd gnd cell_6t
Xbit_r382_c101 bl[101] br[101] wl[382] vdd gnd cell_6t
Xbit_r383_c101 bl[101] br[101] wl[383] vdd gnd cell_6t
Xbit_r384_c101 bl[101] br[101] wl[384] vdd gnd cell_6t
Xbit_r385_c101 bl[101] br[101] wl[385] vdd gnd cell_6t
Xbit_r386_c101 bl[101] br[101] wl[386] vdd gnd cell_6t
Xbit_r387_c101 bl[101] br[101] wl[387] vdd gnd cell_6t
Xbit_r388_c101 bl[101] br[101] wl[388] vdd gnd cell_6t
Xbit_r389_c101 bl[101] br[101] wl[389] vdd gnd cell_6t
Xbit_r390_c101 bl[101] br[101] wl[390] vdd gnd cell_6t
Xbit_r391_c101 bl[101] br[101] wl[391] vdd gnd cell_6t
Xbit_r392_c101 bl[101] br[101] wl[392] vdd gnd cell_6t
Xbit_r393_c101 bl[101] br[101] wl[393] vdd gnd cell_6t
Xbit_r394_c101 bl[101] br[101] wl[394] vdd gnd cell_6t
Xbit_r395_c101 bl[101] br[101] wl[395] vdd gnd cell_6t
Xbit_r396_c101 bl[101] br[101] wl[396] vdd gnd cell_6t
Xbit_r397_c101 bl[101] br[101] wl[397] vdd gnd cell_6t
Xbit_r398_c101 bl[101] br[101] wl[398] vdd gnd cell_6t
Xbit_r399_c101 bl[101] br[101] wl[399] vdd gnd cell_6t
Xbit_r400_c101 bl[101] br[101] wl[400] vdd gnd cell_6t
Xbit_r401_c101 bl[101] br[101] wl[401] vdd gnd cell_6t
Xbit_r402_c101 bl[101] br[101] wl[402] vdd gnd cell_6t
Xbit_r403_c101 bl[101] br[101] wl[403] vdd gnd cell_6t
Xbit_r404_c101 bl[101] br[101] wl[404] vdd gnd cell_6t
Xbit_r405_c101 bl[101] br[101] wl[405] vdd gnd cell_6t
Xbit_r406_c101 bl[101] br[101] wl[406] vdd gnd cell_6t
Xbit_r407_c101 bl[101] br[101] wl[407] vdd gnd cell_6t
Xbit_r408_c101 bl[101] br[101] wl[408] vdd gnd cell_6t
Xbit_r409_c101 bl[101] br[101] wl[409] vdd gnd cell_6t
Xbit_r410_c101 bl[101] br[101] wl[410] vdd gnd cell_6t
Xbit_r411_c101 bl[101] br[101] wl[411] vdd gnd cell_6t
Xbit_r412_c101 bl[101] br[101] wl[412] vdd gnd cell_6t
Xbit_r413_c101 bl[101] br[101] wl[413] vdd gnd cell_6t
Xbit_r414_c101 bl[101] br[101] wl[414] vdd gnd cell_6t
Xbit_r415_c101 bl[101] br[101] wl[415] vdd gnd cell_6t
Xbit_r416_c101 bl[101] br[101] wl[416] vdd gnd cell_6t
Xbit_r417_c101 bl[101] br[101] wl[417] vdd gnd cell_6t
Xbit_r418_c101 bl[101] br[101] wl[418] vdd gnd cell_6t
Xbit_r419_c101 bl[101] br[101] wl[419] vdd gnd cell_6t
Xbit_r420_c101 bl[101] br[101] wl[420] vdd gnd cell_6t
Xbit_r421_c101 bl[101] br[101] wl[421] vdd gnd cell_6t
Xbit_r422_c101 bl[101] br[101] wl[422] vdd gnd cell_6t
Xbit_r423_c101 bl[101] br[101] wl[423] vdd gnd cell_6t
Xbit_r424_c101 bl[101] br[101] wl[424] vdd gnd cell_6t
Xbit_r425_c101 bl[101] br[101] wl[425] vdd gnd cell_6t
Xbit_r426_c101 bl[101] br[101] wl[426] vdd gnd cell_6t
Xbit_r427_c101 bl[101] br[101] wl[427] vdd gnd cell_6t
Xbit_r428_c101 bl[101] br[101] wl[428] vdd gnd cell_6t
Xbit_r429_c101 bl[101] br[101] wl[429] vdd gnd cell_6t
Xbit_r430_c101 bl[101] br[101] wl[430] vdd gnd cell_6t
Xbit_r431_c101 bl[101] br[101] wl[431] vdd gnd cell_6t
Xbit_r432_c101 bl[101] br[101] wl[432] vdd gnd cell_6t
Xbit_r433_c101 bl[101] br[101] wl[433] vdd gnd cell_6t
Xbit_r434_c101 bl[101] br[101] wl[434] vdd gnd cell_6t
Xbit_r435_c101 bl[101] br[101] wl[435] vdd gnd cell_6t
Xbit_r436_c101 bl[101] br[101] wl[436] vdd gnd cell_6t
Xbit_r437_c101 bl[101] br[101] wl[437] vdd gnd cell_6t
Xbit_r438_c101 bl[101] br[101] wl[438] vdd gnd cell_6t
Xbit_r439_c101 bl[101] br[101] wl[439] vdd gnd cell_6t
Xbit_r440_c101 bl[101] br[101] wl[440] vdd gnd cell_6t
Xbit_r441_c101 bl[101] br[101] wl[441] vdd gnd cell_6t
Xbit_r442_c101 bl[101] br[101] wl[442] vdd gnd cell_6t
Xbit_r443_c101 bl[101] br[101] wl[443] vdd gnd cell_6t
Xbit_r444_c101 bl[101] br[101] wl[444] vdd gnd cell_6t
Xbit_r445_c101 bl[101] br[101] wl[445] vdd gnd cell_6t
Xbit_r446_c101 bl[101] br[101] wl[446] vdd gnd cell_6t
Xbit_r447_c101 bl[101] br[101] wl[447] vdd gnd cell_6t
Xbit_r448_c101 bl[101] br[101] wl[448] vdd gnd cell_6t
Xbit_r449_c101 bl[101] br[101] wl[449] vdd gnd cell_6t
Xbit_r450_c101 bl[101] br[101] wl[450] vdd gnd cell_6t
Xbit_r451_c101 bl[101] br[101] wl[451] vdd gnd cell_6t
Xbit_r452_c101 bl[101] br[101] wl[452] vdd gnd cell_6t
Xbit_r453_c101 bl[101] br[101] wl[453] vdd gnd cell_6t
Xbit_r454_c101 bl[101] br[101] wl[454] vdd gnd cell_6t
Xbit_r455_c101 bl[101] br[101] wl[455] vdd gnd cell_6t
Xbit_r456_c101 bl[101] br[101] wl[456] vdd gnd cell_6t
Xbit_r457_c101 bl[101] br[101] wl[457] vdd gnd cell_6t
Xbit_r458_c101 bl[101] br[101] wl[458] vdd gnd cell_6t
Xbit_r459_c101 bl[101] br[101] wl[459] vdd gnd cell_6t
Xbit_r460_c101 bl[101] br[101] wl[460] vdd gnd cell_6t
Xbit_r461_c101 bl[101] br[101] wl[461] vdd gnd cell_6t
Xbit_r462_c101 bl[101] br[101] wl[462] vdd gnd cell_6t
Xbit_r463_c101 bl[101] br[101] wl[463] vdd gnd cell_6t
Xbit_r464_c101 bl[101] br[101] wl[464] vdd gnd cell_6t
Xbit_r465_c101 bl[101] br[101] wl[465] vdd gnd cell_6t
Xbit_r466_c101 bl[101] br[101] wl[466] vdd gnd cell_6t
Xbit_r467_c101 bl[101] br[101] wl[467] vdd gnd cell_6t
Xbit_r468_c101 bl[101] br[101] wl[468] vdd gnd cell_6t
Xbit_r469_c101 bl[101] br[101] wl[469] vdd gnd cell_6t
Xbit_r470_c101 bl[101] br[101] wl[470] vdd gnd cell_6t
Xbit_r471_c101 bl[101] br[101] wl[471] vdd gnd cell_6t
Xbit_r472_c101 bl[101] br[101] wl[472] vdd gnd cell_6t
Xbit_r473_c101 bl[101] br[101] wl[473] vdd gnd cell_6t
Xbit_r474_c101 bl[101] br[101] wl[474] vdd gnd cell_6t
Xbit_r475_c101 bl[101] br[101] wl[475] vdd gnd cell_6t
Xbit_r476_c101 bl[101] br[101] wl[476] vdd gnd cell_6t
Xbit_r477_c101 bl[101] br[101] wl[477] vdd gnd cell_6t
Xbit_r478_c101 bl[101] br[101] wl[478] vdd gnd cell_6t
Xbit_r479_c101 bl[101] br[101] wl[479] vdd gnd cell_6t
Xbit_r480_c101 bl[101] br[101] wl[480] vdd gnd cell_6t
Xbit_r481_c101 bl[101] br[101] wl[481] vdd gnd cell_6t
Xbit_r482_c101 bl[101] br[101] wl[482] vdd gnd cell_6t
Xbit_r483_c101 bl[101] br[101] wl[483] vdd gnd cell_6t
Xbit_r484_c101 bl[101] br[101] wl[484] vdd gnd cell_6t
Xbit_r485_c101 bl[101] br[101] wl[485] vdd gnd cell_6t
Xbit_r486_c101 bl[101] br[101] wl[486] vdd gnd cell_6t
Xbit_r487_c101 bl[101] br[101] wl[487] vdd gnd cell_6t
Xbit_r488_c101 bl[101] br[101] wl[488] vdd gnd cell_6t
Xbit_r489_c101 bl[101] br[101] wl[489] vdd gnd cell_6t
Xbit_r490_c101 bl[101] br[101] wl[490] vdd gnd cell_6t
Xbit_r491_c101 bl[101] br[101] wl[491] vdd gnd cell_6t
Xbit_r492_c101 bl[101] br[101] wl[492] vdd gnd cell_6t
Xbit_r493_c101 bl[101] br[101] wl[493] vdd gnd cell_6t
Xbit_r494_c101 bl[101] br[101] wl[494] vdd gnd cell_6t
Xbit_r495_c101 bl[101] br[101] wl[495] vdd gnd cell_6t
Xbit_r496_c101 bl[101] br[101] wl[496] vdd gnd cell_6t
Xbit_r497_c101 bl[101] br[101] wl[497] vdd gnd cell_6t
Xbit_r498_c101 bl[101] br[101] wl[498] vdd gnd cell_6t
Xbit_r499_c101 bl[101] br[101] wl[499] vdd gnd cell_6t
Xbit_r500_c101 bl[101] br[101] wl[500] vdd gnd cell_6t
Xbit_r501_c101 bl[101] br[101] wl[501] vdd gnd cell_6t
Xbit_r502_c101 bl[101] br[101] wl[502] vdd gnd cell_6t
Xbit_r503_c101 bl[101] br[101] wl[503] vdd gnd cell_6t
Xbit_r504_c101 bl[101] br[101] wl[504] vdd gnd cell_6t
Xbit_r505_c101 bl[101] br[101] wl[505] vdd gnd cell_6t
Xbit_r506_c101 bl[101] br[101] wl[506] vdd gnd cell_6t
Xbit_r507_c101 bl[101] br[101] wl[507] vdd gnd cell_6t
Xbit_r508_c101 bl[101] br[101] wl[508] vdd gnd cell_6t
Xbit_r509_c101 bl[101] br[101] wl[509] vdd gnd cell_6t
Xbit_r510_c101 bl[101] br[101] wl[510] vdd gnd cell_6t
Xbit_r511_c101 bl[101] br[101] wl[511] vdd gnd cell_6t
Xbit_r0_c102 bl[102] br[102] wl[0] vdd gnd cell_6t
Xbit_r1_c102 bl[102] br[102] wl[1] vdd gnd cell_6t
Xbit_r2_c102 bl[102] br[102] wl[2] vdd gnd cell_6t
Xbit_r3_c102 bl[102] br[102] wl[3] vdd gnd cell_6t
Xbit_r4_c102 bl[102] br[102] wl[4] vdd gnd cell_6t
Xbit_r5_c102 bl[102] br[102] wl[5] vdd gnd cell_6t
Xbit_r6_c102 bl[102] br[102] wl[6] vdd gnd cell_6t
Xbit_r7_c102 bl[102] br[102] wl[7] vdd gnd cell_6t
Xbit_r8_c102 bl[102] br[102] wl[8] vdd gnd cell_6t
Xbit_r9_c102 bl[102] br[102] wl[9] vdd gnd cell_6t
Xbit_r10_c102 bl[102] br[102] wl[10] vdd gnd cell_6t
Xbit_r11_c102 bl[102] br[102] wl[11] vdd gnd cell_6t
Xbit_r12_c102 bl[102] br[102] wl[12] vdd gnd cell_6t
Xbit_r13_c102 bl[102] br[102] wl[13] vdd gnd cell_6t
Xbit_r14_c102 bl[102] br[102] wl[14] vdd gnd cell_6t
Xbit_r15_c102 bl[102] br[102] wl[15] vdd gnd cell_6t
Xbit_r16_c102 bl[102] br[102] wl[16] vdd gnd cell_6t
Xbit_r17_c102 bl[102] br[102] wl[17] vdd gnd cell_6t
Xbit_r18_c102 bl[102] br[102] wl[18] vdd gnd cell_6t
Xbit_r19_c102 bl[102] br[102] wl[19] vdd gnd cell_6t
Xbit_r20_c102 bl[102] br[102] wl[20] vdd gnd cell_6t
Xbit_r21_c102 bl[102] br[102] wl[21] vdd gnd cell_6t
Xbit_r22_c102 bl[102] br[102] wl[22] vdd gnd cell_6t
Xbit_r23_c102 bl[102] br[102] wl[23] vdd gnd cell_6t
Xbit_r24_c102 bl[102] br[102] wl[24] vdd gnd cell_6t
Xbit_r25_c102 bl[102] br[102] wl[25] vdd gnd cell_6t
Xbit_r26_c102 bl[102] br[102] wl[26] vdd gnd cell_6t
Xbit_r27_c102 bl[102] br[102] wl[27] vdd gnd cell_6t
Xbit_r28_c102 bl[102] br[102] wl[28] vdd gnd cell_6t
Xbit_r29_c102 bl[102] br[102] wl[29] vdd gnd cell_6t
Xbit_r30_c102 bl[102] br[102] wl[30] vdd gnd cell_6t
Xbit_r31_c102 bl[102] br[102] wl[31] vdd gnd cell_6t
Xbit_r32_c102 bl[102] br[102] wl[32] vdd gnd cell_6t
Xbit_r33_c102 bl[102] br[102] wl[33] vdd gnd cell_6t
Xbit_r34_c102 bl[102] br[102] wl[34] vdd gnd cell_6t
Xbit_r35_c102 bl[102] br[102] wl[35] vdd gnd cell_6t
Xbit_r36_c102 bl[102] br[102] wl[36] vdd gnd cell_6t
Xbit_r37_c102 bl[102] br[102] wl[37] vdd gnd cell_6t
Xbit_r38_c102 bl[102] br[102] wl[38] vdd gnd cell_6t
Xbit_r39_c102 bl[102] br[102] wl[39] vdd gnd cell_6t
Xbit_r40_c102 bl[102] br[102] wl[40] vdd gnd cell_6t
Xbit_r41_c102 bl[102] br[102] wl[41] vdd gnd cell_6t
Xbit_r42_c102 bl[102] br[102] wl[42] vdd gnd cell_6t
Xbit_r43_c102 bl[102] br[102] wl[43] vdd gnd cell_6t
Xbit_r44_c102 bl[102] br[102] wl[44] vdd gnd cell_6t
Xbit_r45_c102 bl[102] br[102] wl[45] vdd gnd cell_6t
Xbit_r46_c102 bl[102] br[102] wl[46] vdd gnd cell_6t
Xbit_r47_c102 bl[102] br[102] wl[47] vdd gnd cell_6t
Xbit_r48_c102 bl[102] br[102] wl[48] vdd gnd cell_6t
Xbit_r49_c102 bl[102] br[102] wl[49] vdd gnd cell_6t
Xbit_r50_c102 bl[102] br[102] wl[50] vdd gnd cell_6t
Xbit_r51_c102 bl[102] br[102] wl[51] vdd gnd cell_6t
Xbit_r52_c102 bl[102] br[102] wl[52] vdd gnd cell_6t
Xbit_r53_c102 bl[102] br[102] wl[53] vdd gnd cell_6t
Xbit_r54_c102 bl[102] br[102] wl[54] vdd gnd cell_6t
Xbit_r55_c102 bl[102] br[102] wl[55] vdd gnd cell_6t
Xbit_r56_c102 bl[102] br[102] wl[56] vdd gnd cell_6t
Xbit_r57_c102 bl[102] br[102] wl[57] vdd gnd cell_6t
Xbit_r58_c102 bl[102] br[102] wl[58] vdd gnd cell_6t
Xbit_r59_c102 bl[102] br[102] wl[59] vdd gnd cell_6t
Xbit_r60_c102 bl[102] br[102] wl[60] vdd gnd cell_6t
Xbit_r61_c102 bl[102] br[102] wl[61] vdd gnd cell_6t
Xbit_r62_c102 bl[102] br[102] wl[62] vdd gnd cell_6t
Xbit_r63_c102 bl[102] br[102] wl[63] vdd gnd cell_6t
Xbit_r64_c102 bl[102] br[102] wl[64] vdd gnd cell_6t
Xbit_r65_c102 bl[102] br[102] wl[65] vdd gnd cell_6t
Xbit_r66_c102 bl[102] br[102] wl[66] vdd gnd cell_6t
Xbit_r67_c102 bl[102] br[102] wl[67] vdd gnd cell_6t
Xbit_r68_c102 bl[102] br[102] wl[68] vdd gnd cell_6t
Xbit_r69_c102 bl[102] br[102] wl[69] vdd gnd cell_6t
Xbit_r70_c102 bl[102] br[102] wl[70] vdd gnd cell_6t
Xbit_r71_c102 bl[102] br[102] wl[71] vdd gnd cell_6t
Xbit_r72_c102 bl[102] br[102] wl[72] vdd gnd cell_6t
Xbit_r73_c102 bl[102] br[102] wl[73] vdd gnd cell_6t
Xbit_r74_c102 bl[102] br[102] wl[74] vdd gnd cell_6t
Xbit_r75_c102 bl[102] br[102] wl[75] vdd gnd cell_6t
Xbit_r76_c102 bl[102] br[102] wl[76] vdd gnd cell_6t
Xbit_r77_c102 bl[102] br[102] wl[77] vdd gnd cell_6t
Xbit_r78_c102 bl[102] br[102] wl[78] vdd gnd cell_6t
Xbit_r79_c102 bl[102] br[102] wl[79] vdd gnd cell_6t
Xbit_r80_c102 bl[102] br[102] wl[80] vdd gnd cell_6t
Xbit_r81_c102 bl[102] br[102] wl[81] vdd gnd cell_6t
Xbit_r82_c102 bl[102] br[102] wl[82] vdd gnd cell_6t
Xbit_r83_c102 bl[102] br[102] wl[83] vdd gnd cell_6t
Xbit_r84_c102 bl[102] br[102] wl[84] vdd gnd cell_6t
Xbit_r85_c102 bl[102] br[102] wl[85] vdd gnd cell_6t
Xbit_r86_c102 bl[102] br[102] wl[86] vdd gnd cell_6t
Xbit_r87_c102 bl[102] br[102] wl[87] vdd gnd cell_6t
Xbit_r88_c102 bl[102] br[102] wl[88] vdd gnd cell_6t
Xbit_r89_c102 bl[102] br[102] wl[89] vdd gnd cell_6t
Xbit_r90_c102 bl[102] br[102] wl[90] vdd gnd cell_6t
Xbit_r91_c102 bl[102] br[102] wl[91] vdd gnd cell_6t
Xbit_r92_c102 bl[102] br[102] wl[92] vdd gnd cell_6t
Xbit_r93_c102 bl[102] br[102] wl[93] vdd gnd cell_6t
Xbit_r94_c102 bl[102] br[102] wl[94] vdd gnd cell_6t
Xbit_r95_c102 bl[102] br[102] wl[95] vdd gnd cell_6t
Xbit_r96_c102 bl[102] br[102] wl[96] vdd gnd cell_6t
Xbit_r97_c102 bl[102] br[102] wl[97] vdd gnd cell_6t
Xbit_r98_c102 bl[102] br[102] wl[98] vdd gnd cell_6t
Xbit_r99_c102 bl[102] br[102] wl[99] vdd gnd cell_6t
Xbit_r100_c102 bl[102] br[102] wl[100] vdd gnd cell_6t
Xbit_r101_c102 bl[102] br[102] wl[101] vdd gnd cell_6t
Xbit_r102_c102 bl[102] br[102] wl[102] vdd gnd cell_6t
Xbit_r103_c102 bl[102] br[102] wl[103] vdd gnd cell_6t
Xbit_r104_c102 bl[102] br[102] wl[104] vdd gnd cell_6t
Xbit_r105_c102 bl[102] br[102] wl[105] vdd gnd cell_6t
Xbit_r106_c102 bl[102] br[102] wl[106] vdd gnd cell_6t
Xbit_r107_c102 bl[102] br[102] wl[107] vdd gnd cell_6t
Xbit_r108_c102 bl[102] br[102] wl[108] vdd gnd cell_6t
Xbit_r109_c102 bl[102] br[102] wl[109] vdd gnd cell_6t
Xbit_r110_c102 bl[102] br[102] wl[110] vdd gnd cell_6t
Xbit_r111_c102 bl[102] br[102] wl[111] vdd gnd cell_6t
Xbit_r112_c102 bl[102] br[102] wl[112] vdd gnd cell_6t
Xbit_r113_c102 bl[102] br[102] wl[113] vdd gnd cell_6t
Xbit_r114_c102 bl[102] br[102] wl[114] vdd gnd cell_6t
Xbit_r115_c102 bl[102] br[102] wl[115] vdd gnd cell_6t
Xbit_r116_c102 bl[102] br[102] wl[116] vdd gnd cell_6t
Xbit_r117_c102 bl[102] br[102] wl[117] vdd gnd cell_6t
Xbit_r118_c102 bl[102] br[102] wl[118] vdd gnd cell_6t
Xbit_r119_c102 bl[102] br[102] wl[119] vdd gnd cell_6t
Xbit_r120_c102 bl[102] br[102] wl[120] vdd gnd cell_6t
Xbit_r121_c102 bl[102] br[102] wl[121] vdd gnd cell_6t
Xbit_r122_c102 bl[102] br[102] wl[122] vdd gnd cell_6t
Xbit_r123_c102 bl[102] br[102] wl[123] vdd gnd cell_6t
Xbit_r124_c102 bl[102] br[102] wl[124] vdd gnd cell_6t
Xbit_r125_c102 bl[102] br[102] wl[125] vdd gnd cell_6t
Xbit_r126_c102 bl[102] br[102] wl[126] vdd gnd cell_6t
Xbit_r127_c102 bl[102] br[102] wl[127] vdd gnd cell_6t
Xbit_r128_c102 bl[102] br[102] wl[128] vdd gnd cell_6t
Xbit_r129_c102 bl[102] br[102] wl[129] vdd gnd cell_6t
Xbit_r130_c102 bl[102] br[102] wl[130] vdd gnd cell_6t
Xbit_r131_c102 bl[102] br[102] wl[131] vdd gnd cell_6t
Xbit_r132_c102 bl[102] br[102] wl[132] vdd gnd cell_6t
Xbit_r133_c102 bl[102] br[102] wl[133] vdd gnd cell_6t
Xbit_r134_c102 bl[102] br[102] wl[134] vdd gnd cell_6t
Xbit_r135_c102 bl[102] br[102] wl[135] vdd gnd cell_6t
Xbit_r136_c102 bl[102] br[102] wl[136] vdd gnd cell_6t
Xbit_r137_c102 bl[102] br[102] wl[137] vdd gnd cell_6t
Xbit_r138_c102 bl[102] br[102] wl[138] vdd gnd cell_6t
Xbit_r139_c102 bl[102] br[102] wl[139] vdd gnd cell_6t
Xbit_r140_c102 bl[102] br[102] wl[140] vdd gnd cell_6t
Xbit_r141_c102 bl[102] br[102] wl[141] vdd gnd cell_6t
Xbit_r142_c102 bl[102] br[102] wl[142] vdd gnd cell_6t
Xbit_r143_c102 bl[102] br[102] wl[143] vdd gnd cell_6t
Xbit_r144_c102 bl[102] br[102] wl[144] vdd gnd cell_6t
Xbit_r145_c102 bl[102] br[102] wl[145] vdd gnd cell_6t
Xbit_r146_c102 bl[102] br[102] wl[146] vdd gnd cell_6t
Xbit_r147_c102 bl[102] br[102] wl[147] vdd gnd cell_6t
Xbit_r148_c102 bl[102] br[102] wl[148] vdd gnd cell_6t
Xbit_r149_c102 bl[102] br[102] wl[149] vdd gnd cell_6t
Xbit_r150_c102 bl[102] br[102] wl[150] vdd gnd cell_6t
Xbit_r151_c102 bl[102] br[102] wl[151] vdd gnd cell_6t
Xbit_r152_c102 bl[102] br[102] wl[152] vdd gnd cell_6t
Xbit_r153_c102 bl[102] br[102] wl[153] vdd gnd cell_6t
Xbit_r154_c102 bl[102] br[102] wl[154] vdd gnd cell_6t
Xbit_r155_c102 bl[102] br[102] wl[155] vdd gnd cell_6t
Xbit_r156_c102 bl[102] br[102] wl[156] vdd gnd cell_6t
Xbit_r157_c102 bl[102] br[102] wl[157] vdd gnd cell_6t
Xbit_r158_c102 bl[102] br[102] wl[158] vdd gnd cell_6t
Xbit_r159_c102 bl[102] br[102] wl[159] vdd gnd cell_6t
Xbit_r160_c102 bl[102] br[102] wl[160] vdd gnd cell_6t
Xbit_r161_c102 bl[102] br[102] wl[161] vdd gnd cell_6t
Xbit_r162_c102 bl[102] br[102] wl[162] vdd gnd cell_6t
Xbit_r163_c102 bl[102] br[102] wl[163] vdd gnd cell_6t
Xbit_r164_c102 bl[102] br[102] wl[164] vdd gnd cell_6t
Xbit_r165_c102 bl[102] br[102] wl[165] vdd gnd cell_6t
Xbit_r166_c102 bl[102] br[102] wl[166] vdd gnd cell_6t
Xbit_r167_c102 bl[102] br[102] wl[167] vdd gnd cell_6t
Xbit_r168_c102 bl[102] br[102] wl[168] vdd gnd cell_6t
Xbit_r169_c102 bl[102] br[102] wl[169] vdd gnd cell_6t
Xbit_r170_c102 bl[102] br[102] wl[170] vdd gnd cell_6t
Xbit_r171_c102 bl[102] br[102] wl[171] vdd gnd cell_6t
Xbit_r172_c102 bl[102] br[102] wl[172] vdd gnd cell_6t
Xbit_r173_c102 bl[102] br[102] wl[173] vdd gnd cell_6t
Xbit_r174_c102 bl[102] br[102] wl[174] vdd gnd cell_6t
Xbit_r175_c102 bl[102] br[102] wl[175] vdd gnd cell_6t
Xbit_r176_c102 bl[102] br[102] wl[176] vdd gnd cell_6t
Xbit_r177_c102 bl[102] br[102] wl[177] vdd gnd cell_6t
Xbit_r178_c102 bl[102] br[102] wl[178] vdd gnd cell_6t
Xbit_r179_c102 bl[102] br[102] wl[179] vdd gnd cell_6t
Xbit_r180_c102 bl[102] br[102] wl[180] vdd gnd cell_6t
Xbit_r181_c102 bl[102] br[102] wl[181] vdd gnd cell_6t
Xbit_r182_c102 bl[102] br[102] wl[182] vdd gnd cell_6t
Xbit_r183_c102 bl[102] br[102] wl[183] vdd gnd cell_6t
Xbit_r184_c102 bl[102] br[102] wl[184] vdd gnd cell_6t
Xbit_r185_c102 bl[102] br[102] wl[185] vdd gnd cell_6t
Xbit_r186_c102 bl[102] br[102] wl[186] vdd gnd cell_6t
Xbit_r187_c102 bl[102] br[102] wl[187] vdd gnd cell_6t
Xbit_r188_c102 bl[102] br[102] wl[188] vdd gnd cell_6t
Xbit_r189_c102 bl[102] br[102] wl[189] vdd gnd cell_6t
Xbit_r190_c102 bl[102] br[102] wl[190] vdd gnd cell_6t
Xbit_r191_c102 bl[102] br[102] wl[191] vdd gnd cell_6t
Xbit_r192_c102 bl[102] br[102] wl[192] vdd gnd cell_6t
Xbit_r193_c102 bl[102] br[102] wl[193] vdd gnd cell_6t
Xbit_r194_c102 bl[102] br[102] wl[194] vdd gnd cell_6t
Xbit_r195_c102 bl[102] br[102] wl[195] vdd gnd cell_6t
Xbit_r196_c102 bl[102] br[102] wl[196] vdd gnd cell_6t
Xbit_r197_c102 bl[102] br[102] wl[197] vdd gnd cell_6t
Xbit_r198_c102 bl[102] br[102] wl[198] vdd gnd cell_6t
Xbit_r199_c102 bl[102] br[102] wl[199] vdd gnd cell_6t
Xbit_r200_c102 bl[102] br[102] wl[200] vdd gnd cell_6t
Xbit_r201_c102 bl[102] br[102] wl[201] vdd gnd cell_6t
Xbit_r202_c102 bl[102] br[102] wl[202] vdd gnd cell_6t
Xbit_r203_c102 bl[102] br[102] wl[203] vdd gnd cell_6t
Xbit_r204_c102 bl[102] br[102] wl[204] vdd gnd cell_6t
Xbit_r205_c102 bl[102] br[102] wl[205] vdd gnd cell_6t
Xbit_r206_c102 bl[102] br[102] wl[206] vdd gnd cell_6t
Xbit_r207_c102 bl[102] br[102] wl[207] vdd gnd cell_6t
Xbit_r208_c102 bl[102] br[102] wl[208] vdd gnd cell_6t
Xbit_r209_c102 bl[102] br[102] wl[209] vdd gnd cell_6t
Xbit_r210_c102 bl[102] br[102] wl[210] vdd gnd cell_6t
Xbit_r211_c102 bl[102] br[102] wl[211] vdd gnd cell_6t
Xbit_r212_c102 bl[102] br[102] wl[212] vdd gnd cell_6t
Xbit_r213_c102 bl[102] br[102] wl[213] vdd gnd cell_6t
Xbit_r214_c102 bl[102] br[102] wl[214] vdd gnd cell_6t
Xbit_r215_c102 bl[102] br[102] wl[215] vdd gnd cell_6t
Xbit_r216_c102 bl[102] br[102] wl[216] vdd gnd cell_6t
Xbit_r217_c102 bl[102] br[102] wl[217] vdd gnd cell_6t
Xbit_r218_c102 bl[102] br[102] wl[218] vdd gnd cell_6t
Xbit_r219_c102 bl[102] br[102] wl[219] vdd gnd cell_6t
Xbit_r220_c102 bl[102] br[102] wl[220] vdd gnd cell_6t
Xbit_r221_c102 bl[102] br[102] wl[221] vdd gnd cell_6t
Xbit_r222_c102 bl[102] br[102] wl[222] vdd gnd cell_6t
Xbit_r223_c102 bl[102] br[102] wl[223] vdd gnd cell_6t
Xbit_r224_c102 bl[102] br[102] wl[224] vdd gnd cell_6t
Xbit_r225_c102 bl[102] br[102] wl[225] vdd gnd cell_6t
Xbit_r226_c102 bl[102] br[102] wl[226] vdd gnd cell_6t
Xbit_r227_c102 bl[102] br[102] wl[227] vdd gnd cell_6t
Xbit_r228_c102 bl[102] br[102] wl[228] vdd gnd cell_6t
Xbit_r229_c102 bl[102] br[102] wl[229] vdd gnd cell_6t
Xbit_r230_c102 bl[102] br[102] wl[230] vdd gnd cell_6t
Xbit_r231_c102 bl[102] br[102] wl[231] vdd gnd cell_6t
Xbit_r232_c102 bl[102] br[102] wl[232] vdd gnd cell_6t
Xbit_r233_c102 bl[102] br[102] wl[233] vdd gnd cell_6t
Xbit_r234_c102 bl[102] br[102] wl[234] vdd gnd cell_6t
Xbit_r235_c102 bl[102] br[102] wl[235] vdd gnd cell_6t
Xbit_r236_c102 bl[102] br[102] wl[236] vdd gnd cell_6t
Xbit_r237_c102 bl[102] br[102] wl[237] vdd gnd cell_6t
Xbit_r238_c102 bl[102] br[102] wl[238] vdd gnd cell_6t
Xbit_r239_c102 bl[102] br[102] wl[239] vdd gnd cell_6t
Xbit_r240_c102 bl[102] br[102] wl[240] vdd gnd cell_6t
Xbit_r241_c102 bl[102] br[102] wl[241] vdd gnd cell_6t
Xbit_r242_c102 bl[102] br[102] wl[242] vdd gnd cell_6t
Xbit_r243_c102 bl[102] br[102] wl[243] vdd gnd cell_6t
Xbit_r244_c102 bl[102] br[102] wl[244] vdd gnd cell_6t
Xbit_r245_c102 bl[102] br[102] wl[245] vdd gnd cell_6t
Xbit_r246_c102 bl[102] br[102] wl[246] vdd gnd cell_6t
Xbit_r247_c102 bl[102] br[102] wl[247] vdd gnd cell_6t
Xbit_r248_c102 bl[102] br[102] wl[248] vdd gnd cell_6t
Xbit_r249_c102 bl[102] br[102] wl[249] vdd gnd cell_6t
Xbit_r250_c102 bl[102] br[102] wl[250] vdd gnd cell_6t
Xbit_r251_c102 bl[102] br[102] wl[251] vdd gnd cell_6t
Xbit_r252_c102 bl[102] br[102] wl[252] vdd gnd cell_6t
Xbit_r253_c102 bl[102] br[102] wl[253] vdd gnd cell_6t
Xbit_r254_c102 bl[102] br[102] wl[254] vdd gnd cell_6t
Xbit_r255_c102 bl[102] br[102] wl[255] vdd gnd cell_6t
Xbit_r256_c102 bl[102] br[102] wl[256] vdd gnd cell_6t
Xbit_r257_c102 bl[102] br[102] wl[257] vdd gnd cell_6t
Xbit_r258_c102 bl[102] br[102] wl[258] vdd gnd cell_6t
Xbit_r259_c102 bl[102] br[102] wl[259] vdd gnd cell_6t
Xbit_r260_c102 bl[102] br[102] wl[260] vdd gnd cell_6t
Xbit_r261_c102 bl[102] br[102] wl[261] vdd gnd cell_6t
Xbit_r262_c102 bl[102] br[102] wl[262] vdd gnd cell_6t
Xbit_r263_c102 bl[102] br[102] wl[263] vdd gnd cell_6t
Xbit_r264_c102 bl[102] br[102] wl[264] vdd gnd cell_6t
Xbit_r265_c102 bl[102] br[102] wl[265] vdd gnd cell_6t
Xbit_r266_c102 bl[102] br[102] wl[266] vdd gnd cell_6t
Xbit_r267_c102 bl[102] br[102] wl[267] vdd gnd cell_6t
Xbit_r268_c102 bl[102] br[102] wl[268] vdd gnd cell_6t
Xbit_r269_c102 bl[102] br[102] wl[269] vdd gnd cell_6t
Xbit_r270_c102 bl[102] br[102] wl[270] vdd gnd cell_6t
Xbit_r271_c102 bl[102] br[102] wl[271] vdd gnd cell_6t
Xbit_r272_c102 bl[102] br[102] wl[272] vdd gnd cell_6t
Xbit_r273_c102 bl[102] br[102] wl[273] vdd gnd cell_6t
Xbit_r274_c102 bl[102] br[102] wl[274] vdd gnd cell_6t
Xbit_r275_c102 bl[102] br[102] wl[275] vdd gnd cell_6t
Xbit_r276_c102 bl[102] br[102] wl[276] vdd gnd cell_6t
Xbit_r277_c102 bl[102] br[102] wl[277] vdd gnd cell_6t
Xbit_r278_c102 bl[102] br[102] wl[278] vdd gnd cell_6t
Xbit_r279_c102 bl[102] br[102] wl[279] vdd gnd cell_6t
Xbit_r280_c102 bl[102] br[102] wl[280] vdd gnd cell_6t
Xbit_r281_c102 bl[102] br[102] wl[281] vdd gnd cell_6t
Xbit_r282_c102 bl[102] br[102] wl[282] vdd gnd cell_6t
Xbit_r283_c102 bl[102] br[102] wl[283] vdd gnd cell_6t
Xbit_r284_c102 bl[102] br[102] wl[284] vdd gnd cell_6t
Xbit_r285_c102 bl[102] br[102] wl[285] vdd gnd cell_6t
Xbit_r286_c102 bl[102] br[102] wl[286] vdd gnd cell_6t
Xbit_r287_c102 bl[102] br[102] wl[287] vdd gnd cell_6t
Xbit_r288_c102 bl[102] br[102] wl[288] vdd gnd cell_6t
Xbit_r289_c102 bl[102] br[102] wl[289] vdd gnd cell_6t
Xbit_r290_c102 bl[102] br[102] wl[290] vdd gnd cell_6t
Xbit_r291_c102 bl[102] br[102] wl[291] vdd gnd cell_6t
Xbit_r292_c102 bl[102] br[102] wl[292] vdd gnd cell_6t
Xbit_r293_c102 bl[102] br[102] wl[293] vdd gnd cell_6t
Xbit_r294_c102 bl[102] br[102] wl[294] vdd gnd cell_6t
Xbit_r295_c102 bl[102] br[102] wl[295] vdd gnd cell_6t
Xbit_r296_c102 bl[102] br[102] wl[296] vdd gnd cell_6t
Xbit_r297_c102 bl[102] br[102] wl[297] vdd gnd cell_6t
Xbit_r298_c102 bl[102] br[102] wl[298] vdd gnd cell_6t
Xbit_r299_c102 bl[102] br[102] wl[299] vdd gnd cell_6t
Xbit_r300_c102 bl[102] br[102] wl[300] vdd gnd cell_6t
Xbit_r301_c102 bl[102] br[102] wl[301] vdd gnd cell_6t
Xbit_r302_c102 bl[102] br[102] wl[302] vdd gnd cell_6t
Xbit_r303_c102 bl[102] br[102] wl[303] vdd gnd cell_6t
Xbit_r304_c102 bl[102] br[102] wl[304] vdd gnd cell_6t
Xbit_r305_c102 bl[102] br[102] wl[305] vdd gnd cell_6t
Xbit_r306_c102 bl[102] br[102] wl[306] vdd gnd cell_6t
Xbit_r307_c102 bl[102] br[102] wl[307] vdd gnd cell_6t
Xbit_r308_c102 bl[102] br[102] wl[308] vdd gnd cell_6t
Xbit_r309_c102 bl[102] br[102] wl[309] vdd gnd cell_6t
Xbit_r310_c102 bl[102] br[102] wl[310] vdd gnd cell_6t
Xbit_r311_c102 bl[102] br[102] wl[311] vdd gnd cell_6t
Xbit_r312_c102 bl[102] br[102] wl[312] vdd gnd cell_6t
Xbit_r313_c102 bl[102] br[102] wl[313] vdd gnd cell_6t
Xbit_r314_c102 bl[102] br[102] wl[314] vdd gnd cell_6t
Xbit_r315_c102 bl[102] br[102] wl[315] vdd gnd cell_6t
Xbit_r316_c102 bl[102] br[102] wl[316] vdd gnd cell_6t
Xbit_r317_c102 bl[102] br[102] wl[317] vdd gnd cell_6t
Xbit_r318_c102 bl[102] br[102] wl[318] vdd gnd cell_6t
Xbit_r319_c102 bl[102] br[102] wl[319] vdd gnd cell_6t
Xbit_r320_c102 bl[102] br[102] wl[320] vdd gnd cell_6t
Xbit_r321_c102 bl[102] br[102] wl[321] vdd gnd cell_6t
Xbit_r322_c102 bl[102] br[102] wl[322] vdd gnd cell_6t
Xbit_r323_c102 bl[102] br[102] wl[323] vdd gnd cell_6t
Xbit_r324_c102 bl[102] br[102] wl[324] vdd gnd cell_6t
Xbit_r325_c102 bl[102] br[102] wl[325] vdd gnd cell_6t
Xbit_r326_c102 bl[102] br[102] wl[326] vdd gnd cell_6t
Xbit_r327_c102 bl[102] br[102] wl[327] vdd gnd cell_6t
Xbit_r328_c102 bl[102] br[102] wl[328] vdd gnd cell_6t
Xbit_r329_c102 bl[102] br[102] wl[329] vdd gnd cell_6t
Xbit_r330_c102 bl[102] br[102] wl[330] vdd gnd cell_6t
Xbit_r331_c102 bl[102] br[102] wl[331] vdd gnd cell_6t
Xbit_r332_c102 bl[102] br[102] wl[332] vdd gnd cell_6t
Xbit_r333_c102 bl[102] br[102] wl[333] vdd gnd cell_6t
Xbit_r334_c102 bl[102] br[102] wl[334] vdd gnd cell_6t
Xbit_r335_c102 bl[102] br[102] wl[335] vdd gnd cell_6t
Xbit_r336_c102 bl[102] br[102] wl[336] vdd gnd cell_6t
Xbit_r337_c102 bl[102] br[102] wl[337] vdd gnd cell_6t
Xbit_r338_c102 bl[102] br[102] wl[338] vdd gnd cell_6t
Xbit_r339_c102 bl[102] br[102] wl[339] vdd gnd cell_6t
Xbit_r340_c102 bl[102] br[102] wl[340] vdd gnd cell_6t
Xbit_r341_c102 bl[102] br[102] wl[341] vdd gnd cell_6t
Xbit_r342_c102 bl[102] br[102] wl[342] vdd gnd cell_6t
Xbit_r343_c102 bl[102] br[102] wl[343] vdd gnd cell_6t
Xbit_r344_c102 bl[102] br[102] wl[344] vdd gnd cell_6t
Xbit_r345_c102 bl[102] br[102] wl[345] vdd gnd cell_6t
Xbit_r346_c102 bl[102] br[102] wl[346] vdd gnd cell_6t
Xbit_r347_c102 bl[102] br[102] wl[347] vdd gnd cell_6t
Xbit_r348_c102 bl[102] br[102] wl[348] vdd gnd cell_6t
Xbit_r349_c102 bl[102] br[102] wl[349] vdd gnd cell_6t
Xbit_r350_c102 bl[102] br[102] wl[350] vdd gnd cell_6t
Xbit_r351_c102 bl[102] br[102] wl[351] vdd gnd cell_6t
Xbit_r352_c102 bl[102] br[102] wl[352] vdd gnd cell_6t
Xbit_r353_c102 bl[102] br[102] wl[353] vdd gnd cell_6t
Xbit_r354_c102 bl[102] br[102] wl[354] vdd gnd cell_6t
Xbit_r355_c102 bl[102] br[102] wl[355] vdd gnd cell_6t
Xbit_r356_c102 bl[102] br[102] wl[356] vdd gnd cell_6t
Xbit_r357_c102 bl[102] br[102] wl[357] vdd gnd cell_6t
Xbit_r358_c102 bl[102] br[102] wl[358] vdd gnd cell_6t
Xbit_r359_c102 bl[102] br[102] wl[359] vdd gnd cell_6t
Xbit_r360_c102 bl[102] br[102] wl[360] vdd gnd cell_6t
Xbit_r361_c102 bl[102] br[102] wl[361] vdd gnd cell_6t
Xbit_r362_c102 bl[102] br[102] wl[362] vdd gnd cell_6t
Xbit_r363_c102 bl[102] br[102] wl[363] vdd gnd cell_6t
Xbit_r364_c102 bl[102] br[102] wl[364] vdd gnd cell_6t
Xbit_r365_c102 bl[102] br[102] wl[365] vdd gnd cell_6t
Xbit_r366_c102 bl[102] br[102] wl[366] vdd gnd cell_6t
Xbit_r367_c102 bl[102] br[102] wl[367] vdd gnd cell_6t
Xbit_r368_c102 bl[102] br[102] wl[368] vdd gnd cell_6t
Xbit_r369_c102 bl[102] br[102] wl[369] vdd gnd cell_6t
Xbit_r370_c102 bl[102] br[102] wl[370] vdd gnd cell_6t
Xbit_r371_c102 bl[102] br[102] wl[371] vdd gnd cell_6t
Xbit_r372_c102 bl[102] br[102] wl[372] vdd gnd cell_6t
Xbit_r373_c102 bl[102] br[102] wl[373] vdd gnd cell_6t
Xbit_r374_c102 bl[102] br[102] wl[374] vdd gnd cell_6t
Xbit_r375_c102 bl[102] br[102] wl[375] vdd gnd cell_6t
Xbit_r376_c102 bl[102] br[102] wl[376] vdd gnd cell_6t
Xbit_r377_c102 bl[102] br[102] wl[377] vdd gnd cell_6t
Xbit_r378_c102 bl[102] br[102] wl[378] vdd gnd cell_6t
Xbit_r379_c102 bl[102] br[102] wl[379] vdd gnd cell_6t
Xbit_r380_c102 bl[102] br[102] wl[380] vdd gnd cell_6t
Xbit_r381_c102 bl[102] br[102] wl[381] vdd gnd cell_6t
Xbit_r382_c102 bl[102] br[102] wl[382] vdd gnd cell_6t
Xbit_r383_c102 bl[102] br[102] wl[383] vdd gnd cell_6t
Xbit_r384_c102 bl[102] br[102] wl[384] vdd gnd cell_6t
Xbit_r385_c102 bl[102] br[102] wl[385] vdd gnd cell_6t
Xbit_r386_c102 bl[102] br[102] wl[386] vdd gnd cell_6t
Xbit_r387_c102 bl[102] br[102] wl[387] vdd gnd cell_6t
Xbit_r388_c102 bl[102] br[102] wl[388] vdd gnd cell_6t
Xbit_r389_c102 bl[102] br[102] wl[389] vdd gnd cell_6t
Xbit_r390_c102 bl[102] br[102] wl[390] vdd gnd cell_6t
Xbit_r391_c102 bl[102] br[102] wl[391] vdd gnd cell_6t
Xbit_r392_c102 bl[102] br[102] wl[392] vdd gnd cell_6t
Xbit_r393_c102 bl[102] br[102] wl[393] vdd gnd cell_6t
Xbit_r394_c102 bl[102] br[102] wl[394] vdd gnd cell_6t
Xbit_r395_c102 bl[102] br[102] wl[395] vdd gnd cell_6t
Xbit_r396_c102 bl[102] br[102] wl[396] vdd gnd cell_6t
Xbit_r397_c102 bl[102] br[102] wl[397] vdd gnd cell_6t
Xbit_r398_c102 bl[102] br[102] wl[398] vdd gnd cell_6t
Xbit_r399_c102 bl[102] br[102] wl[399] vdd gnd cell_6t
Xbit_r400_c102 bl[102] br[102] wl[400] vdd gnd cell_6t
Xbit_r401_c102 bl[102] br[102] wl[401] vdd gnd cell_6t
Xbit_r402_c102 bl[102] br[102] wl[402] vdd gnd cell_6t
Xbit_r403_c102 bl[102] br[102] wl[403] vdd gnd cell_6t
Xbit_r404_c102 bl[102] br[102] wl[404] vdd gnd cell_6t
Xbit_r405_c102 bl[102] br[102] wl[405] vdd gnd cell_6t
Xbit_r406_c102 bl[102] br[102] wl[406] vdd gnd cell_6t
Xbit_r407_c102 bl[102] br[102] wl[407] vdd gnd cell_6t
Xbit_r408_c102 bl[102] br[102] wl[408] vdd gnd cell_6t
Xbit_r409_c102 bl[102] br[102] wl[409] vdd gnd cell_6t
Xbit_r410_c102 bl[102] br[102] wl[410] vdd gnd cell_6t
Xbit_r411_c102 bl[102] br[102] wl[411] vdd gnd cell_6t
Xbit_r412_c102 bl[102] br[102] wl[412] vdd gnd cell_6t
Xbit_r413_c102 bl[102] br[102] wl[413] vdd gnd cell_6t
Xbit_r414_c102 bl[102] br[102] wl[414] vdd gnd cell_6t
Xbit_r415_c102 bl[102] br[102] wl[415] vdd gnd cell_6t
Xbit_r416_c102 bl[102] br[102] wl[416] vdd gnd cell_6t
Xbit_r417_c102 bl[102] br[102] wl[417] vdd gnd cell_6t
Xbit_r418_c102 bl[102] br[102] wl[418] vdd gnd cell_6t
Xbit_r419_c102 bl[102] br[102] wl[419] vdd gnd cell_6t
Xbit_r420_c102 bl[102] br[102] wl[420] vdd gnd cell_6t
Xbit_r421_c102 bl[102] br[102] wl[421] vdd gnd cell_6t
Xbit_r422_c102 bl[102] br[102] wl[422] vdd gnd cell_6t
Xbit_r423_c102 bl[102] br[102] wl[423] vdd gnd cell_6t
Xbit_r424_c102 bl[102] br[102] wl[424] vdd gnd cell_6t
Xbit_r425_c102 bl[102] br[102] wl[425] vdd gnd cell_6t
Xbit_r426_c102 bl[102] br[102] wl[426] vdd gnd cell_6t
Xbit_r427_c102 bl[102] br[102] wl[427] vdd gnd cell_6t
Xbit_r428_c102 bl[102] br[102] wl[428] vdd gnd cell_6t
Xbit_r429_c102 bl[102] br[102] wl[429] vdd gnd cell_6t
Xbit_r430_c102 bl[102] br[102] wl[430] vdd gnd cell_6t
Xbit_r431_c102 bl[102] br[102] wl[431] vdd gnd cell_6t
Xbit_r432_c102 bl[102] br[102] wl[432] vdd gnd cell_6t
Xbit_r433_c102 bl[102] br[102] wl[433] vdd gnd cell_6t
Xbit_r434_c102 bl[102] br[102] wl[434] vdd gnd cell_6t
Xbit_r435_c102 bl[102] br[102] wl[435] vdd gnd cell_6t
Xbit_r436_c102 bl[102] br[102] wl[436] vdd gnd cell_6t
Xbit_r437_c102 bl[102] br[102] wl[437] vdd gnd cell_6t
Xbit_r438_c102 bl[102] br[102] wl[438] vdd gnd cell_6t
Xbit_r439_c102 bl[102] br[102] wl[439] vdd gnd cell_6t
Xbit_r440_c102 bl[102] br[102] wl[440] vdd gnd cell_6t
Xbit_r441_c102 bl[102] br[102] wl[441] vdd gnd cell_6t
Xbit_r442_c102 bl[102] br[102] wl[442] vdd gnd cell_6t
Xbit_r443_c102 bl[102] br[102] wl[443] vdd gnd cell_6t
Xbit_r444_c102 bl[102] br[102] wl[444] vdd gnd cell_6t
Xbit_r445_c102 bl[102] br[102] wl[445] vdd gnd cell_6t
Xbit_r446_c102 bl[102] br[102] wl[446] vdd gnd cell_6t
Xbit_r447_c102 bl[102] br[102] wl[447] vdd gnd cell_6t
Xbit_r448_c102 bl[102] br[102] wl[448] vdd gnd cell_6t
Xbit_r449_c102 bl[102] br[102] wl[449] vdd gnd cell_6t
Xbit_r450_c102 bl[102] br[102] wl[450] vdd gnd cell_6t
Xbit_r451_c102 bl[102] br[102] wl[451] vdd gnd cell_6t
Xbit_r452_c102 bl[102] br[102] wl[452] vdd gnd cell_6t
Xbit_r453_c102 bl[102] br[102] wl[453] vdd gnd cell_6t
Xbit_r454_c102 bl[102] br[102] wl[454] vdd gnd cell_6t
Xbit_r455_c102 bl[102] br[102] wl[455] vdd gnd cell_6t
Xbit_r456_c102 bl[102] br[102] wl[456] vdd gnd cell_6t
Xbit_r457_c102 bl[102] br[102] wl[457] vdd gnd cell_6t
Xbit_r458_c102 bl[102] br[102] wl[458] vdd gnd cell_6t
Xbit_r459_c102 bl[102] br[102] wl[459] vdd gnd cell_6t
Xbit_r460_c102 bl[102] br[102] wl[460] vdd gnd cell_6t
Xbit_r461_c102 bl[102] br[102] wl[461] vdd gnd cell_6t
Xbit_r462_c102 bl[102] br[102] wl[462] vdd gnd cell_6t
Xbit_r463_c102 bl[102] br[102] wl[463] vdd gnd cell_6t
Xbit_r464_c102 bl[102] br[102] wl[464] vdd gnd cell_6t
Xbit_r465_c102 bl[102] br[102] wl[465] vdd gnd cell_6t
Xbit_r466_c102 bl[102] br[102] wl[466] vdd gnd cell_6t
Xbit_r467_c102 bl[102] br[102] wl[467] vdd gnd cell_6t
Xbit_r468_c102 bl[102] br[102] wl[468] vdd gnd cell_6t
Xbit_r469_c102 bl[102] br[102] wl[469] vdd gnd cell_6t
Xbit_r470_c102 bl[102] br[102] wl[470] vdd gnd cell_6t
Xbit_r471_c102 bl[102] br[102] wl[471] vdd gnd cell_6t
Xbit_r472_c102 bl[102] br[102] wl[472] vdd gnd cell_6t
Xbit_r473_c102 bl[102] br[102] wl[473] vdd gnd cell_6t
Xbit_r474_c102 bl[102] br[102] wl[474] vdd gnd cell_6t
Xbit_r475_c102 bl[102] br[102] wl[475] vdd gnd cell_6t
Xbit_r476_c102 bl[102] br[102] wl[476] vdd gnd cell_6t
Xbit_r477_c102 bl[102] br[102] wl[477] vdd gnd cell_6t
Xbit_r478_c102 bl[102] br[102] wl[478] vdd gnd cell_6t
Xbit_r479_c102 bl[102] br[102] wl[479] vdd gnd cell_6t
Xbit_r480_c102 bl[102] br[102] wl[480] vdd gnd cell_6t
Xbit_r481_c102 bl[102] br[102] wl[481] vdd gnd cell_6t
Xbit_r482_c102 bl[102] br[102] wl[482] vdd gnd cell_6t
Xbit_r483_c102 bl[102] br[102] wl[483] vdd gnd cell_6t
Xbit_r484_c102 bl[102] br[102] wl[484] vdd gnd cell_6t
Xbit_r485_c102 bl[102] br[102] wl[485] vdd gnd cell_6t
Xbit_r486_c102 bl[102] br[102] wl[486] vdd gnd cell_6t
Xbit_r487_c102 bl[102] br[102] wl[487] vdd gnd cell_6t
Xbit_r488_c102 bl[102] br[102] wl[488] vdd gnd cell_6t
Xbit_r489_c102 bl[102] br[102] wl[489] vdd gnd cell_6t
Xbit_r490_c102 bl[102] br[102] wl[490] vdd gnd cell_6t
Xbit_r491_c102 bl[102] br[102] wl[491] vdd gnd cell_6t
Xbit_r492_c102 bl[102] br[102] wl[492] vdd gnd cell_6t
Xbit_r493_c102 bl[102] br[102] wl[493] vdd gnd cell_6t
Xbit_r494_c102 bl[102] br[102] wl[494] vdd gnd cell_6t
Xbit_r495_c102 bl[102] br[102] wl[495] vdd gnd cell_6t
Xbit_r496_c102 bl[102] br[102] wl[496] vdd gnd cell_6t
Xbit_r497_c102 bl[102] br[102] wl[497] vdd gnd cell_6t
Xbit_r498_c102 bl[102] br[102] wl[498] vdd gnd cell_6t
Xbit_r499_c102 bl[102] br[102] wl[499] vdd gnd cell_6t
Xbit_r500_c102 bl[102] br[102] wl[500] vdd gnd cell_6t
Xbit_r501_c102 bl[102] br[102] wl[501] vdd gnd cell_6t
Xbit_r502_c102 bl[102] br[102] wl[502] vdd gnd cell_6t
Xbit_r503_c102 bl[102] br[102] wl[503] vdd gnd cell_6t
Xbit_r504_c102 bl[102] br[102] wl[504] vdd gnd cell_6t
Xbit_r505_c102 bl[102] br[102] wl[505] vdd gnd cell_6t
Xbit_r506_c102 bl[102] br[102] wl[506] vdd gnd cell_6t
Xbit_r507_c102 bl[102] br[102] wl[507] vdd gnd cell_6t
Xbit_r508_c102 bl[102] br[102] wl[508] vdd gnd cell_6t
Xbit_r509_c102 bl[102] br[102] wl[509] vdd gnd cell_6t
Xbit_r510_c102 bl[102] br[102] wl[510] vdd gnd cell_6t
Xbit_r511_c102 bl[102] br[102] wl[511] vdd gnd cell_6t
Xbit_r0_c103 bl[103] br[103] wl[0] vdd gnd cell_6t
Xbit_r1_c103 bl[103] br[103] wl[1] vdd gnd cell_6t
Xbit_r2_c103 bl[103] br[103] wl[2] vdd gnd cell_6t
Xbit_r3_c103 bl[103] br[103] wl[3] vdd gnd cell_6t
Xbit_r4_c103 bl[103] br[103] wl[4] vdd gnd cell_6t
Xbit_r5_c103 bl[103] br[103] wl[5] vdd gnd cell_6t
Xbit_r6_c103 bl[103] br[103] wl[6] vdd gnd cell_6t
Xbit_r7_c103 bl[103] br[103] wl[7] vdd gnd cell_6t
Xbit_r8_c103 bl[103] br[103] wl[8] vdd gnd cell_6t
Xbit_r9_c103 bl[103] br[103] wl[9] vdd gnd cell_6t
Xbit_r10_c103 bl[103] br[103] wl[10] vdd gnd cell_6t
Xbit_r11_c103 bl[103] br[103] wl[11] vdd gnd cell_6t
Xbit_r12_c103 bl[103] br[103] wl[12] vdd gnd cell_6t
Xbit_r13_c103 bl[103] br[103] wl[13] vdd gnd cell_6t
Xbit_r14_c103 bl[103] br[103] wl[14] vdd gnd cell_6t
Xbit_r15_c103 bl[103] br[103] wl[15] vdd gnd cell_6t
Xbit_r16_c103 bl[103] br[103] wl[16] vdd gnd cell_6t
Xbit_r17_c103 bl[103] br[103] wl[17] vdd gnd cell_6t
Xbit_r18_c103 bl[103] br[103] wl[18] vdd gnd cell_6t
Xbit_r19_c103 bl[103] br[103] wl[19] vdd gnd cell_6t
Xbit_r20_c103 bl[103] br[103] wl[20] vdd gnd cell_6t
Xbit_r21_c103 bl[103] br[103] wl[21] vdd gnd cell_6t
Xbit_r22_c103 bl[103] br[103] wl[22] vdd gnd cell_6t
Xbit_r23_c103 bl[103] br[103] wl[23] vdd gnd cell_6t
Xbit_r24_c103 bl[103] br[103] wl[24] vdd gnd cell_6t
Xbit_r25_c103 bl[103] br[103] wl[25] vdd gnd cell_6t
Xbit_r26_c103 bl[103] br[103] wl[26] vdd gnd cell_6t
Xbit_r27_c103 bl[103] br[103] wl[27] vdd gnd cell_6t
Xbit_r28_c103 bl[103] br[103] wl[28] vdd gnd cell_6t
Xbit_r29_c103 bl[103] br[103] wl[29] vdd gnd cell_6t
Xbit_r30_c103 bl[103] br[103] wl[30] vdd gnd cell_6t
Xbit_r31_c103 bl[103] br[103] wl[31] vdd gnd cell_6t
Xbit_r32_c103 bl[103] br[103] wl[32] vdd gnd cell_6t
Xbit_r33_c103 bl[103] br[103] wl[33] vdd gnd cell_6t
Xbit_r34_c103 bl[103] br[103] wl[34] vdd gnd cell_6t
Xbit_r35_c103 bl[103] br[103] wl[35] vdd gnd cell_6t
Xbit_r36_c103 bl[103] br[103] wl[36] vdd gnd cell_6t
Xbit_r37_c103 bl[103] br[103] wl[37] vdd gnd cell_6t
Xbit_r38_c103 bl[103] br[103] wl[38] vdd gnd cell_6t
Xbit_r39_c103 bl[103] br[103] wl[39] vdd gnd cell_6t
Xbit_r40_c103 bl[103] br[103] wl[40] vdd gnd cell_6t
Xbit_r41_c103 bl[103] br[103] wl[41] vdd gnd cell_6t
Xbit_r42_c103 bl[103] br[103] wl[42] vdd gnd cell_6t
Xbit_r43_c103 bl[103] br[103] wl[43] vdd gnd cell_6t
Xbit_r44_c103 bl[103] br[103] wl[44] vdd gnd cell_6t
Xbit_r45_c103 bl[103] br[103] wl[45] vdd gnd cell_6t
Xbit_r46_c103 bl[103] br[103] wl[46] vdd gnd cell_6t
Xbit_r47_c103 bl[103] br[103] wl[47] vdd gnd cell_6t
Xbit_r48_c103 bl[103] br[103] wl[48] vdd gnd cell_6t
Xbit_r49_c103 bl[103] br[103] wl[49] vdd gnd cell_6t
Xbit_r50_c103 bl[103] br[103] wl[50] vdd gnd cell_6t
Xbit_r51_c103 bl[103] br[103] wl[51] vdd gnd cell_6t
Xbit_r52_c103 bl[103] br[103] wl[52] vdd gnd cell_6t
Xbit_r53_c103 bl[103] br[103] wl[53] vdd gnd cell_6t
Xbit_r54_c103 bl[103] br[103] wl[54] vdd gnd cell_6t
Xbit_r55_c103 bl[103] br[103] wl[55] vdd gnd cell_6t
Xbit_r56_c103 bl[103] br[103] wl[56] vdd gnd cell_6t
Xbit_r57_c103 bl[103] br[103] wl[57] vdd gnd cell_6t
Xbit_r58_c103 bl[103] br[103] wl[58] vdd gnd cell_6t
Xbit_r59_c103 bl[103] br[103] wl[59] vdd gnd cell_6t
Xbit_r60_c103 bl[103] br[103] wl[60] vdd gnd cell_6t
Xbit_r61_c103 bl[103] br[103] wl[61] vdd gnd cell_6t
Xbit_r62_c103 bl[103] br[103] wl[62] vdd gnd cell_6t
Xbit_r63_c103 bl[103] br[103] wl[63] vdd gnd cell_6t
Xbit_r64_c103 bl[103] br[103] wl[64] vdd gnd cell_6t
Xbit_r65_c103 bl[103] br[103] wl[65] vdd gnd cell_6t
Xbit_r66_c103 bl[103] br[103] wl[66] vdd gnd cell_6t
Xbit_r67_c103 bl[103] br[103] wl[67] vdd gnd cell_6t
Xbit_r68_c103 bl[103] br[103] wl[68] vdd gnd cell_6t
Xbit_r69_c103 bl[103] br[103] wl[69] vdd gnd cell_6t
Xbit_r70_c103 bl[103] br[103] wl[70] vdd gnd cell_6t
Xbit_r71_c103 bl[103] br[103] wl[71] vdd gnd cell_6t
Xbit_r72_c103 bl[103] br[103] wl[72] vdd gnd cell_6t
Xbit_r73_c103 bl[103] br[103] wl[73] vdd gnd cell_6t
Xbit_r74_c103 bl[103] br[103] wl[74] vdd gnd cell_6t
Xbit_r75_c103 bl[103] br[103] wl[75] vdd gnd cell_6t
Xbit_r76_c103 bl[103] br[103] wl[76] vdd gnd cell_6t
Xbit_r77_c103 bl[103] br[103] wl[77] vdd gnd cell_6t
Xbit_r78_c103 bl[103] br[103] wl[78] vdd gnd cell_6t
Xbit_r79_c103 bl[103] br[103] wl[79] vdd gnd cell_6t
Xbit_r80_c103 bl[103] br[103] wl[80] vdd gnd cell_6t
Xbit_r81_c103 bl[103] br[103] wl[81] vdd gnd cell_6t
Xbit_r82_c103 bl[103] br[103] wl[82] vdd gnd cell_6t
Xbit_r83_c103 bl[103] br[103] wl[83] vdd gnd cell_6t
Xbit_r84_c103 bl[103] br[103] wl[84] vdd gnd cell_6t
Xbit_r85_c103 bl[103] br[103] wl[85] vdd gnd cell_6t
Xbit_r86_c103 bl[103] br[103] wl[86] vdd gnd cell_6t
Xbit_r87_c103 bl[103] br[103] wl[87] vdd gnd cell_6t
Xbit_r88_c103 bl[103] br[103] wl[88] vdd gnd cell_6t
Xbit_r89_c103 bl[103] br[103] wl[89] vdd gnd cell_6t
Xbit_r90_c103 bl[103] br[103] wl[90] vdd gnd cell_6t
Xbit_r91_c103 bl[103] br[103] wl[91] vdd gnd cell_6t
Xbit_r92_c103 bl[103] br[103] wl[92] vdd gnd cell_6t
Xbit_r93_c103 bl[103] br[103] wl[93] vdd gnd cell_6t
Xbit_r94_c103 bl[103] br[103] wl[94] vdd gnd cell_6t
Xbit_r95_c103 bl[103] br[103] wl[95] vdd gnd cell_6t
Xbit_r96_c103 bl[103] br[103] wl[96] vdd gnd cell_6t
Xbit_r97_c103 bl[103] br[103] wl[97] vdd gnd cell_6t
Xbit_r98_c103 bl[103] br[103] wl[98] vdd gnd cell_6t
Xbit_r99_c103 bl[103] br[103] wl[99] vdd gnd cell_6t
Xbit_r100_c103 bl[103] br[103] wl[100] vdd gnd cell_6t
Xbit_r101_c103 bl[103] br[103] wl[101] vdd gnd cell_6t
Xbit_r102_c103 bl[103] br[103] wl[102] vdd gnd cell_6t
Xbit_r103_c103 bl[103] br[103] wl[103] vdd gnd cell_6t
Xbit_r104_c103 bl[103] br[103] wl[104] vdd gnd cell_6t
Xbit_r105_c103 bl[103] br[103] wl[105] vdd gnd cell_6t
Xbit_r106_c103 bl[103] br[103] wl[106] vdd gnd cell_6t
Xbit_r107_c103 bl[103] br[103] wl[107] vdd gnd cell_6t
Xbit_r108_c103 bl[103] br[103] wl[108] vdd gnd cell_6t
Xbit_r109_c103 bl[103] br[103] wl[109] vdd gnd cell_6t
Xbit_r110_c103 bl[103] br[103] wl[110] vdd gnd cell_6t
Xbit_r111_c103 bl[103] br[103] wl[111] vdd gnd cell_6t
Xbit_r112_c103 bl[103] br[103] wl[112] vdd gnd cell_6t
Xbit_r113_c103 bl[103] br[103] wl[113] vdd gnd cell_6t
Xbit_r114_c103 bl[103] br[103] wl[114] vdd gnd cell_6t
Xbit_r115_c103 bl[103] br[103] wl[115] vdd gnd cell_6t
Xbit_r116_c103 bl[103] br[103] wl[116] vdd gnd cell_6t
Xbit_r117_c103 bl[103] br[103] wl[117] vdd gnd cell_6t
Xbit_r118_c103 bl[103] br[103] wl[118] vdd gnd cell_6t
Xbit_r119_c103 bl[103] br[103] wl[119] vdd gnd cell_6t
Xbit_r120_c103 bl[103] br[103] wl[120] vdd gnd cell_6t
Xbit_r121_c103 bl[103] br[103] wl[121] vdd gnd cell_6t
Xbit_r122_c103 bl[103] br[103] wl[122] vdd gnd cell_6t
Xbit_r123_c103 bl[103] br[103] wl[123] vdd gnd cell_6t
Xbit_r124_c103 bl[103] br[103] wl[124] vdd gnd cell_6t
Xbit_r125_c103 bl[103] br[103] wl[125] vdd gnd cell_6t
Xbit_r126_c103 bl[103] br[103] wl[126] vdd gnd cell_6t
Xbit_r127_c103 bl[103] br[103] wl[127] vdd gnd cell_6t
Xbit_r128_c103 bl[103] br[103] wl[128] vdd gnd cell_6t
Xbit_r129_c103 bl[103] br[103] wl[129] vdd gnd cell_6t
Xbit_r130_c103 bl[103] br[103] wl[130] vdd gnd cell_6t
Xbit_r131_c103 bl[103] br[103] wl[131] vdd gnd cell_6t
Xbit_r132_c103 bl[103] br[103] wl[132] vdd gnd cell_6t
Xbit_r133_c103 bl[103] br[103] wl[133] vdd gnd cell_6t
Xbit_r134_c103 bl[103] br[103] wl[134] vdd gnd cell_6t
Xbit_r135_c103 bl[103] br[103] wl[135] vdd gnd cell_6t
Xbit_r136_c103 bl[103] br[103] wl[136] vdd gnd cell_6t
Xbit_r137_c103 bl[103] br[103] wl[137] vdd gnd cell_6t
Xbit_r138_c103 bl[103] br[103] wl[138] vdd gnd cell_6t
Xbit_r139_c103 bl[103] br[103] wl[139] vdd gnd cell_6t
Xbit_r140_c103 bl[103] br[103] wl[140] vdd gnd cell_6t
Xbit_r141_c103 bl[103] br[103] wl[141] vdd gnd cell_6t
Xbit_r142_c103 bl[103] br[103] wl[142] vdd gnd cell_6t
Xbit_r143_c103 bl[103] br[103] wl[143] vdd gnd cell_6t
Xbit_r144_c103 bl[103] br[103] wl[144] vdd gnd cell_6t
Xbit_r145_c103 bl[103] br[103] wl[145] vdd gnd cell_6t
Xbit_r146_c103 bl[103] br[103] wl[146] vdd gnd cell_6t
Xbit_r147_c103 bl[103] br[103] wl[147] vdd gnd cell_6t
Xbit_r148_c103 bl[103] br[103] wl[148] vdd gnd cell_6t
Xbit_r149_c103 bl[103] br[103] wl[149] vdd gnd cell_6t
Xbit_r150_c103 bl[103] br[103] wl[150] vdd gnd cell_6t
Xbit_r151_c103 bl[103] br[103] wl[151] vdd gnd cell_6t
Xbit_r152_c103 bl[103] br[103] wl[152] vdd gnd cell_6t
Xbit_r153_c103 bl[103] br[103] wl[153] vdd gnd cell_6t
Xbit_r154_c103 bl[103] br[103] wl[154] vdd gnd cell_6t
Xbit_r155_c103 bl[103] br[103] wl[155] vdd gnd cell_6t
Xbit_r156_c103 bl[103] br[103] wl[156] vdd gnd cell_6t
Xbit_r157_c103 bl[103] br[103] wl[157] vdd gnd cell_6t
Xbit_r158_c103 bl[103] br[103] wl[158] vdd gnd cell_6t
Xbit_r159_c103 bl[103] br[103] wl[159] vdd gnd cell_6t
Xbit_r160_c103 bl[103] br[103] wl[160] vdd gnd cell_6t
Xbit_r161_c103 bl[103] br[103] wl[161] vdd gnd cell_6t
Xbit_r162_c103 bl[103] br[103] wl[162] vdd gnd cell_6t
Xbit_r163_c103 bl[103] br[103] wl[163] vdd gnd cell_6t
Xbit_r164_c103 bl[103] br[103] wl[164] vdd gnd cell_6t
Xbit_r165_c103 bl[103] br[103] wl[165] vdd gnd cell_6t
Xbit_r166_c103 bl[103] br[103] wl[166] vdd gnd cell_6t
Xbit_r167_c103 bl[103] br[103] wl[167] vdd gnd cell_6t
Xbit_r168_c103 bl[103] br[103] wl[168] vdd gnd cell_6t
Xbit_r169_c103 bl[103] br[103] wl[169] vdd gnd cell_6t
Xbit_r170_c103 bl[103] br[103] wl[170] vdd gnd cell_6t
Xbit_r171_c103 bl[103] br[103] wl[171] vdd gnd cell_6t
Xbit_r172_c103 bl[103] br[103] wl[172] vdd gnd cell_6t
Xbit_r173_c103 bl[103] br[103] wl[173] vdd gnd cell_6t
Xbit_r174_c103 bl[103] br[103] wl[174] vdd gnd cell_6t
Xbit_r175_c103 bl[103] br[103] wl[175] vdd gnd cell_6t
Xbit_r176_c103 bl[103] br[103] wl[176] vdd gnd cell_6t
Xbit_r177_c103 bl[103] br[103] wl[177] vdd gnd cell_6t
Xbit_r178_c103 bl[103] br[103] wl[178] vdd gnd cell_6t
Xbit_r179_c103 bl[103] br[103] wl[179] vdd gnd cell_6t
Xbit_r180_c103 bl[103] br[103] wl[180] vdd gnd cell_6t
Xbit_r181_c103 bl[103] br[103] wl[181] vdd gnd cell_6t
Xbit_r182_c103 bl[103] br[103] wl[182] vdd gnd cell_6t
Xbit_r183_c103 bl[103] br[103] wl[183] vdd gnd cell_6t
Xbit_r184_c103 bl[103] br[103] wl[184] vdd gnd cell_6t
Xbit_r185_c103 bl[103] br[103] wl[185] vdd gnd cell_6t
Xbit_r186_c103 bl[103] br[103] wl[186] vdd gnd cell_6t
Xbit_r187_c103 bl[103] br[103] wl[187] vdd gnd cell_6t
Xbit_r188_c103 bl[103] br[103] wl[188] vdd gnd cell_6t
Xbit_r189_c103 bl[103] br[103] wl[189] vdd gnd cell_6t
Xbit_r190_c103 bl[103] br[103] wl[190] vdd gnd cell_6t
Xbit_r191_c103 bl[103] br[103] wl[191] vdd gnd cell_6t
Xbit_r192_c103 bl[103] br[103] wl[192] vdd gnd cell_6t
Xbit_r193_c103 bl[103] br[103] wl[193] vdd gnd cell_6t
Xbit_r194_c103 bl[103] br[103] wl[194] vdd gnd cell_6t
Xbit_r195_c103 bl[103] br[103] wl[195] vdd gnd cell_6t
Xbit_r196_c103 bl[103] br[103] wl[196] vdd gnd cell_6t
Xbit_r197_c103 bl[103] br[103] wl[197] vdd gnd cell_6t
Xbit_r198_c103 bl[103] br[103] wl[198] vdd gnd cell_6t
Xbit_r199_c103 bl[103] br[103] wl[199] vdd gnd cell_6t
Xbit_r200_c103 bl[103] br[103] wl[200] vdd gnd cell_6t
Xbit_r201_c103 bl[103] br[103] wl[201] vdd gnd cell_6t
Xbit_r202_c103 bl[103] br[103] wl[202] vdd gnd cell_6t
Xbit_r203_c103 bl[103] br[103] wl[203] vdd gnd cell_6t
Xbit_r204_c103 bl[103] br[103] wl[204] vdd gnd cell_6t
Xbit_r205_c103 bl[103] br[103] wl[205] vdd gnd cell_6t
Xbit_r206_c103 bl[103] br[103] wl[206] vdd gnd cell_6t
Xbit_r207_c103 bl[103] br[103] wl[207] vdd gnd cell_6t
Xbit_r208_c103 bl[103] br[103] wl[208] vdd gnd cell_6t
Xbit_r209_c103 bl[103] br[103] wl[209] vdd gnd cell_6t
Xbit_r210_c103 bl[103] br[103] wl[210] vdd gnd cell_6t
Xbit_r211_c103 bl[103] br[103] wl[211] vdd gnd cell_6t
Xbit_r212_c103 bl[103] br[103] wl[212] vdd gnd cell_6t
Xbit_r213_c103 bl[103] br[103] wl[213] vdd gnd cell_6t
Xbit_r214_c103 bl[103] br[103] wl[214] vdd gnd cell_6t
Xbit_r215_c103 bl[103] br[103] wl[215] vdd gnd cell_6t
Xbit_r216_c103 bl[103] br[103] wl[216] vdd gnd cell_6t
Xbit_r217_c103 bl[103] br[103] wl[217] vdd gnd cell_6t
Xbit_r218_c103 bl[103] br[103] wl[218] vdd gnd cell_6t
Xbit_r219_c103 bl[103] br[103] wl[219] vdd gnd cell_6t
Xbit_r220_c103 bl[103] br[103] wl[220] vdd gnd cell_6t
Xbit_r221_c103 bl[103] br[103] wl[221] vdd gnd cell_6t
Xbit_r222_c103 bl[103] br[103] wl[222] vdd gnd cell_6t
Xbit_r223_c103 bl[103] br[103] wl[223] vdd gnd cell_6t
Xbit_r224_c103 bl[103] br[103] wl[224] vdd gnd cell_6t
Xbit_r225_c103 bl[103] br[103] wl[225] vdd gnd cell_6t
Xbit_r226_c103 bl[103] br[103] wl[226] vdd gnd cell_6t
Xbit_r227_c103 bl[103] br[103] wl[227] vdd gnd cell_6t
Xbit_r228_c103 bl[103] br[103] wl[228] vdd gnd cell_6t
Xbit_r229_c103 bl[103] br[103] wl[229] vdd gnd cell_6t
Xbit_r230_c103 bl[103] br[103] wl[230] vdd gnd cell_6t
Xbit_r231_c103 bl[103] br[103] wl[231] vdd gnd cell_6t
Xbit_r232_c103 bl[103] br[103] wl[232] vdd gnd cell_6t
Xbit_r233_c103 bl[103] br[103] wl[233] vdd gnd cell_6t
Xbit_r234_c103 bl[103] br[103] wl[234] vdd gnd cell_6t
Xbit_r235_c103 bl[103] br[103] wl[235] vdd gnd cell_6t
Xbit_r236_c103 bl[103] br[103] wl[236] vdd gnd cell_6t
Xbit_r237_c103 bl[103] br[103] wl[237] vdd gnd cell_6t
Xbit_r238_c103 bl[103] br[103] wl[238] vdd gnd cell_6t
Xbit_r239_c103 bl[103] br[103] wl[239] vdd gnd cell_6t
Xbit_r240_c103 bl[103] br[103] wl[240] vdd gnd cell_6t
Xbit_r241_c103 bl[103] br[103] wl[241] vdd gnd cell_6t
Xbit_r242_c103 bl[103] br[103] wl[242] vdd gnd cell_6t
Xbit_r243_c103 bl[103] br[103] wl[243] vdd gnd cell_6t
Xbit_r244_c103 bl[103] br[103] wl[244] vdd gnd cell_6t
Xbit_r245_c103 bl[103] br[103] wl[245] vdd gnd cell_6t
Xbit_r246_c103 bl[103] br[103] wl[246] vdd gnd cell_6t
Xbit_r247_c103 bl[103] br[103] wl[247] vdd gnd cell_6t
Xbit_r248_c103 bl[103] br[103] wl[248] vdd gnd cell_6t
Xbit_r249_c103 bl[103] br[103] wl[249] vdd gnd cell_6t
Xbit_r250_c103 bl[103] br[103] wl[250] vdd gnd cell_6t
Xbit_r251_c103 bl[103] br[103] wl[251] vdd gnd cell_6t
Xbit_r252_c103 bl[103] br[103] wl[252] vdd gnd cell_6t
Xbit_r253_c103 bl[103] br[103] wl[253] vdd gnd cell_6t
Xbit_r254_c103 bl[103] br[103] wl[254] vdd gnd cell_6t
Xbit_r255_c103 bl[103] br[103] wl[255] vdd gnd cell_6t
Xbit_r256_c103 bl[103] br[103] wl[256] vdd gnd cell_6t
Xbit_r257_c103 bl[103] br[103] wl[257] vdd gnd cell_6t
Xbit_r258_c103 bl[103] br[103] wl[258] vdd gnd cell_6t
Xbit_r259_c103 bl[103] br[103] wl[259] vdd gnd cell_6t
Xbit_r260_c103 bl[103] br[103] wl[260] vdd gnd cell_6t
Xbit_r261_c103 bl[103] br[103] wl[261] vdd gnd cell_6t
Xbit_r262_c103 bl[103] br[103] wl[262] vdd gnd cell_6t
Xbit_r263_c103 bl[103] br[103] wl[263] vdd gnd cell_6t
Xbit_r264_c103 bl[103] br[103] wl[264] vdd gnd cell_6t
Xbit_r265_c103 bl[103] br[103] wl[265] vdd gnd cell_6t
Xbit_r266_c103 bl[103] br[103] wl[266] vdd gnd cell_6t
Xbit_r267_c103 bl[103] br[103] wl[267] vdd gnd cell_6t
Xbit_r268_c103 bl[103] br[103] wl[268] vdd gnd cell_6t
Xbit_r269_c103 bl[103] br[103] wl[269] vdd gnd cell_6t
Xbit_r270_c103 bl[103] br[103] wl[270] vdd gnd cell_6t
Xbit_r271_c103 bl[103] br[103] wl[271] vdd gnd cell_6t
Xbit_r272_c103 bl[103] br[103] wl[272] vdd gnd cell_6t
Xbit_r273_c103 bl[103] br[103] wl[273] vdd gnd cell_6t
Xbit_r274_c103 bl[103] br[103] wl[274] vdd gnd cell_6t
Xbit_r275_c103 bl[103] br[103] wl[275] vdd gnd cell_6t
Xbit_r276_c103 bl[103] br[103] wl[276] vdd gnd cell_6t
Xbit_r277_c103 bl[103] br[103] wl[277] vdd gnd cell_6t
Xbit_r278_c103 bl[103] br[103] wl[278] vdd gnd cell_6t
Xbit_r279_c103 bl[103] br[103] wl[279] vdd gnd cell_6t
Xbit_r280_c103 bl[103] br[103] wl[280] vdd gnd cell_6t
Xbit_r281_c103 bl[103] br[103] wl[281] vdd gnd cell_6t
Xbit_r282_c103 bl[103] br[103] wl[282] vdd gnd cell_6t
Xbit_r283_c103 bl[103] br[103] wl[283] vdd gnd cell_6t
Xbit_r284_c103 bl[103] br[103] wl[284] vdd gnd cell_6t
Xbit_r285_c103 bl[103] br[103] wl[285] vdd gnd cell_6t
Xbit_r286_c103 bl[103] br[103] wl[286] vdd gnd cell_6t
Xbit_r287_c103 bl[103] br[103] wl[287] vdd gnd cell_6t
Xbit_r288_c103 bl[103] br[103] wl[288] vdd gnd cell_6t
Xbit_r289_c103 bl[103] br[103] wl[289] vdd gnd cell_6t
Xbit_r290_c103 bl[103] br[103] wl[290] vdd gnd cell_6t
Xbit_r291_c103 bl[103] br[103] wl[291] vdd gnd cell_6t
Xbit_r292_c103 bl[103] br[103] wl[292] vdd gnd cell_6t
Xbit_r293_c103 bl[103] br[103] wl[293] vdd gnd cell_6t
Xbit_r294_c103 bl[103] br[103] wl[294] vdd gnd cell_6t
Xbit_r295_c103 bl[103] br[103] wl[295] vdd gnd cell_6t
Xbit_r296_c103 bl[103] br[103] wl[296] vdd gnd cell_6t
Xbit_r297_c103 bl[103] br[103] wl[297] vdd gnd cell_6t
Xbit_r298_c103 bl[103] br[103] wl[298] vdd gnd cell_6t
Xbit_r299_c103 bl[103] br[103] wl[299] vdd gnd cell_6t
Xbit_r300_c103 bl[103] br[103] wl[300] vdd gnd cell_6t
Xbit_r301_c103 bl[103] br[103] wl[301] vdd gnd cell_6t
Xbit_r302_c103 bl[103] br[103] wl[302] vdd gnd cell_6t
Xbit_r303_c103 bl[103] br[103] wl[303] vdd gnd cell_6t
Xbit_r304_c103 bl[103] br[103] wl[304] vdd gnd cell_6t
Xbit_r305_c103 bl[103] br[103] wl[305] vdd gnd cell_6t
Xbit_r306_c103 bl[103] br[103] wl[306] vdd gnd cell_6t
Xbit_r307_c103 bl[103] br[103] wl[307] vdd gnd cell_6t
Xbit_r308_c103 bl[103] br[103] wl[308] vdd gnd cell_6t
Xbit_r309_c103 bl[103] br[103] wl[309] vdd gnd cell_6t
Xbit_r310_c103 bl[103] br[103] wl[310] vdd gnd cell_6t
Xbit_r311_c103 bl[103] br[103] wl[311] vdd gnd cell_6t
Xbit_r312_c103 bl[103] br[103] wl[312] vdd gnd cell_6t
Xbit_r313_c103 bl[103] br[103] wl[313] vdd gnd cell_6t
Xbit_r314_c103 bl[103] br[103] wl[314] vdd gnd cell_6t
Xbit_r315_c103 bl[103] br[103] wl[315] vdd gnd cell_6t
Xbit_r316_c103 bl[103] br[103] wl[316] vdd gnd cell_6t
Xbit_r317_c103 bl[103] br[103] wl[317] vdd gnd cell_6t
Xbit_r318_c103 bl[103] br[103] wl[318] vdd gnd cell_6t
Xbit_r319_c103 bl[103] br[103] wl[319] vdd gnd cell_6t
Xbit_r320_c103 bl[103] br[103] wl[320] vdd gnd cell_6t
Xbit_r321_c103 bl[103] br[103] wl[321] vdd gnd cell_6t
Xbit_r322_c103 bl[103] br[103] wl[322] vdd gnd cell_6t
Xbit_r323_c103 bl[103] br[103] wl[323] vdd gnd cell_6t
Xbit_r324_c103 bl[103] br[103] wl[324] vdd gnd cell_6t
Xbit_r325_c103 bl[103] br[103] wl[325] vdd gnd cell_6t
Xbit_r326_c103 bl[103] br[103] wl[326] vdd gnd cell_6t
Xbit_r327_c103 bl[103] br[103] wl[327] vdd gnd cell_6t
Xbit_r328_c103 bl[103] br[103] wl[328] vdd gnd cell_6t
Xbit_r329_c103 bl[103] br[103] wl[329] vdd gnd cell_6t
Xbit_r330_c103 bl[103] br[103] wl[330] vdd gnd cell_6t
Xbit_r331_c103 bl[103] br[103] wl[331] vdd gnd cell_6t
Xbit_r332_c103 bl[103] br[103] wl[332] vdd gnd cell_6t
Xbit_r333_c103 bl[103] br[103] wl[333] vdd gnd cell_6t
Xbit_r334_c103 bl[103] br[103] wl[334] vdd gnd cell_6t
Xbit_r335_c103 bl[103] br[103] wl[335] vdd gnd cell_6t
Xbit_r336_c103 bl[103] br[103] wl[336] vdd gnd cell_6t
Xbit_r337_c103 bl[103] br[103] wl[337] vdd gnd cell_6t
Xbit_r338_c103 bl[103] br[103] wl[338] vdd gnd cell_6t
Xbit_r339_c103 bl[103] br[103] wl[339] vdd gnd cell_6t
Xbit_r340_c103 bl[103] br[103] wl[340] vdd gnd cell_6t
Xbit_r341_c103 bl[103] br[103] wl[341] vdd gnd cell_6t
Xbit_r342_c103 bl[103] br[103] wl[342] vdd gnd cell_6t
Xbit_r343_c103 bl[103] br[103] wl[343] vdd gnd cell_6t
Xbit_r344_c103 bl[103] br[103] wl[344] vdd gnd cell_6t
Xbit_r345_c103 bl[103] br[103] wl[345] vdd gnd cell_6t
Xbit_r346_c103 bl[103] br[103] wl[346] vdd gnd cell_6t
Xbit_r347_c103 bl[103] br[103] wl[347] vdd gnd cell_6t
Xbit_r348_c103 bl[103] br[103] wl[348] vdd gnd cell_6t
Xbit_r349_c103 bl[103] br[103] wl[349] vdd gnd cell_6t
Xbit_r350_c103 bl[103] br[103] wl[350] vdd gnd cell_6t
Xbit_r351_c103 bl[103] br[103] wl[351] vdd gnd cell_6t
Xbit_r352_c103 bl[103] br[103] wl[352] vdd gnd cell_6t
Xbit_r353_c103 bl[103] br[103] wl[353] vdd gnd cell_6t
Xbit_r354_c103 bl[103] br[103] wl[354] vdd gnd cell_6t
Xbit_r355_c103 bl[103] br[103] wl[355] vdd gnd cell_6t
Xbit_r356_c103 bl[103] br[103] wl[356] vdd gnd cell_6t
Xbit_r357_c103 bl[103] br[103] wl[357] vdd gnd cell_6t
Xbit_r358_c103 bl[103] br[103] wl[358] vdd gnd cell_6t
Xbit_r359_c103 bl[103] br[103] wl[359] vdd gnd cell_6t
Xbit_r360_c103 bl[103] br[103] wl[360] vdd gnd cell_6t
Xbit_r361_c103 bl[103] br[103] wl[361] vdd gnd cell_6t
Xbit_r362_c103 bl[103] br[103] wl[362] vdd gnd cell_6t
Xbit_r363_c103 bl[103] br[103] wl[363] vdd gnd cell_6t
Xbit_r364_c103 bl[103] br[103] wl[364] vdd gnd cell_6t
Xbit_r365_c103 bl[103] br[103] wl[365] vdd gnd cell_6t
Xbit_r366_c103 bl[103] br[103] wl[366] vdd gnd cell_6t
Xbit_r367_c103 bl[103] br[103] wl[367] vdd gnd cell_6t
Xbit_r368_c103 bl[103] br[103] wl[368] vdd gnd cell_6t
Xbit_r369_c103 bl[103] br[103] wl[369] vdd gnd cell_6t
Xbit_r370_c103 bl[103] br[103] wl[370] vdd gnd cell_6t
Xbit_r371_c103 bl[103] br[103] wl[371] vdd gnd cell_6t
Xbit_r372_c103 bl[103] br[103] wl[372] vdd gnd cell_6t
Xbit_r373_c103 bl[103] br[103] wl[373] vdd gnd cell_6t
Xbit_r374_c103 bl[103] br[103] wl[374] vdd gnd cell_6t
Xbit_r375_c103 bl[103] br[103] wl[375] vdd gnd cell_6t
Xbit_r376_c103 bl[103] br[103] wl[376] vdd gnd cell_6t
Xbit_r377_c103 bl[103] br[103] wl[377] vdd gnd cell_6t
Xbit_r378_c103 bl[103] br[103] wl[378] vdd gnd cell_6t
Xbit_r379_c103 bl[103] br[103] wl[379] vdd gnd cell_6t
Xbit_r380_c103 bl[103] br[103] wl[380] vdd gnd cell_6t
Xbit_r381_c103 bl[103] br[103] wl[381] vdd gnd cell_6t
Xbit_r382_c103 bl[103] br[103] wl[382] vdd gnd cell_6t
Xbit_r383_c103 bl[103] br[103] wl[383] vdd gnd cell_6t
Xbit_r384_c103 bl[103] br[103] wl[384] vdd gnd cell_6t
Xbit_r385_c103 bl[103] br[103] wl[385] vdd gnd cell_6t
Xbit_r386_c103 bl[103] br[103] wl[386] vdd gnd cell_6t
Xbit_r387_c103 bl[103] br[103] wl[387] vdd gnd cell_6t
Xbit_r388_c103 bl[103] br[103] wl[388] vdd gnd cell_6t
Xbit_r389_c103 bl[103] br[103] wl[389] vdd gnd cell_6t
Xbit_r390_c103 bl[103] br[103] wl[390] vdd gnd cell_6t
Xbit_r391_c103 bl[103] br[103] wl[391] vdd gnd cell_6t
Xbit_r392_c103 bl[103] br[103] wl[392] vdd gnd cell_6t
Xbit_r393_c103 bl[103] br[103] wl[393] vdd gnd cell_6t
Xbit_r394_c103 bl[103] br[103] wl[394] vdd gnd cell_6t
Xbit_r395_c103 bl[103] br[103] wl[395] vdd gnd cell_6t
Xbit_r396_c103 bl[103] br[103] wl[396] vdd gnd cell_6t
Xbit_r397_c103 bl[103] br[103] wl[397] vdd gnd cell_6t
Xbit_r398_c103 bl[103] br[103] wl[398] vdd gnd cell_6t
Xbit_r399_c103 bl[103] br[103] wl[399] vdd gnd cell_6t
Xbit_r400_c103 bl[103] br[103] wl[400] vdd gnd cell_6t
Xbit_r401_c103 bl[103] br[103] wl[401] vdd gnd cell_6t
Xbit_r402_c103 bl[103] br[103] wl[402] vdd gnd cell_6t
Xbit_r403_c103 bl[103] br[103] wl[403] vdd gnd cell_6t
Xbit_r404_c103 bl[103] br[103] wl[404] vdd gnd cell_6t
Xbit_r405_c103 bl[103] br[103] wl[405] vdd gnd cell_6t
Xbit_r406_c103 bl[103] br[103] wl[406] vdd gnd cell_6t
Xbit_r407_c103 bl[103] br[103] wl[407] vdd gnd cell_6t
Xbit_r408_c103 bl[103] br[103] wl[408] vdd gnd cell_6t
Xbit_r409_c103 bl[103] br[103] wl[409] vdd gnd cell_6t
Xbit_r410_c103 bl[103] br[103] wl[410] vdd gnd cell_6t
Xbit_r411_c103 bl[103] br[103] wl[411] vdd gnd cell_6t
Xbit_r412_c103 bl[103] br[103] wl[412] vdd gnd cell_6t
Xbit_r413_c103 bl[103] br[103] wl[413] vdd gnd cell_6t
Xbit_r414_c103 bl[103] br[103] wl[414] vdd gnd cell_6t
Xbit_r415_c103 bl[103] br[103] wl[415] vdd gnd cell_6t
Xbit_r416_c103 bl[103] br[103] wl[416] vdd gnd cell_6t
Xbit_r417_c103 bl[103] br[103] wl[417] vdd gnd cell_6t
Xbit_r418_c103 bl[103] br[103] wl[418] vdd gnd cell_6t
Xbit_r419_c103 bl[103] br[103] wl[419] vdd gnd cell_6t
Xbit_r420_c103 bl[103] br[103] wl[420] vdd gnd cell_6t
Xbit_r421_c103 bl[103] br[103] wl[421] vdd gnd cell_6t
Xbit_r422_c103 bl[103] br[103] wl[422] vdd gnd cell_6t
Xbit_r423_c103 bl[103] br[103] wl[423] vdd gnd cell_6t
Xbit_r424_c103 bl[103] br[103] wl[424] vdd gnd cell_6t
Xbit_r425_c103 bl[103] br[103] wl[425] vdd gnd cell_6t
Xbit_r426_c103 bl[103] br[103] wl[426] vdd gnd cell_6t
Xbit_r427_c103 bl[103] br[103] wl[427] vdd gnd cell_6t
Xbit_r428_c103 bl[103] br[103] wl[428] vdd gnd cell_6t
Xbit_r429_c103 bl[103] br[103] wl[429] vdd gnd cell_6t
Xbit_r430_c103 bl[103] br[103] wl[430] vdd gnd cell_6t
Xbit_r431_c103 bl[103] br[103] wl[431] vdd gnd cell_6t
Xbit_r432_c103 bl[103] br[103] wl[432] vdd gnd cell_6t
Xbit_r433_c103 bl[103] br[103] wl[433] vdd gnd cell_6t
Xbit_r434_c103 bl[103] br[103] wl[434] vdd gnd cell_6t
Xbit_r435_c103 bl[103] br[103] wl[435] vdd gnd cell_6t
Xbit_r436_c103 bl[103] br[103] wl[436] vdd gnd cell_6t
Xbit_r437_c103 bl[103] br[103] wl[437] vdd gnd cell_6t
Xbit_r438_c103 bl[103] br[103] wl[438] vdd gnd cell_6t
Xbit_r439_c103 bl[103] br[103] wl[439] vdd gnd cell_6t
Xbit_r440_c103 bl[103] br[103] wl[440] vdd gnd cell_6t
Xbit_r441_c103 bl[103] br[103] wl[441] vdd gnd cell_6t
Xbit_r442_c103 bl[103] br[103] wl[442] vdd gnd cell_6t
Xbit_r443_c103 bl[103] br[103] wl[443] vdd gnd cell_6t
Xbit_r444_c103 bl[103] br[103] wl[444] vdd gnd cell_6t
Xbit_r445_c103 bl[103] br[103] wl[445] vdd gnd cell_6t
Xbit_r446_c103 bl[103] br[103] wl[446] vdd gnd cell_6t
Xbit_r447_c103 bl[103] br[103] wl[447] vdd gnd cell_6t
Xbit_r448_c103 bl[103] br[103] wl[448] vdd gnd cell_6t
Xbit_r449_c103 bl[103] br[103] wl[449] vdd gnd cell_6t
Xbit_r450_c103 bl[103] br[103] wl[450] vdd gnd cell_6t
Xbit_r451_c103 bl[103] br[103] wl[451] vdd gnd cell_6t
Xbit_r452_c103 bl[103] br[103] wl[452] vdd gnd cell_6t
Xbit_r453_c103 bl[103] br[103] wl[453] vdd gnd cell_6t
Xbit_r454_c103 bl[103] br[103] wl[454] vdd gnd cell_6t
Xbit_r455_c103 bl[103] br[103] wl[455] vdd gnd cell_6t
Xbit_r456_c103 bl[103] br[103] wl[456] vdd gnd cell_6t
Xbit_r457_c103 bl[103] br[103] wl[457] vdd gnd cell_6t
Xbit_r458_c103 bl[103] br[103] wl[458] vdd gnd cell_6t
Xbit_r459_c103 bl[103] br[103] wl[459] vdd gnd cell_6t
Xbit_r460_c103 bl[103] br[103] wl[460] vdd gnd cell_6t
Xbit_r461_c103 bl[103] br[103] wl[461] vdd gnd cell_6t
Xbit_r462_c103 bl[103] br[103] wl[462] vdd gnd cell_6t
Xbit_r463_c103 bl[103] br[103] wl[463] vdd gnd cell_6t
Xbit_r464_c103 bl[103] br[103] wl[464] vdd gnd cell_6t
Xbit_r465_c103 bl[103] br[103] wl[465] vdd gnd cell_6t
Xbit_r466_c103 bl[103] br[103] wl[466] vdd gnd cell_6t
Xbit_r467_c103 bl[103] br[103] wl[467] vdd gnd cell_6t
Xbit_r468_c103 bl[103] br[103] wl[468] vdd gnd cell_6t
Xbit_r469_c103 bl[103] br[103] wl[469] vdd gnd cell_6t
Xbit_r470_c103 bl[103] br[103] wl[470] vdd gnd cell_6t
Xbit_r471_c103 bl[103] br[103] wl[471] vdd gnd cell_6t
Xbit_r472_c103 bl[103] br[103] wl[472] vdd gnd cell_6t
Xbit_r473_c103 bl[103] br[103] wl[473] vdd gnd cell_6t
Xbit_r474_c103 bl[103] br[103] wl[474] vdd gnd cell_6t
Xbit_r475_c103 bl[103] br[103] wl[475] vdd gnd cell_6t
Xbit_r476_c103 bl[103] br[103] wl[476] vdd gnd cell_6t
Xbit_r477_c103 bl[103] br[103] wl[477] vdd gnd cell_6t
Xbit_r478_c103 bl[103] br[103] wl[478] vdd gnd cell_6t
Xbit_r479_c103 bl[103] br[103] wl[479] vdd gnd cell_6t
Xbit_r480_c103 bl[103] br[103] wl[480] vdd gnd cell_6t
Xbit_r481_c103 bl[103] br[103] wl[481] vdd gnd cell_6t
Xbit_r482_c103 bl[103] br[103] wl[482] vdd gnd cell_6t
Xbit_r483_c103 bl[103] br[103] wl[483] vdd gnd cell_6t
Xbit_r484_c103 bl[103] br[103] wl[484] vdd gnd cell_6t
Xbit_r485_c103 bl[103] br[103] wl[485] vdd gnd cell_6t
Xbit_r486_c103 bl[103] br[103] wl[486] vdd gnd cell_6t
Xbit_r487_c103 bl[103] br[103] wl[487] vdd gnd cell_6t
Xbit_r488_c103 bl[103] br[103] wl[488] vdd gnd cell_6t
Xbit_r489_c103 bl[103] br[103] wl[489] vdd gnd cell_6t
Xbit_r490_c103 bl[103] br[103] wl[490] vdd gnd cell_6t
Xbit_r491_c103 bl[103] br[103] wl[491] vdd gnd cell_6t
Xbit_r492_c103 bl[103] br[103] wl[492] vdd gnd cell_6t
Xbit_r493_c103 bl[103] br[103] wl[493] vdd gnd cell_6t
Xbit_r494_c103 bl[103] br[103] wl[494] vdd gnd cell_6t
Xbit_r495_c103 bl[103] br[103] wl[495] vdd gnd cell_6t
Xbit_r496_c103 bl[103] br[103] wl[496] vdd gnd cell_6t
Xbit_r497_c103 bl[103] br[103] wl[497] vdd gnd cell_6t
Xbit_r498_c103 bl[103] br[103] wl[498] vdd gnd cell_6t
Xbit_r499_c103 bl[103] br[103] wl[499] vdd gnd cell_6t
Xbit_r500_c103 bl[103] br[103] wl[500] vdd gnd cell_6t
Xbit_r501_c103 bl[103] br[103] wl[501] vdd gnd cell_6t
Xbit_r502_c103 bl[103] br[103] wl[502] vdd gnd cell_6t
Xbit_r503_c103 bl[103] br[103] wl[503] vdd gnd cell_6t
Xbit_r504_c103 bl[103] br[103] wl[504] vdd gnd cell_6t
Xbit_r505_c103 bl[103] br[103] wl[505] vdd gnd cell_6t
Xbit_r506_c103 bl[103] br[103] wl[506] vdd gnd cell_6t
Xbit_r507_c103 bl[103] br[103] wl[507] vdd gnd cell_6t
Xbit_r508_c103 bl[103] br[103] wl[508] vdd gnd cell_6t
Xbit_r509_c103 bl[103] br[103] wl[509] vdd gnd cell_6t
Xbit_r510_c103 bl[103] br[103] wl[510] vdd gnd cell_6t
Xbit_r511_c103 bl[103] br[103] wl[511] vdd gnd cell_6t
Xbit_r0_c104 bl[104] br[104] wl[0] vdd gnd cell_6t
Xbit_r1_c104 bl[104] br[104] wl[1] vdd gnd cell_6t
Xbit_r2_c104 bl[104] br[104] wl[2] vdd gnd cell_6t
Xbit_r3_c104 bl[104] br[104] wl[3] vdd gnd cell_6t
Xbit_r4_c104 bl[104] br[104] wl[4] vdd gnd cell_6t
Xbit_r5_c104 bl[104] br[104] wl[5] vdd gnd cell_6t
Xbit_r6_c104 bl[104] br[104] wl[6] vdd gnd cell_6t
Xbit_r7_c104 bl[104] br[104] wl[7] vdd gnd cell_6t
Xbit_r8_c104 bl[104] br[104] wl[8] vdd gnd cell_6t
Xbit_r9_c104 bl[104] br[104] wl[9] vdd gnd cell_6t
Xbit_r10_c104 bl[104] br[104] wl[10] vdd gnd cell_6t
Xbit_r11_c104 bl[104] br[104] wl[11] vdd gnd cell_6t
Xbit_r12_c104 bl[104] br[104] wl[12] vdd gnd cell_6t
Xbit_r13_c104 bl[104] br[104] wl[13] vdd gnd cell_6t
Xbit_r14_c104 bl[104] br[104] wl[14] vdd gnd cell_6t
Xbit_r15_c104 bl[104] br[104] wl[15] vdd gnd cell_6t
Xbit_r16_c104 bl[104] br[104] wl[16] vdd gnd cell_6t
Xbit_r17_c104 bl[104] br[104] wl[17] vdd gnd cell_6t
Xbit_r18_c104 bl[104] br[104] wl[18] vdd gnd cell_6t
Xbit_r19_c104 bl[104] br[104] wl[19] vdd gnd cell_6t
Xbit_r20_c104 bl[104] br[104] wl[20] vdd gnd cell_6t
Xbit_r21_c104 bl[104] br[104] wl[21] vdd gnd cell_6t
Xbit_r22_c104 bl[104] br[104] wl[22] vdd gnd cell_6t
Xbit_r23_c104 bl[104] br[104] wl[23] vdd gnd cell_6t
Xbit_r24_c104 bl[104] br[104] wl[24] vdd gnd cell_6t
Xbit_r25_c104 bl[104] br[104] wl[25] vdd gnd cell_6t
Xbit_r26_c104 bl[104] br[104] wl[26] vdd gnd cell_6t
Xbit_r27_c104 bl[104] br[104] wl[27] vdd gnd cell_6t
Xbit_r28_c104 bl[104] br[104] wl[28] vdd gnd cell_6t
Xbit_r29_c104 bl[104] br[104] wl[29] vdd gnd cell_6t
Xbit_r30_c104 bl[104] br[104] wl[30] vdd gnd cell_6t
Xbit_r31_c104 bl[104] br[104] wl[31] vdd gnd cell_6t
Xbit_r32_c104 bl[104] br[104] wl[32] vdd gnd cell_6t
Xbit_r33_c104 bl[104] br[104] wl[33] vdd gnd cell_6t
Xbit_r34_c104 bl[104] br[104] wl[34] vdd gnd cell_6t
Xbit_r35_c104 bl[104] br[104] wl[35] vdd gnd cell_6t
Xbit_r36_c104 bl[104] br[104] wl[36] vdd gnd cell_6t
Xbit_r37_c104 bl[104] br[104] wl[37] vdd gnd cell_6t
Xbit_r38_c104 bl[104] br[104] wl[38] vdd gnd cell_6t
Xbit_r39_c104 bl[104] br[104] wl[39] vdd gnd cell_6t
Xbit_r40_c104 bl[104] br[104] wl[40] vdd gnd cell_6t
Xbit_r41_c104 bl[104] br[104] wl[41] vdd gnd cell_6t
Xbit_r42_c104 bl[104] br[104] wl[42] vdd gnd cell_6t
Xbit_r43_c104 bl[104] br[104] wl[43] vdd gnd cell_6t
Xbit_r44_c104 bl[104] br[104] wl[44] vdd gnd cell_6t
Xbit_r45_c104 bl[104] br[104] wl[45] vdd gnd cell_6t
Xbit_r46_c104 bl[104] br[104] wl[46] vdd gnd cell_6t
Xbit_r47_c104 bl[104] br[104] wl[47] vdd gnd cell_6t
Xbit_r48_c104 bl[104] br[104] wl[48] vdd gnd cell_6t
Xbit_r49_c104 bl[104] br[104] wl[49] vdd gnd cell_6t
Xbit_r50_c104 bl[104] br[104] wl[50] vdd gnd cell_6t
Xbit_r51_c104 bl[104] br[104] wl[51] vdd gnd cell_6t
Xbit_r52_c104 bl[104] br[104] wl[52] vdd gnd cell_6t
Xbit_r53_c104 bl[104] br[104] wl[53] vdd gnd cell_6t
Xbit_r54_c104 bl[104] br[104] wl[54] vdd gnd cell_6t
Xbit_r55_c104 bl[104] br[104] wl[55] vdd gnd cell_6t
Xbit_r56_c104 bl[104] br[104] wl[56] vdd gnd cell_6t
Xbit_r57_c104 bl[104] br[104] wl[57] vdd gnd cell_6t
Xbit_r58_c104 bl[104] br[104] wl[58] vdd gnd cell_6t
Xbit_r59_c104 bl[104] br[104] wl[59] vdd gnd cell_6t
Xbit_r60_c104 bl[104] br[104] wl[60] vdd gnd cell_6t
Xbit_r61_c104 bl[104] br[104] wl[61] vdd gnd cell_6t
Xbit_r62_c104 bl[104] br[104] wl[62] vdd gnd cell_6t
Xbit_r63_c104 bl[104] br[104] wl[63] vdd gnd cell_6t
Xbit_r64_c104 bl[104] br[104] wl[64] vdd gnd cell_6t
Xbit_r65_c104 bl[104] br[104] wl[65] vdd gnd cell_6t
Xbit_r66_c104 bl[104] br[104] wl[66] vdd gnd cell_6t
Xbit_r67_c104 bl[104] br[104] wl[67] vdd gnd cell_6t
Xbit_r68_c104 bl[104] br[104] wl[68] vdd gnd cell_6t
Xbit_r69_c104 bl[104] br[104] wl[69] vdd gnd cell_6t
Xbit_r70_c104 bl[104] br[104] wl[70] vdd gnd cell_6t
Xbit_r71_c104 bl[104] br[104] wl[71] vdd gnd cell_6t
Xbit_r72_c104 bl[104] br[104] wl[72] vdd gnd cell_6t
Xbit_r73_c104 bl[104] br[104] wl[73] vdd gnd cell_6t
Xbit_r74_c104 bl[104] br[104] wl[74] vdd gnd cell_6t
Xbit_r75_c104 bl[104] br[104] wl[75] vdd gnd cell_6t
Xbit_r76_c104 bl[104] br[104] wl[76] vdd gnd cell_6t
Xbit_r77_c104 bl[104] br[104] wl[77] vdd gnd cell_6t
Xbit_r78_c104 bl[104] br[104] wl[78] vdd gnd cell_6t
Xbit_r79_c104 bl[104] br[104] wl[79] vdd gnd cell_6t
Xbit_r80_c104 bl[104] br[104] wl[80] vdd gnd cell_6t
Xbit_r81_c104 bl[104] br[104] wl[81] vdd gnd cell_6t
Xbit_r82_c104 bl[104] br[104] wl[82] vdd gnd cell_6t
Xbit_r83_c104 bl[104] br[104] wl[83] vdd gnd cell_6t
Xbit_r84_c104 bl[104] br[104] wl[84] vdd gnd cell_6t
Xbit_r85_c104 bl[104] br[104] wl[85] vdd gnd cell_6t
Xbit_r86_c104 bl[104] br[104] wl[86] vdd gnd cell_6t
Xbit_r87_c104 bl[104] br[104] wl[87] vdd gnd cell_6t
Xbit_r88_c104 bl[104] br[104] wl[88] vdd gnd cell_6t
Xbit_r89_c104 bl[104] br[104] wl[89] vdd gnd cell_6t
Xbit_r90_c104 bl[104] br[104] wl[90] vdd gnd cell_6t
Xbit_r91_c104 bl[104] br[104] wl[91] vdd gnd cell_6t
Xbit_r92_c104 bl[104] br[104] wl[92] vdd gnd cell_6t
Xbit_r93_c104 bl[104] br[104] wl[93] vdd gnd cell_6t
Xbit_r94_c104 bl[104] br[104] wl[94] vdd gnd cell_6t
Xbit_r95_c104 bl[104] br[104] wl[95] vdd gnd cell_6t
Xbit_r96_c104 bl[104] br[104] wl[96] vdd gnd cell_6t
Xbit_r97_c104 bl[104] br[104] wl[97] vdd gnd cell_6t
Xbit_r98_c104 bl[104] br[104] wl[98] vdd gnd cell_6t
Xbit_r99_c104 bl[104] br[104] wl[99] vdd gnd cell_6t
Xbit_r100_c104 bl[104] br[104] wl[100] vdd gnd cell_6t
Xbit_r101_c104 bl[104] br[104] wl[101] vdd gnd cell_6t
Xbit_r102_c104 bl[104] br[104] wl[102] vdd gnd cell_6t
Xbit_r103_c104 bl[104] br[104] wl[103] vdd gnd cell_6t
Xbit_r104_c104 bl[104] br[104] wl[104] vdd gnd cell_6t
Xbit_r105_c104 bl[104] br[104] wl[105] vdd gnd cell_6t
Xbit_r106_c104 bl[104] br[104] wl[106] vdd gnd cell_6t
Xbit_r107_c104 bl[104] br[104] wl[107] vdd gnd cell_6t
Xbit_r108_c104 bl[104] br[104] wl[108] vdd gnd cell_6t
Xbit_r109_c104 bl[104] br[104] wl[109] vdd gnd cell_6t
Xbit_r110_c104 bl[104] br[104] wl[110] vdd gnd cell_6t
Xbit_r111_c104 bl[104] br[104] wl[111] vdd gnd cell_6t
Xbit_r112_c104 bl[104] br[104] wl[112] vdd gnd cell_6t
Xbit_r113_c104 bl[104] br[104] wl[113] vdd gnd cell_6t
Xbit_r114_c104 bl[104] br[104] wl[114] vdd gnd cell_6t
Xbit_r115_c104 bl[104] br[104] wl[115] vdd gnd cell_6t
Xbit_r116_c104 bl[104] br[104] wl[116] vdd gnd cell_6t
Xbit_r117_c104 bl[104] br[104] wl[117] vdd gnd cell_6t
Xbit_r118_c104 bl[104] br[104] wl[118] vdd gnd cell_6t
Xbit_r119_c104 bl[104] br[104] wl[119] vdd gnd cell_6t
Xbit_r120_c104 bl[104] br[104] wl[120] vdd gnd cell_6t
Xbit_r121_c104 bl[104] br[104] wl[121] vdd gnd cell_6t
Xbit_r122_c104 bl[104] br[104] wl[122] vdd gnd cell_6t
Xbit_r123_c104 bl[104] br[104] wl[123] vdd gnd cell_6t
Xbit_r124_c104 bl[104] br[104] wl[124] vdd gnd cell_6t
Xbit_r125_c104 bl[104] br[104] wl[125] vdd gnd cell_6t
Xbit_r126_c104 bl[104] br[104] wl[126] vdd gnd cell_6t
Xbit_r127_c104 bl[104] br[104] wl[127] vdd gnd cell_6t
Xbit_r128_c104 bl[104] br[104] wl[128] vdd gnd cell_6t
Xbit_r129_c104 bl[104] br[104] wl[129] vdd gnd cell_6t
Xbit_r130_c104 bl[104] br[104] wl[130] vdd gnd cell_6t
Xbit_r131_c104 bl[104] br[104] wl[131] vdd gnd cell_6t
Xbit_r132_c104 bl[104] br[104] wl[132] vdd gnd cell_6t
Xbit_r133_c104 bl[104] br[104] wl[133] vdd gnd cell_6t
Xbit_r134_c104 bl[104] br[104] wl[134] vdd gnd cell_6t
Xbit_r135_c104 bl[104] br[104] wl[135] vdd gnd cell_6t
Xbit_r136_c104 bl[104] br[104] wl[136] vdd gnd cell_6t
Xbit_r137_c104 bl[104] br[104] wl[137] vdd gnd cell_6t
Xbit_r138_c104 bl[104] br[104] wl[138] vdd gnd cell_6t
Xbit_r139_c104 bl[104] br[104] wl[139] vdd gnd cell_6t
Xbit_r140_c104 bl[104] br[104] wl[140] vdd gnd cell_6t
Xbit_r141_c104 bl[104] br[104] wl[141] vdd gnd cell_6t
Xbit_r142_c104 bl[104] br[104] wl[142] vdd gnd cell_6t
Xbit_r143_c104 bl[104] br[104] wl[143] vdd gnd cell_6t
Xbit_r144_c104 bl[104] br[104] wl[144] vdd gnd cell_6t
Xbit_r145_c104 bl[104] br[104] wl[145] vdd gnd cell_6t
Xbit_r146_c104 bl[104] br[104] wl[146] vdd gnd cell_6t
Xbit_r147_c104 bl[104] br[104] wl[147] vdd gnd cell_6t
Xbit_r148_c104 bl[104] br[104] wl[148] vdd gnd cell_6t
Xbit_r149_c104 bl[104] br[104] wl[149] vdd gnd cell_6t
Xbit_r150_c104 bl[104] br[104] wl[150] vdd gnd cell_6t
Xbit_r151_c104 bl[104] br[104] wl[151] vdd gnd cell_6t
Xbit_r152_c104 bl[104] br[104] wl[152] vdd gnd cell_6t
Xbit_r153_c104 bl[104] br[104] wl[153] vdd gnd cell_6t
Xbit_r154_c104 bl[104] br[104] wl[154] vdd gnd cell_6t
Xbit_r155_c104 bl[104] br[104] wl[155] vdd gnd cell_6t
Xbit_r156_c104 bl[104] br[104] wl[156] vdd gnd cell_6t
Xbit_r157_c104 bl[104] br[104] wl[157] vdd gnd cell_6t
Xbit_r158_c104 bl[104] br[104] wl[158] vdd gnd cell_6t
Xbit_r159_c104 bl[104] br[104] wl[159] vdd gnd cell_6t
Xbit_r160_c104 bl[104] br[104] wl[160] vdd gnd cell_6t
Xbit_r161_c104 bl[104] br[104] wl[161] vdd gnd cell_6t
Xbit_r162_c104 bl[104] br[104] wl[162] vdd gnd cell_6t
Xbit_r163_c104 bl[104] br[104] wl[163] vdd gnd cell_6t
Xbit_r164_c104 bl[104] br[104] wl[164] vdd gnd cell_6t
Xbit_r165_c104 bl[104] br[104] wl[165] vdd gnd cell_6t
Xbit_r166_c104 bl[104] br[104] wl[166] vdd gnd cell_6t
Xbit_r167_c104 bl[104] br[104] wl[167] vdd gnd cell_6t
Xbit_r168_c104 bl[104] br[104] wl[168] vdd gnd cell_6t
Xbit_r169_c104 bl[104] br[104] wl[169] vdd gnd cell_6t
Xbit_r170_c104 bl[104] br[104] wl[170] vdd gnd cell_6t
Xbit_r171_c104 bl[104] br[104] wl[171] vdd gnd cell_6t
Xbit_r172_c104 bl[104] br[104] wl[172] vdd gnd cell_6t
Xbit_r173_c104 bl[104] br[104] wl[173] vdd gnd cell_6t
Xbit_r174_c104 bl[104] br[104] wl[174] vdd gnd cell_6t
Xbit_r175_c104 bl[104] br[104] wl[175] vdd gnd cell_6t
Xbit_r176_c104 bl[104] br[104] wl[176] vdd gnd cell_6t
Xbit_r177_c104 bl[104] br[104] wl[177] vdd gnd cell_6t
Xbit_r178_c104 bl[104] br[104] wl[178] vdd gnd cell_6t
Xbit_r179_c104 bl[104] br[104] wl[179] vdd gnd cell_6t
Xbit_r180_c104 bl[104] br[104] wl[180] vdd gnd cell_6t
Xbit_r181_c104 bl[104] br[104] wl[181] vdd gnd cell_6t
Xbit_r182_c104 bl[104] br[104] wl[182] vdd gnd cell_6t
Xbit_r183_c104 bl[104] br[104] wl[183] vdd gnd cell_6t
Xbit_r184_c104 bl[104] br[104] wl[184] vdd gnd cell_6t
Xbit_r185_c104 bl[104] br[104] wl[185] vdd gnd cell_6t
Xbit_r186_c104 bl[104] br[104] wl[186] vdd gnd cell_6t
Xbit_r187_c104 bl[104] br[104] wl[187] vdd gnd cell_6t
Xbit_r188_c104 bl[104] br[104] wl[188] vdd gnd cell_6t
Xbit_r189_c104 bl[104] br[104] wl[189] vdd gnd cell_6t
Xbit_r190_c104 bl[104] br[104] wl[190] vdd gnd cell_6t
Xbit_r191_c104 bl[104] br[104] wl[191] vdd gnd cell_6t
Xbit_r192_c104 bl[104] br[104] wl[192] vdd gnd cell_6t
Xbit_r193_c104 bl[104] br[104] wl[193] vdd gnd cell_6t
Xbit_r194_c104 bl[104] br[104] wl[194] vdd gnd cell_6t
Xbit_r195_c104 bl[104] br[104] wl[195] vdd gnd cell_6t
Xbit_r196_c104 bl[104] br[104] wl[196] vdd gnd cell_6t
Xbit_r197_c104 bl[104] br[104] wl[197] vdd gnd cell_6t
Xbit_r198_c104 bl[104] br[104] wl[198] vdd gnd cell_6t
Xbit_r199_c104 bl[104] br[104] wl[199] vdd gnd cell_6t
Xbit_r200_c104 bl[104] br[104] wl[200] vdd gnd cell_6t
Xbit_r201_c104 bl[104] br[104] wl[201] vdd gnd cell_6t
Xbit_r202_c104 bl[104] br[104] wl[202] vdd gnd cell_6t
Xbit_r203_c104 bl[104] br[104] wl[203] vdd gnd cell_6t
Xbit_r204_c104 bl[104] br[104] wl[204] vdd gnd cell_6t
Xbit_r205_c104 bl[104] br[104] wl[205] vdd gnd cell_6t
Xbit_r206_c104 bl[104] br[104] wl[206] vdd gnd cell_6t
Xbit_r207_c104 bl[104] br[104] wl[207] vdd gnd cell_6t
Xbit_r208_c104 bl[104] br[104] wl[208] vdd gnd cell_6t
Xbit_r209_c104 bl[104] br[104] wl[209] vdd gnd cell_6t
Xbit_r210_c104 bl[104] br[104] wl[210] vdd gnd cell_6t
Xbit_r211_c104 bl[104] br[104] wl[211] vdd gnd cell_6t
Xbit_r212_c104 bl[104] br[104] wl[212] vdd gnd cell_6t
Xbit_r213_c104 bl[104] br[104] wl[213] vdd gnd cell_6t
Xbit_r214_c104 bl[104] br[104] wl[214] vdd gnd cell_6t
Xbit_r215_c104 bl[104] br[104] wl[215] vdd gnd cell_6t
Xbit_r216_c104 bl[104] br[104] wl[216] vdd gnd cell_6t
Xbit_r217_c104 bl[104] br[104] wl[217] vdd gnd cell_6t
Xbit_r218_c104 bl[104] br[104] wl[218] vdd gnd cell_6t
Xbit_r219_c104 bl[104] br[104] wl[219] vdd gnd cell_6t
Xbit_r220_c104 bl[104] br[104] wl[220] vdd gnd cell_6t
Xbit_r221_c104 bl[104] br[104] wl[221] vdd gnd cell_6t
Xbit_r222_c104 bl[104] br[104] wl[222] vdd gnd cell_6t
Xbit_r223_c104 bl[104] br[104] wl[223] vdd gnd cell_6t
Xbit_r224_c104 bl[104] br[104] wl[224] vdd gnd cell_6t
Xbit_r225_c104 bl[104] br[104] wl[225] vdd gnd cell_6t
Xbit_r226_c104 bl[104] br[104] wl[226] vdd gnd cell_6t
Xbit_r227_c104 bl[104] br[104] wl[227] vdd gnd cell_6t
Xbit_r228_c104 bl[104] br[104] wl[228] vdd gnd cell_6t
Xbit_r229_c104 bl[104] br[104] wl[229] vdd gnd cell_6t
Xbit_r230_c104 bl[104] br[104] wl[230] vdd gnd cell_6t
Xbit_r231_c104 bl[104] br[104] wl[231] vdd gnd cell_6t
Xbit_r232_c104 bl[104] br[104] wl[232] vdd gnd cell_6t
Xbit_r233_c104 bl[104] br[104] wl[233] vdd gnd cell_6t
Xbit_r234_c104 bl[104] br[104] wl[234] vdd gnd cell_6t
Xbit_r235_c104 bl[104] br[104] wl[235] vdd gnd cell_6t
Xbit_r236_c104 bl[104] br[104] wl[236] vdd gnd cell_6t
Xbit_r237_c104 bl[104] br[104] wl[237] vdd gnd cell_6t
Xbit_r238_c104 bl[104] br[104] wl[238] vdd gnd cell_6t
Xbit_r239_c104 bl[104] br[104] wl[239] vdd gnd cell_6t
Xbit_r240_c104 bl[104] br[104] wl[240] vdd gnd cell_6t
Xbit_r241_c104 bl[104] br[104] wl[241] vdd gnd cell_6t
Xbit_r242_c104 bl[104] br[104] wl[242] vdd gnd cell_6t
Xbit_r243_c104 bl[104] br[104] wl[243] vdd gnd cell_6t
Xbit_r244_c104 bl[104] br[104] wl[244] vdd gnd cell_6t
Xbit_r245_c104 bl[104] br[104] wl[245] vdd gnd cell_6t
Xbit_r246_c104 bl[104] br[104] wl[246] vdd gnd cell_6t
Xbit_r247_c104 bl[104] br[104] wl[247] vdd gnd cell_6t
Xbit_r248_c104 bl[104] br[104] wl[248] vdd gnd cell_6t
Xbit_r249_c104 bl[104] br[104] wl[249] vdd gnd cell_6t
Xbit_r250_c104 bl[104] br[104] wl[250] vdd gnd cell_6t
Xbit_r251_c104 bl[104] br[104] wl[251] vdd gnd cell_6t
Xbit_r252_c104 bl[104] br[104] wl[252] vdd gnd cell_6t
Xbit_r253_c104 bl[104] br[104] wl[253] vdd gnd cell_6t
Xbit_r254_c104 bl[104] br[104] wl[254] vdd gnd cell_6t
Xbit_r255_c104 bl[104] br[104] wl[255] vdd gnd cell_6t
Xbit_r256_c104 bl[104] br[104] wl[256] vdd gnd cell_6t
Xbit_r257_c104 bl[104] br[104] wl[257] vdd gnd cell_6t
Xbit_r258_c104 bl[104] br[104] wl[258] vdd gnd cell_6t
Xbit_r259_c104 bl[104] br[104] wl[259] vdd gnd cell_6t
Xbit_r260_c104 bl[104] br[104] wl[260] vdd gnd cell_6t
Xbit_r261_c104 bl[104] br[104] wl[261] vdd gnd cell_6t
Xbit_r262_c104 bl[104] br[104] wl[262] vdd gnd cell_6t
Xbit_r263_c104 bl[104] br[104] wl[263] vdd gnd cell_6t
Xbit_r264_c104 bl[104] br[104] wl[264] vdd gnd cell_6t
Xbit_r265_c104 bl[104] br[104] wl[265] vdd gnd cell_6t
Xbit_r266_c104 bl[104] br[104] wl[266] vdd gnd cell_6t
Xbit_r267_c104 bl[104] br[104] wl[267] vdd gnd cell_6t
Xbit_r268_c104 bl[104] br[104] wl[268] vdd gnd cell_6t
Xbit_r269_c104 bl[104] br[104] wl[269] vdd gnd cell_6t
Xbit_r270_c104 bl[104] br[104] wl[270] vdd gnd cell_6t
Xbit_r271_c104 bl[104] br[104] wl[271] vdd gnd cell_6t
Xbit_r272_c104 bl[104] br[104] wl[272] vdd gnd cell_6t
Xbit_r273_c104 bl[104] br[104] wl[273] vdd gnd cell_6t
Xbit_r274_c104 bl[104] br[104] wl[274] vdd gnd cell_6t
Xbit_r275_c104 bl[104] br[104] wl[275] vdd gnd cell_6t
Xbit_r276_c104 bl[104] br[104] wl[276] vdd gnd cell_6t
Xbit_r277_c104 bl[104] br[104] wl[277] vdd gnd cell_6t
Xbit_r278_c104 bl[104] br[104] wl[278] vdd gnd cell_6t
Xbit_r279_c104 bl[104] br[104] wl[279] vdd gnd cell_6t
Xbit_r280_c104 bl[104] br[104] wl[280] vdd gnd cell_6t
Xbit_r281_c104 bl[104] br[104] wl[281] vdd gnd cell_6t
Xbit_r282_c104 bl[104] br[104] wl[282] vdd gnd cell_6t
Xbit_r283_c104 bl[104] br[104] wl[283] vdd gnd cell_6t
Xbit_r284_c104 bl[104] br[104] wl[284] vdd gnd cell_6t
Xbit_r285_c104 bl[104] br[104] wl[285] vdd gnd cell_6t
Xbit_r286_c104 bl[104] br[104] wl[286] vdd gnd cell_6t
Xbit_r287_c104 bl[104] br[104] wl[287] vdd gnd cell_6t
Xbit_r288_c104 bl[104] br[104] wl[288] vdd gnd cell_6t
Xbit_r289_c104 bl[104] br[104] wl[289] vdd gnd cell_6t
Xbit_r290_c104 bl[104] br[104] wl[290] vdd gnd cell_6t
Xbit_r291_c104 bl[104] br[104] wl[291] vdd gnd cell_6t
Xbit_r292_c104 bl[104] br[104] wl[292] vdd gnd cell_6t
Xbit_r293_c104 bl[104] br[104] wl[293] vdd gnd cell_6t
Xbit_r294_c104 bl[104] br[104] wl[294] vdd gnd cell_6t
Xbit_r295_c104 bl[104] br[104] wl[295] vdd gnd cell_6t
Xbit_r296_c104 bl[104] br[104] wl[296] vdd gnd cell_6t
Xbit_r297_c104 bl[104] br[104] wl[297] vdd gnd cell_6t
Xbit_r298_c104 bl[104] br[104] wl[298] vdd gnd cell_6t
Xbit_r299_c104 bl[104] br[104] wl[299] vdd gnd cell_6t
Xbit_r300_c104 bl[104] br[104] wl[300] vdd gnd cell_6t
Xbit_r301_c104 bl[104] br[104] wl[301] vdd gnd cell_6t
Xbit_r302_c104 bl[104] br[104] wl[302] vdd gnd cell_6t
Xbit_r303_c104 bl[104] br[104] wl[303] vdd gnd cell_6t
Xbit_r304_c104 bl[104] br[104] wl[304] vdd gnd cell_6t
Xbit_r305_c104 bl[104] br[104] wl[305] vdd gnd cell_6t
Xbit_r306_c104 bl[104] br[104] wl[306] vdd gnd cell_6t
Xbit_r307_c104 bl[104] br[104] wl[307] vdd gnd cell_6t
Xbit_r308_c104 bl[104] br[104] wl[308] vdd gnd cell_6t
Xbit_r309_c104 bl[104] br[104] wl[309] vdd gnd cell_6t
Xbit_r310_c104 bl[104] br[104] wl[310] vdd gnd cell_6t
Xbit_r311_c104 bl[104] br[104] wl[311] vdd gnd cell_6t
Xbit_r312_c104 bl[104] br[104] wl[312] vdd gnd cell_6t
Xbit_r313_c104 bl[104] br[104] wl[313] vdd gnd cell_6t
Xbit_r314_c104 bl[104] br[104] wl[314] vdd gnd cell_6t
Xbit_r315_c104 bl[104] br[104] wl[315] vdd gnd cell_6t
Xbit_r316_c104 bl[104] br[104] wl[316] vdd gnd cell_6t
Xbit_r317_c104 bl[104] br[104] wl[317] vdd gnd cell_6t
Xbit_r318_c104 bl[104] br[104] wl[318] vdd gnd cell_6t
Xbit_r319_c104 bl[104] br[104] wl[319] vdd gnd cell_6t
Xbit_r320_c104 bl[104] br[104] wl[320] vdd gnd cell_6t
Xbit_r321_c104 bl[104] br[104] wl[321] vdd gnd cell_6t
Xbit_r322_c104 bl[104] br[104] wl[322] vdd gnd cell_6t
Xbit_r323_c104 bl[104] br[104] wl[323] vdd gnd cell_6t
Xbit_r324_c104 bl[104] br[104] wl[324] vdd gnd cell_6t
Xbit_r325_c104 bl[104] br[104] wl[325] vdd gnd cell_6t
Xbit_r326_c104 bl[104] br[104] wl[326] vdd gnd cell_6t
Xbit_r327_c104 bl[104] br[104] wl[327] vdd gnd cell_6t
Xbit_r328_c104 bl[104] br[104] wl[328] vdd gnd cell_6t
Xbit_r329_c104 bl[104] br[104] wl[329] vdd gnd cell_6t
Xbit_r330_c104 bl[104] br[104] wl[330] vdd gnd cell_6t
Xbit_r331_c104 bl[104] br[104] wl[331] vdd gnd cell_6t
Xbit_r332_c104 bl[104] br[104] wl[332] vdd gnd cell_6t
Xbit_r333_c104 bl[104] br[104] wl[333] vdd gnd cell_6t
Xbit_r334_c104 bl[104] br[104] wl[334] vdd gnd cell_6t
Xbit_r335_c104 bl[104] br[104] wl[335] vdd gnd cell_6t
Xbit_r336_c104 bl[104] br[104] wl[336] vdd gnd cell_6t
Xbit_r337_c104 bl[104] br[104] wl[337] vdd gnd cell_6t
Xbit_r338_c104 bl[104] br[104] wl[338] vdd gnd cell_6t
Xbit_r339_c104 bl[104] br[104] wl[339] vdd gnd cell_6t
Xbit_r340_c104 bl[104] br[104] wl[340] vdd gnd cell_6t
Xbit_r341_c104 bl[104] br[104] wl[341] vdd gnd cell_6t
Xbit_r342_c104 bl[104] br[104] wl[342] vdd gnd cell_6t
Xbit_r343_c104 bl[104] br[104] wl[343] vdd gnd cell_6t
Xbit_r344_c104 bl[104] br[104] wl[344] vdd gnd cell_6t
Xbit_r345_c104 bl[104] br[104] wl[345] vdd gnd cell_6t
Xbit_r346_c104 bl[104] br[104] wl[346] vdd gnd cell_6t
Xbit_r347_c104 bl[104] br[104] wl[347] vdd gnd cell_6t
Xbit_r348_c104 bl[104] br[104] wl[348] vdd gnd cell_6t
Xbit_r349_c104 bl[104] br[104] wl[349] vdd gnd cell_6t
Xbit_r350_c104 bl[104] br[104] wl[350] vdd gnd cell_6t
Xbit_r351_c104 bl[104] br[104] wl[351] vdd gnd cell_6t
Xbit_r352_c104 bl[104] br[104] wl[352] vdd gnd cell_6t
Xbit_r353_c104 bl[104] br[104] wl[353] vdd gnd cell_6t
Xbit_r354_c104 bl[104] br[104] wl[354] vdd gnd cell_6t
Xbit_r355_c104 bl[104] br[104] wl[355] vdd gnd cell_6t
Xbit_r356_c104 bl[104] br[104] wl[356] vdd gnd cell_6t
Xbit_r357_c104 bl[104] br[104] wl[357] vdd gnd cell_6t
Xbit_r358_c104 bl[104] br[104] wl[358] vdd gnd cell_6t
Xbit_r359_c104 bl[104] br[104] wl[359] vdd gnd cell_6t
Xbit_r360_c104 bl[104] br[104] wl[360] vdd gnd cell_6t
Xbit_r361_c104 bl[104] br[104] wl[361] vdd gnd cell_6t
Xbit_r362_c104 bl[104] br[104] wl[362] vdd gnd cell_6t
Xbit_r363_c104 bl[104] br[104] wl[363] vdd gnd cell_6t
Xbit_r364_c104 bl[104] br[104] wl[364] vdd gnd cell_6t
Xbit_r365_c104 bl[104] br[104] wl[365] vdd gnd cell_6t
Xbit_r366_c104 bl[104] br[104] wl[366] vdd gnd cell_6t
Xbit_r367_c104 bl[104] br[104] wl[367] vdd gnd cell_6t
Xbit_r368_c104 bl[104] br[104] wl[368] vdd gnd cell_6t
Xbit_r369_c104 bl[104] br[104] wl[369] vdd gnd cell_6t
Xbit_r370_c104 bl[104] br[104] wl[370] vdd gnd cell_6t
Xbit_r371_c104 bl[104] br[104] wl[371] vdd gnd cell_6t
Xbit_r372_c104 bl[104] br[104] wl[372] vdd gnd cell_6t
Xbit_r373_c104 bl[104] br[104] wl[373] vdd gnd cell_6t
Xbit_r374_c104 bl[104] br[104] wl[374] vdd gnd cell_6t
Xbit_r375_c104 bl[104] br[104] wl[375] vdd gnd cell_6t
Xbit_r376_c104 bl[104] br[104] wl[376] vdd gnd cell_6t
Xbit_r377_c104 bl[104] br[104] wl[377] vdd gnd cell_6t
Xbit_r378_c104 bl[104] br[104] wl[378] vdd gnd cell_6t
Xbit_r379_c104 bl[104] br[104] wl[379] vdd gnd cell_6t
Xbit_r380_c104 bl[104] br[104] wl[380] vdd gnd cell_6t
Xbit_r381_c104 bl[104] br[104] wl[381] vdd gnd cell_6t
Xbit_r382_c104 bl[104] br[104] wl[382] vdd gnd cell_6t
Xbit_r383_c104 bl[104] br[104] wl[383] vdd gnd cell_6t
Xbit_r384_c104 bl[104] br[104] wl[384] vdd gnd cell_6t
Xbit_r385_c104 bl[104] br[104] wl[385] vdd gnd cell_6t
Xbit_r386_c104 bl[104] br[104] wl[386] vdd gnd cell_6t
Xbit_r387_c104 bl[104] br[104] wl[387] vdd gnd cell_6t
Xbit_r388_c104 bl[104] br[104] wl[388] vdd gnd cell_6t
Xbit_r389_c104 bl[104] br[104] wl[389] vdd gnd cell_6t
Xbit_r390_c104 bl[104] br[104] wl[390] vdd gnd cell_6t
Xbit_r391_c104 bl[104] br[104] wl[391] vdd gnd cell_6t
Xbit_r392_c104 bl[104] br[104] wl[392] vdd gnd cell_6t
Xbit_r393_c104 bl[104] br[104] wl[393] vdd gnd cell_6t
Xbit_r394_c104 bl[104] br[104] wl[394] vdd gnd cell_6t
Xbit_r395_c104 bl[104] br[104] wl[395] vdd gnd cell_6t
Xbit_r396_c104 bl[104] br[104] wl[396] vdd gnd cell_6t
Xbit_r397_c104 bl[104] br[104] wl[397] vdd gnd cell_6t
Xbit_r398_c104 bl[104] br[104] wl[398] vdd gnd cell_6t
Xbit_r399_c104 bl[104] br[104] wl[399] vdd gnd cell_6t
Xbit_r400_c104 bl[104] br[104] wl[400] vdd gnd cell_6t
Xbit_r401_c104 bl[104] br[104] wl[401] vdd gnd cell_6t
Xbit_r402_c104 bl[104] br[104] wl[402] vdd gnd cell_6t
Xbit_r403_c104 bl[104] br[104] wl[403] vdd gnd cell_6t
Xbit_r404_c104 bl[104] br[104] wl[404] vdd gnd cell_6t
Xbit_r405_c104 bl[104] br[104] wl[405] vdd gnd cell_6t
Xbit_r406_c104 bl[104] br[104] wl[406] vdd gnd cell_6t
Xbit_r407_c104 bl[104] br[104] wl[407] vdd gnd cell_6t
Xbit_r408_c104 bl[104] br[104] wl[408] vdd gnd cell_6t
Xbit_r409_c104 bl[104] br[104] wl[409] vdd gnd cell_6t
Xbit_r410_c104 bl[104] br[104] wl[410] vdd gnd cell_6t
Xbit_r411_c104 bl[104] br[104] wl[411] vdd gnd cell_6t
Xbit_r412_c104 bl[104] br[104] wl[412] vdd gnd cell_6t
Xbit_r413_c104 bl[104] br[104] wl[413] vdd gnd cell_6t
Xbit_r414_c104 bl[104] br[104] wl[414] vdd gnd cell_6t
Xbit_r415_c104 bl[104] br[104] wl[415] vdd gnd cell_6t
Xbit_r416_c104 bl[104] br[104] wl[416] vdd gnd cell_6t
Xbit_r417_c104 bl[104] br[104] wl[417] vdd gnd cell_6t
Xbit_r418_c104 bl[104] br[104] wl[418] vdd gnd cell_6t
Xbit_r419_c104 bl[104] br[104] wl[419] vdd gnd cell_6t
Xbit_r420_c104 bl[104] br[104] wl[420] vdd gnd cell_6t
Xbit_r421_c104 bl[104] br[104] wl[421] vdd gnd cell_6t
Xbit_r422_c104 bl[104] br[104] wl[422] vdd gnd cell_6t
Xbit_r423_c104 bl[104] br[104] wl[423] vdd gnd cell_6t
Xbit_r424_c104 bl[104] br[104] wl[424] vdd gnd cell_6t
Xbit_r425_c104 bl[104] br[104] wl[425] vdd gnd cell_6t
Xbit_r426_c104 bl[104] br[104] wl[426] vdd gnd cell_6t
Xbit_r427_c104 bl[104] br[104] wl[427] vdd gnd cell_6t
Xbit_r428_c104 bl[104] br[104] wl[428] vdd gnd cell_6t
Xbit_r429_c104 bl[104] br[104] wl[429] vdd gnd cell_6t
Xbit_r430_c104 bl[104] br[104] wl[430] vdd gnd cell_6t
Xbit_r431_c104 bl[104] br[104] wl[431] vdd gnd cell_6t
Xbit_r432_c104 bl[104] br[104] wl[432] vdd gnd cell_6t
Xbit_r433_c104 bl[104] br[104] wl[433] vdd gnd cell_6t
Xbit_r434_c104 bl[104] br[104] wl[434] vdd gnd cell_6t
Xbit_r435_c104 bl[104] br[104] wl[435] vdd gnd cell_6t
Xbit_r436_c104 bl[104] br[104] wl[436] vdd gnd cell_6t
Xbit_r437_c104 bl[104] br[104] wl[437] vdd gnd cell_6t
Xbit_r438_c104 bl[104] br[104] wl[438] vdd gnd cell_6t
Xbit_r439_c104 bl[104] br[104] wl[439] vdd gnd cell_6t
Xbit_r440_c104 bl[104] br[104] wl[440] vdd gnd cell_6t
Xbit_r441_c104 bl[104] br[104] wl[441] vdd gnd cell_6t
Xbit_r442_c104 bl[104] br[104] wl[442] vdd gnd cell_6t
Xbit_r443_c104 bl[104] br[104] wl[443] vdd gnd cell_6t
Xbit_r444_c104 bl[104] br[104] wl[444] vdd gnd cell_6t
Xbit_r445_c104 bl[104] br[104] wl[445] vdd gnd cell_6t
Xbit_r446_c104 bl[104] br[104] wl[446] vdd gnd cell_6t
Xbit_r447_c104 bl[104] br[104] wl[447] vdd gnd cell_6t
Xbit_r448_c104 bl[104] br[104] wl[448] vdd gnd cell_6t
Xbit_r449_c104 bl[104] br[104] wl[449] vdd gnd cell_6t
Xbit_r450_c104 bl[104] br[104] wl[450] vdd gnd cell_6t
Xbit_r451_c104 bl[104] br[104] wl[451] vdd gnd cell_6t
Xbit_r452_c104 bl[104] br[104] wl[452] vdd gnd cell_6t
Xbit_r453_c104 bl[104] br[104] wl[453] vdd gnd cell_6t
Xbit_r454_c104 bl[104] br[104] wl[454] vdd gnd cell_6t
Xbit_r455_c104 bl[104] br[104] wl[455] vdd gnd cell_6t
Xbit_r456_c104 bl[104] br[104] wl[456] vdd gnd cell_6t
Xbit_r457_c104 bl[104] br[104] wl[457] vdd gnd cell_6t
Xbit_r458_c104 bl[104] br[104] wl[458] vdd gnd cell_6t
Xbit_r459_c104 bl[104] br[104] wl[459] vdd gnd cell_6t
Xbit_r460_c104 bl[104] br[104] wl[460] vdd gnd cell_6t
Xbit_r461_c104 bl[104] br[104] wl[461] vdd gnd cell_6t
Xbit_r462_c104 bl[104] br[104] wl[462] vdd gnd cell_6t
Xbit_r463_c104 bl[104] br[104] wl[463] vdd gnd cell_6t
Xbit_r464_c104 bl[104] br[104] wl[464] vdd gnd cell_6t
Xbit_r465_c104 bl[104] br[104] wl[465] vdd gnd cell_6t
Xbit_r466_c104 bl[104] br[104] wl[466] vdd gnd cell_6t
Xbit_r467_c104 bl[104] br[104] wl[467] vdd gnd cell_6t
Xbit_r468_c104 bl[104] br[104] wl[468] vdd gnd cell_6t
Xbit_r469_c104 bl[104] br[104] wl[469] vdd gnd cell_6t
Xbit_r470_c104 bl[104] br[104] wl[470] vdd gnd cell_6t
Xbit_r471_c104 bl[104] br[104] wl[471] vdd gnd cell_6t
Xbit_r472_c104 bl[104] br[104] wl[472] vdd gnd cell_6t
Xbit_r473_c104 bl[104] br[104] wl[473] vdd gnd cell_6t
Xbit_r474_c104 bl[104] br[104] wl[474] vdd gnd cell_6t
Xbit_r475_c104 bl[104] br[104] wl[475] vdd gnd cell_6t
Xbit_r476_c104 bl[104] br[104] wl[476] vdd gnd cell_6t
Xbit_r477_c104 bl[104] br[104] wl[477] vdd gnd cell_6t
Xbit_r478_c104 bl[104] br[104] wl[478] vdd gnd cell_6t
Xbit_r479_c104 bl[104] br[104] wl[479] vdd gnd cell_6t
Xbit_r480_c104 bl[104] br[104] wl[480] vdd gnd cell_6t
Xbit_r481_c104 bl[104] br[104] wl[481] vdd gnd cell_6t
Xbit_r482_c104 bl[104] br[104] wl[482] vdd gnd cell_6t
Xbit_r483_c104 bl[104] br[104] wl[483] vdd gnd cell_6t
Xbit_r484_c104 bl[104] br[104] wl[484] vdd gnd cell_6t
Xbit_r485_c104 bl[104] br[104] wl[485] vdd gnd cell_6t
Xbit_r486_c104 bl[104] br[104] wl[486] vdd gnd cell_6t
Xbit_r487_c104 bl[104] br[104] wl[487] vdd gnd cell_6t
Xbit_r488_c104 bl[104] br[104] wl[488] vdd gnd cell_6t
Xbit_r489_c104 bl[104] br[104] wl[489] vdd gnd cell_6t
Xbit_r490_c104 bl[104] br[104] wl[490] vdd gnd cell_6t
Xbit_r491_c104 bl[104] br[104] wl[491] vdd gnd cell_6t
Xbit_r492_c104 bl[104] br[104] wl[492] vdd gnd cell_6t
Xbit_r493_c104 bl[104] br[104] wl[493] vdd gnd cell_6t
Xbit_r494_c104 bl[104] br[104] wl[494] vdd gnd cell_6t
Xbit_r495_c104 bl[104] br[104] wl[495] vdd gnd cell_6t
Xbit_r496_c104 bl[104] br[104] wl[496] vdd gnd cell_6t
Xbit_r497_c104 bl[104] br[104] wl[497] vdd gnd cell_6t
Xbit_r498_c104 bl[104] br[104] wl[498] vdd gnd cell_6t
Xbit_r499_c104 bl[104] br[104] wl[499] vdd gnd cell_6t
Xbit_r500_c104 bl[104] br[104] wl[500] vdd gnd cell_6t
Xbit_r501_c104 bl[104] br[104] wl[501] vdd gnd cell_6t
Xbit_r502_c104 bl[104] br[104] wl[502] vdd gnd cell_6t
Xbit_r503_c104 bl[104] br[104] wl[503] vdd gnd cell_6t
Xbit_r504_c104 bl[104] br[104] wl[504] vdd gnd cell_6t
Xbit_r505_c104 bl[104] br[104] wl[505] vdd gnd cell_6t
Xbit_r506_c104 bl[104] br[104] wl[506] vdd gnd cell_6t
Xbit_r507_c104 bl[104] br[104] wl[507] vdd gnd cell_6t
Xbit_r508_c104 bl[104] br[104] wl[508] vdd gnd cell_6t
Xbit_r509_c104 bl[104] br[104] wl[509] vdd gnd cell_6t
Xbit_r510_c104 bl[104] br[104] wl[510] vdd gnd cell_6t
Xbit_r511_c104 bl[104] br[104] wl[511] vdd gnd cell_6t
Xbit_r0_c105 bl[105] br[105] wl[0] vdd gnd cell_6t
Xbit_r1_c105 bl[105] br[105] wl[1] vdd gnd cell_6t
Xbit_r2_c105 bl[105] br[105] wl[2] vdd gnd cell_6t
Xbit_r3_c105 bl[105] br[105] wl[3] vdd gnd cell_6t
Xbit_r4_c105 bl[105] br[105] wl[4] vdd gnd cell_6t
Xbit_r5_c105 bl[105] br[105] wl[5] vdd gnd cell_6t
Xbit_r6_c105 bl[105] br[105] wl[6] vdd gnd cell_6t
Xbit_r7_c105 bl[105] br[105] wl[7] vdd gnd cell_6t
Xbit_r8_c105 bl[105] br[105] wl[8] vdd gnd cell_6t
Xbit_r9_c105 bl[105] br[105] wl[9] vdd gnd cell_6t
Xbit_r10_c105 bl[105] br[105] wl[10] vdd gnd cell_6t
Xbit_r11_c105 bl[105] br[105] wl[11] vdd gnd cell_6t
Xbit_r12_c105 bl[105] br[105] wl[12] vdd gnd cell_6t
Xbit_r13_c105 bl[105] br[105] wl[13] vdd gnd cell_6t
Xbit_r14_c105 bl[105] br[105] wl[14] vdd gnd cell_6t
Xbit_r15_c105 bl[105] br[105] wl[15] vdd gnd cell_6t
Xbit_r16_c105 bl[105] br[105] wl[16] vdd gnd cell_6t
Xbit_r17_c105 bl[105] br[105] wl[17] vdd gnd cell_6t
Xbit_r18_c105 bl[105] br[105] wl[18] vdd gnd cell_6t
Xbit_r19_c105 bl[105] br[105] wl[19] vdd gnd cell_6t
Xbit_r20_c105 bl[105] br[105] wl[20] vdd gnd cell_6t
Xbit_r21_c105 bl[105] br[105] wl[21] vdd gnd cell_6t
Xbit_r22_c105 bl[105] br[105] wl[22] vdd gnd cell_6t
Xbit_r23_c105 bl[105] br[105] wl[23] vdd gnd cell_6t
Xbit_r24_c105 bl[105] br[105] wl[24] vdd gnd cell_6t
Xbit_r25_c105 bl[105] br[105] wl[25] vdd gnd cell_6t
Xbit_r26_c105 bl[105] br[105] wl[26] vdd gnd cell_6t
Xbit_r27_c105 bl[105] br[105] wl[27] vdd gnd cell_6t
Xbit_r28_c105 bl[105] br[105] wl[28] vdd gnd cell_6t
Xbit_r29_c105 bl[105] br[105] wl[29] vdd gnd cell_6t
Xbit_r30_c105 bl[105] br[105] wl[30] vdd gnd cell_6t
Xbit_r31_c105 bl[105] br[105] wl[31] vdd gnd cell_6t
Xbit_r32_c105 bl[105] br[105] wl[32] vdd gnd cell_6t
Xbit_r33_c105 bl[105] br[105] wl[33] vdd gnd cell_6t
Xbit_r34_c105 bl[105] br[105] wl[34] vdd gnd cell_6t
Xbit_r35_c105 bl[105] br[105] wl[35] vdd gnd cell_6t
Xbit_r36_c105 bl[105] br[105] wl[36] vdd gnd cell_6t
Xbit_r37_c105 bl[105] br[105] wl[37] vdd gnd cell_6t
Xbit_r38_c105 bl[105] br[105] wl[38] vdd gnd cell_6t
Xbit_r39_c105 bl[105] br[105] wl[39] vdd gnd cell_6t
Xbit_r40_c105 bl[105] br[105] wl[40] vdd gnd cell_6t
Xbit_r41_c105 bl[105] br[105] wl[41] vdd gnd cell_6t
Xbit_r42_c105 bl[105] br[105] wl[42] vdd gnd cell_6t
Xbit_r43_c105 bl[105] br[105] wl[43] vdd gnd cell_6t
Xbit_r44_c105 bl[105] br[105] wl[44] vdd gnd cell_6t
Xbit_r45_c105 bl[105] br[105] wl[45] vdd gnd cell_6t
Xbit_r46_c105 bl[105] br[105] wl[46] vdd gnd cell_6t
Xbit_r47_c105 bl[105] br[105] wl[47] vdd gnd cell_6t
Xbit_r48_c105 bl[105] br[105] wl[48] vdd gnd cell_6t
Xbit_r49_c105 bl[105] br[105] wl[49] vdd gnd cell_6t
Xbit_r50_c105 bl[105] br[105] wl[50] vdd gnd cell_6t
Xbit_r51_c105 bl[105] br[105] wl[51] vdd gnd cell_6t
Xbit_r52_c105 bl[105] br[105] wl[52] vdd gnd cell_6t
Xbit_r53_c105 bl[105] br[105] wl[53] vdd gnd cell_6t
Xbit_r54_c105 bl[105] br[105] wl[54] vdd gnd cell_6t
Xbit_r55_c105 bl[105] br[105] wl[55] vdd gnd cell_6t
Xbit_r56_c105 bl[105] br[105] wl[56] vdd gnd cell_6t
Xbit_r57_c105 bl[105] br[105] wl[57] vdd gnd cell_6t
Xbit_r58_c105 bl[105] br[105] wl[58] vdd gnd cell_6t
Xbit_r59_c105 bl[105] br[105] wl[59] vdd gnd cell_6t
Xbit_r60_c105 bl[105] br[105] wl[60] vdd gnd cell_6t
Xbit_r61_c105 bl[105] br[105] wl[61] vdd gnd cell_6t
Xbit_r62_c105 bl[105] br[105] wl[62] vdd gnd cell_6t
Xbit_r63_c105 bl[105] br[105] wl[63] vdd gnd cell_6t
Xbit_r64_c105 bl[105] br[105] wl[64] vdd gnd cell_6t
Xbit_r65_c105 bl[105] br[105] wl[65] vdd gnd cell_6t
Xbit_r66_c105 bl[105] br[105] wl[66] vdd gnd cell_6t
Xbit_r67_c105 bl[105] br[105] wl[67] vdd gnd cell_6t
Xbit_r68_c105 bl[105] br[105] wl[68] vdd gnd cell_6t
Xbit_r69_c105 bl[105] br[105] wl[69] vdd gnd cell_6t
Xbit_r70_c105 bl[105] br[105] wl[70] vdd gnd cell_6t
Xbit_r71_c105 bl[105] br[105] wl[71] vdd gnd cell_6t
Xbit_r72_c105 bl[105] br[105] wl[72] vdd gnd cell_6t
Xbit_r73_c105 bl[105] br[105] wl[73] vdd gnd cell_6t
Xbit_r74_c105 bl[105] br[105] wl[74] vdd gnd cell_6t
Xbit_r75_c105 bl[105] br[105] wl[75] vdd gnd cell_6t
Xbit_r76_c105 bl[105] br[105] wl[76] vdd gnd cell_6t
Xbit_r77_c105 bl[105] br[105] wl[77] vdd gnd cell_6t
Xbit_r78_c105 bl[105] br[105] wl[78] vdd gnd cell_6t
Xbit_r79_c105 bl[105] br[105] wl[79] vdd gnd cell_6t
Xbit_r80_c105 bl[105] br[105] wl[80] vdd gnd cell_6t
Xbit_r81_c105 bl[105] br[105] wl[81] vdd gnd cell_6t
Xbit_r82_c105 bl[105] br[105] wl[82] vdd gnd cell_6t
Xbit_r83_c105 bl[105] br[105] wl[83] vdd gnd cell_6t
Xbit_r84_c105 bl[105] br[105] wl[84] vdd gnd cell_6t
Xbit_r85_c105 bl[105] br[105] wl[85] vdd gnd cell_6t
Xbit_r86_c105 bl[105] br[105] wl[86] vdd gnd cell_6t
Xbit_r87_c105 bl[105] br[105] wl[87] vdd gnd cell_6t
Xbit_r88_c105 bl[105] br[105] wl[88] vdd gnd cell_6t
Xbit_r89_c105 bl[105] br[105] wl[89] vdd gnd cell_6t
Xbit_r90_c105 bl[105] br[105] wl[90] vdd gnd cell_6t
Xbit_r91_c105 bl[105] br[105] wl[91] vdd gnd cell_6t
Xbit_r92_c105 bl[105] br[105] wl[92] vdd gnd cell_6t
Xbit_r93_c105 bl[105] br[105] wl[93] vdd gnd cell_6t
Xbit_r94_c105 bl[105] br[105] wl[94] vdd gnd cell_6t
Xbit_r95_c105 bl[105] br[105] wl[95] vdd gnd cell_6t
Xbit_r96_c105 bl[105] br[105] wl[96] vdd gnd cell_6t
Xbit_r97_c105 bl[105] br[105] wl[97] vdd gnd cell_6t
Xbit_r98_c105 bl[105] br[105] wl[98] vdd gnd cell_6t
Xbit_r99_c105 bl[105] br[105] wl[99] vdd gnd cell_6t
Xbit_r100_c105 bl[105] br[105] wl[100] vdd gnd cell_6t
Xbit_r101_c105 bl[105] br[105] wl[101] vdd gnd cell_6t
Xbit_r102_c105 bl[105] br[105] wl[102] vdd gnd cell_6t
Xbit_r103_c105 bl[105] br[105] wl[103] vdd gnd cell_6t
Xbit_r104_c105 bl[105] br[105] wl[104] vdd gnd cell_6t
Xbit_r105_c105 bl[105] br[105] wl[105] vdd gnd cell_6t
Xbit_r106_c105 bl[105] br[105] wl[106] vdd gnd cell_6t
Xbit_r107_c105 bl[105] br[105] wl[107] vdd gnd cell_6t
Xbit_r108_c105 bl[105] br[105] wl[108] vdd gnd cell_6t
Xbit_r109_c105 bl[105] br[105] wl[109] vdd gnd cell_6t
Xbit_r110_c105 bl[105] br[105] wl[110] vdd gnd cell_6t
Xbit_r111_c105 bl[105] br[105] wl[111] vdd gnd cell_6t
Xbit_r112_c105 bl[105] br[105] wl[112] vdd gnd cell_6t
Xbit_r113_c105 bl[105] br[105] wl[113] vdd gnd cell_6t
Xbit_r114_c105 bl[105] br[105] wl[114] vdd gnd cell_6t
Xbit_r115_c105 bl[105] br[105] wl[115] vdd gnd cell_6t
Xbit_r116_c105 bl[105] br[105] wl[116] vdd gnd cell_6t
Xbit_r117_c105 bl[105] br[105] wl[117] vdd gnd cell_6t
Xbit_r118_c105 bl[105] br[105] wl[118] vdd gnd cell_6t
Xbit_r119_c105 bl[105] br[105] wl[119] vdd gnd cell_6t
Xbit_r120_c105 bl[105] br[105] wl[120] vdd gnd cell_6t
Xbit_r121_c105 bl[105] br[105] wl[121] vdd gnd cell_6t
Xbit_r122_c105 bl[105] br[105] wl[122] vdd gnd cell_6t
Xbit_r123_c105 bl[105] br[105] wl[123] vdd gnd cell_6t
Xbit_r124_c105 bl[105] br[105] wl[124] vdd gnd cell_6t
Xbit_r125_c105 bl[105] br[105] wl[125] vdd gnd cell_6t
Xbit_r126_c105 bl[105] br[105] wl[126] vdd gnd cell_6t
Xbit_r127_c105 bl[105] br[105] wl[127] vdd gnd cell_6t
Xbit_r128_c105 bl[105] br[105] wl[128] vdd gnd cell_6t
Xbit_r129_c105 bl[105] br[105] wl[129] vdd gnd cell_6t
Xbit_r130_c105 bl[105] br[105] wl[130] vdd gnd cell_6t
Xbit_r131_c105 bl[105] br[105] wl[131] vdd gnd cell_6t
Xbit_r132_c105 bl[105] br[105] wl[132] vdd gnd cell_6t
Xbit_r133_c105 bl[105] br[105] wl[133] vdd gnd cell_6t
Xbit_r134_c105 bl[105] br[105] wl[134] vdd gnd cell_6t
Xbit_r135_c105 bl[105] br[105] wl[135] vdd gnd cell_6t
Xbit_r136_c105 bl[105] br[105] wl[136] vdd gnd cell_6t
Xbit_r137_c105 bl[105] br[105] wl[137] vdd gnd cell_6t
Xbit_r138_c105 bl[105] br[105] wl[138] vdd gnd cell_6t
Xbit_r139_c105 bl[105] br[105] wl[139] vdd gnd cell_6t
Xbit_r140_c105 bl[105] br[105] wl[140] vdd gnd cell_6t
Xbit_r141_c105 bl[105] br[105] wl[141] vdd gnd cell_6t
Xbit_r142_c105 bl[105] br[105] wl[142] vdd gnd cell_6t
Xbit_r143_c105 bl[105] br[105] wl[143] vdd gnd cell_6t
Xbit_r144_c105 bl[105] br[105] wl[144] vdd gnd cell_6t
Xbit_r145_c105 bl[105] br[105] wl[145] vdd gnd cell_6t
Xbit_r146_c105 bl[105] br[105] wl[146] vdd gnd cell_6t
Xbit_r147_c105 bl[105] br[105] wl[147] vdd gnd cell_6t
Xbit_r148_c105 bl[105] br[105] wl[148] vdd gnd cell_6t
Xbit_r149_c105 bl[105] br[105] wl[149] vdd gnd cell_6t
Xbit_r150_c105 bl[105] br[105] wl[150] vdd gnd cell_6t
Xbit_r151_c105 bl[105] br[105] wl[151] vdd gnd cell_6t
Xbit_r152_c105 bl[105] br[105] wl[152] vdd gnd cell_6t
Xbit_r153_c105 bl[105] br[105] wl[153] vdd gnd cell_6t
Xbit_r154_c105 bl[105] br[105] wl[154] vdd gnd cell_6t
Xbit_r155_c105 bl[105] br[105] wl[155] vdd gnd cell_6t
Xbit_r156_c105 bl[105] br[105] wl[156] vdd gnd cell_6t
Xbit_r157_c105 bl[105] br[105] wl[157] vdd gnd cell_6t
Xbit_r158_c105 bl[105] br[105] wl[158] vdd gnd cell_6t
Xbit_r159_c105 bl[105] br[105] wl[159] vdd gnd cell_6t
Xbit_r160_c105 bl[105] br[105] wl[160] vdd gnd cell_6t
Xbit_r161_c105 bl[105] br[105] wl[161] vdd gnd cell_6t
Xbit_r162_c105 bl[105] br[105] wl[162] vdd gnd cell_6t
Xbit_r163_c105 bl[105] br[105] wl[163] vdd gnd cell_6t
Xbit_r164_c105 bl[105] br[105] wl[164] vdd gnd cell_6t
Xbit_r165_c105 bl[105] br[105] wl[165] vdd gnd cell_6t
Xbit_r166_c105 bl[105] br[105] wl[166] vdd gnd cell_6t
Xbit_r167_c105 bl[105] br[105] wl[167] vdd gnd cell_6t
Xbit_r168_c105 bl[105] br[105] wl[168] vdd gnd cell_6t
Xbit_r169_c105 bl[105] br[105] wl[169] vdd gnd cell_6t
Xbit_r170_c105 bl[105] br[105] wl[170] vdd gnd cell_6t
Xbit_r171_c105 bl[105] br[105] wl[171] vdd gnd cell_6t
Xbit_r172_c105 bl[105] br[105] wl[172] vdd gnd cell_6t
Xbit_r173_c105 bl[105] br[105] wl[173] vdd gnd cell_6t
Xbit_r174_c105 bl[105] br[105] wl[174] vdd gnd cell_6t
Xbit_r175_c105 bl[105] br[105] wl[175] vdd gnd cell_6t
Xbit_r176_c105 bl[105] br[105] wl[176] vdd gnd cell_6t
Xbit_r177_c105 bl[105] br[105] wl[177] vdd gnd cell_6t
Xbit_r178_c105 bl[105] br[105] wl[178] vdd gnd cell_6t
Xbit_r179_c105 bl[105] br[105] wl[179] vdd gnd cell_6t
Xbit_r180_c105 bl[105] br[105] wl[180] vdd gnd cell_6t
Xbit_r181_c105 bl[105] br[105] wl[181] vdd gnd cell_6t
Xbit_r182_c105 bl[105] br[105] wl[182] vdd gnd cell_6t
Xbit_r183_c105 bl[105] br[105] wl[183] vdd gnd cell_6t
Xbit_r184_c105 bl[105] br[105] wl[184] vdd gnd cell_6t
Xbit_r185_c105 bl[105] br[105] wl[185] vdd gnd cell_6t
Xbit_r186_c105 bl[105] br[105] wl[186] vdd gnd cell_6t
Xbit_r187_c105 bl[105] br[105] wl[187] vdd gnd cell_6t
Xbit_r188_c105 bl[105] br[105] wl[188] vdd gnd cell_6t
Xbit_r189_c105 bl[105] br[105] wl[189] vdd gnd cell_6t
Xbit_r190_c105 bl[105] br[105] wl[190] vdd gnd cell_6t
Xbit_r191_c105 bl[105] br[105] wl[191] vdd gnd cell_6t
Xbit_r192_c105 bl[105] br[105] wl[192] vdd gnd cell_6t
Xbit_r193_c105 bl[105] br[105] wl[193] vdd gnd cell_6t
Xbit_r194_c105 bl[105] br[105] wl[194] vdd gnd cell_6t
Xbit_r195_c105 bl[105] br[105] wl[195] vdd gnd cell_6t
Xbit_r196_c105 bl[105] br[105] wl[196] vdd gnd cell_6t
Xbit_r197_c105 bl[105] br[105] wl[197] vdd gnd cell_6t
Xbit_r198_c105 bl[105] br[105] wl[198] vdd gnd cell_6t
Xbit_r199_c105 bl[105] br[105] wl[199] vdd gnd cell_6t
Xbit_r200_c105 bl[105] br[105] wl[200] vdd gnd cell_6t
Xbit_r201_c105 bl[105] br[105] wl[201] vdd gnd cell_6t
Xbit_r202_c105 bl[105] br[105] wl[202] vdd gnd cell_6t
Xbit_r203_c105 bl[105] br[105] wl[203] vdd gnd cell_6t
Xbit_r204_c105 bl[105] br[105] wl[204] vdd gnd cell_6t
Xbit_r205_c105 bl[105] br[105] wl[205] vdd gnd cell_6t
Xbit_r206_c105 bl[105] br[105] wl[206] vdd gnd cell_6t
Xbit_r207_c105 bl[105] br[105] wl[207] vdd gnd cell_6t
Xbit_r208_c105 bl[105] br[105] wl[208] vdd gnd cell_6t
Xbit_r209_c105 bl[105] br[105] wl[209] vdd gnd cell_6t
Xbit_r210_c105 bl[105] br[105] wl[210] vdd gnd cell_6t
Xbit_r211_c105 bl[105] br[105] wl[211] vdd gnd cell_6t
Xbit_r212_c105 bl[105] br[105] wl[212] vdd gnd cell_6t
Xbit_r213_c105 bl[105] br[105] wl[213] vdd gnd cell_6t
Xbit_r214_c105 bl[105] br[105] wl[214] vdd gnd cell_6t
Xbit_r215_c105 bl[105] br[105] wl[215] vdd gnd cell_6t
Xbit_r216_c105 bl[105] br[105] wl[216] vdd gnd cell_6t
Xbit_r217_c105 bl[105] br[105] wl[217] vdd gnd cell_6t
Xbit_r218_c105 bl[105] br[105] wl[218] vdd gnd cell_6t
Xbit_r219_c105 bl[105] br[105] wl[219] vdd gnd cell_6t
Xbit_r220_c105 bl[105] br[105] wl[220] vdd gnd cell_6t
Xbit_r221_c105 bl[105] br[105] wl[221] vdd gnd cell_6t
Xbit_r222_c105 bl[105] br[105] wl[222] vdd gnd cell_6t
Xbit_r223_c105 bl[105] br[105] wl[223] vdd gnd cell_6t
Xbit_r224_c105 bl[105] br[105] wl[224] vdd gnd cell_6t
Xbit_r225_c105 bl[105] br[105] wl[225] vdd gnd cell_6t
Xbit_r226_c105 bl[105] br[105] wl[226] vdd gnd cell_6t
Xbit_r227_c105 bl[105] br[105] wl[227] vdd gnd cell_6t
Xbit_r228_c105 bl[105] br[105] wl[228] vdd gnd cell_6t
Xbit_r229_c105 bl[105] br[105] wl[229] vdd gnd cell_6t
Xbit_r230_c105 bl[105] br[105] wl[230] vdd gnd cell_6t
Xbit_r231_c105 bl[105] br[105] wl[231] vdd gnd cell_6t
Xbit_r232_c105 bl[105] br[105] wl[232] vdd gnd cell_6t
Xbit_r233_c105 bl[105] br[105] wl[233] vdd gnd cell_6t
Xbit_r234_c105 bl[105] br[105] wl[234] vdd gnd cell_6t
Xbit_r235_c105 bl[105] br[105] wl[235] vdd gnd cell_6t
Xbit_r236_c105 bl[105] br[105] wl[236] vdd gnd cell_6t
Xbit_r237_c105 bl[105] br[105] wl[237] vdd gnd cell_6t
Xbit_r238_c105 bl[105] br[105] wl[238] vdd gnd cell_6t
Xbit_r239_c105 bl[105] br[105] wl[239] vdd gnd cell_6t
Xbit_r240_c105 bl[105] br[105] wl[240] vdd gnd cell_6t
Xbit_r241_c105 bl[105] br[105] wl[241] vdd gnd cell_6t
Xbit_r242_c105 bl[105] br[105] wl[242] vdd gnd cell_6t
Xbit_r243_c105 bl[105] br[105] wl[243] vdd gnd cell_6t
Xbit_r244_c105 bl[105] br[105] wl[244] vdd gnd cell_6t
Xbit_r245_c105 bl[105] br[105] wl[245] vdd gnd cell_6t
Xbit_r246_c105 bl[105] br[105] wl[246] vdd gnd cell_6t
Xbit_r247_c105 bl[105] br[105] wl[247] vdd gnd cell_6t
Xbit_r248_c105 bl[105] br[105] wl[248] vdd gnd cell_6t
Xbit_r249_c105 bl[105] br[105] wl[249] vdd gnd cell_6t
Xbit_r250_c105 bl[105] br[105] wl[250] vdd gnd cell_6t
Xbit_r251_c105 bl[105] br[105] wl[251] vdd gnd cell_6t
Xbit_r252_c105 bl[105] br[105] wl[252] vdd gnd cell_6t
Xbit_r253_c105 bl[105] br[105] wl[253] vdd gnd cell_6t
Xbit_r254_c105 bl[105] br[105] wl[254] vdd gnd cell_6t
Xbit_r255_c105 bl[105] br[105] wl[255] vdd gnd cell_6t
Xbit_r256_c105 bl[105] br[105] wl[256] vdd gnd cell_6t
Xbit_r257_c105 bl[105] br[105] wl[257] vdd gnd cell_6t
Xbit_r258_c105 bl[105] br[105] wl[258] vdd gnd cell_6t
Xbit_r259_c105 bl[105] br[105] wl[259] vdd gnd cell_6t
Xbit_r260_c105 bl[105] br[105] wl[260] vdd gnd cell_6t
Xbit_r261_c105 bl[105] br[105] wl[261] vdd gnd cell_6t
Xbit_r262_c105 bl[105] br[105] wl[262] vdd gnd cell_6t
Xbit_r263_c105 bl[105] br[105] wl[263] vdd gnd cell_6t
Xbit_r264_c105 bl[105] br[105] wl[264] vdd gnd cell_6t
Xbit_r265_c105 bl[105] br[105] wl[265] vdd gnd cell_6t
Xbit_r266_c105 bl[105] br[105] wl[266] vdd gnd cell_6t
Xbit_r267_c105 bl[105] br[105] wl[267] vdd gnd cell_6t
Xbit_r268_c105 bl[105] br[105] wl[268] vdd gnd cell_6t
Xbit_r269_c105 bl[105] br[105] wl[269] vdd gnd cell_6t
Xbit_r270_c105 bl[105] br[105] wl[270] vdd gnd cell_6t
Xbit_r271_c105 bl[105] br[105] wl[271] vdd gnd cell_6t
Xbit_r272_c105 bl[105] br[105] wl[272] vdd gnd cell_6t
Xbit_r273_c105 bl[105] br[105] wl[273] vdd gnd cell_6t
Xbit_r274_c105 bl[105] br[105] wl[274] vdd gnd cell_6t
Xbit_r275_c105 bl[105] br[105] wl[275] vdd gnd cell_6t
Xbit_r276_c105 bl[105] br[105] wl[276] vdd gnd cell_6t
Xbit_r277_c105 bl[105] br[105] wl[277] vdd gnd cell_6t
Xbit_r278_c105 bl[105] br[105] wl[278] vdd gnd cell_6t
Xbit_r279_c105 bl[105] br[105] wl[279] vdd gnd cell_6t
Xbit_r280_c105 bl[105] br[105] wl[280] vdd gnd cell_6t
Xbit_r281_c105 bl[105] br[105] wl[281] vdd gnd cell_6t
Xbit_r282_c105 bl[105] br[105] wl[282] vdd gnd cell_6t
Xbit_r283_c105 bl[105] br[105] wl[283] vdd gnd cell_6t
Xbit_r284_c105 bl[105] br[105] wl[284] vdd gnd cell_6t
Xbit_r285_c105 bl[105] br[105] wl[285] vdd gnd cell_6t
Xbit_r286_c105 bl[105] br[105] wl[286] vdd gnd cell_6t
Xbit_r287_c105 bl[105] br[105] wl[287] vdd gnd cell_6t
Xbit_r288_c105 bl[105] br[105] wl[288] vdd gnd cell_6t
Xbit_r289_c105 bl[105] br[105] wl[289] vdd gnd cell_6t
Xbit_r290_c105 bl[105] br[105] wl[290] vdd gnd cell_6t
Xbit_r291_c105 bl[105] br[105] wl[291] vdd gnd cell_6t
Xbit_r292_c105 bl[105] br[105] wl[292] vdd gnd cell_6t
Xbit_r293_c105 bl[105] br[105] wl[293] vdd gnd cell_6t
Xbit_r294_c105 bl[105] br[105] wl[294] vdd gnd cell_6t
Xbit_r295_c105 bl[105] br[105] wl[295] vdd gnd cell_6t
Xbit_r296_c105 bl[105] br[105] wl[296] vdd gnd cell_6t
Xbit_r297_c105 bl[105] br[105] wl[297] vdd gnd cell_6t
Xbit_r298_c105 bl[105] br[105] wl[298] vdd gnd cell_6t
Xbit_r299_c105 bl[105] br[105] wl[299] vdd gnd cell_6t
Xbit_r300_c105 bl[105] br[105] wl[300] vdd gnd cell_6t
Xbit_r301_c105 bl[105] br[105] wl[301] vdd gnd cell_6t
Xbit_r302_c105 bl[105] br[105] wl[302] vdd gnd cell_6t
Xbit_r303_c105 bl[105] br[105] wl[303] vdd gnd cell_6t
Xbit_r304_c105 bl[105] br[105] wl[304] vdd gnd cell_6t
Xbit_r305_c105 bl[105] br[105] wl[305] vdd gnd cell_6t
Xbit_r306_c105 bl[105] br[105] wl[306] vdd gnd cell_6t
Xbit_r307_c105 bl[105] br[105] wl[307] vdd gnd cell_6t
Xbit_r308_c105 bl[105] br[105] wl[308] vdd gnd cell_6t
Xbit_r309_c105 bl[105] br[105] wl[309] vdd gnd cell_6t
Xbit_r310_c105 bl[105] br[105] wl[310] vdd gnd cell_6t
Xbit_r311_c105 bl[105] br[105] wl[311] vdd gnd cell_6t
Xbit_r312_c105 bl[105] br[105] wl[312] vdd gnd cell_6t
Xbit_r313_c105 bl[105] br[105] wl[313] vdd gnd cell_6t
Xbit_r314_c105 bl[105] br[105] wl[314] vdd gnd cell_6t
Xbit_r315_c105 bl[105] br[105] wl[315] vdd gnd cell_6t
Xbit_r316_c105 bl[105] br[105] wl[316] vdd gnd cell_6t
Xbit_r317_c105 bl[105] br[105] wl[317] vdd gnd cell_6t
Xbit_r318_c105 bl[105] br[105] wl[318] vdd gnd cell_6t
Xbit_r319_c105 bl[105] br[105] wl[319] vdd gnd cell_6t
Xbit_r320_c105 bl[105] br[105] wl[320] vdd gnd cell_6t
Xbit_r321_c105 bl[105] br[105] wl[321] vdd gnd cell_6t
Xbit_r322_c105 bl[105] br[105] wl[322] vdd gnd cell_6t
Xbit_r323_c105 bl[105] br[105] wl[323] vdd gnd cell_6t
Xbit_r324_c105 bl[105] br[105] wl[324] vdd gnd cell_6t
Xbit_r325_c105 bl[105] br[105] wl[325] vdd gnd cell_6t
Xbit_r326_c105 bl[105] br[105] wl[326] vdd gnd cell_6t
Xbit_r327_c105 bl[105] br[105] wl[327] vdd gnd cell_6t
Xbit_r328_c105 bl[105] br[105] wl[328] vdd gnd cell_6t
Xbit_r329_c105 bl[105] br[105] wl[329] vdd gnd cell_6t
Xbit_r330_c105 bl[105] br[105] wl[330] vdd gnd cell_6t
Xbit_r331_c105 bl[105] br[105] wl[331] vdd gnd cell_6t
Xbit_r332_c105 bl[105] br[105] wl[332] vdd gnd cell_6t
Xbit_r333_c105 bl[105] br[105] wl[333] vdd gnd cell_6t
Xbit_r334_c105 bl[105] br[105] wl[334] vdd gnd cell_6t
Xbit_r335_c105 bl[105] br[105] wl[335] vdd gnd cell_6t
Xbit_r336_c105 bl[105] br[105] wl[336] vdd gnd cell_6t
Xbit_r337_c105 bl[105] br[105] wl[337] vdd gnd cell_6t
Xbit_r338_c105 bl[105] br[105] wl[338] vdd gnd cell_6t
Xbit_r339_c105 bl[105] br[105] wl[339] vdd gnd cell_6t
Xbit_r340_c105 bl[105] br[105] wl[340] vdd gnd cell_6t
Xbit_r341_c105 bl[105] br[105] wl[341] vdd gnd cell_6t
Xbit_r342_c105 bl[105] br[105] wl[342] vdd gnd cell_6t
Xbit_r343_c105 bl[105] br[105] wl[343] vdd gnd cell_6t
Xbit_r344_c105 bl[105] br[105] wl[344] vdd gnd cell_6t
Xbit_r345_c105 bl[105] br[105] wl[345] vdd gnd cell_6t
Xbit_r346_c105 bl[105] br[105] wl[346] vdd gnd cell_6t
Xbit_r347_c105 bl[105] br[105] wl[347] vdd gnd cell_6t
Xbit_r348_c105 bl[105] br[105] wl[348] vdd gnd cell_6t
Xbit_r349_c105 bl[105] br[105] wl[349] vdd gnd cell_6t
Xbit_r350_c105 bl[105] br[105] wl[350] vdd gnd cell_6t
Xbit_r351_c105 bl[105] br[105] wl[351] vdd gnd cell_6t
Xbit_r352_c105 bl[105] br[105] wl[352] vdd gnd cell_6t
Xbit_r353_c105 bl[105] br[105] wl[353] vdd gnd cell_6t
Xbit_r354_c105 bl[105] br[105] wl[354] vdd gnd cell_6t
Xbit_r355_c105 bl[105] br[105] wl[355] vdd gnd cell_6t
Xbit_r356_c105 bl[105] br[105] wl[356] vdd gnd cell_6t
Xbit_r357_c105 bl[105] br[105] wl[357] vdd gnd cell_6t
Xbit_r358_c105 bl[105] br[105] wl[358] vdd gnd cell_6t
Xbit_r359_c105 bl[105] br[105] wl[359] vdd gnd cell_6t
Xbit_r360_c105 bl[105] br[105] wl[360] vdd gnd cell_6t
Xbit_r361_c105 bl[105] br[105] wl[361] vdd gnd cell_6t
Xbit_r362_c105 bl[105] br[105] wl[362] vdd gnd cell_6t
Xbit_r363_c105 bl[105] br[105] wl[363] vdd gnd cell_6t
Xbit_r364_c105 bl[105] br[105] wl[364] vdd gnd cell_6t
Xbit_r365_c105 bl[105] br[105] wl[365] vdd gnd cell_6t
Xbit_r366_c105 bl[105] br[105] wl[366] vdd gnd cell_6t
Xbit_r367_c105 bl[105] br[105] wl[367] vdd gnd cell_6t
Xbit_r368_c105 bl[105] br[105] wl[368] vdd gnd cell_6t
Xbit_r369_c105 bl[105] br[105] wl[369] vdd gnd cell_6t
Xbit_r370_c105 bl[105] br[105] wl[370] vdd gnd cell_6t
Xbit_r371_c105 bl[105] br[105] wl[371] vdd gnd cell_6t
Xbit_r372_c105 bl[105] br[105] wl[372] vdd gnd cell_6t
Xbit_r373_c105 bl[105] br[105] wl[373] vdd gnd cell_6t
Xbit_r374_c105 bl[105] br[105] wl[374] vdd gnd cell_6t
Xbit_r375_c105 bl[105] br[105] wl[375] vdd gnd cell_6t
Xbit_r376_c105 bl[105] br[105] wl[376] vdd gnd cell_6t
Xbit_r377_c105 bl[105] br[105] wl[377] vdd gnd cell_6t
Xbit_r378_c105 bl[105] br[105] wl[378] vdd gnd cell_6t
Xbit_r379_c105 bl[105] br[105] wl[379] vdd gnd cell_6t
Xbit_r380_c105 bl[105] br[105] wl[380] vdd gnd cell_6t
Xbit_r381_c105 bl[105] br[105] wl[381] vdd gnd cell_6t
Xbit_r382_c105 bl[105] br[105] wl[382] vdd gnd cell_6t
Xbit_r383_c105 bl[105] br[105] wl[383] vdd gnd cell_6t
Xbit_r384_c105 bl[105] br[105] wl[384] vdd gnd cell_6t
Xbit_r385_c105 bl[105] br[105] wl[385] vdd gnd cell_6t
Xbit_r386_c105 bl[105] br[105] wl[386] vdd gnd cell_6t
Xbit_r387_c105 bl[105] br[105] wl[387] vdd gnd cell_6t
Xbit_r388_c105 bl[105] br[105] wl[388] vdd gnd cell_6t
Xbit_r389_c105 bl[105] br[105] wl[389] vdd gnd cell_6t
Xbit_r390_c105 bl[105] br[105] wl[390] vdd gnd cell_6t
Xbit_r391_c105 bl[105] br[105] wl[391] vdd gnd cell_6t
Xbit_r392_c105 bl[105] br[105] wl[392] vdd gnd cell_6t
Xbit_r393_c105 bl[105] br[105] wl[393] vdd gnd cell_6t
Xbit_r394_c105 bl[105] br[105] wl[394] vdd gnd cell_6t
Xbit_r395_c105 bl[105] br[105] wl[395] vdd gnd cell_6t
Xbit_r396_c105 bl[105] br[105] wl[396] vdd gnd cell_6t
Xbit_r397_c105 bl[105] br[105] wl[397] vdd gnd cell_6t
Xbit_r398_c105 bl[105] br[105] wl[398] vdd gnd cell_6t
Xbit_r399_c105 bl[105] br[105] wl[399] vdd gnd cell_6t
Xbit_r400_c105 bl[105] br[105] wl[400] vdd gnd cell_6t
Xbit_r401_c105 bl[105] br[105] wl[401] vdd gnd cell_6t
Xbit_r402_c105 bl[105] br[105] wl[402] vdd gnd cell_6t
Xbit_r403_c105 bl[105] br[105] wl[403] vdd gnd cell_6t
Xbit_r404_c105 bl[105] br[105] wl[404] vdd gnd cell_6t
Xbit_r405_c105 bl[105] br[105] wl[405] vdd gnd cell_6t
Xbit_r406_c105 bl[105] br[105] wl[406] vdd gnd cell_6t
Xbit_r407_c105 bl[105] br[105] wl[407] vdd gnd cell_6t
Xbit_r408_c105 bl[105] br[105] wl[408] vdd gnd cell_6t
Xbit_r409_c105 bl[105] br[105] wl[409] vdd gnd cell_6t
Xbit_r410_c105 bl[105] br[105] wl[410] vdd gnd cell_6t
Xbit_r411_c105 bl[105] br[105] wl[411] vdd gnd cell_6t
Xbit_r412_c105 bl[105] br[105] wl[412] vdd gnd cell_6t
Xbit_r413_c105 bl[105] br[105] wl[413] vdd gnd cell_6t
Xbit_r414_c105 bl[105] br[105] wl[414] vdd gnd cell_6t
Xbit_r415_c105 bl[105] br[105] wl[415] vdd gnd cell_6t
Xbit_r416_c105 bl[105] br[105] wl[416] vdd gnd cell_6t
Xbit_r417_c105 bl[105] br[105] wl[417] vdd gnd cell_6t
Xbit_r418_c105 bl[105] br[105] wl[418] vdd gnd cell_6t
Xbit_r419_c105 bl[105] br[105] wl[419] vdd gnd cell_6t
Xbit_r420_c105 bl[105] br[105] wl[420] vdd gnd cell_6t
Xbit_r421_c105 bl[105] br[105] wl[421] vdd gnd cell_6t
Xbit_r422_c105 bl[105] br[105] wl[422] vdd gnd cell_6t
Xbit_r423_c105 bl[105] br[105] wl[423] vdd gnd cell_6t
Xbit_r424_c105 bl[105] br[105] wl[424] vdd gnd cell_6t
Xbit_r425_c105 bl[105] br[105] wl[425] vdd gnd cell_6t
Xbit_r426_c105 bl[105] br[105] wl[426] vdd gnd cell_6t
Xbit_r427_c105 bl[105] br[105] wl[427] vdd gnd cell_6t
Xbit_r428_c105 bl[105] br[105] wl[428] vdd gnd cell_6t
Xbit_r429_c105 bl[105] br[105] wl[429] vdd gnd cell_6t
Xbit_r430_c105 bl[105] br[105] wl[430] vdd gnd cell_6t
Xbit_r431_c105 bl[105] br[105] wl[431] vdd gnd cell_6t
Xbit_r432_c105 bl[105] br[105] wl[432] vdd gnd cell_6t
Xbit_r433_c105 bl[105] br[105] wl[433] vdd gnd cell_6t
Xbit_r434_c105 bl[105] br[105] wl[434] vdd gnd cell_6t
Xbit_r435_c105 bl[105] br[105] wl[435] vdd gnd cell_6t
Xbit_r436_c105 bl[105] br[105] wl[436] vdd gnd cell_6t
Xbit_r437_c105 bl[105] br[105] wl[437] vdd gnd cell_6t
Xbit_r438_c105 bl[105] br[105] wl[438] vdd gnd cell_6t
Xbit_r439_c105 bl[105] br[105] wl[439] vdd gnd cell_6t
Xbit_r440_c105 bl[105] br[105] wl[440] vdd gnd cell_6t
Xbit_r441_c105 bl[105] br[105] wl[441] vdd gnd cell_6t
Xbit_r442_c105 bl[105] br[105] wl[442] vdd gnd cell_6t
Xbit_r443_c105 bl[105] br[105] wl[443] vdd gnd cell_6t
Xbit_r444_c105 bl[105] br[105] wl[444] vdd gnd cell_6t
Xbit_r445_c105 bl[105] br[105] wl[445] vdd gnd cell_6t
Xbit_r446_c105 bl[105] br[105] wl[446] vdd gnd cell_6t
Xbit_r447_c105 bl[105] br[105] wl[447] vdd gnd cell_6t
Xbit_r448_c105 bl[105] br[105] wl[448] vdd gnd cell_6t
Xbit_r449_c105 bl[105] br[105] wl[449] vdd gnd cell_6t
Xbit_r450_c105 bl[105] br[105] wl[450] vdd gnd cell_6t
Xbit_r451_c105 bl[105] br[105] wl[451] vdd gnd cell_6t
Xbit_r452_c105 bl[105] br[105] wl[452] vdd gnd cell_6t
Xbit_r453_c105 bl[105] br[105] wl[453] vdd gnd cell_6t
Xbit_r454_c105 bl[105] br[105] wl[454] vdd gnd cell_6t
Xbit_r455_c105 bl[105] br[105] wl[455] vdd gnd cell_6t
Xbit_r456_c105 bl[105] br[105] wl[456] vdd gnd cell_6t
Xbit_r457_c105 bl[105] br[105] wl[457] vdd gnd cell_6t
Xbit_r458_c105 bl[105] br[105] wl[458] vdd gnd cell_6t
Xbit_r459_c105 bl[105] br[105] wl[459] vdd gnd cell_6t
Xbit_r460_c105 bl[105] br[105] wl[460] vdd gnd cell_6t
Xbit_r461_c105 bl[105] br[105] wl[461] vdd gnd cell_6t
Xbit_r462_c105 bl[105] br[105] wl[462] vdd gnd cell_6t
Xbit_r463_c105 bl[105] br[105] wl[463] vdd gnd cell_6t
Xbit_r464_c105 bl[105] br[105] wl[464] vdd gnd cell_6t
Xbit_r465_c105 bl[105] br[105] wl[465] vdd gnd cell_6t
Xbit_r466_c105 bl[105] br[105] wl[466] vdd gnd cell_6t
Xbit_r467_c105 bl[105] br[105] wl[467] vdd gnd cell_6t
Xbit_r468_c105 bl[105] br[105] wl[468] vdd gnd cell_6t
Xbit_r469_c105 bl[105] br[105] wl[469] vdd gnd cell_6t
Xbit_r470_c105 bl[105] br[105] wl[470] vdd gnd cell_6t
Xbit_r471_c105 bl[105] br[105] wl[471] vdd gnd cell_6t
Xbit_r472_c105 bl[105] br[105] wl[472] vdd gnd cell_6t
Xbit_r473_c105 bl[105] br[105] wl[473] vdd gnd cell_6t
Xbit_r474_c105 bl[105] br[105] wl[474] vdd gnd cell_6t
Xbit_r475_c105 bl[105] br[105] wl[475] vdd gnd cell_6t
Xbit_r476_c105 bl[105] br[105] wl[476] vdd gnd cell_6t
Xbit_r477_c105 bl[105] br[105] wl[477] vdd gnd cell_6t
Xbit_r478_c105 bl[105] br[105] wl[478] vdd gnd cell_6t
Xbit_r479_c105 bl[105] br[105] wl[479] vdd gnd cell_6t
Xbit_r480_c105 bl[105] br[105] wl[480] vdd gnd cell_6t
Xbit_r481_c105 bl[105] br[105] wl[481] vdd gnd cell_6t
Xbit_r482_c105 bl[105] br[105] wl[482] vdd gnd cell_6t
Xbit_r483_c105 bl[105] br[105] wl[483] vdd gnd cell_6t
Xbit_r484_c105 bl[105] br[105] wl[484] vdd gnd cell_6t
Xbit_r485_c105 bl[105] br[105] wl[485] vdd gnd cell_6t
Xbit_r486_c105 bl[105] br[105] wl[486] vdd gnd cell_6t
Xbit_r487_c105 bl[105] br[105] wl[487] vdd gnd cell_6t
Xbit_r488_c105 bl[105] br[105] wl[488] vdd gnd cell_6t
Xbit_r489_c105 bl[105] br[105] wl[489] vdd gnd cell_6t
Xbit_r490_c105 bl[105] br[105] wl[490] vdd gnd cell_6t
Xbit_r491_c105 bl[105] br[105] wl[491] vdd gnd cell_6t
Xbit_r492_c105 bl[105] br[105] wl[492] vdd gnd cell_6t
Xbit_r493_c105 bl[105] br[105] wl[493] vdd gnd cell_6t
Xbit_r494_c105 bl[105] br[105] wl[494] vdd gnd cell_6t
Xbit_r495_c105 bl[105] br[105] wl[495] vdd gnd cell_6t
Xbit_r496_c105 bl[105] br[105] wl[496] vdd gnd cell_6t
Xbit_r497_c105 bl[105] br[105] wl[497] vdd gnd cell_6t
Xbit_r498_c105 bl[105] br[105] wl[498] vdd gnd cell_6t
Xbit_r499_c105 bl[105] br[105] wl[499] vdd gnd cell_6t
Xbit_r500_c105 bl[105] br[105] wl[500] vdd gnd cell_6t
Xbit_r501_c105 bl[105] br[105] wl[501] vdd gnd cell_6t
Xbit_r502_c105 bl[105] br[105] wl[502] vdd gnd cell_6t
Xbit_r503_c105 bl[105] br[105] wl[503] vdd gnd cell_6t
Xbit_r504_c105 bl[105] br[105] wl[504] vdd gnd cell_6t
Xbit_r505_c105 bl[105] br[105] wl[505] vdd gnd cell_6t
Xbit_r506_c105 bl[105] br[105] wl[506] vdd gnd cell_6t
Xbit_r507_c105 bl[105] br[105] wl[507] vdd gnd cell_6t
Xbit_r508_c105 bl[105] br[105] wl[508] vdd gnd cell_6t
Xbit_r509_c105 bl[105] br[105] wl[509] vdd gnd cell_6t
Xbit_r510_c105 bl[105] br[105] wl[510] vdd gnd cell_6t
Xbit_r511_c105 bl[105] br[105] wl[511] vdd gnd cell_6t
Xbit_r0_c106 bl[106] br[106] wl[0] vdd gnd cell_6t
Xbit_r1_c106 bl[106] br[106] wl[1] vdd gnd cell_6t
Xbit_r2_c106 bl[106] br[106] wl[2] vdd gnd cell_6t
Xbit_r3_c106 bl[106] br[106] wl[3] vdd gnd cell_6t
Xbit_r4_c106 bl[106] br[106] wl[4] vdd gnd cell_6t
Xbit_r5_c106 bl[106] br[106] wl[5] vdd gnd cell_6t
Xbit_r6_c106 bl[106] br[106] wl[6] vdd gnd cell_6t
Xbit_r7_c106 bl[106] br[106] wl[7] vdd gnd cell_6t
Xbit_r8_c106 bl[106] br[106] wl[8] vdd gnd cell_6t
Xbit_r9_c106 bl[106] br[106] wl[9] vdd gnd cell_6t
Xbit_r10_c106 bl[106] br[106] wl[10] vdd gnd cell_6t
Xbit_r11_c106 bl[106] br[106] wl[11] vdd gnd cell_6t
Xbit_r12_c106 bl[106] br[106] wl[12] vdd gnd cell_6t
Xbit_r13_c106 bl[106] br[106] wl[13] vdd gnd cell_6t
Xbit_r14_c106 bl[106] br[106] wl[14] vdd gnd cell_6t
Xbit_r15_c106 bl[106] br[106] wl[15] vdd gnd cell_6t
Xbit_r16_c106 bl[106] br[106] wl[16] vdd gnd cell_6t
Xbit_r17_c106 bl[106] br[106] wl[17] vdd gnd cell_6t
Xbit_r18_c106 bl[106] br[106] wl[18] vdd gnd cell_6t
Xbit_r19_c106 bl[106] br[106] wl[19] vdd gnd cell_6t
Xbit_r20_c106 bl[106] br[106] wl[20] vdd gnd cell_6t
Xbit_r21_c106 bl[106] br[106] wl[21] vdd gnd cell_6t
Xbit_r22_c106 bl[106] br[106] wl[22] vdd gnd cell_6t
Xbit_r23_c106 bl[106] br[106] wl[23] vdd gnd cell_6t
Xbit_r24_c106 bl[106] br[106] wl[24] vdd gnd cell_6t
Xbit_r25_c106 bl[106] br[106] wl[25] vdd gnd cell_6t
Xbit_r26_c106 bl[106] br[106] wl[26] vdd gnd cell_6t
Xbit_r27_c106 bl[106] br[106] wl[27] vdd gnd cell_6t
Xbit_r28_c106 bl[106] br[106] wl[28] vdd gnd cell_6t
Xbit_r29_c106 bl[106] br[106] wl[29] vdd gnd cell_6t
Xbit_r30_c106 bl[106] br[106] wl[30] vdd gnd cell_6t
Xbit_r31_c106 bl[106] br[106] wl[31] vdd gnd cell_6t
Xbit_r32_c106 bl[106] br[106] wl[32] vdd gnd cell_6t
Xbit_r33_c106 bl[106] br[106] wl[33] vdd gnd cell_6t
Xbit_r34_c106 bl[106] br[106] wl[34] vdd gnd cell_6t
Xbit_r35_c106 bl[106] br[106] wl[35] vdd gnd cell_6t
Xbit_r36_c106 bl[106] br[106] wl[36] vdd gnd cell_6t
Xbit_r37_c106 bl[106] br[106] wl[37] vdd gnd cell_6t
Xbit_r38_c106 bl[106] br[106] wl[38] vdd gnd cell_6t
Xbit_r39_c106 bl[106] br[106] wl[39] vdd gnd cell_6t
Xbit_r40_c106 bl[106] br[106] wl[40] vdd gnd cell_6t
Xbit_r41_c106 bl[106] br[106] wl[41] vdd gnd cell_6t
Xbit_r42_c106 bl[106] br[106] wl[42] vdd gnd cell_6t
Xbit_r43_c106 bl[106] br[106] wl[43] vdd gnd cell_6t
Xbit_r44_c106 bl[106] br[106] wl[44] vdd gnd cell_6t
Xbit_r45_c106 bl[106] br[106] wl[45] vdd gnd cell_6t
Xbit_r46_c106 bl[106] br[106] wl[46] vdd gnd cell_6t
Xbit_r47_c106 bl[106] br[106] wl[47] vdd gnd cell_6t
Xbit_r48_c106 bl[106] br[106] wl[48] vdd gnd cell_6t
Xbit_r49_c106 bl[106] br[106] wl[49] vdd gnd cell_6t
Xbit_r50_c106 bl[106] br[106] wl[50] vdd gnd cell_6t
Xbit_r51_c106 bl[106] br[106] wl[51] vdd gnd cell_6t
Xbit_r52_c106 bl[106] br[106] wl[52] vdd gnd cell_6t
Xbit_r53_c106 bl[106] br[106] wl[53] vdd gnd cell_6t
Xbit_r54_c106 bl[106] br[106] wl[54] vdd gnd cell_6t
Xbit_r55_c106 bl[106] br[106] wl[55] vdd gnd cell_6t
Xbit_r56_c106 bl[106] br[106] wl[56] vdd gnd cell_6t
Xbit_r57_c106 bl[106] br[106] wl[57] vdd gnd cell_6t
Xbit_r58_c106 bl[106] br[106] wl[58] vdd gnd cell_6t
Xbit_r59_c106 bl[106] br[106] wl[59] vdd gnd cell_6t
Xbit_r60_c106 bl[106] br[106] wl[60] vdd gnd cell_6t
Xbit_r61_c106 bl[106] br[106] wl[61] vdd gnd cell_6t
Xbit_r62_c106 bl[106] br[106] wl[62] vdd gnd cell_6t
Xbit_r63_c106 bl[106] br[106] wl[63] vdd gnd cell_6t
Xbit_r64_c106 bl[106] br[106] wl[64] vdd gnd cell_6t
Xbit_r65_c106 bl[106] br[106] wl[65] vdd gnd cell_6t
Xbit_r66_c106 bl[106] br[106] wl[66] vdd gnd cell_6t
Xbit_r67_c106 bl[106] br[106] wl[67] vdd gnd cell_6t
Xbit_r68_c106 bl[106] br[106] wl[68] vdd gnd cell_6t
Xbit_r69_c106 bl[106] br[106] wl[69] vdd gnd cell_6t
Xbit_r70_c106 bl[106] br[106] wl[70] vdd gnd cell_6t
Xbit_r71_c106 bl[106] br[106] wl[71] vdd gnd cell_6t
Xbit_r72_c106 bl[106] br[106] wl[72] vdd gnd cell_6t
Xbit_r73_c106 bl[106] br[106] wl[73] vdd gnd cell_6t
Xbit_r74_c106 bl[106] br[106] wl[74] vdd gnd cell_6t
Xbit_r75_c106 bl[106] br[106] wl[75] vdd gnd cell_6t
Xbit_r76_c106 bl[106] br[106] wl[76] vdd gnd cell_6t
Xbit_r77_c106 bl[106] br[106] wl[77] vdd gnd cell_6t
Xbit_r78_c106 bl[106] br[106] wl[78] vdd gnd cell_6t
Xbit_r79_c106 bl[106] br[106] wl[79] vdd gnd cell_6t
Xbit_r80_c106 bl[106] br[106] wl[80] vdd gnd cell_6t
Xbit_r81_c106 bl[106] br[106] wl[81] vdd gnd cell_6t
Xbit_r82_c106 bl[106] br[106] wl[82] vdd gnd cell_6t
Xbit_r83_c106 bl[106] br[106] wl[83] vdd gnd cell_6t
Xbit_r84_c106 bl[106] br[106] wl[84] vdd gnd cell_6t
Xbit_r85_c106 bl[106] br[106] wl[85] vdd gnd cell_6t
Xbit_r86_c106 bl[106] br[106] wl[86] vdd gnd cell_6t
Xbit_r87_c106 bl[106] br[106] wl[87] vdd gnd cell_6t
Xbit_r88_c106 bl[106] br[106] wl[88] vdd gnd cell_6t
Xbit_r89_c106 bl[106] br[106] wl[89] vdd gnd cell_6t
Xbit_r90_c106 bl[106] br[106] wl[90] vdd gnd cell_6t
Xbit_r91_c106 bl[106] br[106] wl[91] vdd gnd cell_6t
Xbit_r92_c106 bl[106] br[106] wl[92] vdd gnd cell_6t
Xbit_r93_c106 bl[106] br[106] wl[93] vdd gnd cell_6t
Xbit_r94_c106 bl[106] br[106] wl[94] vdd gnd cell_6t
Xbit_r95_c106 bl[106] br[106] wl[95] vdd gnd cell_6t
Xbit_r96_c106 bl[106] br[106] wl[96] vdd gnd cell_6t
Xbit_r97_c106 bl[106] br[106] wl[97] vdd gnd cell_6t
Xbit_r98_c106 bl[106] br[106] wl[98] vdd gnd cell_6t
Xbit_r99_c106 bl[106] br[106] wl[99] vdd gnd cell_6t
Xbit_r100_c106 bl[106] br[106] wl[100] vdd gnd cell_6t
Xbit_r101_c106 bl[106] br[106] wl[101] vdd gnd cell_6t
Xbit_r102_c106 bl[106] br[106] wl[102] vdd gnd cell_6t
Xbit_r103_c106 bl[106] br[106] wl[103] vdd gnd cell_6t
Xbit_r104_c106 bl[106] br[106] wl[104] vdd gnd cell_6t
Xbit_r105_c106 bl[106] br[106] wl[105] vdd gnd cell_6t
Xbit_r106_c106 bl[106] br[106] wl[106] vdd gnd cell_6t
Xbit_r107_c106 bl[106] br[106] wl[107] vdd gnd cell_6t
Xbit_r108_c106 bl[106] br[106] wl[108] vdd gnd cell_6t
Xbit_r109_c106 bl[106] br[106] wl[109] vdd gnd cell_6t
Xbit_r110_c106 bl[106] br[106] wl[110] vdd gnd cell_6t
Xbit_r111_c106 bl[106] br[106] wl[111] vdd gnd cell_6t
Xbit_r112_c106 bl[106] br[106] wl[112] vdd gnd cell_6t
Xbit_r113_c106 bl[106] br[106] wl[113] vdd gnd cell_6t
Xbit_r114_c106 bl[106] br[106] wl[114] vdd gnd cell_6t
Xbit_r115_c106 bl[106] br[106] wl[115] vdd gnd cell_6t
Xbit_r116_c106 bl[106] br[106] wl[116] vdd gnd cell_6t
Xbit_r117_c106 bl[106] br[106] wl[117] vdd gnd cell_6t
Xbit_r118_c106 bl[106] br[106] wl[118] vdd gnd cell_6t
Xbit_r119_c106 bl[106] br[106] wl[119] vdd gnd cell_6t
Xbit_r120_c106 bl[106] br[106] wl[120] vdd gnd cell_6t
Xbit_r121_c106 bl[106] br[106] wl[121] vdd gnd cell_6t
Xbit_r122_c106 bl[106] br[106] wl[122] vdd gnd cell_6t
Xbit_r123_c106 bl[106] br[106] wl[123] vdd gnd cell_6t
Xbit_r124_c106 bl[106] br[106] wl[124] vdd gnd cell_6t
Xbit_r125_c106 bl[106] br[106] wl[125] vdd gnd cell_6t
Xbit_r126_c106 bl[106] br[106] wl[126] vdd gnd cell_6t
Xbit_r127_c106 bl[106] br[106] wl[127] vdd gnd cell_6t
Xbit_r128_c106 bl[106] br[106] wl[128] vdd gnd cell_6t
Xbit_r129_c106 bl[106] br[106] wl[129] vdd gnd cell_6t
Xbit_r130_c106 bl[106] br[106] wl[130] vdd gnd cell_6t
Xbit_r131_c106 bl[106] br[106] wl[131] vdd gnd cell_6t
Xbit_r132_c106 bl[106] br[106] wl[132] vdd gnd cell_6t
Xbit_r133_c106 bl[106] br[106] wl[133] vdd gnd cell_6t
Xbit_r134_c106 bl[106] br[106] wl[134] vdd gnd cell_6t
Xbit_r135_c106 bl[106] br[106] wl[135] vdd gnd cell_6t
Xbit_r136_c106 bl[106] br[106] wl[136] vdd gnd cell_6t
Xbit_r137_c106 bl[106] br[106] wl[137] vdd gnd cell_6t
Xbit_r138_c106 bl[106] br[106] wl[138] vdd gnd cell_6t
Xbit_r139_c106 bl[106] br[106] wl[139] vdd gnd cell_6t
Xbit_r140_c106 bl[106] br[106] wl[140] vdd gnd cell_6t
Xbit_r141_c106 bl[106] br[106] wl[141] vdd gnd cell_6t
Xbit_r142_c106 bl[106] br[106] wl[142] vdd gnd cell_6t
Xbit_r143_c106 bl[106] br[106] wl[143] vdd gnd cell_6t
Xbit_r144_c106 bl[106] br[106] wl[144] vdd gnd cell_6t
Xbit_r145_c106 bl[106] br[106] wl[145] vdd gnd cell_6t
Xbit_r146_c106 bl[106] br[106] wl[146] vdd gnd cell_6t
Xbit_r147_c106 bl[106] br[106] wl[147] vdd gnd cell_6t
Xbit_r148_c106 bl[106] br[106] wl[148] vdd gnd cell_6t
Xbit_r149_c106 bl[106] br[106] wl[149] vdd gnd cell_6t
Xbit_r150_c106 bl[106] br[106] wl[150] vdd gnd cell_6t
Xbit_r151_c106 bl[106] br[106] wl[151] vdd gnd cell_6t
Xbit_r152_c106 bl[106] br[106] wl[152] vdd gnd cell_6t
Xbit_r153_c106 bl[106] br[106] wl[153] vdd gnd cell_6t
Xbit_r154_c106 bl[106] br[106] wl[154] vdd gnd cell_6t
Xbit_r155_c106 bl[106] br[106] wl[155] vdd gnd cell_6t
Xbit_r156_c106 bl[106] br[106] wl[156] vdd gnd cell_6t
Xbit_r157_c106 bl[106] br[106] wl[157] vdd gnd cell_6t
Xbit_r158_c106 bl[106] br[106] wl[158] vdd gnd cell_6t
Xbit_r159_c106 bl[106] br[106] wl[159] vdd gnd cell_6t
Xbit_r160_c106 bl[106] br[106] wl[160] vdd gnd cell_6t
Xbit_r161_c106 bl[106] br[106] wl[161] vdd gnd cell_6t
Xbit_r162_c106 bl[106] br[106] wl[162] vdd gnd cell_6t
Xbit_r163_c106 bl[106] br[106] wl[163] vdd gnd cell_6t
Xbit_r164_c106 bl[106] br[106] wl[164] vdd gnd cell_6t
Xbit_r165_c106 bl[106] br[106] wl[165] vdd gnd cell_6t
Xbit_r166_c106 bl[106] br[106] wl[166] vdd gnd cell_6t
Xbit_r167_c106 bl[106] br[106] wl[167] vdd gnd cell_6t
Xbit_r168_c106 bl[106] br[106] wl[168] vdd gnd cell_6t
Xbit_r169_c106 bl[106] br[106] wl[169] vdd gnd cell_6t
Xbit_r170_c106 bl[106] br[106] wl[170] vdd gnd cell_6t
Xbit_r171_c106 bl[106] br[106] wl[171] vdd gnd cell_6t
Xbit_r172_c106 bl[106] br[106] wl[172] vdd gnd cell_6t
Xbit_r173_c106 bl[106] br[106] wl[173] vdd gnd cell_6t
Xbit_r174_c106 bl[106] br[106] wl[174] vdd gnd cell_6t
Xbit_r175_c106 bl[106] br[106] wl[175] vdd gnd cell_6t
Xbit_r176_c106 bl[106] br[106] wl[176] vdd gnd cell_6t
Xbit_r177_c106 bl[106] br[106] wl[177] vdd gnd cell_6t
Xbit_r178_c106 bl[106] br[106] wl[178] vdd gnd cell_6t
Xbit_r179_c106 bl[106] br[106] wl[179] vdd gnd cell_6t
Xbit_r180_c106 bl[106] br[106] wl[180] vdd gnd cell_6t
Xbit_r181_c106 bl[106] br[106] wl[181] vdd gnd cell_6t
Xbit_r182_c106 bl[106] br[106] wl[182] vdd gnd cell_6t
Xbit_r183_c106 bl[106] br[106] wl[183] vdd gnd cell_6t
Xbit_r184_c106 bl[106] br[106] wl[184] vdd gnd cell_6t
Xbit_r185_c106 bl[106] br[106] wl[185] vdd gnd cell_6t
Xbit_r186_c106 bl[106] br[106] wl[186] vdd gnd cell_6t
Xbit_r187_c106 bl[106] br[106] wl[187] vdd gnd cell_6t
Xbit_r188_c106 bl[106] br[106] wl[188] vdd gnd cell_6t
Xbit_r189_c106 bl[106] br[106] wl[189] vdd gnd cell_6t
Xbit_r190_c106 bl[106] br[106] wl[190] vdd gnd cell_6t
Xbit_r191_c106 bl[106] br[106] wl[191] vdd gnd cell_6t
Xbit_r192_c106 bl[106] br[106] wl[192] vdd gnd cell_6t
Xbit_r193_c106 bl[106] br[106] wl[193] vdd gnd cell_6t
Xbit_r194_c106 bl[106] br[106] wl[194] vdd gnd cell_6t
Xbit_r195_c106 bl[106] br[106] wl[195] vdd gnd cell_6t
Xbit_r196_c106 bl[106] br[106] wl[196] vdd gnd cell_6t
Xbit_r197_c106 bl[106] br[106] wl[197] vdd gnd cell_6t
Xbit_r198_c106 bl[106] br[106] wl[198] vdd gnd cell_6t
Xbit_r199_c106 bl[106] br[106] wl[199] vdd gnd cell_6t
Xbit_r200_c106 bl[106] br[106] wl[200] vdd gnd cell_6t
Xbit_r201_c106 bl[106] br[106] wl[201] vdd gnd cell_6t
Xbit_r202_c106 bl[106] br[106] wl[202] vdd gnd cell_6t
Xbit_r203_c106 bl[106] br[106] wl[203] vdd gnd cell_6t
Xbit_r204_c106 bl[106] br[106] wl[204] vdd gnd cell_6t
Xbit_r205_c106 bl[106] br[106] wl[205] vdd gnd cell_6t
Xbit_r206_c106 bl[106] br[106] wl[206] vdd gnd cell_6t
Xbit_r207_c106 bl[106] br[106] wl[207] vdd gnd cell_6t
Xbit_r208_c106 bl[106] br[106] wl[208] vdd gnd cell_6t
Xbit_r209_c106 bl[106] br[106] wl[209] vdd gnd cell_6t
Xbit_r210_c106 bl[106] br[106] wl[210] vdd gnd cell_6t
Xbit_r211_c106 bl[106] br[106] wl[211] vdd gnd cell_6t
Xbit_r212_c106 bl[106] br[106] wl[212] vdd gnd cell_6t
Xbit_r213_c106 bl[106] br[106] wl[213] vdd gnd cell_6t
Xbit_r214_c106 bl[106] br[106] wl[214] vdd gnd cell_6t
Xbit_r215_c106 bl[106] br[106] wl[215] vdd gnd cell_6t
Xbit_r216_c106 bl[106] br[106] wl[216] vdd gnd cell_6t
Xbit_r217_c106 bl[106] br[106] wl[217] vdd gnd cell_6t
Xbit_r218_c106 bl[106] br[106] wl[218] vdd gnd cell_6t
Xbit_r219_c106 bl[106] br[106] wl[219] vdd gnd cell_6t
Xbit_r220_c106 bl[106] br[106] wl[220] vdd gnd cell_6t
Xbit_r221_c106 bl[106] br[106] wl[221] vdd gnd cell_6t
Xbit_r222_c106 bl[106] br[106] wl[222] vdd gnd cell_6t
Xbit_r223_c106 bl[106] br[106] wl[223] vdd gnd cell_6t
Xbit_r224_c106 bl[106] br[106] wl[224] vdd gnd cell_6t
Xbit_r225_c106 bl[106] br[106] wl[225] vdd gnd cell_6t
Xbit_r226_c106 bl[106] br[106] wl[226] vdd gnd cell_6t
Xbit_r227_c106 bl[106] br[106] wl[227] vdd gnd cell_6t
Xbit_r228_c106 bl[106] br[106] wl[228] vdd gnd cell_6t
Xbit_r229_c106 bl[106] br[106] wl[229] vdd gnd cell_6t
Xbit_r230_c106 bl[106] br[106] wl[230] vdd gnd cell_6t
Xbit_r231_c106 bl[106] br[106] wl[231] vdd gnd cell_6t
Xbit_r232_c106 bl[106] br[106] wl[232] vdd gnd cell_6t
Xbit_r233_c106 bl[106] br[106] wl[233] vdd gnd cell_6t
Xbit_r234_c106 bl[106] br[106] wl[234] vdd gnd cell_6t
Xbit_r235_c106 bl[106] br[106] wl[235] vdd gnd cell_6t
Xbit_r236_c106 bl[106] br[106] wl[236] vdd gnd cell_6t
Xbit_r237_c106 bl[106] br[106] wl[237] vdd gnd cell_6t
Xbit_r238_c106 bl[106] br[106] wl[238] vdd gnd cell_6t
Xbit_r239_c106 bl[106] br[106] wl[239] vdd gnd cell_6t
Xbit_r240_c106 bl[106] br[106] wl[240] vdd gnd cell_6t
Xbit_r241_c106 bl[106] br[106] wl[241] vdd gnd cell_6t
Xbit_r242_c106 bl[106] br[106] wl[242] vdd gnd cell_6t
Xbit_r243_c106 bl[106] br[106] wl[243] vdd gnd cell_6t
Xbit_r244_c106 bl[106] br[106] wl[244] vdd gnd cell_6t
Xbit_r245_c106 bl[106] br[106] wl[245] vdd gnd cell_6t
Xbit_r246_c106 bl[106] br[106] wl[246] vdd gnd cell_6t
Xbit_r247_c106 bl[106] br[106] wl[247] vdd gnd cell_6t
Xbit_r248_c106 bl[106] br[106] wl[248] vdd gnd cell_6t
Xbit_r249_c106 bl[106] br[106] wl[249] vdd gnd cell_6t
Xbit_r250_c106 bl[106] br[106] wl[250] vdd gnd cell_6t
Xbit_r251_c106 bl[106] br[106] wl[251] vdd gnd cell_6t
Xbit_r252_c106 bl[106] br[106] wl[252] vdd gnd cell_6t
Xbit_r253_c106 bl[106] br[106] wl[253] vdd gnd cell_6t
Xbit_r254_c106 bl[106] br[106] wl[254] vdd gnd cell_6t
Xbit_r255_c106 bl[106] br[106] wl[255] vdd gnd cell_6t
Xbit_r256_c106 bl[106] br[106] wl[256] vdd gnd cell_6t
Xbit_r257_c106 bl[106] br[106] wl[257] vdd gnd cell_6t
Xbit_r258_c106 bl[106] br[106] wl[258] vdd gnd cell_6t
Xbit_r259_c106 bl[106] br[106] wl[259] vdd gnd cell_6t
Xbit_r260_c106 bl[106] br[106] wl[260] vdd gnd cell_6t
Xbit_r261_c106 bl[106] br[106] wl[261] vdd gnd cell_6t
Xbit_r262_c106 bl[106] br[106] wl[262] vdd gnd cell_6t
Xbit_r263_c106 bl[106] br[106] wl[263] vdd gnd cell_6t
Xbit_r264_c106 bl[106] br[106] wl[264] vdd gnd cell_6t
Xbit_r265_c106 bl[106] br[106] wl[265] vdd gnd cell_6t
Xbit_r266_c106 bl[106] br[106] wl[266] vdd gnd cell_6t
Xbit_r267_c106 bl[106] br[106] wl[267] vdd gnd cell_6t
Xbit_r268_c106 bl[106] br[106] wl[268] vdd gnd cell_6t
Xbit_r269_c106 bl[106] br[106] wl[269] vdd gnd cell_6t
Xbit_r270_c106 bl[106] br[106] wl[270] vdd gnd cell_6t
Xbit_r271_c106 bl[106] br[106] wl[271] vdd gnd cell_6t
Xbit_r272_c106 bl[106] br[106] wl[272] vdd gnd cell_6t
Xbit_r273_c106 bl[106] br[106] wl[273] vdd gnd cell_6t
Xbit_r274_c106 bl[106] br[106] wl[274] vdd gnd cell_6t
Xbit_r275_c106 bl[106] br[106] wl[275] vdd gnd cell_6t
Xbit_r276_c106 bl[106] br[106] wl[276] vdd gnd cell_6t
Xbit_r277_c106 bl[106] br[106] wl[277] vdd gnd cell_6t
Xbit_r278_c106 bl[106] br[106] wl[278] vdd gnd cell_6t
Xbit_r279_c106 bl[106] br[106] wl[279] vdd gnd cell_6t
Xbit_r280_c106 bl[106] br[106] wl[280] vdd gnd cell_6t
Xbit_r281_c106 bl[106] br[106] wl[281] vdd gnd cell_6t
Xbit_r282_c106 bl[106] br[106] wl[282] vdd gnd cell_6t
Xbit_r283_c106 bl[106] br[106] wl[283] vdd gnd cell_6t
Xbit_r284_c106 bl[106] br[106] wl[284] vdd gnd cell_6t
Xbit_r285_c106 bl[106] br[106] wl[285] vdd gnd cell_6t
Xbit_r286_c106 bl[106] br[106] wl[286] vdd gnd cell_6t
Xbit_r287_c106 bl[106] br[106] wl[287] vdd gnd cell_6t
Xbit_r288_c106 bl[106] br[106] wl[288] vdd gnd cell_6t
Xbit_r289_c106 bl[106] br[106] wl[289] vdd gnd cell_6t
Xbit_r290_c106 bl[106] br[106] wl[290] vdd gnd cell_6t
Xbit_r291_c106 bl[106] br[106] wl[291] vdd gnd cell_6t
Xbit_r292_c106 bl[106] br[106] wl[292] vdd gnd cell_6t
Xbit_r293_c106 bl[106] br[106] wl[293] vdd gnd cell_6t
Xbit_r294_c106 bl[106] br[106] wl[294] vdd gnd cell_6t
Xbit_r295_c106 bl[106] br[106] wl[295] vdd gnd cell_6t
Xbit_r296_c106 bl[106] br[106] wl[296] vdd gnd cell_6t
Xbit_r297_c106 bl[106] br[106] wl[297] vdd gnd cell_6t
Xbit_r298_c106 bl[106] br[106] wl[298] vdd gnd cell_6t
Xbit_r299_c106 bl[106] br[106] wl[299] vdd gnd cell_6t
Xbit_r300_c106 bl[106] br[106] wl[300] vdd gnd cell_6t
Xbit_r301_c106 bl[106] br[106] wl[301] vdd gnd cell_6t
Xbit_r302_c106 bl[106] br[106] wl[302] vdd gnd cell_6t
Xbit_r303_c106 bl[106] br[106] wl[303] vdd gnd cell_6t
Xbit_r304_c106 bl[106] br[106] wl[304] vdd gnd cell_6t
Xbit_r305_c106 bl[106] br[106] wl[305] vdd gnd cell_6t
Xbit_r306_c106 bl[106] br[106] wl[306] vdd gnd cell_6t
Xbit_r307_c106 bl[106] br[106] wl[307] vdd gnd cell_6t
Xbit_r308_c106 bl[106] br[106] wl[308] vdd gnd cell_6t
Xbit_r309_c106 bl[106] br[106] wl[309] vdd gnd cell_6t
Xbit_r310_c106 bl[106] br[106] wl[310] vdd gnd cell_6t
Xbit_r311_c106 bl[106] br[106] wl[311] vdd gnd cell_6t
Xbit_r312_c106 bl[106] br[106] wl[312] vdd gnd cell_6t
Xbit_r313_c106 bl[106] br[106] wl[313] vdd gnd cell_6t
Xbit_r314_c106 bl[106] br[106] wl[314] vdd gnd cell_6t
Xbit_r315_c106 bl[106] br[106] wl[315] vdd gnd cell_6t
Xbit_r316_c106 bl[106] br[106] wl[316] vdd gnd cell_6t
Xbit_r317_c106 bl[106] br[106] wl[317] vdd gnd cell_6t
Xbit_r318_c106 bl[106] br[106] wl[318] vdd gnd cell_6t
Xbit_r319_c106 bl[106] br[106] wl[319] vdd gnd cell_6t
Xbit_r320_c106 bl[106] br[106] wl[320] vdd gnd cell_6t
Xbit_r321_c106 bl[106] br[106] wl[321] vdd gnd cell_6t
Xbit_r322_c106 bl[106] br[106] wl[322] vdd gnd cell_6t
Xbit_r323_c106 bl[106] br[106] wl[323] vdd gnd cell_6t
Xbit_r324_c106 bl[106] br[106] wl[324] vdd gnd cell_6t
Xbit_r325_c106 bl[106] br[106] wl[325] vdd gnd cell_6t
Xbit_r326_c106 bl[106] br[106] wl[326] vdd gnd cell_6t
Xbit_r327_c106 bl[106] br[106] wl[327] vdd gnd cell_6t
Xbit_r328_c106 bl[106] br[106] wl[328] vdd gnd cell_6t
Xbit_r329_c106 bl[106] br[106] wl[329] vdd gnd cell_6t
Xbit_r330_c106 bl[106] br[106] wl[330] vdd gnd cell_6t
Xbit_r331_c106 bl[106] br[106] wl[331] vdd gnd cell_6t
Xbit_r332_c106 bl[106] br[106] wl[332] vdd gnd cell_6t
Xbit_r333_c106 bl[106] br[106] wl[333] vdd gnd cell_6t
Xbit_r334_c106 bl[106] br[106] wl[334] vdd gnd cell_6t
Xbit_r335_c106 bl[106] br[106] wl[335] vdd gnd cell_6t
Xbit_r336_c106 bl[106] br[106] wl[336] vdd gnd cell_6t
Xbit_r337_c106 bl[106] br[106] wl[337] vdd gnd cell_6t
Xbit_r338_c106 bl[106] br[106] wl[338] vdd gnd cell_6t
Xbit_r339_c106 bl[106] br[106] wl[339] vdd gnd cell_6t
Xbit_r340_c106 bl[106] br[106] wl[340] vdd gnd cell_6t
Xbit_r341_c106 bl[106] br[106] wl[341] vdd gnd cell_6t
Xbit_r342_c106 bl[106] br[106] wl[342] vdd gnd cell_6t
Xbit_r343_c106 bl[106] br[106] wl[343] vdd gnd cell_6t
Xbit_r344_c106 bl[106] br[106] wl[344] vdd gnd cell_6t
Xbit_r345_c106 bl[106] br[106] wl[345] vdd gnd cell_6t
Xbit_r346_c106 bl[106] br[106] wl[346] vdd gnd cell_6t
Xbit_r347_c106 bl[106] br[106] wl[347] vdd gnd cell_6t
Xbit_r348_c106 bl[106] br[106] wl[348] vdd gnd cell_6t
Xbit_r349_c106 bl[106] br[106] wl[349] vdd gnd cell_6t
Xbit_r350_c106 bl[106] br[106] wl[350] vdd gnd cell_6t
Xbit_r351_c106 bl[106] br[106] wl[351] vdd gnd cell_6t
Xbit_r352_c106 bl[106] br[106] wl[352] vdd gnd cell_6t
Xbit_r353_c106 bl[106] br[106] wl[353] vdd gnd cell_6t
Xbit_r354_c106 bl[106] br[106] wl[354] vdd gnd cell_6t
Xbit_r355_c106 bl[106] br[106] wl[355] vdd gnd cell_6t
Xbit_r356_c106 bl[106] br[106] wl[356] vdd gnd cell_6t
Xbit_r357_c106 bl[106] br[106] wl[357] vdd gnd cell_6t
Xbit_r358_c106 bl[106] br[106] wl[358] vdd gnd cell_6t
Xbit_r359_c106 bl[106] br[106] wl[359] vdd gnd cell_6t
Xbit_r360_c106 bl[106] br[106] wl[360] vdd gnd cell_6t
Xbit_r361_c106 bl[106] br[106] wl[361] vdd gnd cell_6t
Xbit_r362_c106 bl[106] br[106] wl[362] vdd gnd cell_6t
Xbit_r363_c106 bl[106] br[106] wl[363] vdd gnd cell_6t
Xbit_r364_c106 bl[106] br[106] wl[364] vdd gnd cell_6t
Xbit_r365_c106 bl[106] br[106] wl[365] vdd gnd cell_6t
Xbit_r366_c106 bl[106] br[106] wl[366] vdd gnd cell_6t
Xbit_r367_c106 bl[106] br[106] wl[367] vdd gnd cell_6t
Xbit_r368_c106 bl[106] br[106] wl[368] vdd gnd cell_6t
Xbit_r369_c106 bl[106] br[106] wl[369] vdd gnd cell_6t
Xbit_r370_c106 bl[106] br[106] wl[370] vdd gnd cell_6t
Xbit_r371_c106 bl[106] br[106] wl[371] vdd gnd cell_6t
Xbit_r372_c106 bl[106] br[106] wl[372] vdd gnd cell_6t
Xbit_r373_c106 bl[106] br[106] wl[373] vdd gnd cell_6t
Xbit_r374_c106 bl[106] br[106] wl[374] vdd gnd cell_6t
Xbit_r375_c106 bl[106] br[106] wl[375] vdd gnd cell_6t
Xbit_r376_c106 bl[106] br[106] wl[376] vdd gnd cell_6t
Xbit_r377_c106 bl[106] br[106] wl[377] vdd gnd cell_6t
Xbit_r378_c106 bl[106] br[106] wl[378] vdd gnd cell_6t
Xbit_r379_c106 bl[106] br[106] wl[379] vdd gnd cell_6t
Xbit_r380_c106 bl[106] br[106] wl[380] vdd gnd cell_6t
Xbit_r381_c106 bl[106] br[106] wl[381] vdd gnd cell_6t
Xbit_r382_c106 bl[106] br[106] wl[382] vdd gnd cell_6t
Xbit_r383_c106 bl[106] br[106] wl[383] vdd gnd cell_6t
Xbit_r384_c106 bl[106] br[106] wl[384] vdd gnd cell_6t
Xbit_r385_c106 bl[106] br[106] wl[385] vdd gnd cell_6t
Xbit_r386_c106 bl[106] br[106] wl[386] vdd gnd cell_6t
Xbit_r387_c106 bl[106] br[106] wl[387] vdd gnd cell_6t
Xbit_r388_c106 bl[106] br[106] wl[388] vdd gnd cell_6t
Xbit_r389_c106 bl[106] br[106] wl[389] vdd gnd cell_6t
Xbit_r390_c106 bl[106] br[106] wl[390] vdd gnd cell_6t
Xbit_r391_c106 bl[106] br[106] wl[391] vdd gnd cell_6t
Xbit_r392_c106 bl[106] br[106] wl[392] vdd gnd cell_6t
Xbit_r393_c106 bl[106] br[106] wl[393] vdd gnd cell_6t
Xbit_r394_c106 bl[106] br[106] wl[394] vdd gnd cell_6t
Xbit_r395_c106 bl[106] br[106] wl[395] vdd gnd cell_6t
Xbit_r396_c106 bl[106] br[106] wl[396] vdd gnd cell_6t
Xbit_r397_c106 bl[106] br[106] wl[397] vdd gnd cell_6t
Xbit_r398_c106 bl[106] br[106] wl[398] vdd gnd cell_6t
Xbit_r399_c106 bl[106] br[106] wl[399] vdd gnd cell_6t
Xbit_r400_c106 bl[106] br[106] wl[400] vdd gnd cell_6t
Xbit_r401_c106 bl[106] br[106] wl[401] vdd gnd cell_6t
Xbit_r402_c106 bl[106] br[106] wl[402] vdd gnd cell_6t
Xbit_r403_c106 bl[106] br[106] wl[403] vdd gnd cell_6t
Xbit_r404_c106 bl[106] br[106] wl[404] vdd gnd cell_6t
Xbit_r405_c106 bl[106] br[106] wl[405] vdd gnd cell_6t
Xbit_r406_c106 bl[106] br[106] wl[406] vdd gnd cell_6t
Xbit_r407_c106 bl[106] br[106] wl[407] vdd gnd cell_6t
Xbit_r408_c106 bl[106] br[106] wl[408] vdd gnd cell_6t
Xbit_r409_c106 bl[106] br[106] wl[409] vdd gnd cell_6t
Xbit_r410_c106 bl[106] br[106] wl[410] vdd gnd cell_6t
Xbit_r411_c106 bl[106] br[106] wl[411] vdd gnd cell_6t
Xbit_r412_c106 bl[106] br[106] wl[412] vdd gnd cell_6t
Xbit_r413_c106 bl[106] br[106] wl[413] vdd gnd cell_6t
Xbit_r414_c106 bl[106] br[106] wl[414] vdd gnd cell_6t
Xbit_r415_c106 bl[106] br[106] wl[415] vdd gnd cell_6t
Xbit_r416_c106 bl[106] br[106] wl[416] vdd gnd cell_6t
Xbit_r417_c106 bl[106] br[106] wl[417] vdd gnd cell_6t
Xbit_r418_c106 bl[106] br[106] wl[418] vdd gnd cell_6t
Xbit_r419_c106 bl[106] br[106] wl[419] vdd gnd cell_6t
Xbit_r420_c106 bl[106] br[106] wl[420] vdd gnd cell_6t
Xbit_r421_c106 bl[106] br[106] wl[421] vdd gnd cell_6t
Xbit_r422_c106 bl[106] br[106] wl[422] vdd gnd cell_6t
Xbit_r423_c106 bl[106] br[106] wl[423] vdd gnd cell_6t
Xbit_r424_c106 bl[106] br[106] wl[424] vdd gnd cell_6t
Xbit_r425_c106 bl[106] br[106] wl[425] vdd gnd cell_6t
Xbit_r426_c106 bl[106] br[106] wl[426] vdd gnd cell_6t
Xbit_r427_c106 bl[106] br[106] wl[427] vdd gnd cell_6t
Xbit_r428_c106 bl[106] br[106] wl[428] vdd gnd cell_6t
Xbit_r429_c106 bl[106] br[106] wl[429] vdd gnd cell_6t
Xbit_r430_c106 bl[106] br[106] wl[430] vdd gnd cell_6t
Xbit_r431_c106 bl[106] br[106] wl[431] vdd gnd cell_6t
Xbit_r432_c106 bl[106] br[106] wl[432] vdd gnd cell_6t
Xbit_r433_c106 bl[106] br[106] wl[433] vdd gnd cell_6t
Xbit_r434_c106 bl[106] br[106] wl[434] vdd gnd cell_6t
Xbit_r435_c106 bl[106] br[106] wl[435] vdd gnd cell_6t
Xbit_r436_c106 bl[106] br[106] wl[436] vdd gnd cell_6t
Xbit_r437_c106 bl[106] br[106] wl[437] vdd gnd cell_6t
Xbit_r438_c106 bl[106] br[106] wl[438] vdd gnd cell_6t
Xbit_r439_c106 bl[106] br[106] wl[439] vdd gnd cell_6t
Xbit_r440_c106 bl[106] br[106] wl[440] vdd gnd cell_6t
Xbit_r441_c106 bl[106] br[106] wl[441] vdd gnd cell_6t
Xbit_r442_c106 bl[106] br[106] wl[442] vdd gnd cell_6t
Xbit_r443_c106 bl[106] br[106] wl[443] vdd gnd cell_6t
Xbit_r444_c106 bl[106] br[106] wl[444] vdd gnd cell_6t
Xbit_r445_c106 bl[106] br[106] wl[445] vdd gnd cell_6t
Xbit_r446_c106 bl[106] br[106] wl[446] vdd gnd cell_6t
Xbit_r447_c106 bl[106] br[106] wl[447] vdd gnd cell_6t
Xbit_r448_c106 bl[106] br[106] wl[448] vdd gnd cell_6t
Xbit_r449_c106 bl[106] br[106] wl[449] vdd gnd cell_6t
Xbit_r450_c106 bl[106] br[106] wl[450] vdd gnd cell_6t
Xbit_r451_c106 bl[106] br[106] wl[451] vdd gnd cell_6t
Xbit_r452_c106 bl[106] br[106] wl[452] vdd gnd cell_6t
Xbit_r453_c106 bl[106] br[106] wl[453] vdd gnd cell_6t
Xbit_r454_c106 bl[106] br[106] wl[454] vdd gnd cell_6t
Xbit_r455_c106 bl[106] br[106] wl[455] vdd gnd cell_6t
Xbit_r456_c106 bl[106] br[106] wl[456] vdd gnd cell_6t
Xbit_r457_c106 bl[106] br[106] wl[457] vdd gnd cell_6t
Xbit_r458_c106 bl[106] br[106] wl[458] vdd gnd cell_6t
Xbit_r459_c106 bl[106] br[106] wl[459] vdd gnd cell_6t
Xbit_r460_c106 bl[106] br[106] wl[460] vdd gnd cell_6t
Xbit_r461_c106 bl[106] br[106] wl[461] vdd gnd cell_6t
Xbit_r462_c106 bl[106] br[106] wl[462] vdd gnd cell_6t
Xbit_r463_c106 bl[106] br[106] wl[463] vdd gnd cell_6t
Xbit_r464_c106 bl[106] br[106] wl[464] vdd gnd cell_6t
Xbit_r465_c106 bl[106] br[106] wl[465] vdd gnd cell_6t
Xbit_r466_c106 bl[106] br[106] wl[466] vdd gnd cell_6t
Xbit_r467_c106 bl[106] br[106] wl[467] vdd gnd cell_6t
Xbit_r468_c106 bl[106] br[106] wl[468] vdd gnd cell_6t
Xbit_r469_c106 bl[106] br[106] wl[469] vdd gnd cell_6t
Xbit_r470_c106 bl[106] br[106] wl[470] vdd gnd cell_6t
Xbit_r471_c106 bl[106] br[106] wl[471] vdd gnd cell_6t
Xbit_r472_c106 bl[106] br[106] wl[472] vdd gnd cell_6t
Xbit_r473_c106 bl[106] br[106] wl[473] vdd gnd cell_6t
Xbit_r474_c106 bl[106] br[106] wl[474] vdd gnd cell_6t
Xbit_r475_c106 bl[106] br[106] wl[475] vdd gnd cell_6t
Xbit_r476_c106 bl[106] br[106] wl[476] vdd gnd cell_6t
Xbit_r477_c106 bl[106] br[106] wl[477] vdd gnd cell_6t
Xbit_r478_c106 bl[106] br[106] wl[478] vdd gnd cell_6t
Xbit_r479_c106 bl[106] br[106] wl[479] vdd gnd cell_6t
Xbit_r480_c106 bl[106] br[106] wl[480] vdd gnd cell_6t
Xbit_r481_c106 bl[106] br[106] wl[481] vdd gnd cell_6t
Xbit_r482_c106 bl[106] br[106] wl[482] vdd gnd cell_6t
Xbit_r483_c106 bl[106] br[106] wl[483] vdd gnd cell_6t
Xbit_r484_c106 bl[106] br[106] wl[484] vdd gnd cell_6t
Xbit_r485_c106 bl[106] br[106] wl[485] vdd gnd cell_6t
Xbit_r486_c106 bl[106] br[106] wl[486] vdd gnd cell_6t
Xbit_r487_c106 bl[106] br[106] wl[487] vdd gnd cell_6t
Xbit_r488_c106 bl[106] br[106] wl[488] vdd gnd cell_6t
Xbit_r489_c106 bl[106] br[106] wl[489] vdd gnd cell_6t
Xbit_r490_c106 bl[106] br[106] wl[490] vdd gnd cell_6t
Xbit_r491_c106 bl[106] br[106] wl[491] vdd gnd cell_6t
Xbit_r492_c106 bl[106] br[106] wl[492] vdd gnd cell_6t
Xbit_r493_c106 bl[106] br[106] wl[493] vdd gnd cell_6t
Xbit_r494_c106 bl[106] br[106] wl[494] vdd gnd cell_6t
Xbit_r495_c106 bl[106] br[106] wl[495] vdd gnd cell_6t
Xbit_r496_c106 bl[106] br[106] wl[496] vdd gnd cell_6t
Xbit_r497_c106 bl[106] br[106] wl[497] vdd gnd cell_6t
Xbit_r498_c106 bl[106] br[106] wl[498] vdd gnd cell_6t
Xbit_r499_c106 bl[106] br[106] wl[499] vdd gnd cell_6t
Xbit_r500_c106 bl[106] br[106] wl[500] vdd gnd cell_6t
Xbit_r501_c106 bl[106] br[106] wl[501] vdd gnd cell_6t
Xbit_r502_c106 bl[106] br[106] wl[502] vdd gnd cell_6t
Xbit_r503_c106 bl[106] br[106] wl[503] vdd gnd cell_6t
Xbit_r504_c106 bl[106] br[106] wl[504] vdd gnd cell_6t
Xbit_r505_c106 bl[106] br[106] wl[505] vdd gnd cell_6t
Xbit_r506_c106 bl[106] br[106] wl[506] vdd gnd cell_6t
Xbit_r507_c106 bl[106] br[106] wl[507] vdd gnd cell_6t
Xbit_r508_c106 bl[106] br[106] wl[508] vdd gnd cell_6t
Xbit_r509_c106 bl[106] br[106] wl[509] vdd gnd cell_6t
Xbit_r510_c106 bl[106] br[106] wl[510] vdd gnd cell_6t
Xbit_r511_c106 bl[106] br[106] wl[511] vdd gnd cell_6t
Xbit_r0_c107 bl[107] br[107] wl[0] vdd gnd cell_6t
Xbit_r1_c107 bl[107] br[107] wl[1] vdd gnd cell_6t
Xbit_r2_c107 bl[107] br[107] wl[2] vdd gnd cell_6t
Xbit_r3_c107 bl[107] br[107] wl[3] vdd gnd cell_6t
Xbit_r4_c107 bl[107] br[107] wl[4] vdd gnd cell_6t
Xbit_r5_c107 bl[107] br[107] wl[5] vdd gnd cell_6t
Xbit_r6_c107 bl[107] br[107] wl[6] vdd gnd cell_6t
Xbit_r7_c107 bl[107] br[107] wl[7] vdd gnd cell_6t
Xbit_r8_c107 bl[107] br[107] wl[8] vdd gnd cell_6t
Xbit_r9_c107 bl[107] br[107] wl[9] vdd gnd cell_6t
Xbit_r10_c107 bl[107] br[107] wl[10] vdd gnd cell_6t
Xbit_r11_c107 bl[107] br[107] wl[11] vdd gnd cell_6t
Xbit_r12_c107 bl[107] br[107] wl[12] vdd gnd cell_6t
Xbit_r13_c107 bl[107] br[107] wl[13] vdd gnd cell_6t
Xbit_r14_c107 bl[107] br[107] wl[14] vdd gnd cell_6t
Xbit_r15_c107 bl[107] br[107] wl[15] vdd gnd cell_6t
Xbit_r16_c107 bl[107] br[107] wl[16] vdd gnd cell_6t
Xbit_r17_c107 bl[107] br[107] wl[17] vdd gnd cell_6t
Xbit_r18_c107 bl[107] br[107] wl[18] vdd gnd cell_6t
Xbit_r19_c107 bl[107] br[107] wl[19] vdd gnd cell_6t
Xbit_r20_c107 bl[107] br[107] wl[20] vdd gnd cell_6t
Xbit_r21_c107 bl[107] br[107] wl[21] vdd gnd cell_6t
Xbit_r22_c107 bl[107] br[107] wl[22] vdd gnd cell_6t
Xbit_r23_c107 bl[107] br[107] wl[23] vdd gnd cell_6t
Xbit_r24_c107 bl[107] br[107] wl[24] vdd gnd cell_6t
Xbit_r25_c107 bl[107] br[107] wl[25] vdd gnd cell_6t
Xbit_r26_c107 bl[107] br[107] wl[26] vdd gnd cell_6t
Xbit_r27_c107 bl[107] br[107] wl[27] vdd gnd cell_6t
Xbit_r28_c107 bl[107] br[107] wl[28] vdd gnd cell_6t
Xbit_r29_c107 bl[107] br[107] wl[29] vdd gnd cell_6t
Xbit_r30_c107 bl[107] br[107] wl[30] vdd gnd cell_6t
Xbit_r31_c107 bl[107] br[107] wl[31] vdd gnd cell_6t
Xbit_r32_c107 bl[107] br[107] wl[32] vdd gnd cell_6t
Xbit_r33_c107 bl[107] br[107] wl[33] vdd gnd cell_6t
Xbit_r34_c107 bl[107] br[107] wl[34] vdd gnd cell_6t
Xbit_r35_c107 bl[107] br[107] wl[35] vdd gnd cell_6t
Xbit_r36_c107 bl[107] br[107] wl[36] vdd gnd cell_6t
Xbit_r37_c107 bl[107] br[107] wl[37] vdd gnd cell_6t
Xbit_r38_c107 bl[107] br[107] wl[38] vdd gnd cell_6t
Xbit_r39_c107 bl[107] br[107] wl[39] vdd gnd cell_6t
Xbit_r40_c107 bl[107] br[107] wl[40] vdd gnd cell_6t
Xbit_r41_c107 bl[107] br[107] wl[41] vdd gnd cell_6t
Xbit_r42_c107 bl[107] br[107] wl[42] vdd gnd cell_6t
Xbit_r43_c107 bl[107] br[107] wl[43] vdd gnd cell_6t
Xbit_r44_c107 bl[107] br[107] wl[44] vdd gnd cell_6t
Xbit_r45_c107 bl[107] br[107] wl[45] vdd gnd cell_6t
Xbit_r46_c107 bl[107] br[107] wl[46] vdd gnd cell_6t
Xbit_r47_c107 bl[107] br[107] wl[47] vdd gnd cell_6t
Xbit_r48_c107 bl[107] br[107] wl[48] vdd gnd cell_6t
Xbit_r49_c107 bl[107] br[107] wl[49] vdd gnd cell_6t
Xbit_r50_c107 bl[107] br[107] wl[50] vdd gnd cell_6t
Xbit_r51_c107 bl[107] br[107] wl[51] vdd gnd cell_6t
Xbit_r52_c107 bl[107] br[107] wl[52] vdd gnd cell_6t
Xbit_r53_c107 bl[107] br[107] wl[53] vdd gnd cell_6t
Xbit_r54_c107 bl[107] br[107] wl[54] vdd gnd cell_6t
Xbit_r55_c107 bl[107] br[107] wl[55] vdd gnd cell_6t
Xbit_r56_c107 bl[107] br[107] wl[56] vdd gnd cell_6t
Xbit_r57_c107 bl[107] br[107] wl[57] vdd gnd cell_6t
Xbit_r58_c107 bl[107] br[107] wl[58] vdd gnd cell_6t
Xbit_r59_c107 bl[107] br[107] wl[59] vdd gnd cell_6t
Xbit_r60_c107 bl[107] br[107] wl[60] vdd gnd cell_6t
Xbit_r61_c107 bl[107] br[107] wl[61] vdd gnd cell_6t
Xbit_r62_c107 bl[107] br[107] wl[62] vdd gnd cell_6t
Xbit_r63_c107 bl[107] br[107] wl[63] vdd gnd cell_6t
Xbit_r64_c107 bl[107] br[107] wl[64] vdd gnd cell_6t
Xbit_r65_c107 bl[107] br[107] wl[65] vdd gnd cell_6t
Xbit_r66_c107 bl[107] br[107] wl[66] vdd gnd cell_6t
Xbit_r67_c107 bl[107] br[107] wl[67] vdd gnd cell_6t
Xbit_r68_c107 bl[107] br[107] wl[68] vdd gnd cell_6t
Xbit_r69_c107 bl[107] br[107] wl[69] vdd gnd cell_6t
Xbit_r70_c107 bl[107] br[107] wl[70] vdd gnd cell_6t
Xbit_r71_c107 bl[107] br[107] wl[71] vdd gnd cell_6t
Xbit_r72_c107 bl[107] br[107] wl[72] vdd gnd cell_6t
Xbit_r73_c107 bl[107] br[107] wl[73] vdd gnd cell_6t
Xbit_r74_c107 bl[107] br[107] wl[74] vdd gnd cell_6t
Xbit_r75_c107 bl[107] br[107] wl[75] vdd gnd cell_6t
Xbit_r76_c107 bl[107] br[107] wl[76] vdd gnd cell_6t
Xbit_r77_c107 bl[107] br[107] wl[77] vdd gnd cell_6t
Xbit_r78_c107 bl[107] br[107] wl[78] vdd gnd cell_6t
Xbit_r79_c107 bl[107] br[107] wl[79] vdd gnd cell_6t
Xbit_r80_c107 bl[107] br[107] wl[80] vdd gnd cell_6t
Xbit_r81_c107 bl[107] br[107] wl[81] vdd gnd cell_6t
Xbit_r82_c107 bl[107] br[107] wl[82] vdd gnd cell_6t
Xbit_r83_c107 bl[107] br[107] wl[83] vdd gnd cell_6t
Xbit_r84_c107 bl[107] br[107] wl[84] vdd gnd cell_6t
Xbit_r85_c107 bl[107] br[107] wl[85] vdd gnd cell_6t
Xbit_r86_c107 bl[107] br[107] wl[86] vdd gnd cell_6t
Xbit_r87_c107 bl[107] br[107] wl[87] vdd gnd cell_6t
Xbit_r88_c107 bl[107] br[107] wl[88] vdd gnd cell_6t
Xbit_r89_c107 bl[107] br[107] wl[89] vdd gnd cell_6t
Xbit_r90_c107 bl[107] br[107] wl[90] vdd gnd cell_6t
Xbit_r91_c107 bl[107] br[107] wl[91] vdd gnd cell_6t
Xbit_r92_c107 bl[107] br[107] wl[92] vdd gnd cell_6t
Xbit_r93_c107 bl[107] br[107] wl[93] vdd gnd cell_6t
Xbit_r94_c107 bl[107] br[107] wl[94] vdd gnd cell_6t
Xbit_r95_c107 bl[107] br[107] wl[95] vdd gnd cell_6t
Xbit_r96_c107 bl[107] br[107] wl[96] vdd gnd cell_6t
Xbit_r97_c107 bl[107] br[107] wl[97] vdd gnd cell_6t
Xbit_r98_c107 bl[107] br[107] wl[98] vdd gnd cell_6t
Xbit_r99_c107 bl[107] br[107] wl[99] vdd gnd cell_6t
Xbit_r100_c107 bl[107] br[107] wl[100] vdd gnd cell_6t
Xbit_r101_c107 bl[107] br[107] wl[101] vdd gnd cell_6t
Xbit_r102_c107 bl[107] br[107] wl[102] vdd gnd cell_6t
Xbit_r103_c107 bl[107] br[107] wl[103] vdd gnd cell_6t
Xbit_r104_c107 bl[107] br[107] wl[104] vdd gnd cell_6t
Xbit_r105_c107 bl[107] br[107] wl[105] vdd gnd cell_6t
Xbit_r106_c107 bl[107] br[107] wl[106] vdd gnd cell_6t
Xbit_r107_c107 bl[107] br[107] wl[107] vdd gnd cell_6t
Xbit_r108_c107 bl[107] br[107] wl[108] vdd gnd cell_6t
Xbit_r109_c107 bl[107] br[107] wl[109] vdd gnd cell_6t
Xbit_r110_c107 bl[107] br[107] wl[110] vdd gnd cell_6t
Xbit_r111_c107 bl[107] br[107] wl[111] vdd gnd cell_6t
Xbit_r112_c107 bl[107] br[107] wl[112] vdd gnd cell_6t
Xbit_r113_c107 bl[107] br[107] wl[113] vdd gnd cell_6t
Xbit_r114_c107 bl[107] br[107] wl[114] vdd gnd cell_6t
Xbit_r115_c107 bl[107] br[107] wl[115] vdd gnd cell_6t
Xbit_r116_c107 bl[107] br[107] wl[116] vdd gnd cell_6t
Xbit_r117_c107 bl[107] br[107] wl[117] vdd gnd cell_6t
Xbit_r118_c107 bl[107] br[107] wl[118] vdd gnd cell_6t
Xbit_r119_c107 bl[107] br[107] wl[119] vdd gnd cell_6t
Xbit_r120_c107 bl[107] br[107] wl[120] vdd gnd cell_6t
Xbit_r121_c107 bl[107] br[107] wl[121] vdd gnd cell_6t
Xbit_r122_c107 bl[107] br[107] wl[122] vdd gnd cell_6t
Xbit_r123_c107 bl[107] br[107] wl[123] vdd gnd cell_6t
Xbit_r124_c107 bl[107] br[107] wl[124] vdd gnd cell_6t
Xbit_r125_c107 bl[107] br[107] wl[125] vdd gnd cell_6t
Xbit_r126_c107 bl[107] br[107] wl[126] vdd gnd cell_6t
Xbit_r127_c107 bl[107] br[107] wl[127] vdd gnd cell_6t
Xbit_r128_c107 bl[107] br[107] wl[128] vdd gnd cell_6t
Xbit_r129_c107 bl[107] br[107] wl[129] vdd gnd cell_6t
Xbit_r130_c107 bl[107] br[107] wl[130] vdd gnd cell_6t
Xbit_r131_c107 bl[107] br[107] wl[131] vdd gnd cell_6t
Xbit_r132_c107 bl[107] br[107] wl[132] vdd gnd cell_6t
Xbit_r133_c107 bl[107] br[107] wl[133] vdd gnd cell_6t
Xbit_r134_c107 bl[107] br[107] wl[134] vdd gnd cell_6t
Xbit_r135_c107 bl[107] br[107] wl[135] vdd gnd cell_6t
Xbit_r136_c107 bl[107] br[107] wl[136] vdd gnd cell_6t
Xbit_r137_c107 bl[107] br[107] wl[137] vdd gnd cell_6t
Xbit_r138_c107 bl[107] br[107] wl[138] vdd gnd cell_6t
Xbit_r139_c107 bl[107] br[107] wl[139] vdd gnd cell_6t
Xbit_r140_c107 bl[107] br[107] wl[140] vdd gnd cell_6t
Xbit_r141_c107 bl[107] br[107] wl[141] vdd gnd cell_6t
Xbit_r142_c107 bl[107] br[107] wl[142] vdd gnd cell_6t
Xbit_r143_c107 bl[107] br[107] wl[143] vdd gnd cell_6t
Xbit_r144_c107 bl[107] br[107] wl[144] vdd gnd cell_6t
Xbit_r145_c107 bl[107] br[107] wl[145] vdd gnd cell_6t
Xbit_r146_c107 bl[107] br[107] wl[146] vdd gnd cell_6t
Xbit_r147_c107 bl[107] br[107] wl[147] vdd gnd cell_6t
Xbit_r148_c107 bl[107] br[107] wl[148] vdd gnd cell_6t
Xbit_r149_c107 bl[107] br[107] wl[149] vdd gnd cell_6t
Xbit_r150_c107 bl[107] br[107] wl[150] vdd gnd cell_6t
Xbit_r151_c107 bl[107] br[107] wl[151] vdd gnd cell_6t
Xbit_r152_c107 bl[107] br[107] wl[152] vdd gnd cell_6t
Xbit_r153_c107 bl[107] br[107] wl[153] vdd gnd cell_6t
Xbit_r154_c107 bl[107] br[107] wl[154] vdd gnd cell_6t
Xbit_r155_c107 bl[107] br[107] wl[155] vdd gnd cell_6t
Xbit_r156_c107 bl[107] br[107] wl[156] vdd gnd cell_6t
Xbit_r157_c107 bl[107] br[107] wl[157] vdd gnd cell_6t
Xbit_r158_c107 bl[107] br[107] wl[158] vdd gnd cell_6t
Xbit_r159_c107 bl[107] br[107] wl[159] vdd gnd cell_6t
Xbit_r160_c107 bl[107] br[107] wl[160] vdd gnd cell_6t
Xbit_r161_c107 bl[107] br[107] wl[161] vdd gnd cell_6t
Xbit_r162_c107 bl[107] br[107] wl[162] vdd gnd cell_6t
Xbit_r163_c107 bl[107] br[107] wl[163] vdd gnd cell_6t
Xbit_r164_c107 bl[107] br[107] wl[164] vdd gnd cell_6t
Xbit_r165_c107 bl[107] br[107] wl[165] vdd gnd cell_6t
Xbit_r166_c107 bl[107] br[107] wl[166] vdd gnd cell_6t
Xbit_r167_c107 bl[107] br[107] wl[167] vdd gnd cell_6t
Xbit_r168_c107 bl[107] br[107] wl[168] vdd gnd cell_6t
Xbit_r169_c107 bl[107] br[107] wl[169] vdd gnd cell_6t
Xbit_r170_c107 bl[107] br[107] wl[170] vdd gnd cell_6t
Xbit_r171_c107 bl[107] br[107] wl[171] vdd gnd cell_6t
Xbit_r172_c107 bl[107] br[107] wl[172] vdd gnd cell_6t
Xbit_r173_c107 bl[107] br[107] wl[173] vdd gnd cell_6t
Xbit_r174_c107 bl[107] br[107] wl[174] vdd gnd cell_6t
Xbit_r175_c107 bl[107] br[107] wl[175] vdd gnd cell_6t
Xbit_r176_c107 bl[107] br[107] wl[176] vdd gnd cell_6t
Xbit_r177_c107 bl[107] br[107] wl[177] vdd gnd cell_6t
Xbit_r178_c107 bl[107] br[107] wl[178] vdd gnd cell_6t
Xbit_r179_c107 bl[107] br[107] wl[179] vdd gnd cell_6t
Xbit_r180_c107 bl[107] br[107] wl[180] vdd gnd cell_6t
Xbit_r181_c107 bl[107] br[107] wl[181] vdd gnd cell_6t
Xbit_r182_c107 bl[107] br[107] wl[182] vdd gnd cell_6t
Xbit_r183_c107 bl[107] br[107] wl[183] vdd gnd cell_6t
Xbit_r184_c107 bl[107] br[107] wl[184] vdd gnd cell_6t
Xbit_r185_c107 bl[107] br[107] wl[185] vdd gnd cell_6t
Xbit_r186_c107 bl[107] br[107] wl[186] vdd gnd cell_6t
Xbit_r187_c107 bl[107] br[107] wl[187] vdd gnd cell_6t
Xbit_r188_c107 bl[107] br[107] wl[188] vdd gnd cell_6t
Xbit_r189_c107 bl[107] br[107] wl[189] vdd gnd cell_6t
Xbit_r190_c107 bl[107] br[107] wl[190] vdd gnd cell_6t
Xbit_r191_c107 bl[107] br[107] wl[191] vdd gnd cell_6t
Xbit_r192_c107 bl[107] br[107] wl[192] vdd gnd cell_6t
Xbit_r193_c107 bl[107] br[107] wl[193] vdd gnd cell_6t
Xbit_r194_c107 bl[107] br[107] wl[194] vdd gnd cell_6t
Xbit_r195_c107 bl[107] br[107] wl[195] vdd gnd cell_6t
Xbit_r196_c107 bl[107] br[107] wl[196] vdd gnd cell_6t
Xbit_r197_c107 bl[107] br[107] wl[197] vdd gnd cell_6t
Xbit_r198_c107 bl[107] br[107] wl[198] vdd gnd cell_6t
Xbit_r199_c107 bl[107] br[107] wl[199] vdd gnd cell_6t
Xbit_r200_c107 bl[107] br[107] wl[200] vdd gnd cell_6t
Xbit_r201_c107 bl[107] br[107] wl[201] vdd gnd cell_6t
Xbit_r202_c107 bl[107] br[107] wl[202] vdd gnd cell_6t
Xbit_r203_c107 bl[107] br[107] wl[203] vdd gnd cell_6t
Xbit_r204_c107 bl[107] br[107] wl[204] vdd gnd cell_6t
Xbit_r205_c107 bl[107] br[107] wl[205] vdd gnd cell_6t
Xbit_r206_c107 bl[107] br[107] wl[206] vdd gnd cell_6t
Xbit_r207_c107 bl[107] br[107] wl[207] vdd gnd cell_6t
Xbit_r208_c107 bl[107] br[107] wl[208] vdd gnd cell_6t
Xbit_r209_c107 bl[107] br[107] wl[209] vdd gnd cell_6t
Xbit_r210_c107 bl[107] br[107] wl[210] vdd gnd cell_6t
Xbit_r211_c107 bl[107] br[107] wl[211] vdd gnd cell_6t
Xbit_r212_c107 bl[107] br[107] wl[212] vdd gnd cell_6t
Xbit_r213_c107 bl[107] br[107] wl[213] vdd gnd cell_6t
Xbit_r214_c107 bl[107] br[107] wl[214] vdd gnd cell_6t
Xbit_r215_c107 bl[107] br[107] wl[215] vdd gnd cell_6t
Xbit_r216_c107 bl[107] br[107] wl[216] vdd gnd cell_6t
Xbit_r217_c107 bl[107] br[107] wl[217] vdd gnd cell_6t
Xbit_r218_c107 bl[107] br[107] wl[218] vdd gnd cell_6t
Xbit_r219_c107 bl[107] br[107] wl[219] vdd gnd cell_6t
Xbit_r220_c107 bl[107] br[107] wl[220] vdd gnd cell_6t
Xbit_r221_c107 bl[107] br[107] wl[221] vdd gnd cell_6t
Xbit_r222_c107 bl[107] br[107] wl[222] vdd gnd cell_6t
Xbit_r223_c107 bl[107] br[107] wl[223] vdd gnd cell_6t
Xbit_r224_c107 bl[107] br[107] wl[224] vdd gnd cell_6t
Xbit_r225_c107 bl[107] br[107] wl[225] vdd gnd cell_6t
Xbit_r226_c107 bl[107] br[107] wl[226] vdd gnd cell_6t
Xbit_r227_c107 bl[107] br[107] wl[227] vdd gnd cell_6t
Xbit_r228_c107 bl[107] br[107] wl[228] vdd gnd cell_6t
Xbit_r229_c107 bl[107] br[107] wl[229] vdd gnd cell_6t
Xbit_r230_c107 bl[107] br[107] wl[230] vdd gnd cell_6t
Xbit_r231_c107 bl[107] br[107] wl[231] vdd gnd cell_6t
Xbit_r232_c107 bl[107] br[107] wl[232] vdd gnd cell_6t
Xbit_r233_c107 bl[107] br[107] wl[233] vdd gnd cell_6t
Xbit_r234_c107 bl[107] br[107] wl[234] vdd gnd cell_6t
Xbit_r235_c107 bl[107] br[107] wl[235] vdd gnd cell_6t
Xbit_r236_c107 bl[107] br[107] wl[236] vdd gnd cell_6t
Xbit_r237_c107 bl[107] br[107] wl[237] vdd gnd cell_6t
Xbit_r238_c107 bl[107] br[107] wl[238] vdd gnd cell_6t
Xbit_r239_c107 bl[107] br[107] wl[239] vdd gnd cell_6t
Xbit_r240_c107 bl[107] br[107] wl[240] vdd gnd cell_6t
Xbit_r241_c107 bl[107] br[107] wl[241] vdd gnd cell_6t
Xbit_r242_c107 bl[107] br[107] wl[242] vdd gnd cell_6t
Xbit_r243_c107 bl[107] br[107] wl[243] vdd gnd cell_6t
Xbit_r244_c107 bl[107] br[107] wl[244] vdd gnd cell_6t
Xbit_r245_c107 bl[107] br[107] wl[245] vdd gnd cell_6t
Xbit_r246_c107 bl[107] br[107] wl[246] vdd gnd cell_6t
Xbit_r247_c107 bl[107] br[107] wl[247] vdd gnd cell_6t
Xbit_r248_c107 bl[107] br[107] wl[248] vdd gnd cell_6t
Xbit_r249_c107 bl[107] br[107] wl[249] vdd gnd cell_6t
Xbit_r250_c107 bl[107] br[107] wl[250] vdd gnd cell_6t
Xbit_r251_c107 bl[107] br[107] wl[251] vdd gnd cell_6t
Xbit_r252_c107 bl[107] br[107] wl[252] vdd gnd cell_6t
Xbit_r253_c107 bl[107] br[107] wl[253] vdd gnd cell_6t
Xbit_r254_c107 bl[107] br[107] wl[254] vdd gnd cell_6t
Xbit_r255_c107 bl[107] br[107] wl[255] vdd gnd cell_6t
Xbit_r256_c107 bl[107] br[107] wl[256] vdd gnd cell_6t
Xbit_r257_c107 bl[107] br[107] wl[257] vdd gnd cell_6t
Xbit_r258_c107 bl[107] br[107] wl[258] vdd gnd cell_6t
Xbit_r259_c107 bl[107] br[107] wl[259] vdd gnd cell_6t
Xbit_r260_c107 bl[107] br[107] wl[260] vdd gnd cell_6t
Xbit_r261_c107 bl[107] br[107] wl[261] vdd gnd cell_6t
Xbit_r262_c107 bl[107] br[107] wl[262] vdd gnd cell_6t
Xbit_r263_c107 bl[107] br[107] wl[263] vdd gnd cell_6t
Xbit_r264_c107 bl[107] br[107] wl[264] vdd gnd cell_6t
Xbit_r265_c107 bl[107] br[107] wl[265] vdd gnd cell_6t
Xbit_r266_c107 bl[107] br[107] wl[266] vdd gnd cell_6t
Xbit_r267_c107 bl[107] br[107] wl[267] vdd gnd cell_6t
Xbit_r268_c107 bl[107] br[107] wl[268] vdd gnd cell_6t
Xbit_r269_c107 bl[107] br[107] wl[269] vdd gnd cell_6t
Xbit_r270_c107 bl[107] br[107] wl[270] vdd gnd cell_6t
Xbit_r271_c107 bl[107] br[107] wl[271] vdd gnd cell_6t
Xbit_r272_c107 bl[107] br[107] wl[272] vdd gnd cell_6t
Xbit_r273_c107 bl[107] br[107] wl[273] vdd gnd cell_6t
Xbit_r274_c107 bl[107] br[107] wl[274] vdd gnd cell_6t
Xbit_r275_c107 bl[107] br[107] wl[275] vdd gnd cell_6t
Xbit_r276_c107 bl[107] br[107] wl[276] vdd gnd cell_6t
Xbit_r277_c107 bl[107] br[107] wl[277] vdd gnd cell_6t
Xbit_r278_c107 bl[107] br[107] wl[278] vdd gnd cell_6t
Xbit_r279_c107 bl[107] br[107] wl[279] vdd gnd cell_6t
Xbit_r280_c107 bl[107] br[107] wl[280] vdd gnd cell_6t
Xbit_r281_c107 bl[107] br[107] wl[281] vdd gnd cell_6t
Xbit_r282_c107 bl[107] br[107] wl[282] vdd gnd cell_6t
Xbit_r283_c107 bl[107] br[107] wl[283] vdd gnd cell_6t
Xbit_r284_c107 bl[107] br[107] wl[284] vdd gnd cell_6t
Xbit_r285_c107 bl[107] br[107] wl[285] vdd gnd cell_6t
Xbit_r286_c107 bl[107] br[107] wl[286] vdd gnd cell_6t
Xbit_r287_c107 bl[107] br[107] wl[287] vdd gnd cell_6t
Xbit_r288_c107 bl[107] br[107] wl[288] vdd gnd cell_6t
Xbit_r289_c107 bl[107] br[107] wl[289] vdd gnd cell_6t
Xbit_r290_c107 bl[107] br[107] wl[290] vdd gnd cell_6t
Xbit_r291_c107 bl[107] br[107] wl[291] vdd gnd cell_6t
Xbit_r292_c107 bl[107] br[107] wl[292] vdd gnd cell_6t
Xbit_r293_c107 bl[107] br[107] wl[293] vdd gnd cell_6t
Xbit_r294_c107 bl[107] br[107] wl[294] vdd gnd cell_6t
Xbit_r295_c107 bl[107] br[107] wl[295] vdd gnd cell_6t
Xbit_r296_c107 bl[107] br[107] wl[296] vdd gnd cell_6t
Xbit_r297_c107 bl[107] br[107] wl[297] vdd gnd cell_6t
Xbit_r298_c107 bl[107] br[107] wl[298] vdd gnd cell_6t
Xbit_r299_c107 bl[107] br[107] wl[299] vdd gnd cell_6t
Xbit_r300_c107 bl[107] br[107] wl[300] vdd gnd cell_6t
Xbit_r301_c107 bl[107] br[107] wl[301] vdd gnd cell_6t
Xbit_r302_c107 bl[107] br[107] wl[302] vdd gnd cell_6t
Xbit_r303_c107 bl[107] br[107] wl[303] vdd gnd cell_6t
Xbit_r304_c107 bl[107] br[107] wl[304] vdd gnd cell_6t
Xbit_r305_c107 bl[107] br[107] wl[305] vdd gnd cell_6t
Xbit_r306_c107 bl[107] br[107] wl[306] vdd gnd cell_6t
Xbit_r307_c107 bl[107] br[107] wl[307] vdd gnd cell_6t
Xbit_r308_c107 bl[107] br[107] wl[308] vdd gnd cell_6t
Xbit_r309_c107 bl[107] br[107] wl[309] vdd gnd cell_6t
Xbit_r310_c107 bl[107] br[107] wl[310] vdd gnd cell_6t
Xbit_r311_c107 bl[107] br[107] wl[311] vdd gnd cell_6t
Xbit_r312_c107 bl[107] br[107] wl[312] vdd gnd cell_6t
Xbit_r313_c107 bl[107] br[107] wl[313] vdd gnd cell_6t
Xbit_r314_c107 bl[107] br[107] wl[314] vdd gnd cell_6t
Xbit_r315_c107 bl[107] br[107] wl[315] vdd gnd cell_6t
Xbit_r316_c107 bl[107] br[107] wl[316] vdd gnd cell_6t
Xbit_r317_c107 bl[107] br[107] wl[317] vdd gnd cell_6t
Xbit_r318_c107 bl[107] br[107] wl[318] vdd gnd cell_6t
Xbit_r319_c107 bl[107] br[107] wl[319] vdd gnd cell_6t
Xbit_r320_c107 bl[107] br[107] wl[320] vdd gnd cell_6t
Xbit_r321_c107 bl[107] br[107] wl[321] vdd gnd cell_6t
Xbit_r322_c107 bl[107] br[107] wl[322] vdd gnd cell_6t
Xbit_r323_c107 bl[107] br[107] wl[323] vdd gnd cell_6t
Xbit_r324_c107 bl[107] br[107] wl[324] vdd gnd cell_6t
Xbit_r325_c107 bl[107] br[107] wl[325] vdd gnd cell_6t
Xbit_r326_c107 bl[107] br[107] wl[326] vdd gnd cell_6t
Xbit_r327_c107 bl[107] br[107] wl[327] vdd gnd cell_6t
Xbit_r328_c107 bl[107] br[107] wl[328] vdd gnd cell_6t
Xbit_r329_c107 bl[107] br[107] wl[329] vdd gnd cell_6t
Xbit_r330_c107 bl[107] br[107] wl[330] vdd gnd cell_6t
Xbit_r331_c107 bl[107] br[107] wl[331] vdd gnd cell_6t
Xbit_r332_c107 bl[107] br[107] wl[332] vdd gnd cell_6t
Xbit_r333_c107 bl[107] br[107] wl[333] vdd gnd cell_6t
Xbit_r334_c107 bl[107] br[107] wl[334] vdd gnd cell_6t
Xbit_r335_c107 bl[107] br[107] wl[335] vdd gnd cell_6t
Xbit_r336_c107 bl[107] br[107] wl[336] vdd gnd cell_6t
Xbit_r337_c107 bl[107] br[107] wl[337] vdd gnd cell_6t
Xbit_r338_c107 bl[107] br[107] wl[338] vdd gnd cell_6t
Xbit_r339_c107 bl[107] br[107] wl[339] vdd gnd cell_6t
Xbit_r340_c107 bl[107] br[107] wl[340] vdd gnd cell_6t
Xbit_r341_c107 bl[107] br[107] wl[341] vdd gnd cell_6t
Xbit_r342_c107 bl[107] br[107] wl[342] vdd gnd cell_6t
Xbit_r343_c107 bl[107] br[107] wl[343] vdd gnd cell_6t
Xbit_r344_c107 bl[107] br[107] wl[344] vdd gnd cell_6t
Xbit_r345_c107 bl[107] br[107] wl[345] vdd gnd cell_6t
Xbit_r346_c107 bl[107] br[107] wl[346] vdd gnd cell_6t
Xbit_r347_c107 bl[107] br[107] wl[347] vdd gnd cell_6t
Xbit_r348_c107 bl[107] br[107] wl[348] vdd gnd cell_6t
Xbit_r349_c107 bl[107] br[107] wl[349] vdd gnd cell_6t
Xbit_r350_c107 bl[107] br[107] wl[350] vdd gnd cell_6t
Xbit_r351_c107 bl[107] br[107] wl[351] vdd gnd cell_6t
Xbit_r352_c107 bl[107] br[107] wl[352] vdd gnd cell_6t
Xbit_r353_c107 bl[107] br[107] wl[353] vdd gnd cell_6t
Xbit_r354_c107 bl[107] br[107] wl[354] vdd gnd cell_6t
Xbit_r355_c107 bl[107] br[107] wl[355] vdd gnd cell_6t
Xbit_r356_c107 bl[107] br[107] wl[356] vdd gnd cell_6t
Xbit_r357_c107 bl[107] br[107] wl[357] vdd gnd cell_6t
Xbit_r358_c107 bl[107] br[107] wl[358] vdd gnd cell_6t
Xbit_r359_c107 bl[107] br[107] wl[359] vdd gnd cell_6t
Xbit_r360_c107 bl[107] br[107] wl[360] vdd gnd cell_6t
Xbit_r361_c107 bl[107] br[107] wl[361] vdd gnd cell_6t
Xbit_r362_c107 bl[107] br[107] wl[362] vdd gnd cell_6t
Xbit_r363_c107 bl[107] br[107] wl[363] vdd gnd cell_6t
Xbit_r364_c107 bl[107] br[107] wl[364] vdd gnd cell_6t
Xbit_r365_c107 bl[107] br[107] wl[365] vdd gnd cell_6t
Xbit_r366_c107 bl[107] br[107] wl[366] vdd gnd cell_6t
Xbit_r367_c107 bl[107] br[107] wl[367] vdd gnd cell_6t
Xbit_r368_c107 bl[107] br[107] wl[368] vdd gnd cell_6t
Xbit_r369_c107 bl[107] br[107] wl[369] vdd gnd cell_6t
Xbit_r370_c107 bl[107] br[107] wl[370] vdd gnd cell_6t
Xbit_r371_c107 bl[107] br[107] wl[371] vdd gnd cell_6t
Xbit_r372_c107 bl[107] br[107] wl[372] vdd gnd cell_6t
Xbit_r373_c107 bl[107] br[107] wl[373] vdd gnd cell_6t
Xbit_r374_c107 bl[107] br[107] wl[374] vdd gnd cell_6t
Xbit_r375_c107 bl[107] br[107] wl[375] vdd gnd cell_6t
Xbit_r376_c107 bl[107] br[107] wl[376] vdd gnd cell_6t
Xbit_r377_c107 bl[107] br[107] wl[377] vdd gnd cell_6t
Xbit_r378_c107 bl[107] br[107] wl[378] vdd gnd cell_6t
Xbit_r379_c107 bl[107] br[107] wl[379] vdd gnd cell_6t
Xbit_r380_c107 bl[107] br[107] wl[380] vdd gnd cell_6t
Xbit_r381_c107 bl[107] br[107] wl[381] vdd gnd cell_6t
Xbit_r382_c107 bl[107] br[107] wl[382] vdd gnd cell_6t
Xbit_r383_c107 bl[107] br[107] wl[383] vdd gnd cell_6t
Xbit_r384_c107 bl[107] br[107] wl[384] vdd gnd cell_6t
Xbit_r385_c107 bl[107] br[107] wl[385] vdd gnd cell_6t
Xbit_r386_c107 bl[107] br[107] wl[386] vdd gnd cell_6t
Xbit_r387_c107 bl[107] br[107] wl[387] vdd gnd cell_6t
Xbit_r388_c107 bl[107] br[107] wl[388] vdd gnd cell_6t
Xbit_r389_c107 bl[107] br[107] wl[389] vdd gnd cell_6t
Xbit_r390_c107 bl[107] br[107] wl[390] vdd gnd cell_6t
Xbit_r391_c107 bl[107] br[107] wl[391] vdd gnd cell_6t
Xbit_r392_c107 bl[107] br[107] wl[392] vdd gnd cell_6t
Xbit_r393_c107 bl[107] br[107] wl[393] vdd gnd cell_6t
Xbit_r394_c107 bl[107] br[107] wl[394] vdd gnd cell_6t
Xbit_r395_c107 bl[107] br[107] wl[395] vdd gnd cell_6t
Xbit_r396_c107 bl[107] br[107] wl[396] vdd gnd cell_6t
Xbit_r397_c107 bl[107] br[107] wl[397] vdd gnd cell_6t
Xbit_r398_c107 bl[107] br[107] wl[398] vdd gnd cell_6t
Xbit_r399_c107 bl[107] br[107] wl[399] vdd gnd cell_6t
Xbit_r400_c107 bl[107] br[107] wl[400] vdd gnd cell_6t
Xbit_r401_c107 bl[107] br[107] wl[401] vdd gnd cell_6t
Xbit_r402_c107 bl[107] br[107] wl[402] vdd gnd cell_6t
Xbit_r403_c107 bl[107] br[107] wl[403] vdd gnd cell_6t
Xbit_r404_c107 bl[107] br[107] wl[404] vdd gnd cell_6t
Xbit_r405_c107 bl[107] br[107] wl[405] vdd gnd cell_6t
Xbit_r406_c107 bl[107] br[107] wl[406] vdd gnd cell_6t
Xbit_r407_c107 bl[107] br[107] wl[407] vdd gnd cell_6t
Xbit_r408_c107 bl[107] br[107] wl[408] vdd gnd cell_6t
Xbit_r409_c107 bl[107] br[107] wl[409] vdd gnd cell_6t
Xbit_r410_c107 bl[107] br[107] wl[410] vdd gnd cell_6t
Xbit_r411_c107 bl[107] br[107] wl[411] vdd gnd cell_6t
Xbit_r412_c107 bl[107] br[107] wl[412] vdd gnd cell_6t
Xbit_r413_c107 bl[107] br[107] wl[413] vdd gnd cell_6t
Xbit_r414_c107 bl[107] br[107] wl[414] vdd gnd cell_6t
Xbit_r415_c107 bl[107] br[107] wl[415] vdd gnd cell_6t
Xbit_r416_c107 bl[107] br[107] wl[416] vdd gnd cell_6t
Xbit_r417_c107 bl[107] br[107] wl[417] vdd gnd cell_6t
Xbit_r418_c107 bl[107] br[107] wl[418] vdd gnd cell_6t
Xbit_r419_c107 bl[107] br[107] wl[419] vdd gnd cell_6t
Xbit_r420_c107 bl[107] br[107] wl[420] vdd gnd cell_6t
Xbit_r421_c107 bl[107] br[107] wl[421] vdd gnd cell_6t
Xbit_r422_c107 bl[107] br[107] wl[422] vdd gnd cell_6t
Xbit_r423_c107 bl[107] br[107] wl[423] vdd gnd cell_6t
Xbit_r424_c107 bl[107] br[107] wl[424] vdd gnd cell_6t
Xbit_r425_c107 bl[107] br[107] wl[425] vdd gnd cell_6t
Xbit_r426_c107 bl[107] br[107] wl[426] vdd gnd cell_6t
Xbit_r427_c107 bl[107] br[107] wl[427] vdd gnd cell_6t
Xbit_r428_c107 bl[107] br[107] wl[428] vdd gnd cell_6t
Xbit_r429_c107 bl[107] br[107] wl[429] vdd gnd cell_6t
Xbit_r430_c107 bl[107] br[107] wl[430] vdd gnd cell_6t
Xbit_r431_c107 bl[107] br[107] wl[431] vdd gnd cell_6t
Xbit_r432_c107 bl[107] br[107] wl[432] vdd gnd cell_6t
Xbit_r433_c107 bl[107] br[107] wl[433] vdd gnd cell_6t
Xbit_r434_c107 bl[107] br[107] wl[434] vdd gnd cell_6t
Xbit_r435_c107 bl[107] br[107] wl[435] vdd gnd cell_6t
Xbit_r436_c107 bl[107] br[107] wl[436] vdd gnd cell_6t
Xbit_r437_c107 bl[107] br[107] wl[437] vdd gnd cell_6t
Xbit_r438_c107 bl[107] br[107] wl[438] vdd gnd cell_6t
Xbit_r439_c107 bl[107] br[107] wl[439] vdd gnd cell_6t
Xbit_r440_c107 bl[107] br[107] wl[440] vdd gnd cell_6t
Xbit_r441_c107 bl[107] br[107] wl[441] vdd gnd cell_6t
Xbit_r442_c107 bl[107] br[107] wl[442] vdd gnd cell_6t
Xbit_r443_c107 bl[107] br[107] wl[443] vdd gnd cell_6t
Xbit_r444_c107 bl[107] br[107] wl[444] vdd gnd cell_6t
Xbit_r445_c107 bl[107] br[107] wl[445] vdd gnd cell_6t
Xbit_r446_c107 bl[107] br[107] wl[446] vdd gnd cell_6t
Xbit_r447_c107 bl[107] br[107] wl[447] vdd gnd cell_6t
Xbit_r448_c107 bl[107] br[107] wl[448] vdd gnd cell_6t
Xbit_r449_c107 bl[107] br[107] wl[449] vdd gnd cell_6t
Xbit_r450_c107 bl[107] br[107] wl[450] vdd gnd cell_6t
Xbit_r451_c107 bl[107] br[107] wl[451] vdd gnd cell_6t
Xbit_r452_c107 bl[107] br[107] wl[452] vdd gnd cell_6t
Xbit_r453_c107 bl[107] br[107] wl[453] vdd gnd cell_6t
Xbit_r454_c107 bl[107] br[107] wl[454] vdd gnd cell_6t
Xbit_r455_c107 bl[107] br[107] wl[455] vdd gnd cell_6t
Xbit_r456_c107 bl[107] br[107] wl[456] vdd gnd cell_6t
Xbit_r457_c107 bl[107] br[107] wl[457] vdd gnd cell_6t
Xbit_r458_c107 bl[107] br[107] wl[458] vdd gnd cell_6t
Xbit_r459_c107 bl[107] br[107] wl[459] vdd gnd cell_6t
Xbit_r460_c107 bl[107] br[107] wl[460] vdd gnd cell_6t
Xbit_r461_c107 bl[107] br[107] wl[461] vdd gnd cell_6t
Xbit_r462_c107 bl[107] br[107] wl[462] vdd gnd cell_6t
Xbit_r463_c107 bl[107] br[107] wl[463] vdd gnd cell_6t
Xbit_r464_c107 bl[107] br[107] wl[464] vdd gnd cell_6t
Xbit_r465_c107 bl[107] br[107] wl[465] vdd gnd cell_6t
Xbit_r466_c107 bl[107] br[107] wl[466] vdd gnd cell_6t
Xbit_r467_c107 bl[107] br[107] wl[467] vdd gnd cell_6t
Xbit_r468_c107 bl[107] br[107] wl[468] vdd gnd cell_6t
Xbit_r469_c107 bl[107] br[107] wl[469] vdd gnd cell_6t
Xbit_r470_c107 bl[107] br[107] wl[470] vdd gnd cell_6t
Xbit_r471_c107 bl[107] br[107] wl[471] vdd gnd cell_6t
Xbit_r472_c107 bl[107] br[107] wl[472] vdd gnd cell_6t
Xbit_r473_c107 bl[107] br[107] wl[473] vdd gnd cell_6t
Xbit_r474_c107 bl[107] br[107] wl[474] vdd gnd cell_6t
Xbit_r475_c107 bl[107] br[107] wl[475] vdd gnd cell_6t
Xbit_r476_c107 bl[107] br[107] wl[476] vdd gnd cell_6t
Xbit_r477_c107 bl[107] br[107] wl[477] vdd gnd cell_6t
Xbit_r478_c107 bl[107] br[107] wl[478] vdd gnd cell_6t
Xbit_r479_c107 bl[107] br[107] wl[479] vdd gnd cell_6t
Xbit_r480_c107 bl[107] br[107] wl[480] vdd gnd cell_6t
Xbit_r481_c107 bl[107] br[107] wl[481] vdd gnd cell_6t
Xbit_r482_c107 bl[107] br[107] wl[482] vdd gnd cell_6t
Xbit_r483_c107 bl[107] br[107] wl[483] vdd gnd cell_6t
Xbit_r484_c107 bl[107] br[107] wl[484] vdd gnd cell_6t
Xbit_r485_c107 bl[107] br[107] wl[485] vdd gnd cell_6t
Xbit_r486_c107 bl[107] br[107] wl[486] vdd gnd cell_6t
Xbit_r487_c107 bl[107] br[107] wl[487] vdd gnd cell_6t
Xbit_r488_c107 bl[107] br[107] wl[488] vdd gnd cell_6t
Xbit_r489_c107 bl[107] br[107] wl[489] vdd gnd cell_6t
Xbit_r490_c107 bl[107] br[107] wl[490] vdd gnd cell_6t
Xbit_r491_c107 bl[107] br[107] wl[491] vdd gnd cell_6t
Xbit_r492_c107 bl[107] br[107] wl[492] vdd gnd cell_6t
Xbit_r493_c107 bl[107] br[107] wl[493] vdd gnd cell_6t
Xbit_r494_c107 bl[107] br[107] wl[494] vdd gnd cell_6t
Xbit_r495_c107 bl[107] br[107] wl[495] vdd gnd cell_6t
Xbit_r496_c107 bl[107] br[107] wl[496] vdd gnd cell_6t
Xbit_r497_c107 bl[107] br[107] wl[497] vdd gnd cell_6t
Xbit_r498_c107 bl[107] br[107] wl[498] vdd gnd cell_6t
Xbit_r499_c107 bl[107] br[107] wl[499] vdd gnd cell_6t
Xbit_r500_c107 bl[107] br[107] wl[500] vdd gnd cell_6t
Xbit_r501_c107 bl[107] br[107] wl[501] vdd gnd cell_6t
Xbit_r502_c107 bl[107] br[107] wl[502] vdd gnd cell_6t
Xbit_r503_c107 bl[107] br[107] wl[503] vdd gnd cell_6t
Xbit_r504_c107 bl[107] br[107] wl[504] vdd gnd cell_6t
Xbit_r505_c107 bl[107] br[107] wl[505] vdd gnd cell_6t
Xbit_r506_c107 bl[107] br[107] wl[506] vdd gnd cell_6t
Xbit_r507_c107 bl[107] br[107] wl[507] vdd gnd cell_6t
Xbit_r508_c107 bl[107] br[107] wl[508] vdd gnd cell_6t
Xbit_r509_c107 bl[107] br[107] wl[509] vdd gnd cell_6t
Xbit_r510_c107 bl[107] br[107] wl[510] vdd gnd cell_6t
Xbit_r511_c107 bl[107] br[107] wl[511] vdd gnd cell_6t
Xbit_r0_c108 bl[108] br[108] wl[0] vdd gnd cell_6t
Xbit_r1_c108 bl[108] br[108] wl[1] vdd gnd cell_6t
Xbit_r2_c108 bl[108] br[108] wl[2] vdd gnd cell_6t
Xbit_r3_c108 bl[108] br[108] wl[3] vdd gnd cell_6t
Xbit_r4_c108 bl[108] br[108] wl[4] vdd gnd cell_6t
Xbit_r5_c108 bl[108] br[108] wl[5] vdd gnd cell_6t
Xbit_r6_c108 bl[108] br[108] wl[6] vdd gnd cell_6t
Xbit_r7_c108 bl[108] br[108] wl[7] vdd gnd cell_6t
Xbit_r8_c108 bl[108] br[108] wl[8] vdd gnd cell_6t
Xbit_r9_c108 bl[108] br[108] wl[9] vdd gnd cell_6t
Xbit_r10_c108 bl[108] br[108] wl[10] vdd gnd cell_6t
Xbit_r11_c108 bl[108] br[108] wl[11] vdd gnd cell_6t
Xbit_r12_c108 bl[108] br[108] wl[12] vdd gnd cell_6t
Xbit_r13_c108 bl[108] br[108] wl[13] vdd gnd cell_6t
Xbit_r14_c108 bl[108] br[108] wl[14] vdd gnd cell_6t
Xbit_r15_c108 bl[108] br[108] wl[15] vdd gnd cell_6t
Xbit_r16_c108 bl[108] br[108] wl[16] vdd gnd cell_6t
Xbit_r17_c108 bl[108] br[108] wl[17] vdd gnd cell_6t
Xbit_r18_c108 bl[108] br[108] wl[18] vdd gnd cell_6t
Xbit_r19_c108 bl[108] br[108] wl[19] vdd gnd cell_6t
Xbit_r20_c108 bl[108] br[108] wl[20] vdd gnd cell_6t
Xbit_r21_c108 bl[108] br[108] wl[21] vdd gnd cell_6t
Xbit_r22_c108 bl[108] br[108] wl[22] vdd gnd cell_6t
Xbit_r23_c108 bl[108] br[108] wl[23] vdd gnd cell_6t
Xbit_r24_c108 bl[108] br[108] wl[24] vdd gnd cell_6t
Xbit_r25_c108 bl[108] br[108] wl[25] vdd gnd cell_6t
Xbit_r26_c108 bl[108] br[108] wl[26] vdd gnd cell_6t
Xbit_r27_c108 bl[108] br[108] wl[27] vdd gnd cell_6t
Xbit_r28_c108 bl[108] br[108] wl[28] vdd gnd cell_6t
Xbit_r29_c108 bl[108] br[108] wl[29] vdd gnd cell_6t
Xbit_r30_c108 bl[108] br[108] wl[30] vdd gnd cell_6t
Xbit_r31_c108 bl[108] br[108] wl[31] vdd gnd cell_6t
Xbit_r32_c108 bl[108] br[108] wl[32] vdd gnd cell_6t
Xbit_r33_c108 bl[108] br[108] wl[33] vdd gnd cell_6t
Xbit_r34_c108 bl[108] br[108] wl[34] vdd gnd cell_6t
Xbit_r35_c108 bl[108] br[108] wl[35] vdd gnd cell_6t
Xbit_r36_c108 bl[108] br[108] wl[36] vdd gnd cell_6t
Xbit_r37_c108 bl[108] br[108] wl[37] vdd gnd cell_6t
Xbit_r38_c108 bl[108] br[108] wl[38] vdd gnd cell_6t
Xbit_r39_c108 bl[108] br[108] wl[39] vdd gnd cell_6t
Xbit_r40_c108 bl[108] br[108] wl[40] vdd gnd cell_6t
Xbit_r41_c108 bl[108] br[108] wl[41] vdd gnd cell_6t
Xbit_r42_c108 bl[108] br[108] wl[42] vdd gnd cell_6t
Xbit_r43_c108 bl[108] br[108] wl[43] vdd gnd cell_6t
Xbit_r44_c108 bl[108] br[108] wl[44] vdd gnd cell_6t
Xbit_r45_c108 bl[108] br[108] wl[45] vdd gnd cell_6t
Xbit_r46_c108 bl[108] br[108] wl[46] vdd gnd cell_6t
Xbit_r47_c108 bl[108] br[108] wl[47] vdd gnd cell_6t
Xbit_r48_c108 bl[108] br[108] wl[48] vdd gnd cell_6t
Xbit_r49_c108 bl[108] br[108] wl[49] vdd gnd cell_6t
Xbit_r50_c108 bl[108] br[108] wl[50] vdd gnd cell_6t
Xbit_r51_c108 bl[108] br[108] wl[51] vdd gnd cell_6t
Xbit_r52_c108 bl[108] br[108] wl[52] vdd gnd cell_6t
Xbit_r53_c108 bl[108] br[108] wl[53] vdd gnd cell_6t
Xbit_r54_c108 bl[108] br[108] wl[54] vdd gnd cell_6t
Xbit_r55_c108 bl[108] br[108] wl[55] vdd gnd cell_6t
Xbit_r56_c108 bl[108] br[108] wl[56] vdd gnd cell_6t
Xbit_r57_c108 bl[108] br[108] wl[57] vdd gnd cell_6t
Xbit_r58_c108 bl[108] br[108] wl[58] vdd gnd cell_6t
Xbit_r59_c108 bl[108] br[108] wl[59] vdd gnd cell_6t
Xbit_r60_c108 bl[108] br[108] wl[60] vdd gnd cell_6t
Xbit_r61_c108 bl[108] br[108] wl[61] vdd gnd cell_6t
Xbit_r62_c108 bl[108] br[108] wl[62] vdd gnd cell_6t
Xbit_r63_c108 bl[108] br[108] wl[63] vdd gnd cell_6t
Xbit_r64_c108 bl[108] br[108] wl[64] vdd gnd cell_6t
Xbit_r65_c108 bl[108] br[108] wl[65] vdd gnd cell_6t
Xbit_r66_c108 bl[108] br[108] wl[66] vdd gnd cell_6t
Xbit_r67_c108 bl[108] br[108] wl[67] vdd gnd cell_6t
Xbit_r68_c108 bl[108] br[108] wl[68] vdd gnd cell_6t
Xbit_r69_c108 bl[108] br[108] wl[69] vdd gnd cell_6t
Xbit_r70_c108 bl[108] br[108] wl[70] vdd gnd cell_6t
Xbit_r71_c108 bl[108] br[108] wl[71] vdd gnd cell_6t
Xbit_r72_c108 bl[108] br[108] wl[72] vdd gnd cell_6t
Xbit_r73_c108 bl[108] br[108] wl[73] vdd gnd cell_6t
Xbit_r74_c108 bl[108] br[108] wl[74] vdd gnd cell_6t
Xbit_r75_c108 bl[108] br[108] wl[75] vdd gnd cell_6t
Xbit_r76_c108 bl[108] br[108] wl[76] vdd gnd cell_6t
Xbit_r77_c108 bl[108] br[108] wl[77] vdd gnd cell_6t
Xbit_r78_c108 bl[108] br[108] wl[78] vdd gnd cell_6t
Xbit_r79_c108 bl[108] br[108] wl[79] vdd gnd cell_6t
Xbit_r80_c108 bl[108] br[108] wl[80] vdd gnd cell_6t
Xbit_r81_c108 bl[108] br[108] wl[81] vdd gnd cell_6t
Xbit_r82_c108 bl[108] br[108] wl[82] vdd gnd cell_6t
Xbit_r83_c108 bl[108] br[108] wl[83] vdd gnd cell_6t
Xbit_r84_c108 bl[108] br[108] wl[84] vdd gnd cell_6t
Xbit_r85_c108 bl[108] br[108] wl[85] vdd gnd cell_6t
Xbit_r86_c108 bl[108] br[108] wl[86] vdd gnd cell_6t
Xbit_r87_c108 bl[108] br[108] wl[87] vdd gnd cell_6t
Xbit_r88_c108 bl[108] br[108] wl[88] vdd gnd cell_6t
Xbit_r89_c108 bl[108] br[108] wl[89] vdd gnd cell_6t
Xbit_r90_c108 bl[108] br[108] wl[90] vdd gnd cell_6t
Xbit_r91_c108 bl[108] br[108] wl[91] vdd gnd cell_6t
Xbit_r92_c108 bl[108] br[108] wl[92] vdd gnd cell_6t
Xbit_r93_c108 bl[108] br[108] wl[93] vdd gnd cell_6t
Xbit_r94_c108 bl[108] br[108] wl[94] vdd gnd cell_6t
Xbit_r95_c108 bl[108] br[108] wl[95] vdd gnd cell_6t
Xbit_r96_c108 bl[108] br[108] wl[96] vdd gnd cell_6t
Xbit_r97_c108 bl[108] br[108] wl[97] vdd gnd cell_6t
Xbit_r98_c108 bl[108] br[108] wl[98] vdd gnd cell_6t
Xbit_r99_c108 bl[108] br[108] wl[99] vdd gnd cell_6t
Xbit_r100_c108 bl[108] br[108] wl[100] vdd gnd cell_6t
Xbit_r101_c108 bl[108] br[108] wl[101] vdd gnd cell_6t
Xbit_r102_c108 bl[108] br[108] wl[102] vdd gnd cell_6t
Xbit_r103_c108 bl[108] br[108] wl[103] vdd gnd cell_6t
Xbit_r104_c108 bl[108] br[108] wl[104] vdd gnd cell_6t
Xbit_r105_c108 bl[108] br[108] wl[105] vdd gnd cell_6t
Xbit_r106_c108 bl[108] br[108] wl[106] vdd gnd cell_6t
Xbit_r107_c108 bl[108] br[108] wl[107] vdd gnd cell_6t
Xbit_r108_c108 bl[108] br[108] wl[108] vdd gnd cell_6t
Xbit_r109_c108 bl[108] br[108] wl[109] vdd gnd cell_6t
Xbit_r110_c108 bl[108] br[108] wl[110] vdd gnd cell_6t
Xbit_r111_c108 bl[108] br[108] wl[111] vdd gnd cell_6t
Xbit_r112_c108 bl[108] br[108] wl[112] vdd gnd cell_6t
Xbit_r113_c108 bl[108] br[108] wl[113] vdd gnd cell_6t
Xbit_r114_c108 bl[108] br[108] wl[114] vdd gnd cell_6t
Xbit_r115_c108 bl[108] br[108] wl[115] vdd gnd cell_6t
Xbit_r116_c108 bl[108] br[108] wl[116] vdd gnd cell_6t
Xbit_r117_c108 bl[108] br[108] wl[117] vdd gnd cell_6t
Xbit_r118_c108 bl[108] br[108] wl[118] vdd gnd cell_6t
Xbit_r119_c108 bl[108] br[108] wl[119] vdd gnd cell_6t
Xbit_r120_c108 bl[108] br[108] wl[120] vdd gnd cell_6t
Xbit_r121_c108 bl[108] br[108] wl[121] vdd gnd cell_6t
Xbit_r122_c108 bl[108] br[108] wl[122] vdd gnd cell_6t
Xbit_r123_c108 bl[108] br[108] wl[123] vdd gnd cell_6t
Xbit_r124_c108 bl[108] br[108] wl[124] vdd gnd cell_6t
Xbit_r125_c108 bl[108] br[108] wl[125] vdd gnd cell_6t
Xbit_r126_c108 bl[108] br[108] wl[126] vdd gnd cell_6t
Xbit_r127_c108 bl[108] br[108] wl[127] vdd gnd cell_6t
Xbit_r128_c108 bl[108] br[108] wl[128] vdd gnd cell_6t
Xbit_r129_c108 bl[108] br[108] wl[129] vdd gnd cell_6t
Xbit_r130_c108 bl[108] br[108] wl[130] vdd gnd cell_6t
Xbit_r131_c108 bl[108] br[108] wl[131] vdd gnd cell_6t
Xbit_r132_c108 bl[108] br[108] wl[132] vdd gnd cell_6t
Xbit_r133_c108 bl[108] br[108] wl[133] vdd gnd cell_6t
Xbit_r134_c108 bl[108] br[108] wl[134] vdd gnd cell_6t
Xbit_r135_c108 bl[108] br[108] wl[135] vdd gnd cell_6t
Xbit_r136_c108 bl[108] br[108] wl[136] vdd gnd cell_6t
Xbit_r137_c108 bl[108] br[108] wl[137] vdd gnd cell_6t
Xbit_r138_c108 bl[108] br[108] wl[138] vdd gnd cell_6t
Xbit_r139_c108 bl[108] br[108] wl[139] vdd gnd cell_6t
Xbit_r140_c108 bl[108] br[108] wl[140] vdd gnd cell_6t
Xbit_r141_c108 bl[108] br[108] wl[141] vdd gnd cell_6t
Xbit_r142_c108 bl[108] br[108] wl[142] vdd gnd cell_6t
Xbit_r143_c108 bl[108] br[108] wl[143] vdd gnd cell_6t
Xbit_r144_c108 bl[108] br[108] wl[144] vdd gnd cell_6t
Xbit_r145_c108 bl[108] br[108] wl[145] vdd gnd cell_6t
Xbit_r146_c108 bl[108] br[108] wl[146] vdd gnd cell_6t
Xbit_r147_c108 bl[108] br[108] wl[147] vdd gnd cell_6t
Xbit_r148_c108 bl[108] br[108] wl[148] vdd gnd cell_6t
Xbit_r149_c108 bl[108] br[108] wl[149] vdd gnd cell_6t
Xbit_r150_c108 bl[108] br[108] wl[150] vdd gnd cell_6t
Xbit_r151_c108 bl[108] br[108] wl[151] vdd gnd cell_6t
Xbit_r152_c108 bl[108] br[108] wl[152] vdd gnd cell_6t
Xbit_r153_c108 bl[108] br[108] wl[153] vdd gnd cell_6t
Xbit_r154_c108 bl[108] br[108] wl[154] vdd gnd cell_6t
Xbit_r155_c108 bl[108] br[108] wl[155] vdd gnd cell_6t
Xbit_r156_c108 bl[108] br[108] wl[156] vdd gnd cell_6t
Xbit_r157_c108 bl[108] br[108] wl[157] vdd gnd cell_6t
Xbit_r158_c108 bl[108] br[108] wl[158] vdd gnd cell_6t
Xbit_r159_c108 bl[108] br[108] wl[159] vdd gnd cell_6t
Xbit_r160_c108 bl[108] br[108] wl[160] vdd gnd cell_6t
Xbit_r161_c108 bl[108] br[108] wl[161] vdd gnd cell_6t
Xbit_r162_c108 bl[108] br[108] wl[162] vdd gnd cell_6t
Xbit_r163_c108 bl[108] br[108] wl[163] vdd gnd cell_6t
Xbit_r164_c108 bl[108] br[108] wl[164] vdd gnd cell_6t
Xbit_r165_c108 bl[108] br[108] wl[165] vdd gnd cell_6t
Xbit_r166_c108 bl[108] br[108] wl[166] vdd gnd cell_6t
Xbit_r167_c108 bl[108] br[108] wl[167] vdd gnd cell_6t
Xbit_r168_c108 bl[108] br[108] wl[168] vdd gnd cell_6t
Xbit_r169_c108 bl[108] br[108] wl[169] vdd gnd cell_6t
Xbit_r170_c108 bl[108] br[108] wl[170] vdd gnd cell_6t
Xbit_r171_c108 bl[108] br[108] wl[171] vdd gnd cell_6t
Xbit_r172_c108 bl[108] br[108] wl[172] vdd gnd cell_6t
Xbit_r173_c108 bl[108] br[108] wl[173] vdd gnd cell_6t
Xbit_r174_c108 bl[108] br[108] wl[174] vdd gnd cell_6t
Xbit_r175_c108 bl[108] br[108] wl[175] vdd gnd cell_6t
Xbit_r176_c108 bl[108] br[108] wl[176] vdd gnd cell_6t
Xbit_r177_c108 bl[108] br[108] wl[177] vdd gnd cell_6t
Xbit_r178_c108 bl[108] br[108] wl[178] vdd gnd cell_6t
Xbit_r179_c108 bl[108] br[108] wl[179] vdd gnd cell_6t
Xbit_r180_c108 bl[108] br[108] wl[180] vdd gnd cell_6t
Xbit_r181_c108 bl[108] br[108] wl[181] vdd gnd cell_6t
Xbit_r182_c108 bl[108] br[108] wl[182] vdd gnd cell_6t
Xbit_r183_c108 bl[108] br[108] wl[183] vdd gnd cell_6t
Xbit_r184_c108 bl[108] br[108] wl[184] vdd gnd cell_6t
Xbit_r185_c108 bl[108] br[108] wl[185] vdd gnd cell_6t
Xbit_r186_c108 bl[108] br[108] wl[186] vdd gnd cell_6t
Xbit_r187_c108 bl[108] br[108] wl[187] vdd gnd cell_6t
Xbit_r188_c108 bl[108] br[108] wl[188] vdd gnd cell_6t
Xbit_r189_c108 bl[108] br[108] wl[189] vdd gnd cell_6t
Xbit_r190_c108 bl[108] br[108] wl[190] vdd gnd cell_6t
Xbit_r191_c108 bl[108] br[108] wl[191] vdd gnd cell_6t
Xbit_r192_c108 bl[108] br[108] wl[192] vdd gnd cell_6t
Xbit_r193_c108 bl[108] br[108] wl[193] vdd gnd cell_6t
Xbit_r194_c108 bl[108] br[108] wl[194] vdd gnd cell_6t
Xbit_r195_c108 bl[108] br[108] wl[195] vdd gnd cell_6t
Xbit_r196_c108 bl[108] br[108] wl[196] vdd gnd cell_6t
Xbit_r197_c108 bl[108] br[108] wl[197] vdd gnd cell_6t
Xbit_r198_c108 bl[108] br[108] wl[198] vdd gnd cell_6t
Xbit_r199_c108 bl[108] br[108] wl[199] vdd gnd cell_6t
Xbit_r200_c108 bl[108] br[108] wl[200] vdd gnd cell_6t
Xbit_r201_c108 bl[108] br[108] wl[201] vdd gnd cell_6t
Xbit_r202_c108 bl[108] br[108] wl[202] vdd gnd cell_6t
Xbit_r203_c108 bl[108] br[108] wl[203] vdd gnd cell_6t
Xbit_r204_c108 bl[108] br[108] wl[204] vdd gnd cell_6t
Xbit_r205_c108 bl[108] br[108] wl[205] vdd gnd cell_6t
Xbit_r206_c108 bl[108] br[108] wl[206] vdd gnd cell_6t
Xbit_r207_c108 bl[108] br[108] wl[207] vdd gnd cell_6t
Xbit_r208_c108 bl[108] br[108] wl[208] vdd gnd cell_6t
Xbit_r209_c108 bl[108] br[108] wl[209] vdd gnd cell_6t
Xbit_r210_c108 bl[108] br[108] wl[210] vdd gnd cell_6t
Xbit_r211_c108 bl[108] br[108] wl[211] vdd gnd cell_6t
Xbit_r212_c108 bl[108] br[108] wl[212] vdd gnd cell_6t
Xbit_r213_c108 bl[108] br[108] wl[213] vdd gnd cell_6t
Xbit_r214_c108 bl[108] br[108] wl[214] vdd gnd cell_6t
Xbit_r215_c108 bl[108] br[108] wl[215] vdd gnd cell_6t
Xbit_r216_c108 bl[108] br[108] wl[216] vdd gnd cell_6t
Xbit_r217_c108 bl[108] br[108] wl[217] vdd gnd cell_6t
Xbit_r218_c108 bl[108] br[108] wl[218] vdd gnd cell_6t
Xbit_r219_c108 bl[108] br[108] wl[219] vdd gnd cell_6t
Xbit_r220_c108 bl[108] br[108] wl[220] vdd gnd cell_6t
Xbit_r221_c108 bl[108] br[108] wl[221] vdd gnd cell_6t
Xbit_r222_c108 bl[108] br[108] wl[222] vdd gnd cell_6t
Xbit_r223_c108 bl[108] br[108] wl[223] vdd gnd cell_6t
Xbit_r224_c108 bl[108] br[108] wl[224] vdd gnd cell_6t
Xbit_r225_c108 bl[108] br[108] wl[225] vdd gnd cell_6t
Xbit_r226_c108 bl[108] br[108] wl[226] vdd gnd cell_6t
Xbit_r227_c108 bl[108] br[108] wl[227] vdd gnd cell_6t
Xbit_r228_c108 bl[108] br[108] wl[228] vdd gnd cell_6t
Xbit_r229_c108 bl[108] br[108] wl[229] vdd gnd cell_6t
Xbit_r230_c108 bl[108] br[108] wl[230] vdd gnd cell_6t
Xbit_r231_c108 bl[108] br[108] wl[231] vdd gnd cell_6t
Xbit_r232_c108 bl[108] br[108] wl[232] vdd gnd cell_6t
Xbit_r233_c108 bl[108] br[108] wl[233] vdd gnd cell_6t
Xbit_r234_c108 bl[108] br[108] wl[234] vdd gnd cell_6t
Xbit_r235_c108 bl[108] br[108] wl[235] vdd gnd cell_6t
Xbit_r236_c108 bl[108] br[108] wl[236] vdd gnd cell_6t
Xbit_r237_c108 bl[108] br[108] wl[237] vdd gnd cell_6t
Xbit_r238_c108 bl[108] br[108] wl[238] vdd gnd cell_6t
Xbit_r239_c108 bl[108] br[108] wl[239] vdd gnd cell_6t
Xbit_r240_c108 bl[108] br[108] wl[240] vdd gnd cell_6t
Xbit_r241_c108 bl[108] br[108] wl[241] vdd gnd cell_6t
Xbit_r242_c108 bl[108] br[108] wl[242] vdd gnd cell_6t
Xbit_r243_c108 bl[108] br[108] wl[243] vdd gnd cell_6t
Xbit_r244_c108 bl[108] br[108] wl[244] vdd gnd cell_6t
Xbit_r245_c108 bl[108] br[108] wl[245] vdd gnd cell_6t
Xbit_r246_c108 bl[108] br[108] wl[246] vdd gnd cell_6t
Xbit_r247_c108 bl[108] br[108] wl[247] vdd gnd cell_6t
Xbit_r248_c108 bl[108] br[108] wl[248] vdd gnd cell_6t
Xbit_r249_c108 bl[108] br[108] wl[249] vdd gnd cell_6t
Xbit_r250_c108 bl[108] br[108] wl[250] vdd gnd cell_6t
Xbit_r251_c108 bl[108] br[108] wl[251] vdd gnd cell_6t
Xbit_r252_c108 bl[108] br[108] wl[252] vdd gnd cell_6t
Xbit_r253_c108 bl[108] br[108] wl[253] vdd gnd cell_6t
Xbit_r254_c108 bl[108] br[108] wl[254] vdd gnd cell_6t
Xbit_r255_c108 bl[108] br[108] wl[255] vdd gnd cell_6t
Xbit_r256_c108 bl[108] br[108] wl[256] vdd gnd cell_6t
Xbit_r257_c108 bl[108] br[108] wl[257] vdd gnd cell_6t
Xbit_r258_c108 bl[108] br[108] wl[258] vdd gnd cell_6t
Xbit_r259_c108 bl[108] br[108] wl[259] vdd gnd cell_6t
Xbit_r260_c108 bl[108] br[108] wl[260] vdd gnd cell_6t
Xbit_r261_c108 bl[108] br[108] wl[261] vdd gnd cell_6t
Xbit_r262_c108 bl[108] br[108] wl[262] vdd gnd cell_6t
Xbit_r263_c108 bl[108] br[108] wl[263] vdd gnd cell_6t
Xbit_r264_c108 bl[108] br[108] wl[264] vdd gnd cell_6t
Xbit_r265_c108 bl[108] br[108] wl[265] vdd gnd cell_6t
Xbit_r266_c108 bl[108] br[108] wl[266] vdd gnd cell_6t
Xbit_r267_c108 bl[108] br[108] wl[267] vdd gnd cell_6t
Xbit_r268_c108 bl[108] br[108] wl[268] vdd gnd cell_6t
Xbit_r269_c108 bl[108] br[108] wl[269] vdd gnd cell_6t
Xbit_r270_c108 bl[108] br[108] wl[270] vdd gnd cell_6t
Xbit_r271_c108 bl[108] br[108] wl[271] vdd gnd cell_6t
Xbit_r272_c108 bl[108] br[108] wl[272] vdd gnd cell_6t
Xbit_r273_c108 bl[108] br[108] wl[273] vdd gnd cell_6t
Xbit_r274_c108 bl[108] br[108] wl[274] vdd gnd cell_6t
Xbit_r275_c108 bl[108] br[108] wl[275] vdd gnd cell_6t
Xbit_r276_c108 bl[108] br[108] wl[276] vdd gnd cell_6t
Xbit_r277_c108 bl[108] br[108] wl[277] vdd gnd cell_6t
Xbit_r278_c108 bl[108] br[108] wl[278] vdd gnd cell_6t
Xbit_r279_c108 bl[108] br[108] wl[279] vdd gnd cell_6t
Xbit_r280_c108 bl[108] br[108] wl[280] vdd gnd cell_6t
Xbit_r281_c108 bl[108] br[108] wl[281] vdd gnd cell_6t
Xbit_r282_c108 bl[108] br[108] wl[282] vdd gnd cell_6t
Xbit_r283_c108 bl[108] br[108] wl[283] vdd gnd cell_6t
Xbit_r284_c108 bl[108] br[108] wl[284] vdd gnd cell_6t
Xbit_r285_c108 bl[108] br[108] wl[285] vdd gnd cell_6t
Xbit_r286_c108 bl[108] br[108] wl[286] vdd gnd cell_6t
Xbit_r287_c108 bl[108] br[108] wl[287] vdd gnd cell_6t
Xbit_r288_c108 bl[108] br[108] wl[288] vdd gnd cell_6t
Xbit_r289_c108 bl[108] br[108] wl[289] vdd gnd cell_6t
Xbit_r290_c108 bl[108] br[108] wl[290] vdd gnd cell_6t
Xbit_r291_c108 bl[108] br[108] wl[291] vdd gnd cell_6t
Xbit_r292_c108 bl[108] br[108] wl[292] vdd gnd cell_6t
Xbit_r293_c108 bl[108] br[108] wl[293] vdd gnd cell_6t
Xbit_r294_c108 bl[108] br[108] wl[294] vdd gnd cell_6t
Xbit_r295_c108 bl[108] br[108] wl[295] vdd gnd cell_6t
Xbit_r296_c108 bl[108] br[108] wl[296] vdd gnd cell_6t
Xbit_r297_c108 bl[108] br[108] wl[297] vdd gnd cell_6t
Xbit_r298_c108 bl[108] br[108] wl[298] vdd gnd cell_6t
Xbit_r299_c108 bl[108] br[108] wl[299] vdd gnd cell_6t
Xbit_r300_c108 bl[108] br[108] wl[300] vdd gnd cell_6t
Xbit_r301_c108 bl[108] br[108] wl[301] vdd gnd cell_6t
Xbit_r302_c108 bl[108] br[108] wl[302] vdd gnd cell_6t
Xbit_r303_c108 bl[108] br[108] wl[303] vdd gnd cell_6t
Xbit_r304_c108 bl[108] br[108] wl[304] vdd gnd cell_6t
Xbit_r305_c108 bl[108] br[108] wl[305] vdd gnd cell_6t
Xbit_r306_c108 bl[108] br[108] wl[306] vdd gnd cell_6t
Xbit_r307_c108 bl[108] br[108] wl[307] vdd gnd cell_6t
Xbit_r308_c108 bl[108] br[108] wl[308] vdd gnd cell_6t
Xbit_r309_c108 bl[108] br[108] wl[309] vdd gnd cell_6t
Xbit_r310_c108 bl[108] br[108] wl[310] vdd gnd cell_6t
Xbit_r311_c108 bl[108] br[108] wl[311] vdd gnd cell_6t
Xbit_r312_c108 bl[108] br[108] wl[312] vdd gnd cell_6t
Xbit_r313_c108 bl[108] br[108] wl[313] vdd gnd cell_6t
Xbit_r314_c108 bl[108] br[108] wl[314] vdd gnd cell_6t
Xbit_r315_c108 bl[108] br[108] wl[315] vdd gnd cell_6t
Xbit_r316_c108 bl[108] br[108] wl[316] vdd gnd cell_6t
Xbit_r317_c108 bl[108] br[108] wl[317] vdd gnd cell_6t
Xbit_r318_c108 bl[108] br[108] wl[318] vdd gnd cell_6t
Xbit_r319_c108 bl[108] br[108] wl[319] vdd gnd cell_6t
Xbit_r320_c108 bl[108] br[108] wl[320] vdd gnd cell_6t
Xbit_r321_c108 bl[108] br[108] wl[321] vdd gnd cell_6t
Xbit_r322_c108 bl[108] br[108] wl[322] vdd gnd cell_6t
Xbit_r323_c108 bl[108] br[108] wl[323] vdd gnd cell_6t
Xbit_r324_c108 bl[108] br[108] wl[324] vdd gnd cell_6t
Xbit_r325_c108 bl[108] br[108] wl[325] vdd gnd cell_6t
Xbit_r326_c108 bl[108] br[108] wl[326] vdd gnd cell_6t
Xbit_r327_c108 bl[108] br[108] wl[327] vdd gnd cell_6t
Xbit_r328_c108 bl[108] br[108] wl[328] vdd gnd cell_6t
Xbit_r329_c108 bl[108] br[108] wl[329] vdd gnd cell_6t
Xbit_r330_c108 bl[108] br[108] wl[330] vdd gnd cell_6t
Xbit_r331_c108 bl[108] br[108] wl[331] vdd gnd cell_6t
Xbit_r332_c108 bl[108] br[108] wl[332] vdd gnd cell_6t
Xbit_r333_c108 bl[108] br[108] wl[333] vdd gnd cell_6t
Xbit_r334_c108 bl[108] br[108] wl[334] vdd gnd cell_6t
Xbit_r335_c108 bl[108] br[108] wl[335] vdd gnd cell_6t
Xbit_r336_c108 bl[108] br[108] wl[336] vdd gnd cell_6t
Xbit_r337_c108 bl[108] br[108] wl[337] vdd gnd cell_6t
Xbit_r338_c108 bl[108] br[108] wl[338] vdd gnd cell_6t
Xbit_r339_c108 bl[108] br[108] wl[339] vdd gnd cell_6t
Xbit_r340_c108 bl[108] br[108] wl[340] vdd gnd cell_6t
Xbit_r341_c108 bl[108] br[108] wl[341] vdd gnd cell_6t
Xbit_r342_c108 bl[108] br[108] wl[342] vdd gnd cell_6t
Xbit_r343_c108 bl[108] br[108] wl[343] vdd gnd cell_6t
Xbit_r344_c108 bl[108] br[108] wl[344] vdd gnd cell_6t
Xbit_r345_c108 bl[108] br[108] wl[345] vdd gnd cell_6t
Xbit_r346_c108 bl[108] br[108] wl[346] vdd gnd cell_6t
Xbit_r347_c108 bl[108] br[108] wl[347] vdd gnd cell_6t
Xbit_r348_c108 bl[108] br[108] wl[348] vdd gnd cell_6t
Xbit_r349_c108 bl[108] br[108] wl[349] vdd gnd cell_6t
Xbit_r350_c108 bl[108] br[108] wl[350] vdd gnd cell_6t
Xbit_r351_c108 bl[108] br[108] wl[351] vdd gnd cell_6t
Xbit_r352_c108 bl[108] br[108] wl[352] vdd gnd cell_6t
Xbit_r353_c108 bl[108] br[108] wl[353] vdd gnd cell_6t
Xbit_r354_c108 bl[108] br[108] wl[354] vdd gnd cell_6t
Xbit_r355_c108 bl[108] br[108] wl[355] vdd gnd cell_6t
Xbit_r356_c108 bl[108] br[108] wl[356] vdd gnd cell_6t
Xbit_r357_c108 bl[108] br[108] wl[357] vdd gnd cell_6t
Xbit_r358_c108 bl[108] br[108] wl[358] vdd gnd cell_6t
Xbit_r359_c108 bl[108] br[108] wl[359] vdd gnd cell_6t
Xbit_r360_c108 bl[108] br[108] wl[360] vdd gnd cell_6t
Xbit_r361_c108 bl[108] br[108] wl[361] vdd gnd cell_6t
Xbit_r362_c108 bl[108] br[108] wl[362] vdd gnd cell_6t
Xbit_r363_c108 bl[108] br[108] wl[363] vdd gnd cell_6t
Xbit_r364_c108 bl[108] br[108] wl[364] vdd gnd cell_6t
Xbit_r365_c108 bl[108] br[108] wl[365] vdd gnd cell_6t
Xbit_r366_c108 bl[108] br[108] wl[366] vdd gnd cell_6t
Xbit_r367_c108 bl[108] br[108] wl[367] vdd gnd cell_6t
Xbit_r368_c108 bl[108] br[108] wl[368] vdd gnd cell_6t
Xbit_r369_c108 bl[108] br[108] wl[369] vdd gnd cell_6t
Xbit_r370_c108 bl[108] br[108] wl[370] vdd gnd cell_6t
Xbit_r371_c108 bl[108] br[108] wl[371] vdd gnd cell_6t
Xbit_r372_c108 bl[108] br[108] wl[372] vdd gnd cell_6t
Xbit_r373_c108 bl[108] br[108] wl[373] vdd gnd cell_6t
Xbit_r374_c108 bl[108] br[108] wl[374] vdd gnd cell_6t
Xbit_r375_c108 bl[108] br[108] wl[375] vdd gnd cell_6t
Xbit_r376_c108 bl[108] br[108] wl[376] vdd gnd cell_6t
Xbit_r377_c108 bl[108] br[108] wl[377] vdd gnd cell_6t
Xbit_r378_c108 bl[108] br[108] wl[378] vdd gnd cell_6t
Xbit_r379_c108 bl[108] br[108] wl[379] vdd gnd cell_6t
Xbit_r380_c108 bl[108] br[108] wl[380] vdd gnd cell_6t
Xbit_r381_c108 bl[108] br[108] wl[381] vdd gnd cell_6t
Xbit_r382_c108 bl[108] br[108] wl[382] vdd gnd cell_6t
Xbit_r383_c108 bl[108] br[108] wl[383] vdd gnd cell_6t
Xbit_r384_c108 bl[108] br[108] wl[384] vdd gnd cell_6t
Xbit_r385_c108 bl[108] br[108] wl[385] vdd gnd cell_6t
Xbit_r386_c108 bl[108] br[108] wl[386] vdd gnd cell_6t
Xbit_r387_c108 bl[108] br[108] wl[387] vdd gnd cell_6t
Xbit_r388_c108 bl[108] br[108] wl[388] vdd gnd cell_6t
Xbit_r389_c108 bl[108] br[108] wl[389] vdd gnd cell_6t
Xbit_r390_c108 bl[108] br[108] wl[390] vdd gnd cell_6t
Xbit_r391_c108 bl[108] br[108] wl[391] vdd gnd cell_6t
Xbit_r392_c108 bl[108] br[108] wl[392] vdd gnd cell_6t
Xbit_r393_c108 bl[108] br[108] wl[393] vdd gnd cell_6t
Xbit_r394_c108 bl[108] br[108] wl[394] vdd gnd cell_6t
Xbit_r395_c108 bl[108] br[108] wl[395] vdd gnd cell_6t
Xbit_r396_c108 bl[108] br[108] wl[396] vdd gnd cell_6t
Xbit_r397_c108 bl[108] br[108] wl[397] vdd gnd cell_6t
Xbit_r398_c108 bl[108] br[108] wl[398] vdd gnd cell_6t
Xbit_r399_c108 bl[108] br[108] wl[399] vdd gnd cell_6t
Xbit_r400_c108 bl[108] br[108] wl[400] vdd gnd cell_6t
Xbit_r401_c108 bl[108] br[108] wl[401] vdd gnd cell_6t
Xbit_r402_c108 bl[108] br[108] wl[402] vdd gnd cell_6t
Xbit_r403_c108 bl[108] br[108] wl[403] vdd gnd cell_6t
Xbit_r404_c108 bl[108] br[108] wl[404] vdd gnd cell_6t
Xbit_r405_c108 bl[108] br[108] wl[405] vdd gnd cell_6t
Xbit_r406_c108 bl[108] br[108] wl[406] vdd gnd cell_6t
Xbit_r407_c108 bl[108] br[108] wl[407] vdd gnd cell_6t
Xbit_r408_c108 bl[108] br[108] wl[408] vdd gnd cell_6t
Xbit_r409_c108 bl[108] br[108] wl[409] vdd gnd cell_6t
Xbit_r410_c108 bl[108] br[108] wl[410] vdd gnd cell_6t
Xbit_r411_c108 bl[108] br[108] wl[411] vdd gnd cell_6t
Xbit_r412_c108 bl[108] br[108] wl[412] vdd gnd cell_6t
Xbit_r413_c108 bl[108] br[108] wl[413] vdd gnd cell_6t
Xbit_r414_c108 bl[108] br[108] wl[414] vdd gnd cell_6t
Xbit_r415_c108 bl[108] br[108] wl[415] vdd gnd cell_6t
Xbit_r416_c108 bl[108] br[108] wl[416] vdd gnd cell_6t
Xbit_r417_c108 bl[108] br[108] wl[417] vdd gnd cell_6t
Xbit_r418_c108 bl[108] br[108] wl[418] vdd gnd cell_6t
Xbit_r419_c108 bl[108] br[108] wl[419] vdd gnd cell_6t
Xbit_r420_c108 bl[108] br[108] wl[420] vdd gnd cell_6t
Xbit_r421_c108 bl[108] br[108] wl[421] vdd gnd cell_6t
Xbit_r422_c108 bl[108] br[108] wl[422] vdd gnd cell_6t
Xbit_r423_c108 bl[108] br[108] wl[423] vdd gnd cell_6t
Xbit_r424_c108 bl[108] br[108] wl[424] vdd gnd cell_6t
Xbit_r425_c108 bl[108] br[108] wl[425] vdd gnd cell_6t
Xbit_r426_c108 bl[108] br[108] wl[426] vdd gnd cell_6t
Xbit_r427_c108 bl[108] br[108] wl[427] vdd gnd cell_6t
Xbit_r428_c108 bl[108] br[108] wl[428] vdd gnd cell_6t
Xbit_r429_c108 bl[108] br[108] wl[429] vdd gnd cell_6t
Xbit_r430_c108 bl[108] br[108] wl[430] vdd gnd cell_6t
Xbit_r431_c108 bl[108] br[108] wl[431] vdd gnd cell_6t
Xbit_r432_c108 bl[108] br[108] wl[432] vdd gnd cell_6t
Xbit_r433_c108 bl[108] br[108] wl[433] vdd gnd cell_6t
Xbit_r434_c108 bl[108] br[108] wl[434] vdd gnd cell_6t
Xbit_r435_c108 bl[108] br[108] wl[435] vdd gnd cell_6t
Xbit_r436_c108 bl[108] br[108] wl[436] vdd gnd cell_6t
Xbit_r437_c108 bl[108] br[108] wl[437] vdd gnd cell_6t
Xbit_r438_c108 bl[108] br[108] wl[438] vdd gnd cell_6t
Xbit_r439_c108 bl[108] br[108] wl[439] vdd gnd cell_6t
Xbit_r440_c108 bl[108] br[108] wl[440] vdd gnd cell_6t
Xbit_r441_c108 bl[108] br[108] wl[441] vdd gnd cell_6t
Xbit_r442_c108 bl[108] br[108] wl[442] vdd gnd cell_6t
Xbit_r443_c108 bl[108] br[108] wl[443] vdd gnd cell_6t
Xbit_r444_c108 bl[108] br[108] wl[444] vdd gnd cell_6t
Xbit_r445_c108 bl[108] br[108] wl[445] vdd gnd cell_6t
Xbit_r446_c108 bl[108] br[108] wl[446] vdd gnd cell_6t
Xbit_r447_c108 bl[108] br[108] wl[447] vdd gnd cell_6t
Xbit_r448_c108 bl[108] br[108] wl[448] vdd gnd cell_6t
Xbit_r449_c108 bl[108] br[108] wl[449] vdd gnd cell_6t
Xbit_r450_c108 bl[108] br[108] wl[450] vdd gnd cell_6t
Xbit_r451_c108 bl[108] br[108] wl[451] vdd gnd cell_6t
Xbit_r452_c108 bl[108] br[108] wl[452] vdd gnd cell_6t
Xbit_r453_c108 bl[108] br[108] wl[453] vdd gnd cell_6t
Xbit_r454_c108 bl[108] br[108] wl[454] vdd gnd cell_6t
Xbit_r455_c108 bl[108] br[108] wl[455] vdd gnd cell_6t
Xbit_r456_c108 bl[108] br[108] wl[456] vdd gnd cell_6t
Xbit_r457_c108 bl[108] br[108] wl[457] vdd gnd cell_6t
Xbit_r458_c108 bl[108] br[108] wl[458] vdd gnd cell_6t
Xbit_r459_c108 bl[108] br[108] wl[459] vdd gnd cell_6t
Xbit_r460_c108 bl[108] br[108] wl[460] vdd gnd cell_6t
Xbit_r461_c108 bl[108] br[108] wl[461] vdd gnd cell_6t
Xbit_r462_c108 bl[108] br[108] wl[462] vdd gnd cell_6t
Xbit_r463_c108 bl[108] br[108] wl[463] vdd gnd cell_6t
Xbit_r464_c108 bl[108] br[108] wl[464] vdd gnd cell_6t
Xbit_r465_c108 bl[108] br[108] wl[465] vdd gnd cell_6t
Xbit_r466_c108 bl[108] br[108] wl[466] vdd gnd cell_6t
Xbit_r467_c108 bl[108] br[108] wl[467] vdd gnd cell_6t
Xbit_r468_c108 bl[108] br[108] wl[468] vdd gnd cell_6t
Xbit_r469_c108 bl[108] br[108] wl[469] vdd gnd cell_6t
Xbit_r470_c108 bl[108] br[108] wl[470] vdd gnd cell_6t
Xbit_r471_c108 bl[108] br[108] wl[471] vdd gnd cell_6t
Xbit_r472_c108 bl[108] br[108] wl[472] vdd gnd cell_6t
Xbit_r473_c108 bl[108] br[108] wl[473] vdd gnd cell_6t
Xbit_r474_c108 bl[108] br[108] wl[474] vdd gnd cell_6t
Xbit_r475_c108 bl[108] br[108] wl[475] vdd gnd cell_6t
Xbit_r476_c108 bl[108] br[108] wl[476] vdd gnd cell_6t
Xbit_r477_c108 bl[108] br[108] wl[477] vdd gnd cell_6t
Xbit_r478_c108 bl[108] br[108] wl[478] vdd gnd cell_6t
Xbit_r479_c108 bl[108] br[108] wl[479] vdd gnd cell_6t
Xbit_r480_c108 bl[108] br[108] wl[480] vdd gnd cell_6t
Xbit_r481_c108 bl[108] br[108] wl[481] vdd gnd cell_6t
Xbit_r482_c108 bl[108] br[108] wl[482] vdd gnd cell_6t
Xbit_r483_c108 bl[108] br[108] wl[483] vdd gnd cell_6t
Xbit_r484_c108 bl[108] br[108] wl[484] vdd gnd cell_6t
Xbit_r485_c108 bl[108] br[108] wl[485] vdd gnd cell_6t
Xbit_r486_c108 bl[108] br[108] wl[486] vdd gnd cell_6t
Xbit_r487_c108 bl[108] br[108] wl[487] vdd gnd cell_6t
Xbit_r488_c108 bl[108] br[108] wl[488] vdd gnd cell_6t
Xbit_r489_c108 bl[108] br[108] wl[489] vdd gnd cell_6t
Xbit_r490_c108 bl[108] br[108] wl[490] vdd gnd cell_6t
Xbit_r491_c108 bl[108] br[108] wl[491] vdd gnd cell_6t
Xbit_r492_c108 bl[108] br[108] wl[492] vdd gnd cell_6t
Xbit_r493_c108 bl[108] br[108] wl[493] vdd gnd cell_6t
Xbit_r494_c108 bl[108] br[108] wl[494] vdd gnd cell_6t
Xbit_r495_c108 bl[108] br[108] wl[495] vdd gnd cell_6t
Xbit_r496_c108 bl[108] br[108] wl[496] vdd gnd cell_6t
Xbit_r497_c108 bl[108] br[108] wl[497] vdd gnd cell_6t
Xbit_r498_c108 bl[108] br[108] wl[498] vdd gnd cell_6t
Xbit_r499_c108 bl[108] br[108] wl[499] vdd gnd cell_6t
Xbit_r500_c108 bl[108] br[108] wl[500] vdd gnd cell_6t
Xbit_r501_c108 bl[108] br[108] wl[501] vdd gnd cell_6t
Xbit_r502_c108 bl[108] br[108] wl[502] vdd gnd cell_6t
Xbit_r503_c108 bl[108] br[108] wl[503] vdd gnd cell_6t
Xbit_r504_c108 bl[108] br[108] wl[504] vdd gnd cell_6t
Xbit_r505_c108 bl[108] br[108] wl[505] vdd gnd cell_6t
Xbit_r506_c108 bl[108] br[108] wl[506] vdd gnd cell_6t
Xbit_r507_c108 bl[108] br[108] wl[507] vdd gnd cell_6t
Xbit_r508_c108 bl[108] br[108] wl[508] vdd gnd cell_6t
Xbit_r509_c108 bl[108] br[108] wl[509] vdd gnd cell_6t
Xbit_r510_c108 bl[108] br[108] wl[510] vdd gnd cell_6t
Xbit_r511_c108 bl[108] br[108] wl[511] vdd gnd cell_6t
Xbit_r0_c109 bl[109] br[109] wl[0] vdd gnd cell_6t
Xbit_r1_c109 bl[109] br[109] wl[1] vdd gnd cell_6t
Xbit_r2_c109 bl[109] br[109] wl[2] vdd gnd cell_6t
Xbit_r3_c109 bl[109] br[109] wl[3] vdd gnd cell_6t
Xbit_r4_c109 bl[109] br[109] wl[4] vdd gnd cell_6t
Xbit_r5_c109 bl[109] br[109] wl[5] vdd gnd cell_6t
Xbit_r6_c109 bl[109] br[109] wl[6] vdd gnd cell_6t
Xbit_r7_c109 bl[109] br[109] wl[7] vdd gnd cell_6t
Xbit_r8_c109 bl[109] br[109] wl[8] vdd gnd cell_6t
Xbit_r9_c109 bl[109] br[109] wl[9] vdd gnd cell_6t
Xbit_r10_c109 bl[109] br[109] wl[10] vdd gnd cell_6t
Xbit_r11_c109 bl[109] br[109] wl[11] vdd gnd cell_6t
Xbit_r12_c109 bl[109] br[109] wl[12] vdd gnd cell_6t
Xbit_r13_c109 bl[109] br[109] wl[13] vdd gnd cell_6t
Xbit_r14_c109 bl[109] br[109] wl[14] vdd gnd cell_6t
Xbit_r15_c109 bl[109] br[109] wl[15] vdd gnd cell_6t
Xbit_r16_c109 bl[109] br[109] wl[16] vdd gnd cell_6t
Xbit_r17_c109 bl[109] br[109] wl[17] vdd gnd cell_6t
Xbit_r18_c109 bl[109] br[109] wl[18] vdd gnd cell_6t
Xbit_r19_c109 bl[109] br[109] wl[19] vdd gnd cell_6t
Xbit_r20_c109 bl[109] br[109] wl[20] vdd gnd cell_6t
Xbit_r21_c109 bl[109] br[109] wl[21] vdd gnd cell_6t
Xbit_r22_c109 bl[109] br[109] wl[22] vdd gnd cell_6t
Xbit_r23_c109 bl[109] br[109] wl[23] vdd gnd cell_6t
Xbit_r24_c109 bl[109] br[109] wl[24] vdd gnd cell_6t
Xbit_r25_c109 bl[109] br[109] wl[25] vdd gnd cell_6t
Xbit_r26_c109 bl[109] br[109] wl[26] vdd gnd cell_6t
Xbit_r27_c109 bl[109] br[109] wl[27] vdd gnd cell_6t
Xbit_r28_c109 bl[109] br[109] wl[28] vdd gnd cell_6t
Xbit_r29_c109 bl[109] br[109] wl[29] vdd gnd cell_6t
Xbit_r30_c109 bl[109] br[109] wl[30] vdd gnd cell_6t
Xbit_r31_c109 bl[109] br[109] wl[31] vdd gnd cell_6t
Xbit_r32_c109 bl[109] br[109] wl[32] vdd gnd cell_6t
Xbit_r33_c109 bl[109] br[109] wl[33] vdd gnd cell_6t
Xbit_r34_c109 bl[109] br[109] wl[34] vdd gnd cell_6t
Xbit_r35_c109 bl[109] br[109] wl[35] vdd gnd cell_6t
Xbit_r36_c109 bl[109] br[109] wl[36] vdd gnd cell_6t
Xbit_r37_c109 bl[109] br[109] wl[37] vdd gnd cell_6t
Xbit_r38_c109 bl[109] br[109] wl[38] vdd gnd cell_6t
Xbit_r39_c109 bl[109] br[109] wl[39] vdd gnd cell_6t
Xbit_r40_c109 bl[109] br[109] wl[40] vdd gnd cell_6t
Xbit_r41_c109 bl[109] br[109] wl[41] vdd gnd cell_6t
Xbit_r42_c109 bl[109] br[109] wl[42] vdd gnd cell_6t
Xbit_r43_c109 bl[109] br[109] wl[43] vdd gnd cell_6t
Xbit_r44_c109 bl[109] br[109] wl[44] vdd gnd cell_6t
Xbit_r45_c109 bl[109] br[109] wl[45] vdd gnd cell_6t
Xbit_r46_c109 bl[109] br[109] wl[46] vdd gnd cell_6t
Xbit_r47_c109 bl[109] br[109] wl[47] vdd gnd cell_6t
Xbit_r48_c109 bl[109] br[109] wl[48] vdd gnd cell_6t
Xbit_r49_c109 bl[109] br[109] wl[49] vdd gnd cell_6t
Xbit_r50_c109 bl[109] br[109] wl[50] vdd gnd cell_6t
Xbit_r51_c109 bl[109] br[109] wl[51] vdd gnd cell_6t
Xbit_r52_c109 bl[109] br[109] wl[52] vdd gnd cell_6t
Xbit_r53_c109 bl[109] br[109] wl[53] vdd gnd cell_6t
Xbit_r54_c109 bl[109] br[109] wl[54] vdd gnd cell_6t
Xbit_r55_c109 bl[109] br[109] wl[55] vdd gnd cell_6t
Xbit_r56_c109 bl[109] br[109] wl[56] vdd gnd cell_6t
Xbit_r57_c109 bl[109] br[109] wl[57] vdd gnd cell_6t
Xbit_r58_c109 bl[109] br[109] wl[58] vdd gnd cell_6t
Xbit_r59_c109 bl[109] br[109] wl[59] vdd gnd cell_6t
Xbit_r60_c109 bl[109] br[109] wl[60] vdd gnd cell_6t
Xbit_r61_c109 bl[109] br[109] wl[61] vdd gnd cell_6t
Xbit_r62_c109 bl[109] br[109] wl[62] vdd gnd cell_6t
Xbit_r63_c109 bl[109] br[109] wl[63] vdd gnd cell_6t
Xbit_r64_c109 bl[109] br[109] wl[64] vdd gnd cell_6t
Xbit_r65_c109 bl[109] br[109] wl[65] vdd gnd cell_6t
Xbit_r66_c109 bl[109] br[109] wl[66] vdd gnd cell_6t
Xbit_r67_c109 bl[109] br[109] wl[67] vdd gnd cell_6t
Xbit_r68_c109 bl[109] br[109] wl[68] vdd gnd cell_6t
Xbit_r69_c109 bl[109] br[109] wl[69] vdd gnd cell_6t
Xbit_r70_c109 bl[109] br[109] wl[70] vdd gnd cell_6t
Xbit_r71_c109 bl[109] br[109] wl[71] vdd gnd cell_6t
Xbit_r72_c109 bl[109] br[109] wl[72] vdd gnd cell_6t
Xbit_r73_c109 bl[109] br[109] wl[73] vdd gnd cell_6t
Xbit_r74_c109 bl[109] br[109] wl[74] vdd gnd cell_6t
Xbit_r75_c109 bl[109] br[109] wl[75] vdd gnd cell_6t
Xbit_r76_c109 bl[109] br[109] wl[76] vdd gnd cell_6t
Xbit_r77_c109 bl[109] br[109] wl[77] vdd gnd cell_6t
Xbit_r78_c109 bl[109] br[109] wl[78] vdd gnd cell_6t
Xbit_r79_c109 bl[109] br[109] wl[79] vdd gnd cell_6t
Xbit_r80_c109 bl[109] br[109] wl[80] vdd gnd cell_6t
Xbit_r81_c109 bl[109] br[109] wl[81] vdd gnd cell_6t
Xbit_r82_c109 bl[109] br[109] wl[82] vdd gnd cell_6t
Xbit_r83_c109 bl[109] br[109] wl[83] vdd gnd cell_6t
Xbit_r84_c109 bl[109] br[109] wl[84] vdd gnd cell_6t
Xbit_r85_c109 bl[109] br[109] wl[85] vdd gnd cell_6t
Xbit_r86_c109 bl[109] br[109] wl[86] vdd gnd cell_6t
Xbit_r87_c109 bl[109] br[109] wl[87] vdd gnd cell_6t
Xbit_r88_c109 bl[109] br[109] wl[88] vdd gnd cell_6t
Xbit_r89_c109 bl[109] br[109] wl[89] vdd gnd cell_6t
Xbit_r90_c109 bl[109] br[109] wl[90] vdd gnd cell_6t
Xbit_r91_c109 bl[109] br[109] wl[91] vdd gnd cell_6t
Xbit_r92_c109 bl[109] br[109] wl[92] vdd gnd cell_6t
Xbit_r93_c109 bl[109] br[109] wl[93] vdd gnd cell_6t
Xbit_r94_c109 bl[109] br[109] wl[94] vdd gnd cell_6t
Xbit_r95_c109 bl[109] br[109] wl[95] vdd gnd cell_6t
Xbit_r96_c109 bl[109] br[109] wl[96] vdd gnd cell_6t
Xbit_r97_c109 bl[109] br[109] wl[97] vdd gnd cell_6t
Xbit_r98_c109 bl[109] br[109] wl[98] vdd gnd cell_6t
Xbit_r99_c109 bl[109] br[109] wl[99] vdd gnd cell_6t
Xbit_r100_c109 bl[109] br[109] wl[100] vdd gnd cell_6t
Xbit_r101_c109 bl[109] br[109] wl[101] vdd gnd cell_6t
Xbit_r102_c109 bl[109] br[109] wl[102] vdd gnd cell_6t
Xbit_r103_c109 bl[109] br[109] wl[103] vdd gnd cell_6t
Xbit_r104_c109 bl[109] br[109] wl[104] vdd gnd cell_6t
Xbit_r105_c109 bl[109] br[109] wl[105] vdd gnd cell_6t
Xbit_r106_c109 bl[109] br[109] wl[106] vdd gnd cell_6t
Xbit_r107_c109 bl[109] br[109] wl[107] vdd gnd cell_6t
Xbit_r108_c109 bl[109] br[109] wl[108] vdd gnd cell_6t
Xbit_r109_c109 bl[109] br[109] wl[109] vdd gnd cell_6t
Xbit_r110_c109 bl[109] br[109] wl[110] vdd gnd cell_6t
Xbit_r111_c109 bl[109] br[109] wl[111] vdd gnd cell_6t
Xbit_r112_c109 bl[109] br[109] wl[112] vdd gnd cell_6t
Xbit_r113_c109 bl[109] br[109] wl[113] vdd gnd cell_6t
Xbit_r114_c109 bl[109] br[109] wl[114] vdd gnd cell_6t
Xbit_r115_c109 bl[109] br[109] wl[115] vdd gnd cell_6t
Xbit_r116_c109 bl[109] br[109] wl[116] vdd gnd cell_6t
Xbit_r117_c109 bl[109] br[109] wl[117] vdd gnd cell_6t
Xbit_r118_c109 bl[109] br[109] wl[118] vdd gnd cell_6t
Xbit_r119_c109 bl[109] br[109] wl[119] vdd gnd cell_6t
Xbit_r120_c109 bl[109] br[109] wl[120] vdd gnd cell_6t
Xbit_r121_c109 bl[109] br[109] wl[121] vdd gnd cell_6t
Xbit_r122_c109 bl[109] br[109] wl[122] vdd gnd cell_6t
Xbit_r123_c109 bl[109] br[109] wl[123] vdd gnd cell_6t
Xbit_r124_c109 bl[109] br[109] wl[124] vdd gnd cell_6t
Xbit_r125_c109 bl[109] br[109] wl[125] vdd gnd cell_6t
Xbit_r126_c109 bl[109] br[109] wl[126] vdd gnd cell_6t
Xbit_r127_c109 bl[109] br[109] wl[127] vdd gnd cell_6t
Xbit_r128_c109 bl[109] br[109] wl[128] vdd gnd cell_6t
Xbit_r129_c109 bl[109] br[109] wl[129] vdd gnd cell_6t
Xbit_r130_c109 bl[109] br[109] wl[130] vdd gnd cell_6t
Xbit_r131_c109 bl[109] br[109] wl[131] vdd gnd cell_6t
Xbit_r132_c109 bl[109] br[109] wl[132] vdd gnd cell_6t
Xbit_r133_c109 bl[109] br[109] wl[133] vdd gnd cell_6t
Xbit_r134_c109 bl[109] br[109] wl[134] vdd gnd cell_6t
Xbit_r135_c109 bl[109] br[109] wl[135] vdd gnd cell_6t
Xbit_r136_c109 bl[109] br[109] wl[136] vdd gnd cell_6t
Xbit_r137_c109 bl[109] br[109] wl[137] vdd gnd cell_6t
Xbit_r138_c109 bl[109] br[109] wl[138] vdd gnd cell_6t
Xbit_r139_c109 bl[109] br[109] wl[139] vdd gnd cell_6t
Xbit_r140_c109 bl[109] br[109] wl[140] vdd gnd cell_6t
Xbit_r141_c109 bl[109] br[109] wl[141] vdd gnd cell_6t
Xbit_r142_c109 bl[109] br[109] wl[142] vdd gnd cell_6t
Xbit_r143_c109 bl[109] br[109] wl[143] vdd gnd cell_6t
Xbit_r144_c109 bl[109] br[109] wl[144] vdd gnd cell_6t
Xbit_r145_c109 bl[109] br[109] wl[145] vdd gnd cell_6t
Xbit_r146_c109 bl[109] br[109] wl[146] vdd gnd cell_6t
Xbit_r147_c109 bl[109] br[109] wl[147] vdd gnd cell_6t
Xbit_r148_c109 bl[109] br[109] wl[148] vdd gnd cell_6t
Xbit_r149_c109 bl[109] br[109] wl[149] vdd gnd cell_6t
Xbit_r150_c109 bl[109] br[109] wl[150] vdd gnd cell_6t
Xbit_r151_c109 bl[109] br[109] wl[151] vdd gnd cell_6t
Xbit_r152_c109 bl[109] br[109] wl[152] vdd gnd cell_6t
Xbit_r153_c109 bl[109] br[109] wl[153] vdd gnd cell_6t
Xbit_r154_c109 bl[109] br[109] wl[154] vdd gnd cell_6t
Xbit_r155_c109 bl[109] br[109] wl[155] vdd gnd cell_6t
Xbit_r156_c109 bl[109] br[109] wl[156] vdd gnd cell_6t
Xbit_r157_c109 bl[109] br[109] wl[157] vdd gnd cell_6t
Xbit_r158_c109 bl[109] br[109] wl[158] vdd gnd cell_6t
Xbit_r159_c109 bl[109] br[109] wl[159] vdd gnd cell_6t
Xbit_r160_c109 bl[109] br[109] wl[160] vdd gnd cell_6t
Xbit_r161_c109 bl[109] br[109] wl[161] vdd gnd cell_6t
Xbit_r162_c109 bl[109] br[109] wl[162] vdd gnd cell_6t
Xbit_r163_c109 bl[109] br[109] wl[163] vdd gnd cell_6t
Xbit_r164_c109 bl[109] br[109] wl[164] vdd gnd cell_6t
Xbit_r165_c109 bl[109] br[109] wl[165] vdd gnd cell_6t
Xbit_r166_c109 bl[109] br[109] wl[166] vdd gnd cell_6t
Xbit_r167_c109 bl[109] br[109] wl[167] vdd gnd cell_6t
Xbit_r168_c109 bl[109] br[109] wl[168] vdd gnd cell_6t
Xbit_r169_c109 bl[109] br[109] wl[169] vdd gnd cell_6t
Xbit_r170_c109 bl[109] br[109] wl[170] vdd gnd cell_6t
Xbit_r171_c109 bl[109] br[109] wl[171] vdd gnd cell_6t
Xbit_r172_c109 bl[109] br[109] wl[172] vdd gnd cell_6t
Xbit_r173_c109 bl[109] br[109] wl[173] vdd gnd cell_6t
Xbit_r174_c109 bl[109] br[109] wl[174] vdd gnd cell_6t
Xbit_r175_c109 bl[109] br[109] wl[175] vdd gnd cell_6t
Xbit_r176_c109 bl[109] br[109] wl[176] vdd gnd cell_6t
Xbit_r177_c109 bl[109] br[109] wl[177] vdd gnd cell_6t
Xbit_r178_c109 bl[109] br[109] wl[178] vdd gnd cell_6t
Xbit_r179_c109 bl[109] br[109] wl[179] vdd gnd cell_6t
Xbit_r180_c109 bl[109] br[109] wl[180] vdd gnd cell_6t
Xbit_r181_c109 bl[109] br[109] wl[181] vdd gnd cell_6t
Xbit_r182_c109 bl[109] br[109] wl[182] vdd gnd cell_6t
Xbit_r183_c109 bl[109] br[109] wl[183] vdd gnd cell_6t
Xbit_r184_c109 bl[109] br[109] wl[184] vdd gnd cell_6t
Xbit_r185_c109 bl[109] br[109] wl[185] vdd gnd cell_6t
Xbit_r186_c109 bl[109] br[109] wl[186] vdd gnd cell_6t
Xbit_r187_c109 bl[109] br[109] wl[187] vdd gnd cell_6t
Xbit_r188_c109 bl[109] br[109] wl[188] vdd gnd cell_6t
Xbit_r189_c109 bl[109] br[109] wl[189] vdd gnd cell_6t
Xbit_r190_c109 bl[109] br[109] wl[190] vdd gnd cell_6t
Xbit_r191_c109 bl[109] br[109] wl[191] vdd gnd cell_6t
Xbit_r192_c109 bl[109] br[109] wl[192] vdd gnd cell_6t
Xbit_r193_c109 bl[109] br[109] wl[193] vdd gnd cell_6t
Xbit_r194_c109 bl[109] br[109] wl[194] vdd gnd cell_6t
Xbit_r195_c109 bl[109] br[109] wl[195] vdd gnd cell_6t
Xbit_r196_c109 bl[109] br[109] wl[196] vdd gnd cell_6t
Xbit_r197_c109 bl[109] br[109] wl[197] vdd gnd cell_6t
Xbit_r198_c109 bl[109] br[109] wl[198] vdd gnd cell_6t
Xbit_r199_c109 bl[109] br[109] wl[199] vdd gnd cell_6t
Xbit_r200_c109 bl[109] br[109] wl[200] vdd gnd cell_6t
Xbit_r201_c109 bl[109] br[109] wl[201] vdd gnd cell_6t
Xbit_r202_c109 bl[109] br[109] wl[202] vdd gnd cell_6t
Xbit_r203_c109 bl[109] br[109] wl[203] vdd gnd cell_6t
Xbit_r204_c109 bl[109] br[109] wl[204] vdd gnd cell_6t
Xbit_r205_c109 bl[109] br[109] wl[205] vdd gnd cell_6t
Xbit_r206_c109 bl[109] br[109] wl[206] vdd gnd cell_6t
Xbit_r207_c109 bl[109] br[109] wl[207] vdd gnd cell_6t
Xbit_r208_c109 bl[109] br[109] wl[208] vdd gnd cell_6t
Xbit_r209_c109 bl[109] br[109] wl[209] vdd gnd cell_6t
Xbit_r210_c109 bl[109] br[109] wl[210] vdd gnd cell_6t
Xbit_r211_c109 bl[109] br[109] wl[211] vdd gnd cell_6t
Xbit_r212_c109 bl[109] br[109] wl[212] vdd gnd cell_6t
Xbit_r213_c109 bl[109] br[109] wl[213] vdd gnd cell_6t
Xbit_r214_c109 bl[109] br[109] wl[214] vdd gnd cell_6t
Xbit_r215_c109 bl[109] br[109] wl[215] vdd gnd cell_6t
Xbit_r216_c109 bl[109] br[109] wl[216] vdd gnd cell_6t
Xbit_r217_c109 bl[109] br[109] wl[217] vdd gnd cell_6t
Xbit_r218_c109 bl[109] br[109] wl[218] vdd gnd cell_6t
Xbit_r219_c109 bl[109] br[109] wl[219] vdd gnd cell_6t
Xbit_r220_c109 bl[109] br[109] wl[220] vdd gnd cell_6t
Xbit_r221_c109 bl[109] br[109] wl[221] vdd gnd cell_6t
Xbit_r222_c109 bl[109] br[109] wl[222] vdd gnd cell_6t
Xbit_r223_c109 bl[109] br[109] wl[223] vdd gnd cell_6t
Xbit_r224_c109 bl[109] br[109] wl[224] vdd gnd cell_6t
Xbit_r225_c109 bl[109] br[109] wl[225] vdd gnd cell_6t
Xbit_r226_c109 bl[109] br[109] wl[226] vdd gnd cell_6t
Xbit_r227_c109 bl[109] br[109] wl[227] vdd gnd cell_6t
Xbit_r228_c109 bl[109] br[109] wl[228] vdd gnd cell_6t
Xbit_r229_c109 bl[109] br[109] wl[229] vdd gnd cell_6t
Xbit_r230_c109 bl[109] br[109] wl[230] vdd gnd cell_6t
Xbit_r231_c109 bl[109] br[109] wl[231] vdd gnd cell_6t
Xbit_r232_c109 bl[109] br[109] wl[232] vdd gnd cell_6t
Xbit_r233_c109 bl[109] br[109] wl[233] vdd gnd cell_6t
Xbit_r234_c109 bl[109] br[109] wl[234] vdd gnd cell_6t
Xbit_r235_c109 bl[109] br[109] wl[235] vdd gnd cell_6t
Xbit_r236_c109 bl[109] br[109] wl[236] vdd gnd cell_6t
Xbit_r237_c109 bl[109] br[109] wl[237] vdd gnd cell_6t
Xbit_r238_c109 bl[109] br[109] wl[238] vdd gnd cell_6t
Xbit_r239_c109 bl[109] br[109] wl[239] vdd gnd cell_6t
Xbit_r240_c109 bl[109] br[109] wl[240] vdd gnd cell_6t
Xbit_r241_c109 bl[109] br[109] wl[241] vdd gnd cell_6t
Xbit_r242_c109 bl[109] br[109] wl[242] vdd gnd cell_6t
Xbit_r243_c109 bl[109] br[109] wl[243] vdd gnd cell_6t
Xbit_r244_c109 bl[109] br[109] wl[244] vdd gnd cell_6t
Xbit_r245_c109 bl[109] br[109] wl[245] vdd gnd cell_6t
Xbit_r246_c109 bl[109] br[109] wl[246] vdd gnd cell_6t
Xbit_r247_c109 bl[109] br[109] wl[247] vdd gnd cell_6t
Xbit_r248_c109 bl[109] br[109] wl[248] vdd gnd cell_6t
Xbit_r249_c109 bl[109] br[109] wl[249] vdd gnd cell_6t
Xbit_r250_c109 bl[109] br[109] wl[250] vdd gnd cell_6t
Xbit_r251_c109 bl[109] br[109] wl[251] vdd gnd cell_6t
Xbit_r252_c109 bl[109] br[109] wl[252] vdd gnd cell_6t
Xbit_r253_c109 bl[109] br[109] wl[253] vdd gnd cell_6t
Xbit_r254_c109 bl[109] br[109] wl[254] vdd gnd cell_6t
Xbit_r255_c109 bl[109] br[109] wl[255] vdd gnd cell_6t
Xbit_r256_c109 bl[109] br[109] wl[256] vdd gnd cell_6t
Xbit_r257_c109 bl[109] br[109] wl[257] vdd gnd cell_6t
Xbit_r258_c109 bl[109] br[109] wl[258] vdd gnd cell_6t
Xbit_r259_c109 bl[109] br[109] wl[259] vdd gnd cell_6t
Xbit_r260_c109 bl[109] br[109] wl[260] vdd gnd cell_6t
Xbit_r261_c109 bl[109] br[109] wl[261] vdd gnd cell_6t
Xbit_r262_c109 bl[109] br[109] wl[262] vdd gnd cell_6t
Xbit_r263_c109 bl[109] br[109] wl[263] vdd gnd cell_6t
Xbit_r264_c109 bl[109] br[109] wl[264] vdd gnd cell_6t
Xbit_r265_c109 bl[109] br[109] wl[265] vdd gnd cell_6t
Xbit_r266_c109 bl[109] br[109] wl[266] vdd gnd cell_6t
Xbit_r267_c109 bl[109] br[109] wl[267] vdd gnd cell_6t
Xbit_r268_c109 bl[109] br[109] wl[268] vdd gnd cell_6t
Xbit_r269_c109 bl[109] br[109] wl[269] vdd gnd cell_6t
Xbit_r270_c109 bl[109] br[109] wl[270] vdd gnd cell_6t
Xbit_r271_c109 bl[109] br[109] wl[271] vdd gnd cell_6t
Xbit_r272_c109 bl[109] br[109] wl[272] vdd gnd cell_6t
Xbit_r273_c109 bl[109] br[109] wl[273] vdd gnd cell_6t
Xbit_r274_c109 bl[109] br[109] wl[274] vdd gnd cell_6t
Xbit_r275_c109 bl[109] br[109] wl[275] vdd gnd cell_6t
Xbit_r276_c109 bl[109] br[109] wl[276] vdd gnd cell_6t
Xbit_r277_c109 bl[109] br[109] wl[277] vdd gnd cell_6t
Xbit_r278_c109 bl[109] br[109] wl[278] vdd gnd cell_6t
Xbit_r279_c109 bl[109] br[109] wl[279] vdd gnd cell_6t
Xbit_r280_c109 bl[109] br[109] wl[280] vdd gnd cell_6t
Xbit_r281_c109 bl[109] br[109] wl[281] vdd gnd cell_6t
Xbit_r282_c109 bl[109] br[109] wl[282] vdd gnd cell_6t
Xbit_r283_c109 bl[109] br[109] wl[283] vdd gnd cell_6t
Xbit_r284_c109 bl[109] br[109] wl[284] vdd gnd cell_6t
Xbit_r285_c109 bl[109] br[109] wl[285] vdd gnd cell_6t
Xbit_r286_c109 bl[109] br[109] wl[286] vdd gnd cell_6t
Xbit_r287_c109 bl[109] br[109] wl[287] vdd gnd cell_6t
Xbit_r288_c109 bl[109] br[109] wl[288] vdd gnd cell_6t
Xbit_r289_c109 bl[109] br[109] wl[289] vdd gnd cell_6t
Xbit_r290_c109 bl[109] br[109] wl[290] vdd gnd cell_6t
Xbit_r291_c109 bl[109] br[109] wl[291] vdd gnd cell_6t
Xbit_r292_c109 bl[109] br[109] wl[292] vdd gnd cell_6t
Xbit_r293_c109 bl[109] br[109] wl[293] vdd gnd cell_6t
Xbit_r294_c109 bl[109] br[109] wl[294] vdd gnd cell_6t
Xbit_r295_c109 bl[109] br[109] wl[295] vdd gnd cell_6t
Xbit_r296_c109 bl[109] br[109] wl[296] vdd gnd cell_6t
Xbit_r297_c109 bl[109] br[109] wl[297] vdd gnd cell_6t
Xbit_r298_c109 bl[109] br[109] wl[298] vdd gnd cell_6t
Xbit_r299_c109 bl[109] br[109] wl[299] vdd gnd cell_6t
Xbit_r300_c109 bl[109] br[109] wl[300] vdd gnd cell_6t
Xbit_r301_c109 bl[109] br[109] wl[301] vdd gnd cell_6t
Xbit_r302_c109 bl[109] br[109] wl[302] vdd gnd cell_6t
Xbit_r303_c109 bl[109] br[109] wl[303] vdd gnd cell_6t
Xbit_r304_c109 bl[109] br[109] wl[304] vdd gnd cell_6t
Xbit_r305_c109 bl[109] br[109] wl[305] vdd gnd cell_6t
Xbit_r306_c109 bl[109] br[109] wl[306] vdd gnd cell_6t
Xbit_r307_c109 bl[109] br[109] wl[307] vdd gnd cell_6t
Xbit_r308_c109 bl[109] br[109] wl[308] vdd gnd cell_6t
Xbit_r309_c109 bl[109] br[109] wl[309] vdd gnd cell_6t
Xbit_r310_c109 bl[109] br[109] wl[310] vdd gnd cell_6t
Xbit_r311_c109 bl[109] br[109] wl[311] vdd gnd cell_6t
Xbit_r312_c109 bl[109] br[109] wl[312] vdd gnd cell_6t
Xbit_r313_c109 bl[109] br[109] wl[313] vdd gnd cell_6t
Xbit_r314_c109 bl[109] br[109] wl[314] vdd gnd cell_6t
Xbit_r315_c109 bl[109] br[109] wl[315] vdd gnd cell_6t
Xbit_r316_c109 bl[109] br[109] wl[316] vdd gnd cell_6t
Xbit_r317_c109 bl[109] br[109] wl[317] vdd gnd cell_6t
Xbit_r318_c109 bl[109] br[109] wl[318] vdd gnd cell_6t
Xbit_r319_c109 bl[109] br[109] wl[319] vdd gnd cell_6t
Xbit_r320_c109 bl[109] br[109] wl[320] vdd gnd cell_6t
Xbit_r321_c109 bl[109] br[109] wl[321] vdd gnd cell_6t
Xbit_r322_c109 bl[109] br[109] wl[322] vdd gnd cell_6t
Xbit_r323_c109 bl[109] br[109] wl[323] vdd gnd cell_6t
Xbit_r324_c109 bl[109] br[109] wl[324] vdd gnd cell_6t
Xbit_r325_c109 bl[109] br[109] wl[325] vdd gnd cell_6t
Xbit_r326_c109 bl[109] br[109] wl[326] vdd gnd cell_6t
Xbit_r327_c109 bl[109] br[109] wl[327] vdd gnd cell_6t
Xbit_r328_c109 bl[109] br[109] wl[328] vdd gnd cell_6t
Xbit_r329_c109 bl[109] br[109] wl[329] vdd gnd cell_6t
Xbit_r330_c109 bl[109] br[109] wl[330] vdd gnd cell_6t
Xbit_r331_c109 bl[109] br[109] wl[331] vdd gnd cell_6t
Xbit_r332_c109 bl[109] br[109] wl[332] vdd gnd cell_6t
Xbit_r333_c109 bl[109] br[109] wl[333] vdd gnd cell_6t
Xbit_r334_c109 bl[109] br[109] wl[334] vdd gnd cell_6t
Xbit_r335_c109 bl[109] br[109] wl[335] vdd gnd cell_6t
Xbit_r336_c109 bl[109] br[109] wl[336] vdd gnd cell_6t
Xbit_r337_c109 bl[109] br[109] wl[337] vdd gnd cell_6t
Xbit_r338_c109 bl[109] br[109] wl[338] vdd gnd cell_6t
Xbit_r339_c109 bl[109] br[109] wl[339] vdd gnd cell_6t
Xbit_r340_c109 bl[109] br[109] wl[340] vdd gnd cell_6t
Xbit_r341_c109 bl[109] br[109] wl[341] vdd gnd cell_6t
Xbit_r342_c109 bl[109] br[109] wl[342] vdd gnd cell_6t
Xbit_r343_c109 bl[109] br[109] wl[343] vdd gnd cell_6t
Xbit_r344_c109 bl[109] br[109] wl[344] vdd gnd cell_6t
Xbit_r345_c109 bl[109] br[109] wl[345] vdd gnd cell_6t
Xbit_r346_c109 bl[109] br[109] wl[346] vdd gnd cell_6t
Xbit_r347_c109 bl[109] br[109] wl[347] vdd gnd cell_6t
Xbit_r348_c109 bl[109] br[109] wl[348] vdd gnd cell_6t
Xbit_r349_c109 bl[109] br[109] wl[349] vdd gnd cell_6t
Xbit_r350_c109 bl[109] br[109] wl[350] vdd gnd cell_6t
Xbit_r351_c109 bl[109] br[109] wl[351] vdd gnd cell_6t
Xbit_r352_c109 bl[109] br[109] wl[352] vdd gnd cell_6t
Xbit_r353_c109 bl[109] br[109] wl[353] vdd gnd cell_6t
Xbit_r354_c109 bl[109] br[109] wl[354] vdd gnd cell_6t
Xbit_r355_c109 bl[109] br[109] wl[355] vdd gnd cell_6t
Xbit_r356_c109 bl[109] br[109] wl[356] vdd gnd cell_6t
Xbit_r357_c109 bl[109] br[109] wl[357] vdd gnd cell_6t
Xbit_r358_c109 bl[109] br[109] wl[358] vdd gnd cell_6t
Xbit_r359_c109 bl[109] br[109] wl[359] vdd gnd cell_6t
Xbit_r360_c109 bl[109] br[109] wl[360] vdd gnd cell_6t
Xbit_r361_c109 bl[109] br[109] wl[361] vdd gnd cell_6t
Xbit_r362_c109 bl[109] br[109] wl[362] vdd gnd cell_6t
Xbit_r363_c109 bl[109] br[109] wl[363] vdd gnd cell_6t
Xbit_r364_c109 bl[109] br[109] wl[364] vdd gnd cell_6t
Xbit_r365_c109 bl[109] br[109] wl[365] vdd gnd cell_6t
Xbit_r366_c109 bl[109] br[109] wl[366] vdd gnd cell_6t
Xbit_r367_c109 bl[109] br[109] wl[367] vdd gnd cell_6t
Xbit_r368_c109 bl[109] br[109] wl[368] vdd gnd cell_6t
Xbit_r369_c109 bl[109] br[109] wl[369] vdd gnd cell_6t
Xbit_r370_c109 bl[109] br[109] wl[370] vdd gnd cell_6t
Xbit_r371_c109 bl[109] br[109] wl[371] vdd gnd cell_6t
Xbit_r372_c109 bl[109] br[109] wl[372] vdd gnd cell_6t
Xbit_r373_c109 bl[109] br[109] wl[373] vdd gnd cell_6t
Xbit_r374_c109 bl[109] br[109] wl[374] vdd gnd cell_6t
Xbit_r375_c109 bl[109] br[109] wl[375] vdd gnd cell_6t
Xbit_r376_c109 bl[109] br[109] wl[376] vdd gnd cell_6t
Xbit_r377_c109 bl[109] br[109] wl[377] vdd gnd cell_6t
Xbit_r378_c109 bl[109] br[109] wl[378] vdd gnd cell_6t
Xbit_r379_c109 bl[109] br[109] wl[379] vdd gnd cell_6t
Xbit_r380_c109 bl[109] br[109] wl[380] vdd gnd cell_6t
Xbit_r381_c109 bl[109] br[109] wl[381] vdd gnd cell_6t
Xbit_r382_c109 bl[109] br[109] wl[382] vdd gnd cell_6t
Xbit_r383_c109 bl[109] br[109] wl[383] vdd gnd cell_6t
Xbit_r384_c109 bl[109] br[109] wl[384] vdd gnd cell_6t
Xbit_r385_c109 bl[109] br[109] wl[385] vdd gnd cell_6t
Xbit_r386_c109 bl[109] br[109] wl[386] vdd gnd cell_6t
Xbit_r387_c109 bl[109] br[109] wl[387] vdd gnd cell_6t
Xbit_r388_c109 bl[109] br[109] wl[388] vdd gnd cell_6t
Xbit_r389_c109 bl[109] br[109] wl[389] vdd gnd cell_6t
Xbit_r390_c109 bl[109] br[109] wl[390] vdd gnd cell_6t
Xbit_r391_c109 bl[109] br[109] wl[391] vdd gnd cell_6t
Xbit_r392_c109 bl[109] br[109] wl[392] vdd gnd cell_6t
Xbit_r393_c109 bl[109] br[109] wl[393] vdd gnd cell_6t
Xbit_r394_c109 bl[109] br[109] wl[394] vdd gnd cell_6t
Xbit_r395_c109 bl[109] br[109] wl[395] vdd gnd cell_6t
Xbit_r396_c109 bl[109] br[109] wl[396] vdd gnd cell_6t
Xbit_r397_c109 bl[109] br[109] wl[397] vdd gnd cell_6t
Xbit_r398_c109 bl[109] br[109] wl[398] vdd gnd cell_6t
Xbit_r399_c109 bl[109] br[109] wl[399] vdd gnd cell_6t
Xbit_r400_c109 bl[109] br[109] wl[400] vdd gnd cell_6t
Xbit_r401_c109 bl[109] br[109] wl[401] vdd gnd cell_6t
Xbit_r402_c109 bl[109] br[109] wl[402] vdd gnd cell_6t
Xbit_r403_c109 bl[109] br[109] wl[403] vdd gnd cell_6t
Xbit_r404_c109 bl[109] br[109] wl[404] vdd gnd cell_6t
Xbit_r405_c109 bl[109] br[109] wl[405] vdd gnd cell_6t
Xbit_r406_c109 bl[109] br[109] wl[406] vdd gnd cell_6t
Xbit_r407_c109 bl[109] br[109] wl[407] vdd gnd cell_6t
Xbit_r408_c109 bl[109] br[109] wl[408] vdd gnd cell_6t
Xbit_r409_c109 bl[109] br[109] wl[409] vdd gnd cell_6t
Xbit_r410_c109 bl[109] br[109] wl[410] vdd gnd cell_6t
Xbit_r411_c109 bl[109] br[109] wl[411] vdd gnd cell_6t
Xbit_r412_c109 bl[109] br[109] wl[412] vdd gnd cell_6t
Xbit_r413_c109 bl[109] br[109] wl[413] vdd gnd cell_6t
Xbit_r414_c109 bl[109] br[109] wl[414] vdd gnd cell_6t
Xbit_r415_c109 bl[109] br[109] wl[415] vdd gnd cell_6t
Xbit_r416_c109 bl[109] br[109] wl[416] vdd gnd cell_6t
Xbit_r417_c109 bl[109] br[109] wl[417] vdd gnd cell_6t
Xbit_r418_c109 bl[109] br[109] wl[418] vdd gnd cell_6t
Xbit_r419_c109 bl[109] br[109] wl[419] vdd gnd cell_6t
Xbit_r420_c109 bl[109] br[109] wl[420] vdd gnd cell_6t
Xbit_r421_c109 bl[109] br[109] wl[421] vdd gnd cell_6t
Xbit_r422_c109 bl[109] br[109] wl[422] vdd gnd cell_6t
Xbit_r423_c109 bl[109] br[109] wl[423] vdd gnd cell_6t
Xbit_r424_c109 bl[109] br[109] wl[424] vdd gnd cell_6t
Xbit_r425_c109 bl[109] br[109] wl[425] vdd gnd cell_6t
Xbit_r426_c109 bl[109] br[109] wl[426] vdd gnd cell_6t
Xbit_r427_c109 bl[109] br[109] wl[427] vdd gnd cell_6t
Xbit_r428_c109 bl[109] br[109] wl[428] vdd gnd cell_6t
Xbit_r429_c109 bl[109] br[109] wl[429] vdd gnd cell_6t
Xbit_r430_c109 bl[109] br[109] wl[430] vdd gnd cell_6t
Xbit_r431_c109 bl[109] br[109] wl[431] vdd gnd cell_6t
Xbit_r432_c109 bl[109] br[109] wl[432] vdd gnd cell_6t
Xbit_r433_c109 bl[109] br[109] wl[433] vdd gnd cell_6t
Xbit_r434_c109 bl[109] br[109] wl[434] vdd gnd cell_6t
Xbit_r435_c109 bl[109] br[109] wl[435] vdd gnd cell_6t
Xbit_r436_c109 bl[109] br[109] wl[436] vdd gnd cell_6t
Xbit_r437_c109 bl[109] br[109] wl[437] vdd gnd cell_6t
Xbit_r438_c109 bl[109] br[109] wl[438] vdd gnd cell_6t
Xbit_r439_c109 bl[109] br[109] wl[439] vdd gnd cell_6t
Xbit_r440_c109 bl[109] br[109] wl[440] vdd gnd cell_6t
Xbit_r441_c109 bl[109] br[109] wl[441] vdd gnd cell_6t
Xbit_r442_c109 bl[109] br[109] wl[442] vdd gnd cell_6t
Xbit_r443_c109 bl[109] br[109] wl[443] vdd gnd cell_6t
Xbit_r444_c109 bl[109] br[109] wl[444] vdd gnd cell_6t
Xbit_r445_c109 bl[109] br[109] wl[445] vdd gnd cell_6t
Xbit_r446_c109 bl[109] br[109] wl[446] vdd gnd cell_6t
Xbit_r447_c109 bl[109] br[109] wl[447] vdd gnd cell_6t
Xbit_r448_c109 bl[109] br[109] wl[448] vdd gnd cell_6t
Xbit_r449_c109 bl[109] br[109] wl[449] vdd gnd cell_6t
Xbit_r450_c109 bl[109] br[109] wl[450] vdd gnd cell_6t
Xbit_r451_c109 bl[109] br[109] wl[451] vdd gnd cell_6t
Xbit_r452_c109 bl[109] br[109] wl[452] vdd gnd cell_6t
Xbit_r453_c109 bl[109] br[109] wl[453] vdd gnd cell_6t
Xbit_r454_c109 bl[109] br[109] wl[454] vdd gnd cell_6t
Xbit_r455_c109 bl[109] br[109] wl[455] vdd gnd cell_6t
Xbit_r456_c109 bl[109] br[109] wl[456] vdd gnd cell_6t
Xbit_r457_c109 bl[109] br[109] wl[457] vdd gnd cell_6t
Xbit_r458_c109 bl[109] br[109] wl[458] vdd gnd cell_6t
Xbit_r459_c109 bl[109] br[109] wl[459] vdd gnd cell_6t
Xbit_r460_c109 bl[109] br[109] wl[460] vdd gnd cell_6t
Xbit_r461_c109 bl[109] br[109] wl[461] vdd gnd cell_6t
Xbit_r462_c109 bl[109] br[109] wl[462] vdd gnd cell_6t
Xbit_r463_c109 bl[109] br[109] wl[463] vdd gnd cell_6t
Xbit_r464_c109 bl[109] br[109] wl[464] vdd gnd cell_6t
Xbit_r465_c109 bl[109] br[109] wl[465] vdd gnd cell_6t
Xbit_r466_c109 bl[109] br[109] wl[466] vdd gnd cell_6t
Xbit_r467_c109 bl[109] br[109] wl[467] vdd gnd cell_6t
Xbit_r468_c109 bl[109] br[109] wl[468] vdd gnd cell_6t
Xbit_r469_c109 bl[109] br[109] wl[469] vdd gnd cell_6t
Xbit_r470_c109 bl[109] br[109] wl[470] vdd gnd cell_6t
Xbit_r471_c109 bl[109] br[109] wl[471] vdd gnd cell_6t
Xbit_r472_c109 bl[109] br[109] wl[472] vdd gnd cell_6t
Xbit_r473_c109 bl[109] br[109] wl[473] vdd gnd cell_6t
Xbit_r474_c109 bl[109] br[109] wl[474] vdd gnd cell_6t
Xbit_r475_c109 bl[109] br[109] wl[475] vdd gnd cell_6t
Xbit_r476_c109 bl[109] br[109] wl[476] vdd gnd cell_6t
Xbit_r477_c109 bl[109] br[109] wl[477] vdd gnd cell_6t
Xbit_r478_c109 bl[109] br[109] wl[478] vdd gnd cell_6t
Xbit_r479_c109 bl[109] br[109] wl[479] vdd gnd cell_6t
Xbit_r480_c109 bl[109] br[109] wl[480] vdd gnd cell_6t
Xbit_r481_c109 bl[109] br[109] wl[481] vdd gnd cell_6t
Xbit_r482_c109 bl[109] br[109] wl[482] vdd gnd cell_6t
Xbit_r483_c109 bl[109] br[109] wl[483] vdd gnd cell_6t
Xbit_r484_c109 bl[109] br[109] wl[484] vdd gnd cell_6t
Xbit_r485_c109 bl[109] br[109] wl[485] vdd gnd cell_6t
Xbit_r486_c109 bl[109] br[109] wl[486] vdd gnd cell_6t
Xbit_r487_c109 bl[109] br[109] wl[487] vdd gnd cell_6t
Xbit_r488_c109 bl[109] br[109] wl[488] vdd gnd cell_6t
Xbit_r489_c109 bl[109] br[109] wl[489] vdd gnd cell_6t
Xbit_r490_c109 bl[109] br[109] wl[490] vdd gnd cell_6t
Xbit_r491_c109 bl[109] br[109] wl[491] vdd gnd cell_6t
Xbit_r492_c109 bl[109] br[109] wl[492] vdd gnd cell_6t
Xbit_r493_c109 bl[109] br[109] wl[493] vdd gnd cell_6t
Xbit_r494_c109 bl[109] br[109] wl[494] vdd gnd cell_6t
Xbit_r495_c109 bl[109] br[109] wl[495] vdd gnd cell_6t
Xbit_r496_c109 bl[109] br[109] wl[496] vdd gnd cell_6t
Xbit_r497_c109 bl[109] br[109] wl[497] vdd gnd cell_6t
Xbit_r498_c109 bl[109] br[109] wl[498] vdd gnd cell_6t
Xbit_r499_c109 bl[109] br[109] wl[499] vdd gnd cell_6t
Xbit_r500_c109 bl[109] br[109] wl[500] vdd gnd cell_6t
Xbit_r501_c109 bl[109] br[109] wl[501] vdd gnd cell_6t
Xbit_r502_c109 bl[109] br[109] wl[502] vdd gnd cell_6t
Xbit_r503_c109 bl[109] br[109] wl[503] vdd gnd cell_6t
Xbit_r504_c109 bl[109] br[109] wl[504] vdd gnd cell_6t
Xbit_r505_c109 bl[109] br[109] wl[505] vdd gnd cell_6t
Xbit_r506_c109 bl[109] br[109] wl[506] vdd gnd cell_6t
Xbit_r507_c109 bl[109] br[109] wl[507] vdd gnd cell_6t
Xbit_r508_c109 bl[109] br[109] wl[508] vdd gnd cell_6t
Xbit_r509_c109 bl[109] br[109] wl[509] vdd gnd cell_6t
Xbit_r510_c109 bl[109] br[109] wl[510] vdd gnd cell_6t
Xbit_r511_c109 bl[109] br[109] wl[511] vdd gnd cell_6t
Xbit_r0_c110 bl[110] br[110] wl[0] vdd gnd cell_6t
Xbit_r1_c110 bl[110] br[110] wl[1] vdd gnd cell_6t
Xbit_r2_c110 bl[110] br[110] wl[2] vdd gnd cell_6t
Xbit_r3_c110 bl[110] br[110] wl[3] vdd gnd cell_6t
Xbit_r4_c110 bl[110] br[110] wl[4] vdd gnd cell_6t
Xbit_r5_c110 bl[110] br[110] wl[5] vdd gnd cell_6t
Xbit_r6_c110 bl[110] br[110] wl[6] vdd gnd cell_6t
Xbit_r7_c110 bl[110] br[110] wl[7] vdd gnd cell_6t
Xbit_r8_c110 bl[110] br[110] wl[8] vdd gnd cell_6t
Xbit_r9_c110 bl[110] br[110] wl[9] vdd gnd cell_6t
Xbit_r10_c110 bl[110] br[110] wl[10] vdd gnd cell_6t
Xbit_r11_c110 bl[110] br[110] wl[11] vdd gnd cell_6t
Xbit_r12_c110 bl[110] br[110] wl[12] vdd gnd cell_6t
Xbit_r13_c110 bl[110] br[110] wl[13] vdd gnd cell_6t
Xbit_r14_c110 bl[110] br[110] wl[14] vdd gnd cell_6t
Xbit_r15_c110 bl[110] br[110] wl[15] vdd gnd cell_6t
Xbit_r16_c110 bl[110] br[110] wl[16] vdd gnd cell_6t
Xbit_r17_c110 bl[110] br[110] wl[17] vdd gnd cell_6t
Xbit_r18_c110 bl[110] br[110] wl[18] vdd gnd cell_6t
Xbit_r19_c110 bl[110] br[110] wl[19] vdd gnd cell_6t
Xbit_r20_c110 bl[110] br[110] wl[20] vdd gnd cell_6t
Xbit_r21_c110 bl[110] br[110] wl[21] vdd gnd cell_6t
Xbit_r22_c110 bl[110] br[110] wl[22] vdd gnd cell_6t
Xbit_r23_c110 bl[110] br[110] wl[23] vdd gnd cell_6t
Xbit_r24_c110 bl[110] br[110] wl[24] vdd gnd cell_6t
Xbit_r25_c110 bl[110] br[110] wl[25] vdd gnd cell_6t
Xbit_r26_c110 bl[110] br[110] wl[26] vdd gnd cell_6t
Xbit_r27_c110 bl[110] br[110] wl[27] vdd gnd cell_6t
Xbit_r28_c110 bl[110] br[110] wl[28] vdd gnd cell_6t
Xbit_r29_c110 bl[110] br[110] wl[29] vdd gnd cell_6t
Xbit_r30_c110 bl[110] br[110] wl[30] vdd gnd cell_6t
Xbit_r31_c110 bl[110] br[110] wl[31] vdd gnd cell_6t
Xbit_r32_c110 bl[110] br[110] wl[32] vdd gnd cell_6t
Xbit_r33_c110 bl[110] br[110] wl[33] vdd gnd cell_6t
Xbit_r34_c110 bl[110] br[110] wl[34] vdd gnd cell_6t
Xbit_r35_c110 bl[110] br[110] wl[35] vdd gnd cell_6t
Xbit_r36_c110 bl[110] br[110] wl[36] vdd gnd cell_6t
Xbit_r37_c110 bl[110] br[110] wl[37] vdd gnd cell_6t
Xbit_r38_c110 bl[110] br[110] wl[38] vdd gnd cell_6t
Xbit_r39_c110 bl[110] br[110] wl[39] vdd gnd cell_6t
Xbit_r40_c110 bl[110] br[110] wl[40] vdd gnd cell_6t
Xbit_r41_c110 bl[110] br[110] wl[41] vdd gnd cell_6t
Xbit_r42_c110 bl[110] br[110] wl[42] vdd gnd cell_6t
Xbit_r43_c110 bl[110] br[110] wl[43] vdd gnd cell_6t
Xbit_r44_c110 bl[110] br[110] wl[44] vdd gnd cell_6t
Xbit_r45_c110 bl[110] br[110] wl[45] vdd gnd cell_6t
Xbit_r46_c110 bl[110] br[110] wl[46] vdd gnd cell_6t
Xbit_r47_c110 bl[110] br[110] wl[47] vdd gnd cell_6t
Xbit_r48_c110 bl[110] br[110] wl[48] vdd gnd cell_6t
Xbit_r49_c110 bl[110] br[110] wl[49] vdd gnd cell_6t
Xbit_r50_c110 bl[110] br[110] wl[50] vdd gnd cell_6t
Xbit_r51_c110 bl[110] br[110] wl[51] vdd gnd cell_6t
Xbit_r52_c110 bl[110] br[110] wl[52] vdd gnd cell_6t
Xbit_r53_c110 bl[110] br[110] wl[53] vdd gnd cell_6t
Xbit_r54_c110 bl[110] br[110] wl[54] vdd gnd cell_6t
Xbit_r55_c110 bl[110] br[110] wl[55] vdd gnd cell_6t
Xbit_r56_c110 bl[110] br[110] wl[56] vdd gnd cell_6t
Xbit_r57_c110 bl[110] br[110] wl[57] vdd gnd cell_6t
Xbit_r58_c110 bl[110] br[110] wl[58] vdd gnd cell_6t
Xbit_r59_c110 bl[110] br[110] wl[59] vdd gnd cell_6t
Xbit_r60_c110 bl[110] br[110] wl[60] vdd gnd cell_6t
Xbit_r61_c110 bl[110] br[110] wl[61] vdd gnd cell_6t
Xbit_r62_c110 bl[110] br[110] wl[62] vdd gnd cell_6t
Xbit_r63_c110 bl[110] br[110] wl[63] vdd gnd cell_6t
Xbit_r64_c110 bl[110] br[110] wl[64] vdd gnd cell_6t
Xbit_r65_c110 bl[110] br[110] wl[65] vdd gnd cell_6t
Xbit_r66_c110 bl[110] br[110] wl[66] vdd gnd cell_6t
Xbit_r67_c110 bl[110] br[110] wl[67] vdd gnd cell_6t
Xbit_r68_c110 bl[110] br[110] wl[68] vdd gnd cell_6t
Xbit_r69_c110 bl[110] br[110] wl[69] vdd gnd cell_6t
Xbit_r70_c110 bl[110] br[110] wl[70] vdd gnd cell_6t
Xbit_r71_c110 bl[110] br[110] wl[71] vdd gnd cell_6t
Xbit_r72_c110 bl[110] br[110] wl[72] vdd gnd cell_6t
Xbit_r73_c110 bl[110] br[110] wl[73] vdd gnd cell_6t
Xbit_r74_c110 bl[110] br[110] wl[74] vdd gnd cell_6t
Xbit_r75_c110 bl[110] br[110] wl[75] vdd gnd cell_6t
Xbit_r76_c110 bl[110] br[110] wl[76] vdd gnd cell_6t
Xbit_r77_c110 bl[110] br[110] wl[77] vdd gnd cell_6t
Xbit_r78_c110 bl[110] br[110] wl[78] vdd gnd cell_6t
Xbit_r79_c110 bl[110] br[110] wl[79] vdd gnd cell_6t
Xbit_r80_c110 bl[110] br[110] wl[80] vdd gnd cell_6t
Xbit_r81_c110 bl[110] br[110] wl[81] vdd gnd cell_6t
Xbit_r82_c110 bl[110] br[110] wl[82] vdd gnd cell_6t
Xbit_r83_c110 bl[110] br[110] wl[83] vdd gnd cell_6t
Xbit_r84_c110 bl[110] br[110] wl[84] vdd gnd cell_6t
Xbit_r85_c110 bl[110] br[110] wl[85] vdd gnd cell_6t
Xbit_r86_c110 bl[110] br[110] wl[86] vdd gnd cell_6t
Xbit_r87_c110 bl[110] br[110] wl[87] vdd gnd cell_6t
Xbit_r88_c110 bl[110] br[110] wl[88] vdd gnd cell_6t
Xbit_r89_c110 bl[110] br[110] wl[89] vdd gnd cell_6t
Xbit_r90_c110 bl[110] br[110] wl[90] vdd gnd cell_6t
Xbit_r91_c110 bl[110] br[110] wl[91] vdd gnd cell_6t
Xbit_r92_c110 bl[110] br[110] wl[92] vdd gnd cell_6t
Xbit_r93_c110 bl[110] br[110] wl[93] vdd gnd cell_6t
Xbit_r94_c110 bl[110] br[110] wl[94] vdd gnd cell_6t
Xbit_r95_c110 bl[110] br[110] wl[95] vdd gnd cell_6t
Xbit_r96_c110 bl[110] br[110] wl[96] vdd gnd cell_6t
Xbit_r97_c110 bl[110] br[110] wl[97] vdd gnd cell_6t
Xbit_r98_c110 bl[110] br[110] wl[98] vdd gnd cell_6t
Xbit_r99_c110 bl[110] br[110] wl[99] vdd gnd cell_6t
Xbit_r100_c110 bl[110] br[110] wl[100] vdd gnd cell_6t
Xbit_r101_c110 bl[110] br[110] wl[101] vdd gnd cell_6t
Xbit_r102_c110 bl[110] br[110] wl[102] vdd gnd cell_6t
Xbit_r103_c110 bl[110] br[110] wl[103] vdd gnd cell_6t
Xbit_r104_c110 bl[110] br[110] wl[104] vdd gnd cell_6t
Xbit_r105_c110 bl[110] br[110] wl[105] vdd gnd cell_6t
Xbit_r106_c110 bl[110] br[110] wl[106] vdd gnd cell_6t
Xbit_r107_c110 bl[110] br[110] wl[107] vdd gnd cell_6t
Xbit_r108_c110 bl[110] br[110] wl[108] vdd gnd cell_6t
Xbit_r109_c110 bl[110] br[110] wl[109] vdd gnd cell_6t
Xbit_r110_c110 bl[110] br[110] wl[110] vdd gnd cell_6t
Xbit_r111_c110 bl[110] br[110] wl[111] vdd gnd cell_6t
Xbit_r112_c110 bl[110] br[110] wl[112] vdd gnd cell_6t
Xbit_r113_c110 bl[110] br[110] wl[113] vdd gnd cell_6t
Xbit_r114_c110 bl[110] br[110] wl[114] vdd gnd cell_6t
Xbit_r115_c110 bl[110] br[110] wl[115] vdd gnd cell_6t
Xbit_r116_c110 bl[110] br[110] wl[116] vdd gnd cell_6t
Xbit_r117_c110 bl[110] br[110] wl[117] vdd gnd cell_6t
Xbit_r118_c110 bl[110] br[110] wl[118] vdd gnd cell_6t
Xbit_r119_c110 bl[110] br[110] wl[119] vdd gnd cell_6t
Xbit_r120_c110 bl[110] br[110] wl[120] vdd gnd cell_6t
Xbit_r121_c110 bl[110] br[110] wl[121] vdd gnd cell_6t
Xbit_r122_c110 bl[110] br[110] wl[122] vdd gnd cell_6t
Xbit_r123_c110 bl[110] br[110] wl[123] vdd gnd cell_6t
Xbit_r124_c110 bl[110] br[110] wl[124] vdd gnd cell_6t
Xbit_r125_c110 bl[110] br[110] wl[125] vdd gnd cell_6t
Xbit_r126_c110 bl[110] br[110] wl[126] vdd gnd cell_6t
Xbit_r127_c110 bl[110] br[110] wl[127] vdd gnd cell_6t
Xbit_r128_c110 bl[110] br[110] wl[128] vdd gnd cell_6t
Xbit_r129_c110 bl[110] br[110] wl[129] vdd gnd cell_6t
Xbit_r130_c110 bl[110] br[110] wl[130] vdd gnd cell_6t
Xbit_r131_c110 bl[110] br[110] wl[131] vdd gnd cell_6t
Xbit_r132_c110 bl[110] br[110] wl[132] vdd gnd cell_6t
Xbit_r133_c110 bl[110] br[110] wl[133] vdd gnd cell_6t
Xbit_r134_c110 bl[110] br[110] wl[134] vdd gnd cell_6t
Xbit_r135_c110 bl[110] br[110] wl[135] vdd gnd cell_6t
Xbit_r136_c110 bl[110] br[110] wl[136] vdd gnd cell_6t
Xbit_r137_c110 bl[110] br[110] wl[137] vdd gnd cell_6t
Xbit_r138_c110 bl[110] br[110] wl[138] vdd gnd cell_6t
Xbit_r139_c110 bl[110] br[110] wl[139] vdd gnd cell_6t
Xbit_r140_c110 bl[110] br[110] wl[140] vdd gnd cell_6t
Xbit_r141_c110 bl[110] br[110] wl[141] vdd gnd cell_6t
Xbit_r142_c110 bl[110] br[110] wl[142] vdd gnd cell_6t
Xbit_r143_c110 bl[110] br[110] wl[143] vdd gnd cell_6t
Xbit_r144_c110 bl[110] br[110] wl[144] vdd gnd cell_6t
Xbit_r145_c110 bl[110] br[110] wl[145] vdd gnd cell_6t
Xbit_r146_c110 bl[110] br[110] wl[146] vdd gnd cell_6t
Xbit_r147_c110 bl[110] br[110] wl[147] vdd gnd cell_6t
Xbit_r148_c110 bl[110] br[110] wl[148] vdd gnd cell_6t
Xbit_r149_c110 bl[110] br[110] wl[149] vdd gnd cell_6t
Xbit_r150_c110 bl[110] br[110] wl[150] vdd gnd cell_6t
Xbit_r151_c110 bl[110] br[110] wl[151] vdd gnd cell_6t
Xbit_r152_c110 bl[110] br[110] wl[152] vdd gnd cell_6t
Xbit_r153_c110 bl[110] br[110] wl[153] vdd gnd cell_6t
Xbit_r154_c110 bl[110] br[110] wl[154] vdd gnd cell_6t
Xbit_r155_c110 bl[110] br[110] wl[155] vdd gnd cell_6t
Xbit_r156_c110 bl[110] br[110] wl[156] vdd gnd cell_6t
Xbit_r157_c110 bl[110] br[110] wl[157] vdd gnd cell_6t
Xbit_r158_c110 bl[110] br[110] wl[158] vdd gnd cell_6t
Xbit_r159_c110 bl[110] br[110] wl[159] vdd gnd cell_6t
Xbit_r160_c110 bl[110] br[110] wl[160] vdd gnd cell_6t
Xbit_r161_c110 bl[110] br[110] wl[161] vdd gnd cell_6t
Xbit_r162_c110 bl[110] br[110] wl[162] vdd gnd cell_6t
Xbit_r163_c110 bl[110] br[110] wl[163] vdd gnd cell_6t
Xbit_r164_c110 bl[110] br[110] wl[164] vdd gnd cell_6t
Xbit_r165_c110 bl[110] br[110] wl[165] vdd gnd cell_6t
Xbit_r166_c110 bl[110] br[110] wl[166] vdd gnd cell_6t
Xbit_r167_c110 bl[110] br[110] wl[167] vdd gnd cell_6t
Xbit_r168_c110 bl[110] br[110] wl[168] vdd gnd cell_6t
Xbit_r169_c110 bl[110] br[110] wl[169] vdd gnd cell_6t
Xbit_r170_c110 bl[110] br[110] wl[170] vdd gnd cell_6t
Xbit_r171_c110 bl[110] br[110] wl[171] vdd gnd cell_6t
Xbit_r172_c110 bl[110] br[110] wl[172] vdd gnd cell_6t
Xbit_r173_c110 bl[110] br[110] wl[173] vdd gnd cell_6t
Xbit_r174_c110 bl[110] br[110] wl[174] vdd gnd cell_6t
Xbit_r175_c110 bl[110] br[110] wl[175] vdd gnd cell_6t
Xbit_r176_c110 bl[110] br[110] wl[176] vdd gnd cell_6t
Xbit_r177_c110 bl[110] br[110] wl[177] vdd gnd cell_6t
Xbit_r178_c110 bl[110] br[110] wl[178] vdd gnd cell_6t
Xbit_r179_c110 bl[110] br[110] wl[179] vdd gnd cell_6t
Xbit_r180_c110 bl[110] br[110] wl[180] vdd gnd cell_6t
Xbit_r181_c110 bl[110] br[110] wl[181] vdd gnd cell_6t
Xbit_r182_c110 bl[110] br[110] wl[182] vdd gnd cell_6t
Xbit_r183_c110 bl[110] br[110] wl[183] vdd gnd cell_6t
Xbit_r184_c110 bl[110] br[110] wl[184] vdd gnd cell_6t
Xbit_r185_c110 bl[110] br[110] wl[185] vdd gnd cell_6t
Xbit_r186_c110 bl[110] br[110] wl[186] vdd gnd cell_6t
Xbit_r187_c110 bl[110] br[110] wl[187] vdd gnd cell_6t
Xbit_r188_c110 bl[110] br[110] wl[188] vdd gnd cell_6t
Xbit_r189_c110 bl[110] br[110] wl[189] vdd gnd cell_6t
Xbit_r190_c110 bl[110] br[110] wl[190] vdd gnd cell_6t
Xbit_r191_c110 bl[110] br[110] wl[191] vdd gnd cell_6t
Xbit_r192_c110 bl[110] br[110] wl[192] vdd gnd cell_6t
Xbit_r193_c110 bl[110] br[110] wl[193] vdd gnd cell_6t
Xbit_r194_c110 bl[110] br[110] wl[194] vdd gnd cell_6t
Xbit_r195_c110 bl[110] br[110] wl[195] vdd gnd cell_6t
Xbit_r196_c110 bl[110] br[110] wl[196] vdd gnd cell_6t
Xbit_r197_c110 bl[110] br[110] wl[197] vdd gnd cell_6t
Xbit_r198_c110 bl[110] br[110] wl[198] vdd gnd cell_6t
Xbit_r199_c110 bl[110] br[110] wl[199] vdd gnd cell_6t
Xbit_r200_c110 bl[110] br[110] wl[200] vdd gnd cell_6t
Xbit_r201_c110 bl[110] br[110] wl[201] vdd gnd cell_6t
Xbit_r202_c110 bl[110] br[110] wl[202] vdd gnd cell_6t
Xbit_r203_c110 bl[110] br[110] wl[203] vdd gnd cell_6t
Xbit_r204_c110 bl[110] br[110] wl[204] vdd gnd cell_6t
Xbit_r205_c110 bl[110] br[110] wl[205] vdd gnd cell_6t
Xbit_r206_c110 bl[110] br[110] wl[206] vdd gnd cell_6t
Xbit_r207_c110 bl[110] br[110] wl[207] vdd gnd cell_6t
Xbit_r208_c110 bl[110] br[110] wl[208] vdd gnd cell_6t
Xbit_r209_c110 bl[110] br[110] wl[209] vdd gnd cell_6t
Xbit_r210_c110 bl[110] br[110] wl[210] vdd gnd cell_6t
Xbit_r211_c110 bl[110] br[110] wl[211] vdd gnd cell_6t
Xbit_r212_c110 bl[110] br[110] wl[212] vdd gnd cell_6t
Xbit_r213_c110 bl[110] br[110] wl[213] vdd gnd cell_6t
Xbit_r214_c110 bl[110] br[110] wl[214] vdd gnd cell_6t
Xbit_r215_c110 bl[110] br[110] wl[215] vdd gnd cell_6t
Xbit_r216_c110 bl[110] br[110] wl[216] vdd gnd cell_6t
Xbit_r217_c110 bl[110] br[110] wl[217] vdd gnd cell_6t
Xbit_r218_c110 bl[110] br[110] wl[218] vdd gnd cell_6t
Xbit_r219_c110 bl[110] br[110] wl[219] vdd gnd cell_6t
Xbit_r220_c110 bl[110] br[110] wl[220] vdd gnd cell_6t
Xbit_r221_c110 bl[110] br[110] wl[221] vdd gnd cell_6t
Xbit_r222_c110 bl[110] br[110] wl[222] vdd gnd cell_6t
Xbit_r223_c110 bl[110] br[110] wl[223] vdd gnd cell_6t
Xbit_r224_c110 bl[110] br[110] wl[224] vdd gnd cell_6t
Xbit_r225_c110 bl[110] br[110] wl[225] vdd gnd cell_6t
Xbit_r226_c110 bl[110] br[110] wl[226] vdd gnd cell_6t
Xbit_r227_c110 bl[110] br[110] wl[227] vdd gnd cell_6t
Xbit_r228_c110 bl[110] br[110] wl[228] vdd gnd cell_6t
Xbit_r229_c110 bl[110] br[110] wl[229] vdd gnd cell_6t
Xbit_r230_c110 bl[110] br[110] wl[230] vdd gnd cell_6t
Xbit_r231_c110 bl[110] br[110] wl[231] vdd gnd cell_6t
Xbit_r232_c110 bl[110] br[110] wl[232] vdd gnd cell_6t
Xbit_r233_c110 bl[110] br[110] wl[233] vdd gnd cell_6t
Xbit_r234_c110 bl[110] br[110] wl[234] vdd gnd cell_6t
Xbit_r235_c110 bl[110] br[110] wl[235] vdd gnd cell_6t
Xbit_r236_c110 bl[110] br[110] wl[236] vdd gnd cell_6t
Xbit_r237_c110 bl[110] br[110] wl[237] vdd gnd cell_6t
Xbit_r238_c110 bl[110] br[110] wl[238] vdd gnd cell_6t
Xbit_r239_c110 bl[110] br[110] wl[239] vdd gnd cell_6t
Xbit_r240_c110 bl[110] br[110] wl[240] vdd gnd cell_6t
Xbit_r241_c110 bl[110] br[110] wl[241] vdd gnd cell_6t
Xbit_r242_c110 bl[110] br[110] wl[242] vdd gnd cell_6t
Xbit_r243_c110 bl[110] br[110] wl[243] vdd gnd cell_6t
Xbit_r244_c110 bl[110] br[110] wl[244] vdd gnd cell_6t
Xbit_r245_c110 bl[110] br[110] wl[245] vdd gnd cell_6t
Xbit_r246_c110 bl[110] br[110] wl[246] vdd gnd cell_6t
Xbit_r247_c110 bl[110] br[110] wl[247] vdd gnd cell_6t
Xbit_r248_c110 bl[110] br[110] wl[248] vdd gnd cell_6t
Xbit_r249_c110 bl[110] br[110] wl[249] vdd gnd cell_6t
Xbit_r250_c110 bl[110] br[110] wl[250] vdd gnd cell_6t
Xbit_r251_c110 bl[110] br[110] wl[251] vdd gnd cell_6t
Xbit_r252_c110 bl[110] br[110] wl[252] vdd gnd cell_6t
Xbit_r253_c110 bl[110] br[110] wl[253] vdd gnd cell_6t
Xbit_r254_c110 bl[110] br[110] wl[254] vdd gnd cell_6t
Xbit_r255_c110 bl[110] br[110] wl[255] vdd gnd cell_6t
Xbit_r256_c110 bl[110] br[110] wl[256] vdd gnd cell_6t
Xbit_r257_c110 bl[110] br[110] wl[257] vdd gnd cell_6t
Xbit_r258_c110 bl[110] br[110] wl[258] vdd gnd cell_6t
Xbit_r259_c110 bl[110] br[110] wl[259] vdd gnd cell_6t
Xbit_r260_c110 bl[110] br[110] wl[260] vdd gnd cell_6t
Xbit_r261_c110 bl[110] br[110] wl[261] vdd gnd cell_6t
Xbit_r262_c110 bl[110] br[110] wl[262] vdd gnd cell_6t
Xbit_r263_c110 bl[110] br[110] wl[263] vdd gnd cell_6t
Xbit_r264_c110 bl[110] br[110] wl[264] vdd gnd cell_6t
Xbit_r265_c110 bl[110] br[110] wl[265] vdd gnd cell_6t
Xbit_r266_c110 bl[110] br[110] wl[266] vdd gnd cell_6t
Xbit_r267_c110 bl[110] br[110] wl[267] vdd gnd cell_6t
Xbit_r268_c110 bl[110] br[110] wl[268] vdd gnd cell_6t
Xbit_r269_c110 bl[110] br[110] wl[269] vdd gnd cell_6t
Xbit_r270_c110 bl[110] br[110] wl[270] vdd gnd cell_6t
Xbit_r271_c110 bl[110] br[110] wl[271] vdd gnd cell_6t
Xbit_r272_c110 bl[110] br[110] wl[272] vdd gnd cell_6t
Xbit_r273_c110 bl[110] br[110] wl[273] vdd gnd cell_6t
Xbit_r274_c110 bl[110] br[110] wl[274] vdd gnd cell_6t
Xbit_r275_c110 bl[110] br[110] wl[275] vdd gnd cell_6t
Xbit_r276_c110 bl[110] br[110] wl[276] vdd gnd cell_6t
Xbit_r277_c110 bl[110] br[110] wl[277] vdd gnd cell_6t
Xbit_r278_c110 bl[110] br[110] wl[278] vdd gnd cell_6t
Xbit_r279_c110 bl[110] br[110] wl[279] vdd gnd cell_6t
Xbit_r280_c110 bl[110] br[110] wl[280] vdd gnd cell_6t
Xbit_r281_c110 bl[110] br[110] wl[281] vdd gnd cell_6t
Xbit_r282_c110 bl[110] br[110] wl[282] vdd gnd cell_6t
Xbit_r283_c110 bl[110] br[110] wl[283] vdd gnd cell_6t
Xbit_r284_c110 bl[110] br[110] wl[284] vdd gnd cell_6t
Xbit_r285_c110 bl[110] br[110] wl[285] vdd gnd cell_6t
Xbit_r286_c110 bl[110] br[110] wl[286] vdd gnd cell_6t
Xbit_r287_c110 bl[110] br[110] wl[287] vdd gnd cell_6t
Xbit_r288_c110 bl[110] br[110] wl[288] vdd gnd cell_6t
Xbit_r289_c110 bl[110] br[110] wl[289] vdd gnd cell_6t
Xbit_r290_c110 bl[110] br[110] wl[290] vdd gnd cell_6t
Xbit_r291_c110 bl[110] br[110] wl[291] vdd gnd cell_6t
Xbit_r292_c110 bl[110] br[110] wl[292] vdd gnd cell_6t
Xbit_r293_c110 bl[110] br[110] wl[293] vdd gnd cell_6t
Xbit_r294_c110 bl[110] br[110] wl[294] vdd gnd cell_6t
Xbit_r295_c110 bl[110] br[110] wl[295] vdd gnd cell_6t
Xbit_r296_c110 bl[110] br[110] wl[296] vdd gnd cell_6t
Xbit_r297_c110 bl[110] br[110] wl[297] vdd gnd cell_6t
Xbit_r298_c110 bl[110] br[110] wl[298] vdd gnd cell_6t
Xbit_r299_c110 bl[110] br[110] wl[299] vdd gnd cell_6t
Xbit_r300_c110 bl[110] br[110] wl[300] vdd gnd cell_6t
Xbit_r301_c110 bl[110] br[110] wl[301] vdd gnd cell_6t
Xbit_r302_c110 bl[110] br[110] wl[302] vdd gnd cell_6t
Xbit_r303_c110 bl[110] br[110] wl[303] vdd gnd cell_6t
Xbit_r304_c110 bl[110] br[110] wl[304] vdd gnd cell_6t
Xbit_r305_c110 bl[110] br[110] wl[305] vdd gnd cell_6t
Xbit_r306_c110 bl[110] br[110] wl[306] vdd gnd cell_6t
Xbit_r307_c110 bl[110] br[110] wl[307] vdd gnd cell_6t
Xbit_r308_c110 bl[110] br[110] wl[308] vdd gnd cell_6t
Xbit_r309_c110 bl[110] br[110] wl[309] vdd gnd cell_6t
Xbit_r310_c110 bl[110] br[110] wl[310] vdd gnd cell_6t
Xbit_r311_c110 bl[110] br[110] wl[311] vdd gnd cell_6t
Xbit_r312_c110 bl[110] br[110] wl[312] vdd gnd cell_6t
Xbit_r313_c110 bl[110] br[110] wl[313] vdd gnd cell_6t
Xbit_r314_c110 bl[110] br[110] wl[314] vdd gnd cell_6t
Xbit_r315_c110 bl[110] br[110] wl[315] vdd gnd cell_6t
Xbit_r316_c110 bl[110] br[110] wl[316] vdd gnd cell_6t
Xbit_r317_c110 bl[110] br[110] wl[317] vdd gnd cell_6t
Xbit_r318_c110 bl[110] br[110] wl[318] vdd gnd cell_6t
Xbit_r319_c110 bl[110] br[110] wl[319] vdd gnd cell_6t
Xbit_r320_c110 bl[110] br[110] wl[320] vdd gnd cell_6t
Xbit_r321_c110 bl[110] br[110] wl[321] vdd gnd cell_6t
Xbit_r322_c110 bl[110] br[110] wl[322] vdd gnd cell_6t
Xbit_r323_c110 bl[110] br[110] wl[323] vdd gnd cell_6t
Xbit_r324_c110 bl[110] br[110] wl[324] vdd gnd cell_6t
Xbit_r325_c110 bl[110] br[110] wl[325] vdd gnd cell_6t
Xbit_r326_c110 bl[110] br[110] wl[326] vdd gnd cell_6t
Xbit_r327_c110 bl[110] br[110] wl[327] vdd gnd cell_6t
Xbit_r328_c110 bl[110] br[110] wl[328] vdd gnd cell_6t
Xbit_r329_c110 bl[110] br[110] wl[329] vdd gnd cell_6t
Xbit_r330_c110 bl[110] br[110] wl[330] vdd gnd cell_6t
Xbit_r331_c110 bl[110] br[110] wl[331] vdd gnd cell_6t
Xbit_r332_c110 bl[110] br[110] wl[332] vdd gnd cell_6t
Xbit_r333_c110 bl[110] br[110] wl[333] vdd gnd cell_6t
Xbit_r334_c110 bl[110] br[110] wl[334] vdd gnd cell_6t
Xbit_r335_c110 bl[110] br[110] wl[335] vdd gnd cell_6t
Xbit_r336_c110 bl[110] br[110] wl[336] vdd gnd cell_6t
Xbit_r337_c110 bl[110] br[110] wl[337] vdd gnd cell_6t
Xbit_r338_c110 bl[110] br[110] wl[338] vdd gnd cell_6t
Xbit_r339_c110 bl[110] br[110] wl[339] vdd gnd cell_6t
Xbit_r340_c110 bl[110] br[110] wl[340] vdd gnd cell_6t
Xbit_r341_c110 bl[110] br[110] wl[341] vdd gnd cell_6t
Xbit_r342_c110 bl[110] br[110] wl[342] vdd gnd cell_6t
Xbit_r343_c110 bl[110] br[110] wl[343] vdd gnd cell_6t
Xbit_r344_c110 bl[110] br[110] wl[344] vdd gnd cell_6t
Xbit_r345_c110 bl[110] br[110] wl[345] vdd gnd cell_6t
Xbit_r346_c110 bl[110] br[110] wl[346] vdd gnd cell_6t
Xbit_r347_c110 bl[110] br[110] wl[347] vdd gnd cell_6t
Xbit_r348_c110 bl[110] br[110] wl[348] vdd gnd cell_6t
Xbit_r349_c110 bl[110] br[110] wl[349] vdd gnd cell_6t
Xbit_r350_c110 bl[110] br[110] wl[350] vdd gnd cell_6t
Xbit_r351_c110 bl[110] br[110] wl[351] vdd gnd cell_6t
Xbit_r352_c110 bl[110] br[110] wl[352] vdd gnd cell_6t
Xbit_r353_c110 bl[110] br[110] wl[353] vdd gnd cell_6t
Xbit_r354_c110 bl[110] br[110] wl[354] vdd gnd cell_6t
Xbit_r355_c110 bl[110] br[110] wl[355] vdd gnd cell_6t
Xbit_r356_c110 bl[110] br[110] wl[356] vdd gnd cell_6t
Xbit_r357_c110 bl[110] br[110] wl[357] vdd gnd cell_6t
Xbit_r358_c110 bl[110] br[110] wl[358] vdd gnd cell_6t
Xbit_r359_c110 bl[110] br[110] wl[359] vdd gnd cell_6t
Xbit_r360_c110 bl[110] br[110] wl[360] vdd gnd cell_6t
Xbit_r361_c110 bl[110] br[110] wl[361] vdd gnd cell_6t
Xbit_r362_c110 bl[110] br[110] wl[362] vdd gnd cell_6t
Xbit_r363_c110 bl[110] br[110] wl[363] vdd gnd cell_6t
Xbit_r364_c110 bl[110] br[110] wl[364] vdd gnd cell_6t
Xbit_r365_c110 bl[110] br[110] wl[365] vdd gnd cell_6t
Xbit_r366_c110 bl[110] br[110] wl[366] vdd gnd cell_6t
Xbit_r367_c110 bl[110] br[110] wl[367] vdd gnd cell_6t
Xbit_r368_c110 bl[110] br[110] wl[368] vdd gnd cell_6t
Xbit_r369_c110 bl[110] br[110] wl[369] vdd gnd cell_6t
Xbit_r370_c110 bl[110] br[110] wl[370] vdd gnd cell_6t
Xbit_r371_c110 bl[110] br[110] wl[371] vdd gnd cell_6t
Xbit_r372_c110 bl[110] br[110] wl[372] vdd gnd cell_6t
Xbit_r373_c110 bl[110] br[110] wl[373] vdd gnd cell_6t
Xbit_r374_c110 bl[110] br[110] wl[374] vdd gnd cell_6t
Xbit_r375_c110 bl[110] br[110] wl[375] vdd gnd cell_6t
Xbit_r376_c110 bl[110] br[110] wl[376] vdd gnd cell_6t
Xbit_r377_c110 bl[110] br[110] wl[377] vdd gnd cell_6t
Xbit_r378_c110 bl[110] br[110] wl[378] vdd gnd cell_6t
Xbit_r379_c110 bl[110] br[110] wl[379] vdd gnd cell_6t
Xbit_r380_c110 bl[110] br[110] wl[380] vdd gnd cell_6t
Xbit_r381_c110 bl[110] br[110] wl[381] vdd gnd cell_6t
Xbit_r382_c110 bl[110] br[110] wl[382] vdd gnd cell_6t
Xbit_r383_c110 bl[110] br[110] wl[383] vdd gnd cell_6t
Xbit_r384_c110 bl[110] br[110] wl[384] vdd gnd cell_6t
Xbit_r385_c110 bl[110] br[110] wl[385] vdd gnd cell_6t
Xbit_r386_c110 bl[110] br[110] wl[386] vdd gnd cell_6t
Xbit_r387_c110 bl[110] br[110] wl[387] vdd gnd cell_6t
Xbit_r388_c110 bl[110] br[110] wl[388] vdd gnd cell_6t
Xbit_r389_c110 bl[110] br[110] wl[389] vdd gnd cell_6t
Xbit_r390_c110 bl[110] br[110] wl[390] vdd gnd cell_6t
Xbit_r391_c110 bl[110] br[110] wl[391] vdd gnd cell_6t
Xbit_r392_c110 bl[110] br[110] wl[392] vdd gnd cell_6t
Xbit_r393_c110 bl[110] br[110] wl[393] vdd gnd cell_6t
Xbit_r394_c110 bl[110] br[110] wl[394] vdd gnd cell_6t
Xbit_r395_c110 bl[110] br[110] wl[395] vdd gnd cell_6t
Xbit_r396_c110 bl[110] br[110] wl[396] vdd gnd cell_6t
Xbit_r397_c110 bl[110] br[110] wl[397] vdd gnd cell_6t
Xbit_r398_c110 bl[110] br[110] wl[398] vdd gnd cell_6t
Xbit_r399_c110 bl[110] br[110] wl[399] vdd gnd cell_6t
Xbit_r400_c110 bl[110] br[110] wl[400] vdd gnd cell_6t
Xbit_r401_c110 bl[110] br[110] wl[401] vdd gnd cell_6t
Xbit_r402_c110 bl[110] br[110] wl[402] vdd gnd cell_6t
Xbit_r403_c110 bl[110] br[110] wl[403] vdd gnd cell_6t
Xbit_r404_c110 bl[110] br[110] wl[404] vdd gnd cell_6t
Xbit_r405_c110 bl[110] br[110] wl[405] vdd gnd cell_6t
Xbit_r406_c110 bl[110] br[110] wl[406] vdd gnd cell_6t
Xbit_r407_c110 bl[110] br[110] wl[407] vdd gnd cell_6t
Xbit_r408_c110 bl[110] br[110] wl[408] vdd gnd cell_6t
Xbit_r409_c110 bl[110] br[110] wl[409] vdd gnd cell_6t
Xbit_r410_c110 bl[110] br[110] wl[410] vdd gnd cell_6t
Xbit_r411_c110 bl[110] br[110] wl[411] vdd gnd cell_6t
Xbit_r412_c110 bl[110] br[110] wl[412] vdd gnd cell_6t
Xbit_r413_c110 bl[110] br[110] wl[413] vdd gnd cell_6t
Xbit_r414_c110 bl[110] br[110] wl[414] vdd gnd cell_6t
Xbit_r415_c110 bl[110] br[110] wl[415] vdd gnd cell_6t
Xbit_r416_c110 bl[110] br[110] wl[416] vdd gnd cell_6t
Xbit_r417_c110 bl[110] br[110] wl[417] vdd gnd cell_6t
Xbit_r418_c110 bl[110] br[110] wl[418] vdd gnd cell_6t
Xbit_r419_c110 bl[110] br[110] wl[419] vdd gnd cell_6t
Xbit_r420_c110 bl[110] br[110] wl[420] vdd gnd cell_6t
Xbit_r421_c110 bl[110] br[110] wl[421] vdd gnd cell_6t
Xbit_r422_c110 bl[110] br[110] wl[422] vdd gnd cell_6t
Xbit_r423_c110 bl[110] br[110] wl[423] vdd gnd cell_6t
Xbit_r424_c110 bl[110] br[110] wl[424] vdd gnd cell_6t
Xbit_r425_c110 bl[110] br[110] wl[425] vdd gnd cell_6t
Xbit_r426_c110 bl[110] br[110] wl[426] vdd gnd cell_6t
Xbit_r427_c110 bl[110] br[110] wl[427] vdd gnd cell_6t
Xbit_r428_c110 bl[110] br[110] wl[428] vdd gnd cell_6t
Xbit_r429_c110 bl[110] br[110] wl[429] vdd gnd cell_6t
Xbit_r430_c110 bl[110] br[110] wl[430] vdd gnd cell_6t
Xbit_r431_c110 bl[110] br[110] wl[431] vdd gnd cell_6t
Xbit_r432_c110 bl[110] br[110] wl[432] vdd gnd cell_6t
Xbit_r433_c110 bl[110] br[110] wl[433] vdd gnd cell_6t
Xbit_r434_c110 bl[110] br[110] wl[434] vdd gnd cell_6t
Xbit_r435_c110 bl[110] br[110] wl[435] vdd gnd cell_6t
Xbit_r436_c110 bl[110] br[110] wl[436] vdd gnd cell_6t
Xbit_r437_c110 bl[110] br[110] wl[437] vdd gnd cell_6t
Xbit_r438_c110 bl[110] br[110] wl[438] vdd gnd cell_6t
Xbit_r439_c110 bl[110] br[110] wl[439] vdd gnd cell_6t
Xbit_r440_c110 bl[110] br[110] wl[440] vdd gnd cell_6t
Xbit_r441_c110 bl[110] br[110] wl[441] vdd gnd cell_6t
Xbit_r442_c110 bl[110] br[110] wl[442] vdd gnd cell_6t
Xbit_r443_c110 bl[110] br[110] wl[443] vdd gnd cell_6t
Xbit_r444_c110 bl[110] br[110] wl[444] vdd gnd cell_6t
Xbit_r445_c110 bl[110] br[110] wl[445] vdd gnd cell_6t
Xbit_r446_c110 bl[110] br[110] wl[446] vdd gnd cell_6t
Xbit_r447_c110 bl[110] br[110] wl[447] vdd gnd cell_6t
Xbit_r448_c110 bl[110] br[110] wl[448] vdd gnd cell_6t
Xbit_r449_c110 bl[110] br[110] wl[449] vdd gnd cell_6t
Xbit_r450_c110 bl[110] br[110] wl[450] vdd gnd cell_6t
Xbit_r451_c110 bl[110] br[110] wl[451] vdd gnd cell_6t
Xbit_r452_c110 bl[110] br[110] wl[452] vdd gnd cell_6t
Xbit_r453_c110 bl[110] br[110] wl[453] vdd gnd cell_6t
Xbit_r454_c110 bl[110] br[110] wl[454] vdd gnd cell_6t
Xbit_r455_c110 bl[110] br[110] wl[455] vdd gnd cell_6t
Xbit_r456_c110 bl[110] br[110] wl[456] vdd gnd cell_6t
Xbit_r457_c110 bl[110] br[110] wl[457] vdd gnd cell_6t
Xbit_r458_c110 bl[110] br[110] wl[458] vdd gnd cell_6t
Xbit_r459_c110 bl[110] br[110] wl[459] vdd gnd cell_6t
Xbit_r460_c110 bl[110] br[110] wl[460] vdd gnd cell_6t
Xbit_r461_c110 bl[110] br[110] wl[461] vdd gnd cell_6t
Xbit_r462_c110 bl[110] br[110] wl[462] vdd gnd cell_6t
Xbit_r463_c110 bl[110] br[110] wl[463] vdd gnd cell_6t
Xbit_r464_c110 bl[110] br[110] wl[464] vdd gnd cell_6t
Xbit_r465_c110 bl[110] br[110] wl[465] vdd gnd cell_6t
Xbit_r466_c110 bl[110] br[110] wl[466] vdd gnd cell_6t
Xbit_r467_c110 bl[110] br[110] wl[467] vdd gnd cell_6t
Xbit_r468_c110 bl[110] br[110] wl[468] vdd gnd cell_6t
Xbit_r469_c110 bl[110] br[110] wl[469] vdd gnd cell_6t
Xbit_r470_c110 bl[110] br[110] wl[470] vdd gnd cell_6t
Xbit_r471_c110 bl[110] br[110] wl[471] vdd gnd cell_6t
Xbit_r472_c110 bl[110] br[110] wl[472] vdd gnd cell_6t
Xbit_r473_c110 bl[110] br[110] wl[473] vdd gnd cell_6t
Xbit_r474_c110 bl[110] br[110] wl[474] vdd gnd cell_6t
Xbit_r475_c110 bl[110] br[110] wl[475] vdd gnd cell_6t
Xbit_r476_c110 bl[110] br[110] wl[476] vdd gnd cell_6t
Xbit_r477_c110 bl[110] br[110] wl[477] vdd gnd cell_6t
Xbit_r478_c110 bl[110] br[110] wl[478] vdd gnd cell_6t
Xbit_r479_c110 bl[110] br[110] wl[479] vdd gnd cell_6t
Xbit_r480_c110 bl[110] br[110] wl[480] vdd gnd cell_6t
Xbit_r481_c110 bl[110] br[110] wl[481] vdd gnd cell_6t
Xbit_r482_c110 bl[110] br[110] wl[482] vdd gnd cell_6t
Xbit_r483_c110 bl[110] br[110] wl[483] vdd gnd cell_6t
Xbit_r484_c110 bl[110] br[110] wl[484] vdd gnd cell_6t
Xbit_r485_c110 bl[110] br[110] wl[485] vdd gnd cell_6t
Xbit_r486_c110 bl[110] br[110] wl[486] vdd gnd cell_6t
Xbit_r487_c110 bl[110] br[110] wl[487] vdd gnd cell_6t
Xbit_r488_c110 bl[110] br[110] wl[488] vdd gnd cell_6t
Xbit_r489_c110 bl[110] br[110] wl[489] vdd gnd cell_6t
Xbit_r490_c110 bl[110] br[110] wl[490] vdd gnd cell_6t
Xbit_r491_c110 bl[110] br[110] wl[491] vdd gnd cell_6t
Xbit_r492_c110 bl[110] br[110] wl[492] vdd gnd cell_6t
Xbit_r493_c110 bl[110] br[110] wl[493] vdd gnd cell_6t
Xbit_r494_c110 bl[110] br[110] wl[494] vdd gnd cell_6t
Xbit_r495_c110 bl[110] br[110] wl[495] vdd gnd cell_6t
Xbit_r496_c110 bl[110] br[110] wl[496] vdd gnd cell_6t
Xbit_r497_c110 bl[110] br[110] wl[497] vdd gnd cell_6t
Xbit_r498_c110 bl[110] br[110] wl[498] vdd gnd cell_6t
Xbit_r499_c110 bl[110] br[110] wl[499] vdd gnd cell_6t
Xbit_r500_c110 bl[110] br[110] wl[500] vdd gnd cell_6t
Xbit_r501_c110 bl[110] br[110] wl[501] vdd gnd cell_6t
Xbit_r502_c110 bl[110] br[110] wl[502] vdd gnd cell_6t
Xbit_r503_c110 bl[110] br[110] wl[503] vdd gnd cell_6t
Xbit_r504_c110 bl[110] br[110] wl[504] vdd gnd cell_6t
Xbit_r505_c110 bl[110] br[110] wl[505] vdd gnd cell_6t
Xbit_r506_c110 bl[110] br[110] wl[506] vdd gnd cell_6t
Xbit_r507_c110 bl[110] br[110] wl[507] vdd gnd cell_6t
Xbit_r508_c110 bl[110] br[110] wl[508] vdd gnd cell_6t
Xbit_r509_c110 bl[110] br[110] wl[509] vdd gnd cell_6t
Xbit_r510_c110 bl[110] br[110] wl[510] vdd gnd cell_6t
Xbit_r511_c110 bl[110] br[110] wl[511] vdd gnd cell_6t
Xbit_r0_c111 bl[111] br[111] wl[0] vdd gnd cell_6t
Xbit_r1_c111 bl[111] br[111] wl[1] vdd gnd cell_6t
Xbit_r2_c111 bl[111] br[111] wl[2] vdd gnd cell_6t
Xbit_r3_c111 bl[111] br[111] wl[3] vdd gnd cell_6t
Xbit_r4_c111 bl[111] br[111] wl[4] vdd gnd cell_6t
Xbit_r5_c111 bl[111] br[111] wl[5] vdd gnd cell_6t
Xbit_r6_c111 bl[111] br[111] wl[6] vdd gnd cell_6t
Xbit_r7_c111 bl[111] br[111] wl[7] vdd gnd cell_6t
Xbit_r8_c111 bl[111] br[111] wl[8] vdd gnd cell_6t
Xbit_r9_c111 bl[111] br[111] wl[9] vdd gnd cell_6t
Xbit_r10_c111 bl[111] br[111] wl[10] vdd gnd cell_6t
Xbit_r11_c111 bl[111] br[111] wl[11] vdd gnd cell_6t
Xbit_r12_c111 bl[111] br[111] wl[12] vdd gnd cell_6t
Xbit_r13_c111 bl[111] br[111] wl[13] vdd gnd cell_6t
Xbit_r14_c111 bl[111] br[111] wl[14] vdd gnd cell_6t
Xbit_r15_c111 bl[111] br[111] wl[15] vdd gnd cell_6t
Xbit_r16_c111 bl[111] br[111] wl[16] vdd gnd cell_6t
Xbit_r17_c111 bl[111] br[111] wl[17] vdd gnd cell_6t
Xbit_r18_c111 bl[111] br[111] wl[18] vdd gnd cell_6t
Xbit_r19_c111 bl[111] br[111] wl[19] vdd gnd cell_6t
Xbit_r20_c111 bl[111] br[111] wl[20] vdd gnd cell_6t
Xbit_r21_c111 bl[111] br[111] wl[21] vdd gnd cell_6t
Xbit_r22_c111 bl[111] br[111] wl[22] vdd gnd cell_6t
Xbit_r23_c111 bl[111] br[111] wl[23] vdd gnd cell_6t
Xbit_r24_c111 bl[111] br[111] wl[24] vdd gnd cell_6t
Xbit_r25_c111 bl[111] br[111] wl[25] vdd gnd cell_6t
Xbit_r26_c111 bl[111] br[111] wl[26] vdd gnd cell_6t
Xbit_r27_c111 bl[111] br[111] wl[27] vdd gnd cell_6t
Xbit_r28_c111 bl[111] br[111] wl[28] vdd gnd cell_6t
Xbit_r29_c111 bl[111] br[111] wl[29] vdd gnd cell_6t
Xbit_r30_c111 bl[111] br[111] wl[30] vdd gnd cell_6t
Xbit_r31_c111 bl[111] br[111] wl[31] vdd gnd cell_6t
Xbit_r32_c111 bl[111] br[111] wl[32] vdd gnd cell_6t
Xbit_r33_c111 bl[111] br[111] wl[33] vdd gnd cell_6t
Xbit_r34_c111 bl[111] br[111] wl[34] vdd gnd cell_6t
Xbit_r35_c111 bl[111] br[111] wl[35] vdd gnd cell_6t
Xbit_r36_c111 bl[111] br[111] wl[36] vdd gnd cell_6t
Xbit_r37_c111 bl[111] br[111] wl[37] vdd gnd cell_6t
Xbit_r38_c111 bl[111] br[111] wl[38] vdd gnd cell_6t
Xbit_r39_c111 bl[111] br[111] wl[39] vdd gnd cell_6t
Xbit_r40_c111 bl[111] br[111] wl[40] vdd gnd cell_6t
Xbit_r41_c111 bl[111] br[111] wl[41] vdd gnd cell_6t
Xbit_r42_c111 bl[111] br[111] wl[42] vdd gnd cell_6t
Xbit_r43_c111 bl[111] br[111] wl[43] vdd gnd cell_6t
Xbit_r44_c111 bl[111] br[111] wl[44] vdd gnd cell_6t
Xbit_r45_c111 bl[111] br[111] wl[45] vdd gnd cell_6t
Xbit_r46_c111 bl[111] br[111] wl[46] vdd gnd cell_6t
Xbit_r47_c111 bl[111] br[111] wl[47] vdd gnd cell_6t
Xbit_r48_c111 bl[111] br[111] wl[48] vdd gnd cell_6t
Xbit_r49_c111 bl[111] br[111] wl[49] vdd gnd cell_6t
Xbit_r50_c111 bl[111] br[111] wl[50] vdd gnd cell_6t
Xbit_r51_c111 bl[111] br[111] wl[51] vdd gnd cell_6t
Xbit_r52_c111 bl[111] br[111] wl[52] vdd gnd cell_6t
Xbit_r53_c111 bl[111] br[111] wl[53] vdd gnd cell_6t
Xbit_r54_c111 bl[111] br[111] wl[54] vdd gnd cell_6t
Xbit_r55_c111 bl[111] br[111] wl[55] vdd gnd cell_6t
Xbit_r56_c111 bl[111] br[111] wl[56] vdd gnd cell_6t
Xbit_r57_c111 bl[111] br[111] wl[57] vdd gnd cell_6t
Xbit_r58_c111 bl[111] br[111] wl[58] vdd gnd cell_6t
Xbit_r59_c111 bl[111] br[111] wl[59] vdd gnd cell_6t
Xbit_r60_c111 bl[111] br[111] wl[60] vdd gnd cell_6t
Xbit_r61_c111 bl[111] br[111] wl[61] vdd gnd cell_6t
Xbit_r62_c111 bl[111] br[111] wl[62] vdd gnd cell_6t
Xbit_r63_c111 bl[111] br[111] wl[63] vdd gnd cell_6t
Xbit_r64_c111 bl[111] br[111] wl[64] vdd gnd cell_6t
Xbit_r65_c111 bl[111] br[111] wl[65] vdd gnd cell_6t
Xbit_r66_c111 bl[111] br[111] wl[66] vdd gnd cell_6t
Xbit_r67_c111 bl[111] br[111] wl[67] vdd gnd cell_6t
Xbit_r68_c111 bl[111] br[111] wl[68] vdd gnd cell_6t
Xbit_r69_c111 bl[111] br[111] wl[69] vdd gnd cell_6t
Xbit_r70_c111 bl[111] br[111] wl[70] vdd gnd cell_6t
Xbit_r71_c111 bl[111] br[111] wl[71] vdd gnd cell_6t
Xbit_r72_c111 bl[111] br[111] wl[72] vdd gnd cell_6t
Xbit_r73_c111 bl[111] br[111] wl[73] vdd gnd cell_6t
Xbit_r74_c111 bl[111] br[111] wl[74] vdd gnd cell_6t
Xbit_r75_c111 bl[111] br[111] wl[75] vdd gnd cell_6t
Xbit_r76_c111 bl[111] br[111] wl[76] vdd gnd cell_6t
Xbit_r77_c111 bl[111] br[111] wl[77] vdd gnd cell_6t
Xbit_r78_c111 bl[111] br[111] wl[78] vdd gnd cell_6t
Xbit_r79_c111 bl[111] br[111] wl[79] vdd gnd cell_6t
Xbit_r80_c111 bl[111] br[111] wl[80] vdd gnd cell_6t
Xbit_r81_c111 bl[111] br[111] wl[81] vdd gnd cell_6t
Xbit_r82_c111 bl[111] br[111] wl[82] vdd gnd cell_6t
Xbit_r83_c111 bl[111] br[111] wl[83] vdd gnd cell_6t
Xbit_r84_c111 bl[111] br[111] wl[84] vdd gnd cell_6t
Xbit_r85_c111 bl[111] br[111] wl[85] vdd gnd cell_6t
Xbit_r86_c111 bl[111] br[111] wl[86] vdd gnd cell_6t
Xbit_r87_c111 bl[111] br[111] wl[87] vdd gnd cell_6t
Xbit_r88_c111 bl[111] br[111] wl[88] vdd gnd cell_6t
Xbit_r89_c111 bl[111] br[111] wl[89] vdd gnd cell_6t
Xbit_r90_c111 bl[111] br[111] wl[90] vdd gnd cell_6t
Xbit_r91_c111 bl[111] br[111] wl[91] vdd gnd cell_6t
Xbit_r92_c111 bl[111] br[111] wl[92] vdd gnd cell_6t
Xbit_r93_c111 bl[111] br[111] wl[93] vdd gnd cell_6t
Xbit_r94_c111 bl[111] br[111] wl[94] vdd gnd cell_6t
Xbit_r95_c111 bl[111] br[111] wl[95] vdd gnd cell_6t
Xbit_r96_c111 bl[111] br[111] wl[96] vdd gnd cell_6t
Xbit_r97_c111 bl[111] br[111] wl[97] vdd gnd cell_6t
Xbit_r98_c111 bl[111] br[111] wl[98] vdd gnd cell_6t
Xbit_r99_c111 bl[111] br[111] wl[99] vdd gnd cell_6t
Xbit_r100_c111 bl[111] br[111] wl[100] vdd gnd cell_6t
Xbit_r101_c111 bl[111] br[111] wl[101] vdd gnd cell_6t
Xbit_r102_c111 bl[111] br[111] wl[102] vdd gnd cell_6t
Xbit_r103_c111 bl[111] br[111] wl[103] vdd gnd cell_6t
Xbit_r104_c111 bl[111] br[111] wl[104] vdd gnd cell_6t
Xbit_r105_c111 bl[111] br[111] wl[105] vdd gnd cell_6t
Xbit_r106_c111 bl[111] br[111] wl[106] vdd gnd cell_6t
Xbit_r107_c111 bl[111] br[111] wl[107] vdd gnd cell_6t
Xbit_r108_c111 bl[111] br[111] wl[108] vdd gnd cell_6t
Xbit_r109_c111 bl[111] br[111] wl[109] vdd gnd cell_6t
Xbit_r110_c111 bl[111] br[111] wl[110] vdd gnd cell_6t
Xbit_r111_c111 bl[111] br[111] wl[111] vdd gnd cell_6t
Xbit_r112_c111 bl[111] br[111] wl[112] vdd gnd cell_6t
Xbit_r113_c111 bl[111] br[111] wl[113] vdd gnd cell_6t
Xbit_r114_c111 bl[111] br[111] wl[114] vdd gnd cell_6t
Xbit_r115_c111 bl[111] br[111] wl[115] vdd gnd cell_6t
Xbit_r116_c111 bl[111] br[111] wl[116] vdd gnd cell_6t
Xbit_r117_c111 bl[111] br[111] wl[117] vdd gnd cell_6t
Xbit_r118_c111 bl[111] br[111] wl[118] vdd gnd cell_6t
Xbit_r119_c111 bl[111] br[111] wl[119] vdd gnd cell_6t
Xbit_r120_c111 bl[111] br[111] wl[120] vdd gnd cell_6t
Xbit_r121_c111 bl[111] br[111] wl[121] vdd gnd cell_6t
Xbit_r122_c111 bl[111] br[111] wl[122] vdd gnd cell_6t
Xbit_r123_c111 bl[111] br[111] wl[123] vdd gnd cell_6t
Xbit_r124_c111 bl[111] br[111] wl[124] vdd gnd cell_6t
Xbit_r125_c111 bl[111] br[111] wl[125] vdd gnd cell_6t
Xbit_r126_c111 bl[111] br[111] wl[126] vdd gnd cell_6t
Xbit_r127_c111 bl[111] br[111] wl[127] vdd gnd cell_6t
Xbit_r128_c111 bl[111] br[111] wl[128] vdd gnd cell_6t
Xbit_r129_c111 bl[111] br[111] wl[129] vdd gnd cell_6t
Xbit_r130_c111 bl[111] br[111] wl[130] vdd gnd cell_6t
Xbit_r131_c111 bl[111] br[111] wl[131] vdd gnd cell_6t
Xbit_r132_c111 bl[111] br[111] wl[132] vdd gnd cell_6t
Xbit_r133_c111 bl[111] br[111] wl[133] vdd gnd cell_6t
Xbit_r134_c111 bl[111] br[111] wl[134] vdd gnd cell_6t
Xbit_r135_c111 bl[111] br[111] wl[135] vdd gnd cell_6t
Xbit_r136_c111 bl[111] br[111] wl[136] vdd gnd cell_6t
Xbit_r137_c111 bl[111] br[111] wl[137] vdd gnd cell_6t
Xbit_r138_c111 bl[111] br[111] wl[138] vdd gnd cell_6t
Xbit_r139_c111 bl[111] br[111] wl[139] vdd gnd cell_6t
Xbit_r140_c111 bl[111] br[111] wl[140] vdd gnd cell_6t
Xbit_r141_c111 bl[111] br[111] wl[141] vdd gnd cell_6t
Xbit_r142_c111 bl[111] br[111] wl[142] vdd gnd cell_6t
Xbit_r143_c111 bl[111] br[111] wl[143] vdd gnd cell_6t
Xbit_r144_c111 bl[111] br[111] wl[144] vdd gnd cell_6t
Xbit_r145_c111 bl[111] br[111] wl[145] vdd gnd cell_6t
Xbit_r146_c111 bl[111] br[111] wl[146] vdd gnd cell_6t
Xbit_r147_c111 bl[111] br[111] wl[147] vdd gnd cell_6t
Xbit_r148_c111 bl[111] br[111] wl[148] vdd gnd cell_6t
Xbit_r149_c111 bl[111] br[111] wl[149] vdd gnd cell_6t
Xbit_r150_c111 bl[111] br[111] wl[150] vdd gnd cell_6t
Xbit_r151_c111 bl[111] br[111] wl[151] vdd gnd cell_6t
Xbit_r152_c111 bl[111] br[111] wl[152] vdd gnd cell_6t
Xbit_r153_c111 bl[111] br[111] wl[153] vdd gnd cell_6t
Xbit_r154_c111 bl[111] br[111] wl[154] vdd gnd cell_6t
Xbit_r155_c111 bl[111] br[111] wl[155] vdd gnd cell_6t
Xbit_r156_c111 bl[111] br[111] wl[156] vdd gnd cell_6t
Xbit_r157_c111 bl[111] br[111] wl[157] vdd gnd cell_6t
Xbit_r158_c111 bl[111] br[111] wl[158] vdd gnd cell_6t
Xbit_r159_c111 bl[111] br[111] wl[159] vdd gnd cell_6t
Xbit_r160_c111 bl[111] br[111] wl[160] vdd gnd cell_6t
Xbit_r161_c111 bl[111] br[111] wl[161] vdd gnd cell_6t
Xbit_r162_c111 bl[111] br[111] wl[162] vdd gnd cell_6t
Xbit_r163_c111 bl[111] br[111] wl[163] vdd gnd cell_6t
Xbit_r164_c111 bl[111] br[111] wl[164] vdd gnd cell_6t
Xbit_r165_c111 bl[111] br[111] wl[165] vdd gnd cell_6t
Xbit_r166_c111 bl[111] br[111] wl[166] vdd gnd cell_6t
Xbit_r167_c111 bl[111] br[111] wl[167] vdd gnd cell_6t
Xbit_r168_c111 bl[111] br[111] wl[168] vdd gnd cell_6t
Xbit_r169_c111 bl[111] br[111] wl[169] vdd gnd cell_6t
Xbit_r170_c111 bl[111] br[111] wl[170] vdd gnd cell_6t
Xbit_r171_c111 bl[111] br[111] wl[171] vdd gnd cell_6t
Xbit_r172_c111 bl[111] br[111] wl[172] vdd gnd cell_6t
Xbit_r173_c111 bl[111] br[111] wl[173] vdd gnd cell_6t
Xbit_r174_c111 bl[111] br[111] wl[174] vdd gnd cell_6t
Xbit_r175_c111 bl[111] br[111] wl[175] vdd gnd cell_6t
Xbit_r176_c111 bl[111] br[111] wl[176] vdd gnd cell_6t
Xbit_r177_c111 bl[111] br[111] wl[177] vdd gnd cell_6t
Xbit_r178_c111 bl[111] br[111] wl[178] vdd gnd cell_6t
Xbit_r179_c111 bl[111] br[111] wl[179] vdd gnd cell_6t
Xbit_r180_c111 bl[111] br[111] wl[180] vdd gnd cell_6t
Xbit_r181_c111 bl[111] br[111] wl[181] vdd gnd cell_6t
Xbit_r182_c111 bl[111] br[111] wl[182] vdd gnd cell_6t
Xbit_r183_c111 bl[111] br[111] wl[183] vdd gnd cell_6t
Xbit_r184_c111 bl[111] br[111] wl[184] vdd gnd cell_6t
Xbit_r185_c111 bl[111] br[111] wl[185] vdd gnd cell_6t
Xbit_r186_c111 bl[111] br[111] wl[186] vdd gnd cell_6t
Xbit_r187_c111 bl[111] br[111] wl[187] vdd gnd cell_6t
Xbit_r188_c111 bl[111] br[111] wl[188] vdd gnd cell_6t
Xbit_r189_c111 bl[111] br[111] wl[189] vdd gnd cell_6t
Xbit_r190_c111 bl[111] br[111] wl[190] vdd gnd cell_6t
Xbit_r191_c111 bl[111] br[111] wl[191] vdd gnd cell_6t
Xbit_r192_c111 bl[111] br[111] wl[192] vdd gnd cell_6t
Xbit_r193_c111 bl[111] br[111] wl[193] vdd gnd cell_6t
Xbit_r194_c111 bl[111] br[111] wl[194] vdd gnd cell_6t
Xbit_r195_c111 bl[111] br[111] wl[195] vdd gnd cell_6t
Xbit_r196_c111 bl[111] br[111] wl[196] vdd gnd cell_6t
Xbit_r197_c111 bl[111] br[111] wl[197] vdd gnd cell_6t
Xbit_r198_c111 bl[111] br[111] wl[198] vdd gnd cell_6t
Xbit_r199_c111 bl[111] br[111] wl[199] vdd gnd cell_6t
Xbit_r200_c111 bl[111] br[111] wl[200] vdd gnd cell_6t
Xbit_r201_c111 bl[111] br[111] wl[201] vdd gnd cell_6t
Xbit_r202_c111 bl[111] br[111] wl[202] vdd gnd cell_6t
Xbit_r203_c111 bl[111] br[111] wl[203] vdd gnd cell_6t
Xbit_r204_c111 bl[111] br[111] wl[204] vdd gnd cell_6t
Xbit_r205_c111 bl[111] br[111] wl[205] vdd gnd cell_6t
Xbit_r206_c111 bl[111] br[111] wl[206] vdd gnd cell_6t
Xbit_r207_c111 bl[111] br[111] wl[207] vdd gnd cell_6t
Xbit_r208_c111 bl[111] br[111] wl[208] vdd gnd cell_6t
Xbit_r209_c111 bl[111] br[111] wl[209] vdd gnd cell_6t
Xbit_r210_c111 bl[111] br[111] wl[210] vdd gnd cell_6t
Xbit_r211_c111 bl[111] br[111] wl[211] vdd gnd cell_6t
Xbit_r212_c111 bl[111] br[111] wl[212] vdd gnd cell_6t
Xbit_r213_c111 bl[111] br[111] wl[213] vdd gnd cell_6t
Xbit_r214_c111 bl[111] br[111] wl[214] vdd gnd cell_6t
Xbit_r215_c111 bl[111] br[111] wl[215] vdd gnd cell_6t
Xbit_r216_c111 bl[111] br[111] wl[216] vdd gnd cell_6t
Xbit_r217_c111 bl[111] br[111] wl[217] vdd gnd cell_6t
Xbit_r218_c111 bl[111] br[111] wl[218] vdd gnd cell_6t
Xbit_r219_c111 bl[111] br[111] wl[219] vdd gnd cell_6t
Xbit_r220_c111 bl[111] br[111] wl[220] vdd gnd cell_6t
Xbit_r221_c111 bl[111] br[111] wl[221] vdd gnd cell_6t
Xbit_r222_c111 bl[111] br[111] wl[222] vdd gnd cell_6t
Xbit_r223_c111 bl[111] br[111] wl[223] vdd gnd cell_6t
Xbit_r224_c111 bl[111] br[111] wl[224] vdd gnd cell_6t
Xbit_r225_c111 bl[111] br[111] wl[225] vdd gnd cell_6t
Xbit_r226_c111 bl[111] br[111] wl[226] vdd gnd cell_6t
Xbit_r227_c111 bl[111] br[111] wl[227] vdd gnd cell_6t
Xbit_r228_c111 bl[111] br[111] wl[228] vdd gnd cell_6t
Xbit_r229_c111 bl[111] br[111] wl[229] vdd gnd cell_6t
Xbit_r230_c111 bl[111] br[111] wl[230] vdd gnd cell_6t
Xbit_r231_c111 bl[111] br[111] wl[231] vdd gnd cell_6t
Xbit_r232_c111 bl[111] br[111] wl[232] vdd gnd cell_6t
Xbit_r233_c111 bl[111] br[111] wl[233] vdd gnd cell_6t
Xbit_r234_c111 bl[111] br[111] wl[234] vdd gnd cell_6t
Xbit_r235_c111 bl[111] br[111] wl[235] vdd gnd cell_6t
Xbit_r236_c111 bl[111] br[111] wl[236] vdd gnd cell_6t
Xbit_r237_c111 bl[111] br[111] wl[237] vdd gnd cell_6t
Xbit_r238_c111 bl[111] br[111] wl[238] vdd gnd cell_6t
Xbit_r239_c111 bl[111] br[111] wl[239] vdd gnd cell_6t
Xbit_r240_c111 bl[111] br[111] wl[240] vdd gnd cell_6t
Xbit_r241_c111 bl[111] br[111] wl[241] vdd gnd cell_6t
Xbit_r242_c111 bl[111] br[111] wl[242] vdd gnd cell_6t
Xbit_r243_c111 bl[111] br[111] wl[243] vdd gnd cell_6t
Xbit_r244_c111 bl[111] br[111] wl[244] vdd gnd cell_6t
Xbit_r245_c111 bl[111] br[111] wl[245] vdd gnd cell_6t
Xbit_r246_c111 bl[111] br[111] wl[246] vdd gnd cell_6t
Xbit_r247_c111 bl[111] br[111] wl[247] vdd gnd cell_6t
Xbit_r248_c111 bl[111] br[111] wl[248] vdd gnd cell_6t
Xbit_r249_c111 bl[111] br[111] wl[249] vdd gnd cell_6t
Xbit_r250_c111 bl[111] br[111] wl[250] vdd gnd cell_6t
Xbit_r251_c111 bl[111] br[111] wl[251] vdd gnd cell_6t
Xbit_r252_c111 bl[111] br[111] wl[252] vdd gnd cell_6t
Xbit_r253_c111 bl[111] br[111] wl[253] vdd gnd cell_6t
Xbit_r254_c111 bl[111] br[111] wl[254] vdd gnd cell_6t
Xbit_r255_c111 bl[111] br[111] wl[255] vdd gnd cell_6t
Xbit_r256_c111 bl[111] br[111] wl[256] vdd gnd cell_6t
Xbit_r257_c111 bl[111] br[111] wl[257] vdd gnd cell_6t
Xbit_r258_c111 bl[111] br[111] wl[258] vdd gnd cell_6t
Xbit_r259_c111 bl[111] br[111] wl[259] vdd gnd cell_6t
Xbit_r260_c111 bl[111] br[111] wl[260] vdd gnd cell_6t
Xbit_r261_c111 bl[111] br[111] wl[261] vdd gnd cell_6t
Xbit_r262_c111 bl[111] br[111] wl[262] vdd gnd cell_6t
Xbit_r263_c111 bl[111] br[111] wl[263] vdd gnd cell_6t
Xbit_r264_c111 bl[111] br[111] wl[264] vdd gnd cell_6t
Xbit_r265_c111 bl[111] br[111] wl[265] vdd gnd cell_6t
Xbit_r266_c111 bl[111] br[111] wl[266] vdd gnd cell_6t
Xbit_r267_c111 bl[111] br[111] wl[267] vdd gnd cell_6t
Xbit_r268_c111 bl[111] br[111] wl[268] vdd gnd cell_6t
Xbit_r269_c111 bl[111] br[111] wl[269] vdd gnd cell_6t
Xbit_r270_c111 bl[111] br[111] wl[270] vdd gnd cell_6t
Xbit_r271_c111 bl[111] br[111] wl[271] vdd gnd cell_6t
Xbit_r272_c111 bl[111] br[111] wl[272] vdd gnd cell_6t
Xbit_r273_c111 bl[111] br[111] wl[273] vdd gnd cell_6t
Xbit_r274_c111 bl[111] br[111] wl[274] vdd gnd cell_6t
Xbit_r275_c111 bl[111] br[111] wl[275] vdd gnd cell_6t
Xbit_r276_c111 bl[111] br[111] wl[276] vdd gnd cell_6t
Xbit_r277_c111 bl[111] br[111] wl[277] vdd gnd cell_6t
Xbit_r278_c111 bl[111] br[111] wl[278] vdd gnd cell_6t
Xbit_r279_c111 bl[111] br[111] wl[279] vdd gnd cell_6t
Xbit_r280_c111 bl[111] br[111] wl[280] vdd gnd cell_6t
Xbit_r281_c111 bl[111] br[111] wl[281] vdd gnd cell_6t
Xbit_r282_c111 bl[111] br[111] wl[282] vdd gnd cell_6t
Xbit_r283_c111 bl[111] br[111] wl[283] vdd gnd cell_6t
Xbit_r284_c111 bl[111] br[111] wl[284] vdd gnd cell_6t
Xbit_r285_c111 bl[111] br[111] wl[285] vdd gnd cell_6t
Xbit_r286_c111 bl[111] br[111] wl[286] vdd gnd cell_6t
Xbit_r287_c111 bl[111] br[111] wl[287] vdd gnd cell_6t
Xbit_r288_c111 bl[111] br[111] wl[288] vdd gnd cell_6t
Xbit_r289_c111 bl[111] br[111] wl[289] vdd gnd cell_6t
Xbit_r290_c111 bl[111] br[111] wl[290] vdd gnd cell_6t
Xbit_r291_c111 bl[111] br[111] wl[291] vdd gnd cell_6t
Xbit_r292_c111 bl[111] br[111] wl[292] vdd gnd cell_6t
Xbit_r293_c111 bl[111] br[111] wl[293] vdd gnd cell_6t
Xbit_r294_c111 bl[111] br[111] wl[294] vdd gnd cell_6t
Xbit_r295_c111 bl[111] br[111] wl[295] vdd gnd cell_6t
Xbit_r296_c111 bl[111] br[111] wl[296] vdd gnd cell_6t
Xbit_r297_c111 bl[111] br[111] wl[297] vdd gnd cell_6t
Xbit_r298_c111 bl[111] br[111] wl[298] vdd gnd cell_6t
Xbit_r299_c111 bl[111] br[111] wl[299] vdd gnd cell_6t
Xbit_r300_c111 bl[111] br[111] wl[300] vdd gnd cell_6t
Xbit_r301_c111 bl[111] br[111] wl[301] vdd gnd cell_6t
Xbit_r302_c111 bl[111] br[111] wl[302] vdd gnd cell_6t
Xbit_r303_c111 bl[111] br[111] wl[303] vdd gnd cell_6t
Xbit_r304_c111 bl[111] br[111] wl[304] vdd gnd cell_6t
Xbit_r305_c111 bl[111] br[111] wl[305] vdd gnd cell_6t
Xbit_r306_c111 bl[111] br[111] wl[306] vdd gnd cell_6t
Xbit_r307_c111 bl[111] br[111] wl[307] vdd gnd cell_6t
Xbit_r308_c111 bl[111] br[111] wl[308] vdd gnd cell_6t
Xbit_r309_c111 bl[111] br[111] wl[309] vdd gnd cell_6t
Xbit_r310_c111 bl[111] br[111] wl[310] vdd gnd cell_6t
Xbit_r311_c111 bl[111] br[111] wl[311] vdd gnd cell_6t
Xbit_r312_c111 bl[111] br[111] wl[312] vdd gnd cell_6t
Xbit_r313_c111 bl[111] br[111] wl[313] vdd gnd cell_6t
Xbit_r314_c111 bl[111] br[111] wl[314] vdd gnd cell_6t
Xbit_r315_c111 bl[111] br[111] wl[315] vdd gnd cell_6t
Xbit_r316_c111 bl[111] br[111] wl[316] vdd gnd cell_6t
Xbit_r317_c111 bl[111] br[111] wl[317] vdd gnd cell_6t
Xbit_r318_c111 bl[111] br[111] wl[318] vdd gnd cell_6t
Xbit_r319_c111 bl[111] br[111] wl[319] vdd gnd cell_6t
Xbit_r320_c111 bl[111] br[111] wl[320] vdd gnd cell_6t
Xbit_r321_c111 bl[111] br[111] wl[321] vdd gnd cell_6t
Xbit_r322_c111 bl[111] br[111] wl[322] vdd gnd cell_6t
Xbit_r323_c111 bl[111] br[111] wl[323] vdd gnd cell_6t
Xbit_r324_c111 bl[111] br[111] wl[324] vdd gnd cell_6t
Xbit_r325_c111 bl[111] br[111] wl[325] vdd gnd cell_6t
Xbit_r326_c111 bl[111] br[111] wl[326] vdd gnd cell_6t
Xbit_r327_c111 bl[111] br[111] wl[327] vdd gnd cell_6t
Xbit_r328_c111 bl[111] br[111] wl[328] vdd gnd cell_6t
Xbit_r329_c111 bl[111] br[111] wl[329] vdd gnd cell_6t
Xbit_r330_c111 bl[111] br[111] wl[330] vdd gnd cell_6t
Xbit_r331_c111 bl[111] br[111] wl[331] vdd gnd cell_6t
Xbit_r332_c111 bl[111] br[111] wl[332] vdd gnd cell_6t
Xbit_r333_c111 bl[111] br[111] wl[333] vdd gnd cell_6t
Xbit_r334_c111 bl[111] br[111] wl[334] vdd gnd cell_6t
Xbit_r335_c111 bl[111] br[111] wl[335] vdd gnd cell_6t
Xbit_r336_c111 bl[111] br[111] wl[336] vdd gnd cell_6t
Xbit_r337_c111 bl[111] br[111] wl[337] vdd gnd cell_6t
Xbit_r338_c111 bl[111] br[111] wl[338] vdd gnd cell_6t
Xbit_r339_c111 bl[111] br[111] wl[339] vdd gnd cell_6t
Xbit_r340_c111 bl[111] br[111] wl[340] vdd gnd cell_6t
Xbit_r341_c111 bl[111] br[111] wl[341] vdd gnd cell_6t
Xbit_r342_c111 bl[111] br[111] wl[342] vdd gnd cell_6t
Xbit_r343_c111 bl[111] br[111] wl[343] vdd gnd cell_6t
Xbit_r344_c111 bl[111] br[111] wl[344] vdd gnd cell_6t
Xbit_r345_c111 bl[111] br[111] wl[345] vdd gnd cell_6t
Xbit_r346_c111 bl[111] br[111] wl[346] vdd gnd cell_6t
Xbit_r347_c111 bl[111] br[111] wl[347] vdd gnd cell_6t
Xbit_r348_c111 bl[111] br[111] wl[348] vdd gnd cell_6t
Xbit_r349_c111 bl[111] br[111] wl[349] vdd gnd cell_6t
Xbit_r350_c111 bl[111] br[111] wl[350] vdd gnd cell_6t
Xbit_r351_c111 bl[111] br[111] wl[351] vdd gnd cell_6t
Xbit_r352_c111 bl[111] br[111] wl[352] vdd gnd cell_6t
Xbit_r353_c111 bl[111] br[111] wl[353] vdd gnd cell_6t
Xbit_r354_c111 bl[111] br[111] wl[354] vdd gnd cell_6t
Xbit_r355_c111 bl[111] br[111] wl[355] vdd gnd cell_6t
Xbit_r356_c111 bl[111] br[111] wl[356] vdd gnd cell_6t
Xbit_r357_c111 bl[111] br[111] wl[357] vdd gnd cell_6t
Xbit_r358_c111 bl[111] br[111] wl[358] vdd gnd cell_6t
Xbit_r359_c111 bl[111] br[111] wl[359] vdd gnd cell_6t
Xbit_r360_c111 bl[111] br[111] wl[360] vdd gnd cell_6t
Xbit_r361_c111 bl[111] br[111] wl[361] vdd gnd cell_6t
Xbit_r362_c111 bl[111] br[111] wl[362] vdd gnd cell_6t
Xbit_r363_c111 bl[111] br[111] wl[363] vdd gnd cell_6t
Xbit_r364_c111 bl[111] br[111] wl[364] vdd gnd cell_6t
Xbit_r365_c111 bl[111] br[111] wl[365] vdd gnd cell_6t
Xbit_r366_c111 bl[111] br[111] wl[366] vdd gnd cell_6t
Xbit_r367_c111 bl[111] br[111] wl[367] vdd gnd cell_6t
Xbit_r368_c111 bl[111] br[111] wl[368] vdd gnd cell_6t
Xbit_r369_c111 bl[111] br[111] wl[369] vdd gnd cell_6t
Xbit_r370_c111 bl[111] br[111] wl[370] vdd gnd cell_6t
Xbit_r371_c111 bl[111] br[111] wl[371] vdd gnd cell_6t
Xbit_r372_c111 bl[111] br[111] wl[372] vdd gnd cell_6t
Xbit_r373_c111 bl[111] br[111] wl[373] vdd gnd cell_6t
Xbit_r374_c111 bl[111] br[111] wl[374] vdd gnd cell_6t
Xbit_r375_c111 bl[111] br[111] wl[375] vdd gnd cell_6t
Xbit_r376_c111 bl[111] br[111] wl[376] vdd gnd cell_6t
Xbit_r377_c111 bl[111] br[111] wl[377] vdd gnd cell_6t
Xbit_r378_c111 bl[111] br[111] wl[378] vdd gnd cell_6t
Xbit_r379_c111 bl[111] br[111] wl[379] vdd gnd cell_6t
Xbit_r380_c111 bl[111] br[111] wl[380] vdd gnd cell_6t
Xbit_r381_c111 bl[111] br[111] wl[381] vdd gnd cell_6t
Xbit_r382_c111 bl[111] br[111] wl[382] vdd gnd cell_6t
Xbit_r383_c111 bl[111] br[111] wl[383] vdd gnd cell_6t
Xbit_r384_c111 bl[111] br[111] wl[384] vdd gnd cell_6t
Xbit_r385_c111 bl[111] br[111] wl[385] vdd gnd cell_6t
Xbit_r386_c111 bl[111] br[111] wl[386] vdd gnd cell_6t
Xbit_r387_c111 bl[111] br[111] wl[387] vdd gnd cell_6t
Xbit_r388_c111 bl[111] br[111] wl[388] vdd gnd cell_6t
Xbit_r389_c111 bl[111] br[111] wl[389] vdd gnd cell_6t
Xbit_r390_c111 bl[111] br[111] wl[390] vdd gnd cell_6t
Xbit_r391_c111 bl[111] br[111] wl[391] vdd gnd cell_6t
Xbit_r392_c111 bl[111] br[111] wl[392] vdd gnd cell_6t
Xbit_r393_c111 bl[111] br[111] wl[393] vdd gnd cell_6t
Xbit_r394_c111 bl[111] br[111] wl[394] vdd gnd cell_6t
Xbit_r395_c111 bl[111] br[111] wl[395] vdd gnd cell_6t
Xbit_r396_c111 bl[111] br[111] wl[396] vdd gnd cell_6t
Xbit_r397_c111 bl[111] br[111] wl[397] vdd gnd cell_6t
Xbit_r398_c111 bl[111] br[111] wl[398] vdd gnd cell_6t
Xbit_r399_c111 bl[111] br[111] wl[399] vdd gnd cell_6t
Xbit_r400_c111 bl[111] br[111] wl[400] vdd gnd cell_6t
Xbit_r401_c111 bl[111] br[111] wl[401] vdd gnd cell_6t
Xbit_r402_c111 bl[111] br[111] wl[402] vdd gnd cell_6t
Xbit_r403_c111 bl[111] br[111] wl[403] vdd gnd cell_6t
Xbit_r404_c111 bl[111] br[111] wl[404] vdd gnd cell_6t
Xbit_r405_c111 bl[111] br[111] wl[405] vdd gnd cell_6t
Xbit_r406_c111 bl[111] br[111] wl[406] vdd gnd cell_6t
Xbit_r407_c111 bl[111] br[111] wl[407] vdd gnd cell_6t
Xbit_r408_c111 bl[111] br[111] wl[408] vdd gnd cell_6t
Xbit_r409_c111 bl[111] br[111] wl[409] vdd gnd cell_6t
Xbit_r410_c111 bl[111] br[111] wl[410] vdd gnd cell_6t
Xbit_r411_c111 bl[111] br[111] wl[411] vdd gnd cell_6t
Xbit_r412_c111 bl[111] br[111] wl[412] vdd gnd cell_6t
Xbit_r413_c111 bl[111] br[111] wl[413] vdd gnd cell_6t
Xbit_r414_c111 bl[111] br[111] wl[414] vdd gnd cell_6t
Xbit_r415_c111 bl[111] br[111] wl[415] vdd gnd cell_6t
Xbit_r416_c111 bl[111] br[111] wl[416] vdd gnd cell_6t
Xbit_r417_c111 bl[111] br[111] wl[417] vdd gnd cell_6t
Xbit_r418_c111 bl[111] br[111] wl[418] vdd gnd cell_6t
Xbit_r419_c111 bl[111] br[111] wl[419] vdd gnd cell_6t
Xbit_r420_c111 bl[111] br[111] wl[420] vdd gnd cell_6t
Xbit_r421_c111 bl[111] br[111] wl[421] vdd gnd cell_6t
Xbit_r422_c111 bl[111] br[111] wl[422] vdd gnd cell_6t
Xbit_r423_c111 bl[111] br[111] wl[423] vdd gnd cell_6t
Xbit_r424_c111 bl[111] br[111] wl[424] vdd gnd cell_6t
Xbit_r425_c111 bl[111] br[111] wl[425] vdd gnd cell_6t
Xbit_r426_c111 bl[111] br[111] wl[426] vdd gnd cell_6t
Xbit_r427_c111 bl[111] br[111] wl[427] vdd gnd cell_6t
Xbit_r428_c111 bl[111] br[111] wl[428] vdd gnd cell_6t
Xbit_r429_c111 bl[111] br[111] wl[429] vdd gnd cell_6t
Xbit_r430_c111 bl[111] br[111] wl[430] vdd gnd cell_6t
Xbit_r431_c111 bl[111] br[111] wl[431] vdd gnd cell_6t
Xbit_r432_c111 bl[111] br[111] wl[432] vdd gnd cell_6t
Xbit_r433_c111 bl[111] br[111] wl[433] vdd gnd cell_6t
Xbit_r434_c111 bl[111] br[111] wl[434] vdd gnd cell_6t
Xbit_r435_c111 bl[111] br[111] wl[435] vdd gnd cell_6t
Xbit_r436_c111 bl[111] br[111] wl[436] vdd gnd cell_6t
Xbit_r437_c111 bl[111] br[111] wl[437] vdd gnd cell_6t
Xbit_r438_c111 bl[111] br[111] wl[438] vdd gnd cell_6t
Xbit_r439_c111 bl[111] br[111] wl[439] vdd gnd cell_6t
Xbit_r440_c111 bl[111] br[111] wl[440] vdd gnd cell_6t
Xbit_r441_c111 bl[111] br[111] wl[441] vdd gnd cell_6t
Xbit_r442_c111 bl[111] br[111] wl[442] vdd gnd cell_6t
Xbit_r443_c111 bl[111] br[111] wl[443] vdd gnd cell_6t
Xbit_r444_c111 bl[111] br[111] wl[444] vdd gnd cell_6t
Xbit_r445_c111 bl[111] br[111] wl[445] vdd gnd cell_6t
Xbit_r446_c111 bl[111] br[111] wl[446] vdd gnd cell_6t
Xbit_r447_c111 bl[111] br[111] wl[447] vdd gnd cell_6t
Xbit_r448_c111 bl[111] br[111] wl[448] vdd gnd cell_6t
Xbit_r449_c111 bl[111] br[111] wl[449] vdd gnd cell_6t
Xbit_r450_c111 bl[111] br[111] wl[450] vdd gnd cell_6t
Xbit_r451_c111 bl[111] br[111] wl[451] vdd gnd cell_6t
Xbit_r452_c111 bl[111] br[111] wl[452] vdd gnd cell_6t
Xbit_r453_c111 bl[111] br[111] wl[453] vdd gnd cell_6t
Xbit_r454_c111 bl[111] br[111] wl[454] vdd gnd cell_6t
Xbit_r455_c111 bl[111] br[111] wl[455] vdd gnd cell_6t
Xbit_r456_c111 bl[111] br[111] wl[456] vdd gnd cell_6t
Xbit_r457_c111 bl[111] br[111] wl[457] vdd gnd cell_6t
Xbit_r458_c111 bl[111] br[111] wl[458] vdd gnd cell_6t
Xbit_r459_c111 bl[111] br[111] wl[459] vdd gnd cell_6t
Xbit_r460_c111 bl[111] br[111] wl[460] vdd gnd cell_6t
Xbit_r461_c111 bl[111] br[111] wl[461] vdd gnd cell_6t
Xbit_r462_c111 bl[111] br[111] wl[462] vdd gnd cell_6t
Xbit_r463_c111 bl[111] br[111] wl[463] vdd gnd cell_6t
Xbit_r464_c111 bl[111] br[111] wl[464] vdd gnd cell_6t
Xbit_r465_c111 bl[111] br[111] wl[465] vdd gnd cell_6t
Xbit_r466_c111 bl[111] br[111] wl[466] vdd gnd cell_6t
Xbit_r467_c111 bl[111] br[111] wl[467] vdd gnd cell_6t
Xbit_r468_c111 bl[111] br[111] wl[468] vdd gnd cell_6t
Xbit_r469_c111 bl[111] br[111] wl[469] vdd gnd cell_6t
Xbit_r470_c111 bl[111] br[111] wl[470] vdd gnd cell_6t
Xbit_r471_c111 bl[111] br[111] wl[471] vdd gnd cell_6t
Xbit_r472_c111 bl[111] br[111] wl[472] vdd gnd cell_6t
Xbit_r473_c111 bl[111] br[111] wl[473] vdd gnd cell_6t
Xbit_r474_c111 bl[111] br[111] wl[474] vdd gnd cell_6t
Xbit_r475_c111 bl[111] br[111] wl[475] vdd gnd cell_6t
Xbit_r476_c111 bl[111] br[111] wl[476] vdd gnd cell_6t
Xbit_r477_c111 bl[111] br[111] wl[477] vdd gnd cell_6t
Xbit_r478_c111 bl[111] br[111] wl[478] vdd gnd cell_6t
Xbit_r479_c111 bl[111] br[111] wl[479] vdd gnd cell_6t
Xbit_r480_c111 bl[111] br[111] wl[480] vdd gnd cell_6t
Xbit_r481_c111 bl[111] br[111] wl[481] vdd gnd cell_6t
Xbit_r482_c111 bl[111] br[111] wl[482] vdd gnd cell_6t
Xbit_r483_c111 bl[111] br[111] wl[483] vdd gnd cell_6t
Xbit_r484_c111 bl[111] br[111] wl[484] vdd gnd cell_6t
Xbit_r485_c111 bl[111] br[111] wl[485] vdd gnd cell_6t
Xbit_r486_c111 bl[111] br[111] wl[486] vdd gnd cell_6t
Xbit_r487_c111 bl[111] br[111] wl[487] vdd gnd cell_6t
Xbit_r488_c111 bl[111] br[111] wl[488] vdd gnd cell_6t
Xbit_r489_c111 bl[111] br[111] wl[489] vdd gnd cell_6t
Xbit_r490_c111 bl[111] br[111] wl[490] vdd gnd cell_6t
Xbit_r491_c111 bl[111] br[111] wl[491] vdd gnd cell_6t
Xbit_r492_c111 bl[111] br[111] wl[492] vdd gnd cell_6t
Xbit_r493_c111 bl[111] br[111] wl[493] vdd gnd cell_6t
Xbit_r494_c111 bl[111] br[111] wl[494] vdd gnd cell_6t
Xbit_r495_c111 bl[111] br[111] wl[495] vdd gnd cell_6t
Xbit_r496_c111 bl[111] br[111] wl[496] vdd gnd cell_6t
Xbit_r497_c111 bl[111] br[111] wl[497] vdd gnd cell_6t
Xbit_r498_c111 bl[111] br[111] wl[498] vdd gnd cell_6t
Xbit_r499_c111 bl[111] br[111] wl[499] vdd gnd cell_6t
Xbit_r500_c111 bl[111] br[111] wl[500] vdd gnd cell_6t
Xbit_r501_c111 bl[111] br[111] wl[501] vdd gnd cell_6t
Xbit_r502_c111 bl[111] br[111] wl[502] vdd gnd cell_6t
Xbit_r503_c111 bl[111] br[111] wl[503] vdd gnd cell_6t
Xbit_r504_c111 bl[111] br[111] wl[504] vdd gnd cell_6t
Xbit_r505_c111 bl[111] br[111] wl[505] vdd gnd cell_6t
Xbit_r506_c111 bl[111] br[111] wl[506] vdd gnd cell_6t
Xbit_r507_c111 bl[111] br[111] wl[507] vdd gnd cell_6t
Xbit_r508_c111 bl[111] br[111] wl[508] vdd gnd cell_6t
Xbit_r509_c111 bl[111] br[111] wl[509] vdd gnd cell_6t
Xbit_r510_c111 bl[111] br[111] wl[510] vdd gnd cell_6t
Xbit_r511_c111 bl[111] br[111] wl[511] vdd gnd cell_6t
Xbit_r0_c112 bl[112] br[112] wl[0] vdd gnd cell_6t
Xbit_r1_c112 bl[112] br[112] wl[1] vdd gnd cell_6t
Xbit_r2_c112 bl[112] br[112] wl[2] vdd gnd cell_6t
Xbit_r3_c112 bl[112] br[112] wl[3] vdd gnd cell_6t
Xbit_r4_c112 bl[112] br[112] wl[4] vdd gnd cell_6t
Xbit_r5_c112 bl[112] br[112] wl[5] vdd gnd cell_6t
Xbit_r6_c112 bl[112] br[112] wl[6] vdd gnd cell_6t
Xbit_r7_c112 bl[112] br[112] wl[7] vdd gnd cell_6t
Xbit_r8_c112 bl[112] br[112] wl[8] vdd gnd cell_6t
Xbit_r9_c112 bl[112] br[112] wl[9] vdd gnd cell_6t
Xbit_r10_c112 bl[112] br[112] wl[10] vdd gnd cell_6t
Xbit_r11_c112 bl[112] br[112] wl[11] vdd gnd cell_6t
Xbit_r12_c112 bl[112] br[112] wl[12] vdd gnd cell_6t
Xbit_r13_c112 bl[112] br[112] wl[13] vdd gnd cell_6t
Xbit_r14_c112 bl[112] br[112] wl[14] vdd gnd cell_6t
Xbit_r15_c112 bl[112] br[112] wl[15] vdd gnd cell_6t
Xbit_r16_c112 bl[112] br[112] wl[16] vdd gnd cell_6t
Xbit_r17_c112 bl[112] br[112] wl[17] vdd gnd cell_6t
Xbit_r18_c112 bl[112] br[112] wl[18] vdd gnd cell_6t
Xbit_r19_c112 bl[112] br[112] wl[19] vdd gnd cell_6t
Xbit_r20_c112 bl[112] br[112] wl[20] vdd gnd cell_6t
Xbit_r21_c112 bl[112] br[112] wl[21] vdd gnd cell_6t
Xbit_r22_c112 bl[112] br[112] wl[22] vdd gnd cell_6t
Xbit_r23_c112 bl[112] br[112] wl[23] vdd gnd cell_6t
Xbit_r24_c112 bl[112] br[112] wl[24] vdd gnd cell_6t
Xbit_r25_c112 bl[112] br[112] wl[25] vdd gnd cell_6t
Xbit_r26_c112 bl[112] br[112] wl[26] vdd gnd cell_6t
Xbit_r27_c112 bl[112] br[112] wl[27] vdd gnd cell_6t
Xbit_r28_c112 bl[112] br[112] wl[28] vdd gnd cell_6t
Xbit_r29_c112 bl[112] br[112] wl[29] vdd gnd cell_6t
Xbit_r30_c112 bl[112] br[112] wl[30] vdd gnd cell_6t
Xbit_r31_c112 bl[112] br[112] wl[31] vdd gnd cell_6t
Xbit_r32_c112 bl[112] br[112] wl[32] vdd gnd cell_6t
Xbit_r33_c112 bl[112] br[112] wl[33] vdd gnd cell_6t
Xbit_r34_c112 bl[112] br[112] wl[34] vdd gnd cell_6t
Xbit_r35_c112 bl[112] br[112] wl[35] vdd gnd cell_6t
Xbit_r36_c112 bl[112] br[112] wl[36] vdd gnd cell_6t
Xbit_r37_c112 bl[112] br[112] wl[37] vdd gnd cell_6t
Xbit_r38_c112 bl[112] br[112] wl[38] vdd gnd cell_6t
Xbit_r39_c112 bl[112] br[112] wl[39] vdd gnd cell_6t
Xbit_r40_c112 bl[112] br[112] wl[40] vdd gnd cell_6t
Xbit_r41_c112 bl[112] br[112] wl[41] vdd gnd cell_6t
Xbit_r42_c112 bl[112] br[112] wl[42] vdd gnd cell_6t
Xbit_r43_c112 bl[112] br[112] wl[43] vdd gnd cell_6t
Xbit_r44_c112 bl[112] br[112] wl[44] vdd gnd cell_6t
Xbit_r45_c112 bl[112] br[112] wl[45] vdd gnd cell_6t
Xbit_r46_c112 bl[112] br[112] wl[46] vdd gnd cell_6t
Xbit_r47_c112 bl[112] br[112] wl[47] vdd gnd cell_6t
Xbit_r48_c112 bl[112] br[112] wl[48] vdd gnd cell_6t
Xbit_r49_c112 bl[112] br[112] wl[49] vdd gnd cell_6t
Xbit_r50_c112 bl[112] br[112] wl[50] vdd gnd cell_6t
Xbit_r51_c112 bl[112] br[112] wl[51] vdd gnd cell_6t
Xbit_r52_c112 bl[112] br[112] wl[52] vdd gnd cell_6t
Xbit_r53_c112 bl[112] br[112] wl[53] vdd gnd cell_6t
Xbit_r54_c112 bl[112] br[112] wl[54] vdd gnd cell_6t
Xbit_r55_c112 bl[112] br[112] wl[55] vdd gnd cell_6t
Xbit_r56_c112 bl[112] br[112] wl[56] vdd gnd cell_6t
Xbit_r57_c112 bl[112] br[112] wl[57] vdd gnd cell_6t
Xbit_r58_c112 bl[112] br[112] wl[58] vdd gnd cell_6t
Xbit_r59_c112 bl[112] br[112] wl[59] vdd gnd cell_6t
Xbit_r60_c112 bl[112] br[112] wl[60] vdd gnd cell_6t
Xbit_r61_c112 bl[112] br[112] wl[61] vdd gnd cell_6t
Xbit_r62_c112 bl[112] br[112] wl[62] vdd gnd cell_6t
Xbit_r63_c112 bl[112] br[112] wl[63] vdd gnd cell_6t
Xbit_r64_c112 bl[112] br[112] wl[64] vdd gnd cell_6t
Xbit_r65_c112 bl[112] br[112] wl[65] vdd gnd cell_6t
Xbit_r66_c112 bl[112] br[112] wl[66] vdd gnd cell_6t
Xbit_r67_c112 bl[112] br[112] wl[67] vdd gnd cell_6t
Xbit_r68_c112 bl[112] br[112] wl[68] vdd gnd cell_6t
Xbit_r69_c112 bl[112] br[112] wl[69] vdd gnd cell_6t
Xbit_r70_c112 bl[112] br[112] wl[70] vdd gnd cell_6t
Xbit_r71_c112 bl[112] br[112] wl[71] vdd gnd cell_6t
Xbit_r72_c112 bl[112] br[112] wl[72] vdd gnd cell_6t
Xbit_r73_c112 bl[112] br[112] wl[73] vdd gnd cell_6t
Xbit_r74_c112 bl[112] br[112] wl[74] vdd gnd cell_6t
Xbit_r75_c112 bl[112] br[112] wl[75] vdd gnd cell_6t
Xbit_r76_c112 bl[112] br[112] wl[76] vdd gnd cell_6t
Xbit_r77_c112 bl[112] br[112] wl[77] vdd gnd cell_6t
Xbit_r78_c112 bl[112] br[112] wl[78] vdd gnd cell_6t
Xbit_r79_c112 bl[112] br[112] wl[79] vdd gnd cell_6t
Xbit_r80_c112 bl[112] br[112] wl[80] vdd gnd cell_6t
Xbit_r81_c112 bl[112] br[112] wl[81] vdd gnd cell_6t
Xbit_r82_c112 bl[112] br[112] wl[82] vdd gnd cell_6t
Xbit_r83_c112 bl[112] br[112] wl[83] vdd gnd cell_6t
Xbit_r84_c112 bl[112] br[112] wl[84] vdd gnd cell_6t
Xbit_r85_c112 bl[112] br[112] wl[85] vdd gnd cell_6t
Xbit_r86_c112 bl[112] br[112] wl[86] vdd gnd cell_6t
Xbit_r87_c112 bl[112] br[112] wl[87] vdd gnd cell_6t
Xbit_r88_c112 bl[112] br[112] wl[88] vdd gnd cell_6t
Xbit_r89_c112 bl[112] br[112] wl[89] vdd gnd cell_6t
Xbit_r90_c112 bl[112] br[112] wl[90] vdd gnd cell_6t
Xbit_r91_c112 bl[112] br[112] wl[91] vdd gnd cell_6t
Xbit_r92_c112 bl[112] br[112] wl[92] vdd gnd cell_6t
Xbit_r93_c112 bl[112] br[112] wl[93] vdd gnd cell_6t
Xbit_r94_c112 bl[112] br[112] wl[94] vdd gnd cell_6t
Xbit_r95_c112 bl[112] br[112] wl[95] vdd gnd cell_6t
Xbit_r96_c112 bl[112] br[112] wl[96] vdd gnd cell_6t
Xbit_r97_c112 bl[112] br[112] wl[97] vdd gnd cell_6t
Xbit_r98_c112 bl[112] br[112] wl[98] vdd gnd cell_6t
Xbit_r99_c112 bl[112] br[112] wl[99] vdd gnd cell_6t
Xbit_r100_c112 bl[112] br[112] wl[100] vdd gnd cell_6t
Xbit_r101_c112 bl[112] br[112] wl[101] vdd gnd cell_6t
Xbit_r102_c112 bl[112] br[112] wl[102] vdd gnd cell_6t
Xbit_r103_c112 bl[112] br[112] wl[103] vdd gnd cell_6t
Xbit_r104_c112 bl[112] br[112] wl[104] vdd gnd cell_6t
Xbit_r105_c112 bl[112] br[112] wl[105] vdd gnd cell_6t
Xbit_r106_c112 bl[112] br[112] wl[106] vdd gnd cell_6t
Xbit_r107_c112 bl[112] br[112] wl[107] vdd gnd cell_6t
Xbit_r108_c112 bl[112] br[112] wl[108] vdd gnd cell_6t
Xbit_r109_c112 bl[112] br[112] wl[109] vdd gnd cell_6t
Xbit_r110_c112 bl[112] br[112] wl[110] vdd gnd cell_6t
Xbit_r111_c112 bl[112] br[112] wl[111] vdd gnd cell_6t
Xbit_r112_c112 bl[112] br[112] wl[112] vdd gnd cell_6t
Xbit_r113_c112 bl[112] br[112] wl[113] vdd gnd cell_6t
Xbit_r114_c112 bl[112] br[112] wl[114] vdd gnd cell_6t
Xbit_r115_c112 bl[112] br[112] wl[115] vdd gnd cell_6t
Xbit_r116_c112 bl[112] br[112] wl[116] vdd gnd cell_6t
Xbit_r117_c112 bl[112] br[112] wl[117] vdd gnd cell_6t
Xbit_r118_c112 bl[112] br[112] wl[118] vdd gnd cell_6t
Xbit_r119_c112 bl[112] br[112] wl[119] vdd gnd cell_6t
Xbit_r120_c112 bl[112] br[112] wl[120] vdd gnd cell_6t
Xbit_r121_c112 bl[112] br[112] wl[121] vdd gnd cell_6t
Xbit_r122_c112 bl[112] br[112] wl[122] vdd gnd cell_6t
Xbit_r123_c112 bl[112] br[112] wl[123] vdd gnd cell_6t
Xbit_r124_c112 bl[112] br[112] wl[124] vdd gnd cell_6t
Xbit_r125_c112 bl[112] br[112] wl[125] vdd gnd cell_6t
Xbit_r126_c112 bl[112] br[112] wl[126] vdd gnd cell_6t
Xbit_r127_c112 bl[112] br[112] wl[127] vdd gnd cell_6t
Xbit_r128_c112 bl[112] br[112] wl[128] vdd gnd cell_6t
Xbit_r129_c112 bl[112] br[112] wl[129] vdd gnd cell_6t
Xbit_r130_c112 bl[112] br[112] wl[130] vdd gnd cell_6t
Xbit_r131_c112 bl[112] br[112] wl[131] vdd gnd cell_6t
Xbit_r132_c112 bl[112] br[112] wl[132] vdd gnd cell_6t
Xbit_r133_c112 bl[112] br[112] wl[133] vdd gnd cell_6t
Xbit_r134_c112 bl[112] br[112] wl[134] vdd gnd cell_6t
Xbit_r135_c112 bl[112] br[112] wl[135] vdd gnd cell_6t
Xbit_r136_c112 bl[112] br[112] wl[136] vdd gnd cell_6t
Xbit_r137_c112 bl[112] br[112] wl[137] vdd gnd cell_6t
Xbit_r138_c112 bl[112] br[112] wl[138] vdd gnd cell_6t
Xbit_r139_c112 bl[112] br[112] wl[139] vdd gnd cell_6t
Xbit_r140_c112 bl[112] br[112] wl[140] vdd gnd cell_6t
Xbit_r141_c112 bl[112] br[112] wl[141] vdd gnd cell_6t
Xbit_r142_c112 bl[112] br[112] wl[142] vdd gnd cell_6t
Xbit_r143_c112 bl[112] br[112] wl[143] vdd gnd cell_6t
Xbit_r144_c112 bl[112] br[112] wl[144] vdd gnd cell_6t
Xbit_r145_c112 bl[112] br[112] wl[145] vdd gnd cell_6t
Xbit_r146_c112 bl[112] br[112] wl[146] vdd gnd cell_6t
Xbit_r147_c112 bl[112] br[112] wl[147] vdd gnd cell_6t
Xbit_r148_c112 bl[112] br[112] wl[148] vdd gnd cell_6t
Xbit_r149_c112 bl[112] br[112] wl[149] vdd gnd cell_6t
Xbit_r150_c112 bl[112] br[112] wl[150] vdd gnd cell_6t
Xbit_r151_c112 bl[112] br[112] wl[151] vdd gnd cell_6t
Xbit_r152_c112 bl[112] br[112] wl[152] vdd gnd cell_6t
Xbit_r153_c112 bl[112] br[112] wl[153] vdd gnd cell_6t
Xbit_r154_c112 bl[112] br[112] wl[154] vdd gnd cell_6t
Xbit_r155_c112 bl[112] br[112] wl[155] vdd gnd cell_6t
Xbit_r156_c112 bl[112] br[112] wl[156] vdd gnd cell_6t
Xbit_r157_c112 bl[112] br[112] wl[157] vdd gnd cell_6t
Xbit_r158_c112 bl[112] br[112] wl[158] vdd gnd cell_6t
Xbit_r159_c112 bl[112] br[112] wl[159] vdd gnd cell_6t
Xbit_r160_c112 bl[112] br[112] wl[160] vdd gnd cell_6t
Xbit_r161_c112 bl[112] br[112] wl[161] vdd gnd cell_6t
Xbit_r162_c112 bl[112] br[112] wl[162] vdd gnd cell_6t
Xbit_r163_c112 bl[112] br[112] wl[163] vdd gnd cell_6t
Xbit_r164_c112 bl[112] br[112] wl[164] vdd gnd cell_6t
Xbit_r165_c112 bl[112] br[112] wl[165] vdd gnd cell_6t
Xbit_r166_c112 bl[112] br[112] wl[166] vdd gnd cell_6t
Xbit_r167_c112 bl[112] br[112] wl[167] vdd gnd cell_6t
Xbit_r168_c112 bl[112] br[112] wl[168] vdd gnd cell_6t
Xbit_r169_c112 bl[112] br[112] wl[169] vdd gnd cell_6t
Xbit_r170_c112 bl[112] br[112] wl[170] vdd gnd cell_6t
Xbit_r171_c112 bl[112] br[112] wl[171] vdd gnd cell_6t
Xbit_r172_c112 bl[112] br[112] wl[172] vdd gnd cell_6t
Xbit_r173_c112 bl[112] br[112] wl[173] vdd gnd cell_6t
Xbit_r174_c112 bl[112] br[112] wl[174] vdd gnd cell_6t
Xbit_r175_c112 bl[112] br[112] wl[175] vdd gnd cell_6t
Xbit_r176_c112 bl[112] br[112] wl[176] vdd gnd cell_6t
Xbit_r177_c112 bl[112] br[112] wl[177] vdd gnd cell_6t
Xbit_r178_c112 bl[112] br[112] wl[178] vdd gnd cell_6t
Xbit_r179_c112 bl[112] br[112] wl[179] vdd gnd cell_6t
Xbit_r180_c112 bl[112] br[112] wl[180] vdd gnd cell_6t
Xbit_r181_c112 bl[112] br[112] wl[181] vdd gnd cell_6t
Xbit_r182_c112 bl[112] br[112] wl[182] vdd gnd cell_6t
Xbit_r183_c112 bl[112] br[112] wl[183] vdd gnd cell_6t
Xbit_r184_c112 bl[112] br[112] wl[184] vdd gnd cell_6t
Xbit_r185_c112 bl[112] br[112] wl[185] vdd gnd cell_6t
Xbit_r186_c112 bl[112] br[112] wl[186] vdd gnd cell_6t
Xbit_r187_c112 bl[112] br[112] wl[187] vdd gnd cell_6t
Xbit_r188_c112 bl[112] br[112] wl[188] vdd gnd cell_6t
Xbit_r189_c112 bl[112] br[112] wl[189] vdd gnd cell_6t
Xbit_r190_c112 bl[112] br[112] wl[190] vdd gnd cell_6t
Xbit_r191_c112 bl[112] br[112] wl[191] vdd gnd cell_6t
Xbit_r192_c112 bl[112] br[112] wl[192] vdd gnd cell_6t
Xbit_r193_c112 bl[112] br[112] wl[193] vdd gnd cell_6t
Xbit_r194_c112 bl[112] br[112] wl[194] vdd gnd cell_6t
Xbit_r195_c112 bl[112] br[112] wl[195] vdd gnd cell_6t
Xbit_r196_c112 bl[112] br[112] wl[196] vdd gnd cell_6t
Xbit_r197_c112 bl[112] br[112] wl[197] vdd gnd cell_6t
Xbit_r198_c112 bl[112] br[112] wl[198] vdd gnd cell_6t
Xbit_r199_c112 bl[112] br[112] wl[199] vdd gnd cell_6t
Xbit_r200_c112 bl[112] br[112] wl[200] vdd gnd cell_6t
Xbit_r201_c112 bl[112] br[112] wl[201] vdd gnd cell_6t
Xbit_r202_c112 bl[112] br[112] wl[202] vdd gnd cell_6t
Xbit_r203_c112 bl[112] br[112] wl[203] vdd gnd cell_6t
Xbit_r204_c112 bl[112] br[112] wl[204] vdd gnd cell_6t
Xbit_r205_c112 bl[112] br[112] wl[205] vdd gnd cell_6t
Xbit_r206_c112 bl[112] br[112] wl[206] vdd gnd cell_6t
Xbit_r207_c112 bl[112] br[112] wl[207] vdd gnd cell_6t
Xbit_r208_c112 bl[112] br[112] wl[208] vdd gnd cell_6t
Xbit_r209_c112 bl[112] br[112] wl[209] vdd gnd cell_6t
Xbit_r210_c112 bl[112] br[112] wl[210] vdd gnd cell_6t
Xbit_r211_c112 bl[112] br[112] wl[211] vdd gnd cell_6t
Xbit_r212_c112 bl[112] br[112] wl[212] vdd gnd cell_6t
Xbit_r213_c112 bl[112] br[112] wl[213] vdd gnd cell_6t
Xbit_r214_c112 bl[112] br[112] wl[214] vdd gnd cell_6t
Xbit_r215_c112 bl[112] br[112] wl[215] vdd gnd cell_6t
Xbit_r216_c112 bl[112] br[112] wl[216] vdd gnd cell_6t
Xbit_r217_c112 bl[112] br[112] wl[217] vdd gnd cell_6t
Xbit_r218_c112 bl[112] br[112] wl[218] vdd gnd cell_6t
Xbit_r219_c112 bl[112] br[112] wl[219] vdd gnd cell_6t
Xbit_r220_c112 bl[112] br[112] wl[220] vdd gnd cell_6t
Xbit_r221_c112 bl[112] br[112] wl[221] vdd gnd cell_6t
Xbit_r222_c112 bl[112] br[112] wl[222] vdd gnd cell_6t
Xbit_r223_c112 bl[112] br[112] wl[223] vdd gnd cell_6t
Xbit_r224_c112 bl[112] br[112] wl[224] vdd gnd cell_6t
Xbit_r225_c112 bl[112] br[112] wl[225] vdd gnd cell_6t
Xbit_r226_c112 bl[112] br[112] wl[226] vdd gnd cell_6t
Xbit_r227_c112 bl[112] br[112] wl[227] vdd gnd cell_6t
Xbit_r228_c112 bl[112] br[112] wl[228] vdd gnd cell_6t
Xbit_r229_c112 bl[112] br[112] wl[229] vdd gnd cell_6t
Xbit_r230_c112 bl[112] br[112] wl[230] vdd gnd cell_6t
Xbit_r231_c112 bl[112] br[112] wl[231] vdd gnd cell_6t
Xbit_r232_c112 bl[112] br[112] wl[232] vdd gnd cell_6t
Xbit_r233_c112 bl[112] br[112] wl[233] vdd gnd cell_6t
Xbit_r234_c112 bl[112] br[112] wl[234] vdd gnd cell_6t
Xbit_r235_c112 bl[112] br[112] wl[235] vdd gnd cell_6t
Xbit_r236_c112 bl[112] br[112] wl[236] vdd gnd cell_6t
Xbit_r237_c112 bl[112] br[112] wl[237] vdd gnd cell_6t
Xbit_r238_c112 bl[112] br[112] wl[238] vdd gnd cell_6t
Xbit_r239_c112 bl[112] br[112] wl[239] vdd gnd cell_6t
Xbit_r240_c112 bl[112] br[112] wl[240] vdd gnd cell_6t
Xbit_r241_c112 bl[112] br[112] wl[241] vdd gnd cell_6t
Xbit_r242_c112 bl[112] br[112] wl[242] vdd gnd cell_6t
Xbit_r243_c112 bl[112] br[112] wl[243] vdd gnd cell_6t
Xbit_r244_c112 bl[112] br[112] wl[244] vdd gnd cell_6t
Xbit_r245_c112 bl[112] br[112] wl[245] vdd gnd cell_6t
Xbit_r246_c112 bl[112] br[112] wl[246] vdd gnd cell_6t
Xbit_r247_c112 bl[112] br[112] wl[247] vdd gnd cell_6t
Xbit_r248_c112 bl[112] br[112] wl[248] vdd gnd cell_6t
Xbit_r249_c112 bl[112] br[112] wl[249] vdd gnd cell_6t
Xbit_r250_c112 bl[112] br[112] wl[250] vdd gnd cell_6t
Xbit_r251_c112 bl[112] br[112] wl[251] vdd gnd cell_6t
Xbit_r252_c112 bl[112] br[112] wl[252] vdd gnd cell_6t
Xbit_r253_c112 bl[112] br[112] wl[253] vdd gnd cell_6t
Xbit_r254_c112 bl[112] br[112] wl[254] vdd gnd cell_6t
Xbit_r255_c112 bl[112] br[112] wl[255] vdd gnd cell_6t
Xbit_r256_c112 bl[112] br[112] wl[256] vdd gnd cell_6t
Xbit_r257_c112 bl[112] br[112] wl[257] vdd gnd cell_6t
Xbit_r258_c112 bl[112] br[112] wl[258] vdd gnd cell_6t
Xbit_r259_c112 bl[112] br[112] wl[259] vdd gnd cell_6t
Xbit_r260_c112 bl[112] br[112] wl[260] vdd gnd cell_6t
Xbit_r261_c112 bl[112] br[112] wl[261] vdd gnd cell_6t
Xbit_r262_c112 bl[112] br[112] wl[262] vdd gnd cell_6t
Xbit_r263_c112 bl[112] br[112] wl[263] vdd gnd cell_6t
Xbit_r264_c112 bl[112] br[112] wl[264] vdd gnd cell_6t
Xbit_r265_c112 bl[112] br[112] wl[265] vdd gnd cell_6t
Xbit_r266_c112 bl[112] br[112] wl[266] vdd gnd cell_6t
Xbit_r267_c112 bl[112] br[112] wl[267] vdd gnd cell_6t
Xbit_r268_c112 bl[112] br[112] wl[268] vdd gnd cell_6t
Xbit_r269_c112 bl[112] br[112] wl[269] vdd gnd cell_6t
Xbit_r270_c112 bl[112] br[112] wl[270] vdd gnd cell_6t
Xbit_r271_c112 bl[112] br[112] wl[271] vdd gnd cell_6t
Xbit_r272_c112 bl[112] br[112] wl[272] vdd gnd cell_6t
Xbit_r273_c112 bl[112] br[112] wl[273] vdd gnd cell_6t
Xbit_r274_c112 bl[112] br[112] wl[274] vdd gnd cell_6t
Xbit_r275_c112 bl[112] br[112] wl[275] vdd gnd cell_6t
Xbit_r276_c112 bl[112] br[112] wl[276] vdd gnd cell_6t
Xbit_r277_c112 bl[112] br[112] wl[277] vdd gnd cell_6t
Xbit_r278_c112 bl[112] br[112] wl[278] vdd gnd cell_6t
Xbit_r279_c112 bl[112] br[112] wl[279] vdd gnd cell_6t
Xbit_r280_c112 bl[112] br[112] wl[280] vdd gnd cell_6t
Xbit_r281_c112 bl[112] br[112] wl[281] vdd gnd cell_6t
Xbit_r282_c112 bl[112] br[112] wl[282] vdd gnd cell_6t
Xbit_r283_c112 bl[112] br[112] wl[283] vdd gnd cell_6t
Xbit_r284_c112 bl[112] br[112] wl[284] vdd gnd cell_6t
Xbit_r285_c112 bl[112] br[112] wl[285] vdd gnd cell_6t
Xbit_r286_c112 bl[112] br[112] wl[286] vdd gnd cell_6t
Xbit_r287_c112 bl[112] br[112] wl[287] vdd gnd cell_6t
Xbit_r288_c112 bl[112] br[112] wl[288] vdd gnd cell_6t
Xbit_r289_c112 bl[112] br[112] wl[289] vdd gnd cell_6t
Xbit_r290_c112 bl[112] br[112] wl[290] vdd gnd cell_6t
Xbit_r291_c112 bl[112] br[112] wl[291] vdd gnd cell_6t
Xbit_r292_c112 bl[112] br[112] wl[292] vdd gnd cell_6t
Xbit_r293_c112 bl[112] br[112] wl[293] vdd gnd cell_6t
Xbit_r294_c112 bl[112] br[112] wl[294] vdd gnd cell_6t
Xbit_r295_c112 bl[112] br[112] wl[295] vdd gnd cell_6t
Xbit_r296_c112 bl[112] br[112] wl[296] vdd gnd cell_6t
Xbit_r297_c112 bl[112] br[112] wl[297] vdd gnd cell_6t
Xbit_r298_c112 bl[112] br[112] wl[298] vdd gnd cell_6t
Xbit_r299_c112 bl[112] br[112] wl[299] vdd gnd cell_6t
Xbit_r300_c112 bl[112] br[112] wl[300] vdd gnd cell_6t
Xbit_r301_c112 bl[112] br[112] wl[301] vdd gnd cell_6t
Xbit_r302_c112 bl[112] br[112] wl[302] vdd gnd cell_6t
Xbit_r303_c112 bl[112] br[112] wl[303] vdd gnd cell_6t
Xbit_r304_c112 bl[112] br[112] wl[304] vdd gnd cell_6t
Xbit_r305_c112 bl[112] br[112] wl[305] vdd gnd cell_6t
Xbit_r306_c112 bl[112] br[112] wl[306] vdd gnd cell_6t
Xbit_r307_c112 bl[112] br[112] wl[307] vdd gnd cell_6t
Xbit_r308_c112 bl[112] br[112] wl[308] vdd gnd cell_6t
Xbit_r309_c112 bl[112] br[112] wl[309] vdd gnd cell_6t
Xbit_r310_c112 bl[112] br[112] wl[310] vdd gnd cell_6t
Xbit_r311_c112 bl[112] br[112] wl[311] vdd gnd cell_6t
Xbit_r312_c112 bl[112] br[112] wl[312] vdd gnd cell_6t
Xbit_r313_c112 bl[112] br[112] wl[313] vdd gnd cell_6t
Xbit_r314_c112 bl[112] br[112] wl[314] vdd gnd cell_6t
Xbit_r315_c112 bl[112] br[112] wl[315] vdd gnd cell_6t
Xbit_r316_c112 bl[112] br[112] wl[316] vdd gnd cell_6t
Xbit_r317_c112 bl[112] br[112] wl[317] vdd gnd cell_6t
Xbit_r318_c112 bl[112] br[112] wl[318] vdd gnd cell_6t
Xbit_r319_c112 bl[112] br[112] wl[319] vdd gnd cell_6t
Xbit_r320_c112 bl[112] br[112] wl[320] vdd gnd cell_6t
Xbit_r321_c112 bl[112] br[112] wl[321] vdd gnd cell_6t
Xbit_r322_c112 bl[112] br[112] wl[322] vdd gnd cell_6t
Xbit_r323_c112 bl[112] br[112] wl[323] vdd gnd cell_6t
Xbit_r324_c112 bl[112] br[112] wl[324] vdd gnd cell_6t
Xbit_r325_c112 bl[112] br[112] wl[325] vdd gnd cell_6t
Xbit_r326_c112 bl[112] br[112] wl[326] vdd gnd cell_6t
Xbit_r327_c112 bl[112] br[112] wl[327] vdd gnd cell_6t
Xbit_r328_c112 bl[112] br[112] wl[328] vdd gnd cell_6t
Xbit_r329_c112 bl[112] br[112] wl[329] vdd gnd cell_6t
Xbit_r330_c112 bl[112] br[112] wl[330] vdd gnd cell_6t
Xbit_r331_c112 bl[112] br[112] wl[331] vdd gnd cell_6t
Xbit_r332_c112 bl[112] br[112] wl[332] vdd gnd cell_6t
Xbit_r333_c112 bl[112] br[112] wl[333] vdd gnd cell_6t
Xbit_r334_c112 bl[112] br[112] wl[334] vdd gnd cell_6t
Xbit_r335_c112 bl[112] br[112] wl[335] vdd gnd cell_6t
Xbit_r336_c112 bl[112] br[112] wl[336] vdd gnd cell_6t
Xbit_r337_c112 bl[112] br[112] wl[337] vdd gnd cell_6t
Xbit_r338_c112 bl[112] br[112] wl[338] vdd gnd cell_6t
Xbit_r339_c112 bl[112] br[112] wl[339] vdd gnd cell_6t
Xbit_r340_c112 bl[112] br[112] wl[340] vdd gnd cell_6t
Xbit_r341_c112 bl[112] br[112] wl[341] vdd gnd cell_6t
Xbit_r342_c112 bl[112] br[112] wl[342] vdd gnd cell_6t
Xbit_r343_c112 bl[112] br[112] wl[343] vdd gnd cell_6t
Xbit_r344_c112 bl[112] br[112] wl[344] vdd gnd cell_6t
Xbit_r345_c112 bl[112] br[112] wl[345] vdd gnd cell_6t
Xbit_r346_c112 bl[112] br[112] wl[346] vdd gnd cell_6t
Xbit_r347_c112 bl[112] br[112] wl[347] vdd gnd cell_6t
Xbit_r348_c112 bl[112] br[112] wl[348] vdd gnd cell_6t
Xbit_r349_c112 bl[112] br[112] wl[349] vdd gnd cell_6t
Xbit_r350_c112 bl[112] br[112] wl[350] vdd gnd cell_6t
Xbit_r351_c112 bl[112] br[112] wl[351] vdd gnd cell_6t
Xbit_r352_c112 bl[112] br[112] wl[352] vdd gnd cell_6t
Xbit_r353_c112 bl[112] br[112] wl[353] vdd gnd cell_6t
Xbit_r354_c112 bl[112] br[112] wl[354] vdd gnd cell_6t
Xbit_r355_c112 bl[112] br[112] wl[355] vdd gnd cell_6t
Xbit_r356_c112 bl[112] br[112] wl[356] vdd gnd cell_6t
Xbit_r357_c112 bl[112] br[112] wl[357] vdd gnd cell_6t
Xbit_r358_c112 bl[112] br[112] wl[358] vdd gnd cell_6t
Xbit_r359_c112 bl[112] br[112] wl[359] vdd gnd cell_6t
Xbit_r360_c112 bl[112] br[112] wl[360] vdd gnd cell_6t
Xbit_r361_c112 bl[112] br[112] wl[361] vdd gnd cell_6t
Xbit_r362_c112 bl[112] br[112] wl[362] vdd gnd cell_6t
Xbit_r363_c112 bl[112] br[112] wl[363] vdd gnd cell_6t
Xbit_r364_c112 bl[112] br[112] wl[364] vdd gnd cell_6t
Xbit_r365_c112 bl[112] br[112] wl[365] vdd gnd cell_6t
Xbit_r366_c112 bl[112] br[112] wl[366] vdd gnd cell_6t
Xbit_r367_c112 bl[112] br[112] wl[367] vdd gnd cell_6t
Xbit_r368_c112 bl[112] br[112] wl[368] vdd gnd cell_6t
Xbit_r369_c112 bl[112] br[112] wl[369] vdd gnd cell_6t
Xbit_r370_c112 bl[112] br[112] wl[370] vdd gnd cell_6t
Xbit_r371_c112 bl[112] br[112] wl[371] vdd gnd cell_6t
Xbit_r372_c112 bl[112] br[112] wl[372] vdd gnd cell_6t
Xbit_r373_c112 bl[112] br[112] wl[373] vdd gnd cell_6t
Xbit_r374_c112 bl[112] br[112] wl[374] vdd gnd cell_6t
Xbit_r375_c112 bl[112] br[112] wl[375] vdd gnd cell_6t
Xbit_r376_c112 bl[112] br[112] wl[376] vdd gnd cell_6t
Xbit_r377_c112 bl[112] br[112] wl[377] vdd gnd cell_6t
Xbit_r378_c112 bl[112] br[112] wl[378] vdd gnd cell_6t
Xbit_r379_c112 bl[112] br[112] wl[379] vdd gnd cell_6t
Xbit_r380_c112 bl[112] br[112] wl[380] vdd gnd cell_6t
Xbit_r381_c112 bl[112] br[112] wl[381] vdd gnd cell_6t
Xbit_r382_c112 bl[112] br[112] wl[382] vdd gnd cell_6t
Xbit_r383_c112 bl[112] br[112] wl[383] vdd gnd cell_6t
Xbit_r384_c112 bl[112] br[112] wl[384] vdd gnd cell_6t
Xbit_r385_c112 bl[112] br[112] wl[385] vdd gnd cell_6t
Xbit_r386_c112 bl[112] br[112] wl[386] vdd gnd cell_6t
Xbit_r387_c112 bl[112] br[112] wl[387] vdd gnd cell_6t
Xbit_r388_c112 bl[112] br[112] wl[388] vdd gnd cell_6t
Xbit_r389_c112 bl[112] br[112] wl[389] vdd gnd cell_6t
Xbit_r390_c112 bl[112] br[112] wl[390] vdd gnd cell_6t
Xbit_r391_c112 bl[112] br[112] wl[391] vdd gnd cell_6t
Xbit_r392_c112 bl[112] br[112] wl[392] vdd gnd cell_6t
Xbit_r393_c112 bl[112] br[112] wl[393] vdd gnd cell_6t
Xbit_r394_c112 bl[112] br[112] wl[394] vdd gnd cell_6t
Xbit_r395_c112 bl[112] br[112] wl[395] vdd gnd cell_6t
Xbit_r396_c112 bl[112] br[112] wl[396] vdd gnd cell_6t
Xbit_r397_c112 bl[112] br[112] wl[397] vdd gnd cell_6t
Xbit_r398_c112 bl[112] br[112] wl[398] vdd gnd cell_6t
Xbit_r399_c112 bl[112] br[112] wl[399] vdd gnd cell_6t
Xbit_r400_c112 bl[112] br[112] wl[400] vdd gnd cell_6t
Xbit_r401_c112 bl[112] br[112] wl[401] vdd gnd cell_6t
Xbit_r402_c112 bl[112] br[112] wl[402] vdd gnd cell_6t
Xbit_r403_c112 bl[112] br[112] wl[403] vdd gnd cell_6t
Xbit_r404_c112 bl[112] br[112] wl[404] vdd gnd cell_6t
Xbit_r405_c112 bl[112] br[112] wl[405] vdd gnd cell_6t
Xbit_r406_c112 bl[112] br[112] wl[406] vdd gnd cell_6t
Xbit_r407_c112 bl[112] br[112] wl[407] vdd gnd cell_6t
Xbit_r408_c112 bl[112] br[112] wl[408] vdd gnd cell_6t
Xbit_r409_c112 bl[112] br[112] wl[409] vdd gnd cell_6t
Xbit_r410_c112 bl[112] br[112] wl[410] vdd gnd cell_6t
Xbit_r411_c112 bl[112] br[112] wl[411] vdd gnd cell_6t
Xbit_r412_c112 bl[112] br[112] wl[412] vdd gnd cell_6t
Xbit_r413_c112 bl[112] br[112] wl[413] vdd gnd cell_6t
Xbit_r414_c112 bl[112] br[112] wl[414] vdd gnd cell_6t
Xbit_r415_c112 bl[112] br[112] wl[415] vdd gnd cell_6t
Xbit_r416_c112 bl[112] br[112] wl[416] vdd gnd cell_6t
Xbit_r417_c112 bl[112] br[112] wl[417] vdd gnd cell_6t
Xbit_r418_c112 bl[112] br[112] wl[418] vdd gnd cell_6t
Xbit_r419_c112 bl[112] br[112] wl[419] vdd gnd cell_6t
Xbit_r420_c112 bl[112] br[112] wl[420] vdd gnd cell_6t
Xbit_r421_c112 bl[112] br[112] wl[421] vdd gnd cell_6t
Xbit_r422_c112 bl[112] br[112] wl[422] vdd gnd cell_6t
Xbit_r423_c112 bl[112] br[112] wl[423] vdd gnd cell_6t
Xbit_r424_c112 bl[112] br[112] wl[424] vdd gnd cell_6t
Xbit_r425_c112 bl[112] br[112] wl[425] vdd gnd cell_6t
Xbit_r426_c112 bl[112] br[112] wl[426] vdd gnd cell_6t
Xbit_r427_c112 bl[112] br[112] wl[427] vdd gnd cell_6t
Xbit_r428_c112 bl[112] br[112] wl[428] vdd gnd cell_6t
Xbit_r429_c112 bl[112] br[112] wl[429] vdd gnd cell_6t
Xbit_r430_c112 bl[112] br[112] wl[430] vdd gnd cell_6t
Xbit_r431_c112 bl[112] br[112] wl[431] vdd gnd cell_6t
Xbit_r432_c112 bl[112] br[112] wl[432] vdd gnd cell_6t
Xbit_r433_c112 bl[112] br[112] wl[433] vdd gnd cell_6t
Xbit_r434_c112 bl[112] br[112] wl[434] vdd gnd cell_6t
Xbit_r435_c112 bl[112] br[112] wl[435] vdd gnd cell_6t
Xbit_r436_c112 bl[112] br[112] wl[436] vdd gnd cell_6t
Xbit_r437_c112 bl[112] br[112] wl[437] vdd gnd cell_6t
Xbit_r438_c112 bl[112] br[112] wl[438] vdd gnd cell_6t
Xbit_r439_c112 bl[112] br[112] wl[439] vdd gnd cell_6t
Xbit_r440_c112 bl[112] br[112] wl[440] vdd gnd cell_6t
Xbit_r441_c112 bl[112] br[112] wl[441] vdd gnd cell_6t
Xbit_r442_c112 bl[112] br[112] wl[442] vdd gnd cell_6t
Xbit_r443_c112 bl[112] br[112] wl[443] vdd gnd cell_6t
Xbit_r444_c112 bl[112] br[112] wl[444] vdd gnd cell_6t
Xbit_r445_c112 bl[112] br[112] wl[445] vdd gnd cell_6t
Xbit_r446_c112 bl[112] br[112] wl[446] vdd gnd cell_6t
Xbit_r447_c112 bl[112] br[112] wl[447] vdd gnd cell_6t
Xbit_r448_c112 bl[112] br[112] wl[448] vdd gnd cell_6t
Xbit_r449_c112 bl[112] br[112] wl[449] vdd gnd cell_6t
Xbit_r450_c112 bl[112] br[112] wl[450] vdd gnd cell_6t
Xbit_r451_c112 bl[112] br[112] wl[451] vdd gnd cell_6t
Xbit_r452_c112 bl[112] br[112] wl[452] vdd gnd cell_6t
Xbit_r453_c112 bl[112] br[112] wl[453] vdd gnd cell_6t
Xbit_r454_c112 bl[112] br[112] wl[454] vdd gnd cell_6t
Xbit_r455_c112 bl[112] br[112] wl[455] vdd gnd cell_6t
Xbit_r456_c112 bl[112] br[112] wl[456] vdd gnd cell_6t
Xbit_r457_c112 bl[112] br[112] wl[457] vdd gnd cell_6t
Xbit_r458_c112 bl[112] br[112] wl[458] vdd gnd cell_6t
Xbit_r459_c112 bl[112] br[112] wl[459] vdd gnd cell_6t
Xbit_r460_c112 bl[112] br[112] wl[460] vdd gnd cell_6t
Xbit_r461_c112 bl[112] br[112] wl[461] vdd gnd cell_6t
Xbit_r462_c112 bl[112] br[112] wl[462] vdd gnd cell_6t
Xbit_r463_c112 bl[112] br[112] wl[463] vdd gnd cell_6t
Xbit_r464_c112 bl[112] br[112] wl[464] vdd gnd cell_6t
Xbit_r465_c112 bl[112] br[112] wl[465] vdd gnd cell_6t
Xbit_r466_c112 bl[112] br[112] wl[466] vdd gnd cell_6t
Xbit_r467_c112 bl[112] br[112] wl[467] vdd gnd cell_6t
Xbit_r468_c112 bl[112] br[112] wl[468] vdd gnd cell_6t
Xbit_r469_c112 bl[112] br[112] wl[469] vdd gnd cell_6t
Xbit_r470_c112 bl[112] br[112] wl[470] vdd gnd cell_6t
Xbit_r471_c112 bl[112] br[112] wl[471] vdd gnd cell_6t
Xbit_r472_c112 bl[112] br[112] wl[472] vdd gnd cell_6t
Xbit_r473_c112 bl[112] br[112] wl[473] vdd gnd cell_6t
Xbit_r474_c112 bl[112] br[112] wl[474] vdd gnd cell_6t
Xbit_r475_c112 bl[112] br[112] wl[475] vdd gnd cell_6t
Xbit_r476_c112 bl[112] br[112] wl[476] vdd gnd cell_6t
Xbit_r477_c112 bl[112] br[112] wl[477] vdd gnd cell_6t
Xbit_r478_c112 bl[112] br[112] wl[478] vdd gnd cell_6t
Xbit_r479_c112 bl[112] br[112] wl[479] vdd gnd cell_6t
Xbit_r480_c112 bl[112] br[112] wl[480] vdd gnd cell_6t
Xbit_r481_c112 bl[112] br[112] wl[481] vdd gnd cell_6t
Xbit_r482_c112 bl[112] br[112] wl[482] vdd gnd cell_6t
Xbit_r483_c112 bl[112] br[112] wl[483] vdd gnd cell_6t
Xbit_r484_c112 bl[112] br[112] wl[484] vdd gnd cell_6t
Xbit_r485_c112 bl[112] br[112] wl[485] vdd gnd cell_6t
Xbit_r486_c112 bl[112] br[112] wl[486] vdd gnd cell_6t
Xbit_r487_c112 bl[112] br[112] wl[487] vdd gnd cell_6t
Xbit_r488_c112 bl[112] br[112] wl[488] vdd gnd cell_6t
Xbit_r489_c112 bl[112] br[112] wl[489] vdd gnd cell_6t
Xbit_r490_c112 bl[112] br[112] wl[490] vdd gnd cell_6t
Xbit_r491_c112 bl[112] br[112] wl[491] vdd gnd cell_6t
Xbit_r492_c112 bl[112] br[112] wl[492] vdd gnd cell_6t
Xbit_r493_c112 bl[112] br[112] wl[493] vdd gnd cell_6t
Xbit_r494_c112 bl[112] br[112] wl[494] vdd gnd cell_6t
Xbit_r495_c112 bl[112] br[112] wl[495] vdd gnd cell_6t
Xbit_r496_c112 bl[112] br[112] wl[496] vdd gnd cell_6t
Xbit_r497_c112 bl[112] br[112] wl[497] vdd gnd cell_6t
Xbit_r498_c112 bl[112] br[112] wl[498] vdd gnd cell_6t
Xbit_r499_c112 bl[112] br[112] wl[499] vdd gnd cell_6t
Xbit_r500_c112 bl[112] br[112] wl[500] vdd gnd cell_6t
Xbit_r501_c112 bl[112] br[112] wl[501] vdd gnd cell_6t
Xbit_r502_c112 bl[112] br[112] wl[502] vdd gnd cell_6t
Xbit_r503_c112 bl[112] br[112] wl[503] vdd gnd cell_6t
Xbit_r504_c112 bl[112] br[112] wl[504] vdd gnd cell_6t
Xbit_r505_c112 bl[112] br[112] wl[505] vdd gnd cell_6t
Xbit_r506_c112 bl[112] br[112] wl[506] vdd gnd cell_6t
Xbit_r507_c112 bl[112] br[112] wl[507] vdd gnd cell_6t
Xbit_r508_c112 bl[112] br[112] wl[508] vdd gnd cell_6t
Xbit_r509_c112 bl[112] br[112] wl[509] vdd gnd cell_6t
Xbit_r510_c112 bl[112] br[112] wl[510] vdd gnd cell_6t
Xbit_r511_c112 bl[112] br[112] wl[511] vdd gnd cell_6t
Xbit_r0_c113 bl[113] br[113] wl[0] vdd gnd cell_6t
Xbit_r1_c113 bl[113] br[113] wl[1] vdd gnd cell_6t
Xbit_r2_c113 bl[113] br[113] wl[2] vdd gnd cell_6t
Xbit_r3_c113 bl[113] br[113] wl[3] vdd gnd cell_6t
Xbit_r4_c113 bl[113] br[113] wl[4] vdd gnd cell_6t
Xbit_r5_c113 bl[113] br[113] wl[5] vdd gnd cell_6t
Xbit_r6_c113 bl[113] br[113] wl[6] vdd gnd cell_6t
Xbit_r7_c113 bl[113] br[113] wl[7] vdd gnd cell_6t
Xbit_r8_c113 bl[113] br[113] wl[8] vdd gnd cell_6t
Xbit_r9_c113 bl[113] br[113] wl[9] vdd gnd cell_6t
Xbit_r10_c113 bl[113] br[113] wl[10] vdd gnd cell_6t
Xbit_r11_c113 bl[113] br[113] wl[11] vdd gnd cell_6t
Xbit_r12_c113 bl[113] br[113] wl[12] vdd gnd cell_6t
Xbit_r13_c113 bl[113] br[113] wl[13] vdd gnd cell_6t
Xbit_r14_c113 bl[113] br[113] wl[14] vdd gnd cell_6t
Xbit_r15_c113 bl[113] br[113] wl[15] vdd gnd cell_6t
Xbit_r16_c113 bl[113] br[113] wl[16] vdd gnd cell_6t
Xbit_r17_c113 bl[113] br[113] wl[17] vdd gnd cell_6t
Xbit_r18_c113 bl[113] br[113] wl[18] vdd gnd cell_6t
Xbit_r19_c113 bl[113] br[113] wl[19] vdd gnd cell_6t
Xbit_r20_c113 bl[113] br[113] wl[20] vdd gnd cell_6t
Xbit_r21_c113 bl[113] br[113] wl[21] vdd gnd cell_6t
Xbit_r22_c113 bl[113] br[113] wl[22] vdd gnd cell_6t
Xbit_r23_c113 bl[113] br[113] wl[23] vdd gnd cell_6t
Xbit_r24_c113 bl[113] br[113] wl[24] vdd gnd cell_6t
Xbit_r25_c113 bl[113] br[113] wl[25] vdd gnd cell_6t
Xbit_r26_c113 bl[113] br[113] wl[26] vdd gnd cell_6t
Xbit_r27_c113 bl[113] br[113] wl[27] vdd gnd cell_6t
Xbit_r28_c113 bl[113] br[113] wl[28] vdd gnd cell_6t
Xbit_r29_c113 bl[113] br[113] wl[29] vdd gnd cell_6t
Xbit_r30_c113 bl[113] br[113] wl[30] vdd gnd cell_6t
Xbit_r31_c113 bl[113] br[113] wl[31] vdd gnd cell_6t
Xbit_r32_c113 bl[113] br[113] wl[32] vdd gnd cell_6t
Xbit_r33_c113 bl[113] br[113] wl[33] vdd gnd cell_6t
Xbit_r34_c113 bl[113] br[113] wl[34] vdd gnd cell_6t
Xbit_r35_c113 bl[113] br[113] wl[35] vdd gnd cell_6t
Xbit_r36_c113 bl[113] br[113] wl[36] vdd gnd cell_6t
Xbit_r37_c113 bl[113] br[113] wl[37] vdd gnd cell_6t
Xbit_r38_c113 bl[113] br[113] wl[38] vdd gnd cell_6t
Xbit_r39_c113 bl[113] br[113] wl[39] vdd gnd cell_6t
Xbit_r40_c113 bl[113] br[113] wl[40] vdd gnd cell_6t
Xbit_r41_c113 bl[113] br[113] wl[41] vdd gnd cell_6t
Xbit_r42_c113 bl[113] br[113] wl[42] vdd gnd cell_6t
Xbit_r43_c113 bl[113] br[113] wl[43] vdd gnd cell_6t
Xbit_r44_c113 bl[113] br[113] wl[44] vdd gnd cell_6t
Xbit_r45_c113 bl[113] br[113] wl[45] vdd gnd cell_6t
Xbit_r46_c113 bl[113] br[113] wl[46] vdd gnd cell_6t
Xbit_r47_c113 bl[113] br[113] wl[47] vdd gnd cell_6t
Xbit_r48_c113 bl[113] br[113] wl[48] vdd gnd cell_6t
Xbit_r49_c113 bl[113] br[113] wl[49] vdd gnd cell_6t
Xbit_r50_c113 bl[113] br[113] wl[50] vdd gnd cell_6t
Xbit_r51_c113 bl[113] br[113] wl[51] vdd gnd cell_6t
Xbit_r52_c113 bl[113] br[113] wl[52] vdd gnd cell_6t
Xbit_r53_c113 bl[113] br[113] wl[53] vdd gnd cell_6t
Xbit_r54_c113 bl[113] br[113] wl[54] vdd gnd cell_6t
Xbit_r55_c113 bl[113] br[113] wl[55] vdd gnd cell_6t
Xbit_r56_c113 bl[113] br[113] wl[56] vdd gnd cell_6t
Xbit_r57_c113 bl[113] br[113] wl[57] vdd gnd cell_6t
Xbit_r58_c113 bl[113] br[113] wl[58] vdd gnd cell_6t
Xbit_r59_c113 bl[113] br[113] wl[59] vdd gnd cell_6t
Xbit_r60_c113 bl[113] br[113] wl[60] vdd gnd cell_6t
Xbit_r61_c113 bl[113] br[113] wl[61] vdd gnd cell_6t
Xbit_r62_c113 bl[113] br[113] wl[62] vdd gnd cell_6t
Xbit_r63_c113 bl[113] br[113] wl[63] vdd gnd cell_6t
Xbit_r64_c113 bl[113] br[113] wl[64] vdd gnd cell_6t
Xbit_r65_c113 bl[113] br[113] wl[65] vdd gnd cell_6t
Xbit_r66_c113 bl[113] br[113] wl[66] vdd gnd cell_6t
Xbit_r67_c113 bl[113] br[113] wl[67] vdd gnd cell_6t
Xbit_r68_c113 bl[113] br[113] wl[68] vdd gnd cell_6t
Xbit_r69_c113 bl[113] br[113] wl[69] vdd gnd cell_6t
Xbit_r70_c113 bl[113] br[113] wl[70] vdd gnd cell_6t
Xbit_r71_c113 bl[113] br[113] wl[71] vdd gnd cell_6t
Xbit_r72_c113 bl[113] br[113] wl[72] vdd gnd cell_6t
Xbit_r73_c113 bl[113] br[113] wl[73] vdd gnd cell_6t
Xbit_r74_c113 bl[113] br[113] wl[74] vdd gnd cell_6t
Xbit_r75_c113 bl[113] br[113] wl[75] vdd gnd cell_6t
Xbit_r76_c113 bl[113] br[113] wl[76] vdd gnd cell_6t
Xbit_r77_c113 bl[113] br[113] wl[77] vdd gnd cell_6t
Xbit_r78_c113 bl[113] br[113] wl[78] vdd gnd cell_6t
Xbit_r79_c113 bl[113] br[113] wl[79] vdd gnd cell_6t
Xbit_r80_c113 bl[113] br[113] wl[80] vdd gnd cell_6t
Xbit_r81_c113 bl[113] br[113] wl[81] vdd gnd cell_6t
Xbit_r82_c113 bl[113] br[113] wl[82] vdd gnd cell_6t
Xbit_r83_c113 bl[113] br[113] wl[83] vdd gnd cell_6t
Xbit_r84_c113 bl[113] br[113] wl[84] vdd gnd cell_6t
Xbit_r85_c113 bl[113] br[113] wl[85] vdd gnd cell_6t
Xbit_r86_c113 bl[113] br[113] wl[86] vdd gnd cell_6t
Xbit_r87_c113 bl[113] br[113] wl[87] vdd gnd cell_6t
Xbit_r88_c113 bl[113] br[113] wl[88] vdd gnd cell_6t
Xbit_r89_c113 bl[113] br[113] wl[89] vdd gnd cell_6t
Xbit_r90_c113 bl[113] br[113] wl[90] vdd gnd cell_6t
Xbit_r91_c113 bl[113] br[113] wl[91] vdd gnd cell_6t
Xbit_r92_c113 bl[113] br[113] wl[92] vdd gnd cell_6t
Xbit_r93_c113 bl[113] br[113] wl[93] vdd gnd cell_6t
Xbit_r94_c113 bl[113] br[113] wl[94] vdd gnd cell_6t
Xbit_r95_c113 bl[113] br[113] wl[95] vdd gnd cell_6t
Xbit_r96_c113 bl[113] br[113] wl[96] vdd gnd cell_6t
Xbit_r97_c113 bl[113] br[113] wl[97] vdd gnd cell_6t
Xbit_r98_c113 bl[113] br[113] wl[98] vdd gnd cell_6t
Xbit_r99_c113 bl[113] br[113] wl[99] vdd gnd cell_6t
Xbit_r100_c113 bl[113] br[113] wl[100] vdd gnd cell_6t
Xbit_r101_c113 bl[113] br[113] wl[101] vdd gnd cell_6t
Xbit_r102_c113 bl[113] br[113] wl[102] vdd gnd cell_6t
Xbit_r103_c113 bl[113] br[113] wl[103] vdd gnd cell_6t
Xbit_r104_c113 bl[113] br[113] wl[104] vdd gnd cell_6t
Xbit_r105_c113 bl[113] br[113] wl[105] vdd gnd cell_6t
Xbit_r106_c113 bl[113] br[113] wl[106] vdd gnd cell_6t
Xbit_r107_c113 bl[113] br[113] wl[107] vdd gnd cell_6t
Xbit_r108_c113 bl[113] br[113] wl[108] vdd gnd cell_6t
Xbit_r109_c113 bl[113] br[113] wl[109] vdd gnd cell_6t
Xbit_r110_c113 bl[113] br[113] wl[110] vdd gnd cell_6t
Xbit_r111_c113 bl[113] br[113] wl[111] vdd gnd cell_6t
Xbit_r112_c113 bl[113] br[113] wl[112] vdd gnd cell_6t
Xbit_r113_c113 bl[113] br[113] wl[113] vdd gnd cell_6t
Xbit_r114_c113 bl[113] br[113] wl[114] vdd gnd cell_6t
Xbit_r115_c113 bl[113] br[113] wl[115] vdd gnd cell_6t
Xbit_r116_c113 bl[113] br[113] wl[116] vdd gnd cell_6t
Xbit_r117_c113 bl[113] br[113] wl[117] vdd gnd cell_6t
Xbit_r118_c113 bl[113] br[113] wl[118] vdd gnd cell_6t
Xbit_r119_c113 bl[113] br[113] wl[119] vdd gnd cell_6t
Xbit_r120_c113 bl[113] br[113] wl[120] vdd gnd cell_6t
Xbit_r121_c113 bl[113] br[113] wl[121] vdd gnd cell_6t
Xbit_r122_c113 bl[113] br[113] wl[122] vdd gnd cell_6t
Xbit_r123_c113 bl[113] br[113] wl[123] vdd gnd cell_6t
Xbit_r124_c113 bl[113] br[113] wl[124] vdd gnd cell_6t
Xbit_r125_c113 bl[113] br[113] wl[125] vdd gnd cell_6t
Xbit_r126_c113 bl[113] br[113] wl[126] vdd gnd cell_6t
Xbit_r127_c113 bl[113] br[113] wl[127] vdd gnd cell_6t
Xbit_r128_c113 bl[113] br[113] wl[128] vdd gnd cell_6t
Xbit_r129_c113 bl[113] br[113] wl[129] vdd gnd cell_6t
Xbit_r130_c113 bl[113] br[113] wl[130] vdd gnd cell_6t
Xbit_r131_c113 bl[113] br[113] wl[131] vdd gnd cell_6t
Xbit_r132_c113 bl[113] br[113] wl[132] vdd gnd cell_6t
Xbit_r133_c113 bl[113] br[113] wl[133] vdd gnd cell_6t
Xbit_r134_c113 bl[113] br[113] wl[134] vdd gnd cell_6t
Xbit_r135_c113 bl[113] br[113] wl[135] vdd gnd cell_6t
Xbit_r136_c113 bl[113] br[113] wl[136] vdd gnd cell_6t
Xbit_r137_c113 bl[113] br[113] wl[137] vdd gnd cell_6t
Xbit_r138_c113 bl[113] br[113] wl[138] vdd gnd cell_6t
Xbit_r139_c113 bl[113] br[113] wl[139] vdd gnd cell_6t
Xbit_r140_c113 bl[113] br[113] wl[140] vdd gnd cell_6t
Xbit_r141_c113 bl[113] br[113] wl[141] vdd gnd cell_6t
Xbit_r142_c113 bl[113] br[113] wl[142] vdd gnd cell_6t
Xbit_r143_c113 bl[113] br[113] wl[143] vdd gnd cell_6t
Xbit_r144_c113 bl[113] br[113] wl[144] vdd gnd cell_6t
Xbit_r145_c113 bl[113] br[113] wl[145] vdd gnd cell_6t
Xbit_r146_c113 bl[113] br[113] wl[146] vdd gnd cell_6t
Xbit_r147_c113 bl[113] br[113] wl[147] vdd gnd cell_6t
Xbit_r148_c113 bl[113] br[113] wl[148] vdd gnd cell_6t
Xbit_r149_c113 bl[113] br[113] wl[149] vdd gnd cell_6t
Xbit_r150_c113 bl[113] br[113] wl[150] vdd gnd cell_6t
Xbit_r151_c113 bl[113] br[113] wl[151] vdd gnd cell_6t
Xbit_r152_c113 bl[113] br[113] wl[152] vdd gnd cell_6t
Xbit_r153_c113 bl[113] br[113] wl[153] vdd gnd cell_6t
Xbit_r154_c113 bl[113] br[113] wl[154] vdd gnd cell_6t
Xbit_r155_c113 bl[113] br[113] wl[155] vdd gnd cell_6t
Xbit_r156_c113 bl[113] br[113] wl[156] vdd gnd cell_6t
Xbit_r157_c113 bl[113] br[113] wl[157] vdd gnd cell_6t
Xbit_r158_c113 bl[113] br[113] wl[158] vdd gnd cell_6t
Xbit_r159_c113 bl[113] br[113] wl[159] vdd gnd cell_6t
Xbit_r160_c113 bl[113] br[113] wl[160] vdd gnd cell_6t
Xbit_r161_c113 bl[113] br[113] wl[161] vdd gnd cell_6t
Xbit_r162_c113 bl[113] br[113] wl[162] vdd gnd cell_6t
Xbit_r163_c113 bl[113] br[113] wl[163] vdd gnd cell_6t
Xbit_r164_c113 bl[113] br[113] wl[164] vdd gnd cell_6t
Xbit_r165_c113 bl[113] br[113] wl[165] vdd gnd cell_6t
Xbit_r166_c113 bl[113] br[113] wl[166] vdd gnd cell_6t
Xbit_r167_c113 bl[113] br[113] wl[167] vdd gnd cell_6t
Xbit_r168_c113 bl[113] br[113] wl[168] vdd gnd cell_6t
Xbit_r169_c113 bl[113] br[113] wl[169] vdd gnd cell_6t
Xbit_r170_c113 bl[113] br[113] wl[170] vdd gnd cell_6t
Xbit_r171_c113 bl[113] br[113] wl[171] vdd gnd cell_6t
Xbit_r172_c113 bl[113] br[113] wl[172] vdd gnd cell_6t
Xbit_r173_c113 bl[113] br[113] wl[173] vdd gnd cell_6t
Xbit_r174_c113 bl[113] br[113] wl[174] vdd gnd cell_6t
Xbit_r175_c113 bl[113] br[113] wl[175] vdd gnd cell_6t
Xbit_r176_c113 bl[113] br[113] wl[176] vdd gnd cell_6t
Xbit_r177_c113 bl[113] br[113] wl[177] vdd gnd cell_6t
Xbit_r178_c113 bl[113] br[113] wl[178] vdd gnd cell_6t
Xbit_r179_c113 bl[113] br[113] wl[179] vdd gnd cell_6t
Xbit_r180_c113 bl[113] br[113] wl[180] vdd gnd cell_6t
Xbit_r181_c113 bl[113] br[113] wl[181] vdd gnd cell_6t
Xbit_r182_c113 bl[113] br[113] wl[182] vdd gnd cell_6t
Xbit_r183_c113 bl[113] br[113] wl[183] vdd gnd cell_6t
Xbit_r184_c113 bl[113] br[113] wl[184] vdd gnd cell_6t
Xbit_r185_c113 bl[113] br[113] wl[185] vdd gnd cell_6t
Xbit_r186_c113 bl[113] br[113] wl[186] vdd gnd cell_6t
Xbit_r187_c113 bl[113] br[113] wl[187] vdd gnd cell_6t
Xbit_r188_c113 bl[113] br[113] wl[188] vdd gnd cell_6t
Xbit_r189_c113 bl[113] br[113] wl[189] vdd gnd cell_6t
Xbit_r190_c113 bl[113] br[113] wl[190] vdd gnd cell_6t
Xbit_r191_c113 bl[113] br[113] wl[191] vdd gnd cell_6t
Xbit_r192_c113 bl[113] br[113] wl[192] vdd gnd cell_6t
Xbit_r193_c113 bl[113] br[113] wl[193] vdd gnd cell_6t
Xbit_r194_c113 bl[113] br[113] wl[194] vdd gnd cell_6t
Xbit_r195_c113 bl[113] br[113] wl[195] vdd gnd cell_6t
Xbit_r196_c113 bl[113] br[113] wl[196] vdd gnd cell_6t
Xbit_r197_c113 bl[113] br[113] wl[197] vdd gnd cell_6t
Xbit_r198_c113 bl[113] br[113] wl[198] vdd gnd cell_6t
Xbit_r199_c113 bl[113] br[113] wl[199] vdd gnd cell_6t
Xbit_r200_c113 bl[113] br[113] wl[200] vdd gnd cell_6t
Xbit_r201_c113 bl[113] br[113] wl[201] vdd gnd cell_6t
Xbit_r202_c113 bl[113] br[113] wl[202] vdd gnd cell_6t
Xbit_r203_c113 bl[113] br[113] wl[203] vdd gnd cell_6t
Xbit_r204_c113 bl[113] br[113] wl[204] vdd gnd cell_6t
Xbit_r205_c113 bl[113] br[113] wl[205] vdd gnd cell_6t
Xbit_r206_c113 bl[113] br[113] wl[206] vdd gnd cell_6t
Xbit_r207_c113 bl[113] br[113] wl[207] vdd gnd cell_6t
Xbit_r208_c113 bl[113] br[113] wl[208] vdd gnd cell_6t
Xbit_r209_c113 bl[113] br[113] wl[209] vdd gnd cell_6t
Xbit_r210_c113 bl[113] br[113] wl[210] vdd gnd cell_6t
Xbit_r211_c113 bl[113] br[113] wl[211] vdd gnd cell_6t
Xbit_r212_c113 bl[113] br[113] wl[212] vdd gnd cell_6t
Xbit_r213_c113 bl[113] br[113] wl[213] vdd gnd cell_6t
Xbit_r214_c113 bl[113] br[113] wl[214] vdd gnd cell_6t
Xbit_r215_c113 bl[113] br[113] wl[215] vdd gnd cell_6t
Xbit_r216_c113 bl[113] br[113] wl[216] vdd gnd cell_6t
Xbit_r217_c113 bl[113] br[113] wl[217] vdd gnd cell_6t
Xbit_r218_c113 bl[113] br[113] wl[218] vdd gnd cell_6t
Xbit_r219_c113 bl[113] br[113] wl[219] vdd gnd cell_6t
Xbit_r220_c113 bl[113] br[113] wl[220] vdd gnd cell_6t
Xbit_r221_c113 bl[113] br[113] wl[221] vdd gnd cell_6t
Xbit_r222_c113 bl[113] br[113] wl[222] vdd gnd cell_6t
Xbit_r223_c113 bl[113] br[113] wl[223] vdd gnd cell_6t
Xbit_r224_c113 bl[113] br[113] wl[224] vdd gnd cell_6t
Xbit_r225_c113 bl[113] br[113] wl[225] vdd gnd cell_6t
Xbit_r226_c113 bl[113] br[113] wl[226] vdd gnd cell_6t
Xbit_r227_c113 bl[113] br[113] wl[227] vdd gnd cell_6t
Xbit_r228_c113 bl[113] br[113] wl[228] vdd gnd cell_6t
Xbit_r229_c113 bl[113] br[113] wl[229] vdd gnd cell_6t
Xbit_r230_c113 bl[113] br[113] wl[230] vdd gnd cell_6t
Xbit_r231_c113 bl[113] br[113] wl[231] vdd gnd cell_6t
Xbit_r232_c113 bl[113] br[113] wl[232] vdd gnd cell_6t
Xbit_r233_c113 bl[113] br[113] wl[233] vdd gnd cell_6t
Xbit_r234_c113 bl[113] br[113] wl[234] vdd gnd cell_6t
Xbit_r235_c113 bl[113] br[113] wl[235] vdd gnd cell_6t
Xbit_r236_c113 bl[113] br[113] wl[236] vdd gnd cell_6t
Xbit_r237_c113 bl[113] br[113] wl[237] vdd gnd cell_6t
Xbit_r238_c113 bl[113] br[113] wl[238] vdd gnd cell_6t
Xbit_r239_c113 bl[113] br[113] wl[239] vdd gnd cell_6t
Xbit_r240_c113 bl[113] br[113] wl[240] vdd gnd cell_6t
Xbit_r241_c113 bl[113] br[113] wl[241] vdd gnd cell_6t
Xbit_r242_c113 bl[113] br[113] wl[242] vdd gnd cell_6t
Xbit_r243_c113 bl[113] br[113] wl[243] vdd gnd cell_6t
Xbit_r244_c113 bl[113] br[113] wl[244] vdd gnd cell_6t
Xbit_r245_c113 bl[113] br[113] wl[245] vdd gnd cell_6t
Xbit_r246_c113 bl[113] br[113] wl[246] vdd gnd cell_6t
Xbit_r247_c113 bl[113] br[113] wl[247] vdd gnd cell_6t
Xbit_r248_c113 bl[113] br[113] wl[248] vdd gnd cell_6t
Xbit_r249_c113 bl[113] br[113] wl[249] vdd gnd cell_6t
Xbit_r250_c113 bl[113] br[113] wl[250] vdd gnd cell_6t
Xbit_r251_c113 bl[113] br[113] wl[251] vdd gnd cell_6t
Xbit_r252_c113 bl[113] br[113] wl[252] vdd gnd cell_6t
Xbit_r253_c113 bl[113] br[113] wl[253] vdd gnd cell_6t
Xbit_r254_c113 bl[113] br[113] wl[254] vdd gnd cell_6t
Xbit_r255_c113 bl[113] br[113] wl[255] vdd gnd cell_6t
Xbit_r256_c113 bl[113] br[113] wl[256] vdd gnd cell_6t
Xbit_r257_c113 bl[113] br[113] wl[257] vdd gnd cell_6t
Xbit_r258_c113 bl[113] br[113] wl[258] vdd gnd cell_6t
Xbit_r259_c113 bl[113] br[113] wl[259] vdd gnd cell_6t
Xbit_r260_c113 bl[113] br[113] wl[260] vdd gnd cell_6t
Xbit_r261_c113 bl[113] br[113] wl[261] vdd gnd cell_6t
Xbit_r262_c113 bl[113] br[113] wl[262] vdd gnd cell_6t
Xbit_r263_c113 bl[113] br[113] wl[263] vdd gnd cell_6t
Xbit_r264_c113 bl[113] br[113] wl[264] vdd gnd cell_6t
Xbit_r265_c113 bl[113] br[113] wl[265] vdd gnd cell_6t
Xbit_r266_c113 bl[113] br[113] wl[266] vdd gnd cell_6t
Xbit_r267_c113 bl[113] br[113] wl[267] vdd gnd cell_6t
Xbit_r268_c113 bl[113] br[113] wl[268] vdd gnd cell_6t
Xbit_r269_c113 bl[113] br[113] wl[269] vdd gnd cell_6t
Xbit_r270_c113 bl[113] br[113] wl[270] vdd gnd cell_6t
Xbit_r271_c113 bl[113] br[113] wl[271] vdd gnd cell_6t
Xbit_r272_c113 bl[113] br[113] wl[272] vdd gnd cell_6t
Xbit_r273_c113 bl[113] br[113] wl[273] vdd gnd cell_6t
Xbit_r274_c113 bl[113] br[113] wl[274] vdd gnd cell_6t
Xbit_r275_c113 bl[113] br[113] wl[275] vdd gnd cell_6t
Xbit_r276_c113 bl[113] br[113] wl[276] vdd gnd cell_6t
Xbit_r277_c113 bl[113] br[113] wl[277] vdd gnd cell_6t
Xbit_r278_c113 bl[113] br[113] wl[278] vdd gnd cell_6t
Xbit_r279_c113 bl[113] br[113] wl[279] vdd gnd cell_6t
Xbit_r280_c113 bl[113] br[113] wl[280] vdd gnd cell_6t
Xbit_r281_c113 bl[113] br[113] wl[281] vdd gnd cell_6t
Xbit_r282_c113 bl[113] br[113] wl[282] vdd gnd cell_6t
Xbit_r283_c113 bl[113] br[113] wl[283] vdd gnd cell_6t
Xbit_r284_c113 bl[113] br[113] wl[284] vdd gnd cell_6t
Xbit_r285_c113 bl[113] br[113] wl[285] vdd gnd cell_6t
Xbit_r286_c113 bl[113] br[113] wl[286] vdd gnd cell_6t
Xbit_r287_c113 bl[113] br[113] wl[287] vdd gnd cell_6t
Xbit_r288_c113 bl[113] br[113] wl[288] vdd gnd cell_6t
Xbit_r289_c113 bl[113] br[113] wl[289] vdd gnd cell_6t
Xbit_r290_c113 bl[113] br[113] wl[290] vdd gnd cell_6t
Xbit_r291_c113 bl[113] br[113] wl[291] vdd gnd cell_6t
Xbit_r292_c113 bl[113] br[113] wl[292] vdd gnd cell_6t
Xbit_r293_c113 bl[113] br[113] wl[293] vdd gnd cell_6t
Xbit_r294_c113 bl[113] br[113] wl[294] vdd gnd cell_6t
Xbit_r295_c113 bl[113] br[113] wl[295] vdd gnd cell_6t
Xbit_r296_c113 bl[113] br[113] wl[296] vdd gnd cell_6t
Xbit_r297_c113 bl[113] br[113] wl[297] vdd gnd cell_6t
Xbit_r298_c113 bl[113] br[113] wl[298] vdd gnd cell_6t
Xbit_r299_c113 bl[113] br[113] wl[299] vdd gnd cell_6t
Xbit_r300_c113 bl[113] br[113] wl[300] vdd gnd cell_6t
Xbit_r301_c113 bl[113] br[113] wl[301] vdd gnd cell_6t
Xbit_r302_c113 bl[113] br[113] wl[302] vdd gnd cell_6t
Xbit_r303_c113 bl[113] br[113] wl[303] vdd gnd cell_6t
Xbit_r304_c113 bl[113] br[113] wl[304] vdd gnd cell_6t
Xbit_r305_c113 bl[113] br[113] wl[305] vdd gnd cell_6t
Xbit_r306_c113 bl[113] br[113] wl[306] vdd gnd cell_6t
Xbit_r307_c113 bl[113] br[113] wl[307] vdd gnd cell_6t
Xbit_r308_c113 bl[113] br[113] wl[308] vdd gnd cell_6t
Xbit_r309_c113 bl[113] br[113] wl[309] vdd gnd cell_6t
Xbit_r310_c113 bl[113] br[113] wl[310] vdd gnd cell_6t
Xbit_r311_c113 bl[113] br[113] wl[311] vdd gnd cell_6t
Xbit_r312_c113 bl[113] br[113] wl[312] vdd gnd cell_6t
Xbit_r313_c113 bl[113] br[113] wl[313] vdd gnd cell_6t
Xbit_r314_c113 bl[113] br[113] wl[314] vdd gnd cell_6t
Xbit_r315_c113 bl[113] br[113] wl[315] vdd gnd cell_6t
Xbit_r316_c113 bl[113] br[113] wl[316] vdd gnd cell_6t
Xbit_r317_c113 bl[113] br[113] wl[317] vdd gnd cell_6t
Xbit_r318_c113 bl[113] br[113] wl[318] vdd gnd cell_6t
Xbit_r319_c113 bl[113] br[113] wl[319] vdd gnd cell_6t
Xbit_r320_c113 bl[113] br[113] wl[320] vdd gnd cell_6t
Xbit_r321_c113 bl[113] br[113] wl[321] vdd gnd cell_6t
Xbit_r322_c113 bl[113] br[113] wl[322] vdd gnd cell_6t
Xbit_r323_c113 bl[113] br[113] wl[323] vdd gnd cell_6t
Xbit_r324_c113 bl[113] br[113] wl[324] vdd gnd cell_6t
Xbit_r325_c113 bl[113] br[113] wl[325] vdd gnd cell_6t
Xbit_r326_c113 bl[113] br[113] wl[326] vdd gnd cell_6t
Xbit_r327_c113 bl[113] br[113] wl[327] vdd gnd cell_6t
Xbit_r328_c113 bl[113] br[113] wl[328] vdd gnd cell_6t
Xbit_r329_c113 bl[113] br[113] wl[329] vdd gnd cell_6t
Xbit_r330_c113 bl[113] br[113] wl[330] vdd gnd cell_6t
Xbit_r331_c113 bl[113] br[113] wl[331] vdd gnd cell_6t
Xbit_r332_c113 bl[113] br[113] wl[332] vdd gnd cell_6t
Xbit_r333_c113 bl[113] br[113] wl[333] vdd gnd cell_6t
Xbit_r334_c113 bl[113] br[113] wl[334] vdd gnd cell_6t
Xbit_r335_c113 bl[113] br[113] wl[335] vdd gnd cell_6t
Xbit_r336_c113 bl[113] br[113] wl[336] vdd gnd cell_6t
Xbit_r337_c113 bl[113] br[113] wl[337] vdd gnd cell_6t
Xbit_r338_c113 bl[113] br[113] wl[338] vdd gnd cell_6t
Xbit_r339_c113 bl[113] br[113] wl[339] vdd gnd cell_6t
Xbit_r340_c113 bl[113] br[113] wl[340] vdd gnd cell_6t
Xbit_r341_c113 bl[113] br[113] wl[341] vdd gnd cell_6t
Xbit_r342_c113 bl[113] br[113] wl[342] vdd gnd cell_6t
Xbit_r343_c113 bl[113] br[113] wl[343] vdd gnd cell_6t
Xbit_r344_c113 bl[113] br[113] wl[344] vdd gnd cell_6t
Xbit_r345_c113 bl[113] br[113] wl[345] vdd gnd cell_6t
Xbit_r346_c113 bl[113] br[113] wl[346] vdd gnd cell_6t
Xbit_r347_c113 bl[113] br[113] wl[347] vdd gnd cell_6t
Xbit_r348_c113 bl[113] br[113] wl[348] vdd gnd cell_6t
Xbit_r349_c113 bl[113] br[113] wl[349] vdd gnd cell_6t
Xbit_r350_c113 bl[113] br[113] wl[350] vdd gnd cell_6t
Xbit_r351_c113 bl[113] br[113] wl[351] vdd gnd cell_6t
Xbit_r352_c113 bl[113] br[113] wl[352] vdd gnd cell_6t
Xbit_r353_c113 bl[113] br[113] wl[353] vdd gnd cell_6t
Xbit_r354_c113 bl[113] br[113] wl[354] vdd gnd cell_6t
Xbit_r355_c113 bl[113] br[113] wl[355] vdd gnd cell_6t
Xbit_r356_c113 bl[113] br[113] wl[356] vdd gnd cell_6t
Xbit_r357_c113 bl[113] br[113] wl[357] vdd gnd cell_6t
Xbit_r358_c113 bl[113] br[113] wl[358] vdd gnd cell_6t
Xbit_r359_c113 bl[113] br[113] wl[359] vdd gnd cell_6t
Xbit_r360_c113 bl[113] br[113] wl[360] vdd gnd cell_6t
Xbit_r361_c113 bl[113] br[113] wl[361] vdd gnd cell_6t
Xbit_r362_c113 bl[113] br[113] wl[362] vdd gnd cell_6t
Xbit_r363_c113 bl[113] br[113] wl[363] vdd gnd cell_6t
Xbit_r364_c113 bl[113] br[113] wl[364] vdd gnd cell_6t
Xbit_r365_c113 bl[113] br[113] wl[365] vdd gnd cell_6t
Xbit_r366_c113 bl[113] br[113] wl[366] vdd gnd cell_6t
Xbit_r367_c113 bl[113] br[113] wl[367] vdd gnd cell_6t
Xbit_r368_c113 bl[113] br[113] wl[368] vdd gnd cell_6t
Xbit_r369_c113 bl[113] br[113] wl[369] vdd gnd cell_6t
Xbit_r370_c113 bl[113] br[113] wl[370] vdd gnd cell_6t
Xbit_r371_c113 bl[113] br[113] wl[371] vdd gnd cell_6t
Xbit_r372_c113 bl[113] br[113] wl[372] vdd gnd cell_6t
Xbit_r373_c113 bl[113] br[113] wl[373] vdd gnd cell_6t
Xbit_r374_c113 bl[113] br[113] wl[374] vdd gnd cell_6t
Xbit_r375_c113 bl[113] br[113] wl[375] vdd gnd cell_6t
Xbit_r376_c113 bl[113] br[113] wl[376] vdd gnd cell_6t
Xbit_r377_c113 bl[113] br[113] wl[377] vdd gnd cell_6t
Xbit_r378_c113 bl[113] br[113] wl[378] vdd gnd cell_6t
Xbit_r379_c113 bl[113] br[113] wl[379] vdd gnd cell_6t
Xbit_r380_c113 bl[113] br[113] wl[380] vdd gnd cell_6t
Xbit_r381_c113 bl[113] br[113] wl[381] vdd gnd cell_6t
Xbit_r382_c113 bl[113] br[113] wl[382] vdd gnd cell_6t
Xbit_r383_c113 bl[113] br[113] wl[383] vdd gnd cell_6t
Xbit_r384_c113 bl[113] br[113] wl[384] vdd gnd cell_6t
Xbit_r385_c113 bl[113] br[113] wl[385] vdd gnd cell_6t
Xbit_r386_c113 bl[113] br[113] wl[386] vdd gnd cell_6t
Xbit_r387_c113 bl[113] br[113] wl[387] vdd gnd cell_6t
Xbit_r388_c113 bl[113] br[113] wl[388] vdd gnd cell_6t
Xbit_r389_c113 bl[113] br[113] wl[389] vdd gnd cell_6t
Xbit_r390_c113 bl[113] br[113] wl[390] vdd gnd cell_6t
Xbit_r391_c113 bl[113] br[113] wl[391] vdd gnd cell_6t
Xbit_r392_c113 bl[113] br[113] wl[392] vdd gnd cell_6t
Xbit_r393_c113 bl[113] br[113] wl[393] vdd gnd cell_6t
Xbit_r394_c113 bl[113] br[113] wl[394] vdd gnd cell_6t
Xbit_r395_c113 bl[113] br[113] wl[395] vdd gnd cell_6t
Xbit_r396_c113 bl[113] br[113] wl[396] vdd gnd cell_6t
Xbit_r397_c113 bl[113] br[113] wl[397] vdd gnd cell_6t
Xbit_r398_c113 bl[113] br[113] wl[398] vdd gnd cell_6t
Xbit_r399_c113 bl[113] br[113] wl[399] vdd gnd cell_6t
Xbit_r400_c113 bl[113] br[113] wl[400] vdd gnd cell_6t
Xbit_r401_c113 bl[113] br[113] wl[401] vdd gnd cell_6t
Xbit_r402_c113 bl[113] br[113] wl[402] vdd gnd cell_6t
Xbit_r403_c113 bl[113] br[113] wl[403] vdd gnd cell_6t
Xbit_r404_c113 bl[113] br[113] wl[404] vdd gnd cell_6t
Xbit_r405_c113 bl[113] br[113] wl[405] vdd gnd cell_6t
Xbit_r406_c113 bl[113] br[113] wl[406] vdd gnd cell_6t
Xbit_r407_c113 bl[113] br[113] wl[407] vdd gnd cell_6t
Xbit_r408_c113 bl[113] br[113] wl[408] vdd gnd cell_6t
Xbit_r409_c113 bl[113] br[113] wl[409] vdd gnd cell_6t
Xbit_r410_c113 bl[113] br[113] wl[410] vdd gnd cell_6t
Xbit_r411_c113 bl[113] br[113] wl[411] vdd gnd cell_6t
Xbit_r412_c113 bl[113] br[113] wl[412] vdd gnd cell_6t
Xbit_r413_c113 bl[113] br[113] wl[413] vdd gnd cell_6t
Xbit_r414_c113 bl[113] br[113] wl[414] vdd gnd cell_6t
Xbit_r415_c113 bl[113] br[113] wl[415] vdd gnd cell_6t
Xbit_r416_c113 bl[113] br[113] wl[416] vdd gnd cell_6t
Xbit_r417_c113 bl[113] br[113] wl[417] vdd gnd cell_6t
Xbit_r418_c113 bl[113] br[113] wl[418] vdd gnd cell_6t
Xbit_r419_c113 bl[113] br[113] wl[419] vdd gnd cell_6t
Xbit_r420_c113 bl[113] br[113] wl[420] vdd gnd cell_6t
Xbit_r421_c113 bl[113] br[113] wl[421] vdd gnd cell_6t
Xbit_r422_c113 bl[113] br[113] wl[422] vdd gnd cell_6t
Xbit_r423_c113 bl[113] br[113] wl[423] vdd gnd cell_6t
Xbit_r424_c113 bl[113] br[113] wl[424] vdd gnd cell_6t
Xbit_r425_c113 bl[113] br[113] wl[425] vdd gnd cell_6t
Xbit_r426_c113 bl[113] br[113] wl[426] vdd gnd cell_6t
Xbit_r427_c113 bl[113] br[113] wl[427] vdd gnd cell_6t
Xbit_r428_c113 bl[113] br[113] wl[428] vdd gnd cell_6t
Xbit_r429_c113 bl[113] br[113] wl[429] vdd gnd cell_6t
Xbit_r430_c113 bl[113] br[113] wl[430] vdd gnd cell_6t
Xbit_r431_c113 bl[113] br[113] wl[431] vdd gnd cell_6t
Xbit_r432_c113 bl[113] br[113] wl[432] vdd gnd cell_6t
Xbit_r433_c113 bl[113] br[113] wl[433] vdd gnd cell_6t
Xbit_r434_c113 bl[113] br[113] wl[434] vdd gnd cell_6t
Xbit_r435_c113 bl[113] br[113] wl[435] vdd gnd cell_6t
Xbit_r436_c113 bl[113] br[113] wl[436] vdd gnd cell_6t
Xbit_r437_c113 bl[113] br[113] wl[437] vdd gnd cell_6t
Xbit_r438_c113 bl[113] br[113] wl[438] vdd gnd cell_6t
Xbit_r439_c113 bl[113] br[113] wl[439] vdd gnd cell_6t
Xbit_r440_c113 bl[113] br[113] wl[440] vdd gnd cell_6t
Xbit_r441_c113 bl[113] br[113] wl[441] vdd gnd cell_6t
Xbit_r442_c113 bl[113] br[113] wl[442] vdd gnd cell_6t
Xbit_r443_c113 bl[113] br[113] wl[443] vdd gnd cell_6t
Xbit_r444_c113 bl[113] br[113] wl[444] vdd gnd cell_6t
Xbit_r445_c113 bl[113] br[113] wl[445] vdd gnd cell_6t
Xbit_r446_c113 bl[113] br[113] wl[446] vdd gnd cell_6t
Xbit_r447_c113 bl[113] br[113] wl[447] vdd gnd cell_6t
Xbit_r448_c113 bl[113] br[113] wl[448] vdd gnd cell_6t
Xbit_r449_c113 bl[113] br[113] wl[449] vdd gnd cell_6t
Xbit_r450_c113 bl[113] br[113] wl[450] vdd gnd cell_6t
Xbit_r451_c113 bl[113] br[113] wl[451] vdd gnd cell_6t
Xbit_r452_c113 bl[113] br[113] wl[452] vdd gnd cell_6t
Xbit_r453_c113 bl[113] br[113] wl[453] vdd gnd cell_6t
Xbit_r454_c113 bl[113] br[113] wl[454] vdd gnd cell_6t
Xbit_r455_c113 bl[113] br[113] wl[455] vdd gnd cell_6t
Xbit_r456_c113 bl[113] br[113] wl[456] vdd gnd cell_6t
Xbit_r457_c113 bl[113] br[113] wl[457] vdd gnd cell_6t
Xbit_r458_c113 bl[113] br[113] wl[458] vdd gnd cell_6t
Xbit_r459_c113 bl[113] br[113] wl[459] vdd gnd cell_6t
Xbit_r460_c113 bl[113] br[113] wl[460] vdd gnd cell_6t
Xbit_r461_c113 bl[113] br[113] wl[461] vdd gnd cell_6t
Xbit_r462_c113 bl[113] br[113] wl[462] vdd gnd cell_6t
Xbit_r463_c113 bl[113] br[113] wl[463] vdd gnd cell_6t
Xbit_r464_c113 bl[113] br[113] wl[464] vdd gnd cell_6t
Xbit_r465_c113 bl[113] br[113] wl[465] vdd gnd cell_6t
Xbit_r466_c113 bl[113] br[113] wl[466] vdd gnd cell_6t
Xbit_r467_c113 bl[113] br[113] wl[467] vdd gnd cell_6t
Xbit_r468_c113 bl[113] br[113] wl[468] vdd gnd cell_6t
Xbit_r469_c113 bl[113] br[113] wl[469] vdd gnd cell_6t
Xbit_r470_c113 bl[113] br[113] wl[470] vdd gnd cell_6t
Xbit_r471_c113 bl[113] br[113] wl[471] vdd gnd cell_6t
Xbit_r472_c113 bl[113] br[113] wl[472] vdd gnd cell_6t
Xbit_r473_c113 bl[113] br[113] wl[473] vdd gnd cell_6t
Xbit_r474_c113 bl[113] br[113] wl[474] vdd gnd cell_6t
Xbit_r475_c113 bl[113] br[113] wl[475] vdd gnd cell_6t
Xbit_r476_c113 bl[113] br[113] wl[476] vdd gnd cell_6t
Xbit_r477_c113 bl[113] br[113] wl[477] vdd gnd cell_6t
Xbit_r478_c113 bl[113] br[113] wl[478] vdd gnd cell_6t
Xbit_r479_c113 bl[113] br[113] wl[479] vdd gnd cell_6t
Xbit_r480_c113 bl[113] br[113] wl[480] vdd gnd cell_6t
Xbit_r481_c113 bl[113] br[113] wl[481] vdd gnd cell_6t
Xbit_r482_c113 bl[113] br[113] wl[482] vdd gnd cell_6t
Xbit_r483_c113 bl[113] br[113] wl[483] vdd gnd cell_6t
Xbit_r484_c113 bl[113] br[113] wl[484] vdd gnd cell_6t
Xbit_r485_c113 bl[113] br[113] wl[485] vdd gnd cell_6t
Xbit_r486_c113 bl[113] br[113] wl[486] vdd gnd cell_6t
Xbit_r487_c113 bl[113] br[113] wl[487] vdd gnd cell_6t
Xbit_r488_c113 bl[113] br[113] wl[488] vdd gnd cell_6t
Xbit_r489_c113 bl[113] br[113] wl[489] vdd gnd cell_6t
Xbit_r490_c113 bl[113] br[113] wl[490] vdd gnd cell_6t
Xbit_r491_c113 bl[113] br[113] wl[491] vdd gnd cell_6t
Xbit_r492_c113 bl[113] br[113] wl[492] vdd gnd cell_6t
Xbit_r493_c113 bl[113] br[113] wl[493] vdd gnd cell_6t
Xbit_r494_c113 bl[113] br[113] wl[494] vdd gnd cell_6t
Xbit_r495_c113 bl[113] br[113] wl[495] vdd gnd cell_6t
Xbit_r496_c113 bl[113] br[113] wl[496] vdd gnd cell_6t
Xbit_r497_c113 bl[113] br[113] wl[497] vdd gnd cell_6t
Xbit_r498_c113 bl[113] br[113] wl[498] vdd gnd cell_6t
Xbit_r499_c113 bl[113] br[113] wl[499] vdd gnd cell_6t
Xbit_r500_c113 bl[113] br[113] wl[500] vdd gnd cell_6t
Xbit_r501_c113 bl[113] br[113] wl[501] vdd gnd cell_6t
Xbit_r502_c113 bl[113] br[113] wl[502] vdd gnd cell_6t
Xbit_r503_c113 bl[113] br[113] wl[503] vdd gnd cell_6t
Xbit_r504_c113 bl[113] br[113] wl[504] vdd gnd cell_6t
Xbit_r505_c113 bl[113] br[113] wl[505] vdd gnd cell_6t
Xbit_r506_c113 bl[113] br[113] wl[506] vdd gnd cell_6t
Xbit_r507_c113 bl[113] br[113] wl[507] vdd gnd cell_6t
Xbit_r508_c113 bl[113] br[113] wl[508] vdd gnd cell_6t
Xbit_r509_c113 bl[113] br[113] wl[509] vdd gnd cell_6t
Xbit_r510_c113 bl[113] br[113] wl[510] vdd gnd cell_6t
Xbit_r511_c113 bl[113] br[113] wl[511] vdd gnd cell_6t
Xbit_r0_c114 bl[114] br[114] wl[0] vdd gnd cell_6t
Xbit_r1_c114 bl[114] br[114] wl[1] vdd gnd cell_6t
Xbit_r2_c114 bl[114] br[114] wl[2] vdd gnd cell_6t
Xbit_r3_c114 bl[114] br[114] wl[3] vdd gnd cell_6t
Xbit_r4_c114 bl[114] br[114] wl[4] vdd gnd cell_6t
Xbit_r5_c114 bl[114] br[114] wl[5] vdd gnd cell_6t
Xbit_r6_c114 bl[114] br[114] wl[6] vdd gnd cell_6t
Xbit_r7_c114 bl[114] br[114] wl[7] vdd gnd cell_6t
Xbit_r8_c114 bl[114] br[114] wl[8] vdd gnd cell_6t
Xbit_r9_c114 bl[114] br[114] wl[9] vdd gnd cell_6t
Xbit_r10_c114 bl[114] br[114] wl[10] vdd gnd cell_6t
Xbit_r11_c114 bl[114] br[114] wl[11] vdd gnd cell_6t
Xbit_r12_c114 bl[114] br[114] wl[12] vdd gnd cell_6t
Xbit_r13_c114 bl[114] br[114] wl[13] vdd gnd cell_6t
Xbit_r14_c114 bl[114] br[114] wl[14] vdd gnd cell_6t
Xbit_r15_c114 bl[114] br[114] wl[15] vdd gnd cell_6t
Xbit_r16_c114 bl[114] br[114] wl[16] vdd gnd cell_6t
Xbit_r17_c114 bl[114] br[114] wl[17] vdd gnd cell_6t
Xbit_r18_c114 bl[114] br[114] wl[18] vdd gnd cell_6t
Xbit_r19_c114 bl[114] br[114] wl[19] vdd gnd cell_6t
Xbit_r20_c114 bl[114] br[114] wl[20] vdd gnd cell_6t
Xbit_r21_c114 bl[114] br[114] wl[21] vdd gnd cell_6t
Xbit_r22_c114 bl[114] br[114] wl[22] vdd gnd cell_6t
Xbit_r23_c114 bl[114] br[114] wl[23] vdd gnd cell_6t
Xbit_r24_c114 bl[114] br[114] wl[24] vdd gnd cell_6t
Xbit_r25_c114 bl[114] br[114] wl[25] vdd gnd cell_6t
Xbit_r26_c114 bl[114] br[114] wl[26] vdd gnd cell_6t
Xbit_r27_c114 bl[114] br[114] wl[27] vdd gnd cell_6t
Xbit_r28_c114 bl[114] br[114] wl[28] vdd gnd cell_6t
Xbit_r29_c114 bl[114] br[114] wl[29] vdd gnd cell_6t
Xbit_r30_c114 bl[114] br[114] wl[30] vdd gnd cell_6t
Xbit_r31_c114 bl[114] br[114] wl[31] vdd gnd cell_6t
Xbit_r32_c114 bl[114] br[114] wl[32] vdd gnd cell_6t
Xbit_r33_c114 bl[114] br[114] wl[33] vdd gnd cell_6t
Xbit_r34_c114 bl[114] br[114] wl[34] vdd gnd cell_6t
Xbit_r35_c114 bl[114] br[114] wl[35] vdd gnd cell_6t
Xbit_r36_c114 bl[114] br[114] wl[36] vdd gnd cell_6t
Xbit_r37_c114 bl[114] br[114] wl[37] vdd gnd cell_6t
Xbit_r38_c114 bl[114] br[114] wl[38] vdd gnd cell_6t
Xbit_r39_c114 bl[114] br[114] wl[39] vdd gnd cell_6t
Xbit_r40_c114 bl[114] br[114] wl[40] vdd gnd cell_6t
Xbit_r41_c114 bl[114] br[114] wl[41] vdd gnd cell_6t
Xbit_r42_c114 bl[114] br[114] wl[42] vdd gnd cell_6t
Xbit_r43_c114 bl[114] br[114] wl[43] vdd gnd cell_6t
Xbit_r44_c114 bl[114] br[114] wl[44] vdd gnd cell_6t
Xbit_r45_c114 bl[114] br[114] wl[45] vdd gnd cell_6t
Xbit_r46_c114 bl[114] br[114] wl[46] vdd gnd cell_6t
Xbit_r47_c114 bl[114] br[114] wl[47] vdd gnd cell_6t
Xbit_r48_c114 bl[114] br[114] wl[48] vdd gnd cell_6t
Xbit_r49_c114 bl[114] br[114] wl[49] vdd gnd cell_6t
Xbit_r50_c114 bl[114] br[114] wl[50] vdd gnd cell_6t
Xbit_r51_c114 bl[114] br[114] wl[51] vdd gnd cell_6t
Xbit_r52_c114 bl[114] br[114] wl[52] vdd gnd cell_6t
Xbit_r53_c114 bl[114] br[114] wl[53] vdd gnd cell_6t
Xbit_r54_c114 bl[114] br[114] wl[54] vdd gnd cell_6t
Xbit_r55_c114 bl[114] br[114] wl[55] vdd gnd cell_6t
Xbit_r56_c114 bl[114] br[114] wl[56] vdd gnd cell_6t
Xbit_r57_c114 bl[114] br[114] wl[57] vdd gnd cell_6t
Xbit_r58_c114 bl[114] br[114] wl[58] vdd gnd cell_6t
Xbit_r59_c114 bl[114] br[114] wl[59] vdd gnd cell_6t
Xbit_r60_c114 bl[114] br[114] wl[60] vdd gnd cell_6t
Xbit_r61_c114 bl[114] br[114] wl[61] vdd gnd cell_6t
Xbit_r62_c114 bl[114] br[114] wl[62] vdd gnd cell_6t
Xbit_r63_c114 bl[114] br[114] wl[63] vdd gnd cell_6t
Xbit_r64_c114 bl[114] br[114] wl[64] vdd gnd cell_6t
Xbit_r65_c114 bl[114] br[114] wl[65] vdd gnd cell_6t
Xbit_r66_c114 bl[114] br[114] wl[66] vdd gnd cell_6t
Xbit_r67_c114 bl[114] br[114] wl[67] vdd gnd cell_6t
Xbit_r68_c114 bl[114] br[114] wl[68] vdd gnd cell_6t
Xbit_r69_c114 bl[114] br[114] wl[69] vdd gnd cell_6t
Xbit_r70_c114 bl[114] br[114] wl[70] vdd gnd cell_6t
Xbit_r71_c114 bl[114] br[114] wl[71] vdd gnd cell_6t
Xbit_r72_c114 bl[114] br[114] wl[72] vdd gnd cell_6t
Xbit_r73_c114 bl[114] br[114] wl[73] vdd gnd cell_6t
Xbit_r74_c114 bl[114] br[114] wl[74] vdd gnd cell_6t
Xbit_r75_c114 bl[114] br[114] wl[75] vdd gnd cell_6t
Xbit_r76_c114 bl[114] br[114] wl[76] vdd gnd cell_6t
Xbit_r77_c114 bl[114] br[114] wl[77] vdd gnd cell_6t
Xbit_r78_c114 bl[114] br[114] wl[78] vdd gnd cell_6t
Xbit_r79_c114 bl[114] br[114] wl[79] vdd gnd cell_6t
Xbit_r80_c114 bl[114] br[114] wl[80] vdd gnd cell_6t
Xbit_r81_c114 bl[114] br[114] wl[81] vdd gnd cell_6t
Xbit_r82_c114 bl[114] br[114] wl[82] vdd gnd cell_6t
Xbit_r83_c114 bl[114] br[114] wl[83] vdd gnd cell_6t
Xbit_r84_c114 bl[114] br[114] wl[84] vdd gnd cell_6t
Xbit_r85_c114 bl[114] br[114] wl[85] vdd gnd cell_6t
Xbit_r86_c114 bl[114] br[114] wl[86] vdd gnd cell_6t
Xbit_r87_c114 bl[114] br[114] wl[87] vdd gnd cell_6t
Xbit_r88_c114 bl[114] br[114] wl[88] vdd gnd cell_6t
Xbit_r89_c114 bl[114] br[114] wl[89] vdd gnd cell_6t
Xbit_r90_c114 bl[114] br[114] wl[90] vdd gnd cell_6t
Xbit_r91_c114 bl[114] br[114] wl[91] vdd gnd cell_6t
Xbit_r92_c114 bl[114] br[114] wl[92] vdd gnd cell_6t
Xbit_r93_c114 bl[114] br[114] wl[93] vdd gnd cell_6t
Xbit_r94_c114 bl[114] br[114] wl[94] vdd gnd cell_6t
Xbit_r95_c114 bl[114] br[114] wl[95] vdd gnd cell_6t
Xbit_r96_c114 bl[114] br[114] wl[96] vdd gnd cell_6t
Xbit_r97_c114 bl[114] br[114] wl[97] vdd gnd cell_6t
Xbit_r98_c114 bl[114] br[114] wl[98] vdd gnd cell_6t
Xbit_r99_c114 bl[114] br[114] wl[99] vdd gnd cell_6t
Xbit_r100_c114 bl[114] br[114] wl[100] vdd gnd cell_6t
Xbit_r101_c114 bl[114] br[114] wl[101] vdd gnd cell_6t
Xbit_r102_c114 bl[114] br[114] wl[102] vdd gnd cell_6t
Xbit_r103_c114 bl[114] br[114] wl[103] vdd gnd cell_6t
Xbit_r104_c114 bl[114] br[114] wl[104] vdd gnd cell_6t
Xbit_r105_c114 bl[114] br[114] wl[105] vdd gnd cell_6t
Xbit_r106_c114 bl[114] br[114] wl[106] vdd gnd cell_6t
Xbit_r107_c114 bl[114] br[114] wl[107] vdd gnd cell_6t
Xbit_r108_c114 bl[114] br[114] wl[108] vdd gnd cell_6t
Xbit_r109_c114 bl[114] br[114] wl[109] vdd gnd cell_6t
Xbit_r110_c114 bl[114] br[114] wl[110] vdd gnd cell_6t
Xbit_r111_c114 bl[114] br[114] wl[111] vdd gnd cell_6t
Xbit_r112_c114 bl[114] br[114] wl[112] vdd gnd cell_6t
Xbit_r113_c114 bl[114] br[114] wl[113] vdd gnd cell_6t
Xbit_r114_c114 bl[114] br[114] wl[114] vdd gnd cell_6t
Xbit_r115_c114 bl[114] br[114] wl[115] vdd gnd cell_6t
Xbit_r116_c114 bl[114] br[114] wl[116] vdd gnd cell_6t
Xbit_r117_c114 bl[114] br[114] wl[117] vdd gnd cell_6t
Xbit_r118_c114 bl[114] br[114] wl[118] vdd gnd cell_6t
Xbit_r119_c114 bl[114] br[114] wl[119] vdd gnd cell_6t
Xbit_r120_c114 bl[114] br[114] wl[120] vdd gnd cell_6t
Xbit_r121_c114 bl[114] br[114] wl[121] vdd gnd cell_6t
Xbit_r122_c114 bl[114] br[114] wl[122] vdd gnd cell_6t
Xbit_r123_c114 bl[114] br[114] wl[123] vdd gnd cell_6t
Xbit_r124_c114 bl[114] br[114] wl[124] vdd gnd cell_6t
Xbit_r125_c114 bl[114] br[114] wl[125] vdd gnd cell_6t
Xbit_r126_c114 bl[114] br[114] wl[126] vdd gnd cell_6t
Xbit_r127_c114 bl[114] br[114] wl[127] vdd gnd cell_6t
Xbit_r128_c114 bl[114] br[114] wl[128] vdd gnd cell_6t
Xbit_r129_c114 bl[114] br[114] wl[129] vdd gnd cell_6t
Xbit_r130_c114 bl[114] br[114] wl[130] vdd gnd cell_6t
Xbit_r131_c114 bl[114] br[114] wl[131] vdd gnd cell_6t
Xbit_r132_c114 bl[114] br[114] wl[132] vdd gnd cell_6t
Xbit_r133_c114 bl[114] br[114] wl[133] vdd gnd cell_6t
Xbit_r134_c114 bl[114] br[114] wl[134] vdd gnd cell_6t
Xbit_r135_c114 bl[114] br[114] wl[135] vdd gnd cell_6t
Xbit_r136_c114 bl[114] br[114] wl[136] vdd gnd cell_6t
Xbit_r137_c114 bl[114] br[114] wl[137] vdd gnd cell_6t
Xbit_r138_c114 bl[114] br[114] wl[138] vdd gnd cell_6t
Xbit_r139_c114 bl[114] br[114] wl[139] vdd gnd cell_6t
Xbit_r140_c114 bl[114] br[114] wl[140] vdd gnd cell_6t
Xbit_r141_c114 bl[114] br[114] wl[141] vdd gnd cell_6t
Xbit_r142_c114 bl[114] br[114] wl[142] vdd gnd cell_6t
Xbit_r143_c114 bl[114] br[114] wl[143] vdd gnd cell_6t
Xbit_r144_c114 bl[114] br[114] wl[144] vdd gnd cell_6t
Xbit_r145_c114 bl[114] br[114] wl[145] vdd gnd cell_6t
Xbit_r146_c114 bl[114] br[114] wl[146] vdd gnd cell_6t
Xbit_r147_c114 bl[114] br[114] wl[147] vdd gnd cell_6t
Xbit_r148_c114 bl[114] br[114] wl[148] vdd gnd cell_6t
Xbit_r149_c114 bl[114] br[114] wl[149] vdd gnd cell_6t
Xbit_r150_c114 bl[114] br[114] wl[150] vdd gnd cell_6t
Xbit_r151_c114 bl[114] br[114] wl[151] vdd gnd cell_6t
Xbit_r152_c114 bl[114] br[114] wl[152] vdd gnd cell_6t
Xbit_r153_c114 bl[114] br[114] wl[153] vdd gnd cell_6t
Xbit_r154_c114 bl[114] br[114] wl[154] vdd gnd cell_6t
Xbit_r155_c114 bl[114] br[114] wl[155] vdd gnd cell_6t
Xbit_r156_c114 bl[114] br[114] wl[156] vdd gnd cell_6t
Xbit_r157_c114 bl[114] br[114] wl[157] vdd gnd cell_6t
Xbit_r158_c114 bl[114] br[114] wl[158] vdd gnd cell_6t
Xbit_r159_c114 bl[114] br[114] wl[159] vdd gnd cell_6t
Xbit_r160_c114 bl[114] br[114] wl[160] vdd gnd cell_6t
Xbit_r161_c114 bl[114] br[114] wl[161] vdd gnd cell_6t
Xbit_r162_c114 bl[114] br[114] wl[162] vdd gnd cell_6t
Xbit_r163_c114 bl[114] br[114] wl[163] vdd gnd cell_6t
Xbit_r164_c114 bl[114] br[114] wl[164] vdd gnd cell_6t
Xbit_r165_c114 bl[114] br[114] wl[165] vdd gnd cell_6t
Xbit_r166_c114 bl[114] br[114] wl[166] vdd gnd cell_6t
Xbit_r167_c114 bl[114] br[114] wl[167] vdd gnd cell_6t
Xbit_r168_c114 bl[114] br[114] wl[168] vdd gnd cell_6t
Xbit_r169_c114 bl[114] br[114] wl[169] vdd gnd cell_6t
Xbit_r170_c114 bl[114] br[114] wl[170] vdd gnd cell_6t
Xbit_r171_c114 bl[114] br[114] wl[171] vdd gnd cell_6t
Xbit_r172_c114 bl[114] br[114] wl[172] vdd gnd cell_6t
Xbit_r173_c114 bl[114] br[114] wl[173] vdd gnd cell_6t
Xbit_r174_c114 bl[114] br[114] wl[174] vdd gnd cell_6t
Xbit_r175_c114 bl[114] br[114] wl[175] vdd gnd cell_6t
Xbit_r176_c114 bl[114] br[114] wl[176] vdd gnd cell_6t
Xbit_r177_c114 bl[114] br[114] wl[177] vdd gnd cell_6t
Xbit_r178_c114 bl[114] br[114] wl[178] vdd gnd cell_6t
Xbit_r179_c114 bl[114] br[114] wl[179] vdd gnd cell_6t
Xbit_r180_c114 bl[114] br[114] wl[180] vdd gnd cell_6t
Xbit_r181_c114 bl[114] br[114] wl[181] vdd gnd cell_6t
Xbit_r182_c114 bl[114] br[114] wl[182] vdd gnd cell_6t
Xbit_r183_c114 bl[114] br[114] wl[183] vdd gnd cell_6t
Xbit_r184_c114 bl[114] br[114] wl[184] vdd gnd cell_6t
Xbit_r185_c114 bl[114] br[114] wl[185] vdd gnd cell_6t
Xbit_r186_c114 bl[114] br[114] wl[186] vdd gnd cell_6t
Xbit_r187_c114 bl[114] br[114] wl[187] vdd gnd cell_6t
Xbit_r188_c114 bl[114] br[114] wl[188] vdd gnd cell_6t
Xbit_r189_c114 bl[114] br[114] wl[189] vdd gnd cell_6t
Xbit_r190_c114 bl[114] br[114] wl[190] vdd gnd cell_6t
Xbit_r191_c114 bl[114] br[114] wl[191] vdd gnd cell_6t
Xbit_r192_c114 bl[114] br[114] wl[192] vdd gnd cell_6t
Xbit_r193_c114 bl[114] br[114] wl[193] vdd gnd cell_6t
Xbit_r194_c114 bl[114] br[114] wl[194] vdd gnd cell_6t
Xbit_r195_c114 bl[114] br[114] wl[195] vdd gnd cell_6t
Xbit_r196_c114 bl[114] br[114] wl[196] vdd gnd cell_6t
Xbit_r197_c114 bl[114] br[114] wl[197] vdd gnd cell_6t
Xbit_r198_c114 bl[114] br[114] wl[198] vdd gnd cell_6t
Xbit_r199_c114 bl[114] br[114] wl[199] vdd gnd cell_6t
Xbit_r200_c114 bl[114] br[114] wl[200] vdd gnd cell_6t
Xbit_r201_c114 bl[114] br[114] wl[201] vdd gnd cell_6t
Xbit_r202_c114 bl[114] br[114] wl[202] vdd gnd cell_6t
Xbit_r203_c114 bl[114] br[114] wl[203] vdd gnd cell_6t
Xbit_r204_c114 bl[114] br[114] wl[204] vdd gnd cell_6t
Xbit_r205_c114 bl[114] br[114] wl[205] vdd gnd cell_6t
Xbit_r206_c114 bl[114] br[114] wl[206] vdd gnd cell_6t
Xbit_r207_c114 bl[114] br[114] wl[207] vdd gnd cell_6t
Xbit_r208_c114 bl[114] br[114] wl[208] vdd gnd cell_6t
Xbit_r209_c114 bl[114] br[114] wl[209] vdd gnd cell_6t
Xbit_r210_c114 bl[114] br[114] wl[210] vdd gnd cell_6t
Xbit_r211_c114 bl[114] br[114] wl[211] vdd gnd cell_6t
Xbit_r212_c114 bl[114] br[114] wl[212] vdd gnd cell_6t
Xbit_r213_c114 bl[114] br[114] wl[213] vdd gnd cell_6t
Xbit_r214_c114 bl[114] br[114] wl[214] vdd gnd cell_6t
Xbit_r215_c114 bl[114] br[114] wl[215] vdd gnd cell_6t
Xbit_r216_c114 bl[114] br[114] wl[216] vdd gnd cell_6t
Xbit_r217_c114 bl[114] br[114] wl[217] vdd gnd cell_6t
Xbit_r218_c114 bl[114] br[114] wl[218] vdd gnd cell_6t
Xbit_r219_c114 bl[114] br[114] wl[219] vdd gnd cell_6t
Xbit_r220_c114 bl[114] br[114] wl[220] vdd gnd cell_6t
Xbit_r221_c114 bl[114] br[114] wl[221] vdd gnd cell_6t
Xbit_r222_c114 bl[114] br[114] wl[222] vdd gnd cell_6t
Xbit_r223_c114 bl[114] br[114] wl[223] vdd gnd cell_6t
Xbit_r224_c114 bl[114] br[114] wl[224] vdd gnd cell_6t
Xbit_r225_c114 bl[114] br[114] wl[225] vdd gnd cell_6t
Xbit_r226_c114 bl[114] br[114] wl[226] vdd gnd cell_6t
Xbit_r227_c114 bl[114] br[114] wl[227] vdd gnd cell_6t
Xbit_r228_c114 bl[114] br[114] wl[228] vdd gnd cell_6t
Xbit_r229_c114 bl[114] br[114] wl[229] vdd gnd cell_6t
Xbit_r230_c114 bl[114] br[114] wl[230] vdd gnd cell_6t
Xbit_r231_c114 bl[114] br[114] wl[231] vdd gnd cell_6t
Xbit_r232_c114 bl[114] br[114] wl[232] vdd gnd cell_6t
Xbit_r233_c114 bl[114] br[114] wl[233] vdd gnd cell_6t
Xbit_r234_c114 bl[114] br[114] wl[234] vdd gnd cell_6t
Xbit_r235_c114 bl[114] br[114] wl[235] vdd gnd cell_6t
Xbit_r236_c114 bl[114] br[114] wl[236] vdd gnd cell_6t
Xbit_r237_c114 bl[114] br[114] wl[237] vdd gnd cell_6t
Xbit_r238_c114 bl[114] br[114] wl[238] vdd gnd cell_6t
Xbit_r239_c114 bl[114] br[114] wl[239] vdd gnd cell_6t
Xbit_r240_c114 bl[114] br[114] wl[240] vdd gnd cell_6t
Xbit_r241_c114 bl[114] br[114] wl[241] vdd gnd cell_6t
Xbit_r242_c114 bl[114] br[114] wl[242] vdd gnd cell_6t
Xbit_r243_c114 bl[114] br[114] wl[243] vdd gnd cell_6t
Xbit_r244_c114 bl[114] br[114] wl[244] vdd gnd cell_6t
Xbit_r245_c114 bl[114] br[114] wl[245] vdd gnd cell_6t
Xbit_r246_c114 bl[114] br[114] wl[246] vdd gnd cell_6t
Xbit_r247_c114 bl[114] br[114] wl[247] vdd gnd cell_6t
Xbit_r248_c114 bl[114] br[114] wl[248] vdd gnd cell_6t
Xbit_r249_c114 bl[114] br[114] wl[249] vdd gnd cell_6t
Xbit_r250_c114 bl[114] br[114] wl[250] vdd gnd cell_6t
Xbit_r251_c114 bl[114] br[114] wl[251] vdd gnd cell_6t
Xbit_r252_c114 bl[114] br[114] wl[252] vdd gnd cell_6t
Xbit_r253_c114 bl[114] br[114] wl[253] vdd gnd cell_6t
Xbit_r254_c114 bl[114] br[114] wl[254] vdd gnd cell_6t
Xbit_r255_c114 bl[114] br[114] wl[255] vdd gnd cell_6t
Xbit_r256_c114 bl[114] br[114] wl[256] vdd gnd cell_6t
Xbit_r257_c114 bl[114] br[114] wl[257] vdd gnd cell_6t
Xbit_r258_c114 bl[114] br[114] wl[258] vdd gnd cell_6t
Xbit_r259_c114 bl[114] br[114] wl[259] vdd gnd cell_6t
Xbit_r260_c114 bl[114] br[114] wl[260] vdd gnd cell_6t
Xbit_r261_c114 bl[114] br[114] wl[261] vdd gnd cell_6t
Xbit_r262_c114 bl[114] br[114] wl[262] vdd gnd cell_6t
Xbit_r263_c114 bl[114] br[114] wl[263] vdd gnd cell_6t
Xbit_r264_c114 bl[114] br[114] wl[264] vdd gnd cell_6t
Xbit_r265_c114 bl[114] br[114] wl[265] vdd gnd cell_6t
Xbit_r266_c114 bl[114] br[114] wl[266] vdd gnd cell_6t
Xbit_r267_c114 bl[114] br[114] wl[267] vdd gnd cell_6t
Xbit_r268_c114 bl[114] br[114] wl[268] vdd gnd cell_6t
Xbit_r269_c114 bl[114] br[114] wl[269] vdd gnd cell_6t
Xbit_r270_c114 bl[114] br[114] wl[270] vdd gnd cell_6t
Xbit_r271_c114 bl[114] br[114] wl[271] vdd gnd cell_6t
Xbit_r272_c114 bl[114] br[114] wl[272] vdd gnd cell_6t
Xbit_r273_c114 bl[114] br[114] wl[273] vdd gnd cell_6t
Xbit_r274_c114 bl[114] br[114] wl[274] vdd gnd cell_6t
Xbit_r275_c114 bl[114] br[114] wl[275] vdd gnd cell_6t
Xbit_r276_c114 bl[114] br[114] wl[276] vdd gnd cell_6t
Xbit_r277_c114 bl[114] br[114] wl[277] vdd gnd cell_6t
Xbit_r278_c114 bl[114] br[114] wl[278] vdd gnd cell_6t
Xbit_r279_c114 bl[114] br[114] wl[279] vdd gnd cell_6t
Xbit_r280_c114 bl[114] br[114] wl[280] vdd gnd cell_6t
Xbit_r281_c114 bl[114] br[114] wl[281] vdd gnd cell_6t
Xbit_r282_c114 bl[114] br[114] wl[282] vdd gnd cell_6t
Xbit_r283_c114 bl[114] br[114] wl[283] vdd gnd cell_6t
Xbit_r284_c114 bl[114] br[114] wl[284] vdd gnd cell_6t
Xbit_r285_c114 bl[114] br[114] wl[285] vdd gnd cell_6t
Xbit_r286_c114 bl[114] br[114] wl[286] vdd gnd cell_6t
Xbit_r287_c114 bl[114] br[114] wl[287] vdd gnd cell_6t
Xbit_r288_c114 bl[114] br[114] wl[288] vdd gnd cell_6t
Xbit_r289_c114 bl[114] br[114] wl[289] vdd gnd cell_6t
Xbit_r290_c114 bl[114] br[114] wl[290] vdd gnd cell_6t
Xbit_r291_c114 bl[114] br[114] wl[291] vdd gnd cell_6t
Xbit_r292_c114 bl[114] br[114] wl[292] vdd gnd cell_6t
Xbit_r293_c114 bl[114] br[114] wl[293] vdd gnd cell_6t
Xbit_r294_c114 bl[114] br[114] wl[294] vdd gnd cell_6t
Xbit_r295_c114 bl[114] br[114] wl[295] vdd gnd cell_6t
Xbit_r296_c114 bl[114] br[114] wl[296] vdd gnd cell_6t
Xbit_r297_c114 bl[114] br[114] wl[297] vdd gnd cell_6t
Xbit_r298_c114 bl[114] br[114] wl[298] vdd gnd cell_6t
Xbit_r299_c114 bl[114] br[114] wl[299] vdd gnd cell_6t
Xbit_r300_c114 bl[114] br[114] wl[300] vdd gnd cell_6t
Xbit_r301_c114 bl[114] br[114] wl[301] vdd gnd cell_6t
Xbit_r302_c114 bl[114] br[114] wl[302] vdd gnd cell_6t
Xbit_r303_c114 bl[114] br[114] wl[303] vdd gnd cell_6t
Xbit_r304_c114 bl[114] br[114] wl[304] vdd gnd cell_6t
Xbit_r305_c114 bl[114] br[114] wl[305] vdd gnd cell_6t
Xbit_r306_c114 bl[114] br[114] wl[306] vdd gnd cell_6t
Xbit_r307_c114 bl[114] br[114] wl[307] vdd gnd cell_6t
Xbit_r308_c114 bl[114] br[114] wl[308] vdd gnd cell_6t
Xbit_r309_c114 bl[114] br[114] wl[309] vdd gnd cell_6t
Xbit_r310_c114 bl[114] br[114] wl[310] vdd gnd cell_6t
Xbit_r311_c114 bl[114] br[114] wl[311] vdd gnd cell_6t
Xbit_r312_c114 bl[114] br[114] wl[312] vdd gnd cell_6t
Xbit_r313_c114 bl[114] br[114] wl[313] vdd gnd cell_6t
Xbit_r314_c114 bl[114] br[114] wl[314] vdd gnd cell_6t
Xbit_r315_c114 bl[114] br[114] wl[315] vdd gnd cell_6t
Xbit_r316_c114 bl[114] br[114] wl[316] vdd gnd cell_6t
Xbit_r317_c114 bl[114] br[114] wl[317] vdd gnd cell_6t
Xbit_r318_c114 bl[114] br[114] wl[318] vdd gnd cell_6t
Xbit_r319_c114 bl[114] br[114] wl[319] vdd gnd cell_6t
Xbit_r320_c114 bl[114] br[114] wl[320] vdd gnd cell_6t
Xbit_r321_c114 bl[114] br[114] wl[321] vdd gnd cell_6t
Xbit_r322_c114 bl[114] br[114] wl[322] vdd gnd cell_6t
Xbit_r323_c114 bl[114] br[114] wl[323] vdd gnd cell_6t
Xbit_r324_c114 bl[114] br[114] wl[324] vdd gnd cell_6t
Xbit_r325_c114 bl[114] br[114] wl[325] vdd gnd cell_6t
Xbit_r326_c114 bl[114] br[114] wl[326] vdd gnd cell_6t
Xbit_r327_c114 bl[114] br[114] wl[327] vdd gnd cell_6t
Xbit_r328_c114 bl[114] br[114] wl[328] vdd gnd cell_6t
Xbit_r329_c114 bl[114] br[114] wl[329] vdd gnd cell_6t
Xbit_r330_c114 bl[114] br[114] wl[330] vdd gnd cell_6t
Xbit_r331_c114 bl[114] br[114] wl[331] vdd gnd cell_6t
Xbit_r332_c114 bl[114] br[114] wl[332] vdd gnd cell_6t
Xbit_r333_c114 bl[114] br[114] wl[333] vdd gnd cell_6t
Xbit_r334_c114 bl[114] br[114] wl[334] vdd gnd cell_6t
Xbit_r335_c114 bl[114] br[114] wl[335] vdd gnd cell_6t
Xbit_r336_c114 bl[114] br[114] wl[336] vdd gnd cell_6t
Xbit_r337_c114 bl[114] br[114] wl[337] vdd gnd cell_6t
Xbit_r338_c114 bl[114] br[114] wl[338] vdd gnd cell_6t
Xbit_r339_c114 bl[114] br[114] wl[339] vdd gnd cell_6t
Xbit_r340_c114 bl[114] br[114] wl[340] vdd gnd cell_6t
Xbit_r341_c114 bl[114] br[114] wl[341] vdd gnd cell_6t
Xbit_r342_c114 bl[114] br[114] wl[342] vdd gnd cell_6t
Xbit_r343_c114 bl[114] br[114] wl[343] vdd gnd cell_6t
Xbit_r344_c114 bl[114] br[114] wl[344] vdd gnd cell_6t
Xbit_r345_c114 bl[114] br[114] wl[345] vdd gnd cell_6t
Xbit_r346_c114 bl[114] br[114] wl[346] vdd gnd cell_6t
Xbit_r347_c114 bl[114] br[114] wl[347] vdd gnd cell_6t
Xbit_r348_c114 bl[114] br[114] wl[348] vdd gnd cell_6t
Xbit_r349_c114 bl[114] br[114] wl[349] vdd gnd cell_6t
Xbit_r350_c114 bl[114] br[114] wl[350] vdd gnd cell_6t
Xbit_r351_c114 bl[114] br[114] wl[351] vdd gnd cell_6t
Xbit_r352_c114 bl[114] br[114] wl[352] vdd gnd cell_6t
Xbit_r353_c114 bl[114] br[114] wl[353] vdd gnd cell_6t
Xbit_r354_c114 bl[114] br[114] wl[354] vdd gnd cell_6t
Xbit_r355_c114 bl[114] br[114] wl[355] vdd gnd cell_6t
Xbit_r356_c114 bl[114] br[114] wl[356] vdd gnd cell_6t
Xbit_r357_c114 bl[114] br[114] wl[357] vdd gnd cell_6t
Xbit_r358_c114 bl[114] br[114] wl[358] vdd gnd cell_6t
Xbit_r359_c114 bl[114] br[114] wl[359] vdd gnd cell_6t
Xbit_r360_c114 bl[114] br[114] wl[360] vdd gnd cell_6t
Xbit_r361_c114 bl[114] br[114] wl[361] vdd gnd cell_6t
Xbit_r362_c114 bl[114] br[114] wl[362] vdd gnd cell_6t
Xbit_r363_c114 bl[114] br[114] wl[363] vdd gnd cell_6t
Xbit_r364_c114 bl[114] br[114] wl[364] vdd gnd cell_6t
Xbit_r365_c114 bl[114] br[114] wl[365] vdd gnd cell_6t
Xbit_r366_c114 bl[114] br[114] wl[366] vdd gnd cell_6t
Xbit_r367_c114 bl[114] br[114] wl[367] vdd gnd cell_6t
Xbit_r368_c114 bl[114] br[114] wl[368] vdd gnd cell_6t
Xbit_r369_c114 bl[114] br[114] wl[369] vdd gnd cell_6t
Xbit_r370_c114 bl[114] br[114] wl[370] vdd gnd cell_6t
Xbit_r371_c114 bl[114] br[114] wl[371] vdd gnd cell_6t
Xbit_r372_c114 bl[114] br[114] wl[372] vdd gnd cell_6t
Xbit_r373_c114 bl[114] br[114] wl[373] vdd gnd cell_6t
Xbit_r374_c114 bl[114] br[114] wl[374] vdd gnd cell_6t
Xbit_r375_c114 bl[114] br[114] wl[375] vdd gnd cell_6t
Xbit_r376_c114 bl[114] br[114] wl[376] vdd gnd cell_6t
Xbit_r377_c114 bl[114] br[114] wl[377] vdd gnd cell_6t
Xbit_r378_c114 bl[114] br[114] wl[378] vdd gnd cell_6t
Xbit_r379_c114 bl[114] br[114] wl[379] vdd gnd cell_6t
Xbit_r380_c114 bl[114] br[114] wl[380] vdd gnd cell_6t
Xbit_r381_c114 bl[114] br[114] wl[381] vdd gnd cell_6t
Xbit_r382_c114 bl[114] br[114] wl[382] vdd gnd cell_6t
Xbit_r383_c114 bl[114] br[114] wl[383] vdd gnd cell_6t
Xbit_r384_c114 bl[114] br[114] wl[384] vdd gnd cell_6t
Xbit_r385_c114 bl[114] br[114] wl[385] vdd gnd cell_6t
Xbit_r386_c114 bl[114] br[114] wl[386] vdd gnd cell_6t
Xbit_r387_c114 bl[114] br[114] wl[387] vdd gnd cell_6t
Xbit_r388_c114 bl[114] br[114] wl[388] vdd gnd cell_6t
Xbit_r389_c114 bl[114] br[114] wl[389] vdd gnd cell_6t
Xbit_r390_c114 bl[114] br[114] wl[390] vdd gnd cell_6t
Xbit_r391_c114 bl[114] br[114] wl[391] vdd gnd cell_6t
Xbit_r392_c114 bl[114] br[114] wl[392] vdd gnd cell_6t
Xbit_r393_c114 bl[114] br[114] wl[393] vdd gnd cell_6t
Xbit_r394_c114 bl[114] br[114] wl[394] vdd gnd cell_6t
Xbit_r395_c114 bl[114] br[114] wl[395] vdd gnd cell_6t
Xbit_r396_c114 bl[114] br[114] wl[396] vdd gnd cell_6t
Xbit_r397_c114 bl[114] br[114] wl[397] vdd gnd cell_6t
Xbit_r398_c114 bl[114] br[114] wl[398] vdd gnd cell_6t
Xbit_r399_c114 bl[114] br[114] wl[399] vdd gnd cell_6t
Xbit_r400_c114 bl[114] br[114] wl[400] vdd gnd cell_6t
Xbit_r401_c114 bl[114] br[114] wl[401] vdd gnd cell_6t
Xbit_r402_c114 bl[114] br[114] wl[402] vdd gnd cell_6t
Xbit_r403_c114 bl[114] br[114] wl[403] vdd gnd cell_6t
Xbit_r404_c114 bl[114] br[114] wl[404] vdd gnd cell_6t
Xbit_r405_c114 bl[114] br[114] wl[405] vdd gnd cell_6t
Xbit_r406_c114 bl[114] br[114] wl[406] vdd gnd cell_6t
Xbit_r407_c114 bl[114] br[114] wl[407] vdd gnd cell_6t
Xbit_r408_c114 bl[114] br[114] wl[408] vdd gnd cell_6t
Xbit_r409_c114 bl[114] br[114] wl[409] vdd gnd cell_6t
Xbit_r410_c114 bl[114] br[114] wl[410] vdd gnd cell_6t
Xbit_r411_c114 bl[114] br[114] wl[411] vdd gnd cell_6t
Xbit_r412_c114 bl[114] br[114] wl[412] vdd gnd cell_6t
Xbit_r413_c114 bl[114] br[114] wl[413] vdd gnd cell_6t
Xbit_r414_c114 bl[114] br[114] wl[414] vdd gnd cell_6t
Xbit_r415_c114 bl[114] br[114] wl[415] vdd gnd cell_6t
Xbit_r416_c114 bl[114] br[114] wl[416] vdd gnd cell_6t
Xbit_r417_c114 bl[114] br[114] wl[417] vdd gnd cell_6t
Xbit_r418_c114 bl[114] br[114] wl[418] vdd gnd cell_6t
Xbit_r419_c114 bl[114] br[114] wl[419] vdd gnd cell_6t
Xbit_r420_c114 bl[114] br[114] wl[420] vdd gnd cell_6t
Xbit_r421_c114 bl[114] br[114] wl[421] vdd gnd cell_6t
Xbit_r422_c114 bl[114] br[114] wl[422] vdd gnd cell_6t
Xbit_r423_c114 bl[114] br[114] wl[423] vdd gnd cell_6t
Xbit_r424_c114 bl[114] br[114] wl[424] vdd gnd cell_6t
Xbit_r425_c114 bl[114] br[114] wl[425] vdd gnd cell_6t
Xbit_r426_c114 bl[114] br[114] wl[426] vdd gnd cell_6t
Xbit_r427_c114 bl[114] br[114] wl[427] vdd gnd cell_6t
Xbit_r428_c114 bl[114] br[114] wl[428] vdd gnd cell_6t
Xbit_r429_c114 bl[114] br[114] wl[429] vdd gnd cell_6t
Xbit_r430_c114 bl[114] br[114] wl[430] vdd gnd cell_6t
Xbit_r431_c114 bl[114] br[114] wl[431] vdd gnd cell_6t
Xbit_r432_c114 bl[114] br[114] wl[432] vdd gnd cell_6t
Xbit_r433_c114 bl[114] br[114] wl[433] vdd gnd cell_6t
Xbit_r434_c114 bl[114] br[114] wl[434] vdd gnd cell_6t
Xbit_r435_c114 bl[114] br[114] wl[435] vdd gnd cell_6t
Xbit_r436_c114 bl[114] br[114] wl[436] vdd gnd cell_6t
Xbit_r437_c114 bl[114] br[114] wl[437] vdd gnd cell_6t
Xbit_r438_c114 bl[114] br[114] wl[438] vdd gnd cell_6t
Xbit_r439_c114 bl[114] br[114] wl[439] vdd gnd cell_6t
Xbit_r440_c114 bl[114] br[114] wl[440] vdd gnd cell_6t
Xbit_r441_c114 bl[114] br[114] wl[441] vdd gnd cell_6t
Xbit_r442_c114 bl[114] br[114] wl[442] vdd gnd cell_6t
Xbit_r443_c114 bl[114] br[114] wl[443] vdd gnd cell_6t
Xbit_r444_c114 bl[114] br[114] wl[444] vdd gnd cell_6t
Xbit_r445_c114 bl[114] br[114] wl[445] vdd gnd cell_6t
Xbit_r446_c114 bl[114] br[114] wl[446] vdd gnd cell_6t
Xbit_r447_c114 bl[114] br[114] wl[447] vdd gnd cell_6t
Xbit_r448_c114 bl[114] br[114] wl[448] vdd gnd cell_6t
Xbit_r449_c114 bl[114] br[114] wl[449] vdd gnd cell_6t
Xbit_r450_c114 bl[114] br[114] wl[450] vdd gnd cell_6t
Xbit_r451_c114 bl[114] br[114] wl[451] vdd gnd cell_6t
Xbit_r452_c114 bl[114] br[114] wl[452] vdd gnd cell_6t
Xbit_r453_c114 bl[114] br[114] wl[453] vdd gnd cell_6t
Xbit_r454_c114 bl[114] br[114] wl[454] vdd gnd cell_6t
Xbit_r455_c114 bl[114] br[114] wl[455] vdd gnd cell_6t
Xbit_r456_c114 bl[114] br[114] wl[456] vdd gnd cell_6t
Xbit_r457_c114 bl[114] br[114] wl[457] vdd gnd cell_6t
Xbit_r458_c114 bl[114] br[114] wl[458] vdd gnd cell_6t
Xbit_r459_c114 bl[114] br[114] wl[459] vdd gnd cell_6t
Xbit_r460_c114 bl[114] br[114] wl[460] vdd gnd cell_6t
Xbit_r461_c114 bl[114] br[114] wl[461] vdd gnd cell_6t
Xbit_r462_c114 bl[114] br[114] wl[462] vdd gnd cell_6t
Xbit_r463_c114 bl[114] br[114] wl[463] vdd gnd cell_6t
Xbit_r464_c114 bl[114] br[114] wl[464] vdd gnd cell_6t
Xbit_r465_c114 bl[114] br[114] wl[465] vdd gnd cell_6t
Xbit_r466_c114 bl[114] br[114] wl[466] vdd gnd cell_6t
Xbit_r467_c114 bl[114] br[114] wl[467] vdd gnd cell_6t
Xbit_r468_c114 bl[114] br[114] wl[468] vdd gnd cell_6t
Xbit_r469_c114 bl[114] br[114] wl[469] vdd gnd cell_6t
Xbit_r470_c114 bl[114] br[114] wl[470] vdd gnd cell_6t
Xbit_r471_c114 bl[114] br[114] wl[471] vdd gnd cell_6t
Xbit_r472_c114 bl[114] br[114] wl[472] vdd gnd cell_6t
Xbit_r473_c114 bl[114] br[114] wl[473] vdd gnd cell_6t
Xbit_r474_c114 bl[114] br[114] wl[474] vdd gnd cell_6t
Xbit_r475_c114 bl[114] br[114] wl[475] vdd gnd cell_6t
Xbit_r476_c114 bl[114] br[114] wl[476] vdd gnd cell_6t
Xbit_r477_c114 bl[114] br[114] wl[477] vdd gnd cell_6t
Xbit_r478_c114 bl[114] br[114] wl[478] vdd gnd cell_6t
Xbit_r479_c114 bl[114] br[114] wl[479] vdd gnd cell_6t
Xbit_r480_c114 bl[114] br[114] wl[480] vdd gnd cell_6t
Xbit_r481_c114 bl[114] br[114] wl[481] vdd gnd cell_6t
Xbit_r482_c114 bl[114] br[114] wl[482] vdd gnd cell_6t
Xbit_r483_c114 bl[114] br[114] wl[483] vdd gnd cell_6t
Xbit_r484_c114 bl[114] br[114] wl[484] vdd gnd cell_6t
Xbit_r485_c114 bl[114] br[114] wl[485] vdd gnd cell_6t
Xbit_r486_c114 bl[114] br[114] wl[486] vdd gnd cell_6t
Xbit_r487_c114 bl[114] br[114] wl[487] vdd gnd cell_6t
Xbit_r488_c114 bl[114] br[114] wl[488] vdd gnd cell_6t
Xbit_r489_c114 bl[114] br[114] wl[489] vdd gnd cell_6t
Xbit_r490_c114 bl[114] br[114] wl[490] vdd gnd cell_6t
Xbit_r491_c114 bl[114] br[114] wl[491] vdd gnd cell_6t
Xbit_r492_c114 bl[114] br[114] wl[492] vdd gnd cell_6t
Xbit_r493_c114 bl[114] br[114] wl[493] vdd gnd cell_6t
Xbit_r494_c114 bl[114] br[114] wl[494] vdd gnd cell_6t
Xbit_r495_c114 bl[114] br[114] wl[495] vdd gnd cell_6t
Xbit_r496_c114 bl[114] br[114] wl[496] vdd gnd cell_6t
Xbit_r497_c114 bl[114] br[114] wl[497] vdd gnd cell_6t
Xbit_r498_c114 bl[114] br[114] wl[498] vdd gnd cell_6t
Xbit_r499_c114 bl[114] br[114] wl[499] vdd gnd cell_6t
Xbit_r500_c114 bl[114] br[114] wl[500] vdd gnd cell_6t
Xbit_r501_c114 bl[114] br[114] wl[501] vdd gnd cell_6t
Xbit_r502_c114 bl[114] br[114] wl[502] vdd gnd cell_6t
Xbit_r503_c114 bl[114] br[114] wl[503] vdd gnd cell_6t
Xbit_r504_c114 bl[114] br[114] wl[504] vdd gnd cell_6t
Xbit_r505_c114 bl[114] br[114] wl[505] vdd gnd cell_6t
Xbit_r506_c114 bl[114] br[114] wl[506] vdd gnd cell_6t
Xbit_r507_c114 bl[114] br[114] wl[507] vdd gnd cell_6t
Xbit_r508_c114 bl[114] br[114] wl[508] vdd gnd cell_6t
Xbit_r509_c114 bl[114] br[114] wl[509] vdd gnd cell_6t
Xbit_r510_c114 bl[114] br[114] wl[510] vdd gnd cell_6t
Xbit_r511_c114 bl[114] br[114] wl[511] vdd gnd cell_6t
Xbit_r0_c115 bl[115] br[115] wl[0] vdd gnd cell_6t
Xbit_r1_c115 bl[115] br[115] wl[1] vdd gnd cell_6t
Xbit_r2_c115 bl[115] br[115] wl[2] vdd gnd cell_6t
Xbit_r3_c115 bl[115] br[115] wl[3] vdd gnd cell_6t
Xbit_r4_c115 bl[115] br[115] wl[4] vdd gnd cell_6t
Xbit_r5_c115 bl[115] br[115] wl[5] vdd gnd cell_6t
Xbit_r6_c115 bl[115] br[115] wl[6] vdd gnd cell_6t
Xbit_r7_c115 bl[115] br[115] wl[7] vdd gnd cell_6t
Xbit_r8_c115 bl[115] br[115] wl[8] vdd gnd cell_6t
Xbit_r9_c115 bl[115] br[115] wl[9] vdd gnd cell_6t
Xbit_r10_c115 bl[115] br[115] wl[10] vdd gnd cell_6t
Xbit_r11_c115 bl[115] br[115] wl[11] vdd gnd cell_6t
Xbit_r12_c115 bl[115] br[115] wl[12] vdd gnd cell_6t
Xbit_r13_c115 bl[115] br[115] wl[13] vdd gnd cell_6t
Xbit_r14_c115 bl[115] br[115] wl[14] vdd gnd cell_6t
Xbit_r15_c115 bl[115] br[115] wl[15] vdd gnd cell_6t
Xbit_r16_c115 bl[115] br[115] wl[16] vdd gnd cell_6t
Xbit_r17_c115 bl[115] br[115] wl[17] vdd gnd cell_6t
Xbit_r18_c115 bl[115] br[115] wl[18] vdd gnd cell_6t
Xbit_r19_c115 bl[115] br[115] wl[19] vdd gnd cell_6t
Xbit_r20_c115 bl[115] br[115] wl[20] vdd gnd cell_6t
Xbit_r21_c115 bl[115] br[115] wl[21] vdd gnd cell_6t
Xbit_r22_c115 bl[115] br[115] wl[22] vdd gnd cell_6t
Xbit_r23_c115 bl[115] br[115] wl[23] vdd gnd cell_6t
Xbit_r24_c115 bl[115] br[115] wl[24] vdd gnd cell_6t
Xbit_r25_c115 bl[115] br[115] wl[25] vdd gnd cell_6t
Xbit_r26_c115 bl[115] br[115] wl[26] vdd gnd cell_6t
Xbit_r27_c115 bl[115] br[115] wl[27] vdd gnd cell_6t
Xbit_r28_c115 bl[115] br[115] wl[28] vdd gnd cell_6t
Xbit_r29_c115 bl[115] br[115] wl[29] vdd gnd cell_6t
Xbit_r30_c115 bl[115] br[115] wl[30] vdd gnd cell_6t
Xbit_r31_c115 bl[115] br[115] wl[31] vdd gnd cell_6t
Xbit_r32_c115 bl[115] br[115] wl[32] vdd gnd cell_6t
Xbit_r33_c115 bl[115] br[115] wl[33] vdd gnd cell_6t
Xbit_r34_c115 bl[115] br[115] wl[34] vdd gnd cell_6t
Xbit_r35_c115 bl[115] br[115] wl[35] vdd gnd cell_6t
Xbit_r36_c115 bl[115] br[115] wl[36] vdd gnd cell_6t
Xbit_r37_c115 bl[115] br[115] wl[37] vdd gnd cell_6t
Xbit_r38_c115 bl[115] br[115] wl[38] vdd gnd cell_6t
Xbit_r39_c115 bl[115] br[115] wl[39] vdd gnd cell_6t
Xbit_r40_c115 bl[115] br[115] wl[40] vdd gnd cell_6t
Xbit_r41_c115 bl[115] br[115] wl[41] vdd gnd cell_6t
Xbit_r42_c115 bl[115] br[115] wl[42] vdd gnd cell_6t
Xbit_r43_c115 bl[115] br[115] wl[43] vdd gnd cell_6t
Xbit_r44_c115 bl[115] br[115] wl[44] vdd gnd cell_6t
Xbit_r45_c115 bl[115] br[115] wl[45] vdd gnd cell_6t
Xbit_r46_c115 bl[115] br[115] wl[46] vdd gnd cell_6t
Xbit_r47_c115 bl[115] br[115] wl[47] vdd gnd cell_6t
Xbit_r48_c115 bl[115] br[115] wl[48] vdd gnd cell_6t
Xbit_r49_c115 bl[115] br[115] wl[49] vdd gnd cell_6t
Xbit_r50_c115 bl[115] br[115] wl[50] vdd gnd cell_6t
Xbit_r51_c115 bl[115] br[115] wl[51] vdd gnd cell_6t
Xbit_r52_c115 bl[115] br[115] wl[52] vdd gnd cell_6t
Xbit_r53_c115 bl[115] br[115] wl[53] vdd gnd cell_6t
Xbit_r54_c115 bl[115] br[115] wl[54] vdd gnd cell_6t
Xbit_r55_c115 bl[115] br[115] wl[55] vdd gnd cell_6t
Xbit_r56_c115 bl[115] br[115] wl[56] vdd gnd cell_6t
Xbit_r57_c115 bl[115] br[115] wl[57] vdd gnd cell_6t
Xbit_r58_c115 bl[115] br[115] wl[58] vdd gnd cell_6t
Xbit_r59_c115 bl[115] br[115] wl[59] vdd gnd cell_6t
Xbit_r60_c115 bl[115] br[115] wl[60] vdd gnd cell_6t
Xbit_r61_c115 bl[115] br[115] wl[61] vdd gnd cell_6t
Xbit_r62_c115 bl[115] br[115] wl[62] vdd gnd cell_6t
Xbit_r63_c115 bl[115] br[115] wl[63] vdd gnd cell_6t
Xbit_r64_c115 bl[115] br[115] wl[64] vdd gnd cell_6t
Xbit_r65_c115 bl[115] br[115] wl[65] vdd gnd cell_6t
Xbit_r66_c115 bl[115] br[115] wl[66] vdd gnd cell_6t
Xbit_r67_c115 bl[115] br[115] wl[67] vdd gnd cell_6t
Xbit_r68_c115 bl[115] br[115] wl[68] vdd gnd cell_6t
Xbit_r69_c115 bl[115] br[115] wl[69] vdd gnd cell_6t
Xbit_r70_c115 bl[115] br[115] wl[70] vdd gnd cell_6t
Xbit_r71_c115 bl[115] br[115] wl[71] vdd gnd cell_6t
Xbit_r72_c115 bl[115] br[115] wl[72] vdd gnd cell_6t
Xbit_r73_c115 bl[115] br[115] wl[73] vdd gnd cell_6t
Xbit_r74_c115 bl[115] br[115] wl[74] vdd gnd cell_6t
Xbit_r75_c115 bl[115] br[115] wl[75] vdd gnd cell_6t
Xbit_r76_c115 bl[115] br[115] wl[76] vdd gnd cell_6t
Xbit_r77_c115 bl[115] br[115] wl[77] vdd gnd cell_6t
Xbit_r78_c115 bl[115] br[115] wl[78] vdd gnd cell_6t
Xbit_r79_c115 bl[115] br[115] wl[79] vdd gnd cell_6t
Xbit_r80_c115 bl[115] br[115] wl[80] vdd gnd cell_6t
Xbit_r81_c115 bl[115] br[115] wl[81] vdd gnd cell_6t
Xbit_r82_c115 bl[115] br[115] wl[82] vdd gnd cell_6t
Xbit_r83_c115 bl[115] br[115] wl[83] vdd gnd cell_6t
Xbit_r84_c115 bl[115] br[115] wl[84] vdd gnd cell_6t
Xbit_r85_c115 bl[115] br[115] wl[85] vdd gnd cell_6t
Xbit_r86_c115 bl[115] br[115] wl[86] vdd gnd cell_6t
Xbit_r87_c115 bl[115] br[115] wl[87] vdd gnd cell_6t
Xbit_r88_c115 bl[115] br[115] wl[88] vdd gnd cell_6t
Xbit_r89_c115 bl[115] br[115] wl[89] vdd gnd cell_6t
Xbit_r90_c115 bl[115] br[115] wl[90] vdd gnd cell_6t
Xbit_r91_c115 bl[115] br[115] wl[91] vdd gnd cell_6t
Xbit_r92_c115 bl[115] br[115] wl[92] vdd gnd cell_6t
Xbit_r93_c115 bl[115] br[115] wl[93] vdd gnd cell_6t
Xbit_r94_c115 bl[115] br[115] wl[94] vdd gnd cell_6t
Xbit_r95_c115 bl[115] br[115] wl[95] vdd gnd cell_6t
Xbit_r96_c115 bl[115] br[115] wl[96] vdd gnd cell_6t
Xbit_r97_c115 bl[115] br[115] wl[97] vdd gnd cell_6t
Xbit_r98_c115 bl[115] br[115] wl[98] vdd gnd cell_6t
Xbit_r99_c115 bl[115] br[115] wl[99] vdd gnd cell_6t
Xbit_r100_c115 bl[115] br[115] wl[100] vdd gnd cell_6t
Xbit_r101_c115 bl[115] br[115] wl[101] vdd gnd cell_6t
Xbit_r102_c115 bl[115] br[115] wl[102] vdd gnd cell_6t
Xbit_r103_c115 bl[115] br[115] wl[103] vdd gnd cell_6t
Xbit_r104_c115 bl[115] br[115] wl[104] vdd gnd cell_6t
Xbit_r105_c115 bl[115] br[115] wl[105] vdd gnd cell_6t
Xbit_r106_c115 bl[115] br[115] wl[106] vdd gnd cell_6t
Xbit_r107_c115 bl[115] br[115] wl[107] vdd gnd cell_6t
Xbit_r108_c115 bl[115] br[115] wl[108] vdd gnd cell_6t
Xbit_r109_c115 bl[115] br[115] wl[109] vdd gnd cell_6t
Xbit_r110_c115 bl[115] br[115] wl[110] vdd gnd cell_6t
Xbit_r111_c115 bl[115] br[115] wl[111] vdd gnd cell_6t
Xbit_r112_c115 bl[115] br[115] wl[112] vdd gnd cell_6t
Xbit_r113_c115 bl[115] br[115] wl[113] vdd gnd cell_6t
Xbit_r114_c115 bl[115] br[115] wl[114] vdd gnd cell_6t
Xbit_r115_c115 bl[115] br[115] wl[115] vdd gnd cell_6t
Xbit_r116_c115 bl[115] br[115] wl[116] vdd gnd cell_6t
Xbit_r117_c115 bl[115] br[115] wl[117] vdd gnd cell_6t
Xbit_r118_c115 bl[115] br[115] wl[118] vdd gnd cell_6t
Xbit_r119_c115 bl[115] br[115] wl[119] vdd gnd cell_6t
Xbit_r120_c115 bl[115] br[115] wl[120] vdd gnd cell_6t
Xbit_r121_c115 bl[115] br[115] wl[121] vdd gnd cell_6t
Xbit_r122_c115 bl[115] br[115] wl[122] vdd gnd cell_6t
Xbit_r123_c115 bl[115] br[115] wl[123] vdd gnd cell_6t
Xbit_r124_c115 bl[115] br[115] wl[124] vdd gnd cell_6t
Xbit_r125_c115 bl[115] br[115] wl[125] vdd gnd cell_6t
Xbit_r126_c115 bl[115] br[115] wl[126] vdd gnd cell_6t
Xbit_r127_c115 bl[115] br[115] wl[127] vdd gnd cell_6t
Xbit_r128_c115 bl[115] br[115] wl[128] vdd gnd cell_6t
Xbit_r129_c115 bl[115] br[115] wl[129] vdd gnd cell_6t
Xbit_r130_c115 bl[115] br[115] wl[130] vdd gnd cell_6t
Xbit_r131_c115 bl[115] br[115] wl[131] vdd gnd cell_6t
Xbit_r132_c115 bl[115] br[115] wl[132] vdd gnd cell_6t
Xbit_r133_c115 bl[115] br[115] wl[133] vdd gnd cell_6t
Xbit_r134_c115 bl[115] br[115] wl[134] vdd gnd cell_6t
Xbit_r135_c115 bl[115] br[115] wl[135] vdd gnd cell_6t
Xbit_r136_c115 bl[115] br[115] wl[136] vdd gnd cell_6t
Xbit_r137_c115 bl[115] br[115] wl[137] vdd gnd cell_6t
Xbit_r138_c115 bl[115] br[115] wl[138] vdd gnd cell_6t
Xbit_r139_c115 bl[115] br[115] wl[139] vdd gnd cell_6t
Xbit_r140_c115 bl[115] br[115] wl[140] vdd gnd cell_6t
Xbit_r141_c115 bl[115] br[115] wl[141] vdd gnd cell_6t
Xbit_r142_c115 bl[115] br[115] wl[142] vdd gnd cell_6t
Xbit_r143_c115 bl[115] br[115] wl[143] vdd gnd cell_6t
Xbit_r144_c115 bl[115] br[115] wl[144] vdd gnd cell_6t
Xbit_r145_c115 bl[115] br[115] wl[145] vdd gnd cell_6t
Xbit_r146_c115 bl[115] br[115] wl[146] vdd gnd cell_6t
Xbit_r147_c115 bl[115] br[115] wl[147] vdd gnd cell_6t
Xbit_r148_c115 bl[115] br[115] wl[148] vdd gnd cell_6t
Xbit_r149_c115 bl[115] br[115] wl[149] vdd gnd cell_6t
Xbit_r150_c115 bl[115] br[115] wl[150] vdd gnd cell_6t
Xbit_r151_c115 bl[115] br[115] wl[151] vdd gnd cell_6t
Xbit_r152_c115 bl[115] br[115] wl[152] vdd gnd cell_6t
Xbit_r153_c115 bl[115] br[115] wl[153] vdd gnd cell_6t
Xbit_r154_c115 bl[115] br[115] wl[154] vdd gnd cell_6t
Xbit_r155_c115 bl[115] br[115] wl[155] vdd gnd cell_6t
Xbit_r156_c115 bl[115] br[115] wl[156] vdd gnd cell_6t
Xbit_r157_c115 bl[115] br[115] wl[157] vdd gnd cell_6t
Xbit_r158_c115 bl[115] br[115] wl[158] vdd gnd cell_6t
Xbit_r159_c115 bl[115] br[115] wl[159] vdd gnd cell_6t
Xbit_r160_c115 bl[115] br[115] wl[160] vdd gnd cell_6t
Xbit_r161_c115 bl[115] br[115] wl[161] vdd gnd cell_6t
Xbit_r162_c115 bl[115] br[115] wl[162] vdd gnd cell_6t
Xbit_r163_c115 bl[115] br[115] wl[163] vdd gnd cell_6t
Xbit_r164_c115 bl[115] br[115] wl[164] vdd gnd cell_6t
Xbit_r165_c115 bl[115] br[115] wl[165] vdd gnd cell_6t
Xbit_r166_c115 bl[115] br[115] wl[166] vdd gnd cell_6t
Xbit_r167_c115 bl[115] br[115] wl[167] vdd gnd cell_6t
Xbit_r168_c115 bl[115] br[115] wl[168] vdd gnd cell_6t
Xbit_r169_c115 bl[115] br[115] wl[169] vdd gnd cell_6t
Xbit_r170_c115 bl[115] br[115] wl[170] vdd gnd cell_6t
Xbit_r171_c115 bl[115] br[115] wl[171] vdd gnd cell_6t
Xbit_r172_c115 bl[115] br[115] wl[172] vdd gnd cell_6t
Xbit_r173_c115 bl[115] br[115] wl[173] vdd gnd cell_6t
Xbit_r174_c115 bl[115] br[115] wl[174] vdd gnd cell_6t
Xbit_r175_c115 bl[115] br[115] wl[175] vdd gnd cell_6t
Xbit_r176_c115 bl[115] br[115] wl[176] vdd gnd cell_6t
Xbit_r177_c115 bl[115] br[115] wl[177] vdd gnd cell_6t
Xbit_r178_c115 bl[115] br[115] wl[178] vdd gnd cell_6t
Xbit_r179_c115 bl[115] br[115] wl[179] vdd gnd cell_6t
Xbit_r180_c115 bl[115] br[115] wl[180] vdd gnd cell_6t
Xbit_r181_c115 bl[115] br[115] wl[181] vdd gnd cell_6t
Xbit_r182_c115 bl[115] br[115] wl[182] vdd gnd cell_6t
Xbit_r183_c115 bl[115] br[115] wl[183] vdd gnd cell_6t
Xbit_r184_c115 bl[115] br[115] wl[184] vdd gnd cell_6t
Xbit_r185_c115 bl[115] br[115] wl[185] vdd gnd cell_6t
Xbit_r186_c115 bl[115] br[115] wl[186] vdd gnd cell_6t
Xbit_r187_c115 bl[115] br[115] wl[187] vdd gnd cell_6t
Xbit_r188_c115 bl[115] br[115] wl[188] vdd gnd cell_6t
Xbit_r189_c115 bl[115] br[115] wl[189] vdd gnd cell_6t
Xbit_r190_c115 bl[115] br[115] wl[190] vdd gnd cell_6t
Xbit_r191_c115 bl[115] br[115] wl[191] vdd gnd cell_6t
Xbit_r192_c115 bl[115] br[115] wl[192] vdd gnd cell_6t
Xbit_r193_c115 bl[115] br[115] wl[193] vdd gnd cell_6t
Xbit_r194_c115 bl[115] br[115] wl[194] vdd gnd cell_6t
Xbit_r195_c115 bl[115] br[115] wl[195] vdd gnd cell_6t
Xbit_r196_c115 bl[115] br[115] wl[196] vdd gnd cell_6t
Xbit_r197_c115 bl[115] br[115] wl[197] vdd gnd cell_6t
Xbit_r198_c115 bl[115] br[115] wl[198] vdd gnd cell_6t
Xbit_r199_c115 bl[115] br[115] wl[199] vdd gnd cell_6t
Xbit_r200_c115 bl[115] br[115] wl[200] vdd gnd cell_6t
Xbit_r201_c115 bl[115] br[115] wl[201] vdd gnd cell_6t
Xbit_r202_c115 bl[115] br[115] wl[202] vdd gnd cell_6t
Xbit_r203_c115 bl[115] br[115] wl[203] vdd gnd cell_6t
Xbit_r204_c115 bl[115] br[115] wl[204] vdd gnd cell_6t
Xbit_r205_c115 bl[115] br[115] wl[205] vdd gnd cell_6t
Xbit_r206_c115 bl[115] br[115] wl[206] vdd gnd cell_6t
Xbit_r207_c115 bl[115] br[115] wl[207] vdd gnd cell_6t
Xbit_r208_c115 bl[115] br[115] wl[208] vdd gnd cell_6t
Xbit_r209_c115 bl[115] br[115] wl[209] vdd gnd cell_6t
Xbit_r210_c115 bl[115] br[115] wl[210] vdd gnd cell_6t
Xbit_r211_c115 bl[115] br[115] wl[211] vdd gnd cell_6t
Xbit_r212_c115 bl[115] br[115] wl[212] vdd gnd cell_6t
Xbit_r213_c115 bl[115] br[115] wl[213] vdd gnd cell_6t
Xbit_r214_c115 bl[115] br[115] wl[214] vdd gnd cell_6t
Xbit_r215_c115 bl[115] br[115] wl[215] vdd gnd cell_6t
Xbit_r216_c115 bl[115] br[115] wl[216] vdd gnd cell_6t
Xbit_r217_c115 bl[115] br[115] wl[217] vdd gnd cell_6t
Xbit_r218_c115 bl[115] br[115] wl[218] vdd gnd cell_6t
Xbit_r219_c115 bl[115] br[115] wl[219] vdd gnd cell_6t
Xbit_r220_c115 bl[115] br[115] wl[220] vdd gnd cell_6t
Xbit_r221_c115 bl[115] br[115] wl[221] vdd gnd cell_6t
Xbit_r222_c115 bl[115] br[115] wl[222] vdd gnd cell_6t
Xbit_r223_c115 bl[115] br[115] wl[223] vdd gnd cell_6t
Xbit_r224_c115 bl[115] br[115] wl[224] vdd gnd cell_6t
Xbit_r225_c115 bl[115] br[115] wl[225] vdd gnd cell_6t
Xbit_r226_c115 bl[115] br[115] wl[226] vdd gnd cell_6t
Xbit_r227_c115 bl[115] br[115] wl[227] vdd gnd cell_6t
Xbit_r228_c115 bl[115] br[115] wl[228] vdd gnd cell_6t
Xbit_r229_c115 bl[115] br[115] wl[229] vdd gnd cell_6t
Xbit_r230_c115 bl[115] br[115] wl[230] vdd gnd cell_6t
Xbit_r231_c115 bl[115] br[115] wl[231] vdd gnd cell_6t
Xbit_r232_c115 bl[115] br[115] wl[232] vdd gnd cell_6t
Xbit_r233_c115 bl[115] br[115] wl[233] vdd gnd cell_6t
Xbit_r234_c115 bl[115] br[115] wl[234] vdd gnd cell_6t
Xbit_r235_c115 bl[115] br[115] wl[235] vdd gnd cell_6t
Xbit_r236_c115 bl[115] br[115] wl[236] vdd gnd cell_6t
Xbit_r237_c115 bl[115] br[115] wl[237] vdd gnd cell_6t
Xbit_r238_c115 bl[115] br[115] wl[238] vdd gnd cell_6t
Xbit_r239_c115 bl[115] br[115] wl[239] vdd gnd cell_6t
Xbit_r240_c115 bl[115] br[115] wl[240] vdd gnd cell_6t
Xbit_r241_c115 bl[115] br[115] wl[241] vdd gnd cell_6t
Xbit_r242_c115 bl[115] br[115] wl[242] vdd gnd cell_6t
Xbit_r243_c115 bl[115] br[115] wl[243] vdd gnd cell_6t
Xbit_r244_c115 bl[115] br[115] wl[244] vdd gnd cell_6t
Xbit_r245_c115 bl[115] br[115] wl[245] vdd gnd cell_6t
Xbit_r246_c115 bl[115] br[115] wl[246] vdd gnd cell_6t
Xbit_r247_c115 bl[115] br[115] wl[247] vdd gnd cell_6t
Xbit_r248_c115 bl[115] br[115] wl[248] vdd gnd cell_6t
Xbit_r249_c115 bl[115] br[115] wl[249] vdd gnd cell_6t
Xbit_r250_c115 bl[115] br[115] wl[250] vdd gnd cell_6t
Xbit_r251_c115 bl[115] br[115] wl[251] vdd gnd cell_6t
Xbit_r252_c115 bl[115] br[115] wl[252] vdd gnd cell_6t
Xbit_r253_c115 bl[115] br[115] wl[253] vdd gnd cell_6t
Xbit_r254_c115 bl[115] br[115] wl[254] vdd gnd cell_6t
Xbit_r255_c115 bl[115] br[115] wl[255] vdd gnd cell_6t
Xbit_r256_c115 bl[115] br[115] wl[256] vdd gnd cell_6t
Xbit_r257_c115 bl[115] br[115] wl[257] vdd gnd cell_6t
Xbit_r258_c115 bl[115] br[115] wl[258] vdd gnd cell_6t
Xbit_r259_c115 bl[115] br[115] wl[259] vdd gnd cell_6t
Xbit_r260_c115 bl[115] br[115] wl[260] vdd gnd cell_6t
Xbit_r261_c115 bl[115] br[115] wl[261] vdd gnd cell_6t
Xbit_r262_c115 bl[115] br[115] wl[262] vdd gnd cell_6t
Xbit_r263_c115 bl[115] br[115] wl[263] vdd gnd cell_6t
Xbit_r264_c115 bl[115] br[115] wl[264] vdd gnd cell_6t
Xbit_r265_c115 bl[115] br[115] wl[265] vdd gnd cell_6t
Xbit_r266_c115 bl[115] br[115] wl[266] vdd gnd cell_6t
Xbit_r267_c115 bl[115] br[115] wl[267] vdd gnd cell_6t
Xbit_r268_c115 bl[115] br[115] wl[268] vdd gnd cell_6t
Xbit_r269_c115 bl[115] br[115] wl[269] vdd gnd cell_6t
Xbit_r270_c115 bl[115] br[115] wl[270] vdd gnd cell_6t
Xbit_r271_c115 bl[115] br[115] wl[271] vdd gnd cell_6t
Xbit_r272_c115 bl[115] br[115] wl[272] vdd gnd cell_6t
Xbit_r273_c115 bl[115] br[115] wl[273] vdd gnd cell_6t
Xbit_r274_c115 bl[115] br[115] wl[274] vdd gnd cell_6t
Xbit_r275_c115 bl[115] br[115] wl[275] vdd gnd cell_6t
Xbit_r276_c115 bl[115] br[115] wl[276] vdd gnd cell_6t
Xbit_r277_c115 bl[115] br[115] wl[277] vdd gnd cell_6t
Xbit_r278_c115 bl[115] br[115] wl[278] vdd gnd cell_6t
Xbit_r279_c115 bl[115] br[115] wl[279] vdd gnd cell_6t
Xbit_r280_c115 bl[115] br[115] wl[280] vdd gnd cell_6t
Xbit_r281_c115 bl[115] br[115] wl[281] vdd gnd cell_6t
Xbit_r282_c115 bl[115] br[115] wl[282] vdd gnd cell_6t
Xbit_r283_c115 bl[115] br[115] wl[283] vdd gnd cell_6t
Xbit_r284_c115 bl[115] br[115] wl[284] vdd gnd cell_6t
Xbit_r285_c115 bl[115] br[115] wl[285] vdd gnd cell_6t
Xbit_r286_c115 bl[115] br[115] wl[286] vdd gnd cell_6t
Xbit_r287_c115 bl[115] br[115] wl[287] vdd gnd cell_6t
Xbit_r288_c115 bl[115] br[115] wl[288] vdd gnd cell_6t
Xbit_r289_c115 bl[115] br[115] wl[289] vdd gnd cell_6t
Xbit_r290_c115 bl[115] br[115] wl[290] vdd gnd cell_6t
Xbit_r291_c115 bl[115] br[115] wl[291] vdd gnd cell_6t
Xbit_r292_c115 bl[115] br[115] wl[292] vdd gnd cell_6t
Xbit_r293_c115 bl[115] br[115] wl[293] vdd gnd cell_6t
Xbit_r294_c115 bl[115] br[115] wl[294] vdd gnd cell_6t
Xbit_r295_c115 bl[115] br[115] wl[295] vdd gnd cell_6t
Xbit_r296_c115 bl[115] br[115] wl[296] vdd gnd cell_6t
Xbit_r297_c115 bl[115] br[115] wl[297] vdd gnd cell_6t
Xbit_r298_c115 bl[115] br[115] wl[298] vdd gnd cell_6t
Xbit_r299_c115 bl[115] br[115] wl[299] vdd gnd cell_6t
Xbit_r300_c115 bl[115] br[115] wl[300] vdd gnd cell_6t
Xbit_r301_c115 bl[115] br[115] wl[301] vdd gnd cell_6t
Xbit_r302_c115 bl[115] br[115] wl[302] vdd gnd cell_6t
Xbit_r303_c115 bl[115] br[115] wl[303] vdd gnd cell_6t
Xbit_r304_c115 bl[115] br[115] wl[304] vdd gnd cell_6t
Xbit_r305_c115 bl[115] br[115] wl[305] vdd gnd cell_6t
Xbit_r306_c115 bl[115] br[115] wl[306] vdd gnd cell_6t
Xbit_r307_c115 bl[115] br[115] wl[307] vdd gnd cell_6t
Xbit_r308_c115 bl[115] br[115] wl[308] vdd gnd cell_6t
Xbit_r309_c115 bl[115] br[115] wl[309] vdd gnd cell_6t
Xbit_r310_c115 bl[115] br[115] wl[310] vdd gnd cell_6t
Xbit_r311_c115 bl[115] br[115] wl[311] vdd gnd cell_6t
Xbit_r312_c115 bl[115] br[115] wl[312] vdd gnd cell_6t
Xbit_r313_c115 bl[115] br[115] wl[313] vdd gnd cell_6t
Xbit_r314_c115 bl[115] br[115] wl[314] vdd gnd cell_6t
Xbit_r315_c115 bl[115] br[115] wl[315] vdd gnd cell_6t
Xbit_r316_c115 bl[115] br[115] wl[316] vdd gnd cell_6t
Xbit_r317_c115 bl[115] br[115] wl[317] vdd gnd cell_6t
Xbit_r318_c115 bl[115] br[115] wl[318] vdd gnd cell_6t
Xbit_r319_c115 bl[115] br[115] wl[319] vdd gnd cell_6t
Xbit_r320_c115 bl[115] br[115] wl[320] vdd gnd cell_6t
Xbit_r321_c115 bl[115] br[115] wl[321] vdd gnd cell_6t
Xbit_r322_c115 bl[115] br[115] wl[322] vdd gnd cell_6t
Xbit_r323_c115 bl[115] br[115] wl[323] vdd gnd cell_6t
Xbit_r324_c115 bl[115] br[115] wl[324] vdd gnd cell_6t
Xbit_r325_c115 bl[115] br[115] wl[325] vdd gnd cell_6t
Xbit_r326_c115 bl[115] br[115] wl[326] vdd gnd cell_6t
Xbit_r327_c115 bl[115] br[115] wl[327] vdd gnd cell_6t
Xbit_r328_c115 bl[115] br[115] wl[328] vdd gnd cell_6t
Xbit_r329_c115 bl[115] br[115] wl[329] vdd gnd cell_6t
Xbit_r330_c115 bl[115] br[115] wl[330] vdd gnd cell_6t
Xbit_r331_c115 bl[115] br[115] wl[331] vdd gnd cell_6t
Xbit_r332_c115 bl[115] br[115] wl[332] vdd gnd cell_6t
Xbit_r333_c115 bl[115] br[115] wl[333] vdd gnd cell_6t
Xbit_r334_c115 bl[115] br[115] wl[334] vdd gnd cell_6t
Xbit_r335_c115 bl[115] br[115] wl[335] vdd gnd cell_6t
Xbit_r336_c115 bl[115] br[115] wl[336] vdd gnd cell_6t
Xbit_r337_c115 bl[115] br[115] wl[337] vdd gnd cell_6t
Xbit_r338_c115 bl[115] br[115] wl[338] vdd gnd cell_6t
Xbit_r339_c115 bl[115] br[115] wl[339] vdd gnd cell_6t
Xbit_r340_c115 bl[115] br[115] wl[340] vdd gnd cell_6t
Xbit_r341_c115 bl[115] br[115] wl[341] vdd gnd cell_6t
Xbit_r342_c115 bl[115] br[115] wl[342] vdd gnd cell_6t
Xbit_r343_c115 bl[115] br[115] wl[343] vdd gnd cell_6t
Xbit_r344_c115 bl[115] br[115] wl[344] vdd gnd cell_6t
Xbit_r345_c115 bl[115] br[115] wl[345] vdd gnd cell_6t
Xbit_r346_c115 bl[115] br[115] wl[346] vdd gnd cell_6t
Xbit_r347_c115 bl[115] br[115] wl[347] vdd gnd cell_6t
Xbit_r348_c115 bl[115] br[115] wl[348] vdd gnd cell_6t
Xbit_r349_c115 bl[115] br[115] wl[349] vdd gnd cell_6t
Xbit_r350_c115 bl[115] br[115] wl[350] vdd gnd cell_6t
Xbit_r351_c115 bl[115] br[115] wl[351] vdd gnd cell_6t
Xbit_r352_c115 bl[115] br[115] wl[352] vdd gnd cell_6t
Xbit_r353_c115 bl[115] br[115] wl[353] vdd gnd cell_6t
Xbit_r354_c115 bl[115] br[115] wl[354] vdd gnd cell_6t
Xbit_r355_c115 bl[115] br[115] wl[355] vdd gnd cell_6t
Xbit_r356_c115 bl[115] br[115] wl[356] vdd gnd cell_6t
Xbit_r357_c115 bl[115] br[115] wl[357] vdd gnd cell_6t
Xbit_r358_c115 bl[115] br[115] wl[358] vdd gnd cell_6t
Xbit_r359_c115 bl[115] br[115] wl[359] vdd gnd cell_6t
Xbit_r360_c115 bl[115] br[115] wl[360] vdd gnd cell_6t
Xbit_r361_c115 bl[115] br[115] wl[361] vdd gnd cell_6t
Xbit_r362_c115 bl[115] br[115] wl[362] vdd gnd cell_6t
Xbit_r363_c115 bl[115] br[115] wl[363] vdd gnd cell_6t
Xbit_r364_c115 bl[115] br[115] wl[364] vdd gnd cell_6t
Xbit_r365_c115 bl[115] br[115] wl[365] vdd gnd cell_6t
Xbit_r366_c115 bl[115] br[115] wl[366] vdd gnd cell_6t
Xbit_r367_c115 bl[115] br[115] wl[367] vdd gnd cell_6t
Xbit_r368_c115 bl[115] br[115] wl[368] vdd gnd cell_6t
Xbit_r369_c115 bl[115] br[115] wl[369] vdd gnd cell_6t
Xbit_r370_c115 bl[115] br[115] wl[370] vdd gnd cell_6t
Xbit_r371_c115 bl[115] br[115] wl[371] vdd gnd cell_6t
Xbit_r372_c115 bl[115] br[115] wl[372] vdd gnd cell_6t
Xbit_r373_c115 bl[115] br[115] wl[373] vdd gnd cell_6t
Xbit_r374_c115 bl[115] br[115] wl[374] vdd gnd cell_6t
Xbit_r375_c115 bl[115] br[115] wl[375] vdd gnd cell_6t
Xbit_r376_c115 bl[115] br[115] wl[376] vdd gnd cell_6t
Xbit_r377_c115 bl[115] br[115] wl[377] vdd gnd cell_6t
Xbit_r378_c115 bl[115] br[115] wl[378] vdd gnd cell_6t
Xbit_r379_c115 bl[115] br[115] wl[379] vdd gnd cell_6t
Xbit_r380_c115 bl[115] br[115] wl[380] vdd gnd cell_6t
Xbit_r381_c115 bl[115] br[115] wl[381] vdd gnd cell_6t
Xbit_r382_c115 bl[115] br[115] wl[382] vdd gnd cell_6t
Xbit_r383_c115 bl[115] br[115] wl[383] vdd gnd cell_6t
Xbit_r384_c115 bl[115] br[115] wl[384] vdd gnd cell_6t
Xbit_r385_c115 bl[115] br[115] wl[385] vdd gnd cell_6t
Xbit_r386_c115 bl[115] br[115] wl[386] vdd gnd cell_6t
Xbit_r387_c115 bl[115] br[115] wl[387] vdd gnd cell_6t
Xbit_r388_c115 bl[115] br[115] wl[388] vdd gnd cell_6t
Xbit_r389_c115 bl[115] br[115] wl[389] vdd gnd cell_6t
Xbit_r390_c115 bl[115] br[115] wl[390] vdd gnd cell_6t
Xbit_r391_c115 bl[115] br[115] wl[391] vdd gnd cell_6t
Xbit_r392_c115 bl[115] br[115] wl[392] vdd gnd cell_6t
Xbit_r393_c115 bl[115] br[115] wl[393] vdd gnd cell_6t
Xbit_r394_c115 bl[115] br[115] wl[394] vdd gnd cell_6t
Xbit_r395_c115 bl[115] br[115] wl[395] vdd gnd cell_6t
Xbit_r396_c115 bl[115] br[115] wl[396] vdd gnd cell_6t
Xbit_r397_c115 bl[115] br[115] wl[397] vdd gnd cell_6t
Xbit_r398_c115 bl[115] br[115] wl[398] vdd gnd cell_6t
Xbit_r399_c115 bl[115] br[115] wl[399] vdd gnd cell_6t
Xbit_r400_c115 bl[115] br[115] wl[400] vdd gnd cell_6t
Xbit_r401_c115 bl[115] br[115] wl[401] vdd gnd cell_6t
Xbit_r402_c115 bl[115] br[115] wl[402] vdd gnd cell_6t
Xbit_r403_c115 bl[115] br[115] wl[403] vdd gnd cell_6t
Xbit_r404_c115 bl[115] br[115] wl[404] vdd gnd cell_6t
Xbit_r405_c115 bl[115] br[115] wl[405] vdd gnd cell_6t
Xbit_r406_c115 bl[115] br[115] wl[406] vdd gnd cell_6t
Xbit_r407_c115 bl[115] br[115] wl[407] vdd gnd cell_6t
Xbit_r408_c115 bl[115] br[115] wl[408] vdd gnd cell_6t
Xbit_r409_c115 bl[115] br[115] wl[409] vdd gnd cell_6t
Xbit_r410_c115 bl[115] br[115] wl[410] vdd gnd cell_6t
Xbit_r411_c115 bl[115] br[115] wl[411] vdd gnd cell_6t
Xbit_r412_c115 bl[115] br[115] wl[412] vdd gnd cell_6t
Xbit_r413_c115 bl[115] br[115] wl[413] vdd gnd cell_6t
Xbit_r414_c115 bl[115] br[115] wl[414] vdd gnd cell_6t
Xbit_r415_c115 bl[115] br[115] wl[415] vdd gnd cell_6t
Xbit_r416_c115 bl[115] br[115] wl[416] vdd gnd cell_6t
Xbit_r417_c115 bl[115] br[115] wl[417] vdd gnd cell_6t
Xbit_r418_c115 bl[115] br[115] wl[418] vdd gnd cell_6t
Xbit_r419_c115 bl[115] br[115] wl[419] vdd gnd cell_6t
Xbit_r420_c115 bl[115] br[115] wl[420] vdd gnd cell_6t
Xbit_r421_c115 bl[115] br[115] wl[421] vdd gnd cell_6t
Xbit_r422_c115 bl[115] br[115] wl[422] vdd gnd cell_6t
Xbit_r423_c115 bl[115] br[115] wl[423] vdd gnd cell_6t
Xbit_r424_c115 bl[115] br[115] wl[424] vdd gnd cell_6t
Xbit_r425_c115 bl[115] br[115] wl[425] vdd gnd cell_6t
Xbit_r426_c115 bl[115] br[115] wl[426] vdd gnd cell_6t
Xbit_r427_c115 bl[115] br[115] wl[427] vdd gnd cell_6t
Xbit_r428_c115 bl[115] br[115] wl[428] vdd gnd cell_6t
Xbit_r429_c115 bl[115] br[115] wl[429] vdd gnd cell_6t
Xbit_r430_c115 bl[115] br[115] wl[430] vdd gnd cell_6t
Xbit_r431_c115 bl[115] br[115] wl[431] vdd gnd cell_6t
Xbit_r432_c115 bl[115] br[115] wl[432] vdd gnd cell_6t
Xbit_r433_c115 bl[115] br[115] wl[433] vdd gnd cell_6t
Xbit_r434_c115 bl[115] br[115] wl[434] vdd gnd cell_6t
Xbit_r435_c115 bl[115] br[115] wl[435] vdd gnd cell_6t
Xbit_r436_c115 bl[115] br[115] wl[436] vdd gnd cell_6t
Xbit_r437_c115 bl[115] br[115] wl[437] vdd gnd cell_6t
Xbit_r438_c115 bl[115] br[115] wl[438] vdd gnd cell_6t
Xbit_r439_c115 bl[115] br[115] wl[439] vdd gnd cell_6t
Xbit_r440_c115 bl[115] br[115] wl[440] vdd gnd cell_6t
Xbit_r441_c115 bl[115] br[115] wl[441] vdd gnd cell_6t
Xbit_r442_c115 bl[115] br[115] wl[442] vdd gnd cell_6t
Xbit_r443_c115 bl[115] br[115] wl[443] vdd gnd cell_6t
Xbit_r444_c115 bl[115] br[115] wl[444] vdd gnd cell_6t
Xbit_r445_c115 bl[115] br[115] wl[445] vdd gnd cell_6t
Xbit_r446_c115 bl[115] br[115] wl[446] vdd gnd cell_6t
Xbit_r447_c115 bl[115] br[115] wl[447] vdd gnd cell_6t
Xbit_r448_c115 bl[115] br[115] wl[448] vdd gnd cell_6t
Xbit_r449_c115 bl[115] br[115] wl[449] vdd gnd cell_6t
Xbit_r450_c115 bl[115] br[115] wl[450] vdd gnd cell_6t
Xbit_r451_c115 bl[115] br[115] wl[451] vdd gnd cell_6t
Xbit_r452_c115 bl[115] br[115] wl[452] vdd gnd cell_6t
Xbit_r453_c115 bl[115] br[115] wl[453] vdd gnd cell_6t
Xbit_r454_c115 bl[115] br[115] wl[454] vdd gnd cell_6t
Xbit_r455_c115 bl[115] br[115] wl[455] vdd gnd cell_6t
Xbit_r456_c115 bl[115] br[115] wl[456] vdd gnd cell_6t
Xbit_r457_c115 bl[115] br[115] wl[457] vdd gnd cell_6t
Xbit_r458_c115 bl[115] br[115] wl[458] vdd gnd cell_6t
Xbit_r459_c115 bl[115] br[115] wl[459] vdd gnd cell_6t
Xbit_r460_c115 bl[115] br[115] wl[460] vdd gnd cell_6t
Xbit_r461_c115 bl[115] br[115] wl[461] vdd gnd cell_6t
Xbit_r462_c115 bl[115] br[115] wl[462] vdd gnd cell_6t
Xbit_r463_c115 bl[115] br[115] wl[463] vdd gnd cell_6t
Xbit_r464_c115 bl[115] br[115] wl[464] vdd gnd cell_6t
Xbit_r465_c115 bl[115] br[115] wl[465] vdd gnd cell_6t
Xbit_r466_c115 bl[115] br[115] wl[466] vdd gnd cell_6t
Xbit_r467_c115 bl[115] br[115] wl[467] vdd gnd cell_6t
Xbit_r468_c115 bl[115] br[115] wl[468] vdd gnd cell_6t
Xbit_r469_c115 bl[115] br[115] wl[469] vdd gnd cell_6t
Xbit_r470_c115 bl[115] br[115] wl[470] vdd gnd cell_6t
Xbit_r471_c115 bl[115] br[115] wl[471] vdd gnd cell_6t
Xbit_r472_c115 bl[115] br[115] wl[472] vdd gnd cell_6t
Xbit_r473_c115 bl[115] br[115] wl[473] vdd gnd cell_6t
Xbit_r474_c115 bl[115] br[115] wl[474] vdd gnd cell_6t
Xbit_r475_c115 bl[115] br[115] wl[475] vdd gnd cell_6t
Xbit_r476_c115 bl[115] br[115] wl[476] vdd gnd cell_6t
Xbit_r477_c115 bl[115] br[115] wl[477] vdd gnd cell_6t
Xbit_r478_c115 bl[115] br[115] wl[478] vdd gnd cell_6t
Xbit_r479_c115 bl[115] br[115] wl[479] vdd gnd cell_6t
Xbit_r480_c115 bl[115] br[115] wl[480] vdd gnd cell_6t
Xbit_r481_c115 bl[115] br[115] wl[481] vdd gnd cell_6t
Xbit_r482_c115 bl[115] br[115] wl[482] vdd gnd cell_6t
Xbit_r483_c115 bl[115] br[115] wl[483] vdd gnd cell_6t
Xbit_r484_c115 bl[115] br[115] wl[484] vdd gnd cell_6t
Xbit_r485_c115 bl[115] br[115] wl[485] vdd gnd cell_6t
Xbit_r486_c115 bl[115] br[115] wl[486] vdd gnd cell_6t
Xbit_r487_c115 bl[115] br[115] wl[487] vdd gnd cell_6t
Xbit_r488_c115 bl[115] br[115] wl[488] vdd gnd cell_6t
Xbit_r489_c115 bl[115] br[115] wl[489] vdd gnd cell_6t
Xbit_r490_c115 bl[115] br[115] wl[490] vdd gnd cell_6t
Xbit_r491_c115 bl[115] br[115] wl[491] vdd gnd cell_6t
Xbit_r492_c115 bl[115] br[115] wl[492] vdd gnd cell_6t
Xbit_r493_c115 bl[115] br[115] wl[493] vdd gnd cell_6t
Xbit_r494_c115 bl[115] br[115] wl[494] vdd gnd cell_6t
Xbit_r495_c115 bl[115] br[115] wl[495] vdd gnd cell_6t
Xbit_r496_c115 bl[115] br[115] wl[496] vdd gnd cell_6t
Xbit_r497_c115 bl[115] br[115] wl[497] vdd gnd cell_6t
Xbit_r498_c115 bl[115] br[115] wl[498] vdd gnd cell_6t
Xbit_r499_c115 bl[115] br[115] wl[499] vdd gnd cell_6t
Xbit_r500_c115 bl[115] br[115] wl[500] vdd gnd cell_6t
Xbit_r501_c115 bl[115] br[115] wl[501] vdd gnd cell_6t
Xbit_r502_c115 bl[115] br[115] wl[502] vdd gnd cell_6t
Xbit_r503_c115 bl[115] br[115] wl[503] vdd gnd cell_6t
Xbit_r504_c115 bl[115] br[115] wl[504] vdd gnd cell_6t
Xbit_r505_c115 bl[115] br[115] wl[505] vdd gnd cell_6t
Xbit_r506_c115 bl[115] br[115] wl[506] vdd gnd cell_6t
Xbit_r507_c115 bl[115] br[115] wl[507] vdd gnd cell_6t
Xbit_r508_c115 bl[115] br[115] wl[508] vdd gnd cell_6t
Xbit_r509_c115 bl[115] br[115] wl[509] vdd gnd cell_6t
Xbit_r510_c115 bl[115] br[115] wl[510] vdd gnd cell_6t
Xbit_r511_c115 bl[115] br[115] wl[511] vdd gnd cell_6t
Xbit_r0_c116 bl[116] br[116] wl[0] vdd gnd cell_6t
Xbit_r1_c116 bl[116] br[116] wl[1] vdd gnd cell_6t
Xbit_r2_c116 bl[116] br[116] wl[2] vdd gnd cell_6t
Xbit_r3_c116 bl[116] br[116] wl[3] vdd gnd cell_6t
Xbit_r4_c116 bl[116] br[116] wl[4] vdd gnd cell_6t
Xbit_r5_c116 bl[116] br[116] wl[5] vdd gnd cell_6t
Xbit_r6_c116 bl[116] br[116] wl[6] vdd gnd cell_6t
Xbit_r7_c116 bl[116] br[116] wl[7] vdd gnd cell_6t
Xbit_r8_c116 bl[116] br[116] wl[8] vdd gnd cell_6t
Xbit_r9_c116 bl[116] br[116] wl[9] vdd gnd cell_6t
Xbit_r10_c116 bl[116] br[116] wl[10] vdd gnd cell_6t
Xbit_r11_c116 bl[116] br[116] wl[11] vdd gnd cell_6t
Xbit_r12_c116 bl[116] br[116] wl[12] vdd gnd cell_6t
Xbit_r13_c116 bl[116] br[116] wl[13] vdd gnd cell_6t
Xbit_r14_c116 bl[116] br[116] wl[14] vdd gnd cell_6t
Xbit_r15_c116 bl[116] br[116] wl[15] vdd gnd cell_6t
Xbit_r16_c116 bl[116] br[116] wl[16] vdd gnd cell_6t
Xbit_r17_c116 bl[116] br[116] wl[17] vdd gnd cell_6t
Xbit_r18_c116 bl[116] br[116] wl[18] vdd gnd cell_6t
Xbit_r19_c116 bl[116] br[116] wl[19] vdd gnd cell_6t
Xbit_r20_c116 bl[116] br[116] wl[20] vdd gnd cell_6t
Xbit_r21_c116 bl[116] br[116] wl[21] vdd gnd cell_6t
Xbit_r22_c116 bl[116] br[116] wl[22] vdd gnd cell_6t
Xbit_r23_c116 bl[116] br[116] wl[23] vdd gnd cell_6t
Xbit_r24_c116 bl[116] br[116] wl[24] vdd gnd cell_6t
Xbit_r25_c116 bl[116] br[116] wl[25] vdd gnd cell_6t
Xbit_r26_c116 bl[116] br[116] wl[26] vdd gnd cell_6t
Xbit_r27_c116 bl[116] br[116] wl[27] vdd gnd cell_6t
Xbit_r28_c116 bl[116] br[116] wl[28] vdd gnd cell_6t
Xbit_r29_c116 bl[116] br[116] wl[29] vdd gnd cell_6t
Xbit_r30_c116 bl[116] br[116] wl[30] vdd gnd cell_6t
Xbit_r31_c116 bl[116] br[116] wl[31] vdd gnd cell_6t
Xbit_r32_c116 bl[116] br[116] wl[32] vdd gnd cell_6t
Xbit_r33_c116 bl[116] br[116] wl[33] vdd gnd cell_6t
Xbit_r34_c116 bl[116] br[116] wl[34] vdd gnd cell_6t
Xbit_r35_c116 bl[116] br[116] wl[35] vdd gnd cell_6t
Xbit_r36_c116 bl[116] br[116] wl[36] vdd gnd cell_6t
Xbit_r37_c116 bl[116] br[116] wl[37] vdd gnd cell_6t
Xbit_r38_c116 bl[116] br[116] wl[38] vdd gnd cell_6t
Xbit_r39_c116 bl[116] br[116] wl[39] vdd gnd cell_6t
Xbit_r40_c116 bl[116] br[116] wl[40] vdd gnd cell_6t
Xbit_r41_c116 bl[116] br[116] wl[41] vdd gnd cell_6t
Xbit_r42_c116 bl[116] br[116] wl[42] vdd gnd cell_6t
Xbit_r43_c116 bl[116] br[116] wl[43] vdd gnd cell_6t
Xbit_r44_c116 bl[116] br[116] wl[44] vdd gnd cell_6t
Xbit_r45_c116 bl[116] br[116] wl[45] vdd gnd cell_6t
Xbit_r46_c116 bl[116] br[116] wl[46] vdd gnd cell_6t
Xbit_r47_c116 bl[116] br[116] wl[47] vdd gnd cell_6t
Xbit_r48_c116 bl[116] br[116] wl[48] vdd gnd cell_6t
Xbit_r49_c116 bl[116] br[116] wl[49] vdd gnd cell_6t
Xbit_r50_c116 bl[116] br[116] wl[50] vdd gnd cell_6t
Xbit_r51_c116 bl[116] br[116] wl[51] vdd gnd cell_6t
Xbit_r52_c116 bl[116] br[116] wl[52] vdd gnd cell_6t
Xbit_r53_c116 bl[116] br[116] wl[53] vdd gnd cell_6t
Xbit_r54_c116 bl[116] br[116] wl[54] vdd gnd cell_6t
Xbit_r55_c116 bl[116] br[116] wl[55] vdd gnd cell_6t
Xbit_r56_c116 bl[116] br[116] wl[56] vdd gnd cell_6t
Xbit_r57_c116 bl[116] br[116] wl[57] vdd gnd cell_6t
Xbit_r58_c116 bl[116] br[116] wl[58] vdd gnd cell_6t
Xbit_r59_c116 bl[116] br[116] wl[59] vdd gnd cell_6t
Xbit_r60_c116 bl[116] br[116] wl[60] vdd gnd cell_6t
Xbit_r61_c116 bl[116] br[116] wl[61] vdd gnd cell_6t
Xbit_r62_c116 bl[116] br[116] wl[62] vdd gnd cell_6t
Xbit_r63_c116 bl[116] br[116] wl[63] vdd gnd cell_6t
Xbit_r64_c116 bl[116] br[116] wl[64] vdd gnd cell_6t
Xbit_r65_c116 bl[116] br[116] wl[65] vdd gnd cell_6t
Xbit_r66_c116 bl[116] br[116] wl[66] vdd gnd cell_6t
Xbit_r67_c116 bl[116] br[116] wl[67] vdd gnd cell_6t
Xbit_r68_c116 bl[116] br[116] wl[68] vdd gnd cell_6t
Xbit_r69_c116 bl[116] br[116] wl[69] vdd gnd cell_6t
Xbit_r70_c116 bl[116] br[116] wl[70] vdd gnd cell_6t
Xbit_r71_c116 bl[116] br[116] wl[71] vdd gnd cell_6t
Xbit_r72_c116 bl[116] br[116] wl[72] vdd gnd cell_6t
Xbit_r73_c116 bl[116] br[116] wl[73] vdd gnd cell_6t
Xbit_r74_c116 bl[116] br[116] wl[74] vdd gnd cell_6t
Xbit_r75_c116 bl[116] br[116] wl[75] vdd gnd cell_6t
Xbit_r76_c116 bl[116] br[116] wl[76] vdd gnd cell_6t
Xbit_r77_c116 bl[116] br[116] wl[77] vdd gnd cell_6t
Xbit_r78_c116 bl[116] br[116] wl[78] vdd gnd cell_6t
Xbit_r79_c116 bl[116] br[116] wl[79] vdd gnd cell_6t
Xbit_r80_c116 bl[116] br[116] wl[80] vdd gnd cell_6t
Xbit_r81_c116 bl[116] br[116] wl[81] vdd gnd cell_6t
Xbit_r82_c116 bl[116] br[116] wl[82] vdd gnd cell_6t
Xbit_r83_c116 bl[116] br[116] wl[83] vdd gnd cell_6t
Xbit_r84_c116 bl[116] br[116] wl[84] vdd gnd cell_6t
Xbit_r85_c116 bl[116] br[116] wl[85] vdd gnd cell_6t
Xbit_r86_c116 bl[116] br[116] wl[86] vdd gnd cell_6t
Xbit_r87_c116 bl[116] br[116] wl[87] vdd gnd cell_6t
Xbit_r88_c116 bl[116] br[116] wl[88] vdd gnd cell_6t
Xbit_r89_c116 bl[116] br[116] wl[89] vdd gnd cell_6t
Xbit_r90_c116 bl[116] br[116] wl[90] vdd gnd cell_6t
Xbit_r91_c116 bl[116] br[116] wl[91] vdd gnd cell_6t
Xbit_r92_c116 bl[116] br[116] wl[92] vdd gnd cell_6t
Xbit_r93_c116 bl[116] br[116] wl[93] vdd gnd cell_6t
Xbit_r94_c116 bl[116] br[116] wl[94] vdd gnd cell_6t
Xbit_r95_c116 bl[116] br[116] wl[95] vdd gnd cell_6t
Xbit_r96_c116 bl[116] br[116] wl[96] vdd gnd cell_6t
Xbit_r97_c116 bl[116] br[116] wl[97] vdd gnd cell_6t
Xbit_r98_c116 bl[116] br[116] wl[98] vdd gnd cell_6t
Xbit_r99_c116 bl[116] br[116] wl[99] vdd gnd cell_6t
Xbit_r100_c116 bl[116] br[116] wl[100] vdd gnd cell_6t
Xbit_r101_c116 bl[116] br[116] wl[101] vdd gnd cell_6t
Xbit_r102_c116 bl[116] br[116] wl[102] vdd gnd cell_6t
Xbit_r103_c116 bl[116] br[116] wl[103] vdd gnd cell_6t
Xbit_r104_c116 bl[116] br[116] wl[104] vdd gnd cell_6t
Xbit_r105_c116 bl[116] br[116] wl[105] vdd gnd cell_6t
Xbit_r106_c116 bl[116] br[116] wl[106] vdd gnd cell_6t
Xbit_r107_c116 bl[116] br[116] wl[107] vdd gnd cell_6t
Xbit_r108_c116 bl[116] br[116] wl[108] vdd gnd cell_6t
Xbit_r109_c116 bl[116] br[116] wl[109] vdd gnd cell_6t
Xbit_r110_c116 bl[116] br[116] wl[110] vdd gnd cell_6t
Xbit_r111_c116 bl[116] br[116] wl[111] vdd gnd cell_6t
Xbit_r112_c116 bl[116] br[116] wl[112] vdd gnd cell_6t
Xbit_r113_c116 bl[116] br[116] wl[113] vdd gnd cell_6t
Xbit_r114_c116 bl[116] br[116] wl[114] vdd gnd cell_6t
Xbit_r115_c116 bl[116] br[116] wl[115] vdd gnd cell_6t
Xbit_r116_c116 bl[116] br[116] wl[116] vdd gnd cell_6t
Xbit_r117_c116 bl[116] br[116] wl[117] vdd gnd cell_6t
Xbit_r118_c116 bl[116] br[116] wl[118] vdd gnd cell_6t
Xbit_r119_c116 bl[116] br[116] wl[119] vdd gnd cell_6t
Xbit_r120_c116 bl[116] br[116] wl[120] vdd gnd cell_6t
Xbit_r121_c116 bl[116] br[116] wl[121] vdd gnd cell_6t
Xbit_r122_c116 bl[116] br[116] wl[122] vdd gnd cell_6t
Xbit_r123_c116 bl[116] br[116] wl[123] vdd gnd cell_6t
Xbit_r124_c116 bl[116] br[116] wl[124] vdd gnd cell_6t
Xbit_r125_c116 bl[116] br[116] wl[125] vdd gnd cell_6t
Xbit_r126_c116 bl[116] br[116] wl[126] vdd gnd cell_6t
Xbit_r127_c116 bl[116] br[116] wl[127] vdd gnd cell_6t
Xbit_r128_c116 bl[116] br[116] wl[128] vdd gnd cell_6t
Xbit_r129_c116 bl[116] br[116] wl[129] vdd gnd cell_6t
Xbit_r130_c116 bl[116] br[116] wl[130] vdd gnd cell_6t
Xbit_r131_c116 bl[116] br[116] wl[131] vdd gnd cell_6t
Xbit_r132_c116 bl[116] br[116] wl[132] vdd gnd cell_6t
Xbit_r133_c116 bl[116] br[116] wl[133] vdd gnd cell_6t
Xbit_r134_c116 bl[116] br[116] wl[134] vdd gnd cell_6t
Xbit_r135_c116 bl[116] br[116] wl[135] vdd gnd cell_6t
Xbit_r136_c116 bl[116] br[116] wl[136] vdd gnd cell_6t
Xbit_r137_c116 bl[116] br[116] wl[137] vdd gnd cell_6t
Xbit_r138_c116 bl[116] br[116] wl[138] vdd gnd cell_6t
Xbit_r139_c116 bl[116] br[116] wl[139] vdd gnd cell_6t
Xbit_r140_c116 bl[116] br[116] wl[140] vdd gnd cell_6t
Xbit_r141_c116 bl[116] br[116] wl[141] vdd gnd cell_6t
Xbit_r142_c116 bl[116] br[116] wl[142] vdd gnd cell_6t
Xbit_r143_c116 bl[116] br[116] wl[143] vdd gnd cell_6t
Xbit_r144_c116 bl[116] br[116] wl[144] vdd gnd cell_6t
Xbit_r145_c116 bl[116] br[116] wl[145] vdd gnd cell_6t
Xbit_r146_c116 bl[116] br[116] wl[146] vdd gnd cell_6t
Xbit_r147_c116 bl[116] br[116] wl[147] vdd gnd cell_6t
Xbit_r148_c116 bl[116] br[116] wl[148] vdd gnd cell_6t
Xbit_r149_c116 bl[116] br[116] wl[149] vdd gnd cell_6t
Xbit_r150_c116 bl[116] br[116] wl[150] vdd gnd cell_6t
Xbit_r151_c116 bl[116] br[116] wl[151] vdd gnd cell_6t
Xbit_r152_c116 bl[116] br[116] wl[152] vdd gnd cell_6t
Xbit_r153_c116 bl[116] br[116] wl[153] vdd gnd cell_6t
Xbit_r154_c116 bl[116] br[116] wl[154] vdd gnd cell_6t
Xbit_r155_c116 bl[116] br[116] wl[155] vdd gnd cell_6t
Xbit_r156_c116 bl[116] br[116] wl[156] vdd gnd cell_6t
Xbit_r157_c116 bl[116] br[116] wl[157] vdd gnd cell_6t
Xbit_r158_c116 bl[116] br[116] wl[158] vdd gnd cell_6t
Xbit_r159_c116 bl[116] br[116] wl[159] vdd gnd cell_6t
Xbit_r160_c116 bl[116] br[116] wl[160] vdd gnd cell_6t
Xbit_r161_c116 bl[116] br[116] wl[161] vdd gnd cell_6t
Xbit_r162_c116 bl[116] br[116] wl[162] vdd gnd cell_6t
Xbit_r163_c116 bl[116] br[116] wl[163] vdd gnd cell_6t
Xbit_r164_c116 bl[116] br[116] wl[164] vdd gnd cell_6t
Xbit_r165_c116 bl[116] br[116] wl[165] vdd gnd cell_6t
Xbit_r166_c116 bl[116] br[116] wl[166] vdd gnd cell_6t
Xbit_r167_c116 bl[116] br[116] wl[167] vdd gnd cell_6t
Xbit_r168_c116 bl[116] br[116] wl[168] vdd gnd cell_6t
Xbit_r169_c116 bl[116] br[116] wl[169] vdd gnd cell_6t
Xbit_r170_c116 bl[116] br[116] wl[170] vdd gnd cell_6t
Xbit_r171_c116 bl[116] br[116] wl[171] vdd gnd cell_6t
Xbit_r172_c116 bl[116] br[116] wl[172] vdd gnd cell_6t
Xbit_r173_c116 bl[116] br[116] wl[173] vdd gnd cell_6t
Xbit_r174_c116 bl[116] br[116] wl[174] vdd gnd cell_6t
Xbit_r175_c116 bl[116] br[116] wl[175] vdd gnd cell_6t
Xbit_r176_c116 bl[116] br[116] wl[176] vdd gnd cell_6t
Xbit_r177_c116 bl[116] br[116] wl[177] vdd gnd cell_6t
Xbit_r178_c116 bl[116] br[116] wl[178] vdd gnd cell_6t
Xbit_r179_c116 bl[116] br[116] wl[179] vdd gnd cell_6t
Xbit_r180_c116 bl[116] br[116] wl[180] vdd gnd cell_6t
Xbit_r181_c116 bl[116] br[116] wl[181] vdd gnd cell_6t
Xbit_r182_c116 bl[116] br[116] wl[182] vdd gnd cell_6t
Xbit_r183_c116 bl[116] br[116] wl[183] vdd gnd cell_6t
Xbit_r184_c116 bl[116] br[116] wl[184] vdd gnd cell_6t
Xbit_r185_c116 bl[116] br[116] wl[185] vdd gnd cell_6t
Xbit_r186_c116 bl[116] br[116] wl[186] vdd gnd cell_6t
Xbit_r187_c116 bl[116] br[116] wl[187] vdd gnd cell_6t
Xbit_r188_c116 bl[116] br[116] wl[188] vdd gnd cell_6t
Xbit_r189_c116 bl[116] br[116] wl[189] vdd gnd cell_6t
Xbit_r190_c116 bl[116] br[116] wl[190] vdd gnd cell_6t
Xbit_r191_c116 bl[116] br[116] wl[191] vdd gnd cell_6t
Xbit_r192_c116 bl[116] br[116] wl[192] vdd gnd cell_6t
Xbit_r193_c116 bl[116] br[116] wl[193] vdd gnd cell_6t
Xbit_r194_c116 bl[116] br[116] wl[194] vdd gnd cell_6t
Xbit_r195_c116 bl[116] br[116] wl[195] vdd gnd cell_6t
Xbit_r196_c116 bl[116] br[116] wl[196] vdd gnd cell_6t
Xbit_r197_c116 bl[116] br[116] wl[197] vdd gnd cell_6t
Xbit_r198_c116 bl[116] br[116] wl[198] vdd gnd cell_6t
Xbit_r199_c116 bl[116] br[116] wl[199] vdd gnd cell_6t
Xbit_r200_c116 bl[116] br[116] wl[200] vdd gnd cell_6t
Xbit_r201_c116 bl[116] br[116] wl[201] vdd gnd cell_6t
Xbit_r202_c116 bl[116] br[116] wl[202] vdd gnd cell_6t
Xbit_r203_c116 bl[116] br[116] wl[203] vdd gnd cell_6t
Xbit_r204_c116 bl[116] br[116] wl[204] vdd gnd cell_6t
Xbit_r205_c116 bl[116] br[116] wl[205] vdd gnd cell_6t
Xbit_r206_c116 bl[116] br[116] wl[206] vdd gnd cell_6t
Xbit_r207_c116 bl[116] br[116] wl[207] vdd gnd cell_6t
Xbit_r208_c116 bl[116] br[116] wl[208] vdd gnd cell_6t
Xbit_r209_c116 bl[116] br[116] wl[209] vdd gnd cell_6t
Xbit_r210_c116 bl[116] br[116] wl[210] vdd gnd cell_6t
Xbit_r211_c116 bl[116] br[116] wl[211] vdd gnd cell_6t
Xbit_r212_c116 bl[116] br[116] wl[212] vdd gnd cell_6t
Xbit_r213_c116 bl[116] br[116] wl[213] vdd gnd cell_6t
Xbit_r214_c116 bl[116] br[116] wl[214] vdd gnd cell_6t
Xbit_r215_c116 bl[116] br[116] wl[215] vdd gnd cell_6t
Xbit_r216_c116 bl[116] br[116] wl[216] vdd gnd cell_6t
Xbit_r217_c116 bl[116] br[116] wl[217] vdd gnd cell_6t
Xbit_r218_c116 bl[116] br[116] wl[218] vdd gnd cell_6t
Xbit_r219_c116 bl[116] br[116] wl[219] vdd gnd cell_6t
Xbit_r220_c116 bl[116] br[116] wl[220] vdd gnd cell_6t
Xbit_r221_c116 bl[116] br[116] wl[221] vdd gnd cell_6t
Xbit_r222_c116 bl[116] br[116] wl[222] vdd gnd cell_6t
Xbit_r223_c116 bl[116] br[116] wl[223] vdd gnd cell_6t
Xbit_r224_c116 bl[116] br[116] wl[224] vdd gnd cell_6t
Xbit_r225_c116 bl[116] br[116] wl[225] vdd gnd cell_6t
Xbit_r226_c116 bl[116] br[116] wl[226] vdd gnd cell_6t
Xbit_r227_c116 bl[116] br[116] wl[227] vdd gnd cell_6t
Xbit_r228_c116 bl[116] br[116] wl[228] vdd gnd cell_6t
Xbit_r229_c116 bl[116] br[116] wl[229] vdd gnd cell_6t
Xbit_r230_c116 bl[116] br[116] wl[230] vdd gnd cell_6t
Xbit_r231_c116 bl[116] br[116] wl[231] vdd gnd cell_6t
Xbit_r232_c116 bl[116] br[116] wl[232] vdd gnd cell_6t
Xbit_r233_c116 bl[116] br[116] wl[233] vdd gnd cell_6t
Xbit_r234_c116 bl[116] br[116] wl[234] vdd gnd cell_6t
Xbit_r235_c116 bl[116] br[116] wl[235] vdd gnd cell_6t
Xbit_r236_c116 bl[116] br[116] wl[236] vdd gnd cell_6t
Xbit_r237_c116 bl[116] br[116] wl[237] vdd gnd cell_6t
Xbit_r238_c116 bl[116] br[116] wl[238] vdd gnd cell_6t
Xbit_r239_c116 bl[116] br[116] wl[239] vdd gnd cell_6t
Xbit_r240_c116 bl[116] br[116] wl[240] vdd gnd cell_6t
Xbit_r241_c116 bl[116] br[116] wl[241] vdd gnd cell_6t
Xbit_r242_c116 bl[116] br[116] wl[242] vdd gnd cell_6t
Xbit_r243_c116 bl[116] br[116] wl[243] vdd gnd cell_6t
Xbit_r244_c116 bl[116] br[116] wl[244] vdd gnd cell_6t
Xbit_r245_c116 bl[116] br[116] wl[245] vdd gnd cell_6t
Xbit_r246_c116 bl[116] br[116] wl[246] vdd gnd cell_6t
Xbit_r247_c116 bl[116] br[116] wl[247] vdd gnd cell_6t
Xbit_r248_c116 bl[116] br[116] wl[248] vdd gnd cell_6t
Xbit_r249_c116 bl[116] br[116] wl[249] vdd gnd cell_6t
Xbit_r250_c116 bl[116] br[116] wl[250] vdd gnd cell_6t
Xbit_r251_c116 bl[116] br[116] wl[251] vdd gnd cell_6t
Xbit_r252_c116 bl[116] br[116] wl[252] vdd gnd cell_6t
Xbit_r253_c116 bl[116] br[116] wl[253] vdd gnd cell_6t
Xbit_r254_c116 bl[116] br[116] wl[254] vdd gnd cell_6t
Xbit_r255_c116 bl[116] br[116] wl[255] vdd gnd cell_6t
Xbit_r256_c116 bl[116] br[116] wl[256] vdd gnd cell_6t
Xbit_r257_c116 bl[116] br[116] wl[257] vdd gnd cell_6t
Xbit_r258_c116 bl[116] br[116] wl[258] vdd gnd cell_6t
Xbit_r259_c116 bl[116] br[116] wl[259] vdd gnd cell_6t
Xbit_r260_c116 bl[116] br[116] wl[260] vdd gnd cell_6t
Xbit_r261_c116 bl[116] br[116] wl[261] vdd gnd cell_6t
Xbit_r262_c116 bl[116] br[116] wl[262] vdd gnd cell_6t
Xbit_r263_c116 bl[116] br[116] wl[263] vdd gnd cell_6t
Xbit_r264_c116 bl[116] br[116] wl[264] vdd gnd cell_6t
Xbit_r265_c116 bl[116] br[116] wl[265] vdd gnd cell_6t
Xbit_r266_c116 bl[116] br[116] wl[266] vdd gnd cell_6t
Xbit_r267_c116 bl[116] br[116] wl[267] vdd gnd cell_6t
Xbit_r268_c116 bl[116] br[116] wl[268] vdd gnd cell_6t
Xbit_r269_c116 bl[116] br[116] wl[269] vdd gnd cell_6t
Xbit_r270_c116 bl[116] br[116] wl[270] vdd gnd cell_6t
Xbit_r271_c116 bl[116] br[116] wl[271] vdd gnd cell_6t
Xbit_r272_c116 bl[116] br[116] wl[272] vdd gnd cell_6t
Xbit_r273_c116 bl[116] br[116] wl[273] vdd gnd cell_6t
Xbit_r274_c116 bl[116] br[116] wl[274] vdd gnd cell_6t
Xbit_r275_c116 bl[116] br[116] wl[275] vdd gnd cell_6t
Xbit_r276_c116 bl[116] br[116] wl[276] vdd gnd cell_6t
Xbit_r277_c116 bl[116] br[116] wl[277] vdd gnd cell_6t
Xbit_r278_c116 bl[116] br[116] wl[278] vdd gnd cell_6t
Xbit_r279_c116 bl[116] br[116] wl[279] vdd gnd cell_6t
Xbit_r280_c116 bl[116] br[116] wl[280] vdd gnd cell_6t
Xbit_r281_c116 bl[116] br[116] wl[281] vdd gnd cell_6t
Xbit_r282_c116 bl[116] br[116] wl[282] vdd gnd cell_6t
Xbit_r283_c116 bl[116] br[116] wl[283] vdd gnd cell_6t
Xbit_r284_c116 bl[116] br[116] wl[284] vdd gnd cell_6t
Xbit_r285_c116 bl[116] br[116] wl[285] vdd gnd cell_6t
Xbit_r286_c116 bl[116] br[116] wl[286] vdd gnd cell_6t
Xbit_r287_c116 bl[116] br[116] wl[287] vdd gnd cell_6t
Xbit_r288_c116 bl[116] br[116] wl[288] vdd gnd cell_6t
Xbit_r289_c116 bl[116] br[116] wl[289] vdd gnd cell_6t
Xbit_r290_c116 bl[116] br[116] wl[290] vdd gnd cell_6t
Xbit_r291_c116 bl[116] br[116] wl[291] vdd gnd cell_6t
Xbit_r292_c116 bl[116] br[116] wl[292] vdd gnd cell_6t
Xbit_r293_c116 bl[116] br[116] wl[293] vdd gnd cell_6t
Xbit_r294_c116 bl[116] br[116] wl[294] vdd gnd cell_6t
Xbit_r295_c116 bl[116] br[116] wl[295] vdd gnd cell_6t
Xbit_r296_c116 bl[116] br[116] wl[296] vdd gnd cell_6t
Xbit_r297_c116 bl[116] br[116] wl[297] vdd gnd cell_6t
Xbit_r298_c116 bl[116] br[116] wl[298] vdd gnd cell_6t
Xbit_r299_c116 bl[116] br[116] wl[299] vdd gnd cell_6t
Xbit_r300_c116 bl[116] br[116] wl[300] vdd gnd cell_6t
Xbit_r301_c116 bl[116] br[116] wl[301] vdd gnd cell_6t
Xbit_r302_c116 bl[116] br[116] wl[302] vdd gnd cell_6t
Xbit_r303_c116 bl[116] br[116] wl[303] vdd gnd cell_6t
Xbit_r304_c116 bl[116] br[116] wl[304] vdd gnd cell_6t
Xbit_r305_c116 bl[116] br[116] wl[305] vdd gnd cell_6t
Xbit_r306_c116 bl[116] br[116] wl[306] vdd gnd cell_6t
Xbit_r307_c116 bl[116] br[116] wl[307] vdd gnd cell_6t
Xbit_r308_c116 bl[116] br[116] wl[308] vdd gnd cell_6t
Xbit_r309_c116 bl[116] br[116] wl[309] vdd gnd cell_6t
Xbit_r310_c116 bl[116] br[116] wl[310] vdd gnd cell_6t
Xbit_r311_c116 bl[116] br[116] wl[311] vdd gnd cell_6t
Xbit_r312_c116 bl[116] br[116] wl[312] vdd gnd cell_6t
Xbit_r313_c116 bl[116] br[116] wl[313] vdd gnd cell_6t
Xbit_r314_c116 bl[116] br[116] wl[314] vdd gnd cell_6t
Xbit_r315_c116 bl[116] br[116] wl[315] vdd gnd cell_6t
Xbit_r316_c116 bl[116] br[116] wl[316] vdd gnd cell_6t
Xbit_r317_c116 bl[116] br[116] wl[317] vdd gnd cell_6t
Xbit_r318_c116 bl[116] br[116] wl[318] vdd gnd cell_6t
Xbit_r319_c116 bl[116] br[116] wl[319] vdd gnd cell_6t
Xbit_r320_c116 bl[116] br[116] wl[320] vdd gnd cell_6t
Xbit_r321_c116 bl[116] br[116] wl[321] vdd gnd cell_6t
Xbit_r322_c116 bl[116] br[116] wl[322] vdd gnd cell_6t
Xbit_r323_c116 bl[116] br[116] wl[323] vdd gnd cell_6t
Xbit_r324_c116 bl[116] br[116] wl[324] vdd gnd cell_6t
Xbit_r325_c116 bl[116] br[116] wl[325] vdd gnd cell_6t
Xbit_r326_c116 bl[116] br[116] wl[326] vdd gnd cell_6t
Xbit_r327_c116 bl[116] br[116] wl[327] vdd gnd cell_6t
Xbit_r328_c116 bl[116] br[116] wl[328] vdd gnd cell_6t
Xbit_r329_c116 bl[116] br[116] wl[329] vdd gnd cell_6t
Xbit_r330_c116 bl[116] br[116] wl[330] vdd gnd cell_6t
Xbit_r331_c116 bl[116] br[116] wl[331] vdd gnd cell_6t
Xbit_r332_c116 bl[116] br[116] wl[332] vdd gnd cell_6t
Xbit_r333_c116 bl[116] br[116] wl[333] vdd gnd cell_6t
Xbit_r334_c116 bl[116] br[116] wl[334] vdd gnd cell_6t
Xbit_r335_c116 bl[116] br[116] wl[335] vdd gnd cell_6t
Xbit_r336_c116 bl[116] br[116] wl[336] vdd gnd cell_6t
Xbit_r337_c116 bl[116] br[116] wl[337] vdd gnd cell_6t
Xbit_r338_c116 bl[116] br[116] wl[338] vdd gnd cell_6t
Xbit_r339_c116 bl[116] br[116] wl[339] vdd gnd cell_6t
Xbit_r340_c116 bl[116] br[116] wl[340] vdd gnd cell_6t
Xbit_r341_c116 bl[116] br[116] wl[341] vdd gnd cell_6t
Xbit_r342_c116 bl[116] br[116] wl[342] vdd gnd cell_6t
Xbit_r343_c116 bl[116] br[116] wl[343] vdd gnd cell_6t
Xbit_r344_c116 bl[116] br[116] wl[344] vdd gnd cell_6t
Xbit_r345_c116 bl[116] br[116] wl[345] vdd gnd cell_6t
Xbit_r346_c116 bl[116] br[116] wl[346] vdd gnd cell_6t
Xbit_r347_c116 bl[116] br[116] wl[347] vdd gnd cell_6t
Xbit_r348_c116 bl[116] br[116] wl[348] vdd gnd cell_6t
Xbit_r349_c116 bl[116] br[116] wl[349] vdd gnd cell_6t
Xbit_r350_c116 bl[116] br[116] wl[350] vdd gnd cell_6t
Xbit_r351_c116 bl[116] br[116] wl[351] vdd gnd cell_6t
Xbit_r352_c116 bl[116] br[116] wl[352] vdd gnd cell_6t
Xbit_r353_c116 bl[116] br[116] wl[353] vdd gnd cell_6t
Xbit_r354_c116 bl[116] br[116] wl[354] vdd gnd cell_6t
Xbit_r355_c116 bl[116] br[116] wl[355] vdd gnd cell_6t
Xbit_r356_c116 bl[116] br[116] wl[356] vdd gnd cell_6t
Xbit_r357_c116 bl[116] br[116] wl[357] vdd gnd cell_6t
Xbit_r358_c116 bl[116] br[116] wl[358] vdd gnd cell_6t
Xbit_r359_c116 bl[116] br[116] wl[359] vdd gnd cell_6t
Xbit_r360_c116 bl[116] br[116] wl[360] vdd gnd cell_6t
Xbit_r361_c116 bl[116] br[116] wl[361] vdd gnd cell_6t
Xbit_r362_c116 bl[116] br[116] wl[362] vdd gnd cell_6t
Xbit_r363_c116 bl[116] br[116] wl[363] vdd gnd cell_6t
Xbit_r364_c116 bl[116] br[116] wl[364] vdd gnd cell_6t
Xbit_r365_c116 bl[116] br[116] wl[365] vdd gnd cell_6t
Xbit_r366_c116 bl[116] br[116] wl[366] vdd gnd cell_6t
Xbit_r367_c116 bl[116] br[116] wl[367] vdd gnd cell_6t
Xbit_r368_c116 bl[116] br[116] wl[368] vdd gnd cell_6t
Xbit_r369_c116 bl[116] br[116] wl[369] vdd gnd cell_6t
Xbit_r370_c116 bl[116] br[116] wl[370] vdd gnd cell_6t
Xbit_r371_c116 bl[116] br[116] wl[371] vdd gnd cell_6t
Xbit_r372_c116 bl[116] br[116] wl[372] vdd gnd cell_6t
Xbit_r373_c116 bl[116] br[116] wl[373] vdd gnd cell_6t
Xbit_r374_c116 bl[116] br[116] wl[374] vdd gnd cell_6t
Xbit_r375_c116 bl[116] br[116] wl[375] vdd gnd cell_6t
Xbit_r376_c116 bl[116] br[116] wl[376] vdd gnd cell_6t
Xbit_r377_c116 bl[116] br[116] wl[377] vdd gnd cell_6t
Xbit_r378_c116 bl[116] br[116] wl[378] vdd gnd cell_6t
Xbit_r379_c116 bl[116] br[116] wl[379] vdd gnd cell_6t
Xbit_r380_c116 bl[116] br[116] wl[380] vdd gnd cell_6t
Xbit_r381_c116 bl[116] br[116] wl[381] vdd gnd cell_6t
Xbit_r382_c116 bl[116] br[116] wl[382] vdd gnd cell_6t
Xbit_r383_c116 bl[116] br[116] wl[383] vdd gnd cell_6t
Xbit_r384_c116 bl[116] br[116] wl[384] vdd gnd cell_6t
Xbit_r385_c116 bl[116] br[116] wl[385] vdd gnd cell_6t
Xbit_r386_c116 bl[116] br[116] wl[386] vdd gnd cell_6t
Xbit_r387_c116 bl[116] br[116] wl[387] vdd gnd cell_6t
Xbit_r388_c116 bl[116] br[116] wl[388] vdd gnd cell_6t
Xbit_r389_c116 bl[116] br[116] wl[389] vdd gnd cell_6t
Xbit_r390_c116 bl[116] br[116] wl[390] vdd gnd cell_6t
Xbit_r391_c116 bl[116] br[116] wl[391] vdd gnd cell_6t
Xbit_r392_c116 bl[116] br[116] wl[392] vdd gnd cell_6t
Xbit_r393_c116 bl[116] br[116] wl[393] vdd gnd cell_6t
Xbit_r394_c116 bl[116] br[116] wl[394] vdd gnd cell_6t
Xbit_r395_c116 bl[116] br[116] wl[395] vdd gnd cell_6t
Xbit_r396_c116 bl[116] br[116] wl[396] vdd gnd cell_6t
Xbit_r397_c116 bl[116] br[116] wl[397] vdd gnd cell_6t
Xbit_r398_c116 bl[116] br[116] wl[398] vdd gnd cell_6t
Xbit_r399_c116 bl[116] br[116] wl[399] vdd gnd cell_6t
Xbit_r400_c116 bl[116] br[116] wl[400] vdd gnd cell_6t
Xbit_r401_c116 bl[116] br[116] wl[401] vdd gnd cell_6t
Xbit_r402_c116 bl[116] br[116] wl[402] vdd gnd cell_6t
Xbit_r403_c116 bl[116] br[116] wl[403] vdd gnd cell_6t
Xbit_r404_c116 bl[116] br[116] wl[404] vdd gnd cell_6t
Xbit_r405_c116 bl[116] br[116] wl[405] vdd gnd cell_6t
Xbit_r406_c116 bl[116] br[116] wl[406] vdd gnd cell_6t
Xbit_r407_c116 bl[116] br[116] wl[407] vdd gnd cell_6t
Xbit_r408_c116 bl[116] br[116] wl[408] vdd gnd cell_6t
Xbit_r409_c116 bl[116] br[116] wl[409] vdd gnd cell_6t
Xbit_r410_c116 bl[116] br[116] wl[410] vdd gnd cell_6t
Xbit_r411_c116 bl[116] br[116] wl[411] vdd gnd cell_6t
Xbit_r412_c116 bl[116] br[116] wl[412] vdd gnd cell_6t
Xbit_r413_c116 bl[116] br[116] wl[413] vdd gnd cell_6t
Xbit_r414_c116 bl[116] br[116] wl[414] vdd gnd cell_6t
Xbit_r415_c116 bl[116] br[116] wl[415] vdd gnd cell_6t
Xbit_r416_c116 bl[116] br[116] wl[416] vdd gnd cell_6t
Xbit_r417_c116 bl[116] br[116] wl[417] vdd gnd cell_6t
Xbit_r418_c116 bl[116] br[116] wl[418] vdd gnd cell_6t
Xbit_r419_c116 bl[116] br[116] wl[419] vdd gnd cell_6t
Xbit_r420_c116 bl[116] br[116] wl[420] vdd gnd cell_6t
Xbit_r421_c116 bl[116] br[116] wl[421] vdd gnd cell_6t
Xbit_r422_c116 bl[116] br[116] wl[422] vdd gnd cell_6t
Xbit_r423_c116 bl[116] br[116] wl[423] vdd gnd cell_6t
Xbit_r424_c116 bl[116] br[116] wl[424] vdd gnd cell_6t
Xbit_r425_c116 bl[116] br[116] wl[425] vdd gnd cell_6t
Xbit_r426_c116 bl[116] br[116] wl[426] vdd gnd cell_6t
Xbit_r427_c116 bl[116] br[116] wl[427] vdd gnd cell_6t
Xbit_r428_c116 bl[116] br[116] wl[428] vdd gnd cell_6t
Xbit_r429_c116 bl[116] br[116] wl[429] vdd gnd cell_6t
Xbit_r430_c116 bl[116] br[116] wl[430] vdd gnd cell_6t
Xbit_r431_c116 bl[116] br[116] wl[431] vdd gnd cell_6t
Xbit_r432_c116 bl[116] br[116] wl[432] vdd gnd cell_6t
Xbit_r433_c116 bl[116] br[116] wl[433] vdd gnd cell_6t
Xbit_r434_c116 bl[116] br[116] wl[434] vdd gnd cell_6t
Xbit_r435_c116 bl[116] br[116] wl[435] vdd gnd cell_6t
Xbit_r436_c116 bl[116] br[116] wl[436] vdd gnd cell_6t
Xbit_r437_c116 bl[116] br[116] wl[437] vdd gnd cell_6t
Xbit_r438_c116 bl[116] br[116] wl[438] vdd gnd cell_6t
Xbit_r439_c116 bl[116] br[116] wl[439] vdd gnd cell_6t
Xbit_r440_c116 bl[116] br[116] wl[440] vdd gnd cell_6t
Xbit_r441_c116 bl[116] br[116] wl[441] vdd gnd cell_6t
Xbit_r442_c116 bl[116] br[116] wl[442] vdd gnd cell_6t
Xbit_r443_c116 bl[116] br[116] wl[443] vdd gnd cell_6t
Xbit_r444_c116 bl[116] br[116] wl[444] vdd gnd cell_6t
Xbit_r445_c116 bl[116] br[116] wl[445] vdd gnd cell_6t
Xbit_r446_c116 bl[116] br[116] wl[446] vdd gnd cell_6t
Xbit_r447_c116 bl[116] br[116] wl[447] vdd gnd cell_6t
Xbit_r448_c116 bl[116] br[116] wl[448] vdd gnd cell_6t
Xbit_r449_c116 bl[116] br[116] wl[449] vdd gnd cell_6t
Xbit_r450_c116 bl[116] br[116] wl[450] vdd gnd cell_6t
Xbit_r451_c116 bl[116] br[116] wl[451] vdd gnd cell_6t
Xbit_r452_c116 bl[116] br[116] wl[452] vdd gnd cell_6t
Xbit_r453_c116 bl[116] br[116] wl[453] vdd gnd cell_6t
Xbit_r454_c116 bl[116] br[116] wl[454] vdd gnd cell_6t
Xbit_r455_c116 bl[116] br[116] wl[455] vdd gnd cell_6t
Xbit_r456_c116 bl[116] br[116] wl[456] vdd gnd cell_6t
Xbit_r457_c116 bl[116] br[116] wl[457] vdd gnd cell_6t
Xbit_r458_c116 bl[116] br[116] wl[458] vdd gnd cell_6t
Xbit_r459_c116 bl[116] br[116] wl[459] vdd gnd cell_6t
Xbit_r460_c116 bl[116] br[116] wl[460] vdd gnd cell_6t
Xbit_r461_c116 bl[116] br[116] wl[461] vdd gnd cell_6t
Xbit_r462_c116 bl[116] br[116] wl[462] vdd gnd cell_6t
Xbit_r463_c116 bl[116] br[116] wl[463] vdd gnd cell_6t
Xbit_r464_c116 bl[116] br[116] wl[464] vdd gnd cell_6t
Xbit_r465_c116 bl[116] br[116] wl[465] vdd gnd cell_6t
Xbit_r466_c116 bl[116] br[116] wl[466] vdd gnd cell_6t
Xbit_r467_c116 bl[116] br[116] wl[467] vdd gnd cell_6t
Xbit_r468_c116 bl[116] br[116] wl[468] vdd gnd cell_6t
Xbit_r469_c116 bl[116] br[116] wl[469] vdd gnd cell_6t
Xbit_r470_c116 bl[116] br[116] wl[470] vdd gnd cell_6t
Xbit_r471_c116 bl[116] br[116] wl[471] vdd gnd cell_6t
Xbit_r472_c116 bl[116] br[116] wl[472] vdd gnd cell_6t
Xbit_r473_c116 bl[116] br[116] wl[473] vdd gnd cell_6t
Xbit_r474_c116 bl[116] br[116] wl[474] vdd gnd cell_6t
Xbit_r475_c116 bl[116] br[116] wl[475] vdd gnd cell_6t
Xbit_r476_c116 bl[116] br[116] wl[476] vdd gnd cell_6t
Xbit_r477_c116 bl[116] br[116] wl[477] vdd gnd cell_6t
Xbit_r478_c116 bl[116] br[116] wl[478] vdd gnd cell_6t
Xbit_r479_c116 bl[116] br[116] wl[479] vdd gnd cell_6t
Xbit_r480_c116 bl[116] br[116] wl[480] vdd gnd cell_6t
Xbit_r481_c116 bl[116] br[116] wl[481] vdd gnd cell_6t
Xbit_r482_c116 bl[116] br[116] wl[482] vdd gnd cell_6t
Xbit_r483_c116 bl[116] br[116] wl[483] vdd gnd cell_6t
Xbit_r484_c116 bl[116] br[116] wl[484] vdd gnd cell_6t
Xbit_r485_c116 bl[116] br[116] wl[485] vdd gnd cell_6t
Xbit_r486_c116 bl[116] br[116] wl[486] vdd gnd cell_6t
Xbit_r487_c116 bl[116] br[116] wl[487] vdd gnd cell_6t
Xbit_r488_c116 bl[116] br[116] wl[488] vdd gnd cell_6t
Xbit_r489_c116 bl[116] br[116] wl[489] vdd gnd cell_6t
Xbit_r490_c116 bl[116] br[116] wl[490] vdd gnd cell_6t
Xbit_r491_c116 bl[116] br[116] wl[491] vdd gnd cell_6t
Xbit_r492_c116 bl[116] br[116] wl[492] vdd gnd cell_6t
Xbit_r493_c116 bl[116] br[116] wl[493] vdd gnd cell_6t
Xbit_r494_c116 bl[116] br[116] wl[494] vdd gnd cell_6t
Xbit_r495_c116 bl[116] br[116] wl[495] vdd gnd cell_6t
Xbit_r496_c116 bl[116] br[116] wl[496] vdd gnd cell_6t
Xbit_r497_c116 bl[116] br[116] wl[497] vdd gnd cell_6t
Xbit_r498_c116 bl[116] br[116] wl[498] vdd gnd cell_6t
Xbit_r499_c116 bl[116] br[116] wl[499] vdd gnd cell_6t
Xbit_r500_c116 bl[116] br[116] wl[500] vdd gnd cell_6t
Xbit_r501_c116 bl[116] br[116] wl[501] vdd gnd cell_6t
Xbit_r502_c116 bl[116] br[116] wl[502] vdd gnd cell_6t
Xbit_r503_c116 bl[116] br[116] wl[503] vdd gnd cell_6t
Xbit_r504_c116 bl[116] br[116] wl[504] vdd gnd cell_6t
Xbit_r505_c116 bl[116] br[116] wl[505] vdd gnd cell_6t
Xbit_r506_c116 bl[116] br[116] wl[506] vdd gnd cell_6t
Xbit_r507_c116 bl[116] br[116] wl[507] vdd gnd cell_6t
Xbit_r508_c116 bl[116] br[116] wl[508] vdd gnd cell_6t
Xbit_r509_c116 bl[116] br[116] wl[509] vdd gnd cell_6t
Xbit_r510_c116 bl[116] br[116] wl[510] vdd gnd cell_6t
Xbit_r511_c116 bl[116] br[116] wl[511] vdd gnd cell_6t
Xbit_r0_c117 bl[117] br[117] wl[0] vdd gnd cell_6t
Xbit_r1_c117 bl[117] br[117] wl[1] vdd gnd cell_6t
Xbit_r2_c117 bl[117] br[117] wl[2] vdd gnd cell_6t
Xbit_r3_c117 bl[117] br[117] wl[3] vdd gnd cell_6t
Xbit_r4_c117 bl[117] br[117] wl[4] vdd gnd cell_6t
Xbit_r5_c117 bl[117] br[117] wl[5] vdd gnd cell_6t
Xbit_r6_c117 bl[117] br[117] wl[6] vdd gnd cell_6t
Xbit_r7_c117 bl[117] br[117] wl[7] vdd gnd cell_6t
Xbit_r8_c117 bl[117] br[117] wl[8] vdd gnd cell_6t
Xbit_r9_c117 bl[117] br[117] wl[9] vdd gnd cell_6t
Xbit_r10_c117 bl[117] br[117] wl[10] vdd gnd cell_6t
Xbit_r11_c117 bl[117] br[117] wl[11] vdd gnd cell_6t
Xbit_r12_c117 bl[117] br[117] wl[12] vdd gnd cell_6t
Xbit_r13_c117 bl[117] br[117] wl[13] vdd gnd cell_6t
Xbit_r14_c117 bl[117] br[117] wl[14] vdd gnd cell_6t
Xbit_r15_c117 bl[117] br[117] wl[15] vdd gnd cell_6t
Xbit_r16_c117 bl[117] br[117] wl[16] vdd gnd cell_6t
Xbit_r17_c117 bl[117] br[117] wl[17] vdd gnd cell_6t
Xbit_r18_c117 bl[117] br[117] wl[18] vdd gnd cell_6t
Xbit_r19_c117 bl[117] br[117] wl[19] vdd gnd cell_6t
Xbit_r20_c117 bl[117] br[117] wl[20] vdd gnd cell_6t
Xbit_r21_c117 bl[117] br[117] wl[21] vdd gnd cell_6t
Xbit_r22_c117 bl[117] br[117] wl[22] vdd gnd cell_6t
Xbit_r23_c117 bl[117] br[117] wl[23] vdd gnd cell_6t
Xbit_r24_c117 bl[117] br[117] wl[24] vdd gnd cell_6t
Xbit_r25_c117 bl[117] br[117] wl[25] vdd gnd cell_6t
Xbit_r26_c117 bl[117] br[117] wl[26] vdd gnd cell_6t
Xbit_r27_c117 bl[117] br[117] wl[27] vdd gnd cell_6t
Xbit_r28_c117 bl[117] br[117] wl[28] vdd gnd cell_6t
Xbit_r29_c117 bl[117] br[117] wl[29] vdd gnd cell_6t
Xbit_r30_c117 bl[117] br[117] wl[30] vdd gnd cell_6t
Xbit_r31_c117 bl[117] br[117] wl[31] vdd gnd cell_6t
Xbit_r32_c117 bl[117] br[117] wl[32] vdd gnd cell_6t
Xbit_r33_c117 bl[117] br[117] wl[33] vdd gnd cell_6t
Xbit_r34_c117 bl[117] br[117] wl[34] vdd gnd cell_6t
Xbit_r35_c117 bl[117] br[117] wl[35] vdd gnd cell_6t
Xbit_r36_c117 bl[117] br[117] wl[36] vdd gnd cell_6t
Xbit_r37_c117 bl[117] br[117] wl[37] vdd gnd cell_6t
Xbit_r38_c117 bl[117] br[117] wl[38] vdd gnd cell_6t
Xbit_r39_c117 bl[117] br[117] wl[39] vdd gnd cell_6t
Xbit_r40_c117 bl[117] br[117] wl[40] vdd gnd cell_6t
Xbit_r41_c117 bl[117] br[117] wl[41] vdd gnd cell_6t
Xbit_r42_c117 bl[117] br[117] wl[42] vdd gnd cell_6t
Xbit_r43_c117 bl[117] br[117] wl[43] vdd gnd cell_6t
Xbit_r44_c117 bl[117] br[117] wl[44] vdd gnd cell_6t
Xbit_r45_c117 bl[117] br[117] wl[45] vdd gnd cell_6t
Xbit_r46_c117 bl[117] br[117] wl[46] vdd gnd cell_6t
Xbit_r47_c117 bl[117] br[117] wl[47] vdd gnd cell_6t
Xbit_r48_c117 bl[117] br[117] wl[48] vdd gnd cell_6t
Xbit_r49_c117 bl[117] br[117] wl[49] vdd gnd cell_6t
Xbit_r50_c117 bl[117] br[117] wl[50] vdd gnd cell_6t
Xbit_r51_c117 bl[117] br[117] wl[51] vdd gnd cell_6t
Xbit_r52_c117 bl[117] br[117] wl[52] vdd gnd cell_6t
Xbit_r53_c117 bl[117] br[117] wl[53] vdd gnd cell_6t
Xbit_r54_c117 bl[117] br[117] wl[54] vdd gnd cell_6t
Xbit_r55_c117 bl[117] br[117] wl[55] vdd gnd cell_6t
Xbit_r56_c117 bl[117] br[117] wl[56] vdd gnd cell_6t
Xbit_r57_c117 bl[117] br[117] wl[57] vdd gnd cell_6t
Xbit_r58_c117 bl[117] br[117] wl[58] vdd gnd cell_6t
Xbit_r59_c117 bl[117] br[117] wl[59] vdd gnd cell_6t
Xbit_r60_c117 bl[117] br[117] wl[60] vdd gnd cell_6t
Xbit_r61_c117 bl[117] br[117] wl[61] vdd gnd cell_6t
Xbit_r62_c117 bl[117] br[117] wl[62] vdd gnd cell_6t
Xbit_r63_c117 bl[117] br[117] wl[63] vdd gnd cell_6t
Xbit_r64_c117 bl[117] br[117] wl[64] vdd gnd cell_6t
Xbit_r65_c117 bl[117] br[117] wl[65] vdd gnd cell_6t
Xbit_r66_c117 bl[117] br[117] wl[66] vdd gnd cell_6t
Xbit_r67_c117 bl[117] br[117] wl[67] vdd gnd cell_6t
Xbit_r68_c117 bl[117] br[117] wl[68] vdd gnd cell_6t
Xbit_r69_c117 bl[117] br[117] wl[69] vdd gnd cell_6t
Xbit_r70_c117 bl[117] br[117] wl[70] vdd gnd cell_6t
Xbit_r71_c117 bl[117] br[117] wl[71] vdd gnd cell_6t
Xbit_r72_c117 bl[117] br[117] wl[72] vdd gnd cell_6t
Xbit_r73_c117 bl[117] br[117] wl[73] vdd gnd cell_6t
Xbit_r74_c117 bl[117] br[117] wl[74] vdd gnd cell_6t
Xbit_r75_c117 bl[117] br[117] wl[75] vdd gnd cell_6t
Xbit_r76_c117 bl[117] br[117] wl[76] vdd gnd cell_6t
Xbit_r77_c117 bl[117] br[117] wl[77] vdd gnd cell_6t
Xbit_r78_c117 bl[117] br[117] wl[78] vdd gnd cell_6t
Xbit_r79_c117 bl[117] br[117] wl[79] vdd gnd cell_6t
Xbit_r80_c117 bl[117] br[117] wl[80] vdd gnd cell_6t
Xbit_r81_c117 bl[117] br[117] wl[81] vdd gnd cell_6t
Xbit_r82_c117 bl[117] br[117] wl[82] vdd gnd cell_6t
Xbit_r83_c117 bl[117] br[117] wl[83] vdd gnd cell_6t
Xbit_r84_c117 bl[117] br[117] wl[84] vdd gnd cell_6t
Xbit_r85_c117 bl[117] br[117] wl[85] vdd gnd cell_6t
Xbit_r86_c117 bl[117] br[117] wl[86] vdd gnd cell_6t
Xbit_r87_c117 bl[117] br[117] wl[87] vdd gnd cell_6t
Xbit_r88_c117 bl[117] br[117] wl[88] vdd gnd cell_6t
Xbit_r89_c117 bl[117] br[117] wl[89] vdd gnd cell_6t
Xbit_r90_c117 bl[117] br[117] wl[90] vdd gnd cell_6t
Xbit_r91_c117 bl[117] br[117] wl[91] vdd gnd cell_6t
Xbit_r92_c117 bl[117] br[117] wl[92] vdd gnd cell_6t
Xbit_r93_c117 bl[117] br[117] wl[93] vdd gnd cell_6t
Xbit_r94_c117 bl[117] br[117] wl[94] vdd gnd cell_6t
Xbit_r95_c117 bl[117] br[117] wl[95] vdd gnd cell_6t
Xbit_r96_c117 bl[117] br[117] wl[96] vdd gnd cell_6t
Xbit_r97_c117 bl[117] br[117] wl[97] vdd gnd cell_6t
Xbit_r98_c117 bl[117] br[117] wl[98] vdd gnd cell_6t
Xbit_r99_c117 bl[117] br[117] wl[99] vdd gnd cell_6t
Xbit_r100_c117 bl[117] br[117] wl[100] vdd gnd cell_6t
Xbit_r101_c117 bl[117] br[117] wl[101] vdd gnd cell_6t
Xbit_r102_c117 bl[117] br[117] wl[102] vdd gnd cell_6t
Xbit_r103_c117 bl[117] br[117] wl[103] vdd gnd cell_6t
Xbit_r104_c117 bl[117] br[117] wl[104] vdd gnd cell_6t
Xbit_r105_c117 bl[117] br[117] wl[105] vdd gnd cell_6t
Xbit_r106_c117 bl[117] br[117] wl[106] vdd gnd cell_6t
Xbit_r107_c117 bl[117] br[117] wl[107] vdd gnd cell_6t
Xbit_r108_c117 bl[117] br[117] wl[108] vdd gnd cell_6t
Xbit_r109_c117 bl[117] br[117] wl[109] vdd gnd cell_6t
Xbit_r110_c117 bl[117] br[117] wl[110] vdd gnd cell_6t
Xbit_r111_c117 bl[117] br[117] wl[111] vdd gnd cell_6t
Xbit_r112_c117 bl[117] br[117] wl[112] vdd gnd cell_6t
Xbit_r113_c117 bl[117] br[117] wl[113] vdd gnd cell_6t
Xbit_r114_c117 bl[117] br[117] wl[114] vdd gnd cell_6t
Xbit_r115_c117 bl[117] br[117] wl[115] vdd gnd cell_6t
Xbit_r116_c117 bl[117] br[117] wl[116] vdd gnd cell_6t
Xbit_r117_c117 bl[117] br[117] wl[117] vdd gnd cell_6t
Xbit_r118_c117 bl[117] br[117] wl[118] vdd gnd cell_6t
Xbit_r119_c117 bl[117] br[117] wl[119] vdd gnd cell_6t
Xbit_r120_c117 bl[117] br[117] wl[120] vdd gnd cell_6t
Xbit_r121_c117 bl[117] br[117] wl[121] vdd gnd cell_6t
Xbit_r122_c117 bl[117] br[117] wl[122] vdd gnd cell_6t
Xbit_r123_c117 bl[117] br[117] wl[123] vdd gnd cell_6t
Xbit_r124_c117 bl[117] br[117] wl[124] vdd gnd cell_6t
Xbit_r125_c117 bl[117] br[117] wl[125] vdd gnd cell_6t
Xbit_r126_c117 bl[117] br[117] wl[126] vdd gnd cell_6t
Xbit_r127_c117 bl[117] br[117] wl[127] vdd gnd cell_6t
Xbit_r128_c117 bl[117] br[117] wl[128] vdd gnd cell_6t
Xbit_r129_c117 bl[117] br[117] wl[129] vdd gnd cell_6t
Xbit_r130_c117 bl[117] br[117] wl[130] vdd gnd cell_6t
Xbit_r131_c117 bl[117] br[117] wl[131] vdd gnd cell_6t
Xbit_r132_c117 bl[117] br[117] wl[132] vdd gnd cell_6t
Xbit_r133_c117 bl[117] br[117] wl[133] vdd gnd cell_6t
Xbit_r134_c117 bl[117] br[117] wl[134] vdd gnd cell_6t
Xbit_r135_c117 bl[117] br[117] wl[135] vdd gnd cell_6t
Xbit_r136_c117 bl[117] br[117] wl[136] vdd gnd cell_6t
Xbit_r137_c117 bl[117] br[117] wl[137] vdd gnd cell_6t
Xbit_r138_c117 bl[117] br[117] wl[138] vdd gnd cell_6t
Xbit_r139_c117 bl[117] br[117] wl[139] vdd gnd cell_6t
Xbit_r140_c117 bl[117] br[117] wl[140] vdd gnd cell_6t
Xbit_r141_c117 bl[117] br[117] wl[141] vdd gnd cell_6t
Xbit_r142_c117 bl[117] br[117] wl[142] vdd gnd cell_6t
Xbit_r143_c117 bl[117] br[117] wl[143] vdd gnd cell_6t
Xbit_r144_c117 bl[117] br[117] wl[144] vdd gnd cell_6t
Xbit_r145_c117 bl[117] br[117] wl[145] vdd gnd cell_6t
Xbit_r146_c117 bl[117] br[117] wl[146] vdd gnd cell_6t
Xbit_r147_c117 bl[117] br[117] wl[147] vdd gnd cell_6t
Xbit_r148_c117 bl[117] br[117] wl[148] vdd gnd cell_6t
Xbit_r149_c117 bl[117] br[117] wl[149] vdd gnd cell_6t
Xbit_r150_c117 bl[117] br[117] wl[150] vdd gnd cell_6t
Xbit_r151_c117 bl[117] br[117] wl[151] vdd gnd cell_6t
Xbit_r152_c117 bl[117] br[117] wl[152] vdd gnd cell_6t
Xbit_r153_c117 bl[117] br[117] wl[153] vdd gnd cell_6t
Xbit_r154_c117 bl[117] br[117] wl[154] vdd gnd cell_6t
Xbit_r155_c117 bl[117] br[117] wl[155] vdd gnd cell_6t
Xbit_r156_c117 bl[117] br[117] wl[156] vdd gnd cell_6t
Xbit_r157_c117 bl[117] br[117] wl[157] vdd gnd cell_6t
Xbit_r158_c117 bl[117] br[117] wl[158] vdd gnd cell_6t
Xbit_r159_c117 bl[117] br[117] wl[159] vdd gnd cell_6t
Xbit_r160_c117 bl[117] br[117] wl[160] vdd gnd cell_6t
Xbit_r161_c117 bl[117] br[117] wl[161] vdd gnd cell_6t
Xbit_r162_c117 bl[117] br[117] wl[162] vdd gnd cell_6t
Xbit_r163_c117 bl[117] br[117] wl[163] vdd gnd cell_6t
Xbit_r164_c117 bl[117] br[117] wl[164] vdd gnd cell_6t
Xbit_r165_c117 bl[117] br[117] wl[165] vdd gnd cell_6t
Xbit_r166_c117 bl[117] br[117] wl[166] vdd gnd cell_6t
Xbit_r167_c117 bl[117] br[117] wl[167] vdd gnd cell_6t
Xbit_r168_c117 bl[117] br[117] wl[168] vdd gnd cell_6t
Xbit_r169_c117 bl[117] br[117] wl[169] vdd gnd cell_6t
Xbit_r170_c117 bl[117] br[117] wl[170] vdd gnd cell_6t
Xbit_r171_c117 bl[117] br[117] wl[171] vdd gnd cell_6t
Xbit_r172_c117 bl[117] br[117] wl[172] vdd gnd cell_6t
Xbit_r173_c117 bl[117] br[117] wl[173] vdd gnd cell_6t
Xbit_r174_c117 bl[117] br[117] wl[174] vdd gnd cell_6t
Xbit_r175_c117 bl[117] br[117] wl[175] vdd gnd cell_6t
Xbit_r176_c117 bl[117] br[117] wl[176] vdd gnd cell_6t
Xbit_r177_c117 bl[117] br[117] wl[177] vdd gnd cell_6t
Xbit_r178_c117 bl[117] br[117] wl[178] vdd gnd cell_6t
Xbit_r179_c117 bl[117] br[117] wl[179] vdd gnd cell_6t
Xbit_r180_c117 bl[117] br[117] wl[180] vdd gnd cell_6t
Xbit_r181_c117 bl[117] br[117] wl[181] vdd gnd cell_6t
Xbit_r182_c117 bl[117] br[117] wl[182] vdd gnd cell_6t
Xbit_r183_c117 bl[117] br[117] wl[183] vdd gnd cell_6t
Xbit_r184_c117 bl[117] br[117] wl[184] vdd gnd cell_6t
Xbit_r185_c117 bl[117] br[117] wl[185] vdd gnd cell_6t
Xbit_r186_c117 bl[117] br[117] wl[186] vdd gnd cell_6t
Xbit_r187_c117 bl[117] br[117] wl[187] vdd gnd cell_6t
Xbit_r188_c117 bl[117] br[117] wl[188] vdd gnd cell_6t
Xbit_r189_c117 bl[117] br[117] wl[189] vdd gnd cell_6t
Xbit_r190_c117 bl[117] br[117] wl[190] vdd gnd cell_6t
Xbit_r191_c117 bl[117] br[117] wl[191] vdd gnd cell_6t
Xbit_r192_c117 bl[117] br[117] wl[192] vdd gnd cell_6t
Xbit_r193_c117 bl[117] br[117] wl[193] vdd gnd cell_6t
Xbit_r194_c117 bl[117] br[117] wl[194] vdd gnd cell_6t
Xbit_r195_c117 bl[117] br[117] wl[195] vdd gnd cell_6t
Xbit_r196_c117 bl[117] br[117] wl[196] vdd gnd cell_6t
Xbit_r197_c117 bl[117] br[117] wl[197] vdd gnd cell_6t
Xbit_r198_c117 bl[117] br[117] wl[198] vdd gnd cell_6t
Xbit_r199_c117 bl[117] br[117] wl[199] vdd gnd cell_6t
Xbit_r200_c117 bl[117] br[117] wl[200] vdd gnd cell_6t
Xbit_r201_c117 bl[117] br[117] wl[201] vdd gnd cell_6t
Xbit_r202_c117 bl[117] br[117] wl[202] vdd gnd cell_6t
Xbit_r203_c117 bl[117] br[117] wl[203] vdd gnd cell_6t
Xbit_r204_c117 bl[117] br[117] wl[204] vdd gnd cell_6t
Xbit_r205_c117 bl[117] br[117] wl[205] vdd gnd cell_6t
Xbit_r206_c117 bl[117] br[117] wl[206] vdd gnd cell_6t
Xbit_r207_c117 bl[117] br[117] wl[207] vdd gnd cell_6t
Xbit_r208_c117 bl[117] br[117] wl[208] vdd gnd cell_6t
Xbit_r209_c117 bl[117] br[117] wl[209] vdd gnd cell_6t
Xbit_r210_c117 bl[117] br[117] wl[210] vdd gnd cell_6t
Xbit_r211_c117 bl[117] br[117] wl[211] vdd gnd cell_6t
Xbit_r212_c117 bl[117] br[117] wl[212] vdd gnd cell_6t
Xbit_r213_c117 bl[117] br[117] wl[213] vdd gnd cell_6t
Xbit_r214_c117 bl[117] br[117] wl[214] vdd gnd cell_6t
Xbit_r215_c117 bl[117] br[117] wl[215] vdd gnd cell_6t
Xbit_r216_c117 bl[117] br[117] wl[216] vdd gnd cell_6t
Xbit_r217_c117 bl[117] br[117] wl[217] vdd gnd cell_6t
Xbit_r218_c117 bl[117] br[117] wl[218] vdd gnd cell_6t
Xbit_r219_c117 bl[117] br[117] wl[219] vdd gnd cell_6t
Xbit_r220_c117 bl[117] br[117] wl[220] vdd gnd cell_6t
Xbit_r221_c117 bl[117] br[117] wl[221] vdd gnd cell_6t
Xbit_r222_c117 bl[117] br[117] wl[222] vdd gnd cell_6t
Xbit_r223_c117 bl[117] br[117] wl[223] vdd gnd cell_6t
Xbit_r224_c117 bl[117] br[117] wl[224] vdd gnd cell_6t
Xbit_r225_c117 bl[117] br[117] wl[225] vdd gnd cell_6t
Xbit_r226_c117 bl[117] br[117] wl[226] vdd gnd cell_6t
Xbit_r227_c117 bl[117] br[117] wl[227] vdd gnd cell_6t
Xbit_r228_c117 bl[117] br[117] wl[228] vdd gnd cell_6t
Xbit_r229_c117 bl[117] br[117] wl[229] vdd gnd cell_6t
Xbit_r230_c117 bl[117] br[117] wl[230] vdd gnd cell_6t
Xbit_r231_c117 bl[117] br[117] wl[231] vdd gnd cell_6t
Xbit_r232_c117 bl[117] br[117] wl[232] vdd gnd cell_6t
Xbit_r233_c117 bl[117] br[117] wl[233] vdd gnd cell_6t
Xbit_r234_c117 bl[117] br[117] wl[234] vdd gnd cell_6t
Xbit_r235_c117 bl[117] br[117] wl[235] vdd gnd cell_6t
Xbit_r236_c117 bl[117] br[117] wl[236] vdd gnd cell_6t
Xbit_r237_c117 bl[117] br[117] wl[237] vdd gnd cell_6t
Xbit_r238_c117 bl[117] br[117] wl[238] vdd gnd cell_6t
Xbit_r239_c117 bl[117] br[117] wl[239] vdd gnd cell_6t
Xbit_r240_c117 bl[117] br[117] wl[240] vdd gnd cell_6t
Xbit_r241_c117 bl[117] br[117] wl[241] vdd gnd cell_6t
Xbit_r242_c117 bl[117] br[117] wl[242] vdd gnd cell_6t
Xbit_r243_c117 bl[117] br[117] wl[243] vdd gnd cell_6t
Xbit_r244_c117 bl[117] br[117] wl[244] vdd gnd cell_6t
Xbit_r245_c117 bl[117] br[117] wl[245] vdd gnd cell_6t
Xbit_r246_c117 bl[117] br[117] wl[246] vdd gnd cell_6t
Xbit_r247_c117 bl[117] br[117] wl[247] vdd gnd cell_6t
Xbit_r248_c117 bl[117] br[117] wl[248] vdd gnd cell_6t
Xbit_r249_c117 bl[117] br[117] wl[249] vdd gnd cell_6t
Xbit_r250_c117 bl[117] br[117] wl[250] vdd gnd cell_6t
Xbit_r251_c117 bl[117] br[117] wl[251] vdd gnd cell_6t
Xbit_r252_c117 bl[117] br[117] wl[252] vdd gnd cell_6t
Xbit_r253_c117 bl[117] br[117] wl[253] vdd gnd cell_6t
Xbit_r254_c117 bl[117] br[117] wl[254] vdd gnd cell_6t
Xbit_r255_c117 bl[117] br[117] wl[255] vdd gnd cell_6t
Xbit_r256_c117 bl[117] br[117] wl[256] vdd gnd cell_6t
Xbit_r257_c117 bl[117] br[117] wl[257] vdd gnd cell_6t
Xbit_r258_c117 bl[117] br[117] wl[258] vdd gnd cell_6t
Xbit_r259_c117 bl[117] br[117] wl[259] vdd gnd cell_6t
Xbit_r260_c117 bl[117] br[117] wl[260] vdd gnd cell_6t
Xbit_r261_c117 bl[117] br[117] wl[261] vdd gnd cell_6t
Xbit_r262_c117 bl[117] br[117] wl[262] vdd gnd cell_6t
Xbit_r263_c117 bl[117] br[117] wl[263] vdd gnd cell_6t
Xbit_r264_c117 bl[117] br[117] wl[264] vdd gnd cell_6t
Xbit_r265_c117 bl[117] br[117] wl[265] vdd gnd cell_6t
Xbit_r266_c117 bl[117] br[117] wl[266] vdd gnd cell_6t
Xbit_r267_c117 bl[117] br[117] wl[267] vdd gnd cell_6t
Xbit_r268_c117 bl[117] br[117] wl[268] vdd gnd cell_6t
Xbit_r269_c117 bl[117] br[117] wl[269] vdd gnd cell_6t
Xbit_r270_c117 bl[117] br[117] wl[270] vdd gnd cell_6t
Xbit_r271_c117 bl[117] br[117] wl[271] vdd gnd cell_6t
Xbit_r272_c117 bl[117] br[117] wl[272] vdd gnd cell_6t
Xbit_r273_c117 bl[117] br[117] wl[273] vdd gnd cell_6t
Xbit_r274_c117 bl[117] br[117] wl[274] vdd gnd cell_6t
Xbit_r275_c117 bl[117] br[117] wl[275] vdd gnd cell_6t
Xbit_r276_c117 bl[117] br[117] wl[276] vdd gnd cell_6t
Xbit_r277_c117 bl[117] br[117] wl[277] vdd gnd cell_6t
Xbit_r278_c117 bl[117] br[117] wl[278] vdd gnd cell_6t
Xbit_r279_c117 bl[117] br[117] wl[279] vdd gnd cell_6t
Xbit_r280_c117 bl[117] br[117] wl[280] vdd gnd cell_6t
Xbit_r281_c117 bl[117] br[117] wl[281] vdd gnd cell_6t
Xbit_r282_c117 bl[117] br[117] wl[282] vdd gnd cell_6t
Xbit_r283_c117 bl[117] br[117] wl[283] vdd gnd cell_6t
Xbit_r284_c117 bl[117] br[117] wl[284] vdd gnd cell_6t
Xbit_r285_c117 bl[117] br[117] wl[285] vdd gnd cell_6t
Xbit_r286_c117 bl[117] br[117] wl[286] vdd gnd cell_6t
Xbit_r287_c117 bl[117] br[117] wl[287] vdd gnd cell_6t
Xbit_r288_c117 bl[117] br[117] wl[288] vdd gnd cell_6t
Xbit_r289_c117 bl[117] br[117] wl[289] vdd gnd cell_6t
Xbit_r290_c117 bl[117] br[117] wl[290] vdd gnd cell_6t
Xbit_r291_c117 bl[117] br[117] wl[291] vdd gnd cell_6t
Xbit_r292_c117 bl[117] br[117] wl[292] vdd gnd cell_6t
Xbit_r293_c117 bl[117] br[117] wl[293] vdd gnd cell_6t
Xbit_r294_c117 bl[117] br[117] wl[294] vdd gnd cell_6t
Xbit_r295_c117 bl[117] br[117] wl[295] vdd gnd cell_6t
Xbit_r296_c117 bl[117] br[117] wl[296] vdd gnd cell_6t
Xbit_r297_c117 bl[117] br[117] wl[297] vdd gnd cell_6t
Xbit_r298_c117 bl[117] br[117] wl[298] vdd gnd cell_6t
Xbit_r299_c117 bl[117] br[117] wl[299] vdd gnd cell_6t
Xbit_r300_c117 bl[117] br[117] wl[300] vdd gnd cell_6t
Xbit_r301_c117 bl[117] br[117] wl[301] vdd gnd cell_6t
Xbit_r302_c117 bl[117] br[117] wl[302] vdd gnd cell_6t
Xbit_r303_c117 bl[117] br[117] wl[303] vdd gnd cell_6t
Xbit_r304_c117 bl[117] br[117] wl[304] vdd gnd cell_6t
Xbit_r305_c117 bl[117] br[117] wl[305] vdd gnd cell_6t
Xbit_r306_c117 bl[117] br[117] wl[306] vdd gnd cell_6t
Xbit_r307_c117 bl[117] br[117] wl[307] vdd gnd cell_6t
Xbit_r308_c117 bl[117] br[117] wl[308] vdd gnd cell_6t
Xbit_r309_c117 bl[117] br[117] wl[309] vdd gnd cell_6t
Xbit_r310_c117 bl[117] br[117] wl[310] vdd gnd cell_6t
Xbit_r311_c117 bl[117] br[117] wl[311] vdd gnd cell_6t
Xbit_r312_c117 bl[117] br[117] wl[312] vdd gnd cell_6t
Xbit_r313_c117 bl[117] br[117] wl[313] vdd gnd cell_6t
Xbit_r314_c117 bl[117] br[117] wl[314] vdd gnd cell_6t
Xbit_r315_c117 bl[117] br[117] wl[315] vdd gnd cell_6t
Xbit_r316_c117 bl[117] br[117] wl[316] vdd gnd cell_6t
Xbit_r317_c117 bl[117] br[117] wl[317] vdd gnd cell_6t
Xbit_r318_c117 bl[117] br[117] wl[318] vdd gnd cell_6t
Xbit_r319_c117 bl[117] br[117] wl[319] vdd gnd cell_6t
Xbit_r320_c117 bl[117] br[117] wl[320] vdd gnd cell_6t
Xbit_r321_c117 bl[117] br[117] wl[321] vdd gnd cell_6t
Xbit_r322_c117 bl[117] br[117] wl[322] vdd gnd cell_6t
Xbit_r323_c117 bl[117] br[117] wl[323] vdd gnd cell_6t
Xbit_r324_c117 bl[117] br[117] wl[324] vdd gnd cell_6t
Xbit_r325_c117 bl[117] br[117] wl[325] vdd gnd cell_6t
Xbit_r326_c117 bl[117] br[117] wl[326] vdd gnd cell_6t
Xbit_r327_c117 bl[117] br[117] wl[327] vdd gnd cell_6t
Xbit_r328_c117 bl[117] br[117] wl[328] vdd gnd cell_6t
Xbit_r329_c117 bl[117] br[117] wl[329] vdd gnd cell_6t
Xbit_r330_c117 bl[117] br[117] wl[330] vdd gnd cell_6t
Xbit_r331_c117 bl[117] br[117] wl[331] vdd gnd cell_6t
Xbit_r332_c117 bl[117] br[117] wl[332] vdd gnd cell_6t
Xbit_r333_c117 bl[117] br[117] wl[333] vdd gnd cell_6t
Xbit_r334_c117 bl[117] br[117] wl[334] vdd gnd cell_6t
Xbit_r335_c117 bl[117] br[117] wl[335] vdd gnd cell_6t
Xbit_r336_c117 bl[117] br[117] wl[336] vdd gnd cell_6t
Xbit_r337_c117 bl[117] br[117] wl[337] vdd gnd cell_6t
Xbit_r338_c117 bl[117] br[117] wl[338] vdd gnd cell_6t
Xbit_r339_c117 bl[117] br[117] wl[339] vdd gnd cell_6t
Xbit_r340_c117 bl[117] br[117] wl[340] vdd gnd cell_6t
Xbit_r341_c117 bl[117] br[117] wl[341] vdd gnd cell_6t
Xbit_r342_c117 bl[117] br[117] wl[342] vdd gnd cell_6t
Xbit_r343_c117 bl[117] br[117] wl[343] vdd gnd cell_6t
Xbit_r344_c117 bl[117] br[117] wl[344] vdd gnd cell_6t
Xbit_r345_c117 bl[117] br[117] wl[345] vdd gnd cell_6t
Xbit_r346_c117 bl[117] br[117] wl[346] vdd gnd cell_6t
Xbit_r347_c117 bl[117] br[117] wl[347] vdd gnd cell_6t
Xbit_r348_c117 bl[117] br[117] wl[348] vdd gnd cell_6t
Xbit_r349_c117 bl[117] br[117] wl[349] vdd gnd cell_6t
Xbit_r350_c117 bl[117] br[117] wl[350] vdd gnd cell_6t
Xbit_r351_c117 bl[117] br[117] wl[351] vdd gnd cell_6t
Xbit_r352_c117 bl[117] br[117] wl[352] vdd gnd cell_6t
Xbit_r353_c117 bl[117] br[117] wl[353] vdd gnd cell_6t
Xbit_r354_c117 bl[117] br[117] wl[354] vdd gnd cell_6t
Xbit_r355_c117 bl[117] br[117] wl[355] vdd gnd cell_6t
Xbit_r356_c117 bl[117] br[117] wl[356] vdd gnd cell_6t
Xbit_r357_c117 bl[117] br[117] wl[357] vdd gnd cell_6t
Xbit_r358_c117 bl[117] br[117] wl[358] vdd gnd cell_6t
Xbit_r359_c117 bl[117] br[117] wl[359] vdd gnd cell_6t
Xbit_r360_c117 bl[117] br[117] wl[360] vdd gnd cell_6t
Xbit_r361_c117 bl[117] br[117] wl[361] vdd gnd cell_6t
Xbit_r362_c117 bl[117] br[117] wl[362] vdd gnd cell_6t
Xbit_r363_c117 bl[117] br[117] wl[363] vdd gnd cell_6t
Xbit_r364_c117 bl[117] br[117] wl[364] vdd gnd cell_6t
Xbit_r365_c117 bl[117] br[117] wl[365] vdd gnd cell_6t
Xbit_r366_c117 bl[117] br[117] wl[366] vdd gnd cell_6t
Xbit_r367_c117 bl[117] br[117] wl[367] vdd gnd cell_6t
Xbit_r368_c117 bl[117] br[117] wl[368] vdd gnd cell_6t
Xbit_r369_c117 bl[117] br[117] wl[369] vdd gnd cell_6t
Xbit_r370_c117 bl[117] br[117] wl[370] vdd gnd cell_6t
Xbit_r371_c117 bl[117] br[117] wl[371] vdd gnd cell_6t
Xbit_r372_c117 bl[117] br[117] wl[372] vdd gnd cell_6t
Xbit_r373_c117 bl[117] br[117] wl[373] vdd gnd cell_6t
Xbit_r374_c117 bl[117] br[117] wl[374] vdd gnd cell_6t
Xbit_r375_c117 bl[117] br[117] wl[375] vdd gnd cell_6t
Xbit_r376_c117 bl[117] br[117] wl[376] vdd gnd cell_6t
Xbit_r377_c117 bl[117] br[117] wl[377] vdd gnd cell_6t
Xbit_r378_c117 bl[117] br[117] wl[378] vdd gnd cell_6t
Xbit_r379_c117 bl[117] br[117] wl[379] vdd gnd cell_6t
Xbit_r380_c117 bl[117] br[117] wl[380] vdd gnd cell_6t
Xbit_r381_c117 bl[117] br[117] wl[381] vdd gnd cell_6t
Xbit_r382_c117 bl[117] br[117] wl[382] vdd gnd cell_6t
Xbit_r383_c117 bl[117] br[117] wl[383] vdd gnd cell_6t
Xbit_r384_c117 bl[117] br[117] wl[384] vdd gnd cell_6t
Xbit_r385_c117 bl[117] br[117] wl[385] vdd gnd cell_6t
Xbit_r386_c117 bl[117] br[117] wl[386] vdd gnd cell_6t
Xbit_r387_c117 bl[117] br[117] wl[387] vdd gnd cell_6t
Xbit_r388_c117 bl[117] br[117] wl[388] vdd gnd cell_6t
Xbit_r389_c117 bl[117] br[117] wl[389] vdd gnd cell_6t
Xbit_r390_c117 bl[117] br[117] wl[390] vdd gnd cell_6t
Xbit_r391_c117 bl[117] br[117] wl[391] vdd gnd cell_6t
Xbit_r392_c117 bl[117] br[117] wl[392] vdd gnd cell_6t
Xbit_r393_c117 bl[117] br[117] wl[393] vdd gnd cell_6t
Xbit_r394_c117 bl[117] br[117] wl[394] vdd gnd cell_6t
Xbit_r395_c117 bl[117] br[117] wl[395] vdd gnd cell_6t
Xbit_r396_c117 bl[117] br[117] wl[396] vdd gnd cell_6t
Xbit_r397_c117 bl[117] br[117] wl[397] vdd gnd cell_6t
Xbit_r398_c117 bl[117] br[117] wl[398] vdd gnd cell_6t
Xbit_r399_c117 bl[117] br[117] wl[399] vdd gnd cell_6t
Xbit_r400_c117 bl[117] br[117] wl[400] vdd gnd cell_6t
Xbit_r401_c117 bl[117] br[117] wl[401] vdd gnd cell_6t
Xbit_r402_c117 bl[117] br[117] wl[402] vdd gnd cell_6t
Xbit_r403_c117 bl[117] br[117] wl[403] vdd gnd cell_6t
Xbit_r404_c117 bl[117] br[117] wl[404] vdd gnd cell_6t
Xbit_r405_c117 bl[117] br[117] wl[405] vdd gnd cell_6t
Xbit_r406_c117 bl[117] br[117] wl[406] vdd gnd cell_6t
Xbit_r407_c117 bl[117] br[117] wl[407] vdd gnd cell_6t
Xbit_r408_c117 bl[117] br[117] wl[408] vdd gnd cell_6t
Xbit_r409_c117 bl[117] br[117] wl[409] vdd gnd cell_6t
Xbit_r410_c117 bl[117] br[117] wl[410] vdd gnd cell_6t
Xbit_r411_c117 bl[117] br[117] wl[411] vdd gnd cell_6t
Xbit_r412_c117 bl[117] br[117] wl[412] vdd gnd cell_6t
Xbit_r413_c117 bl[117] br[117] wl[413] vdd gnd cell_6t
Xbit_r414_c117 bl[117] br[117] wl[414] vdd gnd cell_6t
Xbit_r415_c117 bl[117] br[117] wl[415] vdd gnd cell_6t
Xbit_r416_c117 bl[117] br[117] wl[416] vdd gnd cell_6t
Xbit_r417_c117 bl[117] br[117] wl[417] vdd gnd cell_6t
Xbit_r418_c117 bl[117] br[117] wl[418] vdd gnd cell_6t
Xbit_r419_c117 bl[117] br[117] wl[419] vdd gnd cell_6t
Xbit_r420_c117 bl[117] br[117] wl[420] vdd gnd cell_6t
Xbit_r421_c117 bl[117] br[117] wl[421] vdd gnd cell_6t
Xbit_r422_c117 bl[117] br[117] wl[422] vdd gnd cell_6t
Xbit_r423_c117 bl[117] br[117] wl[423] vdd gnd cell_6t
Xbit_r424_c117 bl[117] br[117] wl[424] vdd gnd cell_6t
Xbit_r425_c117 bl[117] br[117] wl[425] vdd gnd cell_6t
Xbit_r426_c117 bl[117] br[117] wl[426] vdd gnd cell_6t
Xbit_r427_c117 bl[117] br[117] wl[427] vdd gnd cell_6t
Xbit_r428_c117 bl[117] br[117] wl[428] vdd gnd cell_6t
Xbit_r429_c117 bl[117] br[117] wl[429] vdd gnd cell_6t
Xbit_r430_c117 bl[117] br[117] wl[430] vdd gnd cell_6t
Xbit_r431_c117 bl[117] br[117] wl[431] vdd gnd cell_6t
Xbit_r432_c117 bl[117] br[117] wl[432] vdd gnd cell_6t
Xbit_r433_c117 bl[117] br[117] wl[433] vdd gnd cell_6t
Xbit_r434_c117 bl[117] br[117] wl[434] vdd gnd cell_6t
Xbit_r435_c117 bl[117] br[117] wl[435] vdd gnd cell_6t
Xbit_r436_c117 bl[117] br[117] wl[436] vdd gnd cell_6t
Xbit_r437_c117 bl[117] br[117] wl[437] vdd gnd cell_6t
Xbit_r438_c117 bl[117] br[117] wl[438] vdd gnd cell_6t
Xbit_r439_c117 bl[117] br[117] wl[439] vdd gnd cell_6t
Xbit_r440_c117 bl[117] br[117] wl[440] vdd gnd cell_6t
Xbit_r441_c117 bl[117] br[117] wl[441] vdd gnd cell_6t
Xbit_r442_c117 bl[117] br[117] wl[442] vdd gnd cell_6t
Xbit_r443_c117 bl[117] br[117] wl[443] vdd gnd cell_6t
Xbit_r444_c117 bl[117] br[117] wl[444] vdd gnd cell_6t
Xbit_r445_c117 bl[117] br[117] wl[445] vdd gnd cell_6t
Xbit_r446_c117 bl[117] br[117] wl[446] vdd gnd cell_6t
Xbit_r447_c117 bl[117] br[117] wl[447] vdd gnd cell_6t
Xbit_r448_c117 bl[117] br[117] wl[448] vdd gnd cell_6t
Xbit_r449_c117 bl[117] br[117] wl[449] vdd gnd cell_6t
Xbit_r450_c117 bl[117] br[117] wl[450] vdd gnd cell_6t
Xbit_r451_c117 bl[117] br[117] wl[451] vdd gnd cell_6t
Xbit_r452_c117 bl[117] br[117] wl[452] vdd gnd cell_6t
Xbit_r453_c117 bl[117] br[117] wl[453] vdd gnd cell_6t
Xbit_r454_c117 bl[117] br[117] wl[454] vdd gnd cell_6t
Xbit_r455_c117 bl[117] br[117] wl[455] vdd gnd cell_6t
Xbit_r456_c117 bl[117] br[117] wl[456] vdd gnd cell_6t
Xbit_r457_c117 bl[117] br[117] wl[457] vdd gnd cell_6t
Xbit_r458_c117 bl[117] br[117] wl[458] vdd gnd cell_6t
Xbit_r459_c117 bl[117] br[117] wl[459] vdd gnd cell_6t
Xbit_r460_c117 bl[117] br[117] wl[460] vdd gnd cell_6t
Xbit_r461_c117 bl[117] br[117] wl[461] vdd gnd cell_6t
Xbit_r462_c117 bl[117] br[117] wl[462] vdd gnd cell_6t
Xbit_r463_c117 bl[117] br[117] wl[463] vdd gnd cell_6t
Xbit_r464_c117 bl[117] br[117] wl[464] vdd gnd cell_6t
Xbit_r465_c117 bl[117] br[117] wl[465] vdd gnd cell_6t
Xbit_r466_c117 bl[117] br[117] wl[466] vdd gnd cell_6t
Xbit_r467_c117 bl[117] br[117] wl[467] vdd gnd cell_6t
Xbit_r468_c117 bl[117] br[117] wl[468] vdd gnd cell_6t
Xbit_r469_c117 bl[117] br[117] wl[469] vdd gnd cell_6t
Xbit_r470_c117 bl[117] br[117] wl[470] vdd gnd cell_6t
Xbit_r471_c117 bl[117] br[117] wl[471] vdd gnd cell_6t
Xbit_r472_c117 bl[117] br[117] wl[472] vdd gnd cell_6t
Xbit_r473_c117 bl[117] br[117] wl[473] vdd gnd cell_6t
Xbit_r474_c117 bl[117] br[117] wl[474] vdd gnd cell_6t
Xbit_r475_c117 bl[117] br[117] wl[475] vdd gnd cell_6t
Xbit_r476_c117 bl[117] br[117] wl[476] vdd gnd cell_6t
Xbit_r477_c117 bl[117] br[117] wl[477] vdd gnd cell_6t
Xbit_r478_c117 bl[117] br[117] wl[478] vdd gnd cell_6t
Xbit_r479_c117 bl[117] br[117] wl[479] vdd gnd cell_6t
Xbit_r480_c117 bl[117] br[117] wl[480] vdd gnd cell_6t
Xbit_r481_c117 bl[117] br[117] wl[481] vdd gnd cell_6t
Xbit_r482_c117 bl[117] br[117] wl[482] vdd gnd cell_6t
Xbit_r483_c117 bl[117] br[117] wl[483] vdd gnd cell_6t
Xbit_r484_c117 bl[117] br[117] wl[484] vdd gnd cell_6t
Xbit_r485_c117 bl[117] br[117] wl[485] vdd gnd cell_6t
Xbit_r486_c117 bl[117] br[117] wl[486] vdd gnd cell_6t
Xbit_r487_c117 bl[117] br[117] wl[487] vdd gnd cell_6t
Xbit_r488_c117 bl[117] br[117] wl[488] vdd gnd cell_6t
Xbit_r489_c117 bl[117] br[117] wl[489] vdd gnd cell_6t
Xbit_r490_c117 bl[117] br[117] wl[490] vdd gnd cell_6t
Xbit_r491_c117 bl[117] br[117] wl[491] vdd gnd cell_6t
Xbit_r492_c117 bl[117] br[117] wl[492] vdd gnd cell_6t
Xbit_r493_c117 bl[117] br[117] wl[493] vdd gnd cell_6t
Xbit_r494_c117 bl[117] br[117] wl[494] vdd gnd cell_6t
Xbit_r495_c117 bl[117] br[117] wl[495] vdd gnd cell_6t
Xbit_r496_c117 bl[117] br[117] wl[496] vdd gnd cell_6t
Xbit_r497_c117 bl[117] br[117] wl[497] vdd gnd cell_6t
Xbit_r498_c117 bl[117] br[117] wl[498] vdd gnd cell_6t
Xbit_r499_c117 bl[117] br[117] wl[499] vdd gnd cell_6t
Xbit_r500_c117 bl[117] br[117] wl[500] vdd gnd cell_6t
Xbit_r501_c117 bl[117] br[117] wl[501] vdd gnd cell_6t
Xbit_r502_c117 bl[117] br[117] wl[502] vdd gnd cell_6t
Xbit_r503_c117 bl[117] br[117] wl[503] vdd gnd cell_6t
Xbit_r504_c117 bl[117] br[117] wl[504] vdd gnd cell_6t
Xbit_r505_c117 bl[117] br[117] wl[505] vdd gnd cell_6t
Xbit_r506_c117 bl[117] br[117] wl[506] vdd gnd cell_6t
Xbit_r507_c117 bl[117] br[117] wl[507] vdd gnd cell_6t
Xbit_r508_c117 bl[117] br[117] wl[508] vdd gnd cell_6t
Xbit_r509_c117 bl[117] br[117] wl[509] vdd gnd cell_6t
Xbit_r510_c117 bl[117] br[117] wl[510] vdd gnd cell_6t
Xbit_r511_c117 bl[117] br[117] wl[511] vdd gnd cell_6t
Xbit_r0_c118 bl[118] br[118] wl[0] vdd gnd cell_6t
Xbit_r1_c118 bl[118] br[118] wl[1] vdd gnd cell_6t
Xbit_r2_c118 bl[118] br[118] wl[2] vdd gnd cell_6t
Xbit_r3_c118 bl[118] br[118] wl[3] vdd gnd cell_6t
Xbit_r4_c118 bl[118] br[118] wl[4] vdd gnd cell_6t
Xbit_r5_c118 bl[118] br[118] wl[5] vdd gnd cell_6t
Xbit_r6_c118 bl[118] br[118] wl[6] vdd gnd cell_6t
Xbit_r7_c118 bl[118] br[118] wl[7] vdd gnd cell_6t
Xbit_r8_c118 bl[118] br[118] wl[8] vdd gnd cell_6t
Xbit_r9_c118 bl[118] br[118] wl[9] vdd gnd cell_6t
Xbit_r10_c118 bl[118] br[118] wl[10] vdd gnd cell_6t
Xbit_r11_c118 bl[118] br[118] wl[11] vdd gnd cell_6t
Xbit_r12_c118 bl[118] br[118] wl[12] vdd gnd cell_6t
Xbit_r13_c118 bl[118] br[118] wl[13] vdd gnd cell_6t
Xbit_r14_c118 bl[118] br[118] wl[14] vdd gnd cell_6t
Xbit_r15_c118 bl[118] br[118] wl[15] vdd gnd cell_6t
Xbit_r16_c118 bl[118] br[118] wl[16] vdd gnd cell_6t
Xbit_r17_c118 bl[118] br[118] wl[17] vdd gnd cell_6t
Xbit_r18_c118 bl[118] br[118] wl[18] vdd gnd cell_6t
Xbit_r19_c118 bl[118] br[118] wl[19] vdd gnd cell_6t
Xbit_r20_c118 bl[118] br[118] wl[20] vdd gnd cell_6t
Xbit_r21_c118 bl[118] br[118] wl[21] vdd gnd cell_6t
Xbit_r22_c118 bl[118] br[118] wl[22] vdd gnd cell_6t
Xbit_r23_c118 bl[118] br[118] wl[23] vdd gnd cell_6t
Xbit_r24_c118 bl[118] br[118] wl[24] vdd gnd cell_6t
Xbit_r25_c118 bl[118] br[118] wl[25] vdd gnd cell_6t
Xbit_r26_c118 bl[118] br[118] wl[26] vdd gnd cell_6t
Xbit_r27_c118 bl[118] br[118] wl[27] vdd gnd cell_6t
Xbit_r28_c118 bl[118] br[118] wl[28] vdd gnd cell_6t
Xbit_r29_c118 bl[118] br[118] wl[29] vdd gnd cell_6t
Xbit_r30_c118 bl[118] br[118] wl[30] vdd gnd cell_6t
Xbit_r31_c118 bl[118] br[118] wl[31] vdd gnd cell_6t
Xbit_r32_c118 bl[118] br[118] wl[32] vdd gnd cell_6t
Xbit_r33_c118 bl[118] br[118] wl[33] vdd gnd cell_6t
Xbit_r34_c118 bl[118] br[118] wl[34] vdd gnd cell_6t
Xbit_r35_c118 bl[118] br[118] wl[35] vdd gnd cell_6t
Xbit_r36_c118 bl[118] br[118] wl[36] vdd gnd cell_6t
Xbit_r37_c118 bl[118] br[118] wl[37] vdd gnd cell_6t
Xbit_r38_c118 bl[118] br[118] wl[38] vdd gnd cell_6t
Xbit_r39_c118 bl[118] br[118] wl[39] vdd gnd cell_6t
Xbit_r40_c118 bl[118] br[118] wl[40] vdd gnd cell_6t
Xbit_r41_c118 bl[118] br[118] wl[41] vdd gnd cell_6t
Xbit_r42_c118 bl[118] br[118] wl[42] vdd gnd cell_6t
Xbit_r43_c118 bl[118] br[118] wl[43] vdd gnd cell_6t
Xbit_r44_c118 bl[118] br[118] wl[44] vdd gnd cell_6t
Xbit_r45_c118 bl[118] br[118] wl[45] vdd gnd cell_6t
Xbit_r46_c118 bl[118] br[118] wl[46] vdd gnd cell_6t
Xbit_r47_c118 bl[118] br[118] wl[47] vdd gnd cell_6t
Xbit_r48_c118 bl[118] br[118] wl[48] vdd gnd cell_6t
Xbit_r49_c118 bl[118] br[118] wl[49] vdd gnd cell_6t
Xbit_r50_c118 bl[118] br[118] wl[50] vdd gnd cell_6t
Xbit_r51_c118 bl[118] br[118] wl[51] vdd gnd cell_6t
Xbit_r52_c118 bl[118] br[118] wl[52] vdd gnd cell_6t
Xbit_r53_c118 bl[118] br[118] wl[53] vdd gnd cell_6t
Xbit_r54_c118 bl[118] br[118] wl[54] vdd gnd cell_6t
Xbit_r55_c118 bl[118] br[118] wl[55] vdd gnd cell_6t
Xbit_r56_c118 bl[118] br[118] wl[56] vdd gnd cell_6t
Xbit_r57_c118 bl[118] br[118] wl[57] vdd gnd cell_6t
Xbit_r58_c118 bl[118] br[118] wl[58] vdd gnd cell_6t
Xbit_r59_c118 bl[118] br[118] wl[59] vdd gnd cell_6t
Xbit_r60_c118 bl[118] br[118] wl[60] vdd gnd cell_6t
Xbit_r61_c118 bl[118] br[118] wl[61] vdd gnd cell_6t
Xbit_r62_c118 bl[118] br[118] wl[62] vdd gnd cell_6t
Xbit_r63_c118 bl[118] br[118] wl[63] vdd gnd cell_6t
Xbit_r64_c118 bl[118] br[118] wl[64] vdd gnd cell_6t
Xbit_r65_c118 bl[118] br[118] wl[65] vdd gnd cell_6t
Xbit_r66_c118 bl[118] br[118] wl[66] vdd gnd cell_6t
Xbit_r67_c118 bl[118] br[118] wl[67] vdd gnd cell_6t
Xbit_r68_c118 bl[118] br[118] wl[68] vdd gnd cell_6t
Xbit_r69_c118 bl[118] br[118] wl[69] vdd gnd cell_6t
Xbit_r70_c118 bl[118] br[118] wl[70] vdd gnd cell_6t
Xbit_r71_c118 bl[118] br[118] wl[71] vdd gnd cell_6t
Xbit_r72_c118 bl[118] br[118] wl[72] vdd gnd cell_6t
Xbit_r73_c118 bl[118] br[118] wl[73] vdd gnd cell_6t
Xbit_r74_c118 bl[118] br[118] wl[74] vdd gnd cell_6t
Xbit_r75_c118 bl[118] br[118] wl[75] vdd gnd cell_6t
Xbit_r76_c118 bl[118] br[118] wl[76] vdd gnd cell_6t
Xbit_r77_c118 bl[118] br[118] wl[77] vdd gnd cell_6t
Xbit_r78_c118 bl[118] br[118] wl[78] vdd gnd cell_6t
Xbit_r79_c118 bl[118] br[118] wl[79] vdd gnd cell_6t
Xbit_r80_c118 bl[118] br[118] wl[80] vdd gnd cell_6t
Xbit_r81_c118 bl[118] br[118] wl[81] vdd gnd cell_6t
Xbit_r82_c118 bl[118] br[118] wl[82] vdd gnd cell_6t
Xbit_r83_c118 bl[118] br[118] wl[83] vdd gnd cell_6t
Xbit_r84_c118 bl[118] br[118] wl[84] vdd gnd cell_6t
Xbit_r85_c118 bl[118] br[118] wl[85] vdd gnd cell_6t
Xbit_r86_c118 bl[118] br[118] wl[86] vdd gnd cell_6t
Xbit_r87_c118 bl[118] br[118] wl[87] vdd gnd cell_6t
Xbit_r88_c118 bl[118] br[118] wl[88] vdd gnd cell_6t
Xbit_r89_c118 bl[118] br[118] wl[89] vdd gnd cell_6t
Xbit_r90_c118 bl[118] br[118] wl[90] vdd gnd cell_6t
Xbit_r91_c118 bl[118] br[118] wl[91] vdd gnd cell_6t
Xbit_r92_c118 bl[118] br[118] wl[92] vdd gnd cell_6t
Xbit_r93_c118 bl[118] br[118] wl[93] vdd gnd cell_6t
Xbit_r94_c118 bl[118] br[118] wl[94] vdd gnd cell_6t
Xbit_r95_c118 bl[118] br[118] wl[95] vdd gnd cell_6t
Xbit_r96_c118 bl[118] br[118] wl[96] vdd gnd cell_6t
Xbit_r97_c118 bl[118] br[118] wl[97] vdd gnd cell_6t
Xbit_r98_c118 bl[118] br[118] wl[98] vdd gnd cell_6t
Xbit_r99_c118 bl[118] br[118] wl[99] vdd gnd cell_6t
Xbit_r100_c118 bl[118] br[118] wl[100] vdd gnd cell_6t
Xbit_r101_c118 bl[118] br[118] wl[101] vdd gnd cell_6t
Xbit_r102_c118 bl[118] br[118] wl[102] vdd gnd cell_6t
Xbit_r103_c118 bl[118] br[118] wl[103] vdd gnd cell_6t
Xbit_r104_c118 bl[118] br[118] wl[104] vdd gnd cell_6t
Xbit_r105_c118 bl[118] br[118] wl[105] vdd gnd cell_6t
Xbit_r106_c118 bl[118] br[118] wl[106] vdd gnd cell_6t
Xbit_r107_c118 bl[118] br[118] wl[107] vdd gnd cell_6t
Xbit_r108_c118 bl[118] br[118] wl[108] vdd gnd cell_6t
Xbit_r109_c118 bl[118] br[118] wl[109] vdd gnd cell_6t
Xbit_r110_c118 bl[118] br[118] wl[110] vdd gnd cell_6t
Xbit_r111_c118 bl[118] br[118] wl[111] vdd gnd cell_6t
Xbit_r112_c118 bl[118] br[118] wl[112] vdd gnd cell_6t
Xbit_r113_c118 bl[118] br[118] wl[113] vdd gnd cell_6t
Xbit_r114_c118 bl[118] br[118] wl[114] vdd gnd cell_6t
Xbit_r115_c118 bl[118] br[118] wl[115] vdd gnd cell_6t
Xbit_r116_c118 bl[118] br[118] wl[116] vdd gnd cell_6t
Xbit_r117_c118 bl[118] br[118] wl[117] vdd gnd cell_6t
Xbit_r118_c118 bl[118] br[118] wl[118] vdd gnd cell_6t
Xbit_r119_c118 bl[118] br[118] wl[119] vdd gnd cell_6t
Xbit_r120_c118 bl[118] br[118] wl[120] vdd gnd cell_6t
Xbit_r121_c118 bl[118] br[118] wl[121] vdd gnd cell_6t
Xbit_r122_c118 bl[118] br[118] wl[122] vdd gnd cell_6t
Xbit_r123_c118 bl[118] br[118] wl[123] vdd gnd cell_6t
Xbit_r124_c118 bl[118] br[118] wl[124] vdd gnd cell_6t
Xbit_r125_c118 bl[118] br[118] wl[125] vdd gnd cell_6t
Xbit_r126_c118 bl[118] br[118] wl[126] vdd gnd cell_6t
Xbit_r127_c118 bl[118] br[118] wl[127] vdd gnd cell_6t
Xbit_r128_c118 bl[118] br[118] wl[128] vdd gnd cell_6t
Xbit_r129_c118 bl[118] br[118] wl[129] vdd gnd cell_6t
Xbit_r130_c118 bl[118] br[118] wl[130] vdd gnd cell_6t
Xbit_r131_c118 bl[118] br[118] wl[131] vdd gnd cell_6t
Xbit_r132_c118 bl[118] br[118] wl[132] vdd gnd cell_6t
Xbit_r133_c118 bl[118] br[118] wl[133] vdd gnd cell_6t
Xbit_r134_c118 bl[118] br[118] wl[134] vdd gnd cell_6t
Xbit_r135_c118 bl[118] br[118] wl[135] vdd gnd cell_6t
Xbit_r136_c118 bl[118] br[118] wl[136] vdd gnd cell_6t
Xbit_r137_c118 bl[118] br[118] wl[137] vdd gnd cell_6t
Xbit_r138_c118 bl[118] br[118] wl[138] vdd gnd cell_6t
Xbit_r139_c118 bl[118] br[118] wl[139] vdd gnd cell_6t
Xbit_r140_c118 bl[118] br[118] wl[140] vdd gnd cell_6t
Xbit_r141_c118 bl[118] br[118] wl[141] vdd gnd cell_6t
Xbit_r142_c118 bl[118] br[118] wl[142] vdd gnd cell_6t
Xbit_r143_c118 bl[118] br[118] wl[143] vdd gnd cell_6t
Xbit_r144_c118 bl[118] br[118] wl[144] vdd gnd cell_6t
Xbit_r145_c118 bl[118] br[118] wl[145] vdd gnd cell_6t
Xbit_r146_c118 bl[118] br[118] wl[146] vdd gnd cell_6t
Xbit_r147_c118 bl[118] br[118] wl[147] vdd gnd cell_6t
Xbit_r148_c118 bl[118] br[118] wl[148] vdd gnd cell_6t
Xbit_r149_c118 bl[118] br[118] wl[149] vdd gnd cell_6t
Xbit_r150_c118 bl[118] br[118] wl[150] vdd gnd cell_6t
Xbit_r151_c118 bl[118] br[118] wl[151] vdd gnd cell_6t
Xbit_r152_c118 bl[118] br[118] wl[152] vdd gnd cell_6t
Xbit_r153_c118 bl[118] br[118] wl[153] vdd gnd cell_6t
Xbit_r154_c118 bl[118] br[118] wl[154] vdd gnd cell_6t
Xbit_r155_c118 bl[118] br[118] wl[155] vdd gnd cell_6t
Xbit_r156_c118 bl[118] br[118] wl[156] vdd gnd cell_6t
Xbit_r157_c118 bl[118] br[118] wl[157] vdd gnd cell_6t
Xbit_r158_c118 bl[118] br[118] wl[158] vdd gnd cell_6t
Xbit_r159_c118 bl[118] br[118] wl[159] vdd gnd cell_6t
Xbit_r160_c118 bl[118] br[118] wl[160] vdd gnd cell_6t
Xbit_r161_c118 bl[118] br[118] wl[161] vdd gnd cell_6t
Xbit_r162_c118 bl[118] br[118] wl[162] vdd gnd cell_6t
Xbit_r163_c118 bl[118] br[118] wl[163] vdd gnd cell_6t
Xbit_r164_c118 bl[118] br[118] wl[164] vdd gnd cell_6t
Xbit_r165_c118 bl[118] br[118] wl[165] vdd gnd cell_6t
Xbit_r166_c118 bl[118] br[118] wl[166] vdd gnd cell_6t
Xbit_r167_c118 bl[118] br[118] wl[167] vdd gnd cell_6t
Xbit_r168_c118 bl[118] br[118] wl[168] vdd gnd cell_6t
Xbit_r169_c118 bl[118] br[118] wl[169] vdd gnd cell_6t
Xbit_r170_c118 bl[118] br[118] wl[170] vdd gnd cell_6t
Xbit_r171_c118 bl[118] br[118] wl[171] vdd gnd cell_6t
Xbit_r172_c118 bl[118] br[118] wl[172] vdd gnd cell_6t
Xbit_r173_c118 bl[118] br[118] wl[173] vdd gnd cell_6t
Xbit_r174_c118 bl[118] br[118] wl[174] vdd gnd cell_6t
Xbit_r175_c118 bl[118] br[118] wl[175] vdd gnd cell_6t
Xbit_r176_c118 bl[118] br[118] wl[176] vdd gnd cell_6t
Xbit_r177_c118 bl[118] br[118] wl[177] vdd gnd cell_6t
Xbit_r178_c118 bl[118] br[118] wl[178] vdd gnd cell_6t
Xbit_r179_c118 bl[118] br[118] wl[179] vdd gnd cell_6t
Xbit_r180_c118 bl[118] br[118] wl[180] vdd gnd cell_6t
Xbit_r181_c118 bl[118] br[118] wl[181] vdd gnd cell_6t
Xbit_r182_c118 bl[118] br[118] wl[182] vdd gnd cell_6t
Xbit_r183_c118 bl[118] br[118] wl[183] vdd gnd cell_6t
Xbit_r184_c118 bl[118] br[118] wl[184] vdd gnd cell_6t
Xbit_r185_c118 bl[118] br[118] wl[185] vdd gnd cell_6t
Xbit_r186_c118 bl[118] br[118] wl[186] vdd gnd cell_6t
Xbit_r187_c118 bl[118] br[118] wl[187] vdd gnd cell_6t
Xbit_r188_c118 bl[118] br[118] wl[188] vdd gnd cell_6t
Xbit_r189_c118 bl[118] br[118] wl[189] vdd gnd cell_6t
Xbit_r190_c118 bl[118] br[118] wl[190] vdd gnd cell_6t
Xbit_r191_c118 bl[118] br[118] wl[191] vdd gnd cell_6t
Xbit_r192_c118 bl[118] br[118] wl[192] vdd gnd cell_6t
Xbit_r193_c118 bl[118] br[118] wl[193] vdd gnd cell_6t
Xbit_r194_c118 bl[118] br[118] wl[194] vdd gnd cell_6t
Xbit_r195_c118 bl[118] br[118] wl[195] vdd gnd cell_6t
Xbit_r196_c118 bl[118] br[118] wl[196] vdd gnd cell_6t
Xbit_r197_c118 bl[118] br[118] wl[197] vdd gnd cell_6t
Xbit_r198_c118 bl[118] br[118] wl[198] vdd gnd cell_6t
Xbit_r199_c118 bl[118] br[118] wl[199] vdd gnd cell_6t
Xbit_r200_c118 bl[118] br[118] wl[200] vdd gnd cell_6t
Xbit_r201_c118 bl[118] br[118] wl[201] vdd gnd cell_6t
Xbit_r202_c118 bl[118] br[118] wl[202] vdd gnd cell_6t
Xbit_r203_c118 bl[118] br[118] wl[203] vdd gnd cell_6t
Xbit_r204_c118 bl[118] br[118] wl[204] vdd gnd cell_6t
Xbit_r205_c118 bl[118] br[118] wl[205] vdd gnd cell_6t
Xbit_r206_c118 bl[118] br[118] wl[206] vdd gnd cell_6t
Xbit_r207_c118 bl[118] br[118] wl[207] vdd gnd cell_6t
Xbit_r208_c118 bl[118] br[118] wl[208] vdd gnd cell_6t
Xbit_r209_c118 bl[118] br[118] wl[209] vdd gnd cell_6t
Xbit_r210_c118 bl[118] br[118] wl[210] vdd gnd cell_6t
Xbit_r211_c118 bl[118] br[118] wl[211] vdd gnd cell_6t
Xbit_r212_c118 bl[118] br[118] wl[212] vdd gnd cell_6t
Xbit_r213_c118 bl[118] br[118] wl[213] vdd gnd cell_6t
Xbit_r214_c118 bl[118] br[118] wl[214] vdd gnd cell_6t
Xbit_r215_c118 bl[118] br[118] wl[215] vdd gnd cell_6t
Xbit_r216_c118 bl[118] br[118] wl[216] vdd gnd cell_6t
Xbit_r217_c118 bl[118] br[118] wl[217] vdd gnd cell_6t
Xbit_r218_c118 bl[118] br[118] wl[218] vdd gnd cell_6t
Xbit_r219_c118 bl[118] br[118] wl[219] vdd gnd cell_6t
Xbit_r220_c118 bl[118] br[118] wl[220] vdd gnd cell_6t
Xbit_r221_c118 bl[118] br[118] wl[221] vdd gnd cell_6t
Xbit_r222_c118 bl[118] br[118] wl[222] vdd gnd cell_6t
Xbit_r223_c118 bl[118] br[118] wl[223] vdd gnd cell_6t
Xbit_r224_c118 bl[118] br[118] wl[224] vdd gnd cell_6t
Xbit_r225_c118 bl[118] br[118] wl[225] vdd gnd cell_6t
Xbit_r226_c118 bl[118] br[118] wl[226] vdd gnd cell_6t
Xbit_r227_c118 bl[118] br[118] wl[227] vdd gnd cell_6t
Xbit_r228_c118 bl[118] br[118] wl[228] vdd gnd cell_6t
Xbit_r229_c118 bl[118] br[118] wl[229] vdd gnd cell_6t
Xbit_r230_c118 bl[118] br[118] wl[230] vdd gnd cell_6t
Xbit_r231_c118 bl[118] br[118] wl[231] vdd gnd cell_6t
Xbit_r232_c118 bl[118] br[118] wl[232] vdd gnd cell_6t
Xbit_r233_c118 bl[118] br[118] wl[233] vdd gnd cell_6t
Xbit_r234_c118 bl[118] br[118] wl[234] vdd gnd cell_6t
Xbit_r235_c118 bl[118] br[118] wl[235] vdd gnd cell_6t
Xbit_r236_c118 bl[118] br[118] wl[236] vdd gnd cell_6t
Xbit_r237_c118 bl[118] br[118] wl[237] vdd gnd cell_6t
Xbit_r238_c118 bl[118] br[118] wl[238] vdd gnd cell_6t
Xbit_r239_c118 bl[118] br[118] wl[239] vdd gnd cell_6t
Xbit_r240_c118 bl[118] br[118] wl[240] vdd gnd cell_6t
Xbit_r241_c118 bl[118] br[118] wl[241] vdd gnd cell_6t
Xbit_r242_c118 bl[118] br[118] wl[242] vdd gnd cell_6t
Xbit_r243_c118 bl[118] br[118] wl[243] vdd gnd cell_6t
Xbit_r244_c118 bl[118] br[118] wl[244] vdd gnd cell_6t
Xbit_r245_c118 bl[118] br[118] wl[245] vdd gnd cell_6t
Xbit_r246_c118 bl[118] br[118] wl[246] vdd gnd cell_6t
Xbit_r247_c118 bl[118] br[118] wl[247] vdd gnd cell_6t
Xbit_r248_c118 bl[118] br[118] wl[248] vdd gnd cell_6t
Xbit_r249_c118 bl[118] br[118] wl[249] vdd gnd cell_6t
Xbit_r250_c118 bl[118] br[118] wl[250] vdd gnd cell_6t
Xbit_r251_c118 bl[118] br[118] wl[251] vdd gnd cell_6t
Xbit_r252_c118 bl[118] br[118] wl[252] vdd gnd cell_6t
Xbit_r253_c118 bl[118] br[118] wl[253] vdd gnd cell_6t
Xbit_r254_c118 bl[118] br[118] wl[254] vdd gnd cell_6t
Xbit_r255_c118 bl[118] br[118] wl[255] vdd gnd cell_6t
Xbit_r256_c118 bl[118] br[118] wl[256] vdd gnd cell_6t
Xbit_r257_c118 bl[118] br[118] wl[257] vdd gnd cell_6t
Xbit_r258_c118 bl[118] br[118] wl[258] vdd gnd cell_6t
Xbit_r259_c118 bl[118] br[118] wl[259] vdd gnd cell_6t
Xbit_r260_c118 bl[118] br[118] wl[260] vdd gnd cell_6t
Xbit_r261_c118 bl[118] br[118] wl[261] vdd gnd cell_6t
Xbit_r262_c118 bl[118] br[118] wl[262] vdd gnd cell_6t
Xbit_r263_c118 bl[118] br[118] wl[263] vdd gnd cell_6t
Xbit_r264_c118 bl[118] br[118] wl[264] vdd gnd cell_6t
Xbit_r265_c118 bl[118] br[118] wl[265] vdd gnd cell_6t
Xbit_r266_c118 bl[118] br[118] wl[266] vdd gnd cell_6t
Xbit_r267_c118 bl[118] br[118] wl[267] vdd gnd cell_6t
Xbit_r268_c118 bl[118] br[118] wl[268] vdd gnd cell_6t
Xbit_r269_c118 bl[118] br[118] wl[269] vdd gnd cell_6t
Xbit_r270_c118 bl[118] br[118] wl[270] vdd gnd cell_6t
Xbit_r271_c118 bl[118] br[118] wl[271] vdd gnd cell_6t
Xbit_r272_c118 bl[118] br[118] wl[272] vdd gnd cell_6t
Xbit_r273_c118 bl[118] br[118] wl[273] vdd gnd cell_6t
Xbit_r274_c118 bl[118] br[118] wl[274] vdd gnd cell_6t
Xbit_r275_c118 bl[118] br[118] wl[275] vdd gnd cell_6t
Xbit_r276_c118 bl[118] br[118] wl[276] vdd gnd cell_6t
Xbit_r277_c118 bl[118] br[118] wl[277] vdd gnd cell_6t
Xbit_r278_c118 bl[118] br[118] wl[278] vdd gnd cell_6t
Xbit_r279_c118 bl[118] br[118] wl[279] vdd gnd cell_6t
Xbit_r280_c118 bl[118] br[118] wl[280] vdd gnd cell_6t
Xbit_r281_c118 bl[118] br[118] wl[281] vdd gnd cell_6t
Xbit_r282_c118 bl[118] br[118] wl[282] vdd gnd cell_6t
Xbit_r283_c118 bl[118] br[118] wl[283] vdd gnd cell_6t
Xbit_r284_c118 bl[118] br[118] wl[284] vdd gnd cell_6t
Xbit_r285_c118 bl[118] br[118] wl[285] vdd gnd cell_6t
Xbit_r286_c118 bl[118] br[118] wl[286] vdd gnd cell_6t
Xbit_r287_c118 bl[118] br[118] wl[287] vdd gnd cell_6t
Xbit_r288_c118 bl[118] br[118] wl[288] vdd gnd cell_6t
Xbit_r289_c118 bl[118] br[118] wl[289] vdd gnd cell_6t
Xbit_r290_c118 bl[118] br[118] wl[290] vdd gnd cell_6t
Xbit_r291_c118 bl[118] br[118] wl[291] vdd gnd cell_6t
Xbit_r292_c118 bl[118] br[118] wl[292] vdd gnd cell_6t
Xbit_r293_c118 bl[118] br[118] wl[293] vdd gnd cell_6t
Xbit_r294_c118 bl[118] br[118] wl[294] vdd gnd cell_6t
Xbit_r295_c118 bl[118] br[118] wl[295] vdd gnd cell_6t
Xbit_r296_c118 bl[118] br[118] wl[296] vdd gnd cell_6t
Xbit_r297_c118 bl[118] br[118] wl[297] vdd gnd cell_6t
Xbit_r298_c118 bl[118] br[118] wl[298] vdd gnd cell_6t
Xbit_r299_c118 bl[118] br[118] wl[299] vdd gnd cell_6t
Xbit_r300_c118 bl[118] br[118] wl[300] vdd gnd cell_6t
Xbit_r301_c118 bl[118] br[118] wl[301] vdd gnd cell_6t
Xbit_r302_c118 bl[118] br[118] wl[302] vdd gnd cell_6t
Xbit_r303_c118 bl[118] br[118] wl[303] vdd gnd cell_6t
Xbit_r304_c118 bl[118] br[118] wl[304] vdd gnd cell_6t
Xbit_r305_c118 bl[118] br[118] wl[305] vdd gnd cell_6t
Xbit_r306_c118 bl[118] br[118] wl[306] vdd gnd cell_6t
Xbit_r307_c118 bl[118] br[118] wl[307] vdd gnd cell_6t
Xbit_r308_c118 bl[118] br[118] wl[308] vdd gnd cell_6t
Xbit_r309_c118 bl[118] br[118] wl[309] vdd gnd cell_6t
Xbit_r310_c118 bl[118] br[118] wl[310] vdd gnd cell_6t
Xbit_r311_c118 bl[118] br[118] wl[311] vdd gnd cell_6t
Xbit_r312_c118 bl[118] br[118] wl[312] vdd gnd cell_6t
Xbit_r313_c118 bl[118] br[118] wl[313] vdd gnd cell_6t
Xbit_r314_c118 bl[118] br[118] wl[314] vdd gnd cell_6t
Xbit_r315_c118 bl[118] br[118] wl[315] vdd gnd cell_6t
Xbit_r316_c118 bl[118] br[118] wl[316] vdd gnd cell_6t
Xbit_r317_c118 bl[118] br[118] wl[317] vdd gnd cell_6t
Xbit_r318_c118 bl[118] br[118] wl[318] vdd gnd cell_6t
Xbit_r319_c118 bl[118] br[118] wl[319] vdd gnd cell_6t
Xbit_r320_c118 bl[118] br[118] wl[320] vdd gnd cell_6t
Xbit_r321_c118 bl[118] br[118] wl[321] vdd gnd cell_6t
Xbit_r322_c118 bl[118] br[118] wl[322] vdd gnd cell_6t
Xbit_r323_c118 bl[118] br[118] wl[323] vdd gnd cell_6t
Xbit_r324_c118 bl[118] br[118] wl[324] vdd gnd cell_6t
Xbit_r325_c118 bl[118] br[118] wl[325] vdd gnd cell_6t
Xbit_r326_c118 bl[118] br[118] wl[326] vdd gnd cell_6t
Xbit_r327_c118 bl[118] br[118] wl[327] vdd gnd cell_6t
Xbit_r328_c118 bl[118] br[118] wl[328] vdd gnd cell_6t
Xbit_r329_c118 bl[118] br[118] wl[329] vdd gnd cell_6t
Xbit_r330_c118 bl[118] br[118] wl[330] vdd gnd cell_6t
Xbit_r331_c118 bl[118] br[118] wl[331] vdd gnd cell_6t
Xbit_r332_c118 bl[118] br[118] wl[332] vdd gnd cell_6t
Xbit_r333_c118 bl[118] br[118] wl[333] vdd gnd cell_6t
Xbit_r334_c118 bl[118] br[118] wl[334] vdd gnd cell_6t
Xbit_r335_c118 bl[118] br[118] wl[335] vdd gnd cell_6t
Xbit_r336_c118 bl[118] br[118] wl[336] vdd gnd cell_6t
Xbit_r337_c118 bl[118] br[118] wl[337] vdd gnd cell_6t
Xbit_r338_c118 bl[118] br[118] wl[338] vdd gnd cell_6t
Xbit_r339_c118 bl[118] br[118] wl[339] vdd gnd cell_6t
Xbit_r340_c118 bl[118] br[118] wl[340] vdd gnd cell_6t
Xbit_r341_c118 bl[118] br[118] wl[341] vdd gnd cell_6t
Xbit_r342_c118 bl[118] br[118] wl[342] vdd gnd cell_6t
Xbit_r343_c118 bl[118] br[118] wl[343] vdd gnd cell_6t
Xbit_r344_c118 bl[118] br[118] wl[344] vdd gnd cell_6t
Xbit_r345_c118 bl[118] br[118] wl[345] vdd gnd cell_6t
Xbit_r346_c118 bl[118] br[118] wl[346] vdd gnd cell_6t
Xbit_r347_c118 bl[118] br[118] wl[347] vdd gnd cell_6t
Xbit_r348_c118 bl[118] br[118] wl[348] vdd gnd cell_6t
Xbit_r349_c118 bl[118] br[118] wl[349] vdd gnd cell_6t
Xbit_r350_c118 bl[118] br[118] wl[350] vdd gnd cell_6t
Xbit_r351_c118 bl[118] br[118] wl[351] vdd gnd cell_6t
Xbit_r352_c118 bl[118] br[118] wl[352] vdd gnd cell_6t
Xbit_r353_c118 bl[118] br[118] wl[353] vdd gnd cell_6t
Xbit_r354_c118 bl[118] br[118] wl[354] vdd gnd cell_6t
Xbit_r355_c118 bl[118] br[118] wl[355] vdd gnd cell_6t
Xbit_r356_c118 bl[118] br[118] wl[356] vdd gnd cell_6t
Xbit_r357_c118 bl[118] br[118] wl[357] vdd gnd cell_6t
Xbit_r358_c118 bl[118] br[118] wl[358] vdd gnd cell_6t
Xbit_r359_c118 bl[118] br[118] wl[359] vdd gnd cell_6t
Xbit_r360_c118 bl[118] br[118] wl[360] vdd gnd cell_6t
Xbit_r361_c118 bl[118] br[118] wl[361] vdd gnd cell_6t
Xbit_r362_c118 bl[118] br[118] wl[362] vdd gnd cell_6t
Xbit_r363_c118 bl[118] br[118] wl[363] vdd gnd cell_6t
Xbit_r364_c118 bl[118] br[118] wl[364] vdd gnd cell_6t
Xbit_r365_c118 bl[118] br[118] wl[365] vdd gnd cell_6t
Xbit_r366_c118 bl[118] br[118] wl[366] vdd gnd cell_6t
Xbit_r367_c118 bl[118] br[118] wl[367] vdd gnd cell_6t
Xbit_r368_c118 bl[118] br[118] wl[368] vdd gnd cell_6t
Xbit_r369_c118 bl[118] br[118] wl[369] vdd gnd cell_6t
Xbit_r370_c118 bl[118] br[118] wl[370] vdd gnd cell_6t
Xbit_r371_c118 bl[118] br[118] wl[371] vdd gnd cell_6t
Xbit_r372_c118 bl[118] br[118] wl[372] vdd gnd cell_6t
Xbit_r373_c118 bl[118] br[118] wl[373] vdd gnd cell_6t
Xbit_r374_c118 bl[118] br[118] wl[374] vdd gnd cell_6t
Xbit_r375_c118 bl[118] br[118] wl[375] vdd gnd cell_6t
Xbit_r376_c118 bl[118] br[118] wl[376] vdd gnd cell_6t
Xbit_r377_c118 bl[118] br[118] wl[377] vdd gnd cell_6t
Xbit_r378_c118 bl[118] br[118] wl[378] vdd gnd cell_6t
Xbit_r379_c118 bl[118] br[118] wl[379] vdd gnd cell_6t
Xbit_r380_c118 bl[118] br[118] wl[380] vdd gnd cell_6t
Xbit_r381_c118 bl[118] br[118] wl[381] vdd gnd cell_6t
Xbit_r382_c118 bl[118] br[118] wl[382] vdd gnd cell_6t
Xbit_r383_c118 bl[118] br[118] wl[383] vdd gnd cell_6t
Xbit_r384_c118 bl[118] br[118] wl[384] vdd gnd cell_6t
Xbit_r385_c118 bl[118] br[118] wl[385] vdd gnd cell_6t
Xbit_r386_c118 bl[118] br[118] wl[386] vdd gnd cell_6t
Xbit_r387_c118 bl[118] br[118] wl[387] vdd gnd cell_6t
Xbit_r388_c118 bl[118] br[118] wl[388] vdd gnd cell_6t
Xbit_r389_c118 bl[118] br[118] wl[389] vdd gnd cell_6t
Xbit_r390_c118 bl[118] br[118] wl[390] vdd gnd cell_6t
Xbit_r391_c118 bl[118] br[118] wl[391] vdd gnd cell_6t
Xbit_r392_c118 bl[118] br[118] wl[392] vdd gnd cell_6t
Xbit_r393_c118 bl[118] br[118] wl[393] vdd gnd cell_6t
Xbit_r394_c118 bl[118] br[118] wl[394] vdd gnd cell_6t
Xbit_r395_c118 bl[118] br[118] wl[395] vdd gnd cell_6t
Xbit_r396_c118 bl[118] br[118] wl[396] vdd gnd cell_6t
Xbit_r397_c118 bl[118] br[118] wl[397] vdd gnd cell_6t
Xbit_r398_c118 bl[118] br[118] wl[398] vdd gnd cell_6t
Xbit_r399_c118 bl[118] br[118] wl[399] vdd gnd cell_6t
Xbit_r400_c118 bl[118] br[118] wl[400] vdd gnd cell_6t
Xbit_r401_c118 bl[118] br[118] wl[401] vdd gnd cell_6t
Xbit_r402_c118 bl[118] br[118] wl[402] vdd gnd cell_6t
Xbit_r403_c118 bl[118] br[118] wl[403] vdd gnd cell_6t
Xbit_r404_c118 bl[118] br[118] wl[404] vdd gnd cell_6t
Xbit_r405_c118 bl[118] br[118] wl[405] vdd gnd cell_6t
Xbit_r406_c118 bl[118] br[118] wl[406] vdd gnd cell_6t
Xbit_r407_c118 bl[118] br[118] wl[407] vdd gnd cell_6t
Xbit_r408_c118 bl[118] br[118] wl[408] vdd gnd cell_6t
Xbit_r409_c118 bl[118] br[118] wl[409] vdd gnd cell_6t
Xbit_r410_c118 bl[118] br[118] wl[410] vdd gnd cell_6t
Xbit_r411_c118 bl[118] br[118] wl[411] vdd gnd cell_6t
Xbit_r412_c118 bl[118] br[118] wl[412] vdd gnd cell_6t
Xbit_r413_c118 bl[118] br[118] wl[413] vdd gnd cell_6t
Xbit_r414_c118 bl[118] br[118] wl[414] vdd gnd cell_6t
Xbit_r415_c118 bl[118] br[118] wl[415] vdd gnd cell_6t
Xbit_r416_c118 bl[118] br[118] wl[416] vdd gnd cell_6t
Xbit_r417_c118 bl[118] br[118] wl[417] vdd gnd cell_6t
Xbit_r418_c118 bl[118] br[118] wl[418] vdd gnd cell_6t
Xbit_r419_c118 bl[118] br[118] wl[419] vdd gnd cell_6t
Xbit_r420_c118 bl[118] br[118] wl[420] vdd gnd cell_6t
Xbit_r421_c118 bl[118] br[118] wl[421] vdd gnd cell_6t
Xbit_r422_c118 bl[118] br[118] wl[422] vdd gnd cell_6t
Xbit_r423_c118 bl[118] br[118] wl[423] vdd gnd cell_6t
Xbit_r424_c118 bl[118] br[118] wl[424] vdd gnd cell_6t
Xbit_r425_c118 bl[118] br[118] wl[425] vdd gnd cell_6t
Xbit_r426_c118 bl[118] br[118] wl[426] vdd gnd cell_6t
Xbit_r427_c118 bl[118] br[118] wl[427] vdd gnd cell_6t
Xbit_r428_c118 bl[118] br[118] wl[428] vdd gnd cell_6t
Xbit_r429_c118 bl[118] br[118] wl[429] vdd gnd cell_6t
Xbit_r430_c118 bl[118] br[118] wl[430] vdd gnd cell_6t
Xbit_r431_c118 bl[118] br[118] wl[431] vdd gnd cell_6t
Xbit_r432_c118 bl[118] br[118] wl[432] vdd gnd cell_6t
Xbit_r433_c118 bl[118] br[118] wl[433] vdd gnd cell_6t
Xbit_r434_c118 bl[118] br[118] wl[434] vdd gnd cell_6t
Xbit_r435_c118 bl[118] br[118] wl[435] vdd gnd cell_6t
Xbit_r436_c118 bl[118] br[118] wl[436] vdd gnd cell_6t
Xbit_r437_c118 bl[118] br[118] wl[437] vdd gnd cell_6t
Xbit_r438_c118 bl[118] br[118] wl[438] vdd gnd cell_6t
Xbit_r439_c118 bl[118] br[118] wl[439] vdd gnd cell_6t
Xbit_r440_c118 bl[118] br[118] wl[440] vdd gnd cell_6t
Xbit_r441_c118 bl[118] br[118] wl[441] vdd gnd cell_6t
Xbit_r442_c118 bl[118] br[118] wl[442] vdd gnd cell_6t
Xbit_r443_c118 bl[118] br[118] wl[443] vdd gnd cell_6t
Xbit_r444_c118 bl[118] br[118] wl[444] vdd gnd cell_6t
Xbit_r445_c118 bl[118] br[118] wl[445] vdd gnd cell_6t
Xbit_r446_c118 bl[118] br[118] wl[446] vdd gnd cell_6t
Xbit_r447_c118 bl[118] br[118] wl[447] vdd gnd cell_6t
Xbit_r448_c118 bl[118] br[118] wl[448] vdd gnd cell_6t
Xbit_r449_c118 bl[118] br[118] wl[449] vdd gnd cell_6t
Xbit_r450_c118 bl[118] br[118] wl[450] vdd gnd cell_6t
Xbit_r451_c118 bl[118] br[118] wl[451] vdd gnd cell_6t
Xbit_r452_c118 bl[118] br[118] wl[452] vdd gnd cell_6t
Xbit_r453_c118 bl[118] br[118] wl[453] vdd gnd cell_6t
Xbit_r454_c118 bl[118] br[118] wl[454] vdd gnd cell_6t
Xbit_r455_c118 bl[118] br[118] wl[455] vdd gnd cell_6t
Xbit_r456_c118 bl[118] br[118] wl[456] vdd gnd cell_6t
Xbit_r457_c118 bl[118] br[118] wl[457] vdd gnd cell_6t
Xbit_r458_c118 bl[118] br[118] wl[458] vdd gnd cell_6t
Xbit_r459_c118 bl[118] br[118] wl[459] vdd gnd cell_6t
Xbit_r460_c118 bl[118] br[118] wl[460] vdd gnd cell_6t
Xbit_r461_c118 bl[118] br[118] wl[461] vdd gnd cell_6t
Xbit_r462_c118 bl[118] br[118] wl[462] vdd gnd cell_6t
Xbit_r463_c118 bl[118] br[118] wl[463] vdd gnd cell_6t
Xbit_r464_c118 bl[118] br[118] wl[464] vdd gnd cell_6t
Xbit_r465_c118 bl[118] br[118] wl[465] vdd gnd cell_6t
Xbit_r466_c118 bl[118] br[118] wl[466] vdd gnd cell_6t
Xbit_r467_c118 bl[118] br[118] wl[467] vdd gnd cell_6t
Xbit_r468_c118 bl[118] br[118] wl[468] vdd gnd cell_6t
Xbit_r469_c118 bl[118] br[118] wl[469] vdd gnd cell_6t
Xbit_r470_c118 bl[118] br[118] wl[470] vdd gnd cell_6t
Xbit_r471_c118 bl[118] br[118] wl[471] vdd gnd cell_6t
Xbit_r472_c118 bl[118] br[118] wl[472] vdd gnd cell_6t
Xbit_r473_c118 bl[118] br[118] wl[473] vdd gnd cell_6t
Xbit_r474_c118 bl[118] br[118] wl[474] vdd gnd cell_6t
Xbit_r475_c118 bl[118] br[118] wl[475] vdd gnd cell_6t
Xbit_r476_c118 bl[118] br[118] wl[476] vdd gnd cell_6t
Xbit_r477_c118 bl[118] br[118] wl[477] vdd gnd cell_6t
Xbit_r478_c118 bl[118] br[118] wl[478] vdd gnd cell_6t
Xbit_r479_c118 bl[118] br[118] wl[479] vdd gnd cell_6t
Xbit_r480_c118 bl[118] br[118] wl[480] vdd gnd cell_6t
Xbit_r481_c118 bl[118] br[118] wl[481] vdd gnd cell_6t
Xbit_r482_c118 bl[118] br[118] wl[482] vdd gnd cell_6t
Xbit_r483_c118 bl[118] br[118] wl[483] vdd gnd cell_6t
Xbit_r484_c118 bl[118] br[118] wl[484] vdd gnd cell_6t
Xbit_r485_c118 bl[118] br[118] wl[485] vdd gnd cell_6t
Xbit_r486_c118 bl[118] br[118] wl[486] vdd gnd cell_6t
Xbit_r487_c118 bl[118] br[118] wl[487] vdd gnd cell_6t
Xbit_r488_c118 bl[118] br[118] wl[488] vdd gnd cell_6t
Xbit_r489_c118 bl[118] br[118] wl[489] vdd gnd cell_6t
Xbit_r490_c118 bl[118] br[118] wl[490] vdd gnd cell_6t
Xbit_r491_c118 bl[118] br[118] wl[491] vdd gnd cell_6t
Xbit_r492_c118 bl[118] br[118] wl[492] vdd gnd cell_6t
Xbit_r493_c118 bl[118] br[118] wl[493] vdd gnd cell_6t
Xbit_r494_c118 bl[118] br[118] wl[494] vdd gnd cell_6t
Xbit_r495_c118 bl[118] br[118] wl[495] vdd gnd cell_6t
Xbit_r496_c118 bl[118] br[118] wl[496] vdd gnd cell_6t
Xbit_r497_c118 bl[118] br[118] wl[497] vdd gnd cell_6t
Xbit_r498_c118 bl[118] br[118] wl[498] vdd gnd cell_6t
Xbit_r499_c118 bl[118] br[118] wl[499] vdd gnd cell_6t
Xbit_r500_c118 bl[118] br[118] wl[500] vdd gnd cell_6t
Xbit_r501_c118 bl[118] br[118] wl[501] vdd gnd cell_6t
Xbit_r502_c118 bl[118] br[118] wl[502] vdd gnd cell_6t
Xbit_r503_c118 bl[118] br[118] wl[503] vdd gnd cell_6t
Xbit_r504_c118 bl[118] br[118] wl[504] vdd gnd cell_6t
Xbit_r505_c118 bl[118] br[118] wl[505] vdd gnd cell_6t
Xbit_r506_c118 bl[118] br[118] wl[506] vdd gnd cell_6t
Xbit_r507_c118 bl[118] br[118] wl[507] vdd gnd cell_6t
Xbit_r508_c118 bl[118] br[118] wl[508] vdd gnd cell_6t
Xbit_r509_c118 bl[118] br[118] wl[509] vdd gnd cell_6t
Xbit_r510_c118 bl[118] br[118] wl[510] vdd gnd cell_6t
Xbit_r511_c118 bl[118] br[118] wl[511] vdd gnd cell_6t
Xbit_r0_c119 bl[119] br[119] wl[0] vdd gnd cell_6t
Xbit_r1_c119 bl[119] br[119] wl[1] vdd gnd cell_6t
Xbit_r2_c119 bl[119] br[119] wl[2] vdd gnd cell_6t
Xbit_r3_c119 bl[119] br[119] wl[3] vdd gnd cell_6t
Xbit_r4_c119 bl[119] br[119] wl[4] vdd gnd cell_6t
Xbit_r5_c119 bl[119] br[119] wl[5] vdd gnd cell_6t
Xbit_r6_c119 bl[119] br[119] wl[6] vdd gnd cell_6t
Xbit_r7_c119 bl[119] br[119] wl[7] vdd gnd cell_6t
Xbit_r8_c119 bl[119] br[119] wl[8] vdd gnd cell_6t
Xbit_r9_c119 bl[119] br[119] wl[9] vdd gnd cell_6t
Xbit_r10_c119 bl[119] br[119] wl[10] vdd gnd cell_6t
Xbit_r11_c119 bl[119] br[119] wl[11] vdd gnd cell_6t
Xbit_r12_c119 bl[119] br[119] wl[12] vdd gnd cell_6t
Xbit_r13_c119 bl[119] br[119] wl[13] vdd gnd cell_6t
Xbit_r14_c119 bl[119] br[119] wl[14] vdd gnd cell_6t
Xbit_r15_c119 bl[119] br[119] wl[15] vdd gnd cell_6t
Xbit_r16_c119 bl[119] br[119] wl[16] vdd gnd cell_6t
Xbit_r17_c119 bl[119] br[119] wl[17] vdd gnd cell_6t
Xbit_r18_c119 bl[119] br[119] wl[18] vdd gnd cell_6t
Xbit_r19_c119 bl[119] br[119] wl[19] vdd gnd cell_6t
Xbit_r20_c119 bl[119] br[119] wl[20] vdd gnd cell_6t
Xbit_r21_c119 bl[119] br[119] wl[21] vdd gnd cell_6t
Xbit_r22_c119 bl[119] br[119] wl[22] vdd gnd cell_6t
Xbit_r23_c119 bl[119] br[119] wl[23] vdd gnd cell_6t
Xbit_r24_c119 bl[119] br[119] wl[24] vdd gnd cell_6t
Xbit_r25_c119 bl[119] br[119] wl[25] vdd gnd cell_6t
Xbit_r26_c119 bl[119] br[119] wl[26] vdd gnd cell_6t
Xbit_r27_c119 bl[119] br[119] wl[27] vdd gnd cell_6t
Xbit_r28_c119 bl[119] br[119] wl[28] vdd gnd cell_6t
Xbit_r29_c119 bl[119] br[119] wl[29] vdd gnd cell_6t
Xbit_r30_c119 bl[119] br[119] wl[30] vdd gnd cell_6t
Xbit_r31_c119 bl[119] br[119] wl[31] vdd gnd cell_6t
Xbit_r32_c119 bl[119] br[119] wl[32] vdd gnd cell_6t
Xbit_r33_c119 bl[119] br[119] wl[33] vdd gnd cell_6t
Xbit_r34_c119 bl[119] br[119] wl[34] vdd gnd cell_6t
Xbit_r35_c119 bl[119] br[119] wl[35] vdd gnd cell_6t
Xbit_r36_c119 bl[119] br[119] wl[36] vdd gnd cell_6t
Xbit_r37_c119 bl[119] br[119] wl[37] vdd gnd cell_6t
Xbit_r38_c119 bl[119] br[119] wl[38] vdd gnd cell_6t
Xbit_r39_c119 bl[119] br[119] wl[39] vdd gnd cell_6t
Xbit_r40_c119 bl[119] br[119] wl[40] vdd gnd cell_6t
Xbit_r41_c119 bl[119] br[119] wl[41] vdd gnd cell_6t
Xbit_r42_c119 bl[119] br[119] wl[42] vdd gnd cell_6t
Xbit_r43_c119 bl[119] br[119] wl[43] vdd gnd cell_6t
Xbit_r44_c119 bl[119] br[119] wl[44] vdd gnd cell_6t
Xbit_r45_c119 bl[119] br[119] wl[45] vdd gnd cell_6t
Xbit_r46_c119 bl[119] br[119] wl[46] vdd gnd cell_6t
Xbit_r47_c119 bl[119] br[119] wl[47] vdd gnd cell_6t
Xbit_r48_c119 bl[119] br[119] wl[48] vdd gnd cell_6t
Xbit_r49_c119 bl[119] br[119] wl[49] vdd gnd cell_6t
Xbit_r50_c119 bl[119] br[119] wl[50] vdd gnd cell_6t
Xbit_r51_c119 bl[119] br[119] wl[51] vdd gnd cell_6t
Xbit_r52_c119 bl[119] br[119] wl[52] vdd gnd cell_6t
Xbit_r53_c119 bl[119] br[119] wl[53] vdd gnd cell_6t
Xbit_r54_c119 bl[119] br[119] wl[54] vdd gnd cell_6t
Xbit_r55_c119 bl[119] br[119] wl[55] vdd gnd cell_6t
Xbit_r56_c119 bl[119] br[119] wl[56] vdd gnd cell_6t
Xbit_r57_c119 bl[119] br[119] wl[57] vdd gnd cell_6t
Xbit_r58_c119 bl[119] br[119] wl[58] vdd gnd cell_6t
Xbit_r59_c119 bl[119] br[119] wl[59] vdd gnd cell_6t
Xbit_r60_c119 bl[119] br[119] wl[60] vdd gnd cell_6t
Xbit_r61_c119 bl[119] br[119] wl[61] vdd gnd cell_6t
Xbit_r62_c119 bl[119] br[119] wl[62] vdd gnd cell_6t
Xbit_r63_c119 bl[119] br[119] wl[63] vdd gnd cell_6t
Xbit_r64_c119 bl[119] br[119] wl[64] vdd gnd cell_6t
Xbit_r65_c119 bl[119] br[119] wl[65] vdd gnd cell_6t
Xbit_r66_c119 bl[119] br[119] wl[66] vdd gnd cell_6t
Xbit_r67_c119 bl[119] br[119] wl[67] vdd gnd cell_6t
Xbit_r68_c119 bl[119] br[119] wl[68] vdd gnd cell_6t
Xbit_r69_c119 bl[119] br[119] wl[69] vdd gnd cell_6t
Xbit_r70_c119 bl[119] br[119] wl[70] vdd gnd cell_6t
Xbit_r71_c119 bl[119] br[119] wl[71] vdd gnd cell_6t
Xbit_r72_c119 bl[119] br[119] wl[72] vdd gnd cell_6t
Xbit_r73_c119 bl[119] br[119] wl[73] vdd gnd cell_6t
Xbit_r74_c119 bl[119] br[119] wl[74] vdd gnd cell_6t
Xbit_r75_c119 bl[119] br[119] wl[75] vdd gnd cell_6t
Xbit_r76_c119 bl[119] br[119] wl[76] vdd gnd cell_6t
Xbit_r77_c119 bl[119] br[119] wl[77] vdd gnd cell_6t
Xbit_r78_c119 bl[119] br[119] wl[78] vdd gnd cell_6t
Xbit_r79_c119 bl[119] br[119] wl[79] vdd gnd cell_6t
Xbit_r80_c119 bl[119] br[119] wl[80] vdd gnd cell_6t
Xbit_r81_c119 bl[119] br[119] wl[81] vdd gnd cell_6t
Xbit_r82_c119 bl[119] br[119] wl[82] vdd gnd cell_6t
Xbit_r83_c119 bl[119] br[119] wl[83] vdd gnd cell_6t
Xbit_r84_c119 bl[119] br[119] wl[84] vdd gnd cell_6t
Xbit_r85_c119 bl[119] br[119] wl[85] vdd gnd cell_6t
Xbit_r86_c119 bl[119] br[119] wl[86] vdd gnd cell_6t
Xbit_r87_c119 bl[119] br[119] wl[87] vdd gnd cell_6t
Xbit_r88_c119 bl[119] br[119] wl[88] vdd gnd cell_6t
Xbit_r89_c119 bl[119] br[119] wl[89] vdd gnd cell_6t
Xbit_r90_c119 bl[119] br[119] wl[90] vdd gnd cell_6t
Xbit_r91_c119 bl[119] br[119] wl[91] vdd gnd cell_6t
Xbit_r92_c119 bl[119] br[119] wl[92] vdd gnd cell_6t
Xbit_r93_c119 bl[119] br[119] wl[93] vdd gnd cell_6t
Xbit_r94_c119 bl[119] br[119] wl[94] vdd gnd cell_6t
Xbit_r95_c119 bl[119] br[119] wl[95] vdd gnd cell_6t
Xbit_r96_c119 bl[119] br[119] wl[96] vdd gnd cell_6t
Xbit_r97_c119 bl[119] br[119] wl[97] vdd gnd cell_6t
Xbit_r98_c119 bl[119] br[119] wl[98] vdd gnd cell_6t
Xbit_r99_c119 bl[119] br[119] wl[99] vdd gnd cell_6t
Xbit_r100_c119 bl[119] br[119] wl[100] vdd gnd cell_6t
Xbit_r101_c119 bl[119] br[119] wl[101] vdd gnd cell_6t
Xbit_r102_c119 bl[119] br[119] wl[102] vdd gnd cell_6t
Xbit_r103_c119 bl[119] br[119] wl[103] vdd gnd cell_6t
Xbit_r104_c119 bl[119] br[119] wl[104] vdd gnd cell_6t
Xbit_r105_c119 bl[119] br[119] wl[105] vdd gnd cell_6t
Xbit_r106_c119 bl[119] br[119] wl[106] vdd gnd cell_6t
Xbit_r107_c119 bl[119] br[119] wl[107] vdd gnd cell_6t
Xbit_r108_c119 bl[119] br[119] wl[108] vdd gnd cell_6t
Xbit_r109_c119 bl[119] br[119] wl[109] vdd gnd cell_6t
Xbit_r110_c119 bl[119] br[119] wl[110] vdd gnd cell_6t
Xbit_r111_c119 bl[119] br[119] wl[111] vdd gnd cell_6t
Xbit_r112_c119 bl[119] br[119] wl[112] vdd gnd cell_6t
Xbit_r113_c119 bl[119] br[119] wl[113] vdd gnd cell_6t
Xbit_r114_c119 bl[119] br[119] wl[114] vdd gnd cell_6t
Xbit_r115_c119 bl[119] br[119] wl[115] vdd gnd cell_6t
Xbit_r116_c119 bl[119] br[119] wl[116] vdd gnd cell_6t
Xbit_r117_c119 bl[119] br[119] wl[117] vdd gnd cell_6t
Xbit_r118_c119 bl[119] br[119] wl[118] vdd gnd cell_6t
Xbit_r119_c119 bl[119] br[119] wl[119] vdd gnd cell_6t
Xbit_r120_c119 bl[119] br[119] wl[120] vdd gnd cell_6t
Xbit_r121_c119 bl[119] br[119] wl[121] vdd gnd cell_6t
Xbit_r122_c119 bl[119] br[119] wl[122] vdd gnd cell_6t
Xbit_r123_c119 bl[119] br[119] wl[123] vdd gnd cell_6t
Xbit_r124_c119 bl[119] br[119] wl[124] vdd gnd cell_6t
Xbit_r125_c119 bl[119] br[119] wl[125] vdd gnd cell_6t
Xbit_r126_c119 bl[119] br[119] wl[126] vdd gnd cell_6t
Xbit_r127_c119 bl[119] br[119] wl[127] vdd gnd cell_6t
Xbit_r128_c119 bl[119] br[119] wl[128] vdd gnd cell_6t
Xbit_r129_c119 bl[119] br[119] wl[129] vdd gnd cell_6t
Xbit_r130_c119 bl[119] br[119] wl[130] vdd gnd cell_6t
Xbit_r131_c119 bl[119] br[119] wl[131] vdd gnd cell_6t
Xbit_r132_c119 bl[119] br[119] wl[132] vdd gnd cell_6t
Xbit_r133_c119 bl[119] br[119] wl[133] vdd gnd cell_6t
Xbit_r134_c119 bl[119] br[119] wl[134] vdd gnd cell_6t
Xbit_r135_c119 bl[119] br[119] wl[135] vdd gnd cell_6t
Xbit_r136_c119 bl[119] br[119] wl[136] vdd gnd cell_6t
Xbit_r137_c119 bl[119] br[119] wl[137] vdd gnd cell_6t
Xbit_r138_c119 bl[119] br[119] wl[138] vdd gnd cell_6t
Xbit_r139_c119 bl[119] br[119] wl[139] vdd gnd cell_6t
Xbit_r140_c119 bl[119] br[119] wl[140] vdd gnd cell_6t
Xbit_r141_c119 bl[119] br[119] wl[141] vdd gnd cell_6t
Xbit_r142_c119 bl[119] br[119] wl[142] vdd gnd cell_6t
Xbit_r143_c119 bl[119] br[119] wl[143] vdd gnd cell_6t
Xbit_r144_c119 bl[119] br[119] wl[144] vdd gnd cell_6t
Xbit_r145_c119 bl[119] br[119] wl[145] vdd gnd cell_6t
Xbit_r146_c119 bl[119] br[119] wl[146] vdd gnd cell_6t
Xbit_r147_c119 bl[119] br[119] wl[147] vdd gnd cell_6t
Xbit_r148_c119 bl[119] br[119] wl[148] vdd gnd cell_6t
Xbit_r149_c119 bl[119] br[119] wl[149] vdd gnd cell_6t
Xbit_r150_c119 bl[119] br[119] wl[150] vdd gnd cell_6t
Xbit_r151_c119 bl[119] br[119] wl[151] vdd gnd cell_6t
Xbit_r152_c119 bl[119] br[119] wl[152] vdd gnd cell_6t
Xbit_r153_c119 bl[119] br[119] wl[153] vdd gnd cell_6t
Xbit_r154_c119 bl[119] br[119] wl[154] vdd gnd cell_6t
Xbit_r155_c119 bl[119] br[119] wl[155] vdd gnd cell_6t
Xbit_r156_c119 bl[119] br[119] wl[156] vdd gnd cell_6t
Xbit_r157_c119 bl[119] br[119] wl[157] vdd gnd cell_6t
Xbit_r158_c119 bl[119] br[119] wl[158] vdd gnd cell_6t
Xbit_r159_c119 bl[119] br[119] wl[159] vdd gnd cell_6t
Xbit_r160_c119 bl[119] br[119] wl[160] vdd gnd cell_6t
Xbit_r161_c119 bl[119] br[119] wl[161] vdd gnd cell_6t
Xbit_r162_c119 bl[119] br[119] wl[162] vdd gnd cell_6t
Xbit_r163_c119 bl[119] br[119] wl[163] vdd gnd cell_6t
Xbit_r164_c119 bl[119] br[119] wl[164] vdd gnd cell_6t
Xbit_r165_c119 bl[119] br[119] wl[165] vdd gnd cell_6t
Xbit_r166_c119 bl[119] br[119] wl[166] vdd gnd cell_6t
Xbit_r167_c119 bl[119] br[119] wl[167] vdd gnd cell_6t
Xbit_r168_c119 bl[119] br[119] wl[168] vdd gnd cell_6t
Xbit_r169_c119 bl[119] br[119] wl[169] vdd gnd cell_6t
Xbit_r170_c119 bl[119] br[119] wl[170] vdd gnd cell_6t
Xbit_r171_c119 bl[119] br[119] wl[171] vdd gnd cell_6t
Xbit_r172_c119 bl[119] br[119] wl[172] vdd gnd cell_6t
Xbit_r173_c119 bl[119] br[119] wl[173] vdd gnd cell_6t
Xbit_r174_c119 bl[119] br[119] wl[174] vdd gnd cell_6t
Xbit_r175_c119 bl[119] br[119] wl[175] vdd gnd cell_6t
Xbit_r176_c119 bl[119] br[119] wl[176] vdd gnd cell_6t
Xbit_r177_c119 bl[119] br[119] wl[177] vdd gnd cell_6t
Xbit_r178_c119 bl[119] br[119] wl[178] vdd gnd cell_6t
Xbit_r179_c119 bl[119] br[119] wl[179] vdd gnd cell_6t
Xbit_r180_c119 bl[119] br[119] wl[180] vdd gnd cell_6t
Xbit_r181_c119 bl[119] br[119] wl[181] vdd gnd cell_6t
Xbit_r182_c119 bl[119] br[119] wl[182] vdd gnd cell_6t
Xbit_r183_c119 bl[119] br[119] wl[183] vdd gnd cell_6t
Xbit_r184_c119 bl[119] br[119] wl[184] vdd gnd cell_6t
Xbit_r185_c119 bl[119] br[119] wl[185] vdd gnd cell_6t
Xbit_r186_c119 bl[119] br[119] wl[186] vdd gnd cell_6t
Xbit_r187_c119 bl[119] br[119] wl[187] vdd gnd cell_6t
Xbit_r188_c119 bl[119] br[119] wl[188] vdd gnd cell_6t
Xbit_r189_c119 bl[119] br[119] wl[189] vdd gnd cell_6t
Xbit_r190_c119 bl[119] br[119] wl[190] vdd gnd cell_6t
Xbit_r191_c119 bl[119] br[119] wl[191] vdd gnd cell_6t
Xbit_r192_c119 bl[119] br[119] wl[192] vdd gnd cell_6t
Xbit_r193_c119 bl[119] br[119] wl[193] vdd gnd cell_6t
Xbit_r194_c119 bl[119] br[119] wl[194] vdd gnd cell_6t
Xbit_r195_c119 bl[119] br[119] wl[195] vdd gnd cell_6t
Xbit_r196_c119 bl[119] br[119] wl[196] vdd gnd cell_6t
Xbit_r197_c119 bl[119] br[119] wl[197] vdd gnd cell_6t
Xbit_r198_c119 bl[119] br[119] wl[198] vdd gnd cell_6t
Xbit_r199_c119 bl[119] br[119] wl[199] vdd gnd cell_6t
Xbit_r200_c119 bl[119] br[119] wl[200] vdd gnd cell_6t
Xbit_r201_c119 bl[119] br[119] wl[201] vdd gnd cell_6t
Xbit_r202_c119 bl[119] br[119] wl[202] vdd gnd cell_6t
Xbit_r203_c119 bl[119] br[119] wl[203] vdd gnd cell_6t
Xbit_r204_c119 bl[119] br[119] wl[204] vdd gnd cell_6t
Xbit_r205_c119 bl[119] br[119] wl[205] vdd gnd cell_6t
Xbit_r206_c119 bl[119] br[119] wl[206] vdd gnd cell_6t
Xbit_r207_c119 bl[119] br[119] wl[207] vdd gnd cell_6t
Xbit_r208_c119 bl[119] br[119] wl[208] vdd gnd cell_6t
Xbit_r209_c119 bl[119] br[119] wl[209] vdd gnd cell_6t
Xbit_r210_c119 bl[119] br[119] wl[210] vdd gnd cell_6t
Xbit_r211_c119 bl[119] br[119] wl[211] vdd gnd cell_6t
Xbit_r212_c119 bl[119] br[119] wl[212] vdd gnd cell_6t
Xbit_r213_c119 bl[119] br[119] wl[213] vdd gnd cell_6t
Xbit_r214_c119 bl[119] br[119] wl[214] vdd gnd cell_6t
Xbit_r215_c119 bl[119] br[119] wl[215] vdd gnd cell_6t
Xbit_r216_c119 bl[119] br[119] wl[216] vdd gnd cell_6t
Xbit_r217_c119 bl[119] br[119] wl[217] vdd gnd cell_6t
Xbit_r218_c119 bl[119] br[119] wl[218] vdd gnd cell_6t
Xbit_r219_c119 bl[119] br[119] wl[219] vdd gnd cell_6t
Xbit_r220_c119 bl[119] br[119] wl[220] vdd gnd cell_6t
Xbit_r221_c119 bl[119] br[119] wl[221] vdd gnd cell_6t
Xbit_r222_c119 bl[119] br[119] wl[222] vdd gnd cell_6t
Xbit_r223_c119 bl[119] br[119] wl[223] vdd gnd cell_6t
Xbit_r224_c119 bl[119] br[119] wl[224] vdd gnd cell_6t
Xbit_r225_c119 bl[119] br[119] wl[225] vdd gnd cell_6t
Xbit_r226_c119 bl[119] br[119] wl[226] vdd gnd cell_6t
Xbit_r227_c119 bl[119] br[119] wl[227] vdd gnd cell_6t
Xbit_r228_c119 bl[119] br[119] wl[228] vdd gnd cell_6t
Xbit_r229_c119 bl[119] br[119] wl[229] vdd gnd cell_6t
Xbit_r230_c119 bl[119] br[119] wl[230] vdd gnd cell_6t
Xbit_r231_c119 bl[119] br[119] wl[231] vdd gnd cell_6t
Xbit_r232_c119 bl[119] br[119] wl[232] vdd gnd cell_6t
Xbit_r233_c119 bl[119] br[119] wl[233] vdd gnd cell_6t
Xbit_r234_c119 bl[119] br[119] wl[234] vdd gnd cell_6t
Xbit_r235_c119 bl[119] br[119] wl[235] vdd gnd cell_6t
Xbit_r236_c119 bl[119] br[119] wl[236] vdd gnd cell_6t
Xbit_r237_c119 bl[119] br[119] wl[237] vdd gnd cell_6t
Xbit_r238_c119 bl[119] br[119] wl[238] vdd gnd cell_6t
Xbit_r239_c119 bl[119] br[119] wl[239] vdd gnd cell_6t
Xbit_r240_c119 bl[119] br[119] wl[240] vdd gnd cell_6t
Xbit_r241_c119 bl[119] br[119] wl[241] vdd gnd cell_6t
Xbit_r242_c119 bl[119] br[119] wl[242] vdd gnd cell_6t
Xbit_r243_c119 bl[119] br[119] wl[243] vdd gnd cell_6t
Xbit_r244_c119 bl[119] br[119] wl[244] vdd gnd cell_6t
Xbit_r245_c119 bl[119] br[119] wl[245] vdd gnd cell_6t
Xbit_r246_c119 bl[119] br[119] wl[246] vdd gnd cell_6t
Xbit_r247_c119 bl[119] br[119] wl[247] vdd gnd cell_6t
Xbit_r248_c119 bl[119] br[119] wl[248] vdd gnd cell_6t
Xbit_r249_c119 bl[119] br[119] wl[249] vdd gnd cell_6t
Xbit_r250_c119 bl[119] br[119] wl[250] vdd gnd cell_6t
Xbit_r251_c119 bl[119] br[119] wl[251] vdd gnd cell_6t
Xbit_r252_c119 bl[119] br[119] wl[252] vdd gnd cell_6t
Xbit_r253_c119 bl[119] br[119] wl[253] vdd gnd cell_6t
Xbit_r254_c119 bl[119] br[119] wl[254] vdd gnd cell_6t
Xbit_r255_c119 bl[119] br[119] wl[255] vdd gnd cell_6t
Xbit_r256_c119 bl[119] br[119] wl[256] vdd gnd cell_6t
Xbit_r257_c119 bl[119] br[119] wl[257] vdd gnd cell_6t
Xbit_r258_c119 bl[119] br[119] wl[258] vdd gnd cell_6t
Xbit_r259_c119 bl[119] br[119] wl[259] vdd gnd cell_6t
Xbit_r260_c119 bl[119] br[119] wl[260] vdd gnd cell_6t
Xbit_r261_c119 bl[119] br[119] wl[261] vdd gnd cell_6t
Xbit_r262_c119 bl[119] br[119] wl[262] vdd gnd cell_6t
Xbit_r263_c119 bl[119] br[119] wl[263] vdd gnd cell_6t
Xbit_r264_c119 bl[119] br[119] wl[264] vdd gnd cell_6t
Xbit_r265_c119 bl[119] br[119] wl[265] vdd gnd cell_6t
Xbit_r266_c119 bl[119] br[119] wl[266] vdd gnd cell_6t
Xbit_r267_c119 bl[119] br[119] wl[267] vdd gnd cell_6t
Xbit_r268_c119 bl[119] br[119] wl[268] vdd gnd cell_6t
Xbit_r269_c119 bl[119] br[119] wl[269] vdd gnd cell_6t
Xbit_r270_c119 bl[119] br[119] wl[270] vdd gnd cell_6t
Xbit_r271_c119 bl[119] br[119] wl[271] vdd gnd cell_6t
Xbit_r272_c119 bl[119] br[119] wl[272] vdd gnd cell_6t
Xbit_r273_c119 bl[119] br[119] wl[273] vdd gnd cell_6t
Xbit_r274_c119 bl[119] br[119] wl[274] vdd gnd cell_6t
Xbit_r275_c119 bl[119] br[119] wl[275] vdd gnd cell_6t
Xbit_r276_c119 bl[119] br[119] wl[276] vdd gnd cell_6t
Xbit_r277_c119 bl[119] br[119] wl[277] vdd gnd cell_6t
Xbit_r278_c119 bl[119] br[119] wl[278] vdd gnd cell_6t
Xbit_r279_c119 bl[119] br[119] wl[279] vdd gnd cell_6t
Xbit_r280_c119 bl[119] br[119] wl[280] vdd gnd cell_6t
Xbit_r281_c119 bl[119] br[119] wl[281] vdd gnd cell_6t
Xbit_r282_c119 bl[119] br[119] wl[282] vdd gnd cell_6t
Xbit_r283_c119 bl[119] br[119] wl[283] vdd gnd cell_6t
Xbit_r284_c119 bl[119] br[119] wl[284] vdd gnd cell_6t
Xbit_r285_c119 bl[119] br[119] wl[285] vdd gnd cell_6t
Xbit_r286_c119 bl[119] br[119] wl[286] vdd gnd cell_6t
Xbit_r287_c119 bl[119] br[119] wl[287] vdd gnd cell_6t
Xbit_r288_c119 bl[119] br[119] wl[288] vdd gnd cell_6t
Xbit_r289_c119 bl[119] br[119] wl[289] vdd gnd cell_6t
Xbit_r290_c119 bl[119] br[119] wl[290] vdd gnd cell_6t
Xbit_r291_c119 bl[119] br[119] wl[291] vdd gnd cell_6t
Xbit_r292_c119 bl[119] br[119] wl[292] vdd gnd cell_6t
Xbit_r293_c119 bl[119] br[119] wl[293] vdd gnd cell_6t
Xbit_r294_c119 bl[119] br[119] wl[294] vdd gnd cell_6t
Xbit_r295_c119 bl[119] br[119] wl[295] vdd gnd cell_6t
Xbit_r296_c119 bl[119] br[119] wl[296] vdd gnd cell_6t
Xbit_r297_c119 bl[119] br[119] wl[297] vdd gnd cell_6t
Xbit_r298_c119 bl[119] br[119] wl[298] vdd gnd cell_6t
Xbit_r299_c119 bl[119] br[119] wl[299] vdd gnd cell_6t
Xbit_r300_c119 bl[119] br[119] wl[300] vdd gnd cell_6t
Xbit_r301_c119 bl[119] br[119] wl[301] vdd gnd cell_6t
Xbit_r302_c119 bl[119] br[119] wl[302] vdd gnd cell_6t
Xbit_r303_c119 bl[119] br[119] wl[303] vdd gnd cell_6t
Xbit_r304_c119 bl[119] br[119] wl[304] vdd gnd cell_6t
Xbit_r305_c119 bl[119] br[119] wl[305] vdd gnd cell_6t
Xbit_r306_c119 bl[119] br[119] wl[306] vdd gnd cell_6t
Xbit_r307_c119 bl[119] br[119] wl[307] vdd gnd cell_6t
Xbit_r308_c119 bl[119] br[119] wl[308] vdd gnd cell_6t
Xbit_r309_c119 bl[119] br[119] wl[309] vdd gnd cell_6t
Xbit_r310_c119 bl[119] br[119] wl[310] vdd gnd cell_6t
Xbit_r311_c119 bl[119] br[119] wl[311] vdd gnd cell_6t
Xbit_r312_c119 bl[119] br[119] wl[312] vdd gnd cell_6t
Xbit_r313_c119 bl[119] br[119] wl[313] vdd gnd cell_6t
Xbit_r314_c119 bl[119] br[119] wl[314] vdd gnd cell_6t
Xbit_r315_c119 bl[119] br[119] wl[315] vdd gnd cell_6t
Xbit_r316_c119 bl[119] br[119] wl[316] vdd gnd cell_6t
Xbit_r317_c119 bl[119] br[119] wl[317] vdd gnd cell_6t
Xbit_r318_c119 bl[119] br[119] wl[318] vdd gnd cell_6t
Xbit_r319_c119 bl[119] br[119] wl[319] vdd gnd cell_6t
Xbit_r320_c119 bl[119] br[119] wl[320] vdd gnd cell_6t
Xbit_r321_c119 bl[119] br[119] wl[321] vdd gnd cell_6t
Xbit_r322_c119 bl[119] br[119] wl[322] vdd gnd cell_6t
Xbit_r323_c119 bl[119] br[119] wl[323] vdd gnd cell_6t
Xbit_r324_c119 bl[119] br[119] wl[324] vdd gnd cell_6t
Xbit_r325_c119 bl[119] br[119] wl[325] vdd gnd cell_6t
Xbit_r326_c119 bl[119] br[119] wl[326] vdd gnd cell_6t
Xbit_r327_c119 bl[119] br[119] wl[327] vdd gnd cell_6t
Xbit_r328_c119 bl[119] br[119] wl[328] vdd gnd cell_6t
Xbit_r329_c119 bl[119] br[119] wl[329] vdd gnd cell_6t
Xbit_r330_c119 bl[119] br[119] wl[330] vdd gnd cell_6t
Xbit_r331_c119 bl[119] br[119] wl[331] vdd gnd cell_6t
Xbit_r332_c119 bl[119] br[119] wl[332] vdd gnd cell_6t
Xbit_r333_c119 bl[119] br[119] wl[333] vdd gnd cell_6t
Xbit_r334_c119 bl[119] br[119] wl[334] vdd gnd cell_6t
Xbit_r335_c119 bl[119] br[119] wl[335] vdd gnd cell_6t
Xbit_r336_c119 bl[119] br[119] wl[336] vdd gnd cell_6t
Xbit_r337_c119 bl[119] br[119] wl[337] vdd gnd cell_6t
Xbit_r338_c119 bl[119] br[119] wl[338] vdd gnd cell_6t
Xbit_r339_c119 bl[119] br[119] wl[339] vdd gnd cell_6t
Xbit_r340_c119 bl[119] br[119] wl[340] vdd gnd cell_6t
Xbit_r341_c119 bl[119] br[119] wl[341] vdd gnd cell_6t
Xbit_r342_c119 bl[119] br[119] wl[342] vdd gnd cell_6t
Xbit_r343_c119 bl[119] br[119] wl[343] vdd gnd cell_6t
Xbit_r344_c119 bl[119] br[119] wl[344] vdd gnd cell_6t
Xbit_r345_c119 bl[119] br[119] wl[345] vdd gnd cell_6t
Xbit_r346_c119 bl[119] br[119] wl[346] vdd gnd cell_6t
Xbit_r347_c119 bl[119] br[119] wl[347] vdd gnd cell_6t
Xbit_r348_c119 bl[119] br[119] wl[348] vdd gnd cell_6t
Xbit_r349_c119 bl[119] br[119] wl[349] vdd gnd cell_6t
Xbit_r350_c119 bl[119] br[119] wl[350] vdd gnd cell_6t
Xbit_r351_c119 bl[119] br[119] wl[351] vdd gnd cell_6t
Xbit_r352_c119 bl[119] br[119] wl[352] vdd gnd cell_6t
Xbit_r353_c119 bl[119] br[119] wl[353] vdd gnd cell_6t
Xbit_r354_c119 bl[119] br[119] wl[354] vdd gnd cell_6t
Xbit_r355_c119 bl[119] br[119] wl[355] vdd gnd cell_6t
Xbit_r356_c119 bl[119] br[119] wl[356] vdd gnd cell_6t
Xbit_r357_c119 bl[119] br[119] wl[357] vdd gnd cell_6t
Xbit_r358_c119 bl[119] br[119] wl[358] vdd gnd cell_6t
Xbit_r359_c119 bl[119] br[119] wl[359] vdd gnd cell_6t
Xbit_r360_c119 bl[119] br[119] wl[360] vdd gnd cell_6t
Xbit_r361_c119 bl[119] br[119] wl[361] vdd gnd cell_6t
Xbit_r362_c119 bl[119] br[119] wl[362] vdd gnd cell_6t
Xbit_r363_c119 bl[119] br[119] wl[363] vdd gnd cell_6t
Xbit_r364_c119 bl[119] br[119] wl[364] vdd gnd cell_6t
Xbit_r365_c119 bl[119] br[119] wl[365] vdd gnd cell_6t
Xbit_r366_c119 bl[119] br[119] wl[366] vdd gnd cell_6t
Xbit_r367_c119 bl[119] br[119] wl[367] vdd gnd cell_6t
Xbit_r368_c119 bl[119] br[119] wl[368] vdd gnd cell_6t
Xbit_r369_c119 bl[119] br[119] wl[369] vdd gnd cell_6t
Xbit_r370_c119 bl[119] br[119] wl[370] vdd gnd cell_6t
Xbit_r371_c119 bl[119] br[119] wl[371] vdd gnd cell_6t
Xbit_r372_c119 bl[119] br[119] wl[372] vdd gnd cell_6t
Xbit_r373_c119 bl[119] br[119] wl[373] vdd gnd cell_6t
Xbit_r374_c119 bl[119] br[119] wl[374] vdd gnd cell_6t
Xbit_r375_c119 bl[119] br[119] wl[375] vdd gnd cell_6t
Xbit_r376_c119 bl[119] br[119] wl[376] vdd gnd cell_6t
Xbit_r377_c119 bl[119] br[119] wl[377] vdd gnd cell_6t
Xbit_r378_c119 bl[119] br[119] wl[378] vdd gnd cell_6t
Xbit_r379_c119 bl[119] br[119] wl[379] vdd gnd cell_6t
Xbit_r380_c119 bl[119] br[119] wl[380] vdd gnd cell_6t
Xbit_r381_c119 bl[119] br[119] wl[381] vdd gnd cell_6t
Xbit_r382_c119 bl[119] br[119] wl[382] vdd gnd cell_6t
Xbit_r383_c119 bl[119] br[119] wl[383] vdd gnd cell_6t
Xbit_r384_c119 bl[119] br[119] wl[384] vdd gnd cell_6t
Xbit_r385_c119 bl[119] br[119] wl[385] vdd gnd cell_6t
Xbit_r386_c119 bl[119] br[119] wl[386] vdd gnd cell_6t
Xbit_r387_c119 bl[119] br[119] wl[387] vdd gnd cell_6t
Xbit_r388_c119 bl[119] br[119] wl[388] vdd gnd cell_6t
Xbit_r389_c119 bl[119] br[119] wl[389] vdd gnd cell_6t
Xbit_r390_c119 bl[119] br[119] wl[390] vdd gnd cell_6t
Xbit_r391_c119 bl[119] br[119] wl[391] vdd gnd cell_6t
Xbit_r392_c119 bl[119] br[119] wl[392] vdd gnd cell_6t
Xbit_r393_c119 bl[119] br[119] wl[393] vdd gnd cell_6t
Xbit_r394_c119 bl[119] br[119] wl[394] vdd gnd cell_6t
Xbit_r395_c119 bl[119] br[119] wl[395] vdd gnd cell_6t
Xbit_r396_c119 bl[119] br[119] wl[396] vdd gnd cell_6t
Xbit_r397_c119 bl[119] br[119] wl[397] vdd gnd cell_6t
Xbit_r398_c119 bl[119] br[119] wl[398] vdd gnd cell_6t
Xbit_r399_c119 bl[119] br[119] wl[399] vdd gnd cell_6t
Xbit_r400_c119 bl[119] br[119] wl[400] vdd gnd cell_6t
Xbit_r401_c119 bl[119] br[119] wl[401] vdd gnd cell_6t
Xbit_r402_c119 bl[119] br[119] wl[402] vdd gnd cell_6t
Xbit_r403_c119 bl[119] br[119] wl[403] vdd gnd cell_6t
Xbit_r404_c119 bl[119] br[119] wl[404] vdd gnd cell_6t
Xbit_r405_c119 bl[119] br[119] wl[405] vdd gnd cell_6t
Xbit_r406_c119 bl[119] br[119] wl[406] vdd gnd cell_6t
Xbit_r407_c119 bl[119] br[119] wl[407] vdd gnd cell_6t
Xbit_r408_c119 bl[119] br[119] wl[408] vdd gnd cell_6t
Xbit_r409_c119 bl[119] br[119] wl[409] vdd gnd cell_6t
Xbit_r410_c119 bl[119] br[119] wl[410] vdd gnd cell_6t
Xbit_r411_c119 bl[119] br[119] wl[411] vdd gnd cell_6t
Xbit_r412_c119 bl[119] br[119] wl[412] vdd gnd cell_6t
Xbit_r413_c119 bl[119] br[119] wl[413] vdd gnd cell_6t
Xbit_r414_c119 bl[119] br[119] wl[414] vdd gnd cell_6t
Xbit_r415_c119 bl[119] br[119] wl[415] vdd gnd cell_6t
Xbit_r416_c119 bl[119] br[119] wl[416] vdd gnd cell_6t
Xbit_r417_c119 bl[119] br[119] wl[417] vdd gnd cell_6t
Xbit_r418_c119 bl[119] br[119] wl[418] vdd gnd cell_6t
Xbit_r419_c119 bl[119] br[119] wl[419] vdd gnd cell_6t
Xbit_r420_c119 bl[119] br[119] wl[420] vdd gnd cell_6t
Xbit_r421_c119 bl[119] br[119] wl[421] vdd gnd cell_6t
Xbit_r422_c119 bl[119] br[119] wl[422] vdd gnd cell_6t
Xbit_r423_c119 bl[119] br[119] wl[423] vdd gnd cell_6t
Xbit_r424_c119 bl[119] br[119] wl[424] vdd gnd cell_6t
Xbit_r425_c119 bl[119] br[119] wl[425] vdd gnd cell_6t
Xbit_r426_c119 bl[119] br[119] wl[426] vdd gnd cell_6t
Xbit_r427_c119 bl[119] br[119] wl[427] vdd gnd cell_6t
Xbit_r428_c119 bl[119] br[119] wl[428] vdd gnd cell_6t
Xbit_r429_c119 bl[119] br[119] wl[429] vdd gnd cell_6t
Xbit_r430_c119 bl[119] br[119] wl[430] vdd gnd cell_6t
Xbit_r431_c119 bl[119] br[119] wl[431] vdd gnd cell_6t
Xbit_r432_c119 bl[119] br[119] wl[432] vdd gnd cell_6t
Xbit_r433_c119 bl[119] br[119] wl[433] vdd gnd cell_6t
Xbit_r434_c119 bl[119] br[119] wl[434] vdd gnd cell_6t
Xbit_r435_c119 bl[119] br[119] wl[435] vdd gnd cell_6t
Xbit_r436_c119 bl[119] br[119] wl[436] vdd gnd cell_6t
Xbit_r437_c119 bl[119] br[119] wl[437] vdd gnd cell_6t
Xbit_r438_c119 bl[119] br[119] wl[438] vdd gnd cell_6t
Xbit_r439_c119 bl[119] br[119] wl[439] vdd gnd cell_6t
Xbit_r440_c119 bl[119] br[119] wl[440] vdd gnd cell_6t
Xbit_r441_c119 bl[119] br[119] wl[441] vdd gnd cell_6t
Xbit_r442_c119 bl[119] br[119] wl[442] vdd gnd cell_6t
Xbit_r443_c119 bl[119] br[119] wl[443] vdd gnd cell_6t
Xbit_r444_c119 bl[119] br[119] wl[444] vdd gnd cell_6t
Xbit_r445_c119 bl[119] br[119] wl[445] vdd gnd cell_6t
Xbit_r446_c119 bl[119] br[119] wl[446] vdd gnd cell_6t
Xbit_r447_c119 bl[119] br[119] wl[447] vdd gnd cell_6t
Xbit_r448_c119 bl[119] br[119] wl[448] vdd gnd cell_6t
Xbit_r449_c119 bl[119] br[119] wl[449] vdd gnd cell_6t
Xbit_r450_c119 bl[119] br[119] wl[450] vdd gnd cell_6t
Xbit_r451_c119 bl[119] br[119] wl[451] vdd gnd cell_6t
Xbit_r452_c119 bl[119] br[119] wl[452] vdd gnd cell_6t
Xbit_r453_c119 bl[119] br[119] wl[453] vdd gnd cell_6t
Xbit_r454_c119 bl[119] br[119] wl[454] vdd gnd cell_6t
Xbit_r455_c119 bl[119] br[119] wl[455] vdd gnd cell_6t
Xbit_r456_c119 bl[119] br[119] wl[456] vdd gnd cell_6t
Xbit_r457_c119 bl[119] br[119] wl[457] vdd gnd cell_6t
Xbit_r458_c119 bl[119] br[119] wl[458] vdd gnd cell_6t
Xbit_r459_c119 bl[119] br[119] wl[459] vdd gnd cell_6t
Xbit_r460_c119 bl[119] br[119] wl[460] vdd gnd cell_6t
Xbit_r461_c119 bl[119] br[119] wl[461] vdd gnd cell_6t
Xbit_r462_c119 bl[119] br[119] wl[462] vdd gnd cell_6t
Xbit_r463_c119 bl[119] br[119] wl[463] vdd gnd cell_6t
Xbit_r464_c119 bl[119] br[119] wl[464] vdd gnd cell_6t
Xbit_r465_c119 bl[119] br[119] wl[465] vdd gnd cell_6t
Xbit_r466_c119 bl[119] br[119] wl[466] vdd gnd cell_6t
Xbit_r467_c119 bl[119] br[119] wl[467] vdd gnd cell_6t
Xbit_r468_c119 bl[119] br[119] wl[468] vdd gnd cell_6t
Xbit_r469_c119 bl[119] br[119] wl[469] vdd gnd cell_6t
Xbit_r470_c119 bl[119] br[119] wl[470] vdd gnd cell_6t
Xbit_r471_c119 bl[119] br[119] wl[471] vdd gnd cell_6t
Xbit_r472_c119 bl[119] br[119] wl[472] vdd gnd cell_6t
Xbit_r473_c119 bl[119] br[119] wl[473] vdd gnd cell_6t
Xbit_r474_c119 bl[119] br[119] wl[474] vdd gnd cell_6t
Xbit_r475_c119 bl[119] br[119] wl[475] vdd gnd cell_6t
Xbit_r476_c119 bl[119] br[119] wl[476] vdd gnd cell_6t
Xbit_r477_c119 bl[119] br[119] wl[477] vdd gnd cell_6t
Xbit_r478_c119 bl[119] br[119] wl[478] vdd gnd cell_6t
Xbit_r479_c119 bl[119] br[119] wl[479] vdd gnd cell_6t
Xbit_r480_c119 bl[119] br[119] wl[480] vdd gnd cell_6t
Xbit_r481_c119 bl[119] br[119] wl[481] vdd gnd cell_6t
Xbit_r482_c119 bl[119] br[119] wl[482] vdd gnd cell_6t
Xbit_r483_c119 bl[119] br[119] wl[483] vdd gnd cell_6t
Xbit_r484_c119 bl[119] br[119] wl[484] vdd gnd cell_6t
Xbit_r485_c119 bl[119] br[119] wl[485] vdd gnd cell_6t
Xbit_r486_c119 bl[119] br[119] wl[486] vdd gnd cell_6t
Xbit_r487_c119 bl[119] br[119] wl[487] vdd gnd cell_6t
Xbit_r488_c119 bl[119] br[119] wl[488] vdd gnd cell_6t
Xbit_r489_c119 bl[119] br[119] wl[489] vdd gnd cell_6t
Xbit_r490_c119 bl[119] br[119] wl[490] vdd gnd cell_6t
Xbit_r491_c119 bl[119] br[119] wl[491] vdd gnd cell_6t
Xbit_r492_c119 bl[119] br[119] wl[492] vdd gnd cell_6t
Xbit_r493_c119 bl[119] br[119] wl[493] vdd gnd cell_6t
Xbit_r494_c119 bl[119] br[119] wl[494] vdd gnd cell_6t
Xbit_r495_c119 bl[119] br[119] wl[495] vdd gnd cell_6t
Xbit_r496_c119 bl[119] br[119] wl[496] vdd gnd cell_6t
Xbit_r497_c119 bl[119] br[119] wl[497] vdd gnd cell_6t
Xbit_r498_c119 bl[119] br[119] wl[498] vdd gnd cell_6t
Xbit_r499_c119 bl[119] br[119] wl[499] vdd gnd cell_6t
Xbit_r500_c119 bl[119] br[119] wl[500] vdd gnd cell_6t
Xbit_r501_c119 bl[119] br[119] wl[501] vdd gnd cell_6t
Xbit_r502_c119 bl[119] br[119] wl[502] vdd gnd cell_6t
Xbit_r503_c119 bl[119] br[119] wl[503] vdd gnd cell_6t
Xbit_r504_c119 bl[119] br[119] wl[504] vdd gnd cell_6t
Xbit_r505_c119 bl[119] br[119] wl[505] vdd gnd cell_6t
Xbit_r506_c119 bl[119] br[119] wl[506] vdd gnd cell_6t
Xbit_r507_c119 bl[119] br[119] wl[507] vdd gnd cell_6t
Xbit_r508_c119 bl[119] br[119] wl[508] vdd gnd cell_6t
Xbit_r509_c119 bl[119] br[119] wl[509] vdd gnd cell_6t
Xbit_r510_c119 bl[119] br[119] wl[510] vdd gnd cell_6t
Xbit_r511_c119 bl[119] br[119] wl[511] vdd gnd cell_6t
Xbit_r0_c120 bl[120] br[120] wl[0] vdd gnd cell_6t
Xbit_r1_c120 bl[120] br[120] wl[1] vdd gnd cell_6t
Xbit_r2_c120 bl[120] br[120] wl[2] vdd gnd cell_6t
Xbit_r3_c120 bl[120] br[120] wl[3] vdd gnd cell_6t
Xbit_r4_c120 bl[120] br[120] wl[4] vdd gnd cell_6t
Xbit_r5_c120 bl[120] br[120] wl[5] vdd gnd cell_6t
Xbit_r6_c120 bl[120] br[120] wl[6] vdd gnd cell_6t
Xbit_r7_c120 bl[120] br[120] wl[7] vdd gnd cell_6t
Xbit_r8_c120 bl[120] br[120] wl[8] vdd gnd cell_6t
Xbit_r9_c120 bl[120] br[120] wl[9] vdd gnd cell_6t
Xbit_r10_c120 bl[120] br[120] wl[10] vdd gnd cell_6t
Xbit_r11_c120 bl[120] br[120] wl[11] vdd gnd cell_6t
Xbit_r12_c120 bl[120] br[120] wl[12] vdd gnd cell_6t
Xbit_r13_c120 bl[120] br[120] wl[13] vdd gnd cell_6t
Xbit_r14_c120 bl[120] br[120] wl[14] vdd gnd cell_6t
Xbit_r15_c120 bl[120] br[120] wl[15] vdd gnd cell_6t
Xbit_r16_c120 bl[120] br[120] wl[16] vdd gnd cell_6t
Xbit_r17_c120 bl[120] br[120] wl[17] vdd gnd cell_6t
Xbit_r18_c120 bl[120] br[120] wl[18] vdd gnd cell_6t
Xbit_r19_c120 bl[120] br[120] wl[19] vdd gnd cell_6t
Xbit_r20_c120 bl[120] br[120] wl[20] vdd gnd cell_6t
Xbit_r21_c120 bl[120] br[120] wl[21] vdd gnd cell_6t
Xbit_r22_c120 bl[120] br[120] wl[22] vdd gnd cell_6t
Xbit_r23_c120 bl[120] br[120] wl[23] vdd gnd cell_6t
Xbit_r24_c120 bl[120] br[120] wl[24] vdd gnd cell_6t
Xbit_r25_c120 bl[120] br[120] wl[25] vdd gnd cell_6t
Xbit_r26_c120 bl[120] br[120] wl[26] vdd gnd cell_6t
Xbit_r27_c120 bl[120] br[120] wl[27] vdd gnd cell_6t
Xbit_r28_c120 bl[120] br[120] wl[28] vdd gnd cell_6t
Xbit_r29_c120 bl[120] br[120] wl[29] vdd gnd cell_6t
Xbit_r30_c120 bl[120] br[120] wl[30] vdd gnd cell_6t
Xbit_r31_c120 bl[120] br[120] wl[31] vdd gnd cell_6t
Xbit_r32_c120 bl[120] br[120] wl[32] vdd gnd cell_6t
Xbit_r33_c120 bl[120] br[120] wl[33] vdd gnd cell_6t
Xbit_r34_c120 bl[120] br[120] wl[34] vdd gnd cell_6t
Xbit_r35_c120 bl[120] br[120] wl[35] vdd gnd cell_6t
Xbit_r36_c120 bl[120] br[120] wl[36] vdd gnd cell_6t
Xbit_r37_c120 bl[120] br[120] wl[37] vdd gnd cell_6t
Xbit_r38_c120 bl[120] br[120] wl[38] vdd gnd cell_6t
Xbit_r39_c120 bl[120] br[120] wl[39] vdd gnd cell_6t
Xbit_r40_c120 bl[120] br[120] wl[40] vdd gnd cell_6t
Xbit_r41_c120 bl[120] br[120] wl[41] vdd gnd cell_6t
Xbit_r42_c120 bl[120] br[120] wl[42] vdd gnd cell_6t
Xbit_r43_c120 bl[120] br[120] wl[43] vdd gnd cell_6t
Xbit_r44_c120 bl[120] br[120] wl[44] vdd gnd cell_6t
Xbit_r45_c120 bl[120] br[120] wl[45] vdd gnd cell_6t
Xbit_r46_c120 bl[120] br[120] wl[46] vdd gnd cell_6t
Xbit_r47_c120 bl[120] br[120] wl[47] vdd gnd cell_6t
Xbit_r48_c120 bl[120] br[120] wl[48] vdd gnd cell_6t
Xbit_r49_c120 bl[120] br[120] wl[49] vdd gnd cell_6t
Xbit_r50_c120 bl[120] br[120] wl[50] vdd gnd cell_6t
Xbit_r51_c120 bl[120] br[120] wl[51] vdd gnd cell_6t
Xbit_r52_c120 bl[120] br[120] wl[52] vdd gnd cell_6t
Xbit_r53_c120 bl[120] br[120] wl[53] vdd gnd cell_6t
Xbit_r54_c120 bl[120] br[120] wl[54] vdd gnd cell_6t
Xbit_r55_c120 bl[120] br[120] wl[55] vdd gnd cell_6t
Xbit_r56_c120 bl[120] br[120] wl[56] vdd gnd cell_6t
Xbit_r57_c120 bl[120] br[120] wl[57] vdd gnd cell_6t
Xbit_r58_c120 bl[120] br[120] wl[58] vdd gnd cell_6t
Xbit_r59_c120 bl[120] br[120] wl[59] vdd gnd cell_6t
Xbit_r60_c120 bl[120] br[120] wl[60] vdd gnd cell_6t
Xbit_r61_c120 bl[120] br[120] wl[61] vdd gnd cell_6t
Xbit_r62_c120 bl[120] br[120] wl[62] vdd gnd cell_6t
Xbit_r63_c120 bl[120] br[120] wl[63] vdd gnd cell_6t
Xbit_r64_c120 bl[120] br[120] wl[64] vdd gnd cell_6t
Xbit_r65_c120 bl[120] br[120] wl[65] vdd gnd cell_6t
Xbit_r66_c120 bl[120] br[120] wl[66] vdd gnd cell_6t
Xbit_r67_c120 bl[120] br[120] wl[67] vdd gnd cell_6t
Xbit_r68_c120 bl[120] br[120] wl[68] vdd gnd cell_6t
Xbit_r69_c120 bl[120] br[120] wl[69] vdd gnd cell_6t
Xbit_r70_c120 bl[120] br[120] wl[70] vdd gnd cell_6t
Xbit_r71_c120 bl[120] br[120] wl[71] vdd gnd cell_6t
Xbit_r72_c120 bl[120] br[120] wl[72] vdd gnd cell_6t
Xbit_r73_c120 bl[120] br[120] wl[73] vdd gnd cell_6t
Xbit_r74_c120 bl[120] br[120] wl[74] vdd gnd cell_6t
Xbit_r75_c120 bl[120] br[120] wl[75] vdd gnd cell_6t
Xbit_r76_c120 bl[120] br[120] wl[76] vdd gnd cell_6t
Xbit_r77_c120 bl[120] br[120] wl[77] vdd gnd cell_6t
Xbit_r78_c120 bl[120] br[120] wl[78] vdd gnd cell_6t
Xbit_r79_c120 bl[120] br[120] wl[79] vdd gnd cell_6t
Xbit_r80_c120 bl[120] br[120] wl[80] vdd gnd cell_6t
Xbit_r81_c120 bl[120] br[120] wl[81] vdd gnd cell_6t
Xbit_r82_c120 bl[120] br[120] wl[82] vdd gnd cell_6t
Xbit_r83_c120 bl[120] br[120] wl[83] vdd gnd cell_6t
Xbit_r84_c120 bl[120] br[120] wl[84] vdd gnd cell_6t
Xbit_r85_c120 bl[120] br[120] wl[85] vdd gnd cell_6t
Xbit_r86_c120 bl[120] br[120] wl[86] vdd gnd cell_6t
Xbit_r87_c120 bl[120] br[120] wl[87] vdd gnd cell_6t
Xbit_r88_c120 bl[120] br[120] wl[88] vdd gnd cell_6t
Xbit_r89_c120 bl[120] br[120] wl[89] vdd gnd cell_6t
Xbit_r90_c120 bl[120] br[120] wl[90] vdd gnd cell_6t
Xbit_r91_c120 bl[120] br[120] wl[91] vdd gnd cell_6t
Xbit_r92_c120 bl[120] br[120] wl[92] vdd gnd cell_6t
Xbit_r93_c120 bl[120] br[120] wl[93] vdd gnd cell_6t
Xbit_r94_c120 bl[120] br[120] wl[94] vdd gnd cell_6t
Xbit_r95_c120 bl[120] br[120] wl[95] vdd gnd cell_6t
Xbit_r96_c120 bl[120] br[120] wl[96] vdd gnd cell_6t
Xbit_r97_c120 bl[120] br[120] wl[97] vdd gnd cell_6t
Xbit_r98_c120 bl[120] br[120] wl[98] vdd gnd cell_6t
Xbit_r99_c120 bl[120] br[120] wl[99] vdd gnd cell_6t
Xbit_r100_c120 bl[120] br[120] wl[100] vdd gnd cell_6t
Xbit_r101_c120 bl[120] br[120] wl[101] vdd gnd cell_6t
Xbit_r102_c120 bl[120] br[120] wl[102] vdd gnd cell_6t
Xbit_r103_c120 bl[120] br[120] wl[103] vdd gnd cell_6t
Xbit_r104_c120 bl[120] br[120] wl[104] vdd gnd cell_6t
Xbit_r105_c120 bl[120] br[120] wl[105] vdd gnd cell_6t
Xbit_r106_c120 bl[120] br[120] wl[106] vdd gnd cell_6t
Xbit_r107_c120 bl[120] br[120] wl[107] vdd gnd cell_6t
Xbit_r108_c120 bl[120] br[120] wl[108] vdd gnd cell_6t
Xbit_r109_c120 bl[120] br[120] wl[109] vdd gnd cell_6t
Xbit_r110_c120 bl[120] br[120] wl[110] vdd gnd cell_6t
Xbit_r111_c120 bl[120] br[120] wl[111] vdd gnd cell_6t
Xbit_r112_c120 bl[120] br[120] wl[112] vdd gnd cell_6t
Xbit_r113_c120 bl[120] br[120] wl[113] vdd gnd cell_6t
Xbit_r114_c120 bl[120] br[120] wl[114] vdd gnd cell_6t
Xbit_r115_c120 bl[120] br[120] wl[115] vdd gnd cell_6t
Xbit_r116_c120 bl[120] br[120] wl[116] vdd gnd cell_6t
Xbit_r117_c120 bl[120] br[120] wl[117] vdd gnd cell_6t
Xbit_r118_c120 bl[120] br[120] wl[118] vdd gnd cell_6t
Xbit_r119_c120 bl[120] br[120] wl[119] vdd gnd cell_6t
Xbit_r120_c120 bl[120] br[120] wl[120] vdd gnd cell_6t
Xbit_r121_c120 bl[120] br[120] wl[121] vdd gnd cell_6t
Xbit_r122_c120 bl[120] br[120] wl[122] vdd gnd cell_6t
Xbit_r123_c120 bl[120] br[120] wl[123] vdd gnd cell_6t
Xbit_r124_c120 bl[120] br[120] wl[124] vdd gnd cell_6t
Xbit_r125_c120 bl[120] br[120] wl[125] vdd gnd cell_6t
Xbit_r126_c120 bl[120] br[120] wl[126] vdd gnd cell_6t
Xbit_r127_c120 bl[120] br[120] wl[127] vdd gnd cell_6t
Xbit_r128_c120 bl[120] br[120] wl[128] vdd gnd cell_6t
Xbit_r129_c120 bl[120] br[120] wl[129] vdd gnd cell_6t
Xbit_r130_c120 bl[120] br[120] wl[130] vdd gnd cell_6t
Xbit_r131_c120 bl[120] br[120] wl[131] vdd gnd cell_6t
Xbit_r132_c120 bl[120] br[120] wl[132] vdd gnd cell_6t
Xbit_r133_c120 bl[120] br[120] wl[133] vdd gnd cell_6t
Xbit_r134_c120 bl[120] br[120] wl[134] vdd gnd cell_6t
Xbit_r135_c120 bl[120] br[120] wl[135] vdd gnd cell_6t
Xbit_r136_c120 bl[120] br[120] wl[136] vdd gnd cell_6t
Xbit_r137_c120 bl[120] br[120] wl[137] vdd gnd cell_6t
Xbit_r138_c120 bl[120] br[120] wl[138] vdd gnd cell_6t
Xbit_r139_c120 bl[120] br[120] wl[139] vdd gnd cell_6t
Xbit_r140_c120 bl[120] br[120] wl[140] vdd gnd cell_6t
Xbit_r141_c120 bl[120] br[120] wl[141] vdd gnd cell_6t
Xbit_r142_c120 bl[120] br[120] wl[142] vdd gnd cell_6t
Xbit_r143_c120 bl[120] br[120] wl[143] vdd gnd cell_6t
Xbit_r144_c120 bl[120] br[120] wl[144] vdd gnd cell_6t
Xbit_r145_c120 bl[120] br[120] wl[145] vdd gnd cell_6t
Xbit_r146_c120 bl[120] br[120] wl[146] vdd gnd cell_6t
Xbit_r147_c120 bl[120] br[120] wl[147] vdd gnd cell_6t
Xbit_r148_c120 bl[120] br[120] wl[148] vdd gnd cell_6t
Xbit_r149_c120 bl[120] br[120] wl[149] vdd gnd cell_6t
Xbit_r150_c120 bl[120] br[120] wl[150] vdd gnd cell_6t
Xbit_r151_c120 bl[120] br[120] wl[151] vdd gnd cell_6t
Xbit_r152_c120 bl[120] br[120] wl[152] vdd gnd cell_6t
Xbit_r153_c120 bl[120] br[120] wl[153] vdd gnd cell_6t
Xbit_r154_c120 bl[120] br[120] wl[154] vdd gnd cell_6t
Xbit_r155_c120 bl[120] br[120] wl[155] vdd gnd cell_6t
Xbit_r156_c120 bl[120] br[120] wl[156] vdd gnd cell_6t
Xbit_r157_c120 bl[120] br[120] wl[157] vdd gnd cell_6t
Xbit_r158_c120 bl[120] br[120] wl[158] vdd gnd cell_6t
Xbit_r159_c120 bl[120] br[120] wl[159] vdd gnd cell_6t
Xbit_r160_c120 bl[120] br[120] wl[160] vdd gnd cell_6t
Xbit_r161_c120 bl[120] br[120] wl[161] vdd gnd cell_6t
Xbit_r162_c120 bl[120] br[120] wl[162] vdd gnd cell_6t
Xbit_r163_c120 bl[120] br[120] wl[163] vdd gnd cell_6t
Xbit_r164_c120 bl[120] br[120] wl[164] vdd gnd cell_6t
Xbit_r165_c120 bl[120] br[120] wl[165] vdd gnd cell_6t
Xbit_r166_c120 bl[120] br[120] wl[166] vdd gnd cell_6t
Xbit_r167_c120 bl[120] br[120] wl[167] vdd gnd cell_6t
Xbit_r168_c120 bl[120] br[120] wl[168] vdd gnd cell_6t
Xbit_r169_c120 bl[120] br[120] wl[169] vdd gnd cell_6t
Xbit_r170_c120 bl[120] br[120] wl[170] vdd gnd cell_6t
Xbit_r171_c120 bl[120] br[120] wl[171] vdd gnd cell_6t
Xbit_r172_c120 bl[120] br[120] wl[172] vdd gnd cell_6t
Xbit_r173_c120 bl[120] br[120] wl[173] vdd gnd cell_6t
Xbit_r174_c120 bl[120] br[120] wl[174] vdd gnd cell_6t
Xbit_r175_c120 bl[120] br[120] wl[175] vdd gnd cell_6t
Xbit_r176_c120 bl[120] br[120] wl[176] vdd gnd cell_6t
Xbit_r177_c120 bl[120] br[120] wl[177] vdd gnd cell_6t
Xbit_r178_c120 bl[120] br[120] wl[178] vdd gnd cell_6t
Xbit_r179_c120 bl[120] br[120] wl[179] vdd gnd cell_6t
Xbit_r180_c120 bl[120] br[120] wl[180] vdd gnd cell_6t
Xbit_r181_c120 bl[120] br[120] wl[181] vdd gnd cell_6t
Xbit_r182_c120 bl[120] br[120] wl[182] vdd gnd cell_6t
Xbit_r183_c120 bl[120] br[120] wl[183] vdd gnd cell_6t
Xbit_r184_c120 bl[120] br[120] wl[184] vdd gnd cell_6t
Xbit_r185_c120 bl[120] br[120] wl[185] vdd gnd cell_6t
Xbit_r186_c120 bl[120] br[120] wl[186] vdd gnd cell_6t
Xbit_r187_c120 bl[120] br[120] wl[187] vdd gnd cell_6t
Xbit_r188_c120 bl[120] br[120] wl[188] vdd gnd cell_6t
Xbit_r189_c120 bl[120] br[120] wl[189] vdd gnd cell_6t
Xbit_r190_c120 bl[120] br[120] wl[190] vdd gnd cell_6t
Xbit_r191_c120 bl[120] br[120] wl[191] vdd gnd cell_6t
Xbit_r192_c120 bl[120] br[120] wl[192] vdd gnd cell_6t
Xbit_r193_c120 bl[120] br[120] wl[193] vdd gnd cell_6t
Xbit_r194_c120 bl[120] br[120] wl[194] vdd gnd cell_6t
Xbit_r195_c120 bl[120] br[120] wl[195] vdd gnd cell_6t
Xbit_r196_c120 bl[120] br[120] wl[196] vdd gnd cell_6t
Xbit_r197_c120 bl[120] br[120] wl[197] vdd gnd cell_6t
Xbit_r198_c120 bl[120] br[120] wl[198] vdd gnd cell_6t
Xbit_r199_c120 bl[120] br[120] wl[199] vdd gnd cell_6t
Xbit_r200_c120 bl[120] br[120] wl[200] vdd gnd cell_6t
Xbit_r201_c120 bl[120] br[120] wl[201] vdd gnd cell_6t
Xbit_r202_c120 bl[120] br[120] wl[202] vdd gnd cell_6t
Xbit_r203_c120 bl[120] br[120] wl[203] vdd gnd cell_6t
Xbit_r204_c120 bl[120] br[120] wl[204] vdd gnd cell_6t
Xbit_r205_c120 bl[120] br[120] wl[205] vdd gnd cell_6t
Xbit_r206_c120 bl[120] br[120] wl[206] vdd gnd cell_6t
Xbit_r207_c120 bl[120] br[120] wl[207] vdd gnd cell_6t
Xbit_r208_c120 bl[120] br[120] wl[208] vdd gnd cell_6t
Xbit_r209_c120 bl[120] br[120] wl[209] vdd gnd cell_6t
Xbit_r210_c120 bl[120] br[120] wl[210] vdd gnd cell_6t
Xbit_r211_c120 bl[120] br[120] wl[211] vdd gnd cell_6t
Xbit_r212_c120 bl[120] br[120] wl[212] vdd gnd cell_6t
Xbit_r213_c120 bl[120] br[120] wl[213] vdd gnd cell_6t
Xbit_r214_c120 bl[120] br[120] wl[214] vdd gnd cell_6t
Xbit_r215_c120 bl[120] br[120] wl[215] vdd gnd cell_6t
Xbit_r216_c120 bl[120] br[120] wl[216] vdd gnd cell_6t
Xbit_r217_c120 bl[120] br[120] wl[217] vdd gnd cell_6t
Xbit_r218_c120 bl[120] br[120] wl[218] vdd gnd cell_6t
Xbit_r219_c120 bl[120] br[120] wl[219] vdd gnd cell_6t
Xbit_r220_c120 bl[120] br[120] wl[220] vdd gnd cell_6t
Xbit_r221_c120 bl[120] br[120] wl[221] vdd gnd cell_6t
Xbit_r222_c120 bl[120] br[120] wl[222] vdd gnd cell_6t
Xbit_r223_c120 bl[120] br[120] wl[223] vdd gnd cell_6t
Xbit_r224_c120 bl[120] br[120] wl[224] vdd gnd cell_6t
Xbit_r225_c120 bl[120] br[120] wl[225] vdd gnd cell_6t
Xbit_r226_c120 bl[120] br[120] wl[226] vdd gnd cell_6t
Xbit_r227_c120 bl[120] br[120] wl[227] vdd gnd cell_6t
Xbit_r228_c120 bl[120] br[120] wl[228] vdd gnd cell_6t
Xbit_r229_c120 bl[120] br[120] wl[229] vdd gnd cell_6t
Xbit_r230_c120 bl[120] br[120] wl[230] vdd gnd cell_6t
Xbit_r231_c120 bl[120] br[120] wl[231] vdd gnd cell_6t
Xbit_r232_c120 bl[120] br[120] wl[232] vdd gnd cell_6t
Xbit_r233_c120 bl[120] br[120] wl[233] vdd gnd cell_6t
Xbit_r234_c120 bl[120] br[120] wl[234] vdd gnd cell_6t
Xbit_r235_c120 bl[120] br[120] wl[235] vdd gnd cell_6t
Xbit_r236_c120 bl[120] br[120] wl[236] vdd gnd cell_6t
Xbit_r237_c120 bl[120] br[120] wl[237] vdd gnd cell_6t
Xbit_r238_c120 bl[120] br[120] wl[238] vdd gnd cell_6t
Xbit_r239_c120 bl[120] br[120] wl[239] vdd gnd cell_6t
Xbit_r240_c120 bl[120] br[120] wl[240] vdd gnd cell_6t
Xbit_r241_c120 bl[120] br[120] wl[241] vdd gnd cell_6t
Xbit_r242_c120 bl[120] br[120] wl[242] vdd gnd cell_6t
Xbit_r243_c120 bl[120] br[120] wl[243] vdd gnd cell_6t
Xbit_r244_c120 bl[120] br[120] wl[244] vdd gnd cell_6t
Xbit_r245_c120 bl[120] br[120] wl[245] vdd gnd cell_6t
Xbit_r246_c120 bl[120] br[120] wl[246] vdd gnd cell_6t
Xbit_r247_c120 bl[120] br[120] wl[247] vdd gnd cell_6t
Xbit_r248_c120 bl[120] br[120] wl[248] vdd gnd cell_6t
Xbit_r249_c120 bl[120] br[120] wl[249] vdd gnd cell_6t
Xbit_r250_c120 bl[120] br[120] wl[250] vdd gnd cell_6t
Xbit_r251_c120 bl[120] br[120] wl[251] vdd gnd cell_6t
Xbit_r252_c120 bl[120] br[120] wl[252] vdd gnd cell_6t
Xbit_r253_c120 bl[120] br[120] wl[253] vdd gnd cell_6t
Xbit_r254_c120 bl[120] br[120] wl[254] vdd gnd cell_6t
Xbit_r255_c120 bl[120] br[120] wl[255] vdd gnd cell_6t
Xbit_r256_c120 bl[120] br[120] wl[256] vdd gnd cell_6t
Xbit_r257_c120 bl[120] br[120] wl[257] vdd gnd cell_6t
Xbit_r258_c120 bl[120] br[120] wl[258] vdd gnd cell_6t
Xbit_r259_c120 bl[120] br[120] wl[259] vdd gnd cell_6t
Xbit_r260_c120 bl[120] br[120] wl[260] vdd gnd cell_6t
Xbit_r261_c120 bl[120] br[120] wl[261] vdd gnd cell_6t
Xbit_r262_c120 bl[120] br[120] wl[262] vdd gnd cell_6t
Xbit_r263_c120 bl[120] br[120] wl[263] vdd gnd cell_6t
Xbit_r264_c120 bl[120] br[120] wl[264] vdd gnd cell_6t
Xbit_r265_c120 bl[120] br[120] wl[265] vdd gnd cell_6t
Xbit_r266_c120 bl[120] br[120] wl[266] vdd gnd cell_6t
Xbit_r267_c120 bl[120] br[120] wl[267] vdd gnd cell_6t
Xbit_r268_c120 bl[120] br[120] wl[268] vdd gnd cell_6t
Xbit_r269_c120 bl[120] br[120] wl[269] vdd gnd cell_6t
Xbit_r270_c120 bl[120] br[120] wl[270] vdd gnd cell_6t
Xbit_r271_c120 bl[120] br[120] wl[271] vdd gnd cell_6t
Xbit_r272_c120 bl[120] br[120] wl[272] vdd gnd cell_6t
Xbit_r273_c120 bl[120] br[120] wl[273] vdd gnd cell_6t
Xbit_r274_c120 bl[120] br[120] wl[274] vdd gnd cell_6t
Xbit_r275_c120 bl[120] br[120] wl[275] vdd gnd cell_6t
Xbit_r276_c120 bl[120] br[120] wl[276] vdd gnd cell_6t
Xbit_r277_c120 bl[120] br[120] wl[277] vdd gnd cell_6t
Xbit_r278_c120 bl[120] br[120] wl[278] vdd gnd cell_6t
Xbit_r279_c120 bl[120] br[120] wl[279] vdd gnd cell_6t
Xbit_r280_c120 bl[120] br[120] wl[280] vdd gnd cell_6t
Xbit_r281_c120 bl[120] br[120] wl[281] vdd gnd cell_6t
Xbit_r282_c120 bl[120] br[120] wl[282] vdd gnd cell_6t
Xbit_r283_c120 bl[120] br[120] wl[283] vdd gnd cell_6t
Xbit_r284_c120 bl[120] br[120] wl[284] vdd gnd cell_6t
Xbit_r285_c120 bl[120] br[120] wl[285] vdd gnd cell_6t
Xbit_r286_c120 bl[120] br[120] wl[286] vdd gnd cell_6t
Xbit_r287_c120 bl[120] br[120] wl[287] vdd gnd cell_6t
Xbit_r288_c120 bl[120] br[120] wl[288] vdd gnd cell_6t
Xbit_r289_c120 bl[120] br[120] wl[289] vdd gnd cell_6t
Xbit_r290_c120 bl[120] br[120] wl[290] vdd gnd cell_6t
Xbit_r291_c120 bl[120] br[120] wl[291] vdd gnd cell_6t
Xbit_r292_c120 bl[120] br[120] wl[292] vdd gnd cell_6t
Xbit_r293_c120 bl[120] br[120] wl[293] vdd gnd cell_6t
Xbit_r294_c120 bl[120] br[120] wl[294] vdd gnd cell_6t
Xbit_r295_c120 bl[120] br[120] wl[295] vdd gnd cell_6t
Xbit_r296_c120 bl[120] br[120] wl[296] vdd gnd cell_6t
Xbit_r297_c120 bl[120] br[120] wl[297] vdd gnd cell_6t
Xbit_r298_c120 bl[120] br[120] wl[298] vdd gnd cell_6t
Xbit_r299_c120 bl[120] br[120] wl[299] vdd gnd cell_6t
Xbit_r300_c120 bl[120] br[120] wl[300] vdd gnd cell_6t
Xbit_r301_c120 bl[120] br[120] wl[301] vdd gnd cell_6t
Xbit_r302_c120 bl[120] br[120] wl[302] vdd gnd cell_6t
Xbit_r303_c120 bl[120] br[120] wl[303] vdd gnd cell_6t
Xbit_r304_c120 bl[120] br[120] wl[304] vdd gnd cell_6t
Xbit_r305_c120 bl[120] br[120] wl[305] vdd gnd cell_6t
Xbit_r306_c120 bl[120] br[120] wl[306] vdd gnd cell_6t
Xbit_r307_c120 bl[120] br[120] wl[307] vdd gnd cell_6t
Xbit_r308_c120 bl[120] br[120] wl[308] vdd gnd cell_6t
Xbit_r309_c120 bl[120] br[120] wl[309] vdd gnd cell_6t
Xbit_r310_c120 bl[120] br[120] wl[310] vdd gnd cell_6t
Xbit_r311_c120 bl[120] br[120] wl[311] vdd gnd cell_6t
Xbit_r312_c120 bl[120] br[120] wl[312] vdd gnd cell_6t
Xbit_r313_c120 bl[120] br[120] wl[313] vdd gnd cell_6t
Xbit_r314_c120 bl[120] br[120] wl[314] vdd gnd cell_6t
Xbit_r315_c120 bl[120] br[120] wl[315] vdd gnd cell_6t
Xbit_r316_c120 bl[120] br[120] wl[316] vdd gnd cell_6t
Xbit_r317_c120 bl[120] br[120] wl[317] vdd gnd cell_6t
Xbit_r318_c120 bl[120] br[120] wl[318] vdd gnd cell_6t
Xbit_r319_c120 bl[120] br[120] wl[319] vdd gnd cell_6t
Xbit_r320_c120 bl[120] br[120] wl[320] vdd gnd cell_6t
Xbit_r321_c120 bl[120] br[120] wl[321] vdd gnd cell_6t
Xbit_r322_c120 bl[120] br[120] wl[322] vdd gnd cell_6t
Xbit_r323_c120 bl[120] br[120] wl[323] vdd gnd cell_6t
Xbit_r324_c120 bl[120] br[120] wl[324] vdd gnd cell_6t
Xbit_r325_c120 bl[120] br[120] wl[325] vdd gnd cell_6t
Xbit_r326_c120 bl[120] br[120] wl[326] vdd gnd cell_6t
Xbit_r327_c120 bl[120] br[120] wl[327] vdd gnd cell_6t
Xbit_r328_c120 bl[120] br[120] wl[328] vdd gnd cell_6t
Xbit_r329_c120 bl[120] br[120] wl[329] vdd gnd cell_6t
Xbit_r330_c120 bl[120] br[120] wl[330] vdd gnd cell_6t
Xbit_r331_c120 bl[120] br[120] wl[331] vdd gnd cell_6t
Xbit_r332_c120 bl[120] br[120] wl[332] vdd gnd cell_6t
Xbit_r333_c120 bl[120] br[120] wl[333] vdd gnd cell_6t
Xbit_r334_c120 bl[120] br[120] wl[334] vdd gnd cell_6t
Xbit_r335_c120 bl[120] br[120] wl[335] vdd gnd cell_6t
Xbit_r336_c120 bl[120] br[120] wl[336] vdd gnd cell_6t
Xbit_r337_c120 bl[120] br[120] wl[337] vdd gnd cell_6t
Xbit_r338_c120 bl[120] br[120] wl[338] vdd gnd cell_6t
Xbit_r339_c120 bl[120] br[120] wl[339] vdd gnd cell_6t
Xbit_r340_c120 bl[120] br[120] wl[340] vdd gnd cell_6t
Xbit_r341_c120 bl[120] br[120] wl[341] vdd gnd cell_6t
Xbit_r342_c120 bl[120] br[120] wl[342] vdd gnd cell_6t
Xbit_r343_c120 bl[120] br[120] wl[343] vdd gnd cell_6t
Xbit_r344_c120 bl[120] br[120] wl[344] vdd gnd cell_6t
Xbit_r345_c120 bl[120] br[120] wl[345] vdd gnd cell_6t
Xbit_r346_c120 bl[120] br[120] wl[346] vdd gnd cell_6t
Xbit_r347_c120 bl[120] br[120] wl[347] vdd gnd cell_6t
Xbit_r348_c120 bl[120] br[120] wl[348] vdd gnd cell_6t
Xbit_r349_c120 bl[120] br[120] wl[349] vdd gnd cell_6t
Xbit_r350_c120 bl[120] br[120] wl[350] vdd gnd cell_6t
Xbit_r351_c120 bl[120] br[120] wl[351] vdd gnd cell_6t
Xbit_r352_c120 bl[120] br[120] wl[352] vdd gnd cell_6t
Xbit_r353_c120 bl[120] br[120] wl[353] vdd gnd cell_6t
Xbit_r354_c120 bl[120] br[120] wl[354] vdd gnd cell_6t
Xbit_r355_c120 bl[120] br[120] wl[355] vdd gnd cell_6t
Xbit_r356_c120 bl[120] br[120] wl[356] vdd gnd cell_6t
Xbit_r357_c120 bl[120] br[120] wl[357] vdd gnd cell_6t
Xbit_r358_c120 bl[120] br[120] wl[358] vdd gnd cell_6t
Xbit_r359_c120 bl[120] br[120] wl[359] vdd gnd cell_6t
Xbit_r360_c120 bl[120] br[120] wl[360] vdd gnd cell_6t
Xbit_r361_c120 bl[120] br[120] wl[361] vdd gnd cell_6t
Xbit_r362_c120 bl[120] br[120] wl[362] vdd gnd cell_6t
Xbit_r363_c120 bl[120] br[120] wl[363] vdd gnd cell_6t
Xbit_r364_c120 bl[120] br[120] wl[364] vdd gnd cell_6t
Xbit_r365_c120 bl[120] br[120] wl[365] vdd gnd cell_6t
Xbit_r366_c120 bl[120] br[120] wl[366] vdd gnd cell_6t
Xbit_r367_c120 bl[120] br[120] wl[367] vdd gnd cell_6t
Xbit_r368_c120 bl[120] br[120] wl[368] vdd gnd cell_6t
Xbit_r369_c120 bl[120] br[120] wl[369] vdd gnd cell_6t
Xbit_r370_c120 bl[120] br[120] wl[370] vdd gnd cell_6t
Xbit_r371_c120 bl[120] br[120] wl[371] vdd gnd cell_6t
Xbit_r372_c120 bl[120] br[120] wl[372] vdd gnd cell_6t
Xbit_r373_c120 bl[120] br[120] wl[373] vdd gnd cell_6t
Xbit_r374_c120 bl[120] br[120] wl[374] vdd gnd cell_6t
Xbit_r375_c120 bl[120] br[120] wl[375] vdd gnd cell_6t
Xbit_r376_c120 bl[120] br[120] wl[376] vdd gnd cell_6t
Xbit_r377_c120 bl[120] br[120] wl[377] vdd gnd cell_6t
Xbit_r378_c120 bl[120] br[120] wl[378] vdd gnd cell_6t
Xbit_r379_c120 bl[120] br[120] wl[379] vdd gnd cell_6t
Xbit_r380_c120 bl[120] br[120] wl[380] vdd gnd cell_6t
Xbit_r381_c120 bl[120] br[120] wl[381] vdd gnd cell_6t
Xbit_r382_c120 bl[120] br[120] wl[382] vdd gnd cell_6t
Xbit_r383_c120 bl[120] br[120] wl[383] vdd gnd cell_6t
Xbit_r384_c120 bl[120] br[120] wl[384] vdd gnd cell_6t
Xbit_r385_c120 bl[120] br[120] wl[385] vdd gnd cell_6t
Xbit_r386_c120 bl[120] br[120] wl[386] vdd gnd cell_6t
Xbit_r387_c120 bl[120] br[120] wl[387] vdd gnd cell_6t
Xbit_r388_c120 bl[120] br[120] wl[388] vdd gnd cell_6t
Xbit_r389_c120 bl[120] br[120] wl[389] vdd gnd cell_6t
Xbit_r390_c120 bl[120] br[120] wl[390] vdd gnd cell_6t
Xbit_r391_c120 bl[120] br[120] wl[391] vdd gnd cell_6t
Xbit_r392_c120 bl[120] br[120] wl[392] vdd gnd cell_6t
Xbit_r393_c120 bl[120] br[120] wl[393] vdd gnd cell_6t
Xbit_r394_c120 bl[120] br[120] wl[394] vdd gnd cell_6t
Xbit_r395_c120 bl[120] br[120] wl[395] vdd gnd cell_6t
Xbit_r396_c120 bl[120] br[120] wl[396] vdd gnd cell_6t
Xbit_r397_c120 bl[120] br[120] wl[397] vdd gnd cell_6t
Xbit_r398_c120 bl[120] br[120] wl[398] vdd gnd cell_6t
Xbit_r399_c120 bl[120] br[120] wl[399] vdd gnd cell_6t
Xbit_r400_c120 bl[120] br[120] wl[400] vdd gnd cell_6t
Xbit_r401_c120 bl[120] br[120] wl[401] vdd gnd cell_6t
Xbit_r402_c120 bl[120] br[120] wl[402] vdd gnd cell_6t
Xbit_r403_c120 bl[120] br[120] wl[403] vdd gnd cell_6t
Xbit_r404_c120 bl[120] br[120] wl[404] vdd gnd cell_6t
Xbit_r405_c120 bl[120] br[120] wl[405] vdd gnd cell_6t
Xbit_r406_c120 bl[120] br[120] wl[406] vdd gnd cell_6t
Xbit_r407_c120 bl[120] br[120] wl[407] vdd gnd cell_6t
Xbit_r408_c120 bl[120] br[120] wl[408] vdd gnd cell_6t
Xbit_r409_c120 bl[120] br[120] wl[409] vdd gnd cell_6t
Xbit_r410_c120 bl[120] br[120] wl[410] vdd gnd cell_6t
Xbit_r411_c120 bl[120] br[120] wl[411] vdd gnd cell_6t
Xbit_r412_c120 bl[120] br[120] wl[412] vdd gnd cell_6t
Xbit_r413_c120 bl[120] br[120] wl[413] vdd gnd cell_6t
Xbit_r414_c120 bl[120] br[120] wl[414] vdd gnd cell_6t
Xbit_r415_c120 bl[120] br[120] wl[415] vdd gnd cell_6t
Xbit_r416_c120 bl[120] br[120] wl[416] vdd gnd cell_6t
Xbit_r417_c120 bl[120] br[120] wl[417] vdd gnd cell_6t
Xbit_r418_c120 bl[120] br[120] wl[418] vdd gnd cell_6t
Xbit_r419_c120 bl[120] br[120] wl[419] vdd gnd cell_6t
Xbit_r420_c120 bl[120] br[120] wl[420] vdd gnd cell_6t
Xbit_r421_c120 bl[120] br[120] wl[421] vdd gnd cell_6t
Xbit_r422_c120 bl[120] br[120] wl[422] vdd gnd cell_6t
Xbit_r423_c120 bl[120] br[120] wl[423] vdd gnd cell_6t
Xbit_r424_c120 bl[120] br[120] wl[424] vdd gnd cell_6t
Xbit_r425_c120 bl[120] br[120] wl[425] vdd gnd cell_6t
Xbit_r426_c120 bl[120] br[120] wl[426] vdd gnd cell_6t
Xbit_r427_c120 bl[120] br[120] wl[427] vdd gnd cell_6t
Xbit_r428_c120 bl[120] br[120] wl[428] vdd gnd cell_6t
Xbit_r429_c120 bl[120] br[120] wl[429] vdd gnd cell_6t
Xbit_r430_c120 bl[120] br[120] wl[430] vdd gnd cell_6t
Xbit_r431_c120 bl[120] br[120] wl[431] vdd gnd cell_6t
Xbit_r432_c120 bl[120] br[120] wl[432] vdd gnd cell_6t
Xbit_r433_c120 bl[120] br[120] wl[433] vdd gnd cell_6t
Xbit_r434_c120 bl[120] br[120] wl[434] vdd gnd cell_6t
Xbit_r435_c120 bl[120] br[120] wl[435] vdd gnd cell_6t
Xbit_r436_c120 bl[120] br[120] wl[436] vdd gnd cell_6t
Xbit_r437_c120 bl[120] br[120] wl[437] vdd gnd cell_6t
Xbit_r438_c120 bl[120] br[120] wl[438] vdd gnd cell_6t
Xbit_r439_c120 bl[120] br[120] wl[439] vdd gnd cell_6t
Xbit_r440_c120 bl[120] br[120] wl[440] vdd gnd cell_6t
Xbit_r441_c120 bl[120] br[120] wl[441] vdd gnd cell_6t
Xbit_r442_c120 bl[120] br[120] wl[442] vdd gnd cell_6t
Xbit_r443_c120 bl[120] br[120] wl[443] vdd gnd cell_6t
Xbit_r444_c120 bl[120] br[120] wl[444] vdd gnd cell_6t
Xbit_r445_c120 bl[120] br[120] wl[445] vdd gnd cell_6t
Xbit_r446_c120 bl[120] br[120] wl[446] vdd gnd cell_6t
Xbit_r447_c120 bl[120] br[120] wl[447] vdd gnd cell_6t
Xbit_r448_c120 bl[120] br[120] wl[448] vdd gnd cell_6t
Xbit_r449_c120 bl[120] br[120] wl[449] vdd gnd cell_6t
Xbit_r450_c120 bl[120] br[120] wl[450] vdd gnd cell_6t
Xbit_r451_c120 bl[120] br[120] wl[451] vdd gnd cell_6t
Xbit_r452_c120 bl[120] br[120] wl[452] vdd gnd cell_6t
Xbit_r453_c120 bl[120] br[120] wl[453] vdd gnd cell_6t
Xbit_r454_c120 bl[120] br[120] wl[454] vdd gnd cell_6t
Xbit_r455_c120 bl[120] br[120] wl[455] vdd gnd cell_6t
Xbit_r456_c120 bl[120] br[120] wl[456] vdd gnd cell_6t
Xbit_r457_c120 bl[120] br[120] wl[457] vdd gnd cell_6t
Xbit_r458_c120 bl[120] br[120] wl[458] vdd gnd cell_6t
Xbit_r459_c120 bl[120] br[120] wl[459] vdd gnd cell_6t
Xbit_r460_c120 bl[120] br[120] wl[460] vdd gnd cell_6t
Xbit_r461_c120 bl[120] br[120] wl[461] vdd gnd cell_6t
Xbit_r462_c120 bl[120] br[120] wl[462] vdd gnd cell_6t
Xbit_r463_c120 bl[120] br[120] wl[463] vdd gnd cell_6t
Xbit_r464_c120 bl[120] br[120] wl[464] vdd gnd cell_6t
Xbit_r465_c120 bl[120] br[120] wl[465] vdd gnd cell_6t
Xbit_r466_c120 bl[120] br[120] wl[466] vdd gnd cell_6t
Xbit_r467_c120 bl[120] br[120] wl[467] vdd gnd cell_6t
Xbit_r468_c120 bl[120] br[120] wl[468] vdd gnd cell_6t
Xbit_r469_c120 bl[120] br[120] wl[469] vdd gnd cell_6t
Xbit_r470_c120 bl[120] br[120] wl[470] vdd gnd cell_6t
Xbit_r471_c120 bl[120] br[120] wl[471] vdd gnd cell_6t
Xbit_r472_c120 bl[120] br[120] wl[472] vdd gnd cell_6t
Xbit_r473_c120 bl[120] br[120] wl[473] vdd gnd cell_6t
Xbit_r474_c120 bl[120] br[120] wl[474] vdd gnd cell_6t
Xbit_r475_c120 bl[120] br[120] wl[475] vdd gnd cell_6t
Xbit_r476_c120 bl[120] br[120] wl[476] vdd gnd cell_6t
Xbit_r477_c120 bl[120] br[120] wl[477] vdd gnd cell_6t
Xbit_r478_c120 bl[120] br[120] wl[478] vdd gnd cell_6t
Xbit_r479_c120 bl[120] br[120] wl[479] vdd gnd cell_6t
Xbit_r480_c120 bl[120] br[120] wl[480] vdd gnd cell_6t
Xbit_r481_c120 bl[120] br[120] wl[481] vdd gnd cell_6t
Xbit_r482_c120 bl[120] br[120] wl[482] vdd gnd cell_6t
Xbit_r483_c120 bl[120] br[120] wl[483] vdd gnd cell_6t
Xbit_r484_c120 bl[120] br[120] wl[484] vdd gnd cell_6t
Xbit_r485_c120 bl[120] br[120] wl[485] vdd gnd cell_6t
Xbit_r486_c120 bl[120] br[120] wl[486] vdd gnd cell_6t
Xbit_r487_c120 bl[120] br[120] wl[487] vdd gnd cell_6t
Xbit_r488_c120 bl[120] br[120] wl[488] vdd gnd cell_6t
Xbit_r489_c120 bl[120] br[120] wl[489] vdd gnd cell_6t
Xbit_r490_c120 bl[120] br[120] wl[490] vdd gnd cell_6t
Xbit_r491_c120 bl[120] br[120] wl[491] vdd gnd cell_6t
Xbit_r492_c120 bl[120] br[120] wl[492] vdd gnd cell_6t
Xbit_r493_c120 bl[120] br[120] wl[493] vdd gnd cell_6t
Xbit_r494_c120 bl[120] br[120] wl[494] vdd gnd cell_6t
Xbit_r495_c120 bl[120] br[120] wl[495] vdd gnd cell_6t
Xbit_r496_c120 bl[120] br[120] wl[496] vdd gnd cell_6t
Xbit_r497_c120 bl[120] br[120] wl[497] vdd gnd cell_6t
Xbit_r498_c120 bl[120] br[120] wl[498] vdd gnd cell_6t
Xbit_r499_c120 bl[120] br[120] wl[499] vdd gnd cell_6t
Xbit_r500_c120 bl[120] br[120] wl[500] vdd gnd cell_6t
Xbit_r501_c120 bl[120] br[120] wl[501] vdd gnd cell_6t
Xbit_r502_c120 bl[120] br[120] wl[502] vdd gnd cell_6t
Xbit_r503_c120 bl[120] br[120] wl[503] vdd gnd cell_6t
Xbit_r504_c120 bl[120] br[120] wl[504] vdd gnd cell_6t
Xbit_r505_c120 bl[120] br[120] wl[505] vdd gnd cell_6t
Xbit_r506_c120 bl[120] br[120] wl[506] vdd gnd cell_6t
Xbit_r507_c120 bl[120] br[120] wl[507] vdd gnd cell_6t
Xbit_r508_c120 bl[120] br[120] wl[508] vdd gnd cell_6t
Xbit_r509_c120 bl[120] br[120] wl[509] vdd gnd cell_6t
Xbit_r510_c120 bl[120] br[120] wl[510] vdd gnd cell_6t
Xbit_r511_c120 bl[120] br[120] wl[511] vdd gnd cell_6t
Xbit_r0_c121 bl[121] br[121] wl[0] vdd gnd cell_6t
Xbit_r1_c121 bl[121] br[121] wl[1] vdd gnd cell_6t
Xbit_r2_c121 bl[121] br[121] wl[2] vdd gnd cell_6t
Xbit_r3_c121 bl[121] br[121] wl[3] vdd gnd cell_6t
Xbit_r4_c121 bl[121] br[121] wl[4] vdd gnd cell_6t
Xbit_r5_c121 bl[121] br[121] wl[5] vdd gnd cell_6t
Xbit_r6_c121 bl[121] br[121] wl[6] vdd gnd cell_6t
Xbit_r7_c121 bl[121] br[121] wl[7] vdd gnd cell_6t
Xbit_r8_c121 bl[121] br[121] wl[8] vdd gnd cell_6t
Xbit_r9_c121 bl[121] br[121] wl[9] vdd gnd cell_6t
Xbit_r10_c121 bl[121] br[121] wl[10] vdd gnd cell_6t
Xbit_r11_c121 bl[121] br[121] wl[11] vdd gnd cell_6t
Xbit_r12_c121 bl[121] br[121] wl[12] vdd gnd cell_6t
Xbit_r13_c121 bl[121] br[121] wl[13] vdd gnd cell_6t
Xbit_r14_c121 bl[121] br[121] wl[14] vdd gnd cell_6t
Xbit_r15_c121 bl[121] br[121] wl[15] vdd gnd cell_6t
Xbit_r16_c121 bl[121] br[121] wl[16] vdd gnd cell_6t
Xbit_r17_c121 bl[121] br[121] wl[17] vdd gnd cell_6t
Xbit_r18_c121 bl[121] br[121] wl[18] vdd gnd cell_6t
Xbit_r19_c121 bl[121] br[121] wl[19] vdd gnd cell_6t
Xbit_r20_c121 bl[121] br[121] wl[20] vdd gnd cell_6t
Xbit_r21_c121 bl[121] br[121] wl[21] vdd gnd cell_6t
Xbit_r22_c121 bl[121] br[121] wl[22] vdd gnd cell_6t
Xbit_r23_c121 bl[121] br[121] wl[23] vdd gnd cell_6t
Xbit_r24_c121 bl[121] br[121] wl[24] vdd gnd cell_6t
Xbit_r25_c121 bl[121] br[121] wl[25] vdd gnd cell_6t
Xbit_r26_c121 bl[121] br[121] wl[26] vdd gnd cell_6t
Xbit_r27_c121 bl[121] br[121] wl[27] vdd gnd cell_6t
Xbit_r28_c121 bl[121] br[121] wl[28] vdd gnd cell_6t
Xbit_r29_c121 bl[121] br[121] wl[29] vdd gnd cell_6t
Xbit_r30_c121 bl[121] br[121] wl[30] vdd gnd cell_6t
Xbit_r31_c121 bl[121] br[121] wl[31] vdd gnd cell_6t
Xbit_r32_c121 bl[121] br[121] wl[32] vdd gnd cell_6t
Xbit_r33_c121 bl[121] br[121] wl[33] vdd gnd cell_6t
Xbit_r34_c121 bl[121] br[121] wl[34] vdd gnd cell_6t
Xbit_r35_c121 bl[121] br[121] wl[35] vdd gnd cell_6t
Xbit_r36_c121 bl[121] br[121] wl[36] vdd gnd cell_6t
Xbit_r37_c121 bl[121] br[121] wl[37] vdd gnd cell_6t
Xbit_r38_c121 bl[121] br[121] wl[38] vdd gnd cell_6t
Xbit_r39_c121 bl[121] br[121] wl[39] vdd gnd cell_6t
Xbit_r40_c121 bl[121] br[121] wl[40] vdd gnd cell_6t
Xbit_r41_c121 bl[121] br[121] wl[41] vdd gnd cell_6t
Xbit_r42_c121 bl[121] br[121] wl[42] vdd gnd cell_6t
Xbit_r43_c121 bl[121] br[121] wl[43] vdd gnd cell_6t
Xbit_r44_c121 bl[121] br[121] wl[44] vdd gnd cell_6t
Xbit_r45_c121 bl[121] br[121] wl[45] vdd gnd cell_6t
Xbit_r46_c121 bl[121] br[121] wl[46] vdd gnd cell_6t
Xbit_r47_c121 bl[121] br[121] wl[47] vdd gnd cell_6t
Xbit_r48_c121 bl[121] br[121] wl[48] vdd gnd cell_6t
Xbit_r49_c121 bl[121] br[121] wl[49] vdd gnd cell_6t
Xbit_r50_c121 bl[121] br[121] wl[50] vdd gnd cell_6t
Xbit_r51_c121 bl[121] br[121] wl[51] vdd gnd cell_6t
Xbit_r52_c121 bl[121] br[121] wl[52] vdd gnd cell_6t
Xbit_r53_c121 bl[121] br[121] wl[53] vdd gnd cell_6t
Xbit_r54_c121 bl[121] br[121] wl[54] vdd gnd cell_6t
Xbit_r55_c121 bl[121] br[121] wl[55] vdd gnd cell_6t
Xbit_r56_c121 bl[121] br[121] wl[56] vdd gnd cell_6t
Xbit_r57_c121 bl[121] br[121] wl[57] vdd gnd cell_6t
Xbit_r58_c121 bl[121] br[121] wl[58] vdd gnd cell_6t
Xbit_r59_c121 bl[121] br[121] wl[59] vdd gnd cell_6t
Xbit_r60_c121 bl[121] br[121] wl[60] vdd gnd cell_6t
Xbit_r61_c121 bl[121] br[121] wl[61] vdd gnd cell_6t
Xbit_r62_c121 bl[121] br[121] wl[62] vdd gnd cell_6t
Xbit_r63_c121 bl[121] br[121] wl[63] vdd gnd cell_6t
Xbit_r64_c121 bl[121] br[121] wl[64] vdd gnd cell_6t
Xbit_r65_c121 bl[121] br[121] wl[65] vdd gnd cell_6t
Xbit_r66_c121 bl[121] br[121] wl[66] vdd gnd cell_6t
Xbit_r67_c121 bl[121] br[121] wl[67] vdd gnd cell_6t
Xbit_r68_c121 bl[121] br[121] wl[68] vdd gnd cell_6t
Xbit_r69_c121 bl[121] br[121] wl[69] vdd gnd cell_6t
Xbit_r70_c121 bl[121] br[121] wl[70] vdd gnd cell_6t
Xbit_r71_c121 bl[121] br[121] wl[71] vdd gnd cell_6t
Xbit_r72_c121 bl[121] br[121] wl[72] vdd gnd cell_6t
Xbit_r73_c121 bl[121] br[121] wl[73] vdd gnd cell_6t
Xbit_r74_c121 bl[121] br[121] wl[74] vdd gnd cell_6t
Xbit_r75_c121 bl[121] br[121] wl[75] vdd gnd cell_6t
Xbit_r76_c121 bl[121] br[121] wl[76] vdd gnd cell_6t
Xbit_r77_c121 bl[121] br[121] wl[77] vdd gnd cell_6t
Xbit_r78_c121 bl[121] br[121] wl[78] vdd gnd cell_6t
Xbit_r79_c121 bl[121] br[121] wl[79] vdd gnd cell_6t
Xbit_r80_c121 bl[121] br[121] wl[80] vdd gnd cell_6t
Xbit_r81_c121 bl[121] br[121] wl[81] vdd gnd cell_6t
Xbit_r82_c121 bl[121] br[121] wl[82] vdd gnd cell_6t
Xbit_r83_c121 bl[121] br[121] wl[83] vdd gnd cell_6t
Xbit_r84_c121 bl[121] br[121] wl[84] vdd gnd cell_6t
Xbit_r85_c121 bl[121] br[121] wl[85] vdd gnd cell_6t
Xbit_r86_c121 bl[121] br[121] wl[86] vdd gnd cell_6t
Xbit_r87_c121 bl[121] br[121] wl[87] vdd gnd cell_6t
Xbit_r88_c121 bl[121] br[121] wl[88] vdd gnd cell_6t
Xbit_r89_c121 bl[121] br[121] wl[89] vdd gnd cell_6t
Xbit_r90_c121 bl[121] br[121] wl[90] vdd gnd cell_6t
Xbit_r91_c121 bl[121] br[121] wl[91] vdd gnd cell_6t
Xbit_r92_c121 bl[121] br[121] wl[92] vdd gnd cell_6t
Xbit_r93_c121 bl[121] br[121] wl[93] vdd gnd cell_6t
Xbit_r94_c121 bl[121] br[121] wl[94] vdd gnd cell_6t
Xbit_r95_c121 bl[121] br[121] wl[95] vdd gnd cell_6t
Xbit_r96_c121 bl[121] br[121] wl[96] vdd gnd cell_6t
Xbit_r97_c121 bl[121] br[121] wl[97] vdd gnd cell_6t
Xbit_r98_c121 bl[121] br[121] wl[98] vdd gnd cell_6t
Xbit_r99_c121 bl[121] br[121] wl[99] vdd gnd cell_6t
Xbit_r100_c121 bl[121] br[121] wl[100] vdd gnd cell_6t
Xbit_r101_c121 bl[121] br[121] wl[101] vdd gnd cell_6t
Xbit_r102_c121 bl[121] br[121] wl[102] vdd gnd cell_6t
Xbit_r103_c121 bl[121] br[121] wl[103] vdd gnd cell_6t
Xbit_r104_c121 bl[121] br[121] wl[104] vdd gnd cell_6t
Xbit_r105_c121 bl[121] br[121] wl[105] vdd gnd cell_6t
Xbit_r106_c121 bl[121] br[121] wl[106] vdd gnd cell_6t
Xbit_r107_c121 bl[121] br[121] wl[107] vdd gnd cell_6t
Xbit_r108_c121 bl[121] br[121] wl[108] vdd gnd cell_6t
Xbit_r109_c121 bl[121] br[121] wl[109] vdd gnd cell_6t
Xbit_r110_c121 bl[121] br[121] wl[110] vdd gnd cell_6t
Xbit_r111_c121 bl[121] br[121] wl[111] vdd gnd cell_6t
Xbit_r112_c121 bl[121] br[121] wl[112] vdd gnd cell_6t
Xbit_r113_c121 bl[121] br[121] wl[113] vdd gnd cell_6t
Xbit_r114_c121 bl[121] br[121] wl[114] vdd gnd cell_6t
Xbit_r115_c121 bl[121] br[121] wl[115] vdd gnd cell_6t
Xbit_r116_c121 bl[121] br[121] wl[116] vdd gnd cell_6t
Xbit_r117_c121 bl[121] br[121] wl[117] vdd gnd cell_6t
Xbit_r118_c121 bl[121] br[121] wl[118] vdd gnd cell_6t
Xbit_r119_c121 bl[121] br[121] wl[119] vdd gnd cell_6t
Xbit_r120_c121 bl[121] br[121] wl[120] vdd gnd cell_6t
Xbit_r121_c121 bl[121] br[121] wl[121] vdd gnd cell_6t
Xbit_r122_c121 bl[121] br[121] wl[122] vdd gnd cell_6t
Xbit_r123_c121 bl[121] br[121] wl[123] vdd gnd cell_6t
Xbit_r124_c121 bl[121] br[121] wl[124] vdd gnd cell_6t
Xbit_r125_c121 bl[121] br[121] wl[125] vdd gnd cell_6t
Xbit_r126_c121 bl[121] br[121] wl[126] vdd gnd cell_6t
Xbit_r127_c121 bl[121] br[121] wl[127] vdd gnd cell_6t
Xbit_r128_c121 bl[121] br[121] wl[128] vdd gnd cell_6t
Xbit_r129_c121 bl[121] br[121] wl[129] vdd gnd cell_6t
Xbit_r130_c121 bl[121] br[121] wl[130] vdd gnd cell_6t
Xbit_r131_c121 bl[121] br[121] wl[131] vdd gnd cell_6t
Xbit_r132_c121 bl[121] br[121] wl[132] vdd gnd cell_6t
Xbit_r133_c121 bl[121] br[121] wl[133] vdd gnd cell_6t
Xbit_r134_c121 bl[121] br[121] wl[134] vdd gnd cell_6t
Xbit_r135_c121 bl[121] br[121] wl[135] vdd gnd cell_6t
Xbit_r136_c121 bl[121] br[121] wl[136] vdd gnd cell_6t
Xbit_r137_c121 bl[121] br[121] wl[137] vdd gnd cell_6t
Xbit_r138_c121 bl[121] br[121] wl[138] vdd gnd cell_6t
Xbit_r139_c121 bl[121] br[121] wl[139] vdd gnd cell_6t
Xbit_r140_c121 bl[121] br[121] wl[140] vdd gnd cell_6t
Xbit_r141_c121 bl[121] br[121] wl[141] vdd gnd cell_6t
Xbit_r142_c121 bl[121] br[121] wl[142] vdd gnd cell_6t
Xbit_r143_c121 bl[121] br[121] wl[143] vdd gnd cell_6t
Xbit_r144_c121 bl[121] br[121] wl[144] vdd gnd cell_6t
Xbit_r145_c121 bl[121] br[121] wl[145] vdd gnd cell_6t
Xbit_r146_c121 bl[121] br[121] wl[146] vdd gnd cell_6t
Xbit_r147_c121 bl[121] br[121] wl[147] vdd gnd cell_6t
Xbit_r148_c121 bl[121] br[121] wl[148] vdd gnd cell_6t
Xbit_r149_c121 bl[121] br[121] wl[149] vdd gnd cell_6t
Xbit_r150_c121 bl[121] br[121] wl[150] vdd gnd cell_6t
Xbit_r151_c121 bl[121] br[121] wl[151] vdd gnd cell_6t
Xbit_r152_c121 bl[121] br[121] wl[152] vdd gnd cell_6t
Xbit_r153_c121 bl[121] br[121] wl[153] vdd gnd cell_6t
Xbit_r154_c121 bl[121] br[121] wl[154] vdd gnd cell_6t
Xbit_r155_c121 bl[121] br[121] wl[155] vdd gnd cell_6t
Xbit_r156_c121 bl[121] br[121] wl[156] vdd gnd cell_6t
Xbit_r157_c121 bl[121] br[121] wl[157] vdd gnd cell_6t
Xbit_r158_c121 bl[121] br[121] wl[158] vdd gnd cell_6t
Xbit_r159_c121 bl[121] br[121] wl[159] vdd gnd cell_6t
Xbit_r160_c121 bl[121] br[121] wl[160] vdd gnd cell_6t
Xbit_r161_c121 bl[121] br[121] wl[161] vdd gnd cell_6t
Xbit_r162_c121 bl[121] br[121] wl[162] vdd gnd cell_6t
Xbit_r163_c121 bl[121] br[121] wl[163] vdd gnd cell_6t
Xbit_r164_c121 bl[121] br[121] wl[164] vdd gnd cell_6t
Xbit_r165_c121 bl[121] br[121] wl[165] vdd gnd cell_6t
Xbit_r166_c121 bl[121] br[121] wl[166] vdd gnd cell_6t
Xbit_r167_c121 bl[121] br[121] wl[167] vdd gnd cell_6t
Xbit_r168_c121 bl[121] br[121] wl[168] vdd gnd cell_6t
Xbit_r169_c121 bl[121] br[121] wl[169] vdd gnd cell_6t
Xbit_r170_c121 bl[121] br[121] wl[170] vdd gnd cell_6t
Xbit_r171_c121 bl[121] br[121] wl[171] vdd gnd cell_6t
Xbit_r172_c121 bl[121] br[121] wl[172] vdd gnd cell_6t
Xbit_r173_c121 bl[121] br[121] wl[173] vdd gnd cell_6t
Xbit_r174_c121 bl[121] br[121] wl[174] vdd gnd cell_6t
Xbit_r175_c121 bl[121] br[121] wl[175] vdd gnd cell_6t
Xbit_r176_c121 bl[121] br[121] wl[176] vdd gnd cell_6t
Xbit_r177_c121 bl[121] br[121] wl[177] vdd gnd cell_6t
Xbit_r178_c121 bl[121] br[121] wl[178] vdd gnd cell_6t
Xbit_r179_c121 bl[121] br[121] wl[179] vdd gnd cell_6t
Xbit_r180_c121 bl[121] br[121] wl[180] vdd gnd cell_6t
Xbit_r181_c121 bl[121] br[121] wl[181] vdd gnd cell_6t
Xbit_r182_c121 bl[121] br[121] wl[182] vdd gnd cell_6t
Xbit_r183_c121 bl[121] br[121] wl[183] vdd gnd cell_6t
Xbit_r184_c121 bl[121] br[121] wl[184] vdd gnd cell_6t
Xbit_r185_c121 bl[121] br[121] wl[185] vdd gnd cell_6t
Xbit_r186_c121 bl[121] br[121] wl[186] vdd gnd cell_6t
Xbit_r187_c121 bl[121] br[121] wl[187] vdd gnd cell_6t
Xbit_r188_c121 bl[121] br[121] wl[188] vdd gnd cell_6t
Xbit_r189_c121 bl[121] br[121] wl[189] vdd gnd cell_6t
Xbit_r190_c121 bl[121] br[121] wl[190] vdd gnd cell_6t
Xbit_r191_c121 bl[121] br[121] wl[191] vdd gnd cell_6t
Xbit_r192_c121 bl[121] br[121] wl[192] vdd gnd cell_6t
Xbit_r193_c121 bl[121] br[121] wl[193] vdd gnd cell_6t
Xbit_r194_c121 bl[121] br[121] wl[194] vdd gnd cell_6t
Xbit_r195_c121 bl[121] br[121] wl[195] vdd gnd cell_6t
Xbit_r196_c121 bl[121] br[121] wl[196] vdd gnd cell_6t
Xbit_r197_c121 bl[121] br[121] wl[197] vdd gnd cell_6t
Xbit_r198_c121 bl[121] br[121] wl[198] vdd gnd cell_6t
Xbit_r199_c121 bl[121] br[121] wl[199] vdd gnd cell_6t
Xbit_r200_c121 bl[121] br[121] wl[200] vdd gnd cell_6t
Xbit_r201_c121 bl[121] br[121] wl[201] vdd gnd cell_6t
Xbit_r202_c121 bl[121] br[121] wl[202] vdd gnd cell_6t
Xbit_r203_c121 bl[121] br[121] wl[203] vdd gnd cell_6t
Xbit_r204_c121 bl[121] br[121] wl[204] vdd gnd cell_6t
Xbit_r205_c121 bl[121] br[121] wl[205] vdd gnd cell_6t
Xbit_r206_c121 bl[121] br[121] wl[206] vdd gnd cell_6t
Xbit_r207_c121 bl[121] br[121] wl[207] vdd gnd cell_6t
Xbit_r208_c121 bl[121] br[121] wl[208] vdd gnd cell_6t
Xbit_r209_c121 bl[121] br[121] wl[209] vdd gnd cell_6t
Xbit_r210_c121 bl[121] br[121] wl[210] vdd gnd cell_6t
Xbit_r211_c121 bl[121] br[121] wl[211] vdd gnd cell_6t
Xbit_r212_c121 bl[121] br[121] wl[212] vdd gnd cell_6t
Xbit_r213_c121 bl[121] br[121] wl[213] vdd gnd cell_6t
Xbit_r214_c121 bl[121] br[121] wl[214] vdd gnd cell_6t
Xbit_r215_c121 bl[121] br[121] wl[215] vdd gnd cell_6t
Xbit_r216_c121 bl[121] br[121] wl[216] vdd gnd cell_6t
Xbit_r217_c121 bl[121] br[121] wl[217] vdd gnd cell_6t
Xbit_r218_c121 bl[121] br[121] wl[218] vdd gnd cell_6t
Xbit_r219_c121 bl[121] br[121] wl[219] vdd gnd cell_6t
Xbit_r220_c121 bl[121] br[121] wl[220] vdd gnd cell_6t
Xbit_r221_c121 bl[121] br[121] wl[221] vdd gnd cell_6t
Xbit_r222_c121 bl[121] br[121] wl[222] vdd gnd cell_6t
Xbit_r223_c121 bl[121] br[121] wl[223] vdd gnd cell_6t
Xbit_r224_c121 bl[121] br[121] wl[224] vdd gnd cell_6t
Xbit_r225_c121 bl[121] br[121] wl[225] vdd gnd cell_6t
Xbit_r226_c121 bl[121] br[121] wl[226] vdd gnd cell_6t
Xbit_r227_c121 bl[121] br[121] wl[227] vdd gnd cell_6t
Xbit_r228_c121 bl[121] br[121] wl[228] vdd gnd cell_6t
Xbit_r229_c121 bl[121] br[121] wl[229] vdd gnd cell_6t
Xbit_r230_c121 bl[121] br[121] wl[230] vdd gnd cell_6t
Xbit_r231_c121 bl[121] br[121] wl[231] vdd gnd cell_6t
Xbit_r232_c121 bl[121] br[121] wl[232] vdd gnd cell_6t
Xbit_r233_c121 bl[121] br[121] wl[233] vdd gnd cell_6t
Xbit_r234_c121 bl[121] br[121] wl[234] vdd gnd cell_6t
Xbit_r235_c121 bl[121] br[121] wl[235] vdd gnd cell_6t
Xbit_r236_c121 bl[121] br[121] wl[236] vdd gnd cell_6t
Xbit_r237_c121 bl[121] br[121] wl[237] vdd gnd cell_6t
Xbit_r238_c121 bl[121] br[121] wl[238] vdd gnd cell_6t
Xbit_r239_c121 bl[121] br[121] wl[239] vdd gnd cell_6t
Xbit_r240_c121 bl[121] br[121] wl[240] vdd gnd cell_6t
Xbit_r241_c121 bl[121] br[121] wl[241] vdd gnd cell_6t
Xbit_r242_c121 bl[121] br[121] wl[242] vdd gnd cell_6t
Xbit_r243_c121 bl[121] br[121] wl[243] vdd gnd cell_6t
Xbit_r244_c121 bl[121] br[121] wl[244] vdd gnd cell_6t
Xbit_r245_c121 bl[121] br[121] wl[245] vdd gnd cell_6t
Xbit_r246_c121 bl[121] br[121] wl[246] vdd gnd cell_6t
Xbit_r247_c121 bl[121] br[121] wl[247] vdd gnd cell_6t
Xbit_r248_c121 bl[121] br[121] wl[248] vdd gnd cell_6t
Xbit_r249_c121 bl[121] br[121] wl[249] vdd gnd cell_6t
Xbit_r250_c121 bl[121] br[121] wl[250] vdd gnd cell_6t
Xbit_r251_c121 bl[121] br[121] wl[251] vdd gnd cell_6t
Xbit_r252_c121 bl[121] br[121] wl[252] vdd gnd cell_6t
Xbit_r253_c121 bl[121] br[121] wl[253] vdd gnd cell_6t
Xbit_r254_c121 bl[121] br[121] wl[254] vdd gnd cell_6t
Xbit_r255_c121 bl[121] br[121] wl[255] vdd gnd cell_6t
Xbit_r256_c121 bl[121] br[121] wl[256] vdd gnd cell_6t
Xbit_r257_c121 bl[121] br[121] wl[257] vdd gnd cell_6t
Xbit_r258_c121 bl[121] br[121] wl[258] vdd gnd cell_6t
Xbit_r259_c121 bl[121] br[121] wl[259] vdd gnd cell_6t
Xbit_r260_c121 bl[121] br[121] wl[260] vdd gnd cell_6t
Xbit_r261_c121 bl[121] br[121] wl[261] vdd gnd cell_6t
Xbit_r262_c121 bl[121] br[121] wl[262] vdd gnd cell_6t
Xbit_r263_c121 bl[121] br[121] wl[263] vdd gnd cell_6t
Xbit_r264_c121 bl[121] br[121] wl[264] vdd gnd cell_6t
Xbit_r265_c121 bl[121] br[121] wl[265] vdd gnd cell_6t
Xbit_r266_c121 bl[121] br[121] wl[266] vdd gnd cell_6t
Xbit_r267_c121 bl[121] br[121] wl[267] vdd gnd cell_6t
Xbit_r268_c121 bl[121] br[121] wl[268] vdd gnd cell_6t
Xbit_r269_c121 bl[121] br[121] wl[269] vdd gnd cell_6t
Xbit_r270_c121 bl[121] br[121] wl[270] vdd gnd cell_6t
Xbit_r271_c121 bl[121] br[121] wl[271] vdd gnd cell_6t
Xbit_r272_c121 bl[121] br[121] wl[272] vdd gnd cell_6t
Xbit_r273_c121 bl[121] br[121] wl[273] vdd gnd cell_6t
Xbit_r274_c121 bl[121] br[121] wl[274] vdd gnd cell_6t
Xbit_r275_c121 bl[121] br[121] wl[275] vdd gnd cell_6t
Xbit_r276_c121 bl[121] br[121] wl[276] vdd gnd cell_6t
Xbit_r277_c121 bl[121] br[121] wl[277] vdd gnd cell_6t
Xbit_r278_c121 bl[121] br[121] wl[278] vdd gnd cell_6t
Xbit_r279_c121 bl[121] br[121] wl[279] vdd gnd cell_6t
Xbit_r280_c121 bl[121] br[121] wl[280] vdd gnd cell_6t
Xbit_r281_c121 bl[121] br[121] wl[281] vdd gnd cell_6t
Xbit_r282_c121 bl[121] br[121] wl[282] vdd gnd cell_6t
Xbit_r283_c121 bl[121] br[121] wl[283] vdd gnd cell_6t
Xbit_r284_c121 bl[121] br[121] wl[284] vdd gnd cell_6t
Xbit_r285_c121 bl[121] br[121] wl[285] vdd gnd cell_6t
Xbit_r286_c121 bl[121] br[121] wl[286] vdd gnd cell_6t
Xbit_r287_c121 bl[121] br[121] wl[287] vdd gnd cell_6t
Xbit_r288_c121 bl[121] br[121] wl[288] vdd gnd cell_6t
Xbit_r289_c121 bl[121] br[121] wl[289] vdd gnd cell_6t
Xbit_r290_c121 bl[121] br[121] wl[290] vdd gnd cell_6t
Xbit_r291_c121 bl[121] br[121] wl[291] vdd gnd cell_6t
Xbit_r292_c121 bl[121] br[121] wl[292] vdd gnd cell_6t
Xbit_r293_c121 bl[121] br[121] wl[293] vdd gnd cell_6t
Xbit_r294_c121 bl[121] br[121] wl[294] vdd gnd cell_6t
Xbit_r295_c121 bl[121] br[121] wl[295] vdd gnd cell_6t
Xbit_r296_c121 bl[121] br[121] wl[296] vdd gnd cell_6t
Xbit_r297_c121 bl[121] br[121] wl[297] vdd gnd cell_6t
Xbit_r298_c121 bl[121] br[121] wl[298] vdd gnd cell_6t
Xbit_r299_c121 bl[121] br[121] wl[299] vdd gnd cell_6t
Xbit_r300_c121 bl[121] br[121] wl[300] vdd gnd cell_6t
Xbit_r301_c121 bl[121] br[121] wl[301] vdd gnd cell_6t
Xbit_r302_c121 bl[121] br[121] wl[302] vdd gnd cell_6t
Xbit_r303_c121 bl[121] br[121] wl[303] vdd gnd cell_6t
Xbit_r304_c121 bl[121] br[121] wl[304] vdd gnd cell_6t
Xbit_r305_c121 bl[121] br[121] wl[305] vdd gnd cell_6t
Xbit_r306_c121 bl[121] br[121] wl[306] vdd gnd cell_6t
Xbit_r307_c121 bl[121] br[121] wl[307] vdd gnd cell_6t
Xbit_r308_c121 bl[121] br[121] wl[308] vdd gnd cell_6t
Xbit_r309_c121 bl[121] br[121] wl[309] vdd gnd cell_6t
Xbit_r310_c121 bl[121] br[121] wl[310] vdd gnd cell_6t
Xbit_r311_c121 bl[121] br[121] wl[311] vdd gnd cell_6t
Xbit_r312_c121 bl[121] br[121] wl[312] vdd gnd cell_6t
Xbit_r313_c121 bl[121] br[121] wl[313] vdd gnd cell_6t
Xbit_r314_c121 bl[121] br[121] wl[314] vdd gnd cell_6t
Xbit_r315_c121 bl[121] br[121] wl[315] vdd gnd cell_6t
Xbit_r316_c121 bl[121] br[121] wl[316] vdd gnd cell_6t
Xbit_r317_c121 bl[121] br[121] wl[317] vdd gnd cell_6t
Xbit_r318_c121 bl[121] br[121] wl[318] vdd gnd cell_6t
Xbit_r319_c121 bl[121] br[121] wl[319] vdd gnd cell_6t
Xbit_r320_c121 bl[121] br[121] wl[320] vdd gnd cell_6t
Xbit_r321_c121 bl[121] br[121] wl[321] vdd gnd cell_6t
Xbit_r322_c121 bl[121] br[121] wl[322] vdd gnd cell_6t
Xbit_r323_c121 bl[121] br[121] wl[323] vdd gnd cell_6t
Xbit_r324_c121 bl[121] br[121] wl[324] vdd gnd cell_6t
Xbit_r325_c121 bl[121] br[121] wl[325] vdd gnd cell_6t
Xbit_r326_c121 bl[121] br[121] wl[326] vdd gnd cell_6t
Xbit_r327_c121 bl[121] br[121] wl[327] vdd gnd cell_6t
Xbit_r328_c121 bl[121] br[121] wl[328] vdd gnd cell_6t
Xbit_r329_c121 bl[121] br[121] wl[329] vdd gnd cell_6t
Xbit_r330_c121 bl[121] br[121] wl[330] vdd gnd cell_6t
Xbit_r331_c121 bl[121] br[121] wl[331] vdd gnd cell_6t
Xbit_r332_c121 bl[121] br[121] wl[332] vdd gnd cell_6t
Xbit_r333_c121 bl[121] br[121] wl[333] vdd gnd cell_6t
Xbit_r334_c121 bl[121] br[121] wl[334] vdd gnd cell_6t
Xbit_r335_c121 bl[121] br[121] wl[335] vdd gnd cell_6t
Xbit_r336_c121 bl[121] br[121] wl[336] vdd gnd cell_6t
Xbit_r337_c121 bl[121] br[121] wl[337] vdd gnd cell_6t
Xbit_r338_c121 bl[121] br[121] wl[338] vdd gnd cell_6t
Xbit_r339_c121 bl[121] br[121] wl[339] vdd gnd cell_6t
Xbit_r340_c121 bl[121] br[121] wl[340] vdd gnd cell_6t
Xbit_r341_c121 bl[121] br[121] wl[341] vdd gnd cell_6t
Xbit_r342_c121 bl[121] br[121] wl[342] vdd gnd cell_6t
Xbit_r343_c121 bl[121] br[121] wl[343] vdd gnd cell_6t
Xbit_r344_c121 bl[121] br[121] wl[344] vdd gnd cell_6t
Xbit_r345_c121 bl[121] br[121] wl[345] vdd gnd cell_6t
Xbit_r346_c121 bl[121] br[121] wl[346] vdd gnd cell_6t
Xbit_r347_c121 bl[121] br[121] wl[347] vdd gnd cell_6t
Xbit_r348_c121 bl[121] br[121] wl[348] vdd gnd cell_6t
Xbit_r349_c121 bl[121] br[121] wl[349] vdd gnd cell_6t
Xbit_r350_c121 bl[121] br[121] wl[350] vdd gnd cell_6t
Xbit_r351_c121 bl[121] br[121] wl[351] vdd gnd cell_6t
Xbit_r352_c121 bl[121] br[121] wl[352] vdd gnd cell_6t
Xbit_r353_c121 bl[121] br[121] wl[353] vdd gnd cell_6t
Xbit_r354_c121 bl[121] br[121] wl[354] vdd gnd cell_6t
Xbit_r355_c121 bl[121] br[121] wl[355] vdd gnd cell_6t
Xbit_r356_c121 bl[121] br[121] wl[356] vdd gnd cell_6t
Xbit_r357_c121 bl[121] br[121] wl[357] vdd gnd cell_6t
Xbit_r358_c121 bl[121] br[121] wl[358] vdd gnd cell_6t
Xbit_r359_c121 bl[121] br[121] wl[359] vdd gnd cell_6t
Xbit_r360_c121 bl[121] br[121] wl[360] vdd gnd cell_6t
Xbit_r361_c121 bl[121] br[121] wl[361] vdd gnd cell_6t
Xbit_r362_c121 bl[121] br[121] wl[362] vdd gnd cell_6t
Xbit_r363_c121 bl[121] br[121] wl[363] vdd gnd cell_6t
Xbit_r364_c121 bl[121] br[121] wl[364] vdd gnd cell_6t
Xbit_r365_c121 bl[121] br[121] wl[365] vdd gnd cell_6t
Xbit_r366_c121 bl[121] br[121] wl[366] vdd gnd cell_6t
Xbit_r367_c121 bl[121] br[121] wl[367] vdd gnd cell_6t
Xbit_r368_c121 bl[121] br[121] wl[368] vdd gnd cell_6t
Xbit_r369_c121 bl[121] br[121] wl[369] vdd gnd cell_6t
Xbit_r370_c121 bl[121] br[121] wl[370] vdd gnd cell_6t
Xbit_r371_c121 bl[121] br[121] wl[371] vdd gnd cell_6t
Xbit_r372_c121 bl[121] br[121] wl[372] vdd gnd cell_6t
Xbit_r373_c121 bl[121] br[121] wl[373] vdd gnd cell_6t
Xbit_r374_c121 bl[121] br[121] wl[374] vdd gnd cell_6t
Xbit_r375_c121 bl[121] br[121] wl[375] vdd gnd cell_6t
Xbit_r376_c121 bl[121] br[121] wl[376] vdd gnd cell_6t
Xbit_r377_c121 bl[121] br[121] wl[377] vdd gnd cell_6t
Xbit_r378_c121 bl[121] br[121] wl[378] vdd gnd cell_6t
Xbit_r379_c121 bl[121] br[121] wl[379] vdd gnd cell_6t
Xbit_r380_c121 bl[121] br[121] wl[380] vdd gnd cell_6t
Xbit_r381_c121 bl[121] br[121] wl[381] vdd gnd cell_6t
Xbit_r382_c121 bl[121] br[121] wl[382] vdd gnd cell_6t
Xbit_r383_c121 bl[121] br[121] wl[383] vdd gnd cell_6t
Xbit_r384_c121 bl[121] br[121] wl[384] vdd gnd cell_6t
Xbit_r385_c121 bl[121] br[121] wl[385] vdd gnd cell_6t
Xbit_r386_c121 bl[121] br[121] wl[386] vdd gnd cell_6t
Xbit_r387_c121 bl[121] br[121] wl[387] vdd gnd cell_6t
Xbit_r388_c121 bl[121] br[121] wl[388] vdd gnd cell_6t
Xbit_r389_c121 bl[121] br[121] wl[389] vdd gnd cell_6t
Xbit_r390_c121 bl[121] br[121] wl[390] vdd gnd cell_6t
Xbit_r391_c121 bl[121] br[121] wl[391] vdd gnd cell_6t
Xbit_r392_c121 bl[121] br[121] wl[392] vdd gnd cell_6t
Xbit_r393_c121 bl[121] br[121] wl[393] vdd gnd cell_6t
Xbit_r394_c121 bl[121] br[121] wl[394] vdd gnd cell_6t
Xbit_r395_c121 bl[121] br[121] wl[395] vdd gnd cell_6t
Xbit_r396_c121 bl[121] br[121] wl[396] vdd gnd cell_6t
Xbit_r397_c121 bl[121] br[121] wl[397] vdd gnd cell_6t
Xbit_r398_c121 bl[121] br[121] wl[398] vdd gnd cell_6t
Xbit_r399_c121 bl[121] br[121] wl[399] vdd gnd cell_6t
Xbit_r400_c121 bl[121] br[121] wl[400] vdd gnd cell_6t
Xbit_r401_c121 bl[121] br[121] wl[401] vdd gnd cell_6t
Xbit_r402_c121 bl[121] br[121] wl[402] vdd gnd cell_6t
Xbit_r403_c121 bl[121] br[121] wl[403] vdd gnd cell_6t
Xbit_r404_c121 bl[121] br[121] wl[404] vdd gnd cell_6t
Xbit_r405_c121 bl[121] br[121] wl[405] vdd gnd cell_6t
Xbit_r406_c121 bl[121] br[121] wl[406] vdd gnd cell_6t
Xbit_r407_c121 bl[121] br[121] wl[407] vdd gnd cell_6t
Xbit_r408_c121 bl[121] br[121] wl[408] vdd gnd cell_6t
Xbit_r409_c121 bl[121] br[121] wl[409] vdd gnd cell_6t
Xbit_r410_c121 bl[121] br[121] wl[410] vdd gnd cell_6t
Xbit_r411_c121 bl[121] br[121] wl[411] vdd gnd cell_6t
Xbit_r412_c121 bl[121] br[121] wl[412] vdd gnd cell_6t
Xbit_r413_c121 bl[121] br[121] wl[413] vdd gnd cell_6t
Xbit_r414_c121 bl[121] br[121] wl[414] vdd gnd cell_6t
Xbit_r415_c121 bl[121] br[121] wl[415] vdd gnd cell_6t
Xbit_r416_c121 bl[121] br[121] wl[416] vdd gnd cell_6t
Xbit_r417_c121 bl[121] br[121] wl[417] vdd gnd cell_6t
Xbit_r418_c121 bl[121] br[121] wl[418] vdd gnd cell_6t
Xbit_r419_c121 bl[121] br[121] wl[419] vdd gnd cell_6t
Xbit_r420_c121 bl[121] br[121] wl[420] vdd gnd cell_6t
Xbit_r421_c121 bl[121] br[121] wl[421] vdd gnd cell_6t
Xbit_r422_c121 bl[121] br[121] wl[422] vdd gnd cell_6t
Xbit_r423_c121 bl[121] br[121] wl[423] vdd gnd cell_6t
Xbit_r424_c121 bl[121] br[121] wl[424] vdd gnd cell_6t
Xbit_r425_c121 bl[121] br[121] wl[425] vdd gnd cell_6t
Xbit_r426_c121 bl[121] br[121] wl[426] vdd gnd cell_6t
Xbit_r427_c121 bl[121] br[121] wl[427] vdd gnd cell_6t
Xbit_r428_c121 bl[121] br[121] wl[428] vdd gnd cell_6t
Xbit_r429_c121 bl[121] br[121] wl[429] vdd gnd cell_6t
Xbit_r430_c121 bl[121] br[121] wl[430] vdd gnd cell_6t
Xbit_r431_c121 bl[121] br[121] wl[431] vdd gnd cell_6t
Xbit_r432_c121 bl[121] br[121] wl[432] vdd gnd cell_6t
Xbit_r433_c121 bl[121] br[121] wl[433] vdd gnd cell_6t
Xbit_r434_c121 bl[121] br[121] wl[434] vdd gnd cell_6t
Xbit_r435_c121 bl[121] br[121] wl[435] vdd gnd cell_6t
Xbit_r436_c121 bl[121] br[121] wl[436] vdd gnd cell_6t
Xbit_r437_c121 bl[121] br[121] wl[437] vdd gnd cell_6t
Xbit_r438_c121 bl[121] br[121] wl[438] vdd gnd cell_6t
Xbit_r439_c121 bl[121] br[121] wl[439] vdd gnd cell_6t
Xbit_r440_c121 bl[121] br[121] wl[440] vdd gnd cell_6t
Xbit_r441_c121 bl[121] br[121] wl[441] vdd gnd cell_6t
Xbit_r442_c121 bl[121] br[121] wl[442] vdd gnd cell_6t
Xbit_r443_c121 bl[121] br[121] wl[443] vdd gnd cell_6t
Xbit_r444_c121 bl[121] br[121] wl[444] vdd gnd cell_6t
Xbit_r445_c121 bl[121] br[121] wl[445] vdd gnd cell_6t
Xbit_r446_c121 bl[121] br[121] wl[446] vdd gnd cell_6t
Xbit_r447_c121 bl[121] br[121] wl[447] vdd gnd cell_6t
Xbit_r448_c121 bl[121] br[121] wl[448] vdd gnd cell_6t
Xbit_r449_c121 bl[121] br[121] wl[449] vdd gnd cell_6t
Xbit_r450_c121 bl[121] br[121] wl[450] vdd gnd cell_6t
Xbit_r451_c121 bl[121] br[121] wl[451] vdd gnd cell_6t
Xbit_r452_c121 bl[121] br[121] wl[452] vdd gnd cell_6t
Xbit_r453_c121 bl[121] br[121] wl[453] vdd gnd cell_6t
Xbit_r454_c121 bl[121] br[121] wl[454] vdd gnd cell_6t
Xbit_r455_c121 bl[121] br[121] wl[455] vdd gnd cell_6t
Xbit_r456_c121 bl[121] br[121] wl[456] vdd gnd cell_6t
Xbit_r457_c121 bl[121] br[121] wl[457] vdd gnd cell_6t
Xbit_r458_c121 bl[121] br[121] wl[458] vdd gnd cell_6t
Xbit_r459_c121 bl[121] br[121] wl[459] vdd gnd cell_6t
Xbit_r460_c121 bl[121] br[121] wl[460] vdd gnd cell_6t
Xbit_r461_c121 bl[121] br[121] wl[461] vdd gnd cell_6t
Xbit_r462_c121 bl[121] br[121] wl[462] vdd gnd cell_6t
Xbit_r463_c121 bl[121] br[121] wl[463] vdd gnd cell_6t
Xbit_r464_c121 bl[121] br[121] wl[464] vdd gnd cell_6t
Xbit_r465_c121 bl[121] br[121] wl[465] vdd gnd cell_6t
Xbit_r466_c121 bl[121] br[121] wl[466] vdd gnd cell_6t
Xbit_r467_c121 bl[121] br[121] wl[467] vdd gnd cell_6t
Xbit_r468_c121 bl[121] br[121] wl[468] vdd gnd cell_6t
Xbit_r469_c121 bl[121] br[121] wl[469] vdd gnd cell_6t
Xbit_r470_c121 bl[121] br[121] wl[470] vdd gnd cell_6t
Xbit_r471_c121 bl[121] br[121] wl[471] vdd gnd cell_6t
Xbit_r472_c121 bl[121] br[121] wl[472] vdd gnd cell_6t
Xbit_r473_c121 bl[121] br[121] wl[473] vdd gnd cell_6t
Xbit_r474_c121 bl[121] br[121] wl[474] vdd gnd cell_6t
Xbit_r475_c121 bl[121] br[121] wl[475] vdd gnd cell_6t
Xbit_r476_c121 bl[121] br[121] wl[476] vdd gnd cell_6t
Xbit_r477_c121 bl[121] br[121] wl[477] vdd gnd cell_6t
Xbit_r478_c121 bl[121] br[121] wl[478] vdd gnd cell_6t
Xbit_r479_c121 bl[121] br[121] wl[479] vdd gnd cell_6t
Xbit_r480_c121 bl[121] br[121] wl[480] vdd gnd cell_6t
Xbit_r481_c121 bl[121] br[121] wl[481] vdd gnd cell_6t
Xbit_r482_c121 bl[121] br[121] wl[482] vdd gnd cell_6t
Xbit_r483_c121 bl[121] br[121] wl[483] vdd gnd cell_6t
Xbit_r484_c121 bl[121] br[121] wl[484] vdd gnd cell_6t
Xbit_r485_c121 bl[121] br[121] wl[485] vdd gnd cell_6t
Xbit_r486_c121 bl[121] br[121] wl[486] vdd gnd cell_6t
Xbit_r487_c121 bl[121] br[121] wl[487] vdd gnd cell_6t
Xbit_r488_c121 bl[121] br[121] wl[488] vdd gnd cell_6t
Xbit_r489_c121 bl[121] br[121] wl[489] vdd gnd cell_6t
Xbit_r490_c121 bl[121] br[121] wl[490] vdd gnd cell_6t
Xbit_r491_c121 bl[121] br[121] wl[491] vdd gnd cell_6t
Xbit_r492_c121 bl[121] br[121] wl[492] vdd gnd cell_6t
Xbit_r493_c121 bl[121] br[121] wl[493] vdd gnd cell_6t
Xbit_r494_c121 bl[121] br[121] wl[494] vdd gnd cell_6t
Xbit_r495_c121 bl[121] br[121] wl[495] vdd gnd cell_6t
Xbit_r496_c121 bl[121] br[121] wl[496] vdd gnd cell_6t
Xbit_r497_c121 bl[121] br[121] wl[497] vdd gnd cell_6t
Xbit_r498_c121 bl[121] br[121] wl[498] vdd gnd cell_6t
Xbit_r499_c121 bl[121] br[121] wl[499] vdd gnd cell_6t
Xbit_r500_c121 bl[121] br[121] wl[500] vdd gnd cell_6t
Xbit_r501_c121 bl[121] br[121] wl[501] vdd gnd cell_6t
Xbit_r502_c121 bl[121] br[121] wl[502] vdd gnd cell_6t
Xbit_r503_c121 bl[121] br[121] wl[503] vdd gnd cell_6t
Xbit_r504_c121 bl[121] br[121] wl[504] vdd gnd cell_6t
Xbit_r505_c121 bl[121] br[121] wl[505] vdd gnd cell_6t
Xbit_r506_c121 bl[121] br[121] wl[506] vdd gnd cell_6t
Xbit_r507_c121 bl[121] br[121] wl[507] vdd gnd cell_6t
Xbit_r508_c121 bl[121] br[121] wl[508] vdd gnd cell_6t
Xbit_r509_c121 bl[121] br[121] wl[509] vdd gnd cell_6t
Xbit_r510_c121 bl[121] br[121] wl[510] vdd gnd cell_6t
Xbit_r511_c121 bl[121] br[121] wl[511] vdd gnd cell_6t
Xbit_r0_c122 bl[122] br[122] wl[0] vdd gnd cell_6t
Xbit_r1_c122 bl[122] br[122] wl[1] vdd gnd cell_6t
Xbit_r2_c122 bl[122] br[122] wl[2] vdd gnd cell_6t
Xbit_r3_c122 bl[122] br[122] wl[3] vdd gnd cell_6t
Xbit_r4_c122 bl[122] br[122] wl[4] vdd gnd cell_6t
Xbit_r5_c122 bl[122] br[122] wl[5] vdd gnd cell_6t
Xbit_r6_c122 bl[122] br[122] wl[6] vdd gnd cell_6t
Xbit_r7_c122 bl[122] br[122] wl[7] vdd gnd cell_6t
Xbit_r8_c122 bl[122] br[122] wl[8] vdd gnd cell_6t
Xbit_r9_c122 bl[122] br[122] wl[9] vdd gnd cell_6t
Xbit_r10_c122 bl[122] br[122] wl[10] vdd gnd cell_6t
Xbit_r11_c122 bl[122] br[122] wl[11] vdd gnd cell_6t
Xbit_r12_c122 bl[122] br[122] wl[12] vdd gnd cell_6t
Xbit_r13_c122 bl[122] br[122] wl[13] vdd gnd cell_6t
Xbit_r14_c122 bl[122] br[122] wl[14] vdd gnd cell_6t
Xbit_r15_c122 bl[122] br[122] wl[15] vdd gnd cell_6t
Xbit_r16_c122 bl[122] br[122] wl[16] vdd gnd cell_6t
Xbit_r17_c122 bl[122] br[122] wl[17] vdd gnd cell_6t
Xbit_r18_c122 bl[122] br[122] wl[18] vdd gnd cell_6t
Xbit_r19_c122 bl[122] br[122] wl[19] vdd gnd cell_6t
Xbit_r20_c122 bl[122] br[122] wl[20] vdd gnd cell_6t
Xbit_r21_c122 bl[122] br[122] wl[21] vdd gnd cell_6t
Xbit_r22_c122 bl[122] br[122] wl[22] vdd gnd cell_6t
Xbit_r23_c122 bl[122] br[122] wl[23] vdd gnd cell_6t
Xbit_r24_c122 bl[122] br[122] wl[24] vdd gnd cell_6t
Xbit_r25_c122 bl[122] br[122] wl[25] vdd gnd cell_6t
Xbit_r26_c122 bl[122] br[122] wl[26] vdd gnd cell_6t
Xbit_r27_c122 bl[122] br[122] wl[27] vdd gnd cell_6t
Xbit_r28_c122 bl[122] br[122] wl[28] vdd gnd cell_6t
Xbit_r29_c122 bl[122] br[122] wl[29] vdd gnd cell_6t
Xbit_r30_c122 bl[122] br[122] wl[30] vdd gnd cell_6t
Xbit_r31_c122 bl[122] br[122] wl[31] vdd gnd cell_6t
Xbit_r32_c122 bl[122] br[122] wl[32] vdd gnd cell_6t
Xbit_r33_c122 bl[122] br[122] wl[33] vdd gnd cell_6t
Xbit_r34_c122 bl[122] br[122] wl[34] vdd gnd cell_6t
Xbit_r35_c122 bl[122] br[122] wl[35] vdd gnd cell_6t
Xbit_r36_c122 bl[122] br[122] wl[36] vdd gnd cell_6t
Xbit_r37_c122 bl[122] br[122] wl[37] vdd gnd cell_6t
Xbit_r38_c122 bl[122] br[122] wl[38] vdd gnd cell_6t
Xbit_r39_c122 bl[122] br[122] wl[39] vdd gnd cell_6t
Xbit_r40_c122 bl[122] br[122] wl[40] vdd gnd cell_6t
Xbit_r41_c122 bl[122] br[122] wl[41] vdd gnd cell_6t
Xbit_r42_c122 bl[122] br[122] wl[42] vdd gnd cell_6t
Xbit_r43_c122 bl[122] br[122] wl[43] vdd gnd cell_6t
Xbit_r44_c122 bl[122] br[122] wl[44] vdd gnd cell_6t
Xbit_r45_c122 bl[122] br[122] wl[45] vdd gnd cell_6t
Xbit_r46_c122 bl[122] br[122] wl[46] vdd gnd cell_6t
Xbit_r47_c122 bl[122] br[122] wl[47] vdd gnd cell_6t
Xbit_r48_c122 bl[122] br[122] wl[48] vdd gnd cell_6t
Xbit_r49_c122 bl[122] br[122] wl[49] vdd gnd cell_6t
Xbit_r50_c122 bl[122] br[122] wl[50] vdd gnd cell_6t
Xbit_r51_c122 bl[122] br[122] wl[51] vdd gnd cell_6t
Xbit_r52_c122 bl[122] br[122] wl[52] vdd gnd cell_6t
Xbit_r53_c122 bl[122] br[122] wl[53] vdd gnd cell_6t
Xbit_r54_c122 bl[122] br[122] wl[54] vdd gnd cell_6t
Xbit_r55_c122 bl[122] br[122] wl[55] vdd gnd cell_6t
Xbit_r56_c122 bl[122] br[122] wl[56] vdd gnd cell_6t
Xbit_r57_c122 bl[122] br[122] wl[57] vdd gnd cell_6t
Xbit_r58_c122 bl[122] br[122] wl[58] vdd gnd cell_6t
Xbit_r59_c122 bl[122] br[122] wl[59] vdd gnd cell_6t
Xbit_r60_c122 bl[122] br[122] wl[60] vdd gnd cell_6t
Xbit_r61_c122 bl[122] br[122] wl[61] vdd gnd cell_6t
Xbit_r62_c122 bl[122] br[122] wl[62] vdd gnd cell_6t
Xbit_r63_c122 bl[122] br[122] wl[63] vdd gnd cell_6t
Xbit_r64_c122 bl[122] br[122] wl[64] vdd gnd cell_6t
Xbit_r65_c122 bl[122] br[122] wl[65] vdd gnd cell_6t
Xbit_r66_c122 bl[122] br[122] wl[66] vdd gnd cell_6t
Xbit_r67_c122 bl[122] br[122] wl[67] vdd gnd cell_6t
Xbit_r68_c122 bl[122] br[122] wl[68] vdd gnd cell_6t
Xbit_r69_c122 bl[122] br[122] wl[69] vdd gnd cell_6t
Xbit_r70_c122 bl[122] br[122] wl[70] vdd gnd cell_6t
Xbit_r71_c122 bl[122] br[122] wl[71] vdd gnd cell_6t
Xbit_r72_c122 bl[122] br[122] wl[72] vdd gnd cell_6t
Xbit_r73_c122 bl[122] br[122] wl[73] vdd gnd cell_6t
Xbit_r74_c122 bl[122] br[122] wl[74] vdd gnd cell_6t
Xbit_r75_c122 bl[122] br[122] wl[75] vdd gnd cell_6t
Xbit_r76_c122 bl[122] br[122] wl[76] vdd gnd cell_6t
Xbit_r77_c122 bl[122] br[122] wl[77] vdd gnd cell_6t
Xbit_r78_c122 bl[122] br[122] wl[78] vdd gnd cell_6t
Xbit_r79_c122 bl[122] br[122] wl[79] vdd gnd cell_6t
Xbit_r80_c122 bl[122] br[122] wl[80] vdd gnd cell_6t
Xbit_r81_c122 bl[122] br[122] wl[81] vdd gnd cell_6t
Xbit_r82_c122 bl[122] br[122] wl[82] vdd gnd cell_6t
Xbit_r83_c122 bl[122] br[122] wl[83] vdd gnd cell_6t
Xbit_r84_c122 bl[122] br[122] wl[84] vdd gnd cell_6t
Xbit_r85_c122 bl[122] br[122] wl[85] vdd gnd cell_6t
Xbit_r86_c122 bl[122] br[122] wl[86] vdd gnd cell_6t
Xbit_r87_c122 bl[122] br[122] wl[87] vdd gnd cell_6t
Xbit_r88_c122 bl[122] br[122] wl[88] vdd gnd cell_6t
Xbit_r89_c122 bl[122] br[122] wl[89] vdd gnd cell_6t
Xbit_r90_c122 bl[122] br[122] wl[90] vdd gnd cell_6t
Xbit_r91_c122 bl[122] br[122] wl[91] vdd gnd cell_6t
Xbit_r92_c122 bl[122] br[122] wl[92] vdd gnd cell_6t
Xbit_r93_c122 bl[122] br[122] wl[93] vdd gnd cell_6t
Xbit_r94_c122 bl[122] br[122] wl[94] vdd gnd cell_6t
Xbit_r95_c122 bl[122] br[122] wl[95] vdd gnd cell_6t
Xbit_r96_c122 bl[122] br[122] wl[96] vdd gnd cell_6t
Xbit_r97_c122 bl[122] br[122] wl[97] vdd gnd cell_6t
Xbit_r98_c122 bl[122] br[122] wl[98] vdd gnd cell_6t
Xbit_r99_c122 bl[122] br[122] wl[99] vdd gnd cell_6t
Xbit_r100_c122 bl[122] br[122] wl[100] vdd gnd cell_6t
Xbit_r101_c122 bl[122] br[122] wl[101] vdd gnd cell_6t
Xbit_r102_c122 bl[122] br[122] wl[102] vdd gnd cell_6t
Xbit_r103_c122 bl[122] br[122] wl[103] vdd gnd cell_6t
Xbit_r104_c122 bl[122] br[122] wl[104] vdd gnd cell_6t
Xbit_r105_c122 bl[122] br[122] wl[105] vdd gnd cell_6t
Xbit_r106_c122 bl[122] br[122] wl[106] vdd gnd cell_6t
Xbit_r107_c122 bl[122] br[122] wl[107] vdd gnd cell_6t
Xbit_r108_c122 bl[122] br[122] wl[108] vdd gnd cell_6t
Xbit_r109_c122 bl[122] br[122] wl[109] vdd gnd cell_6t
Xbit_r110_c122 bl[122] br[122] wl[110] vdd gnd cell_6t
Xbit_r111_c122 bl[122] br[122] wl[111] vdd gnd cell_6t
Xbit_r112_c122 bl[122] br[122] wl[112] vdd gnd cell_6t
Xbit_r113_c122 bl[122] br[122] wl[113] vdd gnd cell_6t
Xbit_r114_c122 bl[122] br[122] wl[114] vdd gnd cell_6t
Xbit_r115_c122 bl[122] br[122] wl[115] vdd gnd cell_6t
Xbit_r116_c122 bl[122] br[122] wl[116] vdd gnd cell_6t
Xbit_r117_c122 bl[122] br[122] wl[117] vdd gnd cell_6t
Xbit_r118_c122 bl[122] br[122] wl[118] vdd gnd cell_6t
Xbit_r119_c122 bl[122] br[122] wl[119] vdd gnd cell_6t
Xbit_r120_c122 bl[122] br[122] wl[120] vdd gnd cell_6t
Xbit_r121_c122 bl[122] br[122] wl[121] vdd gnd cell_6t
Xbit_r122_c122 bl[122] br[122] wl[122] vdd gnd cell_6t
Xbit_r123_c122 bl[122] br[122] wl[123] vdd gnd cell_6t
Xbit_r124_c122 bl[122] br[122] wl[124] vdd gnd cell_6t
Xbit_r125_c122 bl[122] br[122] wl[125] vdd gnd cell_6t
Xbit_r126_c122 bl[122] br[122] wl[126] vdd gnd cell_6t
Xbit_r127_c122 bl[122] br[122] wl[127] vdd gnd cell_6t
Xbit_r128_c122 bl[122] br[122] wl[128] vdd gnd cell_6t
Xbit_r129_c122 bl[122] br[122] wl[129] vdd gnd cell_6t
Xbit_r130_c122 bl[122] br[122] wl[130] vdd gnd cell_6t
Xbit_r131_c122 bl[122] br[122] wl[131] vdd gnd cell_6t
Xbit_r132_c122 bl[122] br[122] wl[132] vdd gnd cell_6t
Xbit_r133_c122 bl[122] br[122] wl[133] vdd gnd cell_6t
Xbit_r134_c122 bl[122] br[122] wl[134] vdd gnd cell_6t
Xbit_r135_c122 bl[122] br[122] wl[135] vdd gnd cell_6t
Xbit_r136_c122 bl[122] br[122] wl[136] vdd gnd cell_6t
Xbit_r137_c122 bl[122] br[122] wl[137] vdd gnd cell_6t
Xbit_r138_c122 bl[122] br[122] wl[138] vdd gnd cell_6t
Xbit_r139_c122 bl[122] br[122] wl[139] vdd gnd cell_6t
Xbit_r140_c122 bl[122] br[122] wl[140] vdd gnd cell_6t
Xbit_r141_c122 bl[122] br[122] wl[141] vdd gnd cell_6t
Xbit_r142_c122 bl[122] br[122] wl[142] vdd gnd cell_6t
Xbit_r143_c122 bl[122] br[122] wl[143] vdd gnd cell_6t
Xbit_r144_c122 bl[122] br[122] wl[144] vdd gnd cell_6t
Xbit_r145_c122 bl[122] br[122] wl[145] vdd gnd cell_6t
Xbit_r146_c122 bl[122] br[122] wl[146] vdd gnd cell_6t
Xbit_r147_c122 bl[122] br[122] wl[147] vdd gnd cell_6t
Xbit_r148_c122 bl[122] br[122] wl[148] vdd gnd cell_6t
Xbit_r149_c122 bl[122] br[122] wl[149] vdd gnd cell_6t
Xbit_r150_c122 bl[122] br[122] wl[150] vdd gnd cell_6t
Xbit_r151_c122 bl[122] br[122] wl[151] vdd gnd cell_6t
Xbit_r152_c122 bl[122] br[122] wl[152] vdd gnd cell_6t
Xbit_r153_c122 bl[122] br[122] wl[153] vdd gnd cell_6t
Xbit_r154_c122 bl[122] br[122] wl[154] vdd gnd cell_6t
Xbit_r155_c122 bl[122] br[122] wl[155] vdd gnd cell_6t
Xbit_r156_c122 bl[122] br[122] wl[156] vdd gnd cell_6t
Xbit_r157_c122 bl[122] br[122] wl[157] vdd gnd cell_6t
Xbit_r158_c122 bl[122] br[122] wl[158] vdd gnd cell_6t
Xbit_r159_c122 bl[122] br[122] wl[159] vdd gnd cell_6t
Xbit_r160_c122 bl[122] br[122] wl[160] vdd gnd cell_6t
Xbit_r161_c122 bl[122] br[122] wl[161] vdd gnd cell_6t
Xbit_r162_c122 bl[122] br[122] wl[162] vdd gnd cell_6t
Xbit_r163_c122 bl[122] br[122] wl[163] vdd gnd cell_6t
Xbit_r164_c122 bl[122] br[122] wl[164] vdd gnd cell_6t
Xbit_r165_c122 bl[122] br[122] wl[165] vdd gnd cell_6t
Xbit_r166_c122 bl[122] br[122] wl[166] vdd gnd cell_6t
Xbit_r167_c122 bl[122] br[122] wl[167] vdd gnd cell_6t
Xbit_r168_c122 bl[122] br[122] wl[168] vdd gnd cell_6t
Xbit_r169_c122 bl[122] br[122] wl[169] vdd gnd cell_6t
Xbit_r170_c122 bl[122] br[122] wl[170] vdd gnd cell_6t
Xbit_r171_c122 bl[122] br[122] wl[171] vdd gnd cell_6t
Xbit_r172_c122 bl[122] br[122] wl[172] vdd gnd cell_6t
Xbit_r173_c122 bl[122] br[122] wl[173] vdd gnd cell_6t
Xbit_r174_c122 bl[122] br[122] wl[174] vdd gnd cell_6t
Xbit_r175_c122 bl[122] br[122] wl[175] vdd gnd cell_6t
Xbit_r176_c122 bl[122] br[122] wl[176] vdd gnd cell_6t
Xbit_r177_c122 bl[122] br[122] wl[177] vdd gnd cell_6t
Xbit_r178_c122 bl[122] br[122] wl[178] vdd gnd cell_6t
Xbit_r179_c122 bl[122] br[122] wl[179] vdd gnd cell_6t
Xbit_r180_c122 bl[122] br[122] wl[180] vdd gnd cell_6t
Xbit_r181_c122 bl[122] br[122] wl[181] vdd gnd cell_6t
Xbit_r182_c122 bl[122] br[122] wl[182] vdd gnd cell_6t
Xbit_r183_c122 bl[122] br[122] wl[183] vdd gnd cell_6t
Xbit_r184_c122 bl[122] br[122] wl[184] vdd gnd cell_6t
Xbit_r185_c122 bl[122] br[122] wl[185] vdd gnd cell_6t
Xbit_r186_c122 bl[122] br[122] wl[186] vdd gnd cell_6t
Xbit_r187_c122 bl[122] br[122] wl[187] vdd gnd cell_6t
Xbit_r188_c122 bl[122] br[122] wl[188] vdd gnd cell_6t
Xbit_r189_c122 bl[122] br[122] wl[189] vdd gnd cell_6t
Xbit_r190_c122 bl[122] br[122] wl[190] vdd gnd cell_6t
Xbit_r191_c122 bl[122] br[122] wl[191] vdd gnd cell_6t
Xbit_r192_c122 bl[122] br[122] wl[192] vdd gnd cell_6t
Xbit_r193_c122 bl[122] br[122] wl[193] vdd gnd cell_6t
Xbit_r194_c122 bl[122] br[122] wl[194] vdd gnd cell_6t
Xbit_r195_c122 bl[122] br[122] wl[195] vdd gnd cell_6t
Xbit_r196_c122 bl[122] br[122] wl[196] vdd gnd cell_6t
Xbit_r197_c122 bl[122] br[122] wl[197] vdd gnd cell_6t
Xbit_r198_c122 bl[122] br[122] wl[198] vdd gnd cell_6t
Xbit_r199_c122 bl[122] br[122] wl[199] vdd gnd cell_6t
Xbit_r200_c122 bl[122] br[122] wl[200] vdd gnd cell_6t
Xbit_r201_c122 bl[122] br[122] wl[201] vdd gnd cell_6t
Xbit_r202_c122 bl[122] br[122] wl[202] vdd gnd cell_6t
Xbit_r203_c122 bl[122] br[122] wl[203] vdd gnd cell_6t
Xbit_r204_c122 bl[122] br[122] wl[204] vdd gnd cell_6t
Xbit_r205_c122 bl[122] br[122] wl[205] vdd gnd cell_6t
Xbit_r206_c122 bl[122] br[122] wl[206] vdd gnd cell_6t
Xbit_r207_c122 bl[122] br[122] wl[207] vdd gnd cell_6t
Xbit_r208_c122 bl[122] br[122] wl[208] vdd gnd cell_6t
Xbit_r209_c122 bl[122] br[122] wl[209] vdd gnd cell_6t
Xbit_r210_c122 bl[122] br[122] wl[210] vdd gnd cell_6t
Xbit_r211_c122 bl[122] br[122] wl[211] vdd gnd cell_6t
Xbit_r212_c122 bl[122] br[122] wl[212] vdd gnd cell_6t
Xbit_r213_c122 bl[122] br[122] wl[213] vdd gnd cell_6t
Xbit_r214_c122 bl[122] br[122] wl[214] vdd gnd cell_6t
Xbit_r215_c122 bl[122] br[122] wl[215] vdd gnd cell_6t
Xbit_r216_c122 bl[122] br[122] wl[216] vdd gnd cell_6t
Xbit_r217_c122 bl[122] br[122] wl[217] vdd gnd cell_6t
Xbit_r218_c122 bl[122] br[122] wl[218] vdd gnd cell_6t
Xbit_r219_c122 bl[122] br[122] wl[219] vdd gnd cell_6t
Xbit_r220_c122 bl[122] br[122] wl[220] vdd gnd cell_6t
Xbit_r221_c122 bl[122] br[122] wl[221] vdd gnd cell_6t
Xbit_r222_c122 bl[122] br[122] wl[222] vdd gnd cell_6t
Xbit_r223_c122 bl[122] br[122] wl[223] vdd gnd cell_6t
Xbit_r224_c122 bl[122] br[122] wl[224] vdd gnd cell_6t
Xbit_r225_c122 bl[122] br[122] wl[225] vdd gnd cell_6t
Xbit_r226_c122 bl[122] br[122] wl[226] vdd gnd cell_6t
Xbit_r227_c122 bl[122] br[122] wl[227] vdd gnd cell_6t
Xbit_r228_c122 bl[122] br[122] wl[228] vdd gnd cell_6t
Xbit_r229_c122 bl[122] br[122] wl[229] vdd gnd cell_6t
Xbit_r230_c122 bl[122] br[122] wl[230] vdd gnd cell_6t
Xbit_r231_c122 bl[122] br[122] wl[231] vdd gnd cell_6t
Xbit_r232_c122 bl[122] br[122] wl[232] vdd gnd cell_6t
Xbit_r233_c122 bl[122] br[122] wl[233] vdd gnd cell_6t
Xbit_r234_c122 bl[122] br[122] wl[234] vdd gnd cell_6t
Xbit_r235_c122 bl[122] br[122] wl[235] vdd gnd cell_6t
Xbit_r236_c122 bl[122] br[122] wl[236] vdd gnd cell_6t
Xbit_r237_c122 bl[122] br[122] wl[237] vdd gnd cell_6t
Xbit_r238_c122 bl[122] br[122] wl[238] vdd gnd cell_6t
Xbit_r239_c122 bl[122] br[122] wl[239] vdd gnd cell_6t
Xbit_r240_c122 bl[122] br[122] wl[240] vdd gnd cell_6t
Xbit_r241_c122 bl[122] br[122] wl[241] vdd gnd cell_6t
Xbit_r242_c122 bl[122] br[122] wl[242] vdd gnd cell_6t
Xbit_r243_c122 bl[122] br[122] wl[243] vdd gnd cell_6t
Xbit_r244_c122 bl[122] br[122] wl[244] vdd gnd cell_6t
Xbit_r245_c122 bl[122] br[122] wl[245] vdd gnd cell_6t
Xbit_r246_c122 bl[122] br[122] wl[246] vdd gnd cell_6t
Xbit_r247_c122 bl[122] br[122] wl[247] vdd gnd cell_6t
Xbit_r248_c122 bl[122] br[122] wl[248] vdd gnd cell_6t
Xbit_r249_c122 bl[122] br[122] wl[249] vdd gnd cell_6t
Xbit_r250_c122 bl[122] br[122] wl[250] vdd gnd cell_6t
Xbit_r251_c122 bl[122] br[122] wl[251] vdd gnd cell_6t
Xbit_r252_c122 bl[122] br[122] wl[252] vdd gnd cell_6t
Xbit_r253_c122 bl[122] br[122] wl[253] vdd gnd cell_6t
Xbit_r254_c122 bl[122] br[122] wl[254] vdd gnd cell_6t
Xbit_r255_c122 bl[122] br[122] wl[255] vdd gnd cell_6t
Xbit_r256_c122 bl[122] br[122] wl[256] vdd gnd cell_6t
Xbit_r257_c122 bl[122] br[122] wl[257] vdd gnd cell_6t
Xbit_r258_c122 bl[122] br[122] wl[258] vdd gnd cell_6t
Xbit_r259_c122 bl[122] br[122] wl[259] vdd gnd cell_6t
Xbit_r260_c122 bl[122] br[122] wl[260] vdd gnd cell_6t
Xbit_r261_c122 bl[122] br[122] wl[261] vdd gnd cell_6t
Xbit_r262_c122 bl[122] br[122] wl[262] vdd gnd cell_6t
Xbit_r263_c122 bl[122] br[122] wl[263] vdd gnd cell_6t
Xbit_r264_c122 bl[122] br[122] wl[264] vdd gnd cell_6t
Xbit_r265_c122 bl[122] br[122] wl[265] vdd gnd cell_6t
Xbit_r266_c122 bl[122] br[122] wl[266] vdd gnd cell_6t
Xbit_r267_c122 bl[122] br[122] wl[267] vdd gnd cell_6t
Xbit_r268_c122 bl[122] br[122] wl[268] vdd gnd cell_6t
Xbit_r269_c122 bl[122] br[122] wl[269] vdd gnd cell_6t
Xbit_r270_c122 bl[122] br[122] wl[270] vdd gnd cell_6t
Xbit_r271_c122 bl[122] br[122] wl[271] vdd gnd cell_6t
Xbit_r272_c122 bl[122] br[122] wl[272] vdd gnd cell_6t
Xbit_r273_c122 bl[122] br[122] wl[273] vdd gnd cell_6t
Xbit_r274_c122 bl[122] br[122] wl[274] vdd gnd cell_6t
Xbit_r275_c122 bl[122] br[122] wl[275] vdd gnd cell_6t
Xbit_r276_c122 bl[122] br[122] wl[276] vdd gnd cell_6t
Xbit_r277_c122 bl[122] br[122] wl[277] vdd gnd cell_6t
Xbit_r278_c122 bl[122] br[122] wl[278] vdd gnd cell_6t
Xbit_r279_c122 bl[122] br[122] wl[279] vdd gnd cell_6t
Xbit_r280_c122 bl[122] br[122] wl[280] vdd gnd cell_6t
Xbit_r281_c122 bl[122] br[122] wl[281] vdd gnd cell_6t
Xbit_r282_c122 bl[122] br[122] wl[282] vdd gnd cell_6t
Xbit_r283_c122 bl[122] br[122] wl[283] vdd gnd cell_6t
Xbit_r284_c122 bl[122] br[122] wl[284] vdd gnd cell_6t
Xbit_r285_c122 bl[122] br[122] wl[285] vdd gnd cell_6t
Xbit_r286_c122 bl[122] br[122] wl[286] vdd gnd cell_6t
Xbit_r287_c122 bl[122] br[122] wl[287] vdd gnd cell_6t
Xbit_r288_c122 bl[122] br[122] wl[288] vdd gnd cell_6t
Xbit_r289_c122 bl[122] br[122] wl[289] vdd gnd cell_6t
Xbit_r290_c122 bl[122] br[122] wl[290] vdd gnd cell_6t
Xbit_r291_c122 bl[122] br[122] wl[291] vdd gnd cell_6t
Xbit_r292_c122 bl[122] br[122] wl[292] vdd gnd cell_6t
Xbit_r293_c122 bl[122] br[122] wl[293] vdd gnd cell_6t
Xbit_r294_c122 bl[122] br[122] wl[294] vdd gnd cell_6t
Xbit_r295_c122 bl[122] br[122] wl[295] vdd gnd cell_6t
Xbit_r296_c122 bl[122] br[122] wl[296] vdd gnd cell_6t
Xbit_r297_c122 bl[122] br[122] wl[297] vdd gnd cell_6t
Xbit_r298_c122 bl[122] br[122] wl[298] vdd gnd cell_6t
Xbit_r299_c122 bl[122] br[122] wl[299] vdd gnd cell_6t
Xbit_r300_c122 bl[122] br[122] wl[300] vdd gnd cell_6t
Xbit_r301_c122 bl[122] br[122] wl[301] vdd gnd cell_6t
Xbit_r302_c122 bl[122] br[122] wl[302] vdd gnd cell_6t
Xbit_r303_c122 bl[122] br[122] wl[303] vdd gnd cell_6t
Xbit_r304_c122 bl[122] br[122] wl[304] vdd gnd cell_6t
Xbit_r305_c122 bl[122] br[122] wl[305] vdd gnd cell_6t
Xbit_r306_c122 bl[122] br[122] wl[306] vdd gnd cell_6t
Xbit_r307_c122 bl[122] br[122] wl[307] vdd gnd cell_6t
Xbit_r308_c122 bl[122] br[122] wl[308] vdd gnd cell_6t
Xbit_r309_c122 bl[122] br[122] wl[309] vdd gnd cell_6t
Xbit_r310_c122 bl[122] br[122] wl[310] vdd gnd cell_6t
Xbit_r311_c122 bl[122] br[122] wl[311] vdd gnd cell_6t
Xbit_r312_c122 bl[122] br[122] wl[312] vdd gnd cell_6t
Xbit_r313_c122 bl[122] br[122] wl[313] vdd gnd cell_6t
Xbit_r314_c122 bl[122] br[122] wl[314] vdd gnd cell_6t
Xbit_r315_c122 bl[122] br[122] wl[315] vdd gnd cell_6t
Xbit_r316_c122 bl[122] br[122] wl[316] vdd gnd cell_6t
Xbit_r317_c122 bl[122] br[122] wl[317] vdd gnd cell_6t
Xbit_r318_c122 bl[122] br[122] wl[318] vdd gnd cell_6t
Xbit_r319_c122 bl[122] br[122] wl[319] vdd gnd cell_6t
Xbit_r320_c122 bl[122] br[122] wl[320] vdd gnd cell_6t
Xbit_r321_c122 bl[122] br[122] wl[321] vdd gnd cell_6t
Xbit_r322_c122 bl[122] br[122] wl[322] vdd gnd cell_6t
Xbit_r323_c122 bl[122] br[122] wl[323] vdd gnd cell_6t
Xbit_r324_c122 bl[122] br[122] wl[324] vdd gnd cell_6t
Xbit_r325_c122 bl[122] br[122] wl[325] vdd gnd cell_6t
Xbit_r326_c122 bl[122] br[122] wl[326] vdd gnd cell_6t
Xbit_r327_c122 bl[122] br[122] wl[327] vdd gnd cell_6t
Xbit_r328_c122 bl[122] br[122] wl[328] vdd gnd cell_6t
Xbit_r329_c122 bl[122] br[122] wl[329] vdd gnd cell_6t
Xbit_r330_c122 bl[122] br[122] wl[330] vdd gnd cell_6t
Xbit_r331_c122 bl[122] br[122] wl[331] vdd gnd cell_6t
Xbit_r332_c122 bl[122] br[122] wl[332] vdd gnd cell_6t
Xbit_r333_c122 bl[122] br[122] wl[333] vdd gnd cell_6t
Xbit_r334_c122 bl[122] br[122] wl[334] vdd gnd cell_6t
Xbit_r335_c122 bl[122] br[122] wl[335] vdd gnd cell_6t
Xbit_r336_c122 bl[122] br[122] wl[336] vdd gnd cell_6t
Xbit_r337_c122 bl[122] br[122] wl[337] vdd gnd cell_6t
Xbit_r338_c122 bl[122] br[122] wl[338] vdd gnd cell_6t
Xbit_r339_c122 bl[122] br[122] wl[339] vdd gnd cell_6t
Xbit_r340_c122 bl[122] br[122] wl[340] vdd gnd cell_6t
Xbit_r341_c122 bl[122] br[122] wl[341] vdd gnd cell_6t
Xbit_r342_c122 bl[122] br[122] wl[342] vdd gnd cell_6t
Xbit_r343_c122 bl[122] br[122] wl[343] vdd gnd cell_6t
Xbit_r344_c122 bl[122] br[122] wl[344] vdd gnd cell_6t
Xbit_r345_c122 bl[122] br[122] wl[345] vdd gnd cell_6t
Xbit_r346_c122 bl[122] br[122] wl[346] vdd gnd cell_6t
Xbit_r347_c122 bl[122] br[122] wl[347] vdd gnd cell_6t
Xbit_r348_c122 bl[122] br[122] wl[348] vdd gnd cell_6t
Xbit_r349_c122 bl[122] br[122] wl[349] vdd gnd cell_6t
Xbit_r350_c122 bl[122] br[122] wl[350] vdd gnd cell_6t
Xbit_r351_c122 bl[122] br[122] wl[351] vdd gnd cell_6t
Xbit_r352_c122 bl[122] br[122] wl[352] vdd gnd cell_6t
Xbit_r353_c122 bl[122] br[122] wl[353] vdd gnd cell_6t
Xbit_r354_c122 bl[122] br[122] wl[354] vdd gnd cell_6t
Xbit_r355_c122 bl[122] br[122] wl[355] vdd gnd cell_6t
Xbit_r356_c122 bl[122] br[122] wl[356] vdd gnd cell_6t
Xbit_r357_c122 bl[122] br[122] wl[357] vdd gnd cell_6t
Xbit_r358_c122 bl[122] br[122] wl[358] vdd gnd cell_6t
Xbit_r359_c122 bl[122] br[122] wl[359] vdd gnd cell_6t
Xbit_r360_c122 bl[122] br[122] wl[360] vdd gnd cell_6t
Xbit_r361_c122 bl[122] br[122] wl[361] vdd gnd cell_6t
Xbit_r362_c122 bl[122] br[122] wl[362] vdd gnd cell_6t
Xbit_r363_c122 bl[122] br[122] wl[363] vdd gnd cell_6t
Xbit_r364_c122 bl[122] br[122] wl[364] vdd gnd cell_6t
Xbit_r365_c122 bl[122] br[122] wl[365] vdd gnd cell_6t
Xbit_r366_c122 bl[122] br[122] wl[366] vdd gnd cell_6t
Xbit_r367_c122 bl[122] br[122] wl[367] vdd gnd cell_6t
Xbit_r368_c122 bl[122] br[122] wl[368] vdd gnd cell_6t
Xbit_r369_c122 bl[122] br[122] wl[369] vdd gnd cell_6t
Xbit_r370_c122 bl[122] br[122] wl[370] vdd gnd cell_6t
Xbit_r371_c122 bl[122] br[122] wl[371] vdd gnd cell_6t
Xbit_r372_c122 bl[122] br[122] wl[372] vdd gnd cell_6t
Xbit_r373_c122 bl[122] br[122] wl[373] vdd gnd cell_6t
Xbit_r374_c122 bl[122] br[122] wl[374] vdd gnd cell_6t
Xbit_r375_c122 bl[122] br[122] wl[375] vdd gnd cell_6t
Xbit_r376_c122 bl[122] br[122] wl[376] vdd gnd cell_6t
Xbit_r377_c122 bl[122] br[122] wl[377] vdd gnd cell_6t
Xbit_r378_c122 bl[122] br[122] wl[378] vdd gnd cell_6t
Xbit_r379_c122 bl[122] br[122] wl[379] vdd gnd cell_6t
Xbit_r380_c122 bl[122] br[122] wl[380] vdd gnd cell_6t
Xbit_r381_c122 bl[122] br[122] wl[381] vdd gnd cell_6t
Xbit_r382_c122 bl[122] br[122] wl[382] vdd gnd cell_6t
Xbit_r383_c122 bl[122] br[122] wl[383] vdd gnd cell_6t
Xbit_r384_c122 bl[122] br[122] wl[384] vdd gnd cell_6t
Xbit_r385_c122 bl[122] br[122] wl[385] vdd gnd cell_6t
Xbit_r386_c122 bl[122] br[122] wl[386] vdd gnd cell_6t
Xbit_r387_c122 bl[122] br[122] wl[387] vdd gnd cell_6t
Xbit_r388_c122 bl[122] br[122] wl[388] vdd gnd cell_6t
Xbit_r389_c122 bl[122] br[122] wl[389] vdd gnd cell_6t
Xbit_r390_c122 bl[122] br[122] wl[390] vdd gnd cell_6t
Xbit_r391_c122 bl[122] br[122] wl[391] vdd gnd cell_6t
Xbit_r392_c122 bl[122] br[122] wl[392] vdd gnd cell_6t
Xbit_r393_c122 bl[122] br[122] wl[393] vdd gnd cell_6t
Xbit_r394_c122 bl[122] br[122] wl[394] vdd gnd cell_6t
Xbit_r395_c122 bl[122] br[122] wl[395] vdd gnd cell_6t
Xbit_r396_c122 bl[122] br[122] wl[396] vdd gnd cell_6t
Xbit_r397_c122 bl[122] br[122] wl[397] vdd gnd cell_6t
Xbit_r398_c122 bl[122] br[122] wl[398] vdd gnd cell_6t
Xbit_r399_c122 bl[122] br[122] wl[399] vdd gnd cell_6t
Xbit_r400_c122 bl[122] br[122] wl[400] vdd gnd cell_6t
Xbit_r401_c122 bl[122] br[122] wl[401] vdd gnd cell_6t
Xbit_r402_c122 bl[122] br[122] wl[402] vdd gnd cell_6t
Xbit_r403_c122 bl[122] br[122] wl[403] vdd gnd cell_6t
Xbit_r404_c122 bl[122] br[122] wl[404] vdd gnd cell_6t
Xbit_r405_c122 bl[122] br[122] wl[405] vdd gnd cell_6t
Xbit_r406_c122 bl[122] br[122] wl[406] vdd gnd cell_6t
Xbit_r407_c122 bl[122] br[122] wl[407] vdd gnd cell_6t
Xbit_r408_c122 bl[122] br[122] wl[408] vdd gnd cell_6t
Xbit_r409_c122 bl[122] br[122] wl[409] vdd gnd cell_6t
Xbit_r410_c122 bl[122] br[122] wl[410] vdd gnd cell_6t
Xbit_r411_c122 bl[122] br[122] wl[411] vdd gnd cell_6t
Xbit_r412_c122 bl[122] br[122] wl[412] vdd gnd cell_6t
Xbit_r413_c122 bl[122] br[122] wl[413] vdd gnd cell_6t
Xbit_r414_c122 bl[122] br[122] wl[414] vdd gnd cell_6t
Xbit_r415_c122 bl[122] br[122] wl[415] vdd gnd cell_6t
Xbit_r416_c122 bl[122] br[122] wl[416] vdd gnd cell_6t
Xbit_r417_c122 bl[122] br[122] wl[417] vdd gnd cell_6t
Xbit_r418_c122 bl[122] br[122] wl[418] vdd gnd cell_6t
Xbit_r419_c122 bl[122] br[122] wl[419] vdd gnd cell_6t
Xbit_r420_c122 bl[122] br[122] wl[420] vdd gnd cell_6t
Xbit_r421_c122 bl[122] br[122] wl[421] vdd gnd cell_6t
Xbit_r422_c122 bl[122] br[122] wl[422] vdd gnd cell_6t
Xbit_r423_c122 bl[122] br[122] wl[423] vdd gnd cell_6t
Xbit_r424_c122 bl[122] br[122] wl[424] vdd gnd cell_6t
Xbit_r425_c122 bl[122] br[122] wl[425] vdd gnd cell_6t
Xbit_r426_c122 bl[122] br[122] wl[426] vdd gnd cell_6t
Xbit_r427_c122 bl[122] br[122] wl[427] vdd gnd cell_6t
Xbit_r428_c122 bl[122] br[122] wl[428] vdd gnd cell_6t
Xbit_r429_c122 bl[122] br[122] wl[429] vdd gnd cell_6t
Xbit_r430_c122 bl[122] br[122] wl[430] vdd gnd cell_6t
Xbit_r431_c122 bl[122] br[122] wl[431] vdd gnd cell_6t
Xbit_r432_c122 bl[122] br[122] wl[432] vdd gnd cell_6t
Xbit_r433_c122 bl[122] br[122] wl[433] vdd gnd cell_6t
Xbit_r434_c122 bl[122] br[122] wl[434] vdd gnd cell_6t
Xbit_r435_c122 bl[122] br[122] wl[435] vdd gnd cell_6t
Xbit_r436_c122 bl[122] br[122] wl[436] vdd gnd cell_6t
Xbit_r437_c122 bl[122] br[122] wl[437] vdd gnd cell_6t
Xbit_r438_c122 bl[122] br[122] wl[438] vdd gnd cell_6t
Xbit_r439_c122 bl[122] br[122] wl[439] vdd gnd cell_6t
Xbit_r440_c122 bl[122] br[122] wl[440] vdd gnd cell_6t
Xbit_r441_c122 bl[122] br[122] wl[441] vdd gnd cell_6t
Xbit_r442_c122 bl[122] br[122] wl[442] vdd gnd cell_6t
Xbit_r443_c122 bl[122] br[122] wl[443] vdd gnd cell_6t
Xbit_r444_c122 bl[122] br[122] wl[444] vdd gnd cell_6t
Xbit_r445_c122 bl[122] br[122] wl[445] vdd gnd cell_6t
Xbit_r446_c122 bl[122] br[122] wl[446] vdd gnd cell_6t
Xbit_r447_c122 bl[122] br[122] wl[447] vdd gnd cell_6t
Xbit_r448_c122 bl[122] br[122] wl[448] vdd gnd cell_6t
Xbit_r449_c122 bl[122] br[122] wl[449] vdd gnd cell_6t
Xbit_r450_c122 bl[122] br[122] wl[450] vdd gnd cell_6t
Xbit_r451_c122 bl[122] br[122] wl[451] vdd gnd cell_6t
Xbit_r452_c122 bl[122] br[122] wl[452] vdd gnd cell_6t
Xbit_r453_c122 bl[122] br[122] wl[453] vdd gnd cell_6t
Xbit_r454_c122 bl[122] br[122] wl[454] vdd gnd cell_6t
Xbit_r455_c122 bl[122] br[122] wl[455] vdd gnd cell_6t
Xbit_r456_c122 bl[122] br[122] wl[456] vdd gnd cell_6t
Xbit_r457_c122 bl[122] br[122] wl[457] vdd gnd cell_6t
Xbit_r458_c122 bl[122] br[122] wl[458] vdd gnd cell_6t
Xbit_r459_c122 bl[122] br[122] wl[459] vdd gnd cell_6t
Xbit_r460_c122 bl[122] br[122] wl[460] vdd gnd cell_6t
Xbit_r461_c122 bl[122] br[122] wl[461] vdd gnd cell_6t
Xbit_r462_c122 bl[122] br[122] wl[462] vdd gnd cell_6t
Xbit_r463_c122 bl[122] br[122] wl[463] vdd gnd cell_6t
Xbit_r464_c122 bl[122] br[122] wl[464] vdd gnd cell_6t
Xbit_r465_c122 bl[122] br[122] wl[465] vdd gnd cell_6t
Xbit_r466_c122 bl[122] br[122] wl[466] vdd gnd cell_6t
Xbit_r467_c122 bl[122] br[122] wl[467] vdd gnd cell_6t
Xbit_r468_c122 bl[122] br[122] wl[468] vdd gnd cell_6t
Xbit_r469_c122 bl[122] br[122] wl[469] vdd gnd cell_6t
Xbit_r470_c122 bl[122] br[122] wl[470] vdd gnd cell_6t
Xbit_r471_c122 bl[122] br[122] wl[471] vdd gnd cell_6t
Xbit_r472_c122 bl[122] br[122] wl[472] vdd gnd cell_6t
Xbit_r473_c122 bl[122] br[122] wl[473] vdd gnd cell_6t
Xbit_r474_c122 bl[122] br[122] wl[474] vdd gnd cell_6t
Xbit_r475_c122 bl[122] br[122] wl[475] vdd gnd cell_6t
Xbit_r476_c122 bl[122] br[122] wl[476] vdd gnd cell_6t
Xbit_r477_c122 bl[122] br[122] wl[477] vdd gnd cell_6t
Xbit_r478_c122 bl[122] br[122] wl[478] vdd gnd cell_6t
Xbit_r479_c122 bl[122] br[122] wl[479] vdd gnd cell_6t
Xbit_r480_c122 bl[122] br[122] wl[480] vdd gnd cell_6t
Xbit_r481_c122 bl[122] br[122] wl[481] vdd gnd cell_6t
Xbit_r482_c122 bl[122] br[122] wl[482] vdd gnd cell_6t
Xbit_r483_c122 bl[122] br[122] wl[483] vdd gnd cell_6t
Xbit_r484_c122 bl[122] br[122] wl[484] vdd gnd cell_6t
Xbit_r485_c122 bl[122] br[122] wl[485] vdd gnd cell_6t
Xbit_r486_c122 bl[122] br[122] wl[486] vdd gnd cell_6t
Xbit_r487_c122 bl[122] br[122] wl[487] vdd gnd cell_6t
Xbit_r488_c122 bl[122] br[122] wl[488] vdd gnd cell_6t
Xbit_r489_c122 bl[122] br[122] wl[489] vdd gnd cell_6t
Xbit_r490_c122 bl[122] br[122] wl[490] vdd gnd cell_6t
Xbit_r491_c122 bl[122] br[122] wl[491] vdd gnd cell_6t
Xbit_r492_c122 bl[122] br[122] wl[492] vdd gnd cell_6t
Xbit_r493_c122 bl[122] br[122] wl[493] vdd gnd cell_6t
Xbit_r494_c122 bl[122] br[122] wl[494] vdd gnd cell_6t
Xbit_r495_c122 bl[122] br[122] wl[495] vdd gnd cell_6t
Xbit_r496_c122 bl[122] br[122] wl[496] vdd gnd cell_6t
Xbit_r497_c122 bl[122] br[122] wl[497] vdd gnd cell_6t
Xbit_r498_c122 bl[122] br[122] wl[498] vdd gnd cell_6t
Xbit_r499_c122 bl[122] br[122] wl[499] vdd gnd cell_6t
Xbit_r500_c122 bl[122] br[122] wl[500] vdd gnd cell_6t
Xbit_r501_c122 bl[122] br[122] wl[501] vdd gnd cell_6t
Xbit_r502_c122 bl[122] br[122] wl[502] vdd gnd cell_6t
Xbit_r503_c122 bl[122] br[122] wl[503] vdd gnd cell_6t
Xbit_r504_c122 bl[122] br[122] wl[504] vdd gnd cell_6t
Xbit_r505_c122 bl[122] br[122] wl[505] vdd gnd cell_6t
Xbit_r506_c122 bl[122] br[122] wl[506] vdd gnd cell_6t
Xbit_r507_c122 bl[122] br[122] wl[507] vdd gnd cell_6t
Xbit_r508_c122 bl[122] br[122] wl[508] vdd gnd cell_6t
Xbit_r509_c122 bl[122] br[122] wl[509] vdd gnd cell_6t
Xbit_r510_c122 bl[122] br[122] wl[510] vdd gnd cell_6t
Xbit_r511_c122 bl[122] br[122] wl[511] vdd gnd cell_6t
Xbit_r0_c123 bl[123] br[123] wl[0] vdd gnd cell_6t
Xbit_r1_c123 bl[123] br[123] wl[1] vdd gnd cell_6t
Xbit_r2_c123 bl[123] br[123] wl[2] vdd gnd cell_6t
Xbit_r3_c123 bl[123] br[123] wl[3] vdd gnd cell_6t
Xbit_r4_c123 bl[123] br[123] wl[4] vdd gnd cell_6t
Xbit_r5_c123 bl[123] br[123] wl[5] vdd gnd cell_6t
Xbit_r6_c123 bl[123] br[123] wl[6] vdd gnd cell_6t
Xbit_r7_c123 bl[123] br[123] wl[7] vdd gnd cell_6t
Xbit_r8_c123 bl[123] br[123] wl[8] vdd gnd cell_6t
Xbit_r9_c123 bl[123] br[123] wl[9] vdd gnd cell_6t
Xbit_r10_c123 bl[123] br[123] wl[10] vdd gnd cell_6t
Xbit_r11_c123 bl[123] br[123] wl[11] vdd gnd cell_6t
Xbit_r12_c123 bl[123] br[123] wl[12] vdd gnd cell_6t
Xbit_r13_c123 bl[123] br[123] wl[13] vdd gnd cell_6t
Xbit_r14_c123 bl[123] br[123] wl[14] vdd gnd cell_6t
Xbit_r15_c123 bl[123] br[123] wl[15] vdd gnd cell_6t
Xbit_r16_c123 bl[123] br[123] wl[16] vdd gnd cell_6t
Xbit_r17_c123 bl[123] br[123] wl[17] vdd gnd cell_6t
Xbit_r18_c123 bl[123] br[123] wl[18] vdd gnd cell_6t
Xbit_r19_c123 bl[123] br[123] wl[19] vdd gnd cell_6t
Xbit_r20_c123 bl[123] br[123] wl[20] vdd gnd cell_6t
Xbit_r21_c123 bl[123] br[123] wl[21] vdd gnd cell_6t
Xbit_r22_c123 bl[123] br[123] wl[22] vdd gnd cell_6t
Xbit_r23_c123 bl[123] br[123] wl[23] vdd gnd cell_6t
Xbit_r24_c123 bl[123] br[123] wl[24] vdd gnd cell_6t
Xbit_r25_c123 bl[123] br[123] wl[25] vdd gnd cell_6t
Xbit_r26_c123 bl[123] br[123] wl[26] vdd gnd cell_6t
Xbit_r27_c123 bl[123] br[123] wl[27] vdd gnd cell_6t
Xbit_r28_c123 bl[123] br[123] wl[28] vdd gnd cell_6t
Xbit_r29_c123 bl[123] br[123] wl[29] vdd gnd cell_6t
Xbit_r30_c123 bl[123] br[123] wl[30] vdd gnd cell_6t
Xbit_r31_c123 bl[123] br[123] wl[31] vdd gnd cell_6t
Xbit_r32_c123 bl[123] br[123] wl[32] vdd gnd cell_6t
Xbit_r33_c123 bl[123] br[123] wl[33] vdd gnd cell_6t
Xbit_r34_c123 bl[123] br[123] wl[34] vdd gnd cell_6t
Xbit_r35_c123 bl[123] br[123] wl[35] vdd gnd cell_6t
Xbit_r36_c123 bl[123] br[123] wl[36] vdd gnd cell_6t
Xbit_r37_c123 bl[123] br[123] wl[37] vdd gnd cell_6t
Xbit_r38_c123 bl[123] br[123] wl[38] vdd gnd cell_6t
Xbit_r39_c123 bl[123] br[123] wl[39] vdd gnd cell_6t
Xbit_r40_c123 bl[123] br[123] wl[40] vdd gnd cell_6t
Xbit_r41_c123 bl[123] br[123] wl[41] vdd gnd cell_6t
Xbit_r42_c123 bl[123] br[123] wl[42] vdd gnd cell_6t
Xbit_r43_c123 bl[123] br[123] wl[43] vdd gnd cell_6t
Xbit_r44_c123 bl[123] br[123] wl[44] vdd gnd cell_6t
Xbit_r45_c123 bl[123] br[123] wl[45] vdd gnd cell_6t
Xbit_r46_c123 bl[123] br[123] wl[46] vdd gnd cell_6t
Xbit_r47_c123 bl[123] br[123] wl[47] vdd gnd cell_6t
Xbit_r48_c123 bl[123] br[123] wl[48] vdd gnd cell_6t
Xbit_r49_c123 bl[123] br[123] wl[49] vdd gnd cell_6t
Xbit_r50_c123 bl[123] br[123] wl[50] vdd gnd cell_6t
Xbit_r51_c123 bl[123] br[123] wl[51] vdd gnd cell_6t
Xbit_r52_c123 bl[123] br[123] wl[52] vdd gnd cell_6t
Xbit_r53_c123 bl[123] br[123] wl[53] vdd gnd cell_6t
Xbit_r54_c123 bl[123] br[123] wl[54] vdd gnd cell_6t
Xbit_r55_c123 bl[123] br[123] wl[55] vdd gnd cell_6t
Xbit_r56_c123 bl[123] br[123] wl[56] vdd gnd cell_6t
Xbit_r57_c123 bl[123] br[123] wl[57] vdd gnd cell_6t
Xbit_r58_c123 bl[123] br[123] wl[58] vdd gnd cell_6t
Xbit_r59_c123 bl[123] br[123] wl[59] vdd gnd cell_6t
Xbit_r60_c123 bl[123] br[123] wl[60] vdd gnd cell_6t
Xbit_r61_c123 bl[123] br[123] wl[61] vdd gnd cell_6t
Xbit_r62_c123 bl[123] br[123] wl[62] vdd gnd cell_6t
Xbit_r63_c123 bl[123] br[123] wl[63] vdd gnd cell_6t
Xbit_r64_c123 bl[123] br[123] wl[64] vdd gnd cell_6t
Xbit_r65_c123 bl[123] br[123] wl[65] vdd gnd cell_6t
Xbit_r66_c123 bl[123] br[123] wl[66] vdd gnd cell_6t
Xbit_r67_c123 bl[123] br[123] wl[67] vdd gnd cell_6t
Xbit_r68_c123 bl[123] br[123] wl[68] vdd gnd cell_6t
Xbit_r69_c123 bl[123] br[123] wl[69] vdd gnd cell_6t
Xbit_r70_c123 bl[123] br[123] wl[70] vdd gnd cell_6t
Xbit_r71_c123 bl[123] br[123] wl[71] vdd gnd cell_6t
Xbit_r72_c123 bl[123] br[123] wl[72] vdd gnd cell_6t
Xbit_r73_c123 bl[123] br[123] wl[73] vdd gnd cell_6t
Xbit_r74_c123 bl[123] br[123] wl[74] vdd gnd cell_6t
Xbit_r75_c123 bl[123] br[123] wl[75] vdd gnd cell_6t
Xbit_r76_c123 bl[123] br[123] wl[76] vdd gnd cell_6t
Xbit_r77_c123 bl[123] br[123] wl[77] vdd gnd cell_6t
Xbit_r78_c123 bl[123] br[123] wl[78] vdd gnd cell_6t
Xbit_r79_c123 bl[123] br[123] wl[79] vdd gnd cell_6t
Xbit_r80_c123 bl[123] br[123] wl[80] vdd gnd cell_6t
Xbit_r81_c123 bl[123] br[123] wl[81] vdd gnd cell_6t
Xbit_r82_c123 bl[123] br[123] wl[82] vdd gnd cell_6t
Xbit_r83_c123 bl[123] br[123] wl[83] vdd gnd cell_6t
Xbit_r84_c123 bl[123] br[123] wl[84] vdd gnd cell_6t
Xbit_r85_c123 bl[123] br[123] wl[85] vdd gnd cell_6t
Xbit_r86_c123 bl[123] br[123] wl[86] vdd gnd cell_6t
Xbit_r87_c123 bl[123] br[123] wl[87] vdd gnd cell_6t
Xbit_r88_c123 bl[123] br[123] wl[88] vdd gnd cell_6t
Xbit_r89_c123 bl[123] br[123] wl[89] vdd gnd cell_6t
Xbit_r90_c123 bl[123] br[123] wl[90] vdd gnd cell_6t
Xbit_r91_c123 bl[123] br[123] wl[91] vdd gnd cell_6t
Xbit_r92_c123 bl[123] br[123] wl[92] vdd gnd cell_6t
Xbit_r93_c123 bl[123] br[123] wl[93] vdd gnd cell_6t
Xbit_r94_c123 bl[123] br[123] wl[94] vdd gnd cell_6t
Xbit_r95_c123 bl[123] br[123] wl[95] vdd gnd cell_6t
Xbit_r96_c123 bl[123] br[123] wl[96] vdd gnd cell_6t
Xbit_r97_c123 bl[123] br[123] wl[97] vdd gnd cell_6t
Xbit_r98_c123 bl[123] br[123] wl[98] vdd gnd cell_6t
Xbit_r99_c123 bl[123] br[123] wl[99] vdd gnd cell_6t
Xbit_r100_c123 bl[123] br[123] wl[100] vdd gnd cell_6t
Xbit_r101_c123 bl[123] br[123] wl[101] vdd gnd cell_6t
Xbit_r102_c123 bl[123] br[123] wl[102] vdd gnd cell_6t
Xbit_r103_c123 bl[123] br[123] wl[103] vdd gnd cell_6t
Xbit_r104_c123 bl[123] br[123] wl[104] vdd gnd cell_6t
Xbit_r105_c123 bl[123] br[123] wl[105] vdd gnd cell_6t
Xbit_r106_c123 bl[123] br[123] wl[106] vdd gnd cell_6t
Xbit_r107_c123 bl[123] br[123] wl[107] vdd gnd cell_6t
Xbit_r108_c123 bl[123] br[123] wl[108] vdd gnd cell_6t
Xbit_r109_c123 bl[123] br[123] wl[109] vdd gnd cell_6t
Xbit_r110_c123 bl[123] br[123] wl[110] vdd gnd cell_6t
Xbit_r111_c123 bl[123] br[123] wl[111] vdd gnd cell_6t
Xbit_r112_c123 bl[123] br[123] wl[112] vdd gnd cell_6t
Xbit_r113_c123 bl[123] br[123] wl[113] vdd gnd cell_6t
Xbit_r114_c123 bl[123] br[123] wl[114] vdd gnd cell_6t
Xbit_r115_c123 bl[123] br[123] wl[115] vdd gnd cell_6t
Xbit_r116_c123 bl[123] br[123] wl[116] vdd gnd cell_6t
Xbit_r117_c123 bl[123] br[123] wl[117] vdd gnd cell_6t
Xbit_r118_c123 bl[123] br[123] wl[118] vdd gnd cell_6t
Xbit_r119_c123 bl[123] br[123] wl[119] vdd gnd cell_6t
Xbit_r120_c123 bl[123] br[123] wl[120] vdd gnd cell_6t
Xbit_r121_c123 bl[123] br[123] wl[121] vdd gnd cell_6t
Xbit_r122_c123 bl[123] br[123] wl[122] vdd gnd cell_6t
Xbit_r123_c123 bl[123] br[123] wl[123] vdd gnd cell_6t
Xbit_r124_c123 bl[123] br[123] wl[124] vdd gnd cell_6t
Xbit_r125_c123 bl[123] br[123] wl[125] vdd gnd cell_6t
Xbit_r126_c123 bl[123] br[123] wl[126] vdd gnd cell_6t
Xbit_r127_c123 bl[123] br[123] wl[127] vdd gnd cell_6t
Xbit_r128_c123 bl[123] br[123] wl[128] vdd gnd cell_6t
Xbit_r129_c123 bl[123] br[123] wl[129] vdd gnd cell_6t
Xbit_r130_c123 bl[123] br[123] wl[130] vdd gnd cell_6t
Xbit_r131_c123 bl[123] br[123] wl[131] vdd gnd cell_6t
Xbit_r132_c123 bl[123] br[123] wl[132] vdd gnd cell_6t
Xbit_r133_c123 bl[123] br[123] wl[133] vdd gnd cell_6t
Xbit_r134_c123 bl[123] br[123] wl[134] vdd gnd cell_6t
Xbit_r135_c123 bl[123] br[123] wl[135] vdd gnd cell_6t
Xbit_r136_c123 bl[123] br[123] wl[136] vdd gnd cell_6t
Xbit_r137_c123 bl[123] br[123] wl[137] vdd gnd cell_6t
Xbit_r138_c123 bl[123] br[123] wl[138] vdd gnd cell_6t
Xbit_r139_c123 bl[123] br[123] wl[139] vdd gnd cell_6t
Xbit_r140_c123 bl[123] br[123] wl[140] vdd gnd cell_6t
Xbit_r141_c123 bl[123] br[123] wl[141] vdd gnd cell_6t
Xbit_r142_c123 bl[123] br[123] wl[142] vdd gnd cell_6t
Xbit_r143_c123 bl[123] br[123] wl[143] vdd gnd cell_6t
Xbit_r144_c123 bl[123] br[123] wl[144] vdd gnd cell_6t
Xbit_r145_c123 bl[123] br[123] wl[145] vdd gnd cell_6t
Xbit_r146_c123 bl[123] br[123] wl[146] vdd gnd cell_6t
Xbit_r147_c123 bl[123] br[123] wl[147] vdd gnd cell_6t
Xbit_r148_c123 bl[123] br[123] wl[148] vdd gnd cell_6t
Xbit_r149_c123 bl[123] br[123] wl[149] vdd gnd cell_6t
Xbit_r150_c123 bl[123] br[123] wl[150] vdd gnd cell_6t
Xbit_r151_c123 bl[123] br[123] wl[151] vdd gnd cell_6t
Xbit_r152_c123 bl[123] br[123] wl[152] vdd gnd cell_6t
Xbit_r153_c123 bl[123] br[123] wl[153] vdd gnd cell_6t
Xbit_r154_c123 bl[123] br[123] wl[154] vdd gnd cell_6t
Xbit_r155_c123 bl[123] br[123] wl[155] vdd gnd cell_6t
Xbit_r156_c123 bl[123] br[123] wl[156] vdd gnd cell_6t
Xbit_r157_c123 bl[123] br[123] wl[157] vdd gnd cell_6t
Xbit_r158_c123 bl[123] br[123] wl[158] vdd gnd cell_6t
Xbit_r159_c123 bl[123] br[123] wl[159] vdd gnd cell_6t
Xbit_r160_c123 bl[123] br[123] wl[160] vdd gnd cell_6t
Xbit_r161_c123 bl[123] br[123] wl[161] vdd gnd cell_6t
Xbit_r162_c123 bl[123] br[123] wl[162] vdd gnd cell_6t
Xbit_r163_c123 bl[123] br[123] wl[163] vdd gnd cell_6t
Xbit_r164_c123 bl[123] br[123] wl[164] vdd gnd cell_6t
Xbit_r165_c123 bl[123] br[123] wl[165] vdd gnd cell_6t
Xbit_r166_c123 bl[123] br[123] wl[166] vdd gnd cell_6t
Xbit_r167_c123 bl[123] br[123] wl[167] vdd gnd cell_6t
Xbit_r168_c123 bl[123] br[123] wl[168] vdd gnd cell_6t
Xbit_r169_c123 bl[123] br[123] wl[169] vdd gnd cell_6t
Xbit_r170_c123 bl[123] br[123] wl[170] vdd gnd cell_6t
Xbit_r171_c123 bl[123] br[123] wl[171] vdd gnd cell_6t
Xbit_r172_c123 bl[123] br[123] wl[172] vdd gnd cell_6t
Xbit_r173_c123 bl[123] br[123] wl[173] vdd gnd cell_6t
Xbit_r174_c123 bl[123] br[123] wl[174] vdd gnd cell_6t
Xbit_r175_c123 bl[123] br[123] wl[175] vdd gnd cell_6t
Xbit_r176_c123 bl[123] br[123] wl[176] vdd gnd cell_6t
Xbit_r177_c123 bl[123] br[123] wl[177] vdd gnd cell_6t
Xbit_r178_c123 bl[123] br[123] wl[178] vdd gnd cell_6t
Xbit_r179_c123 bl[123] br[123] wl[179] vdd gnd cell_6t
Xbit_r180_c123 bl[123] br[123] wl[180] vdd gnd cell_6t
Xbit_r181_c123 bl[123] br[123] wl[181] vdd gnd cell_6t
Xbit_r182_c123 bl[123] br[123] wl[182] vdd gnd cell_6t
Xbit_r183_c123 bl[123] br[123] wl[183] vdd gnd cell_6t
Xbit_r184_c123 bl[123] br[123] wl[184] vdd gnd cell_6t
Xbit_r185_c123 bl[123] br[123] wl[185] vdd gnd cell_6t
Xbit_r186_c123 bl[123] br[123] wl[186] vdd gnd cell_6t
Xbit_r187_c123 bl[123] br[123] wl[187] vdd gnd cell_6t
Xbit_r188_c123 bl[123] br[123] wl[188] vdd gnd cell_6t
Xbit_r189_c123 bl[123] br[123] wl[189] vdd gnd cell_6t
Xbit_r190_c123 bl[123] br[123] wl[190] vdd gnd cell_6t
Xbit_r191_c123 bl[123] br[123] wl[191] vdd gnd cell_6t
Xbit_r192_c123 bl[123] br[123] wl[192] vdd gnd cell_6t
Xbit_r193_c123 bl[123] br[123] wl[193] vdd gnd cell_6t
Xbit_r194_c123 bl[123] br[123] wl[194] vdd gnd cell_6t
Xbit_r195_c123 bl[123] br[123] wl[195] vdd gnd cell_6t
Xbit_r196_c123 bl[123] br[123] wl[196] vdd gnd cell_6t
Xbit_r197_c123 bl[123] br[123] wl[197] vdd gnd cell_6t
Xbit_r198_c123 bl[123] br[123] wl[198] vdd gnd cell_6t
Xbit_r199_c123 bl[123] br[123] wl[199] vdd gnd cell_6t
Xbit_r200_c123 bl[123] br[123] wl[200] vdd gnd cell_6t
Xbit_r201_c123 bl[123] br[123] wl[201] vdd gnd cell_6t
Xbit_r202_c123 bl[123] br[123] wl[202] vdd gnd cell_6t
Xbit_r203_c123 bl[123] br[123] wl[203] vdd gnd cell_6t
Xbit_r204_c123 bl[123] br[123] wl[204] vdd gnd cell_6t
Xbit_r205_c123 bl[123] br[123] wl[205] vdd gnd cell_6t
Xbit_r206_c123 bl[123] br[123] wl[206] vdd gnd cell_6t
Xbit_r207_c123 bl[123] br[123] wl[207] vdd gnd cell_6t
Xbit_r208_c123 bl[123] br[123] wl[208] vdd gnd cell_6t
Xbit_r209_c123 bl[123] br[123] wl[209] vdd gnd cell_6t
Xbit_r210_c123 bl[123] br[123] wl[210] vdd gnd cell_6t
Xbit_r211_c123 bl[123] br[123] wl[211] vdd gnd cell_6t
Xbit_r212_c123 bl[123] br[123] wl[212] vdd gnd cell_6t
Xbit_r213_c123 bl[123] br[123] wl[213] vdd gnd cell_6t
Xbit_r214_c123 bl[123] br[123] wl[214] vdd gnd cell_6t
Xbit_r215_c123 bl[123] br[123] wl[215] vdd gnd cell_6t
Xbit_r216_c123 bl[123] br[123] wl[216] vdd gnd cell_6t
Xbit_r217_c123 bl[123] br[123] wl[217] vdd gnd cell_6t
Xbit_r218_c123 bl[123] br[123] wl[218] vdd gnd cell_6t
Xbit_r219_c123 bl[123] br[123] wl[219] vdd gnd cell_6t
Xbit_r220_c123 bl[123] br[123] wl[220] vdd gnd cell_6t
Xbit_r221_c123 bl[123] br[123] wl[221] vdd gnd cell_6t
Xbit_r222_c123 bl[123] br[123] wl[222] vdd gnd cell_6t
Xbit_r223_c123 bl[123] br[123] wl[223] vdd gnd cell_6t
Xbit_r224_c123 bl[123] br[123] wl[224] vdd gnd cell_6t
Xbit_r225_c123 bl[123] br[123] wl[225] vdd gnd cell_6t
Xbit_r226_c123 bl[123] br[123] wl[226] vdd gnd cell_6t
Xbit_r227_c123 bl[123] br[123] wl[227] vdd gnd cell_6t
Xbit_r228_c123 bl[123] br[123] wl[228] vdd gnd cell_6t
Xbit_r229_c123 bl[123] br[123] wl[229] vdd gnd cell_6t
Xbit_r230_c123 bl[123] br[123] wl[230] vdd gnd cell_6t
Xbit_r231_c123 bl[123] br[123] wl[231] vdd gnd cell_6t
Xbit_r232_c123 bl[123] br[123] wl[232] vdd gnd cell_6t
Xbit_r233_c123 bl[123] br[123] wl[233] vdd gnd cell_6t
Xbit_r234_c123 bl[123] br[123] wl[234] vdd gnd cell_6t
Xbit_r235_c123 bl[123] br[123] wl[235] vdd gnd cell_6t
Xbit_r236_c123 bl[123] br[123] wl[236] vdd gnd cell_6t
Xbit_r237_c123 bl[123] br[123] wl[237] vdd gnd cell_6t
Xbit_r238_c123 bl[123] br[123] wl[238] vdd gnd cell_6t
Xbit_r239_c123 bl[123] br[123] wl[239] vdd gnd cell_6t
Xbit_r240_c123 bl[123] br[123] wl[240] vdd gnd cell_6t
Xbit_r241_c123 bl[123] br[123] wl[241] vdd gnd cell_6t
Xbit_r242_c123 bl[123] br[123] wl[242] vdd gnd cell_6t
Xbit_r243_c123 bl[123] br[123] wl[243] vdd gnd cell_6t
Xbit_r244_c123 bl[123] br[123] wl[244] vdd gnd cell_6t
Xbit_r245_c123 bl[123] br[123] wl[245] vdd gnd cell_6t
Xbit_r246_c123 bl[123] br[123] wl[246] vdd gnd cell_6t
Xbit_r247_c123 bl[123] br[123] wl[247] vdd gnd cell_6t
Xbit_r248_c123 bl[123] br[123] wl[248] vdd gnd cell_6t
Xbit_r249_c123 bl[123] br[123] wl[249] vdd gnd cell_6t
Xbit_r250_c123 bl[123] br[123] wl[250] vdd gnd cell_6t
Xbit_r251_c123 bl[123] br[123] wl[251] vdd gnd cell_6t
Xbit_r252_c123 bl[123] br[123] wl[252] vdd gnd cell_6t
Xbit_r253_c123 bl[123] br[123] wl[253] vdd gnd cell_6t
Xbit_r254_c123 bl[123] br[123] wl[254] vdd gnd cell_6t
Xbit_r255_c123 bl[123] br[123] wl[255] vdd gnd cell_6t
Xbit_r256_c123 bl[123] br[123] wl[256] vdd gnd cell_6t
Xbit_r257_c123 bl[123] br[123] wl[257] vdd gnd cell_6t
Xbit_r258_c123 bl[123] br[123] wl[258] vdd gnd cell_6t
Xbit_r259_c123 bl[123] br[123] wl[259] vdd gnd cell_6t
Xbit_r260_c123 bl[123] br[123] wl[260] vdd gnd cell_6t
Xbit_r261_c123 bl[123] br[123] wl[261] vdd gnd cell_6t
Xbit_r262_c123 bl[123] br[123] wl[262] vdd gnd cell_6t
Xbit_r263_c123 bl[123] br[123] wl[263] vdd gnd cell_6t
Xbit_r264_c123 bl[123] br[123] wl[264] vdd gnd cell_6t
Xbit_r265_c123 bl[123] br[123] wl[265] vdd gnd cell_6t
Xbit_r266_c123 bl[123] br[123] wl[266] vdd gnd cell_6t
Xbit_r267_c123 bl[123] br[123] wl[267] vdd gnd cell_6t
Xbit_r268_c123 bl[123] br[123] wl[268] vdd gnd cell_6t
Xbit_r269_c123 bl[123] br[123] wl[269] vdd gnd cell_6t
Xbit_r270_c123 bl[123] br[123] wl[270] vdd gnd cell_6t
Xbit_r271_c123 bl[123] br[123] wl[271] vdd gnd cell_6t
Xbit_r272_c123 bl[123] br[123] wl[272] vdd gnd cell_6t
Xbit_r273_c123 bl[123] br[123] wl[273] vdd gnd cell_6t
Xbit_r274_c123 bl[123] br[123] wl[274] vdd gnd cell_6t
Xbit_r275_c123 bl[123] br[123] wl[275] vdd gnd cell_6t
Xbit_r276_c123 bl[123] br[123] wl[276] vdd gnd cell_6t
Xbit_r277_c123 bl[123] br[123] wl[277] vdd gnd cell_6t
Xbit_r278_c123 bl[123] br[123] wl[278] vdd gnd cell_6t
Xbit_r279_c123 bl[123] br[123] wl[279] vdd gnd cell_6t
Xbit_r280_c123 bl[123] br[123] wl[280] vdd gnd cell_6t
Xbit_r281_c123 bl[123] br[123] wl[281] vdd gnd cell_6t
Xbit_r282_c123 bl[123] br[123] wl[282] vdd gnd cell_6t
Xbit_r283_c123 bl[123] br[123] wl[283] vdd gnd cell_6t
Xbit_r284_c123 bl[123] br[123] wl[284] vdd gnd cell_6t
Xbit_r285_c123 bl[123] br[123] wl[285] vdd gnd cell_6t
Xbit_r286_c123 bl[123] br[123] wl[286] vdd gnd cell_6t
Xbit_r287_c123 bl[123] br[123] wl[287] vdd gnd cell_6t
Xbit_r288_c123 bl[123] br[123] wl[288] vdd gnd cell_6t
Xbit_r289_c123 bl[123] br[123] wl[289] vdd gnd cell_6t
Xbit_r290_c123 bl[123] br[123] wl[290] vdd gnd cell_6t
Xbit_r291_c123 bl[123] br[123] wl[291] vdd gnd cell_6t
Xbit_r292_c123 bl[123] br[123] wl[292] vdd gnd cell_6t
Xbit_r293_c123 bl[123] br[123] wl[293] vdd gnd cell_6t
Xbit_r294_c123 bl[123] br[123] wl[294] vdd gnd cell_6t
Xbit_r295_c123 bl[123] br[123] wl[295] vdd gnd cell_6t
Xbit_r296_c123 bl[123] br[123] wl[296] vdd gnd cell_6t
Xbit_r297_c123 bl[123] br[123] wl[297] vdd gnd cell_6t
Xbit_r298_c123 bl[123] br[123] wl[298] vdd gnd cell_6t
Xbit_r299_c123 bl[123] br[123] wl[299] vdd gnd cell_6t
Xbit_r300_c123 bl[123] br[123] wl[300] vdd gnd cell_6t
Xbit_r301_c123 bl[123] br[123] wl[301] vdd gnd cell_6t
Xbit_r302_c123 bl[123] br[123] wl[302] vdd gnd cell_6t
Xbit_r303_c123 bl[123] br[123] wl[303] vdd gnd cell_6t
Xbit_r304_c123 bl[123] br[123] wl[304] vdd gnd cell_6t
Xbit_r305_c123 bl[123] br[123] wl[305] vdd gnd cell_6t
Xbit_r306_c123 bl[123] br[123] wl[306] vdd gnd cell_6t
Xbit_r307_c123 bl[123] br[123] wl[307] vdd gnd cell_6t
Xbit_r308_c123 bl[123] br[123] wl[308] vdd gnd cell_6t
Xbit_r309_c123 bl[123] br[123] wl[309] vdd gnd cell_6t
Xbit_r310_c123 bl[123] br[123] wl[310] vdd gnd cell_6t
Xbit_r311_c123 bl[123] br[123] wl[311] vdd gnd cell_6t
Xbit_r312_c123 bl[123] br[123] wl[312] vdd gnd cell_6t
Xbit_r313_c123 bl[123] br[123] wl[313] vdd gnd cell_6t
Xbit_r314_c123 bl[123] br[123] wl[314] vdd gnd cell_6t
Xbit_r315_c123 bl[123] br[123] wl[315] vdd gnd cell_6t
Xbit_r316_c123 bl[123] br[123] wl[316] vdd gnd cell_6t
Xbit_r317_c123 bl[123] br[123] wl[317] vdd gnd cell_6t
Xbit_r318_c123 bl[123] br[123] wl[318] vdd gnd cell_6t
Xbit_r319_c123 bl[123] br[123] wl[319] vdd gnd cell_6t
Xbit_r320_c123 bl[123] br[123] wl[320] vdd gnd cell_6t
Xbit_r321_c123 bl[123] br[123] wl[321] vdd gnd cell_6t
Xbit_r322_c123 bl[123] br[123] wl[322] vdd gnd cell_6t
Xbit_r323_c123 bl[123] br[123] wl[323] vdd gnd cell_6t
Xbit_r324_c123 bl[123] br[123] wl[324] vdd gnd cell_6t
Xbit_r325_c123 bl[123] br[123] wl[325] vdd gnd cell_6t
Xbit_r326_c123 bl[123] br[123] wl[326] vdd gnd cell_6t
Xbit_r327_c123 bl[123] br[123] wl[327] vdd gnd cell_6t
Xbit_r328_c123 bl[123] br[123] wl[328] vdd gnd cell_6t
Xbit_r329_c123 bl[123] br[123] wl[329] vdd gnd cell_6t
Xbit_r330_c123 bl[123] br[123] wl[330] vdd gnd cell_6t
Xbit_r331_c123 bl[123] br[123] wl[331] vdd gnd cell_6t
Xbit_r332_c123 bl[123] br[123] wl[332] vdd gnd cell_6t
Xbit_r333_c123 bl[123] br[123] wl[333] vdd gnd cell_6t
Xbit_r334_c123 bl[123] br[123] wl[334] vdd gnd cell_6t
Xbit_r335_c123 bl[123] br[123] wl[335] vdd gnd cell_6t
Xbit_r336_c123 bl[123] br[123] wl[336] vdd gnd cell_6t
Xbit_r337_c123 bl[123] br[123] wl[337] vdd gnd cell_6t
Xbit_r338_c123 bl[123] br[123] wl[338] vdd gnd cell_6t
Xbit_r339_c123 bl[123] br[123] wl[339] vdd gnd cell_6t
Xbit_r340_c123 bl[123] br[123] wl[340] vdd gnd cell_6t
Xbit_r341_c123 bl[123] br[123] wl[341] vdd gnd cell_6t
Xbit_r342_c123 bl[123] br[123] wl[342] vdd gnd cell_6t
Xbit_r343_c123 bl[123] br[123] wl[343] vdd gnd cell_6t
Xbit_r344_c123 bl[123] br[123] wl[344] vdd gnd cell_6t
Xbit_r345_c123 bl[123] br[123] wl[345] vdd gnd cell_6t
Xbit_r346_c123 bl[123] br[123] wl[346] vdd gnd cell_6t
Xbit_r347_c123 bl[123] br[123] wl[347] vdd gnd cell_6t
Xbit_r348_c123 bl[123] br[123] wl[348] vdd gnd cell_6t
Xbit_r349_c123 bl[123] br[123] wl[349] vdd gnd cell_6t
Xbit_r350_c123 bl[123] br[123] wl[350] vdd gnd cell_6t
Xbit_r351_c123 bl[123] br[123] wl[351] vdd gnd cell_6t
Xbit_r352_c123 bl[123] br[123] wl[352] vdd gnd cell_6t
Xbit_r353_c123 bl[123] br[123] wl[353] vdd gnd cell_6t
Xbit_r354_c123 bl[123] br[123] wl[354] vdd gnd cell_6t
Xbit_r355_c123 bl[123] br[123] wl[355] vdd gnd cell_6t
Xbit_r356_c123 bl[123] br[123] wl[356] vdd gnd cell_6t
Xbit_r357_c123 bl[123] br[123] wl[357] vdd gnd cell_6t
Xbit_r358_c123 bl[123] br[123] wl[358] vdd gnd cell_6t
Xbit_r359_c123 bl[123] br[123] wl[359] vdd gnd cell_6t
Xbit_r360_c123 bl[123] br[123] wl[360] vdd gnd cell_6t
Xbit_r361_c123 bl[123] br[123] wl[361] vdd gnd cell_6t
Xbit_r362_c123 bl[123] br[123] wl[362] vdd gnd cell_6t
Xbit_r363_c123 bl[123] br[123] wl[363] vdd gnd cell_6t
Xbit_r364_c123 bl[123] br[123] wl[364] vdd gnd cell_6t
Xbit_r365_c123 bl[123] br[123] wl[365] vdd gnd cell_6t
Xbit_r366_c123 bl[123] br[123] wl[366] vdd gnd cell_6t
Xbit_r367_c123 bl[123] br[123] wl[367] vdd gnd cell_6t
Xbit_r368_c123 bl[123] br[123] wl[368] vdd gnd cell_6t
Xbit_r369_c123 bl[123] br[123] wl[369] vdd gnd cell_6t
Xbit_r370_c123 bl[123] br[123] wl[370] vdd gnd cell_6t
Xbit_r371_c123 bl[123] br[123] wl[371] vdd gnd cell_6t
Xbit_r372_c123 bl[123] br[123] wl[372] vdd gnd cell_6t
Xbit_r373_c123 bl[123] br[123] wl[373] vdd gnd cell_6t
Xbit_r374_c123 bl[123] br[123] wl[374] vdd gnd cell_6t
Xbit_r375_c123 bl[123] br[123] wl[375] vdd gnd cell_6t
Xbit_r376_c123 bl[123] br[123] wl[376] vdd gnd cell_6t
Xbit_r377_c123 bl[123] br[123] wl[377] vdd gnd cell_6t
Xbit_r378_c123 bl[123] br[123] wl[378] vdd gnd cell_6t
Xbit_r379_c123 bl[123] br[123] wl[379] vdd gnd cell_6t
Xbit_r380_c123 bl[123] br[123] wl[380] vdd gnd cell_6t
Xbit_r381_c123 bl[123] br[123] wl[381] vdd gnd cell_6t
Xbit_r382_c123 bl[123] br[123] wl[382] vdd gnd cell_6t
Xbit_r383_c123 bl[123] br[123] wl[383] vdd gnd cell_6t
Xbit_r384_c123 bl[123] br[123] wl[384] vdd gnd cell_6t
Xbit_r385_c123 bl[123] br[123] wl[385] vdd gnd cell_6t
Xbit_r386_c123 bl[123] br[123] wl[386] vdd gnd cell_6t
Xbit_r387_c123 bl[123] br[123] wl[387] vdd gnd cell_6t
Xbit_r388_c123 bl[123] br[123] wl[388] vdd gnd cell_6t
Xbit_r389_c123 bl[123] br[123] wl[389] vdd gnd cell_6t
Xbit_r390_c123 bl[123] br[123] wl[390] vdd gnd cell_6t
Xbit_r391_c123 bl[123] br[123] wl[391] vdd gnd cell_6t
Xbit_r392_c123 bl[123] br[123] wl[392] vdd gnd cell_6t
Xbit_r393_c123 bl[123] br[123] wl[393] vdd gnd cell_6t
Xbit_r394_c123 bl[123] br[123] wl[394] vdd gnd cell_6t
Xbit_r395_c123 bl[123] br[123] wl[395] vdd gnd cell_6t
Xbit_r396_c123 bl[123] br[123] wl[396] vdd gnd cell_6t
Xbit_r397_c123 bl[123] br[123] wl[397] vdd gnd cell_6t
Xbit_r398_c123 bl[123] br[123] wl[398] vdd gnd cell_6t
Xbit_r399_c123 bl[123] br[123] wl[399] vdd gnd cell_6t
Xbit_r400_c123 bl[123] br[123] wl[400] vdd gnd cell_6t
Xbit_r401_c123 bl[123] br[123] wl[401] vdd gnd cell_6t
Xbit_r402_c123 bl[123] br[123] wl[402] vdd gnd cell_6t
Xbit_r403_c123 bl[123] br[123] wl[403] vdd gnd cell_6t
Xbit_r404_c123 bl[123] br[123] wl[404] vdd gnd cell_6t
Xbit_r405_c123 bl[123] br[123] wl[405] vdd gnd cell_6t
Xbit_r406_c123 bl[123] br[123] wl[406] vdd gnd cell_6t
Xbit_r407_c123 bl[123] br[123] wl[407] vdd gnd cell_6t
Xbit_r408_c123 bl[123] br[123] wl[408] vdd gnd cell_6t
Xbit_r409_c123 bl[123] br[123] wl[409] vdd gnd cell_6t
Xbit_r410_c123 bl[123] br[123] wl[410] vdd gnd cell_6t
Xbit_r411_c123 bl[123] br[123] wl[411] vdd gnd cell_6t
Xbit_r412_c123 bl[123] br[123] wl[412] vdd gnd cell_6t
Xbit_r413_c123 bl[123] br[123] wl[413] vdd gnd cell_6t
Xbit_r414_c123 bl[123] br[123] wl[414] vdd gnd cell_6t
Xbit_r415_c123 bl[123] br[123] wl[415] vdd gnd cell_6t
Xbit_r416_c123 bl[123] br[123] wl[416] vdd gnd cell_6t
Xbit_r417_c123 bl[123] br[123] wl[417] vdd gnd cell_6t
Xbit_r418_c123 bl[123] br[123] wl[418] vdd gnd cell_6t
Xbit_r419_c123 bl[123] br[123] wl[419] vdd gnd cell_6t
Xbit_r420_c123 bl[123] br[123] wl[420] vdd gnd cell_6t
Xbit_r421_c123 bl[123] br[123] wl[421] vdd gnd cell_6t
Xbit_r422_c123 bl[123] br[123] wl[422] vdd gnd cell_6t
Xbit_r423_c123 bl[123] br[123] wl[423] vdd gnd cell_6t
Xbit_r424_c123 bl[123] br[123] wl[424] vdd gnd cell_6t
Xbit_r425_c123 bl[123] br[123] wl[425] vdd gnd cell_6t
Xbit_r426_c123 bl[123] br[123] wl[426] vdd gnd cell_6t
Xbit_r427_c123 bl[123] br[123] wl[427] vdd gnd cell_6t
Xbit_r428_c123 bl[123] br[123] wl[428] vdd gnd cell_6t
Xbit_r429_c123 bl[123] br[123] wl[429] vdd gnd cell_6t
Xbit_r430_c123 bl[123] br[123] wl[430] vdd gnd cell_6t
Xbit_r431_c123 bl[123] br[123] wl[431] vdd gnd cell_6t
Xbit_r432_c123 bl[123] br[123] wl[432] vdd gnd cell_6t
Xbit_r433_c123 bl[123] br[123] wl[433] vdd gnd cell_6t
Xbit_r434_c123 bl[123] br[123] wl[434] vdd gnd cell_6t
Xbit_r435_c123 bl[123] br[123] wl[435] vdd gnd cell_6t
Xbit_r436_c123 bl[123] br[123] wl[436] vdd gnd cell_6t
Xbit_r437_c123 bl[123] br[123] wl[437] vdd gnd cell_6t
Xbit_r438_c123 bl[123] br[123] wl[438] vdd gnd cell_6t
Xbit_r439_c123 bl[123] br[123] wl[439] vdd gnd cell_6t
Xbit_r440_c123 bl[123] br[123] wl[440] vdd gnd cell_6t
Xbit_r441_c123 bl[123] br[123] wl[441] vdd gnd cell_6t
Xbit_r442_c123 bl[123] br[123] wl[442] vdd gnd cell_6t
Xbit_r443_c123 bl[123] br[123] wl[443] vdd gnd cell_6t
Xbit_r444_c123 bl[123] br[123] wl[444] vdd gnd cell_6t
Xbit_r445_c123 bl[123] br[123] wl[445] vdd gnd cell_6t
Xbit_r446_c123 bl[123] br[123] wl[446] vdd gnd cell_6t
Xbit_r447_c123 bl[123] br[123] wl[447] vdd gnd cell_6t
Xbit_r448_c123 bl[123] br[123] wl[448] vdd gnd cell_6t
Xbit_r449_c123 bl[123] br[123] wl[449] vdd gnd cell_6t
Xbit_r450_c123 bl[123] br[123] wl[450] vdd gnd cell_6t
Xbit_r451_c123 bl[123] br[123] wl[451] vdd gnd cell_6t
Xbit_r452_c123 bl[123] br[123] wl[452] vdd gnd cell_6t
Xbit_r453_c123 bl[123] br[123] wl[453] vdd gnd cell_6t
Xbit_r454_c123 bl[123] br[123] wl[454] vdd gnd cell_6t
Xbit_r455_c123 bl[123] br[123] wl[455] vdd gnd cell_6t
Xbit_r456_c123 bl[123] br[123] wl[456] vdd gnd cell_6t
Xbit_r457_c123 bl[123] br[123] wl[457] vdd gnd cell_6t
Xbit_r458_c123 bl[123] br[123] wl[458] vdd gnd cell_6t
Xbit_r459_c123 bl[123] br[123] wl[459] vdd gnd cell_6t
Xbit_r460_c123 bl[123] br[123] wl[460] vdd gnd cell_6t
Xbit_r461_c123 bl[123] br[123] wl[461] vdd gnd cell_6t
Xbit_r462_c123 bl[123] br[123] wl[462] vdd gnd cell_6t
Xbit_r463_c123 bl[123] br[123] wl[463] vdd gnd cell_6t
Xbit_r464_c123 bl[123] br[123] wl[464] vdd gnd cell_6t
Xbit_r465_c123 bl[123] br[123] wl[465] vdd gnd cell_6t
Xbit_r466_c123 bl[123] br[123] wl[466] vdd gnd cell_6t
Xbit_r467_c123 bl[123] br[123] wl[467] vdd gnd cell_6t
Xbit_r468_c123 bl[123] br[123] wl[468] vdd gnd cell_6t
Xbit_r469_c123 bl[123] br[123] wl[469] vdd gnd cell_6t
Xbit_r470_c123 bl[123] br[123] wl[470] vdd gnd cell_6t
Xbit_r471_c123 bl[123] br[123] wl[471] vdd gnd cell_6t
Xbit_r472_c123 bl[123] br[123] wl[472] vdd gnd cell_6t
Xbit_r473_c123 bl[123] br[123] wl[473] vdd gnd cell_6t
Xbit_r474_c123 bl[123] br[123] wl[474] vdd gnd cell_6t
Xbit_r475_c123 bl[123] br[123] wl[475] vdd gnd cell_6t
Xbit_r476_c123 bl[123] br[123] wl[476] vdd gnd cell_6t
Xbit_r477_c123 bl[123] br[123] wl[477] vdd gnd cell_6t
Xbit_r478_c123 bl[123] br[123] wl[478] vdd gnd cell_6t
Xbit_r479_c123 bl[123] br[123] wl[479] vdd gnd cell_6t
Xbit_r480_c123 bl[123] br[123] wl[480] vdd gnd cell_6t
Xbit_r481_c123 bl[123] br[123] wl[481] vdd gnd cell_6t
Xbit_r482_c123 bl[123] br[123] wl[482] vdd gnd cell_6t
Xbit_r483_c123 bl[123] br[123] wl[483] vdd gnd cell_6t
Xbit_r484_c123 bl[123] br[123] wl[484] vdd gnd cell_6t
Xbit_r485_c123 bl[123] br[123] wl[485] vdd gnd cell_6t
Xbit_r486_c123 bl[123] br[123] wl[486] vdd gnd cell_6t
Xbit_r487_c123 bl[123] br[123] wl[487] vdd gnd cell_6t
Xbit_r488_c123 bl[123] br[123] wl[488] vdd gnd cell_6t
Xbit_r489_c123 bl[123] br[123] wl[489] vdd gnd cell_6t
Xbit_r490_c123 bl[123] br[123] wl[490] vdd gnd cell_6t
Xbit_r491_c123 bl[123] br[123] wl[491] vdd gnd cell_6t
Xbit_r492_c123 bl[123] br[123] wl[492] vdd gnd cell_6t
Xbit_r493_c123 bl[123] br[123] wl[493] vdd gnd cell_6t
Xbit_r494_c123 bl[123] br[123] wl[494] vdd gnd cell_6t
Xbit_r495_c123 bl[123] br[123] wl[495] vdd gnd cell_6t
Xbit_r496_c123 bl[123] br[123] wl[496] vdd gnd cell_6t
Xbit_r497_c123 bl[123] br[123] wl[497] vdd gnd cell_6t
Xbit_r498_c123 bl[123] br[123] wl[498] vdd gnd cell_6t
Xbit_r499_c123 bl[123] br[123] wl[499] vdd gnd cell_6t
Xbit_r500_c123 bl[123] br[123] wl[500] vdd gnd cell_6t
Xbit_r501_c123 bl[123] br[123] wl[501] vdd gnd cell_6t
Xbit_r502_c123 bl[123] br[123] wl[502] vdd gnd cell_6t
Xbit_r503_c123 bl[123] br[123] wl[503] vdd gnd cell_6t
Xbit_r504_c123 bl[123] br[123] wl[504] vdd gnd cell_6t
Xbit_r505_c123 bl[123] br[123] wl[505] vdd gnd cell_6t
Xbit_r506_c123 bl[123] br[123] wl[506] vdd gnd cell_6t
Xbit_r507_c123 bl[123] br[123] wl[507] vdd gnd cell_6t
Xbit_r508_c123 bl[123] br[123] wl[508] vdd gnd cell_6t
Xbit_r509_c123 bl[123] br[123] wl[509] vdd gnd cell_6t
Xbit_r510_c123 bl[123] br[123] wl[510] vdd gnd cell_6t
Xbit_r511_c123 bl[123] br[123] wl[511] vdd gnd cell_6t
Xbit_r0_c124 bl[124] br[124] wl[0] vdd gnd cell_6t
Xbit_r1_c124 bl[124] br[124] wl[1] vdd gnd cell_6t
Xbit_r2_c124 bl[124] br[124] wl[2] vdd gnd cell_6t
Xbit_r3_c124 bl[124] br[124] wl[3] vdd gnd cell_6t
Xbit_r4_c124 bl[124] br[124] wl[4] vdd gnd cell_6t
Xbit_r5_c124 bl[124] br[124] wl[5] vdd gnd cell_6t
Xbit_r6_c124 bl[124] br[124] wl[6] vdd gnd cell_6t
Xbit_r7_c124 bl[124] br[124] wl[7] vdd gnd cell_6t
Xbit_r8_c124 bl[124] br[124] wl[8] vdd gnd cell_6t
Xbit_r9_c124 bl[124] br[124] wl[9] vdd gnd cell_6t
Xbit_r10_c124 bl[124] br[124] wl[10] vdd gnd cell_6t
Xbit_r11_c124 bl[124] br[124] wl[11] vdd gnd cell_6t
Xbit_r12_c124 bl[124] br[124] wl[12] vdd gnd cell_6t
Xbit_r13_c124 bl[124] br[124] wl[13] vdd gnd cell_6t
Xbit_r14_c124 bl[124] br[124] wl[14] vdd gnd cell_6t
Xbit_r15_c124 bl[124] br[124] wl[15] vdd gnd cell_6t
Xbit_r16_c124 bl[124] br[124] wl[16] vdd gnd cell_6t
Xbit_r17_c124 bl[124] br[124] wl[17] vdd gnd cell_6t
Xbit_r18_c124 bl[124] br[124] wl[18] vdd gnd cell_6t
Xbit_r19_c124 bl[124] br[124] wl[19] vdd gnd cell_6t
Xbit_r20_c124 bl[124] br[124] wl[20] vdd gnd cell_6t
Xbit_r21_c124 bl[124] br[124] wl[21] vdd gnd cell_6t
Xbit_r22_c124 bl[124] br[124] wl[22] vdd gnd cell_6t
Xbit_r23_c124 bl[124] br[124] wl[23] vdd gnd cell_6t
Xbit_r24_c124 bl[124] br[124] wl[24] vdd gnd cell_6t
Xbit_r25_c124 bl[124] br[124] wl[25] vdd gnd cell_6t
Xbit_r26_c124 bl[124] br[124] wl[26] vdd gnd cell_6t
Xbit_r27_c124 bl[124] br[124] wl[27] vdd gnd cell_6t
Xbit_r28_c124 bl[124] br[124] wl[28] vdd gnd cell_6t
Xbit_r29_c124 bl[124] br[124] wl[29] vdd gnd cell_6t
Xbit_r30_c124 bl[124] br[124] wl[30] vdd gnd cell_6t
Xbit_r31_c124 bl[124] br[124] wl[31] vdd gnd cell_6t
Xbit_r32_c124 bl[124] br[124] wl[32] vdd gnd cell_6t
Xbit_r33_c124 bl[124] br[124] wl[33] vdd gnd cell_6t
Xbit_r34_c124 bl[124] br[124] wl[34] vdd gnd cell_6t
Xbit_r35_c124 bl[124] br[124] wl[35] vdd gnd cell_6t
Xbit_r36_c124 bl[124] br[124] wl[36] vdd gnd cell_6t
Xbit_r37_c124 bl[124] br[124] wl[37] vdd gnd cell_6t
Xbit_r38_c124 bl[124] br[124] wl[38] vdd gnd cell_6t
Xbit_r39_c124 bl[124] br[124] wl[39] vdd gnd cell_6t
Xbit_r40_c124 bl[124] br[124] wl[40] vdd gnd cell_6t
Xbit_r41_c124 bl[124] br[124] wl[41] vdd gnd cell_6t
Xbit_r42_c124 bl[124] br[124] wl[42] vdd gnd cell_6t
Xbit_r43_c124 bl[124] br[124] wl[43] vdd gnd cell_6t
Xbit_r44_c124 bl[124] br[124] wl[44] vdd gnd cell_6t
Xbit_r45_c124 bl[124] br[124] wl[45] vdd gnd cell_6t
Xbit_r46_c124 bl[124] br[124] wl[46] vdd gnd cell_6t
Xbit_r47_c124 bl[124] br[124] wl[47] vdd gnd cell_6t
Xbit_r48_c124 bl[124] br[124] wl[48] vdd gnd cell_6t
Xbit_r49_c124 bl[124] br[124] wl[49] vdd gnd cell_6t
Xbit_r50_c124 bl[124] br[124] wl[50] vdd gnd cell_6t
Xbit_r51_c124 bl[124] br[124] wl[51] vdd gnd cell_6t
Xbit_r52_c124 bl[124] br[124] wl[52] vdd gnd cell_6t
Xbit_r53_c124 bl[124] br[124] wl[53] vdd gnd cell_6t
Xbit_r54_c124 bl[124] br[124] wl[54] vdd gnd cell_6t
Xbit_r55_c124 bl[124] br[124] wl[55] vdd gnd cell_6t
Xbit_r56_c124 bl[124] br[124] wl[56] vdd gnd cell_6t
Xbit_r57_c124 bl[124] br[124] wl[57] vdd gnd cell_6t
Xbit_r58_c124 bl[124] br[124] wl[58] vdd gnd cell_6t
Xbit_r59_c124 bl[124] br[124] wl[59] vdd gnd cell_6t
Xbit_r60_c124 bl[124] br[124] wl[60] vdd gnd cell_6t
Xbit_r61_c124 bl[124] br[124] wl[61] vdd gnd cell_6t
Xbit_r62_c124 bl[124] br[124] wl[62] vdd gnd cell_6t
Xbit_r63_c124 bl[124] br[124] wl[63] vdd gnd cell_6t
Xbit_r64_c124 bl[124] br[124] wl[64] vdd gnd cell_6t
Xbit_r65_c124 bl[124] br[124] wl[65] vdd gnd cell_6t
Xbit_r66_c124 bl[124] br[124] wl[66] vdd gnd cell_6t
Xbit_r67_c124 bl[124] br[124] wl[67] vdd gnd cell_6t
Xbit_r68_c124 bl[124] br[124] wl[68] vdd gnd cell_6t
Xbit_r69_c124 bl[124] br[124] wl[69] vdd gnd cell_6t
Xbit_r70_c124 bl[124] br[124] wl[70] vdd gnd cell_6t
Xbit_r71_c124 bl[124] br[124] wl[71] vdd gnd cell_6t
Xbit_r72_c124 bl[124] br[124] wl[72] vdd gnd cell_6t
Xbit_r73_c124 bl[124] br[124] wl[73] vdd gnd cell_6t
Xbit_r74_c124 bl[124] br[124] wl[74] vdd gnd cell_6t
Xbit_r75_c124 bl[124] br[124] wl[75] vdd gnd cell_6t
Xbit_r76_c124 bl[124] br[124] wl[76] vdd gnd cell_6t
Xbit_r77_c124 bl[124] br[124] wl[77] vdd gnd cell_6t
Xbit_r78_c124 bl[124] br[124] wl[78] vdd gnd cell_6t
Xbit_r79_c124 bl[124] br[124] wl[79] vdd gnd cell_6t
Xbit_r80_c124 bl[124] br[124] wl[80] vdd gnd cell_6t
Xbit_r81_c124 bl[124] br[124] wl[81] vdd gnd cell_6t
Xbit_r82_c124 bl[124] br[124] wl[82] vdd gnd cell_6t
Xbit_r83_c124 bl[124] br[124] wl[83] vdd gnd cell_6t
Xbit_r84_c124 bl[124] br[124] wl[84] vdd gnd cell_6t
Xbit_r85_c124 bl[124] br[124] wl[85] vdd gnd cell_6t
Xbit_r86_c124 bl[124] br[124] wl[86] vdd gnd cell_6t
Xbit_r87_c124 bl[124] br[124] wl[87] vdd gnd cell_6t
Xbit_r88_c124 bl[124] br[124] wl[88] vdd gnd cell_6t
Xbit_r89_c124 bl[124] br[124] wl[89] vdd gnd cell_6t
Xbit_r90_c124 bl[124] br[124] wl[90] vdd gnd cell_6t
Xbit_r91_c124 bl[124] br[124] wl[91] vdd gnd cell_6t
Xbit_r92_c124 bl[124] br[124] wl[92] vdd gnd cell_6t
Xbit_r93_c124 bl[124] br[124] wl[93] vdd gnd cell_6t
Xbit_r94_c124 bl[124] br[124] wl[94] vdd gnd cell_6t
Xbit_r95_c124 bl[124] br[124] wl[95] vdd gnd cell_6t
Xbit_r96_c124 bl[124] br[124] wl[96] vdd gnd cell_6t
Xbit_r97_c124 bl[124] br[124] wl[97] vdd gnd cell_6t
Xbit_r98_c124 bl[124] br[124] wl[98] vdd gnd cell_6t
Xbit_r99_c124 bl[124] br[124] wl[99] vdd gnd cell_6t
Xbit_r100_c124 bl[124] br[124] wl[100] vdd gnd cell_6t
Xbit_r101_c124 bl[124] br[124] wl[101] vdd gnd cell_6t
Xbit_r102_c124 bl[124] br[124] wl[102] vdd gnd cell_6t
Xbit_r103_c124 bl[124] br[124] wl[103] vdd gnd cell_6t
Xbit_r104_c124 bl[124] br[124] wl[104] vdd gnd cell_6t
Xbit_r105_c124 bl[124] br[124] wl[105] vdd gnd cell_6t
Xbit_r106_c124 bl[124] br[124] wl[106] vdd gnd cell_6t
Xbit_r107_c124 bl[124] br[124] wl[107] vdd gnd cell_6t
Xbit_r108_c124 bl[124] br[124] wl[108] vdd gnd cell_6t
Xbit_r109_c124 bl[124] br[124] wl[109] vdd gnd cell_6t
Xbit_r110_c124 bl[124] br[124] wl[110] vdd gnd cell_6t
Xbit_r111_c124 bl[124] br[124] wl[111] vdd gnd cell_6t
Xbit_r112_c124 bl[124] br[124] wl[112] vdd gnd cell_6t
Xbit_r113_c124 bl[124] br[124] wl[113] vdd gnd cell_6t
Xbit_r114_c124 bl[124] br[124] wl[114] vdd gnd cell_6t
Xbit_r115_c124 bl[124] br[124] wl[115] vdd gnd cell_6t
Xbit_r116_c124 bl[124] br[124] wl[116] vdd gnd cell_6t
Xbit_r117_c124 bl[124] br[124] wl[117] vdd gnd cell_6t
Xbit_r118_c124 bl[124] br[124] wl[118] vdd gnd cell_6t
Xbit_r119_c124 bl[124] br[124] wl[119] vdd gnd cell_6t
Xbit_r120_c124 bl[124] br[124] wl[120] vdd gnd cell_6t
Xbit_r121_c124 bl[124] br[124] wl[121] vdd gnd cell_6t
Xbit_r122_c124 bl[124] br[124] wl[122] vdd gnd cell_6t
Xbit_r123_c124 bl[124] br[124] wl[123] vdd gnd cell_6t
Xbit_r124_c124 bl[124] br[124] wl[124] vdd gnd cell_6t
Xbit_r125_c124 bl[124] br[124] wl[125] vdd gnd cell_6t
Xbit_r126_c124 bl[124] br[124] wl[126] vdd gnd cell_6t
Xbit_r127_c124 bl[124] br[124] wl[127] vdd gnd cell_6t
Xbit_r128_c124 bl[124] br[124] wl[128] vdd gnd cell_6t
Xbit_r129_c124 bl[124] br[124] wl[129] vdd gnd cell_6t
Xbit_r130_c124 bl[124] br[124] wl[130] vdd gnd cell_6t
Xbit_r131_c124 bl[124] br[124] wl[131] vdd gnd cell_6t
Xbit_r132_c124 bl[124] br[124] wl[132] vdd gnd cell_6t
Xbit_r133_c124 bl[124] br[124] wl[133] vdd gnd cell_6t
Xbit_r134_c124 bl[124] br[124] wl[134] vdd gnd cell_6t
Xbit_r135_c124 bl[124] br[124] wl[135] vdd gnd cell_6t
Xbit_r136_c124 bl[124] br[124] wl[136] vdd gnd cell_6t
Xbit_r137_c124 bl[124] br[124] wl[137] vdd gnd cell_6t
Xbit_r138_c124 bl[124] br[124] wl[138] vdd gnd cell_6t
Xbit_r139_c124 bl[124] br[124] wl[139] vdd gnd cell_6t
Xbit_r140_c124 bl[124] br[124] wl[140] vdd gnd cell_6t
Xbit_r141_c124 bl[124] br[124] wl[141] vdd gnd cell_6t
Xbit_r142_c124 bl[124] br[124] wl[142] vdd gnd cell_6t
Xbit_r143_c124 bl[124] br[124] wl[143] vdd gnd cell_6t
Xbit_r144_c124 bl[124] br[124] wl[144] vdd gnd cell_6t
Xbit_r145_c124 bl[124] br[124] wl[145] vdd gnd cell_6t
Xbit_r146_c124 bl[124] br[124] wl[146] vdd gnd cell_6t
Xbit_r147_c124 bl[124] br[124] wl[147] vdd gnd cell_6t
Xbit_r148_c124 bl[124] br[124] wl[148] vdd gnd cell_6t
Xbit_r149_c124 bl[124] br[124] wl[149] vdd gnd cell_6t
Xbit_r150_c124 bl[124] br[124] wl[150] vdd gnd cell_6t
Xbit_r151_c124 bl[124] br[124] wl[151] vdd gnd cell_6t
Xbit_r152_c124 bl[124] br[124] wl[152] vdd gnd cell_6t
Xbit_r153_c124 bl[124] br[124] wl[153] vdd gnd cell_6t
Xbit_r154_c124 bl[124] br[124] wl[154] vdd gnd cell_6t
Xbit_r155_c124 bl[124] br[124] wl[155] vdd gnd cell_6t
Xbit_r156_c124 bl[124] br[124] wl[156] vdd gnd cell_6t
Xbit_r157_c124 bl[124] br[124] wl[157] vdd gnd cell_6t
Xbit_r158_c124 bl[124] br[124] wl[158] vdd gnd cell_6t
Xbit_r159_c124 bl[124] br[124] wl[159] vdd gnd cell_6t
Xbit_r160_c124 bl[124] br[124] wl[160] vdd gnd cell_6t
Xbit_r161_c124 bl[124] br[124] wl[161] vdd gnd cell_6t
Xbit_r162_c124 bl[124] br[124] wl[162] vdd gnd cell_6t
Xbit_r163_c124 bl[124] br[124] wl[163] vdd gnd cell_6t
Xbit_r164_c124 bl[124] br[124] wl[164] vdd gnd cell_6t
Xbit_r165_c124 bl[124] br[124] wl[165] vdd gnd cell_6t
Xbit_r166_c124 bl[124] br[124] wl[166] vdd gnd cell_6t
Xbit_r167_c124 bl[124] br[124] wl[167] vdd gnd cell_6t
Xbit_r168_c124 bl[124] br[124] wl[168] vdd gnd cell_6t
Xbit_r169_c124 bl[124] br[124] wl[169] vdd gnd cell_6t
Xbit_r170_c124 bl[124] br[124] wl[170] vdd gnd cell_6t
Xbit_r171_c124 bl[124] br[124] wl[171] vdd gnd cell_6t
Xbit_r172_c124 bl[124] br[124] wl[172] vdd gnd cell_6t
Xbit_r173_c124 bl[124] br[124] wl[173] vdd gnd cell_6t
Xbit_r174_c124 bl[124] br[124] wl[174] vdd gnd cell_6t
Xbit_r175_c124 bl[124] br[124] wl[175] vdd gnd cell_6t
Xbit_r176_c124 bl[124] br[124] wl[176] vdd gnd cell_6t
Xbit_r177_c124 bl[124] br[124] wl[177] vdd gnd cell_6t
Xbit_r178_c124 bl[124] br[124] wl[178] vdd gnd cell_6t
Xbit_r179_c124 bl[124] br[124] wl[179] vdd gnd cell_6t
Xbit_r180_c124 bl[124] br[124] wl[180] vdd gnd cell_6t
Xbit_r181_c124 bl[124] br[124] wl[181] vdd gnd cell_6t
Xbit_r182_c124 bl[124] br[124] wl[182] vdd gnd cell_6t
Xbit_r183_c124 bl[124] br[124] wl[183] vdd gnd cell_6t
Xbit_r184_c124 bl[124] br[124] wl[184] vdd gnd cell_6t
Xbit_r185_c124 bl[124] br[124] wl[185] vdd gnd cell_6t
Xbit_r186_c124 bl[124] br[124] wl[186] vdd gnd cell_6t
Xbit_r187_c124 bl[124] br[124] wl[187] vdd gnd cell_6t
Xbit_r188_c124 bl[124] br[124] wl[188] vdd gnd cell_6t
Xbit_r189_c124 bl[124] br[124] wl[189] vdd gnd cell_6t
Xbit_r190_c124 bl[124] br[124] wl[190] vdd gnd cell_6t
Xbit_r191_c124 bl[124] br[124] wl[191] vdd gnd cell_6t
Xbit_r192_c124 bl[124] br[124] wl[192] vdd gnd cell_6t
Xbit_r193_c124 bl[124] br[124] wl[193] vdd gnd cell_6t
Xbit_r194_c124 bl[124] br[124] wl[194] vdd gnd cell_6t
Xbit_r195_c124 bl[124] br[124] wl[195] vdd gnd cell_6t
Xbit_r196_c124 bl[124] br[124] wl[196] vdd gnd cell_6t
Xbit_r197_c124 bl[124] br[124] wl[197] vdd gnd cell_6t
Xbit_r198_c124 bl[124] br[124] wl[198] vdd gnd cell_6t
Xbit_r199_c124 bl[124] br[124] wl[199] vdd gnd cell_6t
Xbit_r200_c124 bl[124] br[124] wl[200] vdd gnd cell_6t
Xbit_r201_c124 bl[124] br[124] wl[201] vdd gnd cell_6t
Xbit_r202_c124 bl[124] br[124] wl[202] vdd gnd cell_6t
Xbit_r203_c124 bl[124] br[124] wl[203] vdd gnd cell_6t
Xbit_r204_c124 bl[124] br[124] wl[204] vdd gnd cell_6t
Xbit_r205_c124 bl[124] br[124] wl[205] vdd gnd cell_6t
Xbit_r206_c124 bl[124] br[124] wl[206] vdd gnd cell_6t
Xbit_r207_c124 bl[124] br[124] wl[207] vdd gnd cell_6t
Xbit_r208_c124 bl[124] br[124] wl[208] vdd gnd cell_6t
Xbit_r209_c124 bl[124] br[124] wl[209] vdd gnd cell_6t
Xbit_r210_c124 bl[124] br[124] wl[210] vdd gnd cell_6t
Xbit_r211_c124 bl[124] br[124] wl[211] vdd gnd cell_6t
Xbit_r212_c124 bl[124] br[124] wl[212] vdd gnd cell_6t
Xbit_r213_c124 bl[124] br[124] wl[213] vdd gnd cell_6t
Xbit_r214_c124 bl[124] br[124] wl[214] vdd gnd cell_6t
Xbit_r215_c124 bl[124] br[124] wl[215] vdd gnd cell_6t
Xbit_r216_c124 bl[124] br[124] wl[216] vdd gnd cell_6t
Xbit_r217_c124 bl[124] br[124] wl[217] vdd gnd cell_6t
Xbit_r218_c124 bl[124] br[124] wl[218] vdd gnd cell_6t
Xbit_r219_c124 bl[124] br[124] wl[219] vdd gnd cell_6t
Xbit_r220_c124 bl[124] br[124] wl[220] vdd gnd cell_6t
Xbit_r221_c124 bl[124] br[124] wl[221] vdd gnd cell_6t
Xbit_r222_c124 bl[124] br[124] wl[222] vdd gnd cell_6t
Xbit_r223_c124 bl[124] br[124] wl[223] vdd gnd cell_6t
Xbit_r224_c124 bl[124] br[124] wl[224] vdd gnd cell_6t
Xbit_r225_c124 bl[124] br[124] wl[225] vdd gnd cell_6t
Xbit_r226_c124 bl[124] br[124] wl[226] vdd gnd cell_6t
Xbit_r227_c124 bl[124] br[124] wl[227] vdd gnd cell_6t
Xbit_r228_c124 bl[124] br[124] wl[228] vdd gnd cell_6t
Xbit_r229_c124 bl[124] br[124] wl[229] vdd gnd cell_6t
Xbit_r230_c124 bl[124] br[124] wl[230] vdd gnd cell_6t
Xbit_r231_c124 bl[124] br[124] wl[231] vdd gnd cell_6t
Xbit_r232_c124 bl[124] br[124] wl[232] vdd gnd cell_6t
Xbit_r233_c124 bl[124] br[124] wl[233] vdd gnd cell_6t
Xbit_r234_c124 bl[124] br[124] wl[234] vdd gnd cell_6t
Xbit_r235_c124 bl[124] br[124] wl[235] vdd gnd cell_6t
Xbit_r236_c124 bl[124] br[124] wl[236] vdd gnd cell_6t
Xbit_r237_c124 bl[124] br[124] wl[237] vdd gnd cell_6t
Xbit_r238_c124 bl[124] br[124] wl[238] vdd gnd cell_6t
Xbit_r239_c124 bl[124] br[124] wl[239] vdd gnd cell_6t
Xbit_r240_c124 bl[124] br[124] wl[240] vdd gnd cell_6t
Xbit_r241_c124 bl[124] br[124] wl[241] vdd gnd cell_6t
Xbit_r242_c124 bl[124] br[124] wl[242] vdd gnd cell_6t
Xbit_r243_c124 bl[124] br[124] wl[243] vdd gnd cell_6t
Xbit_r244_c124 bl[124] br[124] wl[244] vdd gnd cell_6t
Xbit_r245_c124 bl[124] br[124] wl[245] vdd gnd cell_6t
Xbit_r246_c124 bl[124] br[124] wl[246] vdd gnd cell_6t
Xbit_r247_c124 bl[124] br[124] wl[247] vdd gnd cell_6t
Xbit_r248_c124 bl[124] br[124] wl[248] vdd gnd cell_6t
Xbit_r249_c124 bl[124] br[124] wl[249] vdd gnd cell_6t
Xbit_r250_c124 bl[124] br[124] wl[250] vdd gnd cell_6t
Xbit_r251_c124 bl[124] br[124] wl[251] vdd gnd cell_6t
Xbit_r252_c124 bl[124] br[124] wl[252] vdd gnd cell_6t
Xbit_r253_c124 bl[124] br[124] wl[253] vdd gnd cell_6t
Xbit_r254_c124 bl[124] br[124] wl[254] vdd gnd cell_6t
Xbit_r255_c124 bl[124] br[124] wl[255] vdd gnd cell_6t
Xbit_r256_c124 bl[124] br[124] wl[256] vdd gnd cell_6t
Xbit_r257_c124 bl[124] br[124] wl[257] vdd gnd cell_6t
Xbit_r258_c124 bl[124] br[124] wl[258] vdd gnd cell_6t
Xbit_r259_c124 bl[124] br[124] wl[259] vdd gnd cell_6t
Xbit_r260_c124 bl[124] br[124] wl[260] vdd gnd cell_6t
Xbit_r261_c124 bl[124] br[124] wl[261] vdd gnd cell_6t
Xbit_r262_c124 bl[124] br[124] wl[262] vdd gnd cell_6t
Xbit_r263_c124 bl[124] br[124] wl[263] vdd gnd cell_6t
Xbit_r264_c124 bl[124] br[124] wl[264] vdd gnd cell_6t
Xbit_r265_c124 bl[124] br[124] wl[265] vdd gnd cell_6t
Xbit_r266_c124 bl[124] br[124] wl[266] vdd gnd cell_6t
Xbit_r267_c124 bl[124] br[124] wl[267] vdd gnd cell_6t
Xbit_r268_c124 bl[124] br[124] wl[268] vdd gnd cell_6t
Xbit_r269_c124 bl[124] br[124] wl[269] vdd gnd cell_6t
Xbit_r270_c124 bl[124] br[124] wl[270] vdd gnd cell_6t
Xbit_r271_c124 bl[124] br[124] wl[271] vdd gnd cell_6t
Xbit_r272_c124 bl[124] br[124] wl[272] vdd gnd cell_6t
Xbit_r273_c124 bl[124] br[124] wl[273] vdd gnd cell_6t
Xbit_r274_c124 bl[124] br[124] wl[274] vdd gnd cell_6t
Xbit_r275_c124 bl[124] br[124] wl[275] vdd gnd cell_6t
Xbit_r276_c124 bl[124] br[124] wl[276] vdd gnd cell_6t
Xbit_r277_c124 bl[124] br[124] wl[277] vdd gnd cell_6t
Xbit_r278_c124 bl[124] br[124] wl[278] vdd gnd cell_6t
Xbit_r279_c124 bl[124] br[124] wl[279] vdd gnd cell_6t
Xbit_r280_c124 bl[124] br[124] wl[280] vdd gnd cell_6t
Xbit_r281_c124 bl[124] br[124] wl[281] vdd gnd cell_6t
Xbit_r282_c124 bl[124] br[124] wl[282] vdd gnd cell_6t
Xbit_r283_c124 bl[124] br[124] wl[283] vdd gnd cell_6t
Xbit_r284_c124 bl[124] br[124] wl[284] vdd gnd cell_6t
Xbit_r285_c124 bl[124] br[124] wl[285] vdd gnd cell_6t
Xbit_r286_c124 bl[124] br[124] wl[286] vdd gnd cell_6t
Xbit_r287_c124 bl[124] br[124] wl[287] vdd gnd cell_6t
Xbit_r288_c124 bl[124] br[124] wl[288] vdd gnd cell_6t
Xbit_r289_c124 bl[124] br[124] wl[289] vdd gnd cell_6t
Xbit_r290_c124 bl[124] br[124] wl[290] vdd gnd cell_6t
Xbit_r291_c124 bl[124] br[124] wl[291] vdd gnd cell_6t
Xbit_r292_c124 bl[124] br[124] wl[292] vdd gnd cell_6t
Xbit_r293_c124 bl[124] br[124] wl[293] vdd gnd cell_6t
Xbit_r294_c124 bl[124] br[124] wl[294] vdd gnd cell_6t
Xbit_r295_c124 bl[124] br[124] wl[295] vdd gnd cell_6t
Xbit_r296_c124 bl[124] br[124] wl[296] vdd gnd cell_6t
Xbit_r297_c124 bl[124] br[124] wl[297] vdd gnd cell_6t
Xbit_r298_c124 bl[124] br[124] wl[298] vdd gnd cell_6t
Xbit_r299_c124 bl[124] br[124] wl[299] vdd gnd cell_6t
Xbit_r300_c124 bl[124] br[124] wl[300] vdd gnd cell_6t
Xbit_r301_c124 bl[124] br[124] wl[301] vdd gnd cell_6t
Xbit_r302_c124 bl[124] br[124] wl[302] vdd gnd cell_6t
Xbit_r303_c124 bl[124] br[124] wl[303] vdd gnd cell_6t
Xbit_r304_c124 bl[124] br[124] wl[304] vdd gnd cell_6t
Xbit_r305_c124 bl[124] br[124] wl[305] vdd gnd cell_6t
Xbit_r306_c124 bl[124] br[124] wl[306] vdd gnd cell_6t
Xbit_r307_c124 bl[124] br[124] wl[307] vdd gnd cell_6t
Xbit_r308_c124 bl[124] br[124] wl[308] vdd gnd cell_6t
Xbit_r309_c124 bl[124] br[124] wl[309] vdd gnd cell_6t
Xbit_r310_c124 bl[124] br[124] wl[310] vdd gnd cell_6t
Xbit_r311_c124 bl[124] br[124] wl[311] vdd gnd cell_6t
Xbit_r312_c124 bl[124] br[124] wl[312] vdd gnd cell_6t
Xbit_r313_c124 bl[124] br[124] wl[313] vdd gnd cell_6t
Xbit_r314_c124 bl[124] br[124] wl[314] vdd gnd cell_6t
Xbit_r315_c124 bl[124] br[124] wl[315] vdd gnd cell_6t
Xbit_r316_c124 bl[124] br[124] wl[316] vdd gnd cell_6t
Xbit_r317_c124 bl[124] br[124] wl[317] vdd gnd cell_6t
Xbit_r318_c124 bl[124] br[124] wl[318] vdd gnd cell_6t
Xbit_r319_c124 bl[124] br[124] wl[319] vdd gnd cell_6t
Xbit_r320_c124 bl[124] br[124] wl[320] vdd gnd cell_6t
Xbit_r321_c124 bl[124] br[124] wl[321] vdd gnd cell_6t
Xbit_r322_c124 bl[124] br[124] wl[322] vdd gnd cell_6t
Xbit_r323_c124 bl[124] br[124] wl[323] vdd gnd cell_6t
Xbit_r324_c124 bl[124] br[124] wl[324] vdd gnd cell_6t
Xbit_r325_c124 bl[124] br[124] wl[325] vdd gnd cell_6t
Xbit_r326_c124 bl[124] br[124] wl[326] vdd gnd cell_6t
Xbit_r327_c124 bl[124] br[124] wl[327] vdd gnd cell_6t
Xbit_r328_c124 bl[124] br[124] wl[328] vdd gnd cell_6t
Xbit_r329_c124 bl[124] br[124] wl[329] vdd gnd cell_6t
Xbit_r330_c124 bl[124] br[124] wl[330] vdd gnd cell_6t
Xbit_r331_c124 bl[124] br[124] wl[331] vdd gnd cell_6t
Xbit_r332_c124 bl[124] br[124] wl[332] vdd gnd cell_6t
Xbit_r333_c124 bl[124] br[124] wl[333] vdd gnd cell_6t
Xbit_r334_c124 bl[124] br[124] wl[334] vdd gnd cell_6t
Xbit_r335_c124 bl[124] br[124] wl[335] vdd gnd cell_6t
Xbit_r336_c124 bl[124] br[124] wl[336] vdd gnd cell_6t
Xbit_r337_c124 bl[124] br[124] wl[337] vdd gnd cell_6t
Xbit_r338_c124 bl[124] br[124] wl[338] vdd gnd cell_6t
Xbit_r339_c124 bl[124] br[124] wl[339] vdd gnd cell_6t
Xbit_r340_c124 bl[124] br[124] wl[340] vdd gnd cell_6t
Xbit_r341_c124 bl[124] br[124] wl[341] vdd gnd cell_6t
Xbit_r342_c124 bl[124] br[124] wl[342] vdd gnd cell_6t
Xbit_r343_c124 bl[124] br[124] wl[343] vdd gnd cell_6t
Xbit_r344_c124 bl[124] br[124] wl[344] vdd gnd cell_6t
Xbit_r345_c124 bl[124] br[124] wl[345] vdd gnd cell_6t
Xbit_r346_c124 bl[124] br[124] wl[346] vdd gnd cell_6t
Xbit_r347_c124 bl[124] br[124] wl[347] vdd gnd cell_6t
Xbit_r348_c124 bl[124] br[124] wl[348] vdd gnd cell_6t
Xbit_r349_c124 bl[124] br[124] wl[349] vdd gnd cell_6t
Xbit_r350_c124 bl[124] br[124] wl[350] vdd gnd cell_6t
Xbit_r351_c124 bl[124] br[124] wl[351] vdd gnd cell_6t
Xbit_r352_c124 bl[124] br[124] wl[352] vdd gnd cell_6t
Xbit_r353_c124 bl[124] br[124] wl[353] vdd gnd cell_6t
Xbit_r354_c124 bl[124] br[124] wl[354] vdd gnd cell_6t
Xbit_r355_c124 bl[124] br[124] wl[355] vdd gnd cell_6t
Xbit_r356_c124 bl[124] br[124] wl[356] vdd gnd cell_6t
Xbit_r357_c124 bl[124] br[124] wl[357] vdd gnd cell_6t
Xbit_r358_c124 bl[124] br[124] wl[358] vdd gnd cell_6t
Xbit_r359_c124 bl[124] br[124] wl[359] vdd gnd cell_6t
Xbit_r360_c124 bl[124] br[124] wl[360] vdd gnd cell_6t
Xbit_r361_c124 bl[124] br[124] wl[361] vdd gnd cell_6t
Xbit_r362_c124 bl[124] br[124] wl[362] vdd gnd cell_6t
Xbit_r363_c124 bl[124] br[124] wl[363] vdd gnd cell_6t
Xbit_r364_c124 bl[124] br[124] wl[364] vdd gnd cell_6t
Xbit_r365_c124 bl[124] br[124] wl[365] vdd gnd cell_6t
Xbit_r366_c124 bl[124] br[124] wl[366] vdd gnd cell_6t
Xbit_r367_c124 bl[124] br[124] wl[367] vdd gnd cell_6t
Xbit_r368_c124 bl[124] br[124] wl[368] vdd gnd cell_6t
Xbit_r369_c124 bl[124] br[124] wl[369] vdd gnd cell_6t
Xbit_r370_c124 bl[124] br[124] wl[370] vdd gnd cell_6t
Xbit_r371_c124 bl[124] br[124] wl[371] vdd gnd cell_6t
Xbit_r372_c124 bl[124] br[124] wl[372] vdd gnd cell_6t
Xbit_r373_c124 bl[124] br[124] wl[373] vdd gnd cell_6t
Xbit_r374_c124 bl[124] br[124] wl[374] vdd gnd cell_6t
Xbit_r375_c124 bl[124] br[124] wl[375] vdd gnd cell_6t
Xbit_r376_c124 bl[124] br[124] wl[376] vdd gnd cell_6t
Xbit_r377_c124 bl[124] br[124] wl[377] vdd gnd cell_6t
Xbit_r378_c124 bl[124] br[124] wl[378] vdd gnd cell_6t
Xbit_r379_c124 bl[124] br[124] wl[379] vdd gnd cell_6t
Xbit_r380_c124 bl[124] br[124] wl[380] vdd gnd cell_6t
Xbit_r381_c124 bl[124] br[124] wl[381] vdd gnd cell_6t
Xbit_r382_c124 bl[124] br[124] wl[382] vdd gnd cell_6t
Xbit_r383_c124 bl[124] br[124] wl[383] vdd gnd cell_6t
Xbit_r384_c124 bl[124] br[124] wl[384] vdd gnd cell_6t
Xbit_r385_c124 bl[124] br[124] wl[385] vdd gnd cell_6t
Xbit_r386_c124 bl[124] br[124] wl[386] vdd gnd cell_6t
Xbit_r387_c124 bl[124] br[124] wl[387] vdd gnd cell_6t
Xbit_r388_c124 bl[124] br[124] wl[388] vdd gnd cell_6t
Xbit_r389_c124 bl[124] br[124] wl[389] vdd gnd cell_6t
Xbit_r390_c124 bl[124] br[124] wl[390] vdd gnd cell_6t
Xbit_r391_c124 bl[124] br[124] wl[391] vdd gnd cell_6t
Xbit_r392_c124 bl[124] br[124] wl[392] vdd gnd cell_6t
Xbit_r393_c124 bl[124] br[124] wl[393] vdd gnd cell_6t
Xbit_r394_c124 bl[124] br[124] wl[394] vdd gnd cell_6t
Xbit_r395_c124 bl[124] br[124] wl[395] vdd gnd cell_6t
Xbit_r396_c124 bl[124] br[124] wl[396] vdd gnd cell_6t
Xbit_r397_c124 bl[124] br[124] wl[397] vdd gnd cell_6t
Xbit_r398_c124 bl[124] br[124] wl[398] vdd gnd cell_6t
Xbit_r399_c124 bl[124] br[124] wl[399] vdd gnd cell_6t
Xbit_r400_c124 bl[124] br[124] wl[400] vdd gnd cell_6t
Xbit_r401_c124 bl[124] br[124] wl[401] vdd gnd cell_6t
Xbit_r402_c124 bl[124] br[124] wl[402] vdd gnd cell_6t
Xbit_r403_c124 bl[124] br[124] wl[403] vdd gnd cell_6t
Xbit_r404_c124 bl[124] br[124] wl[404] vdd gnd cell_6t
Xbit_r405_c124 bl[124] br[124] wl[405] vdd gnd cell_6t
Xbit_r406_c124 bl[124] br[124] wl[406] vdd gnd cell_6t
Xbit_r407_c124 bl[124] br[124] wl[407] vdd gnd cell_6t
Xbit_r408_c124 bl[124] br[124] wl[408] vdd gnd cell_6t
Xbit_r409_c124 bl[124] br[124] wl[409] vdd gnd cell_6t
Xbit_r410_c124 bl[124] br[124] wl[410] vdd gnd cell_6t
Xbit_r411_c124 bl[124] br[124] wl[411] vdd gnd cell_6t
Xbit_r412_c124 bl[124] br[124] wl[412] vdd gnd cell_6t
Xbit_r413_c124 bl[124] br[124] wl[413] vdd gnd cell_6t
Xbit_r414_c124 bl[124] br[124] wl[414] vdd gnd cell_6t
Xbit_r415_c124 bl[124] br[124] wl[415] vdd gnd cell_6t
Xbit_r416_c124 bl[124] br[124] wl[416] vdd gnd cell_6t
Xbit_r417_c124 bl[124] br[124] wl[417] vdd gnd cell_6t
Xbit_r418_c124 bl[124] br[124] wl[418] vdd gnd cell_6t
Xbit_r419_c124 bl[124] br[124] wl[419] vdd gnd cell_6t
Xbit_r420_c124 bl[124] br[124] wl[420] vdd gnd cell_6t
Xbit_r421_c124 bl[124] br[124] wl[421] vdd gnd cell_6t
Xbit_r422_c124 bl[124] br[124] wl[422] vdd gnd cell_6t
Xbit_r423_c124 bl[124] br[124] wl[423] vdd gnd cell_6t
Xbit_r424_c124 bl[124] br[124] wl[424] vdd gnd cell_6t
Xbit_r425_c124 bl[124] br[124] wl[425] vdd gnd cell_6t
Xbit_r426_c124 bl[124] br[124] wl[426] vdd gnd cell_6t
Xbit_r427_c124 bl[124] br[124] wl[427] vdd gnd cell_6t
Xbit_r428_c124 bl[124] br[124] wl[428] vdd gnd cell_6t
Xbit_r429_c124 bl[124] br[124] wl[429] vdd gnd cell_6t
Xbit_r430_c124 bl[124] br[124] wl[430] vdd gnd cell_6t
Xbit_r431_c124 bl[124] br[124] wl[431] vdd gnd cell_6t
Xbit_r432_c124 bl[124] br[124] wl[432] vdd gnd cell_6t
Xbit_r433_c124 bl[124] br[124] wl[433] vdd gnd cell_6t
Xbit_r434_c124 bl[124] br[124] wl[434] vdd gnd cell_6t
Xbit_r435_c124 bl[124] br[124] wl[435] vdd gnd cell_6t
Xbit_r436_c124 bl[124] br[124] wl[436] vdd gnd cell_6t
Xbit_r437_c124 bl[124] br[124] wl[437] vdd gnd cell_6t
Xbit_r438_c124 bl[124] br[124] wl[438] vdd gnd cell_6t
Xbit_r439_c124 bl[124] br[124] wl[439] vdd gnd cell_6t
Xbit_r440_c124 bl[124] br[124] wl[440] vdd gnd cell_6t
Xbit_r441_c124 bl[124] br[124] wl[441] vdd gnd cell_6t
Xbit_r442_c124 bl[124] br[124] wl[442] vdd gnd cell_6t
Xbit_r443_c124 bl[124] br[124] wl[443] vdd gnd cell_6t
Xbit_r444_c124 bl[124] br[124] wl[444] vdd gnd cell_6t
Xbit_r445_c124 bl[124] br[124] wl[445] vdd gnd cell_6t
Xbit_r446_c124 bl[124] br[124] wl[446] vdd gnd cell_6t
Xbit_r447_c124 bl[124] br[124] wl[447] vdd gnd cell_6t
Xbit_r448_c124 bl[124] br[124] wl[448] vdd gnd cell_6t
Xbit_r449_c124 bl[124] br[124] wl[449] vdd gnd cell_6t
Xbit_r450_c124 bl[124] br[124] wl[450] vdd gnd cell_6t
Xbit_r451_c124 bl[124] br[124] wl[451] vdd gnd cell_6t
Xbit_r452_c124 bl[124] br[124] wl[452] vdd gnd cell_6t
Xbit_r453_c124 bl[124] br[124] wl[453] vdd gnd cell_6t
Xbit_r454_c124 bl[124] br[124] wl[454] vdd gnd cell_6t
Xbit_r455_c124 bl[124] br[124] wl[455] vdd gnd cell_6t
Xbit_r456_c124 bl[124] br[124] wl[456] vdd gnd cell_6t
Xbit_r457_c124 bl[124] br[124] wl[457] vdd gnd cell_6t
Xbit_r458_c124 bl[124] br[124] wl[458] vdd gnd cell_6t
Xbit_r459_c124 bl[124] br[124] wl[459] vdd gnd cell_6t
Xbit_r460_c124 bl[124] br[124] wl[460] vdd gnd cell_6t
Xbit_r461_c124 bl[124] br[124] wl[461] vdd gnd cell_6t
Xbit_r462_c124 bl[124] br[124] wl[462] vdd gnd cell_6t
Xbit_r463_c124 bl[124] br[124] wl[463] vdd gnd cell_6t
Xbit_r464_c124 bl[124] br[124] wl[464] vdd gnd cell_6t
Xbit_r465_c124 bl[124] br[124] wl[465] vdd gnd cell_6t
Xbit_r466_c124 bl[124] br[124] wl[466] vdd gnd cell_6t
Xbit_r467_c124 bl[124] br[124] wl[467] vdd gnd cell_6t
Xbit_r468_c124 bl[124] br[124] wl[468] vdd gnd cell_6t
Xbit_r469_c124 bl[124] br[124] wl[469] vdd gnd cell_6t
Xbit_r470_c124 bl[124] br[124] wl[470] vdd gnd cell_6t
Xbit_r471_c124 bl[124] br[124] wl[471] vdd gnd cell_6t
Xbit_r472_c124 bl[124] br[124] wl[472] vdd gnd cell_6t
Xbit_r473_c124 bl[124] br[124] wl[473] vdd gnd cell_6t
Xbit_r474_c124 bl[124] br[124] wl[474] vdd gnd cell_6t
Xbit_r475_c124 bl[124] br[124] wl[475] vdd gnd cell_6t
Xbit_r476_c124 bl[124] br[124] wl[476] vdd gnd cell_6t
Xbit_r477_c124 bl[124] br[124] wl[477] vdd gnd cell_6t
Xbit_r478_c124 bl[124] br[124] wl[478] vdd gnd cell_6t
Xbit_r479_c124 bl[124] br[124] wl[479] vdd gnd cell_6t
Xbit_r480_c124 bl[124] br[124] wl[480] vdd gnd cell_6t
Xbit_r481_c124 bl[124] br[124] wl[481] vdd gnd cell_6t
Xbit_r482_c124 bl[124] br[124] wl[482] vdd gnd cell_6t
Xbit_r483_c124 bl[124] br[124] wl[483] vdd gnd cell_6t
Xbit_r484_c124 bl[124] br[124] wl[484] vdd gnd cell_6t
Xbit_r485_c124 bl[124] br[124] wl[485] vdd gnd cell_6t
Xbit_r486_c124 bl[124] br[124] wl[486] vdd gnd cell_6t
Xbit_r487_c124 bl[124] br[124] wl[487] vdd gnd cell_6t
Xbit_r488_c124 bl[124] br[124] wl[488] vdd gnd cell_6t
Xbit_r489_c124 bl[124] br[124] wl[489] vdd gnd cell_6t
Xbit_r490_c124 bl[124] br[124] wl[490] vdd gnd cell_6t
Xbit_r491_c124 bl[124] br[124] wl[491] vdd gnd cell_6t
Xbit_r492_c124 bl[124] br[124] wl[492] vdd gnd cell_6t
Xbit_r493_c124 bl[124] br[124] wl[493] vdd gnd cell_6t
Xbit_r494_c124 bl[124] br[124] wl[494] vdd gnd cell_6t
Xbit_r495_c124 bl[124] br[124] wl[495] vdd gnd cell_6t
Xbit_r496_c124 bl[124] br[124] wl[496] vdd gnd cell_6t
Xbit_r497_c124 bl[124] br[124] wl[497] vdd gnd cell_6t
Xbit_r498_c124 bl[124] br[124] wl[498] vdd gnd cell_6t
Xbit_r499_c124 bl[124] br[124] wl[499] vdd gnd cell_6t
Xbit_r500_c124 bl[124] br[124] wl[500] vdd gnd cell_6t
Xbit_r501_c124 bl[124] br[124] wl[501] vdd gnd cell_6t
Xbit_r502_c124 bl[124] br[124] wl[502] vdd gnd cell_6t
Xbit_r503_c124 bl[124] br[124] wl[503] vdd gnd cell_6t
Xbit_r504_c124 bl[124] br[124] wl[504] vdd gnd cell_6t
Xbit_r505_c124 bl[124] br[124] wl[505] vdd gnd cell_6t
Xbit_r506_c124 bl[124] br[124] wl[506] vdd gnd cell_6t
Xbit_r507_c124 bl[124] br[124] wl[507] vdd gnd cell_6t
Xbit_r508_c124 bl[124] br[124] wl[508] vdd gnd cell_6t
Xbit_r509_c124 bl[124] br[124] wl[509] vdd gnd cell_6t
Xbit_r510_c124 bl[124] br[124] wl[510] vdd gnd cell_6t
Xbit_r511_c124 bl[124] br[124] wl[511] vdd gnd cell_6t
Xbit_r0_c125 bl[125] br[125] wl[0] vdd gnd cell_6t
Xbit_r1_c125 bl[125] br[125] wl[1] vdd gnd cell_6t
Xbit_r2_c125 bl[125] br[125] wl[2] vdd gnd cell_6t
Xbit_r3_c125 bl[125] br[125] wl[3] vdd gnd cell_6t
Xbit_r4_c125 bl[125] br[125] wl[4] vdd gnd cell_6t
Xbit_r5_c125 bl[125] br[125] wl[5] vdd gnd cell_6t
Xbit_r6_c125 bl[125] br[125] wl[6] vdd gnd cell_6t
Xbit_r7_c125 bl[125] br[125] wl[7] vdd gnd cell_6t
Xbit_r8_c125 bl[125] br[125] wl[8] vdd gnd cell_6t
Xbit_r9_c125 bl[125] br[125] wl[9] vdd gnd cell_6t
Xbit_r10_c125 bl[125] br[125] wl[10] vdd gnd cell_6t
Xbit_r11_c125 bl[125] br[125] wl[11] vdd gnd cell_6t
Xbit_r12_c125 bl[125] br[125] wl[12] vdd gnd cell_6t
Xbit_r13_c125 bl[125] br[125] wl[13] vdd gnd cell_6t
Xbit_r14_c125 bl[125] br[125] wl[14] vdd gnd cell_6t
Xbit_r15_c125 bl[125] br[125] wl[15] vdd gnd cell_6t
Xbit_r16_c125 bl[125] br[125] wl[16] vdd gnd cell_6t
Xbit_r17_c125 bl[125] br[125] wl[17] vdd gnd cell_6t
Xbit_r18_c125 bl[125] br[125] wl[18] vdd gnd cell_6t
Xbit_r19_c125 bl[125] br[125] wl[19] vdd gnd cell_6t
Xbit_r20_c125 bl[125] br[125] wl[20] vdd gnd cell_6t
Xbit_r21_c125 bl[125] br[125] wl[21] vdd gnd cell_6t
Xbit_r22_c125 bl[125] br[125] wl[22] vdd gnd cell_6t
Xbit_r23_c125 bl[125] br[125] wl[23] vdd gnd cell_6t
Xbit_r24_c125 bl[125] br[125] wl[24] vdd gnd cell_6t
Xbit_r25_c125 bl[125] br[125] wl[25] vdd gnd cell_6t
Xbit_r26_c125 bl[125] br[125] wl[26] vdd gnd cell_6t
Xbit_r27_c125 bl[125] br[125] wl[27] vdd gnd cell_6t
Xbit_r28_c125 bl[125] br[125] wl[28] vdd gnd cell_6t
Xbit_r29_c125 bl[125] br[125] wl[29] vdd gnd cell_6t
Xbit_r30_c125 bl[125] br[125] wl[30] vdd gnd cell_6t
Xbit_r31_c125 bl[125] br[125] wl[31] vdd gnd cell_6t
Xbit_r32_c125 bl[125] br[125] wl[32] vdd gnd cell_6t
Xbit_r33_c125 bl[125] br[125] wl[33] vdd gnd cell_6t
Xbit_r34_c125 bl[125] br[125] wl[34] vdd gnd cell_6t
Xbit_r35_c125 bl[125] br[125] wl[35] vdd gnd cell_6t
Xbit_r36_c125 bl[125] br[125] wl[36] vdd gnd cell_6t
Xbit_r37_c125 bl[125] br[125] wl[37] vdd gnd cell_6t
Xbit_r38_c125 bl[125] br[125] wl[38] vdd gnd cell_6t
Xbit_r39_c125 bl[125] br[125] wl[39] vdd gnd cell_6t
Xbit_r40_c125 bl[125] br[125] wl[40] vdd gnd cell_6t
Xbit_r41_c125 bl[125] br[125] wl[41] vdd gnd cell_6t
Xbit_r42_c125 bl[125] br[125] wl[42] vdd gnd cell_6t
Xbit_r43_c125 bl[125] br[125] wl[43] vdd gnd cell_6t
Xbit_r44_c125 bl[125] br[125] wl[44] vdd gnd cell_6t
Xbit_r45_c125 bl[125] br[125] wl[45] vdd gnd cell_6t
Xbit_r46_c125 bl[125] br[125] wl[46] vdd gnd cell_6t
Xbit_r47_c125 bl[125] br[125] wl[47] vdd gnd cell_6t
Xbit_r48_c125 bl[125] br[125] wl[48] vdd gnd cell_6t
Xbit_r49_c125 bl[125] br[125] wl[49] vdd gnd cell_6t
Xbit_r50_c125 bl[125] br[125] wl[50] vdd gnd cell_6t
Xbit_r51_c125 bl[125] br[125] wl[51] vdd gnd cell_6t
Xbit_r52_c125 bl[125] br[125] wl[52] vdd gnd cell_6t
Xbit_r53_c125 bl[125] br[125] wl[53] vdd gnd cell_6t
Xbit_r54_c125 bl[125] br[125] wl[54] vdd gnd cell_6t
Xbit_r55_c125 bl[125] br[125] wl[55] vdd gnd cell_6t
Xbit_r56_c125 bl[125] br[125] wl[56] vdd gnd cell_6t
Xbit_r57_c125 bl[125] br[125] wl[57] vdd gnd cell_6t
Xbit_r58_c125 bl[125] br[125] wl[58] vdd gnd cell_6t
Xbit_r59_c125 bl[125] br[125] wl[59] vdd gnd cell_6t
Xbit_r60_c125 bl[125] br[125] wl[60] vdd gnd cell_6t
Xbit_r61_c125 bl[125] br[125] wl[61] vdd gnd cell_6t
Xbit_r62_c125 bl[125] br[125] wl[62] vdd gnd cell_6t
Xbit_r63_c125 bl[125] br[125] wl[63] vdd gnd cell_6t
Xbit_r64_c125 bl[125] br[125] wl[64] vdd gnd cell_6t
Xbit_r65_c125 bl[125] br[125] wl[65] vdd gnd cell_6t
Xbit_r66_c125 bl[125] br[125] wl[66] vdd gnd cell_6t
Xbit_r67_c125 bl[125] br[125] wl[67] vdd gnd cell_6t
Xbit_r68_c125 bl[125] br[125] wl[68] vdd gnd cell_6t
Xbit_r69_c125 bl[125] br[125] wl[69] vdd gnd cell_6t
Xbit_r70_c125 bl[125] br[125] wl[70] vdd gnd cell_6t
Xbit_r71_c125 bl[125] br[125] wl[71] vdd gnd cell_6t
Xbit_r72_c125 bl[125] br[125] wl[72] vdd gnd cell_6t
Xbit_r73_c125 bl[125] br[125] wl[73] vdd gnd cell_6t
Xbit_r74_c125 bl[125] br[125] wl[74] vdd gnd cell_6t
Xbit_r75_c125 bl[125] br[125] wl[75] vdd gnd cell_6t
Xbit_r76_c125 bl[125] br[125] wl[76] vdd gnd cell_6t
Xbit_r77_c125 bl[125] br[125] wl[77] vdd gnd cell_6t
Xbit_r78_c125 bl[125] br[125] wl[78] vdd gnd cell_6t
Xbit_r79_c125 bl[125] br[125] wl[79] vdd gnd cell_6t
Xbit_r80_c125 bl[125] br[125] wl[80] vdd gnd cell_6t
Xbit_r81_c125 bl[125] br[125] wl[81] vdd gnd cell_6t
Xbit_r82_c125 bl[125] br[125] wl[82] vdd gnd cell_6t
Xbit_r83_c125 bl[125] br[125] wl[83] vdd gnd cell_6t
Xbit_r84_c125 bl[125] br[125] wl[84] vdd gnd cell_6t
Xbit_r85_c125 bl[125] br[125] wl[85] vdd gnd cell_6t
Xbit_r86_c125 bl[125] br[125] wl[86] vdd gnd cell_6t
Xbit_r87_c125 bl[125] br[125] wl[87] vdd gnd cell_6t
Xbit_r88_c125 bl[125] br[125] wl[88] vdd gnd cell_6t
Xbit_r89_c125 bl[125] br[125] wl[89] vdd gnd cell_6t
Xbit_r90_c125 bl[125] br[125] wl[90] vdd gnd cell_6t
Xbit_r91_c125 bl[125] br[125] wl[91] vdd gnd cell_6t
Xbit_r92_c125 bl[125] br[125] wl[92] vdd gnd cell_6t
Xbit_r93_c125 bl[125] br[125] wl[93] vdd gnd cell_6t
Xbit_r94_c125 bl[125] br[125] wl[94] vdd gnd cell_6t
Xbit_r95_c125 bl[125] br[125] wl[95] vdd gnd cell_6t
Xbit_r96_c125 bl[125] br[125] wl[96] vdd gnd cell_6t
Xbit_r97_c125 bl[125] br[125] wl[97] vdd gnd cell_6t
Xbit_r98_c125 bl[125] br[125] wl[98] vdd gnd cell_6t
Xbit_r99_c125 bl[125] br[125] wl[99] vdd gnd cell_6t
Xbit_r100_c125 bl[125] br[125] wl[100] vdd gnd cell_6t
Xbit_r101_c125 bl[125] br[125] wl[101] vdd gnd cell_6t
Xbit_r102_c125 bl[125] br[125] wl[102] vdd gnd cell_6t
Xbit_r103_c125 bl[125] br[125] wl[103] vdd gnd cell_6t
Xbit_r104_c125 bl[125] br[125] wl[104] vdd gnd cell_6t
Xbit_r105_c125 bl[125] br[125] wl[105] vdd gnd cell_6t
Xbit_r106_c125 bl[125] br[125] wl[106] vdd gnd cell_6t
Xbit_r107_c125 bl[125] br[125] wl[107] vdd gnd cell_6t
Xbit_r108_c125 bl[125] br[125] wl[108] vdd gnd cell_6t
Xbit_r109_c125 bl[125] br[125] wl[109] vdd gnd cell_6t
Xbit_r110_c125 bl[125] br[125] wl[110] vdd gnd cell_6t
Xbit_r111_c125 bl[125] br[125] wl[111] vdd gnd cell_6t
Xbit_r112_c125 bl[125] br[125] wl[112] vdd gnd cell_6t
Xbit_r113_c125 bl[125] br[125] wl[113] vdd gnd cell_6t
Xbit_r114_c125 bl[125] br[125] wl[114] vdd gnd cell_6t
Xbit_r115_c125 bl[125] br[125] wl[115] vdd gnd cell_6t
Xbit_r116_c125 bl[125] br[125] wl[116] vdd gnd cell_6t
Xbit_r117_c125 bl[125] br[125] wl[117] vdd gnd cell_6t
Xbit_r118_c125 bl[125] br[125] wl[118] vdd gnd cell_6t
Xbit_r119_c125 bl[125] br[125] wl[119] vdd gnd cell_6t
Xbit_r120_c125 bl[125] br[125] wl[120] vdd gnd cell_6t
Xbit_r121_c125 bl[125] br[125] wl[121] vdd gnd cell_6t
Xbit_r122_c125 bl[125] br[125] wl[122] vdd gnd cell_6t
Xbit_r123_c125 bl[125] br[125] wl[123] vdd gnd cell_6t
Xbit_r124_c125 bl[125] br[125] wl[124] vdd gnd cell_6t
Xbit_r125_c125 bl[125] br[125] wl[125] vdd gnd cell_6t
Xbit_r126_c125 bl[125] br[125] wl[126] vdd gnd cell_6t
Xbit_r127_c125 bl[125] br[125] wl[127] vdd gnd cell_6t
Xbit_r128_c125 bl[125] br[125] wl[128] vdd gnd cell_6t
Xbit_r129_c125 bl[125] br[125] wl[129] vdd gnd cell_6t
Xbit_r130_c125 bl[125] br[125] wl[130] vdd gnd cell_6t
Xbit_r131_c125 bl[125] br[125] wl[131] vdd gnd cell_6t
Xbit_r132_c125 bl[125] br[125] wl[132] vdd gnd cell_6t
Xbit_r133_c125 bl[125] br[125] wl[133] vdd gnd cell_6t
Xbit_r134_c125 bl[125] br[125] wl[134] vdd gnd cell_6t
Xbit_r135_c125 bl[125] br[125] wl[135] vdd gnd cell_6t
Xbit_r136_c125 bl[125] br[125] wl[136] vdd gnd cell_6t
Xbit_r137_c125 bl[125] br[125] wl[137] vdd gnd cell_6t
Xbit_r138_c125 bl[125] br[125] wl[138] vdd gnd cell_6t
Xbit_r139_c125 bl[125] br[125] wl[139] vdd gnd cell_6t
Xbit_r140_c125 bl[125] br[125] wl[140] vdd gnd cell_6t
Xbit_r141_c125 bl[125] br[125] wl[141] vdd gnd cell_6t
Xbit_r142_c125 bl[125] br[125] wl[142] vdd gnd cell_6t
Xbit_r143_c125 bl[125] br[125] wl[143] vdd gnd cell_6t
Xbit_r144_c125 bl[125] br[125] wl[144] vdd gnd cell_6t
Xbit_r145_c125 bl[125] br[125] wl[145] vdd gnd cell_6t
Xbit_r146_c125 bl[125] br[125] wl[146] vdd gnd cell_6t
Xbit_r147_c125 bl[125] br[125] wl[147] vdd gnd cell_6t
Xbit_r148_c125 bl[125] br[125] wl[148] vdd gnd cell_6t
Xbit_r149_c125 bl[125] br[125] wl[149] vdd gnd cell_6t
Xbit_r150_c125 bl[125] br[125] wl[150] vdd gnd cell_6t
Xbit_r151_c125 bl[125] br[125] wl[151] vdd gnd cell_6t
Xbit_r152_c125 bl[125] br[125] wl[152] vdd gnd cell_6t
Xbit_r153_c125 bl[125] br[125] wl[153] vdd gnd cell_6t
Xbit_r154_c125 bl[125] br[125] wl[154] vdd gnd cell_6t
Xbit_r155_c125 bl[125] br[125] wl[155] vdd gnd cell_6t
Xbit_r156_c125 bl[125] br[125] wl[156] vdd gnd cell_6t
Xbit_r157_c125 bl[125] br[125] wl[157] vdd gnd cell_6t
Xbit_r158_c125 bl[125] br[125] wl[158] vdd gnd cell_6t
Xbit_r159_c125 bl[125] br[125] wl[159] vdd gnd cell_6t
Xbit_r160_c125 bl[125] br[125] wl[160] vdd gnd cell_6t
Xbit_r161_c125 bl[125] br[125] wl[161] vdd gnd cell_6t
Xbit_r162_c125 bl[125] br[125] wl[162] vdd gnd cell_6t
Xbit_r163_c125 bl[125] br[125] wl[163] vdd gnd cell_6t
Xbit_r164_c125 bl[125] br[125] wl[164] vdd gnd cell_6t
Xbit_r165_c125 bl[125] br[125] wl[165] vdd gnd cell_6t
Xbit_r166_c125 bl[125] br[125] wl[166] vdd gnd cell_6t
Xbit_r167_c125 bl[125] br[125] wl[167] vdd gnd cell_6t
Xbit_r168_c125 bl[125] br[125] wl[168] vdd gnd cell_6t
Xbit_r169_c125 bl[125] br[125] wl[169] vdd gnd cell_6t
Xbit_r170_c125 bl[125] br[125] wl[170] vdd gnd cell_6t
Xbit_r171_c125 bl[125] br[125] wl[171] vdd gnd cell_6t
Xbit_r172_c125 bl[125] br[125] wl[172] vdd gnd cell_6t
Xbit_r173_c125 bl[125] br[125] wl[173] vdd gnd cell_6t
Xbit_r174_c125 bl[125] br[125] wl[174] vdd gnd cell_6t
Xbit_r175_c125 bl[125] br[125] wl[175] vdd gnd cell_6t
Xbit_r176_c125 bl[125] br[125] wl[176] vdd gnd cell_6t
Xbit_r177_c125 bl[125] br[125] wl[177] vdd gnd cell_6t
Xbit_r178_c125 bl[125] br[125] wl[178] vdd gnd cell_6t
Xbit_r179_c125 bl[125] br[125] wl[179] vdd gnd cell_6t
Xbit_r180_c125 bl[125] br[125] wl[180] vdd gnd cell_6t
Xbit_r181_c125 bl[125] br[125] wl[181] vdd gnd cell_6t
Xbit_r182_c125 bl[125] br[125] wl[182] vdd gnd cell_6t
Xbit_r183_c125 bl[125] br[125] wl[183] vdd gnd cell_6t
Xbit_r184_c125 bl[125] br[125] wl[184] vdd gnd cell_6t
Xbit_r185_c125 bl[125] br[125] wl[185] vdd gnd cell_6t
Xbit_r186_c125 bl[125] br[125] wl[186] vdd gnd cell_6t
Xbit_r187_c125 bl[125] br[125] wl[187] vdd gnd cell_6t
Xbit_r188_c125 bl[125] br[125] wl[188] vdd gnd cell_6t
Xbit_r189_c125 bl[125] br[125] wl[189] vdd gnd cell_6t
Xbit_r190_c125 bl[125] br[125] wl[190] vdd gnd cell_6t
Xbit_r191_c125 bl[125] br[125] wl[191] vdd gnd cell_6t
Xbit_r192_c125 bl[125] br[125] wl[192] vdd gnd cell_6t
Xbit_r193_c125 bl[125] br[125] wl[193] vdd gnd cell_6t
Xbit_r194_c125 bl[125] br[125] wl[194] vdd gnd cell_6t
Xbit_r195_c125 bl[125] br[125] wl[195] vdd gnd cell_6t
Xbit_r196_c125 bl[125] br[125] wl[196] vdd gnd cell_6t
Xbit_r197_c125 bl[125] br[125] wl[197] vdd gnd cell_6t
Xbit_r198_c125 bl[125] br[125] wl[198] vdd gnd cell_6t
Xbit_r199_c125 bl[125] br[125] wl[199] vdd gnd cell_6t
Xbit_r200_c125 bl[125] br[125] wl[200] vdd gnd cell_6t
Xbit_r201_c125 bl[125] br[125] wl[201] vdd gnd cell_6t
Xbit_r202_c125 bl[125] br[125] wl[202] vdd gnd cell_6t
Xbit_r203_c125 bl[125] br[125] wl[203] vdd gnd cell_6t
Xbit_r204_c125 bl[125] br[125] wl[204] vdd gnd cell_6t
Xbit_r205_c125 bl[125] br[125] wl[205] vdd gnd cell_6t
Xbit_r206_c125 bl[125] br[125] wl[206] vdd gnd cell_6t
Xbit_r207_c125 bl[125] br[125] wl[207] vdd gnd cell_6t
Xbit_r208_c125 bl[125] br[125] wl[208] vdd gnd cell_6t
Xbit_r209_c125 bl[125] br[125] wl[209] vdd gnd cell_6t
Xbit_r210_c125 bl[125] br[125] wl[210] vdd gnd cell_6t
Xbit_r211_c125 bl[125] br[125] wl[211] vdd gnd cell_6t
Xbit_r212_c125 bl[125] br[125] wl[212] vdd gnd cell_6t
Xbit_r213_c125 bl[125] br[125] wl[213] vdd gnd cell_6t
Xbit_r214_c125 bl[125] br[125] wl[214] vdd gnd cell_6t
Xbit_r215_c125 bl[125] br[125] wl[215] vdd gnd cell_6t
Xbit_r216_c125 bl[125] br[125] wl[216] vdd gnd cell_6t
Xbit_r217_c125 bl[125] br[125] wl[217] vdd gnd cell_6t
Xbit_r218_c125 bl[125] br[125] wl[218] vdd gnd cell_6t
Xbit_r219_c125 bl[125] br[125] wl[219] vdd gnd cell_6t
Xbit_r220_c125 bl[125] br[125] wl[220] vdd gnd cell_6t
Xbit_r221_c125 bl[125] br[125] wl[221] vdd gnd cell_6t
Xbit_r222_c125 bl[125] br[125] wl[222] vdd gnd cell_6t
Xbit_r223_c125 bl[125] br[125] wl[223] vdd gnd cell_6t
Xbit_r224_c125 bl[125] br[125] wl[224] vdd gnd cell_6t
Xbit_r225_c125 bl[125] br[125] wl[225] vdd gnd cell_6t
Xbit_r226_c125 bl[125] br[125] wl[226] vdd gnd cell_6t
Xbit_r227_c125 bl[125] br[125] wl[227] vdd gnd cell_6t
Xbit_r228_c125 bl[125] br[125] wl[228] vdd gnd cell_6t
Xbit_r229_c125 bl[125] br[125] wl[229] vdd gnd cell_6t
Xbit_r230_c125 bl[125] br[125] wl[230] vdd gnd cell_6t
Xbit_r231_c125 bl[125] br[125] wl[231] vdd gnd cell_6t
Xbit_r232_c125 bl[125] br[125] wl[232] vdd gnd cell_6t
Xbit_r233_c125 bl[125] br[125] wl[233] vdd gnd cell_6t
Xbit_r234_c125 bl[125] br[125] wl[234] vdd gnd cell_6t
Xbit_r235_c125 bl[125] br[125] wl[235] vdd gnd cell_6t
Xbit_r236_c125 bl[125] br[125] wl[236] vdd gnd cell_6t
Xbit_r237_c125 bl[125] br[125] wl[237] vdd gnd cell_6t
Xbit_r238_c125 bl[125] br[125] wl[238] vdd gnd cell_6t
Xbit_r239_c125 bl[125] br[125] wl[239] vdd gnd cell_6t
Xbit_r240_c125 bl[125] br[125] wl[240] vdd gnd cell_6t
Xbit_r241_c125 bl[125] br[125] wl[241] vdd gnd cell_6t
Xbit_r242_c125 bl[125] br[125] wl[242] vdd gnd cell_6t
Xbit_r243_c125 bl[125] br[125] wl[243] vdd gnd cell_6t
Xbit_r244_c125 bl[125] br[125] wl[244] vdd gnd cell_6t
Xbit_r245_c125 bl[125] br[125] wl[245] vdd gnd cell_6t
Xbit_r246_c125 bl[125] br[125] wl[246] vdd gnd cell_6t
Xbit_r247_c125 bl[125] br[125] wl[247] vdd gnd cell_6t
Xbit_r248_c125 bl[125] br[125] wl[248] vdd gnd cell_6t
Xbit_r249_c125 bl[125] br[125] wl[249] vdd gnd cell_6t
Xbit_r250_c125 bl[125] br[125] wl[250] vdd gnd cell_6t
Xbit_r251_c125 bl[125] br[125] wl[251] vdd gnd cell_6t
Xbit_r252_c125 bl[125] br[125] wl[252] vdd gnd cell_6t
Xbit_r253_c125 bl[125] br[125] wl[253] vdd gnd cell_6t
Xbit_r254_c125 bl[125] br[125] wl[254] vdd gnd cell_6t
Xbit_r255_c125 bl[125] br[125] wl[255] vdd gnd cell_6t
Xbit_r256_c125 bl[125] br[125] wl[256] vdd gnd cell_6t
Xbit_r257_c125 bl[125] br[125] wl[257] vdd gnd cell_6t
Xbit_r258_c125 bl[125] br[125] wl[258] vdd gnd cell_6t
Xbit_r259_c125 bl[125] br[125] wl[259] vdd gnd cell_6t
Xbit_r260_c125 bl[125] br[125] wl[260] vdd gnd cell_6t
Xbit_r261_c125 bl[125] br[125] wl[261] vdd gnd cell_6t
Xbit_r262_c125 bl[125] br[125] wl[262] vdd gnd cell_6t
Xbit_r263_c125 bl[125] br[125] wl[263] vdd gnd cell_6t
Xbit_r264_c125 bl[125] br[125] wl[264] vdd gnd cell_6t
Xbit_r265_c125 bl[125] br[125] wl[265] vdd gnd cell_6t
Xbit_r266_c125 bl[125] br[125] wl[266] vdd gnd cell_6t
Xbit_r267_c125 bl[125] br[125] wl[267] vdd gnd cell_6t
Xbit_r268_c125 bl[125] br[125] wl[268] vdd gnd cell_6t
Xbit_r269_c125 bl[125] br[125] wl[269] vdd gnd cell_6t
Xbit_r270_c125 bl[125] br[125] wl[270] vdd gnd cell_6t
Xbit_r271_c125 bl[125] br[125] wl[271] vdd gnd cell_6t
Xbit_r272_c125 bl[125] br[125] wl[272] vdd gnd cell_6t
Xbit_r273_c125 bl[125] br[125] wl[273] vdd gnd cell_6t
Xbit_r274_c125 bl[125] br[125] wl[274] vdd gnd cell_6t
Xbit_r275_c125 bl[125] br[125] wl[275] vdd gnd cell_6t
Xbit_r276_c125 bl[125] br[125] wl[276] vdd gnd cell_6t
Xbit_r277_c125 bl[125] br[125] wl[277] vdd gnd cell_6t
Xbit_r278_c125 bl[125] br[125] wl[278] vdd gnd cell_6t
Xbit_r279_c125 bl[125] br[125] wl[279] vdd gnd cell_6t
Xbit_r280_c125 bl[125] br[125] wl[280] vdd gnd cell_6t
Xbit_r281_c125 bl[125] br[125] wl[281] vdd gnd cell_6t
Xbit_r282_c125 bl[125] br[125] wl[282] vdd gnd cell_6t
Xbit_r283_c125 bl[125] br[125] wl[283] vdd gnd cell_6t
Xbit_r284_c125 bl[125] br[125] wl[284] vdd gnd cell_6t
Xbit_r285_c125 bl[125] br[125] wl[285] vdd gnd cell_6t
Xbit_r286_c125 bl[125] br[125] wl[286] vdd gnd cell_6t
Xbit_r287_c125 bl[125] br[125] wl[287] vdd gnd cell_6t
Xbit_r288_c125 bl[125] br[125] wl[288] vdd gnd cell_6t
Xbit_r289_c125 bl[125] br[125] wl[289] vdd gnd cell_6t
Xbit_r290_c125 bl[125] br[125] wl[290] vdd gnd cell_6t
Xbit_r291_c125 bl[125] br[125] wl[291] vdd gnd cell_6t
Xbit_r292_c125 bl[125] br[125] wl[292] vdd gnd cell_6t
Xbit_r293_c125 bl[125] br[125] wl[293] vdd gnd cell_6t
Xbit_r294_c125 bl[125] br[125] wl[294] vdd gnd cell_6t
Xbit_r295_c125 bl[125] br[125] wl[295] vdd gnd cell_6t
Xbit_r296_c125 bl[125] br[125] wl[296] vdd gnd cell_6t
Xbit_r297_c125 bl[125] br[125] wl[297] vdd gnd cell_6t
Xbit_r298_c125 bl[125] br[125] wl[298] vdd gnd cell_6t
Xbit_r299_c125 bl[125] br[125] wl[299] vdd gnd cell_6t
Xbit_r300_c125 bl[125] br[125] wl[300] vdd gnd cell_6t
Xbit_r301_c125 bl[125] br[125] wl[301] vdd gnd cell_6t
Xbit_r302_c125 bl[125] br[125] wl[302] vdd gnd cell_6t
Xbit_r303_c125 bl[125] br[125] wl[303] vdd gnd cell_6t
Xbit_r304_c125 bl[125] br[125] wl[304] vdd gnd cell_6t
Xbit_r305_c125 bl[125] br[125] wl[305] vdd gnd cell_6t
Xbit_r306_c125 bl[125] br[125] wl[306] vdd gnd cell_6t
Xbit_r307_c125 bl[125] br[125] wl[307] vdd gnd cell_6t
Xbit_r308_c125 bl[125] br[125] wl[308] vdd gnd cell_6t
Xbit_r309_c125 bl[125] br[125] wl[309] vdd gnd cell_6t
Xbit_r310_c125 bl[125] br[125] wl[310] vdd gnd cell_6t
Xbit_r311_c125 bl[125] br[125] wl[311] vdd gnd cell_6t
Xbit_r312_c125 bl[125] br[125] wl[312] vdd gnd cell_6t
Xbit_r313_c125 bl[125] br[125] wl[313] vdd gnd cell_6t
Xbit_r314_c125 bl[125] br[125] wl[314] vdd gnd cell_6t
Xbit_r315_c125 bl[125] br[125] wl[315] vdd gnd cell_6t
Xbit_r316_c125 bl[125] br[125] wl[316] vdd gnd cell_6t
Xbit_r317_c125 bl[125] br[125] wl[317] vdd gnd cell_6t
Xbit_r318_c125 bl[125] br[125] wl[318] vdd gnd cell_6t
Xbit_r319_c125 bl[125] br[125] wl[319] vdd gnd cell_6t
Xbit_r320_c125 bl[125] br[125] wl[320] vdd gnd cell_6t
Xbit_r321_c125 bl[125] br[125] wl[321] vdd gnd cell_6t
Xbit_r322_c125 bl[125] br[125] wl[322] vdd gnd cell_6t
Xbit_r323_c125 bl[125] br[125] wl[323] vdd gnd cell_6t
Xbit_r324_c125 bl[125] br[125] wl[324] vdd gnd cell_6t
Xbit_r325_c125 bl[125] br[125] wl[325] vdd gnd cell_6t
Xbit_r326_c125 bl[125] br[125] wl[326] vdd gnd cell_6t
Xbit_r327_c125 bl[125] br[125] wl[327] vdd gnd cell_6t
Xbit_r328_c125 bl[125] br[125] wl[328] vdd gnd cell_6t
Xbit_r329_c125 bl[125] br[125] wl[329] vdd gnd cell_6t
Xbit_r330_c125 bl[125] br[125] wl[330] vdd gnd cell_6t
Xbit_r331_c125 bl[125] br[125] wl[331] vdd gnd cell_6t
Xbit_r332_c125 bl[125] br[125] wl[332] vdd gnd cell_6t
Xbit_r333_c125 bl[125] br[125] wl[333] vdd gnd cell_6t
Xbit_r334_c125 bl[125] br[125] wl[334] vdd gnd cell_6t
Xbit_r335_c125 bl[125] br[125] wl[335] vdd gnd cell_6t
Xbit_r336_c125 bl[125] br[125] wl[336] vdd gnd cell_6t
Xbit_r337_c125 bl[125] br[125] wl[337] vdd gnd cell_6t
Xbit_r338_c125 bl[125] br[125] wl[338] vdd gnd cell_6t
Xbit_r339_c125 bl[125] br[125] wl[339] vdd gnd cell_6t
Xbit_r340_c125 bl[125] br[125] wl[340] vdd gnd cell_6t
Xbit_r341_c125 bl[125] br[125] wl[341] vdd gnd cell_6t
Xbit_r342_c125 bl[125] br[125] wl[342] vdd gnd cell_6t
Xbit_r343_c125 bl[125] br[125] wl[343] vdd gnd cell_6t
Xbit_r344_c125 bl[125] br[125] wl[344] vdd gnd cell_6t
Xbit_r345_c125 bl[125] br[125] wl[345] vdd gnd cell_6t
Xbit_r346_c125 bl[125] br[125] wl[346] vdd gnd cell_6t
Xbit_r347_c125 bl[125] br[125] wl[347] vdd gnd cell_6t
Xbit_r348_c125 bl[125] br[125] wl[348] vdd gnd cell_6t
Xbit_r349_c125 bl[125] br[125] wl[349] vdd gnd cell_6t
Xbit_r350_c125 bl[125] br[125] wl[350] vdd gnd cell_6t
Xbit_r351_c125 bl[125] br[125] wl[351] vdd gnd cell_6t
Xbit_r352_c125 bl[125] br[125] wl[352] vdd gnd cell_6t
Xbit_r353_c125 bl[125] br[125] wl[353] vdd gnd cell_6t
Xbit_r354_c125 bl[125] br[125] wl[354] vdd gnd cell_6t
Xbit_r355_c125 bl[125] br[125] wl[355] vdd gnd cell_6t
Xbit_r356_c125 bl[125] br[125] wl[356] vdd gnd cell_6t
Xbit_r357_c125 bl[125] br[125] wl[357] vdd gnd cell_6t
Xbit_r358_c125 bl[125] br[125] wl[358] vdd gnd cell_6t
Xbit_r359_c125 bl[125] br[125] wl[359] vdd gnd cell_6t
Xbit_r360_c125 bl[125] br[125] wl[360] vdd gnd cell_6t
Xbit_r361_c125 bl[125] br[125] wl[361] vdd gnd cell_6t
Xbit_r362_c125 bl[125] br[125] wl[362] vdd gnd cell_6t
Xbit_r363_c125 bl[125] br[125] wl[363] vdd gnd cell_6t
Xbit_r364_c125 bl[125] br[125] wl[364] vdd gnd cell_6t
Xbit_r365_c125 bl[125] br[125] wl[365] vdd gnd cell_6t
Xbit_r366_c125 bl[125] br[125] wl[366] vdd gnd cell_6t
Xbit_r367_c125 bl[125] br[125] wl[367] vdd gnd cell_6t
Xbit_r368_c125 bl[125] br[125] wl[368] vdd gnd cell_6t
Xbit_r369_c125 bl[125] br[125] wl[369] vdd gnd cell_6t
Xbit_r370_c125 bl[125] br[125] wl[370] vdd gnd cell_6t
Xbit_r371_c125 bl[125] br[125] wl[371] vdd gnd cell_6t
Xbit_r372_c125 bl[125] br[125] wl[372] vdd gnd cell_6t
Xbit_r373_c125 bl[125] br[125] wl[373] vdd gnd cell_6t
Xbit_r374_c125 bl[125] br[125] wl[374] vdd gnd cell_6t
Xbit_r375_c125 bl[125] br[125] wl[375] vdd gnd cell_6t
Xbit_r376_c125 bl[125] br[125] wl[376] vdd gnd cell_6t
Xbit_r377_c125 bl[125] br[125] wl[377] vdd gnd cell_6t
Xbit_r378_c125 bl[125] br[125] wl[378] vdd gnd cell_6t
Xbit_r379_c125 bl[125] br[125] wl[379] vdd gnd cell_6t
Xbit_r380_c125 bl[125] br[125] wl[380] vdd gnd cell_6t
Xbit_r381_c125 bl[125] br[125] wl[381] vdd gnd cell_6t
Xbit_r382_c125 bl[125] br[125] wl[382] vdd gnd cell_6t
Xbit_r383_c125 bl[125] br[125] wl[383] vdd gnd cell_6t
Xbit_r384_c125 bl[125] br[125] wl[384] vdd gnd cell_6t
Xbit_r385_c125 bl[125] br[125] wl[385] vdd gnd cell_6t
Xbit_r386_c125 bl[125] br[125] wl[386] vdd gnd cell_6t
Xbit_r387_c125 bl[125] br[125] wl[387] vdd gnd cell_6t
Xbit_r388_c125 bl[125] br[125] wl[388] vdd gnd cell_6t
Xbit_r389_c125 bl[125] br[125] wl[389] vdd gnd cell_6t
Xbit_r390_c125 bl[125] br[125] wl[390] vdd gnd cell_6t
Xbit_r391_c125 bl[125] br[125] wl[391] vdd gnd cell_6t
Xbit_r392_c125 bl[125] br[125] wl[392] vdd gnd cell_6t
Xbit_r393_c125 bl[125] br[125] wl[393] vdd gnd cell_6t
Xbit_r394_c125 bl[125] br[125] wl[394] vdd gnd cell_6t
Xbit_r395_c125 bl[125] br[125] wl[395] vdd gnd cell_6t
Xbit_r396_c125 bl[125] br[125] wl[396] vdd gnd cell_6t
Xbit_r397_c125 bl[125] br[125] wl[397] vdd gnd cell_6t
Xbit_r398_c125 bl[125] br[125] wl[398] vdd gnd cell_6t
Xbit_r399_c125 bl[125] br[125] wl[399] vdd gnd cell_6t
Xbit_r400_c125 bl[125] br[125] wl[400] vdd gnd cell_6t
Xbit_r401_c125 bl[125] br[125] wl[401] vdd gnd cell_6t
Xbit_r402_c125 bl[125] br[125] wl[402] vdd gnd cell_6t
Xbit_r403_c125 bl[125] br[125] wl[403] vdd gnd cell_6t
Xbit_r404_c125 bl[125] br[125] wl[404] vdd gnd cell_6t
Xbit_r405_c125 bl[125] br[125] wl[405] vdd gnd cell_6t
Xbit_r406_c125 bl[125] br[125] wl[406] vdd gnd cell_6t
Xbit_r407_c125 bl[125] br[125] wl[407] vdd gnd cell_6t
Xbit_r408_c125 bl[125] br[125] wl[408] vdd gnd cell_6t
Xbit_r409_c125 bl[125] br[125] wl[409] vdd gnd cell_6t
Xbit_r410_c125 bl[125] br[125] wl[410] vdd gnd cell_6t
Xbit_r411_c125 bl[125] br[125] wl[411] vdd gnd cell_6t
Xbit_r412_c125 bl[125] br[125] wl[412] vdd gnd cell_6t
Xbit_r413_c125 bl[125] br[125] wl[413] vdd gnd cell_6t
Xbit_r414_c125 bl[125] br[125] wl[414] vdd gnd cell_6t
Xbit_r415_c125 bl[125] br[125] wl[415] vdd gnd cell_6t
Xbit_r416_c125 bl[125] br[125] wl[416] vdd gnd cell_6t
Xbit_r417_c125 bl[125] br[125] wl[417] vdd gnd cell_6t
Xbit_r418_c125 bl[125] br[125] wl[418] vdd gnd cell_6t
Xbit_r419_c125 bl[125] br[125] wl[419] vdd gnd cell_6t
Xbit_r420_c125 bl[125] br[125] wl[420] vdd gnd cell_6t
Xbit_r421_c125 bl[125] br[125] wl[421] vdd gnd cell_6t
Xbit_r422_c125 bl[125] br[125] wl[422] vdd gnd cell_6t
Xbit_r423_c125 bl[125] br[125] wl[423] vdd gnd cell_6t
Xbit_r424_c125 bl[125] br[125] wl[424] vdd gnd cell_6t
Xbit_r425_c125 bl[125] br[125] wl[425] vdd gnd cell_6t
Xbit_r426_c125 bl[125] br[125] wl[426] vdd gnd cell_6t
Xbit_r427_c125 bl[125] br[125] wl[427] vdd gnd cell_6t
Xbit_r428_c125 bl[125] br[125] wl[428] vdd gnd cell_6t
Xbit_r429_c125 bl[125] br[125] wl[429] vdd gnd cell_6t
Xbit_r430_c125 bl[125] br[125] wl[430] vdd gnd cell_6t
Xbit_r431_c125 bl[125] br[125] wl[431] vdd gnd cell_6t
Xbit_r432_c125 bl[125] br[125] wl[432] vdd gnd cell_6t
Xbit_r433_c125 bl[125] br[125] wl[433] vdd gnd cell_6t
Xbit_r434_c125 bl[125] br[125] wl[434] vdd gnd cell_6t
Xbit_r435_c125 bl[125] br[125] wl[435] vdd gnd cell_6t
Xbit_r436_c125 bl[125] br[125] wl[436] vdd gnd cell_6t
Xbit_r437_c125 bl[125] br[125] wl[437] vdd gnd cell_6t
Xbit_r438_c125 bl[125] br[125] wl[438] vdd gnd cell_6t
Xbit_r439_c125 bl[125] br[125] wl[439] vdd gnd cell_6t
Xbit_r440_c125 bl[125] br[125] wl[440] vdd gnd cell_6t
Xbit_r441_c125 bl[125] br[125] wl[441] vdd gnd cell_6t
Xbit_r442_c125 bl[125] br[125] wl[442] vdd gnd cell_6t
Xbit_r443_c125 bl[125] br[125] wl[443] vdd gnd cell_6t
Xbit_r444_c125 bl[125] br[125] wl[444] vdd gnd cell_6t
Xbit_r445_c125 bl[125] br[125] wl[445] vdd gnd cell_6t
Xbit_r446_c125 bl[125] br[125] wl[446] vdd gnd cell_6t
Xbit_r447_c125 bl[125] br[125] wl[447] vdd gnd cell_6t
Xbit_r448_c125 bl[125] br[125] wl[448] vdd gnd cell_6t
Xbit_r449_c125 bl[125] br[125] wl[449] vdd gnd cell_6t
Xbit_r450_c125 bl[125] br[125] wl[450] vdd gnd cell_6t
Xbit_r451_c125 bl[125] br[125] wl[451] vdd gnd cell_6t
Xbit_r452_c125 bl[125] br[125] wl[452] vdd gnd cell_6t
Xbit_r453_c125 bl[125] br[125] wl[453] vdd gnd cell_6t
Xbit_r454_c125 bl[125] br[125] wl[454] vdd gnd cell_6t
Xbit_r455_c125 bl[125] br[125] wl[455] vdd gnd cell_6t
Xbit_r456_c125 bl[125] br[125] wl[456] vdd gnd cell_6t
Xbit_r457_c125 bl[125] br[125] wl[457] vdd gnd cell_6t
Xbit_r458_c125 bl[125] br[125] wl[458] vdd gnd cell_6t
Xbit_r459_c125 bl[125] br[125] wl[459] vdd gnd cell_6t
Xbit_r460_c125 bl[125] br[125] wl[460] vdd gnd cell_6t
Xbit_r461_c125 bl[125] br[125] wl[461] vdd gnd cell_6t
Xbit_r462_c125 bl[125] br[125] wl[462] vdd gnd cell_6t
Xbit_r463_c125 bl[125] br[125] wl[463] vdd gnd cell_6t
Xbit_r464_c125 bl[125] br[125] wl[464] vdd gnd cell_6t
Xbit_r465_c125 bl[125] br[125] wl[465] vdd gnd cell_6t
Xbit_r466_c125 bl[125] br[125] wl[466] vdd gnd cell_6t
Xbit_r467_c125 bl[125] br[125] wl[467] vdd gnd cell_6t
Xbit_r468_c125 bl[125] br[125] wl[468] vdd gnd cell_6t
Xbit_r469_c125 bl[125] br[125] wl[469] vdd gnd cell_6t
Xbit_r470_c125 bl[125] br[125] wl[470] vdd gnd cell_6t
Xbit_r471_c125 bl[125] br[125] wl[471] vdd gnd cell_6t
Xbit_r472_c125 bl[125] br[125] wl[472] vdd gnd cell_6t
Xbit_r473_c125 bl[125] br[125] wl[473] vdd gnd cell_6t
Xbit_r474_c125 bl[125] br[125] wl[474] vdd gnd cell_6t
Xbit_r475_c125 bl[125] br[125] wl[475] vdd gnd cell_6t
Xbit_r476_c125 bl[125] br[125] wl[476] vdd gnd cell_6t
Xbit_r477_c125 bl[125] br[125] wl[477] vdd gnd cell_6t
Xbit_r478_c125 bl[125] br[125] wl[478] vdd gnd cell_6t
Xbit_r479_c125 bl[125] br[125] wl[479] vdd gnd cell_6t
Xbit_r480_c125 bl[125] br[125] wl[480] vdd gnd cell_6t
Xbit_r481_c125 bl[125] br[125] wl[481] vdd gnd cell_6t
Xbit_r482_c125 bl[125] br[125] wl[482] vdd gnd cell_6t
Xbit_r483_c125 bl[125] br[125] wl[483] vdd gnd cell_6t
Xbit_r484_c125 bl[125] br[125] wl[484] vdd gnd cell_6t
Xbit_r485_c125 bl[125] br[125] wl[485] vdd gnd cell_6t
Xbit_r486_c125 bl[125] br[125] wl[486] vdd gnd cell_6t
Xbit_r487_c125 bl[125] br[125] wl[487] vdd gnd cell_6t
Xbit_r488_c125 bl[125] br[125] wl[488] vdd gnd cell_6t
Xbit_r489_c125 bl[125] br[125] wl[489] vdd gnd cell_6t
Xbit_r490_c125 bl[125] br[125] wl[490] vdd gnd cell_6t
Xbit_r491_c125 bl[125] br[125] wl[491] vdd gnd cell_6t
Xbit_r492_c125 bl[125] br[125] wl[492] vdd gnd cell_6t
Xbit_r493_c125 bl[125] br[125] wl[493] vdd gnd cell_6t
Xbit_r494_c125 bl[125] br[125] wl[494] vdd gnd cell_6t
Xbit_r495_c125 bl[125] br[125] wl[495] vdd gnd cell_6t
Xbit_r496_c125 bl[125] br[125] wl[496] vdd gnd cell_6t
Xbit_r497_c125 bl[125] br[125] wl[497] vdd gnd cell_6t
Xbit_r498_c125 bl[125] br[125] wl[498] vdd gnd cell_6t
Xbit_r499_c125 bl[125] br[125] wl[499] vdd gnd cell_6t
Xbit_r500_c125 bl[125] br[125] wl[500] vdd gnd cell_6t
Xbit_r501_c125 bl[125] br[125] wl[501] vdd gnd cell_6t
Xbit_r502_c125 bl[125] br[125] wl[502] vdd gnd cell_6t
Xbit_r503_c125 bl[125] br[125] wl[503] vdd gnd cell_6t
Xbit_r504_c125 bl[125] br[125] wl[504] vdd gnd cell_6t
Xbit_r505_c125 bl[125] br[125] wl[505] vdd gnd cell_6t
Xbit_r506_c125 bl[125] br[125] wl[506] vdd gnd cell_6t
Xbit_r507_c125 bl[125] br[125] wl[507] vdd gnd cell_6t
Xbit_r508_c125 bl[125] br[125] wl[508] vdd gnd cell_6t
Xbit_r509_c125 bl[125] br[125] wl[509] vdd gnd cell_6t
Xbit_r510_c125 bl[125] br[125] wl[510] vdd gnd cell_6t
Xbit_r511_c125 bl[125] br[125] wl[511] vdd gnd cell_6t
Xbit_r0_c126 bl[126] br[126] wl[0] vdd gnd cell_6t
Xbit_r1_c126 bl[126] br[126] wl[1] vdd gnd cell_6t
Xbit_r2_c126 bl[126] br[126] wl[2] vdd gnd cell_6t
Xbit_r3_c126 bl[126] br[126] wl[3] vdd gnd cell_6t
Xbit_r4_c126 bl[126] br[126] wl[4] vdd gnd cell_6t
Xbit_r5_c126 bl[126] br[126] wl[5] vdd gnd cell_6t
Xbit_r6_c126 bl[126] br[126] wl[6] vdd gnd cell_6t
Xbit_r7_c126 bl[126] br[126] wl[7] vdd gnd cell_6t
Xbit_r8_c126 bl[126] br[126] wl[8] vdd gnd cell_6t
Xbit_r9_c126 bl[126] br[126] wl[9] vdd gnd cell_6t
Xbit_r10_c126 bl[126] br[126] wl[10] vdd gnd cell_6t
Xbit_r11_c126 bl[126] br[126] wl[11] vdd gnd cell_6t
Xbit_r12_c126 bl[126] br[126] wl[12] vdd gnd cell_6t
Xbit_r13_c126 bl[126] br[126] wl[13] vdd gnd cell_6t
Xbit_r14_c126 bl[126] br[126] wl[14] vdd gnd cell_6t
Xbit_r15_c126 bl[126] br[126] wl[15] vdd gnd cell_6t
Xbit_r16_c126 bl[126] br[126] wl[16] vdd gnd cell_6t
Xbit_r17_c126 bl[126] br[126] wl[17] vdd gnd cell_6t
Xbit_r18_c126 bl[126] br[126] wl[18] vdd gnd cell_6t
Xbit_r19_c126 bl[126] br[126] wl[19] vdd gnd cell_6t
Xbit_r20_c126 bl[126] br[126] wl[20] vdd gnd cell_6t
Xbit_r21_c126 bl[126] br[126] wl[21] vdd gnd cell_6t
Xbit_r22_c126 bl[126] br[126] wl[22] vdd gnd cell_6t
Xbit_r23_c126 bl[126] br[126] wl[23] vdd gnd cell_6t
Xbit_r24_c126 bl[126] br[126] wl[24] vdd gnd cell_6t
Xbit_r25_c126 bl[126] br[126] wl[25] vdd gnd cell_6t
Xbit_r26_c126 bl[126] br[126] wl[26] vdd gnd cell_6t
Xbit_r27_c126 bl[126] br[126] wl[27] vdd gnd cell_6t
Xbit_r28_c126 bl[126] br[126] wl[28] vdd gnd cell_6t
Xbit_r29_c126 bl[126] br[126] wl[29] vdd gnd cell_6t
Xbit_r30_c126 bl[126] br[126] wl[30] vdd gnd cell_6t
Xbit_r31_c126 bl[126] br[126] wl[31] vdd gnd cell_6t
Xbit_r32_c126 bl[126] br[126] wl[32] vdd gnd cell_6t
Xbit_r33_c126 bl[126] br[126] wl[33] vdd gnd cell_6t
Xbit_r34_c126 bl[126] br[126] wl[34] vdd gnd cell_6t
Xbit_r35_c126 bl[126] br[126] wl[35] vdd gnd cell_6t
Xbit_r36_c126 bl[126] br[126] wl[36] vdd gnd cell_6t
Xbit_r37_c126 bl[126] br[126] wl[37] vdd gnd cell_6t
Xbit_r38_c126 bl[126] br[126] wl[38] vdd gnd cell_6t
Xbit_r39_c126 bl[126] br[126] wl[39] vdd gnd cell_6t
Xbit_r40_c126 bl[126] br[126] wl[40] vdd gnd cell_6t
Xbit_r41_c126 bl[126] br[126] wl[41] vdd gnd cell_6t
Xbit_r42_c126 bl[126] br[126] wl[42] vdd gnd cell_6t
Xbit_r43_c126 bl[126] br[126] wl[43] vdd gnd cell_6t
Xbit_r44_c126 bl[126] br[126] wl[44] vdd gnd cell_6t
Xbit_r45_c126 bl[126] br[126] wl[45] vdd gnd cell_6t
Xbit_r46_c126 bl[126] br[126] wl[46] vdd gnd cell_6t
Xbit_r47_c126 bl[126] br[126] wl[47] vdd gnd cell_6t
Xbit_r48_c126 bl[126] br[126] wl[48] vdd gnd cell_6t
Xbit_r49_c126 bl[126] br[126] wl[49] vdd gnd cell_6t
Xbit_r50_c126 bl[126] br[126] wl[50] vdd gnd cell_6t
Xbit_r51_c126 bl[126] br[126] wl[51] vdd gnd cell_6t
Xbit_r52_c126 bl[126] br[126] wl[52] vdd gnd cell_6t
Xbit_r53_c126 bl[126] br[126] wl[53] vdd gnd cell_6t
Xbit_r54_c126 bl[126] br[126] wl[54] vdd gnd cell_6t
Xbit_r55_c126 bl[126] br[126] wl[55] vdd gnd cell_6t
Xbit_r56_c126 bl[126] br[126] wl[56] vdd gnd cell_6t
Xbit_r57_c126 bl[126] br[126] wl[57] vdd gnd cell_6t
Xbit_r58_c126 bl[126] br[126] wl[58] vdd gnd cell_6t
Xbit_r59_c126 bl[126] br[126] wl[59] vdd gnd cell_6t
Xbit_r60_c126 bl[126] br[126] wl[60] vdd gnd cell_6t
Xbit_r61_c126 bl[126] br[126] wl[61] vdd gnd cell_6t
Xbit_r62_c126 bl[126] br[126] wl[62] vdd gnd cell_6t
Xbit_r63_c126 bl[126] br[126] wl[63] vdd gnd cell_6t
Xbit_r64_c126 bl[126] br[126] wl[64] vdd gnd cell_6t
Xbit_r65_c126 bl[126] br[126] wl[65] vdd gnd cell_6t
Xbit_r66_c126 bl[126] br[126] wl[66] vdd gnd cell_6t
Xbit_r67_c126 bl[126] br[126] wl[67] vdd gnd cell_6t
Xbit_r68_c126 bl[126] br[126] wl[68] vdd gnd cell_6t
Xbit_r69_c126 bl[126] br[126] wl[69] vdd gnd cell_6t
Xbit_r70_c126 bl[126] br[126] wl[70] vdd gnd cell_6t
Xbit_r71_c126 bl[126] br[126] wl[71] vdd gnd cell_6t
Xbit_r72_c126 bl[126] br[126] wl[72] vdd gnd cell_6t
Xbit_r73_c126 bl[126] br[126] wl[73] vdd gnd cell_6t
Xbit_r74_c126 bl[126] br[126] wl[74] vdd gnd cell_6t
Xbit_r75_c126 bl[126] br[126] wl[75] vdd gnd cell_6t
Xbit_r76_c126 bl[126] br[126] wl[76] vdd gnd cell_6t
Xbit_r77_c126 bl[126] br[126] wl[77] vdd gnd cell_6t
Xbit_r78_c126 bl[126] br[126] wl[78] vdd gnd cell_6t
Xbit_r79_c126 bl[126] br[126] wl[79] vdd gnd cell_6t
Xbit_r80_c126 bl[126] br[126] wl[80] vdd gnd cell_6t
Xbit_r81_c126 bl[126] br[126] wl[81] vdd gnd cell_6t
Xbit_r82_c126 bl[126] br[126] wl[82] vdd gnd cell_6t
Xbit_r83_c126 bl[126] br[126] wl[83] vdd gnd cell_6t
Xbit_r84_c126 bl[126] br[126] wl[84] vdd gnd cell_6t
Xbit_r85_c126 bl[126] br[126] wl[85] vdd gnd cell_6t
Xbit_r86_c126 bl[126] br[126] wl[86] vdd gnd cell_6t
Xbit_r87_c126 bl[126] br[126] wl[87] vdd gnd cell_6t
Xbit_r88_c126 bl[126] br[126] wl[88] vdd gnd cell_6t
Xbit_r89_c126 bl[126] br[126] wl[89] vdd gnd cell_6t
Xbit_r90_c126 bl[126] br[126] wl[90] vdd gnd cell_6t
Xbit_r91_c126 bl[126] br[126] wl[91] vdd gnd cell_6t
Xbit_r92_c126 bl[126] br[126] wl[92] vdd gnd cell_6t
Xbit_r93_c126 bl[126] br[126] wl[93] vdd gnd cell_6t
Xbit_r94_c126 bl[126] br[126] wl[94] vdd gnd cell_6t
Xbit_r95_c126 bl[126] br[126] wl[95] vdd gnd cell_6t
Xbit_r96_c126 bl[126] br[126] wl[96] vdd gnd cell_6t
Xbit_r97_c126 bl[126] br[126] wl[97] vdd gnd cell_6t
Xbit_r98_c126 bl[126] br[126] wl[98] vdd gnd cell_6t
Xbit_r99_c126 bl[126] br[126] wl[99] vdd gnd cell_6t
Xbit_r100_c126 bl[126] br[126] wl[100] vdd gnd cell_6t
Xbit_r101_c126 bl[126] br[126] wl[101] vdd gnd cell_6t
Xbit_r102_c126 bl[126] br[126] wl[102] vdd gnd cell_6t
Xbit_r103_c126 bl[126] br[126] wl[103] vdd gnd cell_6t
Xbit_r104_c126 bl[126] br[126] wl[104] vdd gnd cell_6t
Xbit_r105_c126 bl[126] br[126] wl[105] vdd gnd cell_6t
Xbit_r106_c126 bl[126] br[126] wl[106] vdd gnd cell_6t
Xbit_r107_c126 bl[126] br[126] wl[107] vdd gnd cell_6t
Xbit_r108_c126 bl[126] br[126] wl[108] vdd gnd cell_6t
Xbit_r109_c126 bl[126] br[126] wl[109] vdd gnd cell_6t
Xbit_r110_c126 bl[126] br[126] wl[110] vdd gnd cell_6t
Xbit_r111_c126 bl[126] br[126] wl[111] vdd gnd cell_6t
Xbit_r112_c126 bl[126] br[126] wl[112] vdd gnd cell_6t
Xbit_r113_c126 bl[126] br[126] wl[113] vdd gnd cell_6t
Xbit_r114_c126 bl[126] br[126] wl[114] vdd gnd cell_6t
Xbit_r115_c126 bl[126] br[126] wl[115] vdd gnd cell_6t
Xbit_r116_c126 bl[126] br[126] wl[116] vdd gnd cell_6t
Xbit_r117_c126 bl[126] br[126] wl[117] vdd gnd cell_6t
Xbit_r118_c126 bl[126] br[126] wl[118] vdd gnd cell_6t
Xbit_r119_c126 bl[126] br[126] wl[119] vdd gnd cell_6t
Xbit_r120_c126 bl[126] br[126] wl[120] vdd gnd cell_6t
Xbit_r121_c126 bl[126] br[126] wl[121] vdd gnd cell_6t
Xbit_r122_c126 bl[126] br[126] wl[122] vdd gnd cell_6t
Xbit_r123_c126 bl[126] br[126] wl[123] vdd gnd cell_6t
Xbit_r124_c126 bl[126] br[126] wl[124] vdd gnd cell_6t
Xbit_r125_c126 bl[126] br[126] wl[125] vdd gnd cell_6t
Xbit_r126_c126 bl[126] br[126] wl[126] vdd gnd cell_6t
Xbit_r127_c126 bl[126] br[126] wl[127] vdd gnd cell_6t
Xbit_r128_c126 bl[126] br[126] wl[128] vdd gnd cell_6t
Xbit_r129_c126 bl[126] br[126] wl[129] vdd gnd cell_6t
Xbit_r130_c126 bl[126] br[126] wl[130] vdd gnd cell_6t
Xbit_r131_c126 bl[126] br[126] wl[131] vdd gnd cell_6t
Xbit_r132_c126 bl[126] br[126] wl[132] vdd gnd cell_6t
Xbit_r133_c126 bl[126] br[126] wl[133] vdd gnd cell_6t
Xbit_r134_c126 bl[126] br[126] wl[134] vdd gnd cell_6t
Xbit_r135_c126 bl[126] br[126] wl[135] vdd gnd cell_6t
Xbit_r136_c126 bl[126] br[126] wl[136] vdd gnd cell_6t
Xbit_r137_c126 bl[126] br[126] wl[137] vdd gnd cell_6t
Xbit_r138_c126 bl[126] br[126] wl[138] vdd gnd cell_6t
Xbit_r139_c126 bl[126] br[126] wl[139] vdd gnd cell_6t
Xbit_r140_c126 bl[126] br[126] wl[140] vdd gnd cell_6t
Xbit_r141_c126 bl[126] br[126] wl[141] vdd gnd cell_6t
Xbit_r142_c126 bl[126] br[126] wl[142] vdd gnd cell_6t
Xbit_r143_c126 bl[126] br[126] wl[143] vdd gnd cell_6t
Xbit_r144_c126 bl[126] br[126] wl[144] vdd gnd cell_6t
Xbit_r145_c126 bl[126] br[126] wl[145] vdd gnd cell_6t
Xbit_r146_c126 bl[126] br[126] wl[146] vdd gnd cell_6t
Xbit_r147_c126 bl[126] br[126] wl[147] vdd gnd cell_6t
Xbit_r148_c126 bl[126] br[126] wl[148] vdd gnd cell_6t
Xbit_r149_c126 bl[126] br[126] wl[149] vdd gnd cell_6t
Xbit_r150_c126 bl[126] br[126] wl[150] vdd gnd cell_6t
Xbit_r151_c126 bl[126] br[126] wl[151] vdd gnd cell_6t
Xbit_r152_c126 bl[126] br[126] wl[152] vdd gnd cell_6t
Xbit_r153_c126 bl[126] br[126] wl[153] vdd gnd cell_6t
Xbit_r154_c126 bl[126] br[126] wl[154] vdd gnd cell_6t
Xbit_r155_c126 bl[126] br[126] wl[155] vdd gnd cell_6t
Xbit_r156_c126 bl[126] br[126] wl[156] vdd gnd cell_6t
Xbit_r157_c126 bl[126] br[126] wl[157] vdd gnd cell_6t
Xbit_r158_c126 bl[126] br[126] wl[158] vdd gnd cell_6t
Xbit_r159_c126 bl[126] br[126] wl[159] vdd gnd cell_6t
Xbit_r160_c126 bl[126] br[126] wl[160] vdd gnd cell_6t
Xbit_r161_c126 bl[126] br[126] wl[161] vdd gnd cell_6t
Xbit_r162_c126 bl[126] br[126] wl[162] vdd gnd cell_6t
Xbit_r163_c126 bl[126] br[126] wl[163] vdd gnd cell_6t
Xbit_r164_c126 bl[126] br[126] wl[164] vdd gnd cell_6t
Xbit_r165_c126 bl[126] br[126] wl[165] vdd gnd cell_6t
Xbit_r166_c126 bl[126] br[126] wl[166] vdd gnd cell_6t
Xbit_r167_c126 bl[126] br[126] wl[167] vdd gnd cell_6t
Xbit_r168_c126 bl[126] br[126] wl[168] vdd gnd cell_6t
Xbit_r169_c126 bl[126] br[126] wl[169] vdd gnd cell_6t
Xbit_r170_c126 bl[126] br[126] wl[170] vdd gnd cell_6t
Xbit_r171_c126 bl[126] br[126] wl[171] vdd gnd cell_6t
Xbit_r172_c126 bl[126] br[126] wl[172] vdd gnd cell_6t
Xbit_r173_c126 bl[126] br[126] wl[173] vdd gnd cell_6t
Xbit_r174_c126 bl[126] br[126] wl[174] vdd gnd cell_6t
Xbit_r175_c126 bl[126] br[126] wl[175] vdd gnd cell_6t
Xbit_r176_c126 bl[126] br[126] wl[176] vdd gnd cell_6t
Xbit_r177_c126 bl[126] br[126] wl[177] vdd gnd cell_6t
Xbit_r178_c126 bl[126] br[126] wl[178] vdd gnd cell_6t
Xbit_r179_c126 bl[126] br[126] wl[179] vdd gnd cell_6t
Xbit_r180_c126 bl[126] br[126] wl[180] vdd gnd cell_6t
Xbit_r181_c126 bl[126] br[126] wl[181] vdd gnd cell_6t
Xbit_r182_c126 bl[126] br[126] wl[182] vdd gnd cell_6t
Xbit_r183_c126 bl[126] br[126] wl[183] vdd gnd cell_6t
Xbit_r184_c126 bl[126] br[126] wl[184] vdd gnd cell_6t
Xbit_r185_c126 bl[126] br[126] wl[185] vdd gnd cell_6t
Xbit_r186_c126 bl[126] br[126] wl[186] vdd gnd cell_6t
Xbit_r187_c126 bl[126] br[126] wl[187] vdd gnd cell_6t
Xbit_r188_c126 bl[126] br[126] wl[188] vdd gnd cell_6t
Xbit_r189_c126 bl[126] br[126] wl[189] vdd gnd cell_6t
Xbit_r190_c126 bl[126] br[126] wl[190] vdd gnd cell_6t
Xbit_r191_c126 bl[126] br[126] wl[191] vdd gnd cell_6t
Xbit_r192_c126 bl[126] br[126] wl[192] vdd gnd cell_6t
Xbit_r193_c126 bl[126] br[126] wl[193] vdd gnd cell_6t
Xbit_r194_c126 bl[126] br[126] wl[194] vdd gnd cell_6t
Xbit_r195_c126 bl[126] br[126] wl[195] vdd gnd cell_6t
Xbit_r196_c126 bl[126] br[126] wl[196] vdd gnd cell_6t
Xbit_r197_c126 bl[126] br[126] wl[197] vdd gnd cell_6t
Xbit_r198_c126 bl[126] br[126] wl[198] vdd gnd cell_6t
Xbit_r199_c126 bl[126] br[126] wl[199] vdd gnd cell_6t
Xbit_r200_c126 bl[126] br[126] wl[200] vdd gnd cell_6t
Xbit_r201_c126 bl[126] br[126] wl[201] vdd gnd cell_6t
Xbit_r202_c126 bl[126] br[126] wl[202] vdd gnd cell_6t
Xbit_r203_c126 bl[126] br[126] wl[203] vdd gnd cell_6t
Xbit_r204_c126 bl[126] br[126] wl[204] vdd gnd cell_6t
Xbit_r205_c126 bl[126] br[126] wl[205] vdd gnd cell_6t
Xbit_r206_c126 bl[126] br[126] wl[206] vdd gnd cell_6t
Xbit_r207_c126 bl[126] br[126] wl[207] vdd gnd cell_6t
Xbit_r208_c126 bl[126] br[126] wl[208] vdd gnd cell_6t
Xbit_r209_c126 bl[126] br[126] wl[209] vdd gnd cell_6t
Xbit_r210_c126 bl[126] br[126] wl[210] vdd gnd cell_6t
Xbit_r211_c126 bl[126] br[126] wl[211] vdd gnd cell_6t
Xbit_r212_c126 bl[126] br[126] wl[212] vdd gnd cell_6t
Xbit_r213_c126 bl[126] br[126] wl[213] vdd gnd cell_6t
Xbit_r214_c126 bl[126] br[126] wl[214] vdd gnd cell_6t
Xbit_r215_c126 bl[126] br[126] wl[215] vdd gnd cell_6t
Xbit_r216_c126 bl[126] br[126] wl[216] vdd gnd cell_6t
Xbit_r217_c126 bl[126] br[126] wl[217] vdd gnd cell_6t
Xbit_r218_c126 bl[126] br[126] wl[218] vdd gnd cell_6t
Xbit_r219_c126 bl[126] br[126] wl[219] vdd gnd cell_6t
Xbit_r220_c126 bl[126] br[126] wl[220] vdd gnd cell_6t
Xbit_r221_c126 bl[126] br[126] wl[221] vdd gnd cell_6t
Xbit_r222_c126 bl[126] br[126] wl[222] vdd gnd cell_6t
Xbit_r223_c126 bl[126] br[126] wl[223] vdd gnd cell_6t
Xbit_r224_c126 bl[126] br[126] wl[224] vdd gnd cell_6t
Xbit_r225_c126 bl[126] br[126] wl[225] vdd gnd cell_6t
Xbit_r226_c126 bl[126] br[126] wl[226] vdd gnd cell_6t
Xbit_r227_c126 bl[126] br[126] wl[227] vdd gnd cell_6t
Xbit_r228_c126 bl[126] br[126] wl[228] vdd gnd cell_6t
Xbit_r229_c126 bl[126] br[126] wl[229] vdd gnd cell_6t
Xbit_r230_c126 bl[126] br[126] wl[230] vdd gnd cell_6t
Xbit_r231_c126 bl[126] br[126] wl[231] vdd gnd cell_6t
Xbit_r232_c126 bl[126] br[126] wl[232] vdd gnd cell_6t
Xbit_r233_c126 bl[126] br[126] wl[233] vdd gnd cell_6t
Xbit_r234_c126 bl[126] br[126] wl[234] vdd gnd cell_6t
Xbit_r235_c126 bl[126] br[126] wl[235] vdd gnd cell_6t
Xbit_r236_c126 bl[126] br[126] wl[236] vdd gnd cell_6t
Xbit_r237_c126 bl[126] br[126] wl[237] vdd gnd cell_6t
Xbit_r238_c126 bl[126] br[126] wl[238] vdd gnd cell_6t
Xbit_r239_c126 bl[126] br[126] wl[239] vdd gnd cell_6t
Xbit_r240_c126 bl[126] br[126] wl[240] vdd gnd cell_6t
Xbit_r241_c126 bl[126] br[126] wl[241] vdd gnd cell_6t
Xbit_r242_c126 bl[126] br[126] wl[242] vdd gnd cell_6t
Xbit_r243_c126 bl[126] br[126] wl[243] vdd gnd cell_6t
Xbit_r244_c126 bl[126] br[126] wl[244] vdd gnd cell_6t
Xbit_r245_c126 bl[126] br[126] wl[245] vdd gnd cell_6t
Xbit_r246_c126 bl[126] br[126] wl[246] vdd gnd cell_6t
Xbit_r247_c126 bl[126] br[126] wl[247] vdd gnd cell_6t
Xbit_r248_c126 bl[126] br[126] wl[248] vdd gnd cell_6t
Xbit_r249_c126 bl[126] br[126] wl[249] vdd gnd cell_6t
Xbit_r250_c126 bl[126] br[126] wl[250] vdd gnd cell_6t
Xbit_r251_c126 bl[126] br[126] wl[251] vdd gnd cell_6t
Xbit_r252_c126 bl[126] br[126] wl[252] vdd gnd cell_6t
Xbit_r253_c126 bl[126] br[126] wl[253] vdd gnd cell_6t
Xbit_r254_c126 bl[126] br[126] wl[254] vdd gnd cell_6t
Xbit_r255_c126 bl[126] br[126] wl[255] vdd gnd cell_6t
Xbit_r256_c126 bl[126] br[126] wl[256] vdd gnd cell_6t
Xbit_r257_c126 bl[126] br[126] wl[257] vdd gnd cell_6t
Xbit_r258_c126 bl[126] br[126] wl[258] vdd gnd cell_6t
Xbit_r259_c126 bl[126] br[126] wl[259] vdd gnd cell_6t
Xbit_r260_c126 bl[126] br[126] wl[260] vdd gnd cell_6t
Xbit_r261_c126 bl[126] br[126] wl[261] vdd gnd cell_6t
Xbit_r262_c126 bl[126] br[126] wl[262] vdd gnd cell_6t
Xbit_r263_c126 bl[126] br[126] wl[263] vdd gnd cell_6t
Xbit_r264_c126 bl[126] br[126] wl[264] vdd gnd cell_6t
Xbit_r265_c126 bl[126] br[126] wl[265] vdd gnd cell_6t
Xbit_r266_c126 bl[126] br[126] wl[266] vdd gnd cell_6t
Xbit_r267_c126 bl[126] br[126] wl[267] vdd gnd cell_6t
Xbit_r268_c126 bl[126] br[126] wl[268] vdd gnd cell_6t
Xbit_r269_c126 bl[126] br[126] wl[269] vdd gnd cell_6t
Xbit_r270_c126 bl[126] br[126] wl[270] vdd gnd cell_6t
Xbit_r271_c126 bl[126] br[126] wl[271] vdd gnd cell_6t
Xbit_r272_c126 bl[126] br[126] wl[272] vdd gnd cell_6t
Xbit_r273_c126 bl[126] br[126] wl[273] vdd gnd cell_6t
Xbit_r274_c126 bl[126] br[126] wl[274] vdd gnd cell_6t
Xbit_r275_c126 bl[126] br[126] wl[275] vdd gnd cell_6t
Xbit_r276_c126 bl[126] br[126] wl[276] vdd gnd cell_6t
Xbit_r277_c126 bl[126] br[126] wl[277] vdd gnd cell_6t
Xbit_r278_c126 bl[126] br[126] wl[278] vdd gnd cell_6t
Xbit_r279_c126 bl[126] br[126] wl[279] vdd gnd cell_6t
Xbit_r280_c126 bl[126] br[126] wl[280] vdd gnd cell_6t
Xbit_r281_c126 bl[126] br[126] wl[281] vdd gnd cell_6t
Xbit_r282_c126 bl[126] br[126] wl[282] vdd gnd cell_6t
Xbit_r283_c126 bl[126] br[126] wl[283] vdd gnd cell_6t
Xbit_r284_c126 bl[126] br[126] wl[284] vdd gnd cell_6t
Xbit_r285_c126 bl[126] br[126] wl[285] vdd gnd cell_6t
Xbit_r286_c126 bl[126] br[126] wl[286] vdd gnd cell_6t
Xbit_r287_c126 bl[126] br[126] wl[287] vdd gnd cell_6t
Xbit_r288_c126 bl[126] br[126] wl[288] vdd gnd cell_6t
Xbit_r289_c126 bl[126] br[126] wl[289] vdd gnd cell_6t
Xbit_r290_c126 bl[126] br[126] wl[290] vdd gnd cell_6t
Xbit_r291_c126 bl[126] br[126] wl[291] vdd gnd cell_6t
Xbit_r292_c126 bl[126] br[126] wl[292] vdd gnd cell_6t
Xbit_r293_c126 bl[126] br[126] wl[293] vdd gnd cell_6t
Xbit_r294_c126 bl[126] br[126] wl[294] vdd gnd cell_6t
Xbit_r295_c126 bl[126] br[126] wl[295] vdd gnd cell_6t
Xbit_r296_c126 bl[126] br[126] wl[296] vdd gnd cell_6t
Xbit_r297_c126 bl[126] br[126] wl[297] vdd gnd cell_6t
Xbit_r298_c126 bl[126] br[126] wl[298] vdd gnd cell_6t
Xbit_r299_c126 bl[126] br[126] wl[299] vdd gnd cell_6t
Xbit_r300_c126 bl[126] br[126] wl[300] vdd gnd cell_6t
Xbit_r301_c126 bl[126] br[126] wl[301] vdd gnd cell_6t
Xbit_r302_c126 bl[126] br[126] wl[302] vdd gnd cell_6t
Xbit_r303_c126 bl[126] br[126] wl[303] vdd gnd cell_6t
Xbit_r304_c126 bl[126] br[126] wl[304] vdd gnd cell_6t
Xbit_r305_c126 bl[126] br[126] wl[305] vdd gnd cell_6t
Xbit_r306_c126 bl[126] br[126] wl[306] vdd gnd cell_6t
Xbit_r307_c126 bl[126] br[126] wl[307] vdd gnd cell_6t
Xbit_r308_c126 bl[126] br[126] wl[308] vdd gnd cell_6t
Xbit_r309_c126 bl[126] br[126] wl[309] vdd gnd cell_6t
Xbit_r310_c126 bl[126] br[126] wl[310] vdd gnd cell_6t
Xbit_r311_c126 bl[126] br[126] wl[311] vdd gnd cell_6t
Xbit_r312_c126 bl[126] br[126] wl[312] vdd gnd cell_6t
Xbit_r313_c126 bl[126] br[126] wl[313] vdd gnd cell_6t
Xbit_r314_c126 bl[126] br[126] wl[314] vdd gnd cell_6t
Xbit_r315_c126 bl[126] br[126] wl[315] vdd gnd cell_6t
Xbit_r316_c126 bl[126] br[126] wl[316] vdd gnd cell_6t
Xbit_r317_c126 bl[126] br[126] wl[317] vdd gnd cell_6t
Xbit_r318_c126 bl[126] br[126] wl[318] vdd gnd cell_6t
Xbit_r319_c126 bl[126] br[126] wl[319] vdd gnd cell_6t
Xbit_r320_c126 bl[126] br[126] wl[320] vdd gnd cell_6t
Xbit_r321_c126 bl[126] br[126] wl[321] vdd gnd cell_6t
Xbit_r322_c126 bl[126] br[126] wl[322] vdd gnd cell_6t
Xbit_r323_c126 bl[126] br[126] wl[323] vdd gnd cell_6t
Xbit_r324_c126 bl[126] br[126] wl[324] vdd gnd cell_6t
Xbit_r325_c126 bl[126] br[126] wl[325] vdd gnd cell_6t
Xbit_r326_c126 bl[126] br[126] wl[326] vdd gnd cell_6t
Xbit_r327_c126 bl[126] br[126] wl[327] vdd gnd cell_6t
Xbit_r328_c126 bl[126] br[126] wl[328] vdd gnd cell_6t
Xbit_r329_c126 bl[126] br[126] wl[329] vdd gnd cell_6t
Xbit_r330_c126 bl[126] br[126] wl[330] vdd gnd cell_6t
Xbit_r331_c126 bl[126] br[126] wl[331] vdd gnd cell_6t
Xbit_r332_c126 bl[126] br[126] wl[332] vdd gnd cell_6t
Xbit_r333_c126 bl[126] br[126] wl[333] vdd gnd cell_6t
Xbit_r334_c126 bl[126] br[126] wl[334] vdd gnd cell_6t
Xbit_r335_c126 bl[126] br[126] wl[335] vdd gnd cell_6t
Xbit_r336_c126 bl[126] br[126] wl[336] vdd gnd cell_6t
Xbit_r337_c126 bl[126] br[126] wl[337] vdd gnd cell_6t
Xbit_r338_c126 bl[126] br[126] wl[338] vdd gnd cell_6t
Xbit_r339_c126 bl[126] br[126] wl[339] vdd gnd cell_6t
Xbit_r340_c126 bl[126] br[126] wl[340] vdd gnd cell_6t
Xbit_r341_c126 bl[126] br[126] wl[341] vdd gnd cell_6t
Xbit_r342_c126 bl[126] br[126] wl[342] vdd gnd cell_6t
Xbit_r343_c126 bl[126] br[126] wl[343] vdd gnd cell_6t
Xbit_r344_c126 bl[126] br[126] wl[344] vdd gnd cell_6t
Xbit_r345_c126 bl[126] br[126] wl[345] vdd gnd cell_6t
Xbit_r346_c126 bl[126] br[126] wl[346] vdd gnd cell_6t
Xbit_r347_c126 bl[126] br[126] wl[347] vdd gnd cell_6t
Xbit_r348_c126 bl[126] br[126] wl[348] vdd gnd cell_6t
Xbit_r349_c126 bl[126] br[126] wl[349] vdd gnd cell_6t
Xbit_r350_c126 bl[126] br[126] wl[350] vdd gnd cell_6t
Xbit_r351_c126 bl[126] br[126] wl[351] vdd gnd cell_6t
Xbit_r352_c126 bl[126] br[126] wl[352] vdd gnd cell_6t
Xbit_r353_c126 bl[126] br[126] wl[353] vdd gnd cell_6t
Xbit_r354_c126 bl[126] br[126] wl[354] vdd gnd cell_6t
Xbit_r355_c126 bl[126] br[126] wl[355] vdd gnd cell_6t
Xbit_r356_c126 bl[126] br[126] wl[356] vdd gnd cell_6t
Xbit_r357_c126 bl[126] br[126] wl[357] vdd gnd cell_6t
Xbit_r358_c126 bl[126] br[126] wl[358] vdd gnd cell_6t
Xbit_r359_c126 bl[126] br[126] wl[359] vdd gnd cell_6t
Xbit_r360_c126 bl[126] br[126] wl[360] vdd gnd cell_6t
Xbit_r361_c126 bl[126] br[126] wl[361] vdd gnd cell_6t
Xbit_r362_c126 bl[126] br[126] wl[362] vdd gnd cell_6t
Xbit_r363_c126 bl[126] br[126] wl[363] vdd gnd cell_6t
Xbit_r364_c126 bl[126] br[126] wl[364] vdd gnd cell_6t
Xbit_r365_c126 bl[126] br[126] wl[365] vdd gnd cell_6t
Xbit_r366_c126 bl[126] br[126] wl[366] vdd gnd cell_6t
Xbit_r367_c126 bl[126] br[126] wl[367] vdd gnd cell_6t
Xbit_r368_c126 bl[126] br[126] wl[368] vdd gnd cell_6t
Xbit_r369_c126 bl[126] br[126] wl[369] vdd gnd cell_6t
Xbit_r370_c126 bl[126] br[126] wl[370] vdd gnd cell_6t
Xbit_r371_c126 bl[126] br[126] wl[371] vdd gnd cell_6t
Xbit_r372_c126 bl[126] br[126] wl[372] vdd gnd cell_6t
Xbit_r373_c126 bl[126] br[126] wl[373] vdd gnd cell_6t
Xbit_r374_c126 bl[126] br[126] wl[374] vdd gnd cell_6t
Xbit_r375_c126 bl[126] br[126] wl[375] vdd gnd cell_6t
Xbit_r376_c126 bl[126] br[126] wl[376] vdd gnd cell_6t
Xbit_r377_c126 bl[126] br[126] wl[377] vdd gnd cell_6t
Xbit_r378_c126 bl[126] br[126] wl[378] vdd gnd cell_6t
Xbit_r379_c126 bl[126] br[126] wl[379] vdd gnd cell_6t
Xbit_r380_c126 bl[126] br[126] wl[380] vdd gnd cell_6t
Xbit_r381_c126 bl[126] br[126] wl[381] vdd gnd cell_6t
Xbit_r382_c126 bl[126] br[126] wl[382] vdd gnd cell_6t
Xbit_r383_c126 bl[126] br[126] wl[383] vdd gnd cell_6t
Xbit_r384_c126 bl[126] br[126] wl[384] vdd gnd cell_6t
Xbit_r385_c126 bl[126] br[126] wl[385] vdd gnd cell_6t
Xbit_r386_c126 bl[126] br[126] wl[386] vdd gnd cell_6t
Xbit_r387_c126 bl[126] br[126] wl[387] vdd gnd cell_6t
Xbit_r388_c126 bl[126] br[126] wl[388] vdd gnd cell_6t
Xbit_r389_c126 bl[126] br[126] wl[389] vdd gnd cell_6t
Xbit_r390_c126 bl[126] br[126] wl[390] vdd gnd cell_6t
Xbit_r391_c126 bl[126] br[126] wl[391] vdd gnd cell_6t
Xbit_r392_c126 bl[126] br[126] wl[392] vdd gnd cell_6t
Xbit_r393_c126 bl[126] br[126] wl[393] vdd gnd cell_6t
Xbit_r394_c126 bl[126] br[126] wl[394] vdd gnd cell_6t
Xbit_r395_c126 bl[126] br[126] wl[395] vdd gnd cell_6t
Xbit_r396_c126 bl[126] br[126] wl[396] vdd gnd cell_6t
Xbit_r397_c126 bl[126] br[126] wl[397] vdd gnd cell_6t
Xbit_r398_c126 bl[126] br[126] wl[398] vdd gnd cell_6t
Xbit_r399_c126 bl[126] br[126] wl[399] vdd gnd cell_6t
Xbit_r400_c126 bl[126] br[126] wl[400] vdd gnd cell_6t
Xbit_r401_c126 bl[126] br[126] wl[401] vdd gnd cell_6t
Xbit_r402_c126 bl[126] br[126] wl[402] vdd gnd cell_6t
Xbit_r403_c126 bl[126] br[126] wl[403] vdd gnd cell_6t
Xbit_r404_c126 bl[126] br[126] wl[404] vdd gnd cell_6t
Xbit_r405_c126 bl[126] br[126] wl[405] vdd gnd cell_6t
Xbit_r406_c126 bl[126] br[126] wl[406] vdd gnd cell_6t
Xbit_r407_c126 bl[126] br[126] wl[407] vdd gnd cell_6t
Xbit_r408_c126 bl[126] br[126] wl[408] vdd gnd cell_6t
Xbit_r409_c126 bl[126] br[126] wl[409] vdd gnd cell_6t
Xbit_r410_c126 bl[126] br[126] wl[410] vdd gnd cell_6t
Xbit_r411_c126 bl[126] br[126] wl[411] vdd gnd cell_6t
Xbit_r412_c126 bl[126] br[126] wl[412] vdd gnd cell_6t
Xbit_r413_c126 bl[126] br[126] wl[413] vdd gnd cell_6t
Xbit_r414_c126 bl[126] br[126] wl[414] vdd gnd cell_6t
Xbit_r415_c126 bl[126] br[126] wl[415] vdd gnd cell_6t
Xbit_r416_c126 bl[126] br[126] wl[416] vdd gnd cell_6t
Xbit_r417_c126 bl[126] br[126] wl[417] vdd gnd cell_6t
Xbit_r418_c126 bl[126] br[126] wl[418] vdd gnd cell_6t
Xbit_r419_c126 bl[126] br[126] wl[419] vdd gnd cell_6t
Xbit_r420_c126 bl[126] br[126] wl[420] vdd gnd cell_6t
Xbit_r421_c126 bl[126] br[126] wl[421] vdd gnd cell_6t
Xbit_r422_c126 bl[126] br[126] wl[422] vdd gnd cell_6t
Xbit_r423_c126 bl[126] br[126] wl[423] vdd gnd cell_6t
Xbit_r424_c126 bl[126] br[126] wl[424] vdd gnd cell_6t
Xbit_r425_c126 bl[126] br[126] wl[425] vdd gnd cell_6t
Xbit_r426_c126 bl[126] br[126] wl[426] vdd gnd cell_6t
Xbit_r427_c126 bl[126] br[126] wl[427] vdd gnd cell_6t
Xbit_r428_c126 bl[126] br[126] wl[428] vdd gnd cell_6t
Xbit_r429_c126 bl[126] br[126] wl[429] vdd gnd cell_6t
Xbit_r430_c126 bl[126] br[126] wl[430] vdd gnd cell_6t
Xbit_r431_c126 bl[126] br[126] wl[431] vdd gnd cell_6t
Xbit_r432_c126 bl[126] br[126] wl[432] vdd gnd cell_6t
Xbit_r433_c126 bl[126] br[126] wl[433] vdd gnd cell_6t
Xbit_r434_c126 bl[126] br[126] wl[434] vdd gnd cell_6t
Xbit_r435_c126 bl[126] br[126] wl[435] vdd gnd cell_6t
Xbit_r436_c126 bl[126] br[126] wl[436] vdd gnd cell_6t
Xbit_r437_c126 bl[126] br[126] wl[437] vdd gnd cell_6t
Xbit_r438_c126 bl[126] br[126] wl[438] vdd gnd cell_6t
Xbit_r439_c126 bl[126] br[126] wl[439] vdd gnd cell_6t
Xbit_r440_c126 bl[126] br[126] wl[440] vdd gnd cell_6t
Xbit_r441_c126 bl[126] br[126] wl[441] vdd gnd cell_6t
Xbit_r442_c126 bl[126] br[126] wl[442] vdd gnd cell_6t
Xbit_r443_c126 bl[126] br[126] wl[443] vdd gnd cell_6t
Xbit_r444_c126 bl[126] br[126] wl[444] vdd gnd cell_6t
Xbit_r445_c126 bl[126] br[126] wl[445] vdd gnd cell_6t
Xbit_r446_c126 bl[126] br[126] wl[446] vdd gnd cell_6t
Xbit_r447_c126 bl[126] br[126] wl[447] vdd gnd cell_6t
Xbit_r448_c126 bl[126] br[126] wl[448] vdd gnd cell_6t
Xbit_r449_c126 bl[126] br[126] wl[449] vdd gnd cell_6t
Xbit_r450_c126 bl[126] br[126] wl[450] vdd gnd cell_6t
Xbit_r451_c126 bl[126] br[126] wl[451] vdd gnd cell_6t
Xbit_r452_c126 bl[126] br[126] wl[452] vdd gnd cell_6t
Xbit_r453_c126 bl[126] br[126] wl[453] vdd gnd cell_6t
Xbit_r454_c126 bl[126] br[126] wl[454] vdd gnd cell_6t
Xbit_r455_c126 bl[126] br[126] wl[455] vdd gnd cell_6t
Xbit_r456_c126 bl[126] br[126] wl[456] vdd gnd cell_6t
Xbit_r457_c126 bl[126] br[126] wl[457] vdd gnd cell_6t
Xbit_r458_c126 bl[126] br[126] wl[458] vdd gnd cell_6t
Xbit_r459_c126 bl[126] br[126] wl[459] vdd gnd cell_6t
Xbit_r460_c126 bl[126] br[126] wl[460] vdd gnd cell_6t
Xbit_r461_c126 bl[126] br[126] wl[461] vdd gnd cell_6t
Xbit_r462_c126 bl[126] br[126] wl[462] vdd gnd cell_6t
Xbit_r463_c126 bl[126] br[126] wl[463] vdd gnd cell_6t
Xbit_r464_c126 bl[126] br[126] wl[464] vdd gnd cell_6t
Xbit_r465_c126 bl[126] br[126] wl[465] vdd gnd cell_6t
Xbit_r466_c126 bl[126] br[126] wl[466] vdd gnd cell_6t
Xbit_r467_c126 bl[126] br[126] wl[467] vdd gnd cell_6t
Xbit_r468_c126 bl[126] br[126] wl[468] vdd gnd cell_6t
Xbit_r469_c126 bl[126] br[126] wl[469] vdd gnd cell_6t
Xbit_r470_c126 bl[126] br[126] wl[470] vdd gnd cell_6t
Xbit_r471_c126 bl[126] br[126] wl[471] vdd gnd cell_6t
Xbit_r472_c126 bl[126] br[126] wl[472] vdd gnd cell_6t
Xbit_r473_c126 bl[126] br[126] wl[473] vdd gnd cell_6t
Xbit_r474_c126 bl[126] br[126] wl[474] vdd gnd cell_6t
Xbit_r475_c126 bl[126] br[126] wl[475] vdd gnd cell_6t
Xbit_r476_c126 bl[126] br[126] wl[476] vdd gnd cell_6t
Xbit_r477_c126 bl[126] br[126] wl[477] vdd gnd cell_6t
Xbit_r478_c126 bl[126] br[126] wl[478] vdd gnd cell_6t
Xbit_r479_c126 bl[126] br[126] wl[479] vdd gnd cell_6t
Xbit_r480_c126 bl[126] br[126] wl[480] vdd gnd cell_6t
Xbit_r481_c126 bl[126] br[126] wl[481] vdd gnd cell_6t
Xbit_r482_c126 bl[126] br[126] wl[482] vdd gnd cell_6t
Xbit_r483_c126 bl[126] br[126] wl[483] vdd gnd cell_6t
Xbit_r484_c126 bl[126] br[126] wl[484] vdd gnd cell_6t
Xbit_r485_c126 bl[126] br[126] wl[485] vdd gnd cell_6t
Xbit_r486_c126 bl[126] br[126] wl[486] vdd gnd cell_6t
Xbit_r487_c126 bl[126] br[126] wl[487] vdd gnd cell_6t
Xbit_r488_c126 bl[126] br[126] wl[488] vdd gnd cell_6t
Xbit_r489_c126 bl[126] br[126] wl[489] vdd gnd cell_6t
Xbit_r490_c126 bl[126] br[126] wl[490] vdd gnd cell_6t
Xbit_r491_c126 bl[126] br[126] wl[491] vdd gnd cell_6t
Xbit_r492_c126 bl[126] br[126] wl[492] vdd gnd cell_6t
Xbit_r493_c126 bl[126] br[126] wl[493] vdd gnd cell_6t
Xbit_r494_c126 bl[126] br[126] wl[494] vdd gnd cell_6t
Xbit_r495_c126 bl[126] br[126] wl[495] vdd gnd cell_6t
Xbit_r496_c126 bl[126] br[126] wl[496] vdd gnd cell_6t
Xbit_r497_c126 bl[126] br[126] wl[497] vdd gnd cell_6t
Xbit_r498_c126 bl[126] br[126] wl[498] vdd gnd cell_6t
Xbit_r499_c126 bl[126] br[126] wl[499] vdd gnd cell_6t
Xbit_r500_c126 bl[126] br[126] wl[500] vdd gnd cell_6t
Xbit_r501_c126 bl[126] br[126] wl[501] vdd gnd cell_6t
Xbit_r502_c126 bl[126] br[126] wl[502] vdd gnd cell_6t
Xbit_r503_c126 bl[126] br[126] wl[503] vdd gnd cell_6t
Xbit_r504_c126 bl[126] br[126] wl[504] vdd gnd cell_6t
Xbit_r505_c126 bl[126] br[126] wl[505] vdd gnd cell_6t
Xbit_r506_c126 bl[126] br[126] wl[506] vdd gnd cell_6t
Xbit_r507_c126 bl[126] br[126] wl[507] vdd gnd cell_6t
Xbit_r508_c126 bl[126] br[126] wl[508] vdd gnd cell_6t
Xbit_r509_c126 bl[126] br[126] wl[509] vdd gnd cell_6t
Xbit_r510_c126 bl[126] br[126] wl[510] vdd gnd cell_6t
Xbit_r511_c126 bl[126] br[126] wl[511] vdd gnd cell_6t
Xbit_r0_c127 bl[127] br[127] wl[0] vdd gnd cell_6t
Xbit_r1_c127 bl[127] br[127] wl[1] vdd gnd cell_6t
Xbit_r2_c127 bl[127] br[127] wl[2] vdd gnd cell_6t
Xbit_r3_c127 bl[127] br[127] wl[3] vdd gnd cell_6t
Xbit_r4_c127 bl[127] br[127] wl[4] vdd gnd cell_6t
Xbit_r5_c127 bl[127] br[127] wl[5] vdd gnd cell_6t
Xbit_r6_c127 bl[127] br[127] wl[6] vdd gnd cell_6t
Xbit_r7_c127 bl[127] br[127] wl[7] vdd gnd cell_6t
Xbit_r8_c127 bl[127] br[127] wl[8] vdd gnd cell_6t
Xbit_r9_c127 bl[127] br[127] wl[9] vdd gnd cell_6t
Xbit_r10_c127 bl[127] br[127] wl[10] vdd gnd cell_6t
Xbit_r11_c127 bl[127] br[127] wl[11] vdd gnd cell_6t
Xbit_r12_c127 bl[127] br[127] wl[12] vdd gnd cell_6t
Xbit_r13_c127 bl[127] br[127] wl[13] vdd gnd cell_6t
Xbit_r14_c127 bl[127] br[127] wl[14] vdd gnd cell_6t
Xbit_r15_c127 bl[127] br[127] wl[15] vdd gnd cell_6t
Xbit_r16_c127 bl[127] br[127] wl[16] vdd gnd cell_6t
Xbit_r17_c127 bl[127] br[127] wl[17] vdd gnd cell_6t
Xbit_r18_c127 bl[127] br[127] wl[18] vdd gnd cell_6t
Xbit_r19_c127 bl[127] br[127] wl[19] vdd gnd cell_6t
Xbit_r20_c127 bl[127] br[127] wl[20] vdd gnd cell_6t
Xbit_r21_c127 bl[127] br[127] wl[21] vdd gnd cell_6t
Xbit_r22_c127 bl[127] br[127] wl[22] vdd gnd cell_6t
Xbit_r23_c127 bl[127] br[127] wl[23] vdd gnd cell_6t
Xbit_r24_c127 bl[127] br[127] wl[24] vdd gnd cell_6t
Xbit_r25_c127 bl[127] br[127] wl[25] vdd gnd cell_6t
Xbit_r26_c127 bl[127] br[127] wl[26] vdd gnd cell_6t
Xbit_r27_c127 bl[127] br[127] wl[27] vdd gnd cell_6t
Xbit_r28_c127 bl[127] br[127] wl[28] vdd gnd cell_6t
Xbit_r29_c127 bl[127] br[127] wl[29] vdd gnd cell_6t
Xbit_r30_c127 bl[127] br[127] wl[30] vdd gnd cell_6t
Xbit_r31_c127 bl[127] br[127] wl[31] vdd gnd cell_6t
Xbit_r32_c127 bl[127] br[127] wl[32] vdd gnd cell_6t
Xbit_r33_c127 bl[127] br[127] wl[33] vdd gnd cell_6t
Xbit_r34_c127 bl[127] br[127] wl[34] vdd gnd cell_6t
Xbit_r35_c127 bl[127] br[127] wl[35] vdd gnd cell_6t
Xbit_r36_c127 bl[127] br[127] wl[36] vdd gnd cell_6t
Xbit_r37_c127 bl[127] br[127] wl[37] vdd gnd cell_6t
Xbit_r38_c127 bl[127] br[127] wl[38] vdd gnd cell_6t
Xbit_r39_c127 bl[127] br[127] wl[39] vdd gnd cell_6t
Xbit_r40_c127 bl[127] br[127] wl[40] vdd gnd cell_6t
Xbit_r41_c127 bl[127] br[127] wl[41] vdd gnd cell_6t
Xbit_r42_c127 bl[127] br[127] wl[42] vdd gnd cell_6t
Xbit_r43_c127 bl[127] br[127] wl[43] vdd gnd cell_6t
Xbit_r44_c127 bl[127] br[127] wl[44] vdd gnd cell_6t
Xbit_r45_c127 bl[127] br[127] wl[45] vdd gnd cell_6t
Xbit_r46_c127 bl[127] br[127] wl[46] vdd gnd cell_6t
Xbit_r47_c127 bl[127] br[127] wl[47] vdd gnd cell_6t
Xbit_r48_c127 bl[127] br[127] wl[48] vdd gnd cell_6t
Xbit_r49_c127 bl[127] br[127] wl[49] vdd gnd cell_6t
Xbit_r50_c127 bl[127] br[127] wl[50] vdd gnd cell_6t
Xbit_r51_c127 bl[127] br[127] wl[51] vdd gnd cell_6t
Xbit_r52_c127 bl[127] br[127] wl[52] vdd gnd cell_6t
Xbit_r53_c127 bl[127] br[127] wl[53] vdd gnd cell_6t
Xbit_r54_c127 bl[127] br[127] wl[54] vdd gnd cell_6t
Xbit_r55_c127 bl[127] br[127] wl[55] vdd gnd cell_6t
Xbit_r56_c127 bl[127] br[127] wl[56] vdd gnd cell_6t
Xbit_r57_c127 bl[127] br[127] wl[57] vdd gnd cell_6t
Xbit_r58_c127 bl[127] br[127] wl[58] vdd gnd cell_6t
Xbit_r59_c127 bl[127] br[127] wl[59] vdd gnd cell_6t
Xbit_r60_c127 bl[127] br[127] wl[60] vdd gnd cell_6t
Xbit_r61_c127 bl[127] br[127] wl[61] vdd gnd cell_6t
Xbit_r62_c127 bl[127] br[127] wl[62] vdd gnd cell_6t
Xbit_r63_c127 bl[127] br[127] wl[63] vdd gnd cell_6t
Xbit_r64_c127 bl[127] br[127] wl[64] vdd gnd cell_6t
Xbit_r65_c127 bl[127] br[127] wl[65] vdd gnd cell_6t
Xbit_r66_c127 bl[127] br[127] wl[66] vdd gnd cell_6t
Xbit_r67_c127 bl[127] br[127] wl[67] vdd gnd cell_6t
Xbit_r68_c127 bl[127] br[127] wl[68] vdd gnd cell_6t
Xbit_r69_c127 bl[127] br[127] wl[69] vdd gnd cell_6t
Xbit_r70_c127 bl[127] br[127] wl[70] vdd gnd cell_6t
Xbit_r71_c127 bl[127] br[127] wl[71] vdd gnd cell_6t
Xbit_r72_c127 bl[127] br[127] wl[72] vdd gnd cell_6t
Xbit_r73_c127 bl[127] br[127] wl[73] vdd gnd cell_6t
Xbit_r74_c127 bl[127] br[127] wl[74] vdd gnd cell_6t
Xbit_r75_c127 bl[127] br[127] wl[75] vdd gnd cell_6t
Xbit_r76_c127 bl[127] br[127] wl[76] vdd gnd cell_6t
Xbit_r77_c127 bl[127] br[127] wl[77] vdd gnd cell_6t
Xbit_r78_c127 bl[127] br[127] wl[78] vdd gnd cell_6t
Xbit_r79_c127 bl[127] br[127] wl[79] vdd gnd cell_6t
Xbit_r80_c127 bl[127] br[127] wl[80] vdd gnd cell_6t
Xbit_r81_c127 bl[127] br[127] wl[81] vdd gnd cell_6t
Xbit_r82_c127 bl[127] br[127] wl[82] vdd gnd cell_6t
Xbit_r83_c127 bl[127] br[127] wl[83] vdd gnd cell_6t
Xbit_r84_c127 bl[127] br[127] wl[84] vdd gnd cell_6t
Xbit_r85_c127 bl[127] br[127] wl[85] vdd gnd cell_6t
Xbit_r86_c127 bl[127] br[127] wl[86] vdd gnd cell_6t
Xbit_r87_c127 bl[127] br[127] wl[87] vdd gnd cell_6t
Xbit_r88_c127 bl[127] br[127] wl[88] vdd gnd cell_6t
Xbit_r89_c127 bl[127] br[127] wl[89] vdd gnd cell_6t
Xbit_r90_c127 bl[127] br[127] wl[90] vdd gnd cell_6t
Xbit_r91_c127 bl[127] br[127] wl[91] vdd gnd cell_6t
Xbit_r92_c127 bl[127] br[127] wl[92] vdd gnd cell_6t
Xbit_r93_c127 bl[127] br[127] wl[93] vdd gnd cell_6t
Xbit_r94_c127 bl[127] br[127] wl[94] vdd gnd cell_6t
Xbit_r95_c127 bl[127] br[127] wl[95] vdd gnd cell_6t
Xbit_r96_c127 bl[127] br[127] wl[96] vdd gnd cell_6t
Xbit_r97_c127 bl[127] br[127] wl[97] vdd gnd cell_6t
Xbit_r98_c127 bl[127] br[127] wl[98] vdd gnd cell_6t
Xbit_r99_c127 bl[127] br[127] wl[99] vdd gnd cell_6t
Xbit_r100_c127 bl[127] br[127] wl[100] vdd gnd cell_6t
Xbit_r101_c127 bl[127] br[127] wl[101] vdd gnd cell_6t
Xbit_r102_c127 bl[127] br[127] wl[102] vdd gnd cell_6t
Xbit_r103_c127 bl[127] br[127] wl[103] vdd gnd cell_6t
Xbit_r104_c127 bl[127] br[127] wl[104] vdd gnd cell_6t
Xbit_r105_c127 bl[127] br[127] wl[105] vdd gnd cell_6t
Xbit_r106_c127 bl[127] br[127] wl[106] vdd gnd cell_6t
Xbit_r107_c127 bl[127] br[127] wl[107] vdd gnd cell_6t
Xbit_r108_c127 bl[127] br[127] wl[108] vdd gnd cell_6t
Xbit_r109_c127 bl[127] br[127] wl[109] vdd gnd cell_6t
Xbit_r110_c127 bl[127] br[127] wl[110] vdd gnd cell_6t
Xbit_r111_c127 bl[127] br[127] wl[111] vdd gnd cell_6t
Xbit_r112_c127 bl[127] br[127] wl[112] vdd gnd cell_6t
Xbit_r113_c127 bl[127] br[127] wl[113] vdd gnd cell_6t
Xbit_r114_c127 bl[127] br[127] wl[114] vdd gnd cell_6t
Xbit_r115_c127 bl[127] br[127] wl[115] vdd gnd cell_6t
Xbit_r116_c127 bl[127] br[127] wl[116] vdd gnd cell_6t
Xbit_r117_c127 bl[127] br[127] wl[117] vdd gnd cell_6t
Xbit_r118_c127 bl[127] br[127] wl[118] vdd gnd cell_6t
Xbit_r119_c127 bl[127] br[127] wl[119] vdd gnd cell_6t
Xbit_r120_c127 bl[127] br[127] wl[120] vdd gnd cell_6t
Xbit_r121_c127 bl[127] br[127] wl[121] vdd gnd cell_6t
Xbit_r122_c127 bl[127] br[127] wl[122] vdd gnd cell_6t
Xbit_r123_c127 bl[127] br[127] wl[123] vdd gnd cell_6t
Xbit_r124_c127 bl[127] br[127] wl[124] vdd gnd cell_6t
Xbit_r125_c127 bl[127] br[127] wl[125] vdd gnd cell_6t
Xbit_r126_c127 bl[127] br[127] wl[126] vdd gnd cell_6t
Xbit_r127_c127 bl[127] br[127] wl[127] vdd gnd cell_6t
Xbit_r128_c127 bl[127] br[127] wl[128] vdd gnd cell_6t
Xbit_r129_c127 bl[127] br[127] wl[129] vdd gnd cell_6t
Xbit_r130_c127 bl[127] br[127] wl[130] vdd gnd cell_6t
Xbit_r131_c127 bl[127] br[127] wl[131] vdd gnd cell_6t
Xbit_r132_c127 bl[127] br[127] wl[132] vdd gnd cell_6t
Xbit_r133_c127 bl[127] br[127] wl[133] vdd gnd cell_6t
Xbit_r134_c127 bl[127] br[127] wl[134] vdd gnd cell_6t
Xbit_r135_c127 bl[127] br[127] wl[135] vdd gnd cell_6t
Xbit_r136_c127 bl[127] br[127] wl[136] vdd gnd cell_6t
Xbit_r137_c127 bl[127] br[127] wl[137] vdd gnd cell_6t
Xbit_r138_c127 bl[127] br[127] wl[138] vdd gnd cell_6t
Xbit_r139_c127 bl[127] br[127] wl[139] vdd gnd cell_6t
Xbit_r140_c127 bl[127] br[127] wl[140] vdd gnd cell_6t
Xbit_r141_c127 bl[127] br[127] wl[141] vdd gnd cell_6t
Xbit_r142_c127 bl[127] br[127] wl[142] vdd gnd cell_6t
Xbit_r143_c127 bl[127] br[127] wl[143] vdd gnd cell_6t
Xbit_r144_c127 bl[127] br[127] wl[144] vdd gnd cell_6t
Xbit_r145_c127 bl[127] br[127] wl[145] vdd gnd cell_6t
Xbit_r146_c127 bl[127] br[127] wl[146] vdd gnd cell_6t
Xbit_r147_c127 bl[127] br[127] wl[147] vdd gnd cell_6t
Xbit_r148_c127 bl[127] br[127] wl[148] vdd gnd cell_6t
Xbit_r149_c127 bl[127] br[127] wl[149] vdd gnd cell_6t
Xbit_r150_c127 bl[127] br[127] wl[150] vdd gnd cell_6t
Xbit_r151_c127 bl[127] br[127] wl[151] vdd gnd cell_6t
Xbit_r152_c127 bl[127] br[127] wl[152] vdd gnd cell_6t
Xbit_r153_c127 bl[127] br[127] wl[153] vdd gnd cell_6t
Xbit_r154_c127 bl[127] br[127] wl[154] vdd gnd cell_6t
Xbit_r155_c127 bl[127] br[127] wl[155] vdd gnd cell_6t
Xbit_r156_c127 bl[127] br[127] wl[156] vdd gnd cell_6t
Xbit_r157_c127 bl[127] br[127] wl[157] vdd gnd cell_6t
Xbit_r158_c127 bl[127] br[127] wl[158] vdd gnd cell_6t
Xbit_r159_c127 bl[127] br[127] wl[159] vdd gnd cell_6t
Xbit_r160_c127 bl[127] br[127] wl[160] vdd gnd cell_6t
Xbit_r161_c127 bl[127] br[127] wl[161] vdd gnd cell_6t
Xbit_r162_c127 bl[127] br[127] wl[162] vdd gnd cell_6t
Xbit_r163_c127 bl[127] br[127] wl[163] vdd gnd cell_6t
Xbit_r164_c127 bl[127] br[127] wl[164] vdd gnd cell_6t
Xbit_r165_c127 bl[127] br[127] wl[165] vdd gnd cell_6t
Xbit_r166_c127 bl[127] br[127] wl[166] vdd gnd cell_6t
Xbit_r167_c127 bl[127] br[127] wl[167] vdd gnd cell_6t
Xbit_r168_c127 bl[127] br[127] wl[168] vdd gnd cell_6t
Xbit_r169_c127 bl[127] br[127] wl[169] vdd gnd cell_6t
Xbit_r170_c127 bl[127] br[127] wl[170] vdd gnd cell_6t
Xbit_r171_c127 bl[127] br[127] wl[171] vdd gnd cell_6t
Xbit_r172_c127 bl[127] br[127] wl[172] vdd gnd cell_6t
Xbit_r173_c127 bl[127] br[127] wl[173] vdd gnd cell_6t
Xbit_r174_c127 bl[127] br[127] wl[174] vdd gnd cell_6t
Xbit_r175_c127 bl[127] br[127] wl[175] vdd gnd cell_6t
Xbit_r176_c127 bl[127] br[127] wl[176] vdd gnd cell_6t
Xbit_r177_c127 bl[127] br[127] wl[177] vdd gnd cell_6t
Xbit_r178_c127 bl[127] br[127] wl[178] vdd gnd cell_6t
Xbit_r179_c127 bl[127] br[127] wl[179] vdd gnd cell_6t
Xbit_r180_c127 bl[127] br[127] wl[180] vdd gnd cell_6t
Xbit_r181_c127 bl[127] br[127] wl[181] vdd gnd cell_6t
Xbit_r182_c127 bl[127] br[127] wl[182] vdd gnd cell_6t
Xbit_r183_c127 bl[127] br[127] wl[183] vdd gnd cell_6t
Xbit_r184_c127 bl[127] br[127] wl[184] vdd gnd cell_6t
Xbit_r185_c127 bl[127] br[127] wl[185] vdd gnd cell_6t
Xbit_r186_c127 bl[127] br[127] wl[186] vdd gnd cell_6t
Xbit_r187_c127 bl[127] br[127] wl[187] vdd gnd cell_6t
Xbit_r188_c127 bl[127] br[127] wl[188] vdd gnd cell_6t
Xbit_r189_c127 bl[127] br[127] wl[189] vdd gnd cell_6t
Xbit_r190_c127 bl[127] br[127] wl[190] vdd gnd cell_6t
Xbit_r191_c127 bl[127] br[127] wl[191] vdd gnd cell_6t
Xbit_r192_c127 bl[127] br[127] wl[192] vdd gnd cell_6t
Xbit_r193_c127 bl[127] br[127] wl[193] vdd gnd cell_6t
Xbit_r194_c127 bl[127] br[127] wl[194] vdd gnd cell_6t
Xbit_r195_c127 bl[127] br[127] wl[195] vdd gnd cell_6t
Xbit_r196_c127 bl[127] br[127] wl[196] vdd gnd cell_6t
Xbit_r197_c127 bl[127] br[127] wl[197] vdd gnd cell_6t
Xbit_r198_c127 bl[127] br[127] wl[198] vdd gnd cell_6t
Xbit_r199_c127 bl[127] br[127] wl[199] vdd gnd cell_6t
Xbit_r200_c127 bl[127] br[127] wl[200] vdd gnd cell_6t
Xbit_r201_c127 bl[127] br[127] wl[201] vdd gnd cell_6t
Xbit_r202_c127 bl[127] br[127] wl[202] vdd gnd cell_6t
Xbit_r203_c127 bl[127] br[127] wl[203] vdd gnd cell_6t
Xbit_r204_c127 bl[127] br[127] wl[204] vdd gnd cell_6t
Xbit_r205_c127 bl[127] br[127] wl[205] vdd gnd cell_6t
Xbit_r206_c127 bl[127] br[127] wl[206] vdd gnd cell_6t
Xbit_r207_c127 bl[127] br[127] wl[207] vdd gnd cell_6t
Xbit_r208_c127 bl[127] br[127] wl[208] vdd gnd cell_6t
Xbit_r209_c127 bl[127] br[127] wl[209] vdd gnd cell_6t
Xbit_r210_c127 bl[127] br[127] wl[210] vdd gnd cell_6t
Xbit_r211_c127 bl[127] br[127] wl[211] vdd gnd cell_6t
Xbit_r212_c127 bl[127] br[127] wl[212] vdd gnd cell_6t
Xbit_r213_c127 bl[127] br[127] wl[213] vdd gnd cell_6t
Xbit_r214_c127 bl[127] br[127] wl[214] vdd gnd cell_6t
Xbit_r215_c127 bl[127] br[127] wl[215] vdd gnd cell_6t
Xbit_r216_c127 bl[127] br[127] wl[216] vdd gnd cell_6t
Xbit_r217_c127 bl[127] br[127] wl[217] vdd gnd cell_6t
Xbit_r218_c127 bl[127] br[127] wl[218] vdd gnd cell_6t
Xbit_r219_c127 bl[127] br[127] wl[219] vdd gnd cell_6t
Xbit_r220_c127 bl[127] br[127] wl[220] vdd gnd cell_6t
Xbit_r221_c127 bl[127] br[127] wl[221] vdd gnd cell_6t
Xbit_r222_c127 bl[127] br[127] wl[222] vdd gnd cell_6t
Xbit_r223_c127 bl[127] br[127] wl[223] vdd gnd cell_6t
Xbit_r224_c127 bl[127] br[127] wl[224] vdd gnd cell_6t
Xbit_r225_c127 bl[127] br[127] wl[225] vdd gnd cell_6t
Xbit_r226_c127 bl[127] br[127] wl[226] vdd gnd cell_6t
Xbit_r227_c127 bl[127] br[127] wl[227] vdd gnd cell_6t
Xbit_r228_c127 bl[127] br[127] wl[228] vdd gnd cell_6t
Xbit_r229_c127 bl[127] br[127] wl[229] vdd gnd cell_6t
Xbit_r230_c127 bl[127] br[127] wl[230] vdd gnd cell_6t
Xbit_r231_c127 bl[127] br[127] wl[231] vdd gnd cell_6t
Xbit_r232_c127 bl[127] br[127] wl[232] vdd gnd cell_6t
Xbit_r233_c127 bl[127] br[127] wl[233] vdd gnd cell_6t
Xbit_r234_c127 bl[127] br[127] wl[234] vdd gnd cell_6t
Xbit_r235_c127 bl[127] br[127] wl[235] vdd gnd cell_6t
Xbit_r236_c127 bl[127] br[127] wl[236] vdd gnd cell_6t
Xbit_r237_c127 bl[127] br[127] wl[237] vdd gnd cell_6t
Xbit_r238_c127 bl[127] br[127] wl[238] vdd gnd cell_6t
Xbit_r239_c127 bl[127] br[127] wl[239] vdd gnd cell_6t
Xbit_r240_c127 bl[127] br[127] wl[240] vdd gnd cell_6t
Xbit_r241_c127 bl[127] br[127] wl[241] vdd gnd cell_6t
Xbit_r242_c127 bl[127] br[127] wl[242] vdd gnd cell_6t
Xbit_r243_c127 bl[127] br[127] wl[243] vdd gnd cell_6t
Xbit_r244_c127 bl[127] br[127] wl[244] vdd gnd cell_6t
Xbit_r245_c127 bl[127] br[127] wl[245] vdd gnd cell_6t
Xbit_r246_c127 bl[127] br[127] wl[246] vdd gnd cell_6t
Xbit_r247_c127 bl[127] br[127] wl[247] vdd gnd cell_6t
Xbit_r248_c127 bl[127] br[127] wl[248] vdd gnd cell_6t
Xbit_r249_c127 bl[127] br[127] wl[249] vdd gnd cell_6t
Xbit_r250_c127 bl[127] br[127] wl[250] vdd gnd cell_6t
Xbit_r251_c127 bl[127] br[127] wl[251] vdd gnd cell_6t
Xbit_r252_c127 bl[127] br[127] wl[252] vdd gnd cell_6t
Xbit_r253_c127 bl[127] br[127] wl[253] vdd gnd cell_6t
Xbit_r254_c127 bl[127] br[127] wl[254] vdd gnd cell_6t
Xbit_r255_c127 bl[127] br[127] wl[255] vdd gnd cell_6t
Xbit_r256_c127 bl[127] br[127] wl[256] vdd gnd cell_6t
Xbit_r257_c127 bl[127] br[127] wl[257] vdd gnd cell_6t
Xbit_r258_c127 bl[127] br[127] wl[258] vdd gnd cell_6t
Xbit_r259_c127 bl[127] br[127] wl[259] vdd gnd cell_6t
Xbit_r260_c127 bl[127] br[127] wl[260] vdd gnd cell_6t
Xbit_r261_c127 bl[127] br[127] wl[261] vdd gnd cell_6t
Xbit_r262_c127 bl[127] br[127] wl[262] vdd gnd cell_6t
Xbit_r263_c127 bl[127] br[127] wl[263] vdd gnd cell_6t
Xbit_r264_c127 bl[127] br[127] wl[264] vdd gnd cell_6t
Xbit_r265_c127 bl[127] br[127] wl[265] vdd gnd cell_6t
Xbit_r266_c127 bl[127] br[127] wl[266] vdd gnd cell_6t
Xbit_r267_c127 bl[127] br[127] wl[267] vdd gnd cell_6t
Xbit_r268_c127 bl[127] br[127] wl[268] vdd gnd cell_6t
Xbit_r269_c127 bl[127] br[127] wl[269] vdd gnd cell_6t
Xbit_r270_c127 bl[127] br[127] wl[270] vdd gnd cell_6t
Xbit_r271_c127 bl[127] br[127] wl[271] vdd gnd cell_6t
Xbit_r272_c127 bl[127] br[127] wl[272] vdd gnd cell_6t
Xbit_r273_c127 bl[127] br[127] wl[273] vdd gnd cell_6t
Xbit_r274_c127 bl[127] br[127] wl[274] vdd gnd cell_6t
Xbit_r275_c127 bl[127] br[127] wl[275] vdd gnd cell_6t
Xbit_r276_c127 bl[127] br[127] wl[276] vdd gnd cell_6t
Xbit_r277_c127 bl[127] br[127] wl[277] vdd gnd cell_6t
Xbit_r278_c127 bl[127] br[127] wl[278] vdd gnd cell_6t
Xbit_r279_c127 bl[127] br[127] wl[279] vdd gnd cell_6t
Xbit_r280_c127 bl[127] br[127] wl[280] vdd gnd cell_6t
Xbit_r281_c127 bl[127] br[127] wl[281] vdd gnd cell_6t
Xbit_r282_c127 bl[127] br[127] wl[282] vdd gnd cell_6t
Xbit_r283_c127 bl[127] br[127] wl[283] vdd gnd cell_6t
Xbit_r284_c127 bl[127] br[127] wl[284] vdd gnd cell_6t
Xbit_r285_c127 bl[127] br[127] wl[285] vdd gnd cell_6t
Xbit_r286_c127 bl[127] br[127] wl[286] vdd gnd cell_6t
Xbit_r287_c127 bl[127] br[127] wl[287] vdd gnd cell_6t
Xbit_r288_c127 bl[127] br[127] wl[288] vdd gnd cell_6t
Xbit_r289_c127 bl[127] br[127] wl[289] vdd gnd cell_6t
Xbit_r290_c127 bl[127] br[127] wl[290] vdd gnd cell_6t
Xbit_r291_c127 bl[127] br[127] wl[291] vdd gnd cell_6t
Xbit_r292_c127 bl[127] br[127] wl[292] vdd gnd cell_6t
Xbit_r293_c127 bl[127] br[127] wl[293] vdd gnd cell_6t
Xbit_r294_c127 bl[127] br[127] wl[294] vdd gnd cell_6t
Xbit_r295_c127 bl[127] br[127] wl[295] vdd gnd cell_6t
Xbit_r296_c127 bl[127] br[127] wl[296] vdd gnd cell_6t
Xbit_r297_c127 bl[127] br[127] wl[297] vdd gnd cell_6t
Xbit_r298_c127 bl[127] br[127] wl[298] vdd gnd cell_6t
Xbit_r299_c127 bl[127] br[127] wl[299] vdd gnd cell_6t
Xbit_r300_c127 bl[127] br[127] wl[300] vdd gnd cell_6t
Xbit_r301_c127 bl[127] br[127] wl[301] vdd gnd cell_6t
Xbit_r302_c127 bl[127] br[127] wl[302] vdd gnd cell_6t
Xbit_r303_c127 bl[127] br[127] wl[303] vdd gnd cell_6t
Xbit_r304_c127 bl[127] br[127] wl[304] vdd gnd cell_6t
Xbit_r305_c127 bl[127] br[127] wl[305] vdd gnd cell_6t
Xbit_r306_c127 bl[127] br[127] wl[306] vdd gnd cell_6t
Xbit_r307_c127 bl[127] br[127] wl[307] vdd gnd cell_6t
Xbit_r308_c127 bl[127] br[127] wl[308] vdd gnd cell_6t
Xbit_r309_c127 bl[127] br[127] wl[309] vdd gnd cell_6t
Xbit_r310_c127 bl[127] br[127] wl[310] vdd gnd cell_6t
Xbit_r311_c127 bl[127] br[127] wl[311] vdd gnd cell_6t
Xbit_r312_c127 bl[127] br[127] wl[312] vdd gnd cell_6t
Xbit_r313_c127 bl[127] br[127] wl[313] vdd gnd cell_6t
Xbit_r314_c127 bl[127] br[127] wl[314] vdd gnd cell_6t
Xbit_r315_c127 bl[127] br[127] wl[315] vdd gnd cell_6t
Xbit_r316_c127 bl[127] br[127] wl[316] vdd gnd cell_6t
Xbit_r317_c127 bl[127] br[127] wl[317] vdd gnd cell_6t
Xbit_r318_c127 bl[127] br[127] wl[318] vdd gnd cell_6t
Xbit_r319_c127 bl[127] br[127] wl[319] vdd gnd cell_6t
Xbit_r320_c127 bl[127] br[127] wl[320] vdd gnd cell_6t
Xbit_r321_c127 bl[127] br[127] wl[321] vdd gnd cell_6t
Xbit_r322_c127 bl[127] br[127] wl[322] vdd gnd cell_6t
Xbit_r323_c127 bl[127] br[127] wl[323] vdd gnd cell_6t
Xbit_r324_c127 bl[127] br[127] wl[324] vdd gnd cell_6t
Xbit_r325_c127 bl[127] br[127] wl[325] vdd gnd cell_6t
Xbit_r326_c127 bl[127] br[127] wl[326] vdd gnd cell_6t
Xbit_r327_c127 bl[127] br[127] wl[327] vdd gnd cell_6t
Xbit_r328_c127 bl[127] br[127] wl[328] vdd gnd cell_6t
Xbit_r329_c127 bl[127] br[127] wl[329] vdd gnd cell_6t
Xbit_r330_c127 bl[127] br[127] wl[330] vdd gnd cell_6t
Xbit_r331_c127 bl[127] br[127] wl[331] vdd gnd cell_6t
Xbit_r332_c127 bl[127] br[127] wl[332] vdd gnd cell_6t
Xbit_r333_c127 bl[127] br[127] wl[333] vdd gnd cell_6t
Xbit_r334_c127 bl[127] br[127] wl[334] vdd gnd cell_6t
Xbit_r335_c127 bl[127] br[127] wl[335] vdd gnd cell_6t
Xbit_r336_c127 bl[127] br[127] wl[336] vdd gnd cell_6t
Xbit_r337_c127 bl[127] br[127] wl[337] vdd gnd cell_6t
Xbit_r338_c127 bl[127] br[127] wl[338] vdd gnd cell_6t
Xbit_r339_c127 bl[127] br[127] wl[339] vdd gnd cell_6t
Xbit_r340_c127 bl[127] br[127] wl[340] vdd gnd cell_6t
Xbit_r341_c127 bl[127] br[127] wl[341] vdd gnd cell_6t
Xbit_r342_c127 bl[127] br[127] wl[342] vdd gnd cell_6t
Xbit_r343_c127 bl[127] br[127] wl[343] vdd gnd cell_6t
Xbit_r344_c127 bl[127] br[127] wl[344] vdd gnd cell_6t
Xbit_r345_c127 bl[127] br[127] wl[345] vdd gnd cell_6t
Xbit_r346_c127 bl[127] br[127] wl[346] vdd gnd cell_6t
Xbit_r347_c127 bl[127] br[127] wl[347] vdd gnd cell_6t
Xbit_r348_c127 bl[127] br[127] wl[348] vdd gnd cell_6t
Xbit_r349_c127 bl[127] br[127] wl[349] vdd gnd cell_6t
Xbit_r350_c127 bl[127] br[127] wl[350] vdd gnd cell_6t
Xbit_r351_c127 bl[127] br[127] wl[351] vdd gnd cell_6t
Xbit_r352_c127 bl[127] br[127] wl[352] vdd gnd cell_6t
Xbit_r353_c127 bl[127] br[127] wl[353] vdd gnd cell_6t
Xbit_r354_c127 bl[127] br[127] wl[354] vdd gnd cell_6t
Xbit_r355_c127 bl[127] br[127] wl[355] vdd gnd cell_6t
Xbit_r356_c127 bl[127] br[127] wl[356] vdd gnd cell_6t
Xbit_r357_c127 bl[127] br[127] wl[357] vdd gnd cell_6t
Xbit_r358_c127 bl[127] br[127] wl[358] vdd gnd cell_6t
Xbit_r359_c127 bl[127] br[127] wl[359] vdd gnd cell_6t
Xbit_r360_c127 bl[127] br[127] wl[360] vdd gnd cell_6t
Xbit_r361_c127 bl[127] br[127] wl[361] vdd gnd cell_6t
Xbit_r362_c127 bl[127] br[127] wl[362] vdd gnd cell_6t
Xbit_r363_c127 bl[127] br[127] wl[363] vdd gnd cell_6t
Xbit_r364_c127 bl[127] br[127] wl[364] vdd gnd cell_6t
Xbit_r365_c127 bl[127] br[127] wl[365] vdd gnd cell_6t
Xbit_r366_c127 bl[127] br[127] wl[366] vdd gnd cell_6t
Xbit_r367_c127 bl[127] br[127] wl[367] vdd gnd cell_6t
Xbit_r368_c127 bl[127] br[127] wl[368] vdd gnd cell_6t
Xbit_r369_c127 bl[127] br[127] wl[369] vdd gnd cell_6t
Xbit_r370_c127 bl[127] br[127] wl[370] vdd gnd cell_6t
Xbit_r371_c127 bl[127] br[127] wl[371] vdd gnd cell_6t
Xbit_r372_c127 bl[127] br[127] wl[372] vdd gnd cell_6t
Xbit_r373_c127 bl[127] br[127] wl[373] vdd gnd cell_6t
Xbit_r374_c127 bl[127] br[127] wl[374] vdd gnd cell_6t
Xbit_r375_c127 bl[127] br[127] wl[375] vdd gnd cell_6t
Xbit_r376_c127 bl[127] br[127] wl[376] vdd gnd cell_6t
Xbit_r377_c127 bl[127] br[127] wl[377] vdd gnd cell_6t
Xbit_r378_c127 bl[127] br[127] wl[378] vdd gnd cell_6t
Xbit_r379_c127 bl[127] br[127] wl[379] vdd gnd cell_6t
Xbit_r380_c127 bl[127] br[127] wl[380] vdd gnd cell_6t
Xbit_r381_c127 bl[127] br[127] wl[381] vdd gnd cell_6t
Xbit_r382_c127 bl[127] br[127] wl[382] vdd gnd cell_6t
Xbit_r383_c127 bl[127] br[127] wl[383] vdd gnd cell_6t
Xbit_r384_c127 bl[127] br[127] wl[384] vdd gnd cell_6t
Xbit_r385_c127 bl[127] br[127] wl[385] vdd gnd cell_6t
Xbit_r386_c127 bl[127] br[127] wl[386] vdd gnd cell_6t
Xbit_r387_c127 bl[127] br[127] wl[387] vdd gnd cell_6t
Xbit_r388_c127 bl[127] br[127] wl[388] vdd gnd cell_6t
Xbit_r389_c127 bl[127] br[127] wl[389] vdd gnd cell_6t
Xbit_r390_c127 bl[127] br[127] wl[390] vdd gnd cell_6t
Xbit_r391_c127 bl[127] br[127] wl[391] vdd gnd cell_6t
Xbit_r392_c127 bl[127] br[127] wl[392] vdd gnd cell_6t
Xbit_r393_c127 bl[127] br[127] wl[393] vdd gnd cell_6t
Xbit_r394_c127 bl[127] br[127] wl[394] vdd gnd cell_6t
Xbit_r395_c127 bl[127] br[127] wl[395] vdd gnd cell_6t
Xbit_r396_c127 bl[127] br[127] wl[396] vdd gnd cell_6t
Xbit_r397_c127 bl[127] br[127] wl[397] vdd gnd cell_6t
Xbit_r398_c127 bl[127] br[127] wl[398] vdd gnd cell_6t
Xbit_r399_c127 bl[127] br[127] wl[399] vdd gnd cell_6t
Xbit_r400_c127 bl[127] br[127] wl[400] vdd gnd cell_6t
Xbit_r401_c127 bl[127] br[127] wl[401] vdd gnd cell_6t
Xbit_r402_c127 bl[127] br[127] wl[402] vdd gnd cell_6t
Xbit_r403_c127 bl[127] br[127] wl[403] vdd gnd cell_6t
Xbit_r404_c127 bl[127] br[127] wl[404] vdd gnd cell_6t
Xbit_r405_c127 bl[127] br[127] wl[405] vdd gnd cell_6t
Xbit_r406_c127 bl[127] br[127] wl[406] vdd gnd cell_6t
Xbit_r407_c127 bl[127] br[127] wl[407] vdd gnd cell_6t
Xbit_r408_c127 bl[127] br[127] wl[408] vdd gnd cell_6t
Xbit_r409_c127 bl[127] br[127] wl[409] vdd gnd cell_6t
Xbit_r410_c127 bl[127] br[127] wl[410] vdd gnd cell_6t
Xbit_r411_c127 bl[127] br[127] wl[411] vdd gnd cell_6t
Xbit_r412_c127 bl[127] br[127] wl[412] vdd gnd cell_6t
Xbit_r413_c127 bl[127] br[127] wl[413] vdd gnd cell_6t
Xbit_r414_c127 bl[127] br[127] wl[414] vdd gnd cell_6t
Xbit_r415_c127 bl[127] br[127] wl[415] vdd gnd cell_6t
Xbit_r416_c127 bl[127] br[127] wl[416] vdd gnd cell_6t
Xbit_r417_c127 bl[127] br[127] wl[417] vdd gnd cell_6t
Xbit_r418_c127 bl[127] br[127] wl[418] vdd gnd cell_6t
Xbit_r419_c127 bl[127] br[127] wl[419] vdd gnd cell_6t
Xbit_r420_c127 bl[127] br[127] wl[420] vdd gnd cell_6t
Xbit_r421_c127 bl[127] br[127] wl[421] vdd gnd cell_6t
Xbit_r422_c127 bl[127] br[127] wl[422] vdd gnd cell_6t
Xbit_r423_c127 bl[127] br[127] wl[423] vdd gnd cell_6t
Xbit_r424_c127 bl[127] br[127] wl[424] vdd gnd cell_6t
Xbit_r425_c127 bl[127] br[127] wl[425] vdd gnd cell_6t
Xbit_r426_c127 bl[127] br[127] wl[426] vdd gnd cell_6t
Xbit_r427_c127 bl[127] br[127] wl[427] vdd gnd cell_6t
Xbit_r428_c127 bl[127] br[127] wl[428] vdd gnd cell_6t
Xbit_r429_c127 bl[127] br[127] wl[429] vdd gnd cell_6t
Xbit_r430_c127 bl[127] br[127] wl[430] vdd gnd cell_6t
Xbit_r431_c127 bl[127] br[127] wl[431] vdd gnd cell_6t
Xbit_r432_c127 bl[127] br[127] wl[432] vdd gnd cell_6t
Xbit_r433_c127 bl[127] br[127] wl[433] vdd gnd cell_6t
Xbit_r434_c127 bl[127] br[127] wl[434] vdd gnd cell_6t
Xbit_r435_c127 bl[127] br[127] wl[435] vdd gnd cell_6t
Xbit_r436_c127 bl[127] br[127] wl[436] vdd gnd cell_6t
Xbit_r437_c127 bl[127] br[127] wl[437] vdd gnd cell_6t
Xbit_r438_c127 bl[127] br[127] wl[438] vdd gnd cell_6t
Xbit_r439_c127 bl[127] br[127] wl[439] vdd gnd cell_6t
Xbit_r440_c127 bl[127] br[127] wl[440] vdd gnd cell_6t
Xbit_r441_c127 bl[127] br[127] wl[441] vdd gnd cell_6t
Xbit_r442_c127 bl[127] br[127] wl[442] vdd gnd cell_6t
Xbit_r443_c127 bl[127] br[127] wl[443] vdd gnd cell_6t
Xbit_r444_c127 bl[127] br[127] wl[444] vdd gnd cell_6t
Xbit_r445_c127 bl[127] br[127] wl[445] vdd gnd cell_6t
Xbit_r446_c127 bl[127] br[127] wl[446] vdd gnd cell_6t
Xbit_r447_c127 bl[127] br[127] wl[447] vdd gnd cell_6t
Xbit_r448_c127 bl[127] br[127] wl[448] vdd gnd cell_6t
Xbit_r449_c127 bl[127] br[127] wl[449] vdd gnd cell_6t
Xbit_r450_c127 bl[127] br[127] wl[450] vdd gnd cell_6t
Xbit_r451_c127 bl[127] br[127] wl[451] vdd gnd cell_6t
Xbit_r452_c127 bl[127] br[127] wl[452] vdd gnd cell_6t
Xbit_r453_c127 bl[127] br[127] wl[453] vdd gnd cell_6t
Xbit_r454_c127 bl[127] br[127] wl[454] vdd gnd cell_6t
Xbit_r455_c127 bl[127] br[127] wl[455] vdd gnd cell_6t
Xbit_r456_c127 bl[127] br[127] wl[456] vdd gnd cell_6t
Xbit_r457_c127 bl[127] br[127] wl[457] vdd gnd cell_6t
Xbit_r458_c127 bl[127] br[127] wl[458] vdd gnd cell_6t
Xbit_r459_c127 bl[127] br[127] wl[459] vdd gnd cell_6t
Xbit_r460_c127 bl[127] br[127] wl[460] vdd gnd cell_6t
Xbit_r461_c127 bl[127] br[127] wl[461] vdd gnd cell_6t
Xbit_r462_c127 bl[127] br[127] wl[462] vdd gnd cell_6t
Xbit_r463_c127 bl[127] br[127] wl[463] vdd gnd cell_6t
Xbit_r464_c127 bl[127] br[127] wl[464] vdd gnd cell_6t
Xbit_r465_c127 bl[127] br[127] wl[465] vdd gnd cell_6t
Xbit_r466_c127 bl[127] br[127] wl[466] vdd gnd cell_6t
Xbit_r467_c127 bl[127] br[127] wl[467] vdd gnd cell_6t
Xbit_r468_c127 bl[127] br[127] wl[468] vdd gnd cell_6t
Xbit_r469_c127 bl[127] br[127] wl[469] vdd gnd cell_6t
Xbit_r470_c127 bl[127] br[127] wl[470] vdd gnd cell_6t
Xbit_r471_c127 bl[127] br[127] wl[471] vdd gnd cell_6t
Xbit_r472_c127 bl[127] br[127] wl[472] vdd gnd cell_6t
Xbit_r473_c127 bl[127] br[127] wl[473] vdd gnd cell_6t
Xbit_r474_c127 bl[127] br[127] wl[474] vdd gnd cell_6t
Xbit_r475_c127 bl[127] br[127] wl[475] vdd gnd cell_6t
Xbit_r476_c127 bl[127] br[127] wl[476] vdd gnd cell_6t
Xbit_r477_c127 bl[127] br[127] wl[477] vdd gnd cell_6t
Xbit_r478_c127 bl[127] br[127] wl[478] vdd gnd cell_6t
Xbit_r479_c127 bl[127] br[127] wl[479] vdd gnd cell_6t
Xbit_r480_c127 bl[127] br[127] wl[480] vdd gnd cell_6t
Xbit_r481_c127 bl[127] br[127] wl[481] vdd gnd cell_6t
Xbit_r482_c127 bl[127] br[127] wl[482] vdd gnd cell_6t
Xbit_r483_c127 bl[127] br[127] wl[483] vdd gnd cell_6t
Xbit_r484_c127 bl[127] br[127] wl[484] vdd gnd cell_6t
Xbit_r485_c127 bl[127] br[127] wl[485] vdd gnd cell_6t
Xbit_r486_c127 bl[127] br[127] wl[486] vdd gnd cell_6t
Xbit_r487_c127 bl[127] br[127] wl[487] vdd gnd cell_6t
Xbit_r488_c127 bl[127] br[127] wl[488] vdd gnd cell_6t
Xbit_r489_c127 bl[127] br[127] wl[489] vdd gnd cell_6t
Xbit_r490_c127 bl[127] br[127] wl[490] vdd gnd cell_6t
Xbit_r491_c127 bl[127] br[127] wl[491] vdd gnd cell_6t
Xbit_r492_c127 bl[127] br[127] wl[492] vdd gnd cell_6t
Xbit_r493_c127 bl[127] br[127] wl[493] vdd gnd cell_6t
Xbit_r494_c127 bl[127] br[127] wl[494] vdd gnd cell_6t
Xbit_r495_c127 bl[127] br[127] wl[495] vdd gnd cell_6t
Xbit_r496_c127 bl[127] br[127] wl[496] vdd gnd cell_6t
Xbit_r497_c127 bl[127] br[127] wl[497] vdd gnd cell_6t
Xbit_r498_c127 bl[127] br[127] wl[498] vdd gnd cell_6t
Xbit_r499_c127 bl[127] br[127] wl[499] vdd gnd cell_6t
Xbit_r500_c127 bl[127] br[127] wl[500] vdd gnd cell_6t
Xbit_r501_c127 bl[127] br[127] wl[501] vdd gnd cell_6t
Xbit_r502_c127 bl[127] br[127] wl[502] vdd gnd cell_6t
Xbit_r503_c127 bl[127] br[127] wl[503] vdd gnd cell_6t
Xbit_r504_c127 bl[127] br[127] wl[504] vdd gnd cell_6t
Xbit_r505_c127 bl[127] br[127] wl[505] vdd gnd cell_6t
Xbit_r506_c127 bl[127] br[127] wl[506] vdd gnd cell_6t
Xbit_r507_c127 bl[127] br[127] wl[507] vdd gnd cell_6t
Xbit_r508_c127 bl[127] br[127] wl[508] vdd gnd cell_6t
Xbit_r509_c127 bl[127] br[127] wl[509] vdd gnd cell_6t
Xbit_r510_c127 bl[127] br[127] wl[510] vdd gnd cell_6t
Xbit_r511_c127 bl[127] br[127] wl[511] vdd gnd cell_6t
.ENDS bitcell_array

* ptx M{0} {1} pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p

.SUBCKT precharge bl br en vdd
Mlower_pmos bl en BR vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mupper_pmos1 bl en vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mupper_pmos2 br en vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
.ENDS precharge

.SUBCKT precharge_array bl[0] br[0] bl[1] br[1] bl[2] br[2] bl[3] br[3] bl[4] br[4] bl[5] br[5] bl[6] br[6] bl[7] br[7] bl[8] br[8] bl[9] br[9] bl[10] br[10] bl[11] br[11] bl[12] br[12] bl[13] br[13] bl[14] br[14] bl[15] br[15] bl[16] br[16] bl[17] br[17] bl[18] br[18] bl[19] br[19] bl[20] br[20] bl[21] br[21] bl[22] br[22] bl[23] br[23] bl[24] br[24] bl[25] br[25] bl[26] br[26] bl[27] br[27] bl[28] br[28] bl[29] br[29] bl[30] br[30] bl[31] br[31] bl[32] br[32] bl[33] br[33] bl[34] br[34] bl[35] br[35] bl[36] br[36] bl[37] br[37] bl[38] br[38] bl[39] br[39] bl[40] br[40] bl[41] br[41] bl[42] br[42] bl[43] br[43] bl[44] br[44] bl[45] br[45] bl[46] br[46] bl[47] br[47] bl[48] br[48] bl[49] br[49] bl[50] br[50] bl[51] br[51] bl[52] br[52] bl[53] br[53] bl[54] br[54] bl[55] br[55] bl[56] br[56] bl[57] br[57] bl[58] br[58] bl[59] br[59] bl[60] br[60] bl[61] br[61] bl[62] br[62] bl[63] br[63] bl[64] br[64] bl[65] br[65] bl[66] br[66] bl[67] br[67] bl[68] br[68] bl[69] br[69] bl[70] br[70] bl[71] br[71] bl[72] br[72] bl[73] br[73] bl[74] br[74] bl[75] br[75] bl[76] br[76] bl[77] br[77] bl[78] br[78] bl[79] br[79] bl[80] br[80] bl[81] br[81] bl[82] br[82] bl[83] br[83] bl[84] br[84] bl[85] br[85] bl[86] br[86] bl[87] br[87] bl[88] br[88] bl[89] br[89] bl[90] br[90] bl[91] br[91] bl[92] br[92] bl[93] br[93] bl[94] br[94] bl[95] br[95] bl[96] br[96] bl[97] br[97] bl[98] br[98] bl[99] br[99] bl[100] br[100] bl[101] br[101] bl[102] br[102] bl[103] br[103] bl[104] br[104] bl[105] br[105] bl[106] br[106] bl[107] br[107] bl[108] br[108] bl[109] br[109] bl[110] br[110] bl[111] br[111] bl[112] br[112] bl[113] br[113] bl[114] br[114] bl[115] br[115] bl[116] br[116] bl[117] br[117] bl[118] br[118] bl[119] br[119] bl[120] br[120] bl[121] br[121] bl[122] br[122] bl[123] br[123] bl[124] br[124] bl[125] br[125] bl[126] br[126] bl[127] br[127] en vdd
Xpre_column_0 bl[0] br[0] en vdd precharge
Xpre_column_1 bl[1] br[1] en vdd precharge
Xpre_column_2 bl[2] br[2] en vdd precharge
Xpre_column_3 bl[3] br[3] en vdd precharge
Xpre_column_4 bl[4] br[4] en vdd precharge
Xpre_column_5 bl[5] br[5] en vdd precharge
Xpre_column_6 bl[6] br[6] en vdd precharge
Xpre_column_7 bl[7] br[7] en vdd precharge
Xpre_column_8 bl[8] br[8] en vdd precharge
Xpre_column_9 bl[9] br[9] en vdd precharge
Xpre_column_10 bl[10] br[10] en vdd precharge
Xpre_column_11 bl[11] br[11] en vdd precharge
Xpre_column_12 bl[12] br[12] en vdd precharge
Xpre_column_13 bl[13] br[13] en vdd precharge
Xpre_column_14 bl[14] br[14] en vdd precharge
Xpre_column_15 bl[15] br[15] en vdd precharge
Xpre_column_16 bl[16] br[16] en vdd precharge
Xpre_column_17 bl[17] br[17] en vdd precharge
Xpre_column_18 bl[18] br[18] en vdd precharge
Xpre_column_19 bl[19] br[19] en vdd precharge
Xpre_column_20 bl[20] br[20] en vdd precharge
Xpre_column_21 bl[21] br[21] en vdd precharge
Xpre_column_22 bl[22] br[22] en vdd precharge
Xpre_column_23 bl[23] br[23] en vdd precharge
Xpre_column_24 bl[24] br[24] en vdd precharge
Xpre_column_25 bl[25] br[25] en vdd precharge
Xpre_column_26 bl[26] br[26] en vdd precharge
Xpre_column_27 bl[27] br[27] en vdd precharge
Xpre_column_28 bl[28] br[28] en vdd precharge
Xpre_column_29 bl[29] br[29] en vdd precharge
Xpre_column_30 bl[30] br[30] en vdd precharge
Xpre_column_31 bl[31] br[31] en vdd precharge
Xpre_column_32 bl[32] br[32] en vdd precharge
Xpre_column_33 bl[33] br[33] en vdd precharge
Xpre_column_34 bl[34] br[34] en vdd precharge
Xpre_column_35 bl[35] br[35] en vdd precharge
Xpre_column_36 bl[36] br[36] en vdd precharge
Xpre_column_37 bl[37] br[37] en vdd precharge
Xpre_column_38 bl[38] br[38] en vdd precharge
Xpre_column_39 bl[39] br[39] en vdd precharge
Xpre_column_40 bl[40] br[40] en vdd precharge
Xpre_column_41 bl[41] br[41] en vdd precharge
Xpre_column_42 bl[42] br[42] en vdd precharge
Xpre_column_43 bl[43] br[43] en vdd precharge
Xpre_column_44 bl[44] br[44] en vdd precharge
Xpre_column_45 bl[45] br[45] en vdd precharge
Xpre_column_46 bl[46] br[46] en vdd precharge
Xpre_column_47 bl[47] br[47] en vdd precharge
Xpre_column_48 bl[48] br[48] en vdd precharge
Xpre_column_49 bl[49] br[49] en vdd precharge
Xpre_column_50 bl[50] br[50] en vdd precharge
Xpre_column_51 bl[51] br[51] en vdd precharge
Xpre_column_52 bl[52] br[52] en vdd precharge
Xpre_column_53 bl[53] br[53] en vdd precharge
Xpre_column_54 bl[54] br[54] en vdd precharge
Xpre_column_55 bl[55] br[55] en vdd precharge
Xpre_column_56 bl[56] br[56] en vdd precharge
Xpre_column_57 bl[57] br[57] en vdd precharge
Xpre_column_58 bl[58] br[58] en vdd precharge
Xpre_column_59 bl[59] br[59] en vdd precharge
Xpre_column_60 bl[60] br[60] en vdd precharge
Xpre_column_61 bl[61] br[61] en vdd precharge
Xpre_column_62 bl[62] br[62] en vdd precharge
Xpre_column_63 bl[63] br[63] en vdd precharge
Xpre_column_64 bl[64] br[64] en vdd precharge
Xpre_column_65 bl[65] br[65] en vdd precharge
Xpre_column_66 bl[66] br[66] en vdd precharge
Xpre_column_67 bl[67] br[67] en vdd precharge
Xpre_column_68 bl[68] br[68] en vdd precharge
Xpre_column_69 bl[69] br[69] en vdd precharge
Xpre_column_70 bl[70] br[70] en vdd precharge
Xpre_column_71 bl[71] br[71] en vdd precharge
Xpre_column_72 bl[72] br[72] en vdd precharge
Xpre_column_73 bl[73] br[73] en vdd precharge
Xpre_column_74 bl[74] br[74] en vdd precharge
Xpre_column_75 bl[75] br[75] en vdd precharge
Xpre_column_76 bl[76] br[76] en vdd precharge
Xpre_column_77 bl[77] br[77] en vdd precharge
Xpre_column_78 bl[78] br[78] en vdd precharge
Xpre_column_79 bl[79] br[79] en vdd precharge
Xpre_column_80 bl[80] br[80] en vdd precharge
Xpre_column_81 bl[81] br[81] en vdd precharge
Xpre_column_82 bl[82] br[82] en vdd precharge
Xpre_column_83 bl[83] br[83] en vdd precharge
Xpre_column_84 bl[84] br[84] en vdd precharge
Xpre_column_85 bl[85] br[85] en vdd precharge
Xpre_column_86 bl[86] br[86] en vdd precharge
Xpre_column_87 bl[87] br[87] en vdd precharge
Xpre_column_88 bl[88] br[88] en vdd precharge
Xpre_column_89 bl[89] br[89] en vdd precharge
Xpre_column_90 bl[90] br[90] en vdd precharge
Xpre_column_91 bl[91] br[91] en vdd precharge
Xpre_column_92 bl[92] br[92] en vdd precharge
Xpre_column_93 bl[93] br[93] en vdd precharge
Xpre_column_94 bl[94] br[94] en vdd precharge
Xpre_column_95 bl[95] br[95] en vdd precharge
Xpre_column_96 bl[96] br[96] en vdd precharge
Xpre_column_97 bl[97] br[97] en vdd precharge
Xpre_column_98 bl[98] br[98] en vdd precharge
Xpre_column_99 bl[99] br[99] en vdd precharge
Xpre_column_100 bl[100] br[100] en vdd precharge
Xpre_column_101 bl[101] br[101] en vdd precharge
Xpre_column_102 bl[102] br[102] en vdd precharge
Xpre_column_103 bl[103] br[103] en vdd precharge
Xpre_column_104 bl[104] br[104] en vdd precharge
Xpre_column_105 bl[105] br[105] en vdd precharge
Xpre_column_106 bl[106] br[106] en vdd precharge
Xpre_column_107 bl[107] br[107] en vdd precharge
Xpre_column_108 bl[108] br[108] en vdd precharge
Xpre_column_109 bl[109] br[109] en vdd precharge
Xpre_column_110 bl[110] br[110] en vdd precharge
Xpre_column_111 bl[111] br[111] en vdd precharge
Xpre_column_112 bl[112] br[112] en vdd precharge
Xpre_column_113 bl[113] br[113] en vdd precharge
Xpre_column_114 bl[114] br[114] en vdd precharge
Xpre_column_115 bl[115] br[115] en vdd precharge
Xpre_column_116 bl[116] br[116] en vdd precharge
Xpre_column_117 bl[117] br[117] en vdd precharge
Xpre_column_118 bl[118] br[118] en vdd precharge
Xpre_column_119 bl[119] br[119] en vdd precharge
Xpre_column_120 bl[120] br[120] en vdd precharge
Xpre_column_121 bl[121] br[121] en vdd precharge
Xpre_column_122 bl[122] br[122] en vdd precharge
Xpre_column_123 bl[123] br[123] en vdd precharge
Xpre_column_124 bl[124] br[124] en vdd precharge
Xpre_column_125 bl[125] br[125] en vdd precharge
Xpre_column_126 bl[126] br[126] en vdd precharge
Xpre_column_127 bl[127] br[127] en vdd precharge
.ENDS precharge_array

* ptx M{0} {1} nmos_vtg m=1 w=0.72u l=0.05u pd=1.54u ps=1.54u as=0.09p ad=0.09p

.SUBCKT single_level_column_mux_8 bl br bl_out br_out sel gnd
Mmux_tx1 bl sel bl_out gnd nmos_vtg m=1 w=0.72u l=0.05u pd=1.54u ps=1.54u as=0.09p ad=0.09p
Mmux_tx2 br sel br_out gnd nmos_vtg m=1 w=0.72u l=0.05u pd=1.54u ps=1.54u as=0.09p ad=0.09p
.ENDS single_level_column_mux_8

.SUBCKT columnmux_array bl[0] br[0] bl[1] br[1] bl[2] br[2] bl[3] br[3] bl[4] br[4] bl[5] br[5] bl[6] br[6] bl[7] br[7] bl[8] br[8] bl[9] br[9] bl[10] br[10] bl[11] br[11] bl[12] br[12] bl[13] br[13] bl[14] br[14] bl[15] br[15] bl[16] br[16] bl[17] br[17] bl[18] br[18] bl[19] br[19] bl[20] br[20] bl[21] br[21] bl[22] br[22] bl[23] br[23] bl[24] br[24] bl[25] br[25] bl[26] br[26] bl[27] br[27] bl[28] br[28] bl[29] br[29] bl[30] br[30] bl[31] br[31] bl[32] br[32] bl[33] br[33] bl[34] br[34] bl[35] br[35] bl[36] br[36] bl[37] br[37] bl[38] br[38] bl[39] br[39] bl[40] br[40] bl[41] br[41] bl[42] br[42] bl[43] br[43] bl[44] br[44] bl[45] br[45] bl[46] br[46] bl[47] br[47] bl[48] br[48] bl[49] br[49] bl[50] br[50] bl[51] br[51] bl[52] br[52] bl[53] br[53] bl[54] br[54] bl[55] br[55] bl[56] br[56] bl[57] br[57] bl[58] br[58] bl[59] br[59] bl[60] br[60] bl[61] br[61] bl[62] br[62] bl[63] br[63] bl[64] br[64] bl[65] br[65] bl[66] br[66] bl[67] br[67] bl[68] br[68] bl[69] br[69] bl[70] br[70] bl[71] br[71] bl[72] br[72] bl[73] br[73] bl[74] br[74] bl[75] br[75] bl[76] br[76] bl[77] br[77] bl[78] br[78] bl[79] br[79] bl[80] br[80] bl[81] br[81] bl[82] br[82] bl[83] br[83] bl[84] br[84] bl[85] br[85] bl[86] br[86] bl[87] br[87] bl[88] br[88] bl[89] br[89] bl[90] br[90] bl[91] br[91] bl[92] br[92] bl[93] br[93] bl[94] br[94] bl[95] br[95] bl[96] br[96] bl[97] br[97] bl[98] br[98] bl[99] br[99] bl[100] br[100] bl[101] br[101] bl[102] br[102] bl[103] br[103] bl[104] br[104] bl[105] br[105] bl[106] br[106] bl[107] br[107] bl[108] br[108] bl[109] br[109] bl[110] br[110] bl[111] br[111] bl[112] br[112] bl[113] br[113] bl[114] br[114] bl[115] br[115] bl[116] br[116] bl[117] br[117] bl[118] br[118] bl[119] br[119] bl[120] br[120] bl[121] br[121] bl[122] br[122] bl[123] br[123] bl[124] br[124] bl[125] br[125] bl[126] br[126] bl[127] br[127] sel[0] sel[1] sel[2] sel[3] bl_out[0] br_out[0] bl_out[1] br_out[1] bl_out[2] br_out[2] bl_out[3] br_out[3] bl_out[4] br_out[4] bl_out[5] br_out[5] bl_out[6] br_out[6] bl_out[7] br_out[7] bl_out[8] br_out[8] bl_out[9] br_out[9] bl_out[10] br_out[10] bl_out[11] br_out[11] bl_out[12] br_out[12] bl_out[13] br_out[13] bl_out[14] br_out[14] bl_out[15] br_out[15] bl_out[16] br_out[16] bl_out[17] br_out[17] bl_out[18] br_out[18] bl_out[19] br_out[19] bl_out[20] br_out[20] bl_out[21] br_out[21] bl_out[22] br_out[22] bl_out[23] br_out[23] bl_out[24] br_out[24] bl_out[25] br_out[25] bl_out[26] br_out[26] bl_out[27] br_out[27] bl_out[28] br_out[28] bl_out[29] br_out[29] bl_out[30] br_out[30] bl_out[31] br_out[31] gnd
XXMUX0 bl[0] br[0] bl_out[0] br_out[0] sel[0] gnd single_level_column_mux_8
XXMUX1 bl[1] br[1] bl_out[0] br_out[0] sel[1] gnd single_level_column_mux_8
XXMUX2 bl[2] br[2] bl_out[0] br_out[0] sel[2] gnd single_level_column_mux_8
XXMUX3 bl[3] br[3] bl_out[0] br_out[0] sel[3] gnd single_level_column_mux_8
XXMUX4 bl[4] br[4] bl_out[1] br_out[1] sel[0] gnd single_level_column_mux_8
XXMUX5 bl[5] br[5] bl_out[1] br_out[1] sel[1] gnd single_level_column_mux_8
XXMUX6 bl[6] br[6] bl_out[1] br_out[1] sel[2] gnd single_level_column_mux_8
XXMUX7 bl[7] br[7] bl_out[1] br_out[1] sel[3] gnd single_level_column_mux_8
XXMUX8 bl[8] br[8] bl_out[2] br_out[2] sel[0] gnd single_level_column_mux_8
XXMUX9 bl[9] br[9] bl_out[2] br_out[2] sel[1] gnd single_level_column_mux_8
XXMUX10 bl[10] br[10] bl_out[2] br_out[2] sel[2] gnd single_level_column_mux_8
XXMUX11 bl[11] br[11] bl_out[2] br_out[2] sel[3] gnd single_level_column_mux_8
XXMUX12 bl[12] br[12] bl_out[3] br_out[3] sel[0] gnd single_level_column_mux_8
XXMUX13 bl[13] br[13] bl_out[3] br_out[3] sel[1] gnd single_level_column_mux_8
XXMUX14 bl[14] br[14] bl_out[3] br_out[3] sel[2] gnd single_level_column_mux_8
XXMUX15 bl[15] br[15] bl_out[3] br_out[3] sel[3] gnd single_level_column_mux_8
XXMUX16 bl[16] br[16] bl_out[4] br_out[4] sel[0] gnd single_level_column_mux_8
XXMUX17 bl[17] br[17] bl_out[4] br_out[4] sel[1] gnd single_level_column_mux_8
XXMUX18 bl[18] br[18] bl_out[4] br_out[4] sel[2] gnd single_level_column_mux_8
XXMUX19 bl[19] br[19] bl_out[4] br_out[4] sel[3] gnd single_level_column_mux_8
XXMUX20 bl[20] br[20] bl_out[5] br_out[5] sel[0] gnd single_level_column_mux_8
XXMUX21 bl[21] br[21] bl_out[5] br_out[5] sel[1] gnd single_level_column_mux_8
XXMUX22 bl[22] br[22] bl_out[5] br_out[5] sel[2] gnd single_level_column_mux_8
XXMUX23 bl[23] br[23] bl_out[5] br_out[5] sel[3] gnd single_level_column_mux_8
XXMUX24 bl[24] br[24] bl_out[6] br_out[6] sel[0] gnd single_level_column_mux_8
XXMUX25 bl[25] br[25] bl_out[6] br_out[6] sel[1] gnd single_level_column_mux_8
XXMUX26 bl[26] br[26] bl_out[6] br_out[6] sel[2] gnd single_level_column_mux_8
XXMUX27 bl[27] br[27] bl_out[6] br_out[6] sel[3] gnd single_level_column_mux_8
XXMUX28 bl[28] br[28] bl_out[7] br_out[7] sel[0] gnd single_level_column_mux_8
XXMUX29 bl[29] br[29] bl_out[7] br_out[7] sel[1] gnd single_level_column_mux_8
XXMUX30 bl[30] br[30] bl_out[7] br_out[7] sel[2] gnd single_level_column_mux_8
XXMUX31 bl[31] br[31] bl_out[7] br_out[7] sel[3] gnd single_level_column_mux_8
XXMUX32 bl[32] br[32] bl_out[8] br_out[8] sel[0] gnd single_level_column_mux_8
XXMUX33 bl[33] br[33] bl_out[8] br_out[8] sel[1] gnd single_level_column_mux_8
XXMUX34 bl[34] br[34] bl_out[8] br_out[8] sel[2] gnd single_level_column_mux_8
XXMUX35 bl[35] br[35] bl_out[8] br_out[8] sel[3] gnd single_level_column_mux_8
XXMUX36 bl[36] br[36] bl_out[9] br_out[9] sel[0] gnd single_level_column_mux_8
XXMUX37 bl[37] br[37] bl_out[9] br_out[9] sel[1] gnd single_level_column_mux_8
XXMUX38 bl[38] br[38] bl_out[9] br_out[9] sel[2] gnd single_level_column_mux_8
XXMUX39 bl[39] br[39] bl_out[9] br_out[9] sel[3] gnd single_level_column_mux_8
XXMUX40 bl[40] br[40] bl_out[10] br_out[10] sel[0] gnd single_level_column_mux_8
XXMUX41 bl[41] br[41] bl_out[10] br_out[10] sel[1] gnd single_level_column_mux_8
XXMUX42 bl[42] br[42] bl_out[10] br_out[10] sel[2] gnd single_level_column_mux_8
XXMUX43 bl[43] br[43] bl_out[10] br_out[10] sel[3] gnd single_level_column_mux_8
XXMUX44 bl[44] br[44] bl_out[11] br_out[11] sel[0] gnd single_level_column_mux_8
XXMUX45 bl[45] br[45] bl_out[11] br_out[11] sel[1] gnd single_level_column_mux_8
XXMUX46 bl[46] br[46] bl_out[11] br_out[11] sel[2] gnd single_level_column_mux_8
XXMUX47 bl[47] br[47] bl_out[11] br_out[11] sel[3] gnd single_level_column_mux_8
XXMUX48 bl[48] br[48] bl_out[12] br_out[12] sel[0] gnd single_level_column_mux_8
XXMUX49 bl[49] br[49] bl_out[12] br_out[12] sel[1] gnd single_level_column_mux_8
XXMUX50 bl[50] br[50] bl_out[12] br_out[12] sel[2] gnd single_level_column_mux_8
XXMUX51 bl[51] br[51] bl_out[12] br_out[12] sel[3] gnd single_level_column_mux_8
XXMUX52 bl[52] br[52] bl_out[13] br_out[13] sel[0] gnd single_level_column_mux_8
XXMUX53 bl[53] br[53] bl_out[13] br_out[13] sel[1] gnd single_level_column_mux_8
XXMUX54 bl[54] br[54] bl_out[13] br_out[13] sel[2] gnd single_level_column_mux_8
XXMUX55 bl[55] br[55] bl_out[13] br_out[13] sel[3] gnd single_level_column_mux_8
XXMUX56 bl[56] br[56] bl_out[14] br_out[14] sel[0] gnd single_level_column_mux_8
XXMUX57 bl[57] br[57] bl_out[14] br_out[14] sel[1] gnd single_level_column_mux_8
XXMUX58 bl[58] br[58] bl_out[14] br_out[14] sel[2] gnd single_level_column_mux_8
XXMUX59 bl[59] br[59] bl_out[14] br_out[14] sel[3] gnd single_level_column_mux_8
XXMUX60 bl[60] br[60] bl_out[15] br_out[15] sel[0] gnd single_level_column_mux_8
XXMUX61 bl[61] br[61] bl_out[15] br_out[15] sel[1] gnd single_level_column_mux_8
XXMUX62 bl[62] br[62] bl_out[15] br_out[15] sel[2] gnd single_level_column_mux_8
XXMUX63 bl[63] br[63] bl_out[15] br_out[15] sel[3] gnd single_level_column_mux_8
XXMUX64 bl[64] br[64] bl_out[16] br_out[16] sel[0] gnd single_level_column_mux_8
XXMUX65 bl[65] br[65] bl_out[16] br_out[16] sel[1] gnd single_level_column_mux_8
XXMUX66 bl[66] br[66] bl_out[16] br_out[16] sel[2] gnd single_level_column_mux_8
XXMUX67 bl[67] br[67] bl_out[16] br_out[16] sel[3] gnd single_level_column_mux_8
XXMUX68 bl[68] br[68] bl_out[17] br_out[17] sel[0] gnd single_level_column_mux_8
XXMUX69 bl[69] br[69] bl_out[17] br_out[17] sel[1] gnd single_level_column_mux_8
XXMUX70 bl[70] br[70] bl_out[17] br_out[17] sel[2] gnd single_level_column_mux_8
XXMUX71 bl[71] br[71] bl_out[17] br_out[17] sel[3] gnd single_level_column_mux_8
XXMUX72 bl[72] br[72] bl_out[18] br_out[18] sel[0] gnd single_level_column_mux_8
XXMUX73 bl[73] br[73] bl_out[18] br_out[18] sel[1] gnd single_level_column_mux_8
XXMUX74 bl[74] br[74] bl_out[18] br_out[18] sel[2] gnd single_level_column_mux_8
XXMUX75 bl[75] br[75] bl_out[18] br_out[18] sel[3] gnd single_level_column_mux_8
XXMUX76 bl[76] br[76] bl_out[19] br_out[19] sel[0] gnd single_level_column_mux_8
XXMUX77 bl[77] br[77] bl_out[19] br_out[19] sel[1] gnd single_level_column_mux_8
XXMUX78 bl[78] br[78] bl_out[19] br_out[19] sel[2] gnd single_level_column_mux_8
XXMUX79 bl[79] br[79] bl_out[19] br_out[19] sel[3] gnd single_level_column_mux_8
XXMUX80 bl[80] br[80] bl_out[20] br_out[20] sel[0] gnd single_level_column_mux_8
XXMUX81 bl[81] br[81] bl_out[20] br_out[20] sel[1] gnd single_level_column_mux_8
XXMUX82 bl[82] br[82] bl_out[20] br_out[20] sel[2] gnd single_level_column_mux_8
XXMUX83 bl[83] br[83] bl_out[20] br_out[20] sel[3] gnd single_level_column_mux_8
XXMUX84 bl[84] br[84] bl_out[21] br_out[21] sel[0] gnd single_level_column_mux_8
XXMUX85 bl[85] br[85] bl_out[21] br_out[21] sel[1] gnd single_level_column_mux_8
XXMUX86 bl[86] br[86] bl_out[21] br_out[21] sel[2] gnd single_level_column_mux_8
XXMUX87 bl[87] br[87] bl_out[21] br_out[21] sel[3] gnd single_level_column_mux_8
XXMUX88 bl[88] br[88] bl_out[22] br_out[22] sel[0] gnd single_level_column_mux_8
XXMUX89 bl[89] br[89] bl_out[22] br_out[22] sel[1] gnd single_level_column_mux_8
XXMUX90 bl[90] br[90] bl_out[22] br_out[22] sel[2] gnd single_level_column_mux_8
XXMUX91 bl[91] br[91] bl_out[22] br_out[22] sel[3] gnd single_level_column_mux_8
XXMUX92 bl[92] br[92] bl_out[23] br_out[23] sel[0] gnd single_level_column_mux_8
XXMUX93 bl[93] br[93] bl_out[23] br_out[23] sel[1] gnd single_level_column_mux_8
XXMUX94 bl[94] br[94] bl_out[23] br_out[23] sel[2] gnd single_level_column_mux_8
XXMUX95 bl[95] br[95] bl_out[23] br_out[23] sel[3] gnd single_level_column_mux_8
XXMUX96 bl[96] br[96] bl_out[24] br_out[24] sel[0] gnd single_level_column_mux_8
XXMUX97 bl[97] br[97] bl_out[24] br_out[24] sel[1] gnd single_level_column_mux_8
XXMUX98 bl[98] br[98] bl_out[24] br_out[24] sel[2] gnd single_level_column_mux_8
XXMUX99 bl[99] br[99] bl_out[24] br_out[24] sel[3] gnd single_level_column_mux_8
XXMUX100 bl[100] br[100] bl_out[25] br_out[25] sel[0] gnd single_level_column_mux_8
XXMUX101 bl[101] br[101] bl_out[25] br_out[25] sel[1] gnd single_level_column_mux_8
XXMUX102 bl[102] br[102] bl_out[25] br_out[25] sel[2] gnd single_level_column_mux_8
XXMUX103 bl[103] br[103] bl_out[25] br_out[25] sel[3] gnd single_level_column_mux_8
XXMUX104 bl[104] br[104] bl_out[26] br_out[26] sel[0] gnd single_level_column_mux_8
XXMUX105 bl[105] br[105] bl_out[26] br_out[26] sel[1] gnd single_level_column_mux_8
XXMUX106 bl[106] br[106] bl_out[26] br_out[26] sel[2] gnd single_level_column_mux_8
XXMUX107 bl[107] br[107] bl_out[26] br_out[26] sel[3] gnd single_level_column_mux_8
XXMUX108 bl[108] br[108] bl_out[27] br_out[27] sel[0] gnd single_level_column_mux_8
XXMUX109 bl[109] br[109] bl_out[27] br_out[27] sel[1] gnd single_level_column_mux_8
XXMUX110 bl[110] br[110] bl_out[27] br_out[27] sel[2] gnd single_level_column_mux_8
XXMUX111 bl[111] br[111] bl_out[27] br_out[27] sel[3] gnd single_level_column_mux_8
XXMUX112 bl[112] br[112] bl_out[28] br_out[28] sel[0] gnd single_level_column_mux_8
XXMUX113 bl[113] br[113] bl_out[28] br_out[28] sel[1] gnd single_level_column_mux_8
XXMUX114 bl[114] br[114] bl_out[28] br_out[28] sel[2] gnd single_level_column_mux_8
XXMUX115 bl[115] br[115] bl_out[28] br_out[28] sel[3] gnd single_level_column_mux_8
XXMUX116 bl[116] br[116] bl_out[29] br_out[29] sel[0] gnd single_level_column_mux_8
XXMUX117 bl[117] br[117] bl_out[29] br_out[29] sel[1] gnd single_level_column_mux_8
XXMUX118 bl[118] br[118] bl_out[29] br_out[29] sel[2] gnd single_level_column_mux_8
XXMUX119 bl[119] br[119] bl_out[29] br_out[29] sel[3] gnd single_level_column_mux_8
XXMUX120 bl[120] br[120] bl_out[30] br_out[30] sel[0] gnd single_level_column_mux_8
XXMUX121 bl[121] br[121] bl_out[30] br_out[30] sel[1] gnd single_level_column_mux_8
XXMUX122 bl[122] br[122] bl_out[30] br_out[30] sel[2] gnd single_level_column_mux_8
XXMUX123 bl[123] br[123] bl_out[30] br_out[30] sel[3] gnd single_level_column_mux_8
XXMUX124 bl[124] br[124] bl_out[31] br_out[31] sel[0] gnd single_level_column_mux_8
XXMUX125 bl[125] br[125] bl_out[31] br_out[31] sel[1] gnd single_level_column_mux_8
XXMUX126 bl[126] br[126] bl_out[31] br_out[31] sel[2] gnd single_level_column_mux_8
XXMUX127 bl[127] br[127] bl_out[31] br_out[31] sel[3] gnd single_level_column_mux_8
.ENDS columnmux_array

.SUBCKT sense_amp bl br dout en vdd gnd
M_1 dout net_1 vdd vdd pmos_vtg w=540.0n l=50.0n
M_3 net_1 dout vdd vdd pmos_vtg w=540.0n l=50.0n
M_2 dout net_1 net_2 gnd nmos_vtg w=270.0n l=50.0n
M_8 net_1 dout net_2 gnd nmos_vtg w=270.0n l=50.0n
M_5 bl en dout vdd pmos_vtg w=720.0n l=50.0n
M_6 br en net_1 vdd pmos_vtg w=720.0n l=50.0n
M_7 net_2 en gnd gnd nmos_vtg w=270.0n l=50.0n
.ENDS sense_amp


.SUBCKT sense_amp_array data[0] bl[0] br[0] data[1] bl[4] br[4] data[2] bl[8] br[8] data[3] bl[12] br[12] data[4] bl[16] br[16] data[5] bl[20] br[20] data[6] bl[24] br[24] data[7] bl[28] br[28] data[8] bl[32] br[32] data[9] bl[36] br[36] data[10] bl[40] br[40] data[11] bl[44] br[44] data[12] bl[48] br[48] data[13] bl[52] br[52] data[14] bl[56] br[56] data[15] bl[60] br[60] data[16] bl[64] br[64] data[17] bl[68] br[68] data[18] bl[72] br[72] data[19] bl[76] br[76] data[20] bl[80] br[80] data[21] bl[84] br[84] data[22] bl[88] br[88] data[23] bl[92] br[92] data[24] bl[96] br[96] data[25] bl[100] br[100] data[26] bl[104] br[104] data[27] bl[108] br[108] data[28] bl[112] br[112] data[29] bl[116] br[116] data[30] bl[120] br[120] data[31] bl[124] br[124] en vdd gnd
Xsa_d0 bl[0] br[0] data[0] en vdd gnd sense_amp
Xsa_d4 bl[4] br[4] data[1] en vdd gnd sense_amp
Xsa_d8 bl[8] br[8] data[2] en vdd gnd sense_amp
Xsa_d12 bl[12] br[12] data[3] en vdd gnd sense_amp
Xsa_d16 bl[16] br[16] data[4] en vdd gnd sense_amp
Xsa_d20 bl[20] br[20] data[5] en vdd gnd sense_amp
Xsa_d24 bl[24] br[24] data[6] en vdd gnd sense_amp
Xsa_d28 bl[28] br[28] data[7] en vdd gnd sense_amp
Xsa_d32 bl[32] br[32] data[8] en vdd gnd sense_amp
Xsa_d36 bl[36] br[36] data[9] en vdd gnd sense_amp
Xsa_d40 bl[40] br[40] data[10] en vdd gnd sense_amp
Xsa_d44 bl[44] br[44] data[11] en vdd gnd sense_amp
Xsa_d48 bl[48] br[48] data[12] en vdd gnd sense_amp
Xsa_d52 bl[52] br[52] data[13] en vdd gnd sense_amp
Xsa_d56 bl[56] br[56] data[14] en vdd gnd sense_amp
Xsa_d60 bl[60] br[60] data[15] en vdd gnd sense_amp
Xsa_d64 bl[64] br[64] data[16] en vdd gnd sense_amp
Xsa_d68 bl[68] br[68] data[17] en vdd gnd sense_amp
Xsa_d72 bl[72] br[72] data[18] en vdd gnd sense_amp
Xsa_d76 bl[76] br[76] data[19] en vdd gnd sense_amp
Xsa_d80 bl[80] br[80] data[20] en vdd gnd sense_amp
Xsa_d84 bl[84] br[84] data[21] en vdd gnd sense_amp
Xsa_d88 bl[88] br[88] data[22] en vdd gnd sense_amp
Xsa_d92 bl[92] br[92] data[23] en vdd gnd sense_amp
Xsa_d96 bl[96] br[96] data[24] en vdd gnd sense_amp
Xsa_d100 bl[100] br[100] data[25] en vdd gnd sense_amp
Xsa_d104 bl[104] br[104] data[26] en vdd gnd sense_amp
Xsa_d108 bl[108] br[108] data[27] en vdd gnd sense_amp
Xsa_d112 bl[112] br[112] data[28] en vdd gnd sense_amp
Xsa_d116 bl[116] br[116] data[29] en vdd gnd sense_amp
Xsa_d120 bl[120] br[120] data[30] en vdd gnd sense_amp
Xsa_d124 bl[124] br[124] data[31] en vdd gnd sense_amp
.ENDS sense_amp_array

.SUBCKT write_driver din bl br en vdd gnd
*inverters for enable and data input
minP bl_bar din vdd vdd pmos_vtg w=360.000000n l=50.000000n
minN bl_bar din gnd gnd nmos_vtg w=180.000000n l=50.000000n
moutP en_bar en vdd vdd pmos_vtg w=360.000000n l=50.000000n
moutN en_bar en gnd gnd nmos_vtg w=180.000000n l=50.000000n

*tristate for BL
mout0P int1 bl_bar vdd vdd pmos_vtg w=360.000000n l=50.000000n
mout0P2 bl en_bar int1 vdd pmos_vtg w=360.000000n l=50.000000n
mout0N bl en int2 gnd nmos_vtg w=180.000000n l=50.000000n
mout0N2 int2 bl_bar gnd gnd nmos_vtg w=180.000000n l=50.000000n

*tristate for BR
mout1P int3 din vdd vdd pmos_vtg w=360.000000n l=50.000000n
mout1P2 br en_bar int3 vdd pmos_vtg w=360.000000n l=50.000000n
mout1N br en int4 gnd nmos_vtg w=180.000000n l=50.000000n
mout1N2 int4 din gnd gnd nmos_vtg w=180.000000n l=50.000000n
.ENDS write_driver


.SUBCKT write_driver_array data[0] data[1] data[2] data[3] data[4] data[5] data[6] data[7] data[8] data[9] data[10] data[11] data[12] data[13] data[14] data[15] data[16] data[17] data[18] data[19] data[20] data[21] data[22] data[23] data[24] data[25] data[26] data[27] data[28] data[29] data[30] data[31] bl[0] br[0] bl[1] br[1] bl[2] br[2] bl[3] br[3] bl[4] br[4] bl[5] br[5] bl[6] br[6] bl[7] br[7] bl[8] br[8] bl[9] br[9] bl[10] br[10] bl[11] br[11] bl[12] br[12] bl[13] br[13] bl[14] br[14] bl[15] br[15] bl[16] br[16] bl[17] br[17] bl[18] br[18] bl[19] br[19] bl[20] br[20] bl[21] br[21] bl[22] br[22] bl[23] br[23] bl[24] br[24] bl[25] br[25] bl[26] br[26] bl[27] br[27] bl[28] br[28] bl[29] br[29] bl[30] br[30] bl[31] br[31] en vdd gnd
XXwrite_driver0 data[0] bl[0] br[0] en vdd gnd write_driver
XXwrite_driver4 data[1] bl[1] br[1] en vdd gnd write_driver
XXwrite_driver8 data[2] bl[2] br[2] en vdd gnd write_driver
XXwrite_driver12 data[3] bl[3] br[3] en vdd gnd write_driver
XXwrite_driver16 data[4] bl[4] br[4] en vdd gnd write_driver
XXwrite_driver20 data[5] bl[5] br[5] en vdd gnd write_driver
XXwrite_driver24 data[6] bl[6] br[6] en vdd gnd write_driver
XXwrite_driver28 data[7] bl[7] br[7] en vdd gnd write_driver
XXwrite_driver32 data[8] bl[8] br[8] en vdd gnd write_driver
XXwrite_driver36 data[9] bl[9] br[9] en vdd gnd write_driver
XXwrite_driver40 data[10] bl[10] br[10] en vdd gnd write_driver
XXwrite_driver44 data[11] bl[11] br[11] en vdd gnd write_driver
XXwrite_driver48 data[12] bl[12] br[12] en vdd gnd write_driver
XXwrite_driver52 data[13] bl[13] br[13] en vdd gnd write_driver
XXwrite_driver56 data[14] bl[14] br[14] en vdd gnd write_driver
XXwrite_driver60 data[15] bl[15] br[15] en vdd gnd write_driver
XXwrite_driver64 data[16] bl[16] br[16] en vdd gnd write_driver
XXwrite_driver68 data[17] bl[17] br[17] en vdd gnd write_driver
XXwrite_driver72 data[18] bl[18] br[18] en vdd gnd write_driver
XXwrite_driver76 data[19] bl[19] br[19] en vdd gnd write_driver
XXwrite_driver80 data[20] bl[20] br[20] en vdd gnd write_driver
XXwrite_driver84 data[21] bl[21] br[21] en vdd gnd write_driver
XXwrite_driver88 data[22] bl[22] br[22] en vdd gnd write_driver
XXwrite_driver92 data[23] bl[23] br[23] en vdd gnd write_driver
XXwrite_driver96 data[24] bl[24] br[24] en vdd gnd write_driver
XXwrite_driver100 data[25] bl[25] br[25] en vdd gnd write_driver
XXwrite_driver104 data[26] bl[26] br[26] en vdd gnd write_driver
XXwrite_driver108 data[27] bl[27] br[27] en vdd gnd write_driver
XXwrite_driver112 data[28] bl[28] br[28] en vdd gnd write_driver
XXwrite_driver116 data[29] bl[29] br[29] en vdd gnd write_driver
XXwrite_driver120 data[30] bl[30] br[30] en vdd gnd write_driver
XXwrite_driver124 data[31] bl[31] br[31] en vdd gnd write_driver
.ENDS write_driver_array

.SUBCKT pinv_8 A Z vdd gnd
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01125p ad=0.01125p
.ENDS pinv_8

.SUBCKT pnand2_2 A B Z vdd gnd
Mpnand2_pmos1 vdd A Z vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpnand2_pmos2 Z B vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpnand2_nmos1 Z B net1 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.0225p ad=0.0225p
Mpnand2_nmos2 net1 A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.0225p ad=0.0225p
.ENDS pnand2_2

.SUBCKT pnand3_2 A B C Z vdd gnd
Mpnand3_pmos1 vdd A Z vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpnand3_pmos2 Z B vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpnand3_pmos3 Z C vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpnand3_nmos1 Z C net1 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.0225p ad=0.0225p
Mpnand3_nmos2 net1 B net2 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.0225p ad=0.0225p
Mpnand3_nmos3 net2 A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.0225p ad=0.0225p
.ENDS pnand3_2

.SUBCKT pinv_9 A Z vdd gnd
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01125p ad=0.01125p
.ENDS pinv_9

.SUBCKT pnand2_3 A B Z vdd gnd
Mpnand2_pmos1 vdd A Z vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpnand2_pmos2 Z B vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpnand2_nmos1 Z B net1 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.0225p ad=0.0225p
Mpnand2_nmos2 net1 A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.0225p ad=0.0225p
.ENDS pnand2_3

.SUBCKT pre2x4 in[0] in[1] out[0] out[1] out[2] out[3] vdd gnd
XXpre_inv[0] in[0] inbar[0] vdd gnd pinv_9
XXpre_inv[1] in[1] inbar[1] vdd gnd pinv_9
XXpre_nand_inv[0] Z[0] out[0] vdd gnd pinv_9
XXpre_nand_inv[1] Z[1] out[1] vdd gnd pinv_9
XXpre_nand_inv[2] Z[2] out[2] vdd gnd pinv_9
XXpre_nand_inv[3] Z[3] out[3] vdd gnd pinv_9
XXpre2x4_nand[0] inbar[0] inbar[1] Z[0] vdd gnd pnand2_3
XXpre2x4_nand[1] in[0] inbar[1] Z[1] vdd gnd pnand2_3
XXpre2x4_nand[2] inbar[0] in[1] Z[2] vdd gnd pnand2_3
XXpre2x4_nand[3] in[0] in[1] Z[3] vdd gnd pnand2_3
.ENDS pre2x4

.SUBCKT pinv_10 A Z vdd gnd
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01125p ad=0.01125p
.ENDS pinv_10

.SUBCKT pnand3_3 A B C Z vdd gnd
Mpnand3_pmos1 vdd A Z vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpnand3_pmos2 Z B vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpnand3_pmos3 Z C vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpnand3_nmos1 Z C net1 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.0225p ad=0.0225p
Mpnand3_nmos2 net1 B net2 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.0225p ad=0.0225p
Mpnand3_nmos3 net2 A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.0225p ad=0.0225p
.ENDS pnand3_3

.SUBCKT pre3x8 in[0] in[1] in[2] out[0] out[1] out[2] out[3] out[4] out[5] out[6] out[7] vdd gnd
XXpre_inv[0] in[0] inbar[0] vdd gnd pinv_10
XXpre_inv[1] in[1] inbar[1] vdd gnd pinv_10
XXpre_inv[2] in[2] inbar[2] vdd gnd pinv_10
XXpre_nand_inv[0] Z[0] out[0] vdd gnd pinv_10
XXpre_nand_inv[1] Z[1] out[1] vdd gnd pinv_10
XXpre_nand_inv[2] Z[2] out[2] vdd gnd pinv_10
XXpre_nand_inv[3] Z[3] out[3] vdd gnd pinv_10
XXpre_nand_inv[4] Z[4] out[4] vdd gnd pinv_10
XXpre_nand_inv[5] Z[5] out[5] vdd gnd pinv_10
XXpre_nand_inv[6] Z[6] out[6] vdd gnd pinv_10
XXpre_nand_inv[7] Z[7] out[7] vdd gnd pinv_10
XXpre3x8_nand[0] inbar[0] inbar[1] inbar[2] Z[0] vdd gnd pnand3_3
XXpre3x8_nand[1] in[0] inbar[1] inbar[2] Z[1] vdd gnd pnand3_3
XXpre3x8_nand[2] inbar[0] in[1] inbar[2] Z[2] vdd gnd pnand3_3
XXpre3x8_nand[3] in[0] in[1] inbar[2] Z[3] vdd gnd pnand3_3
XXpre3x8_nand[4] inbar[0] inbar[1] in[2] Z[4] vdd gnd pnand3_3
XXpre3x8_nand[5] in[0] inbar[1] in[2] Z[5] vdd gnd pnand3_3
XXpre3x8_nand[6] inbar[0] in[1] in[2] Z[6] vdd gnd pnand3_3
XXpre3x8_nand[7] in[0] in[1] in[2] Z[7] vdd gnd pnand3_3
.ENDS pre3x8

.SUBCKT hierarchical_decoder_512rows A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7] A[8] decode[0] decode[1] decode[2] decode[3] decode[4] decode[5] decode[6] decode[7] decode[8] decode[9] decode[10] decode[11] decode[12] decode[13] decode[14] decode[15] decode[16] decode[17] decode[18] decode[19] decode[20] decode[21] decode[22] decode[23] decode[24] decode[25] decode[26] decode[27] decode[28] decode[29] decode[30] decode[31] decode[32] decode[33] decode[34] decode[35] decode[36] decode[37] decode[38] decode[39] decode[40] decode[41] decode[42] decode[43] decode[44] decode[45] decode[46] decode[47] decode[48] decode[49] decode[50] decode[51] decode[52] decode[53] decode[54] decode[55] decode[56] decode[57] decode[58] decode[59] decode[60] decode[61] decode[62] decode[63] decode[64] decode[65] decode[66] decode[67] decode[68] decode[69] decode[70] decode[71] decode[72] decode[73] decode[74] decode[75] decode[76] decode[77] decode[78] decode[79] decode[80] decode[81] decode[82] decode[83] decode[84] decode[85] decode[86] decode[87] decode[88] decode[89] decode[90] decode[91] decode[92] decode[93] decode[94] decode[95] decode[96] decode[97] decode[98] decode[99] decode[100] decode[101] decode[102] decode[103] decode[104] decode[105] decode[106] decode[107] decode[108] decode[109] decode[110] decode[111] decode[112] decode[113] decode[114] decode[115] decode[116] decode[117] decode[118] decode[119] decode[120] decode[121] decode[122] decode[123] decode[124] decode[125] decode[126] decode[127] decode[128] decode[129] decode[130] decode[131] decode[132] decode[133] decode[134] decode[135] decode[136] decode[137] decode[138] decode[139] decode[140] decode[141] decode[142] decode[143] decode[144] decode[145] decode[146] decode[147] decode[148] decode[149] decode[150] decode[151] decode[152] decode[153] decode[154] decode[155] decode[156] decode[157] decode[158] decode[159] decode[160] decode[161] decode[162] decode[163] decode[164] decode[165] decode[166] decode[167] decode[168] decode[169] decode[170] decode[171] decode[172] decode[173] decode[174] decode[175] decode[176] decode[177] decode[178] decode[179] decode[180] decode[181] decode[182] decode[183] decode[184] decode[185] decode[186] decode[187] decode[188] decode[189] decode[190] decode[191] decode[192] decode[193] decode[194] decode[195] decode[196] decode[197] decode[198] decode[199] decode[200] decode[201] decode[202] decode[203] decode[204] decode[205] decode[206] decode[207] decode[208] decode[209] decode[210] decode[211] decode[212] decode[213] decode[214] decode[215] decode[216] decode[217] decode[218] decode[219] decode[220] decode[221] decode[222] decode[223] decode[224] decode[225] decode[226] decode[227] decode[228] decode[229] decode[230] decode[231] decode[232] decode[233] decode[234] decode[235] decode[236] decode[237] decode[238] decode[239] decode[240] decode[241] decode[242] decode[243] decode[244] decode[245] decode[246] decode[247] decode[248] decode[249] decode[250] decode[251] decode[252] decode[253] decode[254] decode[255] decode[256] decode[257] decode[258] decode[259] decode[260] decode[261] decode[262] decode[263] decode[264] decode[265] decode[266] decode[267] decode[268] decode[269] decode[270] decode[271] decode[272] decode[273] decode[274] decode[275] decode[276] decode[277] decode[278] decode[279] decode[280] decode[281] decode[282] decode[283] decode[284] decode[285] decode[286] decode[287] decode[288] decode[289] decode[290] decode[291] decode[292] decode[293] decode[294] decode[295] decode[296] decode[297] decode[298] decode[299] decode[300] decode[301] decode[302] decode[303] decode[304] decode[305] decode[306] decode[307] decode[308] decode[309] decode[310] decode[311] decode[312] decode[313] decode[314] decode[315] decode[316] decode[317] decode[318] decode[319] decode[320] decode[321] decode[322] decode[323] decode[324] decode[325] decode[326] decode[327] decode[328] decode[329] decode[330] decode[331] decode[332] decode[333] decode[334] decode[335] decode[336] decode[337] decode[338] decode[339] decode[340] decode[341] decode[342] decode[343] decode[344] decode[345] decode[346] decode[347] decode[348] decode[349] decode[350] decode[351] decode[352] decode[353] decode[354] decode[355] decode[356] decode[357] decode[358] decode[359] decode[360] decode[361] decode[362] decode[363] decode[364] decode[365] decode[366] decode[367] decode[368] decode[369] decode[370] decode[371] decode[372] decode[373] decode[374] decode[375] decode[376] decode[377] decode[378] decode[379] decode[380] decode[381] decode[382] decode[383] decode[384] decode[385] decode[386] decode[387] decode[388] decode[389] decode[390] decode[391] decode[392] decode[393] decode[394] decode[395] decode[396] decode[397] decode[398] decode[399] decode[400] decode[401] decode[402] decode[403] decode[404] decode[405] decode[406] decode[407] decode[408] decode[409] decode[410] decode[411] decode[412] decode[413] decode[414] decode[415] decode[416] decode[417] decode[418] decode[419] decode[420] decode[421] decode[422] decode[423] decode[424] decode[425] decode[426] decode[427] decode[428] decode[429] decode[430] decode[431] decode[432] decode[433] decode[434] decode[435] decode[436] decode[437] decode[438] decode[439] decode[440] decode[441] decode[442] decode[443] decode[444] decode[445] decode[446] decode[447] decode[448] decode[449] decode[450] decode[451] decode[452] decode[453] decode[454] decode[455] decode[456] decode[457] decode[458] decode[459] decode[460] decode[461] decode[462] decode[463] decode[464] decode[465] decode[466] decode[467] decode[468] decode[469] decode[470] decode[471] decode[472] decode[473] decode[474] decode[475] decode[476] decode[477] decode[478] decode[479] decode[480] decode[481] decode[482] decode[483] decode[484] decode[485] decode[486] decode[487] decode[488] decode[489] decode[490] decode[491] decode[492] decode[493] decode[494] decode[495] decode[496] decode[497] decode[498] decode[499] decode[500] decode[501] decode[502] decode[503] decode[504] decode[505] decode[506] decode[507] decode[508] decode[509] decode[510] decode[511] vdd gnd
Xpre3x8[0] A[0] A[1] A[2] out[0] out[1] out[2] out[3] out[4] out[5] out[6] out[7] vdd gnd pre3x8
Xpre3x8[1] A[3] A[4] A[5] out[8] out[9] out[10] out[11] out[12] out[13] out[14] out[15] vdd gnd pre3x8
Xpre3x8[2] A[6] A[7] A[8] out[16] out[17] out[18] out[19] out[20] out[21] out[22] out[23] vdd gnd pre3x8
XDEC_NAND[0] out[0] out[8] out[16] Z[0] vdd gnd pnand3_2
XDEC_NAND[1] out[0] out[8] out[17] Z[1] vdd gnd pnand3_2
XDEC_NAND[2] out[0] out[8] out[18] Z[2] vdd gnd pnand3_2
XDEC_NAND[3] out[0] out[8] out[19] Z[3] vdd gnd pnand3_2
XDEC_NAND[4] out[0] out[8] out[20] Z[4] vdd gnd pnand3_2
XDEC_NAND[5] out[0] out[8] out[21] Z[5] vdd gnd pnand3_2
XDEC_NAND[6] out[0] out[8] out[22] Z[6] vdd gnd pnand3_2
XDEC_NAND[7] out[0] out[8] out[23] Z[7] vdd gnd pnand3_2
XDEC_NAND[8] out[0] out[9] out[16] Z[8] vdd gnd pnand3_2
XDEC_NAND[9] out[0] out[9] out[17] Z[9] vdd gnd pnand3_2
XDEC_NAND[10] out[0] out[9] out[18] Z[10] vdd gnd pnand3_2
XDEC_NAND[11] out[0] out[9] out[19] Z[11] vdd gnd pnand3_2
XDEC_NAND[12] out[0] out[9] out[20] Z[12] vdd gnd pnand3_2
XDEC_NAND[13] out[0] out[9] out[21] Z[13] vdd gnd pnand3_2
XDEC_NAND[14] out[0] out[9] out[22] Z[14] vdd gnd pnand3_2
XDEC_NAND[15] out[0] out[9] out[23] Z[15] vdd gnd pnand3_2
XDEC_NAND[16] out[0] out[10] out[16] Z[16] vdd gnd pnand3_2
XDEC_NAND[17] out[0] out[10] out[17] Z[17] vdd gnd pnand3_2
XDEC_NAND[18] out[0] out[10] out[18] Z[18] vdd gnd pnand3_2
XDEC_NAND[19] out[0] out[10] out[19] Z[19] vdd gnd pnand3_2
XDEC_NAND[20] out[0] out[10] out[20] Z[20] vdd gnd pnand3_2
XDEC_NAND[21] out[0] out[10] out[21] Z[21] vdd gnd pnand3_2
XDEC_NAND[22] out[0] out[10] out[22] Z[22] vdd gnd pnand3_2
XDEC_NAND[23] out[0] out[10] out[23] Z[23] vdd gnd pnand3_2
XDEC_NAND[24] out[0] out[11] out[16] Z[24] vdd gnd pnand3_2
XDEC_NAND[25] out[0] out[11] out[17] Z[25] vdd gnd pnand3_2
XDEC_NAND[26] out[0] out[11] out[18] Z[26] vdd gnd pnand3_2
XDEC_NAND[27] out[0] out[11] out[19] Z[27] vdd gnd pnand3_2
XDEC_NAND[28] out[0] out[11] out[20] Z[28] vdd gnd pnand3_2
XDEC_NAND[29] out[0] out[11] out[21] Z[29] vdd gnd pnand3_2
XDEC_NAND[30] out[0] out[11] out[22] Z[30] vdd gnd pnand3_2
XDEC_NAND[31] out[0] out[11] out[23] Z[31] vdd gnd pnand3_2
XDEC_NAND[32] out[0] out[12] out[16] Z[32] vdd gnd pnand3_2
XDEC_NAND[33] out[0] out[12] out[17] Z[33] vdd gnd pnand3_2
XDEC_NAND[34] out[0] out[12] out[18] Z[34] vdd gnd pnand3_2
XDEC_NAND[35] out[0] out[12] out[19] Z[35] vdd gnd pnand3_2
XDEC_NAND[36] out[0] out[12] out[20] Z[36] vdd gnd pnand3_2
XDEC_NAND[37] out[0] out[12] out[21] Z[37] vdd gnd pnand3_2
XDEC_NAND[38] out[0] out[12] out[22] Z[38] vdd gnd pnand3_2
XDEC_NAND[39] out[0] out[12] out[23] Z[39] vdd gnd pnand3_2
XDEC_NAND[40] out[0] out[13] out[16] Z[40] vdd gnd pnand3_2
XDEC_NAND[41] out[0] out[13] out[17] Z[41] vdd gnd pnand3_2
XDEC_NAND[42] out[0] out[13] out[18] Z[42] vdd gnd pnand3_2
XDEC_NAND[43] out[0] out[13] out[19] Z[43] vdd gnd pnand3_2
XDEC_NAND[44] out[0] out[13] out[20] Z[44] vdd gnd pnand3_2
XDEC_NAND[45] out[0] out[13] out[21] Z[45] vdd gnd pnand3_2
XDEC_NAND[46] out[0] out[13] out[22] Z[46] vdd gnd pnand3_2
XDEC_NAND[47] out[0] out[13] out[23] Z[47] vdd gnd pnand3_2
XDEC_NAND[48] out[0] out[14] out[16] Z[48] vdd gnd pnand3_2
XDEC_NAND[49] out[0] out[14] out[17] Z[49] vdd gnd pnand3_2
XDEC_NAND[50] out[0] out[14] out[18] Z[50] vdd gnd pnand3_2
XDEC_NAND[51] out[0] out[14] out[19] Z[51] vdd gnd pnand3_2
XDEC_NAND[52] out[0] out[14] out[20] Z[52] vdd gnd pnand3_2
XDEC_NAND[53] out[0] out[14] out[21] Z[53] vdd gnd pnand3_2
XDEC_NAND[54] out[0] out[14] out[22] Z[54] vdd gnd pnand3_2
XDEC_NAND[55] out[0] out[14] out[23] Z[55] vdd gnd pnand3_2
XDEC_NAND[56] out[0] out[15] out[16] Z[56] vdd gnd pnand3_2
XDEC_NAND[57] out[0] out[15] out[17] Z[57] vdd gnd pnand3_2
XDEC_NAND[58] out[0] out[15] out[18] Z[58] vdd gnd pnand3_2
XDEC_NAND[59] out[0] out[15] out[19] Z[59] vdd gnd pnand3_2
XDEC_NAND[60] out[0] out[15] out[20] Z[60] vdd gnd pnand3_2
XDEC_NAND[61] out[0] out[15] out[21] Z[61] vdd gnd pnand3_2
XDEC_NAND[62] out[0] out[15] out[22] Z[62] vdd gnd pnand3_2
XDEC_NAND[63] out[0] out[15] out[23] Z[63] vdd gnd pnand3_2
XDEC_NAND[64] out[1] out[8] out[16] Z[64] vdd gnd pnand3_2
XDEC_NAND[65] out[1] out[8] out[17] Z[65] vdd gnd pnand3_2
XDEC_NAND[66] out[1] out[8] out[18] Z[66] vdd gnd pnand3_2
XDEC_NAND[67] out[1] out[8] out[19] Z[67] vdd gnd pnand3_2
XDEC_NAND[68] out[1] out[8] out[20] Z[68] vdd gnd pnand3_2
XDEC_NAND[69] out[1] out[8] out[21] Z[69] vdd gnd pnand3_2
XDEC_NAND[70] out[1] out[8] out[22] Z[70] vdd gnd pnand3_2
XDEC_NAND[71] out[1] out[8] out[23] Z[71] vdd gnd pnand3_2
XDEC_NAND[72] out[1] out[9] out[16] Z[72] vdd gnd pnand3_2
XDEC_NAND[73] out[1] out[9] out[17] Z[73] vdd gnd pnand3_2
XDEC_NAND[74] out[1] out[9] out[18] Z[74] vdd gnd pnand3_2
XDEC_NAND[75] out[1] out[9] out[19] Z[75] vdd gnd pnand3_2
XDEC_NAND[76] out[1] out[9] out[20] Z[76] vdd gnd pnand3_2
XDEC_NAND[77] out[1] out[9] out[21] Z[77] vdd gnd pnand3_2
XDEC_NAND[78] out[1] out[9] out[22] Z[78] vdd gnd pnand3_2
XDEC_NAND[79] out[1] out[9] out[23] Z[79] vdd gnd pnand3_2
XDEC_NAND[80] out[1] out[10] out[16] Z[80] vdd gnd pnand3_2
XDEC_NAND[81] out[1] out[10] out[17] Z[81] vdd gnd pnand3_2
XDEC_NAND[82] out[1] out[10] out[18] Z[82] vdd gnd pnand3_2
XDEC_NAND[83] out[1] out[10] out[19] Z[83] vdd gnd pnand3_2
XDEC_NAND[84] out[1] out[10] out[20] Z[84] vdd gnd pnand3_2
XDEC_NAND[85] out[1] out[10] out[21] Z[85] vdd gnd pnand3_2
XDEC_NAND[86] out[1] out[10] out[22] Z[86] vdd gnd pnand3_2
XDEC_NAND[87] out[1] out[10] out[23] Z[87] vdd gnd pnand3_2
XDEC_NAND[88] out[1] out[11] out[16] Z[88] vdd gnd pnand3_2
XDEC_NAND[89] out[1] out[11] out[17] Z[89] vdd gnd pnand3_2
XDEC_NAND[90] out[1] out[11] out[18] Z[90] vdd gnd pnand3_2
XDEC_NAND[91] out[1] out[11] out[19] Z[91] vdd gnd pnand3_2
XDEC_NAND[92] out[1] out[11] out[20] Z[92] vdd gnd pnand3_2
XDEC_NAND[93] out[1] out[11] out[21] Z[93] vdd gnd pnand3_2
XDEC_NAND[94] out[1] out[11] out[22] Z[94] vdd gnd pnand3_2
XDEC_NAND[95] out[1] out[11] out[23] Z[95] vdd gnd pnand3_2
XDEC_NAND[96] out[1] out[12] out[16] Z[96] vdd gnd pnand3_2
XDEC_NAND[97] out[1] out[12] out[17] Z[97] vdd gnd pnand3_2
XDEC_NAND[98] out[1] out[12] out[18] Z[98] vdd gnd pnand3_2
XDEC_NAND[99] out[1] out[12] out[19] Z[99] vdd gnd pnand3_2
XDEC_NAND[100] out[1] out[12] out[20] Z[100] vdd gnd pnand3_2
XDEC_NAND[101] out[1] out[12] out[21] Z[101] vdd gnd pnand3_2
XDEC_NAND[102] out[1] out[12] out[22] Z[102] vdd gnd pnand3_2
XDEC_NAND[103] out[1] out[12] out[23] Z[103] vdd gnd pnand3_2
XDEC_NAND[104] out[1] out[13] out[16] Z[104] vdd gnd pnand3_2
XDEC_NAND[105] out[1] out[13] out[17] Z[105] vdd gnd pnand3_2
XDEC_NAND[106] out[1] out[13] out[18] Z[106] vdd gnd pnand3_2
XDEC_NAND[107] out[1] out[13] out[19] Z[107] vdd gnd pnand3_2
XDEC_NAND[108] out[1] out[13] out[20] Z[108] vdd gnd pnand3_2
XDEC_NAND[109] out[1] out[13] out[21] Z[109] vdd gnd pnand3_2
XDEC_NAND[110] out[1] out[13] out[22] Z[110] vdd gnd pnand3_2
XDEC_NAND[111] out[1] out[13] out[23] Z[111] vdd gnd pnand3_2
XDEC_NAND[112] out[1] out[14] out[16] Z[112] vdd gnd pnand3_2
XDEC_NAND[113] out[1] out[14] out[17] Z[113] vdd gnd pnand3_2
XDEC_NAND[114] out[1] out[14] out[18] Z[114] vdd gnd pnand3_2
XDEC_NAND[115] out[1] out[14] out[19] Z[115] vdd gnd pnand3_2
XDEC_NAND[116] out[1] out[14] out[20] Z[116] vdd gnd pnand3_2
XDEC_NAND[117] out[1] out[14] out[21] Z[117] vdd gnd pnand3_2
XDEC_NAND[118] out[1] out[14] out[22] Z[118] vdd gnd pnand3_2
XDEC_NAND[119] out[1] out[14] out[23] Z[119] vdd gnd pnand3_2
XDEC_NAND[120] out[1] out[15] out[16] Z[120] vdd gnd pnand3_2
XDEC_NAND[121] out[1] out[15] out[17] Z[121] vdd gnd pnand3_2
XDEC_NAND[122] out[1] out[15] out[18] Z[122] vdd gnd pnand3_2
XDEC_NAND[123] out[1] out[15] out[19] Z[123] vdd gnd pnand3_2
XDEC_NAND[124] out[1] out[15] out[20] Z[124] vdd gnd pnand3_2
XDEC_NAND[125] out[1] out[15] out[21] Z[125] vdd gnd pnand3_2
XDEC_NAND[126] out[1] out[15] out[22] Z[126] vdd gnd pnand3_2
XDEC_NAND[127] out[1] out[15] out[23] Z[127] vdd gnd pnand3_2
XDEC_NAND[128] out[2] out[8] out[16] Z[128] vdd gnd pnand3_2
XDEC_NAND[129] out[2] out[8] out[17] Z[129] vdd gnd pnand3_2
XDEC_NAND[130] out[2] out[8] out[18] Z[130] vdd gnd pnand3_2
XDEC_NAND[131] out[2] out[8] out[19] Z[131] vdd gnd pnand3_2
XDEC_NAND[132] out[2] out[8] out[20] Z[132] vdd gnd pnand3_2
XDEC_NAND[133] out[2] out[8] out[21] Z[133] vdd gnd pnand3_2
XDEC_NAND[134] out[2] out[8] out[22] Z[134] vdd gnd pnand3_2
XDEC_NAND[135] out[2] out[8] out[23] Z[135] vdd gnd pnand3_2
XDEC_NAND[136] out[2] out[9] out[16] Z[136] vdd gnd pnand3_2
XDEC_NAND[137] out[2] out[9] out[17] Z[137] vdd gnd pnand3_2
XDEC_NAND[138] out[2] out[9] out[18] Z[138] vdd gnd pnand3_2
XDEC_NAND[139] out[2] out[9] out[19] Z[139] vdd gnd pnand3_2
XDEC_NAND[140] out[2] out[9] out[20] Z[140] vdd gnd pnand3_2
XDEC_NAND[141] out[2] out[9] out[21] Z[141] vdd gnd pnand3_2
XDEC_NAND[142] out[2] out[9] out[22] Z[142] vdd gnd pnand3_2
XDEC_NAND[143] out[2] out[9] out[23] Z[143] vdd gnd pnand3_2
XDEC_NAND[144] out[2] out[10] out[16] Z[144] vdd gnd pnand3_2
XDEC_NAND[145] out[2] out[10] out[17] Z[145] vdd gnd pnand3_2
XDEC_NAND[146] out[2] out[10] out[18] Z[146] vdd gnd pnand3_2
XDEC_NAND[147] out[2] out[10] out[19] Z[147] vdd gnd pnand3_2
XDEC_NAND[148] out[2] out[10] out[20] Z[148] vdd gnd pnand3_2
XDEC_NAND[149] out[2] out[10] out[21] Z[149] vdd gnd pnand3_2
XDEC_NAND[150] out[2] out[10] out[22] Z[150] vdd gnd pnand3_2
XDEC_NAND[151] out[2] out[10] out[23] Z[151] vdd gnd pnand3_2
XDEC_NAND[152] out[2] out[11] out[16] Z[152] vdd gnd pnand3_2
XDEC_NAND[153] out[2] out[11] out[17] Z[153] vdd gnd pnand3_2
XDEC_NAND[154] out[2] out[11] out[18] Z[154] vdd gnd pnand3_2
XDEC_NAND[155] out[2] out[11] out[19] Z[155] vdd gnd pnand3_2
XDEC_NAND[156] out[2] out[11] out[20] Z[156] vdd gnd pnand3_2
XDEC_NAND[157] out[2] out[11] out[21] Z[157] vdd gnd pnand3_2
XDEC_NAND[158] out[2] out[11] out[22] Z[158] vdd gnd pnand3_2
XDEC_NAND[159] out[2] out[11] out[23] Z[159] vdd gnd pnand3_2
XDEC_NAND[160] out[2] out[12] out[16] Z[160] vdd gnd pnand3_2
XDEC_NAND[161] out[2] out[12] out[17] Z[161] vdd gnd pnand3_2
XDEC_NAND[162] out[2] out[12] out[18] Z[162] vdd gnd pnand3_2
XDEC_NAND[163] out[2] out[12] out[19] Z[163] vdd gnd pnand3_2
XDEC_NAND[164] out[2] out[12] out[20] Z[164] vdd gnd pnand3_2
XDEC_NAND[165] out[2] out[12] out[21] Z[165] vdd gnd pnand3_2
XDEC_NAND[166] out[2] out[12] out[22] Z[166] vdd gnd pnand3_2
XDEC_NAND[167] out[2] out[12] out[23] Z[167] vdd gnd pnand3_2
XDEC_NAND[168] out[2] out[13] out[16] Z[168] vdd gnd pnand3_2
XDEC_NAND[169] out[2] out[13] out[17] Z[169] vdd gnd pnand3_2
XDEC_NAND[170] out[2] out[13] out[18] Z[170] vdd gnd pnand3_2
XDEC_NAND[171] out[2] out[13] out[19] Z[171] vdd gnd pnand3_2
XDEC_NAND[172] out[2] out[13] out[20] Z[172] vdd gnd pnand3_2
XDEC_NAND[173] out[2] out[13] out[21] Z[173] vdd gnd pnand3_2
XDEC_NAND[174] out[2] out[13] out[22] Z[174] vdd gnd pnand3_2
XDEC_NAND[175] out[2] out[13] out[23] Z[175] vdd gnd pnand3_2
XDEC_NAND[176] out[2] out[14] out[16] Z[176] vdd gnd pnand3_2
XDEC_NAND[177] out[2] out[14] out[17] Z[177] vdd gnd pnand3_2
XDEC_NAND[178] out[2] out[14] out[18] Z[178] vdd gnd pnand3_2
XDEC_NAND[179] out[2] out[14] out[19] Z[179] vdd gnd pnand3_2
XDEC_NAND[180] out[2] out[14] out[20] Z[180] vdd gnd pnand3_2
XDEC_NAND[181] out[2] out[14] out[21] Z[181] vdd gnd pnand3_2
XDEC_NAND[182] out[2] out[14] out[22] Z[182] vdd gnd pnand3_2
XDEC_NAND[183] out[2] out[14] out[23] Z[183] vdd gnd pnand3_2
XDEC_NAND[184] out[2] out[15] out[16] Z[184] vdd gnd pnand3_2
XDEC_NAND[185] out[2] out[15] out[17] Z[185] vdd gnd pnand3_2
XDEC_NAND[186] out[2] out[15] out[18] Z[186] vdd gnd pnand3_2
XDEC_NAND[187] out[2] out[15] out[19] Z[187] vdd gnd pnand3_2
XDEC_NAND[188] out[2] out[15] out[20] Z[188] vdd gnd pnand3_2
XDEC_NAND[189] out[2] out[15] out[21] Z[189] vdd gnd pnand3_2
XDEC_NAND[190] out[2] out[15] out[22] Z[190] vdd gnd pnand3_2
XDEC_NAND[191] out[2] out[15] out[23] Z[191] vdd gnd pnand3_2
XDEC_NAND[192] out[3] out[8] out[16] Z[192] vdd gnd pnand3_2
XDEC_NAND[193] out[3] out[8] out[17] Z[193] vdd gnd pnand3_2
XDEC_NAND[194] out[3] out[8] out[18] Z[194] vdd gnd pnand3_2
XDEC_NAND[195] out[3] out[8] out[19] Z[195] vdd gnd pnand3_2
XDEC_NAND[196] out[3] out[8] out[20] Z[196] vdd gnd pnand3_2
XDEC_NAND[197] out[3] out[8] out[21] Z[197] vdd gnd pnand3_2
XDEC_NAND[198] out[3] out[8] out[22] Z[198] vdd gnd pnand3_2
XDEC_NAND[199] out[3] out[8] out[23] Z[199] vdd gnd pnand3_2
XDEC_NAND[200] out[3] out[9] out[16] Z[200] vdd gnd pnand3_2
XDEC_NAND[201] out[3] out[9] out[17] Z[201] vdd gnd pnand3_2
XDEC_NAND[202] out[3] out[9] out[18] Z[202] vdd gnd pnand3_2
XDEC_NAND[203] out[3] out[9] out[19] Z[203] vdd gnd pnand3_2
XDEC_NAND[204] out[3] out[9] out[20] Z[204] vdd gnd pnand3_2
XDEC_NAND[205] out[3] out[9] out[21] Z[205] vdd gnd pnand3_2
XDEC_NAND[206] out[3] out[9] out[22] Z[206] vdd gnd pnand3_2
XDEC_NAND[207] out[3] out[9] out[23] Z[207] vdd gnd pnand3_2
XDEC_NAND[208] out[3] out[10] out[16] Z[208] vdd gnd pnand3_2
XDEC_NAND[209] out[3] out[10] out[17] Z[209] vdd gnd pnand3_2
XDEC_NAND[210] out[3] out[10] out[18] Z[210] vdd gnd pnand3_2
XDEC_NAND[211] out[3] out[10] out[19] Z[211] vdd gnd pnand3_2
XDEC_NAND[212] out[3] out[10] out[20] Z[212] vdd gnd pnand3_2
XDEC_NAND[213] out[3] out[10] out[21] Z[213] vdd gnd pnand3_2
XDEC_NAND[214] out[3] out[10] out[22] Z[214] vdd gnd pnand3_2
XDEC_NAND[215] out[3] out[10] out[23] Z[215] vdd gnd pnand3_2
XDEC_NAND[216] out[3] out[11] out[16] Z[216] vdd gnd pnand3_2
XDEC_NAND[217] out[3] out[11] out[17] Z[217] vdd gnd pnand3_2
XDEC_NAND[218] out[3] out[11] out[18] Z[218] vdd gnd pnand3_2
XDEC_NAND[219] out[3] out[11] out[19] Z[219] vdd gnd pnand3_2
XDEC_NAND[220] out[3] out[11] out[20] Z[220] vdd gnd pnand3_2
XDEC_NAND[221] out[3] out[11] out[21] Z[221] vdd gnd pnand3_2
XDEC_NAND[222] out[3] out[11] out[22] Z[222] vdd gnd pnand3_2
XDEC_NAND[223] out[3] out[11] out[23] Z[223] vdd gnd pnand3_2
XDEC_NAND[224] out[3] out[12] out[16] Z[224] vdd gnd pnand3_2
XDEC_NAND[225] out[3] out[12] out[17] Z[225] vdd gnd pnand3_2
XDEC_NAND[226] out[3] out[12] out[18] Z[226] vdd gnd pnand3_2
XDEC_NAND[227] out[3] out[12] out[19] Z[227] vdd gnd pnand3_2
XDEC_NAND[228] out[3] out[12] out[20] Z[228] vdd gnd pnand3_2
XDEC_NAND[229] out[3] out[12] out[21] Z[229] vdd gnd pnand3_2
XDEC_NAND[230] out[3] out[12] out[22] Z[230] vdd gnd pnand3_2
XDEC_NAND[231] out[3] out[12] out[23] Z[231] vdd gnd pnand3_2
XDEC_NAND[232] out[3] out[13] out[16] Z[232] vdd gnd pnand3_2
XDEC_NAND[233] out[3] out[13] out[17] Z[233] vdd gnd pnand3_2
XDEC_NAND[234] out[3] out[13] out[18] Z[234] vdd gnd pnand3_2
XDEC_NAND[235] out[3] out[13] out[19] Z[235] vdd gnd pnand3_2
XDEC_NAND[236] out[3] out[13] out[20] Z[236] vdd gnd pnand3_2
XDEC_NAND[237] out[3] out[13] out[21] Z[237] vdd gnd pnand3_2
XDEC_NAND[238] out[3] out[13] out[22] Z[238] vdd gnd pnand3_2
XDEC_NAND[239] out[3] out[13] out[23] Z[239] vdd gnd pnand3_2
XDEC_NAND[240] out[3] out[14] out[16] Z[240] vdd gnd pnand3_2
XDEC_NAND[241] out[3] out[14] out[17] Z[241] vdd gnd pnand3_2
XDEC_NAND[242] out[3] out[14] out[18] Z[242] vdd gnd pnand3_2
XDEC_NAND[243] out[3] out[14] out[19] Z[243] vdd gnd pnand3_2
XDEC_NAND[244] out[3] out[14] out[20] Z[244] vdd gnd pnand3_2
XDEC_NAND[245] out[3] out[14] out[21] Z[245] vdd gnd pnand3_2
XDEC_NAND[246] out[3] out[14] out[22] Z[246] vdd gnd pnand3_2
XDEC_NAND[247] out[3] out[14] out[23] Z[247] vdd gnd pnand3_2
XDEC_NAND[248] out[3] out[15] out[16] Z[248] vdd gnd pnand3_2
XDEC_NAND[249] out[3] out[15] out[17] Z[249] vdd gnd pnand3_2
XDEC_NAND[250] out[3] out[15] out[18] Z[250] vdd gnd pnand3_2
XDEC_NAND[251] out[3] out[15] out[19] Z[251] vdd gnd pnand3_2
XDEC_NAND[252] out[3] out[15] out[20] Z[252] vdd gnd pnand3_2
XDEC_NAND[253] out[3] out[15] out[21] Z[253] vdd gnd pnand3_2
XDEC_NAND[254] out[3] out[15] out[22] Z[254] vdd gnd pnand3_2
XDEC_NAND[255] out[3] out[15] out[23] Z[255] vdd gnd pnand3_2
XDEC_NAND[256] out[4] out[8] out[16] Z[256] vdd gnd pnand3_2
XDEC_NAND[257] out[4] out[8] out[17] Z[257] vdd gnd pnand3_2
XDEC_NAND[258] out[4] out[8] out[18] Z[258] vdd gnd pnand3_2
XDEC_NAND[259] out[4] out[8] out[19] Z[259] vdd gnd pnand3_2
XDEC_NAND[260] out[4] out[8] out[20] Z[260] vdd gnd pnand3_2
XDEC_NAND[261] out[4] out[8] out[21] Z[261] vdd gnd pnand3_2
XDEC_NAND[262] out[4] out[8] out[22] Z[262] vdd gnd pnand3_2
XDEC_NAND[263] out[4] out[8] out[23] Z[263] vdd gnd pnand3_2
XDEC_NAND[264] out[4] out[9] out[16] Z[264] vdd gnd pnand3_2
XDEC_NAND[265] out[4] out[9] out[17] Z[265] vdd gnd pnand3_2
XDEC_NAND[266] out[4] out[9] out[18] Z[266] vdd gnd pnand3_2
XDEC_NAND[267] out[4] out[9] out[19] Z[267] vdd gnd pnand3_2
XDEC_NAND[268] out[4] out[9] out[20] Z[268] vdd gnd pnand3_2
XDEC_NAND[269] out[4] out[9] out[21] Z[269] vdd gnd pnand3_2
XDEC_NAND[270] out[4] out[9] out[22] Z[270] vdd gnd pnand3_2
XDEC_NAND[271] out[4] out[9] out[23] Z[271] vdd gnd pnand3_2
XDEC_NAND[272] out[4] out[10] out[16] Z[272] vdd gnd pnand3_2
XDEC_NAND[273] out[4] out[10] out[17] Z[273] vdd gnd pnand3_2
XDEC_NAND[274] out[4] out[10] out[18] Z[274] vdd gnd pnand3_2
XDEC_NAND[275] out[4] out[10] out[19] Z[275] vdd gnd pnand3_2
XDEC_NAND[276] out[4] out[10] out[20] Z[276] vdd gnd pnand3_2
XDEC_NAND[277] out[4] out[10] out[21] Z[277] vdd gnd pnand3_2
XDEC_NAND[278] out[4] out[10] out[22] Z[278] vdd gnd pnand3_2
XDEC_NAND[279] out[4] out[10] out[23] Z[279] vdd gnd pnand3_2
XDEC_NAND[280] out[4] out[11] out[16] Z[280] vdd gnd pnand3_2
XDEC_NAND[281] out[4] out[11] out[17] Z[281] vdd gnd pnand3_2
XDEC_NAND[282] out[4] out[11] out[18] Z[282] vdd gnd pnand3_2
XDEC_NAND[283] out[4] out[11] out[19] Z[283] vdd gnd pnand3_2
XDEC_NAND[284] out[4] out[11] out[20] Z[284] vdd gnd pnand3_2
XDEC_NAND[285] out[4] out[11] out[21] Z[285] vdd gnd pnand3_2
XDEC_NAND[286] out[4] out[11] out[22] Z[286] vdd gnd pnand3_2
XDEC_NAND[287] out[4] out[11] out[23] Z[287] vdd gnd pnand3_2
XDEC_NAND[288] out[4] out[12] out[16] Z[288] vdd gnd pnand3_2
XDEC_NAND[289] out[4] out[12] out[17] Z[289] vdd gnd pnand3_2
XDEC_NAND[290] out[4] out[12] out[18] Z[290] vdd gnd pnand3_2
XDEC_NAND[291] out[4] out[12] out[19] Z[291] vdd gnd pnand3_2
XDEC_NAND[292] out[4] out[12] out[20] Z[292] vdd gnd pnand3_2
XDEC_NAND[293] out[4] out[12] out[21] Z[293] vdd gnd pnand3_2
XDEC_NAND[294] out[4] out[12] out[22] Z[294] vdd gnd pnand3_2
XDEC_NAND[295] out[4] out[12] out[23] Z[295] vdd gnd pnand3_2
XDEC_NAND[296] out[4] out[13] out[16] Z[296] vdd gnd pnand3_2
XDEC_NAND[297] out[4] out[13] out[17] Z[297] vdd gnd pnand3_2
XDEC_NAND[298] out[4] out[13] out[18] Z[298] vdd gnd pnand3_2
XDEC_NAND[299] out[4] out[13] out[19] Z[299] vdd gnd pnand3_2
XDEC_NAND[300] out[4] out[13] out[20] Z[300] vdd gnd pnand3_2
XDEC_NAND[301] out[4] out[13] out[21] Z[301] vdd gnd pnand3_2
XDEC_NAND[302] out[4] out[13] out[22] Z[302] vdd gnd pnand3_2
XDEC_NAND[303] out[4] out[13] out[23] Z[303] vdd gnd pnand3_2
XDEC_NAND[304] out[4] out[14] out[16] Z[304] vdd gnd pnand3_2
XDEC_NAND[305] out[4] out[14] out[17] Z[305] vdd gnd pnand3_2
XDEC_NAND[306] out[4] out[14] out[18] Z[306] vdd gnd pnand3_2
XDEC_NAND[307] out[4] out[14] out[19] Z[307] vdd gnd pnand3_2
XDEC_NAND[308] out[4] out[14] out[20] Z[308] vdd gnd pnand3_2
XDEC_NAND[309] out[4] out[14] out[21] Z[309] vdd gnd pnand3_2
XDEC_NAND[310] out[4] out[14] out[22] Z[310] vdd gnd pnand3_2
XDEC_NAND[311] out[4] out[14] out[23] Z[311] vdd gnd pnand3_2
XDEC_NAND[312] out[4] out[15] out[16] Z[312] vdd gnd pnand3_2
XDEC_NAND[313] out[4] out[15] out[17] Z[313] vdd gnd pnand3_2
XDEC_NAND[314] out[4] out[15] out[18] Z[314] vdd gnd pnand3_2
XDEC_NAND[315] out[4] out[15] out[19] Z[315] vdd gnd pnand3_2
XDEC_NAND[316] out[4] out[15] out[20] Z[316] vdd gnd pnand3_2
XDEC_NAND[317] out[4] out[15] out[21] Z[317] vdd gnd pnand3_2
XDEC_NAND[318] out[4] out[15] out[22] Z[318] vdd gnd pnand3_2
XDEC_NAND[319] out[4] out[15] out[23] Z[319] vdd gnd pnand3_2
XDEC_NAND[320] out[5] out[8] out[16] Z[320] vdd gnd pnand3_2
XDEC_NAND[321] out[5] out[8] out[17] Z[321] vdd gnd pnand3_2
XDEC_NAND[322] out[5] out[8] out[18] Z[322] vdd gnd pnand3_2
XDEC_NAND[323] out[5] out[8] out[19] Z[323] vdd gnd pnand3_2
XDEC_NAND[324] out[5] out[8] out[20] Z[324] vdd gnd pnand3_2
XDEC_NAND[325] out[5] out[8] out[21] Z[325] vdd gnd pnand3_2
XDEC_NAND[326] out[5] out[8] out[22] Z[326] vdd gnd pnand3_2
XDEC_NAND[327] out[5] out[8] out[23] Z[327] vdd gnd pnand3_2
XDEC_NAND[328] out[5] out[9] out[16] Z[328] vdd gnd pnand3_2
XDEC_NAND[329] out[5] out[9] out[17] Z[329] vdd gnd pnand3_2
XDEC_NAND[330] out[5] out[9] out[18] Z[330] vdd gnd pnand3_2
XDEC_NAND[331] out[5] out[9] out[19] Z[331] vdd gnd pnand3_2
XDEC_NAND[332] out[5] out[9] out[20] Z[332] vdd gnd pnand3_2
XDEC_NAND[333] out[5] out[9] out[21] Z[333] vdd gnd pnand3_2
XDEC_NAND[334] out[5] out[9] out[22] Z[334] vdd gnd pnand3_2
XDEC_NAND[335] out[5] out[9] out[23] Z[335] vdd gnd pnand3_2
XDEC_NAND[336] out[5] out[10] out[16] Z[336] vdd gnd pnand3_2
XDEC_NAND[337] out[5] out[10] out[17] Z[337] vdd gnd pnand3_2
XDEC_NAND[338] out[5] out[10] out[18] Z[338] vdd gnd pnand3_2
XDEC_NAND[339] out[5] out[10] out[19] Z[339] vdd gnd pnand3_2
XDEC_NAND[340] out[5] out[10] out[20] Z[340] vdd gnd pnand3_2
XDEC_NAND[341] out[5] out[10] out[21] Z[341] vdd gnd pnand3_2
XDEC_NAND[342] out[5] out[10] out[22] Z[342] vdd gnd pnand3_2
XDEC_NAND[343] out[5] out[10] out[23] Z[343] vdd gnd pnand3_2
XDEC_NAND[344] out[5] out[11] out[16] Z[344] vdd gnd pnand3_2
XDEC_NAND[345] out[5] out[11] out[17] Z[345] vdd gnd pnand3_2
XDEC_NAND[346] out[5] out[11] out[18] Z[346] vdd gnd pnand3_2
XDEC_NAND[347] out[5] out[11] out[19] Z[347] vdd gnd pnand3_2
XDEC_NAND[348] out[5] out[11] out[20] Z[348] vdd gnd pnand3_2
XDEC_NAND[349] out[5] out[11] out[21] Z[349] vdd gnd pnand3_2
XDEC_NAND[350] out[5] out[11] out[22] Z[350] vdd gnd pnand3_2
XDEC_NAND[351] out[5] out[11] out[23] Z[351] vdd gnd pnand3_2
XDEC_NAND[352] out[5] out[12] out[16] Z[352] vdd gnd pnand3_2
XDEC_NAND[353] out[5] out[12] out[17] Z[353] vdd gnd pnand3_2
XDEC_NAND[354] out[5] out[12] out[18] Z[354] vdd gnd pnand3_2
XDEC_NAND[355] out[5] out[12] out[19] Z[355] vdd gnd pnand3_2
XDEC_NAND[356] out[5] out[12] out[20] Z[356] vdd gnd pnand3_2
XDEC_NAND[357] out[5] out[12] out[21] Z[357] vdd gnd pnand3_2
XDEC_NAND[358] out[5] out[12] out[22] Z[358] vdd gnd pnand3_2
XDEC_NAND[359] out[5] out[12] out[23] Z[359] vdd gnd pnand3_2
XDEC_NAND[360] out[5] out[13] out[16] Z[360] vdd gnd pnand3_2
XDEC_NAND[361] out[5] out[13] out[17] Z[361] vdd gnd pnand3_2
XDEC_NAND[362] out[5] out[13] out[18] Z[362] vdd gnd pnand3_2
XDEC_NAND[363] out[5] out[13] out[19] Z[363] vdd gnd pnand3_2
XDEC_NAND[364] out[5] out[13] out[20] Z[364] vdd gnd pnand3_2
XDEC_NAND[365] out[5] out[13] out[21] Z[365] vdd gnd pnand3_2
XDEC_NAND[366] out[5] out[13] out[22] Z[366] vdd gnd pnand3_2
XDEC_NAND[367] out[5] out[13] out[23] Z[367] vdd gnd pnand3_2
XDEC_NAND[368] out[5] out[14] out[16] Z[368] vdd gnd pnand3_2
XDEC_NAND[369] out[5] out[14] out[17] Z[369] vdd gnd pnand3_2
XDEC_NAND[370] out[5] out[14] out[18] Z[370] vdd gnd pnand3_2
XDEC_NAND[371] out[5] out[14] out[19] Z[371] vdd gnd pnand3_2
XDEC_NAND[372] out[5] out[14] out[20] Z[372] vdd gnd pnand3_2
XDEC_NAND[373] out[5] out[14] out[21] Z[373] vdd gnd pnand3_2
XDEC_NAND[374] out[5] out[14] out[22] Z[374] vdd gnd pnand3_2
XDEC_NAND[375] out[5] out[14] out[23] Z[375] vdd gnd pnand3_2
XDEC_NAND[376] out[5] out[15] out[16] Z[376] vdd gnd pnand3_2
XDEC_NAND[377] out[5] out[15] out[17] Z[377] vdd gnd pnand3_2
XDEC_NAND[378] out[5] out[15] out[18] Z[378] vdd gnd pnand3_2
XDEC_NAND[379] out[5] out[15] out[19] Z[379] vdd gnd pnand3_2
XDEC_NAND[380] out[5] out[15] out[20] Z[380] vdd gnd pnand3_2
XDEC_NAND[381] out[5] out[15] out[21] Z[381] vdd gnd pnand3_2
XDEC_NAND[382] out[5] out[15] out[22] Z[382] vdd gnd pnand3_2
XDEC_NAND[383] out[5] out[15] out[23] Z[383] vdd gnd pnand3_2
XDEC_NAND[384] out[6] out[8] out[16] Z[384] vdd gnd pnand3_2
XDEC_NAND[385] out[6] out[8] out[17] Z[385] vdd gnd pnand3_2
XDEC_NAND[386] out[6] out[8] out[18] Z[386] vdd gnd pnand3_2
XDEC_NAND[387] out[6] out[8] out[19] Z[387] vdd gnd pnand3_2
XDEC_NAND[388] out[6] out[8] out[20] Z[388] vdd gnd pnand3_2
XDEC_NAND[389] out[6] out[8] out[21] Z[389] vdd gnd pnand3_2
XDEC_NAND[390] out[6] out[8] out[22] Z[390] vdd gnd pnand3_2
XDEC_NAND[391] out[6] out[8] out[23] Z[391] vdd gnd pnand3_2
XDEC_NAND[392] out[6] out[9] out[16] Z[392] vdd gnd pnand3_2
XDEC_NAND[393] out[6] out[9] out[17] Z[393] vdd gnd pnand3_2
XDEC_NAND[394] out[6] out[9] out[18] Z[394] vdd gnd pnand3_2
XDEC_NAND[395] out[6] out[9] out[19] Z[395] vdd gnd pnand3_2
XDEC_NAND[396] out[6] out[9] out[20] Z[396] vdd gnd pnand3_2
XDEC_NAND[397] out[6] out[9] out[21] Z[397] vdd gnd pnand3_2
XDEC_NAND[398] out[6] out[9] out[22] Z[398] vdd gnd pnand3_2
XDEC_NAND[399] out[6] out[9] out[23] Z[399] vdd gnd pnand3_2
XDEC_NAND[400] out[6] out[10] out[16] Z[400] vdd gnd pnand3_2
XDEC_NAND[401] out[6] out[10] out[17] Z[401] vdd gnd pnand3_2
XDEC_NAND[402] out[6] out[10] out[18] Z[402] vdd gnd pnand3_2
XDEC_NAND[403] out[6] out[10] out[19] Z[403] vdd gnd pnand3_2
XDEC_NAND[404] out[6] out[10] out[20] Z[404] vdd gnd pnand3_2
XDEC_NAND[405] out[6] out[10] out[21] Z[405] vdd gnd pnand3_2
XDEC_NAND[406] out[6] out[10] out[22] Z[406] vdd gnd pnand3_2
XDEC_NAND[407] out[6] out[10] out[23] Z[407] vdd gnd pnand3_2
XDEC_NAND[408] out[6] out[11] out[16] Z[408] vdd gnd pnand3_2
XDEC_NAND[409] out[6] out[11] out[17] Z[409] vdd gnd pnand3_2
XDEC_NAND[410] out[6] out[11] out[18] Z[410] vdd gnd pnand3_2
XDEC_NAND[411] out[6] out[11] out[19] Z[411] vdd gnd pnand3_2
XDEC_NAND[412] out[6] out[11] out[20] Z[412] vdd gnd pnand3_2
XDEC_NAND[413] out[6] out[11] out[21] Z[413] vdd gnd pnand3_2
XDEC_NAND[414] out[6] out[11] out[22] Z[414] vdd gnd pnand3_2
XDEC_NAND[415] out[6] out[11] out[23] Z[415] vdd gnd pnand3_2
XDEC_NAND[416] out[6] out[12] out[16] Z[416] vdd gnd pnand3_2
XDEC_NAND[417] out[6] out[12] out[17] Z[417] vdd gnd pnand3_2
XDEC_NAND[418] out[6] out[12] out[18] Z[418] vdd gnd pnand3_2
XDEC_NAND[419] out[6] out[12] out[19] Z[419] vdd gnd pnand3_2
XDEC_NAND[420] out[6] out[12] out[20] Z[420] vdd gnd pnand3_2
XDEC_NAND[421] out[6] out[12] out[21] Z[421] vdd gnd pnand3_2
XDEC_NAND[422] out[6] out[12] out[22] Z[422] vdd gnd pnand3_2
XDEC_NAND[423] out[6] out[12] out[23] Z[423] vdd gnd pnand3_2
XDEC_NAND[424] out[6] out[13] out[16] Z[424] vdd gnd pnand3_2
XDEC_NAND[425] out[6] out[13] out[17] Z[425] vdd gnd pnand3_2
XDEC_NAND[426] out[6] out[13] out[18] Z[426] vdd gnd pnand3_2
XDEC_NAND[427] out[6] out[13] out[19] Z[427] vdd gnd pnand3_2
XDEC_NAND[428] out[6] out[13] out[20] Z[428] vdd gnd pnand3_2
XDEC_NAND[429] out[6] out[13] out[21] Z[429] vdd gnd pnand3_2
XDEC_NAND[430] out[6] out[13] out[22] Z[430] vdd gnd pnand3_2
XDEC_NAND[431] out[6] out[13] out[23] Z[431] vdd gnd pnand3_2
XDEC_NAND[432] out[6] out[14] out[16] Z[432] vdd gnd pnand3_2
XDEC_NAND[433] out[6] out[14] out[17] Z[433] vdd gnd pnand3_2
XDEC_NAND[434] out[6] out[14] out[18] Z[434] vdd gnd pnand3_2
XDEC_NAND[435] out[6] out[14] out[19] Z[435] vdd gnd pnand3_2
XDEC_NAND[436] out[6] out[14] out[20] Z[436] vdd gnd pnand3_2
XDEC_NAND[437] out[6] out[14] out[21] Z[437] vdd gnd pnand3_2
XDEC_NAND[438] out[6] out[14] out[22] Z[438] vdd gnd pnand3_2
XDEC_NAND[439] out[6] out[14] out[23] Z[439] vdd gnd pnand3_2
XDEC_NAND[440] out[6] out[15] out[16] Z[440] vdd gnd pnand3_2
XDEC_NAND[441] out[6] out[15] out[17] Z[441] vdd gnd pnand3_2
XDEC_NAND[442] out[6] out[15] out[18] Z[442] vdd gnd pnand3_2
XDEC_NAND[443] out[6] out[15] out[19] Z[443] vdd gnd pnand3_2
XDEC_NAND[444] out[6] out[15] out[20] Z[444] vdd gnd pnand3_2
XDEC_NAND[445] out[6] out[15] out[21] Z[445] vdd gnd pnand3_2
XDEC_NAND[446] out[6] out[15] out[22] Z[446] vdd gnd pnand3_2
XDEC_NAND[447] out[6] out[15] out[23] Z[447] vdd gnd pnand3_2
XDEC_NAND[448] out[7] out[8] out[16] Z[448] vdd gnd pnand3_2
XDEC_NAND[449] out[7] out[8] out[17] Z[449] vdd gnd pnand3_2
XDEC_NAND[450] out[7] out[8] out[18] Z[450] vdd gnd pnand3_2
XDEC_NAND[451] out[7] out[8] out[19] Z[451] vdd gnd pnand3_2
XDEC_NAND[452] out[7] out[8] out[20] Z[452] vdd gnd pnand3_2
XDEC_NAND[453] out[7] out[8] out[21] Z[453] vdd gnd pnand3_2
XDEC_NAND[454] out[7] out[8] out[22] Z[454] vdd gnd pnand3_2
XDEC_NAND[455] out[7] out[8] out[23] Z[455] vdd gnd pnand3_2
XDEC_NAND[456] out[7] out[9] out[16] Z[456] vdd gnd pnand3_2
XDEC_NAND[457] out[7] out[9] out[17] Z[457] vdd gnd pnand3_2
XDEC_NAND[458] out[7] out[9] out[18] Z[458] vdd gnd pnand3_2
XDEC_NAND[459] out[7] out[9] out[19] Z[459] vdd gnd pnand3_2
XDEC_NAND[460] out[7] out[9] out[20] Z[460] vdd gnd pnand3_2
XDEC_NAND[461] out[7] out[9] out[21] Z[461] vdd gnd pnand3_2
XDEC_NAND[462] out[7] out[9] out[22] Z[462] vdd gnd pnand3_2
XDEC_NAND[463] out[7] out[9] out[23] Z[463] vdd gnd pnand3_2
XDEC_NAND[464] out[7] out[10] out[16] Z[464] vdd gnd pnand3_2
XDEC_NAND[465] out[7] out[10] out[17] Z[465] vdd gnd pnand3_2
XDEC_NAND[466] out[7] out[10] out[18] Z[466] vdd gnd pnand3_2
XDEC_NAND[467] out[7] out[10] out[19] Z[467] vdd gnd pnand3_2
XDEC_NAND[468] out[7] out[10] out[20] Z[468] vdd gnd pnand3_2
XDEC_NAND[469] out[7] out[10] out[21] Z[469] vdd gnd pnand3_2
XDEC_NAND[470] out[7] out[10] out[22] Z[470] vdd gnd pnand3_2
XDEC_NAND[471] out[7] out[10] out[23] Z[471] vdd gnd pnand3_2
XDEC_NAND[472] out[7] out[11] out[16] Z[472] vdd gnd pnand3_2
XDEC_NAND[473] out[7] out[11] out[17] Z[473] vdd gnd pnand3_2
XDEC_NAND[474] out[7] out[11] out[18] Z[474] vdd gnd pnand3_2
XDEC_NAND[475] out[7] out[11] out[19] Z[475] vdd gnd pnand3_2
XDEC_NAND[476] out[7] out[11] out[20] Z[476] vdd gnd pnand3_2
XDEC_NAND[477] out[7] out[11] out[21] Z[477] vdd gnd pnand3_2
XDEC_NAND[478] out[7] out[11] out[22] Z[478] vdd gnd pnand3_2
XDEC_NAND[479] out[7] out[11] out[23] Z[479] vdd gnd pnand3_2
XDEC_NAND[480] out[7] out[12] out[16] Z[480] vdd gnd pnand3_2
XDEC_NAND[481] out[7] out[12] out[17] Z[481] vdd gnd pnand3_2
XDEC_NAND[482] out[7] out[12] out[18] Z[482] vdd gnd pnand3_2
XDEC_NAND[483] out[7] out[12] out[19] Z[483] vdd gnd pnand3_2
XDEC_NAND[484] out[7] out[12] out[20] Z[484] vdd gnd pnand3_2
XDEC_NAND[485] out[7] out[12] out[21] Z[485] vdd gnd pnand3_2
XDEC_NAND[486] out[7] out[12] out[22] Z[486] vdd gnd pnand3_2
XDEC_NAND[487] out[7] out[12] out[23] Z[487] vdd gnd pnand3_2
XDEC_NAND[488] out[7] out[13] out[16] Z[488] vdd gnd pnand3_2
XDEC_NAND[489] out[7] out[13] out[17] Z[489] vdd gnd pnand3_2
XDEC_NAND[490] out[7] out[13] out[18] Z[490] vdd gnd pnand3_2
XDEC_NAND[491] out[7] out[13] out[19] Z[491] vdd gnd pnand3_2
XDEC_NAND[492] out[7] out[13] out[20] Z[492] vdd gnd pnand3_2
XDEC_NAND[493] out[7] out[13] out[21] Z[493] vdd gnd pnand3_2
XDEC_NAND[494] out[7] out[13] out[22] Z[494] vdd gnd pnand3_2
XDEC_NAND[495] out[7] out[13] out[23] Z[495] vdd gnd pnand3_2
XDEC_NAND[496] out[7] out[14] out[16] Z[496] vdd gnd pnand3_2
XDEC_NAND[497] out[7] out[14] out[17] Z[497] vdd gnd pnand3_2
XDEC_NAND[498] out[7] out[14] out[18] Z[498] vdd gnd pnand3_2
XDEC_NAND[499] out[7] out[14] out[19] Z[499] vdd gnd pnand3_2
XDEC_NAND[500] out[7] out[14] out[20] Z[500] vdd gnd pnand3_2
XDEC_NAND[501] out[7] out[14] out[21] Z[501] vdd gnd pnand3_2
XDEC_NAND[502] out[7] out[14] out[22] Z[502] vdd gnd pnand3_2
XDEC_NAND[503] out[7] out[14] out[23] Z[503] vdd gnd pnand3_2
XDEC_NAND[504] out[7] out[15] out[16] Z[504] vdd gnd pnand3_2
XDEC_NAND[505] out[7] out[15] out[17] Z[505] vdd gnd pnand3_2
XDEC_NAND[506] out[7] out[15] out[18] Z[506] vdd gnd pnand3_2
XDEC_NAND[507] out[7] out[15] out[19] Z[507] vdd gnd pnand3_2
XDEC_NAND[508] out[7] out[15] out[20] Z[508] vdd gnd pnand3_2
XDEC_NAND[509] out[7] out[15] out[21] Z[509] vdd gnd pnand3_2
XDEC_NAND[510] out[7] out[15] out[22] Z[510] vdd gnd pnand3_2
XDEC_NAND[511] out[7] out[15] out[23] Z[511] vdd gnd pnand3_2
XDEC_INV_[0] Z[0] decode[0] vdd gnd pinv_8
XDEC_INV_[1] Z[1] decode[1] vdd gnd pinv_8
XDEC_INV_[2] Z[2] decode[2] vdd gnd pinv_8
XDEC_INV_[3] Z[3] decode[3] vdd gnd pinv_8
XDEC_INV_[4] Z[4] decode[4] vdd gnd pinv_8
XDEC_INV_[5] Z[5] decode[5] vdd gnd pinv_8
XDEC_INV_[6] Z[6] decode[6] vdd gnd pinv_8
XDEC_INV_[7] Z[7] decode[7] vdd gnd pinv_8
XDEC_INV_[8] Z[8] decode[8] vdd gnd pinv_8
XDEC_INV_[9] Z[9] decode[9] vdd gnd pinv_8
XDEC_INV_[10] Z[10] decode[10] vdd gnd pinv_8
XDEC_INV_[11] Z[11] decode[11] vdd gnd pinv_8
XDEC_INV_[12] Z[12] decode[12] vdd gnd pinv_8
XDEC_INV_[13] Z[13] decode[13] vdd gnd pinv_8
XDEC_INV_[14] Z[14] decode[14] vdd gnd pinv_8
XDEC_INV_[15] Z[15] decode[15] vdd gnd pinv_8
XDEC_INV_[16] Z[16] decode[16] vdd gnd pinv_8
XDEC_INV_[17] Z[17] decode[17] vdd gnd pinv_8
XDEC_INV_[18] Z[18] decode[18] vdd gnd pinv_8
XDEC_INV_[19] Z[19] decode[19] vdd gnd pinv_8
XDEC_INV_[20] Z[20] decode[20] vdd gnd pinv_8
XDEC_INV_[21] Z[21] decode[21] vdd gnd pinv_8
XDEC_INV_[22] Z[22] decode[22] vdd gnd pinv_8
XDEC_INV_[23] Z[23] decode[23] vdd gnd pinv_8
XDEC_INV_[24] Z[24] decode[24] vdd gnd pinv_8
XDEC_INV_[25] Z[25] decode[25] vdd gnd pinv_8
XDEC_INV_[26] Z[26] decode[26] vdd gnd pinv_8
XDEC_INV_[27] Z[27] decode[27] vdd gnd pinv_8
XDEC_INV_[28] Z[28] decode[28] vdd gnd pinv_8
XDEC_INV_[29] Z[29] decode[29] vdd gnd pinv_8
XDEC_INV_[30] Z[30] decode[30] vdd gnd pinv_8
XDEC_INV_[31] Z[31] decode[31] vdd gnd pinv_8
XDEC_INV_[32] Z[32] decode[32] vdd gnd pinv_8
XDEC_INV_[33] Z[33] decode[33] vdd gnd pinv_8
XDEC_INV_[34] Z[34] decode[34] vdd gnd pinv_8
XDEC_INV_[35] Z[35] decode[35] vdd gnd pinv_8
XDEC_INV_[36] Z[36] decode[36] vdd gnd pinv_8
XDEC_INV_[37] Z[37] decode[37] vdd gnd pinv_8
XDEC_INV_[38] Z[38] decode[38] vdd gnd pinv_8
XDEC_INV_[39] Z[39] decode[39] vdd gnd pinv_8
XDEC_INV_[40] Z[40] decode[40] vdd gnd pinv_8
XDEC_INV_[41] Z[41] decode[41] vdd gnd pinv_8
XDEC_INV_[42] Z[42] decode[42] vdd gnd pinv_8
XDEC_INV_[43] Z[43] decode[43] vdd gnd pinv_8
XDEC_INV_[44] Z[44] decode[44] vdd gnd pinv_8
XDEC_INV_[45] Z[45] decode[45] vdd gnd pinv_8
XDEC_INV_[46] Z[46] decode[46] vdd gnd pinv_8
XDEC_INV_[47] Z[47] decode[47] vdd gnd pinv_8
XDEC_INV_[48] Z[48] decode[48] vdd gnd pinv_8
XDEC_INV_[49] Z[49] decode[49] vdd gnd pinv_8
XDEC_INV_[50] Z[50] decode[50] vdd gnd pinv_8
XDEC_INV_[51] Z[51] decode[51] vdd gnd pinv_8
XDEC_INV_[52] Z[52] decode[52] vdd gnd pinv_8
XDEC_INV_[53] Z[53] decode[53] vdd gnd pinv_8
XDEC_INV_[54] Z[54] decode[54] vdd gnd pinv_8
XDEC_INV_[55] Z[55] decode[55] vdd gnd pinv_8
XDEC_INV_[56] Z[56] decode[56] vdd gnd pinv_8
XDEC_INV_[57] Z[57] decode[57] vdd gnd pinv_8
XDEC_INV_[58] Z[58] decode[58] vdd gnd pinv_8
XDEC_INV_[59] Z[59] decode[59] vdd gnd pinv_8
XDEC_INV_[60] Z[60] decode[60] vdd gnd pinv_8
XDEC_INV_[61] Z[61] decode[61] vdd gnd pinv_8
XDEC_INV_[62] Z[62] decode[62] vdd gnd pinv_8
XDEC_INV_[63] Z[63] decode[63] vdd gnd pinv_8
XDEC_INV_[64] Z[64] decode[64] vdd gnd pinv_8
XDEC_INV_[65] Z[65] decode[65] vdd gnd pinv_8
XDEC_INV_[66] Z[66] decode[66] vdd gnd pinv_8
XDEC_INV_[67] Z[67] decode[67] vdd gnd pinv_8
XDEC_INV_[68] Z[68] decode[68] vdd gnd pinv_8
XDEC_INV_[69] Z[69] decode[69] vdd gnd pinv_8
XDEC_INV_[70] Z[70] decode[70] vdd gnd pinv_8
XDEC_INV_[71] Z[71] decode[71] vdd gnd pinv_8
XDEC_INV_[72] Z[72] decode[72] vdd gnd pinv_8
XDEC_INV_[73] Z[73] decode[73] vdd gnd pinv_8
XDEC_INV_[74] Z[74] decode[74] vdd gnd pinv_8
XDEC_INV_[75] Z[75] decode[75] vdd gnd pinv_8
XDEC_INV_[76] Z[76] decode[76] vdd gnd pinv_8
XDEC_INV_[77] Z[77] decode[77] vdd gnd pinv_8
XDEC_INV_[78] Z[78] decode[78] vdd gnd pinv_8
XDEC_INV_[79] Z[79] decode[79] vdd gnd pinv_8
XDEC_INV_[80] Z[80] decode[80] vdd gnd pinv_8
XDEC_INV_[81] Z[81] decode[81] vdd gnd pinv_8
XDEC_INV_[82] Z[82] decode[82] vdd gnd pinv_8
XDEC_INV_[83] Z[83] decode[83] vdd gnd pinv_8
XDEC_INV_[84] Z[84] decode[84] vdd gnd pinv_8
XDEC_INV_[85] Z[85] decode[85] vdd gnd pinv_8
XDEC_INV_[86] Z[86] decode[86] vdd gnd pinv_8
XDEC_INV_[87] Z[87] decode[87] vdd gnd pinv_8
XDEC_INV_[88] Z[88] decode[88] vdd gnd pinv_8
XDEC_INV_[89] Z[89] decode[89] vdd gnd pinv_8
XDEC_INV_[90] Z[90] decode[90] vdd gnd pinv_8
XDEC_INV_[91] Z[91] decode[91] vdd gnd pinv_8
XDEC_INV_[92] Z[92] decode[92] vdd gnd pinv_8
XDEC_INV_[93] Z[93] decode[93] vdd gnd pinv_8
XDEC_INV_[94] Z[94] decode[94] vdd gnd pinv_8
XDEC_INV_[95] Z[95] decode[95] vdd gnd pinv_8
XDEC_INV_[96] Z[96] decode[96] vdd gnd pinv_8
XDEC_INV_[97] Z[97] decode[97] vdd gnd pinv_8
XDEC_INV_[98] Z[98] decode[98] vdd gnd pinv_8
XDEC_INV_[99] Z[99] decode[99] vdd gnd pinv_8
XDEC_INV_[100] Z[100] decode[100] vdd gnd pinv_8
XDEC_INV_[101] Z[101] decode[101] vdd gnd pinv_8
XDEC_INV_[102] Z[102] decode[102] vdd gnd pinv_8
XDEC_INV_[103] Z[103] decode[103] vdd gnd pinv_8
XDEC_INV_[104] Z[104] decode[104] vdd gnd pinv_8
XDEC_INV_[105] Z[105] decode[105] vdd gnd pinv_8
XDEC_INV_[106] Z[106] decode[106] vdd gnd pinv_8
XDEC_INV_[107] Z[107] decode[107] vdd gnd pinv_8
XDEC_INV_[108] Z[108] decode[108] vdd gnd pinv_8
XDEC_INV_[109] Z[109] decode[109] vdd gnd pinv_8
XDEC_INV_[110] Z[110] decode[110] vdd gnd pinv_8
XDEC_INV_[111] Z[111] decode[111] vdd gnd pinv_8
XDEC_INV_[112] Z[112] decode[112] vdd gnd pinv_8
XDEC_INV_[113] Z[113] decode[113] vdd gnd pinv_8
XDEC_INV_[114] Z[114] decode[114] vdd gnd pinv_8
XDEC_INV_[115] Z[115] decode[115] vdd gnd pinv_8
XDEC_INV_[116] Z[116] decode[116] vdd gnd pinv_8
XDEC_INV_[117] Z[117] decode[117] vdd gnd pinv_8
XDEC_INV_[118] Z[118] decode[118] vdd gnd pinv_8
XDEC_INV_[119] Z[119] decode[119] vdd gnd pinv_8
XDEC_INV_[120] Z[120] decode[120] vdd gnd pinv_8
XDEC_INV_[121] Z[121] decode[121] vdd gnd pinv_8
XDEC_INV_[122] Z[122] decode[122] vdd gnd pinv_8
XDEC_INV_[123] Z[123] decode[123] vdd gnd pinv_8
XDEC_INV_[124] Z[124] decode[124] vdd gnd pinv_8
XDEC_INV_[125] Z[125] decode[125] vdd gnd pinv_8
XDEC_INV_[126] Z[126] decode[126] vdd gnd pinv_8
XDEC_INV_[127] Z[127] decode[127] vdd gnd pinv_8
XDEC_INV_[128] Z[128] decode[128] vdd gnd pinv_8
XDEC_INV_[129] Z[129] decode[129] vdd gnd pinv_8
XDEC_INV_[130] Z[130] decode[130] vdd gnd pinv_8
XDEC_INV_[131] Z[131] decode[131] vdd gnd pinv_8
XDEC_INV_[132] Z[132] decode[132] vdd gnd pinv_8
XDEC_INV_[133] Z[133] decode[133] vdd gnd pinv_8
XDEC_INV_[134] Z[134] decode[134] vdd gnd pinv_8
XDEC_INV_[135] Z[135] decode[135] vdd gnd pinv_8
XDEC_INV_[136] Z[136] decode[136] vdd gnd pinv_8
XDEC_INV_[137] Z[137] decode[137] vdd gnd pinv_8
XDEC_INV_[138] Z[138] decode[138] vdd gnd pinv_8
XDEC_INV_[139] Z[139] decode[139] vdd gnd pinv_8
XDEC_INV_[140] Z[140] decode[140] vdd gnd pinv_8
XDEC_INV_[141] Z[141] decode[141] vdd gnd pinv_8
XDEC_INV_[142] Z[142] decode[142] vdd gnd pinv_8
XDEC_INV_[143] Z[143] decode[143] vdd gnd pinv_8
XDEC_INV_[144] Z[144] decode[144] vdd gnd pinv_8
XDEC_INV_[145] Z[145] decode[145] vdd gnd pinv_8
XDEC_INV_[146] Z[146] decode[146] vdd gnd pinv_8
XDEC_INV_[147] Z[147] decode[147] vdd gnd pinv_8
XDEC_INV_[148] Z[148] decode[148] vdd gnd pinv_8
XDEC_INV_[149] Z[149] decode[149] vdd gnd pinv_8
XDEC_INV_[150] Z[150] decode[150] vdd gnd pinv_8
XDEC_INV_[151] Z[151] decode[151] vdd gnd pinv_8
XDEC_INV_[152] Z[152] decode[152] vdd gnd pinv_8
XDEC_INV_[153] Z[153] decode[153] vdd gnd pinv_8
XDEC_INV_[154] Z[154] decode[154] vdd gnd pinv_8
XDEC_INV_[155] Z[155] decode[155] vdd gnd pinv_8
XDEC_INV_[156] Z[156] decode[156] vdd gnd pinv_8
XDEC_INV_[157] Z[157] decode[157] vdd gnd pinv_8
XDEC_INV_[158] Z[158] decode[158] vdd gnd pinv_8
XDEC_INV_[159] Z[159] decode[159] vdd gnd pinv_8
XDEC_INV_[160] Z[160] decode[160] vdd gnd pinv_8
XDEC_INV_[161] Z[161] decode[161] vdd gnd pinv_8
XDEC_INV_[162] Z[162] decode[162] vdd gnd pinv_8
XDEC_INV_[163] Z[163] decode[163] vdd gnd pinv_8
XDEC_INV_[164] Z[164] decode[164] vdd gnd pinv_8
XDEC_INV_[165] Z[165] decode[165] vdd gnd pinv_8
XDEC_INV_[166] Z[166] decode[166] vdd gnd pinv_8
XDEC_INV_[167] Z[167] decode[167] vdd gnd pinv_8
XDEC_INV_[168] Z[168] decode[168] vdd gnd pinv_8
XDEC_INV_[169] Z[169] decode[169] vdd gnd pinv_8
XDEC_INV_[170] Z[170] decode[170] vdd gnd pinv_8
XDEC_INV_[171] Z[171] decode[171] vdd gnd pinv_8
XDEC_INV_[172] Z[172] decode[172] vdd gnd pinv_8
XDEC_INV_[173] Z[173] decode[173] vdd gnd pinv_8
XDEC_INV_[174] Z[174] decode[174] vdd gnd pinv_8
XDEC_INV_[175] Z[175] decode[175] vdd gnd pinv_8
XDEC_INV_[176] Z[176] decode[176] vdd gnd pinv_8
XDEC_INV_[177] Z[177] decode[177] vdd gnd pinv_8
XDEC_INV_[178] Z[178] decode[178] vdd gnd pinv_8
XDEC_INV_[179] Z[179] decode[179] vdd gnd pinv_8
XDEC_INV_[180] Z[180] decode[180] vdd gnd pinv_8
XDEC_INV_[181] Z[181] decode[181] vdd gnd pinv_8
XDEC_INV_[182] Z[182] decode[182] vdd gnd pinv_8
XDEC_INV_[183] Z[183] decode[183] vdd gnd pinv_8
XDEC_INV_[184] Z[184] decode[184] vdd gnd pinv_8
XDEC_INV_[185] Z[185] decode[185] vdd gnd pinv_8
XDEC_INV_[186] Z[186] decode[186] vdd gnd pinv_8
XDEC_INV_[187] Z[187] decode[187] vdd gnd pinv_8
XDEC_INV_[188] Z[188] decode[188] vdd gnd pinv_8
XDEC_INV_[189] Z[189] decode[189] vdd gnd pinv_8
XDEC_INV_[190] Z[190] decode[190] vdd gnd pinv_8
XDEC_INV_[191] Z[191] decode[191] vdd gnd pinv_8
XDEC_INV_[192] Z[192] decode[192] vdd gnd pinv_8
XDEC_INV_[193] Z[193] decode[193] vdd gnd pinv_8
XDEC_INV_[194] Z[194] decode[194] vdd gnd pinv_8
XDEC_INV_[195] Z[195] decode[195] vdd gnd pinv_8
XDEC_INV_[196] Z[196] decode[196] vdd gnd pinv_8
XDEC_INV_[197] Z[197] decode[197] vdd gnd pinv_8
XDEC_INV_[198] Z[198] decode[198] vdd gnd pinv_8
XDEC_INV_[199] Z[199] decode[199] vdd gnd pinv_8
XDEC_INV_[200] Z[200] decode[200] vdd gnd pinv_8
XDEC_INV_[201] Z[201] decode[201] vdd gnd pinv_8
XDEC_INV_[202] Z[202] decode[202] vdd gnd pinv_8
XDEC_INV_[203] Z[203] decode[203] vdd gnd pinv_8
XDEC_INV_[204] Z[204] decode[204] vdd gnd pinv_8
XDEC_INV_[205] Z[205] decode[205] vdd gnd pinv_8
XDEC_INV_[206] Z[206] decode[206] vdd gnd pinv_8
XDEC_INV_[207] Z[207] decode[207] vdd gnd pinv_8
XDEC_INV_[208] Z[208] decode[208] vdd gnd pinv_8
XDEC_INV_[209] Z[209] decode[209] vdd gnd pinv_8
XDEC_INV_[210] Z[210] decode[210] vdd gnd pinv_8
XDEC_INV_[211] Z[211] decode[211] vdd gnd pinv_8
XDEC_INV_[212] Z[212] decode[212] vdd gnd pinv_8
XDEC_INV_[213] Z[213] decode[213] vdd gnd pinv_8
XDEC_INV_[214] Z[214] decode[214] vdd gnd pinv_8
XDEC_INV_[215] Z[215] decode[215] vdd gnd pinv_8
XDEC_INV_[216] Z[216] decode[216] vdd gnd pinv_8
XDEC_INV_[217] Z[217] decode[217] vdd gnd pinv_8
XDEC_INV_[218] Z[218] decode[218] vdd gnd pinv_8
XDEC_INV_[219] Z[219] decode[219] vdd gnd pinv_8
XDEC_INV_[220] Z[220] decode[220] vdd gnd pinv_8
XDEC_INV_[221] Z[221] decode[221] vdd gnd pinv_8
XDEC_INV_[222] Z[222] decode[222] vdd gnd pinv_8
XDEC_INV_[223] Z[223] decode[223] vdd gnd pinv_8
XDEC_INV_[224] Z[224] decode[224] vdd gnd pinv_8
XDEC_INV_[225] Z[225] decode[225] vdd gnd pinv_8
XDEC_INV_[226] Z[226] decode[226] vdd gnd pinv_8
XDEC_INV_[227] Z[227] decode[227] vdd gnd pinv_8
XDEC_INV_[228] Z[228] decode[228] vdd gnd pinv_8
XDEC_INV_[229] Z[229] decode[229] vdd gnd pinv_8
XDEC_INV_[230] Z[230] decode[230] vdd gnd pinv_8
XDEC_INV_[231] Z[231] decode[231] vdd gnd pinv_8
XDEC_INV_[232] Z[232] decode[232] vdd gnd pinv_8
XDEC_INV_[233] Z[233] decode[233] vdd gnd pinv_8
XDEC_INV_[234] Z[234] decode[234] vdd gnd pinv_8
XDEC_INV_[235] Z[235] decode[235] vdd gnd pinv_8
XDEC_INV_[236] Z[236] decode[236] vdd gnd pinv_8
XDEC_INV_[237] Z[237] decode[237] vdd gnd pinv_8
XDEC_INV_[238] Z[238] decode[238] vdd gnd pinv_8
XDEC_INV_[239] Z[239] decode[239] vdd gnd pinv_8
XDEC_INV_[240] Z[240] decode[240] vdd gnd pinv_8
XDEC_INV_[241] Z[241] decode[241] vdd gnd pinv_8
XDEC_INV_[242] Z[242] decode[242] vdd gnd pinv_8
XDEC_INV_[243] Z[243] decode[243] vdd gnd pinv_8
XDEC_INV_[244] Z[244] decode[244] vdd gnd pinv_8
XDEC_INV_[245] Z[245] decode[245] vdd gnd pinv_8
XDEC_INV_[246] Z[246] decode[246] vdd gnd pinv_8
XDEC_INV_[247] Z[247] decode[247] vdd gnd pinv_8
XDEC_INV_[248] Z[248] decode[248] vdd gnd pinv_8
XDEC_INV_[249] Z[249] decode[249] vdd gnd pinv_8
XDEC_INV_[250] Z[250] decode[250] vdd gnd pinv_8
XDEC_INV_[251] Z[251] decode[251] vdd gnd pinv_8
XDEC_INV_[252] Z[252] decode[252] vdd gnd pinv_8
XDEC_INV_[253] Z[253] decode[253] vdd gnd pinv_8
XDEC_INV_[254] Z[254] decode[254] vdd gnd pinv_8
XDEC_INV_[255] Z[255] decode[255] vdd gnd pinv_8
XDEC_INV_[256] Z[256] decode[256] vdd gnd pinv_8
XDEC_INV_[257] Z[257] decode[257] vdd gnd pinv_8
XDEC_INV_[258] Z[258] decode[258] vdd gnd pinv_8
XDEC_INV_[259] Z[259] decode[259] vdd gnd pinv_8
XDEC_INV_[260] Z[260] decode[260] vdd gnd pinv_8
XDEC_INV_[261] Z[261] decode[261] vdd gnd pinv_8
XDEC_INV_[262] Z[262] decode[262] vdd gnd pinv_8
XDEC_INV_[263] Z[263] decode[263] vdd gnd pinv_8
XDEC_INV_[264] Z[264] decode[264] vdd gnd pinv_8
XDEC_INV_[265] Z[265] decode[265] vdd gnd pinv_8
XDEC_INV_[266] Z[266] decode[266] vdd gnd pinv_8
XDEC_INV_[267] Z[267] decode[267] vdd gnd pinv_8
XDEC_INV_[268] Z[268] decode[268] vdd gnd pinv_8
XDEC_INV_[269] Z[269] decode[269] vdd gnd pinv_8
XDEC_INV_[270] Z[270] decode[270] vdd gnd pinv_8
XDEC_INV_[271] Z[271] decode[271] vdd gnd pinv_8
XDEC_INV_[272] Z[272] decode[272] vdd gnd pinv_8
XDEC_INV_[273] Z[273] decode[273] vdd gnd pinv_8
XDEC_INV_[274] Z[274] decode[274] vdd gnd pinv_8
XDEC_INV_[275] Z[275] decode[275] vdd gnd pinv_8
XDEC_INV_[276] Z[276] decode[276] vdd gnd pinv_8
XDEC_INV_[277] Z[277] decode[277] vdd gnd pinv_8
XDEC_INV_[278] Z[278] decode[278] vdd gnd pinv_8
XDEC_INV_[279] Z[279] decode[279] vdd gnd pinv_8
XDEC_INV_[280] Z[280] decode[280] vdd gnd pinv_8
XDEC_INV_[281] Z[281] decode[281] vdd gnd pinv_8
XDEC_INV_[282] Z[282] decode[282] vdd gnd pinv_8
XDEC_INV_[283] Z[283] decode[283] vdd gnd pinv_8
XDEC_INV_[284] Z[284] decode[284] vdd gnd pinv_8
XDEC_INV_[285] Z[285] decode[285] vdd gnd pinv_8
XDEC_INV_[286] Z[286] decode[286] vdd gnd pinv_8
XDEC_INV_[287] Z[287] decode[287] vdd gnd pinv_8
XDEC_INV_[288] Z[288] decode[288] vdd gnd pinv_8
XDEC_INV_[289] Z[289] decode[289] vdd gnd pinv_8
XDEC_INV_[290] Z[290] decode[290] vdd gnd pinv_8
XDEC_INV_[291] Z[291] decode[291] vdd gnd pinv_8
XDEC_INV_[292] Z[292] decode[292] vdd gnd pinv_8
XDEC_INV_[293] Z[293] decode[293] vdd gnd pinv_8
XDEC_INV_[294] Z[294] decode[294] vdd gnd pinv_8
XDEC_INV_[295] Z[295] decode[295] vdd gnd pinv_8
XDEC_INV_[296] Z[296] decode[296] vdd gnd pinv_8
XDEC_INV_[297] Z[297] decode[297] vdd gnd pinv_8
XDEC_INV_[298] Z[298] decode[298] vdd gnd pinv_8
XDEC_INV_[299] Z[299] decode[299] vdd gnd pinv_8
XDEC_INV_[300] Z[300] decode[300] vdd gnd pinv_8
XDEC_INV_[301] Z[301] decode[301] vdd gnd pinv_8
XDEC_INV_[302] Z[302] decode[302] vdd gnd pinv_8
XDEC_INV_[303] Z[303] decode[303] vdd gnd pinv_8
XDEC_INV_[304] Z[304] decode[304] vdd gnd pinv_8
XDEC_INV_[305] Z[305] decode[305] vdd gnd pinv_8
XDEC_INV_[306] Z[306] decode[306] vdd gnd pinv_8
XDEC_INV_[307] Z[307] decode[307] vdd gnd pinv_8
XDEC_INV_[308] Z[308] decode[308] vdd gnd pinv_8
XDEC_INV_[309] Z[309] decode[309] vdd gnd pinv_8
XDEC_INV_[310] Z[310] decode[310] vdd gnd pinv_8
XDEC_INV_[311] Z[311] decode[311] vdd gnd pinv_8
XDEC_INV_[312] Z[312] decode[312] vdd gnd pinv_8
XDEC_INV_[313] Z[313] decode[313] vdd gnd pinv_8
XDEC_INV_[314] Z[314] decode[314] vdd gnd pinv_8
XDEC_INV_[315] Z[315] decode[315] vdd gnd pinv_8
XDEC_INV_[316] Z[316] decode[316] vdd gnd pinv_8
XDEC_INV_[317] Z[317] decode[317] vdd gnd pinv_8
XDEC_INV_[318] Z[318] decode[318] vdd gnd pinv_8
XDEC_INV_[319] Z[319] decode[319] vdd gnd pinv_8
XDEC_INV_[320] Z[320] decode[320] vdd gnd pinv_8
XDEC_INV_[321] Z[321] decode[321] vdd gnd pinv_8
XDEC_INV_[322] Z[322] decode[322] vdd gnd pinv_8
XDEC_INV_[323] Z[323] decode[323] vdd gnd pinv_8
XDEC_INV_[324] Z[324] decode[324] vdd gnd pinv_8
XDEC_INV_[325] Z[325] decode[325] vdd gnd pinv_8
XDEC_INV_[326] Z[326] decode[326] vdd gnd pinv_8
XDEC_INV_[327] Z[327] decode[327] vdd gnd pinv_8
XDEC_INV_[328] Z[328] decode[328] vdd gnd pinv_8
XDEC_INV_[329] Z[329] decode[329] vdd gnd pinv_8
XDEC_INV_[330] Z[330] decode[330] vdd gnd pinv_8
XDEC_INV_[331] Z[331] decode[331] vdd gnd pinv_8
XDEC_INV_[332] Z[332] decode[332] vdd gnd pinv_8
XDEC_INV_[333] Z[333] decode[333] vdd gnd pinv_8
XDEC_INV_[334] Z[334] decode[334] vdd gnd pinv_8
XDEC_INV_[335] Z[335] decode[335] vdd gnd pinv_8
XDEC_INV_[336] Z[336] decode[336] vdd gnd pinv_8
XDEC_INV_[337] Z[337] decode[337] vdd gnd pinv_8
XDEC_INV_[338] Z[338] decode[338] vdd gnd pinv_8
XDEC_INV_[339] Z[339] decode[339] vdd gnd pinv_8
XDEC_INV_[340] Z[340] decode[340] vdd gnd pinv_8
XDEC_INV_[341] Z[341] decode[341] vdd gnd pinv_8
XDEC_INV_[342] Z[342] decode[342] vdd gnd pinv_8
XDEC_INV_[343] Z[343] decode[343] vdd gnd pinv_8
XDEC_INV_[344] Z[344] decode[344] vdd gnd pinv_8
XDEC_INV_[345] Z[345] decode[345] vdd gnd pinv_8
XDEC_INV_[346] Z[346] decode[346] vdd gnd pinv_8
XDEC_INV_[347] Z[347] decode[347] vdd gnd pinv_8
XDEC_INV_[348] Z[348] decode[348] vdd gnd pinv_8
XDEC_INV_[349] Z[349] decode[349] vdd gnd pinv_8
XDEC_INV_[350] Z[350] decode[350] vdd gnd pinv_8
XDEC_INV_[351] Z[351] decode[351] vdd gnd pinv_8
XDEC_INV_[352] Z[352] decode[352] vdd gnd pinv_8
XDEC_INV_[353] Z[353] decode[353] vdd gnd pinv_8
XDEC_INV_[354] Z[354] decode[354] vdd gnd pinv_8
XDEC_INV_[355] Z[355] decode[355] vdd gnd pinv_8
XDEC_INV_[356] Z[356] decode[356] vdd gnd pinv_8
XDEC_INV_[357] Z[357] decode[357] vdd gnd pinv_8
XDEC_INV_[358] Z[358] decode[358] vdd gnd pinv_8
XDEC_INV_[359] Z[359] decode[359] vdd gnd pinv_8
XDEC_INV_[360] Z[360] decode[360] vdd gnd pinv_8
XDEC_INV_[361] Z[361] decode[361] vdd gnd pinv_8
XDEC_INV_[362] Z[362] decode[362] vdd gnd pinv_8
XDEC_INV_[363] Z[363] decode[363] vdd gnd pinv_8
XDEC_INV_[364] Z[364] decode[364] vdd gnd pinv_8
XDEC_INV_[365] Z[365] decode[365] vdd gnd pinv_8
XDEC_INV_[366] Z[366] decode[366] vdd gnd pinv_8
XDEC_INV_[367] Z[367] decode[367] vdd gnd pinv_8
XDEC_INV_[368] Z[368] decode[368] vdd gnd pinv_8
XDEC_INV_[369] Z[369] decode[369] vdd gnd pinv_8
XDEC_INV_[370] Z[370] decode[370] vdd gnd pinv_8
XDEC_INV_[371] Z[371] decode[371] vdd gnd pinv_8
XDEC_INV_[372] Z[372] decode[372] vdd gnd pinv_8
XDEC_INV_[373] Z[373] decode[373] vdd gnd pinv_8
XDEC_INV_[374] Z[374] decode[374] vdd gnd pinv_8
XDEC_INV_[375] Z[375] decode[375] vdd gnd pinv_8
XDEC_INV_[376] Z[376] decode[376] vdd gnd pinv_8
XDEC_INV_[377] Z[377] decode[377] vdd gnd pinv_8
XDEC_INV_[378] Z[378] decode[378] vdd gnd pinv_8
XDEC_INV_[379] Z[379] decode[379] vdd gnd pinv_8
XDEC_INV_[380] Z[380] decode[380] vdd gnd pinv_8
XDEC_INV_[381] Z[381] decode[381] vdd gnd pinv_8
XDEC_INV_[382] Z[382] decode[382] vdd gnd pinv_8
XDEC_INV_[383] Z[383] decode[383] vdd gnd pinv_8
XDEC_INV_[384] Z[384] decode[384] vdd gnd pinv_8
XDEC_INV_[385] Z[385] decode[385] vdd gnd pinv_8
XDEC_INV_[386] Z[386] decode[386] vdd gnd pinv_8
XDEC_INV_[387] Z[387] decode[387] vdd gnd pinv_8
XDEC_INV_[388] Z[388] decode[388] vdd gnd pinv_8
XDEC_INV_[389] Z[389] decode[389] vdd gnd pinv_8
XDEC_INV_[390] Z[390] decode[390] vdd gnd pinv_8
XDEC_INV_[391] Z[391] decode[391] vdd gnd pinv_8
XDEC_INV_[392] Z[392] decode[392] vdd gnd pinv_8
XDEC_INV_[393] Z[393] decode[393] vdd gnd pinv_8
XDEC_INV_[394] Z[394] decode[394] vdd gnd pinv_8
XDEC_INV_[395] Z[395] decode[395] vdd gnd pinv_8
XDEC_INV_[396] Z[396] decode[396] vdd gnd pinv_8
XDEC_INV_[397] Z[397] decode[397] vdd gnd pinv_8
XDEC_INV_[398] Z[398] decode[398] vdd gnd pinv_8
XDEC_INV_[399] Z[399] decode[399] vdd gnd pinv_8
XDEC_INV_[400] Z[400] decode[400] vdd gnd pinv_8
XDEC_INV_[401] Z[401] decode[401] vdd gnd pinv_8
XDEC_INV_[402] Z[402] decode[402] vdd gnd pinv_8
XDEC_INV_[403] Z[403] decode[403] vdd gnd pinv_8
XDEC_INV_[404] Z[404] decode[404] vdd gnd pinv_8
XDEC_INV_[405] Z[405] decode[405] vdd gnd pinv_8
XDEC_INV_[406] Z[406] decode[406] vdd gnd pinv_8
XDEC_INV_[407] Z[407] decode[407] vdd gnd pinv_8
XDEC_INV_[408] Z[408] decode[408] vdd gnd pinv_8
XDEC_INV_[409] Z[409] decode[409] vdd gnd pinv_8
XDEC_INV_[410] Z[410] decode[410] vdd gnd pinv_8
XDEC_INV_[411] Z[411] decode[411] vdd gnd pinv_8
XDEC_INV_[412] Z[412] decode[412] vdd gnd pinv_8
XDEC_INV_[413] Z[413] decode[413] vdd gnd pinv_8
XDEC_INV_[414] Z[414] decode[414] vdd gnd pinv_8
XDEC_INV_[415] Z[415] decode[415] vdd gnd pinv_8
XDEC_INV_[416] Z[416] decode[416] vdd gnd pinv_8
XDEC_INV_[417] Z[417] decode[417] vdd gnd pinv_8
XDEC_INV_[418] Z[418] decode[418] vdd gnd pinv_8
XDEC_INV_[419] Z[419] decode[419] vdd gnd pinv_8
XDEC_INV_[420] Z[420] decode[420] vdd gnd pinv_8
XDEC_INV_[421] Z[421] decode[421] vdd gnd pinv_8
XDEC_INV_[422] Z[422] decode[422] vdd gnd pinv_8
XDEC_INV_[423] Z[423] decode[423] vdd gnd pinv_8
XDEC_INV_[424] Z[424] decode[424] vdd gnd pinv_8
XDEC_INV_[425] Z[425] decode[425] vdd gnd pinv_8
XDEC_INV_[426] Z[426] decode[426] vdd gnd pinv_8
XDEC_INV_[427] Z[427] decode[427] vdd gnd pinv_8
XDEC_INV_[428] Z[428] decode[428] vdd gnd pinv_8
XDEC_INV_[429] Z[429] decode[429] vdd gnd pinv_8
XDEC_INV_[430] Z[430] decode[430] vdd gnd pinv_8
XDEC_INV_[431] Z[431] decode[431] vdd gnd pinv_8
XDEC_INV_[432] Z[432] decode[432] vdd gnd pinv_8
XDEC_INV_[433] Z[433] decode[433] vdd gnd pinv_8
XDEC_INV_[434] Z[434] decode[434] vdd gnd pinv_8
XDEC_INV_[435] Z[435] decode[435] vdd gnd pinv_8
XDEC_INV_[436] Z[436] decode[436] vdd gnd pinv_8
XDEC_INV_[437] Z[437] decode[437] vdd gnd pinv_8
XDEC_INV_[438] Z[438] decode[438] vdd gnd pinv_8
XDEC_INV_[439] Z[439] decode[439] vdd gnd pinv_8
XDEC_INV_[440] Z[440] decode[440] vdd gnd pinv_8
XDEC_INV_[441] Z[441] decode[441] vdd gnd pinv_8
XDEC_INV_[442] Z[442] decode[442] vdd gnd pinv_8
XDEC_INV_[443] Z[443] decode[443] vdd gnd pinv_8
XDEC_INV_[444] Z[444] decode[444] vdd gnd pinv_8
XDEC_INV_[445] Z[445] decode[445] vdd gnd pinv_8
XDEC_INV_[446] Z[446] decode[446] vdd gnd pinv_8
XDEC_INV_[447] Z[447] decode[447] vdd gnd pinv_8
XDEC_INV_[448] Z[448] decode[448] vdd gnd pinv_8
XDEC_INV_[449] Z[449] decode[449] vdd gnd pinv_8
XDEC_INV_[450] Z[450] decode[450] vdd gnd pinv_8
XDEC_INV_[451] Z[451] decode[451] vdd gnd pinv_8
XDEC_INV_[452] Z[452] decode[452] vdd gnd pinv_8
XDEC_INV_[453] Z[453] decode[453] vdd gnd pinv_8
XDEC_INV_[454] Z[454] decode[454] vdd gnd pinv_8
XDEC_INV_[455] Z[455] decode[455] vdd gnd pinv_8
XDEC_INV_[456] Z[456] decode[456] vdd gnd pinv_8
XDEC_INV_[457] Z[457] decode[457] vdd gnd pinv_8
XDEC_INV_[458] Z[458] decode[458] vdd gnd pinv_8
XDEC_INV_[459] Z[459] decode[459] vdd gnd pinv_8
XDEC_INV_[460] Z[460] decode[460] vdd gnd pinv_8
XDEC_INV_[461] Z[461] decode[461] vdd gnd pinv_8
XDEC_INV_[462] Z[462] decode[462] vdd gnd pinv_8
XDEC_INV_[463] Z[463] decode[463] vdd gnd pinv_8
XDEC_INV_[464] Z[464] decode[464] vdd gnd pinv_8
XDEC_INV_[465] Z[465] decode[465] vdd gnd pinv_8
XDEC_INV_[466] Z[466] decode[466] vdd gnd pinv_8
XDEC_INV_[467] Z[467] decode[467] vdd gnd pinv_8
XDEC_INV_[468] Z[468] decode[468] vdd gnd pinv_8
XDEC_INV_[469] Z[469] decode[469] vdd gnd pinv_8
XDEC_INV_[470] Z[470] decode[470] vdd gnd pinv_8
XDEC_INV_[471] Z[471] decode[471] vdd gnd pinv_8
XDEC_INV_[472] Z[472] decode[472] vdd gnd pinv_8
XDEC_INV_[473] Z[473] decode[473] vdd gnd pinv_8
XDEC_INV_[474] Z[474] decode[474] vdd gnd pinv_8
XDEC_INV_[475] Z[475] decode[475] vdd gnd pinv_8
XDEC_INV_[476] Z[476] decode[476] vdd gnd pinv_8
XDEC_INV_[477] Z[477] decode[477] vdd gnd pinv_8
XDEC_INV_[478] Z[478] decode[478] vdd gnd pinv_8
XDEC_INV_[479] Z[479] decode[479] vdd gnd pinv_8
XDEC_INV_[480] Z[480] decode[480] vdd gnd pinv_8
XDEC_INV_[481] Z[481] decode[481] vdd gnd pinv_8
XDEC_INV_[482] Z[482] decode[482] vdd gnd pinv_8
XDEC_INV_[483] Z[483] decode[483] vdd gnd pinv_8
XDEC_INV_[484] Z[484] decode[484] vdd gnd pinv_8
XDEC_INV_[485] Z[485] decode[485] vdd gnd pinv_8
XDEC_INV_[486] Z[486] decode[486] vdd gnd pinv_8
XDEC_INV_[487] Z[487] decode[487] vdd gnd pinv_8
XDEC_INV_[488] Z[488] decode[488] vdd gnd pinv_8
XDEC_INV_[489] Z[489] decode[489] vdd gnd pinv_8
XDEC_INV_[490] Z[490] decode[490] vdd gnd pinv_8
XDEC_INV_[491] Z[491] decode[491] vdd gnd pinv_8
XDEC_INV_[492] Z[492] decode[492] vdd gnd pinv_8
XDEC_INV_[493] Z[493] decode[493] vdd gnd pinv_8
XDEC_INV_[494] Z[494] decode[494] vdd gnd pinv_8
XDEC_INV_[495] Z[495] decode[495] vdd gnd pinv_8
XDEC_INV_[496] Z[496] decode[496] vdd gnd pinv_8
XDEC_INV_[497] Z[497] decode[497] vdd gnd pinv_8
XDEC_INV_[498] Z[498] decode[498] vdd gnd pinv_8
XDEC_INV_[499] Z[499] decode[499] vdd gnd pinv_8
XDEC_INV_[500] Z[500] decode[500] vdd gnd pinv_8
XDEC_INV_[501] Z[501] decode[501] vdd gnd pinv_8
XDEC_INV_[502] Z[502] decode[502] vdd gnd pinv_8
XDEC_INV_[503] Z[503] decode[503] vdd gnd pinv_8
XDEC_INV_[504] Z[504] decode[504] vdd gnd pinv_8
XDEC_INV_[505] Z[505] decode[505] vdd gnd pinv_8
XDEC_INV_[506] Z[506] decode[506] vdd gnd pinv_8
XDEC_INV_[507] Z[507] decode[507] vdd gnd pinv_8
XDEC_INV_[508] Z[508] decode[508] vdd gnd pinv_8
XDEC_INV_[509] Z[509] decode[509] vdd gnd pinv_8
XDEC_INV_[510] Z[510] decode[510] vdd gnd pinv_8
XDEC_INV_[511] Z[511] decode[511] vdd gnd pinv_8
.ENDS hierarchical_decoder_512rows

.SUBCKT msf_address din[0] din[1] din[2] din[3] din[4] din[5] din[6] din[7] din[8] din[9] din[10] dout[0] dout_bar[0] dout[1] dout_bar[1] dout[2] dout_bar[2] dout[3] dout_bar[3] dout[4] dout_bar[4] dout[5] dout_bar[5] dout[6] dout_bar[6] dout[7] dout_bar[7] dout[8] dout_bar[8] dout[9] dout_bar[9] dout[10] dout_bar[10] clk vdd gnd
XXdff0 din[0] dout[0] dout_bar[0] clk vdd gnd ms_flop
XXdff1 din[1] dout[1] dout_bar[1] clk vdd gnd ms_flop
XXdff2 din[2] dout[2] dout_bar[2] clk vdd gnd ms_flop
XXdff3 din[3] dout[3] dout_bar[3] clk vdd gnd ms_flop
XXdff4 din[4] dout[4] dout_bar[4] clk vdd gnd ms_flop
XXdff5 din[5] dout[5] dout_bar[5] clk vdd gnd ms_flop
XXdff6 din[6] dout[6] dout_bar[6] clk vdd gnd ms_flop
XXdff7 din[7] dout[7] dout_bar[7] clk vdd gnd ms_flop
XXdff8 din[8] dout[8] dout_bar[8] clk vdd gnd ms_flop
XXdff9 din[9] dout[9] dout_bar[9] clk vdd gnd ms_flop
XXdff10 din[10] dout[10] dout_bar[10] clk vdd gnd ms_flop
.ENDS msf_address

.SUBCKT msf_data_in din[0] din[1] din[2] din[3] din[4] din[5] din[6] din[7] din[8] din[9] din[10] din[11] din[12] din[13] din[14] din[15] din[16] din[17] din[18] din[19] din[20] din[21] din[22] din[23] din[24] din[25] din[26] din[27] din[28] din[29] din[30] din[31] dout[0] dout_bar[0] dout[1] dout_bar[1] dout[2] dout_bar[2] dout[3] dout_bar[3] dout[4] dout_bar[4] dout[5] dout_bar[5] dout[6] dout_bar[6] dout[7] dout_bar[7] dout[8] dout_bar[8] dout[9] dout_bar[9] dout[10] dout_bar[10] dout[11] dout_bar[11] dout[12] dout_bar[12] dout[13] dout_bar[13] dout[14] dout_bar[14] dout[15] dout_bar[15] dout[16] dout_bar[16] dout[17] dout_bar[17] dout[18] dout_bar[18] dout[19] dout_bar[19] dout[20] dout_bar[20] dout[21] dout_bar[21] dout[22] dout_bar[22] dout[23] dout_bar[23] dout[24] dout_bar[24] dout[25] dout_bar[25] dout[26] dout_bar[26] dout[27] dout_bar[27] dout[28] dout_bar[28] dout[29] dout_bar[29] dout[30] dout_bar[30] dout[31] dout_bar[31] clk vdd gnd
XXdff0 din[0] dout[0] dout_bar[0] clk vdd gnd ms_flop
XXdff4 din[1] dout[1] dout_bar[1] clk vdd gnd ms_flop
XXdff8 din[2] dout[2] dout_bar[2] clk vdd gnd ms_flop
XXdff12 din[3] dout[3] dout_bar[3] clk vdd gnd ms_flop
XXdff16 din[4] dout[4] dout_bar[4] clk vdd gnd ms_flop
XXdff20 din[5] dout[5] dout_bar[5] clk vdd gnd ms_flop
XXdff24 din[6] dout[6] dout_bar[6] clk vdd gnd ms_flop
XXdff28 din[7] dout[7] dout_bar[7] clk vdd gnd ms_flop
XXdff32 din[8] dout[8] dout_bar[8] clk vdd gnd ms_flop
XXdff36 din[9] dout[9] dout_bar[9] clk vdd gnd ms_flop
XXdff40 din[10] dout[10] dout_bar[10] clk vdd gnd ms_flop
XXdff44 din[11] dout[11] dout_bar[11] clk vdd gnd ms_flop
XXdff48 din[12] dout[12] dout_bar[12] clk vdd gnd ms_flop
XXdff52 din[13] dout[13] dout_bar[13] clk vdd gnd ms_flop
XXdff56 din[14] dout[14] dout_bar[14] clk vdd gnd ms_flop
XXdff60 din[15] dout[15] dout_bar[15] clk vdd gnd ms_flop
XXdff64 din[16] dout[16] dout_bar[16] clk vdd gnd ms_flop
XXdff68 din[17] dout[17] dout_bar[17] clk vdd gnd ms_flop
XXdff72 din[18] dout[18] dout_bar[18] clk vdd gnd ms_flop
XXdff76 din[19] dout[19] dout_bar[19] clk vdd gnd ms_flop
XXdff80 din[20] dout[20] dout_bar[20] clk vdd gnd ms_flop
XXdff84 din[21] dout[21] dout_bar[21] clk vdd gnd ms_flop
XXdff88 din[22] dout[22] dout_bar[22] clk vdd gnd ms_flop
XXdff92 din[23] dout[23] dout_bar[23] clk vdd gnd ms_flop
XXdff96 din[24] dout[24] dout_bar[24] clk vdd gnd ms_flop
XXdff100 din[25] dout[25] dout_bar[25] clk vdd gnd ms_flop
XXdff104 din[26] dout[26] dout_bar[26] clk vdd gnd ms_flop
XXdff108 din[27] dout[27] dout_bar[27] clk vdd gnd ms_flop
XXdff112 din[28] dout[28] dout_bar[28] clk vdd gnd ms_flop
XXdff116 din[29] dout[29] dout_bar[29] clk vdd gnd ms_flop
XXdff120 din[30] dout[30] dout_bar[30] clk vdd gnd ms_flop
XXdff124 din[31] dout[31] dout_bar[31] clk vdd gnd ms_flop
.ENDS msf_data_in

.SUBCKT tri_gate in out en en_bar vdd gnd
M_1 net_2 in_inv gnd gnd NMOS_VTG W=180.000000n L=50.000000n
M_2 out en net_2 gnd NMOS_VTG W=180.000000n L=50.000000n
M_3 net_3 in_inv vdd vdd PMOS_VTG W=360.000000n L=50.000000n
M_4 out en_bar net_3 vdd PMOS_VTG W=360.000000n L=50.000000n
M_5 in_inv in vdd vdd PMOS_VTG W=180.000000n L=50.000000n
M_6 in_inv in gnd gnd NMOS_VTG W=90.000000n L=50.000000n
.ENDS


.SUBCKT tri_gate_array in[0] in[1] in[2] in[3] in[4] in[5] in[6] in[7] in[8] in[9] in[10] in[11] in[12] in[13] in[14] in[15] in[16] in[17] in[18] in[19] in[20] in[21] in[22] in[23] in[24] in[25] in[26] in[27] in[28] in[29] in[30] in[31] out[0] out[1] out[2] out[3] out[4] out[5] out[6] out[7] out[8] out[9] out[10] out[11] out[12] out[13] out[14] out[15] out[16] out[17] out[18] out[19] out[20] out[21] out[22] out[23] out[24] out[25] out[26] out[27] out[28] out[29] out[30] out[31] en en_bar vdd gnd
XXtri_gate0 in[0] out[0] en en_bar vdd gnd tri_gate
XXtri_gate4 in[1] out[1] en en_bar vdd gnd tri_gate
XXtri_gate8 in[2] out[2] en en_bar vdd gnd tri_gate
XXtri_gate12 in[3] out[3] en en_bar vdd gnd tri_gate
XXtri_gate16 in[4] out[4] en en_bar vdd gnd tri_gate
XXtri_gate20 in[5] out[5] en en_bar vdd gnd tri_gate
XXtri_gate24 in[6] out[6] en en_bar vdd gnd tri_gate
XXtri_gate28 in[7] out[7] en en_bar vdd gnd tri_gate
XXtri_gate32 in[8] out[8] en en_bar vdd gnd tri_gate
XXtri_gate36 in[9] out[9] en en_bar vdd gnd tri_gate
XXtri_gate40 in[10] out[10] en en_bar vdd gnd tri_gate
XXtri_gate44 in[11] out[11] en en_bar vdd gnd tri_gate
XXtri_gate48 in[12] out[12] en en_bar vdd gnd tri_gate
XXtri_gate52 in[13] out[13] en en_bar vdd gnd tri_gate
XXtri_gate56 in[14] out[14] en en_bar vdd gnd tri_gate
XXtri_gate60 in[15] out[15] en en_bar vdd gnd tri_gate
XXtri_gate64 in[16] out[16] en en_bar vdd gnd tri_gate
XXtri_gate68 in[17] out[17] en en_bar vdd gnd tri_gate
XXtri_gate72 in[18] out[18] en en_bar vdd gnd tri_gate
XXtri_gate76 in[19] out[19] en en_bar vdd gnd tri_gate
XXtri_gate80 in[20] out[20] en en_bar vdd gnd tri_gate
XXtri_gate84 in[21] out[21] en en_bar vdd gnd tri_gate
XXtri_gate88 in[22] out[22] en en_bar vdd gnd tri_gate
XXtri_gate92 in[23] out[23] en en_bar vdd gnd tri_gate
XXtri_gate96 in[24] out[24] en en_bar vdd gnd tri_gate
XXtri_gate100 in[25] out[25] en en_bar vdd gnd tri_gate
XXtri_gate104 in[26] out[26] en en_bar vdd gnd tri_gate
XXtri_gate108 in[27] out[27] en en_bar vdd gnd tri_gate
XXtri_gate112 in[28] out[28] en en_bar vdd gnd tri_gate
XXtri_gate116 in[29] out[29] en en_bar vdd gnd tri_gate
XXtri_gate120 in[30] out[30] en en_bar vdd gnd tri_gate
XXtri_gate124 in[31] out[31] en en_bar vdd gnd tri_gate
.ENDS tri_gate_array

.SUBCKT pinv_11 A Z vdd gnd
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01125p ad=0.01125p
.ENDS pinv_11

.SUBCKT pinv_12 A Z vdd gnd
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01125p ad=0.01125p
.ENDS pinv_12

.SUBCKT pnand2_4 A B Z vdd gnd
Mpnand2_pmos1 vdd A Z vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpnand2_pmos2 Z B vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpnand2_nmos1 Z B net1 gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.0225p ad=0.0225p
Mpnand2_nmos2 net1 A gnd gnd nmos_vtg m=1 w=0.18u l=0.05u pd=0.46u ps=0.46u as=0.0225p ad=0.0225p
.ENDS pnand2_4

.SUBCKT wordline_driver in[0] in[1] in[2] in[3] in[4] in[5] in[6] in[7] in[8] in[9] in[10] in[11] in[12] in[13] in[14] in[15] in[16] in[17] in[18] in[19] in[20] in[21] in[22] in[23] in[24] in[25] in[26] in[27] in[28] in[29] in[30] in[31] in[32] in[33] in[34] in[35] in[36] in[37] in[38] in[39] in[40] in[41] in[42] in[43] in[44] in[45] in[46] in[47] in[48] in[49] in[50] in[51] in[52] in[53] in[54] in[55] in[56] in[57] in[58] in[59] in[60] in[61] in[62] in[63] in[64] in[65] in[66] in[67] in[68] in[69] in[70] in[71] in[72] in[73] in[74] in[75] in[76] in[77] in[78] in[79] in[80] in[81] in[82] in[83] in[84] in[85] in[86] in[87] in[88] in[89] in[90] in[91] in[92] in[93] in[94] in[95] in[96] in[97] in[98] in[99] in[100] in[101] in[102] in[103] in[104] in[105] in[106] in[107] in[108] in[109] in[110] in[111] in[112] in[113] in[114] in[115] in[116] in[117] in[118] in[119] in[120] in[121] in[122] in[123] in[124] in[125] in[126] in[127] in[128] in[129] in[130] in[131] in[132] in[133] in[134] in[135] in[136] in[137] in[138] in[139] in[140] in[141] in[142] in[143] in[144] in[145] in[146] in[147] in[148] in[149] in[150] in[151] in[152] in[153] in[154] in[155] in[156] in[157] in[158] in[159] in[160] in[161] in[162] in[163] in[164] in[165] in[166] in[167] in[168] in[169] in[170] in[171] in[172] in[173] in[174] in[175] in[176] in[177] in[178] in[179] in[180] in[181] in[182] in[183] in[184] in[185] in[186] in[187] in[188] in[189] in[190] in[191] in[192] in[193] in[194] in[195] in[196] in[197] in[198] in[199] in[200] in[201] in[202] in[203] in[204] in[205] in[206] in[207] in[208] in[209] in[210] in[211] in[212] in[213] in[214] in[215] in[216] in[217] in[218] in[219] in[220] in[221] in[222] in[223] in[224] in[225] in[226] in[227] in[228] in[229] in[230] in[231] in[232] in[233] in[234] in[235] in[236] in[237] in[238] in[239] in[240] in[241] in[242] in[243] in[244] in[245] in[246] in[247] in[248] in[249] in[250] in[251] in[252] in[253] in[254] in[255] in[256] in[257] in[258] in[259] in[260] in[261] in[262] in[263] in[264] in[265] in[266] in[267] in[268] in[269] in[270] in[271] in[272] in[273] in[274] in[275] in[276] in[277] in[278] in[279] in[280] in[281] in[282] in[283] in[284] in[285] in[286] in[287] in[288] in[289] in[290] in[291] in[292] in[293] in[294] in[295] in[296] in[297] in[298] in[299] in[300] in[301] in[302] in[303] in[304] in[305] in[306] in[307] in[308] in[309] in[310] in[311] in[312] in[313] in[314] in[315] in[316] in[317] in[318] in[319] in[320] in[321] in[322] in[323] in[324] in[325] in[326] in[327] in[328] in[329] in[330] in[331] in[332] in[333] in[334] in[335] in[336] in[337] in[338] in[339] in[340] in[341] in[342] in[343] in[344] in[345] in[346] in[347] in[348] in[349] in[350] in[351] in[352] in[353] in[354] in[355] in[356] in[357] in[358] in[359] in[360] in[361] in[362] in[363] in[364] in[365] in[366] in[367] in[368] in[369] in[370] in[371] in[372] in[373] in[374] in[375] in[376] in[377] in[378] in[379] in[380] in[381] in[382] in[383] in[384] in[385] in[386] in[387] in[388] in[389] in[390] in[391] in[392] in[393] in[394] in[395] in[396] in[397] in[398] in[399] in[400] in[401] in[402] in[403] in[404] in[405] in[406] in[407] in[408] in[409] in[410] in[411] in[412] in[413] in[414] in[415] in[416] in[417] in[418] in[419] in[420] in[421] in[422] in[423] in[424] in[425] in[426] in[427] in[428] in[429] in[430] in[431] in[432] in[433] in[434] in[435] in[436] in[437] in[438] in[439] in[440] in[441] in[442] in[443] in[444] in[445] in[446] in[447] in[448] in[449] in[450] in[451] in[452] in[453] in[454] in[455] in[456] in[457] in[458] in[459] in[460] in[461] in[462] in[463] in[464] in[465] in[466] in[467] in[468] in[469] in[470] in[471] in[472] in[473] in[474] in[475] in[476] in[477] in[478] in[479] in[480] in[481] in[482] in[483] in[484] in[485] in[486] in[487] in[488] in[489] in[490] in[491] in[492] in[493] in[494] in[495] in[496] in[497] in[498] in[499] in[500] in[501] in[502] in[503] in[504] in[505] in[506] in[507] in[508] in[509] in[510] in[511] wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] wl[128] wl[129] wl[130] wl[131] wl[132] wl[133] wl[134] wl[135] wl[136] wl[137] wl[138] wl[139] wl[140] wl[141] wl[142] wl[143] wl[144] wl[145] wl[146] wl[147] wl[148] wl[149] wl[150] wl[151] wl[152] wl[153] wl[154] wl[155] wl[156] wl[157] wl[158] wl[159] wl[160] wl[161] wl[162] wl[163] wl[164] wl[165] wl[166] wl[167] wl[168] wl[169] wl[170] wl[171] wl[172] wl[173] wl[174] wl[175] wl[176] wl[177] wl[178] wl[179] wl[180] wl[181] wl[182] wl[183] wl[184] wl[185] wl[186] wl[187] wl[188] wl[189] wl[190] wl[191] wl[192] wl[193] wl[194] wl[195] wl[196] wl[197] wl[198] wl[199] wl[200] wl[201] wl[202] wl[203] wl[204] wl[205] wl[206] wl[207] wl[208] wl[209] wl[210] wl[211] wl[212] wl[213] wl[214] wl[215] wl[216] wl[217] wl[218] wl[219] wl[220] wl[221] wl[222] wl[223] wl[224] wl[225] wl[226] wl[227] wl[228] wl[229] wl[230] wl[231] wl[232] wl[233] wl[234] wl[235] wl[236] wl[237] wl[238] wl[239] wl[240] wl[241] wl[242] wl[243] wl[244] wl[245] wl[246] wl[247] wl[248] wl[249] wl[250] wl[251] wl[252] wl[253] wl[254] wl[255] wl[256] wl[257] wl[258] wl[259] wl[260] wl[261] wl[262] wl[263] wl[264] wl[265] wl[266] wl[267] wl[268] wl[269] wl[270] wl[271] wl[272] wl[273] wl[274] wl[275] wl[276] wl[277] wl[278] wl[279] wl[280] wl[281] wl[282] wl[283] wl[284] wl[285] wl[286] wl[287] wl[288] wl[289] wl[290] wl[291] wl[292] wl[293] wl[294] wl[295] wl[296] wl[297] wl[298] wl[299] wl[300] wl[301] wl[302] wl[303] wl[304] wl[305] wl[306] wl[307] wl[308] wl[309] wl[310] wl[311] wl[312] wl[313] wl[314] wl[315] wl[316] wl[317] wl[318] wl[319] wl[320] wl[321] wl[322] wl[323] wl[324] wl[325] wl[326] wl[327] wl[328] wl[329] wl[330] wl[331] wl[332] wl[333] wl[334] wl[335] wl[336] wl[337] wl[338] wl[339] wl[340] wl[341] wl[342] wl[343] wl[344] wl[345] wl[346] wl[347] wl[348] wl[349] wl[350] wl[351] wl[352] wl[353] wl[354] wl[355] wl[356] wl[357] wl[358] wl[359] wl[360] wl[361] wl[362] wl[363] wl[364] wl[365] wl[366] wl[367] wl[368] wl[369] wl[370] wl[371] wl[372] wl[373] wl[374] wl[375] wl[376] wl[377] wl[378] wl[379] wl[380] wl[381] wl[382] wl[383] wl[384] wl[385] wl[386] wl[387] wl[388] wl[389] wl[390] wl[391] wl[392] wl[393] wl[394] wl[395] wl[396] wl[397] wl[398] wl[399] wl[400] wl[401] wl[402] wl[403] wl[404] wl[405] wl[406] wl[407] wl[408] wl[409] wl[410] wl[411] wl[412] wl[413] wl[414] wl[415] wl[416] wl[417] wl[418] wl[419] wl[420] wl[421] wl[422] wl[423] wl[424] wl[425] wl[426] wl[427] wl[428] wl[429] wl[430] wl[431] wl[432] wl[433] wl[434] wl[435] wl[436] wl[437] wl[438] wl[439] wl[440] wl[441] wl[442] wl[443] wl[444] wl[445] wl[446] wl[447] wl[448] wl[449] wl[450] wl[451] wl[452] wl[453] wl[454] wl[455] wl[456] wl[457] wl[458] wl[459] wl[460] wl[461] wl[462] wl[463] wl[464] wl[465] wl[466] wl[467] wl[468] wl[469] wl[470] wl[471] wl[472] wl[473] wl[474] wl[475] wl[476] wl[477] wl[478] wl[479] wl[480] wl[481] wl[482] wl[483] wl[484] wl[485] wl[486] wl[487] wl[488] wl[489] wl[490] wl[491] wl[492] wl[493] wl[494] wl[495] wl[496] wl[497] wl[498] wl[499] wl[500] wl[501] wl[502] wl[503] wl[504] wl[505] wl[506] wl[507] wl[508] wl[509] wl[510] wl[511] en vdd gnd
Xwl_driver_inv_en0 en en_bar[0] vdd gnd pinv_12
Xwl_driver_nand0 en_bar[0] in[0] net[0] vdd gnd pnand2_4
Xwl_driver_inv0 net[0] wl[0] vdd gnd pinv_11
Xwl_driver_inv_en1 en en_bar[1] vdd gnd pinv_12
Xwl_driver_nand1 en_bar[1] in[1] net[1] vdd gnd pnand2_4
Xwl_driver_inv1 net[1] wl[1] vdd gnd pinv_11
Xwl_driver_inv_en2 en en_bar[2] vdd gnd pinv_12
Xwl_driver_nand2 en_bar[2] in[2] net[2] vdd gnd pnand2_4
Xwl_driver_inv2 net[2] wl[2] vdd gnd pinv_11
Xwl_driver_inv_en3 en en_bar[3] vdd gnd pinv_12
Xwl_driver_nand3 en_bar[3] in[3] net[3] vdd gnd pnand2_4
Xwl_driver_inv3 net[3] wl[3] vdd gnd pinv_11
Xwl_driver_inv_en4 en en_bar[4] vdd gnd pinv_12
Xwl_driver_nand4 en_bar[4] in[4] net[4] vdd gnd pnand2_4
Xwl_driver_inv4 net[4] wl[4] vdd gnd pinv_11
Xwl_driver_inv_en5 en en_bar[5] vdd gnd pinv_12
Xwl_driver_nand5 en_bar[5] in[5] net[5] vdd gnd pnand2_4
Xwl_driver_inv5 net[5] wl[5] vdd gnd pinv_11
Xwl_driver_inv_en6 en en_bar[6] vdd gnd pinv_12
Xwl_driver_nand6 en_bar[6] in[6] net[6] vdd gnd pnand2_4
Xwl_driver_inv6 net[6] wl[6] vdd gnd pinv_11
Xwl_driver_inv_en7 en en_bar[7] vdd gnd pinv_12
Xwl_driver_nand7 en_bar[7] in[7] net[7] vdd gnd pnand2_4
Xwl_driver_inv7 net[7] wl[7] vdd gnd pinv_11
Xwl_driver_inv_en8 en en_bar[8] vdd gnd pinv_12
Xwl_driver_nand8 en_bar[8] in[8] net[8] vdd gnd pnand2_4
Xwl_driver_inv8 net[8] wl[8] vdd gnd pinv_11
Xwl_driver_inv_en9 en en_bar[9] vdd gnd pinv_12
Xwl_driver_nand9 en_bar[9] in[9] net[9] vdd gnd pnand2_4
Xwl_driver_inv9 net[9] wl[9] vdd gnd pinv_11
Xwl_driver_inv_en10 en en_bar[10] vdd gnd pinv_12
Xwl_driver_nand10 en_bar[10] in[10] net[10] vdd gnd pnand2_4
Xwl_driver_inv10 net[10] wl[10] vdd gnd pinv_11
Xwl_driver_inv_en11 en en_bar[11] vdd gnd pinv_12
Xwl_driver_nand11 en_bar[11] in[11] net[11] vdd gnd pnand2_4
Xwl_driver_inv11 net[11] wl[11] vdd gnd pinv_11
Xwl_driver_inv_en12 en en_bar[12] vdd gnd pinv_12
Xwl_driver_nand12 en_bar[12] in[12] net[12] vdd gnd pnand2_4
Xwl_driver_inv12 net[12] wl[12] vdd gnd pinv_11
Xwl_driver_inv_en13 en en_bar[13] vdd gnd pinv_12
Xwl_driver_nand13 en_bar[13] in[13] net[13] vdd gnd pnand2_4
Xwl_driver_inv13 net[13] wl[13] vdd gnd pinv_11
Xwl_driver_inv_en14 en en_bar[14] vdd gnd pinv_12
Xwl_driver_nand14 en_bar[14] in[14] net[14] vdd gnd pnand2_4
Xwl_driver_inv14 net[14] wl[14] vdd gnd pinv_11
Xwl_driver_inv_en15 en en_bar[15] vdd gnd pinv_12
Xwl_driver_nand15 en_bar[15] in[15] net[15] vdd gnd pnand2_4
Xwl_driver_inv15 net[15] wl[15] vdd gnd pinv_11
Xwl_driver_inv_en16 en en_bar[16] vdd gnd pinv_12
Xwl_driver_nand16 en_bar[16] in[16] net[16] vdd gnd pnand2_4
Xwl_driver_inv16 net[16] wl[16] vdd gnd pinv_11
Xwl_driver_inv_en17 en en_bar[17] vdd gnd pinv_12
Xwl_driver_nand17 en_bar[17] in[17] net[17] vdd gnd pnand2_4
Xwl_driver_inv17 net[17] wl[17] vdd gnd pinv_11
Xwl_driver_inv_en18 en en_bar[18] vdd gnd pinv_12
Xwl_driver_nand18 en_bar[18] in[18] net[18] vdd gnd pnand2_4
Xwl_driver_inv18 net[18] wl[18] vdd gnd pinv_11
Xwl_driver_inv_en19 en en_bar[19] vdd gnd pinv_12
Xwl_driver_nand19 en_bar[19] in[19] net[19] vdd gnd pnand2_4
Xwl_driver_inv19 net[19] wl[19] vdd gnd pinv_11
Xwl_driver_inv_en20 en en_bar[20] vdd gnd pinv_12
Xwl_driver_nand20 en_bar[20] in[20] net[20] vdd gnd pnand2_4
Xwl_driver_inv20 net[20] wl[20] vdd gnd pinv_11
Xwl_driver_inv_en21 en en_bar[21] vdd gnd pinv_12
Xwl_driver_nand21 en_bar[21] in[21] net[21] vdd gnd pnand2_4
Xwl_driver_inv21 net[21] wl[21] vdd gnd pinv_11
Xwl_driver_inv_en22 en en_bar[22] vdd gnd pinv_12
Xwl_driver_nand22 en_bar[22] in[22] net[22] vdd gnd pnand2_4
Xwl_driver_inv22 net[22] wl[22] vdd gnd pinv_11
Xwl_driver_inv_en23 en en_bar[23] vdd gnd pinv_12
Xwl_driver_nand23 en_bar[23] in[23] net[23] vdd gnd pnand2_4
Xwl_driver_inv23 net[23] wl[23] vdd gnd pinv_11
Xwl_driver_inv_en24 en en_bar[24] vdd gnd pinv_12
Xwl_driver_nand24 en_bar[24] in[24] net[24] vdd gnd pnand2_4
Xwl_driver_inv24 net[24] wl[24] vdd gnd pinv_11
Xwl_driver_inv_en25 en en_bar[25] vdd gnd pinv_12
Xwl_driver_nand25 en_bar[25] in[25] net[25] vdd gnd pnand2_4
Xwl_driver_inv25 net[25] wl[25] vdd gnd pinv_11
Xwl_driver_inv_en26 en en_bar[26] vdd gnd pinv_12
Xwl_driver_nand26 en_bar[26] in[26] net[26] vdd gnd pnand2_4
Xwl_driver_inv26 net[26] wl[26] vdd gnd pinv_11
Xwl_driver_inv_en27 en en_bar[27] vdd gnd pinv_12
Xwl_driver_nand27 en_bar[27] in[27] net[27] vdd gnd pnand2_4
Xwl_driver_inv27 net[27] wl[27] vdd gnd pinv_11
Xwl_driver_inv_en28 en en_bar[28] vdd gnd pinv_12
Xwl_driver_nand28 en_bar[28] in[28] net[28] vdd gnd pnand2_4
Xwl_driver_inv28 net[28] wl[28] vdd gnd pinv_11
Xwl_driver_inv_en29 en en_bar[29] vdd gnd pinv_12
Xwl_driver_nand29 en_bar[29] in[29] net[29] vdd gnd pnand2_4
Xwl_driver_inv29 net[29] wl[29] vdd gnd pinv_11
Xwl_driver_inv_en30 en en_bar[30] vdd gnd pinv_12
Xwl_driver_nand30 en_bar[30] in[30] net[30] vdd gnd pnand2_4
Xwl_driver_inv30 net[30] wl[30] vdd gnd pinv_11
Xwl_driver_inv_en31 en en_bar[31] vdd gnd pinv_12
Xwl_driver_nand31 en_bar[31] in[31] net[31] vdd gnd pnand2_4
Xwl_driver_inv31 net[31] wl[31] vdd gnd pinv_11
Xwl_driver_inv_en32 en en_bar[32] vdd gnd pinv_12
Xwl_driver_nand32 en_bar[32] in[32] net[32] vdd gnd pnand2_4
Xwl_driver_inv32 net[32] wl[32] vdd gnd pinv_11
Xwl_driver_inv_en33 en en_bar[33] vdd gnd pinv_12
Xwl_driver_nand33 en_bar[33] in[33] net[33] vdd gnd pnand2_4
Xwl_driver_inv33 net[33] wl[33] vdd gnd pinv_11
Xwl_driver_inv_en34 en en_bar[34] vdd gnd pinv_12
Xwl_driver_nand34 en_bar[34] in[34] net[34] vdd gnd pnand2_4
Xwl_driver_inv34 net[34] wl[34] vdd gnd pinv_11
Xwl_driver_inv_en35 en en_bar[35] vdd gnd pinv_12
Xwl_driver_nand35 en_bar[35] in[35] net[35] vdd gnd pnand2_4
Xwl_driver_inv35 net[35] wl[35] vdd gnd pinv_11
Xwl_driver_inv_en36 en en_bar[36] vdd gnd pinv_12
Xwl_driver_nand36 en_bar[36] in[36] net[36] vdd gnd pnand2_4
Xwl_driver_inv36 net[36] wl[36] vdd gnd pinv_11
Xwl_driver_inv_en37 en en_bar[37] vdd gnd pinv_12
Xwl_driver_nand37 en_bar[37] in[37] net[37] vdd gnd pnand2_4
Xwl_driver_inv37 net[37] wl[37] vdd gnd pinv_11
Xwl_driver_inv_en38 en en_bar[38] vdd gnd pinv_12
Xwl_driver_nand38 en_bar[38] in[38] net[38] vdd gnd pnand2_4
Xwl_driver_inv38 net[38] wl[38] vdd gnd pinv_11
Xwl_driver_inv_en39 en en_bar[39] vdd gnd pinv_12
Xwl_driver_nand39 en_bar[39] in[39] net[39] vdd gnd pnand2_4
Xwl_driver_inv39 net[39] wl[39] vdd gnd pinv_11
Xwl_driver_inv_en40 en en_bar[40] vdd gnd pinv_12
Xwl_driver_nand40 en_bar[40] in[40] net[40] vdd gnd pnand2_4
Xwl_driver_inv40 net[40] wl[40] vdd gnd pinv_11
Xwl_driver_inv_en41 en en_bar[41] vdd gnd pinv_12
Xwl_driver_nand41 en_bar[41] in[41] net[41] vdd gnd pnand2_4
Xwl_driver_inv41 net[41] wl[41] vdd gnd pinv_11
Xwl_driver_inv_en42 en en_bar[42] vdd gnd pinv_12
Xwl_driver_nand42 en_bar[42] in[42] net[42] vdd gnd pnand2_4
Xwl_driver_inv42 net[42] wl[42] vdd gnd pinv_11
Xwl_driver_inv_en43 en en_bar[43] vdd gnd pinv_12
Xwl_driver_nand43 en_bar[43] in[43] net[43] vdd gnd pnand2_4
Xwl_driver_inv43 net[43] wl[43] vdd gnd pinv_11
Xwl_driver_inv_en44 en en_bar[44] vdd gnd pinv_12
Xwl_driver_nand44 en_bar[44] in[44] net[44] vdd gnd pnand2_4
Xwl_driver_inv44 net[44] wl[44] vdd gnd pinv_11
Xwl_driver_inv_en45 en en_bar[45] vdd gnd pinv_12
Xwl_driver_nand45 en_bar[45] in[45] net[45] vdd gnd pnand2_4
Xwl_driver_inv45 net[45] wl[45] vdd gnd pinv_11
Xwl_driver_inv_en46 en en_bar[46] vdd gnd pinv_12
Xwl_driver_nand46 en_bar[46] in[46] net[46] vdd gnd pnand2_4
Xwl_driver_inv46 net[46] wl[46] vdd gnd pinv_11
Xwl_driver_inv_en47 en en_bar[47] vdd gnd pinv_12
Xwl_driver_nand47 en_bar[47] in[47] net[47] vdd gnd pnand2_4
Xwl_driver_inv47 net[47] wl[47] vdd gnd pinv_11
Xwl_driver_inv_en48 en en_bar[48] vdd gnd pinv_12
Xwl_driver_nand48 en_bar[48] in[48] net[48] vdd gnd pnand2_4
Xwl_driver_inv48 net[48] wl[48] vdd gnd pinv_11
Xwl_driver_inv_en49 en en_bar[49] vdd gnd pinv_12
Xwl_driver_nand49 en_bar[49] in[49] net[49] vdd gnd pnand2_4
Xwl_driver_inv49 net[49] wl[49] vdd gnd pinv_11
Xwl_driver_inv_en50 en en_bar[50] vdd gnd pinv_12
Xwl_driver_nand50 en_bar[50] in[50] net[50] vdd gnd pnand2_4
Xwl_driver_inv50 net[50] wl[50] vdd gnd pinv_11
Xwl_driver_inv_en51 en en_bar[51] vdd gnd pinv_12
Xwl_driver_nand51 en_bar[51] in[51] net[51] vdd gnd pnand2_4
Xwl_driver_inv51 net[51] wl[51] vdd gnd pinv_11
Xwl_driver_inv_en52 en en_bar[52] vdd gnd pinv_12
Xwl_driver_nand52 en_bar[52] in[52] net[52] vdd gnd pnand2_4
Xwl_driver_inv52 net[52] wl[52] vdd gnd pinv_11
Xwl_driver_inv_en53 en en_bar[53] vdd gnd pinv_12
Xwl_driver_nand53 en_bar[53] in[53] net[53] vdd gnd pnand2_4
Xwl_driver_inv53 net[53] wl[53] vdd gnd pinv_11
Xwl_driver_inv_en54 en en_bar[54] vdd gnd pinv_12
Xwl_driver_nand54 en_bar[54] in[54] net[54] vdd gnd pnand2_4
Xwl_driver_inv54 net[54] wl[54] vdd gnd pinv_11
Xwl_driver_inv_en55 en en_bar[55] vdd gnd pinv_12
Xwl_driver_nand55 en_bar[55] in[55] net[55] vdd gnd pnand2_4
Xwl_driver_inv55 net[55] wl[55] vdd gnd pinv_11
Xwl_driver_inv_en56 en en_bar[56] vdd gnd pinv_12
Xwl_driver_nand56 en_bar[56] in[56] net[56] vdd gnd pnand2_4
Xwl_driver_inv56 net[56] wl[56] vdd gnd pinv_11
Xwl_driver_inv_en57 en en_bar[57] vdd gnd pinv_12
Xwl_driver_nand57 en_bar[57] in[57] net[57] vdd gnd pnand2_4
Xwl_driver_inv57 net[57] wl[57] vdd gnd pinv_11
Xwl_driver_inv_en58 en en_bar[58] vdd gnd pinv_12
Xwl_driver_nand58 en_bar[58] in[58] net[58] vdd gnd pnand2_4
Xwl_driver_inv58 net[58] wl[58] vdd gnd pinv_11
Xwl_driver_inv_en59 en en_bar[59] vdd gnd pinv_12
Xwl_driver_nand59 en_bar[59] in[59] net[59] vdd gnd pnand2_4
Xwl_driver_inv59 net[59] wl[59] vdd gnd pinv_11
Xwl_driver_inv_en60 en en_bar[60] vdd gnd pinv_12
Xwl_driver_nand60 en_bar[60] in[60] net[60] vdd gnd pnand2_4
Xwl_driver_inv60 net[60] wl[60] vdd gnd pinv_11
Xwl_driver_inv_en61 en en_bar[61] vdd gnd pinv_12
Xwl_driver_nand61 en_bar[61] in[61] net[61] vdd gnd pnand2_4
Xwl_driver_inv61 net[61] wl[61] vdd gnd pinv_11
Xwl_driver_inv_en62 en en_bar[62] vdd gnd pinv_12
Xwl_driver_nand62 en_bar[62] in[62] net[62] vdd gnd pnand2_4
Xwl_driver_inv62 net[62] wl[62] vdd gnd pinv_11
Xwl_driver_inv_en63 en en_bar[63] vdd gnd pinv_12
Xwl_driver_nand63 en_bar[63] in[63] net[63] vdd gnd pnand2_4
Xwl_driver_inv63 net[63] wl[63] vdd gnd pinv_11
Xwl_driver_inv_en64 en en_bar[64] vdd gnd pinv_12
Xwl_driver_nand64 en_bar[64] in[64] net[64] vdd gnd pnand2_4
Xwl_driver_inv64 net[64] wl[64] vdd gnd pinv_11
Xwl_driver_inv_en65 en en_bar[65] vdd gnd pinv_12
Xwl_driver_nand65 en_bar[65] in[65] net[65] vdd gnd pnand2_4
Xwl_driver_inv65 net[65] wl[65] vdd gnd pinv_11
Xwl_driver_inv_en66 en en_bar[66] vdd gnd pinv_12
Xwl_driver_nand66 en_bar[66] in[66] net[66] vdd gnd pnand2_4
Xwl_driver_inv66 net[66] wl[66] vdd gnd pinv_11
Xwl_driver_inv_en67 en en_bar[67] vdd gnd pinv_12
Xwl_driver_nand67 en_bar[67] in[67] net[67] vdd gnd pnand2_4
Xwl_driver_inv67 net[67] wl[67] vdd gnd pinv_11
Xwl_driver_inv_en68 en en_bar[68] vdd gnd pinv_12
Xwl_driver_nand68 en_bar[68] in[68] net[68] vdd gnd pnand2_4
Xwl_driver_inv68 net[68] wl[68] vdd gnd pinv_11
Xwl_driver_inv_en69 en en_bar[69] vdd gnd pinv_12
Xwl_driver_nand69 en_bar[69] in[69] net[69] vdd gnd pnand2_4
Xwl_driver_inv69 net[69] wl[69] vdd gnd pinv_11
Xwl_driver_inv_en70 en en_bar[70] vdd gnd pinv_12
Xwl_driver_nand70 en_bar[70] in[70] net[70] vdd gnd pnand2_4
Xwl_driver_inv70 net[70] wl[70] vdd gnd pinv_11
Xwl_driver_inv_en71 en en_bar[71] vdd gnd pinv_12
Xwl_driver_nand71 en_bar[71] in[71] net[71] vdd gnd pnand2_4
Xwl_driver_inv71 net[71] wl[71] vdd gnd pinv_11
Xwl_driver_inv_en72 en en_bar[72] vdd gnd pinv_12
Xwl_driver_nand72 en_bar[72] in[72] net[72] vdd gnd pnand2_4
Xwl_driver_inv72 net[72] wl[72] vdd gnd pinv_11
Xwl_driver_inv_en73 en en_bar[73] vdd gnd pinv_12
Xwl_driver_nand73 en_bar[73] in[73] net[73] vdd gnd pnand2_4
Xwl_driver_inv73 net[73] wl[73] vdd gnd pinv_11
Xwl_driver_inv_en74 en en_bar[74] vdd gnd pinv_12
Xwl_driver_nand74 en_bar[74] in[74] net[74] vdd gnd pnand2_4
Xwl_driver_inv74 net[74] wl[74] vdd gnd pinv_11
Xwl_driver_inv_en75 en en_bar[75] vdd gnd pinv_12
Xwl_driver_nand75 en_bar[75] in[75] net[75] vdd gnd pnand2_4
Xwl_driver_inv75 net[75] wl[75] vdd gnd pinv_11
Xwl_driver_inv_en76 en en_bar[76] vdd gnd pinv_12
Xwl_driver_nand76 en_bar[76] in[76] net[76] vdd gnd pnand2_4
Xwl_driver_inv76 net[76] wl[76] vdd gnd pinv_11
Xwl_driver_inv_en77 en en_bar[77] vdd gnd pinv_12
Xwl_driver_nand77 en_bar[77] in[77] net[77] vdd gnd pnand2_4
Xwl_driver_inv77 net[77] wl[77] vdd gnd pinv_11
Xwl_driver_inv_en78 en en_bar[78] vdd gnd pinv_12
Xwl_driver_nand78 en_bar[78] in[78] net[78] vdd gnd pnand2_4
Xwl_driver_inv78 net[78] wl[78] vdd gnd pinv_11
Xwl_driver_inv_en79 en en_bar[79] vdd gnd pinv_12
Xwl_driver_nand79 en_bar[79] in[79] net[79] vdd gnd pnand2_4
Xwl_driver_inv79 net[79] wl[79] vdd gnd pinv_11
Xwl_driver_inv_en80 en en_bar[80] vdd gnd pinv_12
Xwl_driver_nand80 en_bar[80] in[80] net[80] vdd gnd pnand2_4
Xwl_driver_inv80 net[80] wl[80] vdd gnd pinv_11
Xwl_driver_inv_en81 en en_bar[81] vdd gnd pinv_12
Xwl_driver_nand81 en_bar[81] in[81] net[81] vdd gnd pnand2_4
Xwl_driver_inv81 net[81] wl[81] vdd gnd pinv_11
Xwl_driver_inv_en82 en en_bar[82] vdd gnd pinv_12
Xwl_driver_nand82 en_bar[82] in[82] net[82] vdd gnd pnand2_4
Xwl_driver_inv82 net[82] wl[82] vdd gnd pinv_11
Xwl_driver_inv_en83 en en_bar[83] vdd gnd pinv_12
Xwl_driver_nand83 en_bar[83] in[83] net[83] vdd gnd pnand2_4
Xwl_driver_inv83 net[83] wl[83] vdd gnd pinv_11
Xwl_driver_inv_en84 en en_bar[84] vdd gnd pinv_12
Xwl_driver_nand84 en_bar[84] in[84] net[84] vdd gnd pnand2_4
Xwl_driver_inv84 net[84] wl[84] vdd gnd pinv_11
Xwl_driver_inv_en85 en en_bar[85] vdd gnd pinv_12
Xwl_driver_nand85 en_bar[85] in[85] net[85] vdd gnd pnand2_4
Xwl_driver_inv85 net[85] wl[85] vdd gnd pinv_11
Xwl_driver_inv_en86 en en_bar[86] vdd gnd pinv_12
Xwl_driver_nand86 en_bar[86] in[86] net[86] vdd gnd pnand2_4
Xwl_driver_inv86 net[86] wl[86] vdd gnd pinv_11
Xwl_driver_inv_en87 en en_bar[87] vdd gnd pinv_12
Xwl_driver_nand87 en_bar[87] in[87] net[87] vdd gnd pnand2_4
Xwl_driver_inv87 net[87] wl[87] vdd gnd pinv_11
Xwl_driver_inv_en88 en en_bar[88] vdd gnd pinv_12
Xwl_driver_nand88 en_bar[88] in[88] net[88] vdd gnd pnand2_4
Xwl_driver_inv88 net[88] wl[88] vdd gnd pinv_11
Xwl_driver_inv_en89 en en_bar[89] vdd gnd pinv_12
Xwl_driver_nand89 en_bar[89] in[89] net[89] vdd gnd pnand2_4
Xwl_driver_inv89 net[89] wl[89] vdd gnd pinv_11
Xwl_driver_inv_en90 en en_bar[90] vdd gnd pinv_12
Xwl_driver_nand90 en_bar[90] in[90] net[90] vdd gnd pnand2_4
Xwl_driver_inv90 net[90] wl[90] vdd gnd pinv_11
Xwl_driver_inv_en91 en en_bar[91] vdd gnd pinv_12
Xwl_driver_nand91 en_bar[91] in[91] net[91] vdd gnd pnand2_4
Xwl_driver_inv91 net[91] wl[91] vdd gnd pinv_11
Xwl_driver_inv_en92 en en_bar[92] vdd gnd pinv_12
Xwl_driver_nand92 en_bar[92] in[92] net[92] vdd gnd pnand2_4
Xwl_driver_inv92 net[92] wl[92] vdd gnd pinv_11
Xwl_driver_inv_en93 en en_bar[93] vdd gnd pinv_12
Xwl_driver_nand93 en_bar[93] in[93] net[93] vdd gnd pnand2_4
Xwl_driver_inv93 net[93] wl[93] vdd gnd pinv_11
Xwl_driver_inv_en94 en en_bar[94] vdd gnd pinv_12
Xwl_driver_nand94 en_bar[94] in[94] net[94] vdd gnd pnand2_4
Xwl_driver_inv94 net[94] wl[94] vdd gnd pinv_11
Xwl_driver_inv_en95 en en_bar[95] vdd gnd pinv_12
Xwl_driver_nand95 en_bar[95] in[95] net[95] vdd gnd pnand2_4
Xwl_driver_inv95 net[95] wl[95] vdd gnd pinv_11
Xwl_driver_inv_en96 en en_bar[96] vdd gnd pinv_12
Xwl_driver_nand96 en_bar[96] in[96] net[96] vdd gnd pnand2_4
Xwl_driver_inv96 net[96] wl[96] vdd gnd pinv_11
Xwl_driver_inv_en97 en en_bar[97] vdd gnd pinv_12
Xwl_driver_nand97 en_bar[97] in[97] net[97] vdd gnd pnand2_4
Xwl_driver_inv97 net[97] wl[97] vdd gnd pinv_11
Xwl_driver_inv_en98 en en_bar[98] vdd gnd pinv_12
Xwl_driver_nand98 en_bar[98] in[98] net[98] vdd gnd pnand2_4
Xwl_driver_inv98 net[98] wl[98] vdd gnd pinv_11
Xwl_driver_inv_en99 en en_bar[99] vdd gnd pinv_12
Xwl_driver_nand99 en_bar[99] in[99] net[99] vdd gnd pnand2_4
Xwl_driver_inv99 net[99] wl[99] vdd gnd pinv_11
Xwl_driver_inv_en100 en en_bar[100] vdd gnd pinv_12
Xwl_driver_nand100 en_bar[100] in[100] net[100] vdd gnd pnand2_4
Xwl_driver_inv100 net[100] wl[100] vdd gnd pinv_11
Xwl_driver_inv_en101 en en_bar[101] vdd gnd pinv_12
Xwl_driver_nand101 en_bar[101] in[101] net[101] vdd gnd pnand2_4
Xwl_driver_inv101 net[101] wl[101] vdd gnd pinv_11
Xwl_driver_inv_en102 en en_bar[102] vdd gnd pinv_12
Xwl_driver_nand102 en_bar[102] in[102] net[102] vdd gnd pnand2_4
Xwl_driver_inv102 net[102] wl[102] vdd gnd pinv_11
Xwl_driver_inv_en103 en en_bar[103] vdd gnd pinv_12
Xwl_driver_nand103 en_bar[103] in[103] net[103] vdd gnd pnand2_4
Xwl_driver_inv103 net[103] wl[103] vdd gnd pinv_11
Xwl_driver_inv_en104 en en_bar[104] vdd gnd pinv_12
Xwl_driver_nand104 en_bar[104] in[104] net[104] vdd gnd pnand2_4
Xwl_driver_inv104 net[104] wl[104] vdd gnd pinv_11
Xwl_driver_inv_en105 en en_bar[105] vdd gnd pinv_12
Xwl_driver_nand105 en_bar[105] in[105] net[105] vdd gnd pnand2_4
Xwl_driver_inv105 net[105] wl[105] vdd gnd pinv_11
Xwl_driver_inv_en106 en en_bar[106] vdd gnd pinv_12
Xwl_driver_nand106 en_bar[106] in[106] net[106] vdd gnd pnand2_4
Xwl_driver_inv106 net[106] wl[106] vdd gnd pinv_11
Xwl_driver_inv_en107 en en_bar[107] vdd gnd pinv_12
Xwl_driver_nand107 en_bar[107] in[107] net[107] vdd gnd pnand2_4
Xwl_driver_inv107 net[107] wl[107] vdd gnd pinv_11
Xwl_driver_inv_en108 en en_bar[108] vdd gnd pinv_12
Xwl_driver_nand108 en_bar[108] in[108] net[108] vdd gnd pnand2_4
Xwl_driver_inv108 net[108] wl[108] vdd gnd pinv_11
Xwl_driver_inv_en109 en en_bar[109] vdd gnd pinv_12
Xwl_driver_nand109 en_bar[109] in[109] net[109] vdd gnd pnand2_4
Xwl_driver_inv109 net[109] wl[109] vdd gnd pinv_11
Xwl_driver_inv_en110 en en_bar[110] vdd gnd pinv_12
Xwl_driver_nand110 en_bar[110] in[110] net[110] vdd gnd pnand2_4
Xwl_driver_inv110 net[110] wl[110] vdd gnd pinv_11
Xwl_driver_inv_en111 en en_bar[111] vdd gnd pinv_12
Xwl_driver_nand111 en_bar[111] in[111] net[111] vdd gnd pnand2_4
Xwl_driver_inv111 net[111] wl[111] vdd gnd pinv_11
Xwl_driver_inv_en112 en en_bar[112] vdd gnd pinv_12
Xwl_driver_nand112 en_bar[112] in[112] net[112] vdd gnd pnand2_4
Xwl_driver_inv112 net[112] wl[112] vdd gnd pinv_11
Xwl_driver_inv_en113 en en_bar[113] vdd gnd pinv_12
Xwl_driver_nand113 en_bar[113] in[113] net[113] vdd gnd pnand2_4
Xwl_driver_inv113 net[113] wl[113] vdd gnd pinv_11
Xwl_driver_inv_en114 en en_bar[114] vdd gnd pinv_12
Xwl_driver_nand114 en_bar[114] in[114] net[114] vdd gnd pnand2_4
Xwl_driver_inv114 net[114] wl[114] vdd gnd pinv_11
Xwl_driver_inv_en115 en en_bar[115] vdd gnd pinv_12
Xwl_driver_nand115 en_bar[115] in[115] net[115] vdd gnd pnand2_4
Xwl_driver_inv115 net[115] wl[115] vdd gnd pinv_11
Xwl_driver_inv_en116 en en_bar[116] vdd gnd pinv_12
Xwl_driver_nand116 en_bar[116] in[116] net[116] vdd gnd pnand2_4
Xwl_driver_inv116 net[116] wl[116] vdd gnd pinv_11
Xwl_driver_inv_en117 en en_bar[117] vdd gnd pinv_12
Xwl_driver_nand117 en_bar[117] in[117] net[117] vdd gnd pnand2_4
Xwl_driver_inv117 net[117] wl[117] vdd gnd pinv_11
Xwl_driver_inv_en118 en en_bar[118] vdd gnd pinv_12
Xwl_driver_nand118 en_bar[118] in[118] net[118] vdd gnd pnand2_4
Xwl_driver_inv118 net[118] wl[118] vdd gnd pinv_11
Xwl_driver_inv_en119 en en_bar[119] vdd gnd pinv_12
Xwl_driver_nand119 en_bar[119] in[119] net[119] vdd gnd pnand2_4
Xwl_driver_inv119 net[119] wl[119] vdd gnd pinv_11
Xwl_driver_inv_en120 en en_bar[120] vdd gnd pinv_12
Xwl_driver_nand120 en_bar[120] in[120] net[120] vdd gnd pnand2_4
Xwl_driver_inv120 net[120] wl[120] vdd gnd pinv_11
Xwl_driver_inv_en121 en en_bar[121] vdd gnd pinv_12
Xwl_driver_nand121 en_bar[121] in[121] net[121] vdd gnd pnand2_4
Xwl_driver_inv121 net[121] wl[121] vdd gnd pinv_11
Xwl_driver_inv_en122 en en_bar[122] vdd gnd pinv_12
Xwl_driver_nand122 en_bar[122] in[122] net[122] vdd gnd pnand2_4
Xwl_driver_inv122 net[122] wl[122] vdd gnd pinv_11
Xwl_driver_inv_en123 en en_bar[123] vdd gnd pinv_12
Xwl_driver_nand123 en_bar[123] in[123] net[123] vdd gnd pnand2_4
Xwl_driver_inv123 net[123] wl[123] vdd gnd pinv_11
Xwl_driver_inv_en124 en en_bar[124] vdd gnd pinv_12
Xwl_driver_nand124 en_bar[124] in[124] net[124] vdd gnd pnand2_4
Xwl_driver_inv124 net[124] wl[124] vdd gnd pinv_11
Xwl_driver_inv_en125 en en_bar[125] vdd gnd pinv_12
Xwl_driver_nand125 en_bar[125] in[125] net[125] vdd gnd pnand2_4
Xwl_driver_inv125 net[125] wl[125] vdd gnd pinv_11
Xwl_driver_inv_en126 en en_bar[126] vdd gnd pinv_12
Xwl_driver_nand126 en_bar[126] in[126] net[126] vdd gnd pnand2_4
Xwl_driver_inv126 net[126] wl[126] vdd gnd pinv_11
Xwl_driver_inv_en127 en en_bar[127] vdd gnd pinv_12
Xwl_driver_nand127 en_bar[127] in[127] net[127] vdd gnd pnand2_4
Xwl_driver_inv127 net[127] wl[127] vdd gnd pinv_11
Xwl_driver_inv_en128 en en_bar[128] vdd gnd pinv_12
Xwl_driver_nand128 en_bar[128] in[128] net[128] vdd gnd pnand2_4
Xwl_driver_inv128 net[128] wl[128] vdd gnd pinv_11
Xwl_driver_inv_en129 en en_bar[129] vdd gnd pinv_12
Xwl_driver_nand129 en_bar[129] in[129] net[129] vdd gnd pnand2_4
Xwl_driver_inv129 net[129] wl[129] vdd gnd pinv_11
Xwl_driver_inv_en130 en en_bar[130] vdd gnd pinv_12
Xwl_driver_nand130 en_bar[130] in[130] net[130] vdd gnd pnand2_4
Xwl_driver_inv130 net[130] wl[130] vdd gnd pinv_11
Xwl_driver_inv_en131 en en_bar[131] vdd gnd pinv_12
Xwl_driver_nand131 en_bar[131] in[131] net[131] vdd gnd pnand2_4
Xwl_driver_inv131 net[131] wl[131] vdd gnd pinv_11
Xwl_driver_inv_en132 en en_bar[132] vdd gnd pinv_12
Xwl_driver_nand132 en_bar[132] in[132] net[132] vdd gnd pnand2_4
Xwl_driver_inv132 net[132] wl[132] vdd gnd pinv_11
Xwl_driver_inv_en133 en en_bar[133] vdd gnd pinv_12
Xwl_driver_nand133 en_bar[133] in[133] net[133] vdd gnd pnand2_4
Xwl_driver_inv133 net[133] wl[133] vdd gnd pinv_11
Xwl_driver_inv_en134 en en_bar[134] vdd gnd pinv_12
Xwl_driver_nand134 en_bar[134] in[134] net[134] vdd gnd pnand2_4
Xwl_driver_inv134 net[134] wl[134] vdd gnd pinv_11
Xwl_driver_inv_en135 en en_bar[135] vdd gnd pinv_12
Xwl_driver_nand135 en_bar[135] in[135] net[135] vdd gnd pnand2_4
Xwl_driver_inv135 net[135] wl[135] vdd gnd pinv_11
Xwl_driver_inv_en136 en en_bar[136] vdd gnd pinv_12
Xwl_driver_nand136 en_bar[136] in[136] net[136] vdd gnd pnand2_4
Xwl_driver_inv136 net[136] wl[136] vdd gnd pinv_11
Xwl_driver_inv_en137 en en_bar[137] vdd gnd pinv_12
Xwl_driver_nand137 en_bar[137] in[137] net[137] vdd gnd pnand2_4
Xwl_driver_inv137 net[137] wl[137] vdd gnd pinv_11
Xwl_driver_inv_en138 en en_bar[138] vdd gnd pinv_12
Xwl_driver_nand138 en_bar[138] in[138] net[138] vdd gnd pnand2_4
Xwl_driver_inv138 net[138] wl[138] vdd gnd pinv_11
Xwl_driver_inv_en139 en en_bar[139] vdd gnd pinv_12
Xwl_driver_nand139 en_bar[139] in[139] net[139] vdd gnd pnand2_4
Xwl_driver_inv139 net[139] wl[139] vdd gnd pinv_11
Xwl_driver_inv_en140 en en_bar[140] vdd gnd pinv_12
Xwl_driver_nand140 en_bar[140] in[140] net[140] vdd gnd pnand2_4
Xwl_driver_inv140 net[140] wl[140] vdd gnd pinv_11
Xwl_driver_inv_en141 en en_bar[141] vdd gnd pinv_12
Xwl_driver_nand141 en_bar[141] in[141] net[141] vdd gnd pnand2_4
Xwl_driver_inv141 net[141] wl[141] vdd gnd pinv_11
Xwl_driver_inv_en142 en en_bar[142] vdd gnd pinv_12
Xwl_driver_nand142 en_bar[142] in[142] net[142] vdd gnd pnand2_4
Xwl_driver_inv142 net[142] wl[142] vdd gnd pinv_11
Xwl_driver_inv_en143 en en_bar[143] vdd gnd pinv_12
Xwl_driver_nand143 en_bar[143] in[143] net[143] vdd gnd pnand2_4
Xwl_driver_inv143 net[143] wl[143] vdd gnd pinv_11
Xwl_driver_inv_en144 en en_bar[144] vdd gnd pinv_12
Xwl_driver_nand144 en_bar[144] in[144] net[144] vdd gnd pnand2_4
Xwl_driver_inv144 net[144] wl[144] vdd gnd pinv_11
Xwl_driver_inv_en145 en en_bar[145] vdd gnd pinv_12
Xwl_driver_nand145 en_bar[145] in[145] net[145] vdd gnd pnand2_4
Xwl_driver_inv145 net[145] wl[145] vdd gnd pinv_11
Xwl_driver_inv_en146 en en_bar[146] vdd gnd pinv_12
Xwl_driver_nand146 en_bar[146] in[146] net[146] vdd gnd pnand2_4
Xwl_driver_inv146 net[146] wl[146] vdd gnd pinv_11
Xwl_driver_inv_en147 en en_bar[147] vdd gnd pinv_12
Xwl_driver_nand147 en_bar[147] in[147] net[147] vdd gnd pnand2_4
Xwl_driver_inv147 net[147] wl[147] vdd gnd pinv_11
Xwl_driver_inv_en148 en en_bar[148] vdd gnd pinv_12
Xwl_driver_nand148 en_bar[148] in[148] net[148] vdd gnd pnand2_4
Xwl_driver_inv148 net[148] wl[148] vdd gnd pinv_11
Xwl_driver_inv_en149 en en_bar[149] vdd gnd pinv_12
Xwl_driver_nand149 en_bar[149] in[149] net[149] vdd gnd pnand2_4
Xwl_driver_inv149 net[149] wl[149] vdd gnd pinv_11
Xwl_driver_inv_en150 en en_bar[150] vdd gnd pinv_12
Xwl_driver_nand150 en_bar[150] in[150] net[150] vdd gnd pnand2_4
Xwl_driver_inv150 net[150] wl[150] vdd gnd pinv_11
Xwl_driver_inv_en151 en en_bar[151] vdd gnd pinv_12
Xwl_driver_nand151 en_bar[151] in[151] net[151] vdd gnd pnand2_4
Xwl_driver_inv151 net[151] wl[151] vdd gnd pinv_11
Xwl_driver_inv_en152 en en_bar[152] vdd gnd pinv_12
Xwl_driver_nand152 en_bar[152] in[152] net[152] vdd gnd pnand2_4
Xwl_driver_inv152 net[152] wl[152] vdd gnd pinv_11
Xwl_driver_inv_en153 en en_bar[153] vdd gnd pinv_12
Xwl_driver_nand153 en_bar[153] in[153] net[153] vdd gnd pnand2_4
Xwl_driver_inv153 net[153] wl[153] vdd gnd pinv_11
Xwl_driver_inv_en154 en en_bar[154] vdd gnd pinv_12
Xwl_driver_nand154 en_bar[154] in[154] net[154] vdd gnd pnand2_4
Xwl_driver_inv154 net[154] wl[154] vdd gnd pinv_11
Xwl_driver_inv_en155 en en_bar[155] vdd gnd pinv_12
Xwl_driver_nand155 en_bar[155] in[155] net[155] vdd gnd pnand2_4
Xwl_driver_inv155 net[155] wl[155] vdd gnd pinv_11
Xwl_driver_inv_en156 en en_bar[156] vdd gnd pinv_12
Xwl_driver_nand156 en_bar[156] in[156] net[156] vdd gnd pnand2_4
Xwl_driver_inv156 net[156] wl[156] vdd gnd pinv_11
Xwl_driver_inv_en157 en en_bar[157] vdd gnd pinv_12
Xwl_driver_nand157 en_bar[157] in[157] net[157] vdd gnd pnand2_4
Xwl_driver_inv157 net[157] wl[157] vdd gnd pinv_11
Xwl_driver_inv_en158 en en_bar[158] vdd gnd pinv_12
Xwl_driver_nand158 en_bar[158] in[158] net[158] vdd gnd pnand2_4
Xwl_driver_inv158 net[158] wl[158] vdd gnd pinv_11
Xwl_driver_inv_en159 en en_bar[159] vdd gnd pinv_12
Xwl_driver_nand159 en_bar[159] in[159] net[159] vdd gnd pnand2_4
Xwl_driver_inv159 net[159] wl[159] vdd gnd pinv_11
Xwl_driver_inv_en160 en en_bar[160] vdd gnd pinv_12
Xwl_driver_nand160 en_bar[160] in[160] net[160] vdd gnd pnand2_4
Xwl_driver_inv160 net[160] wl[160] vdd gnd pinv_11
Xwl_driver_inv_en161 en en_bar[161] vdd gnd pinv_12
Xwl_driver_nand161 en_bar[161] in[161] net[161] vdd gnd pnand2_4
Xwl_driver_inv161 net[161] wl[161] vdd gnd pinv_11
Xwl_driver_inv_en162 en en_bar[162] vdd gnd pinv_12
Xwl_driver_nand162 en_bar[162] in[162] net[162] vdd gnd pnand2_4
Xwl_driver_inv162 net[162] wl[162] vdd gnd pinv_11
Xwl_driver_inv_en163 en en_bar[163] vdd gnd pinv_12
Xwl_driver_nand163 en_bar[163] in[163] net[163] vdd gnd pnand2_4
Xwl_driver_inv163 net[163] wl[163] vdd gnd pinv_11
Xwl_driver_inv_en164 en en_bar[164] vdd gnd pinv_12
Xwl_driver_nand164 en_bar[164] in[164] net[164] vdd gnd pnand2_4
Xwl_driver_inv164 net[164] wl[164] vdd gnd pinv_11
Xwl_driver_inv_en165 en en_bar[165] vdd gnd pinv_12
Xwl_driver_nand165 en_bar[165] in[165] net[165] vdd gnd pnand2_4
Xwl_driver_inv165 net[165] wl[165] vdd gnd pinv_11
Xwl_driver_inv_en166 en en_bar[166] vdd gnd pinv_12
Xwl_driver_nand166 en_bar[166] in[166] net[166] vdd gnd pnand2_4
Xwl_driver_inv166 net[166] wl[166] vdd gnd pinv_11
Xwl_driver_inv_en167 en en_bar[167] vdd gnd pinv_12
Xwl_driver_nand167 en_bar[167] in[167] net[167] vdd gnd pnand2_4
Xwl_driver_inv167 net[167] wl[167] vdd gnd pinv_11
Xwl_driver_inv_en168 en en_bar[168] vdd gnd pinv_12
Xwl_driver_nand168 en_bar[168] in[168] net[168] vdd gnd pnand2_4
Xwl_driver_inv168 net[168] wl[168] vdd gnd pinv_11
Xwl_driver_inv_en169 en en_bar[169] vdd gnd pinv_12
Xwl_driver_nand169 en_bar[169] in[169] net[169] vdd gnd pnand2_4
Xwl_driver_inv169 net[169] wl[169] vdd gnd pinv_11
Xwl_driver_inv_en170 en en_bar[170] vdd gnd pinv_12
Xwl_driver_nand170 en_bar[170] in[170] net[170] vdd gnd pnand2_4
Xwl_driver_inv170 net[170] wl[170] vdd gnd pinv_11
Xwl_driver_inv_en171 en en_bar[171] vdd gnd pinv_12
Xwl_driver_nand171 en_bar[171] in[171] net[171] vdd gnd pnand2_4
Xwl_driver_inv171 net[171] wl[171] vdd gnd pinv_11
Xwl_driver_inv_en172 en en_bar[172] vdd gnd pinv_12
Xwl_driver_nand172 en_bar[172] in[172] net[172] vdd gnd pnand2_4
Xwl_driver_inv172 net[172] wl[172] vdd gnd pinv_11
Xwl_driver_inv_en173 en en_bar[173] vdd gnd pinv_12
Xwl_driver_nand173 en_bar[173] in[173] net[173] vdd gnd pnand2_4
Xwl_driver_inv173 net[173] wl[173] vdd gnd pinv_11
Xwl_driver_inv_en174 en en_bar[174] vdd gnd pinv_12
Xwl_driver_nand174 en_bar[174] in[174] net[174] vdd gnd pnand2_4
Xwl_driver_inv174 net[174] wl[174] vdd gnd pinv_11
Xwl_driver_inv_en175 en en_bar[175] vdd gnd pinv_12
Xwl_driver_nand175 en_bar[175] in[175] net[175] vdd gnd pnand2_4
Xwl_driver_inv175 net[175] wl[175] vdd gnd pinv_11
Xwl_driver_inv_en176 en en_bar[176] vdd gnd pinv_12
Xwl_driver_nand176 en_bar[176] in[176] net[176] vdd gnd pnand2_4
Xwl_driver_inv176 net[176] wl[176] vdd gnd pinv_11
Xwl_driver_inv_en177 en en_bar[177] vdd gnd pinv_12
Xwl_driver_nand177 en_bar[177] in[177] net[177] vdd gnd pnand2_4
Xwl_driver_inv177 net[177] wl[177] vdd gnd pinv_11
Xwl_driver_inv_en178 en en_bar[178] vdd gnd pinv_12
Xwl_driver_nand178 en_bar[178] in[178] net[178] vdd gnd pnand2_4
Xwl_driver_inv178 net[178] wl[178] vdd gnd pinv_11
Xwl_driver_inv_en179 en en_bar[179] vdd gnd pinv_12
Xwl_driver_nand179 en_bar[179] in[179] net[179] vdd gnd pnand2_4
Xwl_driver_inv179 net[179] wl[179] vdd gnd pinv_11
Xwl_driver_inv_en180 en en_bar[180] vdd gnd pinv_12
Xwl_driver_nand180 en_bar[180] in[180] net[180] vdd gnd pnand2_4
Xwl_driver_inv180 net[180] wl[180] vdd gnd pinv_11
Xwl_driver_inv_en181 en en_bar[181] vdd gnd pinv_12
Xwl_driver_nand181 en_bar[181] in[181] net[181] vdd gnd pnand2_4
Xwl_driver_inv181 net[181] wl[181] vdd gnd pinv_11
Xwl_driver_inv_en182 en en_bar[182] vdd gnd pinv_12
Xwl_driver_nand182 en_bar[182] in[182] net[182] vdd gnd pnand2_4
Xwl_driver_inv182 net[182] wl[182] vdd gnd pinv_11
Xwl_driver_inv_en183 en en_bar[183] vdd gnd pinv_12
Xwl_driver_nand183 en_bar[183] in[183] net[183] vdd gnd pnand2_4
Xwl_driver_inv183 net[183] wl[183] vdd gnd pinv_11
Xwl_driver_inv_en184 en en_bar[184] vdd gnd pinv_12
Xwl_driver_nand184 en_bar[184] in[184] net[184] vdd gnd pnand2_4
Xwl_driver_inv184 net[184] wl[184] vdd gnd pinv_11
Xwl_driver_inv_en185 en en_bar[185] vdd gnd pinv_12
Xwl_driver_nand185 en_bar[185] in[185] net[185] vdd gnd pnand2_4
Xwl_driver_inv185 net[185] wl[185] vdd gnd pinv_11
Xwl_driver_inv_en186 en en_bar[186] vdd gnd pinv_12
Xwl_driver_nand186 en_bar[186] in[186] net[186] vdd gnd pnand2_4
Xwl_driver_inv186 net[186] wl[186] vdd gnd pinv_11
Xwl_driver_inv_en187 en en_bar[187] vdd gnd pinv_12
Xwl_driver_nand187 en_bar[187] in[187] net[187] vdd gnd pnand2_4
Xwl_driver_inv187 net[187] wl[187] vdd gnd pinv_11
Xwl_driver_inv_en188 en en_bar[188] vdd gnd pinv_12
Xwl_driver_nand188 en_bar[188] in[188] net[188] vdd gnd pnand2_4
Xwl_driver_inv188 net[188] wl[188] vdd gnd pinv_11
Xwl_driver_inv_en189 en en_bar[189] vdd gnd pinv_12
Xwl_driver_nand189 en_bar[189] in[189] net[189] vdd gnd pnand2_4
Xwl_driver_inv189 net[189] wl[189] vdd gnd pinv_11
Xwl_driver_inv_en190 en en_bar[190] vdd gnd pinv_12
Xwl_driver_nand190 en_bar[190] in[190] net[190] vdd gnd pnand2_4
Xwl_driver_inv190 net[190] wl[190] vdd gnd pinv_11
Xwl_driver_inv_en191 en en_bar[191] vdd gnd pinv_12
Xwl_driver_nand191 en_bar[191] in[191] net[191] vdd gnd pnand2_4
Xwl_driver_inv191 net[191] wl[191] vdd gnd pinv_11
Xwl_driver_inv_en192 en en_bar[192] vdd gnd pinv_12
Xwl_driver_nand192 en_bar[192] in[192] net[192] vdd gnd pnand2_4
Xwl_driver_inv192 net[192] wl[192] vdd gnd pinv_11
Xwl_driver_inv_en193 en en_bar[193] vdd gnd pinv_12
Xwl_driver_nand193 en_bar[193] in[193] net[193] vdd gnd pnand2_4
Xwl_driver_inv193 net[193] wl[193] vdd gnd pinv_11
Xwl_driver_inv_en194 en en_bar[194] vdd gnd pinv_12
Xwl_driver_nand194 en_bar[194] in[194] net[194] vdd gnd pnand2_4
Xwl_driver_inv194 net[194] wl[194] vdd gnd pinv_11
Xwl_driver_inv_en195 en en_bar[195] vdd gnd pinv_12
Xwl_driver_nand195 en_bar[195] in[195] net[195] vdd gnd pnand2_4
Xwl_driver_inv195 net[195] wl[195] vdd gnd pinv_11
Xwl_driver_inv_en196 en en_bar[196] vdd gnd pinv_12
Xwl_driver_nand196 en_bar[196] in[196] net[196] vdd gnd pnand2_4
Xwl_driver_inv196 net[196] wl[196] vdd gnd pinv_11
Xwl_driver_inv_en197 en en_bar[197] vdd gnd pinv_12
Xwl_driver_nand197 en_bar[197] in[197] net[197] vdd gnd pnand2_4
Xwl_driver_inv197 net[197] wl[197] vdd gnd pinv_11
Xwl_driver_inv_en198 en en_bar[198] vdd gnd pinv_12
Xwl_driver_nand198 en_bar[198] in[198] net[198] vdd gnd pnand2_4
Xwl_driver_inv198 net[198] wl[198] vdd gnd pinv_11
Xwl_driver_inv_en199 en en_bar[199] vdd gnd pinv_12
Xwl_driver_nand199 en_bar[199] in[199] net[199] vdd gnd pnand2_4
Xwl_driver_inv199 net[199] wl[199] vdd gnd pinv_11
Xwl_driver_inv_en200 en en_bar[200] vdd gnd pinv_12
Xwl_driver_nand200 en_bar[200] in[200] net[200] vdd gnd pnand2_4
Xwl_driver_inv200 net[200] wl[200] vdd gnd pinv_11
Xwl_driver_inv_en201 en en_bar[201] vdd gnd pinv_12
Xwl_driver_nand201 en_bar[201] in[201] net[201] vdd gnd pnand2_4
Xwl_driver_inv201 net[201] wl[201] vdd gnd pinv_11
Xwl_driver_inv_en202 en en_bar[202] vdd gnd pinv_12
Xwl_driver_nand202 en_bar[202] in[202] net[202] vdd gnd pnand2_4
Xwl_driver_inv202 net[202] wl[202] vdd gnd pinv_11
Xwl_driver_inv_en203 en en_bar[203] vdd gnd pinv_12
Xwl_driver_nand203 en_bar[203] in[203] net[203] vdd gnd pnand2_4
Xwl_driver_inv203 net[203] wl[203] vdd gnd pinv_11
Xwl_driver_inv_en204 en en_bar[204] vdd gnd pinv_12
Xwl_driver_nand204 en_bar[204] in[204] net[204] vdd gnd pnand2_4
Xwl_driver_inv204 net[204] wl[204] vdd gnd pinv_11
Xwl_driver_inv_en205 en en_bar[205] vdd gnd pinv_12
Xwl_driver_nand205 en_bar[205] in[205] net[205] vdd gnd pnand2_4
Xwl_driver_inv205 net[205] wl[205] vdd gnd pinv_11
Xwl_driver_inv_en206 en en_bar[206] vdd gnd pinv_12
Xwl_driver_nand206 en_bar[206] in[206] net[206] vdd gnd pnand2_4
Xwl_driver_inv206 net[206] wl[206] vdd gnd pinv_11
Xwl_driver_inv_en207 en en_bar[207] vdd gnd pinv_12
Xwl_driver_nand207 en_bar[207] in[207] net[207] vdd gnd pnand2_4
Xwl_driver_inv207 net[207] wl[207] vdd gnd pinv_11
Xwl_driver_inv_en208 en en_bar[208] vdd gnd pinv_12
Xwl_driver_nand208 en_bar[208] in[208] net[208] vdd gnd pnand2_4
Xwl_driver_inv208 net[208] wl[208] vdd gnd pinv_11
Xwl_driver_inv_en209 en en_bar[209] vdd gnd pinv_12
Xwl_driver_nand209 en_bar[209] in[209] net[209] vdd gnd pnand2_4
Xwl_driver_inv209 net[209] wl[209] vdd gnd pinv_11
Xwl_driver_inv_en210 en en_bar[210] vdd gnd pinv_12
Xwl_driver_nand210 en_bar[210] in[210] net[210] vdd gnd pnand2_4
Xwl_driver_inv210 net[210] wl[210] vdd gnd pinv_11
Xwl_driver_inv_en211 en en_bar[211] vdd gnd pinv_12
Xwl_driver_nand211 en_bar[211] in[211] net[211] vdd gnd pnand2_4
Xwl_driver_inv211 net[211] wl[211] vdd gnd pinv_11
Xwl_driver_inv_en212 en en_bar[212] vdd gnd pinv_12
Xwl_driver_nand212 en_bar[212] in[212] net[212] vdd gnd pnand2_4
Xwl_driver_inv212 net[212] wl[212] vdd gnd pinv_11
Xwl_driver_inv_en213 en en_bar[213] vdd gnd pinv_12
Xwl_driver_nand213 en_bar[213] in[213] net[213] vdd gnd pnand2_4
Xwl_driver_inv213 net[213] wl[213] vdd gnd pinv_11
Xwl_driver_inv_en214 en en_bar[214] vdd gnd pinv_12
Xwl_driver_nand214 en_bar[214] in[214] net[214] vdd gnd pnand2_4
Xwl_driver_inv214 net[214] wl[214] vdd gnd pinv_11
Xwl_driver_inv_en215 en en_bar[215] vdd gnd pinv_12
Xwl_driver_nand215 en_bar[215] in[215] net[215] vdd gnd pnand2_4
Xwl_driver_inv215 net[215] wl[215] vdd gnd pinv_11
Xwl_driver_inv_en216 en en_bar[216] vdd gnd pinv_12
Xwl_driver_nand216 en_bar[216] in[216] net[216] vdd gnd pnand2_4
Xwl_driver_inv216 net[216] wl[216] vdd gnd pinv_11
Xwl_driver_inv_en217 en en_bar[217] vdd gnd pinv_12
Xwl_driver_nand217 en_bar[217] in[217] net[217] vdd gnd pnand2_4
Xwl_driver_inv217 net[217] wl[217] vdd gnd pinv_11
Xwl_driver_inv_en218 en en_bar[218] vdd gnd pinv_12
Xwl_driver_nand218 en_bar[218] in[218] net[218] vdd gnd pnand2_4
Xwl_driver_inv218 net[218] wl[218] vdd gnd pinv_11
Xwl_driver_inv_en219 en en_bar[219] vdd gnd pinv_12
Xwl_driver_nand219 en_bar[219] in[219] net[219] vdd gnd pnand2_4
Xwl_driver_inv219 net[219] wl[219] vdd gnd pinv_11
Xwl_driver_inv_en220 en en_bar[220] vdd gnd pinv_12
Xwl_driver_nand220 en_bar[220] in[220] net[220] vdd gnd pnand2_4
Xwl_driver_inv220 net[220] wl[220] vdd gnd pinv_11
Xwl_driver_inv_en221 en en_bar[221] vdd gnd pinv_12
Xwl_driver_nand221 en_bar[221] in[221] net[221] vdd gnd pnand2_4
Xwl_driver_inv221 net[221] wl[221] vdd gnd pinv_11
Xwl_driver_inv_en222 en en_bar[222] vdd gnd pinv_12
Xwl_driver_nand222 en_bar[222] in[222] net[222] vdd gnd pnand2_4
Xwl_driver_inv222 net[222] wl[222] vdd gnd pinv_11
Xwl_driver_inv_en223 en en_bar[223] vdd gnd pinv_12
Xwl_driver_nand223 en_bar[223] in[223] net[223] vdd gnd pnand2_4
Xwl_driver_inv223 net[223] wl[223] vdd gnd pinv_11
Xwl_driver_inv_en224 en en_bar[224] vdd gnd pinv_12
Xwl_driver_nand224 en_bar[224] in[224] net[224] vdd gnd pnand2_4
Xwl_driver_inv224 net[224] wl[224] vdd gnd pinv_11
Xwl_driver_inv_en225 en en_bar[225] vdd gnd pinv_12
Xwl_driver_nand225 en_bar[225] in[225] net[225] vdd gnd pnand2_4
Xwl_driver_inv225 net[225] wl[225] vdd gnd pinv_11
Xwl_driver_inv_en226 en en_bar[226] vdd gnd pinv_12
Xwl_driver_nand226 en_bar[226] in[226] net[226] vdd gnd pnand2_4
Xwl_driver_inv226 net[226] wl[226] vdd gnd pinv_11
Xwl_driver_inv_en227 en en_bar[227] vdd gnd pinv_12
Xwl_driver_nand227 en_bar[227] in[227] net[227] vdd gnd pnand2_4
Xwl_driver_inv227 net[227] wl[227] vdd gnd pinv_11
Xwl_driver_inv_en228 en en_bar[228] vdd gnd pinv_12
Xwl_driver_nand228 en_bar[228] in[228] net[228] vdd gnd pnand2_4
Xwl_driver_inv228 net[228] wl[228] vdd gnd pinv_11
Xwl_driver_inv_en229 en en_bar[229] vdd gnd pinv_12
Xwl_driver_nand229 en_bar[229] in[229] net[229] vdd gnd pnand2_4
Xwl_driver_inv229 net[229] wl[229] vdd gnd pinv_11
Xwl_driver_inv_en230 en en_bar[230] vdd gnd pinv_12
Xwl_driver_nand230 en_bar[230] in[230] net[230] vdd gnd pnand2_4
Xwl_driver_inv230 net[230] wl[230] vdd gnd pinv_11
Xwl_driver_inv_en231 en en_bar[231] vdd gnd pinv_12
Xwl_driver_nand231 en_bar[231] in[231] net[231] vdd gnd pnand2_4
Xwl_driver_inv231 net[231] wl[231] vdd gnd pinv_11
Xwl_driver_inv_en232 en en_bar[232] vdd gnd pinv_12
Xwl_driver_nand232 en_bar[232] in[232] net[232] vdd gnd pnand2_4
Xwl_driver_inv232 net[232] wl[232] vdd gnd pinv_11
Xwl_driver_inv_en233 en en_bar[233] vdd gnd pinv_12
Xwl_driver_nand233 en_bar[233] in[233] net[233] vdd gnd pnand2_4
Xwl_driver_inv233 net[233] wl[233] vdd gnd pinv_11
Xwl_driver_inv_en234 en en_bar[234] vdd gnd pinv_12
Xwl_driver_nand234 en_bar[234] in[234] net[234] vdd gnd pnand2_4
Xwl_driver_inv234 net[234] wl[234] vdd gnd pinv_11
Xwl_driver_inv_en235 en en_bar[235] vdd gnd pinv_12
Xwl_driver_nand235 en_bar[235] in[235] net[235] vdd gnd pnand2_4
Xwl_driver_inv235 net[235] wl[235] vdd gnd pinv_11
Xwl_driver_inv_en236 en en_bar[236] vdd gnd pinv_12
Xwl_driver_nand236 en_bar[236] in[236] net[236] vdd gnd pnand2_4
Xwl_driver_inv236 net[236] wl[236] vdd gnd pinv_11
Xwl_driver_inv_en237 en en_bar[237] vdd gnd pinv_12
Xwl_driver_nand237 en_bar[237] in[237] net[237] vdd gnd pnand2_4
Xwl_driver_inv237 net[237] wl[237] vdd gnd pinv_11
Xwl_driver_inv_en238 en en_bar[238] vdd gnd pinv_12
Xwl_driver_nand238 en_bar[238] in[238] net[238] vdd gnd pnand2_4
Xwl_driver_inv238 net[238] wl[238] vdd gnd pinv_11
Xwl_driver_inv_en239 en en_bar[239] vdd gnd pinv_12
Xwl_driver_nand239 en_bar[239] in[239] net[239] vdd gnd pnand2_4
Xwl_driver_inv239 net[239] wl[239] vdd gnd pinv_11
Xwl_driver_inv_en240 en en_bar[240] vdd gnd pinv_12
Xwl_driver_nand240 en_bar[240] in[240] net[240] vdd gnd pnand2_4
Xwl_driver_inv240 net[240] wl[240] vdd gnd pinv_11
Xwl_driver_inv_en241 en en_bar[241] vdd gnd pinv_12
Xwl_driver_nand241 en_bar[241] in[241] net[241] vdd gnd pnand2_4
Xwl_driver_inv241 net[241] wl[241] vdd gnd pinv_11
Xwl_driver_inv_en242 en en_bar[242] vdd gnd pinv_12
Xwl_driver_nand242 en_bar[242] in[242] net[242] vdd gnd pnand2_4
Xwl_driver_inv242 net[242] wl[242] vdd gnd pinv_11
Xwl_driver_inv_en243 en en_bar[243] vdd gnd pinv_12
Xwl_driver_nand243 en_bar[243] in[243] net[243] vdd gnd pnand2_4
Xwl_driver_inv243 net[243] wl[243] vdd gnd pinv_11
Xwl_driver_inv_en244 en en_bar[244] vdd gnd pinv_12
Xwl_driver_nand244 en_bar[244] in[244] net[244] vdd gnd pnand2_4
Xwl_driver_inv244 net[244] wl[244] vdd gnd pinv_11
Xwl_driver_inv_en245 en en_bar[245] vdd gnd pinv_12
Xwl_driver_nand245 en_bar[245] in[245] net[245] vdd gnd pnand2_4
Xwl_driver_inv245 net[245] wl[245] vdd gnd pinv_11
Xwl_driver_inv_en246 en en_bar[246] vdd gnd pinv_12
Xwl_driver_nand246 en_bar[246] in[246] net[246] vdd gnd pnand2_4
Xwl_driver_inv246 net[246] wl[246] vdd gnd pinv_11
Xwl_driver_inv_en247 en en_bar[247] vdd gnd pinv_12
Xwl_driver_nand247 en_bar[247] in[247] net[247] vdd gnd pnand2_4
Xwl_driver_inv247 net[247] wl[247] vdd gnd pinv_11
Xwl_driver_inv_en248 en en_bar[248] vdd gnd pinv_12
Xwl_driver_nand248 en_bar[248] in[248] net[248] vdd gnd pnand2_4
Xwl_driver_inv248 net[248] wl[248] vdd gnd pinv_11
Xwl_driver_inv_en249 en en_bar[249] vdd gnd pinv_12
Xwl_driver_nand249 en_bar[249] in[249] net[249] vdd gnd pnand2_4
Xwl_driver_inv249 net[249] wl[249] vdd gnd pinv_11
Xwl_driver_inv_en250 en en_bar[250] vdd gnd pinv_12
Xwl_driver_nand250 en_bar[250] in[250] net[250] vdd gnd pnand2_4
Xwl_driver_inv250 net[250] wl[250] vdd gnd pinv_11
Xwl_driver_inv_en251 en en_bar[251] vdd gnd pinv_12
Xwl_driver_nand251 en_bar[251] in[251] net[251] vdd gnd pnand2_4
Xwl_driver_inv251 net[251] wl[251] vdd gnd pinv_11
Xwl_driver_inv_en252 en en_bar[252] vdd gnd pinv_12
Xwl_driver_nand252 en_bar[252] in[252] net[252] vdd gnd pnand2_4
Xwl_driver_inv252 net[252] wl[252] vdd gnd pinv_11
Xwl_driver_inv_en253 en en_bar[253] vdd gnd pinv_12
Xwl_driver_nand253 en_bar[253] in[253] net[253] vdd gnd pnand2_4
Xwl_driver_inv253 net[253] wl[253] vdd gnd pinv_11
Xwl_driver_inv_en254 en en_bar[254] vdd gnd pinv_12
Xwl_driver_nand254 en_bar[254] in[254] net[254] vdd gnd pnand2_4
Xwl_driver_inv254 net[254] wl[254] vdd gnd pinv_11
Xwl_driver_inv_en255 en en_bar[255] vdd gnd pinv_12
Xwl_driver_nand255 en_bar[255] in[255] net[255] vdd gnd pnand2_4
Xwl_driver_inv255 net[255] wl[255] vdd gnd pinv_11
Xwl_driver_inv_en256 en en_bar[256] vdd gnd pinv_12
Xwl_driver_nand256 en_bar[256] in[256] net[256] vdd gnd pnand2_4
Xwl_driver_inv256 net[256] wl[256] vdd gnd pinv_11
Xwl_driver_inv_en257 en en_bar[257] vdd gnd pinv_12
Xwl_driver_nand257 en_bar[257] in[257] net[257] vdd gnd pnand2_4
Xwl_driver_inv257 net[257] wl[257] vdd gnd pinv_11
Xwl_driver_inv_en258 en en_bar[258] vdd gnd pinv_12
Xwl_driver_nand258 en_bar[258] in[258] net[258] vdd gnd pnand2_4
Xwl_driver_inv258 net[258] wl[258] vdd gnd pinv_11
Xwl_driver_inv_en259 en en_bar[259] vdd gnd pinv_12
Xwl_driver_nand259 en_bar[259] in[259] net[259] vdd gnd pnand2_4
Xwl_driver_inv259 net[259] wl[259] vdd gnd pinv_11
Xwl_driver_inv_en260 en en_bar[260] vdd gnd pinv_12
Xwl_driver_nand260 en_bar[260] in[260] net[260] vdd gnd pnand2_4
Xwl_driver_inv260 net[260] wl[260] vdd gnd pinv_11
Xwl_driver_inv_en261 en en_bar[261] vdd gnd pinv_12
Xwl_driver_nand261 en_bar[261] in[261] net[261] vdd gnd pnand2_4
Xwl_driver_inv261 net[261] wl[261] vdd gnd pinv_11
Xwl_driver_inv_en262 en en_bar[262] vdd gnd pinv_12
Xwl_driver_nand262 en_bar[262] in[262] net[262] vdd gnd pnand2_4
Xwl_driver_inv262 net[262] wl[262] vdd gnd pinv_11
Xwl_driver_inv_en263 en en_bar[263] vdd gnd pinv_12
Xwl_driver_nand263 en_bar[263] in[263] net[263] vdd gnd pnand2_4
Xwl_driver_inv263 net[263] wl[263] vdd gnd pinv_11
Xwl_driver_inv_en264 en en_bar[264] vdd gnd pinv_12
Xwl_driver_nand264 en_bar[264] in[264] net[264] vdd gnd pnand2_4
Xwl_driver_inv264 net[264] wl[264] vdd gnd pinv_11
Xwl_driver_inv_en265 en en_bar[265] vdd gnd pinv_12
Xwl_driver_nand265 en_bar[265] in[265] net[265] vdd gnd pnand2_4
Xwl_driver_inv265 net[265] wl[265] vdd gnd pinv_11
Xwl_driver_inv_en266 en en_bar[266] vdd gnd pinv_12
Xwl_driver_nand266 en_bar[266] in[266] net[266] vdd gnd pnand2_4
Xwl_driver_inv266 net[266] wl[266] vdd gnd pinv_11
Xwl_driver_inv_en267 en en_bar[267] vdd gnd pinv_12
Xwl_driver_nand267 en_bar[267] in[267] net[267] vdd gnd pnand2_4
Xwl_driver_inv267 net[267] wl[267] vdd gnd pinv_11
Xwl_driver_inv_en268 en en_bar[268] vdd gnd pinv_12
Xwl_driver_nand268 en_bar[268] in[268] net[268] vdd gnd pnand2_4
Xwl_driver_inv268 net[268] wl[268] vdd gnd pinv_11
Xwl_driver_inv_en269 en en_bar[269] vdd gnd pinv_12
Xwl_driver_nand269 en_bar[269] in[269] net[269] vdd gnd pnand2_4
Xwl_driver_inv269 net[269] wl[269] vdd gnd pinv_11
Xwl_driver_inv_en270 en en_bar[270] vdd gnd pinv_12
Xwl_driver_nand270 en_bar[270] in[270] net[270] vdd gnd pnand2_4
Xwl_driver_inv270 net[270] wl[270] vdd gnd pinv_11
Xwl_driver_inv_en271 en en_bar[271] vdd gnd pinv_12
Xwl_driver_nand271 en_bar[271] in[271] net[271] vdd gnd pnand2_4
Xwl_driver_inv271 net[271] wl[271] vdd gnd pinv_11
Xwl_driver_inv_en272 en en_bar[272] vdd gnd pinv_12
Xwl_driver_nand272 en_bar[272] in[272] net[272] vdd gnd pnand2_4
Xwl_driver_inv272 net[272] wl[272] vdd gnd pinv_11
Xwl_driver_inv_en273 en en_bar[273] vdd gnd pinv_12
Xwl_driver_nand273 en_bar[273] in[273] net[273] vdd gnd pnand2_4
Xwl_driver_inv273 net[273] wl[273] vdd gnd pinv_11
Xwl_driver_inv_en274 en en_bar[274] vdd gnd pinv_12
Xwl_driver_nand274 en_bar[274] in[274] net[274] vdd gnd pnand2_4
Xwl_driver_inv274 net[274] wl[274] vdd gnd pinv_11
Xwl_driver_inv_en275 en en_bar[275] vdd gnd pinv_12
Xwl_driver_nand275 en_bar[275] in[275] net[275] vdd gnd pnand2_4
Xwl_driver_inv275 net[275] wl[275] vdd gnd pinv_11
Xwl_driver_inv_en276 en en_bar[276] vdd gnd pinv_12
Xwl_driver_nand276 en_bar[276] in[276] net[276] vdd gnd pnand2_4
Xwl_driver_inv276 net[276] wl[276] vdd gnd pinv_11
Xwl_driver_inv_en277 en en_bar[277] vdd gnd pinv_12
Xwl_driver_nand277 en_bar[277] in[277] net[277] vdd gnd pnand2_4
Xwl_driver_inv277 net[277] wl[277] vdd gnd pinv_11
Xwl_driver_inv_en278 en en_bar[278] vdd gnd pinv_12
Xwl_driver_nand278 en_bar[278] in[278] net[278] vdd gnd pnand2_4
Xwl_driver_inv278 net[278] wl[278] vdd gnd pinv_11
Xwl_driver_inv_en279 en en_bar[279] vdd gnd pinv_12
Xwl_driver_nand279 en_bar[279] in[279] net[279] vdd gnd pnand2_4
Xwl_driver_inv279 net[279] wl[279] vdd gnd pinv_11
Xwl_driver_inv_en280 en en_bar[280] vdd gnd pinv_12
Xwl_driver_nand280 en_bar[280] in[280] net[280] vdd gnd pnand2_4
Xwl_driver_inv280 net[280] wl[280] vdd gnd pinv_11
Xwl_driver_inv_en281 en en_bar[281] vdd gnd pinv_12
Xwl_driver_nand281 en_bar[281] in[281] net[281] vdd gnd pnand2_4
Xwl_driver_inv281 net[281] wl[281] vdd gnd pinv_11
Xwl_driver_inv_en282 en en_bar[282] vdd gnd pinv_12
Xwl_driver_nand282 en_bar[282] in[282] net[282] vdd gnd pnand2_4
Xwl_driver_inv282 net[282] wl[282] vdd gnd pinv_11
Xwl_driver_inv_en283 en en_bar[283] vdd gnd pinv_12
Xwl_driver_nand283 en_bar[283] in[283] net[283] vdd gnd pnand2_4
Xwl_driver_inv283 net[283] wl[283] vdd gnd pinv_11
Xwl_driver_inv_en284 en en_bar[284] vdd gnd pinv_12
Xwl_driver_nand284 en_bar[284] in[284] net[284] vdd gnd pnand2_4
Xwl_driver_inv284 net[284] wl[284] vdd gnd pinv_11
Xwl_driver_inv_en285 en en_bar[285] vdd gnd pinv_12
Xwl_driver_nand285 en_bar[285] in[285] net[285] vdd gnd pnand2_4
Xwl_driver_inv285 net[285] wl[285] vdd gnd pinv_11
Xwl_driver_inv_en286 en en_bar[286] vdd gnd pinv_12
Xwl_driver_nand286 en_bar[286] in[286] net[286] vdd gnd pnand2_4
Xwl_driver_inv286 net[286] wl[286] vdd gnd pinv_11
Xwl_driver_inv_en287 en en_bar[287] vdd gnd pinv_12
Xwl_driver_nand287 en_bar[287] in[287] net[287] vdd gnd pnand2_4
Xwl_driver_inv287 net[287] wl[287] vdd gnd pinv_11
Xwl_driver_inv_en288 en en_bar[288] vdd gnd pinv_12
Xwl_driver_nand288 en_bar[288] in[288] net[288] vdd gnd pnand2_4
Xwl_driver_inv288 net[288] wl[288] vdd gnd pinv_11
Xwl_driver_inv_en289 en en_bar[289] vdd gnd pinv_12
Xwl_driver_nand289 en_bar[289] in[289] net[289] vdd gnd pnand2_4
Xwl_driver_inv289 net[289] wl[289] vdd gnd pinv_11
Xwl_driver_inv_en290 en en_bar[290] vdd gnd pinv_12
Xwl_driver_nand290 en_bar[290] in[290] net[290] vdd gnd pnand2_4
Xwl_driver_inv290 net[290] wl[290] vdd gnd pinv_11
Xwl_driver_inv_en291 en en_bar[291] vdd gnd pinv_12
Xwl_driver_nand291 en_bar[291] in[291] net[291] vdd gnd pnand2_4
Xwl_driver_inv291 net[291] wl[291] vdd gnd pinv_11
Xwl_driver_inv_en292 en en_bar[292] vdd gnd pinv_12
Xwl_driver_nand292 en_bar[292] in[292] net[292] vdd gnd pnand2_4
Xwl_driver_inv292 net[292] wl[292] vdd gnd pinv_11
Xwl_driver_inv_en293 en en_bar[293] vdd gnd pinv_12
Xwl_driver_nand293 en_bar[293] in[293] net[293] vdd gnd pnand2_4
Xwl_driver_inv293 net[293] wl[293] vdd gnd pinv_11
Xwl_driver_inv_en294 en en_bar[294] vdd gnd pinv_12
Xwl_driver_nand294 en_bar[294] in[294] net[294] vdd gnd pnand2_4
Xwl_driver_inv294 net[294] wl[294] vdd gnd pinv_11
Xwl_driver_inv_en295 en en_bar[295] vdd gnd pinv_12
Xwl_driver_nand295 en_bar[295] in[295] net[295] vdd gnd pnand2_4
Xwl_driver_inv295 net[295] wl[295] vdd gnd pinv_11
Xwl_driver_inv_en296 en en_bar[296] vdd gnd pinv_12
Xwl_driver_nand296 en_bar[296] in[296] net[296] vdd gnd pnand2_4
Xwl_driver_inv296 net[296] wl[296] vdd gnd pinv_11
Xwl_driver_inv_en297 en en_bar[297] vdd gnd pinv_12
Xwl_driver_nand297 en_bar[297] in[297] net[297] vdd gnd pnand2_4
Xwl_driver_inv297 net[297] wl[297] vdd gnd pinv_11
Xwl_driver_inv_en298 en en_bar[298] vdd gnd pinv_12
Xwl_driver_nand298 en_bar[298] in[298] net[298] vdd gnd pnand2_4
Xwl_driver_inv298 net[298] wl[298] vdd gnd pinv_11
Xwl_driver_inv_en299 en en_bar[299] vdd gnd pinv_12
Xwl_driver_nand299 en_bar[299] in[299] net[299] vdd gnd pnand2_4
Xwl_driver_inv299 net[299] wl[299] vdd gnd pinv_11
Xwl_driver_inv_en300 en en_bar[300] vdd gnd pinv_12
Xwl_driver_nand300 en_bar[300] in[300] net[300] vdd gnd pnand2_4
Xwl_driver_inv300 net[300] wl[300] vdd gnd pinv_11
Xwl_driver_inv_en301 en en_bar[301] vdd gnd pinv_12
Xwl_driver_nand301 en_bar[301] in[301] net[301] vdd gnd pnand2_4
Xwl_driver_inv301 net[301] wl[301] vdd gnd pinv_11
Xwl_driver_inv_en302 en en_bar[302] vdd gnd pinv_12
Xwl_driver_nand302 en_bar[302] in[302] net[302] vdd gnd pnand2_4
Xwl_driver_inv302 net[302] wl[302] vdd gnd pinv_11
Xwl_driver_inv_en303 en en_bar[303] vdd gnd pinv_12
Xwl_driver_nand303 en_bar[303] in[303] net[303] vdd gnd pnand2_4
Xwl_driver_inv303 net[303] wl[303] vdd gnd pinv_11
Xwl_driver_inv_en304 en en_bar[304] vdd gnd pinv_12
Xwl_driver_nand304 en_bar[304] in[304] net[304] vdd gnd pnand2_4
Xwl_driver_inv304 net[304] wl[304] vdd gnd pinv_11
Xwl_driver_inv_en305 en en_bar[305] vdd gnd pinv_12
Xwl_driver_nand305 en_bar[305] in[305] net[305] vdd gnd pnand2_4
Xwl_driver_inv305 net[305] wl[305] vdd gnd pinv_11
Xwl_driver_inv_en306 en en_bar[306] vdd gnd pinv_12
Xwl_driver_nand306 en_bar[306] in[306] net[306] vdd gnd pnand2_4
Xwl_driver_inv306 net[306] wl[306] vdd gnd pinv_11
Xwl_driver_inv_en307 en en_bar[307] vdd gnd pinv_12
Xwl_driver_nand307 en_bar[307] in[307] net[307] vdd gnd pnand2_4
Xwl_driver_inv307 net[307] wl[307] vdd gnd pinv_11
Xwl_driver_inv_en308 en en_bar[308] vdd gnd pinv_12
Xwl_driver_nand308 en_bar[308] in[308] net[308] vdd gnd pnand2_4
Xwl_driver_inv308 net[308] wl[308] vdd gnd pinv_11
Xwl_driver_inv_en309 en en_bar[309] vdd gnd pinv_12
Xwl_driver_nand309 en_bar[309] in[309] net[309] vdd gnd pnand2_4
Xwl_driver_inv309 net[309] wl[309] vdd gnd pinv_11
Xwl_driver_inv_en310 en en_bar[310] vdd gnd pinv_12
Xwl_driver_nand310 en_bar[310] in[310] net[310] vdd gnd pnand2_4
Xwl_driver_inv310 net[310] wl[310] vdd gnd pinv_11
Xwl_driver_inv_en311 en en_bar[311] vdd gnd pinv_12
Xwl_driver_nand311 en_bar[311] in[311] net[311] vdd gnd pnand2_4
Xwl_driver_inv311 net[311] wl[311] vdd gnd pinv_11
Xwl_driver_inv_en312 en en_bar[312] vdd gnd pinv_12
Xwl_driver_nand312 en_bar[312] in[312] net[312] vdd gnd pnand2_4
Xwl_driver_inv312 net[312] wl[312] vdd gnd pinv_11
Xwl_driver_inv_en313 en en_bar[313] vdd gnd pinv_12
Xwl_driver_nand313 en_bar[313] in[313] net[313] vdd gnd pnand2_4
Xwl_driver_inv313 net[313] wl[313] vdd gnd pinv_11
Xwl_driver_inv_en314 en en_bar[314] vdd gnd pinv_12
Xwl_driver_nand314 en_bar[314] in[314] net[314] vdd gnd pnand2_4
Xwl_driver_inv314 net[314] wl[314] vdd gnd pinv_11
Xwl_driver_inv_en315 en en_bar[315] vdd gnd pinv_12
Xwl_driver_nand315 en_bar[315] in[315] net[315] vdd gnd pnand2_4
Xwl_driver_inv315 net[315] wl[315] vdd gnd pinv_11
Xwl_driver_inv_en316 en en_bar[316] vdd gnd pinv_12
Xwl_driver_nand316 en_bar[316] in[316] net[316] vdd gnd pnand2_4
Xwl_driver_inv316 net[316] wl[316] vdd gnd pinv_11
Xwl_driver_inv_en317 en en_bar[317] vdd gnd pinv_12
Xwl_driver_nand317 en_bar[317] in[317] net[317] vdd gnd pnand2_4
Xwl_driver_inv317 net[317] wl[317] vdd gnd pinv_11
Xwl_driver_inv_en318 en en_bar[318] vdd gnd pinv_12
Xwl_driver_nand318 en_bar[318] in[318] net[318] vdd gnd pnand2_4
Xwl_driver_inv318 net[318] wl[318] vdd gnd pinv_11
Xwl_driver_inv_en319 en en_bar[319] vdd gnd pinv_12
Xwl_driver_nand319 en_bar[319] in[319] net[319] vdd gnd pnand2_4
Xwl_driver_inv319 net[319] wl[319] vdd gnd pinv_11
Xwl_driver_inv_en320 en en_bar[320] vdd gnd pinv_12
Xwl_driver_nand320 en_bar[320] in[320] net[320] vdd gnd pnand2_4
Xwl_driver_inv320 net[320] wl[320] vdd gnd pinv_11
Xwl_driver_inv_en321 en en_bar[321] vdd gnd pinv_12
Xwl_driver_nand321 en_bar[321] in[321] net[321] vdd gnd pnand2_4
Xwl_driver_inv321 net[321] wl[321] vdd gnd pinv_11
Xwl_driver_inv_en322 en en_bar[322] vdd gnd pinv_12
Xwl_driver_nand322 en_bar[322] in[322] net[322] vdd gnd pnand2_4
Xwl_driver_inv322 net[322] wl[322] vdd gnd pinv_11
Xwl_driver_inv_en323 en en_bar[323] vdd gnd pinv_12
Xwl_driver_nand323 en_bar[323] in[323] net[323] vdd gnd pnand2_4
Xwl_driver_inv323 net[323] wl[323] vdd gnd pinv_11
Xwl_driver_inv_en324 en en_bar[324] vdd gnd pinv_12
Xwl_driver_nand324 en_bar[324] in[324] net[324] vdd gnd pnand2_4
Xwl_driver_inv324 net[324] wl[324] vdd gnd pinv_11
Xwl_driver_inv_en325 en en_bar[325] vdd gnd pinv_12
Xwl_driver_nand325 en_bar[325] in[325] net[325] vdd gnd pnand2_4
Xwl_driver_inv325 net[325] wl[325] vdd gnd pinv_11
Xwl_driver_inv_en326 en en_bar[326] vdd gnd pinv_12
Xwl_driver_nand326 en_bar[326] in[326] net[326] vdd gnd pnand2_4
Xwl_driver_inv326 net[326] wl[326] vdd gnd pinv_11
Xwl_driver_inv_en327 en en_bar[327] vdd gnd pinv_12
Xwl_driver_nand327 en_bar[327] in[327] net[327] vdd gnd pnand2_4
Xwl_driver_inv327 net[327] wl[327] vdd gnd pinv_11
Xwl_driver_inv_en328 en en_bar[328] vdd gnd pinv_12
Xwl_driver_nand328 en_bar[328] in[328] net[328] vdd gnd pnand2_4
Xwl_driver_inv328 net[328] wl[328] vdd gnd pinv_11
Xwl_driver_inv_en329 en en_bar[329] vdd gnd pinv_12
Xwl_driver_nand329 en_bar[329] in[329] net[329] vdd gnd pnand2_4
Xwl_driver_inv329 net[329] wl[329] vdd gnd pinv_11
Xwl_driver_inv_en330 en en_bar[330] vdd gnd pinv_12
Xwl_driver_nand330 en_bar[330] in[330] net[330] vdd gnd pnand2_4
Xwl_driver_inv330 net[330] wl[330] vdd gnd pinv_11
Xwl_driver_inv_en331 en en_bar[331] vdd gnd pinv_12
Xwl_driver_nand331 en_bar[331] in[331] net[331] vdd gnd pnand2_4
Xwl_driver_inv331 net[331] wl[331] vdd gnd pinv_11
Xwl_driver_inv_en332 en en_bar[332] vdd gnd pinv_12
Xwl_driver_nand332 en_bar[332] in[332] net[332] vdd gnd pnand2_4
Xwl_driver_inv332 net[332] wl[332] vdd gnd pinv_11
Xwl_driver_inv_en333 en en_bar[333] vdd gnd pinv_12
Xwl_driver_nand333 en_bar[333] in[333] net[333] vdd gnd pnand2_4
Xwl_driver_inv333 net[333] wl[333] vdd gnd pinv_11
Xwl_driver_inv_en334 en en_bar[334] vdd gnd pinv_12
Xwl_driver_nand334 en_bar[334] in[334] net[334] vdd gnd pnand2_4
Xwl_driver_inv334 net[334] wl[334] vdd gnd pinv_11
Xwl_driver_inv_en335 en en_bar[335] vdd gnd pinv_12
Xwl_driver_nand335 en_bar[335] in[335] net[335] vdd gnd pnand2_4
Xwl_driver_inv335 net[335] wl[335] vdd gnd pinv_11
Xwl_driver_inv_en336 en en_bar[336] vdd gnd pinv_12
Xwl_driver_nand336 en_bar[336] in[336] net[336] vdd gnd pnand2_4
Xwl_driver_inv336 net[336] wl[336] vdd gnd pinv_11
Xwl_driver_inv_en337 en en_bar[337] vdd gnd pinv_12
Xwl_driver_nand337 en_bar[337] in[337] net[337] vdd gnd pnand2_4
Xwl_driver_inv337 net[337] wl[337] vdd gnd pinv_11
Xwl_driver_inv_en338 en en_bar[338] vdd gnd pinv_12
Xwl_driver_nand338 en_bar[338] in[338] net[338] vdd gnd pnand2_4
Xwl_driver_inv338 net[338] wl[338] vdd gnd pinv_11
Xwl_driver_inv_en339 en en_bar[339] vdd gnd pinv_12
Xwl_driver_nand339 en_bar[339] in[339] net[339] vdd gnd pnand2_4
Xwl_driver_inv339 net[339] wl[339] vdd gnd pinv_11
Xwl_driver_inv_en340 en en_bar[340] vdd gnd pinv_12
Xwl_driver_nand340 en_bar[340] in[340] net[340] vdd gnd pnand2_4
Xwl_driver_inv340 net[340] wl[340] vdd gnd pinv_11
Xwl_driver_inv_en341 en en_bar[341] vdd gnd pinv_12
Xwl_driver_nand341 en_bar[341] in[341] net[341] vdd gnd pnand2_4
Xwl_driver_inv341 net[341] wl[341] vdd gnd pinv_11
Xwl_driver_inv_en342 en en_bar[342] vdd gnd pinv_12
Xwl_driver_nand342 en_bar[342] in[342] net[342] vdd gnd pnand2_4
Xwl_driver_inv342 net[342] wl[342] vdd gnd pinv_11
Xwl_driver_inv_en343 en en_bar[343] vdd gnd pinv_12
Xwl_driver_nand343 en_bar[343] in[343] net[343] vdd gnd pnand2_4
Xwl_driver_inv343 net[343] wl[343] vdd gnd pinv_11
Xwl_driver_inv_en344 en en_bar[344] vdd gnd pinv_12
Xwl_driver_nand344 en_bar[344] in[344] net[344] vdd gnd pnand2_4
Xwl_driver_inv344 net[344] wl[344] vdd gnd pinv_11
Xwl_driver_inv_en345 en en_bar[345] vdd gnd pinv_12
Xwl_driver_nand345 en_bar[345] in[345] net[345] vdd gnd pnand2_4
Xwl_driver_inv345 net[345] wl[345] vdd gnd pinv_11
Xwl_driver_inv_en346 en en_bar[346] vdd gnd pinv_12
Xwl_driver_nand346 en_bar[346] in[346] net[346] vdd gnd pnand2_4
Xwl_driver_inv346 net[346] wl[346] vdd gnd pinv_11
Xwl_driver_inv_en347 en en_bar[347] vdd gnd pinv_12
Xwl_driver_nand347 en_bar[347] in[347] net[347] vdd gnd pnand2_4
Xwl_driver_inv347 net[347] wl[347] vdd gnd pinv_11
Xwl_driver_inv_en348 en en_bar[348] vdd gnd pinv_12
Xwl_driver_nand348 en_bar[348] in[348] net[348] vdd gnd pnand2_4
Xwl_driver_inv348 net[348] wl[348] vdd gnd pinv_11
Xwl_driver_inv_en349 en en_bar[349] vdd gnd pinv_12
Xwl_driver_nand349 en_bar[349] in[349] net[349] vdd gnd pnand2_4
Xwl_driver_inv349 net[349] wl[349] vdd gnd pinv_11
Xwl_driver_inv_en350 en en_bar[350] vdd gnd pinv_12
Xwl_driver_nand350 en_bar[350] in[350] net[350] vdd gnd pnand2_4
Xwl_driver_inv350 net[350] wl[350] vdd gnd pinv_11
Xwl_driver_inv_en351 en en_bar[351] vdd gnd pinv_12
Xwl_driver_nand351 en_bar[351] in[351] net[351] vdd gnd pnand2_4
Xwl_driver_inv351 net[351] wl[351] vdd gnd pinv_11
Xwl_driver_inv_en352 en en_bar[352] vdd gnd pinv_12
Xwl_driver_nand352 en_bar[352] in[352] net[352] vdd gnd pnand2_4
Xwl_driver_inv352 net[352] wl[352] vdd gnd pinv_11
Xwl_driver_inv_en353 en en_bar[353] vdd gnd pinv_12
Xwl_driver_nand353 en_bar[353] in[353] net[353] vdd gnd pnand2_4
Xwl_driver_inv353 net[353] wl[353] vdd gnd pinv_11
Xwl_driver_inv_en354 en en_bar[354] vdd gnd pinv_12
Xwl_driver_nand354 en_bar[354] in[354] net[354] vdd gnd pnand2_4
Xwl_driver_inv354 net[354] wl[354] vdd gnd pinv_11
Xwl_driver_inv_en355 en en_bar[355] vdd gnd pinv_12
Xwl_driver_nand355 en_bar[355] in[355] net[355] vdd gnd pnand2_4
Xwl_driver_inv355 net[355] wl[355] vdd gnd pinv_11
Xwl_driver_inv_en356 en en_bar[356] vdd gnd pinv_12
Xwl_driver_nand356 en_bar[356] in[356] net[356] vdd gnd pnand2_4
Xwl_driver_inv356 net[356] wl[356] vdd gnd pinv_11
Xwl_driver_inv_en357 en en_bar[357] vdd gnd pinv_12
Xwl_driver_nand357 en_bar[357] in[357] net[357] vdd gnd pnand2_4
Xwl_driver_inv357 net[357] wl[357] vdd gnd pinv_11
Xwl_driver_inv_en358 en en_bar[358] vdd gnd pinv_12
Xwl_driver_nand358 en_bar[358] in[358] net[358] vdd gnd pnand2_4
Xwl_driver_inv358 net[358] wl[358] vdd gnd pinv_11
Xwl_driver_inv_en359 en en_bar[359] vdd gnd pinv_12
Xwl_driver_nand359 en_bar[359] in[359] net[359] vdd gnd pnand2_4
Xwl_driver_inv359 net[359] wl[359] vdd gnd pinv_11
Xwl_driver_inv_en360 en en_bar[360] vdd gnd pinv_12
Xwl_driver_nand360 en_bar[360] in[360] net[360] vdd gnd pnand2_4
Xwl_driver_inv360 net[360] wl[360] vdd gnd pinv_11
Xwl_driver_inv_en361 en en_bar[361] vdd gnd pinv_12
Xwl_driver_nand361 en_bar[361] in[361] net[361] vdd gnd pnand2_4
Xwl_driver_inv361 net[361] wl[361] vdd gnd pinv_11
Xwl_driver_inv_en362 en en_bar[362] vdd gnd pinv_12
Xwl_driver_nand362 en_bar[362] in[362] net[362] vdd gnd pnand2_4
Xwl_driver_inv362 net[362] wl[362] vdd gnd pinv_11
Xwl_driver_inv_en363 en en_bar[363] vdd gnd pinv_12
Xwl_driver_nand363 en_bar[363] in[363] net[363] vdd gnd pnand2_4
Xwl_driver_inv363 net[363] wl[363] vdd gnd pinv_11
Xwl_driver_inv_en364 en en_bar[364] vdd gnd pinv_12
Xwl_driver_nand364 en_bar[364] in[364] net[364] vdd gnd pnand2_4
Xwl_driver_inv364 net[364] wl[364] vdd gnd pinv_11
Xwl_driver_inv_en365 en en_bar[365] vdd gnd pinv_12
Xwl_driver_nand365 en_bar[365] in[365] net[365] vdd gnd pnand2_4
Xwl_driver_inv365 net[365] wl[365] vdd gnd pinv_11
Xwl_driver_inv_en366 en en_bar[366] vdd gnd pinv_12
Xwl_driver_nand366 en_bar[366] in[366] net[366] vdd gnd pnand2_4
Xwl_driver_inv366 net[366] wl[366] vdd gnd pinv_11
Xwl_driver_inv_en367 en en_bar[367] vdd gnd pinv_12
Xwl_driver_nand367 en_bar[367] in[367] net[367] vdd gnd pnand2_4
Xwl_driver_inv367 net[367] wl[367] vdd gnd pinv_11
Xwl_driver_inv_en368 en en_bar[368] vdd gnd pinv_12
Xwl_driver_nand368 en_bar[368] in[368] net[368] vdd gnd pnand2_4
Xwl_driver_inv368 net[368] wl[368] vdd gnd pinv_11
Xwl_driver_inv_en369 en en_bar[369] vdd gnd pinv_12
Xwl_driver_nand369 en_bar[369] in[369] net[369] vdd gnd pnand2_4
Xwl_driver_inv369 net[369] wl[369] vdd gnd pinv_11
Xwl_driver_inv_en370 en en_bar[370] vdd gnd pinv_12
Xwl_driver_nand370 en_bar[370] in[370] net[370] vdd gnd pnand2_4
Xwl_driver_inv370 net[370] wl[370] vdd gnd pinv_11
Xwl_driver_inv_en371 en en_bar[371] vdd gnd pinv_12
Xwl_driver_nand371 en_bar[371] in[371] net[371] vdd gnd pnand2_4
Xwl_driver_inv371 net[371] wl[371] vdd gnd pinv_11
Xwl_driver_inv_en372 en en_bar[372] vdd gnd pinv_12
Xwl_driver_nand372 en_bar[372] in[372] net[372] vdd gnd pnand2_4
Xwl_driver_inv372 net[372] wl[372] vdd gnd pinv_11
Xwl_driver_inv_en373 en en_bar[373] vdd gnd pinv_12
Xwl_driver_nand373 en_bar[373] in[373] net[373] vdd gnd pnand2_4
Xwl_driver_inv373 net[373] wl[373] vdd gnd pinv_11
Xwl_driver_inv_en374 en en_bar[374] vdd gnd pinv_12
Xwl_driver_nand374 en_bar[374] in[374] net[374] vdd gnd pnand2_4
Xwl_driver_inv374 net[374] wl[374] vdd gnd pinv_11
Xwl_driver_inv_en375 en en_bar[375] vdd gnd pinv_12
Xwl_driver_nand375 en_bar[375] in[375] net[375] vdd gnd pnand2_4
Xwl_driver_inv375 net[375] wl[375] vdd gnd pinv_11
Xwl_driver_inv_en376 en en_bar[376] vdd gnd pinv_12
Xwl_driver_nand376 en_bar[376] in[376] net[376] vdd gnd pnand2_4
Xwl_driver_inv376 net[376] wl[376] vdd gnd pinv_11
Xwl_driver_inv_en377 en en_bar[377] vdd gnd pinv_12
Xwl_driver_nand377 en_bar[377] in[377] net[377] vdd gnd pnand2_4
Xwl_driver_inv377 net[377] wl[377] vdd gnd pinv_11
Xwl_driver_inv_en378 en en_bar[378] vdd gnd pinv_12
Xwl_driver_nand378 en_bar[378] in[378] net[378] vdd gnd pnand2_4
Xwl_driver_inv378 net[378] wl[378] vdd gnd pinv_11
Xwl_driver_inv_en379 en en_bar[379] vdd gnd pinv_12
Xwl_driver_nand379 en_bar[379] in[379] net[379] vdd gnd pnand2_4
Xwl_driver_inv379 net[379] wl[379] vdd gnd pinv_11
Xwl_driver_inv_en380 en en_bar[380] vdd gnd pinv_12
Xwl_driver_nand380 en_bar[380] in[380] net[380] vdd gnd pnand2_4
Xwl_driver_inv380 net[380] wl[380] vdd gnd pinv_11
Xwl_driver_inv_en381 en en_bar[381] vdd gnd pinv_12
Xwl_driver_nand381 en_bar[381] in[381] net[381] vdd gnd pnand2_4
Xwl_driver_inv381 net[381] wl[381] vdd gnd pinv_11
Xwl_driver_inv_en382 en en_bar[382] vdd gnd pinv_12
Xwl_driver_nand382 en_bar[382] in[382] net[382] vdd gnd pnand2_4
Xwl_driver_inv382 net[382] wl[382] vdd gnd pinv_11
Xwl_driver_inv_en383 en en_bar[383] vdd gnd pinv_12
Xwl_driver_nand383 en_bar[383] in[383] net[383] vdd gnd pnand2_4
Xwl_driver_inv383 net[383] wl[383] vdd gnd pinv_11
Xwl_driver_inv_en384 en en_bar[384] vdd gnd pinv_12
Xwl_driver_nand384 en_bar[384] in[384] net[384] vdd gnd pnand2_4
Xwl_driver_inv384 net[384] wl[384] vdd gnd pinv_11
Xwl_driver_inv_en385 en en_bar[385] vdd gnd pinv_12
Xwl_driver_nand385 en_bar[385] in[385] net[385] vdd gnd pnand2_4
Xwl_driver_inv385 net[385] wl[385] vdd gnd pinv_11
Xwl_driver_inv_en386 en en_bar[386] vdd gnd pinv_12
Xwl_driver_nand386 en_bar[386] in[386] net[386] vdd gnd pnand2_4
Xwl_driver_inv386 net[386] wl[386] vdd gnd pinv_11
Xwl_driver_inv_en387 en en_bar[387] vdd gnd pinv_12
Xwl_driver_nand387 en_bar[387] in[387] net[387] vdd gnd pnand2_4
Xwl_driver_inv387 net[387] wl[387] vdd gnd pinv_11
Xwl_driver_inv_en388 en en_bar[388] vdd gnd pinv_12
Xwl_driver_nand388 en_bar[388] in[388] net[388] vdd gnd pnand2_4
Xwl_driver_inv388 net[388] wl[388] vdd gnd pinv_11
Xwl_driver_inv_en389 en en_bar[389] vdd gnd pinv_12
Xwl_driver_nand389 en_bar[389] in[389] net[389] vdd gnd pnand2_4
Xwl_driver_inv389 net[389] wl[389] vdd gnd pinv_11
Xwl_driver_inv_en390 en en_bar[390] vdd gnd pinv_12
Xwl_driver_nand390 en_bar[390] in[390] net[390] vdd gnd pnand2_4
Xwl_driver_inv390 net[390] wl[390] vdd gnd pinv_11
Xwl_driver_inv_en391 en en_bar[391] vdd gnd pinv_12
Xwl_driver_nand391 en_bar[391] in[391] net[391] vdd gnd pnand2_4
Xwl_driver_inv391 net[391] wl[391] vdd gnd pinv_11
Xwl_driver_inv_en392 en en_bar[392] vdd gnd pinv_12
Xwl_driver_nand392 en_bar[392] in[392] net[392] vdd gnd pnand2_4
Xwl_driver_inv392 net[392] wl[392] vdd gnd pinv_11
Xwl_driver_inv_en393 en en_bar[393] vdd gnd pinv_12
Xwl_driver_nand393 en_bar[393] in[393] net[393] vdd gnd pnand2_4
Xwl_driver_inv393 net[393] wl[393] vdd gnd pinv_11
Xwl_driver_inv_en394 en en_bar[394] vdd gnd pinv_12
Xwl_driver_nand394 en_bar[394] in[394] net[394] vdd gnd pnand2_4
Xwl_driver_inv394 net[394] wl[394] vdd gnd pinv_11
Xwl_driver_inv_en395 en en_bar[395] vdd gnd pinv_12
Xwl_driver_nand395 en_bar[395] in[395] net[395] vdd gnd pnand2_4
Xwl_driver_inv395 net[395] wl[395] vdd gnd pinv_11
Xwl_driver_inv_en396 en en_bar[396] vdd gnd pinv_12
Xwl_driver_nand396 en_bar[396] in[396] net[396] vdd gnd pnand2_4
Xwl_driver_inv396 net[396] wl[396] vdd gnd pinv_11
Xwl_driver_inv_en397 en en_bar[397] vdd gnd pinv_12
Xwl_driver_nand397 en_bar[397] in[397] net[397] vdd gnd pnand2_4
Xwl_driver_inv397 net[397] wl[397] vdd gnd pinv_11
Xwl_driver_inv_en398 en en_bar[398] vdd gnd pinv_12
Xwl_driver_nand398 en_bar[398] in[398] net[398] vdd gnd pnand2_4
Xwl_driver_inv398 net[398] wl[398] vdd gnd pinv_11
Xwl_driver_inv_en399 en en_bar[399] vdd gnd pinv_12
Xwl_driver_nand399 en_bar[399] in[399] net[399] vdd gnd pnand2_4
Xwl_driver_inv399 net[399] wl[399] vdd gnd pinv_11
Xwl_driver_inv_en400 en en_bar[400] vdd gnd pinv_12
Xwl_driver_nand400 en_bar[400] in[400] net[400] vdd gnd pnand2_4
Xwl_driver_inv400 net[400] wl[400] vdd gnd pinv_11
Xwl_driver_inv_en401 en en_bar[401] vdd gnd pinv_12
Xwl_driver_nand401 en_bar[401] in[401] net[401] vdd gnd pnand2_4
Xwl_driver_inv401 net[401] wl[401] vdd gnd pinv_11
Xwl_driver_inv_en402 en en_bar[402] vdd gnd pinv_12
Xwl_driver_nand402 en_bar[402] in[402] net[402] vdd gnd pnand2_4
Xwl_driver_inv402 net[402] wl[402] vdd gnd pinv_11
Xwl_driver_inv_en403 en en_bar[403] vdd gnd pinv_12
Xwl_driver_nand403 en_bar[403] in[403] net[403] vdd gnd pnand2_4
Xwl_driver_inv403 net[403] wl[403] vdd gnd pinv_11
Xwl_driver_inv_en404 en en_bar[404] vdd gnd pinv_12
Xwl_driver_nand404 en_bar[404] in[404] net[404] vdd gnd pnand2_4
Xwl_driver_inv404 net[404] wl[404] vdd gnd pinv_11
Xwl_driver_inv_en405 en en_bar[405] vdd gnd pinv_12
Xwl_driver_nand405 en_bar[405] in[405] net[405] vdd gnd pnand2_4
Xwl_driver_inv405 net[405] wl[405] vdd gnd pinv_11
Xwl_driver_inv_en406 en en_bar[406] vdd gnd pinv_12
Xwl_driver_nand406 en_bar[406] in[406] net[406] vdd gnd pnand2_4
Xwl_driver_inv406 net[406] wl[406] vdd gnd pinv_11
Xwl_driver_inv_en407 en en_bar[407] vdd gnd pinv_12
Xwl_driver_nand407 en_bar[407] in[407] net[407] vdd gnd pnand2_4
Xwl_driver_inv407 net[407] wl[407] vdd gnd pinv_11
Xwl_driver_inv_en408 en en_bar[408] vdd gnd pinv_12
Xwl_driver_nand408 en_bar[408] in[408] net[408] vdd gnd pnand2_4
Xwl_driver_inv408 net[408] wl[408] vdd gnd pinv_11
Xwl_driver_inv_en409 en en_bar[409] vdd gnd pinv_12
Xwl_driver_nand409 en_bar[409] in[409] net[409] vdd gnd pnand2_4
Xwl_driver_inv409 net[409] wl[409] vdd gnd pinv_11
Xwl_driver_inv_en410 en en_bar[410] vdd gnd pinv_12
Xwl_driver_nand410 en_bar[410] in[410] net[410] vdd gnd pnand2_4
Xwl_driver_inv410 net[410] wl[410] vdd gnd pinv_11
Xwl_driver_inv_en411 en en_bar[411] vdd gnd pinv_12
Xwl_driver_nand411 en_bar[411] in[411] net[411] vdd gnd pnand2_4
Xwl_driver_inv411 net[411] wl[411] vdd gnd pinv_11
Xwl_driver_inv_en412 en en_bar[412] vdd gnd pinv_12
Xwl_driver_nand412 en_bar[412] in[412] net[412] vdd gnd pnand2_4
Xwl_driver_inv412 net[412] wl[412] vdd gnd pinv_11
Xwl_driver_inv_en413 en en_bar[413] vdd gnd pinv_12
Xwl_driver_nand413 en_bar[413] in[413] net[413] vdd gnd pnand2_4
Xwl_driver_inv413 net[413] wl[413] vdd gnd pinv_11
Xwl_driver_inv_en414 en en_bar[414] vdd gnd pinv_12
Xwl_driver_nand414 en_bar[414] in[414] net[414] vdd gnd pnand2_4
Xwl_driver_inv414 net[414] wl[414] vdd gnd pinv_11
Xwl_driver_inv_en415 en en_bar[415] vdd gnd pinv_12
Xwl_driver_nand415 en_bar[415] in[415] net[415] vdd gnd pnand2_4
Xwl_driver_inv415 net[415] wl[415] vdd gnd pinv_11
Xwl_driver_inv_en416 en en_bar[416] vdd gnd pinv_12
Xwl_driver_nand416 en_bar[416] in[416] net[416] vdd gnd pnand2_4
Xwl_driver_inv416 net[416] wl[416] vdd gnd pinv_11
Xwl_driver_inv_en417 en en_bar[417] vdd gnd pinv_12
Xwl_driver_nand417 en_bar[417] in[417] net[417] vdd gnd pnand2_4
Xwl_driver_inv417 net[417] wl[417] vdd gnd pinv_11
Xwl_driver_inv_en418 en en_bar[418] vdd gnd pinv_12
Xwl_driver_nand418 en_bar[418] in[418] net[418] vdd gnd pnand2_4
Xwl_driver_inv418 net[418] wl[418] vdd gnd pinv_11
Xwl_driver_inv_en419 en en_bar[419] vdd gnd pinv_12
Xwl_driver_nand419 en_bar[419] in[419] net[419] vdd gnd pnand2_4
Xwl_driver_inv419 net[419] wl[419] vdd gnd pinv_11
Xwl_driver_inv_en420 en en_bar[420] vdd gnd pinv_12
Xwl_driver_nand420 en_bar[420] in[420] net[420] vdd gnd pnand2_4
Xwl_driver_inv420 net[420] wl[420] vdd gnd pinv_11
Xwl_driver_inv_en421 en en_bar[421] vdd gnd pinv_12
Xwl_driver_nand421 en_bar[421] in[421] net[421] vdd gnd pnand2_4
Xwl_driver_inv421 net[421] wl[421] vdd gnd pinv_11
Xwl_driver_inv_en422 en en_bar[422] vdd gnd pinv_12
Xwl_driver_nand422 en_bar[422] in[422] net[422] vdd gnd pnand2_4
Xwl_driver_inv422 net[422] wl[422] vdd gnd pinv_11
Xwl_driver_inv_en423 en en_bar[423] vdd gnd pinv_12
Xwl_driver_nand423 en_bar[423] in[423] net[423] vdd gnd pnand2_4
Xwl_driver_inv423 net[423] wl[423] vdd gnd pinv_11
Xwl_driver_inv_en424 en en_bar[424] vdd gnd pinv_12
Xwl_driver_nand424 en_bar[424] in[424] net[424] vdd gnd pnand2_4
Xwl_driver_inv424 net[424] wl[424] vdd gnd pinv_11
Xwl_driver_inv_en425 en en_bar[425] vdd gnd pinv_12
Xwl_driver_nand425 en_bar[425] in[425] net[425] vdd gnd pnand2_4
Xwl_driver_inv425 net[425] wl[425] vdd gnd pinv_11
Xwl_driver_inv_en426 en en_bar[426] vdd gnd pinv_12
Xwl_driver_nand426 en_bar[426] in[426] net[426] vdd gnd pnand2_4
Xwl_driver_inv426 net[426] wl[426] vdd gnd pinv_11
Xwl_driver_inv_en427 en en_bar[427] vdd gnd pinv_12
Xwl_driver_nand427 en_bar[427] in[427] net[427] vdd gnd pnand2_4
Xwl_driver_inv427 net[427] wl[427] vdd gnd pinv_11
Xwl_driver_inv_en428 en en_bar[428] vdd gnd pinv_12
Xwl_driver_nand428 en_bar[428] in[428] net[428] vdd gnd pnand2_4
Xwl_driver_inv428 net[428] wl[428] vdd gnd pinv_11
Xwl_driver_inv_en429 en en_bar[429] vdd gnd pinv_12
Xwl_driver_nand429 en_bar[429] in[429] net[429] vdd gnd pnand2_4
Xwl_driver_inv429 net[429] wl[429] vdd gnd pinv_11
Xwl_driver_inv_en430 en en_bar[430] vdd gnd pinv_12
Xwl_driver_nand430 en_bar[430] in[430] net[430] vdd gnd pnand2_4
Xwl_driver_inv430 net[430] wl[430] vdd gnd pinv_11
Xwl_driver_inv_en431 en en_bar[431] vdd gnd pinv_12
Xwl_driver_nand431 en_bar[431] in[431] net[431] vdd gnd pnand2_4
Xwl_driver_inv431 net[431] wl[431] vdd gnd pinv_11
Xwl_driver_inv_en432 en en_bar[432] vdd gnd pinv_12
Xwl_driver_nand432 en_bar[432] in[432] net[432] vdd gnd pnand2_4
Xwl_driver_inv432 net[432] wl[432] vdd gnd pinv_11
Xwl_driver_inv_en433 en en_bar[433] vdd gnd pinv_12
Xwl_driver_nand433 en_bar[433] in[433] net[433] vdd gnd pnand2_4
Xwl_driver_inv433 net[433] wl[433] vdd gnd pinv_11
Xwl_driver_inv_en434 en en_bar[434] vdd gnd pinv_12
Xwl_driver_nand434 en_bar[434] in[434] net[434] vdd gnd pnand2_4
Xwl_driver_inv434 net[434] wl[434] vdd gnd pinv_11
Xwl_driver_inv_en435 en en_bar[435] vdd gnd pinv_12
Xwl_driver_nand435 en_bar[435] in[435] net[435] vdd gnd pnand2_4
Xwl_driver_inv435 net[435] wl[435] vdd gnd pinv_11
Xwl_driver_inv_en436 en en_bar[436] vdd gnd pinv_12
Xwl_driver_nand436 en_bar[436] in[436] net[436] vdd gnd pnand2_4
Xwl_driver_inv436 net[436] wl[436] vdd gnd pinv_11
Xwl_driver_inv_en437 en en_bar[437] vdd gnd pinv_12
Xwl_driver_nand437 en_bar[437] in[437] net[437] vdd gnd pnand2_4
Xwl_driver_inv437 net[437] wl[437] vdd gnd pinv_11
Xwl_driver_inv_en438 en en_bar[438] vdd gnd pinv_12
Xwl_driver_nand438 en_bar[438] in[438] net[438] vdd gnd pnand2_4
Xwl_driver_inv438 net[438] wl[438] vdd gnd pinv_11
Xwl_driver_inv_en439 en en_bar[439] vdd gnd pinv_12
Xwl_driver_nand439 en_bar[439] in[439] net[439] vdd gnd pnand2_4
Xwl_driver_inv439 net[439] wl[439] vdd gnd pinv_11
Xwl_driver_inv_en440 en en_bar[440] vdd gnd pinv_12
Xwl_driver_nand440 en_bar[440] in[440] net[440] vdd gnd pnand2_4
Xwl_driver_inv440 net[440] wl[440] vdd gnd pinv_11
Xwl_driver_inv_en441 en en_bar[441] vdd gnd pinv_12
Xwl_driver_nand441 en_bar[441] in[441] net[441] vdd gnd pnand2_4
Xwl_driver_inv441 net[441] wl[441] vdd gnd pinv_11
Xwl_driver_inv_en442 en en_bar[442] vdd gnd pinv_12
Xwl_driver_nand442 en_bar[442] in[442] net[442] vdd gnd pnand2_4
Xwl_driver_inv442 net[442] wl[442] vdd gnd pinv_11
Xwl_driver_inv_en443 en en_bar[443] vdd gnd pinv_12
Xwl_driver_nand443 en_bar[443] in[443] net[443] vdd gnd pnand2_4
Xwl_driver_inv443 net[443] wl[443] vdd gnd pinv_11
Xwl_driver_inv_en444 en en_bar[444] vdd gnd pinv_12
Xwl_driver_nand444 en_bar[444] in[444] net[444] vdd gnd pnand2_4
Xwl_driver_inv444 net[444] wl[444] vdd gnd pinv_11
Xwl_driver_inv_en445 en en_bar[445] vdd gnd pinv_12
Xwl_driver_nand445 en_bar[445] in[445] net[445] vdd gnd pnand2_4
Xwl_driver_inv445 net[445] wl[445] vdd gnd pinv_11
Xwl_driver_inv_en446 en en_bar[446] vdd gnd pinv_12
Xwl_driver_nand446 en_bar[446] in[446] net[446] vdd gnd pnand2_4
Xwl_driver_inv446 net[446] wl[446] vdd gnd pinv_11
Xwl_driver_inv_en447 en en_bar[447] vdd gnd pinv_12
Xwl_driver_nand447 en_bar[447] in[447] net[447] vdd gnd pnand2_4
Xwl_driver_inv447 net[447] wl[447] vdd gnd pinv_11
Xwl_driver_inv_en448 en en_bar[448] vdd gnd pinv_12
Xwl_driver_nand448 en_bar[448] in[448] net[448] vdd gnd pnand2_4
Xwl_driver_inv448 net[448] wl[448] vdd gnd pinv_11
Xwl_driver_inv_en449 en en_bar[449] vdd gnd pinv_12
Xwl_driver_nand449 en_bar[449] in[449] net[449] vdd gnd pnand2_4
Xwl_driver_inv449 net[449] wl[449] vdd gnd pinv_11
Xwl_driver_inv_en450 en en_bar[450] vdd gnd pinv_12
Xwl_driver_nand450 en_bar[450] in[450] net[450] vdd gnd pnand2_4
Xwl_driver_inv450 net[450] wl[450] vdd gnd pinv_11
Xwl_driver_inv_en451 en en_bar[451] vdd gnd pinv_12
Xwl_driver_nand451 en_bar[451] in[451] net[451] vdd gnd pnand2_4
Xwl_driver_inv451 net[451] wl[451] vdd gnd pinv_11
Xwl_driver_inv_en452 en en_bar[452] vdd gnd pinv_12
Xwl_driver_nand452 en_bar[452] in[452] net[452] vdd gnd pnand2_4
Xwl_driver_inv452 net[452] wl[452] vdd gnd pinv_11
Xwl_driver_inv_en453 en en_bar[453] vdd gnd pinv_12
Xwl_driver_nand453 en_bar[453] in[453] net[453] vdd gnd pnand2_4
Xwl_driver_inv453 net[453] wl[453] vdd gnd pinv_11
Xwl_driver_inv_en454 en en_bar[454] vdd gnd pinv_12
Xwl_driver_nand454 en_bar[454] in[454] net[454] vdd gnd pnand2_4
Xwl_driver_inv454 net[454] wl[454] vdd gnd pinv_11
Xwl_driver_inv_en455 en en_bar[455] vdd gnd pinv_12
Xwl_driver_nand455 en_bar[455] in[455] net[455] vdd gnd pnand2_4
Xwl_driver_inv455 net[455] wl[455] vdd gnd pinv_11
Xwl_driver_inv_en456 en en_bar[456] vdd gnd pinv_12
Xwl_driver_nand456 en_bar[456] in[456] net[456] vdd gnd pnand2_4
Xwl_driver_inv456 net[456] wl[456] vdd gnd pinv_11
Xwl_driver_inv_en457 en en_bar[457] vdd gnd pinv_12
Xwl_driver_nand457 en_bar[457] in[457] net[457] vdd gnd pnand2_4
Xwl_driver_inv457 net[457] wl[457] vdd gnd pinv_11
Xwl_driver_inv_en458 en en_bar[458] vdd gnd pinv_12
Xwl_driver_nand458 en_bar[458] in[458] net[458] vdd gnd pnand2_4
Xwl_driver_inv458 net[458] wl[458] vdd gnd pinv_11
Xwl_driver_inv_en459 en en_bar[459] vdd gnd pinv_12
Xwl_driver_nand459 en_bar[459] in[459] net[459] vdd gnd pnand2_4
Xwl_driver_inv459 net[459] wl[459] vdd gnd pinv_11
Xwl_driver_inv_en460 en en_bar[460] vdd gnd pinv_12
Xwl_driver_nand460 en_bar[460] in[460] net[460] vdd gnd pnand2_4
Xwl_driver_inv460 net[460] wl[460] vdd gnd pinv_11
Xwl_driver_inv_en461 en en_bar[461] vdd gnd pinv_12
Xwl_driver_nand461 en_bar[461] in[461] net[461] vdd gnd pnand2_4
Xwl_driver_inv461 net[461] wl[461] vdd gnd pinv_11
Xwl_driver_inv_en462 en en_bar[462] vdd gnd pinv_12
Xwl_driver_nand462 en_bar[462] in[462] net[462] vdd gnd pnand2_4
Xwl_driver_inv462 net[462] wl[462] vdd gnd pinv_11
Xwl_driver_inv_en463 en en_bar[463] vdd gnd pinv_12
Xwl_driver_nand463 en_bar[463] in[463] net[463] vdd gnd pnand2_4
Xwl_driver_inv463 net[463] wl[463] vdd gnd pinv_11
Xwl_driver_inv_en464 en en_bar[464] vdd gnd pinv_12
Xwl_driver_nand464 en_bar[464] in[464] net[464] vdd gnd pnand2_4
Xwl_driver_inv464 net[464] wl[464] vdd gnd pinv_11
Xwl_driver_inv_en465 en en_bar[465] vdd gnd pinv_12
Xwl_driver_nand465 en_bar[465] in[465] net[465] vdd gnd pnand2_4
Xwl_driver_inv465 net[465] wl[465] vdd gnd pinv_11
Xwl_driver_inv_en466 en en_bar[466] vdd gnd pinv_12
Xwl_driver_nand466 en_bar[466] in[466] net[466] vdd gnd pnand2_4
Xwl_driver_inv466 net[466] wl[466] vdd gnd pinv_11
Xwl_driver_inv_en467 en en_bar[467] vdd gnd pinv_12
Xwl_driver_nand467 en_bar[467] in[467] net[467] vdd gnd pnand2_4
Xwl_driver_inv467 net[467] wl[467] vdd gnd pinv_11
Xwl_driver_inv_en468 en en_bar[468] vdd gnd pinv_12
Xwl_driver_nand468 en_bar[468] in[468] net[468] vdd gnd pnand2_4
Xwl_driver_inv468 net[468] wl[468] vdd gnd pinv_11
Xwl_driver_inv_en469 en en_bar[469] vdd gnd pinv_12
Xwl_driver_nand469 en_bar[469] in[469] net[469] vdd gnd pnand2_4
Xwl_driver_inv469 net[469] wl[469] vdd gnd pinv_11
Xwl_driver_inv_en470 en en_bar[470] vdd gnd pinv_12
Xwl_driver_nand470 en_bar[470] in[470] net[470] vdd gnd pnand2_4
Xwl_driver_inv470 net[470] wl[470] vdd gnd pinv_11
Xwl_driver_inv_en471 en en_bar[471] vdd gnd pinv_12
Xwl_driver_nand471 en_bar[471] in[471] net[471] vdd gnd pnand2_4
Xwl_driver_inv471 net[471] wl[471] vdd gnd pinv_11
Xwl_driver_inv_en472 en en_bar[472] vdd gnd pinv_12
Xwl_driver_nand472 en_bar[472] in[472] net[472] vdd gnd pnand2_4
Xwl_driver_inv472 net[472] wl[472] vdd gnd pinv_11
Xwl_driver_inv_en473 en en_bar[473] vdd gnd pinv_12
Xwl_driver_nand473 en_bar[473] in[473] net[473] vdd gnd pnand2_4
Xwl_driver_inv473 net[473] wl[473] vdd gnd pinv_11
Xwl_driver_inv_en474 en en_bar[474] vdd gnd pinv_12
Xwl_driver_nand474 en_bar[474] in[474] net[474] vdd gnd pnand2_4
Xwl_driver_inv474 net[474] wl[474] vdd gnd pinv_11
Xwl_driver_inv_en475 en en_bar[475] vdd gnd pinv_12
Xwl_driver_nand475 en_bar[475] in[475] net[475] vdd gnd pnand2_4
Xwl_driver_inv475 net[475] wl[475] vdd gnd pinv_11
Xwl_driver_inv_en476 en en_bar[476] vdd gnd pinv_12
Xwl_driver_nand476 en_bar[476] in[476] net[476] vdd gnd pnand2_4
Xwl_driver_inv476 net[476] wl[476] vdd gnd pinv_11
Xwl_driver_inv_en477 en en_bar[477] vdd gnd pinv_12
Xwl_driver_nand477 en_bar[477] in[477] net[477] vdd gnd pnand2_4
Xwl_driver_inv477 net[477] wl[477] vdd gnd pinv_11
Xwl_driver_inv_en478 en en_bar[478] vdd gnd pinv_12
Xwl_driver_nand478 en_bar[478] in[478] net[478] vdd gnd pnand2_4
Xwl_driver_inv478 net[478] wl[478] vdd gnd pinv_11
Xwl_driver_inv_en479 en en_bar[479] vdd gnd pinv_12
Xwl_driver_nand479 en_bar[479] in[479] net[479] vdd gnd pnand2_4
Xwl_driver_inv479 net[479] wl[479] vdd gnd pinv_11
Xwl_driver_inv_en480 en en_bar[480] vdd gnd pinv_12
Xwl_driver_nand480 en_bar[480] in[480] net[480] vdd gnd pnand2_4
Xwl_driver_inv480 net[480] wl[480] vdd gnd pinv_11
Xwl_driver_inv_en481 en en_bar[481] vdd gnd pinv_12
Xwl_driver_nand481 en_bar[481] in[481] net[481] vdd gnd pnand2_4
Xwl_driver_inv481 net[481] wl[481] vdd gnd pinv_11
Xwl_driver_inv_en482 en en_bar[482] vdd gnd pinv_12
Xwl_driver_nand482 en_bar[482] in[482] net[482] vdd gnd pnand2_4
Xwl_driver_inv482 net[482] wl[482] vdd gnd pinv_11
Xwl_driver_inv_en483 en en_bar[483] vdd gnd pinv_12
Xwl_driver_nand483 en_bar[483] in[483] net[483] vdd gnd pnand2_4
Xwl_driver_inv483 net[483] wl[483] vdd gnd pinv_11
Xwl_driver_inv_en484 en en_bar[484] vdd gnd pinv_12
Xwl_driver_nand484 en_bar[484] in[484] net[484] vdd gnd pnand2_4
Xwl_driver_inv484 net[484] wl[484] vdd gnd pinv_11
Xwl_driver_inv_en485 en en_bar[485] vdd gnd pinv_12
Xwl_driver_nand485 en_bar[485] in[485] net[485] vdd gnd pnand2_4
Xwl_driver_inv485 net[485] wl[485] vdd gnd pinv_11
Xwl_driver_inv_en486 en en_bar[486] vdd gnd pinv_12
Xwl_driver_nand486 en_bar[486] in[486] net[486] vdd gnd pnand2_4
Xwl_driver_inv486 net[486] wl[486] vdd gnd pinv_11
Xwl_driver_inv_en487 en en_bar[487] vdd gnd pinv_12
Xwl_driver_nand487 en_bar[487] in[487] net[487] vdd gnd pnand2_4
Xwl_driver_inv487 net[487] wl[487] vdd gnd pinv_11
Xwl_driver_inv_en488 en en_bar[488] vdd gnd pinv_12
Xwl_driver_nand488 en_bar[488] in[488] net[488] vdd gnd pnand2_4
Xwl_driver_inv488 net[488] wl[488] vdd gnd pinv_11
Xwl_driver_inv_en489 en en_bar[489] vdd gnd pinv_12
Xwl_driver_nand489 en_bar[489] in[489] net[489] vdd gnd pnand2_4
Xwl_driver_inv489 net[489] wl[489] vdd gnd pinv_11
Xwl_driver_inv_en490 en en_bar[490] vdd gnd pinv_12
Xwl_driver_nand490 en_bar[490] in[490] net[490] vdd gnd pnand2_4
Xwl_driver_inv490 net[490] wl[490] vdd gnd pinv_11
Xwl_driver_inv_en491 en en_bar[491] vdd gnd pinv_12
Xwl_driver_nand491 en_bar[491] in[491] net[491] vdd gnd pnand2_4
Xwl_driver_inv491 net[491] wl[491] vdd gnd pinv_11
Xwl_driver_inv_en492 en en_bar[492] vdd gnd pinv_12
Xwl_driver_nand492 en_bar[492] in[492] net[492] vdd gnd pnand2_4
Xwl_driver_inv492 net[492] wl[492] vdd gnd pinv_11
Xwl_driver_inv_en493 en en_bar[493] vdd gnd pinv_12
Xwl_driver_nand493 en_bar[493] in[493] net[493] vdd gnd pnand2_4
Xwl_driver_inv493 net[493] wl[493] vdd gnd pinv_11
Xwl_driver_inv_en494 en en_bar[494] vdd gnd pinv_12
Xwl_driver_nand494 en_bar[494] in[494] net[494] vdd gnd pnand2_4
Xwl_driver_inv494 net[494] wl[494] vdd gnd pinv_11
Xwl_driver_inv_en495 en en_bar[495] vdd gnd pinv_12
Xwl_driver_nand495 en_bar[495] in[495] net[495] vdd gnd pnand2_4
Xwl_driver_inv495 net[495] wl[495] vdd gnd pinv_11
Xwl_driver_inv_en496 en en_bar[496] vdd gnd pinv_12
Xwl_driver_nand496 en_bar[496] in[496] net[496] vdd gnd pnand2_4
Xwl_driver_inv496 net[496] wl[496] vdd gnd pinv_11
Xwl_driver_inv_en497 en en_bar[497] vdd gnd pinv_12
Xwl_driver_nand497 en_bar[497] in[497] net[497] vdd gnd pnand2_4
Xwl_driver_inv497 net[497] wl[497] vdd gnd pinv_11
Xwl_driver_inv_en498 en en_bar[498] vdd gnd pinv_12
Xwl_driver_nand498 en_bar[498] in[498] net[498] vdd gnd pnand2_4
Xwl_driver_inv498 net[498] wl[498] vdd gnd pinv_11
Xwl_driver_inv_en499 en en_bar[499] vdd gnd pinv_12
Xwl_driver_nand499 en_bar[499] in[499] net[499] vdd gnd pnand2_4
Xwl_driver_inv499 net[499] wl[499] vdd gnd pinv_11
Xwl_driver_inv_en500 en en_bar[500] vdd gnd pinv_12
Xwl_driver_nand500 en_bar[500] in[500] net[500] vdd gnd pnand2_4
Xwl_driver_inv500 net[500] wl[500] vdd gnd pinv_11
Xwl_driver_inv_en501 en en_bar[501] vdd gnd pinv_12
Xwl_driver_nand501 en_bar[501] in[501] net[501] vdd gnd pnand2_4
Xwl_driver_inv501 net[501] wl[501] vdd gnd pinv_11
Xwl_driver_inv_en502 en en_bar[502] vdd gnd pinv_12
Xwl_driver_nand502 en_bar[502] in[502] net[502] vdd gnd pnand2_4
Xwl_driver_inv502 net[502] wl[502] vdd gnd pinv_11
Xwl_driver_inv_en503 en en_bar[503] vdd gnd pinv_12
Xwl_driver_nand503 en_bar[503] in[503] net[503] vdd gnd pnand2_4
Xwl_driver_inv503 net[503] wl[503] vdd gnd pinv_11
Xwl_driver_inv_en504 en en_bar[504] vdd gnd pinv_12
Xwl_driver_nand504 en_bar[504] in[504] net[504] vdd gnd pnand2_4
Xwl_driver_inv504 net[504] wl[504] vdd gnd pinv_11
Xwl_driver_inv_en505 en en_bar[505] vdd gnd pinv_12
Xwl_driver_nand505 en_bar[505] in[505] net[505] vdd gnd pnand2_4
Xwl_driver_inv505 net[505] wl[505] vdd gnd pinv_11
Xwl_driver_inv_en506 en en_bar[506] vdd gnd pinv_12
Xwl_driver_nand506 en_bar[506] in[506] net[506] vdd gnd pnand2_4
Xwl_driver_inv506 net[506] wl[506] vdd gnd pinv_11
Xwl_driver_inv_en507 en en_bar[507] vdd gnd pinv_12
Xwl_driver_nand507 en_bar[507] in[507] net[507] vdd gnd pnand2_4
Xwl_driver_inv507 net[507] wl[507] vdd gnd pinv_11
Xwl_driver_inv_en508 en en_bar[508] vdd gnd pinv_12
Xwl_driver_nand508 en_bar[508] in[508] net[508] vdd gnd pnand2_4
Xwl_driver_inv508 net[508] wl[508] vdd gnd pinv_11
Xwl_driver_inv_en509 en en_bar[509] vdd gnd pinv_12
Xwl_driver_nand509 en_bar[509] in[509] net[509] vdd gnd pnand2_4
Xwl_driver_inv509 net[509] wl[509] vdd gnd pinv_11
Xwl_driver_inv_en510 en en_bar[510] vdd gnd pinv_12
Xwl_driver_nand510 en_bar[510] in[510] net[510] vdd gnd pnand2_4
Xwl_driver_inv510 net[510] wl[510] vdd gnd pinv_11
Xwl_driver_inv_en511 en en_bar[511] vdd gnd pinv_12
Xwl_driver_nand511 en_bar[511] in[511] net[511] vdd gnd pnand2_4
Xwl_driver_inv511 net[511] wl[511] vdd gnd pinv_11
.ENDS wordline_driver

.SUBCKT pinv_13 A Z vdd gnd
Mpinv_pmos Z A vdd vdd pmos_vtg m=1 w=0.27u l=0.05u pd=0.64u ps=0.64u as=0.03375p ad=0.03375p
Mpinv_nmos Z A gnd gnd nmos_vtg m=1 w=0.09u l=0.05u pd=0.28u ps=0.28u as=0.01125p ad=0.01125p
.ENDS pinv_13

.SUBCKT bank DATA[0] DATA[1] DATA[2] DATA[3] DATA[4] DATA[5] DATA[6] DATA[7] DATA[8] DATA[9] DATA[10] DATA[11] DATA[12] DATA[13] DATA[14] DATA[15] DATA[16] DATA[17] DATA[18] DATA[19] DATA[20] DATA[21] DATA[22] DATA[23] DATA[24] DATA[25] DATA[26] DATA[27] DATA[28] DATA[29] DATA[30] DATA[31] ADDR[0] ADDR[1] ADDR[2] ADDR[3] ADDR[4] ADDR[5] ADDR[6] ADDR[7] ADDR[8] ADDR[9] ADDR[10] s_en w_en tri_en_bar tri_en clk_bar clk_buf vdd gnd
Xbitcell_array bl[0] br[0] bl[1] br[1] bl[2] br[2] bl[3] br[3] bl[4] br[4] bl[5] br[5] bl[6] br[6] bl[7] br[7] bl[8] br[8] bl[9] br[9] bl[10] br[10] bl[11] br[11] bl[12] br[12] bl[13] br[13] bl[14] br[14] bl[15] br[15] bl[16] br[16] bl[17] br[17] bl[18] br[18] bl[19] br[19] bl[20] br[20] bl[21] br[21] bl[22] br[22] bl[23] br[23] bl[24] br[24] bl[25] br[25] bl[26] br[26] bl[27] br[27] bl[28] br[28] bl[29] br[29] bl[30] br[30] bl[31] br[31] bl[32] br[32] bl[33] br[33] bl[34] br[34] bl[35] br[35] bl[36] br[36] bl[37] br[37] bl[38] br[38] bl[39] br[39] bl[40] br[40] bl[41] br[41] bl[42] br[42] bl[43] br[43] bl[44] br[44] bl[45] br[45] bl[46] br[46] bl[47] br[47] bl[48] br[48] bl[49] br[49] bl[50] br[50] bl[51] br[51] bl[52] br[52] bl[53] br[53] bl[54] br[54] bl[55] br[55] bl[56] br[56] bl[57] br[57] bl[58] br[58] bl[59] br[59] bl[60] br[60] bl[61] br[61] bl[62] br[62] bl[63] br[63] bl[64] br[64] bl[65] br[65] bl[66] br[66] bl[67] br[67] bl[68] br[68] bl[69] br[69] bl[70] br[70] bl[71] br[71] bl[72] br[72] bl[73] br[73] bl[74] br[74] bl[75] br[75] bl[76] br[76] bl[77] br[77] bl[78] br[78] bl[79] br[79] bl[80] br[80] bl[81] br[81] bl[82] br[82] bl[83] br[83] bl[84] br[84] bl[85] br[85] bl[86] br[86] bl[87] br[87] bl[88] br[88] bl[89] br[89] bl[90] br[90] bl[91] br[91] bl[92] br[92] bl[93] br[93] bl[94] br[94] bl[95] br[95] bl[96] br[96] bl[97] br[97] bl[98] br[98] bl[99] br[99] bl[100] br[100] bl[101] br[101] bl[102] br[102] bl[103] br[103] bl[104] br[104] bl[105] br[105] bl[106] br[106] bl[107] br[107] bl[108] br[108] bl[109] br[109] bl[110] br[110] bl[111] br[111] bl[112] br[112] bl[113] br[113] bl[114] br[114] bl[115] br[115] bl[116] br[116] bl[117] br[117] bl[118] br[118] bl[119] br[119] bl[120] br[120] bl[121] br[121] bl[122] br[122] bl[123] br[123] bl[124] br[124] bl[125] br[125] bl[126] br[126] bl[127] br[127] wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] wl[128] wl[129] wl[130] wl[131] wl[132] wl[133] wl[134] wl[135] wl[136] wl[137] wl[138] wl[139] wl[140] wl[141] wl[142] wl[143] wl[144] wl[145] wl[146] wl[147] wl[148] wl[149] wl[150] wl[151] wl[152] wl[153] wl[154] wl[155] wl[156] wl[157] wl[158] wl[159] wl[160] wl[161] wl[162] wl[163] wl[164] wl[165] wl[166] wl[167] wl[168] wl[169] wl[170] wl[171] wl[172] wl[173] wl[174] wl[175] wl[176] wl[177] wl[178] wl[179] wl[180] wl[181] wl[182] wl[183] wl[184] wl[185] wl[186] wl[187] wl[188] wl[189] wl[190] wl[191] wl[192] wl[193] wl[194] wl[195] wl[196] wl[197] wl[198] wl[199] wl[200] wl[201] wl[202] wl[203] wl[204] wl[205] wl[206] wl[207] wl[208] wl[209] wl[210] wl[211] wl[212] wl[213] wl[214] wl[215] wl[216] wl[217] wl[218] wl[219] wl[220] wl[221] wl[222] wl[223] wl[224] wl[225] wl[226] wl[227] wl[228] wl[229] wl[230] wl[231] wl[232] wl[233] wl[234] wl[235] wl[236] wl[237] wl[238] wl[239] wl[240] wl[241] wl[242] wl[243] wl[244] wl[245] wl[246] wl[247] wl[248] wl[249] wl[250] wl[251] wl[252] wl[253] wl[254] wl[255] wl[256] wl[257] wl[258] wl[259] wl[260] wl[261] wl[262] wl[263] wl[264] wl[265] wl[266] wl[267] wl[268] wl[269] wl[270] wl[271] wl[272] wl[273] wl[274] wl[275] wl[276] wl[277] wl[278] wl[279] wl[280] wl[281] wl[282] wl[283] wl[284] wl[285] wl[286] wl[287] wl[288] wl[289] wl[290] wl[291] wl[292] wl[293] wl[294] wl[295] wl[296] wl[297] wl[298] wl[299] wl[300] wl[301] wl[302] wl[303] wl[304] wl[305] wl[306] wl[307] wl[308] wl[309] wl[310] wl[311] wl[312] wl[313] wl[314] wl[315] wl[316] wl[317] wl[318] wl[319] wl[320] wl[321] wl[322] wl[323] wl[324] wl[325] wl[326] wl[327] wl[328] wl[329] wl[330] wl[331] wl[332] wl[333] wl[334] wl[335] wl[336] wl[337] wl[338] wl[339] wl[340] wl[341] wl[342] wl[343] wl[344] wl[345] wl[346] wl[347] wl[348] wl[349] wl[350] wl[351] wl[352] wl[353] wl[354] wl[355] wl[356] wl[357] wl[358] wl[359] wl[360] wl[361] wl[362] wl[363] wl[364] wl[365] wl[366] wl[367] wl[368] wl[369] wl[370] wl[371] wl[372] wl[373] wl[374] wl[375] wl[376] wl[377] wl[378] wl[379] wl[380] wl[381] wl[382] wl[383] wl[384] wl[385] wl[386] wl[387] wl[388] wl[389] wl[390] wl[391] wl[392] wl[393] wl[394] wl[395] wl[396] wl[397] wl[398] wl[399] wl[400] wl[401] wl[402] wl[403] wl[404] wl[405] wl[406] wl[407] wl[408] wl[409] wl[410] wl[411] wl[412] wl[413] wl[414] wl[415] wl[416] wl[417] wl[418] wl[419] wl[420] wl[421] wl[422] wl[423] wl[424] wl[425] wl[426] wl[427] wl[428] wl[429] wl[430] wl[431] wl[432] wl[433] wl[434] wl[435] wl[436] wl[437] wl[438] wl[439] wl[440] wl[441] wl[442] wl[443] wl[444] wl[445] wl[446] wl[447] wl[448] wl[449] wl[450] wl[451] wl[452] wl[453] wl[454] wl[455] wl[456] wl[457] wl[458] wl[459] wl[460] wl[461] wl[462] wl[463] wl[464] wl[465] wl[466] wl[467] wl[468] wl[469] wl[470] wl[471] wl[472] wl[473] wl[474] wl[475] wl[476] wl[477] wl[478] wl[479] wl[480] wl[481] wl[482] wl[483] wl[484] wl[485] wl[486] wl[487] wl[488] wl[489] wl[490] wl[491] wl[492] wl[493] wl[494] wl[495] wl[496] wl[497] wl[498] wl[499] wl[500] wl[501] wl[502] wl[503] wl[504] wl[505] wl[506] wl[507] wl[508] wl[509] wl[510] wl[511] vdd gnd bitcell_array
Xprecharge_array bl[0] br[0] bl[1] br[1] bl[2] br[2] bl[3] br[3] bl[4] br[4] bl[5] br[5] bl[6] br[6] bl[7] br[7] bl[8] br[8] bl[9] br[9] bl[10] br[10] bl[11] br[11] bl[12] br[12] bl[13] br[13] bl[14] br[14] bl[15] br[15] bl[16] br[16] bl[17] br[17] bl[18] br[18] bl[19] br[19] bl[20] br[20] bl[21] br[21] bl[22] br[22] bl[23] br[23] bl[24] br[24] bl[25] br[25] bl[26] br[26] bl[27] br[27] bl[28] br[28] bl[29] br[29] bl[30] br[30] bl[31] br[31] bl[32] br[32] bl[33] br[33] bl[34] br[34] bl[35] br[35] bl[36] br[36] bl[37] br[37] bl[38] br[38] bl[39] br[39] bl[40] br[40] bl[41] br[41] bl[42] br[42] bl[43] br[43] bl[44] br[44] bl[45] br[45] bl[46] br[46] bl[47] br[47] bl[48] br[48] bl[49] br[49] bl[50] br[50] bl[51] br[51] bl[52] br[52] bl[53] br[53] bl[54] br[54] bl[55] br[55] bl[56] br[56] bl[57] br[57] bl[58] br[58] bl[59] br[59] bl[60] br[60] bl[61] br[61] bl[62] br[62] bl[63] br[63] bl[64] br[64] bl[65] br[65] bl[66] br[66] bl[67] br[67] bl[68] br[68] bl[69] br[69] bl[70] br[70] bl[71] br[71] bl[72] br[72] bl[73] br[73] bl[74] br[74] bl[75] br[75] bl[76] br[76] bl[77] br[77] bl[78] br[78] bl[79] br[79] bl[80] br[80] bl[81] br[81] bl[82] br[82] bl[83] br[83] bl[84] br[84] bl[85] br[85] bl[86] br[86] bl[87] br[87] bl[88] br[88] bl[89] br[89] bl[90] br[90] bl[91] br[91] bl[92] br[92] bl[93] br[93] bl[94] br[94] bl[95] br[95] bl[96] br[96] bl[97] br[97] bl[98] br[98] bl[99] br[99] bl[100] br[100] bl[101] br[101] bl[102] br[102] bl[103] br[103] bl[104] br[104] bl[105] br[105] bl[106] br[106] bl[107] br[107] bl[108] br[108] bl[109] br[109] bl[110] br[110] bl[111] br[111] bl[112] br[112] bl[113] br[113] bl[114] br[114] bl[115] br[115] bl[116] br[116] bl[117] br[117] bl[118] br[118] bl[119] br[119] bl[120] br[120] bl[121] br[121] bl[122] br[122] bl[123] br[123] bl[124] br[124] bl[125] br[125] bl[126] br[126] bl[127] br[127] clk_bar vdd precharge_array
Xcolumn_mux_array bl[0] br[0] bl[1] br[1] bl[2] br[2] bl[3] br[3] bl[4] br[4] bl[5] br[5] bl[6] br[6] bl[7] br[7] bl[8] br[8] bl[9] br[9] bl[10] br[10] bl[11] br[11] bl[12] br[12] bl[13] br[13] bl[14] br[14] bl[15] br[15] bl[16] br[16] bl[17] br[17] bl[18] br[18] bl[19] br[19] bl[20] br[20] bl[21] br[21] bl[22] br[22] bl[23] br[23] bl[24] br[24] bl[25] br[25] bl[26] br[26] bl[27] br[27] bl[28] br[28] bl[29] br[29] bl[30] br[30] bl[31] br[31] bl[32] br[32] bl[33] br[33] bl[34] br[34] bl[35] br[35] bl[36] br[36] bl[37] br[37] bl[38] br[38] bl[39] br[39] bl[40] br[40] bl[41] br[41] bl[42] br[42] bl[43] br[43] bl[44] br[44] bl[45] br[45] bl[46] br[46] bl[47] br[47] bl[48] br[48] bl[49] br[49] bl[50] br[50] bl[51] br[51] bl[52] br[52] bl[53] br[53] bl[54] br[54] bl[55] br[55] bl[56] br[56] bl[57] br[57] bl[58] br[58] bl[59] br[59] bl[60] br[60] bl[61] br[61] bl[62] br[62] bl[63] br[63] bl[64] br[64] bl[65] br[65] bl[66] br[66] bl[67] br[67] bl[68] br[68] bl[69] br[69] bl[70] br[70] bl[71] br[71] bl[72] br[72] bl[73] br[73] bl[74] br[74] bl[75] br[75] bl[76] br[76] bl[77] br[77] bl[78] br[78] bl[79] br[79] bl[80] br[80] bl[81] br[81] bl[82] br[82] bl[83] br[83] bl[84] br[84] bl[85] br[85] bl[86] br[86] bl[87] br[87] bl[88] br[88] bl[89] br[89] bl[90] br[90] bl[91] br[91] bl[92] br[92] bl[93] br[93] bl[94] br[94] bl[95] br[95] bl[96] br[96] bl[97] br[97] bl[98] br[98] bl[99] br[99] bl[100] br[100] bl[101] br[101] bl[102] br[102] bl[103] br[103] bl[104] br[104] bl[105] br[105] bl[106] br[106] bl[107] br[107] bl[108] br[108] bl[109] br[109] bl[110] br[110] bl[111] br[111] bl[112] br[112] bl[113] br[113] bl[114] br[114] bl[115] br[115] bl[116] br[116] bl[117] br[117] bl[118] br[118] bl[119] br[119] bl[120] br[120] bl[121] br[121] bl[122] br[122] bl[123] br[123] bl[124] br[124] bl[125] br[125] bl[126] br[126] bl[127] br[127] sel[0] sel[1] sel[2] sel[3] bl_out[0] br_out[0] bl_out[1] br_out[1] bl_out[2] br_out[2] bl_out[3] br_out[3] bl_out[4] br_out[4] bl_out[5] br_out[5] bl_out[6] br_out[6] bl_out[7] br_out[7] bl_out[8] br_out[8] bl_out[9] br_out[9] bl_out[10] br_out[10] bl_out[11] br_out[11] bl_out[12] br_out[12] bl_out[13] br_out[13] bl_out[14] br_out[14] bl_out[15] br_out[15] bl_out[16] br_out[16] bl_out[17] br_out[17] bl_out[18] br_out[18] bl_out[19] br_out[19] bl_out[20] br_out[20] bl_out[21] br_out[21] bl_out[22] br_out[22] bl_out[23] br_out[23] bl_out[24] br_out[24] bl_out[25] br_out[25] bl_out[26] br_out[26] bl_out[27] br_out[27] bl_out[28] br_out[28] bl_out[29] br_out[29] bl_out[30] br_out[30] bl_out[31] br_out[31] gnd columnmux_array
Xcol_address_decoder A[9] A[10] sel[0] sel[1] sel[2] sel[3] vdd gnd pre2x4
Xsense_amp_array data_out[0] bl_out[0] br_out[0] data_out[1] bl_out[1] br_out[1] data_out[2] bl_out[2] br_out[2] data_out[3] bl_out[3] br_out[3] data_out[4] bl_out[4] br_out[4] data_out[5] bl_out[5] br_out[5] data_out[6] bl_out[6] br_out[6] data_out[7] bl_out[7] br_out[7] data_out[8] bl_out[8] br_out[8] data_out[9] bl_out[9] br_out[9] data_out[10] bl_out[10] br_out[10] data_out[11] bl_out[11] br_out[11] data_out[12] bl_out[12] br_out[12] data_out[13] bl_out[13] br_out[13] data_out[14] bl_out[14] br_out[14] data_out[15] bl_out[15] br_out[15] data_out[16] bl_out[16] br_out[16] data_out[17] bl_out[17] br_out[17] data_out[18] bl_out[18] br_out[18] data_out[19] bl_out[19] br_out[19] data_out[20] bl_out[20] br_out[20] data_out[21] bl_out[21] br_out[21] data_out[22] bl_out[22] br_out[22] data_out[23] bl_out[23] br_out[23] data_out[24] bl_out[24] br_out[24] data_out[25] bl_out[25] br_out[25] data_out[26] bl_out[26] br_out[26] data_out[27] bl_out[27] br_out[27] data_out[28] bl_out[28] br_out[28] data_out[29] bl_out[29] br_out[29] data_out[30] bl_out[30] br_out[30] data_out[31] bl_out[31] br_out[31] s_en vdd gnd sense_amp_array
Xwrite_driver_array data_in[0] data_in[1] data_in[2] data_in[3] data_in[4] data_in[5] data_in[6] data_in[7] data_in[8] data_in[9] data_in[10] data_in[11] data_in[12] data_in[13] data_in[14] data_in[15] data_in[16] data_in[17] data_in[18] data_in[19] data_in[20] data_in[21] data_in[22] data_in[23] data_in[24] data_in[25] data_in[26] data_in[27] data_in[28] data_in[29] data_in[30] data_in[31] bl_out[0] br_out[0] bl_out[1] br_out[1] bl_out[2] br_out[2] bl_out[3] br_out[3] bl_out[4] br_out[4] bl_out[5] br_out[5] bl_out[6] br_out[6] bl_out[7] br_out[7] bl_out[8] br_out[8] bl_out[9] br_out[9] bl_out[10] br_out[10] bl_out[11] br_out[11] bl_out[12] br_out[12] bl_out[13] br_out[13] bl_out[14] br_out[14] bl_out[15] br_out[15] bl_out[16] br_out[16] bl_out[17] br_out[17] bl_out[18] br_out[18] bl_out[19] br_out[19] bl_out[20] br_out[20] bl_out[21] br_out[21] bl_out[22] br_out[22] bl_out[23] br_out[23] bl_out[24] br_out[24] bl_out[25] br_out[25] bl_out[26] br_out[26] bl_out[27] br_out[27] bl_out[28] br_out[28] bl_out[29] br_out[29] bl_out[30] br_out[30] bl_out[31] br_out[31] w_en vdd gnd write_driver_array
Xdata_in_flop_array DATA[0] DATA[1] DATA[2] DATA[3] DATA[4] DATA[5] DATA[6] DATA[7] DATA[8] DATA[9] DATA[10] DATA[11] DATA[12] DATA[13] DATA[14] DATA[15] DATA[16] DATA[17] DATA[18] DATA[19] DATA[20] DATA[21] DATA[22] DATA[23] DATA[24] DATA[25] DATA[26] DATA[27] DATA[28] DATA[29] DATA[30] DATA[31] data_in[0] data_in_bar[0] data_in[1] data_in_bar[1] data_in[2] data_in_bar[2] data_in[3] data_in_bar[3] data_in[4] data_in_bar[4] data_in[5] data_in_bar[5] data_in[6] data_in_bar[6] data_in[7] data_in_bar[7] data_in[8] data_in_bar[8] data_in[9] data_in_bar[9] data_in[10] data_in_bar[10] data_in[11] data_in_bar[11] data_in[12] data_in_bar[12] data_in[13] data_in_bar[13] data_in[14] data_in_bar[14] data_in[15] data_in_bar[15] data_in[16] data_in_bar[16] data_in[17] data_in_bar[17] data_in[18] data_in_bar[18] data_in[19] data_in_bar[19] data_in[20] data_in_bar[20] data_in[21] data_in_bar[21] data_in[22] data_in_bar[22] data_in[23] data_in_bar[23] data_in[24] data_in_bar[24] data_in[25] data_in_bar[25] data_in[26] data_in_bar[26] data_in[27] data_in_bar[27] data_in[28] data_in_bar[28] data_in[29] data_in_bar[29] data_in[30] data_in_bar[30] data_in[31] data_in_bar[31] clk_bar vdd gnd msf_data_in
Xtri_gate_array data_out[0] data_out[1] data_out[2] data_out[3] data_out[4] data_out[5] data_out[6] data_out[7] data_out[8] data_out[9] data_out[10] data_out[11] data_out[12] data_out[13] data_out[14] data_out[15] data_out[16] data_out[17] data_out[18] data_out[19] data_out[20] data_out[21] data_out[22] data_out[23] data_out[24] data_out[25] data_out[26] data_out[27] data_out[28] data_out[29] data_out[30] data_out[31] DATA[0] DATA[1] DATA[2] DATA[3] DATA[4] DATA[5] DATA[6] DATA[7] DATA[8] DATA[9] DATA[10] DATA[11] DATA[12] DATA[13] DATA[14] DATA[15] DATA[16] DATA[17] DATA[18] DATA[19] DATA[20] DATA[21] DATA[22] DATA[23] DATA[24] DATA[25] DATA[26] DATA[27] DATA[28] DATA[29] DATA[30] DATA[31] tri_en tri_en_bar vdd gnd tri_gate_array
Xrow_decoder A[0] A[1] A[2] A[3] A[4] A[5] A[6] A[7] A[8] dec_out[0] dec_out[1] dec_out[2] dec_out[3] dec_out[4] dec_out[5] dec_out[6] dec_out[7] dec_out[8] dec_out[9] dec_out[10] dec_out[11] dec_out[12] dec_out[13] dec_out[14] dec_out[15] dec_out[16] dec_out[17] dec_out[18] dec_out[19] dec_out[20] dec_out[21] dec_out[22] dec_out[23] dec_out[24] dec_out[25] dec_out[26] dec_out[27] dec_out[28] dec_out[29] dec_out[30] dec_out[31] dec_out[32] dec_out[33] dec_out[34] dec_out[35] dec_out[36] dec_out[37] dec_out[38] dec_out[39] dec_out[40] dec_out[41] dec_out[42] dec_out[43] dec_out[44] dec_out[45] dec_out[46] dec_out[47] dec_out[48] dec_out[49] dec_out[50] dec_out[51] dec_out[52] dec_out[53] dec_out[54] dec_out[55] dec_out[56] dec_out[57] dec_out[58] dec_out[59] dec_out[60] dec_out[61] dec_out[62] dec_out[63] dec_out[64] dec_out[65] dec_out[66] dec_out[67] dec_out[68] dec_out[69] dec_out[70] dec_out[71] dec_out[72] dec_out[73] dec_out[74] dec_out[75] dec_out[76] dec_out[77] dec_out[78] dec_out[79] dec_out[80] dec_out[81] dec_out[82] dec_out[83] dec_out[84] dec_out[85] dec_out[86] dec_out[87] dec_out[88] dec_out[89] dec_out[90] dec_out[91] dec_out[92] dec_out[93] dec_out[94] dec_out[95] dec_out[96] dec_out[97] dec_out[98] dec_out[99] dec_out[100] dec_out[101] dec_out[102] dec_out[103] dec_out[104] dec_out[105] dec_out[106] dec_out[107] dec_out[108] dec_out[109] dec_out[110] dec_out[111] dec_out[112] dec_out[113] dec_out[114] dec_out[115] dec_out[116] dec_out[117] dec_out[118] dec_out[119] dec_out[120] dec_out[121] dec_out[122] dec_out[123] dec_out[124] dec_out[125] dec_out[126] dec_out[127] dec_out[128] dec_out[129] dec_out[130] dec_out[131] dec_out[132] dec_out[133] dec_out[134] dec_out[135] dec_out[136] dec_out[137] dec_out[138] dec_out[139] dec_out[140] dec_out[141] dec_out[142] dec_out[143] dec_out[144] dec_out[145] dec_out[146] dec_out[147] dec_out[148] dec_out[149] dec_out[150] dec_out[151] dec_out[152] dec_out[153] dec_out[154] dec_out[155] dec_out[156] dec_out[157] dec_out[158] dec_out[159] dec_out[160] dec_out[161] dec_out[162] dec_out[163] dec_out[164] dec_out[165] dec_out[166] dec_out[167] dec_out[168] dec_out[169] dec_out[170] dec_out[171] dec_out[172] dec_out[173] dec_out[174] dec_out[175] dec_out[176] dec_out[177] dec_out[178] dec_out[179] dec_out[180] dec_out[181] dec_out[182] dec_out[183] dec_out[184] dec_out[185] dec_out[186] dec_out[187] dec_out[188] dec_out[189] dec_out[190] dec_out[191] dec_out[192] dec_out[193] dec_out[194] dec_out[195] dec_out[196] dec_out[197] dec_out[198] dec_out[199] dec_out[200] dec_out[201] dec_out[202] dec_out[203] dec_out[204] dec_out[205] dec_out[206] dec_out[207] dec_out[208] dec_out[209] dec_out[210] dec_out[211] dec_out[212] dec_out[213] dec_out[214] dec_out[215] dec_out[216] dec_out[217] dec_out[218] dec_out[219] dec_out[220] dec_out[221] dec_out[222] dec_out[223] dec_out[224] dec_out[225] dec_out[226] dec_out[227] dec_out[228] dec_out[229] dec_out[230] dec_out[231] dec_out[232] dec_out[233] dec_out[234] dec_out[235] dec_out[236] dec_out[237] dec_out[238] dec_out[239] dec_out[240] dec_out[241] dec_out[242] dec_out[243] dec_out[244] dec_out[245] dec_out[246] dec_out[247] dec_out[248] dec_out[249] dec_out[250] dec_out[251] dec_out[252] dec_out[253] dec_out[254] dec_out[255] dec_out[256] dec_out[257] dec_out[258] dec_out[259] dec_out[260] dec_out[261] dec_out[262] dec_out[263] dec_out[264] dec_out[265] dec_out[266] dec_out[267] dec_out[268] dec_out[269] dec_out[270] dec_out[271] dec_out[272] dec_out[273] dec_out[274] dec_out[275] dec_out[276] dec_out[277] dec_out[278] dec_out[279] dec_out[280] dec_out[281] dec_out[282] dec_out[283] dec_out[284] dec_out[285] dec_out[286] dec_out[287] dec_out[288] dec_out[289] dec_out[290] dec_out[291] dec_out[292] dec_out[293] dec_out[294] dec_out[295] dec_out[296] dec_out[297] dec_out[298] dec_out[299] dec_out[300] dec_out[301] dec_out[302] dec_out[303] dec_out[304] dec_out[305] dec_out[306] dec_out[307] dec_out[308] dec_out[309] dec_out[310] dec_out[311] dec_out[312] dec_out[313] dec_out[314] dec_out[315] dec_out[316] dec_out[317] dec_out[318] dec_out[319] dec_out[320] dec_out[321] dec_out[322] dec_out[323] dec_out[324] dec_out[325] dec_out[326] dec_out[327] dec_out[328] dec_out[329] dec_out[330] dec_out[331] dec_out[332] dec_out[333] dec_out[334] dec_out[335] dec_out[336] dec_out[337] dec_out[338] dec_out[339] dec_out[340] dec_out[341] dec_out[342] dec_out[343] dec_out[344] dec_out[345] dec_out[346] dec_out[347] dec_out[348] dec_out[349] dec_out[350] dec_out[351] dec_out[352] dec_out[353] dec_out[354] dec_out[355] dec_out[356] dec_out[357] dec_out[358] dec_out[359] dec_out[360] dec_out[361] dec_out[362] dec_out[363] dec_out[364] dec_out[365] dec_out[366] dec_out[367] dec_out[368] dec_out[369] dec_out[370] dec_out[371] dec_out[372] dec_out[373] dec_out[374] dec_out[375] dec_out[376] dec_out[377] dec_out[378] dec_out[379] dec_out[380] dec_out[381] dec_out[382] dec_out[383] dec_out[384] dec_out[385] dec_out[386] dec_out[387] dec_out[388] dec_out[389] dec_out[390] dec_out[391] dec_out[392] dec_out[393] dec_out[394] dec_out[395] dec_out[396] dec_out[397] dec_out[398] dec_out[399] dec_out[400] dec_out[401] dec_out[402] dec_out[403] dec_out[404] dec_out[405] dec_out[406] dec_out[407] dec_out[408] dec_out[409] dec_out[410] dec_out[411] dec_out[412] dec_out[413] dec_out[414] dec_out[415] dec_out[416] dec_out[417] dec_out[418] dec_out[419] dec_out[420] dec_out[421] dec_out[422] dec_out[423] dec_out[424] dec_out[425] dec_out[426] dec_out[427] dec_out[428] dec_out[429] dec_out[430] dec_out[431] dec_out[432] dec_out[433] dec_out[434] dec_out[435] dec_out[436] dec_out[437] dec_out[438] dec_out[439] dec_out[440] dec_out[441] dec_out[442] dec_out[443] dec_out[444] dec_out[445] dec_out[446] dec_out[447] dec_out[448] dec_out[449] dec_out[450] dec_out[451] dec_out[452] dec_out[453] dec_out[454] dec_out[455] dec_out[456] dec_out[457] dec_out[458] dec_out[459] dec_out[460] dec_out[461] dec_out[462] dec_out[463] dec_out[464] dec_out[465] dec_out[466] dec_out[467] dec_out[468] dec_out[469] dec_out[470] dec_out[471] dec_out[472] dec_out[473] dec_out[474] dec_out[475] dec_out[476] dec_out[477] dec_out[478] dec_out[479] dec_out[480] dec_out[481] dec_out[482] dec_out[483] dec_out[484] dec_out[485] dec_out[486] dec_out[487] dec_out[488] dec_out[489] dec_out[490] dec_out[491] dec_out[492] dec_out[493] dec_out[494] dec_out[495] dec_out[496] dec_out[497] dec_out[498] dec_out[499] dec_out[500] dec_out[501] dec_out[502] dec_out[503] dec_out[504] dec_out[505] dec_out[506] dec_out[507] dec_out[508] dec_out[509] dec_out[510] dec_out[511] vdd gnd hierarchical_decoder_512rows
Xwordline_driver dec_out[0] dec_out[1] dec_out[2] dec_out[3] dec_out[4] dec_out[5] dec_out[6] dec_out[7] dec_out[8] dec_out[9] dec_out[10] dec_out[11] dec_out[12] dec_out[13] dec_out[14] dec_out[15] dec_out[16] dec_out[17] dec_out[18] dec_out[19] dec_out[20] dec_out[21] dec_out[22] dec_out[23] dec_out[24] dec_out[25] dec_out[26] dec_out[27] dec_out[28] dec_out[29] dec_out[30] dec_out[31] dec_out[32] dec_out[33] dec_out[34] dec_out[35] dec_out[36] dec_out[37] dec_out[38] dec_out[39] dec_out[40] dec_out[41] dec_out[42] dec_out[43] dec_out[44] dec_out[45] dec_out[46] dec_out[47] dec_out[48] dec_out[49] dec_out[50] dec_out[51] dec_out[52] dec_out[53] dec_out[54] dec_out[55] dec_out[56] dec_out[57] dec_out[58] dec_out[59] dec_out[60] dec_out[61] dec_out[62] dec_out[63] dec_out[64] dec_out[65] dec_out[66] dec_out[67] dec_out[68] dec_out[69] dec_out[70] dec_out[71] dec_out[72] dec_out[73] dec_out[74] dec_out[75] dec_out[76] dec_out[77] dec_out[78] dec_out[79] dec_out[80] dec_out[81] dec_out[82] dec_out[83] dec_out[84] dec_out[85] dec_out[86] dec_out[87] dec_out[88] dec_out[89] dec_out[90] dec_out[91] dec_out[92] dec_out[93] dec_out[94] dec_out[95] dec_out[96] dec_out[97] dec_out[98] dec_out[99] dec_out[100] dec_out[101] dec_out[102] dec_out[103] dec_out[104] dec_out[105] dec_out[106] dec_out[107] dec_out[108] dec_out[109] dec_out[110] dec_out[111] dec_out[112] dec_out[113] dec_out[114] dec_out[115] dec_out[116] dec_out[117] dec_out[118] dec_out[119] dec_out[120] dec_out[121] dec_out[122] dec_out[123] dec_out[124] dec_out[125] dec_out[126] dec_out[127] dec_out[128] dec_out[129] dec_out[130] dec_out[131] dec_out[132] dec_out[133] dec_out[134] dec_out[135] dec_out[136] dec_out[137] dec_out[138] dec_out[139] dec_out[140] dec_out[141] dec_out[142] dec_out[143] dec_out[144] dec_out[145] dec_out[146] dec_out[147] dec_out[148] dec_out[149] dec_out[150] dec_out[151] dec_out[152] dec_out[153] dec_out[154] dec_out[155] dec_out[156] dec_out[157] dec_out[158] dec_out[159] dec_out[160] dec_out[161] dec_out[162] dec_out[163] dec_out[164] dec_out[165] dec_out[166] dec_out[167] dec_out[168] dec_out[169] dec_out[170] dec_out[171] dec_out[172] dec_out[173] dec_out[174] dec_out[175] dec_out[176] dec_out[177] dec_out[178] dec_out[179] dec_out[180] dec_out[181] dec_out[182] dec_out[183] dec_out[184] dec_out[185] dec_out[186] dec_out[187] dec_out[188] dec_out[189] dec_out[190] dec_out[191] dec_out[192] dec_out[193] dec_out[194] dec_out[195] dec_out[196] dec_out[197] dec_out[198] dec_out[199] dec_out[200] dec_out[201] dec_out[202] dec_out[203] dec_out[204] dec_out[205] dec_out[206] dec_out[207] dec_out[208] dec_out[209] dec_out[210] dec_out[211] dec_out[212] dec_out[213] dec_out[214] dec_out[215] dec_out[216] dec_out[217] dec_out[218] dec_out[219] dec_out[220] dec_out[221] dec_out[222] dec_out[223] dec_out[224] dec_out[225] dec_out[226] dec_out[227] dec_out[228] dec_out[229] dec_out[230] dec_out[231] dec_out[232] dec_out[233] dec_out[234] dec_out[235] dec_out[236] dec_out[237] dec_out[238] dec_out[239] dec_out[240] dec_out[241] dec_out[242] dec_out[243] dec_out[244] dec_out[245] dec_out[246] dec_out[247] dec_out[248] dec_out[249] dec_out[250] dec_out[251] dec_out[252] dec_out[253] dec_out[254] dec_out[255] dec_out[256] dec_out[257] dec_out[258] dec_out[259] dec_out[260] dec_out[261] dec_out[262] dec_out[263] dec_out[264] dec_out[265] dec_out[266] dec_out[267] dec_out[268] dec_out[269] dec_out[270] dec_out[271] dec_out[272] dec_out[273] dec_out[274] dec_out[275] dec_out[276] dec_out[277] dec_out[278] dec_out[279] dec_out[280] dec_out[281] dec_out[282] dec_out[283] dec_out[284] dec_out[285] dec_out[286] dec_out[287] dec_out[288] dec_out[289] dec_out[290] dec_out[291] dec_out[292] dec_out[293] dec_out[294] dec_out[295] dec_out[296] dec_out[297] dec_out[298] dec_out[299] dec_out[300] dec_out[301] dec_out[302] dec_out[303] dec_out[304] dec_out[305] dec_out[306] dec_out[307] dec_out[308] dec_out[309] dec_out[310] dec_out[311] dec_out[312] dec_out[313] dec_out[314] dec_out[315] dec_out[316] dec_out[317] dec_out[318] dec_out[319] dec_out[320] dec_out[321] dec_out[322] dec_out[323] dec_out[324] dec_out[325] dec_out[326] dec_out[327] dec_out[328] dec_out[329] dec_out[330] dec_out[331] dec_out[332] dec_out[333] dec_out[334] dec_out[335] dec_out[336] dec_out[337] dec_out[338] dec_out[339] dec_out[340] dec_out[341] dec_out[342] dec_out[343] dec_out[344] dec_out[345] dec_out[346] dec_out[347] dec_out[348] dec_out[349] dec_out[350] dec_out[351] dec_out[352] dec_out[353] dec_out[354] dec_out[355] dec_out[356] dec_out[357] dec_out[358] dec_out[359] dec_out[360] dec_out[361] dec_out[362] dec_out[363] dec_out[364] dec_out[365] dec_out[366] dec_out[367] dec_out[368] dec_out[369] dec_out[370] dec_out[371] dec_out[372] dec_out[373] dec_out[374] dec_out[375] dec_out[376] dec_out[377] dec_out[378] dec_out[379] dec_out[380] dec_out[381] dec_out[382] dec_out[383] dec_out[384] dec_out[385] dec_out[386] dec_out[387] dec_out[388] dec_out[389] dec_out[390] dec_out[391] dec_out[392] dec_out[393] dec_out[394] dec_out[395] dec_out[396] dec_out[397] dec_out[398] dec_out[399] dec_out[400] dec_out[401] dec_out[402] dec_out[403] dec_out[404] dec_out[405] dec_out[406] dec_out[407] dec_out[408] dec_out[409] dec_out[410] dec_out[411] dec_out[412] dec_out[413] dec_out[414] dec_out[415] dec_out[416] dec_out[417] dec_out[418] dec_out[419] dec_out[420] dec_out[421] dec_out[422] dec_out[423] dec_out[424] dec_out[425] dec_out[426] dec_out[427] dec_out[428] dec_out[429] dec_out[430] dec_out[431] dec_out[432] dec_out[433] dec_out[434] dec_out[435] dec_out[436] dec_out[437] dec_out[438] dec_out[439] dec_out[440] dec_out[441] dec_out[442] dec_out[443] dec_out[444] dec_out[445] dec_out[446] dec_out[447] dec_out[448] dec_out[449] dec_out[450] dec_out[451] dec_out[452] dec_out[453] dec_out[454] dec_out[455] dec_out[456] dec_out[457] dec_out[458] dec_out[459] dec_out[460] dec_out[461] dec_out[462] dec_out[463] dec_out[464] dec_out[465] dec_out[466] dec_out[467] dec_out[468] dec_out[469] dec_out[470] dec_out[471] dec_out[472] dec_out[473] dec_out[474] dec_out[475] dec_out[476] dec_out[477] dec_out[478] dec_out[479] dec_out[480] dec_out[481] dec_out[482] dec_out[483] dec_out[484] dec_out[485] dec_out[486] dec_out[487] dec_out[488] dec_out[489] dec_out[490] dec_out[491] dec_out[492] dec_out[493] dec_out[494] dec_out[495] dec_out[496] dec_out[497] dec_out[498] dec_out[499] dec_out[500] dec_out[501] dec_out[502] dec_out[503] dec_out[504] dec_out[505] dec_out[506] dec_out[507] dec_out[508] dec_out[509] dec_out[510] dec_out[511] wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] wl[128] wl[129] wl[130] wl[131] wl[132] wl[133] wl[134] wl[135] wl[136] wl[137] wl[138] wl[139] wl[140] wl[141] wl[142] wl[143] wl[144] wl[145] wl[146] wl[147] wl[148] wl[149] wl[150] wl[151] wl[152] wl[153] wl[154] wl[155] wl[156] wl[157] wl[158] wl[159] wl[160] wl[161] wl[162] wl[163] wl[164] wl[165] wl[166] wl[167] wl[168] wl[169] wl[170] wl[171] wl[172] wl[173] wl[174] wl[175] wl[176] wl[177] wl[178] wl[179] wl[180] wl[181] wl[182] wl[183] wl[184] wl[185] wl[186] wl[187] wl[188] wl[189] wl[190] wl[191] wl[192] wl[193] wl[194] wl[195] wl[196] wl[197] wl[198] wl[199] wl[200] wl[201] wl[202] wl[203] wl[204] wl[205] wl[206] wl[207] wl[208] wl[209] wl[210] wl[211] wl[212] wl[213] wl[214] wl[215] wl[216] wl[217] wl[218] wl[219] wl[220] wl[221] wl[222] wl[223] wl[224] wl[225] wl[226] wl[227] wl[228] wl[229] wl[230] wl[231] wl[232] wl[233] wl[234] wl[235] wl[236] wl[237] wl[238] wl[239] wl[240] wl[241] wl[242] wl[243] wl[244] wl[245] wl[246] wl[247] wl[248] wl[249] wl[250] wl[251] wl[252] wl[253] wl[254] wl[255] wl[256] wl[257] wl[258] wl[259] wl[260] wl[261] wl[262] wl[263] wl[264] wl[265] wl[266] wl[267] wl[268] wl[269] wl[270] wl[271] wl[272] wl[273] wl[274] wl[275] wl[276] wl[277] wl[278] wl[279] wl[280] wl[281] wl[282] wl[283] wl[284] wl[285] wl[286] wl[287] wl[288] wl[289] wl[290] wl[291] wl[292] wl[293] wl[294] wl[295] wl[296] wl[297] wl[298] wl[299] wl[300] wl[301] wl[302] wl[303] wl[304] wl[305] wl[306] wl[307] wl[308] wl[309] wl[310] wl[311] wl[312] wl[313] wl[314] wl[315] wl[316] wl[317] wl[318] wl[319] wl[320] wl[321] wl[322] wl[323] wl[324] wl[325] wl[326] wl[327] wl[328] wl[329] wl[330] wl[331] wl[332] wl[333] wl[334] wl[335] wl[336] wl[337] wl[338] wl[339] wl[340] wl[341] wl[342] wl[343] wl[344] wl[345] wl[346] wl[347] wl[348] wl[349] wl[350] wl[351] wl[352] wl[353] wl[354] wl[355] wl[356] wl[357] wl[358] wl[359] wl[360] wl[361] wl[362] wl[363] wl[364] wl[365] wl[366] wl[367] wl[368] wl[369] wl[370] wl[371] wl[372] wl[373] wl[374] wl[375] wl[376] wl[377] wl[378] wl[379] wl[380] wl[381] wl[382] wl[383] wl[384] wl[385] wl[386] wl[387] wl[388] wl[389] wl[390] wl[391] wl[392] wl[393] wl[394] wl[395] wl[396] wl[397] wl[398] wl[399] wl[400] wl[401] wl[402] wl[403] wl[404] wl[405] wl[406] wl[407] wl[408] wl[409] wl[410] wl[411] wl[412] wl[413] wl[414] wl[415] wl[416] wl[417] wl[418] wl[419] wl[420] wl[421] wl[422] wl[423] wl[424] wl[425] wl[426] wl[427] wl[428] wl[429] wl[430] wl[431] wl[432] wl[433] wl[434] wl[435] wl[436] wl[437] wl[438] wl[439] wl[440] wl[441] wl[442] wl[443] wl[444] wl[445] wl[446] wl[447] wl[448] wl[449] wl[450] wl[451] wl[452] wl[453] wl[454] wl[455] wl[456] wl[457] wl[458] wl[459] wl[460] wl[461] wl[462] wl[463] wl[464] wl[465] wl[466] wl[467] wl[468] wl[469] wl[470] wl[471] wl[472] wl[473] wl[474] wl[475] wl[476] wl[477] wl[478] wl[479] wl[480] wl[481] wl[482] wl[483] wl[484] wl[485] wl[486] wl[487] wl[488] wl[489] wl[490] wl[491] wl[492] wl[493] wl[494] wl[495] wl[496] wl[497] wl[498] wl[499] wl[500] wl[501] wl[502] wl[503] wl[504] wl[505] wl[506] wl[507] wl[508] wl[509] wl[510] wl[511] clk_buf vdd gnd wordline_driver
Xaddress_flop_array ADDR[0] ADDR[1] ADDR[2] ADDR[3] ADDR[4] ADDR[5] ADDR[6] ADDR[7] ADDR[8] ADDR[9] ADDR[10] A[0] A_bar[0] A[1] A_bar[1] A[2] A_bar[2] A[3] A_bar[3] A[4] A_bar[4] A[5] A_bar[5] A[6] A_bar[6] A[7] A_bar[7] A[8] A_bar[8] A[9] A_bar[9] A[10] A_bar[10] clk_buf vdd gnd msf_address
.ENDS bank

.SUBCKT sram_1rw_32b_2048w_1bank_freepdk45 DATA[0] DATA[1] DATA[2] DATA[3] DATA[4] DATA[5] DATA[6] DATA[7] DATA[8] DATA[9] DATA[10] DATA[11] DATA[12] DATA[13] DATA[14] DATA[15] DATA[16] DATA[17] DATA[18] DATA[19] DATA[20] DATA[21] DATA[22] DATA[23] DATA[24] DATA[25] DATA[26] DATA[27] DATA[28] DATA[29] DATA[30] DATA[31] ADDR[0] ADDR[1] ADDR[2] ADDR[3] ADDR[4] ADDR[5] ADDR[6] ADDR[7] ADDR[8] ADDR[9] ADDR[10] CSb WEb OEb clk vdd gnd
Xbank0 DATA[0] DATA[1] DATA[2] DATA[3] DATA[4] DATA[5] DATA[6] DATA[7] DATA[8] DATA[9] DATA[10] DATA[11] DATA[12] DATA[13] DATA[14] DATA[15] DATA[16] DATA[17] DATA[18] DATA[19] DATA[20] DATA[21] DATA[22] DATA[23] DATA[24] DATA[25] DATA[26] DATA[27] DATA[28] DATA[29] DATA[30] DATA[31] ADDR[0] ADDR[1] ADDR[2] ADDR[3] ADDR[4] ADDR[5] ADDR[6] ADDR[7] ADDR[8] ADDR[9] ADDR[10] s_en w_en tri_en_bar tri_en clk_bar clk_buf vdd gnd bank
Xcontrol CSb WEb OEb clk s_en w_en tri_en tri_en_bar clk_bar clk_buf vdd gnd control_logic
.ENDS sram_1rw_32b_2048w_1bank_freepdk45
