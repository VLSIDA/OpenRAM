magic
tech gf180mcuD
magscale 1 10
timestamp 1694553776
<< nwell >>
rect 675 -30 1355 650
<< nmos >>
rect 211 310 381 370
rect 211 200 381 260
<< pmos >>
rect 765 340 1106 400
rect 765 170 1106 230
<< ndiff >>
rect 211 448 381 470
rect 211 402 273 448
rect 319 402 381 448
rect 211 370 381 402
rect 211 260 381 310
rect 211 168 381 200
rect 211 122 273 168
rect 319 122 381 168
rect 211 100 381 122
<< pdiff >>
rect 765 478 1106 500
rect 765 432 818 478
rect 1052 432 1106 478
rect 765 400 1106 432
rect 765 308 1106 340
rect 765 262 818 308
rect 1052 262 1106 308
rect 765 230 1106 262
rect 765 138 1106 170
rect 765 92 818 138
rect 1052 92 1106 138
rect 765 70 1106 92
<< ndiffc >>
rect 273 402 319 448
rect 273 122 319 168
<< pdiffc >>
rect 818 432 1052 478
rect 818 262 1052 308
rect 818 92 1052 138
<< psubdiff >>
rect 74 33 181 50
rect 74 -13 114 33
rect 160 -13 181 33
rect 74 -30 181 -13
<< nsubdiff >>
rect 1172 117 1252 154
rect 1172 71 1189 117
rect 1235 71 1252 117
rect 1172 47 1252 71
<< psubdiffcont >>
rect 114 -13 160 33
<< nsubdiffcont >>
rect 1189 71 1235 117
<< polysilicon >>
rect 88 383 171 410
rect 88 337 104 383
rect 150 370 171 383
rect 431 370 765 400
rect 150 337 211 370
rect 88 310 211 337
rect 381 340 765 370
rect 1106 340 1156 400
rect 381 310 471 340
rect 88 244 211 260
rect 88 198 104 244
rect 150 200 211 244
rect 381 230 471 260
rect 381 200 765 230
rect 150 198 171 200
rect 88 160 171 198
rect 431 170 765 200
rect 1106 170 1156 230
<< polycontact >>
rect 104 337 150 383
rect 104 198 150 244
<< metal1 >>
rect 260 448 630 450
rect 101 383 153 435
rect 260 402 273 448
rect 319 402 630 448
rect 807 432 818 478
rect 1052 432 1064 478
rect 903 426 915 432
rect 967 426 979 432
rect 260 400 630 402
rect 101 337 104 383
rect 150 337 153 383
rect 101 323 153 337
rect 580 310 630 400
rect 580 308 1182 310
rect 580 262 818 308
rect 1052 262 1182 308
rect 580 260 1182 262
rect 101 244 153 258
rect 101 198 104 244
rect 150 198 153 244
rect 101 139 153 198
rect 241 116 273 168
rect 325 116 348 168
rect 903 138 915 144
rect 967 138 979 144
rect 241 110 348 116
rect 807 92 818 138
rect 1052 92 1064 138
rect 1139 68 1186 120
rect 1238 68 1250 120
rect 80 36 179 46
rect 80 -16 111 36
rect 163 -16 179 36
rect 80 -24 179 -16
<< via1 >>
rect 915 432 967 478
rect 915 426 967 432
rect 273 122 319 168
rect 319 122 325 168
rect 273 116 325 122
rect 915 138 967 144
rect 915 92 967 138
rect 1186 117 1238 120
rect 1186 71 1189 117
rect 1189 71 1235 117
rect 1235 71 1238 117
rect 1186 68 1238 71
rect 111 33 163 36
rect 111 -13 114 33
rect 114 -13 160 33
rect 160 -13 163 33
rect 111 -16 163 -13
<< metal2 >>
rect 271 168 327 530
rect 271 116 273 168
rect 325 116 327 168
rect 271 38 327 116
rect 89 36 327 38
rect 89 -16 111 36
rect 163 -16 327 36
rect 913 478 969 530
rect 913 426 915 478
rect 967 426 969 478
rect 913 144 969 426
rect 913 92 915 144
rect 967 122 969 144
rect 967 120 1250 122
rect 967 92 1186 120
rect 913 68 1186 92
rect 1238 68 1250 120
rect 913 66 1250 68
rect 913 18 969 66
rect 89 -18 327 -16
<< labels >>
rlabel metal2 s 271 38 327 530 4 GND
port 1 nsew
rlabel metal2 s 941 43 941 43 4 VDD
flabel metal1 s 605 425 605 425 2 FreeSans 368 0 0 0 Z
port 2 nsew
flabel metal1 s 127 360 127 360 2 FreeSans 368 0 0 0 A
port 3 nsew
flabel metal1 s 127 221 127 221 2 FreeSans 368 0 0 0 B
port 4 nsew
<< properties >>
string FIXED_BBOX -17 0 1373 542
<< end >>
