magic
tech gf180mcuD
magscale 1 10
timestamp 1694482220
<< nwell >>
rect 620 -40 1300 580
<< nmos >>
rect 156 300 326 360
rect 156 190 326 250
<< pmos >>
rect 710 330 1051 390
rect 710 160 1051 220
<< ndiff >>
rect 156 438 326 460
rect 156 392 218 438
rect 264 392 326 438
rect 156 360 326 392
rect 156 250 326 300
rect 156 158 326 190
rect 156 112 218 158
rect 264 112 326 158
rect 156 90 326 112
<< pdiff >>
rect 710 468 1051 490
rect 710 422 763 468
rect 997 422 1051 468
rect 710 390 1051 422
rect 710 298 1051 330
rect 710 252 763 298
rect 997 252 1051 298
rect 710 220 1051 252
rect 710 128 1051 160
rect 710 82 763 128
rect 997 82 1051 128
rect 710 60 1051 82
<< ndiffc >>
rect 218 392 264 438
rect 218 112 264 158
<< pdiffc >>
rect 763 422 997 468
rect 763 252 997 298
rect 763 82 997 128
<< psubdiff >>
rect 19 23 126 40
rect 19 -23 59 23
rect 105 -23 126 23
rect 19 -40 126 -23
<< nsubdiff >>
rect 1117 107 1197 144
rect 1117 61 1134 107
rect 1180 61 1197 107
rect 1117 37 1197 61
<< psubdiffcont >>
rect 59 -23 105 23
<< nsubdiffcont >>
rect 1134 61 1180 107
<< polysilicon >>
rect 33 373 116 400
rect 33 327 49 373
rect 95 360 116 373
rect 376 360 710 390
rect 95 327 156 360
rect 33 300 156 327
rect 326 330 710 360
rect 1051 330 1101 390
rect 326 300 416 330
rect 33 234 156 250
rect 33 188 49 234
rect 95 190 156 234
rect 326 220 416 250
rect 326 190 710 220
rect 95 188 116 190
rect 33 150 116 188
rect 376 160 710 190
rect 1051 160 1101 220
<< polycontact >>
rect 49 327 95 373
rect 49 188 95 234
<< metal1 >>
rect 156 438 396 440
rect 46 373 98 425
rect 156 392 218 438
rect 264 392 396 438
rect 752 422 763 468
rect 997 422 1009 468
rect 848 416 860 422
rect 912 416 924 422
rect 156 390 396 392
rect 46 327 49 373
rect 95 327 98 373
rect 46 313 98 327
rect 346 300 396 390
rect 1075 300 1127 463
rect 346 298 1127 300
rect 346 252 763 298
rect 997 252 1127 298
rect 346 250 1127 252
rect 46 234 98 248
rect 46 188 49 234
rect 95 188 98 234
rect 46 129 98 188
rect 186 106 218 158
rect 270 106 293 158
rect 848 128 860 134
rect 912 128 924 134
rect 186 100 293 106
rect 752 82 763 128
rect 997 82 1009 128
rect 1084 58 1131 110
rect 1183 58 1195 110
rect 25 26 124 36
rect 25 -26 56 26
rect 108 -26 124 26
rect 25 -34 124 -26
<< via1 >>
rect 860 422 912 468
rect 860 416 912 422
rect 218 112 264 158
rect 264 112 270 158
rect 218 106 270 112
rect 860 128 912 134
rect 860 82 912 128
rect 1131 107 1183 110
rect 1131 61 1134 107
rect 1134 61 1180 107
rect 1180 61 1183 107
rect 1131 58 1183 61
rect 56 23 108 26
rect 56 -23 59 23
rect 59 -23 105 23
rect 105 -23 108 23
rect 56 -26 108 -23
<< metal2 >>
rect 216 158 272 520
rect 216 106 218 158
rect 270 106 272 158
rect 216 28 272 106
rect 34 26 272 28
rect 34 -26 56 26
rect 108 -26 272 26
rect 858 468 914 520
rect 858 416 860 468
rect 912 416 914 468
rect 858 134 914 416
rect 858 82 860 134
rect 912 112 914 134
rect 912 110 1195 112
rect 912 82 1131 110
rect 858 58 1131 82
rect 1183 58 1195 110
rect 858 56 1195 58
rect 858 8 914 56
rect 34 -28 272 -26
<< labels >>
rlabel metal1 s 73 350 73 350 4 B
rlabel metal1 s 73 211 73 211 4 A
rlabel metal1 s 1101 439 1101 439 4 Y
rlabel metal2 s 886 33 886 33 4 VDD
rlabel metal2 s 245 56 245 56 4 GND
<< properties >>
string FIXED_BBOX 0 0 1300 522
<< end >>
