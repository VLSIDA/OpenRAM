magic
tech sky130A
magscale 1 2
timestamp 1595931502
<< checkpaint >>
rect -1309 -1311 6706 22869
<< locali >>
rect 3974 11295 5362 11329
rect 3388 9881 5362 9915
rect 3388 8467 5362 8501
rect 3552 7350 3586 7832
rect 3367 7316 3586 7350
rect 4114 7053 5362 7087
rect 4406 5639 5362 5673
rect 4414 4225 5362 4259
rect 4414 2811 5362 2845
rect 3349 2541 3534 2575
rect 3349 2176 3383 2541
rect 3216 2142 3383 2176
rect 4782 1397 5362 1431
<< metal1 >>
rect 5330 11286 5394 11338
rect 2362 11028 3116 11056
rect 2446 10904 3249 10932
rect 2698 10780 3382 10808
rect 3666 10605 3730 10657
rect 5330 9872 5394 9924
rect 2362 9139 3101 9167
rect 3184 9127 3248 9179
rect 5330 8458 5394 8510
rect 2530 8200 3149 8228
rect 2362 7952 3249 7980
rect 4020 7789 4084 7841
rect 203 7039 2362 7067
rect 5330 7044 5394 7096
rect 3882 6337 3946 6389
rect 2446 6160 3382 6188
rect 2278 6036 3249 6064
rect 2614 5912 3116 5940
rect 5330 5630 5394 5682
rect 2446 4973 3101 5001
rect 4286 4923 4350 4975
rect 383 4228 2782 4256
rect 5330 4216 5394 4268
rect 3888 3493 3952 3545
rect 2866 3332 3249 3360
rect 2782 3084 3149 3112
rect 5330 2802 5394 2854
rect 3585 2284 3649 2336
rect 2782 2145 3101 2173
rect 4256 2111 4320 2163
rect 5330 1388 5394 1440
rect 3069 643 3133 695
rect 4832 681 4896 733
rect 5330 -26 5394 26
<< metal2 >>
rect 1748 11472 1776 11994
rect 189 7053 217 11472
rect 369 2828 397 4242
rect 137 2238 203 2290
rect 137 538 203 590
rect 2264 0 2292 11388
rect 2348 0 2376 11388
rect 2432 0 2460 11388
rect 2516 0 2544 11388
rect 2600 0 2628 11388
rect 2684 0 2712 11388
rect 2768 0 2796 11388
rect 2852 0 2880 11388
rect 5334 11288 5390 11336
rect 3698 10617 5446 10645
rect 5334 9874 5390 9922
rect 3202 8587 3230 9153
rect 5334 8460 5390 8508
rect 4052 7801 5446 7829
rect 5334 7046 5390 7094
rect 3914 6349 5446 6377
rect 5334 5632 5390 5680
rect 4318 4935 5446 4963
rect 5334 4218 5390 4266
rect 3892 3495 3948 3543
rect 5334 2804 5390 2852
rect 3589 2286 3645 2334
rect 4274 1571 4302 2137
rect 5334 1390 5390 1438
rect 4864 707 5446 721
rect 4850 693 5446 707
rect 3087 655 3115 683
rect 4850 141 4878 693
rect 5334 -24 5390 24
<< metal3 >>
rect 399 21503 497 21601
rect 1135 21503 1233 21601
rect 399 20383 497 20481
rect 1135 20383 1233 20481
rect 399 19263 497 19361
rect 1135 19263 1233 19361
rect 399 18143 497 18241
rect 1135 18143 1233 18241
rect 399 17023 497 17121
rect 1135 17023 1233 17121
rect 399 15903 497 16001
rect 1135 15903 1233 16001
rect 399 14783 497 14881
rect 1135 14783 1233 14881
rect 399 13663 497 13761
rect 1135 13663 1233 13761
rect 399 12543 497 12641
rect 1135 12543 1233 12641
rect 399 11423 497 11521
rect 1135 11423 1233 11521
rect 5313 11263 5411 11361
rect 5313 9849 5411 9947
rect 2278 8557 3216 8617
rect 5313 8435 5411 8533
rect 5313 7021 5411 7119
rect 5313 5607 5411 5705
rect 5313 4193 5411 4291
rect 2530 3489 3920 3549
rect -49 2781 49 2879
rect 5313 2779 5411 2877
rect 2088 2295 2698 2355
rect 2866 2280 3617 2340
rect 1582 1913 2614 1973
rect 2446 1541 4288 1601
rect -49 1365 49 1463
rect 5313 1365 5411 1463
rect 1582 855 2866 915
rect 2782 111 4864 171
rect -49 -51 49 47
rect 5313 -49 5411 49
use pand3_0  pand3_0_0
timestamp 1595931502
transform 1 0 3020 0 -1 11312
box -36 -17 990 1471
use pdriver_4  pdriver_4_0
timestamp 1595931502
transform 1 0 3488 0 -1 8484
box -36 -17 662 1471
use contact_9  contact_9_21
timestamp 1595931502
transform 1 0 1549 0 1 848
box 0 0 66 74
use contact_9  contact_9_20
timestamp 1595931502
transform 1 0 1549 0 1 1906
box 0 0 66 74
use contact_9  contact_9_19
timestamp 1595931502
transform 1 0 2055 0 1 2288
box 0 0 66 74
use contact_9  contact_9_18
timestamp 1595931502
transform 1 0 3584 0 1 2273
box 0 0 66 74
use contact_9  contact_9_17
timestamp 1595931502
transform 1 0 3584 0 1 2273
box 0 0 66 74
use contact_9  contact_9_16
timestamp 1595931502
transform 1 0 3887 0 1 3482
box 0 0 66 74
use contact_9  contact_9_15
timestamp 1595931502
transform 1 0 5329 0 1 1377
box 0 0 66 74
use contact_9  contact_9_14
timestamp 1595931502
transform 1 0 5329 0 1 -37
box 0 0 66 74
use contact_9  contact_9_13
timestamp 1595931502
transform 1 0 5329 0 1 1377
box 0 0 66 74
use contact_9  contact_9_12
timestamp 1595931502
transform 1 0 5329 0 1 2791
box 0 0 66 74
use contact_9  contact_9_11
timestamp 1595931502
transform 1 0 5329 0 1 4205
box 0 0 66 74
use contact_9  contact_9_10
timestamp 1595931502
transform 1 0 5329 0 1 2791
box 0 0 66 74
use contact_9  contact_9_9
timestamp 1595931502
transform 1 0 5329 0 1 4205
box 0 0 66 74
use contact_9  contact_9_8
timestamp 1595931502
transform 1 0 5329 0 1 5619
box 0 0 66 74
use contact_9  contact_9_7
timestamp 1595931502
transform 1 0 5329 0 1 7033
box 0 0 66 74
use contact_9  contact_9_6
timestamp 1595931502
transform 1 0 5329 0 1 5619
box 0 0 66 74
use contact_9  contact_9_5
timestamp 1595931502
transform 1 0 5329 0 1 7033
box 0 0 66 74
use contact_9  contact_9_4
timestamp 1595931502
transform 1 0 5329 0 1 8447
box 0 0 66 74
use contact_9  contact_9_3
timestamp 1595931502
transform 1 0 5329 0 1 9861
box 0 0 66 74
use contact_9  contact_9_2
timestamp 1595931502
transform 1 0 5329 0 1 8447
box 0 0 66 74
use contact_9  contact_9_1
timestamp 1595931502
transform 1 0 5329 0 1 9861
box 0 0 66 74
use contact_9  contact_9_0
timestamp 1595931502
transform 1 0 5329 0 1 11275
box 0 0 66 74
use pdriver_1  pdriver_1_0
timestamp 1595931502
transform 1 0 3020 0 -1 5656
box -36 -17 1508 1471
use pand2  pand2_1
timestamp 1595931502
transform 1 0 3388 0 -1 2828
box -36 -17 1430 1471
use pand2  pand2_0
timestamp 1595931502
transform 1 0 3020 0 1 2828
box -36 -17 1430 1471
use delay_chain  delay_chain_0
timestamp 1595931502
transform -1 0 1840 0 1 11472
box -36 -49 1876 10137
use contact_8  contact_8_0
timestamp 1595931502
transform 1 0 5330 0 1 11280
box 0 0 64 64
use contact_7  contact_7_0
timestamp 1595931502
transform 1 0 5333 0 1 11279
box 0 0 58 66
use contact_8  contact_8_1
timestamp 1595931502
transform 1 0 5330 0 1 9866
box 0 0 64 64
use contact_7  contact_7_1
timestamp 1595931502
transform 1 0 5333 0 1 9865
box 0 0 58 66
use contact_8  contact_8_2
timestamp 1595931502
transform 1 0 5330 0 1 8452
box 0 0 64 64
use contact_7  contact_7_2
timestamp 1595931502
transform 1 0 5333 0 1 8451
box 0 0 58 66
use contact_8  contact_8_3
timestamp 1595931502
transform 1 0 5330 0 1 9866
box 0 0 64 64
use contact_7  contact_7_3
timestamp 1595931502
transform 1 0 5333 0 1 9865
box 0 0 58 66
use contact_8  contact_8_4
timestamp 1595931502
transform 1 0 5330 0 1 8452
box 0 0 64 64
use contact_7  contact_7_4
timestamp 1595931502
transform 1 0 5333 0 1 8451
box 0 0 58 66
use contact_8  contact_8_5
timestamp 1595931502
transform 1 0 5330 0 1 7038
box 0 0 64 64
use contact_7  contact_7_5
timestamp 1595931502
transform 1 0 5333 0 1 7037
box 0 0 58 66
use contact_8  contact_8_6
timestamp 1595931502
transform 1 0 5330 0 1 5624
box 0 0 64 64
use contact_7  contact_7_6
timestamp 1595931502
transform 1 0 5333 0 1 5623
box 0 0 58 66
use contact_8  contact_8_7
timestamp 1595931502
transform 1 0 5330 0 1 7038
box 0 0 64 64
use contact_7  contact_7_7
timestamp 1595931502
transform 1 0 5333 0 1 7037
box 0 0 58 66
use contact_8  contact_8_8
timestamp 1595931502
transform 1 0 5330 0 1 5624
box 0 0 64 64
use contact_7  contact_7_8
timestamp 1595931502
transform 1 0 5333 0 1 5623
box 0 0 58 66
use contact_8  contact_8_9
timestamp 1595931502
transform 1 0 5330 0 1 4210
box 0 0 64 64
use contact_7  contact_7_9
timestamp 1595931502
transform 1 0 5333 0 1 4209
box 0 0 58 66
use contact_8  contact_8_10
timestamp 1595931502
transform 1 0 5330 0 1 2796
box 0 0 64 64
use contact_7  contact_7_10
timestamp 1595931502
transform 1 0 5333 0 1 2795
box 0 0 58 66
use contact_8  contact_8_11
timestamp 1595931502
transform 1 0 5330 0 1 4210
box 0 0 64 64
use contact_7  contact_7_11
timestamp 1595931502
transform 1 0 5333 0 1 4209
box 0 0 58 66
use contact_8  contact_8_12
timestamp 1595931502
transform 1 0 5330 0 1 2796
box 0 0 64 64
use contact_7  contact_7_12
timestamp 1595931502
transform 1 0 5333 0 1 2795
box 0 0 58 66
use contact_8  contact_8_13
timestamp 1595931502
transform 1 0 5330 0 1 1382
box 0 0 64 64
use contact_7  contact_7_13
timestamp 1595931502
transform 1 0 5333 0 1 1381
box 0 0 58 66
use contact_8  contact_8_14
timestamp 1595931502
transform 1 0 5330 0 1 -32
box 0 0 64 64
use contact_7  contact_7_14
timestamp 1595931502
transform 1 0 5333 0 1 -33
box 0 0 58 66
use contact_8  contact_8_15
timestamp 1595931502
transform 1 0 5330 0 1 1382
box 0 0 64 64
use contact_7  contact_7_15
timestamp 1595931502
transform 1 0 5333 0 1 1381
box 0 0 58 66
use contact_8  contact_8_16
timestamp 1595931502
transform 1 0 3888 0 1 3487
box 0 0 64 64
use contact_7  contact_7_16
timestamp 1595931502
transform 1 0 3891 0 1 3486
box 0 0 58 66
use contact_8  contact_8_17
timestamp 1595931502
transform 1 0 3888 0 1 3487
box 0 0 64 64
use contact_7  contact_7_17
timestamp 1595931502
transform 1 0 3891 0 1 3486
box 0 0 58 66
use contact_27  contact_27_0
timestamp 1595931502
transform 1 0 2497 0 1 3482
box 0 0 66 74
use contact_7  contact_7_18
timestamp 1595931502
transform 1 0 3220 0 1 3313
box 0 0 58 66
use contact_8  contact_8_18
timestamp 1595931502
transform 1 0 2834 0 1 3314
box 0 0 64 64
use contact_7  contact_7_19
timestamp 1595931502
transform 1 0 3120 0 1 3065
box 0 0 58 66
use contact_8  contact_8_19
timestamp 1595931502
transform 1 0 2750 0 1 3066
box 0 0 64 64
use contact_8  contact_8_20
timestamp 1595931502
transform 1 0 4256 0 1 2105
box 0 0 64 64
use contact_7  contact_7_20
timestamp 1595931502
transform 1 0 4259 0 1 2104
box 0 0 58 66
use contact_27  contact_27_1
timestamp 1595931502
transform 1 0 2413 0 1 1534
box 0 0 66 74
use contact_27  contact_27_2
timestamp 1595931502
transform 1 0 4255 0 1 1534
box 0 0 66 74
use contact_8  contact_8_21
timestamp 1595931502
transform 1 0 3585 0 1 2278
box 0 0 64 64
use contact_7  contact_7_21
timestamp 1595931502
transform 1 0 3588 0 1 2277
box 0 0 58 66
use contact_8  contact_8_22
timestamp 1595931502
transform 1 0 3585 0 1 2278
box 0 0 64 64
use contact_7  contact_7_22
timestamp 1595931502
transform 1 0 3588 0 1 2277
box 0 0 58 66
use contact_27  contact_27_3
timestamp 1595931502
transform 1 0 2833 0 1 2273
box 0 0 66 74
use contact_7  contact_7_23
timestamp 1595931502
transform 1 0 3072 0 1 2126
box 0 0 58 66
use contact_8  contact_8_23
timestamp 1595931502
transform 1 0 2750 0 1 2127
box 0 0 64 64
use contact_8  contact_8_24
timestamp 1595931502
transform 1 0 4832 0 1 675
box 0 0 64 64
use contact_7  contact_7_24
timestamp 1595931502
transform 1 0 4835 0 1 674
box 0 0 58 66
use contact_8  contact_8_25
timestamp 1595931502
transform 1 0 4832 0 1 675
box 0 0 64 64
use contact_7  contact_7_25
timestamp 1595931502
transform 1 0 4835 0 1 674
box 0 0 58 66
use contact_27  contact_27_4
timestamp 1595931502
transform 1 0 2749 0 1 104
box 0 0 66 74
use contact_27  contact_27_5
timestamp 1595931502
transform 1 0 4831 0 1 104
box 0 0 66 74
use contact_8  contact_8_26
timestamp 1595931502
transform 1 0 3069 0 1 637
box 0 0 64 64
use contact_7  contact_7_26
timestamp 1595931502
transform 1 0 3072 0 1 636
box 0 0 58 66
use contact_8  contact_8_27
timestamp 1595931502
transform 1 0 4020 0 1 7783
box 0 0 64 64
use contact_7  contact_7_27
timestamp 1595931502
transform 1 0 4023 0 1 7782
box 0 0 58 66
use contact_7  contact_7_28
timestamp 1595931502
transform 1 0 3220 0 1 7933
box 0 0 58 66
use contact_8  contact_8_28
timestamp 1595931502
transform 1 0 2330 0 1 7934
box 0 0 64 64
use contact_7  contact_7_29
timestamp 1595931502
transform 1 0 3120 0 1 8181
box 0 0 58 66
use contact_8  contact_8_29
timestamp 1595931502
transform 1 0 2498 0 1 8182
box 0 0 64 64
use contact_8  contact_8_30
timestamp 1595931502
transform 1 0 2330 0 1 7021
box 0 0 64 64
use contact_8  contact_8_31
timestamp 1595931502
transform 1 0 171 0 1 7021
box 0 0 64 64
use contact_8  contact_8_32
timestamp 1595931502
transform 1 0 3666 0 1 10599
box 0 0 64 64
use contact_7  contact_7_30
timestamp 1595931502
transform 1 0 3669 0 1 10598
box 0 0 58 66
use contact_7  contact_7_31
timestamp 1595931502
transform 1 0 3353 0 1 10761
box 0 0 58 66
use contact_8  contact_8_33
timestamp 1595931502
transform 1 0 2666 0 1 10762
box 0 0 64 64
use contact_7  contact_7_32
timestamp 1595931502
transform 1 0 3220 0 1 10885
box 0 0 58 66
use contact_8  contact_8_34
timestamp 1595931502
transform 1 0 2414 0 1 10886
box 0 0 64 64
use contact_7  contact_7_33
timestamp 1595931502
transform 1 0 3087 0 1 11009
box 0 0 58 66
use contact_8  contact_8_35
timestamp 1595931502
transform 1 0 2330 0 1 11010
box 0 0 64 64
use contact_8  contact_8_36
timestamp 1595931502
transform 1 0 3882 0 1 6331
box 0 0 64 64
use contact_7  contact_7_34
timestamp 1595931502
transform 1 0 3885 0 1 6330
box 0 0 58 66
use contact_7  contact_7_35
timestamp 1595931502
transform 1 0 3353 0 1 6141
box 0 0 58 66
use contact_8  contact_8_37
timestamp 1595931502
transform 1 0 2414 0 1 6142
box 0 0 64 64
use contact_7  contact_7_36
timestamp 1595931502
transform 1 0 3220 0 1 6017
box 0 0 58 66
use contact_8  contact_8_38
timestamp 1595931502
transform 1 0 2246 0 1 6018
box 0 0 64 64
use contact_7  contact_7_37
timestamp 1595931502
transform 1 0 3087 0 1 5893
box 0 0 58 66
use contact_8  contact_8_39
timestamp 1595931502
transform 1 0 2582 0 1 5894
box 0 0 64 64
use contact_7  contact_7_38
timestamp 1595931502
transform 1 0 3072 0 1 9120
box 0 0 58 66
use contact_8  contact_8_40
timestamp 1595931502
transform 1 0 2330 0 1 9121
box 0 0 64 64
use contact_8  contact_8_41
timestamp 1595931502
transform 1 0 3184 0 1 9121
box 0 0 64 64
use contact_7  contact_7_39
timestamp 1595931502
transform 1 0 3187 0 1 9120
box 0 0 58 66
use contact_27  contact_27_6
timestamp 1595931502
transform 1 0 2245 0 1 8550
box 0 0 66 74
use contact_27  contact_27_7
timestamp 1595931502
transform 1 0 3183 0 1 8550
box 0 0 66 74
use contact_8  contact_8_42
timestamp 1595931502
transform 1 0 4286 0 1 4917
box 0 0 64 64
use contact_7  contact_7_40
timestamp 1595931502
transform 1 0 4289 0 1 4916
box 0 0 58 66
use contact_7  contact_7_41
timestamp 1595931502
transform 1 0 3072 0 1 4954
box 0 0 58 66
use contact_8  contact_8_43
timestamp 1595931502
transform 1 0 2414 0 1 4955
box 0 0 64 64
use contact_8  contact_8_44
timestamp 1595931502
transform 1 0 2750 0 1 4210
box 0 0 64 64
use contact_8  contact_8_45
timestamp 1595931502
transform 1 0 351 0 1 4210
box 0 0 64 64
use contact_27  contact_27_8
timestamp 1595931502
transform 1 0 2665 0 1 2288
box 0 0 66 74
use contact_27  contact_27_9
timestamp 1595931502
transform 1 0 2581 0 1 1906
box 0 0 66 74
use contact_27  contact_27_10
timestamp 1595931502
transform 1 0 2833 0 1 848
box 0 0 66 74
use pnand2_0  pnand2_0_0
timestamp 1595931502
transform 1 0 3020 0 -1 8484
box -36 -17 504 1471
use pand3  pand3_0
timestamp 1595931502
transform 1 0 3020 0 1 5656
box -36 -17 1422 1471
use pinv_2  pinv_2_0
timestamp 1595931502
transform 1 0 3020 0 1 8484
box -36 -17 404 1471
use pinv_2  pinv_2_1
timestamp 1595931502
transform 1 0 3020 0 -1 2828
box -36 -17 404 1471
use pdriver_0  pdriver_0_0
timestamp 1595931502
transform 1 0 3020 0 1 0
box -36 -17 2378 1471
use dff_buf_array  dff_buf_array_0
timestamp 1595931502
transform 1 0 0 0 1 0
box -49 -51 2300 2879
<< labels >>
rlabel metal2 s 5155 707 5155 707 4 clk_buf
rlabel metal3 s 1184 15952 1184 15952 4 gnd
rlabel metal3 s 5362 0 5362 0 4 gnd
rlabel metal3 s 1184 11472 1184 11472 4 gnd
rlabel metal3 s 5362 5656 5362 5656 4 gnd
rlabel metal3 s 5362 2828 5362 2828 4 gnd
rlabel metal3 s 448 15952 448 15952 4 gnd
rlabel metal3 s 448 18192 448 18192 4 gnd
rlabel metal3 s 448 20432 448 20432 4 gnd
rlabel metal3 s 0 2830 0 2830 4 gnd
rlabel metal3 s 0 -2 0 -2 4 gnd
rlabel metal3 s 5362 8484 5362 8484 4 gnd
rlabel metal3 s 1184 20432 1184 20432 4 gnd
rlabel metal3 s 448 11472 448 11472 4 gnd
rlabel metal3 s 1184 18192 1184 18192 4 gnd
rlabel metal3 s 1184 13712 1184 13712 4 gnd
rlabel metal3 s 5362 11312 5362 11312 4 gnd
rlabel metal3 s 448 13712 448 13712 4 gnd
rlabel metal2 s 170 564 170 564 4 csb
rlabel metal2 s 4882 4949 4882 4949 4 wl_en
rlabel metal2 s 1762 11733 1762 11733 4 rbl_bl
rlabel metal2 s 3101 669 3101 669 4 clk
rlabel metal2 s 170 2264 170 2264 4 web
rlabel metal2 s 4749 7815 4749 7815 4 p_en_bar
rlabel metal2 s 4572 10631 4572 10631 4 s_en
rlabel metal3 s 1184 14832 1184 14832 4 vdd
rlabel metal3 s 5362 4242 5362 4242 4 vdd
rlabel metal3 s 5362 1414 5362 1414 4 vdd
rlabel metal3 s 0 1414 0 1414 4 vdd
rlabel metal3 s 448 12592 448 12592 4 vdd
rlabel metal3 s 448 17072 448 17072 4 vdd
rlabel metal3 s 448 14832 448 14832 4 vdd
rlabel metal3 s 1184 17072 1184 17072 4 vdd
rlabel metal3 s 1184 19312 1184 19312 4 vdd
rlabel metal3 s 448 21552 448 21552 4 vdd
rlabel metal3 s 448 19312 448 19312 4 vdd
rlabel metal3 s 1184 21552 1184 21552 4 vdd
rlabel metal3 s 5362 9898 5362 9898 4 vdd
rlabel metal3 s 1184 12592 1184 12592 4 vdd
rlabel metal3 s 5362 7070 5362 7070 4 vdd
rlabel metal2 s 4680 6363 4680 6363 4 w_en
<< properties >>
string FIXED_BBOX 0 0 5446 21712
<< end >>
