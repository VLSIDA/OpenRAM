VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_2_16_sky130
   CLASS BLOCK ;
   SIZE 151.29 BY 140.08 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  33.755 2.69 34.085 2.95 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  39.595 2.69 39.925 2.95 ;
      END
   END din0[1]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  22.075 111.25 22.405 111.51 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  22.075 119.75 22.405 120.01 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  22.075 125.39 22.405 125.65 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  22.075 133.89 22.405 134.15 ;
      END
   END addr0[3]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  130.415 42.71 130.745 42.97 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  130.415 34.21 130.745 34.47 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  130.415 28.57 130.745 28.83 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  130.415 20.07 130.745 20.33 ;
      END
   END addr1[3]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  0.685 2.69 1.015 2.95 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  150.275 137.13 150.605 137.39 ;
      END
   END csb1
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  0.685 11.19 1.015 11.45 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  15.435 3.275 15.575 3.415 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER m2 ;
         RECT  136.135 136.665 136.275 136.805 ;
      END
   END clk1
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER m1 ;
         RECT  73.6 39.79 73.83 41.06 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER m1 ;
         RECT  77.95 39.79 78.18 41.06 ;
      END
   END dout0[1]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER m1 ;
         RECT  73.6 113.16 73.83 114.43 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER m1 ;
         RECT  77.95 113.16 78.18 114.43 ;
      END
   END dout1[1]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER m3 ;
         RECT  77.075 29.185 77.565 29.675 ;
         LAYER m3 ;
         RECT  74.215 29.185 74.705 29.675 ;
         LAYER m3 ;
         RECT  76.61 45.885 77.1 46.375 ;
         LAYER m3 ;
         RECT  54.545 90.835 55.035 91.325 ;
         LAYER m3 ;
         RECT  125.765 132.765 126.255 133.255 ;
         LAYER m3 ;
         RECT  40.22 63.22 40.71 63.71 ;
         LAYER m3 ;
         RECT  118.305 75.035 118.795 75.525 ;
         LAYER m3 ;
         RECT  77.61 95.565 77.91 95.865 ;
         LAYER m3 ;
         RECT  74.115 33.935 74.605 34.425 ;
         LAYER m3 ;
         RECT  111.69 75.07 112.18 75.56 ;
         LAYER m3 ;
         RECT  148.805 46.215 149.295 46.705 ;
         LAYER m3 ;
         RECT  74.74 112.035 75.23 112.525 ;
         LAYER m3 ;
         RECT  1.995 62.715 2.485 63.205 ;
         LAYER m3 ;
         RECT  148.805 91.015 149.295 91.505 ;
         LAYER m3 ;
         RECT  71.275 95.47 71.765 95.96 ;
         LAYER m3 ;
         RECT  5.675 62.715 6.165 63.205 ;
         LAYER m3 ;
         RECT  71.275 58.26 71.765 58.75 ;
         LAYER m3 ;
         RECT  78.11 98.425 78.6 98.915 ;
         LAYER m3 ;
         RECT  111.69 63.22 112.18 63.71 ;
         LAYER m3 ;
         RECT  40.22 75.07 40.71 75.56 ;
         LAYER m3 ;
         RECT  100.62 75.07 101.11 75.56 ;
         LAYER m3 ;
         RECT  100.62 73.22 101.11 73.71 ;
         LAYER m3 ;
         RECT  1.995 96.315 2.485 96.805 ;
         LAYER m3 ;
         RECT  5.675 96.315 6.165 96.805 ;
         LAYER m3 ;
         RECT  24.065 115.385 24.555 115.875 ;
         LAYER m3 ;
         RECT  78.11 55.305 78.6 55.795 ;
         LAYER m3 ;
         RECT  97.365 84.91 97.855 85.4 ;
         LAYER m3 ;
         RECT  35.745 6.825 36.235 7.315 ;
         LAYER m3 ;
         RECT  100.62 85.07 101.11 85.56 ;
         LAYER m3 ;
         RECT  76.55 41.695 77.04 42.185 ;
         LAYER m3 ;
         RECT  71.87 55.305 72.36 55.795 ;
         LAYER m3 ;
         RECT  54.545 73.06 55.035 73.55 ;
         LAYER m3 ;
         RECT  63.475 76.865 63.965 77.355 ;
         LAYER m3 ;
         RECT  51.29 71.12 51.78 71.61 ;
         LAYER m3 ;
         RECT  97.365 67.135 97.855 67.625 ;
         LAYER m3 ;
         RECT  100.62 67.17 101.11 67.66 ;
         LAYER m3 ;
         RECT  51.29 85.07 51.78 85.56 ;
         LAYER m3 ;
         RECT  100.62 77.17 101.11 77.66 ;
         LAYER m3 ;
         RECT  54.545 67.135 55.035 67.625 ;
         LAYER m3 ;
         RECT  1.995 73.915 2.485 74.405 ;
         LAYER m3 ;
         RECT  145.125 46.215 145.615 46.705 ;
         LAYER m3 ;
         RECT  93.01 76.785 93.5 77.275 ;
         LAYER m3 ;
         RECT  100.62 82.97 101.11 83.46 ;
         LAYER m3 ;
         RECT  100.62 65.32 101.11 65.81 ;
         LAYER m3 ;
         RECT  1.995 85.115 2.485 85.605 ;
         LAYER m3 ;
         RECT  97.365 71.085 97.855 71.575 ;
         LAYER m3 ;
         RECT  54.545 65.16 55.035 65.65 ;
         LAYER m3 ;
         RECT  111.69 67.17 112.18 67.66 ;
         LAYER m3 ;
         RECT  54.545 78.985 55.035 79.475 ;
         LAYER m3 ;
         RECT  97.365 86.885 97.855 87.375 ;
         LAYER m3 ;
         RECT  54.545 82.935 55.035 83.425 ;
         LAYER m3 ;
         RECT  33.605 75.035 34.095 75.525 ;
         LAYER m3 ;
         RECT  97.365 63.185 97.855 63.675 ;
         LAYER m3 ;
         RECT  58.9 76.785 59.39 77.275 ;
         LAYER m3 ;
         RECT  100.62 81.12 101.11 81.61 ;
         LAYER m3 ;
         RECT  148.805 79.815 149.295 80.305 ;
         LAYER m3 ;
         RECT  51.29 73.22 51.78 73.71 ;
         LAYER m3 ;
         RECT  26.565 20.965 27.055 21.455 ;
         LAYER m3 ;
         RECT  54.545 84.91 55.035 85.4 ;
         LAYER m3 ;
         RECT  43.475 75.035 43.965 75.525 ;
         LAYER m3 ;
         RECT  77.61 58.355 77.91 58.655 ;
         LAYER m3 ;
         RECT  108.435 67.135 108.925 67.625 ;
         LAYER m3 ;
         RECT  40.22 79.02 40.71 79.51 ;
         LAYER m3 ;
         RECT  54.545 88.86 55.035 89.35 ;
         LAYER m3 ;
         RECT  73.8 98.425 74.29 98.915 ;
         LAYER m3 ;
         RECT  43.475 78.985 43.965 79.475 ;
         LAYER m3 ;
         RECT  24.065 129.525 24.555 130.015 ;
         LAYER m3 ;
         RECT  76.61 107.845 77.1 108.335 ;
         LAYER m3 ;
         RECT  26.565 49.245 27.055 49.735 ;
         LAYER m3 ;
         RECT  54.545 75.035 55.035 75.525 ;
         LAYER m3 ;
         RECT  76.55 112.035 77.04 112.525 ;
         LAYER m3 ;
         RECT  100.62 86.92 101.11 87.41 ;
         LAYER m3 ;
         RECT  151.045 132.765 151.535 133.255 ;
         LAYER m3 ;
         RECT  5.675 107.515 6.165 108.005 ;
         LAYER m3 ;
         RECT  108.435 78.985 108.925 79.475 ;
         LAYER m3 ;
         RECT  51.29 63.22 51.78 63.71 ;
         LAYER m3 ;
         RECT  80.635 58.26 81.125 58.75 ;
         LAYER m3 ;
         RECT  51.29 82.97 51.78 83.46 ;
         LAYER m3 ;
         RECT  100.62 89.02 101.11 89.51 ;
         LAYER m3 ;
         RECT  41.585 6.825 42.075 7.315 ;
         LAYER m3 ;
         RECT  54.545 71.085 55.035 71.575 ;
         LAYER m3 ;
         RECT  125.765 118.625 126.255 119.115 ;
         LAYER m3 ;
         RECT  128.265 38.345 128.755 38.835 ;
         LAYER m3 ;
         RECT  111.69 79.02 112.18 79.51 ;
         LAYER m3 ;
         RECT  100.62 90.87 101.11 91.36 ;
         LAYER m3 ;
         RECT  100.62 79.02 101.11 79.51 ;
         LAYER m3 ;
         RECT  100.62 71.12 101.11 71.61 ;
         LAYER m3 ;
         RECT  26.565 35.105 27.055 35.595 ;
         LAYER m3 ;
         RECT  148.805 68.615 149.295 69.105 ;
         LAYER m3 ;
         RECT  97.365 69.11 97.855 69.6 ;
         LAYER m3 ;
         RECT  145.125 68.615 145.615 69.105 ;
         LAYER m3 ;
         RECT  97.365 82.935 97.855 83.425 ;
         LAYER m3 ;
         RECT  51.29 89.02 51.78 89.51 ;
         LAYER m3 ;
         RECT  125.765 104.485 126.255 104.975 ;
         LAYER m3 ;
         RECT  97.365 90.835 97.855 91.325 ;
         LAYER m3 ;
         RECT  97.365 88.86 97.855 89.35 ;
         LAYER m3 ;
         RECT  51.29 75.07 51.78 75.56 ;
         LAYER m3 ;
         RECT  145.125 57.415 145.615 57.905 ;
         LAYER m3 ;
         RECT  74.49 95.565 74.79 95.865 ;
         LAYER m3 ;
         RECT  51.29 69.27 51.78 69.76 ;
         LAYER m3 ;
         RECT  74.49 58.355 74.79 58.655 ;
         LAYER m3 ;
         RECT  1.995 107.515 2.485 108.005 ;
         LAYER m3 ;
         RECT  97.365 75.035 97.855 75.525 ;
         LAYER m3 ;
         RECT  88.435 76.865 88.925 77.355 ;
         LAYER m3 ;
         RECT  74.68 45.885 75.17 46.375 ;
         LAYER m3 ;
         RECT  51.29 77.17 51.78 77.66 ;
         LAYER m3 ;
         RECT  5.675 85.115 6.165 85.605 ;
         LAYER m3 ;
         RECT  54.545 69.11 55.035 69.6 ;
         LAYER m3 ;
         RECT  26.565 6.825 27.055 7.315 ;
         LAYER m3 ;
         RECT  73.8 55.305 74.29 55.795 ;
         LAYER m3 ;
         RECT  108.435 75.035 108.925 75.525 ;
         LAYER m3 ;
         RECT  77.175 33.935 77.665 34.425 ;
         LAYER m3 ;
         RECT  100.62 69.27 101.11 69.76 ;
         LAYER m3 ;
         RECT  -0.245 6.825 0.245 7.315 ;
         LAYER m3 ;
         RECT  74.74 41.695 75.23 42.185 ;
         LAYER m3 ;
         RECT  97.365 78.985 97.855 79.475 ;
         LAYER m3 ;
         RECT  145.125 91.015 145.615 91.505 ;
         LAYER m3 ;
         RECT  54.545 77.01 55.035 77.5 ;
         LAYER m3 ;
         RECT  54.545 80.96 55.035 81.45 ;
         LAYER m3 ;
         RECT  97.365 73.06 97.855 73.55 ;
         LAYER m3 ;
         RECT  51.29 65.32 51.78 65.81 ;
         LAYER m3 ;
         RECT  97.365 80.96 97.855 81.45 ;
         LAYER m3 ;
         RECT  97.365 65.16 97.855 65.65 ;
         LAYER m3 ;
         RECT  80.04 98.425 80.53 98.915 ;
         LAYER m3 ;
         RECT  128.265 24.205 128.755 24.695 ;
         LAYER m3 ;
         RECT  100.62 63.22 101.11 63.71 ;
         LAYER m3 ;
         RECT  51.29 79.02 51.78 79.51 ;
         LAYER m3 ;
         RECT  74.68 107.845 75.17 108.335 ;
         LAYER m3 ;
         RECT  5.675 73.915 6.165 74.405 ;
         LAYER m3 ;
         RECT  51.29 90.87 51.78 91.36 ;
         LAYER m3 ;
         RECT  108.435 63.185 108.925 63.675 ;
         LAYER m3 ;
         RECT  51.29 86.92 51.78 87.41 ;
         LAYER m3 ;
         RECT  54.545 86.885 55.035 87.375 ;
         LAYER m3 ;
         RECT  51.29 81.12 51.78 81.61 ;
         LAYER m3 ;
         RECT  80.635 95.47 81.125 95.96 ;
         LAYER m3 ;
         RECT  43.475 63.185 43.965 63.675 ;
         LAYER m3 ;
         RECT  54.545 63.185 55.035 63.675 ;
         LAYER m3 ;
         RECT  97.365 77.01 97.855 77.5 ;
         LAYER m3 ;
         RECT  43.475 67.135 43.965 67.625 ;
         LAYER m3 ;
         RECT  40.22 67.17 40.71 67.66 ;
         LAYER m3 ;
         RECT  33.605 63.185 34.095 63.675 ;
         LAYER m3 ;
         RECT  118.305 63.185 118.795 63.675 ;
         LAYER m3 ;
         RECT  51.29 67.17 51.78 67.66 ;
         LAYER m3 ;
         RECT  148.805 57.415 149.295 57.905 ;
         LAYER m3 ;
         RECT  145.125 79.815 145.615 80.305 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER m3 ;
         RECT  102.745 69.26 103.235 69.75 ;
         LAYER m3 ;
         RECT  5.675 79.515 6.165 80.005 ;
         LAYER m3 ;
         RECT  148.805 63.015 149.295 63.505 ;
         LAYER m3 ;
         RECT  49.165 85.06 49.655 85.55 ;
         LAYER m3 ;
         RECT  32.245 75.035 32.735 75.525 ;
         LAYER m3 ;
         RECT  125.765 125.695 126.255 126.185 ;
         LAYER m3 ;
         RECT  77.12 36.12 77.61 36.61 ;
         LAYER m3 ;
         RECT  5.675 68.315 6.165 68.805 ;
         LAYER m3 ;
         RECT  84.21 80.91 84.51 81.21 ;
         LAYER m3 ;
         RECT  113.815 75.07 114.305 75.56 ;
         LAYER m3 ;
         RECT  26.565 56.315 27.055 56.805 ;
         LAYER m3 ;
         RECT  67.89 70.245 68.19 70.545 ;
         LAYER m3 ;
         RECT  53.185 90.835 53.675 91.325 ;
         LAYER m3 ;
         RECT  1.995 68.315 2.485 68.805 ;
         LAYER m3 ;
         RECT  38.095 67.17 38.585 67.66 ;
         LAYER m3 ;
         RECT  84.21 88.81 84.51 89.11 ;
         LAYER m3 ;
         RECT  67.89 78.145 68.19 78.445 ;
         LAYER m3 ;
         RECT  53.185 69.11 53.675 69.6 ;
         LAYER m3 ;
         RECT  74.17 36.12 74.66 36.61 ;
         LAYER m3 ;
         RECT  49.165 71.12 49.655 71.61 ;
         LAYER m3 ;
         RECT  77.145 31.265 77.635 31.755 ;
         LAYER m3 ;
         RECT  98.725 78.985 99.215 79.475 ;
         LAYER m3 ;
         RECT  109.795 75.035 110.285 75.525 ;
         LAYER m3 ;
         RECT  90.925 76.865 91.415 77.355 ;
         LAYER m3 ;
         RECT  102.745 85.06 103.235 85.55 ;
         LAYER m3 ;
         RECT  84.21 74.195 84.51 74.495 ;
         LAYER m3 ;
         RECT  53.185 75.035 53.675 75.525 ;
         LAYER m3 ;
         RECT  67.89 63.925 68.19 64.225 ;
         LAYER m3 ;
         RECT  49.165 63.22 49.655 63.71 ;
         LAYER m3 ;
         RECT  53.185 86.885 53.675 87.375 ;
         LAYER m3 ;
         RECT  74.72 32.275 75.21 32.765 ;
         LAYER m3 ;
         RECT  76.55 113.645 77.04 114.135 ;
         LAYER m3 ;
         RECT  148.805 74.215 149.295 74.705 ;
         LAYER m3 ;
         RECT  67.89 92.76 68.19 93.06 ;
         LAYER m3 ;
         RECT  38.095 63.22 38.585 63.71 ;
         LAYER m3 ;
         RECT  49.165 65.31 49.655 65.8 ;
         LAYER m3 ;
         RECT  49.165 82.97 49.655 83.46 ;
         LAYER m3 ;
         RECT  84.21 79.725 84.51 80.025 ;
         LAYER m3 ;
         RECT  53.185 67.135 53.675 67.625 ;
         LAYER m3 ;
         RECT  24.065 122.455 24.555 122.945 ;
         LAYER m3 ;
         RECT  76.55 40.085 77.04 40.575 ;
         LAYER m3 ;
         RECT  119.665 63.185 120.155 63.675 ;
         LAYER m3 ;
         RECT  84.21 63.925 84.51 64.225 ;
         LAYER m3 ;
         RECT  84.21 91.575 84.51 91.875 ;
         LAYER m3 ;
         RECT  98.725 77.01 99.215 77.5 ;
         LAYER m3 ;
         RECT  56.775 76.79 57.265 77.28 ;
         LAYER m3 ;
         RECT  67.89 82.095 68.19 82.395 ;
         LAYER m3 ;
         RECT  109.795 67.135 110.285 67.625 ;
         LAYER m3 ;
         RECT  84.21 73.01 84.51 73.31 ;
         LAYER m3 ;
         RECT  102.745 75.07 103.235 75.56 ;
         LAYER m3 ;
         RECT  102.745 65.31 103.235 65.8 ;
         LAYER m3 ;
         RECT  102.745 71.12 103.235 71.61 ;
         LAYER m3 ;
         RECT  84.21 59.975 84.51 60.275 ;
         LAYER m3 ;
         RECT  67.89 86.045 68.19 86.345 ;
         LAYER m3 ;
         RECT  67.89 91.575 68.19 91.875 ;
         LAYER m3 ;
         RECT  98.725 88.86 99.215 89.35 ;
         LAYER m3 ;
         RECT  49.165 67.17 49.655 67.66 ;
         LAYER m3 ;
         RECT  125.765 139.835 126.255 140.325 ;
         LAYER m3 ;
         RECT  102.745 81.11 103.235 81.6 ;
         LAYER m3 ;
         RECT  1.995 101.915 2.485 102.405 ;
         LAYER m3 ;
         RECT  119.665 75.035 120.155 75.525 ;
         LAYER m3 ;
         RECT  53.185 84.91 53.675 85.4 ;
         LAYER m3 ;
         RECT  42.115 67.135 42.605 67.625 ;
         LAYER m3 ;
         RECT  53.185 71.085 53.675 71.575 ;
         LAYER m3 ;
         RECT  67.89 71.825 68.19 72.125 ;
         LAYER m3 ;
         RECT  67.89 76.96 68.19 77.26 ;
         LAYER m3 ;
         RECT  102.745 82.97 103.235 83.46 ;
         LAYER m3 ;
         RECT  75.09 103.975 75.58 104.465 ;
         LAYER m3 ;
         RECT  53.185 63.185 53.675 63.675 ;
         LAYER m3 ;
         RECT  98.725 90.835 99.215 91.325 ;
         LAYER m3 ;
         RECT  84.21 76.96 84.51 77.26 ;
         LAYER m3 ;
         RECT  1.995 79.515 2.485 80.005 ;
         LAYER m3 ;
         RECT  95.135 76.79 95.625 77.28 ;
         LAYER m3 ;
         RECT  98.725 67.135 99.215 67.625 ;
         LAYER m3 ;
         RECT  26.565 28.035 27.055 28.525 ;
         LAYER m3 ;
         RECT  35.745 -0.245 36.235 0.245 ;
         LAYER m3 ;
         RECT  84.21 69.06 84.51 69.36 ;
         LAYER m3 ;
         RECT  38.095 75.07 38.585 75.56 ;
         LAYER m3 ;
         RECT  109.795 78.985 110.285 79.475 ;
         LAYER m3 ;
         RECT  98.725 63.185 99.215 63.675 ;
         LAYER m3 ;
         RECT  125.765 97.415 126.255 97.905 ;
         LAYER m3 ;
         RECT  113.815 79.02 114.305 79.51 ;
         LAYER m3 ;
         RECT  102.745 89.01 103.235 89.5 ;
         LAYER m3 ;
         RECT  84.21 61.16 84.51 61.46 ;
         LAYER m3 ;
         RECT  128.265 17.135 128.755 17.625 ;
         LAYER m3 ;
         RECT  84.21 82.095 84.51 82.395 ;
         LAYER m3 ;
         RECT  49.165 77.16 49.655 77.65 ;
         LAYER m3 ;
         RECT  74.145 31.265 74.635 31.755 ;
         LAYER m3 ;
         RECT  98.725 69.11 99.215 69.6 ;
         LAYER m3 ;
         RECT  102.745 73.21 103.235 73.7 ;
         LAYER m3 ;
         RECT  38.095 79.02 38.585 79.51 ;
         LAYER m3 ;
         RECT  67.89 79.725 68.19 80.025 ;
         LAYER m3 ;
         RECT  84.21 75.775 84.51 76.075 ;
         LAYER m3 ;
         RECT  102.745 67.17 103.235 67.66 ;
         LAYER m3 ;
         RECT  67.89 61.16 68.19 61.46 ;
         LAYER m3 ;
         RECT  145.125 74.215 145.615 74.705 ;
         LAYER m3 ;
         RECT  102.745 90.87 103.235 91.36 ;
         LAYER m3 ;
         RECT  74.74 113.645 75.23 114.135 ;
         LAYER m3 ;
         RECT  53.185 82.935 53.675 83.425 ;
         LAYER m3 ;
         RECT  24.065 108.315 24.555 108.805 ;
         LAYER m3 ;
         RECT  84.21 78.145 84.51 78.445 ;
         LAYER m3 ;
         RECT  98.725 80.96 99.215 81.45 ;
         LAYER m3 ;
         RECT  67.89 73.01 68.19 73.31 ;
         LAYER m3 ;
         RECT  84.21 92.76 84.51 93.06 ;
         LAYER m3 ;
         RECT  1.995 90.715 2.485 91.205 ;
         LAYER m3 ;
         RECT  67.89 69.06 68.19 69.36 ;
         LAYER m3 ;
         RECT  84.21 62.345 84.51 62.645 ;
         LAYER m3 ;
         RECT  98.725 82.935 99.215 83.425 ;
         LAYER m3 ;
         RECT  84.21 87.625 84.51 87.925 ;
         LAYER m3 ;
         RECT  67.89 62.345 68.19 62.645 ;
         LAYER m3 ;
         RECT  113.815 67.17 114.305 67.66 ;
         LAYER m3 ;
         RECT  26.565 -0.245 27.055 0.245 ;
         LAYER m3 ;
         RECT  -0.245 13.905 0.245 14.395 ;
         LAYER m3 ;
         RECT  67.89 93.945 68.19 94.245 ;
         LAYER m3 ;
         RECT  84.21 66.295 84.51 66.595 ;
         LAYER m3 ;
         RECT  42.115 63.185 42.605 63.675 ;
         LAYER m3 ;
         RECT  98.725 71.085 99.215 71.575 ;
         LAYER m3 ;
         RECT  53.185 80.96 53.675 81.45 ;
         LAYER m3 ;
         RECT  151.045 139.845 151.535 140.335 ;
         LAYER m3 ;
         RECT  84.21 93.945 84.51 94.245 ;
         LAYER m3 ;
         RECT  49.165 90.87 49.655 91.36 ;
         LAYER m3 ;
         RECT  67.89 80.91 68.19 81.21 ;
         LAYER m3 ;
         RECT  26.565 13.895 27.055 14.385 ;
         LAYER m3 ;
         RECT  84.21 71.825 84.51 72.125 ;
         LAYER m3 ;
         RECT  125.765 111.555 126.255 112.045 ;
         LAYER m3 ;
         RECT  67.89 83.675 68.19 83.975 ;
         LAYER m3 ;
         RECT  67.89 65.11 68.19 65.41 ;
         LAYER m3 ;
         RECT  148.805 85.415 149.295 85.905 ;
         LAYER m3 ;
         RECT  84.21 70.245 84.51 70.545 ;
         LAYER m3 ;
         RECT  67.89 67.875 68.19 68.175 ;
         LAYER m3 ;
         RECT  60.985 76.865 61.475 77.355 ;
         LAYER m3 ;
         RECT  24.065 136.595 24.555 137.085 ;
         LAYER m3 ;
         RECT  84.21 65.11 84.51 65.41 ;
         LAYER m3 ;
         RECT  5.675 90.715 6.165 91.205 ;
         LAYER m3 ;
         RECT  5.675 101.915 6.165 102.405 ;
         LAYER m3 ;
         RECT  148.805 96.615 149.295 97.105 ;
         LAYER m3 ;
         RECT  128.265 31.275 128.755 31.765 ;
         LAYER m3 ;
         RECT  26.565 42.175 27.055 42.665 ;
         LAYER m3 ;
         RECT  49.165 75.07 49.655 75.56 ;
         LAYER m3 ;
         RECT  67.89 89.995 68.19 90.295 ;
         LAYER m3 ;
         RECT  -0.245 -0.255 0.245 0.235 ;
         LAYER m3 ;
         RECT  98.725 84.91 99.215 85.4 ;
         LAYER m3 ;
         RECT  53.185 77.01 53.675 77.5 ;
         LAYER m3 ;
         RECT  53.185 73.06 53.675 73.55 ;
         LAYER m3 ;
         RECT  76.57 32.275 77.06 32.765 ;
         LAYER m3 ;
         RECT  84.21 83.675 84.51 83.975 ;
         LAYER m3 ;
         RECT  42.115 78.985 42.605 79.475 ;
         LAYER m3 ;
         RECT  128.265 45.415 128.755 45.905 ;
         LAYER m3 ;
         RECT  67.89 84.86 68.19 85.16 ;
         LAYER m3 ;
         RECT  67.89 87.625 68.19 87.925 ;
         LAYER m3 ;
         RECT  145.125 85.415 145.615 85.905 ;
         LAYER m3 ;
         RECT  49.165 69.26 49.655 69.75 ;
         LAYER m3 ;
         RECT  98.725 75.035 99.215 75.525 ;
         LAYER m3 ;
         RECT  49.165 81.11 49.655 81.6 ;
         LAYER m3 ;
         RECT  98.725 65.16 99.215 65.65 ;
         LAYER m3 ;
         RECT  53.185 88.86 53.675 89.35 ;
         LAYER m3 ;
         RECT  84.21 84.86 84.51 85.16 ;
         LAYER m3 ;
         RECT  145.125 51.815 145.615 52.305 ;
         LAYER m3 ;
         RECT  1.995 57.115 2.485 57.605 ;
         LAYER m3 ;
         RECT  145.125 63.015 145.615 63.505 ;
         LAYER m3 ;
         RECT  49.165 73.21 49.655 73.7 ;
         LAYER m3 ;
         RECT  148.805 51.815 149.295 52.305 ;
         LAYER m3 ;
         RECT  84.21 67.875 84.51 68.175 ;
         LAYER m3 ;
         RECT  49.165 89.01 49.655 89.5 ;
         LAYER m3 ;
         RECT  84.21 89.995 84.51 90.295 ;
         LAYER m3 ;
         RECT  49.165 79.02 49.655 79.51 ;
         LAYER m3 ;
         RECT  67.89 74.195 68.19 74.495 ;
         LAYER m3 ;
         RECT  74.74 40.085 75.23 40.575 ;
         LAYER m3 ;
         RECT  67.89 75.775 68.19 76.075 ;
         LAYER m3 ;
         RECT  67.89 59.975 68.19 60.275 ;
         LAYER m3 ;
         RECT  53.185 65.16 53.675 65.65 ;
         LAYER m3 ;
         RECT  41.585 -0.245 42.075 0.245 ;
         LAYER m3 ;
         RECT  84.21 86.045 84.51 86.345 ;
         LAYER m3 ;
         RECT  5.675 57.115 6.165 57.605 ;
         LAYER m3 ;
         RECT  102.745 79.02 103.235 79.51 ;
         LAYER m3 ;
         RECT  109.795 63.185 110.285 63.675 ;
         LAYER m3 ;
         RECT  102.745 63.22 103.235 63.71 ;
         LAYER m3 ;
         RECT  98.725 73.06 99.215 73.55 ;
         LAYER m3 ;
         RECT  67.89 88.81 68.19 89.11 ;
         LAYER m3 ;
         RECT  49.165 86.92 49.655 87.41 ;
         LAYER m3 ;
         RECT  98.725 86.885 99.215 87.375 ;
         LAYER m3 ;
         RECT  67.89 66.295 68.19 66.595 ;
         LAYER m3 ;
         RECT  76.2 49.755 76.69 50.245 ;
         LAYER m3 ;
         RECT  145.125 96.615 145.615 97.105 ;
         LAYER m3 ;
         RECT  53.185 78.985 53.675 79.475 ;
         LAYER m3 ;
         RECT  102.745 77.16 103.235 77.65 ;
         LAYER m3 ;
         RECT  102.745 86.92 103.235 87.41 ;
         LAYER m3 ;
         RECT  32.245 63.185 32.735 63.675 ;
         LAYER m3 ;
         RECT  113.815 63.22 114.305 63.71 ;
         LAYER m3 ;
         RECT  76.2 103.975 76.69 104.465 ;
         LAYER m3 ;
         RECT  75.09 49.755 75.58 50.245 ;
         LAYER m3 ;
         RECT  42.115 75.035 42.605 75.525 ;
      END
   END gnd
   OBS
   LAYER  m1 ;
      RECT  75.915 61.705 75.99 63.41 ;
      RECT  75.99 61.12 76.2 61.5 ;
      RECT  73.83 60.79 74.01 61.705 ;
      POLYGON  75.48 61.795 75.48 62.205 75.655 62.205 75.735 62.125 75.735 61.795 75.48 61.795 ;
      RECT  73.47 61.705 73.65 63.41 ;
      RECT  73.83 61.705 74.01 63.41 ;
      RECT  73.08 61.705 73.29 63.41 ;
      RECT  72.87 61.5 73.08 61.705 ;
      RECT  72.87 61.705 73.08 63.41 ;
      RECT  75.99 61.705 76.2 63.41 ;
      POLYGON  75.48 62.785 75.48 63.195 75.735 63.195 75.735 62.865 75.655 62.785 75.48 62.785 ;
      RECT  73.08 61.12 73.29 61.5 ;
      RECT  75.99 60.79 76.2 61.12 ;
      RECT  74.19 60.79 74.37 61.705 ;
      RECT  75.83 62.29 75.915 62.7 ;
      RECT  74.91 61.705 75.09 63.41 ;
      RECT  75.27 62.785 75.48 63.195 ;
      RECT  73.08 60.79 73.29 61.12 ;
      RECT  75.27 61.795 75.48 62.205 ;
      RECT  75.27 61.12 75.48 61.5 ;
      RECT  72.87 61.12 73.08 61.5 ;
      RECT  74.55 60.79 74.73 61.705 ;
      RECT  74.55 61.705 74.73 63.41 ;
      RECT  75.99 61.5 76.2 61.705 ;
      RECT  73.08 61.5 73.29 61.705 ;
      RECT  72.87 60.79 73.08 61.12 ;
      RECT  74.91 60.79 75.09 61.705 ;
      RECT  73.47 60.79 73.65 61.705 ;
      POLYGON  75.915 60.79 75.915 61.12 75.48 61.12 75.48 61.5 75.915 61.5 75.915 61.705 75.99 61.705 75.99 60.79 75.915 60.79 ;
      RECT  74.19 61.705 74.37 63.41 ;
      RECT  75.915 64.865 75.99 63.16 ;
      RECT  75.99 65.45 76.2 65.07 ;
      RECT  73.83 65.78 74.01 64.865 ;
      POLYGON  75.48 64.775 75.48 64.365 75.655 64.365 75.735 64.445 75.735 64.775 75.48 64.775 ;
      RECT  73.47 64.865 73.65 63.16 ;
      RECT  73.83 64.865 74.01 63.16 ;
      RECT  73.08 64.865 73.29 63.16 ;
      RECT  72.87 65.07 73.08 64.865 ;
      RECT  72.87 64.865 73.08 63.16 ;
      RECT  75.99 64.865 76.2 63.16 ;
      POLYGON  75.48 63.785 75.48 63.375 75.735 63.375 75.735 63.705 75.655 63.785 75.48 63.785 ;
      RECT  73.08 65.45 73.29 65.07 ;
      RECT  75.99 65.78 76.2 65.45 ;
      RECT  74.19 65.78 74.37 64.865 ;
      RECT  75.83 64.28 75.915 63.87 ;
      RECT  74.91 64.865 75.09 63.16 ;
      RECT  75.27 63.785 75.48 63.375 ;
      RECT  73.08 65.78 73.29 65.45 ;
      RECT  75.27 64.775 75.48 64.365 ;
      RECT  75.27 65.45 75.48 65.07 ;
      RECT  72.87 65.45 73.08 65.07 ;
      RECT  74.55 65.78 74.73 64.865 ;
      RECT  74.55 64.865 74.73 63.16 ;
      RECT  75.99 65.07 76.2 64.865 ;
      RECT  73.08 65.07 73.29 64.865 ;
      RECT  72.87 65.78 73.08 65.45 ;
      RECT  74.91 65.78 75.09 64.865 ;
      RECT  73.47 65.78 73.65 64.865 ;
      POLYGON  75.915 65.78 75.915 65.45 75.48 65.45 75.48 65.07 75.915 65.07 75.915 64.865 75.99 64.865 75.99 65.78 75.915 65.78 ;
      RECT  74.19 64.865 74.37 63.16 ;
      RECT  75.915 65.655 75.99 67.36 ;
      RECT  75.99 65.07 76.2 65.45 ;
      RECT  73.83 64.74 74.01 65.655 ;
      POLYGON  75.48 65.745 75.48 66.155 75.655 66.155 75.735 66.075 75.735 65.745 75.48 65.745 ;
      RECT  73.47 65.655 73.65 67.36 ;
      RECT  73.83 65.655 74.01 67.36 ;
      RECT  73.08 65.655 73.29 67.36 ;
      RECT  72.87 65.45 73.08 65.655 ;
      RECT  72.87 65.655 73.08 67.36 ;
      RECT  75.99 65.655 76.2 67.36 ;
      POLYGON  75.48 66.735 75.48 67.145 75.735 67.145 75.735 66.815 75.655 66.735 75.48 66.735 ;
      RECT  73.08 65.07 73.29 65.45 ;
      RECT  75.99 64.74 76.2 65.07 ;
      RECT  74.19 64.74 74.37 65.655 ;
      RECT  75.83 66.24 75.915 66.65 ;
      RECT  74.91 65.655 75.09 67.36 ;
      RECT  75.27 66.735 75.48 67.145 ;
      RECT  73.08 64.74 73.29 65.07 ;
      RECT  75.27 65.745 75.48 66.155 ;
      RECT  75.27 65.07 75.48 65.45 ;
      RECT  72.87 65.07 73.08 65.45 ;
      RECT  74.55 64.74 74.73 65.655 ;
      RECT  74.55 65.655 74.73 67.36 ;
      RECT  75.99 65.45 76.2 65.655 ;
      RECT  73.08 65.45 73.29 65.655 ;
      RECT  72.87 64.74 73.08 65.07 ;
      RECT  74.91 64.74 75.09 65.655 ;
      RECT  73.47 64.74 73.65 65.655 ;
      POLYGON  75.915 64.74 75.915 65.07 75.48 65.07 75.48 65.45 75.915 65.45 75.915 65.655 75.99 65.655 75.99 64.74 75.915 64.74 ;
      RECT  74.19 65.655 74.37 67.36 ;
      RECT  75.915 68.815 75.99 67.11 ;
      RECT  75.99 69.4 76.2 69.02 ;
      RECT  73.83 69.73 74.01 68.815 ;
      POLYGON  75.48 68.725 75.48 68.315 75.655 68.315 75.735 68.395 75.735 68.725 75.48 68.725 ;
      RECT  73.47 68.815 73.65 67.11 ;
      RECT  73.83 68.815 74.01 67.11 ;
      RECT  73.08 68.815 73.29 67.11 ;
      RECT  72.87 69.02 73.08 68.815 ;
      RECT  72.87 68.815 73.08 67.11 ;
      RECT  75.99 68.815 76.2 67.11 ;
      POLYGON  75.48 67.735 75.48 67.325 75.735 67.325 75.735 67.655 75.655 67.735 75.48 67.735 ;
      RECT  73.08 69.4 73.29 69.02 ;
      RECT  75.99 69.73 76.2 69.4 ;
      RECT  74.19 69.73 74.37 68.815 ;
      RECT  75.83 68.23 75.915 67.82 ;
      RECT  74.91 68.815 75.09 67.11 ;
      RECT  75.27 67.735 75.48 67.325 ;
      RECT  73.08 69.73 73.29 69.4 ;
      RECT  75.27 68.725 75.48 68.315 ;
      RECT  75.27 69.4 75.48 69.02 ;
      RECT  72.87 69.4 73.08 69.02 ;
      RECT  74.55 69.73 74.73 68.815 ;
      RECT  74.55 68.815 74.73 67.11 ;
      RECT  75.99 69.02 76.2 68.815 ;
      RECT  73.08 69.02 73.29 68.815 ;
      RECT  72.87 69.73 73.08 69.4 ;
      RECT  74.91 69.73 75.09 68.815 ;
      RECT  73.47 69.73 73.65 68.815 ;
      POLYGON  75.915 69.73 75.915 69.4 75.48 69.4 75.48 69.02 75.915 69.02 75.915 68.815 75.99 68.815 75.99 69.73 75.915 69.73 ;
      RECT  74.19 68.815 74.37 67.11 ;
      RECT  75.915 69.605 75.99 71.31 ;
      RECT  75.99 69.02 76.2 69.4 ;
      RECT  73.83 68.69 74.01 69.605 ;
      POLYGON  75.48 69.695 75.48 70.105 75.655 70.105 75.735 70.025 75.735 69.695 75.48 69.695 ;
      RECT  73.47 69.605 73.65 71.31 ;
      RECT  73.83 69.605 74.01 71.31 ;
      RECT  73.08 69.605 73.29 71.31 ;
      RECT  72.87 69.4 73.08 69.605 ;
      RECT  72.87 69.605 73.08 71.31 ;
      RECT  75.99 69.605 76.2 71.31 ;
      POLYGON  75.48 70.685 75.48 71.095 75.735 71.095 75.735 70.765 75.655 70.685 75.48 70.685 ;
      RECT  73.08 69.02 73.29 69.4 ;
      RECT  75.99 68.69 76.2 69.02 ;
      RECT  74.19 68.69 74.37 69.605 ;
      RECT  75.83 70.19 75.915 70.6 ;
      RECT  74.91 69.605 75.09 71.31 ;
      RECT  75.27 70.685 75.48 71.095 ;
      RECT  73.08 68.69 73.29 69.02 ;
      RECT  75.27 69.695 75.48 70.105 ;
      RECT  75.27 69.02 75.48 69.4 ;
      RECT  72.87 69.02 73.08 69.4 ;
      RECT  74.55 68.69 74.73 69.605 ;
      RECT  74.55 69.605 74.73 71.31 ;
      RECT  75.99 69.4 76.2 69.605 ;
      RECT  73.08 69.4 73.29 69.605 ;
      RECT  72.87 68.69 73.08 69.02 ;
      RECT  74.91 68.69 75.09 69.605 ;
      RECT  73.47 68.69 73.65 69.605 ;
      POLYGON  75.915 68.69 75.915 69.02 75.48 69.02 75.48 69.4 75.915 69.4 75.915 69.605 75.99 69.605 75.99 68.69 75.915 68.69 ;
      RECT  74.19 69.605 74.37 71.31 ;
      RECT  75.915 72.765 75.99 71.06 ;
      RECT  75.99 73.35 76.2 72.97 ;
      RECT  73.83 73.68 74.01 72.765 ;
      POLYGON  75.48 72.675 75.48 72.265 75.655 72.265 75.735 72.345 75.735 72.675 75.48 72.675 ;
      RECT  73.47 72.765 73.65 71.06 ;
      RECT  73.83 72.765 74.01 71.06 ;
      RECT  73.08 72.765 73.29 71.06 ;
      RECT  72.87 72.97 73.08 72.765 ;
      RECT  72.87 72.765 73.08 71.06 ;
      RECT  75.99 72.765 76.2 71.06 ;
      POLYGON  75.48 71.685 75.48 71.275 75.735 71.275 75.735 71.605 75.655 71.685 75.48 71.685 ;
      RECT  73.08 73.35 73.29 72.97 ;
      RECT  75.99 73.68 76.2 73.35 ;
      RECT  74.19 73.68 74.37 72.765 ;
      RECT  75.83 72.18 75.915 71.77 ;
      RECT  74.91 72.765 75.09 71.06 ;
      RECT  75.27 71.685 75.48 71.275 ;
      RECT  73.08 73.68 73.29 73.35 ;
      RECT  75.27 72.675 75.48 72.265 ;
      RECT  75.27 73.35 75.48 72.97 ;
      RECT  72.87 73.35 73.08 72.97 ;
      RECT  74.55 73.68 74.73 72.765 ;
      RECT  74.55 72.765 74.73 71.06 ;
      RECT  75.99 72.97 76.2 72.765 ;
      RECT  73.08 72.97 73.29 72.765 ;
      RECT  72.87 73.68 73.08 73.35 ;
      RECT  74.91 73.68 75.09 72.765 ;
      RECT  73.47 73.68 73.65 72.765 ;
      POLYGON  75.915 73.68 75.915 73.35 75.48 73.35 75.48 72.97 75.915 72.97 75.915 72.765 75.99 72.765 75.99 73.68 75.915 73.68 ;
      RECT  74.19 72.765 74.37 71.06 ;
      RECT  75.915 73.555 75.99 75.26 ;
      RECT  75.99 72.97 76.2 73.35 ;
      RECT  73.83 72.64 74.01 73.555 ;
      POLYGON  75.48 73.645 75.48 74.055 75.655 74.055 75.735 73.975 75.735 73.645 75.48 73.645 ;
      RECT  73.47 73.555 73.65 75.26 ;
      RECT  73.83 73.555 74.01 75.26 ;
      RECT  73.08 73.555 73.29 75.26 ;
      RECT  72.87 73.35 73.08 73.555 ;
      RECT  72.87 73.555 73.08 75.26 ;
      RECT  75.99 73.555 76.2 75.26 ;
      POLYGON  75.48 74.635 75.48 75.045 75.735 75.045 75.735 74.715 75.655 74.635 75.48 74.635 ;
      RECT  73.08 72.97 73.29 73.35 ;
      RECT  75.99 72.64 76.2 72.97 ;
      RECT  74.19 72.64 74.37 73.555 ;
      RECT  75.83 74.14 75.915 74.55 ;
      RECT  74.91 73.555 75.09 75.26 ;
      RECT  75.27 74.635 75.48 75.045 ;
      RECT  73.08 72.64 73.29 72.97 ;
      RECT  75.27 73.645 75.48 74.055 ;
      RECT  75.27 72.97 75.48 73.35 ;
      RECT  72.87 72.97 73.08 73.35 ;
      RECT  74.55 72.64 74.73 73.555 ;
      RECT  74.55 73.555 74.73 75.26 ;
      RECT  75.99 73.35 76.2 73.555 ;
      RECT  73.08 73.35 73.29 73.555 ;
      RECT  72.87 72.64 73.08 72.97 ;
      RECT  74.91 72.64 75.09 73.555 ;
      RECT  73.47 72.64 73.65 73.555 ;
      POLYGON  75.915 72.64 75.915 72.97 75.48 72.97 75.48 73.35 75.915 73.35 75.915 73.555 75.99 73.555 75.99 72.64 75.915 72.64 ;
      RECT  74.19 73.555 74.37 75.26 ;
      RECT  75.915 76.715 75.99 75.01 ;
      RECT  75.99 77.3 76.2 76.92 ;
      RECT  73.83 77.63 74.01 76.715 ;
      POLYGON  75.48 76.625 75.48 76.215 75.655 76.215 75.735 76.295 75.735 76.625 75.48 76.625 ;
      RECT  73.47 76.715 73.65 75.01 ;
      RECT  73.83 76.715 74.01 75.01 ;
      RECT  73.08 76.715 73.29 75.01 ;
      RECT  72.87 76.92 73.08 76.715 ;
      RECT  72.87 76.715 73.08 75.01 ;
      RECT  75.99 76.715 76.2 75.01 ;
      POLYGON  75.48 75.635 75.48 75.225 75.735 75.225 75.735 75.555 75.655 75.635 75.48 75.635 ;
      RECT  73.08 77.3 73.29 76.92 ;
      RECT  75.99 77.63 76.2 77.3 ;
      RECT  74.19 77.63 74.37 76.715 ;
      RECT  75.83 76.13 75.915 75.72 ;
      RECT  74.91 76.715 75.09 75.01 ;
      RECT  75.27 75.635 75.48 75.225 ;
      RECT  73.08 77.63 73.29 77.3 ;
      RECT  75.27 76.625 75.48 76.215 ;
      RECT  75.27 77.3 75.48 76.92 ;
      RECT  72.87 77.3 73.08 76.92 ;
      RECT  74.55 77.63 74.73 76.715 ;
      RECT  74.55 76.715 74.73 75.01 ;
      RECT  75.99 76.92 76.2 76.715 ;
      RECT  73.08 76.92 73.29 76.715 ;
      RECT  72.87 77.63 73.08 77.3 ;
      RECT  74.91 77.63 75.09 76.715 ;
      RECT  73.47 77.63 73.65 76.715 ;
      POLYGON  75.915 77.63 75.915 77.3 75.48 77.3 75.48 76.92 75.915 76.92 75.915 76.715 75.99 76.715 75.99 77.63 75.915 77.63 ;
      RECT  74.19 76.715 74.37 75.01 ;
      RECT  75.915 77.505 75.99 79.21 ;
      RECT  75.99 76.92 76.2 77.3 ;
      RECT  73.83 76.59 74.01 77.505 ;
      POLYGON  75.48 77.595 75.48 78.005 75.655 78.005 75.735 77.925 75.735 77.595 75.48 77.595 ;
      RECT  73.47 77.505 73.65 79.21 ;
      RECT  73.83 77.505 74.01 79.21 ;
      RECT  73.08 77.505 73.29 79.21 ;
      RECT  72.87 77.3 73.08 77.505 ;
      RECT  72.87 77.505 73.08 79.21 ;
      RECT  75.99 77.505 76.2 79.21 ;
      POLYGON  75.48 78.585 75.48 78.995 75.735 78.995 75.735 78.665 75.655 78.585 75.48 78.585 ;
      RECT  73.08 76.92 73.29 77.3 ;
      RECT  75.99 76.59 76.2 76.92 ;
      RECT  74.19 76.59 74.37 77.505 ;
      RECT  75.83 78.09 75.915 78.5 ;
      RECT  74.91 77.505 75.09 79.21 ;
      RECT  75.27 78.585 75.48 78.995 ;
      RECT  73.08 76.59 73.29 76.92 ;
      RECT  75.27 77.595 75.48 78.005 ;
      RECT  75.27 76.92 75.48 77.3 ;
      RECT  72.87 76.92 73.08 77.3 ;
      RECT  74.55 76.59 74.73 77.505 ;
      RECT  74.55 77.505 74.73 79.21 ;
      RECT  75.99 77.3 76.2 77.505 ;
      RECT  73.08 77.3 73.29 77.505 ;
      RECT  72.87 76.59 73.08 76.92 ;
      RECT  74.91 76.59 75.09 77.505 ;
      RECT  73.47 76.59 73.65 77.505 ;
      POLYGON  75.915 76.59 75.915 76.92 75.48 76.92 75.48 77.3 75.915 77.3 75.915 77.505 75.99 77.505 75.99 76.59 75.915 76.59 ;
      RECT  74.19 77.505 74.37 79.21 ;
      RECT  75.915 80.665 75.99 78.96 ;
      RECT  75.99 81.25 76.2 80.87 ;
      RECT  73.83 81.58 74.01 80.665 ;
      POLYGON  75.48 80.575 75.48 80.165 75.655 80.165 75.735 80.245 75.735 80.575 75.48 80.575 ;
      RECT  73.47 80.665 73.65 78.96 ;
      RECT  73.83 80.665 74.01 78.96 ;
      RECT  73.08 80.665 73.29 78.96 ;
      RECT  72.87 80.87 73.08 80.665 ;
      RECT  72.87 80.665 73.08 78.96 ;
      RECT  75.99 80.665 76.2 78.96 ;
      POLYGON  75.48 79.585 75.48 79.175 75.735 79.175 75.735 79.505 75.655 79.585 75.48 79.585 ;
      RECT  73.08 81.25 73.29 80.87 ;
      RECT  75.99 81.58 76.2 81.25 ;
      RECT  74.19 81.58 74.37 80.665 ;
      RECT  75.83 80.08 75.915 79.67 ;
      RECT  74.91 80.665 75.09 78.96 ;
      RECT  75.27 79.585 75.48 79.175 ;
      RECT  73.08 81.58 73.29 81.25 ;
      RECT  75.27 80.575 75.48 80.165 ;
      RECT  75.27 81.25 75.48 80.87 ;
      RECT  72.87 81.25 73.08 80.87 ;
      RECT  74.55 81.58 74.73 80.665 ;
      RECT  74.55 80.665 74.73 78.96 ;
      RECT  75.99 80.87 76.2 80.665 ;
      RECT  73.08 80.87 73.29 80.665 ;
      RECT  72.87 81.58 73.08 81.25 ;
      RECT  74.91 81.58 75.09 80.665 ;
      RECT  73.47 81.58 73.65 80.665 ;
      POLYGON  75.915 81.58 75.915 81.25 75.48 81.25 75.48 80.87 75.915 80.87 75.915 80.665 75.99 80.665 75.99 81.58 75.915 81.58 ;
      RECT  74.19 80.665 74.37 78.96 ;
      RECT  75.915 81.455 75.99 83.16 ;
      RECT  75.99 80.87 76.2 81.25 ;
      RECT  73.83 80.54 74.01 81.455 ;
      POLYGON  75.48 81.545 75.48 81.955 75.655 81.955 75.735 81.875 75.735 81.545 75.48 81.545 ;
      RECT  73.47 81.455 73.65 83.16 ;
      RECT  73.83 81.455 74.01 83.16 ;
      RECT  73.08 81.455 73.29 83.16 ;
      RECT  72.87 81.25 73.08 81.455 ;
      RECT  72.87 81.455 73.08 83.16 ;
      RECT  75.99 81.455 76.2 83.16 ;
      POLYGON  75.48 82.535 75.48 82.945 75.735 82.945 75.735 82.615 75.655 82.535 75.48 82.535 ;
      RECT  73.08 80.87 73.29 81.25 ;
      RECT  75.99 80.54 76.2 80.87 ;
      RECT  74.19 80.54 74.37 81.455 ;
      RECT  75.83 82.04 75.915 82.45 ;
      RECT  74.91 81.455 75.09 83.16 ;
      RECT  75.27 82.535 75.48 82.945 ;
      RECT  73.08 80.54 73.29 80.87 ;
      RECT  75.27 81.545 75.48 81.955 ;
      RECT  75.27 80.87 75.48 81.25 ;
      RECT  72.87 80.87 73.08 81.25 ;
      RECT  74.55 80.54 74.73 81.455 ;
      RECT  74.55 81.455 74.73 83.16 ;
      RECT  75.99 81.25 76.2 81.455 ;
      RECT  73.08 81.25 73.29 81.455 ;
      RECT  72.87 80.54 73.08 80.87 ;
      RECT  74.91 80.54 75.09 81.455 ;
      RECT  73.47 80.54 73.65 81.455 ;
      POLYGON  75.915 80.54 75.915 80.87 75.48 80.87 75.48 81.25 75.915 81.25 75.915 81.455 75.99 81.455 75.99 80.54 75.915 80.54 ;
      RECT  74.19 81.455 74.37 83.16 ;
      RECT  75.915 84.615 75.99 82.91 ;
      RECT  75.99 85.2 76.2 84.82 ;
      RECT  73.83 85.53 74.01 84.615 ;
      POLYGON  75.48 84.525 75.48 84.115 75.655 84.115 75.735 84.195 75.735 84.525 75.48 84.525 ;
      RECT  73.47 84.615 73.65 82.91 ;
      RECT  73.83 84.615 74.01 82.91 ;
      RECT  73.08 84.615 73.29 82.91 ;
      RECT  72.87 84.82 73.08 84.615 ;
      RECT  72.87 84.615 73.08 82.91 ;
      RECT  75.99 84.615 76.2 82.91 ;
      POLYGON  75.48 83.535 75.48 83.125 75.735 83.125 75.735 83.455 75.655 83.535 75.48 83.535 ;
      RECT  73.08 85.2 73.29 84.82 ;
      RECT  75.99 85.53 76.2 85.2 ;
      RECT  74.19 85.53 74.37 84.615 ;
      RECT  75.83 84.03 75.915 83.62 ;
      RECT  74.91 84.615 75.09 82.91 ;
      RECT  75.27 83.535 75.48 83.125 ;
      RECT  73.08 85.53 73.29 85.2 ;
      RECT  75.27 84.525 75.48 84.115 ;
      RECT  75.27 85.2 75.48 84.82 ;
      RECT  72.87 85.2 73.08 84.82 ;
      RECT  74.55 85.53 74.73 84.615 ;
      RECT  74.55 84.615 74.73 82.91 ;
      RECT  75.99 84.82 76.2 84.615 ;
      RECT  73.08 84.82 73.29 84.615 ;
      RECT  72.87 85.53 73.08 85.2 ;
      RECT  74.91 85.53 75.09 84.615 ;
      RECT  73.47 85.53 73.65 84.615 ;
      POLYGON  75.915 85.53 75.915 85.2 75.48 85.2 75.48 84.82 75.915 84.82 75.915 84.615 75.99 84.615 75.99 85.53 75.915 85.53 ;
      RECT  74.19 84.615 74.37 82.91 ;
      RECT  75.915 85.405 75.99 87.11 ;
      RECT  75.99 84.82 76.2 85.2 ;
      RECT  73.83 84.49 74.01 85.405 ;
      POLYGON  75.48 85.495 75.48 85.905 75.655 85.905 75.735 85.825 75.735 85.495 75.48 85.495 ;
      RECT  73.47 85.405 73.65 87.11 ;
      RECT  73.83 85.405 74.01 87.11 ;
      RECT  73.08 85.405 73.29 87.11 ;
      RECT  72.87 85.2 73.08 85.405 ;
      RECT  72.87 85.405 73.08 87.11 ;
      RECT  75.99 85.405 76.2 87.11 ;
      POLYGON  75.48 86.485 75.48 86.895 75.735 86.895 75.735 86.565 75.655 86.485 75.48 86.485 ;
      RECT  73.08 84.82 73.29 85.2 ;
      RECT  75.99 84.49 76.2 84.82 ;
      RECT  74.19 84.49 74.37 85.405 ;
      RECT  75.83 85.99 75.915 86.4 ;
      RECT  74.91 85.405 75.09 87.11 ;
      RECT  75.27 86.485 75.48 86.895 ;
      RECT  73.08 84.49 73.29 84.82 ;
      RECT  75.27 85.495 75.48 85.905 ;
      RECT  75.27 84.82 75.48 85.2 ;
      RECT  72.87 84.82 73.08 85.2 ;
      RECT  74.55 84.49 74.73 85.405 ;
      RECT  74.55 85.405 74.73 87.11 ;
      RECT  75.99 85.2 76.2 85.405 ;
      RECT  73.08 85.2 73.29 85.405 ;
      RECT  72.87 84.49 73.08 84.82 ;
      RECT  74.91 84.49 75.09 85.405 ;
      RECT  73.47 84.49 73.65 85.405 ;
      POLYGON  75.915 84.49 75.915 84.82 75.48 84.82 75.48 85.2 75.915 85.2 75.915 85.405 75.99 85.405 75.99 84.49 75.915 84.49 ;
      RECT  74.19 85.405 74.37 87.11 ;
      RECT  75.915 88.565 75.99 86.86 ;
      RECT  75.99 89.15 76.2 88.77 ;
      RECT  73.83 89.48 74.01 88.565 ;
      POLYGON  75.48 88.475 75.48 88.065 75.655 88.065 75.735 88.145 75.735 88.475 75.48 88.475 ;
      RECT  73.47 88.565 73.65 86.86 ;
      RECT  73.83 88.565 74.01 86.86 ;
      RECT  73.08 88.565 73.29 86.86 ;
      RECT  72.87 88.77 73.08 88.565 ;
      RECT  72.87 88.565 73.08 86.86 ;
      RECT  75.99 88.565 76.2 86.86 ;
      POLYGON  75.48 87.485 75.48 87.075 75.735 87.075 75.735 87.405 75.655 87.485 75.48 87.485 ;
      RECT  73.08 89.15 73.29 88.77 ;
      RECT  75.99 89.48 76.2 89.15 ;
      RECT  74.19 89.48 74.37 88.565 ;
      RECT  75.83 87.98 75.915 87.57 ;
      RECT  74.91 88.565 75.09 86.86 ;
      RECT  75.27 87.485 75.48 87.075 ;
      RECT  73.08 89.48 73.29 89.15 ;
      RECT  75.27 88.475 75.48 88.065 ;
      RECT  75.27 89.15 75.48 88.77 ;
      RECT  72.87 89.15 73.08 88.77 ;
      RECT  74.55 89.48 74.73 88.565 ;
      RECT  74.55 88.565 74.73 86.86 ;
      RECT  75.99 88.77 76.2 88.565 ;
      RECT  73.08 88.77 73.29 88.565 ;
      RECT  72.87 89.48 73.08 89.15 ;
      RECT  74.91 89.48 75.09 88.565 ;
      RECT  73.47 89.48 73.65 88.565 ;
      POLYGON  75.915 89.48 75.915 89.15 75.48 89.15 75.48 88.77 75.915 88.77 75.915 88.565 75.99 88.565 75.99 89.48 75.915 89.48 ;
      RECT  74.19 88.565 74.37 86.86 ;
      RECT  75.915 89.355 75.99 91.06 ;
      RECT  75.99 88.77 76.2 89.15 ;
      RECT  73.83 88.44 74.01 89.355 ;
      POLYGON  75.48 89.445 75.48 89.855 75.655 89.855 75.735 89.775 75.735 89.445 75.48 89.445 ;
      RECT  73.47 89.355 73.65 91.06 ;
      RECT  73.83 89.355 74.01 91.06 ;
      RECT  73.08 89.355 73.29 91.06 ;
      RECT  72.87 89.15 73.08 89.355 ;
      RECT  72.87 89.355 73.08 91.06 ;
      RECT  75.99 89.355 76.2 91.06 ;
      POLYGON  75.48 90.435 75.48 90.845 75.735 90.845 75.735 90.515 75.655 90.435 75.48 90.435 ;
      RECT  73.08 88.77 73.29 89.15 ;
      RECT  75.99 88.44 76.2 88.77 ;
      RECT  74.19 88.44 74.37 89.355 ;
      RECT  75.83 89.94 75.915 90.35 ;
      RECT  74.91 89.355 75.09 91.06 ;
      RECT  75.27 90.435 75.48 90.845 ;
      RECT  73.08 88.44 73.29 88.77 ;
      RECT  75.27 89.445 75.48 89.855 ;
      RECT  75.27 88.77 75.48 89.15 ;
      RECT  72.87 88.77 73.08 89.15 ;
      RECT  74.55 88.44 74.73 89.355 ;
      RECT  74.55 89.355 74.73 91.06 ;
      RECT  75.99 89.15 76.2 89.355 ;
      RECT  73.08 89.15 73.29 89.355 ;
      RECT  72.87 88.44 73.08 88.77 ;
      RECT  74.91 88.44 75.09 89.355 ;
      RECT  73.47 88.44 73.65 89.355 ;
      POLYGON  75.915 88.44 75.915 88.77 75.48 88.77 75.48 89.15 75.915 89.15 75.915 89.355 75.99 89.355 75.99 88.44 75.915 88.44 ;
      RECT  74.19 89.355 74.37 91.06 ;
      RECT  75.915 92.515 75.99 90.81 ;
      RECT  75.99 93.1 76.2 92.72 ;
      RECT  73.83 93.43 74.01 92.515 ;
      POLYGON  75.48 92.425 75.48 92.015 75.655 92.015 75.735 92.095 75.735 92.425 75.48 92.425 ;
      RECT  73.47 92.515 73.65 90.81 ;
      RECT  73.83 92.515 74.01 90.81 ;
      RECT  73.08 92.515 73.29 90.81 ;
      RECT  72.87 92.72 73.08 92.515 ;
      RECT  72.87 92.515 73.08 90.81 ;
      RECT  75.99 92.515 76.2 90.81 ;
      POLYGON  75.48 91.435 75.48 91.025 75.735 91.025 75.735 91.355 75.655 91.435 75.48 91.435 ;
      RECT  73.08 93.1 73.29 92.72 ;
      RECT  75.99 93.43 76.2 93.1 ;
      RECT  74.19 93.43 74.37 92.515 ;
      RECT  75.83 91.93 75.915 91.52 ;
      RECT  74.91 92.515 75.09 90.81 ;
      RECT  75.27 91.435 75.48 91.025 ;
      RECT  73.08 93.43 73.29 93.1 ;
      RECT  75.27 92.425 75.48 92.015 ;
      RECT  75.27 93.1 75.48 92.72 ;
      RECT  72.87 93.1 73.08 92.72 ;
      RECT  74.55 93.43 74.73 92.515 ;
      RECT  74.55 92.515 74.73 90.81 ;
      RECT  75.99 92.72 76.2 92.515 ;
      RECT  73.08 92.72 73.29 92.515 ;
      RECT  72.87 93.43 73.08 93.1 ;
      RECT  74.91 93.43 75.09 92.515 ;
      RECT  73.47 93.43 73.65 92.515 ;
      POLYGON  75.915 93.43 75.915 93.1 75.48 93.1 75.48 92.72 75.915 92.72 75.915 92.515 75.99 92.515 75.99 93.43 75.915 93.43 ;
      RECT  74.19 92.515 74.37 90.81 ;
      RECT  76.485 61.705 76.41 63.41 ;
      RECT  76.41 61.12 76.2 61.5 ;
      RECT  78.57 60.79 78.39 61.705 ;
      POLYGON  76.92 61.795 76.92 62.205 76.745 62.205 76.665 62.125 76.665 61.795 76.92 61.795 ;
      RECT  78.93 61.705 78.75 63.41 ;
      RECT  78.57 61.705 78.39 63.41 ;
      RECT  79.32 61.705 79.11 63.41 ;
      RECT  79.53 61.5 79.32 61.705 ;
      RECT  79.53 61.705 79.32 63.41 ;
      RECT  76.41 61.705 76.2 63.41 ;
      POLYGON  76.92 62.785 76.92 63.195 76.665 63.195 76.665 62.865 76.745 62.785 76.92 62.785 ;
      RECT  79.32 61.12 79.11 61.5 ;
      RECT  76.41 60.79 76.2 61.12 ;
      RECT  78.21 60.79 78.03 61.705 ;
      RECT  76.57 62.29 76.485 62.7 ;
      RECT  77.49 61.705 77.31 63.41 ;
      RECT  77.13 62.785 76.92 63.195 ;
      RECT  79.32 60.79 79.11 61.12 ;
      RECT  77.13 61.795 76.92 62.205 ;
      RECT  77.13 61.12 76.92 61.5 ;
      RECT  79.53 61.12 79.32 61.5 ;
      RECT  77.85 60.79 77.67 61.705 ;
      RECT  77.85 61.705 77.67 63.41 ;
      RECT  76.41 61.5 76.2 61.705 ;
      RECT  79.32 61.5 79.11 61.705 ;
      RECT  79.53 60.79 79.32 61.12 ;
      RECT  77.49 60.79 77.31 61.705 ;
      RECT  78.93 60.79 78.75 61.705 ;
      POLYGON  76.485 60.79 76.485 61.12 76.92 61.12 76.92 61.5 76.485 61.5 76.485 61.705 76.41 61.705 76.41 60.79 76.485 60.79 ;
      RECT  78.21 61.705 78.03 63.41 ;
      RECT  76.485 64.865 76.41 63.16 ;
      RECT  76.41 65.45 76.2 65.07 ;
      RECT  78.57 65.78 78.39 64.865 ;
      POLYGON  76.92 64.775 76.92 64.365 76.745 64.365 76.665 64.445 76.665 64.775 76.92 64.775 ;
      RECT  78.93 64.865 78.75 63.16 ;
      RECT  78.57 64.865 78.39 63.16 ;
      RECT  79.32 64.865 79.11 63.16 ;
      RECT  79.53 65.07 79.32 64.865 ;
      RECT  79.53 64.865 79.32 63.16 ;
      RECT  76.41 64.865 76.2 63.16 ;
      POLYGON  76.92 63.785 76.92 63.375 76.665 63.375 76.665 63.705 76.745 63.785 76.92 63.785 ;
      RECT  79.32 65.45 79.11 65.07 ;
      RECT  76.41 65.78 76.2 65.45 ;
      RECT  78.21 65.78 78.03 64.865 ;
      RECT  76.57 64.28 76.485 63.87 ;
      RECT  77.49 64.865 77.31 63.16 ;
      RECT  77.13 63.785 76.92 63.375 ;
      RECT  79.32 65.78 79.11 65.45 ;
      RECT  77.13 64.775 76.92 64.365 ;
      RECT  77.13 65.45 76.92 65.07 ;
      RECT  79.53 65.45 79.32 65.07 ;
      RECT  77.85 65.78 77.67 64.865 ;
      RECT  77.85 64.865 77.67 63.16 ;
      RECT  76.41 65.07 76.2 64.865 ;
      RECT  79.32 65.07 79.11 64.865 ;
      RECT  79.53 65.78 79.32 65.45 ;
      RECT  77.49 65.78 77.31 64.865 ;
      RECT  78.93 65.78 78.75 64.865 ;
      POLYGON  76.485 65.78 76.485 65.45 76.92 65.45 76.92 65.07 76.485 65.07 76.485 64.865 76.41 64.865 76.41 65.78 76.485 65.78 ;
      RECT  78.21 64.865 78.03 63.16 ;
      RECT  76.485 65.655 76.41 67.36 ;
      RECT  76.41 65.07 76.2 65.45 ;
      RECT  78.57 64.74 78.39 65.655 ;
      POLYGON  76.92 65.745 76.92 66.155 76.745 66.155 76.665 66.075 76.665 65.745 76.92 65.745 ;
      RECT  78.93 65.655 78.75 67.36 ;
      RECT  78.57 65.655 78.39 67.36 ;
      RECT  79.32 65.655 79.11 67.36 ;
      RECT  79.53 65.45 79.32 65.655 ;
      RECT  79.53 65.655 79.32 67.36 ;
      RECT  76.41 65.655 76.2 67.36 ;
      POLYGON  76.92 66.735 76.92 67.145 76.665 67.145 76.665 66.815 76.745 66.735 76.92 66.735 ;
      RECT  79.32 65.07 79.11 65.45 ;
      RECT  76.41 64.74 76.2 65.07 ;
      RECT  78.21 64.74 78.03 65.655 ;
      RECT  76.57 66.24 76.485 66.65 ;
      RECT  77.49 65.655 77.31 67.36 ;
      RECT  77.13 66.735 76.92 67.145 ;
      RECT  79.32 64.74 79.11 65.07 ;
      RECT  77.13 65.745 76.92 66.155 ;
      RECT  77.13 65.07 76.92 65.45 ;
      RECT  79.53 65.07 79.32 65.45 ;
      RECT  77.85 64.74 77.67 65.655 ;
      RECT  77.85 65.655 77.67 67.36 ;
      RECT  76.41 65.45 76.2 65.655 ;
      RECT  79.32 65.45 79.11 65.655 ;
      RECT  79.53 64.74 79.32 65.07 ;
      RECT  77.49 64.74 77.31 65.655 ;
      RECT  78.93 64.74 78.75 65.655 ;
      POLYGON  76.485 64.74 76.485 65.07 76.92 65.07 76.92 65.45 76.485 65.45 76.485 65.655 76.41 65.655 76.41 64.74 76.485 64.74 ;
      RECT  78.21 65.655 78.03 67.36 ;
      RECT  76.485 68.815 76.41 67.11 ;
      RECT  76.41 69.4 76.2 69.02 ;
      RECT  78.57 69.73 78.39 68.815 ;
      POLYGON  76.92 68.725 76.92 68.315 76.745 68.315 76.665 68.395 76.665 68.725 76.92 68.725 ;
      RECT  78.93 68.815 78.75 67.11 ;
      RECT  78.57 68.815 78.39 67.11 ;
      RECT  79.32 68.815 79.11 67.11 ;
      RECT  79.53 69.02 79.32 68.815 ;
      RECT  79.53 68.815 79.32 67.11 ;
      RECT  76.41 68.815 76.2 67.11 ;
      POLYGON  76.92 67.735 76.92 67.325 76.665 67.325 76.665 67.655 76.745 67.735 76.92 67.735 ;
      RECT  79.32 69.4 79.11 69.02 ;
      RECT  76.41 69.73 76.2 69.4 ;
      RECT  78.21 69.73 78.03 68.815 ;
      RECT  76.57 68.23 76.485 67.82 ;
      RECT  77.49 68.815 77.31 67.11 ;
      RECT  77.13 67.735 76.92 67.325 ;
      RECT  79.32 69.73 79.11 69.4 ;
      RECT  77.13 68.725 76.92 68.315 ;
      RECT  77.13 69.4 76.92 69.02 ;
      RECT  79.53 69.4 79.32 69.02 ;
      RECT  77.85 69.73 77.67 68.815 ;
      RECT  77.85 68.815 77.67 67.11 ;
      RECT  76.41 69.02 76.2 68.815 ;
      RECT  79.32 69.02 79.11 68.815 ;
      RECT  79.53 69.73 79.32 69.4 ;
      RECT  77.49 69.73 77.31 68.815 ;
      RECT  78.93 69.73 78.75 68.815 ;
      POLYGON  76.485 69.73 76.485 69.4 76.92 69.4 76.92 69.02 76.485 69.02 76.485 68.815 76.41 68.815 76.41 69.73 76.485 69.73 ;
      RECT  78.21 68.815 78.03 67.11 ;
      RECT  76.485 69.605 76.41 71.31 ;
      RECT  76.41 69.02 76.2 69.4 ;
      RECT  78.57 68.69 78.39 69.605 ;
      POLYGON  76.92 69.695 76.92 70.105 76.745 70.105 76.665 70.025 76.665 69.695 76.92 69.695 ;
      RECT  78.93 69.605 78.75 71.31 ;
      RECT  78.57 69.605 78.39 71.31 ;
      RECT  79.32 69.605 79.11 71.31 ;
      RECT  79.53 69.4 79.32 69.605 ;
      RECT  79.53 69.605 79.32 71.31 ;
      RECT  76.41 69.605 76.2 71.31 ;
      POLYGON  76.92 70.685 76.92 71.095 76.665 71.095 76.665 70.765 76.745 70.685 76.92 70.685 ;
      RECT  79.32 69.02 79.11 69.4 ;
      RECT  76.41 68.69 76.2 69.02 ;
      RECT  78.21 68.69 78.03 69.605 ;
      RECT  76.57 70.19 76.485 70.6 ;
      RECT  77.49 69.605 77.31 71.31 ;
      RECT  77.13 70.685 76.92 71.095 ;
      RECT  79.32 68.69 79.11 69.02 ;
      RECT  77.13 69.695 76.92 70.105 ;
      RECT  77.13 69.02 76.92 69.4 ;
      RECT  79.53 69.02 79.32 69.4 ;
      RECT  77.85 68.69 77.67 69.605 ;
      RECT  77.85 69.605 77.67 71.31 ;
      RECT  76.41 69.4 76.2 69.605 ;
      RECT  79.32 69.4 79.11 69.605 ;
      RECT  79.53 68.69 79.32 69.02 ;
      RECT  77.49 68.69 77.31 69.605 ;
      RECT  78.93 68.69 78.75 69.605 ;
      POLYGON  76.485 68.69 76.485 69.02 76.92 69.02 76.92 69.4 76.485 69.4 76.485 69.605 76.41 69.605 76.41 68.69 76.485 68.69 ;
      RECT  78.21 69.605 78.03 71.31 ;
      RECT  76.485 72.765 76.41 71.06 ;
      RECT  76.41 73.35 76.2 72.97 ;
      RECT  78.57 73.68 78.39 72.765 ;
      POLYGON  76.92 72.675 76.92 72.265 76.745 72.265 76.665 72.345 76.665 72.675 76.92 72.675 ;
      RECT  78.93 72.765 78.75 71.06 ;
      RECT  78.57 72.765 78.39 71.06 ;
      RECT  79.32 72.765 79.11 71.06 ;
      RECT  79.53 72.97 79.32 72.765 ;
      RECT  79.53 72.765 79.32 71.06 ;
      RECT  76.41 72.765 76.2 71.06 ;
      POLYGON  76.92 71.685 76.92 71.275 76.665 71.275 76.665 71.605 76.745 71.685 76.92 71.685 ;
      RECT  79.32 73.35 79.11 72.97 ;
      RECT  76.41 73.68 76.2 73.35 ;
      RECT  78.21 73.68 78.03 72.765 ;
      RECT  76.57 72.18 76.485 71.77 ;
      RECT  77.49 72.765 77.31 71.06 ;
      RECT  77.13 71.685 76.92 71.275 ;
      RECT  79.32 73.68 79.11 73.35 ;
      RECT  77.13 72.675 76.92 72.265 ;
      RECT  77.13 73.35 76.92 72.97 ;
      RECT  79.53 73.35 79.32 72.97 ;
      RECT  77.85 73.68 77.67 72.765 ;
      RECT  77.85 72.765 77.67 71.06 ;
      RECT  76.41 72.97 76.2 72.765 ;
      RECT  79.32 72.97 79.11 72.765 ;
      RECT  79.53 73.68 79.32 73.35 ;
      RECT  77.49 73.68 77.31 72.765 ;
      RECT  78.93 73.68 78.75 72.765 ;
      POLYGON  76.485 73.68 76.485 73.35 76.92 73.35 76.92 72.97 76.485 72.97 76.485 72.765 76.41 72.765 76.41 73.68 76.485 73.68 ;
      RECT  78.21 72.765 78.03 71.06 ;
      RECT  76.485 73.555 76.41 75.26 ;
      RECT  76.41 72.97 76.2 73.35 ;
      RECT  78.57 72.64 78.39 73.555 ;
      POLYGON  76.92 73.645 76.92 74.055 76.745 74.055 76.665 73.975 76.665 73.645 76.92 73.645 ;
      RECT  78.93 73.555 78.75 75.26 ;
      RECT  78.57 73.555 78.39 75.26 ;
      RECT  79.32 73.555 79.11 75.26 ;
      RECT  79.53 73.35 79.32 73.555 ;
      RECT  79.53 73.555 79.32 75.26 ;
      RECT  76.41 73.555 76.2 75.26 ;
      POLYGON  76.92 74.635 76.92 75.045 76.665 75.045 76.665 74.715 76.745 74.635 76.92 74.635 ;
      RECT  79.32 72.97 79.11 73.35 ;
      RECT  76.41 72.64 76.2 72.97 ;
      RECT  78.21 72.64 78.03 73.555 ;
      RECT  76.57 74.14 76.485 74.55 ;
      RECT  77.49 73.555 77.31 75.26 ;
      RECT  77.13 74.635 76.92 75.045 ;
      RECT  79.32 72.64 79.11 72.97 ;
      RECT  77.13 73.645 76.92 74.055 ;
      RECT  77.13 72.97 76.92 73.35 ;
      RECT  79.53 72.97 79.32 73.35 ;
      RECT  77.85 72.64 77.67 73.555 ;
      RECT  77.85 73.555 77.67 75.26 ;
      RECT  76.41 73.35 76.2 73.555 ;
      RECT  79.32 73.35 79.11 73.555 ;
      RECT  79.53 72.64 79.32 72.97 ;
      RECT  77.49 72.64 77.31 73.555 ;
      RECT  78.93 72.64 78.75 73.555 ;
      POLYGON  76.485 72.64 76.485 72.97 76.92 72.97 76.92 73.35 76.485 73.35 76.485 73.555 76.41 73.555 76.41 72.64 76.485 72.64 ;
      RECT  78.21 73.555 78.03 75.26 ;
      RECT  76.485 76.715 76.41 75.01 ;
      RECT  76.41 77.3 76.2 76.92 ;
      RECT  78.57 77.63 78.39 76.715 ;
      POLYGON  76.92 76.625 76.92 76.215 76.745 76.215 76.665 76.295 76.665 76.625 76.92 76.625 ;
      RECT  78.93 76.715 78.75 75.01 ;
      RECT  78.57 76.715 78.39 75.01 ;
      RECT  79.32 76.715 79.11 75.01 ;
      RECT  79.53 76.92 79.32 76.715 ;
      RECT  79.53 76.715 79.32 75.01 ;
      RECT  76.41 76.715 76.2 75.01 ;
      POLYGON  76.92 75.635 76.92 75.225 76.665 75.225 76.665 75.555 76.745 75.635 76.92 75.635 ;
      RECT  79.32 77.3 79.11 76.92 ;
      RECT  76.41 77.63 76.2 77.3 ;
      RECT  78.21 77.63 78.03 76.715 ;
      RECT  76.57 76.13 76.485 75.72 ;
      RECT  77.49 76.715 77.31 75.01 ;
      RECT  77.13 75.635 76.92 75.225 ;
      RECT  79.32 77.63 79.11 77.3 ;
      RECT  77.13 76.625 76.92 76.215 ;
      RECT  77.13 77.3 76.92 76.92 ;
      RECT  79.53 77.3 79.32 76.92 ;
      RECT  77.85 77.63 77.67 76.715 ;
      RECT  77.85 76.715 77.67 75.01 ;
      RECT  76.41 76.92 76.2 76.715 ;
      RECT  79.32 76.92 79.11 76.715 ;
      RECT  79.53 77.63 79.32 77.3 ;
      RECT  77.49 77.63 77.31 76.715 ;
      RECT  78.93 77.63 78.75 76.715 ;
      POLYGON  76.485 77.63 76.485 77.3 76.92 77.3 76.92 76.92 76.485 76.92 76.485 76.715 76.41 76.715 76.41 77.63 76.485 77.63 ;
      RECT  78.21 76.715 78.03 75.01 ;
      RECT  76.485 77.505 76.41 79.21 ;
      RECT  76.41 76.92 76.2 77.3 ;
      RECT  78.57 76.59 78.39 77.505 ;
      POLYGON  76.92 77.595 76.92 78.005 76.745 78.005 76.665 77.925 76.665 77.595 76.92 77.595 ;
      RECT  78.93 77.505 78.75 79.21 ;
      RECT  78.57 77.505 78.39 79.21 ;
      RECT  79.32 77.505 79.11 79.21 ;
      RECT  79.53 77.3 79.32 77.505 ;
      RECT  79.53 77.505 79.32 79.21 ;
      RECT  76.41 77.505 76.2 79.21 ;
      POLYGON  76.92 78.585 76.92 78.995 76.665 78.995 76.665 78.665 76.745 78.585 76.92 78.585 ;
      RECT  79.32 76.92 79.11 77.3 ;
      RECT  76.41 76.59 76.2 76.92 ;
      RECT  78.21 76.59 78.03 77.505 ;
      RECT  76.57 78.09 76.485 78.5 ;
      RECT  77.49 77.505 77.31 79.21 ;
      RECT  77.13 78.585 76.92 78.995 ;
      RECT  79.32 76.59 79.11 76.92 ;
      RECT  77.13 77.595 76.92 78.005 ;
      RECT  77.13 76.92 76.92 77.3 ;
      RECT  79.53 76.92 79.32 77.3 ;
      RECT  77.85 76.59 77.67 77.505 ;
      RECT  77.85 77.505 77.67 79.21 ;
      RECT  76.41 77.3 76.2 77.505 ;
      RECT  79.32 77.3 79.11 77.505 ;
      RECT  79.53 76.59 79.32 76.92 ;
      RECT  77.49 76.59 77.31 77.505 ;
      RECT  78.93 76.59 78.75 77.505 ;
      POLYGON  76.485 76.59 76.485 76.92 76.92 76.92 76.92 77.3 76.485 77.3 76.485 77.505 76.41 77.505 76.41 76.59 76.485 76.59 ;
      RECT  78.21 77.505 78.03 79.21 ;
      RECT  76.485 80.665 76.41 78.96 ;
      RECT  76.41 81.25 76.2 80.87 ;
      RECT  78.57 81.58 78.39 80.665 ;
      POLYGON  76.92 80.575 76.92 80.165 76.745 80.165 76.665 80.245 76.665 80.575 76.92 80.575 ;
      RECT  78.93 80.665 78.75 78.96 ;
      RECT  78.57 80.665 78.39 78.96 ;
      RECT  79.32 80.665 79.11 78.96 ;
      RECT  79.53 80.87 79.32 80.665 ;
      RECT  79.53 80.665 79.32 78.96 ;
      RECT  76.41 80.665 76.2 78.96 ;
      POLYGON  76.92 79.585 76.92 79.175 76.665 79.175 76.665 79.505 76.745 79.585 76.92 79.585 ;
      RECT  79.32 81.25 79.11 80.87 ;
      RECT  76.41 81.58 76.2 81.25 ;
      RECT  78.21 81.58 78.03 80.665 ;
      RECT  76.57 80.08 76.485 79.67 ;
      RECT  77.49 80.665 77.31 78.96 ;
      RECT  77.13 79.585 76.92 79.175 ;
      RECT  79.32 81.58 79.11 81.25 ;
      RECT  77.13 80.575 76.92 80.165 ;
      RECT  77.13 81.25 76.92 80.87 ;
      RECT  79.53 81.25 79.32 80.87 ;
      RECT  77.85 81.58 77.67 80.665 ;
      RECT  77.85 80.665 77.67 78.96 ;
      RECT  76.41 80.87 76.2 80.665 ;
      RECT  79.32 80.87 79.11 80.665 ;
      RECT  79.53 81.58 79.32 81.25 ;
      RECT  77.49 81.58 77.31 80.665 ;
      RECT  78.93 81.58 78.75 80.665 ;
      POLYGON  76.485 81.58 76.485 81.25 76.92 81.25 76.92 80.87 76.485 80.87 76.485 80.665 76.41 80.665 76.41 81.58 76.485 81.58 ;
      RECT  78.21 80.665 78.03 78.96 ;
      RECT  76.485 81.455 76.41 83.16 ;
      RECT  76.41 80.87 76.2 81.25 ;
      RECT  78.57 80.54 78.39 81.455 ;
      POLYGON  76.92 81.545 76.92 81.955 76.745 81.955 76.665 81.875 76.665 81.545 76.92 81.545 ;
      RECT  78.93 81.455 78.75 83.16 ;
      RECT  78.57 81.455 78.39 83.16 ;
      RECT  79.32 81.455 79.11 83.16 ;
      RECT  79.53 81.25 79.32 81.455 ;
      RECT  79.53 81.455 79.32 83.16 ;
      RECT  76.41 81.455 76.2 83.16 ;
      POLYGON  76.92 82.535 76.92 82.945 76.665 82.945 76.665 82.615 76.745 82.535 76.92 82.535 ;
      RECT  79.32 80.87 79.11 81.25 ;
      RECT  76.41 80.54 76.2 80.87 ;
      RECT  78.21 80.54 78.03 81.455 ;
      RECT  76.57 82.04 76.485 82.45 ;
      RECT  77.49 81.455 77.31 83.16 ;
      RECT  77.13 82.535 76.92 82.945 ;
      RECT  79.32 80.54 79.11 80.87 ;
      RECT  77.13 81.545 76.92 81.955 ;
      RECT  77.13 80.87 76.92 81.25 ;
      RECT  79.53 80.87 79.32 81.25 ;
      RECT  77.85 80.54 77.67 81.455 ;
      RECT  77.85 81.455 77.67 83.16 ;
      RECT  76.41 81.25 76.2 81.455 ;
      RECT  79.32 81.25 79.11 81.455 ;
      RECT  79.53 80.54 79.32 80.87 ;
      RECT  77.49 80.54 77.31 81.455 ;
      RECT  78.93 80.54 78.75 81.455 ;
      POLYGON  76.485 80.54 76.485 80.87 76.92 80.87 76.92 81.25 76.485 81.25 76.485 81.455 76.41 81.455 76.41 80.54 76.485 80.54 ;
      RECT  78.21 81.455 78.03 83.16 ;
      RECT  76.485 84.615 76.41 82.91 ;
      RECT  76.41 85.2 76.2 84.82 ;
      RECT  78.57 85.53 78.39 84.615 ;
      POLYGON  76.92 84.525 76.92 84.115 76.745 84.115 76.665 84.195 76.665 84.525 76.92 84.525 ;
      RECT  78.93 84.615 78.75 82.91 ;
      RECT  78.57 84.615 78.39 82.91 ;
      RECT  79.32 84.615 79.11 82.91 ;
      RECT  79.53 84.82 79.32 84.615 ;
      RECT  79.53 84.615 79.32 82.91 ;
      RECT  76.41 84.615 76.2 82.91 ;
      POLYGON  76.92 83.535 76.92 83.125 76.665 83.125 76.665 83.455 76.745 83.535 76.92 83.535 ;
      RECT  79.32 85.2 79.11 84.82 ;
      RECT  76.41 85.53 76.2 85.2 ;
      RECT  78.21 85.53 78.03 84.615 ;
      RECT  76.57 84.03 76.485 83.62 ;
      RECT  77.49 84.615 77.31 82.91 ;
      RECT  77.13 83.535 76.92 83.125 ;
      RECT  79.32 85.53 79.11 85.2 ;
      RECT  77.13 84.525 76.92 84.115 ;
      RECT  77.13 85.2 76.92 84.82 ;
      RECT  79.53 85.2 79.32 84.82 ;
      RECT  77.85 85.53 77.67 84.615 ;
      RECT  77.85 84.615 77.67 82.91 ;
      RECT  76.41 84.82 76.2 84.615 ;
      RECT  79.32 84.82 79.11 84.615 ;
      RECT  79.53 85.53 79.32 85.2 ;
      RECT  77.49 85.53 77.31 84.615 ;
      RECT  78.93 85.53 78.75 84.615 ;
      POLYGON  76.485 85.53 76.485 85.2 76.92 85.2 76.92 84.82 76.485 84.82 76.485 84.615 76.41 84.615 76.41 85.53 76.485 85.53 ;
      RECT  78.21 84.615 78.03 82.91 ;
      RECT  76.485 85.405 76.41 87.11 ;
      RECT  76.41 84.82 76.2 85.2 ;
      RECT  78.57 84.49 78.39 85.405 ;
      POLYGON  76.92 85.495 76.92 85.905 76.745 85.905 76.665 85.825 76.665 85.495 76.92 85.495 ;
      RECT  78.93 85.405 78.75 87.11 ;
      RECT  78.57 85.405 78.39 87.11 ;
      RECT  79.32 85.405 79.11 87.11 ;
      RECT  79.53 85.2 79.32 85.405 ;
      RECT  79.53 85.405 79.32 87.11 ;
      RECT  76.41 85.405 76.2 87.11 ;
      POLYGON  76.92 86.485 76.92 86.895 76.665 86.895 76.665 86.565 76.745 86.485 76.92 86.485 ;
      RECT  79.32 84.82 79.11 85.2 ;
      RECT  76.41 84.49 76.2 84.82 ;
      RECT  78.21 84.49 78.03 85.405 ;
      RECT  76.57 85.99 76.485 86.4 ;
      RECT  77.49 85.405 77.31 87.11 ;
      RECT  77.13 86.485 76.92 86.895 ;
      RECT  79.32 84.49 79.11 84.82 ;
      RECT  77.13 85.495 76.92 85.905 ;
      RECT  77.13 84.82 76.92 85.2 ;
      RECT  79.53 84.82 79.32 85.2 ;
      RECT  77.85 84.49 77.67 85.405 ;
      RECT  77.85 85.405 77.67 87.11 ;
      RECT  76.41 85.2 76.2 85.405 ;
      RECT  79.32 85.2 79.11 85.405 ;
      RECT  79.53 84.49 79.32 84.82 ;
      RECT  77.49 84.49 77.31 85.405 ;
      RECT  78.93 84.49 78.75 85.405 ;
      POLYGON  76.485 84.49 76.485 84.82 76.92 84.82 76.92 85.2 76.485 85.2 76.485 85.405 76.41 85.405 76.41 84.49 76.485 84.49 ;
      RECT  78.21 85.405 78.03 87.11 ;
      RECT  76.485 88.565 76.41 86.86 ;
      RECT  76.41 89.15 76.2 88.77 ;
      RECT  78.57 89.48 78.39 88.565 ;
      POLYGON  76.92 88.475 76.92 88.065 76.745 88.065 76.665 88.145 76.665 88.475 76.92 88.475 ;
      RECT  78.93 88.565 78.75 86.86 ;
      RECT  78.57 88.565 78.39 86.86 ;
      RECT  79.32 88.565 79.11 86.86 ;
      RECT  79.53 88.77 79.32 88.565 ;
      RECT  79.53 88.565 79.32 86.86 ;
      RECT  76.41 88.565 76.2 86.86 ;
      POLYGON  76.92 87.485 76.92 87.075 76.665 87.075 76.665 87.405 76.745 87.485 76.92 87.485 ;
      RECT  79.32 89.15 79.11 88.77 ;
      RECT  76.41 89.48 76.2 89.15 ;
      RECT  78.21 89.48 78.03 88.565 ;
      RECT  76.57 87.98 76.485 87.57 ;
      RECT  77.49 88.565 77.31 86.86 ;
      RECT  77.13 87.485 76.92 87.075 ;
      RECT  79.32 89.48 79.11 89.15 ;
      RECT  77.13 88.475 76.92 88.065 ;
      RECT  77.13 89.15 76.92 88.77 ;
      RECT  79.53 89.15 79.32 88.77 ;
      RECT  77.85 89.48 77.67 88.565 ;
      RECT  77.85 88.565 77.67 86.86 ;
      RECT  76.41 88.77 76.2 88.565 ;
      RECT  79.32 88.77 79.11 88.565 ;
      RECT  79.53 89.48 79.32 89.15 ;
      RECT  77.49 89.48 77.31 88.565 ;
      RECT  78.93 89.48 78.75 88.565 ;
      POLYGON  76.485 89.48 76.485 89.15 76.92 89.15 76.92 88.77 76.485 88.77 76.485 88.565 76.41 88.565 76.41 89.48 76.485 89.48 ;
      RECT  78.21 88.565 78.03 86.86 ;
      RECT  76.485 89.355 76.41 91.06 ;
      RECT  76.41 88.77 76.2 89.15 ;
      RECT  78.57 88.44 78.39 89.355 ;
      POLYGON  76.92 89.445 76.92 89.855 76.745 89.855 76.665 89.775 76.665 89.445 76.92 89.445 ;
      RECT  78.93 89.355 78.75 91.06 ;
      RECT  78.57 89.355 78.39 91.06 ;
      RECT  79.32 89.355 79.11 91.06 ;
      RECT  79.53 89.15 79.32 89.355 ;
      RECT  79.53 89.355 79.32 91.06 ;
      RECT  76.41 89.355 76.2 91.06 ;
      POLYGON  76.92 90.435 76.92 90.845 76.665 90.845 76.665 90.515 76.745 90.435 76.92 90.435 ;
      RECT  79.32 88.77 79.11 89.15 ;
      RECT  76.41 88.44 76.2 88.77 ;
      RECT  78.21 88.44 78.03 89.355 ;
      RECT  76.57 89.94 76.485 90.35 ;
      RECT  77.49 89.355 77.31 91.06 ;
      RECT  77.13 90.435 76.92 90.845 ;
      RECT  79.32 88.44 79.11 88.77 ;
      RECT  77.13 89.445 76.92 89.855 ;
      RECT  77.13 88.77 76.92 89.15 ;
      RECT  79.53 88.77 79.32 89.15 ;
      RECT  77.85 88.44 77.67 89.355 ;
      RECT  77.85 89.355 77.67 91.06 ;
      RECT  76.41 89.15 76.2 89.355 ;
      RECT  79.32 89.15 79.11 89.355 ;
      RECT  79.53 88.44 79.32 88.77 ;
      RECT  77.49 88.44 77.31 89.355 ;
      RECT  78.93 88.44 78.75 89.355 ;
      POLYGON  76.485 88.44 76.485 88.77 76.92 88.77 76.92 89.15 76.485 89.15 76.485 89.355 76.41 89.355 76.41 88.44 76.485 88.44 ;
      RECT  78.21 89.355 78.03 91.06 ;
      RECT  76.485 92.515 76.41 90.81 ;
      RECT  76.41 93.1 76.2 92.72 ;
      RECT  78.57 93.43 78.39 92.515 ;
      POLYGON  76.92 92.425 76.92 92.015 76.745 92.015 76.665 92.095 76.665 92.425 76.92 92.425 ;
      RECT  78.93 92.515 78.75 90.81 ;
      RECT  78.57 92.515 78.39 90.81 ;
      RECT  79.32 92.515 79.11 90.81 ;
      RECT  79.53 92.72 79.32 92.515 ;
      RECT  79.53 92.515 79.32 90.81 ;
      RECT  76.41 92.515 76.2 90.81 ;
      POLYGON  76.92 91.435 76.92 91.025 76.665 91.025 76.665 91.355 76.745 91.435 76.92 91.435 ;
      RECT  79.32 93.1 79.11 92.72 ;
      RECT  76.41 93.43 76.2 93.1 ;
      RECT  78.21 93.43 78.03 92.515 ;
      RECT  76.57 91.93 76.485 91.52 ;
      RECT  77.49 92.515 77.31 90.81 ;
      RECT  77.13 91.435 76.92 91.025 ;
      RECT  79.32 93.43 79.11 93.1 ;
      RECT  77.13 92.425 76.92 92.015 ;
      RECT  77.13 93.1 76.92 92.72 ;
      RECT  79.53 93.1 79.32 92.72 ;
      RECT  77.85 93.43 77.67 92.515 ;
      RECT  77.85 92.515 77.67 90.81 ;
      RECT  76.41 92.72 76.2 92.515 ;
      RECT  79.32 92.72 79.11 92.515 ;
      RECT  79.53 93.43 79.32 93.1 ;
      RECT  77.49 93.43 77.31 92.515 ;
      RECT  78.93 93.43 78.75 92.515 ;
      POLYGON  76.485 93.43 76.485 93.1 76.92 93.1 76.92 92.72 76.485 92.72 76.485 92.515 76.41 92.515 76.41 93.43 76.485 93.43 ;
      RECT  78.21 92.515 78.03 90.81 ;
      RECT  73.47 61.31 73.65 92.91 ;
      RECT  73.83 61.31 74.01 92.91 ;
      RECT  74.55 61.31 74.73 92.91 ;
      RECT  74.91 61.31 75.09 92.91 ;
      RECT  78.75 61.31 78.93 92.91 ;
      RECT  78.39 61.31 78.57 92.91 ;
      RECT  77.67 61.31 77.85 92.91 ;
      RECT  77.31 61.31 77.49 92.91 ;
      RECT  74.19 90.81 74.37 92.515 ;
      RECT  74.19 82.91 74.37 84.615 ;
      RECT  74.19 61.705 74.37 63.41 ;
      RECT  74.19 67.11 74.37 68.815 ;
      RECT  74.19 71.06 74.37 72.765 ;
      RECT  78.03 82.91 78.21 84.615 ;
      RECT  74.19 89.355 74.37 91.06 ;
      RECT  74.19 85.405 74.37 87.11 ;
      RECT  74.19 73.555 74.37 75.26 ;
      RECT  74.19 86.86 74.37 88.565 ;
      RECT  74.19 63.16 74.37 64.865 ;
      RECT  74.19 75.01 74.37 76.715 ;
      RECT  78.03 61.705 78.21 63.41 ;
      RECT  78.03 75.01 78.21 76.715 ;
      RECT  78.03 73.555 78.21 75.26 ;
      RECT  78.03 89.355 78.21 91.06 ;
      RECT  74.19 78.96 74.37 80.665 ;
      RECT  74.19 69.605 74.37 71.31 ;
      RECT  78.03 86.86 78.21 88.565 ;
      RECT  78.03 90.81 78.21 92.515 ;
      RECT  78.03 63.16 78.21 64.865 ;
      RECT  78.03 81.455 78.21 83.16 ;
      RECT  78.03 65.655 78.21 67.36 ;
      RECT  78.03 67.11 78.21 68.815 ;
      RECT  78.03 71.06 78.21 72.765 ;
      RECT  78.03 77.505 78.21 79.21 ;
      RECT  74.19 81.455 74.37 83.16 ;
      RECT  78.03 69.605 78.21 71.31 ;
      RECT  78.03 85.405 78.21 87.11 ;
      RECT  74.19 77.505 74.37 79.21 ;
      RECT  74.19 65.655 74.37 67.36 ;
      RECT  78.03 78.96 78.21 80.665 ;
      RECT  71.97 58.15 71.79 59.73 ;
      RECT  72.33 58.15 72.15 59.73 ;
      RECT  71.88 58.15 71.75 58.86 ;
      RECT  71.61 58.15 71.43 59.73 ;
      RECT  72.01 58.15 71.88 58.86 ;
      RECT  72.33 57.36 72.15 58.15 ;
      RECT  72.69 57.36 72.51 58.15 ;
      RECT  71.25 57.36 71.07 58.15 ;
      RECT  71.97 57.36 71.79 58.15 ;
      RECT  71.61 57.36 71.43 58.15 ;
      RECT  72.69 58.15 72.51 59.73 ;
      RECT  71.25 58.15 71.07 59.73 ;
      RECT  70.245 60.915 70.17 59.21 ;
      RECT  70.17 61.5 69.96 61.12 ;
      RECT  72.33 61.83 72.15 60.915 ;
      POLYGON  70.68 60.825 70.68 60.415 70.505 60.415 70.425 60.495 70.425 60.825 70.68 60.825 ;
      RECT  72.69 60.915 72.51 59.21 ;
      RECT  72.33 60.915 72.15 59.21 ;
      RECT  73.08 60.915 72.87 59.21 ;
      RECT  73.29 61.12 73.08 60.915 ;
      RECT  73.29 60.915 73.08 59.21 ;
      RECT  70.17 60.915 69.96 59.21 ;
      POLYGON  70.68 59.835 70.68 59.425 70.425 59.425 70.425 59.755 70.505 59.835 70.68 59.835 ;
      RECT  73.08 61.5 72.87 61.12 ;
      RECT  70.17 61.83 69.96 61.5 ;
      RECT  71.97 61.83 71.79 60.915 ;
      RECT  70.33 60.33 70.245 59.92 ;
      RECT  71.25 60.915 71.07 59.21 ;
      RECT  70.89 59.835 70.68 59.425 ;
      RECT  73.08 61.83 72.87 61.5 ;
      RECT  70.89 60.825 70.68 60.415 ;
      RECT  70.89 61.5 70.68 61.12 ;
      RECT  73.29 61.5 73.08 61.12 ;
      RECT  71.61 61.83 71.43 60.915 ;
      RECT  71.61 60.915 71.43 59.21 ;
      RECT  70.17 61.12 69.96 60.915 ;
      RECT  73.08 61.12 72.87 60.915 ;
      RECT  73.29 61.83 73.08 61.5 ;
      RECT  71.25 61.83 71.07 60.915 ;
      RECT  72.69 61.83 72.51 60.915 ;
      POLYGON  70.245 61.83 70.245 61.5 70.68 61.5 70.68 61.12 70.245 61.12 70.245 60.915 70.17 60.915 70.17 61.83 70.245 61.83 ;
      RECT  71.97 60.915 71.79 59.21 ;
      RECT  70.245 61.705 70.17 63.41 ;
      RECT  70.17 61.12 69.96 61.5 ;
      RECT  72.33 60.79 72.15 61.705 ;
      POLYGON  70.68 61.795 70.68 62.205 70.505 62.205 70.425 62.125 70.425 61.795 70.68 61.795 ;
      RECT  72.69 61.705 72.51 63.41 ;
      RECT  72.33 61.705 72.15 63.41 ;
      RECT  73.08 61.705 72.87 63.41 ;
      RECT  73.29 61.5 73.08 61.705 ;
      RECT  73.29 61.705 73.08 63.41 ;
      RECT  70.17 61.705 69.96 63.41 ;
      POLYGON  70.68 62.785 70.68 63.195 70.425 63.195 70.425 62.865 70.505 62.785 70.68 62.785 ;
      RECT  73.08 61.12 72.87 61.5 ;
      RECT  70.17 60.79 69.96 61.12 ;
      RECT  71.97 60.79 71.79 61.705 ;
      RECT  70.33 62.29 70.245 62.7 ;
      RECT  71.25 61.705 71.07 63.41 ;
      RECT  70.89 62.785 70.68 63.195 ;
      RECT  73.08 60.79 72.87 61.12 ;
      RECT  70.89 61.795 70.68 62.205 ;
      RECT  70.89 61.12 70.68 61.5 ;
      RECT  73.29 61.12 73.08 61.5 ;
      RECT  71.61 60.79 71.43 61.705 ;
      RECT  71.61 61.705 71.43 63.41 ;
      RECT  70.17 61.5 69.96 61.705 ;
      RECT  73.08 61.5 72.87 61.705 ;
      RECT  73.29 60.79 73.08 61.12 ;
      RECT  71.25 60.79 71.07 61.705 ;
      RECT  72.69 60.79 72.51 61.705 ;
      POLYGON  70.245 60.79 70.245 61.12 70.68 61.12 70.68 61.5 70.245 61.5 70.245 61.705 70.17 61.705 70.17 60.79 70.245 60.79 ;
      RECT  71.97 61.705 71.79 63.41 ;
      RECT  70.245 64.865 70.17 63.16 ;
      RECT  70.17 65.45 69.96 65.07 ;
      RECT  72.33 65.78 72.15 64.865 ;
      POLYGON  70.68 64.775 70.68 64.365 70.505 64.365 70.425 64.445 70.425 64.775 70.68 64.775 ;
      RECT  72.69 64.865 72.51 63.16 ;
      RECT  72.33 64.865 72.15 63.16 ;
      RECT  73.08 64.865 72.87 63.16 ;
      RECT  73.29 65.07 73.08 64.865 ;
      RECT  73.29 64.865 73.08 63.16 ;
      RECT  70.17 64.865 69.96 63.16 ;
      POLYGON  70.68 63.785 70.68 63.375 70.425 63.375 70.425 63.705 70.505 63.785 70.68 63.785 ;
      RECT  73.08 65.45 72.87 65.07 ;
      RECT  70.17 65.78 69.96 65.45 ;
      RECT  71.97 65.78 71.79 64.865 ;
      RECT  70.33 64.28 70.245 63.87 ;
      RECT  71.25 64.865 71.07 63.16 ;
      RECT  70.89 63.785 70.68 63.375 ;
      RECT  73.08 65.78 72.87 65.45 ;
      RECT  70.89 64.775 70.68 64.365 ;
      RECT  70.89 65.45 70.68 65.07 ;
      RECT  73.29 65.45 73.08 65.07 ;
      RECT  71.61 65.78 71.43 64.865 ;
      RECT  71.61 64.865 71.43 63.16 ;
      RECT  70.17 65.07 69.96 64.865 ;
      RECT  73.08 65.07 72.87 64.865 ;
      RECT  73.29 65.78 73.08 65.45 ;
      RECT  71.25 65.78 71.07 64.865 ;
      RECT  72.69 65.78 72.51 64.865 ;
      POLYGON  70.245 65.78 70.245 65.45 70.68 65.45 70.68 65.07 70.245 65.07 70.245 64.865 70.17 64.865 70.17 65.78 70.245 65.78 ;
      RECT  71.97 64.865 71.79 63.16 ;
      RECT  70.245 65.655 70.17 67.36 ;
      RECT  70.17 65.07 69.96 65.45 ;
      RECT  72.33 64.74 72.15 65.655 ;
      POLYGON  70.68 65.745 70.68 66.155 70.505 66.155 70.425 66.075 70.425 65.745 70.68 65.745 ;
      RECT  72.69 65.655 72.51 67.36 ;
      RECT  72.33 65.655 72.15 67.36 ;
      RECT  73.08 65.655 72.87 67.36 ;
      RECT  73.29 65.45 73.08 65.655 ;
      RECT  73.29 65.655 73.08 67.36 ;
      RECT  70.17 65.655 69.96 67.36 ;
      POLYGON  70.68 66.735 70.68 67.145 70.425 67.145 70.425 66.815 70.505 66.735 70.68 66.735 ;
      RECT  73.08 65.07 72.87 65.45 ;
      RECT  70.17 64.74 69.96 65.07 ;
      RECT  71.97 64.74 71.79 65.655 ;
      RECT  70.33 66.24 70.245 66.65 ;
      RECT  71.25 65.655 71.07 67.36 ;
      RECT  70.89 66.735 70.68 67.145 ;
      RECT  73.08 64.74 72.87 65.07 ;
      RECT  70.89 65.745 70.68 66.155 ;
      RECT  70.89 65.07 70.68 65.45 ;
      RECT  73.29 65.07 73.08 65.45 ;
      RECT  71.61 64.74 71.43 65.655 ;
      RECT  71.61 65.655 71.43 67.36 ;
      RECT  70.17 65.45 69.96 65.655 ;
      RECT  73.08 65.45 72.87 65.655 ;
      RECT  73.29 64.74 73.08 65.07 ;
      RECT  71.25 64.74 71.07 65.655 ;
      RECT  72.69 64.74 72.51 65.655 ;
      POLYGON  70.245 64.74 70.245 65.07 70.68 65.07 70.68 65.45 70.245 65.45 70.245 65.655 70.17 65.655 70.17 64.74 70.245 64.74 ;
      RECT  71.97 65.655 71.79 67.36 ;
      RECT  70.245 68.815 70.17 67.11 ;
      RECT  70.17 69.4 69.96 69.02 ;
      RECT  72.33 69.73 72.15 68.815 ;
      POLYGON  70.68 68.725 70.68 68.315 70.505 68.315 70.425 68.395 70.425 68.725 70.68 68.725 ;
      RECT  72.69 68.815 72.51 67.11 ;
      RECT  72.33 68.815 72.15 67.11 ;
      RECT  73.08 68.815 72.87 67.11 ;
      RECT  73.29 69.02 73.08 68.815 ;
      RECT  73.29 68.815 73.08 67.11 ;
      RECT  70.17 68.815 69.96 67.11 ;
      POLYGON  70.68 67.735 70.68 67.325 70.425 67.325 70.425 67.655 70.505 67.735 70.68 67.735 ;
      RECT  73.08 69.4 72.87 69.02 ;
      RECT  70.17 69.73 69.96 69.4 ;
      RECT  71.97 69.73 71.79 68.815 ;
      RECT  70.33 68.23 70.245 67.82 ;
      RECT  71.25 68.815 71.07 67.11 ;
      RECT  70.89 67.735 70.68 67.325 ;
      RECT  73.08 69.73 72.87 69.4 ;
      RECT  70.89 68.725 70.68 68.315 ;
      RECT  70.89 69.4 70.68 69.02 ;
      RECT  73.29 69.4 73.08 69.02 ;
      RECT  71.61 69.73 71.43 68.815 ;
      RECT  71.61 68.815 71.43 67.11 ;
      RECT  70.17 69.02 69.96 68.815 ;
      RECT  73.08 69.02 72.87 68.815 ;
      RECT  73.29 69.73 73.08 69.4 ;
      RECT  71.25 69.73 71.07 68.815 ;
      RECT  72.69 69.73 72.51 68.815 ;
      POLYGON  70.245 69.73 70.245 69.4 70.68 69.4 70.68 69.02 70.245 69.02 70.245 68.815 70.17 68.815 70.17 69.73 70.245 69.73 ;
      RECT  71.97 68.815 71.79 67.11 ;
      RECT  70.245 69.605 70.17 71.31 ;
      RECT  70.17 69.02 69.96 69.4 ;
      RECT  72.33 68.69 72.15 69.605 ;
      POLYGON  70.68 69.695 70.68 70.105 70.505 70.105 70.425 70.025 70.425 69.695 70.68 69.695 ;
      RECT  72.69 69.605 72.51 71.31 ;
      RECT  72.33 69.605 72.15 71.31 ;
      RECT  73.08 69.605 72.87 71.31 ;
      RECT  73.29 69.4 73.08 69.605 ;
      RECT  73.29 69.605 73.08 71.31 ;
      RECT  70.17 69.605 69.96 71.31 ;
      POLYGON  70.68 70.685 70.68 71.095 70.425 71.095 70.425 70.765 70.505 70.685 70.68 70.685 ;
      RECT  73.08 69.02 72.87 69.4 ;
      RECT  70.17 68.69 69.96 69.02 ;
      RECT  71.97 68.69 71.79 69.605 ;
      RECT  70.33 70.19 70.245 70.6 ;
      RECT  71.25 69.605 71.07 71.31 ;
      RECT  70.89 70.685 70.68 71.095 ;
      RECT  73.08 68.69 72.87 69.02 ;
      RECT  70.89 69.695 70.68 70.105 ;
      RECT  70.89 69.02 70.68 69.4 ;
      RECT  73.29 69.02 73.08 69.4 ;
      RECT  71.61 68.69 71.43 69.605 ;
      RECT  71.61 69.605 71.43 71.31 ;
      RECT  70.17 69.4 69.96 69.605 ;
      RECT  73.08 69.4 72.87 69.605 ;
      RECT  73.29 68.69 73.08 69.02 ;
      RECT  71.25 68.69 71.07 69.605 ;
      RECT  72.69 68.69 72.51 69.605 ;
      POLYGON  70.245 68.69 70.245 69.02 70.68 69.02 70.68 69.4 70.245 69.4 70.245 69.605 70.17 69.605 70.17 68.69 70.245 68.69 ;
      RECT  71.97 69.605 71.79 71.31 ;
      RECT  70.245 72.765 70.17 71.06 ;
      RECT  70.17 73.35 69.96 72.97 ;
      RECT  72.33 73.68 72.15 72.765 ;
      POLYGON  70.68 72.675 70.68 72.265 70.505 72.265 70.425 72.345 70.425 72.675 70.68 72.675 ;
      RECT  72.69 72.765 72.51 71.06 ;
      RECT  72.33 72.765 72.15 71.06 ;
      RECT  73.08 72.765 72.87 71.06 ;
      RECT  73.29 72.97 73.08 72.765 ;
      RECT  73.29 72.765 73.08 71.06 ;
      RECT  70.17 72.765 69.96 71.06 ;
      POLYGON  70.68 71.685 70.68 71.275 70.425 71.275 70.425 71.605 70.505 71.685 70.68 71.685 ;
      RECT  73.08 73.35 72.87 72.97 ;
      RECT  70.17 73.68 69.96 73.35 ;
      RECT  71.97 73.68 71.79 72.765 ;
      RECT  70.33 72.18 70.245 71.77 ;
      RECT  71.25 72.765 71.07 71.06 ;
      RECT  70.89 71.685 70.68 71.275 ;
      RECT  73.08 73.68 72.87 73.35 ;
      RECT  70.89 72.675 70.68 72.265 ;
      RECT  70.89 73.35 70.68 72.97 ;
      RECT  73.29 73.35 73.08 72.97 ;
      RECT  71.61 73.68 71.43 72.765 ;
      RECT  71.61 72.765 71.43 71.06 ;
      RECT  70.17 72.97 69.96 72.765 ;
      RECT  73.08 72.97 72.87 72.765 ;
      RECT  73.29 73.68 73.08 73.35 ;
      RECT  71.25 73.68 71.07 72.765 ;
      RECT  72.69 73.68 72.51 72.765 ;
      POLYGON  70.245 73.68 70.245 73.35 70.68 73.35 70.68 72.97 70.245 72.97 70.245 72.765 70.17 72.765 70.17 73.68 70.245 73.68 ;
      RECT  71.97 72.765 71.79 71.06 ;
      RECT  70.245 73.555 70.17 75.26 ;
      RECT  70.17 72.97 69.96 73.35 ;
      RECT  72.33 72.64 72.15 73.555 ;
      POLYGON  70.68 73.645 70.68 74.055 70.505 74.055 70.425 73.975 70.425 73.645 70.68 73.645 ;
      RECT  72.69 73.555 72.51 75.26 ;
      RECT  72.33 73.555 72.15 75.26 ;
      RECT  73.08 73.555 72.87 75.26 ;
      RECT  73.29 73.35 73.08 73.555 ;
      RECT  73.29 73.555 73.08 75.26 ;
      RECT  70.17 73.555 69.96 75.26 ;
      POLYGON  70.68 74.635 70.68 75.045 70.425 75.045 70.425 74.715 70.505 74.635 70.68 74.635 ;
      RECT  73.08 72.97 72.87 73.35 ;
      RECT  70.17 72.64 69.96 72.97 ;
      RECT  71.97 72.64 71.79 73.555 ;
      RECT  70.33 74.14 70.245 74.55 ;
      RECT  71.25 73.555 71.07 75.26 ;
      RECT  70.89 74.635 70.68 75.045 ;
      RECT  73.08 72.64 72.87 72.97 ;
      RECT  70.89 73.645 70.68 74.055 ;
      RECT  70.89 72.97 70.68 73.35 ;
      RECT  73.29 72.97 73.08 73.35 ;
      RECT  71.61 72.64 71.43 73.555 ;
      RECT  71.61 73.555 71.43 75.26 ;
      RECT  70.17 73.35 69.96 73.555 ;
      RECT  73.08 73.35 72.87 73.555 ;
      RECT  73.29 72.64 73.08 72.97 ;
      RECT  71.25 72.64 71.07 73.555 ;
      RECT  72.69 72.64 72.51 73.555 ;
      POLYGON  70.245 72.64 70.245 72.97 70.68 72.97 70.68 73.35 70.245 73.35 70.245 73.555 70.17 73.555 70.17 72.64 70.245 72.64 ;
      RECT  71.97 73.555 71.79 75.26 ;
      RECT  70.245 76.715 70.17 75.01 ;
      RECT  70.17 77.3 69.96 76.92 ;
      RECT  72.33 77.63 72.15 76.715 ;
      POLYGON  70.68 76.625 70.68 76.215 70.505 76.215 70.425 76.295 70.425 76.625 70.68 76.625 ;
      RECT  72.69 76.715 72.51 75.01 ;
      RECT  72.33 76.715 72.15 75.01 ;
      RECT  73.08 76.715 72.87 75.01 ;
      RECT  73.29 76.92 73.08 76.715 ;
      RECT  73.29 76.715 73.08 75.01 ;
      RECT  70.17 76.715 69.96 75.01 ;
      POLYGON  70.68 75.635 70.68 75.225 70.425 75.225 70.425 75.555 70.505 75.635 70.68 75.635 ;
      RECT  73.08 77.3 72.87 76.92 ;
      RECT  70.17 77.63 69.96 77.3 ;
      RECT  71.97 77.63 71.79 76.715 ;
      RECT  70.33 76.13 70.245 75.72 ;
      RECT  71.25 76.715 71.07 75.01 ;
      RECT  70.89 75.635 70.68 75.225 ;
      RECT  73.08 77.63 72.87 77.3 ;
      RECT  70.89 76.625 70.68 76.215 ;
      RECT  70.89 77.3 70.68 76.92 ;
      RECT  73.29 77.3 73.08 76.92 ;
      RECT  71.61 77.63 71.43 76.715 ;
      RECT  71.61 76.715 71.43 75.01 ;
      RECT  70.17 76.92 69.96 76.715 ;
      RECT  73.08 76.92 72.87 76.715 ;
      RECT  73.29 77.63 73.08 77.3 ;
      RECT  71.25 77.63 71.07 76.715 ;
      RECT  72.69 77.63 72.51 76.715 ;
      POLYGON  70.245 77.63 70.245 77.3 70.68 77.3 70.68 76.92 70.245 76.92 70.245 76.715 70.17 76.715 70.17 77.63 70.245 77.63 ;
      RECT  71.97 76.715 71.79 75.01 ;
      RECT  70.245 77.505 70.17 79.21 ;
      RECT  70.17 76.92 69.96 77.3 ;
      RECT  72.33 76.59 72.15 77.505 ;
      POLYGON  70.68 77.595 70.68 78.005 70.505 78.005 70.425 77.925 70.425 77.595 70.68 77.595 ;
      RECT  72.69 77.505 72.51 79.21 ;
      RECT  72.33 77.505 72.15 79.21 ;
      RECT  73.08 77.505 72.87 79.21 ;
      RECT  73.29 77.3 73.08 77.505 ;
      RECT  73.29 77.505 73.08 79.21 ;
      RECT  70.17 77.505 69.96 79.21 ;
      POLYGON  70.68 78.585 70.68 78.995 70.425 78.995 70.425 78.665 70.505 78.585 70.68 78.585 ;
      RECT  73.08 76.92 72.87 77.3 ;
      RECT  70.17 76.59 69.96 76.92 ;
      RECT  71.97 76.59 71.79 77.505 ;
      RECT  70.33 78.09 70.245 78.5 ;
      RECT  71.25 77.505 71.07 79.21 ;
      RECT  70.89 78.585 70.68 78.995 ;
      RECT  73.08 76.59 72.87 76.92 ;
      RECT  70.89 77.595 70.68 78.005 ;
      RECT  70.89 76.92 70.68 77.3 ;
      RECT  73.29 76.92 73.08 77.3 ;
      RECT  71.61 76.59 71.43 77.505 ;
      RECT  71.61 77.505 71.43 79.21 ;
      RECT  70.17 77.3 69.96 77.505 ;
      RECT  73.08 77.3 72.87 77.505 ;
      RECT  73.29 76.59 73.08 76.92 ;
      RECT  71.25 76.59 71.07 77.505 ;
      RECT  72.69 76.59 72.51 77.505 ;
      POLYGON  70.245 76.59 70.245 76.92 70.68 76.92 70.68 77.3 70.245 77.3 70.245 77.505 70.17 77.505 70.17 76.59 70.245 76.59 ;
      RECT  71.97 77.505 71.79 79.21 ;
      RECT  70.245 80.665 70.17 78.96 ;
      RECT  70.17 81.25 69.96 80.87 ;
      RECT  72.33 81.58 72.15 80.665 ;
      POLYGON  70.68 80.575 70.68 80.165 70.505 80.165 70.425 80.245 70.425 80.575 70.68 80.575 ;
      RECT  72.69 80.665 72.51 78.96 ;
      RECT  72.33 80.665 72.15 78.96 ;
      RECT  73.08 80.665 72.87 78.96 ;
      RECT  73.29 80.87 73.08 80.665 ;
      RECT  73.29 80.665 73.08 78.96 ;
      RECT  70.17 80.665 69.96 78.96 ;
      POLYGON  70.68 79.585 70.68 79.175 70.425 79.175 70.425 79.505 70.505 79.585 70.68 79.585 ;
      RECT  73.08 81.25 72.87 80.87 ;
      RECT  70.17 81.58 69.96 81.25 ;
      RECT  71.97 81.58 71.79 80.665 ;
      RECT  70.33 80.08 70.245 79.67 ;
      RECT  71.25 80.665 71.07 78.96 ;
      RECT  70.89 79.585 70.68 79.175 ;
      RECT  73.08 81.58 72.87 81.25 ;
      RECT  70.89 80.575 70.68 80.165 ;
      RECT  70.89 81.25 70.68 80.87 ;
      RECT  73.29 81.25 73.08 80.87 ;
      RECT  71.61 81.58 71.43 80.665 ;
      RECT  71.61 80.665 71.43 78.96 ;
      RECT  70.17 80.87 69.96 80.665 ;
      RECT  73.08 80.87 72.87 80.665 ;
      RECT  73.29 81.58 73.08 81.25 ;
      RECT  71.25 81.58 71.07 80.665 ;
      RECT  72.69 81.58 72.51 80.665 ;
      POLYGON  70.245 81.58 70.245 81.25 70.68 81.25 70.68 80.87 70.245 80.87 70.245 80.665 70.17 80.665 70.17 81.58 70.245 81.58 ;
      RECT  71.97 80.665 71.79 78.96 ;
      RECT  70.245 81.455 70.17 83.16 ;
      RECT  70.17 80.87 69.96 81.25 ;
      RECT  72.33 80.54 72.15 81.455 ;
      POLYGON  70.68 81.545 70.68 81.955 70.505 81.955 70.425 81.875 70.425 81.545 70.68 81.545 ;
      RECT  72.69 81.455 72.51 83.16 ;
      RECT  72.33 81.455 72.15 83.16 ;
      RECT  73.08 81.455 72.87 83.16 ;
      RECT  73.29 81.25 73.08 81.455 ;
      RECT  73.29 81.455 73.08 83.16 ;
      RECT  70.17 81.455 69.96 83.16 ;
      POLYGON  70.68 82.535 70.68 82.945 70.425 82.945 70.425 82.615 70.505 82.535 70.68 82.535 ;
      RECT  73.08 80.87 72.87 81.25 ;
      RECT  70.17 80.54 69.96 80.87 ;
      RECT  71.97 80.54 71.79 81.455 ;
      RECT  70.33 82.04 70.245 82.45 ;
      RECT  71.25 81.455 71.07 83.16 ;
      RECT  70.89 82.535 70.68 82.945 ;
      RECT  73.08 80.54 72.87 80.87 ;
      RECT  70.89 81.545 70.68 81.955 ;
      RECT  70.89 80.87 70.68 81.25 ;
      RECT  73.29 80.87 73.08 81.25 ;
      RECT  71.61 80.54 71.43 81.455 ;
      RECT  71.61 81.455 71.43 83.16 ;
      RECT  70.17 81.25 69.96 81.455 ;
      RECT  73.08 81.25 72.87 81.455 ;
      RECT  73.29 80.54 73.08 80.87 ;
      RECT  71.25 80.54 71.07 81.455 ;
      RECT  72.69 80.54 72.51 81.455 ;
      POLYGON  70.245 80.54 70.245 80.87 70.68 80.87 70.68 81.25 70.245 81.25 70.245 81.455 70.17 81.455 70.17 80.54 70.245 80.54 ;
      RECT  71.97 81.455 71.79 83.16 ;
      RECT  70.245 84.615 70.17 82.91 ;
      RECT  70.17 85.2 69.96 84.82 ;
      RECT  72.33 85.53 72.15 84.615 ;
      POLYGON  70.68 84.525 70.68 84.115 70.505 84.115 70.425 84.195 70.425 84.525 70.68 84.525 ;
      RECT  72.69 84.615 72.51 82.91 ;
      RECT  72.33 84.615 72.15 82.91 ;
      RECT  73.08 84.615 72.87 82.91 ;
      RECT  73.29 84.82 73.08 84.615 ;
      RECT  73.29 84.615 73.08 82.91 ;
      RECT  70.17 84.615 69.96 82.91 ;
      POLYGON  70.68 83.535 70.68 83.125 70.425 83.125 70.425 83.455 70.505 83.535 70.68 83.535 ;
      RECT  73.08 85.2 72.87 84.82 ;
      RECT  70.17 85.53 69.96 85.2 ;
      RECT  71.97 85.53 71.79 84.615 ;
      RECT  70.33 84.03 70.245 83.62 ;
      RECT  71.25 84.615 71.07 82.91 ;
      RECT  70.89 83.535 70.68 83.125 ;
      RECT  73.08 85.53 72.87 85.2 ;
      RECT  70.89 84.525 70.68 84.115 ;
      RECT  70.89 85.2 70.68 84.82 ;
      RECT  73.29 85.2 73.08 84.82 ;
      RECT  71.61 85.53 71.43 84.615 ;
      RECT  71.61 84.615 71.43 82.91 ;
      RECT  70.17 84.82 69.96 84.615 ;
      RECT  73.08 84.82 72.87 84.615 ;
      RECT  73.29 85.53 73.08 85.2 ;
      RECT  71.25 85.53 71.07 84.615 ;
      RECT  72.69 85.53 72.51 84.615 ;
      POLYGON  70.245 85.53 70.245 85.2 70.68 85.2 70.68 84.82 70.245 84.82 70.245 84.615 70.17 84.615 70.17 85.53 70.245 85.53 ;
      RECT  71.97 84.615 71.79 82.91 ;
      RECT  70.245 85.405 70.17 87.11 ;
      RECT  70.17 84.82 69.96 85.2 ;
      RECT  72.33 84.49 72.15 85.405 ;
      POLYGON  70.68 85.495 70.68 85.905 70.505 85.905 70.425 85.825 70.425 85.495 70.68 85.495 ;
      RECT  72.69 85.405 72.51 87.11 ;
      RECT  72.33 85.405 72.15 87.11 ;
      RECT  73.08 85.405 72.87 87.11 ;
      RECT  73.29 85.2 73.08 85.405 ;
      RECT  73.29 85.405 73.08 87.11 ;
      RECT  70.17 85.405 69.96 87.11 ;
      POLYGON  70.68 86.485 70.68 86.895 70.425 86.895 70.425 86.565 70.505 86.485 70.68 86.485 ;
      RECT  73.08 84.82 72.87 85.2 ;
      RECT  70.17 84.49 69.96 84.82 ;
      RECT  71.97 84.49 71.79 85.405 ;
      RECT  70.33 85.99 70.245 86.4 ;
      RECT  71.25 85.405 71.07 87.11 ;
      RECT  70.89 86.485 70.68 86.895 ;
      RECT  73.08 84.49 72.87 84.82 ;
      RECT  70.89 85.495 70.68 85.905 ;
      RECT  70.89 84.82 70.68 85.2 ;
      RECT  73.29 84.82 73.08 85.2 ;
      RECT  71.61 84.49 71.43 85.405 ;
      RECT  71.61 85.405 71.43 87.11 ;
      RECT  70.17 85.2 69.96 85.405 ;
      RECT  73.08 85.2 72.87 85.405 ;
      RECT  73.29 84.49 73.08 84.82 ;
      RECT  71.25 84.49 71.07 85.405 ;
      RECT  72.69 84.49 72.51 85.405 ;
      POLYGON  70.245 84.49 70.245 84.82 70.68 84.82 70.68 85.2 70.245 85.2 70.245 85.405 70.17 85.405 70.17 84.49 70.245 84.49 ;
      RECT  71.97 85.405 71.79 87.11 ;
      RECT  70.245 88.565 70.17 86.86 ;
      RECT  70.17 89.15 69.96 88.77 ;
      RECT  72.33 89.48 72.15 88.565 ;
      POLYGON  70.68 88.475 70.68 88.065 70.505 88.065 70.425 88.145 70.425 88.475 70.68 88.475 ;
      RECT  72.69 88.565 72.51 86.86 ;
      RECT  72.33 88.565 72.15 86.86 ;
      RECT  73.08 88.565 72.87 86.86 ;
      RECT  73.29 88.77 73.08 88.565 ;
      RECT  73.29 88.565 73.08 86.86 ;
      RECT  70.17 88.565 69.96 86.86 ;
      POLYGON  70.68 87.485 70.68 87.075 70.425 87.075 70.425 87.405 70.505 87.485 70.68 87.485 ;
      RECT  73.08 89.15 72.87 88.77 ;
      RECT  70.17 89.48 69.96 89.15 ;
      RECT  71.97 89.48 71.79 88.565 ;
      RECT  70.33 87.98 70.245 87.57 ;
      RECT  71.25 88.565 71.07 86.86 ;
      RECT  70.89 87.485 70.68 87.075 ;
      RECT  73.08 89.48 72.87 89.15 ;
      RECT  70.89 88.475 70.68 88.065 ;
      RECT  70.89 89.15 70.68 88.77 ;
      RECT  73.29 89.15 73.08 88.77 ;
      RECT  71.61 89.48 71.43 88.565 ;
      RECT  71.61 88.565 71.43 86.86 ;
      RECT  70.17 88.77 69.96 88.565 ;
      RECT  73.08 88.77 72.87 88.565 ;
      RECT  73.29 89.48 73.08 89.15 ;
      RECT  71.25 89.48 71.07 88.565 ;
      RECT  72.69 89.48 72.51 88.565 ;
      POLYGON  70.245 89.48 70.245 89.15 70.68 89.15 70.68 88.77 70.245 88.77 70.245 88.565 70.17 88.565 70.17 89.48 70.245 89.48 ;
      RECT  71.97 88.565 71.79 86.86 ;
      RECT  70.245 89.355 70.17 91.06 ;
      RECT  70.17 88.77 69.96 89.15 ;
      RECT  72.33 88.44 72.15 89.355 ;
      POLYGON  70.68 89.445 70.68 89.855 70.505 89.855 70.425 89.775 70.425 89.445 70.68 89.445 ;
      RECT  72.69 89.355 72.51 91.06 ;
      RECT  72.33 89.355 72.15 91.06 ;
      RECT  73.08 89.355 72.87 91.06 ;
      RECT  73.29 89.15 73.08 89.355 ;
      RECT  73.29 89.355 73.08 91.06 ;
      RECT  70.17 89.355 69.96 91.06 ;
      POLYGON  70.68 90.435 70.68 90.845 70.425 90.845 70.425 90.515 70.505 90.435 70.68 90.435 ;
      RECT  73.08 88.77 72.87 89.15 ;
      RECT  70.17 88.44 69.96 88.77 ;
      RECT  71.97 88.44 71.79 89.355 ;
      RECT  70.33 89.94 70.245 90.35 ;
      RECT  71.25 89.355 71.07 91.06 ;
      RECT  70.89 90.435 70.68 90.845 ;
      RECT  73.08 88.44 72.87 88.77 ;
      RECT  70.89 89.445 70.68 89.855 ;
      RECT  70.89 88.77 70.68 89.15 ;
      RECT  73.29 88.77 73.08 89.15 ;
      RECT  71.61 88.44 71.43 89.355 ;
      RECT  71.61 89.355 71.43 91.06 ;
      RECT  70.17 89.15 69.96 89.355 ;
      RECT  73.08 89.15 72.87 89.355 ;
      RECT  73.29 88.44 73.08 88.77 ;
      RECT  71.25 88.44 71.07 89.355 ;
      RECT  72.69 88.44 72.51 89.355 ;
      POLYGON  70.245 88.44 70.245 88.77 70.68 88.77 70.68 89.15 70.245 89.15 70.245 89.355 70.17 89.355 70.17 88.44 70.245 88.44 ;
      RECT  71.97 89.355 71.79 91.06 ;
      RECT  70.245 92.515 70.17 90.81 ;
      RECT  70.17 93.1 69.96 92.72 ;
      RECT  72.33 93.43 72.15 92.515 ;
      POLYGON  70.68 92.425 70.68 92.015 70.505 92.015 70.425 92.095 70.425 92.425 70.68 92.425 ;
      RECT  72.69 92.515 72.51 90.81 ;
      RECT  72.33 92.515 72.15 90.81 ;
      RECT  73.08 92.515 72.87 90.81 ;
      RECT  73.29 92.72 73.08 92.515 ;
      RECT  73.29 92.515 73.08 90.81 ;
      RECT  70.17 92.515 69.96 90.81 ;
      POLYGON  70.68 91.435 70.68 91.025 70.425 91.025 70.425 91.355 70.505 91.435 70.68 91.435 ;
      RECT  73.08 93.1 72.87 92.72 ;
      RECT  70.17 93.43 69.96 93.1 ;
      RECT  71.97 93.43 71.79 92.515 ;
      RECT  70.33 91.93 70.245 91.52 ;
      RECT  71.25 92.515 71.07 90.81 ;
      RECT  70.89 91.435 70.68 91.025 ;
      RECT  73.08 93.43 72.87 93.1 ;
      RECT  70.89 92.425 70.68 92.015 ;
      RECT  70.89 93.1 70.68 92.72 ;
      RECT  73.29 93.1 73.08 92.72 ;
      RECT  71.61 93.43 71.43 92.515 ;
      RECT  71.61 92.515 71.43 90.81 ;
      RECT  70.17 92.72 69.96 92.515 ;
      RECT  73.08 92.72 72.87 92.515 ;
      RECT  73.29 93.43 73.08 93.1 ;
      RECT  71.25 93.43 71.07 92.515 ;
      RECT  72.69 93.43 72.51 92.515 ;
      POLYGON  70.245 93.43 70.245 93.1 70.68 93.1 70.68 92.72 70.245 92.72 70.245 92.515 70.17 92.515 70.17 93.43 70.245 93.43 ;
      RECT  71.97 92.515 71.79 90.81 ;
      RECT  70.245 93.305 70.17 95.01 ;
      RECT  70.17 92.72 69.96 93.1 ;
      RECT  72.33 92.39 72.15 93.305 ;
      POLYGON  70.68 93.395 70.68 93.805 70.505 93.805 70.425 93.725 70.425 93.395 70.68 93.395 ;
      RECT  72.69 93.305 72.51 95.01 ;
      RECT  72.33 93.305 72.15 95.01 ;
      RECT  73.08 93.305 72.87 95.01 ;
      RECT  73.29 93.1 73.08 93.305 ;
      RECT  73.29 93.305 73.08 95.01 ;
      RECT  70.17 93.305 69.96 95.01 ;
      POLYGON  70.68 94.385 70.68 94.795 70.425 94.795 70.425 94.465 70.505 94.385 70.68 94.385 ;
      RECT  73.08 92.72 72.87 93.1 ;
      RECT  70.17 92.39 69.96 92.72 ;
      RECT  71.97 92.39 71.79 93.305 ;
      RECT  70.33 93.89 70.245 94.3 ;
      RECT  71.25 93.305 71.07 95.01 ;
      RECT  70.89 94.385 70.68 94.795 ;
      RECT  73.08 92.39 72.87 92.72 ;
      RECT  70.89 93.395 70.68 93.805 ;
      RECT  70.89 92.72 70.68 93.1 ;
      RECT  73.29 92.72 73.08 93.1 ;
      RECT  71.61 92.39 71.43 93.305 ;
      RECT  71.61 93.305 71.43 95.01 ;
      RECT  70.17 93.1 69.96 93.305 ;
      RECT  73.08 93.1 72.87 93.305 ;
      RECT  73.29 92.39 73.08 92.72 ;
      RECT  71.25 92.39 71.07 93.305 ;
      RECT  72.69 92.39 72.51 93.305 ;
      POLYGON  70.245 92.39 70.245 92.72 70.68 92.72 70.68 93.1 70.245 93.1 70.245 93.305 70.17 93.305 70.17 92.39 70.245 92.39 ;
      RECT  71.97 93.305 71.79 95.01 ;
      RECT  71.97 96.07 71.79 94.49 ;
      RECT  72.33 96.07 72.15 94.49 ;
      RECT  71.88 96.07 71.75 95.36 ;
      RECT  71.61 96.07 71.43 94.49 ;
      RECT  72.01 96.07 71.88 95.36 ;
      RECT  72.33 96.86 72.15 96.07 ;
      RECT  72.69 96.86 72.51 96.07 ;
      RECT  71.25 96.86 71.07 96.07 ;
      RECT  71.97 96.86 71.79 96.07 ;
      RECT  71.61 96.86 71.43 96.07 ;
      RECT  72.69 96.07 72.51 94.49 ;
      RECT  71.25 96.07 71.07 94.49 ;
      RECT  71.79 73.555 71.97 75.26 ;
      RECT  71.79 86.86 71.97 88.565 ;
      RECT  71.79 89.355 71.97 91.06 ;
      RECT  71.79 61.705 71.97 63.41 ;
      RECT  71.79 85.405 71.97 87.11 ;
      RECT  71.79 78.96 71.97 80.665 ;
      RECT  71.79 63.16 71.97 64.865 ;
      RECT  71.79 71.06 71.97 72.765 ;
      RECT  71.79 75.01 71.97 76.715 ;
      RECT  71.79 59.21 71.97 60.915 ;
      RECT  71.79 82.91 71.97 84.615 ;
      RECT  71.79 65.655 71.97 67.36 ;
      RECT  71.79 69.605 71.97 71.31 ;
      RECT  71.79 67.11 71.97 68.815 ;
      RECT  71.79 90.81 71.97 92.515 ;
      RECT  71.79 93.305 71.97 95.01 ;
      RECT  71.79 77.505 71.97 79.21 ;
      RECT  71.79 81.455 71.97 83.16 ;
      RECT  80.43 58.15 80.61 59.73 ;
      RECT  80.07 58.15 80.25 59.73 ;
      RECT  80.52 58.15 80.65 58.86 ;
      RECT  80.79 58.15 80.97 59.73 ;
      RECT  80.39 58.15 80.52 58.86 ;
      RECT  80.07 57.36 80.25 58.15 ;
      RECT  79.71 57.36 79.89 58.15 ;
      RECT  81.15 57.36 81.33 58.15 ;
      RECT  80.43 57.36 80.61 58.15 ;
      RECT  80.79 57.36 80.97 58.15 ;
      RECT  79.71 58.15 79.89 59.73 ;
      RECT  81.15 58.15 81.33 59.73 ;
      RECT  82.155 60.915 82.23 59.21 ;
      RECT  82.23 61.5 82.44 61.12 ;
      RECT  80.07 61.83 80.25 60.915 ;
      POLYGON  81.72 60.825 81.72 60.415 81.895 60.415 81.975 60.495 81.975 60.825 81.72 60.825 ;
      RECT  79.71 60.915 79.89 59.21 ;
      RECT  80.07 60.915 80.25 59.21 ;
      RECT  79.32 60.915 79.53 59.21 ;
      RECT  79.11 61.12 79.32 60.915 ;
      RECT  79.11 60.915 79.32 59.21 ;
      RECT  82.23 60.915 82.44 59.21 ;
      POLYGON  81.72 59.835 81.72 59.425 81.975 59.425 81.975 59.755 81.895 59.835 81.72 59.835 ;
      RECT  79.32 61.5 79.53 61.12 ;
      RECT  82.23 61.83 82.44 61.5 ;
      RECT  80.43 61.83 80.61 60.915 ;
      RECT  82.07 60.33 82.155 59.92 ;
      RECT  81.15 60.915 81.33 59.21 ;
      RECT  81.51 59.835 81.72 59.425 ;
      RECT  79.32 61.83 79.53 61.5 ;
      RECT  81.51 60.825 81.72 60.415 ;
      RECT  81.51 61.5 81.72 61.12 ;
      RECT  79.11 61.5 79.32 61.12 ;
      RECT  80.79 61.83 80.97 60.915 ;
      RECT  80.79 60.915 80.97 59.21 ;
      RECT  82.23 61.12 82.44 60.915 ;
      RECT  79.32 61.12 79.53 60.915 ;
      RECT  79.11 61.83 79.32 61.5 ;
      RECT  81.15 61.83 81.33 60.915 ;
      RECT  79.71 61.83 79.89 60.915 ;
      POLYGON  82.155 61.83 82.155 61.5 81.72 61.5 81.72 61.12 82.155 61.12 82.155 60.915 82.23 60.915 82.23 61.83 82.155 61.83 ;
      RECT  80.43 60.915 80.61 59.21 ;
      RECT  82.155 61.705 82.23 63.41 ;
      RECT  82.23 61.12 82.44 61.5 ;
      RECT  80.07 60.79 80.25 61.705 ;
      POLYGON  81.72 61.795 81.72 62.205 81.895 62.205 81.975 62.125 81.975 61.795 81.72 61.795 ;
      RECT  79.71 61.705 79.89 63.41 ;
      RECT  80.07 61.705 80.25 63.41 ;
      RECT  79.32 61.705 79.53 63.41 ;
      RECT  79.11 61.5 79.32 61.705 ;
      RECT  79.11 61.705 79.32 63.41 ;
      RECT  82.23 61.705 82.44 63.41 ;
      POLYGON  81.72 62.785 81.72 63.195 81.975 63.195 81.975 62.865 81.895 62.785 81.72 62.785 ;
      RECT  79.32 61.12 79.53 61.5 ;
      RECT  82.23 60.79 82.44 61.12 ;
      RECT  80.43 60.79 80.61 61.705 ;
      RECT  82.07 62.29 82.155 62.7 ;
      RECT  81.15 61.705 81.33 63.41 ;
      RECT  81.51 62.785 81.72 63.195 ;
      RECT  79.32 60.79 79.53 61.12 ;
      RECT  81.51 61.795 81.72 62.205 ;
      RECT  81.51 61.12 81.72 61.5 ;
      RECT  79.11 61.12 79.32 61.5 ;
      RECT  80.79 60.79 80.97 61.705 ;
      RECT  80.79 61.705 80.97 63.41 ;
      RECT  82.23 61.5 82.44 61.705 ;
      RECT  79.32 61.5 79.53 61.705 ;
      RECT  79.11 60.79 79.32 61.12 ;
      RECT  81.15 60.79 81.33 61.705 ;
      RECT  79.71 60.79 79.89 61.705 ;
      POLYGON  82.155 60.79 82.155 61.12 81.72 61.12 81.72 61.5 82.155 61.5 82.155 61.705 82.23 61.705 82.23 60.79 82.155 60.79 ;
      RECT  80.43 61.705 80.61 63.41 ;
      RECT  82.155 64.865 82.23 63.16 ;
      RECT  82.23 65.45 82.44 65.07 ;
      RECT  80.07 65.78 80.25 64.865 ;
      POLYGON  81.72 64.775 81.72 64.365 81.895 64.365 81.975 64.445 81.975 64.775 81.72 64.775 ;
      RECT  79.71 64.865 79.89 63.16 ;
      RECT  80.07 64.865 80.25 63.16 ;
      RECT  79.32 64.865 79.53 63.16 ;
      RECT  79.11 65.07 79.32 64.865 ;
      RECT  79.11 64.865 79.32 63.16 ;
      RECT  82.23 64.865 82.44 63.16 ;
      POLYGON  81.72 63.785 81.72 63.375 81.975 63.375 81.975 63.705 81.895 63.785 81.72 63.785 ;
      RECT  79.32 65.45 79.53 65.07 ;
      RECT  82.23 65.78 82.44 65.45 ;
      RECT  80.43 65.78 80.61 64.865 ;
      RECT  82.07 64.28 82.155 63.87 ;
      RECT  81.15 64.865 81.33 63.16 ;
      RECT  81.51 63.785 81.72 63.375 ;
      RECT  79.32 65.78 79.53 65.45 ;
      RECT  81.51 64.775 81.72 64.365 ;
      RECT  81.51 65.45 81.72 65.07 ;
      RECT  79.11 65.45 79.32 65.07 ;
      RECT  80.79 65.78 80.97 64.865 ;
      RECT  80.79 64.865 80.97 63.16 ;
      RECT  82.23 65.07 82.44 64.865 ;
      RECT  79.32 65.07 79.53 64.865 ;
      RECT  79.11 65.78 79.32 65.45 ;
      RECT  81.15 65.78 81.33 64.865 ;
      RECT  79.71 65.78 79.89 64.865 ;
      POLYGON  82.155 65.78 82.155 65.45 81.72 65.45 81.72 65.07 82.155 65.07 82.155 64.865 82.23 64.865 82.23 65.78 82.155 65.78 ;
      RECT  80.43 64.865 80.61 63.16 ;
      RECT  82.155 65.655 82.23 67.36 ;
      RECT  82.23 65.07 82.44 65.45 ;
      RECT  80.07 64.74 80.25 65.655 ;
      POLYGON  81.72 65.745 81.72 66.155 81.895 66.155 81.975 66.075 81.975 65.745 81.72 65.745 ;
      RECT  79.71 65.655 79.89 67.36 ;
      RECT  80.07 65.655 80.25 67.36 ;
      RECT  79.32 65.655 79.53 67.36 ;
      RECT  79.11 65.45 79.32 65.655 ;
      RECT  79.11 65.655 79.32 67.36 ;
      RECT  82.23 65.655 82.44 67.36 ;
      POLYGON  81.72 66.735 81.72 67.145 81.975 67.145 81.975 66.815 81.895 66.735 81.72 66.735 ;
      RECT  79.32 65.07 79.53 65.45 ;
      RECT  82.23 64.74 82.44 65.07 ;
      RECT  80.43 64.74 80.61 65.655 ;
      RECT  82.07 66.24 82.155 66.65 ;
      RECT  81.15 65.655 81.33 67.36 ;
      RECT  81.51 66.735 81.72 67.145 ;
      RECT  79.32 64.74 79.53 65.07 ;
      RECT  81.51 65.745 81.72 66.155 ;
      RECT  81.51 65.07 81.72 65.45 ;
      RECT  79.11 65.07 79.32 65.45 ;
      RECT  80.79 64.74 80.97 65.655 ;
      RECT  80.79 65.655 80.97 67.36 ;
      RECT  82.23 65.45 82.44 65.655 ;
      RECT  79.32 65.45 79.53 65.655 ;
      RECT  79.11 64.74 79.32 65.07 ;
      RECT  81.15 64.74 81.33 65.655 ;
      RECT  79.71 64.74 79.89 65.655 ;
      POLYGON  82.155 64.74 82.155 65.07 81.72 65.07 81.72 65.45 82.155 65.45 82.155 65.655 82.23 65.655 82.23 64.74 82.155 64.74 ;
      RECT  80.43 65.655 80.61 67.36 ;
      RECT  82.155 68.815 82.23 67.11 ;
      RECT  82.23 69.4 82.44 69.02 ;
      RECT  80.07 69.73 80.25 68.815 ;
      POLYGON  81.72 68.725 81.72 68.315 81.895 68.315 81.975 68.395 81.975 68.725 81.72 68.725 ;
      RECT  79.71 68.815 79.89 67.11 ;
      RECT  80.07 68.815 80.25 67.11 ;
      RECT  79.32 68.815 79.53 67.11 ;
      RECT  79.11 69.02 79.32 68.815 ;
      RECT  79.11 68.815 79.32 67.11 ;
      RECT  82.23 68.815 82.44 67.11 ;
      POLYGON  81.72 67.735 81.72 67.325 81.975 67.325 81.975 67.655 81.895 67.735 81.72 67.735 ;
      RECT  79.32 69.4 79.53 69.02 ;
      RECT  82.23 69.73 82.44 69.4 ;
      RECT  80.43 69.73 80.61 68.815 ;
      RECT  82.07 68.23 82.155 67.82 ;
      RECT  81.15 68.815 81.33 67.11 ;
      RECT  81.51 67.735 81.72 67.325 ;
      RECT  79.32 69.73 79.53 69.4 ;
      RECT  81.51 68.725 81.72 68.315 ;
      RECT  81.51 69.4 81.72 69.02 ;
      RECT  79.11 69.4 79.32 69.02 ;
      RECT  80.79 69.73 80.97 68.815 ;
      RECT  80.79 68.815 80.97 67.11 ;
      RECT  82.23 69.02 82.44 68.815 ;
      RECT  79.32 69.02 79.53 68.815 ;
      RECT  79.11 69.73 79.32 69.4 ;
      RECT  81.15 69.73 81.33 68.815 ;
      RECT  79.71 69.73 79.89 68.815 ;
      POLYGON  82.155 69.73 82.155 69.4 81.72 69.4 81.72 69.02 82.155 69.02 82.155 68.815 82.23 68.815 82.23 69.73 82.155 69.73 ;
      RECT  80.43 68.815 80.61 67.11 ;
      RECT  82.155 69.605 82.23 71.31 ;
      RECT  82.23 69.02 82.44 69.4 ;
      RECT  80.07 68.69 80.25 69.605 ;
      POLYGON  81.72 69.695 81.72 70.105 81.895 70.105 81.975 70.025 81.975 69.695 81.72 69.695 ;
      RECT  79.71 69.605 79.89 71.31 ;
      RECT  80.07 69.605 80.25 71.31 ;
      RECT  79.32 69.605 79.53 71.31 ;
      RECT  79.11 69.4 79.32 69.605 ;
      RECT  79.11 69.605 79.32 71.31 ;
      RECT  82.23 69.605 82.44 71.31 ;
      POLYGON  81.72 70.685 81.72 71.095 81.975 71.095 81.975 70.765 81.895 70.685 81.72 70.685 ;
      RECT  79.32 69.02 79.53 69.4 ;
      RECT  82.23 68.69 82.44 69.02 ;
      RECT  80.43 68.69 80.61 69.605 ;
      RECT  82.07 70.19 82.155 70.6 ;
      RECT  81.15 69.605 81.33 71.31 ;
      RECT  81.51 70.685 81.72 71.095 ;
      RECT  79.32 68.69 79.53 69.02 ;
      RECT  81.51 69.695 81.72 70.105 ;
      RECT  81.51 69.02 81.72 69.4 ;
      RECT  79.11 69.02 79.32 69.4 ;
      RECT  80.79 68.69 80.97 69.605 ;
      RECT  80.79 69.605 80.97 71.31 ;
      RECT  82.23 69.4 82.44 69.605 ;
      RECT  79.32 69.4 79.53 69.605 ;
      RECT  79.11 68.69 79.32 69.02 ;
      RECT  81.15 68.69 81.33 69.605 ;
      RECT  79.71 68.69 79.89 69.605 ;
      POLYGON  82.155 68.69 82.155 69.02 81.72 69.02 81.72 69.4 82.155 69.4 82.155 69.605 82.23 69.605 82.23 68.69 82.155 68.69 ;
      RECT  80.43 69.605 80.61 71.31 ;
      RECT  82.155 72.765 82.23 71.06 ;
      RECT  82.23 73.35 82.44 72.97 ;
      RECT  80.07 73.68 80.25 72.765 ;
      POLYGON  81.72 72.675 81.72 72.265 81.895 72.265 81.975 72.345 81.975 72.675 81.72 72.675 ;
      RECT  79.71 72.765 79.89 71.06 ;
      RECT  80.07 72.765 80.25 71.06 ;
      RECT  79.32 72.765 79.53 71.06 ;
      RECT  79.11 72.97 79.32 72.765 ;
      RECT  79.11 72.765 79.32 71.06 ;
      RECT  82.23 72.765 82.44 71.06 ;
      POLYGON  81.72 71.685 81.72 71.275 81.975 71.275 81.975 71.605 81.895 71.685 81.72 71.685 ;
      RECT  79.32 73.35 79.53 72.97 ;
      RECT  82.23 73.68 82.44 73.35 ;
      RECT  80.43 73.68 80.61 72.765 ;
      RECT  82.07 72.18 82.155 71.77 ;
      RECT  81.15 72.765 81.33 71.06 ;
      RECT  81.51 71.685 81.72 71.275 ;
      RECT  79.32 73.68 79.53 73.35 ;
      RECT  81.51 72.675 81.72 72.265 ;
      RECT  81.51 73.35 81.72 72.97 ;
      RECT  79.11 73.35 79.32 72.97 ;
      RECT  80.79 73.68 80.97 72.765 ;
      RECT  80.79 72.765 80.97 71.06 ;
      RECT  82.23 72.97 82.44 72.765 ;
      RECT  79.32 72.97 79.53 72.765 ;
      RECT  79.11 73.68 79.32 73.35 ;
      RECT  81.15 73.68 81.33 72.765 ;
      RECT  79.71 73.68 79.89 72.765 ;
      POLYGON  82.155 73.68 82.155 73.35 81.72 73.35 81.72 72.97 82.155 72.97 82.155 72.765 82.23 72.765 82.23 73.68 82.155 73.68 ;
      RECT  80.43 72.765 80.61 71.06 ;
      RECT  82.155 73.555 82.23 75.26 ;
      RECT  82.23 72.97 82.44 73.35 ;
      RECT  80.07 72.64 80.25 73.555 ;
      POLYGON  81.72 73.645 81.72 74.055 81.895 74.055 81.975 73.975 81.975 73.645 81.72 73.645 ;
      RECT  79.71 73.555 79.89 75.26 ;
      RECT  80.07 73.555 80.25 75.26 ;
      RECT  79.32 73.555 79.53 75.26 ;
      RECT  79.11 73.35 79.32 73.555 ;
      RECT  79.11 73.555 79.32 75.26 ;
      RECT  82.23 73.555 82.44 75.26 ;
      POLYGON  81.72 74.635 81.72 75.045 81.975 75.045 81.975 74.715 81.895 74.635 81.72 74.635 ;
      RECT  79.32 72.97 79.53 73.35 ;
      RECT  82.23 72.64 82.44 72.97 ;
      RECT  80.43 72.64 80.61 73.555 ;
      RECT  82.07 74.14 82.155 74.55 ;
      RECT  81.15 73.555 81.33 75.26 ;
      RECT  81.51 74.635 81.72 75.045 ;
      RECT  79.32 72.64 79.53 72.97 ;
      RECT  81.51 73.645 81.72 74.055 ;
      RECT  81.51 72.97 81.72 73.35 ;
      RECT  79.11 72.97 79.32 73.35 ;
      RECT  80.79 72.64 80.97 73.555 ;
      RECT  80.79 73.555 80.97 75.26 ;
      RECT  82.23 73.35 82.44 73.555 ;
      RECT  79.32 73.35 79.53 73.555 ;
      RECT  79.11 72.64 79.32 72.97 ;
      RECT  81.15 72.64 81.33 73.555 ;
      RECT  79.71 72.64 79.89 73.555 ;
      POLYGON  82.155 72.64 82.155 72.97 81.72 72.97 81.72 73.35 82.155 73.35 82.155 73.555 82.23 73.555 82.23 72.64 82.155 72.64 ;
      RECT  80.43 73.555 80.61 75.26 ;
      RECT  82.155 76.715 82.23 75.01 ;
      RECT  82.23 77.3 82.44 76.92 ;
      RECT  80.07 77.63 80.25 76.715 ;
      POLYGON  81.72 76.625 81.72 76.215 81.895 76.215 81.975 76.295 81.975 76.625 81.72 76.625 ;
      RECT  79.71 76.715 79.89 75.01 ;
      RECT  80.07 76.715 80.25 75.01 ;
      RECT  79.32 76.715 79.53 75.01 ;
      RECT  79.11 76.92 79.32 76.715 ;
      RECT  79.11 76.715 79.32 75.01 ;
      RECT  82.23 76.715 82.44 75.01 ;
      POLYGON  81.72 75.635 81.72 75.225 81.975 75.225 81.975 75.555 81.895 75.635 81.72 75.635 ;
      RECT  79.32 77.3 79.53 76.92 ;
      RECT  82.23 77.63 82.44 77.3 ;
      RECT  80.43 77.63 80.61 76.715 ;
      RECT  82.07 76.13 82.155 75.72 ;
      RECT  81.15 76.715 81.33 75.01 ;
      RECT  81.51 75.635 81.72 75.225 ;
      RECT  79.32 77.63 79.53 77.3 ;
      RECT  81.51 76.625 81.72 76.215 ;
      RECT  81.51 77.3 81.72 76.92 ;
      RECT  79.11 77.3 79.32 76.92 ;
      RECT  80.79 77.63 80.97 76.715 ;
      RECT  80.79 76.715 80.97 75.01 ;
      RECT  82.23 76.92 82.44 76.715 ;
      RECT  79.32 76.92 79.53 76.715 ;
      RECT  79.11 77.63 79.32 77.3 ;
      RECT  81.15 77.63 81.33 76.715 ;
      RECT  79.71 77.63 79.89 76.715 ;
      POLYGON  82.155 77.63 82.155 77.3 81.72 77.3 81.72 76.92 82.155 76.92 82.155 76.715 82.23 76.715 82.23 77.63 82.155 77.63 ;
      RECT  80.43 76.715 80.61 75.01 ;
      RECT  82.155 77.505 82.23 79.21 ;
      RECT  82.23 76.92 82.44 77.3 ;
      RECT  80.07 76.59 80.25 77.505 ;
      POLYGON  81.72 77.595 81.72 78.005 81.895 78.005 81.975 77.925 81.975 77.595 81.72 77.595 ;
      RECT  79.71 77.505 79.89 79.21 ;
      RECT  80.07 77.505 80.25 79.21 ;
      RECT  79.32 77.505 79.53 79.21 ;
      RECT  79.11 77.3 79.32 77.505 ;
      RECT  79.11 77.505 79.32 79.21 ;
      RECT  82.23 77.505 82.44 79.21 ;
      POLYGON  81.72 78.585 81.72 78.995 81.975 78.995 81.975 78.665 81.895 78.585 81.72 78.585 ;
      RECT  79.32 76.92 79.53 77.3 ;
      RECT  82.23 76.59 82.44 76.92 ;
      RECT  80.43 76.59 80.61 77.505 ;
      RECT  82.07 78.09 82.155 78.5 ;
      RECT  81.15 77.505 81.33 79.21 ;
      RECT  81.51 78.585 81.72 78.995 ;
      RECT  79.32 76.59 79.53 76.92 ;
      RECT  81.51 77.595 81.72 78.005 ;
      RECT  81.51 76.92 81.72 77.3 ;
      RECT  79.11 76.92 79.32 77.3 ;
      RECT  80.79 76.59 80.97 77.505 ;
      RECT  80.79 77.505 80.97 79.21 ;
      RECT  82.23 77.3 82.44 77.505 ;
      RECT  79.32 77.3 79.53 77.505 ;
      RECT  79.11 76.59 79.32 76.92 ;
      RECT  81.15 76.59 81.33 77.505 ;
      RECT  79.71 76.59 79.89 77.505 ;
      POLYGON  82.155 76.59 82.155 76.92 81.72 76.92 81.72 77.3 82.155 77.3 82.155 77.505 82.23 77.505 82.23 76.59 82.155 76.59 ;
      RECT  80.43 77.505 80.61 79.21 ;
      RECT  82.155 80.665 82.23 78.96 ;
      RECT  82.23 81.25 82.44 80.87 ;
      RECT  80.07 81.58 80.25 80.665 ;
      POLYGON  81.72 80.575 81.72 80.165 81.895 80.165 81.975 80.245 81.975 80.575 81.72 80.575 ;
      RECT  79.71 80.665 79.89 78.96 ;
      RECT  80.07 80.665 80.25 78.96 ;
      RECT  79.32 80.665 79.53 78.96 ;
      RECT  79.11 80.87 79.32 80.665 ;
      RECT  79.11 80.665 79.32 78.96 ;
      RECT  82.23 80.665 82.44 78.96 ;
      POLYGON  81.72 79.585 81.72 79.175 81.975 79.175 81.975 79.505 81.895 79.585 81.72 79.585 ;
      RECT  79.32 81.25 79.53 80.87 ;
      RECT  82.23 81.58 82.44 81.25 ;
      RECT  80.43 81.58 80.61 80.665 ;
      RECT  82.07 80.08 82.155 79.67 ;
      RECT  81.15 80.665 81.33 78.96 ;
      RECT  81.51 79.585 81.72 79.175 ;
      RECT  79.32 81.58 79.53 81.25 ;
      RECT  81.51 80.575 81.72 80.165 ;
      RECT  81.51 81.25 81.72 80.87 ;
      RECT  79.11 81.25 79.32 80.87 ;
      RECT  80.79 81.58 80.97 80.665 ;
      RECT  80.79 80.665 80.97 78.96 ;
      RECT  82.23 80.87 82.44 80.665 ;
      RECT  79.32 80.87 79.53 80.665 ;
      RECT  79.11 81.58 79.32 81.25 ;
      RECT  81.15 81.58 81.33 80.665 ;
      RECT  79.71 81.58 79.89 80.665 ;
      POLYGON  82.155 81.58 82.155 81.25 81.72 81.25 81.72 80.87 82.155 80.87 82.155 80.665 82.23 80.665 82.23 81.58 82.155 81.58 ;
      RECT  80.43 80.665 80.61 78.96 ;
      RECT  82.155 81.455 82.23 83.16 ;
      RECT  82.23 80.87 82.44 81.25 ;
      RECT  80.07 80.54 80.25 81.455 ;
      POLYGON  81.72 81.545 81.72 81.955 81.895 81.955 81.975 81.875 81.975 81.545 81.72 81.545 ;
      RECT  79.71 81.455 79.89 83.16 ;
      RECT  80.07 81.455 80.25 83.16 ;
      RECT  79.32 81.455 79.53 83.16 ;
      RECT  79.11 81.25 79.32 81.455 ;
      RECT  79.11 81.455 79.32 83.16 ;
      RECT  82.23 81.455 82.44 83.16 ;
      POLYGON  81.72 82.535 81.72 82.945 81.975 82.945 81.975 82.615 81.895 82.535 81.72 82.535 ;
      RECT  79.32 80.87 79.53 81.25 ;
      RECT  82.23 80.54 82.44 80.87 ;
      RECT  80.43 80.54 80.61 81.455 ;
      RECT  82.07 82.04 82.155 82.45 ;
      RECT  81.15 81.455 81.33 83.16 ;
      RECT  81.51 82.535 81.72 82.945 ;
      RECT  79.32 80.54 79.53 80.87 ;
      RECT  81.51 81.545 81.72 81.955 ;
      RECT  81.51 80.87 81.72 81.25 ;
      RECT  79.11 80.87 79.32 81.25 ;
      RECT  80.79 80.54 80.97 81.455 ;
      RECT  80.79 81.455 80.97 83.16 ;
      RECT  82.23 81.25 82.44 81.455 ;
      RECT  79.32 81.25 79.53 81.455 ;
      RECT  79.11 80.54 79.32 80.87 ;
      RECT  81.15 80.54 81.33 81.455 ;
      RECT  79.71 80.54 79.89 81.455 ;
      POLYGON  82.155 80.54 82.155 80.87 81.72 80.87 81.72 81.25 82.155 81.25 82.155 81.455 82.23 81.455 82.23 80.54 82.155 80.54 ;
      RECT  80.43 81.455 80.61 83.16 ;
      RECT  82.155 84.615 82.23 82.91 ;
      RECT  82.23 85.2 82.44 84.82 ;
      RECT  80.07 85.53 80.25 84.615 ;
      POLYGON  81.72 84.525 81.72 84.115 81.895 84.115 81.975 84.195 81.975 84.525 81.72 84.525 ;
      RECT  79.71 84.615 79.89 82.91 ;
      RECT  80.07 84.615 80.25 82.91 ;
      RECT  79.32 84.615 79.53 82.91 ;
      RECT  79.11 84.82 79.32 84.615 ;
      RECT  79.11 84.615 79.32 82.91 ;
      RECT  82.23 84.615 82.44 82.91 ;
      POLYGON  81.72 83.535 81.72 83.125 81.975 83.125 81.975 83.455 81.895 83.535 81.72 83.535 ;
      RECT  79.32 85.2 79.53 84.82 ;
      RECT  82.23 85.53 82.44 85.2 ;
      RECT  80.43 85.53 80.61 84.615 ;
      RECT  82.07 84.03 82.155 83.62 ;
      RECT  81.15 84.615 81.33 82.91 ;
      RECT  81.51 83.535 81.72 83.125 ;
      RECT  79.32 85.53 79.53 85.2 ;
      RECT  81.51 84.525 81.72 84.115 ;
      RECT  81.51 85.2 81.72 84.82 ;
      RECT  79.11 85.2 79.32 84.82 ;
      RECT  80.79 85.53 80.97 84.615 ;
      RECT  80.79 84.615 80.97 82.91 ;
      RECT  82.23 84.82 82.44 84.615 ;
      RECT  79.32 84.82 79.53 84.615 ;
      RECT  79.11 85.53 79.32 85.2 ;
      RECT  81.15 85.53 81.33 84.615 ;
      RECT  79.71 85.53 79.89 84.615 ;
      POLYGON  82.155 85.53 82.155 85.2 81.72 85.2 81.72 84.82 82.155 84.82 82.155 84.615 82.23 84.615 82.23 85.53 82.155 85.53 ;
      RECT  80.43 84.615 80.61 82.91 ;
      RECT  82.155 85.405 82.23 87.11 ;
      RECT  82.23 84.82 82.44 85.2 ;
      RECT  80.07 84.49 80.25 85.405 ;
      POLYGON  81.72 85.495 81.72 85.905 81.895 85.905 81.975 85.825 81.975 85.495 81.72 85.495 ;
      RECT  79.71 85.405 79.89 87.11 ;
      RECT  80.07 85.405 80.25 87.11 ;
      RECT  79.32 85.405 79.53 87.11 ;
      RECT  79.11 85.2 79.32 85.405 ;
      RECT  79.11 85.405 79.32 87.11 ;
      RECT  82.23 85.405 82.44 87.11 ;
      POLYGON  81.72 86.485 81.72 86.895 81.975 86.895 81.975 86.565 81.895 86.485 81.72 86.485 ;
      RECT  79.32 84.82 79.53 85.2 ;
      RECT  82.23 84.49 82.44 84.82 ;
      RECT  80.43 84.49 80.61 85.405 ;
      RECT  82.07 85.99 82.155 86.4 ;
      RECT  81.15 85.405 81.33 87.11 ;
      RECT  81.51 86.485 81.72 86.895 ;
      RECT  79.32 84.49 79.53 84.82 ;
      RECT  81.51 85.495 81.72 85.905 ;
      RECT  81.51 84.82 81.72 85.2 ;
      RECT  79.11 84.82 79.32 85.2 ;
      RECT  80.79 84.49 80.97 85.405 ;
      RECT  80.79 85.405 80.97 87.11 ;
      RECT  82.23 85.2 82.44 85.405 ;
      RECT  79.32 85.2 79.53 85.405 ;
      RECT  79.11 84.49 79.32 84.82 ;
      RECT  81.15 84.49 81.33 85.405 ;
      RECT  79.71 84.49 79.89 85.405 ;
      POLYGON  82.155 84.49 82.155 84.82 81.72 84.82 81.72 85.2 82.155 85.2 82.155 85.405 82.23 85.405 82.23 84.49 82.155 84.49 ;
      RECT  80.43 85.405 80.61 87.11 ;
      RECT  82.155 88.565 82.23 86.86 ;
      RECT  82.23 89.15 82.44 88.77 ;
      RECT  80.07 89.48 80.25 88.565 ;
      POLYGON  81.72 88.475 81.72 88.065 81.895 88.065 81.975 88.145 81.975 88.475 81.72 88.475 ;
      RECT  79.71 88.565 79.89 86.86 ;
      RECT  80.07 88.565 80.25 86.86 ;
      RECT  79.32 88.565 79.53 86.86 ;
      RECT  79.11 88.77 79.32 88.565 ;
      RECT  79.11 88.565 79.32 86.86 ;
      RECT  82.23 88.565 82.44 86.86 ;
      POLYGON  81.72 87.485 81.72 87.075 81.975 87.075 81.975 87.405 81.895 87.485 81.72 87.485 ;
      RECT  79.32 89.15 79.53 88.77 ;
      RECT  82.23 89.48 82.44 89.15 ;
      RECT  80.43 89.48 80.61 88.565 ;
      RECT  82.07 87.98 82.155 87.57 ;
      RECT  81.15 88.565 81.33 86.86 ;
      RECT  81.51 87.485 81.72 87.075 ;
      RECT  79.32 89.48 79.53 89.15 ;
      RECT  81.51 88.475 81.72 88.065 ;
      RECT  81.51 89.15 81.72 88.77 ;
      RECT  79.11 89.15 79.32 88.77 ;
      RECT  80.79 89.48 80.97 88.565 ;
      RECT  80.79 88.565 80.97 86.86 ;
      RECT  82.23 88.77 82.44 88.565 ;
      RECT  79.32 88.77 79.53 88.565 ;
      RECT  79.11 89.48 79.32 89.15 ;
      RECT  81.15 89.48 81.33 88.565 ;
      RECT  79.71 89.48 79.89 88.565 ;
      POLYGON  82.155 89.48 82.155 89.15 81.72 89.15 81.72 88.77 82.155 88.77 82.155 88.565 82.23 88.565 82.23 89.48 82.155 89.48 ;
      RECT  80.43 88.565 80.61 86.86 ;
      RECT  82.155 89.355 82.23 91.06 ;
      RECT  82.23 88.77 82.44 89.15 ;
      RECT  80.07 88.44 80.25 89.355 ;
      POLYGON  81.72 89.445 81.72 89.855 81.895 89.855 81.975 89.775 81.975 89.445 81.72 89.445 ;
      RECT  79.71 89.355 79.89 91.06 ;
      RECT  80.07 89.355 80.25 91.06 ;
      RECT  79.32 89.355 79.53 91.06 ;
      RECT  79.11 89.15 79.32 89.355 ;
      RECT  79.11 89.355 79.32 91.06 ;
      RECT  82.23 89.355 82.44 91.06 ;
      POLYGON  81.72 90.435 81.72 90.845 81.975 90.845 81.975 90.515 81.895 90.435 81.72 90.435 ;
      RECT  79.32 88.77 79.53 89.15 ;
      RECT  82.23 88.44 82.44 88.77 ;
      RECT  80.43 88.44 80.61 89.355 ;
      RECT  82.07 89.94 82.155 90.35 ;
      RECT  81.15 89.355 81.33 91.06 ;
      RECT  81.51 90.435 81.72 90.845 ;
      RECT  79.32 88.44 79.53 88.77 ;
      RECT  81.51 89.445 81.72 89.855 ;
      RECT  81.51 88.77 81.72 89.15 ;
      RECT  79.11 88.77 79.32 89.15 ;
      RECT  80.79 88.44 80.97 89.355 ;
      RECT  80.79 89.355 80.97 91.06 ;
      RECT  82.23 89.15 82.44 89.355 ;
      RECT  79.32 89.15 79.53 89.355 ;
      RECT  79.11 88.44 79.32 88.77 ;
      RECT  81.15 88.44 81.33 89.355 ;
      RECT  79.71 88.44 79.89 89.355 ;
      POLYGON  82.155 88.44 82.155 88.77 81.72 88.77 81.72 89.15 82.155 89.15 82.155 89.355 82.23 89.355 82.23 88.44 82.155 88.44 ;
      RECT  80.43 89.355 80.61 91.06 ;
      RECT  82.155 92.515 82.23 90.81 ;
      RECT  82.23 93.1 82.44 92.72 ;
      RECT  80.07 93.43 80.25 92.515 ;
      POLYGON  81.72 92.425 81.72 92.015 81.895 92.015 81.975 92.095 81.975 92.425 81.72 92.425 ;
      RECT  79.71 92.515 79.89 90.81 ;
      RECT  80.07 92.515 80.25 90.81 ;
      RECT  79.32 92.515 79.53 90.81 ;
      RECT  79.11 92.72 79.32 92.515 ;
      RECT  79.11 92.515 79.32 90.81 ;
      RECT  82.23 92.515 82.44 90.81 ;
      POLYGON  81.72 91.435 81.72 91.025 81.975 91.025 81.975 91.355 81.895 91.435 81.72 91.435 ;
      RECT  79.32 93.1 79.53 92.72 ;
      RECT  82.23 93.43 82.44 93.1 ;
      RECT  80.43 93.43 80.61 92.515 ;
      RECT  82.07 91.93 82.155 91.52 ;
      RECT  81.15 92.515 81.33 90.81 ;
      RECT  81.51 91.435 81.72 91.025 ;
      RECT  79.32 93.43 79.53 93.1 ;
      RECT  81.51 92.425 81.72 92.015 ;
      RECT  81.51 93.1 81.72 92.72 ;
      RECT  79.11 93.1 79.32 92.72 ;
      RECT  80.79 93.43 80.97 92.515 ;
      RECT  80.79 92.515 80.97 90.81 ;
      RECT  82.23 92.72 82.44 92.515 ;
      RECT  79.32 92.72 79.53 92.515 ;
      RECT  79.11 93.43 79.32 93.1 ;
      RECT  81.15 93.43 81.33 92.515 ;
      RECT  79.71 93.43 79.89 92.515 ;
      POLYGON  82.155 93.43 82.155 93.1 81.72 93.1 81.72 92.72 82.155 92.72 82.155 92.515 82.23 92.515 82.23 93.43 82.155 93.43 ;
      RECT  80.43 92.515 80.61 90.81 ;
      RECT  82.155 93.305 82.23 95.01 ;
      RECT  82.23 92.72 82.44 93.1 ;
      RECT  80.07 92.39 80.25 93.305 ;
      POLYGON  81.72 93.395 81.72 93.805 81.895 93.805 81.975 93.725 81.975 93.395 81.72 93.395 ;
      RECT  79.71 93.305 79.89 95.01 ;
      RECT  80.07 93.305 80.25 95.01 ;
      RECT  79.32 93.305 79.53 95.01 ;
      RECT  79.11 93.1 79.32 93.305 ;
      RECT  79.11 93.305 79.32 95.01 ;
      RECT  82.23 93.305 82.44 95.01 ;
      POLYGON  81.72 94.385 81.72 94.795 81.975 94.795 81.975 94.465 81.895 94.385 81.72 94.385 ;
      RECT  79.32 92.72 79.53 93.1 ;
      RECT  82.23 92.39 82.44 92.72 ;
      RECT  80.43 92.39 80.61 93.305 ;
      RECT  82.07 93.89 82.155 94.3 ;
      RECT  81.15 93.305 81.33 95.01 ;
      RECT  81.51 94.385 81.72 94.795 ;
      RECT  79.32 92.39 79.53 92.72 ;
      RECT  81.51 93.395 81.72 93.805 ;
      RECT  81.51 92.72 81.72 93.1 ;
      RECT  79.11 92.72 79.32 93.1 ;
      RECT  80.79 92.39 80.97 93.305 ;
      RECT  80.79 93.305 80.97 95.01 ;
      RECT  82.23 93.1 82.44 93.305 ;
      RECT  79.32 93.1 79.53 93.305 ;
      RECT  79.11 92.39 79.32 92.72 ;
      RECT  81.15 92.39 81.33 93.305 ;
      RECT  79.71 92.39 79.89 93.305 ;
      POLYGON  82.155 92.39 82.155 92.72 81.72 92.72 81.72 93.1 82.155 93.1 82.155 93.305 82.23 93.305 82.23 92.39 82.155 92.39 ;
      RECT  80.43 93.305 80.61 95.01 ;
      RECT  80.43 96.07 80.61 94.49 ;
      RECT  80.07 96.07 80.25 94.49 ;
      RECT  80.52 96.07 80.65 95.36 ;
      RECT  80.79 96.07 80.97 94.49 ;
      RECT  80.39 96.07 80.52 95.36 ;
      RECT  80.07 96.86 80.25 96.07 ;
      RECT  79.71 96.86 79.89 96.07 ;
      RECT  81.15 96.86 81.33 96.07 ;
      RECT  80.43 96.86 80.61 96.07 ;
      RECT  80.79 96.86 80.97 96.07 ;
      RECT  79.71 96.07 79.89 94.49 ;
      RECT  81.15 96.07 81.33 94.49 ;
      RECT  80.43 82.91 80.61 84.615 ;
      RECT  80.43 86.86 80.61 88.565 ;
      RECT  80.43 65.655 80.61 67.36 ;
      RECT  80.43 59.21 80.61 60.915 ;
      RECT  80.43 81.455 80.61 83.16 ;
      RECT  80.43 71.06 80.61 72.765 ;
      RECT  80.43 78.96 80.61 80.665 ;
      RECT  80.43 89.355 80.61 91.06 ;
      RECT  80.43 63.16 80.61 64.865 ;
      RECT  80.43 93.305 80.61 95.01 ;
      RECT  80.43 90.81 80.61 92.515 ;
      RECT  80.43 67.11 80.61 68.815 ;
      RECT  80.43 73.555 80.61 75.26 ;
      RECT  80.43 61.705 80.61 63.41 ;
      RECT  80.43 85.405 80.61 87.11 ;
      RECT  80.43 69.605 80.61 71.31 ;
      RECT  80.43 75.01 80.61 76.715 ;
      RECT  80.43 77.505 80.61 79.21 ;
      RECT  75.915 60.915 75.99 59.21 ;
      RECT  75.99 61.5 76.2 61.12 ;
      RECT  73.83 61.83 74.01 60.915 ;
      POLYGON  75.48 60.825 75.48 60.415 75.655 60.415 75.735 60.495 75.735 60.825 75.48 60.825 ;
      RECT  73.47 60.915 73.65 59.21 ;
      RECT  73.83 60.915 74.01 59.21 ;
      RECT  73.08 60.915 73.29 59.21 ;
      RECT  72.87 61.12 73.08 60.915 ;
      RECT  72.87 60.915 73.08 59.21 ;
      RECT  75.99 60.915 76.2 59.21 ;
      POLYGON  75.48 59.835 75.48 59.425 75.735 59.425 75.735 59.755 75.655 59.835 75.48 59.835 ;
      RECT  73.08 61.5 73.29 61.12 ;
      RECT  75.99 61.83 76.2 61.5 ;
      RECT  74.19 61.83 74.37 60.915 ;
      RECT  75.83 60.33 75.915 59.92 ;
      RECT  74.91 60.915 75.09 59.21 ;
      RECT  75.27 59.835 75.48 59.425 ;
      RECT  73.08 61.83 73.29 61.5 ;
      RECT  75.27 60.825 75.48 60.415 ;
      RECT  75.27 61.5 75.48 61.12 ;
      RECT  72.87 61.5 73.08 61.12 ;
      RECT  74.55 61.83 74.73 60.915 ;
      RECT  74.55 60.915 74.73 59.21 ;
      RECT  75.99 61.12 76.2 60.915 ;
      RECT  73.08 61.12 73.29 60.915 ;
      RECT  72.87 61.83 73.08 61.5 ;
      RECT  74.91 61.83 75.09 60.915 ;
      RECT  73.47 61.83 73.65 60.915 ;
      POLYGON  75.915 61.83 75.915 61.5 75.48 61.5 75.48 61.12 75.915 61.12 75.915 60.915 75.99 60.915 75.99 61.83 75.915 61.83 ;
      RECT  74.19 60.915 74.37 59.21 ;
      RECT  76.485 60.915 76.41 59.21 ;
      RECT  76.41 61.5 76.2 61.12 ;
      RECT  78.57 61.83 78.39 60.915 ;
      POLYGON  76.92 60.825 76.92 60.415 76.745 60.415 76.665 60.495 76.665 60.825 76.92 60.825 ;
      RECT  78.93 60.915 78.75 59.21 ;
      RECT  78.57 60.915 78.39 59.21 ;
      RECT  79.32 60.915 79.11 59.21 ;
      RECT  79.53 61.12 79.32 60.915 ;
      RECT  79.53 60.915 79.32 59.21 ;
      RECT  76.41 60.915 76.2 59.21 ;
      POLYGON  76.92 59.835 76.92 59.425 76.665 59.425 76.665 59.755 76.745 59.835 76.92 59.835 ;
      RECT  79.32 61.5 79.11 61.12 ;
      RECT  76.41 61.83 76.2 61.5 ;
      RECT  78.21 61.83 78.03 60.915 ;
      RECT  76.57 60.33 76.485 59.92 ;
      RECT  77.49 60.915 77.31 59.21 ;
      RECT  77.13 59.835 76.92 59.425 ;
      RECT  79.32 61.83 79.11 61.5 ;
      RECT  77.13 60.825 76.92 60.415 ;
      RECT  77.13 61.5 76.92 61.12 ;
      RECT  79.53 61.5 79.32 61.12 ;
      RECT  77.85 61.83 77.67 60.915 ;
      RECT  77.85 60.915 77.67 59.21 ;
      RECT  76.41 61.12 76.2 60.915 ;
      RECT  79.32 61.12 79.11 60.915 ;
      RECT  79.53 61.83 79.32 61.5 ;
      RECT  77.49 61.83 77.31 60.915 ;
      RECT  78.93 61.83 78.75 60.915 ;
      POLYGON  76.485 61.83 76.485 61.5 76.92 61.5 76.92 61.12 76.485 61.12 76.485 60.915 76.41 60.915 76.41 61.83 76.485 61.83 ;
      RECT  78.21 60.915 78.03 59.21 ;
      RECT  73.47 61.31 73.65 59.335 ;
      RECT  73.83 61.31 74.01 59.335 ;
      RECT  74.55 61.31 74.73 59.335 ;
      RECT  74.91 61.31 75.09 59.335 ;
      RECT  78.75 61.31 78.93 59.335 ;
      RECT  78.39 61.31 78.57 59.335 ;
      RECT  77.67 61.31 77.85 59.335 ;
      RECT  77.31 61.31 77.49 59.335 ;
      RECT  74.19 60.915 74.37 59.21 ;
      RECT  78.03 60.915 78.21 59.21 ;
      RECT  75.915 93.305 75.99 95.01 ;
      RECT  75.99 92.72 76.2 93.1 ;
      RECT  73.83 92.39 74.01 93.305 ;
      POLYGON  75.48 93.395 75.48 93.805 75.655 93.805 75.735 93.725 75.735 93.395 75.48 93.395 ;
      RECT  73.47 93.305 73.65 95.01 ;
      RECT  73.83 93.305 74.01 95.01 ;
      RECT  73.08 93.305 73.29 95.01 ;
      RECT  72.87 93.1 73.08 93.305 ;
      RECT  72.87 93.305 73.08 95.01 ;
      RECT  75.99 93.305 76.2 95.01 ;
      POLYGON  75.48 94.385 75.48 94.795 75.735 94.795 75.735 94.465 75.655 94.385 75.48 94.385 ;
      RECT  73.08 92.72 73.29 93.1 ;
      RECT  75.99 92.39 76.2 92.72 ;
      RECT  74.19 92.39 74.37 93.305 ;
      RECT  75.83 93.89 75.915 94.3 ;
      RECT  74.91 93.305 75.09 95.01 ;
      RECT  75.27 94.385 75.48 94.795 ;
      RECT  73.08 92.39 73.29 92.72 ;
      RECT  75.27 93.395 75.48 93.805 ;
      RECT  75.27 92.72 75.48 93.1 ;
      RECT  72.87 92.72 73.08 93.1 ;
      RECT  74.55 92.39 74.73 93.305 ;
      RECT  74.55 93.305 74.73 95.01 ;
      RECT  75.99 93.1 76.2 93.305 ;
      RECT  73.08 93.1 73.29 93.305 ;
      RECT  72.87 92.39 73.08 92.72 ;
      RECT  74.91 92.39 75.09 93.305 ;
      RECT  73.47 92.39 73.65 93.305 ;
      POLYGON  75.915 92.39 75.915 92.72 75.48 92.72 75.48 93.1 75.915 93.1 75.915 93.305 75.99 93.305 75.99 92.39 75.915 92.39 ;
      RECT  74.19 93.305 74.37 95.01 ;
      RECT  76.485 93.305 76.41 95.01 ;
      RECT  76.41 92.72 76.2 93.1 ;
      RECT  78.57 92.39 78.39 93.305 ;
      POLYGON  76.92 93.395 76.92 93.805 76.745 93.805 76.665 93.725 76.665 93.395 76.92 93.395 ;
      RECT  78.93 93.305 78.75 95.01 ;
      RECT  78.57 93.305 78.39 95.01 ;
      RECT  79.32 93.305 79.11 95.01 ;
      RECT  79.53 93.1 79.32 93.305 ;
      RECT  79.53 93.305 79.32 95.01 ;
      RECT  76.41 93.305 76.2 95.01 ;
      POLYGON  76.92 94.385 76.92 94.795 76.665 94.795 76.665 94.465 76.745 94.385 76.92 94.385 ;
      RECT  79.32 92.72 79.11 93.1 ;
      RECT  76.41 92.39 76.2 92.72 ;
      RECT  78.21 92.39 78.03 93.305 ;
      RECT  76.57 93.89 76.485 94.3 ;
      RECT  77.49 93.305 77.31 95.01 ;
      RECT  77.13 94.385 76.92 94.795 ;
      RECT  79.32 92.39 79.11 92.72 ;
      RECT  77.13 93.395 76.92 93.805 ;
      RECT  77.13 92.72 76.92 93.1 ;
      RECT  79.53 92.72 79.32 93.1 ;
      RECT  77.85 92.39 77.67 93.305 ;
      RECT  77.85 93.305 77.67 95.01 ;
      RECT  76.41 93.1 76.2 93.305 ;
      RECT  79.32 93.1 79.11 93.305 ;
      RECT  79.53 92.39 79.32 92.72 ;
      RECT  77.49 92.39 77.31 93.305 ;
      RECT  78.93 92.39 78.75 93.305 ;
      POLYGON  76.485 92.39 76.485 92.72 76.92 92.72 76.92 93.1 76.485 93.1 76.485 93.305 76.41 93.305 76.41 92.39 76.485 92.39 ;
      RECT  78.21 93.305 78.03 95.01 ;
      RECT  73.47 92.91 73.65 94.885 ;
      RECT  73.83 92.91 74.01 94.885 ;
      RECT  74.55 92.91 74.73 94.885 ;
      RECT  74.91 92.91 75.09 94.885 ;
      RECT  78.75 92.91 78.93 94.885 ;
      RECT  78.39 92.91 78.57 94.885 ;
      RECT  77.67 92.91 77.85 94.885 ;
      RECT  77.31 92.91 77.49 94.885 ;
      RECT  74.19 93.305 74.37 95.01 ;
      RECT  78.03 93.305 78.21 95.01 ;
      RECT  74.19 58.15 74.37 59.73 ;
      RECT  73.83 58.15 74.01 59.73 ;
      RECT  74.28 58.15 74.41 58.86 ;
      RECT  74.55 58.15 74.73 59.73 ;
      RECT  74.15 58.15 74.28 58.86 ;
      RECT  73.83 57.36 74.01 58.15 ;
      RECT  73.47 57.36 73.65 58.15 ;
      RECT  74.91 57.36 75.09 58.15 ;
      RECT  74.19 57.36 74.37 58.15 ;
      RECT  74.55 57.36 74.73 58.15 ;
      RECT  73.47 58.15 73.65 59.73 ;
      RECT  74.91 58.15 75.09 59.73 ;
      RECT  78.21 58.15 78.03 59.73 ;
      RECT  78.57 58.15 78.39 59.73 ;
      RECT  78.12 58.15 77.99 58.86 ;
      RECT  77.85 58.15 77.67 59.73 ;
      RECT  78.25 58.15 78.12 58.86 ;
      RECT  78.57 57.36 78.39 58.15 ;
      RECT  78.93 57.36 78.75 58.15 ;
      RECT  77.49 57.36 77.31 58.15 ;
      RECT  78.21 57.36 78.03 58.15 ;
      RECT  77.85 57.36 77.67 58.15 ;
      RECT  78.93 58.15 78.75 59.73 ;
      RECT  77.49 58.15 77.31 59.73 ;
      RECT  73.47 57.36 73.65 59.335 ;
      RECT  73.83 57.36 74.01 59.335 ;
      RECT  74.55 57.36 74.73 59.335 ;
      RECT  74.91 57.36 75.09 59.335 ;
      RECT  78.75 57.36 78.93 59.335 ;
      RECT  78.39 57.36 78.57 59.335 ;
      RECT  77.67 57.36 77.85 59.335 ;
      RECT  77.31 57.36 77.49 59.335 ;
      RECT  74.19 96.07 74.37 94.49 ;
      RECT  73.83 96.07 74.01 94.49 ;
      RECT  74.28 96.07 74.41 95.36 ;
      RECT  74.55 96.07 74.73 94.49 ;
      RECT  74.15 96.07 74.28 95.36 ;
      RECT  73.83 96.86 74.01 96.07 ;
      RECT  73.47 96.86 73.65 96.07 ;
      RECT  74.91 96.86 75.09 96.07 ;
      RECT  74.19 96.86 74.37 96.07 ;
      RECT  74.55 96.86 74.73 96.07 ;
      RECT  73.47 96.07 73.65 94.49 ;
      RECT  74.91 96.07 75.09 94.49 ;
      RECT  78.21 96.07 78.03 94.49 ;
      RECT  78.57 96.07 78.39 94.49 ;
      RECT  78.12 96.07 77.99 95.36 ;
      RECT  77.85 96.07 77.67 94.49 ;
      RECT  78.25 96.07 78.12 95.36 ;
      RECT  78.57 96.86 78.39 96.07 ;
      RECT  78.93 96.86 78.75 96.07 ;
      RECT  77.49 96.86 77.31 96.07 ;
      RECT  78.21 96.86 78.03 96.07 ;
      RECT  77.85 96.86 77.67 96.07 ;
      RECT  78.93 96.07 78.75 94.49 ;
      RECT  77.49 96.07 77.31 94.49 ;
      RECT  73.47 96.86 73.65 94.885 ;
      RECT  73.83 96.86 74.01 94.885 ;
      RECT  74.55 96.86 74.73 94.885 ;
      RECT  74.91 96.86 75.09 94.885 ;
      RECT  78.75 96.86 78.93 94.885 ;
      RECT  78.39 96.86 78.57 94.885 ;
      RECT  77.67 96.86 77.85 94.885 ;
      RECT  77.31 96.86 77.49 94.885 ;
      RECT  73.47 57.36 73.65 96.86 ;
      RECT  73.83 57.36 74.01 96.86 ;
      RECT  74.55 57.36 74.73 96.86 ;
      RECT  74.91 57.36 75.09 96.86 ;
      RECT  78.75 57.36 78.93 96.86 ;
      RECT  78.39 57.36 78.57 96.86 ;
      RECT  77.67 57.36 77.85 96.86 ;
      RECT  77.31 57.36 77.49 96.86 ;
      RECT  72.51 57.36 72.69 96.86 ;
      RECT  72.15 57.36 72.33 96.86 ;
      RECT  80.79 57.36 80.97 96.86 ;
      RECT  81.15 57.36 81.33 96.86 ;
      RECT  80.43 73.555 80.61 75.26 ;
      RECT  80.43 86.86 80.61 88.565 ;
      RECT  80.43 71.06 80.61 72.765 ;
      RECT  71.79 89.355 71.97 91.06 ;
      RECT  71.79 78.96 71.97 80.665 ;
      RECT  80.43 85.405 80.61 87.11 ;
      RECT  80.43 82.91 80.61 84.615 ;
      RECT  71.79 71.06 71.97 72.765 ;
      RECT  71.79 69.605 71.97 71.31 ;
      RECT  80.43 69.605 80.61 71.31 ;
      RECT  71.79 85.405 71.97 87.11 ;
      RECT  80.43 65.655 80.61 67.36 ;
      RECT  80.43 89.355 80.61 91.06 ;
      RECT  71.79 82.91 71.97 84.615 ;
      RECT  71.79 86.86 71.97 88.565 ;
      RECT  71.79 59.21 71.97 60.915 ;
      RECT  71.79 77.505 71.97 79.21 ;
      RECT  71.79 61.705 71.97 63.41 ;
      RECT  80.43 81.455 80.61 83.16 ;
      RECT  80.43 61.705 80.61 63.41 ;
      RECT  71.79 63.16 71.97 64.865 ;
      RECT  71.79 90.81 71.97 92.515 ;
      RECT  80.43 59.21 80.61 60.915 ;
      RECT  71.79 67.11 71.97 68.815 ;
      RECT  71.79 73.555 71.97 75.26 ;
      RECT  80.43 93.305 80.61 95.01 ;
      RECT  71.79 65.655 71.97 67.36 ;
      RECT  80.43 90.81 80.61 92.515 ;
      RECT  71.79 93.305 71.97 95.01 ;
      RECT  71.79 81.455 71.97 83.16 ;
      RECT  80.43 77.505 80.61 79.21 ;
      RECT  80.43 78.96 80.61 80.665 ;
      RECT  80.43 75.01 80.61 76.715 ;
      RECT  71.79 75.01 71.97 76.715 ;
      RECT  80.43 67.11 80.61 68.815 ;
      RECT  80.43 63.16 80.61 64.865 ;
      RECT  72.75 52.33 72.61 56.1 ;
      RECT  70.43 52.33 70.29 56.1 ;
      RECT  73.41 52.33 73.55 56.1 ;
      RECT  75.73 52.33 75.87 56.1 ;
      RECT  78.99 52.33 78.85 56.1 ;
      RECT  76.67 52.33 76.53 56.1 ;
      RECT  72.61 52.33 72.75 56.1 ;
      RECT  70.29 52.33 70.43 56.1 ;
      RECT  73.41 52.33 73.55 56.1 ;
      RECT  75.73 52.33 75.87 56.1 ;
      RECT  78.85 52.33 78.99 56.1 ;
      RECT  76.53 52.33 76.67 56.1 ;
      RECT  74.06 45.44 74.23 51.07 ;
      RECT  74.44 39.79 74.58 45.21 ;
      RECT  74.87 40.145 75.1 40.515 ;
      RECT  74.87 41.75 75.1 42.13 ;
      RECT  75.22 49.815 75.45 50.185 ;
      RECT  73.6 39.79 73.83 41.06 ;
      RECT  74.44 45.21 74.78 45.5 ;
      RECT  74.06 39.79 74.23 45.21 ;
      RECT  74.0 45.21 74.29 45.44 ;
      RECT  74.77 45.96 75.08 46.3 ;
      RECT  74.44 45.5 74.58 51.07 ;
      RECT  73.55 50.61 73.84 50.91 ;
      RECT  77.72 45.44 77.55 51.07 ;
      RECT  77.34 39.79 77.2 45.21 ;
      RECT  76.91 40.145 76.68 40.515 ;
      RECT  76.91 41.75 76.68 42.13 ;
      RECT  76.56 49.815 76.33 50.185 ;
      RECT  78.18 39.79 77.95 41.06 ;
      RECT  77.34 45.21 77.0 45.5 ;
      RECT  77.72 39.79 77.55 45.21 ;
      RECT  77.78 45.21 77.49 45.44 ;
      RECT  77.01 45.96 76.7 46.3 ;
      RECT  77.34 45.5 77.2 51.07 ;
      RECT  78.23 50.61 77.94 50.91 ;
      RECT  73.6 39.79 73.83 41.06 ;
      RECT  74.06 45.44 74.23 51.07 ;
      RECT  74.44 45.5 74.58 51.07 ;
      RECT  77.95 39.79 78.18 41.06 ;
      RECT  77.55 45.44 77.72 51.07 ;
      RECT  77.2 45.5 77.34 51.07 ;
      RECT  74.145 36.28 74.685 36.45 ;
      RECT  74.245 29.315 74.675 29.545 ;
      RECT  74.59 37.98 74.875 38.27 ;
      RECT  73.575 28.945 75.58 29.115 ;
      RECT  74.72 38.27 74.87 38.53 ;
      RECT  74.355 28.495 74.655 28.775 ;
      RECT  73.575 29.115 73.865 29.255 ;
      RECT  73.71 38.27 73.86 38.53 ;
      RECT  74.145 36.25 74.575 36.28 ;
      RECT  74.145 34.065 74.575 34.295 ;
      RECT  74.75 32.42 75.18 32.625 ;
      RECT  74.145 36.45 74.575 36.48 ;
      RECT  73.705 37.98 73.99 38.27 ;
      RECT  74.175 31.395 74.605 31.625 ;
      RECT  74.815 32.395 75.18 32.42 ;
      RECT  77.635 36.28 77.095 36.45 ;
      RECT  77.535 29.315 77.105 29.545 ;
      RECT  77.19 37.98 76.905 38.27 ;
      RECT  78.205 28.945 76.2 29.115 ;
      RECT  77.06 38.27 76.91 38.53 ;
      RECT  77.425 28.495 77.125 28.775 ;
      RECT  78.205 29.115 77.915 29.255 ;
      RECT  78.07 38.27 77.92 38.53 ;
      RECT  77.635 36.25 77.205 36.28 ;
      RECT  77.635 34.065 77.205 34.295 ;
      RECT  77.03 32.42 76.6 32.625 ;
      RECT  77.635 36.45 77.205 36.48 ;
      RECT  78.075 37.98 77.79 38.27 ;
      RECT  77.605 31.395 77.175 31.625 ;
      RECT  76.965 32.395 76.6 32.42 ;
      RECT  74.355 28.495 74.655 28.775 ;
      RECT  77.125 28.495 77.425 28.775 ;
      RECT  73.71 38.27 73.86 38.53 ;
      RECT  74.72 38.27 74.87 38.53 ;
      RECT  77.92 38.27 78.07 38.53 ;
      RECT  76.91 38.27 77.06 38.53 ;
      RECT  73.08 28.945 79.32 29.085 ;
      RECT  72.61 56.1 72.75 52.33 ;
      RECT  70.29 56.1 70.43 52.33 ;
      RECT  73.6 41.06 73.83 39.79 ;
      RECT  77.95 41.06 78.18 39.79 ;
      RECT  74.355 28.775 74.655 28.495 ;
      RECT  77.125 28.775 77.425 28.495 ;
      RECT  73.08 29.085 79.32 28.945 ;
      RECT  73.41 101.89 73.55 98.12 ;
      RECT  75.73 101.89 75.87 98.12 ;
      RECT  78.99 101.89 78.85 98.12 ;
      RECT  76.67 101.89 76.53 98.12 ;
      RECT  79.65 101.89 79.79 98.12 ;
      RECT  81.97 101.89 82.11 98.12 ;
      RECT  73.41 101.89 73.55 98.12 ;
      RECT  75.73 101.89 75.87 98.12 ;
      RECT  78.85 101.89 78.99 98.12 ;
      RECT  76.53 101.89 76.67 98.12 ;
      RECT  79.65 101.89 79.79 98.12 ;
      RECT  81.97 101.89 82.11 98.12 ;
      RECT  74.06 108.78 74.23 103.15 ;
      RECT  74.44 114.43 74.58 109.01 ;
      RECT  74.87 114.075 75.1 113.705 ;
      RECT  74.87 112.47 75.1 112.09 ;
      RECT  75.22 104.405 75.45 104.035 ;
      RECT  73.6 114.43 73.83 113.16 ;
      RECT  74.44 109.01 74.78 108.72 ;
      RECT  74.06 114.43 74.23 109.01 ;
      RECT  74.0 109.01 74.29 108.78 ;
      RECT  74.77 108.26 75.08 107.92 ;
      RECT  74.44 108.72 74.58 103.15 ;
      RECT  73.55 103.61 73.84 103.31 ;
      RECT  77.72 108.78 77.55 103.15 ;
      RECT  77.34 114.43 77.2 109.01 ;
      RECT  76.91 114.075 76.68 113.705 ;
      RECT  76.91 112.47 76.68 112.09 ;
      RECT  76.56 104.405 76.33 104.035 ;
      RECT  78.18 114.43 77.95 113.16 ;
      RECT  77.34 109.01 77.0 108.72 ;
      RECT  77.72 114.43 77.55 109.01 ;
      RECT  77.78 109.01 77.49 108.78 ;
      RECT  77.01 108.26 76.7 107.92 ;
      RECT  77.34 108.72 77.2 103.15 ;
      RECT  78.23 103.61 77.94 103.31 ;
      RECT  73.6 114.43 73.83 113.16 ;
      RECT  74.06 108.78 74.23 103.15 ;
      RECT  74.44 108.72 74.58 103.15 ;
      RECT  77.95 114.43 78.18 113.16 ;
      RECT  77.55 108.78 77.72 103.15 ;
      RECT  77.2 108.72 77.34 103.15 ;
      RECT  79.65 98.12 79.79 101.89 ;
      RECT  81.97 98.12 82.11 101.89 ;
      RECT  73.6 113.16 73.83 114.43 ;
      RECT  77.95 113.16 78.18 114.43 ;
      RECT  33.78 61.455 33.92 63.43 ;
      RECT  32.42 61.455 32.56 63.43 ;
      RECT  33.78 65.405 33.92 63.43 ;
      RECT  32.42 65.405 32.56 63.43 ;
      RECT  40.34 61.295 40.59 63.465 ;
      RECT  38.22 61.305 38.46 63.465 ;
      RECT  43.65 61.455 43.79 63.43 ;
      RECT  42.29 61.455 42.43 63.43 ;
      RECT  40.34 61.295 40.59 63.465 ;
      RECT  43.65 61.455 43.79 63.43 ;
      RECT  38.22 61.305 38.46 63.465 ;
      RECT  42.29 61.455 42.43 63.43 ;
      RECT  40.34 65.565 40.59 63.395 ;
      RECT  38.22 65.555 38.46 63.395 ;
      RECT  43.65 65.405 43.79 63.43 ;
      RECT  42.29 65.405 42.43 63.43 ;
      RECT  40.34 65.565 40.59 63.395 ;
      RECT  43.65 65.405 43.79 63.43 ;
      RECT  38.22 65.555 38.46 63.395 ;
      RECT  42.29 65.405 42.43 63.43 ;
      RECT  40.34 65.245 40.59 67.415 ;
      RECT  38.22 65.255 38.46 67.415 ;
      RECT  43.65 65.405 43.79 67.38 ;
      RECT  42.29 65.405 42.43 67.38 ;
      RECT  40.34 65.245 40.59 67.415 ;
      RECT  43.65 65.405 43.79 67.38 ;
      RECT  38.22 65.255 38.46 67.415 ;
      RECT  42.29 65.405 42.43 67.38 ;
      RECT  40.34 69.515 40.59 67.345 ;
      RECT  38.22 69.505 38.46 67.345 ;
      RECT  43.65 69.355 43.79 67.38 ;
      RECT  42.29 69.355 42.43 67.38 ;
      RECT  40.34 69.515 40.59 67.345 ;
      RECT  43.65 69.355 43.79 67.38 ;
      RECT  38.22 69.505 38.46 67.345 ;
      RECT  42.29 69.355 42.43 67.38 ;
      RECT  30.24 62.28 30.5 62.6 ;
      RECT  30.64 64.26 30.9 64.58 ;
      RECT  33.78 73.305 33.92 75.28 ;
      RECT  32.42 73.305 32.56 75.28 ;
      RECT  33.78 77.255 33.92 75.28 ;
      RECT  32.42 77.255 32.56 75.28 ;
      RECT  40.34 73.145 40.59 75.315 ;
      RECT  38.22 73.155 38.46 75.315 ;
      RECT  43.65 73.305 43.79 75.28 ;
      RECT  42.29 73.305 42.43 75.28 ;
      RECT  40.34 73.145 40.59 75.315 ;
      RECT  43.65 73.305 43.79 75.28 ;
      RECT  38.22 73.155 38.46 75.315 ;
      RECT  42.29 73.305 42.43 75.28 ;
      RECT  40.34 77.415 40.59 75.245 ;
      RECT  38.22 77.405 38.46 75.245 ;
      RECT  43.65 77.255 43.79 75.28 ;
      RECT  42.29 77.255 42.43 75.28 ;
      RECT  40.34 77.415 40.59 75.245 ;
      RECT  43.65 77.255 43.79 75.28 ;
      RECT  38.22 77.405 38.46 75.245 ;
      RECT  42.29 77.255 42.43 75.28 ;
      RECT  40.34 77.095 40.59 79.265 ;
      RECT  38.22 77.105 38.46 79.265 ;
      RECT  43.65 77.255 43.79 79.23 ;
      RECT  42.29 77.255 42.43 79.23 ;
      RECT  40.34 77.095 40.59 79.265 ;
      RECT  43.65 77.255 43.79 79.23 ;
      RECT  38.22 77.105 38.46 79.265 ;
      RECT  42.29 77.255 42.43 79.23 ;
      RECT  40.34 81.365 40.59 79.195 ;
      RECT  38.22 81.355 38.46 79.195 ;
      RECT  43.65 81.205 43.79 79.23 ;
      RECT  42.29 81.205 42.43 79.23 ;
      RECT  40.34 81.365 40.59 79.195 ;
      RECT  43.65 81.205 43.79 79.23 ;
      RECT  38.22 81.355 38.46 79.195 ;
      RECT  42.29 81.205 42.43 79.23 ;
      RECT  30.24 74.13 30.5 74.45 ;
      RECT  30.64 76.11 30.9 76.43 ;
      RECT  51.41 61.295 51.66 63.465 ;
      RECT  49.29 61.305 49.53 63.465 ;
      RECT  54.72 61.455 54.86 63.43 ;
      RECT  53.36 61.455 53.5 63.43 ;
      RECT  51.41 61.295 51.66 63.465 ;
      RECT  54.72 61.455 54.86 63.43 ;
      RECT  49.29 61.305 49.53 63.465 ;
      RECT  53.36 61.455 53.5 63.43 ;
      RECT  51.41 65.565 51.66 63.395 ;
      RECT  49.29 65.555 49.53 63.395 ;
      RECT  54.72 65.405 54.86 63.43 ;
      RECT  53.36 65.405 53.5 63.43 ;
      RECT  51.41 65.565 51.66 63.395 ;
      RECT  54.72 65.405 54.86 63.43 ;
      RECT  49.29 65.555 49.53 63.395 ;
      RECT  53.36 65.405 53.5 63.43 ;
      RECT  51.41 65.245 51.66 67.415 ;
      RECT  49.29 65.255 49.53 67.415 ;
      RECT  54.72 65.405 54.86 67.38 ;
      RECT  53.36 65.405 53.5 67.38 ;
      RECT  51.41 65.245 51.66 67.415 ;
      RECT  54.72 65.405 54.86 67.38 ;
      RECT  49.29 65.255 49.53 67.415 ;
      RECT  53.36 65.405 53.5 67.38 ;
      RECT  51.41 69.515 51.66 67.345 ;
      RECT  49.29 69.505 49.53 67.345 ;
      RECT  54.72 69.355 54.86 67.38 ;
      RECT  53.36 69.355 53.5 67.38 ;
      RECT  51.41 69.515 51.66 67.345 ;
      RECT  54.72 69.355 54.86 67.38 ;
      RECT  49.29 69.505 49.53 67.345 ;
      RECT  53.36 69.355 53.5 67.38 ;
      RECT  51.41 69.195 51.66 71.365 ;
      RECT  49.29 69.205 49.53 71.365 ;
      RECT  54.72 69.355 54.86 71.33 ;
      RECT  53.36 69.355 53.5 71.33 ;
      RECT  51.41 69.195 51.66 71.365 ;
      RECT  54.72 69.355 54.86 71.33 ;
      RECT  49.29 69.205 49.53 71.365 ;
      RECT  53.36 69.355 53.5 71.33 ;
      RECT  51.41 73.465 51.66 71.295 ;
      RECT  49.29 73.455 49.53 71.295 ;
      RECT  54.72 73.305 54.86 71.33 ;
      RECT  53.36 73.305 53.5 71.33 ;
      RECT  51.41 73.465 51.66 71.295 ;
      RECT  54.72 73.305 54.86 71.33 ;
      RECT  49.29 73.455 49.53 71.295 ;
      RECT  53.36 73.305 53.5 71.33 ;
      RECT  51.41 73.145 51.66 75.315 ;
      RECT  49.29 73.155 49.53 75.315 ;
      RECT  54.72 73.305 54.86 75.28 ;
      RECT  53.36 73.305 53.5 75.28 ;
      RECT  51.41 73.145 51.66 75.315 ;
      RECT  54.72 73.305 54.86 75.28 ;
      RECT  49.29 73.155 49.53 75.315 ;
      RECT  53.36 73.305 53.5 75.28 ;
      RECT  51.41 77.415 51.66 75.245 ;
      RECT  49.29 77.405 49.53 75.245 ;
      RECT  54.72 77.255 54.86 75.28 ;
      RECT  53.36 77.255 53.5 75.28 ;
      RECT  51.41 77.415 51.66 75.245 ;
      RECT  54.72 77.255 54.86 75.28 ;
      RECT  49.29 77.405 49.53 75.245 ;
      RECT  53.36 77.255 53.5 75.28 ;
      RECT  51.41 77.095 51.66 79.265 ;
      RECT  49.29 77.105 49.53 79.265 ;
      RECT  54.72 77.255 54.86 79.23 ;
      RECT  53.36 77.255 53.5 79.23 ;
      RECT  51.41 77.095 51.66 79.265 ;
      RECT  54.72 77.255 54.86 79.23 ;
      RECT  49.29 77.105 49.53 79.265 ;
      RECT  53.36 77.255 53.5 79.23 ;
      RECT  51.41 81.365 51.66 79.195 ;
      RECT  49.29 81.355 49.53 79.195 ;
      RECT  54.72 81.205 54.86 79.23 ;
      RECT  53.36 81.205 53.5 79.23 ;
      RECT  51.41 81.365 51.66 79.195 ;
      RECT  54.72 81.205 54.86 79.23 ;
      RECT  49.29 81.355 49.53 79.195 ;
      RECT  53.36 81.205 53.5 79.23 ;
      RECT  51.41 81.045 51.66 83.215 ;
      RECT  49.29 81.055 49.53 83.215 ;
      RECT  54.72 81.205 54.86 83.18 ;
      RECT  53.36 81.205 53.5 83.18 ;
      RECT  51.41 81.045 51.66 83.215 ;
      RECT  54.72 81.205 54.86 83.18 ;
      RECT  49.29 81.055 49.53 83.215 ;
      RECT  53.36 81.205 53.5 83.18 ;
      RECT  51.41 85.315 51.66 83.145 ;
      RECT  49.29 85.305 49.53 83.145 ;
      RECT  54.72 85.155 54.86 83.18 ;
      RECT  53.36 85.155 53.5 83.18 ;
      RECT  51.41 85.315 51.66 83.145 ;
      RECT  54.72 85.155 54.86 83.18 ;
      RECT  49.29 85.305 49.53 83.145 ;
      RECT  53.36 85.155 53.5 83.18 ;
      RECT  51.41 84.995 51.66 87.165 ;
      RECT  49.29 85.005 49.53 87.165 ;
      RECT  54.72 85.155 54.86 87.13 ;
      RECT  53.36 85.155 53.5 87.13 ;
      RECT  51.41 84.995 51.66 87.165 ;
      RECT  54.72 85.155 54.86 87.13 ;
      RECT  49.29 85.005 49.53 87.165 ;
      RECT  53.36 85.155 53.5 87.13 ;
      RECT  51.41 89.265 51.66 87.095 ;
      RECT  49.29 89.255 49.53 87.095 ;
      RECT  54.72 89.105 54.86 87.13 ;
      RECT  53.36 89.105 53.5 87.13 ;
      RECT  51.41 89.265 51.66 87.095 ;
      RECT  54.72 89.105 54.86 87.13 ;
      RECT  49.29 89.255 49.53 87.095 ;
      RECT  53.36 89.105 53.5 87.13 ;
      RECT  51.41 88.945 51.66 91.115 ;
      RECT  49.29 88.955 49.53 91.115 ;
      RECT  54.72 89.105 54.86 91.08 ;
      RECT  53.36 89.105 53.5 91.08 ;
      RECT  51.41 88.945 51.66 91.115 ;
      RECT  54.72 89.105 54.86 91.08 ;
      RECT  49.29 88.955 49.53 91.115 ;
      RECT  53.36 89.105 53.5 91.08 ;
      RECT  51.41 93.215 51.66 91.045 ;
      RECT  49.29 93.205 49.53 91.045 ;
      RECT  54.72 93.055 54.86 91.08 ;
      RECT  53.36 93.055 53.5 91.08 ;
      RECT  51.41 93.215 51.66 91.045 ;
      RECT  54.72 93.055 54.86 91.08 ;
      RECT  49.29 93.205 49.53 91.045 ;
      RECT  53.36 93.055 53.5 91.08 ;
      RECT  28.16 61.455 28.3 81.205 ;
      RECT  28.56 61.455 28.7 81.205 ;
      RECT  28.96 61.455 29.1 81.205 ;
      RECT  29.36 61.455 29.5 81.205 ;
      RECT  59.02 61.15 59.27 63.32 ;
      RECT  56.9 61.16 57.14 63.32 ;
      RECT  63.65 61.31 63.79 63.285 ;
      RECT  61.16 61.31 61.3 63.285 ;
      RECT  59.02 61.15 59.27 63.32 ;
      RECT  63.65 61.31 63.79 63.285 ;
      RECT  56.9 61.16 57.14 63.32 ;
      RECT  61.16 61.31 61.3 63.285 ;
      RECT  59.02 65.42 59.27 63.25 ;
      RECT  56.9 65.41 57.14 63.25 ;
      RECT  63.65 65.26 63.79 63.285 ;
      RECT  61.16 65.26 61.3 63.285 ;
      RECT  59.02 65.42 59.27 63.25 ;
      RECT  63.65 65.26 63.79 63.285 ;
      RECT  56.9 65.41 57.14 63.25 ;
      RECT  61.16 65.26 61.3 63.285 ;
      RECT  59.02 65.1 59.27 67.27 ;
      RECT  56.9 65.11 57.14 67.27 ;
      RECT  63.65 65.26 63.79 67.235 ;
      RECT  61.16 65.26 61.3 67.235 ;
      RECT  59.02 65.1 59.27 67.27 ;
      RECT  63.65 65.26 63.79 67.235 ;
      RECT  56.9 65.11 57.14 67.27 ;
      RECT  61.16 65.26 61.3 67.235 ;
      RECT  59.02 69.37 59.27 67.2 ;
      RECT  56.9 69.36 57.14 67.2 ;
      RECT  63.65 69.21 63.79 67.235 ;
      RECT  61.16 69.21 61.3 67.235 ;
      RECT  59.02 69.37 59.27 67.2 ;
      RECT  63.65 69.21 63.79 67.235 ;
      RECT  56.9 69.36 57.14 67.2 ;
      RECT  61.16 69.21 61.3 67.235 ;
      RECT  59.02 69.05 59.27 71.22 ;
      RECT  56.9 69.06 57.14 71.22 ;
      RECT  63.65 69.21 63.79 71.185 ;
      RECT  61.16 69.21 61.3 71.185 ;
      RECT  59.02 69.05 59.27 71.22 ;
      RECT  63.65 69.21 63.79 71.185 ;
      RECT  56.9 69.06 57.14 71.22 ;
      RECT  61.16 69.21 61.3 71.185 ;
      RECT  59.02 73.32 59.27 71.15 ;
      RECT  56.9 73.31 57.14 71.15 ;
      RECT  63.65 73.16 63.79 71.185 ;
      RECT  61.16 73.16 61.3 71.185 ;
      RECT  59.02 73.32 59.27 71.15 ;
      RECT  63.65 73.16 63.79 71.185 ;
      RECT  56.9 73.31 57.14 71.15 ;
      RECT  61.16 73.16 61.3 71.185 ;
      RECT  59.02 73.0 59.27 75.17 ;
      RECT  56.9 73.01 57.14 75.17 ;
      RECT  63.65 73.16 63.79 75.135 ;
      RECT  61.16 73.16 61.3 75.135 ;
      RECT  59.02 73.0 59.27 75.17 ;
      RECT  63.65 73.16 63.79 75.135 ;
      RECT  56.9 73.01 57.14 75.17 ;
      RECT  61.16 73.16 61.3 75.135 ;
      RECT  59.02 77.27 59.27 75.1 ;
      RECT  56.9 77.26 57.14 75.1 ;
      RECT  63.65 77.11 63.79 75.135 ;
      RECT  61.16 77.11 61.3 75.135 ;
      RECT  59.02 77.27 59.27 75.1 ;
      RECT  63.65 77.11 63.79 75.135 ;
      RECT  56.9 77.26 57.14 75.1 ;
      RECT  61.16 77.11 61.3 75.135 ;
      RECT  59.02 76.95 59.27 79.12 ;
      RECT  56.9 76.96 57.14 79.12 ;
      RECT  63.65 77.11 63.79 79.085 ;
      RECT  61.16 77.11 61.3 79.085 ;
      RECT  59.02 76.95 59.27 79.12 ;
      RECT  63.65 77.11 63.79 79.085 ;
      RECT  56.9 76.96 57.14 79.12 ;
      RECT  61.16 77.11 61.3 79.085 ;
      RECT  59.02 81.22 59.27 79.05 ;
      RECT  56.9 81.21 57.14 79.05 ;
      RECT  63.65 81.06 63.79 79.085 ;
      RECT  61.16 81.06 61.3 79.085 ;
      RECT  59.02 81.22 59.27 79.05 ;
      RECT  63.65 81.06 63.79 79.085 ;
      RECT  56.9 81.21 57.14 79.05 ;
      RECT  61.16 81.06 61.3 79.085 ;
      RECT  59.02 80.9 59.27 83.07 ;
      RECT  56.9 80.91 57.14 83.07 ;
      RECT  63.65 81.06 63.79 83.035 ;
      RECT  61.16 81.06 61.3 83.035 ;
      RECT  59.02 80.9 59.27 83.07 ;
      RECT  63.65 81.06 63.79 83.035 ;
      RECT  56.9 80.91 57.14 83.07 ;
      RECT  61.16 81.06 61.3 83.035 ;
      RECT  59.02 85.17 59.27 83.0 ;
      RECT  56.9 85.16 57.14 83.0 ;
      RECT  63.65 85.01 63.79 83.035 ;
      RECT  61.16 85.01 61.3 83.035 ;
      RECT  59.02 85.17 59.27 83.0 ;
      RECT  63.65 85.01 63.79 83.035 ;
      RECT  56.9 85.16 57.14 83.0 ;
      RECT  61.16 85.01 61.3 83.035 ;
      RECT  59.02 84.85 59.27 87.02 ;
      RECT  56.9 84.86 57.14 87.02 ;
      RECT  63.65 85.01 63.79 86.985 ;
      RECT  61.16 85.01 61.3 86.985 ;
      RECT  59.02 84.85 59.27 87.02 ;
      RECT  63.65 85.01 63.79 86.985 ;
      RECT  56.9 84.86 57.14 87.02 ;
      RECT  61.16 85.01 61.3 86.985 ;
      RECT  59.02 89.12 59.27 86.95 ;
      RECT  56.9 89.11 57.14 86.95 ;
      RECT  63.65 88.96 63.79 86.985 ;
      RECT  61.16 88.96 61.3 86.985 ;
      RECT  59.02 89.12 59.27 86.95 ;
      RECT  63.65 88.96 63.79 86.985 ;
      RECT  56.9 89.11 57.14 86.95 ;
      RECT  61.16 88.96 61.3 86.985 ;
      RECT  59.02 88.8 59.27 90.97 ;
      RECT  56.9 88.81 57.14 90.97 ;
      RECT  63.65 88.96 63.79 90.935 ;
      RECT  61.16 88.96 61.3 90.935 ;
      RECT  59.02 88.8 59.27 90.97 ;
      RECT  63.65 88.96 63.79 90.935 ;
      RECT  56.9 88.81 57.14 90.97 ;
      RECT  61.16 88.96 61.3 90.935 ;
      RECT  59.02 93.07 59.27 90.9 ;
      RECT  56.9 93.06 57.14 90.9 ;
      RECT  63.65 92.91 63.79 90.935 ;
      RECT  61.16 92.91 61.3 90.935 ;
      RECT  59.02 93.07 59.27 90.9 ;
      RECT  63.65 92.91 63.79 90.935 ;
      RECT  56.9 93.06 57.14 90.9 ;
      RECT  61.16 92.91 61.3 90.935 ;
      RECT  63.65 61.31 63.79 92.91 ;
      RECT  59.075 61.15 59.215 92.91 ;
      RECT  56.95 61.16 57.09 92.91 ;
      RECT  61.16 61.31 61.3 92.91 ;
      RECT  28.16 61.455 28.3 81.205 ;
      RECT  28.56 61.455 28.7 81.205 ;
      RECT  28.96 61.455 29.1 81.205 ;
      RECT  29.36 61.455 29.5 81.205 ;
      RECT  118.62 61.455 118.48 63.43 ;
      RECT  119.98 61.455 119.84 63.43 ;
      RECT  118.62 65.405 118.48 63.43 ;
      RECT  119.98 65.405 119.84 63.43 ;
      RECT  112.06 61.295 111.81 63.465 ;
      RECT  114.18 61.305 113.94 63.465 ;
      RECT  108.75 61.455 108.61 63.43 ;
      RECT  110.11 61.455 109.97 63.43 ;
      RECT  112.06 61.295 111.81 63.465 ;
      RECT  108.75 61.455 108.61 63.43 ;
      RECT  114.18 61.305 113.94 63.465 ;
      RECT  110.11 61.455 109.97 63.43 ;
      RECT  112.06 65.565 111.81 63.395 ;
      RECT  114.18 65.555 113.94 63.395 ;
      RECT  108.75 65.405 108.61 63.43 ;
      RECT  110.11 65.405 109.97 63.43 ;
      RECT  112.06 65.565 111.81 63.395 ;
      RECT  108.75 65.405 108.61 63.43 ;
      RECT  114.18 65.555 113.94 63.395 ;
      RECT  110.11 65.405 109.97 63.43 ;
      RECT  112.06 65.245 111.81 67.415 ;
      RECT  114.18 65.255 113.94 67.415 ;
      RECT  108.75 65.405 108.61 67.38 ;
      RECT  110.11 65.405 109.97 67.38 ;
      RECT  112.06 65.245 111.81 67.415 ;
      RECT  108.75 65.405 108.61 67.38 ;
      RECT  114.18 65.255 113.94 67.415 ;
      RECT  110.11 65.405 109.97 67.38 ;
      RECT  112.06 69.515 111.81 67.345 ;
      RECT  114.18 69.505 113.94 67.345 ;
      RECT  108.75 69.355 108.61 67.38 ;
      RECT  110.11 69.355 109.97 67.38 ;
      RECT  112.06 69.515 111.81 67.345 ;
      RECT  108.75 69.355 108.61 67.38 ;
      RECT  114.18 69.505 113.94 67.345 ;
      RECT  110.11 69.355 109.97 67.38 ;
      RECT  122.16 62.28 121.9 62.6 ;
      RECT  121.76 64.26 121.5 64.58 ;
      RECT  118.62 73.305 118.48 75.28 ;
      RECT  119.98 73.305 119.84 75.28 ;
      RECT  118.62 77.255 118.48 75.28 ;
      RECT  119.98 77.255 119.84 75.28 ;
      RECT  112.06 73.145 111.81 75.315 ;
      RECT  114.18 73.155 113.94 75.315 ;
      RECT  108.75 73.305 108.61 75.28 ;
      RECT  110.11 73.305 109.97 75.28 ;
      RECT  112.06 73.145 111.81 75.315 ;
      RECT  108.75 73.305 108.61 75.28 ;
      RECT  114.18 73.155 113.94 75.315 ;
      RECT  110.11 73.305 109.97 75.28 ;
      RECT  112.06 77.415 111.81 75.245 ;
      RECT  114.18 77.405 113.94 75.245 ;
      RECT  108.75 77.255 108.61 75.28 ;
      RECT  110.11 77.255 109.97 75.28 ;
      RECT  112.06 77.415 111.81 75.245 ;
      RECT  108.75 77.255 108.61 75.28 ;
      RECT  114.18 77.405 113.94 75.245 ;
      RECT  110.11 77.255 109.97 75.28 ;
      RECT  112.06 77.095 111.81 79.265 ;
      RECT  114.18 77.105 113.94 79.265 ;
      RECT  108.75 77.255 108.61 79.23 ;
      RECT  110.11 77.255 109.97 79.23 ;
      RECT  112.06 77.095 111.81 79.265 ;
      RECT  108.75 77.255 108.61 79.23 ;
      RECT  114.18 77.105 113.94 79.265 ;
      RECT  110.11 77.255 109.97 79.23 ;
      RECT  112.06 81.365 111.81 79.195 ;
      RECT  114.18 81.355 113.94 79.195 ;
      RECT  108.75 81.205 108.61 79.23 ;
      RECT  110.11 81.205 109.97 79.23 ;
      RECT  112.06 81.365 111.81 79.195 ;
      RECT  108.75 81.205 108.61 79.23 ;
      RECT  114.18 81.355 113.94 79.195 ;
      RECT  110.11 81.205 109.97 79.23 ;
      RECT  122.16 74.13 121.9 74.45 ;
      RECT  121.76 76.11 121.5 76.43 ;
      RECT  100.99 61.295 100.74 63.465 ;
      RECT  103.11 61.305 102.87 63.465 ;
      RECT  97.68 61.455 97.54 63.43 ;
      RECT  99.04 61.455 98.9 63.43 ;
      RECT  100.99 61.295 100.74 63.465 ;
      RECT  97.68 61.455 97.54 63.43 ;
      RECT  103.11 61.305 102.87 63.465 ;
      RECT  99.04 61.455 98.9 63.43 ;
      RECT  100.99 65.565 100.74 63.395 ;
      RECT  103.11 65.555 102.87 63.395 ;
      RECT  97.68 65.405 97.54 63.43 ;
      RECT  99.04 65.405 98.9 63.43 ;
      RECT  100.99 65.565 100.74 63.395 ;
      RECT  97.68 65.405 97.54 63.43 ;
      RECT  103.11 65.555 102.87 63.395 ;
      RECT  99.04 65.405 98.9 63.43 ;
      RECT  100.99 65.245 100.74 67.415 ;
      RECT  103.11 65.255 102.87 67.415 ;
      RECT  97.68 65.405 97.54 67.38 ;
      RECT  99.04 65.405 98.9 67.38 ;
      RECT  100.99 65.245 100.74 67.415 ;
      RECT  97.68 65.405 97.54 67.38 ;
      RECT  103.11 65.255 102.87 67.415 ;
      RECT  99.04 65.405 98.9 67.38 ;
      RECT  100.99 69.515 100.74 67.345 ;
      RECT  103.11 69.505 102.87 67.345 ;
      RECT  97.68 69.355 97.54 67.38 ;
      RECT  99.04 69.355 98.9 67.38 ;
      RECT  100.99 69.515 100.74 67.345 ;
      RECT  97.68 69.355 97.54 67.38 ;
      RECT  103.11 69.505 102.87 67.345 ;
      RECT  99.04 69.355 98.9 67.38 ;
      RECT  100.99 69.195 100.74 71.365 ;
      RECT  103.11 69.205 102.87 71.365 ;
      RECT  97.68 69.355 97.54 71.33 ;
      RECT  99.04 69.355 98.9 71.33 ;
      RECT  100.99 69.195 100.74 71.365 ;
      RECT  97.68 69.355 97.54 71.33 ;
      RECT  103.11 69.205 102.87 71.365 ;
      RECT  99.04 69.355 98.9 71.33 ;
      RECT  100.99 73.465 100.74 71.295 ;
      RECT  103.11 73.455 102.87 71.295 ;
      RECT  97.68 73.305 97.54 71.33 ;
      RECT  99.04 73.305 98.9 71.33 ;
      RECT  100.99 73.465 100.74 71.295 ;
      RECT  97.68 73.305 97.54 71.33 ;
      RECT  103.11 73.455 102.87 71.295 ;
      RECT  99.04 73.305 98.9 71.33 ;
      RECT  100.99 73.145 100.74 75.315 ;
      RECT  103.11 73.155 102.87 75.315 ;
      RECT  97.68 73.305 97.54 75.28 ;
      RECT  99.04 73.305 98.9 75.28 ;
      RECT  100.99 73.145 100.74 75.315 ;
      RECT  97.68 73.305 97.54 75.28 ;
      RECT  103.11 73.155 102.87 75.315 ;
      RECT  99.04 73.305 98.9 75.28 ;
      RECT  100.99 77.415 100.74 75.245 ;
      RECT  103.11 77.405 102.87 75.245 ;
      RECT  97.68 77.255 97.54 75.28 ;
      RECT  99.04 77.255 98.9 75.28 ;
      RECT  100.99 77.415 100.74 75.245 ;
      RECT  97.68 77.255 97.54 75.28 ;
      RECT  103.11 77.405 102.87 75.245 ;
      RECT  99.04 77.255 98.9 75.28 ;
      RECT  100.99 77.095 100.74 79.265 ;
      RECT  103.11 77.105 102.87 79.265 ;
      RECT  97.68 77.255 97.54 79.23 ;
      RECT  99.04 77.255 98.9 79.23 ;
      RECT  100.99 77.095 100.74 79.265 ;
      RECT  97.68 77.255 97.54 79.23 ;
      RECT  103.11 77.105 102.87 79.265 ;
      RECT  99.04 77.255 98.9 79.23 ;
      RECT  100.99 81.365 100.74 79.195 ;
      RECT  103.11 81.355 102.87 79.195 ;
      RECT  97.68 81.205 97.54 79.23 ;
      RECT  99.04 81.205 98.9 79.23 ;
      RECT  100.99 81.365 100.74 79.195 ;
      RECT  97.68 81.205 97.54 79.23 ;
      RECT  103.11 81.355 102.87 79.195 ;
      RECT  99.04 81.205 98.9 79.23 ;
      RECT  100.99 81.045 100.74 83.215 ;
      RECT  103.11 81.055 102.87 83.215 ;
      RECT  97.68 81.205 97.54 83.18 ;
      RECT  99.04 81.205 98.9 83.18 ;
      RECT  100.99 81.045 100.74 83.215 ;
      RECT  97.68 81.205 97.54 83.18 ;
      RECT  103.11 81.055 102.87 83.215 ;
      RECT  99.04 81.205 98.9 83.18 ;
      RECT  100.99 85.315 100.74 83.145 ;
      RECT  103.11 85.305 102.87 83.145 ;
      RECT  97.68 85.155 97.54 83.18 ;
      RECT  99.04 85.155 98.9 83.18 ;
      RECT  100.99 85.315 100.74 83.145 ;
      RECT  97.68 85.155 97.54 83.18 ;
      RECT  103.11 85.305 102.87 83.145 ;
      RECT  99.04 85.155 98.9 83.18 ;
      RECT  100.99 84.995 100.74 87.165 ;
      RECT  103.11 85.005 102.87 87.165 ;
      RECT  97.68 85.155 97.54 87.13 ;
      RECT  99.04 85.155 98.9 87.13 ;
      RECT  100.99 84.995 100.74 87.165 ;
      RECT  97.68 85.155 97.54 87.13 ;
      RECT  103.11 85.005 102.87 87.165 ;
      RECT  99.04 85.155 98.9 87.13 ;
      RECT  100.99 89.265 100.74 87.095 ;
      RECT  103.11 89.255 102.87 87.095 ;
      RECT  97.68 89.105 97.54 87.13 ;
      RECT  99.04 89.105 98.9 87.13 ;
      RECT  100.99 89.265 100.74 87.095 ;
      RECT  97.68 89.105 97.54 87.13 ;
      RECT  103.11 89.255 102.87 87.095 ;
      RECT  99.04 89.105 98.9 87.13 ;
      RECT  100.99 88.945 100.74 91.115 ;
      RECT  103.11 88.955 102.87 91.115 ;
      RECT  97.68 89.105 97.54 91.08 ;
      RECT  99.04 89.105 98.9 91.08 ;
      RECT  100.99 88.945 100.74 91.115 ;
      RECT  97.68 89.105 97.54 91.08 ;
      RECT  103.11 88.955 102.87 91.115 ;
      RECT  99.04 89.105 98.9 91.08 ;
      RECT  100.99 93.215 100.74 91.045 ;
      RECT  103.11 93.205 102.87 91.045 ;
      RECT  97.68 93.055 97.54 91.08 ;
      RECT  99.04 93.055 98.9 91.08 ;
      RECT  100.99 93.215 100.74 91.045 ;
      RECT  97.68 93.055 97.54 91.08 ;
      RECT  103.11 93.205 102.87 91.045 ;
      RECT  99.04 93.055 98.9 91.08 ;
      RECT  124.24 61.455 124.1 81.205 ;
      RECT  123.84 61.455 123.7 81.205 ;
      RECT  123.44 61.455 123.3 81.205 ;
      RECT  123.04 61.455 122.9 81.205 ;
      RECT  93.38 61.15 93.13 63.32 ;
      RECT  95.5 61.16 95.26 63.32 ;
      RECT  88.75 61.31 88.61 63.285 ;
      RECT  91.24 61.31 91.1 63.285 ;
      RECT  93.38 61.15 93.13 63.32 ;
      RECT  88.75 61.31 88.61 63.285 ;
      RECT  95.5 61.16 95.26 63.32 ;
      RECT  91.24 61.31 91.1 63.285 ;
      RECT  93.38 65.42 93.13 63.25 ;
      RECT  95.5 65.41 95.26 63.25 ;
      RECT  88.75 65.26 88.61 63.285 ;
      RECT  91.24 65.26 91.1 63.285 ;
      RECT  93.38 65.42 93.13 63.25 ;
      RECT  88.75 65.26 88.61 63.285 ;
      RECT  95.5 65.41 95.26 63.25 ;
      RECT  91.24 65.26 91.1 63.285 ;
      RECT  93.38 65.1 93.13 67.27 ;
      RECT  95.5 65.11 95.26 67.27 ;
      RECT  88.75 65.26 88.61 67.235 ;
      RECT  91.24 65.26 91.1 67.235 ;
      RECT  93.38 65.1 93.13 67.27 ;
      RECT  88.75 65.26 88.61 67.235 ;
      RECT  95.5 65.11 95.26 67.27 ;
      RECT  91.24 65.26 91.1 67.235 ;
      RECT  93.38 69.37 93.13 67.2 ;
      RECT  95.5 69.36 95.26 67.2 ;
      RECT  88.75 69.21 88.61 67.235 ;
      RECT  91.24 69.21 91.1 67.235 ;
      RECT  93.38 69.37 93.13 67.2 ;
      RECT  88.75 69.21 88.61 67.235 ;
      RECT  95.5 69.36 95.26 67.2 ;
      RECT  91.24 69.21 91.1 67.235 ;
      RECT  93.38 69.05 93.13 71.22 ;
      RECT  95.5 69.06 95.26 71.22 ;
      RECT  88.75 69.21 88.61 71.185 ;
      RECT  91.24 69.21 91.1 71.185 ;
      RECT  93.38 69.05 93.13 71.22 ;
      RECT  88.75 69.21 88.61 71.185 ;
      RECT  95.5 69.06 95.26 71.22 ;
      RECT  91.24 69.21 91.1 71.185 ;
      RECT  93.38 73.32 93.13 71.15 ;
      RECT  95.5 73.31 95.26 71.15 ;
      RECT  88.75 73.16 88.61 71.185 ;
      RECT  91.24 73.16 91.1 71.185 ;
      RECT  93.38 73.32 93.13 71.15 ;
      RECT  88.75 73.16 88.61 71.185 ;
      RECT  95.5 73.31 95.26 71.15 ;
      RECT  91.24 73.16 91.1 71.185 ;
      RECT  93.38 73.0 93.13 75.17 ;
      RECT  95.5 73.01 95.26 75.17 ;
      RECT  88.75 73.16 88.61 75.135 ;
      RECT  91.24 73.16 91.1 75.135 ;
      RECT  93.38 73.0 93.13 75.17 ;
      RECT  88.75 73.16 88.61 75.135 ;
      RECT  95.5 73.01 95.26 75.17 ;
      RECT  91.24 73.16 91.1 75.135 ;
      RECT  93.38 77.27 93.13 75.1 ;
      RECT  95.5 77.26 95.26 75.1 ;
      RECT  88.75 77.11 88.61 75.135 ;
      RECT  91.24 77.11 91.1 75.135 ;
      RECT  93.38 77.27 93.13 75.1 ;
      RECT  88.75 77.11 88.61 75.135 ;
      RECT  95.5 77.26 95.26 75.1 ;
      RECT  91.24 77.11 91.1 75.135 ;
      RECT  93.38 76.95 93.13 79.12 ;
      RECT  95.5 76.96 95.26 79.12 ;
      RECT  88.75 77.11 88.61 79.085 ;
      RECT  91.24 77.11 91.1 79.085 ;
      RECT  93.38 76.95 93.13 79.12 ;
      RECT  88.75 77.11 88.61 79.085 ;
      RECT  95.5 76.96 95.26 79.12 ;
      RECT  91.24 77.11 91.1 79.085 ;
      RECT  93.38 81.22 93.13 79.05 ;
      RECT  95.5 81.21 95.26 79.05 ;
      RECT  88.75 81.06 88.61 79.085 ;
      RECT  91.24 81.06 91.1 79.085 ;
      RECT  93.38 81.22 93.13 79.05 ;
      RECT  88.75 81.06 88.61 79.085 ;
      RECT  95.5 81.21 95.26 79.05 ;
      RECT  91.24 81.06 91.1 79.085 ;
      RECT  93.38 80.9 93.13 83.07 ;
      RECT  95.5 80.91 95.26 83.07 ;
      RECT  88.75 81.06 88.61 83.035 ;
      RECT  91.24 81.06 91.1 83.035 ;
      RECT  93.38 80.9 93.13 83.07 ;
      RECT  88.75 81.06 88.61 83.035 ;
      RECT  95.5 80.91 95.26 83.07 ;
      RECT  91.24 81.06 91.1 83.035 ;
      RECT  93.38 85.17 93.13 83.0 ;
      RECT  95.5 85.16 95.26 83.0 ;
      RECT  88.75 85.01 88.61 83.035 ;
      RECT  91.24 85.01 91.1 83.035 ;
      RECT  93.38 85.17 93.13 83.0 ;
      RECT  88.75 85.01 88.61 83.035 ;
      RECT  95.5 85.16 95.26 83.0 ;
      RECT  91.24 85.01 91.1 83.035 ;
      RECT  93.38 84.85 93.13 87.02 ;
      RECT  95.5 84.86 95.26 87.02 ;
      RECT  88.75 85.01 88.61 86.985 ;
      RECT  91.24 85.01 91.1 86.985 ;
      RECT  93.38 84.85 93.13 87.02 ;
      RECT  88.75 85.01 88.61 86.985 ;
      RECT  95.5 84.86 95.26 87.02 ;
      RECT  91.24 85.01 91.1 86.985 ;
      RECT  93.38 89.12 93.13 86.95 ;
      RECT  95.5 89.11 95.26 86.95 ;
      RECT  88.75 88.96 88.61 86.985 ;
      RECT  91.24 88.96 91.1 86.985 ;
      RECT  93.38 89.12 93.13 86.95 ;
      RECT  88.75 88.96 88.61 86.985 ;
      RECT  95.5 89.11 95.26 86.95 ;
      RECT  91.24 88.96 91.1 86.985 ;
      RECT  93.38 88.8 93.13 90.97 ;
      RECT  95.5 88.81 95.26 90.97 ;
      RECT  88.75 88.96 88.61 90.935 ;
      RECT  91.24 88.96 91.1 90.935 ;
      RECT  93.38 88.8 93.13 90.97 ;
      RECT  88.75 88.96 88.61 90.935 ;
      RECT  95.5 88.81 95.26 90.97 ;
      RECT  91.24 88.96 91.1 90.935 ;
      RECT  93.38 93.07 93.13 90.9 ;
      RECT  95.5 93.06 95.26 90.9 ;
      RECT  88.75 92.91 88.61 90.935 ;
      RECT  91.24 92.91 91.1 90.935 ;
      RECT  93.38 93.07 93.13 90.9 ;
      RECT  88.75 92.91 88.61 90.935 ;
      RECT  95.5 93.06 95.26 90.9 ;
      RECT  91.24 92.91 91.1 90.935 ;
      RECT  88.75 61.31 88.61 92.91 ;
      RECT  93.325 61.15 93.185 92.91 ;
      RECT  95.45 61.16 95.31 92.91 ;
      RECT  91.24 61.31 91.1 92.91 ;
      RECT  124.24 61.455 124.1 81.205 ;
      RECT  123.84 61.455 123.7 81.205 ;
      RECT  123.44 61.455 123.3 81.205 ;
      RECT  123.04 61.455 122.9 81.205 ;
      RECT  73.6 39.79 73.83 41.06 ;
      RECT  77.95 39.79 78.18 41.06 ;
      RECT  73.6 113.16 73.83 114.43 ;
      RECT  77.95 113.16 78.18 114.43 ;
      RECT  74.355 28.495 74.655 28.775 ;
      RECT  77.125 28.495 77.425 28.775 ;
      RECT  28.16 61.455 28.3 81.205 ;
      RECT  28.56 61.455 28.7 81.205 ;
      RECT  28.96 61.455 29.1 81.205 ;
      RECT  29.36 61.455 29.5 81.205 ;
      RECT  124.1 61.455 124.24 81.205 ;
      RECT  123.7 61.455 123.84 81.205 ;
      RECT  123.3 61.455 123.44 81.205 ;
      RECT  122.9 61.455 123.04 81.205 ;
      RECT  0.505 3.105 0.795 3.135 ;
      RECT  0.18 1.335 0.35 2.305 ;
      RECT  4.48 1.105 4.77 1.335 ;
      RECT  3.175 1.105 3.465 1.335 ;
      RECT  1.895 2.18 2.065 3.46 ;
      RECT  0.12 3.905 0.41 4.135 ;
      RECT  0.12 2.305 0.41 2.535 ;
      RECT  1.845 3.735 2.115 3.78 ;
      RECT  1.845 2.135 2.115 2.18 ;
      RECT  4.48 3.905 4.77 4.135 ;
      RECT  4.48 2.305 4.77 2.535 ;
      RECT  1.425 3.905 1.715 4.135 ;
      RECT  0.18 2.535 0.35 3.905 ;
      RECT  0.12 1.105 0.41 1.335 ;
      RECT  0.505 3.305 0.795 3.335 ;
      RECT  4.54 2.535 4.71 3.905 ;
      RECT  5.41 3.045 5.74 3.305 ;
      RECT  3.235 1.335 3.405 3.905 ;
      RECT  0.505 3.135 1.655 3.305 ;
      RECT  0.685 2.69 1.015 2.95 ;
      RECT  5.43 3.905 5.72 4.135 ;
      RECT  5.02 2.29 5.35 2.55 ;
      RECT  1.485 3.305 1.655 3.905 ;
      RECT  1.845 3.46 2.115 3.505 ;
      RECT  1.845 1.86 2.115 1.905 ;
      RECT  3.175 3.905 3.465 4.135 ;
      RECT  1.835 3.505 2.125 3.735 ;
      RECT  1.835 1.905 2.125 2.135 ;
      RECT  1.425 1.105 1.715 1.335 ;
      RECT  5.49 3.305 5.66 3.905 ;
      RECT  4.54 1.335 4.71 2.305 ;
      RECT  5.49 1.335 5.66 3.045 ;
      RECT  5.43 1.105 5.72 1.335 ;
      RECT  1.485 1.335 1.655 3.135 ;
      RECT  0.505 11.035 0.795 11.005 ;
      RECT  0.18 12.805 0.35 11.835 ;
      RECT  4.48 13.035 4.77 12.805 ;
      RECT  3.175 13.035 3.465 12.805 ;
      RECT  1.895 11.96 2.065 10.68 ;
      RECT  0.12 10.235 0.41 10.005 ;
      RECT  0.12 11.835 0.41 11.605 ;
      RECT  1.845 10.405 2.115 10.36 ;
      RECT  1.845 12.005 2.115 11.96 ;
      RECT  4.48 10.235 4.77 10.005 ;
      RECT  4.48 11.835 4.77 11.605 ;
      RECT  1.425 10.235 1.715 10.005 ;
      RECT  0.18 11.605 0.35 10.235 ;
      RECT  0.12 13.035 0.41 12.805 ;
      RECT  0.505 10.835 0.795 10.805 ;
      RECT  4.54 11.605 4.71 10.235 ;
      RECT  5.41 11.095 5.74 10.835 ;
      RECT  3.235 12.805 3.405 10.235 ;
      RECT  0.505 11.005 1.655 10.835 ;
      RECT  0.685 11.45 1.015 11.19 ;
      RECT  5.43 10.235 5.72 10.005 ;
      RECT  5.02 11.85 5.35 11.59 ;
      RECT  1.485 10.835 1.655 10.235 ;
      RECT  1.845 10.68 2.115 10.635 ;
      RECT  1.845 12.28 2.115 12.235 ;
      RECT  3.175 10.235 3.465 10.005 ;
      RECT  1.835 10.635 2.125 10.405 ;
      RECT  1.835 12.235 2.125 12.005 ;
      RECT  1.425 13.035 1.715 12.805 ;
      RECT  5.49 10.835 5.66 10.235 ;
      RECT  4.54 12.805 4.71 11.835 ;
      RECT  5.49 12.805 5.66 11.095 ;
      RECT  5.43 13.035 5.72 12.805 ;
      RECT  1.485 12.805 1.655 11.005 ;
      RECT  150.785 136.975 150.495 136.945 ;
      RECT  151.11 138.745 150.94 137.775 ;
      RECT  146.81 138.975 146.52 138.745 ;
      RECT  148.115 138.975 147.825 138.745 ;
      RECT  149.395 137.9 149.225 136.62 ;
      RECT  151.17 136.175 150.88 135.945 ;
      RECT  151.17 137.775 150.88 137.545 ;
      RECT  149.445 136.345 149.175 136.3 ;
      RECT  149.445 137.945 149.175 137.9 ;
      RECT  146.81 136.175 146.52 135.945 ;
      RECT  146.81 137.775 146.52 137.545 ;
      RECT  149.865 136.175 149.575 135.945 ;
      RECT  151.11 137.545 150.94 136.175 ;
      RECT  151.17 138.975 150.88 138.745 ;
      RECT  150.785 136.775 150.495 136.745 ;
      RECT  146.75 137.545 146.58 136.175 ;
      RECT  145.88 137.035 145.55 136.775 ;
      RECT  148.055 138.745 147.885 136.175 ;
      RECT  150.785 136.945 149.635 136.775 ;
      RECT  150.605 137.39 150.275 137.13 ;
      RECT  145.86 136.175 145.57 135.945 ;
      RECT  146.27 137.79 145.94 137.53 ;
      RECT  149.805 136.775 149.635 136.175 ;
      RECT  149.445 136.62 149.175 136.575 ;
      RECT  149.445 138.22 149.175 138.175 ;
      RECT  148.115 136.175 147.825 135.945 ;
      RECT  149.455 136.575 149.165 136.345 ;
      RECT  149.455 138.175 149.165 137.945 ;
      RECT  149.865 138.975 149.575 138.745 ;
      RECT  145.8 136.775 145.63 136.175 ;
      RECT  146.75 138.745 146.58 137.775 ;
      RECT  145.8 138.745 145.63 137.035 ;
      RECT  145.86 138.975 145.57 138.745 ;
      RECT  149.805 138.745 149.635 136.945 ;
      RECT  21.895 111.665 22.185 111.695 ;
      RECT  21.57 109.895 21.74 110.865 ;
      RECT  25.87 109.665 26.16 109.895 ;
      RECT  24.565 109.665 24.855 109.895 ;
      RECT  23.285 110.74 23.455 112.02 ;
      RECT  21.51 112.465 21.8 112.695 ;
      RECT  21.51 110.865 21.8 111.095 ;
      RECT  23.235 112.295 23.505 112.34 ;
      RECT  23.235 110.695 23.505 110.74 ;
      RECT  25.87 112.465 26.16 112.695 ;
      RECT  25.87 110.865 26.16 111.095 ;
      RECT  22.815 112.465 23.105 112.695 ;
      RECT  21.57 111.095 21.74 112.465 ;
      RECT  21.51 109.665 21.8 109.895 ;
      RECT  21.895 111.865 22.185 111.895 ;
      RECT  25.93 111.095 26.1 112.465 ;
      RECT  26.8 111.605 27.13 111.865 ;
      RECT  24.625 109.895 24.795 112.465 ;
      RECT  21.895 111.695 23.045 111.865 ;
      RECT  22.075 111.25 22.405 111.51 ;
      RECT  26.82 112.465 27.11 112.695 ;
      RECT  26.41 110.85 26.74 111.11 ;
      RECT  22.875 111.865 23.045 112.465 ;
      RECT  23.235 112.02 23.505 112.065 ;
      RECT  23.235 110.42 23.505 110.465 ;
      RECT  24.565 112.465 24.855 112.695 ;
      RECT  23.225 112.065 23.515 112.295 ;
      RECT  23.225 110.465 23.515 110.695 ;
      RECT  22.815 109.665 23.105 109.895 ;
      RECT  26.88 111.865 27.05 112.465 ;
      RECT  25.93 109.895 26.1 110.865 ;
      RECT  26.88 109.895 27.05 111.605 ;
      RECT  26.82 109.665 27.11 109.895 ;
      RECT  22.875 109.895 23.045 111.695 ;
      RECT  21.895 119.595 22.185 119.565 ;
      RECT  21.57 121.365 21.74 120.395 ;
      RECT  25.87 121.595 26.16 121.365 ;
      RECT  24.565 121.595 24.855 121.365 ;
      RECT  23.285 120.52 23.455 119.24 ;
      RECT  21.51 118.795 21.8 118.565 ;
      RECT  21.51 120.395 21.8 120.165 ;
      RECT  23.235 118.965 23.505 118.92 ;
      RECT  23.235 120.565 23.505 120.52 ;
      RECT  25.87 118.795 26.16 118.565 ;
      RECT  25.87 120.395 26.16 120.165 ;
      RECT  22.815 118.795 23.105 118.565 ;
      RECT  21.57 120.165 21.74 118.795 ;
      RECT  21.51 121.595 21.8 121.365 ;
      RECT  21.895 119.395 22.185 119.365 ;
      RECT  25.93 120.165 26.1 118.795 ;
      RECT  26.8 119.655 27.13 119.395 ;
      RECT  24.625 121.365 24.795 118.795 ;
      RECT  21.895 119.565 23.045 119.395 ;
      RECT  22.075 120.01 22.405 119.75 ;
      RECT  26.82 118.795 27.11 118.565 ;
      RECT  26.41 120.41 26.74 120.15 ;
      RECT  22.875 119.395 23.045 118.795 ;
      RECT  23.235 119.24 23.505 119.195 ;
      RECT  23.235 120.84 23.505 120.795 ;
      RECT  24.565 118.795 24.855 118.565 ;
      RECT  23.225 119.195 23.515 118.965 ;
      RECT  23.225 120.795 23.515 120.565 ;
      RECT  22.815 121.595 23.105 121.365 ;
      RECT  26.88 119.395 27.05 118.795 ;
      RECT  25.93 121.365 26.1 120.395 ;
      RECT  26.88 121.365 27.05 119.655 ;
      RECT  26.82 121.595 27.11 121.365 ;
      RECT  22.875 121.365 23.045 119.565 ;
      RECT  21.895 125.805 22.185 125.835 ;
      RECT  21.57 124.035 21.74 125.005 ;
      RECT  25.87 123.805 26.16 124.035 ;
      RECT  24.565 123.805 24.855 124.035 ;
      RECT  23.285 124.88 23.455 126.16 ;
      RECT  21.51 126.605 21.8 126.835 ;
      RECT  21.51 125.005 21.8 125.235 ;
      RECT  23.235 126.435 23.505 126.48 ;
      RECT  23.235 124.835 23.505 124.88 ;
      RECT  25.87 126.605 26.16 126.835 ;
      RECT  25.87 125.005 26.16 125.235 ;
      RECT  22.815 126.605 23.105 126.835 ;
      RECT  21.57 125.235 21.74 126.605 ;
      RECT  21.51 123.805 21.8 124.035 ;
      RECT  21.895 126.005 22.185 126.035 ;
      RECT  25.93 125.235 26.1 126.605 ;
      RECT  26.8 125.745 27.13 126.005 ;
      RECT  24.625 124.035 24.795 126.605 ;
      RECT  21.895 125.835 23.045 126.005 ;
      RECT  22.075 125.39 22.405 125.65 ;
      RECT  26.82 126.605 27.11 126.835 ;
      RECT  26.41 124.99 26.74 125.25 ;
      RECT  22.875 126.005 23.045 126.605 ;
      RECT  23.235 126.16 23.505 126.205 ;
      RECT  23.235 124.56 23.505 124.605 ;
      RECT  24.565 126.605 24.855 126.835 ;
      RECT  23.225 126.205 23.515 126.435 ;
      RECT  23.225 124.605 23.515 124.835 ;
      RECT  22.815 123.805 23.105 124.035 ;
      RECT  26.88 126.005 27.05 126.605 ;
      RECT  25.93 124.035 26.1 125.005 ;
      RECT  26.88 124.035 27.05 125.745 ;
      RECT  26.82 123.805 27.11 124.035 ;
      RECT  22.875 124.035 23.045 125.835 ;
      RECT  21.895 133.735 22.185 133.705 ;
      RECT  21.57 135.505 21.74 134.535 ;
      RECT  25.87 135.735 26.16 135.505 ;
      RECT  24.565 135.735 24.855 135.505 ;
      RECT  23.285 134.66 23.455 133.38 ;
      RECT  21.51 132.935 21.8 132.705 ;
      RECT  21.51 134.535 21.8 134.305 ;
      RECT  23.235 133.105 23.505 133.06 ;
      RECT  23.235 134.705 23.505 134.66 ;
      RECT  25.87 132.935 26.16 132.705 ;
      RECT  25.87 134.535 26.16 134.305 ;
      RECT  22.815 132.935 23.105 132.705 ;
      RECT  21.57 134.305 21.74 132.935 ;
      RECT  21.51 135.735 21.8 135.505 ;
      RECT  21.895 133.535 22.185 133.505 ;
      RECT  25.93 134.305 26.1 132.935 ;
      RECT  26.8 133.795 27.13 133.535 ;
      RECT  24.625 135.505 24.795 132.935 ;
      RECT  21.895 133.705 23.045 133.535 ;
      RECT  22.075 134.15 22.405 133.89 ;
      RECT  26.82 132.935 27.11 132.705 ;
      RECT  26.41 134.55 26.74 134.29 ;
      RECT  22.875 133.535 23.045 132.935 ;
      RECT  23.235 133.38 23.505 133.335 ;
      RECT  23.235 134.98 23.505 134.935 ;
      RECT  24.565 132.935 24.855 132.705 ;
      RECT  23.225 133.335 23.515 133.105 ;
      RECT  23.225 134.935 23.515 134.705 ;
      RECT  22.815 135.735 23.105 135.505 ;
      RECT  26.88 133.535 27.05 132.935 ;
      RECT  25.93 135.505 26.1 134.535 ;
      RECT  26.88 135.505 27.05 133.795 ;
      RECT  26.82 135.735 27.11 135.505 ;
      RECT  22.875 135.505 23.045 133.705 ;
      RECT  130.925 42.555 130.635 42.525 ;
      RECT  131.25 44.325 131.08 43.355 ;
      RECT  126.95 44.555 126.66 44.325 ;
      RECT  128.255 44.555 127.965 44.325 ;
      RECT  129.535 43.48 129.365 42.2 ;
      RECT  131.31 41.755 131.02 41.525 ;
      RECT  131.31 43.355 131.02 43.125 ;
      RECT  129.585 41.925 129.315 41.88 ;
      RECT  129.585 43.525 129.315 43.48 ;
      RECT  126.95 41.755 126.66 41.525 ;
      RECT  126.95 43.355 126.66 43.125 ;
      RECT  130.005 41.755 129.715 41.525 ;
      RECT  131.25 43.125 131.08 41.755 ;
      RECT  131.31 44.555 131.02 44.325 ;
      RECT  130.925 42.355 130.635 42.325 ;
      RECT  126.89 43.125 126.72 41.755 ;
      RECT  126.02 42.615 125.69 42.355 ;
      RECT  128.195 44.325 128.025 41.755 ;
      RECT  130.925 42.525 129.775 42.355 ;
      RECT  130.745 42.97 130.415 42.71 ;
      RECT  126.0 41.755 125.71 41.525 ;
      RECT  126.41 43.37 126.08 43.11 ;
      RECT  129.945 42.355 129.775 41.755 ;
      RECT  129.585 42.2 129.315 42.155 ;
      RECT  129.585 43.8 129.315 43.755 ;
      RECT  128.255 41.755 127.965 41.525 ;
      RECT  129.595 42.155 129.305 41.925 ;
      RECT  129.595 43.755 129.305 43.525 ;
      RECT  130.005 44.555 129.715 44.325 ;
      RECT  125.94 42.355 125.77 41.755 ;
      RECT  126.89 44.325 126.72 43.355 ;
      RECT  125.94 44.325 125.77 42.615 ;
      RECT  126.0 44.555 125.71 44.325 ;
      RECT  129.945 44.325 129.775 42.525 ;
      RECT  130.925 34.625 130.635 34.655 ;
      RECT  131.25 32.855 131.08 33.825 ;
      RECT  126.95 32.625 126.66 32.855 ;
      RECT  128.255 32.625 127.965 32.855 ;
      RECT  129.535 33.7 129.365 34.98 ;
      RECT  131.31 35.425 131.02 35.655 ;
      RECT  131.31 33.825 131.02 34.055 ;
      RECT  129.585 35.255 129.315 35.3 ;
      RECT  129.585 33.655 129.315 33.7 ;
      RECT  126.95 35.425 126.66 35.655 ;
      RECT  126.95 33.825 126.66 34.055 ;
      RECT  130.005 35.425 129.715 35.655 ;
      RECT  131.25 34.055 131.08 35.425 ;
      RECT  131.31 32.625 131.02 32.855 ;
      RECT  130.925 34.825 130.635 34.855 ;
      RECT  126.89 34.055 126.72 35.425 ;
      RECT  126.02 34.565 125.69 34.825 ;
      RECT  128.195 32.855 128.025 35.425 ;
      RECT  130.925 34.655 129.775 34.825 ;
      RECT  130.745 34.21 130.415 34.47 ;
      RECT  126.0 35.425 125.71 35.655 ;
      RECT  126.41 33.81 126.08 34.07 ;
      RECT  129.945 34.825 129.775 35.425 ;
      RECT  129.585 34.98 129.315 35.025 ;
      RECT  129.585 33.38 129.315 33.425 ;
      RECT  128.255 35.425 127.965 35.655 ;
      RECT  129.595 35.025 129.305 35.255 ;
      RECT  129.595 33.425 129.305 33.655 ;
      RECT  130.005 32.625 129.715 32.855 ;
      RECT  125.94 34.825 125.77 35.425 ;
      RECT  126.89 32.855 126.72 33.825 ;
      RECT  125.94 32.855 125.77 34.565 ;
      RECT  126.0 32.625 125.71 32.855 ;
      RECT  129.945 32.855 129.775 34.655 ;
      RECT  130.925 28.415 130.635 28.385 ;
      RECT  131.25 30.185 131.08 29.215 ;
      RECT  126.95 30.415 126.66 30.185 ;
      RECT  128.255 30.415 127.965 30.185 ;
      RECT  129.535 29.34 129.365 28.06 ;
      RECT  131.31 27.615 131.02 27.385 ;
      RECT  131.31 29.215 131.02 28.985 ;
      RECT  129.585 27.785 129.315 27.74 ;
      RECT  129.585 29.385 129.315 29.34 ;
      RECT  126.95 27.615 126.66 27.385 ;
      RECT  126.95 29.215 126.66 28.985 ;
      RECT  130.005 27.615 129.715 27.385 ;
      RECT  131.25 28.985 131.08 27.615 ;
      RECT  131.31 30.415 131.02 30.185 ;
      RECT  130.925 28.215 130.635 28.185 ;
      RECT  126.89 28.985 126.72 27.615 ;
      RECT  126.02 28.475 125.69 28.215 ;
      RECT  128.195 30.185 128.025 27.615 ;
      RECT  130.925 28.385 129.775 28.215 ;
      RECT  130.745 28.83 130.415 28.57 ;
      RECT  126.0 27.615 125.71 27.385 ;
      RECT  126.41 29.23 126.08 28.97 ;
      RECT  129.945 28.215 129.775 27.615 ;
      RECT  129.585 28.06 129.315 28.015 ;
      RECT  129.585 29.66 129.315 29.615 ;
      RECT  128.255 27.615 127.965 27.385 ;
      RECT  129.595 28.015 129.305 27.785 ;
      RECT  129.595 29.615 129.305 29.385 ;
      RECT  130.005 30.415 129.715 30.185 ;
      RECT  125.94 28.215 125.77 27.615 ;
      RECT  126.89 30.185 126.72 29.215 ;
      RECT  125.94 30.185 125.77 28.475 ;
      RECT  126.0 30.415 125.71 30.185 ;
      RECT  129.945 30.185 129.775 28.385 ;
      RECT  130.925 20.485 130.635 20.515 ;
      RECT  131.25 18.715 131.08 19.685 ;
      RECT  126.95 18.485 126.66 18.715 ;
      RECT  128.255 18.485 127.965 18.715 ;
      RECT  129.535 19.56 129.365 20.84 ;
      RECT  131.31 21.285 131.02 21.515 ;
      RECT  131.31 19.685 131.02 19.915 ;
      RECT  129.585 21.115 129.315 21.16 ;
      RECT  129.585 19.515 129.315 19.56 ;
      RECT  126.95 21.285 126.66 21.515 ;
      RECT  126.95 19.685 126.66 19.915 ;
      RECT  130.005 21.285 129.715 21.515 ;
      RECT  131.25 19.915 131.08 21.285 ;
      RECT  131.31 18.485 131.02 18.715 ;
      RECT  130.925 20.685 130.635 20.715 ;
      RECT  126.89 19.915 126.72 21.285 ;
      RECT  126.02 20.425 125.69 20.685 ;
      RECT  128.195 18.715 128.025 21.285 ;
      RECT  130.925 20.515 129.775 20.685 ;
      RECT  130.745 20.07 130.415 20.33 ;
      RECT  126.0 21.285 125.71 21.515 ;
      RECT  126.41 19.67 126.08 19.93 ;
      RECT  129.945 20.685 129.775 21.285 ;
      RECT  129.585 20.84 129.315 20.885 ;
      RECT  129.585 19.24 129.315 19.285 ;
      RECT  128.255 21.285 127.965 21.515 ;
      RECT  129.595 20.885 129.305 21.115 ;
      RECT  129.595 19.285 129.305 19.515 ;
      RECT  130.005 18.485 129.715 18.715 ;
      RECT  125.94 20.685 125.77 21.285 ;
      RECT  126.89 18.715 126.72 19.685 ;
      RECT  125.94 18.715 125.77 20.425 ;
      RECT  126.0 18.485 125.71 18.715 ;
      RECT  129.945 18.715 129.775 20.515 ;
      RECT  33.575 3.105 33.865 3.135 ;
      RECT  33.25 1.335 33.42 2.305 ;
      RECT  37.55 1.105 37.84 1.335 ;
      RECT  36.245 1.105 36.535 1.335 ;
      RECT  34.965 2.18 35.135 3.46 ;
      RECT  33.19 3.905 33.48 4.135 ;
      RECT  33.19 2.305 33.48 2.535 ;
      RECT  34.915 3.735 35.185 3.78 ;
      RECT  34.915 2.135 35.185 2.18 ;
      RECT  37.55 3.905 37.84 4.135 ;
      RECT  37.55 2.305 37.84 2.535 ;
      RECT  34.495 3.905 34.785 4.135 ;
      RECT  33.25 2.535 33.42 3.905 ;
      RECT  33.19 1.105 33.48 1.335 ;
      RECT  33.575 3.305 33.865 3.335 ;
      RECT  37.61 2.535 37.78 3.905 ;
      RECT  38.48 3.045 38.81 3.305 ;
      RECT  36.305 1.335 36.475 3.905 ;
      RECT  33.575 3.135 34.725 3.305 ;
      RECT  33.755 2.69 34.085 2.95 ;
      RECT  38.5 3.905 38.79 4.135 ;
      RECT  38.09 2.29 38.42 2.55 ;
      RECT  34.555 3.305 34.725 3.905 ;
      RECT  34.915 3.46 35.185 3.505 ;
      RECT  34.915 1.86 35.185 1.905 ;
      RECT  36.245 3.905 36.535 4.135 ;
      RECT  34.905 3.505 35.195 3.735 ;
      RECT  34.905 1.905 35.195 2.135 ;
      RECT  34.495 1.105 34.785 1.335 ;
      RECT  38.56 3.305 38.73 3.905 ;
      RECT  37.61 1.335 37.78 2.305 ;
      RECT  38.56 1.335 38.73 3.045 ;
      RECT  38.5 1.105 38.79 1.335 ;
      RECT  34.555 1.335 34.725 3.135 ;
      RECT  39.415 3.105 39.705 3.135 ;
      RECT  39.09 1.335 39.26 2.305 ;
      RECT  43.39 1.105 43.68 1.335 ;
      RECT  42.085 1.105 42.375 1.335 ;
      RECT  40.805 2.18 40.975 3.46 ;
      RECT  39.03 3.905 39.32 4.135 ;
      RECT  39.03 2.305 39.32 2.535 ;
      RECT  40.755 3.735 41.025 3.78 ;
      RECT  40.755 2.135 41.025 2.18 ;
      RECT  43.39 3.905 43.68 4.135 ;
      RECT  43.39 2.305 43.68 2.535 ;
      RECT  40.335 3.905 40.625 4.135 ;
      RECT  39.09 2.535 39.26 3.905 ;
      RECT  39.03 1.105 39.32 1.335 ;
      RECT  39.415 3.305 39.705 3.335 ;
      RECT  43.45 2.535 43.62 3.905 ;
      RECT  44.32 3.045 44.65 3.305 ;
      RECT  42.145 1.335 42.315 3.905 ;
      RECT  39.415 3.135 40.565 3.305 ;
      RECT  39.595 2.69 39.925 2.95 ;
      RECT  44.34 3.905 44.63 4.135 ;
      RECT  43.93 2.29 44.26 2.55 ;
      RECT  40.395 3.305 40.565 3.905 ;
      RECT  40.755 3.46 41.025 3.505 ;
      RECT  40.755 1.86 41.025 1.905 ;
      RECT  42.085 3.905 42.375 4.135 ;
      RECT  40.745 3.505 41.035 3.735 ;
      RECT  40.745 1.905 41.035 2.135 ;
      RECT  40.335 1.105 40.625 1.335 ;
      RECT  44.4 3.305 44.57 3.905 ;
      RECT  43.45 1.335 43.62 2.305 ;
      RECT  44.4 1.335 44.57 3.045 ;
      RECT  44.34 1.105 44.63 1.335 ;
      RECT  40.395 1.335 40.565 3.135 ;
   LAYER  m2 ;
      RECT  75.48 62.925 75.99 63.165 ;
      RECT  75.48 62.855 75.68 62.925 ;
      RECT  74.01 62.305 74.55 62.685 ;
      RECT  73.08 61.035 74.01 61.585 ;
      RECT  72.87 62.925 73.08 63.165 ;
      RECT  75.99 62.925 76.2 63.165 ;
      RECT  73.08 62.925 75.48 63.165 ;
      RECT  75.27 62.065 75.48 62.135 ;
      RECT  75.99 62.305 76.2 62.685 ;
      RECT  75.27 62.855 75.48 62.925 ;
      RECT  75.48 62.065 75.68 62.135 ;
      RECT  73.08 61.825 75.48 62.065 ;
      RECT  75.99 61.825 76.2 62.065 ;
      RECT  74.01 61.035 74.55 61.585 ;
      RECT  72.87 62.305 74.01 62.685 ;
      RECT  72.87 61.035 73.08 61.585 ;
      POLYGON  75.85 62.305 75.85 62.375 75.48 62.375 75.48 62.615 75.85 62.615 75.85 62.685 75.99 62.685 75.99 62.305 75.85 62.305 ;
      RECT  75.48 61.825 75.99 62.065 ;
      RECT  74.55 61.035 76.2 61.585 ;
      POLYGON  74.55 62.305 74.55 62.685 75.1 62.685 75.1 62.615 75.48 62.615 75.48 62.375 75.1 62.375 75.1 62.305 74.55 62.305 ;
      RECT  72.87 61.825 73.08 62.065 ;
      RECT  75.48 63.645 75.99 63.405 ;
      RECT  75.48 63.715 75.68 63.645 ;
      RECT  74.01 64.265 74.55 63.885 ;
      RECT  73.08 65.535 74.01 64.985 ;
      RECT  72.87 63.645 73.08 63.405 ;
      RECT  75.99 63.645 76.2 63.405 ;
      RECT  73.08 63.645 75.48 63.405 ;
      RECT  75.27 64.505 75.48 64.435 ;
      RECT  75.99 64.265 76.2 63.885 ;
      RECT  75.27 63.715 75.48 63.645 ;
      RECT  75.48 64.505 75.68 64.435 ;
      RECT  73.08 64.745 75.48 64.505 ;
      RECT  75.99 64.745 76.2 64.505 ;
      RECT  74.01 65.535 74.55 64.985 ;
      RECT  72.87 64.265 74.01 63.885 ;
      RECT  72.87 65.535 73.08 64.985 ;
      POLYGON  75.85 64.265 75.85 64.195 75.48 64.195 75.48 63.955 75.85 63.955 75.85 63.885 75.99 63.885 75.99 64.265 75.85 64.265 ;
      RECT  75.48 64.745 75.99 64.505 ;
      RECT  74.55 65.535 76.2 64.985 ;
      POLYGON  74.55 64.265 74.55 63.885 75.1 63.885 75.1 63.955 75.48 63.955 75.48 64.195 75.1 64.195 75.1 64.265 74.55 64.265 ;
      RECT  72.87 64.745 73.08 64.505 ;
      RECT  75.48 66.875 75.99 67.115 ;
      RECT  75.48 66.805 75.68 66.875 ;
      RECT  74.01 66.255 74.55 66.635 ;
      RECT  73.08 64.985 74.01 65.535 ;
      RECT  72.87 66.875 73.08 67.115 ;
      RECT  75.99 66.875 76.2 67.115 ;
      RECT  73.08 66.875 75.48 67.115 ;
      RECT  75.27 66.015 75.48 66.085 ;
      RECT  75.99 66.255 76.2 66.635 ;
      RECT  75.27 66.805 75.48 66.875 ;
      RECT  75.48 66.015 75.68 66.085 ;
      RECT  73.08 65.775 75.48 66.015 ;
      RECT  75.99 65.775 76.2 66.015 ;
      RECT  74.01 64.985 74.55 65.535 ;
      RECT  72.87 66.255 74.01 66.635 ;
      RECT  72.87 64.985 73.08 65.535 ;
      POLYGON  75.85 66.255 75.85 66.325 75.48 66.325 75.48 66.565 75.85 66.565 75.85 66.635 75.99 66.635 75.99 66.255 75.85 66.255 ;
      RECT  75.48 65.775 75.99 66.015 ;
      RECT  74.55 64.985 76.2 65.535 ;
      POLYGON  74.55 66.255 74.55 66.635 75.1 66.635 75.1 66.565 75.48 66.565 75.48 66.325 75.1 66.325 75.1 66.255 74.55 66.255 ;
      RECT  72.87 65.775 73.08 66.015 ;
      RECT  75.48 67.595 75.99 67.355 ;
      RECT  75.48 67.665 75.68 67.595 ;
      RECT  74.01 68.215 74.55 67.835 ;
      RECT  73.08 69.485 74.01 68.935 ;
      RECT  72.87 67.595 73.08 67.355 ;
      RECT  75.99 67.595 76.2 67.355 ;
      RECT  73.08 67.595 75.48 67.355 ;
      RECT  75.27 68.455 75.48 68.385 ;
      RECT  75.99 68.215 76.2 67.835 ;
      RECT  75.27 67.665 75.48 67.595 ;
      RECT  75.48 68.455 75.68 68.385 ;
      RECT  73.08 68.695 75.48 68.455 ;
      RECT  75.99 68.695 76.2 68.455 ;
      RECT  74.01 69.485 74.55 68.935 ;
      RECT  72.87 68.215 74.01 67.835 ;
      RECT  72.87 69.485 73.08 68.935 ;
      POLYGON  75.85 68.215 75.85 68.145 75.48 68.145 75.48 67.905 75.85 67.905 75.85 67.835 75.99 67.835 75.99 68.215 75.85 68.215 ;
      RECT  75.48 68.695 75.99 68.455 ;
      RECT  74.55 69.485 76.2 68.935 ;
      POLYGON  74.55 68.215 74.55 67.835 75.1 67.835 75.1 67.905 75.48 67.905 75.48 68.145 75.1 68.145 75.1 68.215 74.55 68.215 ;
      RECT  72.87 68.695 73.08 68.455 ;
      RECT  75.48 70.825 75.99 71.065 ;
      RECT  75.48 70.755 75.68 70.825 ;
      RECT  74.01 70.205 74.55 70.585 ;
      RECT  73.08 68.935 74.01 69.485 ;
      RECT  72.87 70.825 73.08 71.065 ;
      RECT  75.99 70.825 76.2 71.065 ;
      RECT  73.08 70.825 75.48 71.065 ;
      RECT  75.27 69.965 75.48 70.035 ;
      RECT  75.99 70.205 76.2 70.585 ;
      RECT  75.27 70.755 75.48 70.825 ;
      RECT  75.48 69.965 75.68 70.035 ;
      RECT  73.08 69.725 75.48 69.965 ;
      RECT  75.99 69.725 76.2 69.965 ;
      RECT  74.01 68.935 74.55 69.485 ;
      RECT  72.87 70.205 74.01 70.585 ;
      RECT  72.87 68.935 73.08 69.485 ;
      POLYGON  75.85 70.205 75.85 70.275 75.48 70.275 75.48 70.515 75.85 70.515 75.85 70.585 75.99 70.585 75.99 70.205 75.85 70.205 ;
      RECT  75.48 69.725 75.99 69.965 ;
      RECT  74.55 68.935 76.2 69.485 ;
      POLYGON  74.55 70.205 74.55 70.585 75.1 70.585 75.1 70.515 75.48 70.515 75.48 70.275 75.1 70.275 75.1 70.205 74.55 70.205 ;
      RECT  72.87 69.725 73.08 69.965 ;
      RECT  75.48 71.545 75.99 71.305 ;
      RECT  75.48 71.615 75.68 71.545 ;
      RECT  74.01 72.165 74.55 71.785 ;
      RECT  73.08 73.435 74.01 72.885 ;
      RECT  72.87 71.545 73.08 71.305 ;
      RECT  75.99 71.545 76.2 71.305 ;
      RECT  73.08 71.545 75.48 71.305 ;
      RECT  75.27 72.405 75.48 72.335 ;
      RECT  75.99 72.165 76.2 71.785 ;
      RECT  75.27 71.615 75.48 71.545 ;
      RECT  75.48 72.405 75.68 72.335 ;
      RECT  73.08 72.645 75.48 72.405 ;
      RECT  75.99 72.645 76.2 72.405 ;
      RECT  74.01 73.435 74.55 72.885 ;
      RECT  72.87 72.165 74.01 71.785 ;
      RECT  72.87 73.435 73.08 72.885 ;
      POLYGON  75.85 72.165 75.85 72.095 75.48 72.095 75.48 71.855 75.85 71.855 75.85 71.785 75.99 71.785 75.99 72.165 75.85 72.165 ;
      RECT  75.48 72.645 75.99 72.405 ;
      RECT  74.55 73.435 76.2 72.885 ;
      POLYGON  74.55 72.165 74.55 71.785 75.1 71.785 75.1 71.855 75.48 71.855 75.48 72.095 75.1 72.095 75.1 72.165 74.55 72.165 ;
      RECT  72.87 72.645 73.08 72.405 ;
      RECT  75.48 74.775 75.99 75.015 ;
      RECT  75.48 74.705 75.68 74.775 ;
      RECT  74.01 74.155 74.55 74.535 ;
      RECT  73.08 72.885 74.01 73.435 ;
      RECT  72.87 74.775 73.08 75.015 ;
      RECT  75.99 74.775 76.2 75.015 ;
      RECT  73.08 74.775 75.48 75.015 ;
      RECT  75.27 73.915 75.48 73.985 ;
      RECT  75.99 74.155 76.2 74.535 ;
      RECT  75.27 74.705 75.48 74.775 ;
      RECT  75.48 73.915 75.68 73.985 ;
      RECT  73.08 73.675 75.48 73.915 ;
      RECT  75.99 73.675 76.2 73.915 ;
      RECT  74.01 72.885 74.55 73.435 ;
      RECT  72.87 74.155 74.01 74.535 ;
      RECT  72.87 72.885 73.08 73.435 ;
      POLYGON  75.85 74.155 75.85 74.225 75.48 74.225 75.48 74.465 75.85 74.465 75.85 74.535 75.99 74.535 75.99 74.155 75.85 74.155 ;
      RECT  75.48 73.675 75.99 73.915 ;
      RECT  74.55 72.885 76.2 73.435 ;
      POLYGON  74.55 74.155 74.55 74.535 75.1 74.535 75.1 74.465 75.48 74.465 75.48 74.225 75.1 74.225 75.1 74.155 74.55 74.155 ;
      RECT  72.87 73.675 73.08 73.915 ;
      RECT  75.48 75.495 75.99 75.255 ;
      RECT  75.48 75.565 75.68 75.495 ;
      RECT  74.01 76.115 74.55 75.735 ;
      RECT  73.08 77.385 74.01 76.835 ;
      RECT  72.87 75.495 73.08 75.255 ;
      RECT  75.99 75.495 76.2 75.255 ;
      RECT  73.08 75.495 75.48 75.255 ;
      RECT  75.27 76.355 75.48 76.285 ;
      RECT  75.99 76.115 76.2 75.735 ;
      RECT  75.27 75.565 75.48 75.495 ;
      RECT  75.48 76.355 75.68 76.285 ;
      RECT  73.08 76.595 75.48 76.355 ;
      RECT  75.99 76.595 76.2 76.355 ;
      RECT  74.01 77.385 74.55 76.835 ;
      RECT  72.87 76.115 74.01 75.735 ;
      RECT  72.87 77.385 73.08 76.835 ;
      POLYGON  75.85 76.115 75.85 76.045 75.48 76.045 75.48 75.805 75.85 75.805 75.85 75.735 75.99 75.735 75.99 76.115 75.85 76.115 ;
      RECT  75.48 76.595 75.99 76.355 ;
      RECT  74.55 77.385 76.2 76.835 ;
      POLYGON  74.55 76.115 74.55 75.735 75.1 75.735 75.1 75.805 75.48 75.805 75.48 76.045 75.1 76.045 75.1 76.115 74.55 76.115 ;
      RECT  72.87 76.595 73.08 76.355 ;
      RECT  75.48 78.725 75.99 78.965 ;
      RECT  75.48 78.655 75.68 78.725 ;
      RECT  74.01 78.105 74.55 78.485 ;
      RECT  73.08 76.835 74.01 77.385 ;
      RECT  72.87 78.725 73.08 78.965 ;
      RECT  75.99 78.725 76.2 78.965 ;
      RECT  73.08 78.725 75.48 78.965 ;
      RECT  75.27 77.865 75.48 77.935 ;
      RECT  75.99 78.105 76.2 78.485 ;
      RECT  75.27 78.655 75.48 78.725 ;
      RECT  75.48 77.865 75.68 77.935 ;
      RECT  73.08 77.625 75.48 77.865 ;
      RECT  75.99 77.625 76.2 77.865 ;
      RECT  74.01 76.835 74.55 77.385 ;
      RECT  72.87 78.105 74.01 78.485 ;
      RECT  72.87 76.835 73.08 77.385 ;
      POLYGON  75.85 78.105 75.85 78.175 75.48 78.175 75.48 78.415 75.85 78.415 75.85 78.485 75.99 78.485 75.99 78.105 75.85 78.105 ;
      RECT  75.48 77.625 75.99 77.865 ;
      RECT  74.55 76.835 76.2 77.385 ;
      POLYGON  74.55 78.105 74.55 78.485 75.1 78.485 75.1 78.415 75.48 78.415 75.48 78.175 75.1 78.175 75.1 78.105 74.55 78.105 ;
      RECT  72.87 77.625 73.08 77.865 ;
      RECT  75.48 79.445 75.99 79.205 ;
      RECT  75.48 79.515 75.68 79.445 ;
      RECT  74.01 80.065 74.55 79.685 ;
      RECT  73.08 81.335 74.01 80.785 ;
      RECT  72.87 79.445 73.08 79.205 ;
      RECT  75.99 79.445 76.2 79.205 ;
      RECT  73.08 79.445 75.48 79.205 ;
      RECT  75.27 80.305 75.48 80.235 ;
      RECT  75.99 80.065 76.2 79.685 ;
      RECT  75.27 79.515 75.48 79.445 ;
      RECT  75.48 80.305 75.68 80.235 ;
      RECT  73.08 80.545 75.48 80.305 ;
      RECT  75.99 80.545 76.2 80.305 ;
      RECT  74.01 81.335 74.55 80.785 ;
      RECT  72.87 80.065 74.01 79.685 ;
      RECT  72.87 81.335 73.08 80.785 ;
      POLYGON  75.85 80.065 75.85 79.995 75.48 79.995 75.48 79.755 75.85 79.755 75.85 79.685 75.99 79.685 75.99 80.065 75.85 80.065 ;
      RECT  75.48 80.545 75.99 80.305 ;
      RECT  74.55 81.335 76.2 80.785 ;
      POLYGON  74.55 80.065 74.55 79.685 75.1 79.685 75.1 79.755 75.48 79.755 75.48 79.995 75.1 79.995 75.1 80.065 74.55 80.065 ;
      RECT  72.87 80.545 73.08 80.305 ;
      RECT  75.48 82.675 75.99 82.915 ;
      RECT  75.48 82.605 75.68 82.675 ;
      RECT  74.01 82.055 74.55 82.435 ;
      RECT  73.08 80.785 74.01 81.335 ;
      RECT  72.87 82.675 73.08 82.915 ;
      RECT  75.99 82.675 76.2 82.915 ;
      RECT  73.08 82.675 75.48 82.915 ;
      RECT  75.27 81.815 75.48 81.885 ;
      RECT  75.99 82.055 76.2 82.435 ;
      RECT  75.27 82.605 75.48 82.675 ;
      RECT  75.48 81.815 75.68 81.885 ;
      RECT  73.08 81.575 75.48 81.815 ;
      RECT  75.99 81.575 76.2 81.815 ;
      RECT  74.01 80.785 74.55 81.335 ;
      RECT  72.87 82.055 74.01 82.435 ;
      RECT  72.87 80.785 73.08 81.335 ;
      POLYGON  75.85 82.055 75.85 82.125 75.48 82.125 75.48 82.365 75.85 82.365 75.85 82.435 75.99 82.435 75.99 82.055 75.85 82.055 ;
      RECT  75.48 81.575 75.99 81.815 ;
      RECT  74.55 80.785 76.2 81.335 ;
      POLYGON  74.55 82.055 74.55 82.435 75.1 82.435 75.1 82.365 75.48 82.365 75.48 82.125 75.1 82.125 75.1 82.055 74.55 82.055 ;
      RECT  72.87 81.575 73.08 81.815 ;
      RECT  75.48 83.395 75.99 83.155 ;
      RECT  75.48 83.465 75.68 83.395 ;
      RECT  74.01 84.015 74.55 83.635 ;
      RECT  73.08 85.285 74.01 84.735 ;
      RECT  72.87 83.395 73.08 83.155 ;
      RECT  75.99 83.395 76.2 83.155 ;
      RECT  73.08 83.395 75.48 83.155 ;
      RECT  75.27 84.255 75.48 84.185 ;
      RECT  75.99 84.015 76.2 83.635 ;
      RECT  75.27 83.465 75.48 83.395 ;
      RECT  75.48 84.255 75.68 84.185 ;
      RECT  73.08 84.495 75.48 84.255 ;
      RECT  75.99 84.495 76.2 84.255 ;
      RECT  74.01 85.285 74.55 84.735 ;
      RECT  72.87 84.015 74.01 83.635 ;
      RECT  72.87 85.285 73.08 84.735 ;
      POLYGON  75.85 84.015 75.85 83.945 75.48 83.945 75.48 83.705 75.85 83.705 75.85 83.635 75.99 83.635 75.99 84.015 75.85 84.015 ;
      RECT  75.48 84.495 75.99 84.255 ;
      RECT  74.55 85.285 76.2 84.735 ;
      POLYGON  74.55 84.015 74.55 83.635 75.1 83.635 75.1 83.705 75.48 83.705 75.48 83.945 75.1 83.945 75.1 84.015 74.55 84.015 ;
      RECT  72.87 84.495 73.08 84.255 ;
      RECT  75.48 86.625 75.99 86.865 ;
      RECT  75.48 86.555 75.68 86.625 ;
      RECT  74.01 86.005 74.55 86.385 ;
      RECT  73.08 84.735 74.01 85.285 ;
      RECT  72.87 86.625 73.08 86.865 ;
      RECT  75.99 86.625 76.2 86.865 ;
      RECT  73.08 86.625 75.48 86.865 ;
      RECT  75.27 85.765 75.48 85.835 ;
      RECT  75.99 86.005 76.2 86.385 ;
      RECT  75.27 86.555 75.48 86.625 ;
      RECT  75.48 85.765 75.68 85.835 ;
      RECT  73.08 85.525 75.48 85.765 ;
      RECT  75.99 85.525 76.2 85.765 ;
      RECT  74.01 84.735 74.55 85.285 ;
      RECT  72.87 86.005 74.01 86.385 ;
      RECT  72.87 84.735 73.08 85.285 ;
      POLYGON  75.85 86.005 75.85 86.075 75.48 86.075 75.48 86.315 75.85 86.315 75.85 86.385 75.99 86.385 75.99 86.005 75.85 86.005 ;
      RECT  75.48 85.525 75.99 85.765 ;
      RECT  74.55 84.735 76.2 85.285 ;
      POLYGON  74.55 86.005 74.55 86.385 75.1 86.385 75.1 86.315 75.48 86.315 75.48 86.075 75.1 86.075 75.1 86.005 74.55 86.005 ;
      RECT  72.87 85.525 73.08 85.765 ;
      RECT  75.48 87.345 75.99 87.105 ;
      RECT  75.48 87.415 75.68 87.345 ;
      RECT  74.01 87.965 74.55 87.585 ;
      RECT  73.08 89.235 74.01 88.685 ;
      RECT  72.87 87.345 73.08 87.105 ;
      RECT  75.99 87.345 76.2 87.105 ;
      RECT  73.08 87.345 75.48 87.105 ;
      RECT  75.27 88.205 75.48 88.135 ;
      RECT  75.99 87.965 76.2 87.585 ;
      RECT  75.27 87.415 75.48 87.345 ;
      RECT  75.48 88.205 75.68 88.135 ;
      RECT  73.08 88.445 75.48 88.205 ;
      RECT  75.99 88.445 76.2 88.205 ;
      RECT  74.01 89.235 74.55 88.685 ;
      RECT  72.87 87.965 74.01 87.585 ;
      RECT  72.87 89.235 73.08 88.685 ;
      POLYGON  75.85 87.965 75.85 87.895 75.48 87.895 75.48 87.655 75.85 87.655 75.85 87.585 75.99 87.585 75.99 87.965 75.85 87.965 ;
      RECT  75.48 88.445 75.99 88.205 ;
      RECT  74.55 89.235 76.2 88.685 ;
      POLYGON  74.55 87.965 74.55 87.585 75.1 87.585 75.1 87.655 75.48 87.655 75.48 87.895 75.1 87.895 75.1 87.965 74.55 87.965 ;
      RECT  72.87 88.445 73.08 88.205 ;
      RECT  75.48 90.575 75.99 90.815 ;
      RECT  75.48 90.505 75.68 90.575 ;
      RECT  74.01 89.955 74.55 90.335 ;
      RECT  73.08 88.685 74.01 89.235 ;
      RECT  72.87 90.575 73.08 90.815 ;
      RECT  75.99 90.575 76.2 90.815 ;
      RECT  73.08 90.575 75.48 90.815 ;
      RECT  75.27 89.715 75.48 89.785 ;
      RECT  75.99 89.955 76.2 90.335 ;
      RECT  75.27 90.505 75.48 90.575 ;
      RECT  75.48 89.715 75.68 89.785 ;
      RECT  73.08 89.475 75.48 89.715 ;
      RECT  75.99 89.475 76.2 89.715 ;
      RECT  74.01 88.685 74.55 89.235 ;
      RECT  72.87 89.955 74.01 90.335 ;
      RECT  72.87 88.685 73.08 89.235 ;
      POLYGON  75.85 89.955 75.85 90.025 75.48 90.025 75.48 90.265 75.85 90.265 75.85 90.335 75.99 90.335 75.99 89.955 75.85 89.955 ;
      RECT  75.48 89.475 75.99 89.715 ;
      RECT  74.55 88.685 76.2 89.235 ;
      POLYGON  74.55 89.955 74.55 90.335 75.1 90.335 75.1 90.265 75.48 90.265 75.48 90.025 75.1 90.025 75.1 89.955 74.55 89.955 ;
      RECT  72.87 89.475 73.08 89.715 ;
      RECT  75.48 91.295 75.99 91.055 ;
      RECT  75.48 91.365 75.68 91.295 ;
      RECT  74.01 91.915 74.55 91.535 ;
      RECT  73.08 93.185 74.01 92.635 ;
      RECT  72.87 91.295 73.08 91.055 ;
      RECT  75.99 91.295 76.2 91.055 ;
      RECT  73.08 91.295 75.48 91.055 ;
      RECT  75.27 92.155 75.48 92.085 ;
      RECT  75.99 91.915 76.2 91.535 ;
      RECT  75.27 91.365 75.48 91.295 ;
      RECT  75.48 92.155 75.68 92.085 ;
      RECT  73.08 92.395 75.48 92.155 ;
      RECT  75.99 92.395 76.2 92.155 ;
      RECT  74.01 93.185 74.55 92.635 ;
      RECT  72.87 91.915 74.01 91.535 ;
      RECT  72.87 93.185 73.08 92.635 ;
      POLYGON  75.85 91.915 75.85 91.845 75.48 91.845 75.48 91.605 75.85 91.605 75.85 91.535 75.99 91.535 75.99 91.915 75.85 91.915 ;
      RECT  75.48 92.395 75.99 92.155 ;
      RECT  74.55 93.185 76.2 92.635 ;
      POLYGON  74.55 91.915 74.55 91.535 75.1 91.535 75.1 91.605 75.48 91.605 75.48 91.845 75.1 91.845 75.1 91.915 74.55 91.915 ;
      RECT  72.87 92.395 73.08 92.155 ;
      RECT  76.92 62.925 76.41 63.165 ;
      RECT  76.92 62.855 76.72 62.925 ;
      RECT  78.39 62.305 77.85 62.685 ;
      RECT  79.32 61.035 78.39 61.585 ;
      RECT  79.53 62.925 79.32 63.165 ;
      RECT  76.41 62.925 76.2 63.165 ;
      RECT  79.32 62.925 76.92 63.165 ;
      RECT  77.13 62.065 76.92 62.135 ;
      RECT  76.41 62.305 76.2 62.685 ;
      RECT  77.13 62.855 76.92 62.925 ;
      RECT  76.92 62.065 76.72 62.135 ;
      RECT  79.32 61.825 76.92 62.065 ;
      RECT  76.41 61.825 76.2 62.065 ;
      RECT  78.39 61.035 77.85 61.585 ;
      RECT  79.53 62.305 78.39 62.685 ;
      RECT  79.53 61.035 79.32 61.585 ;
      POLYGON  76.55 62.305 76.55 62.375 76.92 62.375 76.92 62.615 76.55 62.615 76.55 62.685 76.41 62.685 76.41 62.305 76.55 62.305 ;
      RECT  76.92 61.825 76.41 62.065 ;
      RECT  77.85 61.035 76.2 61.585 ;
      POLYGON  77.85 62.305 77.85 62.685 77.3 62.685 77.3 62.615 76.92 62.615 76.92 62.375 77.3 62.375 77.3 62.305 77.85 62.305 ;
      RECT  79.53 61.825 79.32 62.065 ;
      RECT  76.92 63.645 76.41 63.405 ;
      RECT  76.92 63.715 76.72 63.645 ;
      RECT  78.39 64.265 77.85 63.885 ;
      RECT  79.32 65.535 78.39 64.985 ;
      RECT  79.53 63.645 79.32 63.405 ;
      RECT  76.41 63.645 76.2 63.405 ;
      RECT  79.32 63.645 76.92 63.405 ;
      RECT  77.13 64.505 76.92 64.435 ;
      RECT  76.41 64.265 76.2 63.885 ;
      RECT  77.13 63.715 76.92 63.645 ;
      RECT  76.92 64.505 76.72 64.435 ;
      RECT  79.32 64.745 76.92 64.505 ;
      RECT  76.41 64.745 76.2 64.505 ;
      RECT  78.39 65.535 77.85 64.985 ;
      RECT  79.53 64.265 78.39 63.885 ;
      RECT  79.53 65.535 79.32 64.985 ;
      POLYGON  76.55 64.265 76.55 64.195 76.92 64.195 76.92 63.955 76.55 63.955 76.55 63.885 76.41 63.885 76.41 64.265 76.55 64.265 ;
      RECT  76.92 64.745 76.41 64.505 ;
      RECT  77.85 65.535 76.2 64.985 ;
      POLYGON  77.85 64.265 77.85 63.885 77.3 63.885 77.3 63.955 76.92 63.955 76.92 64.195 77.3 64.195 77.3 64.265 77.85 64.265 ;
      RECT  79.53 64.745 79.32 64.505 ;
      RECT  76.92 66.875 76.41 67.115 ;
      RECT  76.92 66.805 76.72 66.875 ;
      RECT  78.39 66.255 77.85 66.635 ;
      RECT  79.32 64.985 78.39 65.535 ;
      RECT  79.53 66.875 79.32 67.115 ;
      RECT  76.41 66.875 76.2 67.115 ;
      RECT  79.32 66.875 76.92 67.115 ;
      RECT  77.13 66.015 76.92 66.085 ;
      RECT  76.41 66.255 76.2 66.635 ;
      RECT  77.13 66.805 76.92 66.875 ;
      RECT  76.92 66.015 76.72 66.085 ;
      RECT  79.32 65.775 76.92 66.015 ;
      RECT  76.41 65.775 76.2 66.015 ;
      RECT  78.39 64.985 77.85 65.535 ;
      RECT  79.53 66.255 78.39 66.635 ;
      RECT  79.53 64.985 79.32 65.535 ;
      POLYGON  76.55 66.255 76.55 66.325 76.92 66.325 76.92 66.565 76.55 66.565 76.55 66.635 76.41 66.635 76.41 66.255 76.55 66.255 ;
      RECT  76.92 65.775 76.41 66.015 ;
      RECT  77.85 64.985 76.2 65.535 ;
      POLYGON  77.85 66.255 77.85 66.635 77.3 66.635 77.3 66.565 76.92 66.565 76.92 66.325 77.3 66.325 77.3 66.255 77.85 66.255 ;
      RECT  79.53 65.775 79.32 66.015 ;
      RECT  76.92 67.595 76.41 67.355 ;
      RECT  76.92 67.665 76.72 67.595 ;
      RECT  78.39 68.215 77.85 67.835 ;
      RECT  79.32 69.485 78.39 68.935 ;
      RECT  79.53 67.595 79.32 67.355 ;
      RECT  76.41 67.595 76.2 67.355 ;
      RECT  79.32 67.595 76.92 67.355 ;
      RECT  77.13 68.455 76.92 68.385 ;
      RECT  76.41 68.215 76.2 67.835 ;
      RECT  77.13 67.665 76.92 67.595 ;
      RECT  76.92 68.455 76.72 68.385 ;
      RECT  79.32 68.695 76.92 68.455 ;
      RECT  76.41 68.695 76.2 68.455 ;
      RECT  78.39 69.485 77.85 68.935 ;
      RECT  79.53 68.215 78.39 67.835 ;
      RECT  79.53 69.485 79.32 68.935 ;
      POLYGON  76.55 68.215 76.55 68.145 76.92 68.145 76.92 67.905 76.55 67.905 76.55 67.835 76.41 67.835 76.41 68.215 76.55 68.215 ;
      RECT  76.92 68.695 76.41 68.455 ;
      RECT  77.85 69.485 76.2 68.935 ;
      POLYGON  77.85 68.215 77.85 67.835 77.3 67.835 77.3 67.905 76.92 67.905 76.92 68.145 77.3 68.145 77.3 68.215 77.85 68.215 ;
      RECT  79.53 68.695 79.32 68.455 ;
      RECT  76.92 70.825 76.41 71.065 ;
      RECT  76.92 70.755 76.72 70.825 ;
      RECT  78.39 70.205 77.85 70.585 ;
      RECT  79.32 68.935 78.39 69.485 ;
      RECT  79.53 70.825 79.32 71.065 ;
      RECT  76.41 70.825 76.2 71.065 ;
      RECT  79.32 70.825 76.92 71.065 ;
      RECT  77.13 69.965 76.92 70.035 ;
      RECT  76.41 70.205 76.2 70.585 ;
      RECT  77.13 70.755 76.92 70.825 ;
      RECT  76.92 69.965 76.72 70.035 ;
      RECT  79.32 69.725 76.92 69.965 ;
      RECT  76.41 69.725 76.2 69.965 ;
      RECT  78.39 68.935 77.85 69.485 ;
      RECT  79.53 70.205 78.39 70.585 ;
      RECT  79.53 68.935 79.32 69.485 ;
      POLYGON  76.55 70.205 76.55 70.275 76.92 70.275 76.92 70.515 76.55 70.515 76.55 70.585 76.41 70.585 76.41 70.205 76.55 70.205 ;
      RECT  76.92 69.725 76.41 69.965 ;
      RECT  77.85 68.935 76.2 69.485 ;
      POLYGON  77.85 70.205 77.85 70.585 77.3 70.585 77.3 70.515 76.92 70.515 76.92 70.275 77.3 70.275 77.3 70.205 77.85 70.205 ;
      RECT  79.53 69.725 79.32 69.965 ;
      RECT  76.92 71.545 76.41 71.305 ;
      RECT  76.92 71.615 76.72 71.545 ;
      RECT  78.39 72.165 77.85 71.785 ;
      RECT  79.32 73.435 78.39 72.885 ;
      RECT  79.53 71.545 79.32 71.305 ;
      RECT  76.41 71.545 76.2 71.305 ;
      RECT  79.32 71.545 76.92 71.305 ;
      RECT  77.13 72.405 76.92 72.335 ;
      RECT  76.41 72.165 76.2 71.785 ;
      RECT  77.13 71.615 76.92 71.545 ;
      RECT  76.92 72.405 76.72 72.335 ;
      RECT  79.32 72.645 76.92 72.405 ;
      RECT  76.41 72.645 76.2 72.405 ;
      RECT  78.39 73.435 77.85 72.885 ;
      RECT  79.53 72.165 78.39 71.785 ;
      RECT  79.53 73.435 79.32 72.885 ;
      POLYGON  76.55 72.165 76.55 72.095 76.92 72.095 76.92 71.855 76.55 71.855 76.55 71.785 76.41 71.785 76.41 72.165 76.55 72.165 ;
      RECT  76.92 72.645 76.41 72.405 ;
      RECT  77.85 73.435 76.2 72.885 ;
      POLYGON  77.85 72.165 77.85 71.785 77.3 71.785 77.3 71.855 76.92 71.855 76.92 72.095 77.3 72.095 77.3 72.165 77.85 72.165 ;
      RECT  79.53 72.645 79.32 72.405 ;
      RECT  76.92 74.775 76.41 75.015 ;
      RECT  76.92 74.705 76.72 74.775 ;
      RECT  78.39 74.155 77.85 74.535 ;
      RECT  79.32 72.885 78.39 73.435 ;
      RECT  79.53 74.775 79.32 75.015 ;
      RECT  76.41 74.775 76.2 75.015 ;
      RECT  79.32 74.775 76.92 75.015 ;
      RECT  77.13 73.915 76.92 73.985 ;
      RECT  76.41 74.155 76.2 74.535 ;
      RECT  77.13 74.705 76.92 74.775 ;
      RECT  76.92 73.915 76.72 73.985 ;
      RECT  79.32 73.675 76.92 73.915 ;
      RECT  76.41 73.675 76.2 73.915 ;
      RECT  78.39 72.885 77.85 73.435 ;
      RECT  79.53 74.155 78.39 74.535 ;
      RECT  79.53 72.885 79.32 73.435 ;
      POLYGON  76.55 74.155 76.55 74.225 76.92 74.225 76.92 74.465 76.55 74.465 76.55 74.535 76.41 74.535 76.41 74.155 76.55 74.155 ;
      RECT  76.92 73.675 76.41 73.915 ;
      RECT  77.85 72.885 76.2 73.435 ;
      POLYGON  77.85 74.155 77.85 74.535 77.3 74.535 77.3 74.465 76.92 74.465 76.92 74.225 77.3 74.225 77.3 74.155 77.85 74.155 ;
      RECT  79.53 73.675 79.32 73.915 ;
      RECT  76.92 75.495 76.41 75.255 ;
      RECT  76.92 75.565 76.72 75.495 ;
      RECT  78.39 76.115 77.85 75.735 ;
      RECT  79.32 77.385 78.39 76.835 ;
      RECT  79.53 75.495 79.32 75.255 ;
      RECT  76.41 75.495 76.2 75.255 ;
      RECT  79.32 75.495 76.92 75.255 ;
      RECT  77.13 76.355 76.92 76.285 ;
      RECT  76.41 76.115 76.2 75.735 ;
      RECT  77.13 75.565 76.92 75.495 ;
      RECT  76.92 76.355 76.72 76.285 ;
      RECT  79.32 76.595 76.92 76.355 ;
      RECT  76.41 76.595 76.2 76.355 ;
      RECT  78.39 77.385 77.85 76.835 ;
      RECT  79.53 76.115 78.39 75.735 ;
      RECT  79.53 77.385 79.32 76.835 ;
      POLYGON  76.55 76.115 76.55 76.045 76.92 76.045 76.92 75.805 76.55 75.805 76.55 75.735 76.41 75.735 76.41 76.115 76.55 76.115 ;
      RECT  76.92 76.595 76.41 76.355 ;
      RECT  77.85 77.385 76.2 76.835 ;
      POLYGON  77.85 76.115 77.85 75.735 77.3 75.735 77.3 75.805 76.92 75.805 76.92 76.045 77.3 76.045 77.3 76.115 77.85 76.115 ;
      RECT  79.53 76.595 79.32 76.355 ;
      RECT  76.92 78.725 76.41 78.965 ;
      RECT  76.92 78.655 76.72 78.725 ;
      RECT  78.39 78.105 77.85 78.485 ;
      RECT  79.32 76.835 78.39 77.385 ;
      RECT  79.53 78.725 79.32 78.965 ;
      RECT  76.41 78.725 76.2 78.965 ;
      RECT  79.32 78.725 76.92 78.965 ;
      RECT  77.13 77.865 76.92 77.935 ;
      RECT  76.41 78.105 76.2 78.485 ;
      RECT  77.13 78.655 76.92 78.725 ;
      RECT  76.92 77.865 76.72 77.935 ;
      RECT  79.32 77.625 76.92 77.865 ;
      RECT  76.41 77.625 76.2 77.865 ;
      RECT  78.39 76.835 77.85 77.385 ;
      RECT  79.53 78.105 78.39 78.485 ;
      RECT  79.53 76.835 79.32 77.385 ;
      POLYGON  76.55 78.105 76.55 78.175 76.92 78.175 76.92 78.415 76.55 78.415 76.55 78.485 76.41 78.485 76.41 78.105 76.55 78.105 ;
      RECT  76.92 77.625 76.41 77.865 ;
      RECT  77.85 76.835 76.2 77.385 ;
      POLYGON  77.85 78.105 77.85 78.485 77.3 78.485 77.3 78.415 76.92 78.415 76.92 78.175 77.3 78.175 77.3 78.105 77.85 78.105 ;
      RECT  79.53 77.625 79.32 77.865 ;
      RECT  76.92 79.445 76.41 79.205 ;
      RECT  76.92 79.515 76.72 79.445 ;
      RECT  78.39 80.065 77.85 79.685 ;
      RECT  79.32 81.335 78.39 80.785 ;
      RECT  79.53 79.445 79.32 79.205 ;
      RECT  76.41 79.445 76.2 79.205 ;
      RECT  79.32 79.445 76.92 79.205 ;
      RECT  77.13 80.305 76.92 80.235 ;
      RECT  76.41 80.065 76.2 79.685 ;
      RECT  77.13 79.515 76.92 79.445 ;
      RECT  76.92 80.305 76.72 80.235 ;
      RECT  79.32 80.545 76.92 80.305 ;
      RECT  76.41 80.545 76.2 80.305 ;
      RECT  78.39 81.335 77.85 80.785 ;
      RECT  79.53 80.065 78.39 79.685 ;
      RECT  79.53 81.335 79.32 80.785 ;
      POLYGON  76.55 80.065 76.55 79.995 76.92 79.995 76.92 79.755 76.55 79.755 76.55 79.685 76.41 79.685 76.41 80.065 76.55 80.065 ;
      RECT  76.92 80.545 76.41 80.305 ;
      RECT  77.85 81.335 76.2 80.785 ;
      POLYGON  77.85 80.065 77.85 79.685 77.3 79.685 77.3 79.755 76.92 79.755 76.92 79.995 77.3 79.995 77.3 80.065 77.85 80.065 ;
      RECT  79.53 80.545 79.32 80.305 ;
      RECT  76.92 82.675 76.41 82.915 ;
      RECT  76.92 82.605 76.72 82.675 ;
      RECT  78.39 82.055 77.85 82.435 ;
      RECT  79.32 80.785 78.39 81.335 ;
      RECT  79.53 82.675 79.32 82.915 ;
      RECT  76.41 82.675 76.2 82.915 ;
      RECT  79.32 82.675 76.92 82.915 ;
      RECT  77.13 81.815 76.92 81.885 ;
      RECT  76.41 82.055 76.2 82.435 ;
      RECT  77.13 82.605 76.92 82.675 ;
      RECT  76.92 81.815 76.72 81.885 ;
      RECT  79.32 81.575 76.92 81.815 ;
      RECT  76.41 81.575 76.2 81.815 ;
      RECT  78.39 80.785 77.85 81.335 ;
      RECT  79.53 82.055 78.39 82.435 ;
      RECT  79.53 80.785 79.32 81.335 ;
      POLYGON  76.55 82.055 76.55 82.125 76.92 82.125 76.92 82.365 76.55 82.365 76.55 82.435 76.41 82.435 76.41 82.055 76.55 82.055 ;
      RECT  76.92 81.575 76.41 81.815 ;
      RECT  77.85 80.785 76.2 81.335 ;
      POLYGON  77.85 82.055 77.85 82.435 77.3 82.435 77.3 82.365 76.92 82.365 76.92 82.125 77.3 82.125 77.3 82.055 77.85 82.055 ;
      RECT  79.53 81.575 79.32 81.815 ;
      RECT  76.92 83.395 76.41 83.155 ;
      RECT  76.92 83.465 76.72 83.395 ;
      RECT  78.39 84.015 77.85 83.635 ;
      RECT  79.32 85.285 78.39 84.735 ;
      RECT  79.53 83.395 79.32 83.155 ;
      RECT  76.41 83.395 76.2 83.155 ;
      RECT  79.32 83.395 76.92 83.155 ;
      RECT  77.13 84.255 76.92 84.185 ;
      RECT  76.41 84.015 76.2 83.635 ;
      RECT  77.13 83.465 76.92 83.395 ;
      RECT  76.92 84.255 76.72 84.185 ;
      RECT  79.32 84.495 76.92 84.255 ;
      RECT  76.41 84.495 76.2 84.255 ;
      RECT  78.39 85.285 77.85 84.735 ;
      RECT  79.53 84.015 78.39 83.635 ;
      RECT  79.53 85.285 79.32 84.735 ;
      POLYGON  76.55 84.015 76.55 83.945 76.92 83.945 76.92 83.705 76.55 83.705 76.55 83.635 76.41 83.635 76.41 84.015 76.55 84.015 ;
      RECT  76.92 84.495 76.41 84.255 ;
      RECT  77.85 85.285 76.2 84.735 ;
      POLYGON  77.85 84.015 77.85 83.635 77.3 83.635 77.3 83.705 76.92 83.705 76.92 83.945 77.3 83.945 77.3 84.015 77.85 84.015 ;
      RECT  79.53 84.495 79.32 84.255 ;
      RECT  76.92 86.625 76.41 86.865 ;
      RECT  76.92 86.555 76.72 86.625 ;
      RECT  78.39 86.005 77.85 86.385 ;
      RECT  79.32 84.735 78.39 85.285 ;
      RECT  79.53 86.625 79.32 86.865 ;
      RECT  76.41 86.625 76.2 86.865 ;
      RECT  79.32 86.625 76.92 86.865 ;
      RECT  77.13 85.765 76.92 85.835 ;
      RECT  76.41 86.005 76.2 86.385 ;
      RECT  77.13 86.555 76.92 86.625 ;
      RECT  76.92 85.765 76.72 85.835 ;
      RECT  79.32 85.525 76.92 85.765 ;
      RECT  76.41 85.525 76.2 85.765 ;
      RECT  78.39 84.735 77.85 85.285 ;
      RECT  79.53 86.005 78.39 86.385 ;
      RECT  79.53 84.735 79.32 85.285 ;
      POLYGON  76.55 86.005 76.55 86.075 76.92 86.075 76.92 86.315 76.55 86.315 76.55 86.385 76.41 86.385 76.41 86.005 76.55 86.005 ;
      RECT  76.92 85.525 76.41 85.765 ;
      RECT  77.85 84.735 76.2 85.285 ;
      POLYGON  77.85 86.005 77.85 86.385 77.3 86.385 77.3 86.315 76.92 86.315 76.92 86.075 77.3 86.075 77.3 86.005 77.85 86.005 ;
      RECT  79.53 85.525 79.32 85.765 ;
      RECT  76.92 87.345 76.41 87.105 ;
      RECT  76.92 87.415 76.72 87.345 ;
      RECT  78.39 87.965 77.85 87.585 ;
      RECT  79.32 89.235 78.39 88.685 ;
      RECT  79.53 87.345 79.32 87.105 ;
      RECT  76.41 87.345 76.2 87.105 ;
      RECT  79.32 87.345 76.92 87.105 ;
      RECT  77.13 88.205 76.92 88.135 ;
      RECT  76.41 87.965 76.2 87.585 ;
      RECT  77.13 87.415 76.92 87.345 ;
      RECT  76.92 88.205 76.72 88.135 ;
      RECT  79.32 88.445 76.92 88.205 ;
      RECT  76.41 88.445 76.2 88.205 ;
      RECT  78.39 89.235 77.85 88.685 ;
      RECT  79.53 87.965 78.39 87.585 ;
      RECT  79.53 89.235 79.32 88.685 ;
      POLYGON  76.55 87.965 76.55 87.895 76.92 87.895 76.92 87.655 76.55 87.655 76.55 87.585 76.41 87.585 76.41 87.965 76.55 87.965 ;
      RECT  76.92 88.445 76.41 88.205 ;
      RECT  77.85 89.235 76.2 88.685 ;
      POLYGON  77.85 87.965 77.85 87.585 77.3 87.585 77.3 87.655 76.92 87.655 76.92 87.895 77.3 87.895 77.3 87.965 77.85 87.965 ;
      RECT  79.53 88.445 79.32 88.205 ;
      RECT  76.92 90.575 76.41 90.815 ;
      RECT  76.92 90.505 76.72 90.575 ;
      RECT  78.39 89.955 77.85 90.335 ;
      RECT  79.32 88.685 78.39 89.235 ;
      RECT  79.53 90.575 79.32 90.815 ;
      RECT  76.41 90.575 76.2 90.815 ;
      RECT  79.32 90.575 76.92 90.815 ;
      RECT  77.13 89.715 76.92 89.785 ;
      RECT  76.41 89.955 76.2 90.335 ;
      RECT  77.13 90.505 76.92 90.575 ;
      RECT  76.92 89.715 76.72 89.785 ;
      RECT  79.32 89.475 76.92 89.715 ;
      RECT  76.41 89.475 76.2 89.715 ;
      RECT  78.39 88.685 77.85 89.235 ;
      RECT  79.53 89.955 78.39 90.335 ;
      RECT  79.53 88.685 79.32 89.235 ;
      POLYGON  76.55 89.955 76.55 90.025 76.92 90.025 76.92 90.265 76.55 90.265 76.55 90.335 76.41 90.335 76.41 89.955 76.55 89.955 ;
      RECT  76.92 89.475 76.41 89.715 ;
      RECT  77.85 88.685 76.2 89.235 ;
      POLYGON  77.85 89.955 77.85 90.335 77.3 90.335 77.3 90.265 76.92 90.265 76.92 90.025 77.3 90.025 77.3 89.955 77.85 89.955 ;
      RECT  79.53 89.475 79.32 89.715 ;
      RECT  76.92 91.295 76.41 91.055 ;
      RECT  76.92 91.365 76.72 91.295 ;
      RECT  78.39 91.915 77.85 91.535 ;
      RECT  79.32 93.185 78.39 92.635 ;
      RECT  79.53 91.295 79.32 91.055 ;
      RECT  76.41 91.295 76.2 91.055 ;
      RECT  79.32 91.295 76.92 91.055 ;
      RECT  77.13 92.155 76.92 92.085 ;
      RECT  76.41 91.915 76.2 91.535 ;
      RECT  77.13 91.365 76.92 91.295 ;
      RECT  76.92 92.155 76.72 92.085 ;
      RECT  79.32 92.395 76.92 92.155 ;
      RECT  76.41 92.395 76.2 92.155 ;
      RECT  78.39 93.185 77.85 92.635 ;
      RECT  79.53 91.915 78.39 91.535 ;
      RECT  79.53 93.185 79.32 92.635 ;
      POLYGON  76.55 91.915 76.55 91.845 76.92 91.845 76.92 91.605 76.55 91.605 76.55 91.535 76.41 91.535 76.41 91.915 76.55 91.915 ;
      RECT  76.92 92.395 76.41 92.155 ;
      RECT  77.85 93.185 76.2 92.635 ;
      POLYGON  77.85 91.915 77.85 91.535 77.3 91.535 77.3 91.605 76.92 91.605 76.92 91.845 77.3 91.845 77.3 91.915 77.85 91.915 ;
      RECT  79.53 92.395 79.32 92.155 ;
      RECT  73.08 62.925 79.32 63.165 ;
      RECT  73.08 61.825 79.32 62.065 ;
      RECT  73.08 63.405 79.32 63.645 ;
      RECT  73.08 64.505 79.32 64.745 ;
      RECT  73.08 66.875 79.32 67.115 ;
      RECT  73.08 65.775 79.32 66.015 ;
      RECT  73.08 67.355 79.32 67.595 ;
      RECT  73.08 68.455 79.32 68.695 ;
      RECT  73.08 70.825 79.32 71.065 ;
      RECT  73.08 69.725 79.32 69.965 ;
      RECT  73.08 71.305 79.32 71.545 ;
      RECT  73.08 72.405 79.32 72.645 ;
      RECT  73.08 74.775 79.32 75.015 ;
      RECT  73.08 73.675 79.32 73.915 ;
      RECT  73.08 75.255 79.32 75.495 ;
      RECT  73.08 76.355 79.32 76.595 ;
      RECT  73.08 78.725 79.32 78.965 ;
      RECT  73.08 77.625 79.32 77.865 ;
      RECT  73.08 79.205 79.32 79.445 ;
      RECT  73.08 80.305 79.32 80.545 ;
      RECT  73.08 82.675 79.32 82.915 ;
      RECT  73.08 81.575 79.32 81.815 ;
      RECT  73.08 83.155 79.32 83.395 ;
      RECT  73.08 84.255 79.32 84.495 ;
      RECT  73.08 86.625 79.32 86.865 ;
      RECT  73.08 85.525 79.32 85.765 ;
      RECT  73.08 87.105 79.32 87.345 ;
      RECT  73.08 88.205 79.32 88.445 ;
      RECT  73.08 90.575 79.32 90.815 ;
      RECT  73.08 89.475 79.32 89.715 ;
      RECT  73.08 91.055 79.32 91.295 ;
      RECT  73.08 92.155 79.32 92.395 ;
      RECT  77.85 61.035 78.39 61.585 ;
      RECT  77.85 82.055 78.39 82.435 ;
      RECT  74.01 78.105 74.55 78.485 ;
      RECT  74.01 89.955 74.55 90.335 ;
      RECT  77.85 74.155 78.39 74.535 ;
      RECT  77.85 76.835 78.39 77.385 ;
      RECT  77.85 91.535 78.39 91.915 ;
      RECT  74.01 67.835 74.55 68.215 ;
      RECT  74.01 87.585 74.55 87.965 ;
      RECT  77.85 63.885 78.39 64.265 ;
      RECT  74.01 86.005 74.55 86.385 ;
      RECT  74.01 62.305 74.55 62.685 ;
      RECT  74.01 72.885 74.55 73.435 ;
      RECT  74.01 61.035 74.55 61.585 ;
      RECT  74.01 66.255 74.55 66.635 ;
      RECT  77.85 86.005 78.39 86.385 ;
      RECT  77.85 87.585 78.39 87.965 ;
      RECT  74.01 80.785 74.55 81.335 ;
      RECT  77.85 71.785 78.39 72.165 ;
      RECT  74.01 91.535 74.55 91.915 ;
      RECT  74.01 83.635 74.55 84.015 ;
      RECT  74.01 79.685 74.55 80.065 ;
      RECT  77.85 67.835 78.39 68.215 ;
      RECT  77.85 92.635 78.39 93.185 ;
      RECT  77.85 83.635 78.39 84.015 ;
      RECT  74.01 75.735 74.55 76.115 ;
      RECT  74.01 82.055 74.55 82.435 ;
      RECT  74.01 84.735 74.55 85.285 ;
      RECT  74.01 64.985 74.55 65.535 ;
      RECT  77.85 62.305 78.39 62.685 ;
      RECT  74.01 92.635 74.55 93.185 ;
      RECT  74.01 74.155 74.55 74.535 ;
      RECT  74.01 71.785 74.55 72.165 ;
      RECT  74.01 63.885 74.55 64.265 ;
      RECT  77.85 80.785 78.39 81.335 ;
      RECT  77.85 89.955 78.39 90.335 ;
      RECT  77.85 78.105 78.39 78.485 ;
      RECT  77.85 72.885 78.39 73.435 ;
      RECT  77.85 68.935 78.39 69.485 ;
      RECT  77.85 75.735 78.39 76.115 ;
      RECT  77.85 64.985 78.39 65.535 ;
      RECT  77.85 84.735 78.39 85.285 ;
      RECT  77.85 66.255 78.39 66.635 ;
      RECT  74.01 68.935 74.55 69.485 ;
      RECT  74.01 76.835 74.55 77.385 ;
      RECT  77.85 79.685 78.39 80.065 ;
      RECT  77.85 88.685 78.39 89.235 ;
      RECT  74.01 88.685 74.55 89.235 ;
      RECT  74.01 70.205 74.55 70.585 ;
      RECT  77.85 70.205 78.39 70.585 ;
      RECT  73.08 58.23 69.96 58.78 ;
      RECT  70.68 59.695 70.17 59.455 ;
      RECT  70.68 59.765 70.48 59.695 ;
      RECT  72.15 60.315 71.61 59.935 ;
      RECT  73.08 61.585 72.15 61.035 ;
      RECT  73.29 59.695 73.08 59.455 ;
      RECT  70.17 59.695 69.96 59.455 ;
      RECT  73.08 59.695 70.68 59.455 ;
      RECT  70.89 60.555 70.68 60.485 ;
      RECT  70.17 60.315 69.96 59.935 ;
      RECT  70.89 59.765 70.68 59.695 ;
      RECT  70.68 60.555 70.48 60.485 ;
      RECT  73.08 60.795 70.68 60.555 ;
      RECT  70.17 60.795 69.96 60.555 ;
      RECT  72.15 61.585 71.61 61.035 ;
      RECT  73.29 60.315 72.15 59.935 ;
      RECT  73.29 61.585 73.08 61.035 ;
      POLYGON  70.31 60.315 70.31 60.245 70.68 60.245 70.68 60.005 70.31 60.005 70.31 59.935 70.17 59.935 70.17 60.315 70.31 60.315 ;
      RECT  70.68 60.795 70.17 60.555 ;
      RECT  71.61 61.585 69.96 61.035 ;
      POLYGON  71.61 60.315 71.61 59.935 71.06 59.935 71.06 60.005 70.68 60.005 70.68 60.245 71.06 60.245 71.06 60.315 71.61 60.315 ;
      RECT  73.29 60.795 73.08 60.555 ;
      RECT  70.68 62.925 70.17 63.165 ;
      RECT  70.68 62.855 70.48 62.925 ;
      RECT  72.15 62.305 71.61 62.685 ;
      RECT  73.08 61.035 72.15 61.585 ;
      RECT  73.29 62.925 73.08 63.165 ;
      RECT  70.17 62.925 69.96 63.165 ;
      RECT  73.08 62.925 70.68 63.165 ;
      RECT  70.89 62.065 70.68 62.135 ;
      RECT  70.17 62.305 69.96 62.685 ;
      RECT  70.89 62.855 70.68 62.925 ;
      RECT  70.68 62.065 70.48 62.135 ;
      RECT  73.08 61.825 70.68 62.065 ;
      RECT  70.17 61.825 69.96 62.065 ;
      RECT  72.15 61.035 71.61 61.585 ;
      RECT  73.29 62.305 72.15 62.685 ;
      RECT  73.29 61.035 73.08 61.585 ;
      POLYGON  70.31 62.305 70.31 62.375 70.68 62.375 70.68 62.615 70.31 62.615 70.31 62.685 70.17 62.685 70.17 62.305 70.31 62.305 ;
      RECT  70.68 61.825 70.17 62.065 ;
      RECT  71.61 61.035 69.96 61.585 ;
      POLYGON  71.61 62.305 71.61 62.685 71.06 62.685 71.06 62.615 70.68 62.615 70.68 62.375 71.06 62.375 71.06 62.305 71.61 62.305 ;
      RECT  73.29 61.825 73.08 62.065 ;
      RECT  70.68 63.645 70.17 63.405 ;
      RECT  70.68 63.715 70.48 63.645 ;
      RECT  72.15 64.265 71.61 63.885 ;
      RECT  73.08 65.535 72.15 64.985 ;
      RECT  73.29 63.645 73.08 63.405 ;
      RECT  70.17 63.645 69.96 63.405 ;
      RECT  73.08 63.645 70.68 63.405 ;
      RECT  70.89 64.505 70.68 64.435 ;
      RECT  70.17 64.265 69.96 63.885 ;
      RECT  70.89 63.715 70.68 63.645 ;
      RECT  70.68 64.505 70.48 64.435 ;
      RECT  73.08 64.745 70.68 64.505 ;
      RECT  70.17 64.745 69.96 64.505 ;
      RECT  72.15 65.535 71.61 64.985 ;
      RECT  73.29 64.265 72.15 63.885 ;
      RECT  73.29 65.535 73.08 64.985 ;
      POLYGON  70.31 64.265 70.31 64.195 70.68 64.195 70.68 63.955 70.31 63.955 70.31 63.885 70.17 63.885 70.17 64.265 70.31 64.265 ;
      RECT  70.68 64.745 70.17 64.505 ;
      RECT  71.61 65.535 69.96 64.985 ;
      POLYGON  71.61 64.265 71.61 63.885 71.06 63.885 71.06 63.955 70.68 63.955 70.68 64.195 71.06 64.195 71.06 64.265 71.61 64.265 ;
      RECT  73.29 64.745 73.08 64.505 ;
      RECT  70.68 66.875 70.17 67.115 ;
      RECT  70.68 66.805 70.48 66.875 ;
      RECT  72.15 66.255 71.61 66.635 ;
      RECT  73.08 64.985 72.15 65.535 ;
      RECT  73.29 66.875 73.08 67.115 ;
      RECT  70.17 66.875 69.96 67.115 ;
      RECT  73.08 66.875 70.68 67.115 ;
      RECT  70.89 66.015 70.68 66.085 ;
      RECT  70.17 66.255 69.96 66.635 ;
      RECT  70.89 66.805 70.68 66.875 ;
      RECT  70.68 66.015 70.48 66.085 ;
      RECT  73.08 65.775 70.68 66.015 ;
      RECT  70.17 65.775 69.96 66.015 ;
      RECT  72.15 64.985 71.61 65.535 ;
      RECT  73.29 66.255 72.15 66.635 ;
      RECT  73.29 64.985 73.08 65.535 ;
      POLYGON  70.31 66.255 70.31 66.325 70.68 66.325 70.68 66.565 70.31 66.565 70.31 66.635 70.17 66.635 70.17 66.255 70.31 66.255 ;
      RECT  70.68 65.775 70.17 66.015 ;
      RECT  71.61 64.985 69.96 65.535 ;
      POLYGON  71.61 66.255 71.61 66.635 71.06 66.635 71.06 66.565 70.68 66.565 70.68 66.325 71.06 66.325 71.06 66.255 71.61 66.255 ;
      RECT  73.29 65.775 73.08 66.015 ;
      RECT  70.68 67.595 70.17 67.355 ;
      RECT  70.68 67.665 70.48 67.595 ;
      RECT  72.15 68.215 71.61 67.835 ;
      RECT  73.08 69.485 72.15 68.935 ;
      RECT  73.29 67.595 73.08 67.355 ;
      RECT  70.17 67.595 69.96 67.355 ;
      RECT  73.08 67.595 70.68 67.355 ;
      RECT  70.89 68.455 70.68 68.385 ;
      RECT  70.17 68.215 69.96 67.835 ;
      RECT  70.89 67.665 70.68 67.595 ;
      RECT  70.68 68.455 70.48 68.385 ;
      RECT  73.08 68.695 70.68 68.455 ;
      RECT  70.17 68.695 69.96 68.455 ;
      RECT  72.15 69.485 71.61 68.935 ;
      RECT  73.29 68.215 72.15 67.835 ;
      RECT  73.29 69.485 73.08 68.935 ;
      POLYGON  70.31 68.215 70.31 68.145 70.68 68.145 70.68 67.905 70.31 67.905 70.31 67.835 70.17 67.835 70.17 68.215 70.31 68.215 ;
      RECT  70.68 68.695 70.17 68.455 ;
      RECT  71.61 69.485 69.96 68.935 ;
      POLYGON  71.61 68.215 71.61 67.835 71.06 67.835 71.06 67.905 70.68 67.905 70.68 68.145 71.06 68.145 71.06 68.215 71.61 68.215 ;
      RECT  73.29 68.695 73.08 68.455 ;
      RECT  70.68 70.825 70.17 71.065 ;
      RECT  70.68 70.755 70.48 70.825 ;
      RECT  72.15 70.205 71.61 70.585 ;
      RECT  73.08 68.935 72.15 69.485 ;
      RECT  73.29 70.825 73.08 71.065 ;
      RECT  70.17 70.825 69.96 71.065 ;
      RECT  73.08 70.825 70.68 71.065 ;
      RECT  70.89 69.965 70.68 70.035 ;
      RECT  70.17 70.205 69.96 70.585 ;
      RECT  70.89 70.755 70.68 70.825 ;
      RECT  70.68 69.965 70.48 70.035 ;
      RECT  73.08 69.725 70.68 69.965 ;
      RECT  70.17 69.725 69.96 69.965 ;
      RECT  72.15 68.935 71.61 69.485 ;
      RECT  73.29 70.205 72.15 70.585 ;
      RECT  73.29 68.935 73.08 69.485 ;
      POLYGON  70.31 70.205 70.31 70.275 70.68 70.275 70.68 70.515 70.31 70.515 70.31 70.585 70.17 70.585 70.17 70.205 70.31 70.205 ;
      RECT  70.68 69.725 70.17 69.965 ;
      RECT  71.61 68.935 69.96 69.485 ;
      POLYGON  71.61 70.205 71.61 70.585 71.06 70.585 71.06 70.515 70.68 70.515 70.68 70.275 71.06 70.275 71.06 70.205 71.61 70.205 ;
      RECT  73.29 69.725 73.08 69.965 ;
      RECT  70.68 71.545 70.17 71.305 ;
      RECT  70.68 71.615 70.48 71.545 ;
      RECT  72.15 72.165 71.61 71.785 ;
      RECT  73.08 73.435 72.15 72.885 ;
      RECT  73.29 71.545 73.08 71.305 ;
      RECT  70.17 71.545 69.96 71.305 ;
      RECT  73.08 71.545 70.68 71.305 ;
      RECT  70.89 72.405 70.68 72.335 ;
      RECT  70.17 72.165 69.96 71.785 ;
      RECT  70.89 71.615 70.68 71.545 ;
      RECT  70.68 72.405 70.48 72.335 ;
      RECT  73.08 72.645 70.68 72.405 ;
      RECT  70.17 72.645 69.96 72.405 ;
      RECT  72.15 73.435 71.61 72.885 ;
      RECT  73.29 72.165 72.15 71.785 ;
      RECT  73.29 73.435 73.08 72.885 ;
      POLYGON  70.31 72.165 70.31 72.095 70.68 72.095 70.68 71.855 70.31 71.855 70.31 71.785 70.17 71.785 70.17 72.165 70.31 72.165 ;
      RECT  70.68 72.645 70.17 72.405 ;
      RECT  71.61 73.435 69.96 72.885 ;
      POLYGON  71.61 72.165 71.61 71.785 71.06 71.785 71.06 71.855 70.68 71.855 70.68 72.095 71.06 72.095 71.06 72.165 71.61 72.165 ;
      RECT  73.29 72.645 73.08 72.405 ;
      RECT  70.68 74.775 70.17 75.015 ;
      RECT  70.68 74.705 70.48 74.775 ;
      RECT  72.15 74.155 71.61 74.535 ;
      RECT  73.08 72.885 72.15 73.435 ;
      RECT  73.29 74.775 73.08 75.015 ;
      RECT  70.17 74.775 69.96 75.015 ;
      RECT  73.08 74.775 70.68 75.015 ;
      RECT  70.89 73.915 70.68 73.985 ;
      RECT  70.17 74.155 69.96 74.535 ;
      RECT  70.89 74.705 70.68 74.775 ;
      RECT  70.68 73.915 70.48 73.985 ;
      RECT  73.08 73.675 70.68 73.915 ;
      RECT  70.17 73.675 69.96 73.915 ;
      RECT  72.15 72.885 71.61 73.435 ;
      RECT  73.29 74.155 72.15 74.535 ;
      RECT  73.29 72.885 73.08 73.435 ;
      POLYGON  70.31 74.155 70.31 74.225 70.68 74.225 70.68 74.465 70.31 74.465 70.31 74.535 70.17 74.535 70.17 74.155 70.31 74.155 ;
      RECT  70.68 73.675 70.17 73.915 ;
      RECT  71.61 72.885 69.96 73.435 ;
      POLYGON  71.61 74.155 71.61 74.535 71.06 74.535 71.06 74.465 70.68 74.465 70.68 74.225 71.06 74.225 71.06 74.155 71.61 74.155 ;
      RECT  73.29 73.675 73.08 73.915 ;
      RECT  70.68 75.495 70.17 75.255 ;
      RECT  70.68 75.565 70.48 75.495 ;
      RECT  72.15 76.115 71.61 75.735 ;
      RECT  73.08 77.385 72.15 76.835 ;
      RECT  73.29 75.495 73.08 75.255 ;
      RECT  70.17 75.495 69.96 75.255 ;
      RECT  73.08 75.495 70.68 75.255 ;
      RECT  70.89 76.355 70.68 76.285 ;
      RECT  70.17 76.115 69.96 75.735 ;
      RECT  70.89 75.565 70.68 75.495 ;
      RECT  70.68 76.355 70.48 76.285 ;
      RECT  73.08 76.595 70.68 76.355 ;
      RECT  70.17 76.595 69.96 76.355 ;
      RECT  72.15 77.385 71.61 76.835 ;
      RECT  73.29 76.115 72.15 75.735 ;
      RECT  73.29 77.385 73.08 76.835 ;
      POLYGON  70.31 76.115 70.31 76.045 70.68 76.045 70.68 75.805 70.31 75.805 70.31 75.735 70.17 75.735 70.17 76.115 70.31 76.115 ;
      RECT  70.68 76.595 70.17 76.355 ;
      RECT  71.61 77.385 69.96 76.835 ;
      POLYGON  71.61 76.115 71.61 75.735 71.06 75.735 71.06 75.805 70.68 75.805 70.68 76.045 71.06 76.045 71.06 76.115 71.61 76.115 ;
      RECT  73.29 76.595 73.08 76.355 ;
      RECT  70.68 78.725 70.17 78.965 ;
      RECT  70.68 78.655 70.48 78.725 ;
      RECT  72.15 78.105 71.61 78.485 ;
      RECT  73.08 76.835 72.15 77.385 ;
      RECT  73.29 78.725 73.08 78.965 ;
      RECT  70.17 78.725 69.96 78.965 ;
      RECT  73.08 78.725 70.68 78.965 ;
      RECT  70.89 77.865 70.68 77.935 ;
      RECT  70.17 78.105 69.96 78.485 ;
      RECT  70.89 78.655 70.68 78.725 ;
      RECT  70.68 77.865 70.48 77.935 ;
      RECT  73.08 77.625 70.68 77.865 ;
      RECT  70.17 77.625 69.96 77.865 ;
      RECT  72.15 76.835 71.61 77.385 ;
      RECT  73.29 78.105 72.15 78.485 ;
      RECT  73.29 76.835 73.08 77.385 ;
      POLYGON  70.31 78.105 70.31 78.175 70.68 78.175 70.68 78.415 70.31 78.415 70.31 78.485 70.17 78.485 70.17 78.105 70.31 78.105 ;
      RECT  70.68 77.625 70.17 77.865 ;
      RECT  71.61 76.835 69.96 77.385 ;
      POLYGON  71.61 78.105 71.61 78.485 71.06 78.485 71.06 78.415 70.68 78.415 70.68 78.175 71.06 78.175 71.06 78.105 71.61 78.105 ;
      RECT  73.29 77.625 73.08 77.865 ;
      RECT  70.68 79.445 70.17 79.205 ;
      RECT  70.68 79.515 70.48 79.445 ;
      RECT  72.15 80.065 71.61 79.685 ;
      RECT  73.08 81.335 72.15 80.785 ;
      RECT  73.29 79.445 73.08 79.205 ;
      RECT  70.17 79.445 69.96 79.205 ;
      RECT  73.08 79.445 70.68 79.205 ;
      RECT  70.89 80.305 70.68 80.235 ;
      RECT  70.17 80.065 69.96 79.685 ;
      RECT  70.89 79.515 70.68 79.445 ;
      RECT  70.68 80.305 70.48 80.235 ;
      RECT  73.08 80.545 70.68 80.305 ;
      RECT  70.17 80.545 69.96 80.305 ;
      RECT  72.15 81.335 71.61 80.785 ;
      RECT  73.29 80.065 72.15 79.685 ;
      RECT  73.29 81.335 73.08 80.785 ;
      POLYGON  70.31 80.065 70.31 79.995 70.68 79.995 70.68 79.755 70.31 79.755 70.31 79.685 70.17 79.685 70.17 80.065 70.31 80.065 ;
      RECT  70.68 80.545 70.17 80.305 ;
      RECT  71.61 81.335 69.96 80.785 ;
      POLYGON  71.61 80.065 71.61 79.685 71.06 79.685 71.06 79.755 70.68 79.755 70.68 79.995 71.06 79.995 71.06 80.065 71.61 80.065 ;
      RECT  73.29 80.545 73.08 80.305 ;
      RECT  70.68 82.675 70.17 82.915 ;
      RECT  70.68 82.605 70.48 82.675 ;
      RECT  72.15 82.055 71.61 82.435 ;
      RECT  73.08 80.785 72.15 81.335 ;
      RECT  73.29 82.675 73.08 82.915 ;
      RECT  70.17 82.675 69.96 82.915 ;
      RECT  73.08 82.675 70.68 82.915 ;
      RECT  70.89 81.815 70.68 81.885 ;
      RECT  70.17 82.055 69.96 82.435 ;
      RECT  70.89 82.605 70.68 82.675 ;
      RECT  70.68 81.815 70.48 81.885 ;
      RECT  73.08 81.575 70.68 81.815 ;
      RECT  70.17 81.575 69.96 81.815 ;
      RECT  72.15 80.785 71.61 81.335 ;
      RECT  73.29 82.055 72.15 82.435 ;
      RECT  73.29 80.785 73.08 81.335 ;
      POLYGON  70.31 82.055 70.31 82.125 70.68 82.125 70.68 82.365 70.31 82.365 70.31 82.435 70.17 82.435 70.17 82.055 70.31 82.055 ;
      RECT  70.68 81.575 70.17 81.815 ;
      RECT  71.61 80.785 69.96 81.335 ;
      POLYGON  71.61 82.055 71.61 82.435 71.06 82.435 71.06 82.365 70.68 82.365 70.68 82.125 71.06 82.125 71.06 82.055 71.61 82.055 ;
      RECT  73.29 81.575 73.08 81.815 ;
      RECT  70.68 83.395 70.17 83.155 ;
      RECT  70.68 83.465 70.48 83.395 ;
      RECT  72.15 84.015 71.61 83.635 ;
      RECT  73.08 85.285 72.15 84.735 ;
      RECT  73.29 83.395 73.08 83.155 ;
      RECT  70.17 83.395 69.96 83.155 ;
      RECT  73.08 83.395 70.68 83.155 ;
      RECT  70.89 84.255 70.68 84.185 ;
      RECT  70.17 84.015 69.96 83.635 ;
      RECT  70.89 83.465 70.68 83.395 ;
      RECT  70.68 84.255 70.48 84.185 ;
      RECT  73.08 84.495 70.68 84.255 ;
      RECT  70.17 84.495 69.96 84.255 ;
      RECT  72.15 85.285 71.61 84.735 ;
      RECT  73.29 84.015 72.15 83.635 ;
      RECT  73.29 85.285 73.08 84.735 ;
      POLYGON  70.31 84.015 70.31 83.945 70.68 83.945 70.68 83.705 70.31 83.705 70.31 83.635 70.17 83.635 70.17 84.015 70.31 84.015 ;
      RECT  70.68 84.495 70.17 84.255 ;
      RECT  71.61 85.285 69.96 84.735 ;
      POLYGON  71.61 84.015 71.61 83.635 71.06 83.635 71.06 83.705 70.68 83.705 70.68 83.945 71.06 83.945 71.06 84.015 71.61 84.015 ;
      RECT  73.29 84.495 73.08 84.255 ;
      RECT  70.68 86.625 70.17 86.865 ;
      RECT  70.68 86.555 70.48 86.625 ;
      RECT  72.15 86.005 71.61 86.385 ;
      RECT  73.08 84.735 72.15 85.285 ;
      RECT  73.29 86.625 73.08 86.865 ;
      RECT  70.17 86.625 69.96 86.865 ;
      RECT  73.08 86.625 70.68 86.865 ;
      RECT  70.89 85.765 70.68 85.835 ;
      RECT  70.17 86.005 69.96 86.385 ;
      RECT  70.89 86.555 70.68 86.625 ;
      RECT  70.68 85.765 70.48 85.835 ;
      RECT  73.08 85.525 70.68 85.765 ;
      RECT  70.17 85.525 69.96 85.765 ;
      RECT  72.15 84.735 71.61 85.285 ;
      RECT  73.29 86.005 72.15 86.385 ;
      RECT  73.29 84.735 73.08 85.285 ;
      POLYGON  70.31 86.005 70.31 86.075 70.68 86.075 70.68 86.315 70.31 86.315 70.31 86.385 70.17 86.385 70.17 86.005 70.31 86.005 ;
      RECT  70.68 85.525 70.17 85.765 ;
      RECT  71.61 84.735 69.96 85.285 ;
      POLYGON  71.61 86.005 71.61 86.385 71.06 86.385 71.06 86.315 70.68 86.315 70.68 86.075 71.06 86.075 71.06 86.005 71.61 86.005 ;
      RECT  73.29 85.525 73.08 85.765 ;
      RECT  70.68 87.345 70.17 87.105 ;
      RECT  70.68 87.415 70.48 87.345 ;
      RECT  72.15 87.965 71.61 87.585 ;
      RECT  73.08 89.235 72.15 88.685 ;
      RECT  73.29 87.345 73.08 87.105 ;
      RECT  70.17 87.345 69.96 87.105 ;
      RECT  73.08 87.345 70.68 87.105 ;
      RECT  70.89 88.205 70.68 88.135 ;
      RECT  70.17 87.965 69.96 87.585 ;
      RECT  70.89 87.415 70.68 87.345 ;
      RECT  70.68 88.205 70.48 88.135 ;
      RECT  73.08 88.445 70.68 88.205 ;
      RECT  70.17 88.445 69.96 88.205 ;
      RECT  72.15 89.235 71.61 88.685 ;
      RECT  73.29 87.965 72.15 87.585 ;
      RECT  73.29 89.235 73.08 88.685 ;
      POLYGON  70.31 87.965 70.31 87.895 70.68 87.895 70.68 87.655 70.31 87.655 70.31 87.585 70.17 87.585 70.17 87.965 70.31 87.965 ;
      RECT  70.68 88.445 70.17 88.205 ;
      RECT  71.61 89.235 69.96 88.685 ;
      POLYGON  71.61 87.965 71.61 87.585 71.06 87.585 71.06 87.655 70.68 87.655 70.68 87.895 71.06 87.895 71.06 87.965 71.61 87.965 ;
      RECT  73.29 88.445 73.08 88.205 ;
      RECT  70.68 90.575 70.17 90.815 ;
      RECT  70.68 90.505 70.48 90.575 ;
      RECT  72.15 89.955 71.61 90.335 ;
      RECT  73.08 88.685 72.15 89.235 ;
      RECT  73.29 90.575 73.08 90.815 ;
      RECT  70.17 90.575 69.96 90.815 ;
      RECT  73.08 90.575 70.68 90.815 ;
      RECT  70.89 89.715 70.68 89.785 ;
      RECT  70.17 89.955 69.96 90.335 ;
      RECT  70.89 90.505 70.68 90.575 ;
      RECT  70.68 89.715 70.48 89.785 ;
      RECT  73.08 89.475 70.68 89.715 ;
      RECT  70.17 89.475 69.96 89.715 ;
      RECT  72.15 88.685 71.61 89.235 ;
      RECT  73.29 89.955 72.15 90.335 ;
      RECT  73.29 88.685 73.08 89.235 ;
      POLYGON  70.31 89.955 70.31 90.025 70.68 90.025 70.68 90.265 70.31 90.265 70.31 90.335 70.17 90.335 70.17 89.955 70.31 89.955 ;
      RECT  70.68 89.475 70.17 89.715 ;
      RECT  71.61 88.685 69.96 89.235 ;
      POLYGON  71.61 89.955 71.61 90.335 71.06 90.335 71.06 90.265 70.68 90.265 70.68 90.025 71.06 90.025 71.06 89.955 71.61 89.955 ;
      RECT  73.29 89.475 73.08 89.715 ;
      RECT  70.68 91.295 70.17 91.055 ;
      RECT  70.68 91.365 70.48 91.295 ;
      RECT  72.15 91.915 71.61 91.535 ;
      RECT  73.08 93.185 72.15 92.635 ;
      RECT  73.29 91.295 73.08 91.055 ;
      RECT  70.17 91.295 69.96 91.055 ;
      RECT  73.08 91.295 70.68 91.055 ;
      RECT  70.89 92.155 70.68 92.085 ;
      RECT  70.17 91.915 69.96 91.535 ;
      RECT  70.89 91.365 70.68 91.295 ;
      RECT  70.68 92.155 70.48 92.085 ;
      RECT  73.08 92.395 70.68 92.155 ;
      RECT  70.17 92.395 69.96 92.155 ;
      RECT  72.15 93.185 71.61 92.635 ;
      RECT  73.29 91.915 72.15 91.535 ;
      RECT  73.29 93.185 73.08 92.635 ;
      POLYGON  70.31 91.915 70.31 91.845 70.68 91.845 70.68 91.605 70.31 91.605 70.31 91.535 70.17 91.535 70.17 91.915 70.31 91.915 ;
      RECT  70.68 92.395 70.17 92.155 ;
      RECT  71.61 93.185 69.96 92.635 ;
      POLYGON  71.61 91.915 71.61 91.535 71.06 91.535 71.06 91.605 70.68 91.605 70.68 91.845 71.06 91.845 71.06 91.915 71.61 91.915 ;
      RECT  73.29 92.395 73.08 92.155 ;
      RECT  70.68 94.525 70.17 94.765 ;
      RECT  70.68 94.455 70.48 94.525 ;
      RECT  72.15 93.905 71.61 94.285 ;
      RECT  73.08 92.635 72.15 93.185 ;
      RECT  73.29 94.525 73.08 94.765 ;
      RECT  70.17 94.525 69.96 94.765 ;
      RECT  73.08 94.525 70.68 94.765 ;
      RECT  70.89 93.665 70.68 93.735 ;
      RECT  70.17 93.905 69.96 94.285 ;
      RECT  70.89 94.455 70.68 94.525 ;
      RECT  70.68 93.665 70.48 93.735 ;
      RECT  73.08 93.425 70.68 93.665 ;
      RECT  70.17 93.425 69.96 93.665 ;
      RECT  72.15 92.635 71.61 93.185 ;
      RECT  73.29 93.905 72.15 94.285 ;
      RECT  73.29 92.635 73.08 93.185 ;
      POLYGON  70.31 93.905 70.31 93.975 70.68 93.975 70.68 94.215 70.31 94.215 70.31 94.285 70.17 94.285 70.17 93.905 70.31 93.905 ;
      RECT  70.68 93.425 70.17 93.665 ;
      RECT  71.61 92.635 69.96 93.185 ;
      POLYGON  71.61 93.905 71.61 94.285 71.06 94.285 71.06 94.215 70.68 94.215 70.68 93.975 71.06 93.975 71.06 93.905 71.61 93.905 ;
      RECT  73.29 93.425 73.08 93.665 ;
      RECT  73.08 95.99 69.96 95.44 ;
      RECT  69.96 59.455 73.08 59.695 ;
      RECT  69.96 60.555 73.08 60.795 ;
      RECT  69.96 62.925 73.08 63.165 ;
      RECT  69.96 61.825 73.08 62.065 ;
      RECT  69.96 63.405 73.08 63.645 ;
      RECT  69.96 64.505 73.08 64.745 ;
      RECT  69.96 66.875 73.08 67.115 ;
      RECT  69.96 65.775 73.08 66.015 ;
      RECT  69.96 67.355 73.08 67.595 ;
      RECT  69.96 68.455 73.08 68.695 ;
      RECT  69.96 70.825 73.08 71.065 ;
      RECT  69.96 69.725 73.08 69.965 ;
      RECT  69.96 71.305 73.08 71.545 ;
      RECT  69.96 72.405 73.08 72.645 ;
      RECT  69.96 74.775 73.08 75.015 ;
      RECT  69.96 73.675 73.08 73.915 ;
      RECT  69.96 75.255 73.08 75.495 ;
      RECT  69.96 76.355 73.08 76.595 ;
      RECT  69.96 78.725 73.08 78.965 ;
      RECT  69.96 77.625 73.08 77.865 ;
      RECT  69.96 79.205 73.08 79.445 ;
      RECT  69.96 80.305 73.08 80.545 ;
      RECT  69.96 82.675 73.08 82.915 ;
      RECT  69.96 81.575 73.08 81.815 ;
      RECT  69.96 83.155 73.08 83.395 ;
      RECT  69.96 84.255 73.08 84.495 ;
      RECT  69.96 86.625 73.08 86.865 ;
      RECT  69.96 85.525 73.08 85.765 ;
      RECT  69.96 87.105 73.08 87.345 ;
      RECT  69.96 88.205 73.08 88.445 ;
      RECT  69.96 90.575 73.08 90.815 ;
      RECT  69.96 89.475 73.08 89.715 ;
      RECT  69.96 91.055 73.08 91.295 ;
      RECT  69.96 92.155 73.08 92.395 ;
      RECT  69.96 94.525 73.08 94.765 ;
      RECT  69.96 93.425 73.08 93.665 ;
      RECT  71.61 63.885 72.15 64.265 ;
      RECT  71.61 66.255 72.15 66.635 ;
      RECT  71.61 91.535 72.15 91.915 ;
      RECT  71.61 68.935 72.15 69.485 ;
      RECT  71.61 64.985 72.15 65.535 ;
      RECT  71.61 67.835 72.15 68.215 ;
      RECT  71.61 83.635 72.15 84.015 ;
      RECT  71.61 89.955 72.15 90.335 ;
      RECT  71.61 75.735 72.15 76.115 ;
      RECT  71.61 59.935 72.15 60.315 ;
      RECT  71.61 70.205 72.15 70.585 ;
      RECT  71.61 79.685 72.15 80.065 ;
      RECT  71.61 80.785 72.15 81.335 ;
      RECT  71.61 72.885 72.15 73.435 ;
      RECT  71.61 78.105 72.15 78.485 ;
      RECT  71.61 76.835 72.15 77.385 ;
      RECT  71.61 93.905 72.15 94.285 ;
      RECT  71.61 87.585 72.15 87.965 ;
      RECT  71.61 82.055 72.15 82.435 ;
      RECT  71.61 92.635 72.15 93.185 ;
      RECT  71.61 84.735 72.15 85.285 ;
      RECT  71.61 86.005 72.15 86.385 ;
      RECT  71.61 88.685 72.15 89.235 ;
      RECT  71.61 74.155 72.15 74.535 ;
      RECT  71.61 62.305 72.15 62.685 ;
      RECT  71.61 61.035 72.15 61.585 ;
      RECT  71.61 71.785 72.15 72.165 ;
      RECT  79.32 58.23 82.44 58.78 ;
      RECT  81.72 59.695 82.23 59.455 ;
      RECT  81.72 59.765 81.92 59.695 ;
      RECT  80.25 60.315 80.79 59.935 ;
      RECT  79.32 61.585 80.25 61.035 ;
      RECT  79.11 59.695 79.32 59.455 ;
      RECT  82.23 59.695 82.44 59.455 ;
      RECT  79.32 59.695 81.72 59.455 ;
      RECT  81.51 60.555 81.72 60.485 ;
      RECT  82.23 60.315 82.44 59.935 ;
      RECT  81.51 59.765 81.72 59.695 ;
      RECT  81.72 60.555 81.92 60.485 ;
      RECT  79.32 60.795 81.72 60.555 ;
      RECT  82.23 60.795 82.44 60.555 ;
      RECT  80.25 61.585 80.79 61.035 ;
      RECT  79.11 60.315 80.25 59.935 ;
      RECT  79.11 61.585 79.32 61.035 ;
      POLYGON  82.09 60.315 82.09 60.245 81.72 60.245 81.72 60.005 82.09 60.005 82.09 59.935 82.23 59.935 82.23 60.315 82.09 60.315 ;
      RECT  81.72 60.795 82.23 60.555 ;
      RECT  80.79 61.585 82.44 61.035 ;
      POLYGON  80.79 60.315 80.79 59.935 81.34 59.935 81.34 60.005 81.72 60.005 81.72 60.245 81.34 60.245 81.34 60.315 80.79 60.315 ;
      RECT  79.11 60.795 79.32 60.555 ;
      RECT  81.72 62.925 82.23 63.165 ;
      RECT  81.72 62.855 81.92 62.925 ;
      RECT  80.25 62.305 80.79 62.685 ;
      RECT  79.32 61.035 80.25 61.585 ;
      RECT  79.11 62.925 79.32 63.165 ;
      RECT  82.23 62.925 82.44 63.165 ;
      RECT  79.32 62.925 81.72 63.165 ;
      RECT  81.51 62.065 81.72 62.135 ;
      RECT  82.23 62.305 82.44 62.685 ;
      RECT  81.51 62.855 81.72 62.925 ;
      RECT  81.72 62.065 81.92 62.135 ;
      RECT  79.32 61.825 81.72 62.065 ;
      RECT  82.23 61.825 82.44 62.065 ;
      RECT  80.25 61.035 80.79 61.585 ;
      RECT  79.11 62.305 80.25 62.685 ;
      RECT  79.11 61.035 79.32 61.585 ;
      POLYGON  82.09 62.305 82.09 62.375 81.72 62.375 81.72 62.615 82.09 62.615 82.09 62.685 82.23 62.685 82.23 62.305 82.09 62.305 ;
      RECT  81.72 61.825 82.23 62.065 ;
      RECT  80.79 61.035 82.44 61.585 ;
      POLYGON  80.79 62.305 80.79 62.685 81.34 62.685 81.34 62.615 81.72 62.615 81.72 62.375 81.34 62.375 81.34 62.305 80.79 62.305 ;
      RECT  79.11 61.825 79.32 62.065 ;
      RECT  81.72 63.645 82.23 63.405 ;
      RECT  81.72 63.715 81.92 63.645 ;
      RECT  80.25 64.265 80.79 63.885 ;
      RECT  79.32 65.535 80.25 64.985 ;
      RECT  79.11 63.645 79.32 63.405 ;
      RECT  82.23 63.645 82.44 63.405 ;
      RECT  79.32 63.645 81.72 63.405 ;
      RECT  81.51 64.505 81.72 64.435 ;
      RECT  82.23 64.265 82.44 63.885 ;
      RECT  81.51 63.715 81.72 63.645 ;
      RECT  81.72 64.505 81.92 64.435 ;
      RECT  79.32 64.745 81.72 64.505 ;
      RECT  82.23 64.745 82.44 64.505 ;
      RECT  80.25 65.535 80.79 64.985 ;
      RECT  79.11 64.265 80.25 63.885 ;
      RECT  79.11 65.535 79.32 64.985 ;
      POLYGON  82.09 64.265 82.09 64.195 81.72 64.195 81.72 63.955 82.09 63.955 82.09 63.885 82.23 63.885 82.23 64.265 82.09 64.265 ;
      RECT  81.72 64.745 82.23 64.505 ;
      RECT  80.79 65.535 82.44 64.985 ;
      POLYGON  80.79 64.265 80.79 63.885 81.34 63.885 81.34 63.955 81.72 63.955 81.72 64.195 81.34 64.195 81.34 64.265 80.79 64.265 ;
      RECT  79.11 64.745 79.32 64.505 ;
      RECT  81.72 66.875 82.23 67.115 ;
      RECT  81.72 66.805 81.92 66.875 ;
      RECT  80.25 66.255 80.79 66.635 ;
      RECT  79.32 64.985 80.25 65.535 ;
      RECT  79.11 66.875 79.32 67.115 ;
      RECT  82.23 66.875 82.44 67.115 ;
      RECT  79.32 66.875 81.72 67.115 ;
      RECT  81.51 66.015 81.72 66.085 ;
      RECT  82.23 66.255 82.44 66.635 ;
      RECT  81.51 66.805 81.72 66.875 ;
      RECT  81.72 66.015 81.92 66.085 ;
      RECT  79.32 65.775 81.72 66.015 ;
      RECT  82.23 65.775 82.44 66.015 ;
      RECT  80.25 64.985 80.79 65.535 ;
      RECT  79.11 66.255 80.25 66.635 ;
      RECT  79.11 64.985 79.32 65.535 ;
      POLYGON  82.09 66.255 82.09 66.325 81.72 66.325 81.72 66.565 82.09 66.565 82.09 66.635 82.23 66.635 82.23 66.255 82.09 66.255 ;
      RECT  81.72 65.775 82.23 66.015 ;
      RECT  80.79 64.985 82.44 65.535 ;
      POLYGON  80.79 66.255 80.79 66.635 81.34 66.635 81.34 66.565 81.72 66.565 81.72 66.325 81.34 66.325 81.34 66.255 80.79 66.255 ;
      RECT  79.11 65.775 79.32 66.015 ;
      RECT  81.72 67.595 82.23 67.355 ;
      RECT  81.72 67.665 81.92 67.595 ;
      RECT  80.25 68.215 80.79 67.835 ;
      RECT  79.32 69.485 80.25 68.935 ;
      RECT  79.11 67.595 79.32 67.355 ;
      RECT  82.23 67.595 82.44 67.355 ;
      RECT  79.32 67.595 81.72 67.355 ;
      RECT  81.51 68.455 81.72 68.385 ;
      RECT  82.23 68.215 82.44 67.835 ;
      RECT  81.51 67.665 81.72 67.595 ;
      RECT  81.72 68.455 81.92 68.385 ;
      RECT  79.32 68.695 81.72 68.455 ;
      RECT  82.23 68.695 82.44 68.455 ;
      RECT  80.25 69.485 80.79 68.935 ;
      RECT  79.11 68.215 80.25 67.835 ;
      RECT  79.11 69.485 79.32 68.935 ;
      POLYGON  82.09 68.215 82.09 68.145 81.72 68.145 81.72 67.905 82.09 67.905 82.09 67.835 82.23 67.835 82.23 68.215 82.09 68.215 ;
      RECT  81.72 68.695 82.23 68.455 ;
      RECT  80.79 69.485 82.44 68.935 ;
      POLYGON  80.79 68.215 80.79 67.835 81.34 67.835 81.34 67.905 81.72 67.905 81.72 68.145 81.34 68.145 81.34 68.215 80.79 68.215 ;
      RECT  79.11 68.695 79.32 68.455 ;
      RECT  81.72 70.825 82.23 71.065 ;
      RECT  81.72 70.755 81.92 70.825 ;
      RECT  80.25 70.205 80.79 70.585 ;
      RECT  79.32 68.935 80.25 69.485 ;
      RECT  79.11 70.825 79.32 71.065 ;
      RECT  82.23 70.825 82.44 71.065 ;
      RECT  79.32 70.825 81.72 71.065 ;
      RECT  81.51 69.965 81.72 70.035 ;
      RECT  82.23 70.205 82.44 70.585 ;
      RECT  81.51 70.755 81.72 70.825 ;
      RECT  81.72 69.965 81.92 70.035 ;
      RECT  79.32 69.725 81.72 69.965 ;
      RECT  82.23 69.725 82.44 69.965 ;
      RECT  80.25 68.935 80.79 69.485 ;
      RECT  79.11 70.205 80.25 70.585 ;
      RECT  79.11 68.935 79.32 69.485 ;
      POLYGON  82.09 70.205 82.09 70.275 81.72 70.275 81.72 70.515 82.09 70.515 82.09 70.585 82.23 70.585 82.23 70.205 82.09 70.205 ;
      RECT  81.72 69.725 82.23 69.965 ;
      RECT  80.79 68.935 82.44 69.485 ;
      POLYGON  80.79 70.205 80.79 70.585 81.34 70.585 81.34 70.515 81.72 70.515 81.72 70.275 81.34 70.275 81.34 70.205 80.79 70.205 ;
      RECT  79.11 69.725 79.32 69.965 ;
      RECT  81.72 71.545 82.23 71.305 ;
      RECT  81.72 71.615 81.92 71.545 ;
      RECT  80.25 72.165 80.79 71.785 ;
      RECT  79.32 73.435 80.25 72.885 ;
      RECT  79.11 71.545 79.32 71.305 ;
      RECT  82.23 71.545 82.44 71.305 ;
      RECT  79.32 71.545 81.72 71.305 ;
      RECT  81.51 72.405 81.72 72.335 ;
      RECT  82.23 72.165 82.44 71.785 ;
      RECT  81.51 71.615 81.72 71.545 ;
      RECT  81.72 72.405 81.92 72.335 ;
      RECT  79.32 72.645 81.72 72.405 ;
      RECT  82.23 72.645 82.44 72.405 ;
      RECT  80.25 73.435 80.79 72.885 ;
      RECT  79.11 72.165 80.25 71.785 ;
      RECT  79.11 73.435 79.32 72.885 ;
      POLYGON  82.09 72.165 82.09 72.095 81.72 72.095 81.72 71.855 82.09 71.855 82.09 71.785 82.23 71.785 82.23 72.165 82.09 72.165 ;
      RECT  81.72 72.645 82.23 72.405 ;
      RECT  80.79 73.435 82.44 72.885 ;
      POLYGON  80.79 72.165 80.79 71.785 81.34 71.785 81.34 71.855 81.72 71.855 81.72 72.095 81.34 72.095 81.34 72.165 80.79 72.165 ;
      RECT  79.11 72.645 79.32 72.405 ;
      RECT  81.72 74.775 82.23 75.015 ;
      RECT  81.72 74.705 81.92 74.775 ;
      RECT  80.25 74.155 80.79 74.535 ;
      RECT  79.32 72.885 80.25 73.435 ;
      RECT  79.11 74.775 79.32 75.015 ;
      RECT  82.23 74.775 82.44 75.015 ;
      RECT  79.32 74.775 81.72 75.015 ;
      RECT  81.51 73.915 81.72 73.985 ;
      RECT  82.23 74.155 82.44 74.535 ;
      RECT  81.51 74.705 81.72 74.775 ;
      RECT  81.72 73.915 81.92 73.985 ;
      RECT  79.32 73.675 81.72 73.915 ;
      RECT  82.23 73.675 82.44 73.915 ;
      RECT  80.25 72.885 80.79 73.435 ;
      RECT  79.11 74.155 80.25 74.535 ;
      RECT  79.11 72.885 79.32 73.435 ;
      POLYGON  82.09 74.155 82.09 74.225 81.72 74.225 81.72 74.465 82.09 74.465 82.09 74.535 82.23 74.535 82.23 74.155 82.09 74.155 ;
      RECT  81.72 73.675 82.23 73.915 ;
      RECT  80.79 72.885 82.44 73.435 ;
      POLYGON  80.79 74.155 80.79 74.535 81.34 74.535 81.34 74.465 81.72 74.465 81.72 74.225 81.34 74.225 81.34 74.155 80.79 74.155 ;
      RECT  79.11 73.675 79.32 73.915 ;
      RECT  81.72 75.495 82.23 75.255 ;
      RECT  81.72 75.565 81.92 75.495 ;
      RECT  80.25 76.115 80.79 75.735 ;
      RECT  79.32 77.385 80.25 76.835 ;
      RECT  79.11 75.495 79.32 75.255 ;
      RECT  82.23 75.495 82.44 75.255 ;
      RECT  79.32 75.495 81.72 75.255 ;
      RECT  81.51 76.355 81.72 76.285 ;
      RECT  82.23 76.115 82.44 75.735 ;
      RECT  81.51 75.565 81.72 75.495 ;
      RECT  81.72 76.355 81.92 76.285 ;
      RECT  79.32 76.595 81.72 76.355 ;
      RECT  82.23 76.595 82.44 76.355 ;
      RECT  80.25 77.385 80.79 76.835 ;
      RECT  79.11 76.115 80.25 75.735 ;
      RECT  79.11 77.385 79.32 76.835 ;
      POLYGON  82.09 76.115 82.09 76.045 81.72 76.045 81.72 75.805 82.09 75.805 82.09 75.735 82.23 75.735 82.23 76.115 82.09 76.115 ;
      RECT  81.72 76.595 82.23 76.355 ;
      RECT  80.79 77.385 82.44 76.835 ;
      POLYGON  80.79 76.115 80.79 75.735 81.34 75.735 81.34 75.805 81.72 75.805 81.72 76.045 81.34 76.045 81.34 76.115 80.79 76.115 ;
      RECT  79.11 76.595 79.32 76.355 ;
      RECT  81.72 78.725 82.23 78.965 ;
      RECT  81.72 78.655 81.92 78.725 ;
      RECT  80.25 78.105 80.79 78.485 ;
      RECT  79.32 76.835 80.25 77.385 ;
      RECT  79.11 78.725 79.32 78.965 ;
      RECT  82.23 78.725 82.44 78.965 ;
      RECT  79.32 78.725 81.72 78.965 ;
      RECT  81.51 77.865 81.72 77.935 ;
      RECT  82.23 78.105 82.44 78.485 ;
      RECT  81.51 78.655 81.72 78.725 ;
      RECT  81.72 77.865 81.92 77.935 ;
      RECT  79.32 77.625 81.72 77.865 ;
      RECT  82.23 77.625 82.44 77.865 ;
      RECT  80.25 76.835 80.79 77.385 ;
      RECT  79.11 78.105 80.25 78.485 ;
      RECT  79.11 76.835 79.32 77.385 ;
      POLYGON  82.09 78.105 82.09 78.175 81.72 78.175 81.72 78.415 82.09 78.415 82.09 78.485 82.23 78.485 82.23 78.105 82.09 78.105 ;
      RECT  81.72 77.625 82.23 77.865 ;
      RECT  80.79 76.835 82.44 77.385 ;
      POLYGON  80.79 78.105 80.79 78.485 81.34 78.485 81.34 78.415 81.72 78.415 81.72 78.175 81.34 78.175 81.34 78.105 80.79 78.105 ;
      RECT  79.11 77.625 79.32 77.865 ;
      RECT  81.72 79.445 82.23 79.205 ;
      RECT  81.72 79.515 81.92 79.445 ;
      RECT  80.25 80.065 80.79 79.685 ;
      RECT  79.32 81.335 80.25 80.785 ;
      RECT  79.11 79.445 79.32 79.205 ;
      RECT  82.23 79.445 82.44 79.205 ;
      RECT  79.32 79.445 81.72 79.205 ;
      RECT  81.51 80.305 81.72 80.235 ;
      RECT  82.23 80.065 82.44 79.685 ;
      RECT  81.51 79.515 81.72 79.445 ;
      RECT  81.72 80.305 81.92 80.235 ;
      RECT  79.32 80.545 81.72 80.305 ;
      RECT  82.23 80.545 82.44 80.305 ;
      RECT  80.25 81.335 80.79 80.785 ;
      RECT  79.11 80.065 80.25 79.685 ;
      RECT  79.11 81.335 79.32 80.785 ;
      POLYGON  82.09 80.065 82.09 79.995 81.72 79.995 81.72 79.755 82.09 79.755 82.09 79.685 82.23 79.685 82.23 80.065 82.09 80.065 ;
      RECT  81.72 80.545 82.23 80.305 ;
      RECT  80.79 81.335 82.44 80.785 ;
      POLYGON  80.79 80.065 80.79 79.685 81.34 79.685 81.34 79.755 81.72 79.755 81.72 79.995 81.34 79.995 81.34 80.065 80.79 80.065 ;
      RECT  79.11 80.545 79.32 80.305 ;
      RECT  81.72 82.675 82.23 82.915 ;
      RECT  81.72 82.605 81.92 82.675 ;
      RECT  80.25 82.055 80.79 82.435 ;
      RECT  79.32 80.785 80.25 81.335 ;
      RECT  79.11 82.675 79.32 82.915 ;
      RECT  82.23 82.675 82.44 82.915 ;
      RECT  79.32 82.675 81.72 82.915 ;
      RECT  81.51 81.815 81.72 81.885 ;
      RECT  82.23 82.055 82.44 82.435 ;
      RECT  81.51 82.605 81.72 82.675 ;
      RECT  81.72 81.815 81.92 81.885 ;
      RECT  79.32 81.575 81.72 81.815 ;
      RECT  82.23 81.575 82.44 81.815 ;
      RECT  80.25 80.785 80.79 81.335 ;
      RECT  79.11 82.055 80.25 82.435 ;
      RECT  79.11 80.785 79.32 81.335 ;
      POLYGON  82.09 82.055 82.09 82.125 81.72 82.125 81.72 82.365 82.09 82.365 82.09 82.435 82.23 82.435 82.23 82.055 82.09 82.055 ;
      RECT  81.72 81.575 82.23 81.815 ;
      RECT  80.79 80.785 82.44 81.335 ;
      POLYGON  80.79 82.055 80.79 82.435 81.34 82.435 81.34 82.365 81.72 82.365 81.72 82.125 81.34 82.125 81.34 82.055 80.79 82.055 ;
      RECT  79.11 81.575 79.32 81.815 ;
      RECT  81.72 83.395 82.23 83.155 ;
      RECT  81.72 83.465 81.92 83.395 ;
      RECT  80.25 84.015 80.79 83.635 ;
      RECT  79.32 85.285 80.25 84.735 ;
      RECT  79.11 83.395 79.32 83.155 ;
      RECT  82.23 83.395 82.44 83.155 ;
      RECT  79.32 83.395 81.72 83.155 ;
      RECT  81.51 84.255 81.72 84.185 ;
      RECT  82.23 84.015 82.44 83.635 ;
      RECT  81.51 83.465 81.72 83.395 ;
      RECT  81.72 84.255 81.92 84.185 ;
      RECT  79.32 84.495 81.72 84.255 ;
      RECT  82.23 84.495 82.44 84.255 ;
      RECT  80.25 85.285 80.79 84.735 ;
      RECT  79.11 84.015 80.25 83.635 ;
      RECT  79.11 85.285 79.32 84.735 ;
      POLYGON  82.09 84.015 82.09 83.945 81.72 83.945 81.72 83.705 82.09 83.705 82.09 83.635 82.23 83.635 82.23 84.015 82.09 84.015 ;
      RECT  81.72 84.495 82.23 84.255 ;
      RECT  80.79 85.285 82.44 84.735 ;
      POLYGON  80.79 84.015 80.79 83.635 81.34 83.635 81.34 83.705 81.72 83.705 81.72 83.945 81.34 83.945 81.34 84.015 80.79 84.015 ;
      RECT  79.11 84.495 79.32 84.255 ;
      RECT  81.72 86.625 82.23 86.865 ;
      RECT  81.72 86.555 81.92 86.625 ;
      RECT  80.25 86.005 80.79 86.385 ;
      RECT  79.32 84.735 80.25 85.285 ;
      RECT  79.11 86.625 79.32 86.865 ;
      RECT  82.23 86.625 82.44 86.865 ;
      RECT  79.32 86.625 81.72 86.865 ;
      RECT  81.51 85.765 81.72 85.835 ;
      RECT  82.23 86.005 82.44 86.385 ;
      RECT  81.51 86.555 81.72 86.625 ;
      RECT  81.72 85.765 81.92 85.835 ;
      RECT  79.32 85.525 81.72 85.765 ;
      RECT  82.23 85.525 82.44 85.765 ;
      RECT  80.25 84.735 80.79 85.285 ;
      RECT  79.11 86.005 80.25 86.385 ;
      RECT  79.11 84.735 79.32 85.285 ;
      POLYGON  82.09 86.005 82.09 86.075 81.72 86.075 81.72 86.315 82.09 86.315 82.09 86.385 82.23 86.385 82.23 86.005 82.09 86.005 ;
      RECT  81.72 85.525 82.23 85.765 ;
      RECT  80.79 84.735 82.44 85.285 ;
      POLYGON  80.79 86.005 80.79 86.385 81.34 86.385 81.34 86.315 81.72 86.315 81.72 86.075 81.34 86.075 81.34 86.005 80.79 86.005 ;
      RECT  79.11 85.525 79.32 85.765 ;
      RECT  81.72 87.345 82.23 87.105 ;
      RECT  81.72 87.415 81.92 87.345 ;
      RECT  80.25 87.965 80.79 87.585 ;
      RECT  79.32 89.235 80.25 88.685 ;
      RECT  79.11 87.345 79.32 87.105 ;
      RECT  82.23 87.345 82.44 87.105 ;
      RECT  79.32 87.345 81.72 87.105 ;
      RECT  81.51 88.205 81.72 88.135 ;
      RECT  82.23 87.965 82.44 87.585 ;
      RECT  81.51 87.415 81.72 87.345 ;
      RECT  81.72 88.205 81.92 88.135 ;
      RECT  79.32 88.445 81.72 88.205 ;
      RECT  82.23 88.445 82.44 88.205 ;
      RECT  80.25 89.235 80.79 88.685 ;
      RECT  79.11 87.965 80.25 87.585 ;
      RECT  79.11 89.235 79.32 88.685 ;
      POLYGON  82.09 87.965 82.09 87.895 81.72 87.895 81.72 87.655 82.09 87.655 82.09 87.585 82.23 87.585 82.23 87.965 82.09 87.965 ;
      RECT  81.72 88.445 82.23 88.205 ;
      RECT  80.79 89.235 82.44 88.685 ;
      POLYGON  80.79 87.965 80.79 87.585 81.34 87.585 81.34 87.655 81.72 87.655 81.72 87.895 81.34 87.895 81.34 87.965 80.79 87.965 ;
      RECT  79.11 88.445 79.32 88.205 ;
      RECT  81.72 90.575 82.23 90.815 ;
      RECT  81.72 90.505 81.92 90.575 ;
      RECT  80.25 89.955 80.79 90.335 ;
      RECT  79.32 88.685 80.25 89.235 ;
      RECT  79.11 90.575 79.32 90.815 ;
      RECT  82.23 90.575 82.44 90.815 ;
      RECT  79.32 90.575 81.72 90.815 ;
      RECT  81.51 89.715 81.72 89.785 ;
      RECT  82.23 89.955 82.44 90.335 ;
      RECT  81.51 90.505 81.72 90.575 ;
      RECT  81.72 89.715 81.92 89.785 ;
      RECT  79.32 89.475 81.72 89.715 ;
      RECT  82.23 89.475 82.44 89.715 ;
      RECT  80.25 88.685 80.79 89.235 ;
      RECT  79.11 89.955 80.25 90.335 ;
      RECT  79.11 88.685 79.32 89.235 ;
      POLYGON  82.09 89.955 82.09 90.025 81.72 90.025 81.72 90.265 82.09 90.265 82.09 90.335 82.23 90.335 82.23 89.955 82.09 89.955 ;
      RECT  81.72 89.475 82.23 89.715 ;
      RECT  80.79 88.685 82.44 89.235 ;
      POLYGON  80.79 89.955 80.79 90.335 81.34 90.335 81.34 90.265 81.72 90.265 81.72 90.025 81.34 90.025 81.34 89.955 80.79 89.955 ;
      RECT  79.11 89.475 79.32 89.715 ;
      RECT  81.72 91.295 82.23 91.055 ;
      RECT  81.72 91.365 81.92 91.295 ;
      RECT  80.25 91.915 80.79 91.535 ;
      RECT  79.32 93.185 80.25 92.635 ;
      RECT  79.11 91.295 79.32 91.055 ;
      RECT  82.23 91.295 82.44 91.055 ;
      RECT  79.32 91.295 81.72 91.055 ;
      RECT  81.51 92.155 81.72 92.085 ;
      RECT  82.23 91.915 82.44 91.535 ;
      RECT  81.51 91.365 81.72 91.295 ;
      RECT  81.72 92.155 81.92 92.085 ;
      RECT  79.32 92.395 81.72 92.155 ;
      RECT  82.23 92.395 82.44 92.155 ;
      RECT  80.25 93.185 80.79 92.635 ;
      RECT  79.11 91.915 80.25 91.535 ;
      RECT  79.11 93.185 79.32 92.635 ;
      POLYGON  82.09 91.915 82.09 91.845 81.72 91.845 81.72 91.605 82.09 91.605 82.09 91.535 82.23 91.535 82.23 91.915 82.09 91.915 ;
      RECT  81.72 92.395 82.23 92.155 ;
      RECT  80.79 93.185 82.44 92.635 ;
      POLYGON  80.79 91.915 80.79 91.535 81.34 91.535 81.34 91.605 81.72 91.605 81.72 91.845 81.34 91.845 81.34 91.915 80.79 91.915 ;
      RECT  79.11 92.395 79.32 92.155 ;
      RECT  81.72 94.525 82.23 94.765 ;
      RECT  81.72 94.455 81.92 94.525 ;
      RECT  80.25 93.905 80.79 94.285 ;
      RECT  79.32 92.635 80.25 93.185 ;
      RECT  79.11 94.525 79.32 94.765 ;
      RECT  82.23 94.525 82.44 94.765 ;
      RECT  79.32 94.525 81.72 94.765 ;
      RECT  81.51 93.665 81.72 93.735 ;
      RECT  82.23 93.905 82.44 94.285 ;
      RECT  81.51 94.455 81.72 94.525 ;
      RECT  81.72 93.665 81.92 93.735 ;
      RECT  79.32 93.425 81.72 93.665 ;
      RECT  82.23 93.425 82.44 93.665 ;
      RECT  80.25 92.635 80.79 93.185 ;
      RECT  79.11 93.905 80.25 94.285 ;
      RECT  79.11 92.635 79.32 93.185 ;
      POLYGON  82.09 93.905 82.09 93.975 81.72 93.975 81.72 94.215 82.09 94.215 82.09 94.285 82.23 94.285 82.23 93.905 82.09 93.905 ;
      RECT  81.72 93.425 82.23 93.665 ;
      RECT  80.79 92.635 82.44 93.185 ;
      POLYGON  80.79 93.905 80.79 94.285 81.34 94.285 81.34 94.215 81.72 94.215 81.72 93.975 81.34 93.975 81.34 93.905 80.79 93.905 ;
      RECT  79.11 93.425 79.32 93.665 ;
      RECT  79.32 95.99 82.44 95.44 ;
      RECT  79.32 59.455 82.44 59.695 ;
      RECT  79.32 60.555 82.44 60.795 ;
      RECT  79.32 62.925 82.44 63.165 ;
      RECT  79.32 61.825 82.44 62.065 ;
      RECT  79.32 63.405 82.44 63.645 ;
      RECT  79.32 64.505 82.44 64.745 ;
      RECT  79.32 66.875 82.44 67.115 ;
      RECT  79.32 65.775 82.44 66.015 ;
      RECT  79.32 67.355 82.44 67.595 ;
      RECT  79.32 68.455 82.44 68.695 ;
      RECT  79.32 70.825 82.44 71.065 ;
      RECT  79.32 69.725 82.44 69.965 ;
      RECT  79.32 71.305 82.44 71.545 ;
      RECT  79.32 72.405 82.44 72.645 ;
      RECT  79.32 74.775 82.44 75.015 ;
      RECT  79.32 73.675 82.44 73.915 ;
      RECT  79.32 75.255 82.44 75.495 ;
      RECT  79.32 76.355 82.44 76.595 ;
      RECT  79.32 78.725 82.44 78.965 ;
      RECT  79.32 77.625 82.44 77.865 ;
      RECT  79.32 79.205 82.44 79.445 ;
      RECT  79.32 80.305 82.44 80.545 ;
      RECT  79.32 82.675 82.44 82.915 ;
      RECT  79.32 81.575 82.44 81.815 ;
      RECT  79.32 83.155 82.44 83.395 ;
      RECT  79.32 84.255 82.44 84.495 ;
      RECT  79.32 86.625 82.44 86.865 ;
      RECT  79.32 85.525 82.44 85.765 ;
      RECT  79.32 87.105 82.44 87.345 ;
      RECT  79.32 88.205 82.44 88.445 ;
      RECT  79.32 90.575 82.44 90.815 ;
      RECT  79.32 89.475 82.44 89.715 ;
      RECT  79.32 91.055 82.44 91.295 ;
      RECT  79.32 92.155 82.44 92.395 ;
      RECT  79.32 94.525 82.44 94.765 ;
      RECT  79.32 93.425 82.44 93.665 ;
      RECT  80.25 74.155 80.79 74.535 ;
      RECT  80.25 86.005 80.79 86.385 ;
      RECT  80.25 63.885 80.79 64.265 ;
      RECT  80.25 83.635 80.79 84.015 ;
      RECT  80.25 91.535 80.79 91.915 ;
      RECT  80.25 82.055 80.79 82.435 ;
      RECT  80.25 68.935 80.79 69.485 ;
      RECT  80.25 62.305 80.79 62.685 ;
      RECT  80.25 76.835 80.79 77.385 ;
      RECT  80.25 87.585 80.79 87.965 ;
      RECT  80.25 79.685 80.79 80.065 ;
      RECT  80.25 75.735 80.79 76.115 ;
      RECT  80.25 71.785 80.79 72.165 ;
      RECT  80.25 78.105 80.79 78.485 ;
      RECT  80.25 93.905 80.79 94.285 ;
      RECT  80.25 80.785 80.79 81.335 ;
      RECT  80.25 61.035 80.79 61.585 ;
      RECT  80.25 88.685 80.79 89.235 ;
      RECT  80.25 70.205 80.79 70.585 ;
      RECT  80.25 67.835 80.79 68.215 ;
      RECT  80.25 59.935 80.79 60.315 ;
      RECT  80.25 92.635 80.79 93.185 ;
      RECT  80.25 64.985 80.79 65.535 ;
      RECT  80.25 72.885 80.79 73.435 ;
      RECT  80.25 89.955 80.79 90.335 ;
      RECT  80.25 84.735 80.79 85.285 ;
      RECT  80.25 66.255 80.79 66.635 ;
      RECT  75.48 59.695 75.99 59.455 ;
      RECT  75.48 59.765 75.68 59.695 ;
      RECT  74.01 60.315 74.55 59.935 ;
      RECT  73.08 61.585 74.01 61.035 ;
      RECT  72.87 59.695 73.08 59.455 ;
      RECT  75.99 59.695 76.2 59.455 ;
      RECT  73.08 59.695 75.48 59.455 ;
      RECT  75.27 60.555 75.48 60.485 ;
      RECT  75.99 60.315 76.2 59.935 ;
      RECT  75.27 59.765 75.48 59.695 ;
      RECT  75.48 60.555 75.68 60.485 ;
      RECT  73.08 60.795 75.48 60.555 ;
      RECT  75.99 60.795 76.2 60.555 ;
      RECT  74.01 61.585 74.55 61.035 ;
      RECT  72.87 60.315 74.01 59.935 ;
      RECT  72.87 61.585 73.08 61.035 ;
      POLYGON  75.85 60.315 75.85 60.245 75.48 60.245 75.48 60.005 75.85 60.005 75.85 59.935 75.99 59.935 75.99 60.315 75.85 60.315 ;
      RECT  75.48 60.795 75.99 60.555 ;
      RECT  74.55 61.585 76.2 61.035 ;
      POLYGON  74.55 60.315 74.55 59.935 75.1 59.935 75.1 60.005 75.48 60.005 75.48 60.245 75.1 60.245 75.1 60.315 74.55 60.315 ;
      RECT  72.87 60.795 73.08 60.555 ;
      RECT  76.92 59.695 76.41 59.455 ;
      RECT  76.92 59.765 76.72 59.695 ;
      RECT  78.39 60.315 77.85 59.935 ;
      RECT  79.32 61.585 78.39 61.035 ;
      RECT  79.53 59.695 79.32 59.455 ;
      RECT  76.41 59.695 76.2 59.455 ;
      RECT  79.32 59.695 76.92 59.455 ;
      RECT  77.13 60.555 76.92 60.485 ;
      RECT  76.41 60.315 76.2 59.935 ;
      RECT  77.13 59.765 76.92 59.695 ;
      RECT  76.92 60.555 76.72 60.485 ;
      RECT  79.32 60.795 76.92 60.555 ;
      RECT  76.41 60.795 76.2 60.555 ;
      RECT  78.39 61.585 77.85 61.035 ;
      RECT  79.53 60.315 78.39 59.935 ;
      RECT  79.53 61.585 79.32 61.035 ;
      POLYGON  76.55 60.315 76.55 60.245 76.92 60.245 76.92 60.005 76.55 60.005 76.55 59.935 76.41 59.935 76.41 60.315 76.55 60.315 ;
      RECT  76.92 60.795 76.41 60.555 ;
      RECT  77.85 61.585 76.2 61.035 ;
      POLYGON  77.85 60.315 77.85 59.935 77.3 59.935 77.3 60.005 76.92 60.005 76.92 60.245 77.3 60.245 77.3 60.315 77.85 60.315 ;
      RECT  79.53 60.795 79.32 60.555 ;
      RECT  73.08 59.695 79.32 59.455 ;
      RECT  73.08 60.795 79.32 60.555 ;
      RECT  77.85 61.585 78.39 61.035 ;
      RECT  74.01 60.315 74.55 59.935 ;
      RECT  74.01 61.585 74.55 61.035 ;
      RECT  77.85 60.315 78.39 59.935 ;
      RECT  75.48 94.525 75.99 94.765 ;
      RECT  75.48 94.455 75.68 94.525 ;
      RECT  74.01 93.905 74.55 94.285 ;
      RECT  73.08 92.635 74.01 93.185 ;
      RECT  72.87 94.525 73.08 94.765 ;
      RECT  75.99 94.525 76.2 94.765 ;
      RECT  73.08 94.525 75.48 94.765 ;
      RECT  75.27 93.665 75.48 93.735 ;
      RECT  75.99 93.905 76.2 94.285 ;
      RECT  75.27 94.455 75.48 94.525 ;
      RECT  75.48 93.665 75.68 93.735 ;
      RECT  73.08 93.425 75.48 93.665 ;
      RECT  75.99 93.425 76.2 93.665 ;
      RECT  74.01 92.635 74.55 93.185 ;
      RECT  72.87 93.905 74.01 94.285 ;
      RECT  72.87 92.635 73.08 93.185 ;
      POLYGON  75.85 93.905 75.85 93.975 75.48 93.975 75.48 94.215 75.85 94.215 75.85 94.285 75.99 94.285 75.99 93.905 75.85 93.905 ;
      RECT  75.48 93.425 75.99 93.665 ;
      RECT  74.55 92.635 76.2 93.185 ;
      POLYGON  74.55 93.905 74.55 94.285 75.1 94.285 75.1 94.215 75.48 94.215 75.48 93.975 75.1 93.975 75.1 93.905 74.55 93.905 ;
      RECT  72.87 93.425 73.08 93.665 ;
      RECT  76.92 94.525 76.41 94.765 ;
      RECT  76.92 94.455 76.72 94.525 ;
      RECT  78.39 93.905 77.85 94.285 ;
      RECT  79.32 92.635 78.39 93.185 ;
      RECT  79.53 94.525 79.32 94.765 ;
      RECT  76.41 94.525 76.2 94.765 ;
      RECT  79.32 94.525 76.92 94.765 ;
      RECT  77.13 93.665 76.92 93.735 ;
      RECT  76.41 93.905 76.2 94.285 ;
      RECT  77.13 94.455 76.92 94.525 ;
      RECT  76.92 93.665 76.72 93.735 ;
      RECT  79.32 93.425 76.92 93.665 ;
      RECT  76.41 93.425 76.2 93.665 ;
      RECT  78.39 92.635 77.85 93.185 ;
      RECT  79.53 93.905 78.39 94.285 ;
      RECT  79.53 92.635 79.32 93.185 ;
      POLYGON  76.55 93.905 76.55 93.975 76.92 93.975 76.92 94.215 76.55 94.215 76.55 94.285 76.41 94.285 76.41 93.905 76.55 93.905 ;
      RECT  76.92 93.425 76.41 93.665 ;
      RECT  77.85 92.635 76.2 93.185 ;
      POLYGON  77.85 93.905 77.85 94.285 77.3 94.285 77.3 94.215 76.92 94.215 76.92 93.975 77.3 93.975 77.3 93.905 77.85 93.905 ;
      RECT  79.53 93.425 79.32 93.665 ;
      RECT  73.08 94.525 79.32 94.765 ;
      RECT  73.08 93.425 79.32 93.665 ;
      RECT  77.85 92.635 78.39 93.185 ;
      RECT  74.01 93.905 74.55 94.285 ;
      RECT  74.01 92.635 74.55 93.185 ;
      RECT  77.85 93.905 78.39 94.285 ;
      RECT  73.08 58.23 76.2 58.78 ;
      RECT  79.32 58.23 76.2 58.78 ;
      RECT  73.08 95.99 76.2 95.44 ;
      RECT  79.32 95.99 76.2 95.44 ;
      RECT  69.24 59.695 69.75 59.455 ;
      RECT  69.24 59.765 69.44 59.695 ;
      RECT  67.77 60.315 68.31 59.935 ;
      RECT  66.84 61.585 67.77 61.035 ;
      RECT  66.63 59.695 66.84 59.455 ;
      RECT  69.75 59.695 69.96 59.455 ;
      RECT  66.84 59.695 69.24 59.455 ;
      RECT  69.03 60.555 69.24 60.485 ;
      RECT  69.75 60.315 69.96 59.935 ;
      RECT  69.03 59.765 69.24 59.695 ;
      RECT  69.24 60.555 69.44 60.485 ;
      RECT  66.84 60.795 69.24 60.555 ;
      RECT  69.75 60.795 69.96 60.555 ;
      RECT  67.77 61.585 68.31 61.035 ;
      RECT  66.63 60.315 67.77 59.935 ;
      RECT  66.63 61.585 66.84 61.035 ;
      POLYGON  69.61 60.315 69.61 60.245 69.24 60.245 69.24 60.005 69.61 60.005 69.61 59.935 69.75 59.935 69.75 60.315 69.61 60.315 ;
      RECT  69.24 60.795 69.75 60.555 ;
      RECT  68.31 61.585 69.96 61.035 ;
      POLYGON  68.31 60.315 68.31 59.935 68.86 59.935 68.86 60.005 69.24 60.005 69.24 60.245 68.86 60.245 68.86 60.315 68.31 60.315 ;
      RECT  66.63 60.795 66.84 60.555 ;
      RECT  69.24 62.925 69.75 63.165 ;
      RECT  69.24 62.855 69.44 62.925 ;
      RECT  67.77 62.305 68.31 62.685 ;
      RECT  66.84 61.035 67.77 61.585 ;
      RECT  66.63 62.925 66.84 63.165 ;
      RECT  69.75 62.925 69.96 63.165 ;
      RECT  66.84 62.925 69.24 63.165 ;
      RECT  69.03 62.065 69.24 62.135 ;
      RECT  69.75 62.305 69.96 62.685 ;
      RECT  69.03 62.855 69.24 62.925 ;
      RECT  69.24 62.065 69.44 62.135 ;
      RECT  66.84 61.825 69.24 62.065 ;
      RECT  69.75 61.825 69.96 62.065 ;
      RECT  67.77 61.035 68.31 61.585 ;
      RECT  66.63 62.305 67.77 62.685 ;
      RECT  66.63 61.035 66.84 61.585 ;
      POLYGON  69.61 62.305 69.61 62.375 69.24 62.375 69.24 62.615 69.61 62.615 69.61 62.685 69.75 62.685 69.75 62.305 69.61 62.305 ;
      RECT  69.24 61.825 69.75 62.065 ;
      RECT  68.31 61.035 69.96 61.585 ;
      POLYGON  68.31 62.305 68.31 62.685 68.86 62.685 68.86 62.615 69.24 62.615 69.24 62.375 68.86 62.375 68.86 62.305 68.31 62.305 ;
      RECT  66.63 61.825 66.84 62.065 ;
      RECT  69.24 63.645 69.75 63.405 ;
      RECT  69.24 63.715 69.44 63.645 ;
      RECT  67.77 64.265 68.31 63.885 ;
      RECT  66.84 65.535 67.77 64.985 ;
      RECT  66.63 63.645 66.84 63.405 ;
      RECT  69.75 63.645 69.96 63.405 ;
      RECT  66.84 63.645 69.24 63.405 ;
      RECT  69.03 64.505 69.24 64.435 ;
      RECT  69.75 64.265 69.96 63.885 ;
      RECT  69.03 63.715 69.24 63.645 ;
      RECT  69.24 64.505 69.44 64.435 ;
      RECT  66.84 64.745 69.24 64.505 ;
      RECT  69.75 64.745 69.96 64.505 ;
      RECT  67.77 65.535 68.31 64.985 ;
      RECT  66.63 64.265 67.77 63.885 ;
      RECT  66.63 65.535 66.84 64.985 ;
      POLYGON  69.61 64.265 69.61 64.195 69.24 64.195 69.24 63.955 69.61 63.955 69.61 63.885 69.75 63.885 69.75 64.265 69.61 64.265 ;
      RECT  69.24 64.745 69.75 64.505 ;
      RECT  68.31 65.535 69.96 64.985 ;
      POLYGON  68.31 64.265 68.31 63.885 68.86 63.885 68.86 63.955 69.24 63.955 69.24 64.195 68.86 64.195 68.86 64.265 68.31 64.265 ;
      RECT  66.63 64.745 66.84 64.505 ;
      RECT  69.24 66.875 69.75 67.115 ;
      RECT  69.24 66.805 69.44 66.875 ;
      RECT  67.77 66.255 68.31 66.635 ;
      RECT  66.84 64.985 67.77 65.535 ;
      RECT  66.63 66.875 66.84 67.115 ;
      RECT  69.75 66.875 69.96 67.115 ;
      RECT  66.84 66.875 69.24 67.115 ;
      RECT  69.03 66.015 69.24 66.085 ;
      RECT  69.75 66.255 69.96 66.635 ;
      RECT  69.03 66.805 69.24 66.875 ;
      RECT  69.24 66.015 69.44 66.085 ;
      RECT  66.84 65.775 69.24 66.015 ;
      RECT  69.75 65.775 69.96 66.015 ;
      RECT  67.77 64.985 68.31 65.535 ;
      RECT  66.63 66.255 67.77 66.635 ;
      RECT  66.63 64.985 66.84 65.535 ;
      POLYGON  69.61 66.255 69.61 66.325 69.24 66.325 69.24 66.565 69.61 66.565 69.61 66.635 69.75 66.635 69.75 66.255 69.61 66.255 ;
      RECT  69.24 65.775 69.75 66.015 ;
      RECT  68.31 64.985 69.96 65.535 ;
      POLYGON  68.31 66.255 68.31 66.635 68.86 66.635 68.86 66.565 69.24 66.565 69.24 66.325 68.86 66.325 68.86 66.255 68.31 66.255 ;
      RECT  66.63 65.775 66.84 66.015 ;
      RECT  69.24 67.595 69.75 67.355 ;
      RECT  69.24 67.665 69.44 67.595 ;
      RECT  67.77 68.215 68.31 67.835 ;
      RECT  66.84 69.485 67.77 68.935 ;
      RECT  66.63 67.595 66.84 67.355 ;
      RECT  69.75 67.595 69.96 67.355 ;
      RECT  66.84 67.595 69.24 67.355 ;
      RECT  69.03 68.455 69.24 68.385 ;
      RECT  69.75 68.215 69.96 67.835 ;
      RECT  69.03 67.665 69.24 67.595 ;
      RECT  69.24 68.455 69.44 68.385 ;
      RECT  66.84 68.695 69.24 68.455 ;
      RECT  69.75 68.695 69.96 68.455 ;
      RECT  67.77 69.485 68.31 68.935 ;
      RECT  66.63 68.215 67.77 67.835 ;
      RECT  66.63 69.485 66.84 68.935 ;
      POLYGON  69.61 68.215 69.61 68.145 69.24 68.145 69.24 67.905 69.61 67.905 69.61 67.835 69.75 67.835 69.75 68.215 69.61 68.215 ;
      RECT  69.24 68.695 69.75 68.455 ;
      RECT  68.31 69.485 69.96 68.935 ;
      POLYGON  68.31 68.215 68.31 67.835 68.86 67.835 68.86 67.905 69.24 67.905 69.24 68.145 68.86 68.145 68.86 68.215 68.31 68.215 ;
      RECT  66.63 68.695 66.84 68.455 ;
      RECT  69.24 70.825 69.75 71.065 ;
      RECT  69.24 70.755 69.44 70.825 ;
      RECT  67.77 70.205 68.31 70.585 ;
      RECT  66.84 68.935 67.77 69.485 ;
      RECT  66.63 70.825 66.84 71.065 ;
      RECT  69.75 70.825 69.96 71.065 ;
      RECT  66.84 70.825 69.24 71.065 ;
      RECT  69.03 69.965 69.24 70.035 ;
      RECT  69.75 70.205 69.96 70.585 ;
      RECT  69.03 70.755 69.24 70.825 ;
      RECT  69.24 69.965 69.44 70.035 ;
      RECT  66.84 69.725 69.24 69.965 ;
      RECT  69.75 69.725 69.96 69.965 ;
      RECT  67.77 68.935 68.31 69.485 ;
      RECT  66.63 70.205 67.77 70.585 ;
      RECT  66.63 68.935 66.84 69.485 ;
      POLYGON  69.61 70.205 69.61 70.275 69.24 70.275 69.24 70.515 69.61 70.515 69.61 70.585 69.75 70.585 69.75 70.205 69.61 70.205 ;
      RECT  69.24 69.725 69.75 69.965 ;
      RECT  68.31 68.935 69.96 69.485 ;
      POLYGON  68.31 70.205 68.31 70.585 68.86 70.585 68.86 70.515 69.24 70.515 69.24 70.275 68.86 70.275 68.86 70.205 68.31 70.205 ;
      RECT  66.63 69.725 66.84 69.965 ;
      RECT  69.24 71.545 69.75 71.305 ;
      RECT  69.24 71.615 69.44 71.545 ;
      RECT  67.77 72.165 68.31 71.785 ;
      RECT  66.84 73.435 67.77 72.885 ;
      RECT  66.63 71.545 66.84 71.305 ;
      RECT  69.75 71.545 69.96 71.305 ;
      RECT  66.84 71.545 69.24 71.305 ;
      RECT  69.03 72.405 69.24 72.335 ;
      RECT  69.75 72.165 69.96 71.785 ;
      RECT  69.03 71.615 69.24 71.545 ;
      RECT  69.24 72.405 69.44 72.335 ;
      RECT  66.84 72.645 69.24 72.405 ;
      RECT  69.75 72.645 69.96 72.405 ;
      RECT  67.77 73.435 68.31 72.885 ;
      RECT  66.63 72.165 67.77 71.785 ;
      RECT  66.63 73.435 66.84 72.885 ;
      POLYGON  69.61 72.165 69.61 72.095 69.24 72.095 69.24 71.855 69.61 71.855 69.61 71.785 69.75 71.785 69.75 72.165 69.61 72.165 ;
      RECT  69.24 72.645 69.75 72.405 ;
      RECT  68.31 73.435 69.96 72.885 ;
      POLYGON  68.31 72.165 68.31 71.785 68.86 71.785 68.86 71.855 69.24 71.855 69.24 72.095 68.86 72.095 68.86 72.165 68.31 72.165 ;
      RECT  66.63 72.645 66.84 72.405 ;
      RECT  69.24 74.775 69.75 75.015 ;
      RECT  69.24 74.705 69.44 74.775 ;
      RECT  67.77 74.155 68.31 74.535 ;
      RECT  66.84 72.885 67.77 73.435 ;
      RECT  66.63 74.775 66.84 75.015 ;
      RECT  69.75 74.775 69.96 75.015 ;
      RECT  66.84 74.775 69.24 75.015 ;
      RECT  69.03 73.915 69.24 73.985 ;
      RECT  69.75 74.155 69.96 74.535 ;
      RECT  69.03 74.705 69.24 74.775 ;
      RECT  69.24 73.915 69.44 73.985 ;
      RECT  66.84 73.675 69.24 73.915 ;
      RECT  69.75 73.675 69.96 73.915 ;
      RECT  67.77 72.885 68.31 73.435 ;
      RECT  66.63 74.155 67.77 74.535 ;
      RECT  66.63 72.885 66.84 73.435 ;
      POLYGON  69.61 74.155 69.61 74.225 69.24 74.225 69.24 74.465 69.61 74.465 69.61 74.535 69.75 74.535 69.75 74.155 69.61 74.155 ;
      RECT  69.24 73.675 69.75 73.915 ;
      RECT  68.31 72.885 69.96 73.435 ;
      POLYGON  68.31 74.155 68.31 74.535 68.86 74.535 68.86 74.465 69.24 74.465 69.24 74.225 68.86 74.225 68.86 74.155 68.31 74.155 ;
      RECT  66.63 73.675 66.84 73.915 ;
      RECT  69.24 75.495 69.75 75.255 ;
      RECT  69.24 75.565 69.44 75.495 ;
      RECT  67.77 76.115 68.31 75.735 ;
      RECT  66.84 77.385 67.77 76.835 ;
      RECT  66.63 75.495 66.84 75.255 ;
      RECT  69.75 75.495 69.96 75.255 ;
      RECT  66.84 75.495 69.24 75.255 ;
      RECT  69.03 76.355 69.24 76.285 ;
      RECT  69.75 76.115 69.96 75.735 ;
      RECT  69.03 75.565 69.24 75.495 ;
      RECT  69.24 76.355 69.44 76.285 ;
      RECT  66.84 76.595 69.24 76.355 ;
      RECT  69.75 76.595 69.96 76.355 ;
      RECT  67.77 77.385 68.31 76.835 ;
      RECT  66.63 76.115 67.77 75.735 ;
      RECT  66.63 77.385 66.84 76.835 ;
      POLYGON  69.61 76.115 69.61 76.045 69.24 76.045 69.24 75.805 69.61 75.805 69.61 75.735 69.75 75.735 69.75 76.115 69.61 76.115 ;
      RECT  69.24 76.595 69.75 76.355 ;
      RECT  68.31 77.385 69.96 76.835 ;
      POLYGON  68.31 76.115 68.31 75.735 68.86 75.735 68.86 75.805 69.24 75.805 69.24 76.045 68.86 76.045 68.86 76.115 68.31 76.115 ;
      RECT  66.63 76.595 66.84 76.355 ;
      RECT  69.24 78.725 69.75 78.965 ;
      RECT  69.24 78.655 69.44 78.725 ;
      RECT  67.77 78.105 68.31 78.485 ;
      RECT  66.84 76.835 67.77 77.385 ;
      RECT  66.63 78.725 66.84 78.965 ;
      RECT  69.75 78.725 69.96 78.965 ;
      RECT  66.84 78.725 69.24 78.965 ;
      RECT  69.03 77.865 69.24 77.935 ;
      RECT  69.75 78.105 69.96 78.485 ;
      RECT  69.03 78.655 69.24 78.725 ;
      RECT  69.24 77.865 69.44 77.935 ;
      RECT  66.84 77.625 69.24 77.865 ;
      RECT  69.75 77.625 69.96 77.865 ;
      RECT  67.77 76.835 68.31 77.385 ;
      RECT  66.63 78.105 67.77 78.485 ;
      RECT  66.63 76.835 66.84 77.385 ;
      POLYGON  69.61 78.105 69.61 78.175 69.24 78.175 69.24 78.415 69.61 78.415 69.61 78.485 69.75 78.485 69.75 78.105 69.61 78.105 ;
      RECT  69.24 77.625 69.75 77.865 ;
      RECT  68.31 76.835 69.96 77.385 ;
      POLYGON  68.31 78.105 68.31 78.485 68.86 78.485 68.86 78.415 69.24 78.415 69.24 78.175 68.86 78.175 68.86 78.105 68.31 78.105 ;
      RECT  66.63 77.625 66.84 77.865 ;
      RECT  69.24 79.445 69.75 79.205 ;
      RECT  69.24 79.515 69.44 79.445 ;
      RECT  67.77 80.065 68.31 79.685 ;
      RECT  66.84 81.335 67.77 80.785 ;
      RECT  66.63 79.445 66.84 79.205 ;
      RECT  69.75 79.445 69.96 79.205 ;
      RECT  66.84 79.445 69.24 79.205 ;
      RECT  69.03 80.305 69.24 80.235 ;
      RECT  69.75 80.065 69.96 79.685 ;
      RECT  69.03 79.515 69.24 79.445 ;
      RECT  69.24 80.305 69.44 80.235 ;
      RECT  66.84 80.545 69.24 80.305 ;
      RECT  69.75 80.545 69.96 80.305 ;
      RECT  67.77 81.335 68.31 80.785 ;
      RECT  66.63 80.065 67.77 79.685 ;
      RECT  66.63 81.335 66.84 80.785 ;
      POLYGON  69.61 80.065 69.61 79.995 69.24 79.995 69.24 79.755 69.61 79.755 69.61 79.685 69.75 79.685 69.75 80.065 69.61 80.065 ;
      RECT  69.24 80.545 69.75 80.305 ;
      RECT  68.31 81.335 69.96 80.785 ;
      POLYGON  68.31 80.065 68.31 79.685 68.86 79.685 68.86 79.755 69.24 79.755 69.24 79.995 68.86 79.995 68.86 80.065 68.31 80.065 ;
      RECT  66.63 80.545 66.84 80.305 ;
      RECT  69.24 82.675 69.75 82.915 ;
      RECT  69.24 82.605 69.44 82.675 ;
      RECT  67.77 82.055 68.31 82.435 ;
      RECT  66.84 80.785 67.77 81.335 ;
      RECT  66.63 82.675 66.84 82.915 ;
      RECT  69.75 82.675 69.96 82.915 ;
      RECT  66.84 82.675 69.24 82.915 ;
      RECT  69.03 81.815 69.24 81.885 ;
      RECT  69.75 82.055 69.96 82.435 ;
      RECT  69.03 82.605 69.24 82.675 ;
      RECT  69.24 81.815 69.44 81.885 ;
      RECT  66.84 81.575 69.24 81.815 ;
      RECT  69.75 81.575 69.96 81.815 ;
      RECT  67.77 80.785 68.31 81.335 ;
      RECT  66.63 82.055 67.77 82.435 ;
      RECT  66.63 80.785 66.84 81.335 ;
      POLYGON  69.61 82.055 69.61 82.125 69.24 82.125 69.24 82.365 69.61 82.365 69.61 82.435 69.75 82.435 69.75 82.055 69.61 82.055 ;
      RECT  69.24 81.575 69.75 81.815 ;
      RECT  68.31 80.785 69.96 81.335 ;
      POLYGON  68.31 82.055 68.31 82.435 68.86 82.435 68.86 82.365 69.24 82.365 69.24 82.125 68.86 82.125 68.86 82.055 68.31 82.055 ;
      RECT  66.63 81.575 66.84 81.815 ;
      RECT  69.24 83.395 69.75 83.155 ;
      RECT  69.24 83.465 69.44 83.395 ;
      RECT  67.77 84.015 68.31 83.635 ;
      RECT  66.84 85.285 67.77 84.735 ;
      RECT  66.63 83.395 66.84 83.155 ;
      RECT  69.75 83.395 69.96 83.155 ;
      RECT  66.84 83.395 69.24 83.155 ;
      RECT  69.03 84.255 69.24 84.185 ;
      RECT  69.75 84.015 69.96 83.635 ;
      RECT  69.03 83.465 69.24 83.395 ;
      RECT  69.24 84.255 69.44 84.185 ;
      RECT  66.84 84.495 69.24 84.255 ;
      RECT  69.75 84.495 69.96 84.255 ;
      RECT  67.77 85.285 68.31 84.735 ;
      RECT  66.63 84.015 67.77 83.635 ;
      RECT  66.63 85.285 66.84 84.735 ;
      POLYGON  69.61 84.015 69.61 83.945 69.24 83.945 69.24 83.705 69.61 83.705 69.61 83.635 69.75 83.635 69.75 84.015 69.61 84.015 ;
      RECT  69.24 84.495 69.75 84.255 ;
      RECT  68.31 85.285 69.96 84.735 ;
      POLYGON  68.31 84.015 68.31 83.635 68.86 83.635 68.86 83.705 69.24 83.705 69.24 83.945 68.86 83.945 68.86 84.015 68.31 84.015 ;
      RECT  66.63 84.495 66.84 84.255 ;
      RECT  69.24 86.625 69.75 86.865 ;
      RECT  69.24 86.555 69.44 86.625 ;
      RECT  67.77 86.005 68.31 86.385 ;
      RECT  66.84 84.735 67.77 85.285 ;
      RECT  66.63 86.625 66.84 86.865 ;
      RECT  69.75 86.625 69.96 86.865 ;
      RECT  66.84 86.625 69.24 86.865 ;
      RECT  69.03 85.765 69.24 85.835 ;
      RECT  69.75 86.005 69.96 86.385 ;
      RECT  69.03 86.555 69.24 86.625 ;
      RECT  69.24 85.765 69.44 85.835 ;
      RECT  66.84 85.525 69.24 85.765 ;
      RECT  69.75 85.525 69.96 85.765 ;
      RECT  67.77 84.735 68.31 85.285 ;
      RECT  66.63 86.005 67.77 86.385 ;
      RECT  66.63 84.735 66.84 85.285 ;
      POLYGON  69.61 86.005 69.61 86.075 69.24 86.075 69.24 86.315 69.61 86.315 69.61 86.385 69.75 86.385 69.75 86.005 69.61 86.005 ;
      RECT  69.24 85.525 69.75 85.765 ;
      RECT  68.31 84.735 69.96 85.285 ;
      POLYGON  68.31 86.005 68.31 86.385 68.86 86.385 68.86 86.315 69.24 86.315 69.24 86.075 68.86 86.075 68.86 86.005 68.31 86.005 ;
      RECT  66.63 85.525 66.84 85.765 ;
      RECT  69.24 87.345 69.75 87.105 ;
      RECT  69.24 87.415 69.44 87.345 ;
      RECT  67.77 87.965 68.31 87.585 ;
      RECT  66.84 89.235 67.77 88.685 ;
      RECT  66.63 87.345 66.84 87.105 ;
      RECT  69.75 87.345 69.96 87.105 ;
      RECT  66.84 87.345 69.24 87.105 ;
      RECT  69.03 88.205 69.24 88.135 ;
      RECT  69.75 87.965 69.96 87.585 ;
      RECT  69.03 87.415 69.24 87.345 ;
      RECT  69.24 88.205 69.44 88.135 ;
      RECT  66.84 88.445 69.24 88.205 ;
      RECT  69.75 88.445 69.96 88.205 ;
      RECT  67.77 89.235 68.31 88.685 ;
      RECT  66.63 87.965 67.77 87.585 ;
      RECT  66.63 89.235 66.84 88.685 ;
      POLYGON  69.61 87.965 69.61 87.895 69.24 87.895 69.24 87.655 69.61 87.655 69.61 87.585 69.75 87.585 69.75 87.965 69.61 87.965 ;
      RECT  69.24 88.445 69.75 88.205 ;
      RECT  68.31 89.235 69.96 88.685 ;
      POLYGON  68.31 87.965 68.31 87.585 68.86 87.585 68.86 87.655 69.24 87.655 69.24 87.895 68.86 87.895 68.86 87.965 68.31 87.965 ;
      RECT  66.63 88.445 66.84 88.205 ;
      RECT  69.24 90.575 69.75 90.815 ;
      RECT  69.24 90.505 69.44 90.575 ;
      RECT  67.77 89.955 68.31 90.335 ;
      RECT  66.84 88.685 67.77 89.235 ;
      RECT  66.63 90.575 66.84 90.815 ;
      RECT  69.75 90.575 69.96 90.815 ;
      RECT  66.84 90.575 69.24 90.815 ;
      RECT  69.03 89.715 69.24 89.785 ;
      RECT  69.75 89.955 69.96 90.335 ;
      RECT  69.03 90.505 69.24 90.575 ;
      RECT  69.24 89.715 69.44 89.785 ;
      RECT  66.84 89.475 69.24 89.715 ;
      RECT  69.75 89.475 69.96 89.715 ;
      RECT  67.77 88.685 68.31 89.235 ;
      RECT  66.63 89.955 67.77 90.335 ;
      RECT  66.63 88.685 66.84 89.235 ;
      POLYGON  69.61 89.955 69.61 90.025 69.24 90.025 69.24 90.265 69.61 90.265 69.61 90.335 69.75 90.335 69.75 89.955 69.61 89.955 ;
      RECT  69.24 89.475 69.75 89.715 ;
      RECT  68.31 88.685 69.96 89.235 ;
      POLYGON  68.31 89.955 68.31 90.335 68.86 90.335 68.86 90.265 69.24 90.265 69.24 90.025 68.86 90.025 68.86 89.955 68.31 89.955 ;
      RECT  66.63 89.475 66.84 89.715 ;
      RECT  69.24 91.295 69.75 91.055 ;
      RECT  69.24 91.365 69.44 91.295 ;
      RECT  67.77 91.915 68.31 91.535 ;
      RECT  66.84 93.185 67.77 92.635 ;
      RECT  66.63 91.295 66.84 91.055 ;
      RECT  69.75 91.295 69.96 91.055 ;
      RECT  66.84 91.295 69.24 91.055 ;
      RECT  69.03 92.155 69.24 92.085 ;
      RECT  69.75 91.915 69.96 91.535 ;
      RECT  69.03 91.365 69.24 91.295 ;
      RECT  69.24 92.155 69.44 92.085 ;
      RECT  66.84 92.395 69.24 92.155 ;
      RECT  69.75 92.395 69.96 92.155 ;
      RECT  67.77 93.185 68.31 92.635 ;
      RECT  66.63 91.915 67.77 91.535 ;
      RECT  66.63 93.185 66.84 92.635 ;
      POLYGON  69.61 91.915 69.61 91.845 69.24 91.845 69.24 91.605 69.61 91.605 69.61 91.535 69.75 91.535 69.75 91.915 69.61 91.915 ;
      RECT  69.24 92.395 69.75 92.155 ;
      RECT  68.31 93.185 69.96 92.635 ;
      POLYGON  68.31 91.915 68.31 91.535 68.86 91.535 68.86 91.605 69.24 91.605 69.24 91.845 68.86 91.845 68.86 91.915 68.31 91.915 ;
      RECT  66.63 92.395 66.84 92.155 ;
      RECT  69.24 94.525 69.75 94.765 ;
      RECT  69.24 94.455 69.44 94.525 ;
      RECT  67.77 93.905 68.31 94.285 ;
      RECT  66.84 92.635 67.77 93.185 ;
      RECT  66.63 94.525 66.84 94.765 ;
      RECT  69.75 94.525 69.96 94.765 ;
      RECT  66.84 94.525 69.24 94.765 ;
      RECT  69.03 93.665 69.24 93.735 ;
      RECT  69.75 93.905 69.96 94.285 ;
      RECT  69.03 94.455 69.24 94.525 ;
      RECT  69.24 93.665 69.44 93.735 ;
      RECT  66.84 93.425 69.24 93.665 ;
      RECT  69.75 93.425 69.96 93.665 ;
      RECT  67.77 92.635 68.31 93.185 ;
      RECT  66.63 93.905 67.77 94.285 ;
      RECT  66.63 92.635 66.84 93.185 ;
      POLYGON  69.61 93.905 69.61 93.975 69.24 93.975 69.24 94.215 69.61 94.215 69.61 94.285 69.75 94.285 69.75 93.905 69.61 93.905 ;
      RECT  69.24 93.425 69.75 93.665 ;
      RECT  68.31 92.635 69.96 93.185 ;
      POLYGON  68.31 93.905 68.31 94.285 68.86 94.285 68.86 94.215 69.24 94.215 69.24 93.975 68.86 93.975 68.86 93.905 68.31 93.905 ;
      RECT  66.63 93.425 66.84 93.665 ;
      RECT  66.84 59.455 69.96 59.695 ;
      RECT  66.84 60.555 69.96 60.795 ;
      RECT  66.84 62.925 69.96 63.165 ;
      RECT  66.84 61.825 69.96 62.065 ;
      RECT  66.84 63.405 69.96 63.645 ;
      RECT  66.84 64.505 69.96 64.745 ;
      RECT  66.84 66.875 69.96 67.115 ;
      RECT  66.84 65.775 69.96 66.015 ;
      RECT  66.84 67.355 69.96 67.595 ;
      RECT  66.84 68.455 69.96 68.695 ;
      RECT  66.84 70.825 69.96 71.065 ;
      RECT  66.84 69.725 69.96 69.965 ;
      RECT  66.84 71.305 69.96 71.545 ;
      RECT  66.84 72.405 69.96 72.645 ;
      RECT  66.84 74.775 69.96 75.015 ;
      RECT  66.84 73.675 69.96 73.915 ;
      RECT  66.84 75.255 69.96 75.495 ;
      RECT  66.84 76.355 69.96 76.595 ;
      RECT  66.84 78.725 69.96 78.965 ;
      RECT  66.84 77.625 69.96 77.865 ;
      RECT  66.84 79.205 69.96 79.445 ;
      RECT  66.84 80.305 69.96 80.545 ;
      RECT  66.84 82.675 69.96 82.915 ;
      RECT  66.84 81.575 69.96 81.815 ;
      RECT  66.84 83.155 69.96 83.395 ;
      RECT  66.84 84.255 69.96 84.495 ;
      RECT  66.84 86.625 69.96 86.865 ;
      RECT  66.84 85.525 69.96 85.765 ;
      RECT  66.84 87.105 69.96 87.345 ;
      RECT  66.84 88.205 69.96 88.445 ;
      RECT  66.84 90.575 69.96 90.815 ;
      RECT  66.84 89.475 69.96 89.715 ;
      RECT  66.84 91.055 69.96 91.295 ;
      RECT  66.84 92.155 69.96 92.395 ;
      RECT  66.84 94.525 69.96 94.765 ;
      RECT  66.84 93.425 69.96 93.665 ;
      RECT  83.16 59.695 82.65 59.455 ;
      RECT  83.16 59.765 82.96 59.695 ;
      RECT  84.63 60.315 84.09 59.935 ;
      RECT  85.56 61.585 84.63 61.035 ;
      RECT  85.77 59.695 85.56 59.455 ;
      RECT  82.65 59.695 82.44 59.455 ;
      RECT  85.56 59.695 83.16 59.455 ;
      RECT  83.37 60.555 83.16 60.485 ;
      RECT  82.65 60.315 82.44 59.935 ;
      RECT  83.37 59.765 83.16 59.695 ;
      RECT  83.16 60.555 82.96 60.485 ;
      RECT  85.56 60.795 83.16 60.555 ;
      RECT  82.65 60.795 82.44 60.555 ;
      RECT  84.63 61.585 84.09 61.035 ;
      RECT  85.77 60.315 84.63 59.935 ;
      RECT  85.77 61.585 85.56 61.035 ;
      POLYGON  82.79 60.315 82.79 60.245 83.16 60.245 83.16 60.005 82.79 60.005 82.79 59.935 82.65 59.935 82.65 60.315 82.79 60.315 ;
      RECT  83.16 60.795 82.65 60.555 ;
      RECT  84.09 61.585 82.44 61.035 ;
      POLYGON  84.09 60.315 84.09 59.935 83.54 59.935 83.54 60.005 83.16 60.005 83.16 60.245 83.54 60.245 83.54 60.315 84.09 60.315 ;
      RECT  85.77 60.795 85.56 60.555 ;
      RECT  83.16 62.925 82.65 63.165 ;
      RECT  83.16 62.855 82.96 62.925 ;
      RECT  84.63 62.305 84.09 62.685 ;
      RECT  85.56 61.035 84.63 61.585 ;
      RECT  85.77 62.925 85.56 63.165 ;
      RECT  82.65 62.925 82.44 63.165 ;
      RECT  85.56 62.925 83.16 63.165 ;
      RECT  83.37 62.065 83.16 62.135 ;
      RECT  82.65 62.305 82.44 62.685 ;
      RECT  83.37 62.855 83.16 62.925 ;
      RECT  83.16 62.065 82.96 62.135 ;
      RECT  85.56 61.825 83.16 62.065 ;
      RECT  82.65 61.825 82.44 62.065 ;
      RECT  84.63 61.035 84.09 61.585 ;
      RECT  85.77 62.305 84.63 62.685 ;
      RECT  85.77 61.035 85.56 61.585 ;
      POLYGON  82.79 62.305 82.79 62.375 83.16 62.375 83.16 62.615 82.79 62.615 82.79 62.685 82.65 62.685 82.65 62.305 82.79 62.305 ;
      RECT  83.16 61.825 82.65 62.065 ;
      RECT  84.09 61.035 82.44 61.585 ;
      POLYGON  84.09 62.305 84.09 62.685 83.54 62.685 83.54 62.615 83.16 62.615 83.16 62.375 83.54 62.375 83.54 62.305 84.09 62.305 ;
      RECT  85.77 61.825 85.56 62.065 ;
      RECT  83.16 63.645 82.65 63.405 ;
      RECT  83.16 63.715 82.96 63.645 ;
      RECT  84.63 64.265 84.09 63.885 ;
      RECT  85.56 65.535 84.63 64.985 ;
      RECT  85.77 63.645 85.56 63.405 ;
      RECT  82.65 63.645 82.44 63.405 ;
      RECT  85.56 63.645 83.16 63.405 ;
      RECT  83.37 64.505 83.16 64.435 ;
      RECT  82.65 64.265 82.44 63.885 ;
      RECT  83.37 63.715 83.16 63.645 ;
      RECT  83.16 64.505 82.96 64.435 ;
      RECT  85.56 64.745 83.16 64.505 ;
      RECT  82.65 64.745 82.44 64.505 ;
      RECT  84.63 65.535 84.09 64.985 ;
      RECT  85.77 64.265 84.63 63.885 ;
      RECT  85.77 65.535 85.56 64.985 ;
      POLYGON  82.79 64.265 82.79 64.195 83.16 64.195 83.16 63.955 82.79 63.955 82.79 63.885 82.65 63.885 82.65 64.265 82.79 64.265 ;
      RECT  83.16 64.745 82.65 64.505 ;
      RECT  84.09 65.535 82.44 64.985 ;
      POLYGON  84.09 64.265 84.09 63.885 83.54 63.885 83.54 63.955 83.16 63.955 83.16 64.195 83.54 64.195 83.54 64.265 84.09 64.265 ;
      RECT  85.77 64.745 85.56 64.505 ;
      RECT  83.16 66.875 82.65 67.115 ;
      RECT  83.16 66.805 82.96 66.875 ;
      RECT  84.63 66.255 84.09 66.635 ;
      RECT  85.56 64.985 84.63 65.535 ;
      RECT  85.77 66.875 85.56 67.115 ;
      RECT  82.65 66.875 82.44 67.115 ;
      RECT  85.56 66.875 83.16 67.115 ;
      RECT  83.37 66.015 83.16 66.085 ;
      RECT  82.65 66.255 82.44 66.635 ;
      RECT  83.37 66.805 83.16 66.875 ;
      RECT  83.16 66.015 82.96 66.085 ;
      RECT  85.56 65.775 83.16 66.015 ;
      RECT  82.65 65.775 82.44 66.015 ;
      RECT  84.63 64.985 84.09 65.535 ;
      RECT  85.77 66.255 84.63 66.635 ;
      RECT  85.77 64.985 85.56 65.535 ;
      POLYGON  82.79 66.255 82.79 66.325 83.16 66.325 83.16 66.565 82.79 66.565 82.79 66.635 82.65 66.635 82.65 66.255 82.79 66.255 ;
      RECT  83.16 65.775 82.65 66.015 ;
      RECT  84.09 64.985 82.44 65.535 ;
      POLYGON  84.09 66.255 84.09 66.635 83.54 66.635 83.54 66.565 83.16 66.565 83.16 66.325 83.54 66.325 83.54 66.255 84.09 66.255 ;
      RECT  85.77 65.775 85.56 66.015 ;
      RECT  83.16 67.595 82.65 67.355 ;
      RECT  83.16 67.665 82.96 67.595 ;
      RECT  84.63 68.215 84.09 67.835 ;
      RECT  85.56 69.485 84.63 68.935 ;
      RECT  85.77 67.595 85.56 67.355 ;
      RECT  82.65 67.595 82.44 67.355 ;
      RECT  85.56 67.595 83.16 67.355 ;
      RECT  83.37 68.455 83.16 68.385 ;
      RECT  82.65 68.215 82.44 67.835 ;
      RECT  83.37 67.665 83.16 67.595 ;
      RECT  83.16 68.455 82.96 68.385 ;
      RECT  85.56 68.695 83.16 68.455 ;
      RECT  82.65 68.695 82.44 68.455 ;
      RECT  84.63 69.485 84.09 68.935 ;
      RECT  85.77 68.215 84.63 67.835 ;
      RECT  85.77 69.485 85.56 68.935 ;
      POLYGON  82.79 68.215 82.79 68.145 83.16 68.145 83.16 67.905 82.79 67.905 82.79 67.835 82.65 67.835 82.65 68.215 82.79 68.215 ;
      RECT  83.16 68.695 82.65 68.455 ;
      RECT  84.09 69.485 82.44 68.935 ;
      POLYGON  84.09 68.215 84.09 67.835 83.54 67.835 83.54 67.905 83.16 67.905 83.16 68.145 83.54 68.145 83.54 68.215 84.09 68.215 ;
      RECT  85.77 68.695 85.56 68.455 ;
      RECT  83.16 70.825 82.65 71.065 ;
      RECT  83.16 70.755 82.96 70.825 ;
      RECT  84.63 70.205 84.09 70.585 ;
      RECT  85.56 68.935 84.63 69.485 ;
      RECT  85.77 70.825 85.56 71.065 ;
      RECT  82.65 70.825 82.44 71.065 ;
      RECT  85.56 70.825 83.16 71.065 ;
      RECT  83.37 69.965 83.16 70.035 ;
      RECT  82.65 70.205 82.44 70.585 ;
      RECT  83.37 70.755 83.16 70.825 ;
      RECT  83.16 69.965 82.96 70.035 ;
      RECT  85.56 69.725 83.16 69.965 ;
      RECT  82.65 69.725 82.44 69.965 ;
      RECT  84.63 68.935 84.09 69.485 ;
      RECT  85.77 70.205 84.63 70.585 ;
      RECT  85.77 68.935 85.56 69.485 ;
      POLYGON  82.79 70.205 82.79 70.275 83.16 70.275 83.16 70.515 82.79 70.515 82.79 70.585 82.65 70.585 82.65 70.205 82.79 70.205 ;
      RECT  83.16 69.725 82.65 69.965 ;
      RECT  84.09 68.935 82.44 69.485 ;
      POLYGON  84.09 70.205 84.09 70.585 83.54 70.585 83.54 70.515 83.16 70.515 83.16 70.275 83.54 70.275 83.54 70.205 84.09 70.205 ;
      RECT  85.77 69.725 85.56 69.965 ;
      RECT  83.16 71.545 82.65 71.305 ;
      RECT  83.16 71.615 82.96 71.545 ;
      RECT  84.63 72.165 84.09 71.785 ;
      RECT  85.56 73.435 84.63 72.885 ;
      RECT  85.77 71.545 85.56 71.305 ;
      RECT  82.65 71.545 82.44 71.305 ;
      RECT  85.56 71.545 83.16 71.305 ;
      RECT  83.37 72.405 83.16 72.335 ;
      RECT  82.65 72.165 82.44 71.785 ;
      RECT  83.37 71.615 83.16 71.545 ;
      RECT  83.16 72.405 82.96 72.335 ;
      RECT  85.56 72.645 83.16 72.405 ;
      RECT  82.65 72.645 82.44 72.405 ;
      RECT  84.63 73.435 84.09 72.885 ;
      RECT  85.77 72.165 84.63 71.785 ;
      RECT  85.77 73.435 85.56 72.885 ;
      POLYGON  82.79 72.165 82.79 72.095 83.16 72.095 83.16 71.855 82.79 71.855 82.79 71.785 82.65 71.785 82.65 72.165 82.79 72.165 ;
      RECT  83.16 72.645 82.65 72.405 ;
      RECT  84.09 73.435 82.44 72.885 ;
      POLYGON  84.09 72.165 84.09 71.785 83.54 71.785 83.54 71.855 83.16 71.855 83.16 72.095 83.54 72.095 83.54 72.165 84.09 72.165 ;
      RECT  85.77 72.645 85.56 72.405 ;
      RECT  83.16 74.775 82.65 75.015 ;
      RECT  83.16 74.705 82.96 74.775 ;
      RECT  84.63 74.155 84.09 74.535 ;
      RECT  85.56 72.885 84.63 73.435 ;
      RECT  85.77 74.775 85.56 75.015 ;
      RECT  82.65 74.775 82.44 75.015 ;
      RECT  85.56 74.775 83.16 75.015 ;
      RECT  83.37 73.915 83.16 73.985 ;
      RECT  82.65 74.155 82.44 74.535 ;
      RECT  83.37 74.705 83.16 74.775 ;
      RECT  83.16 73.915 82.96 73.985 ;
      RECT  85.56 73.675 83.16 73.915 ;
      RECT  82.65 73.675 82.44 73.915 ;
      RECT  84.63 72.885 84.09 73.435 ;
      RECT  85.77 74.155 84.63 74.535 ;
      RECT  85.77 72.885 85.56 73.435 ;
      POLYGON  82.79 74.155 82.79 74.225 83.16 74.225 83.16 74.465 82.79 74.465 82.79 74.535 82.65 74.535 82.65 74.155 82.79 74.155 ;
      RECT  83.16 73.675 82.65 73.915 ;
      RECT  84.09 72.885 82.44 73.435 ;
      POLYGON  84.09 74.155 84.09 74.535 83.54 74.535 83.54 74.465 83.16 74.465 83.16 74.225 83.54 74.225 83.54 74.155 84.09 74.155 ;
      RECT  85.77 73.675 85.56 73.915 ;
      RECT  83.16 75.495 82.65 75.255 ;
      RECT  83.16 75.565 82.96 75.495 ;
      RECT  84.63 76.115 84.09 75.735 ;
      RECT  85.56 77.385 84.63 76.835 ;
      RECT  85.77 75.495 85.56 75.255 ;
      RECT  82.65 75.495 82.44 75.255 ;
      RECT  85.56 75.495 83.16 75.255 ;
      RECT  83.37 76.355 83.16 76.285 ;
      RECT  82.65 76.115 82.44 75.735 ;
      RECT  83.37 75.565 83.16 75.495 ;
      RECT  83.16 76.355 82.96 76.285 ;
      RECT  85.56 76.595 83.16 76.355 ;
      RECT  82.65 76.595 82.44 76.355 ;
      RECT  84.63 77.385 84.09 76.835 ;
      RECT  85.77 76.115 84.63 75.735 ;
      RECT  85.77 77.385 85.56 76.835 ;
      POLYGON  82.79 76.115 82.79 76.045 83.16 76.045 83.16 75.805 82.79 75.805 82.79 75.735 82.65 75.735 82.65 76.115 82.79 76.115 ;
      RECT  83.16 76.595 82.65 76.355 ;
      RECT  84.09 77.385 82.44 76.835 ;
      POLYGON  84.09 76.115 84.09 75.735 83.54 75.735 83.54 75.805 83.16 75.805 83.16 76.045 83.54 76.045 83.54 76.115 84.09 76.115 ;
      RECT  85.77 76.595 85.56 76.355 ;
      RECT  83.16 78.725 82.65 78.965 ;
      RECT  83.16 78.655 82.96 78.725 ;
      RECT  84.63 78.105 84.09 78.485 ;
      RECT  85.56 76.835 84.63 77.385 ;
      RECT  85.77 78.725 85.56 78.965 ;
      RECT  82.65 78.725 82.44 78.965 ;
      RECT  85.56 78.725 83.16 78.965 ;
      RECT  83.37 77.865 83.16 77.935 ;
      RECT  82.65 78.105 82.44 78.485 ;
      RECT  83.37 78.655 83.16 78.725 ;
      RECT  83.16 77.865 82.96 77.935 ;
      RECT  85.56 77.625 83.16 77.865 ;
      RECT  82.65 77.625 82.44 77.865 ;
      RECT  84.63 76.835 84.09 77.385 ;
      RECT  85.77 78.105 84.63 78.485 ;
      RECT  85.77 76.835 85.56 77.385 ;
      POLYGON  82.79 78.105 82.79 78.175 83.16 78.175 83.16 78.415 82.79 78.415 82.79 78.485 82.65 78.485 82.65 78.105 82.79 78.105 ;
      RECT  83.16 77.625 82.65 77.865 ;
      RECT  84.09 76.835 82.44 77.385 ;
      POLYGON  84.09 78.105 84.09 78.485 83.54 78.485 83.54 78.415 83.16 78.415 83.16 78.175 83.54 78.175 83.54 78.105 84.09 78.105 ;
      RECT  85.77 77.625 85.56 77.865 ;
      RECT  83.16 79.445 82.65 79.205 ;
      RECT  83.16 79.515 82.96 79.445 ;
      RECT  84.63 80.065 84.09 79.685 ;
      RECT  85.56 81.335 84.63 80.785 ;
      RECT  85.77 79.445 85.56 79.205 ;
      RECT  82.65 79.445 82.44 79.205 ;
      RECT  85.56 79.445 83.16 79.205 ;
      RECT  83.37 80.305 83.16 80.235 ;
      RECT  82.65 80.065 82.44 79.685 ;
      RECT  83.37 79.515 83.16 79.445 ;
      RECT  83.16 80.305 82.96 80.235 ;
      RECT  85.56 80.545 83.16 80.305 ;
      RECT  82.65 80.545 82.44 80.305 ;
      RECT  84.63 81.335 84.09 80.785 ;
      RECT  85.77 80.065 84.63 79.685 ;
      RECT  85.77 81.335 85.56 80.785 ;
      POLYGON  82.79 80.065 82.79 79.995 83.16 79.995 83.16 79.755 82.79 79.755 82.79 79.685 82.65 79.685 82.65 80.065 82.79 80.065 ;
      RECT  83.16 80.545 82.65 80.305 ;
      RECT  84.09 81.335 82.44 80.785 ;
      POLYGON  84.09 80.065 84.09 79.685 83.54 79.685 83.54 79.755 83.16 79.755 83.16 79.995 83.54 79.995 83.54 80.065 84.09 80.065 ;
      RECT  85.77 80.545 85.56 80.305 ;
      RECT  83.16 82.675 82.65 82.915 ;
      RECT  83.16 82.605 82.96 82.675 ;
      RECT  84.63 82.055 84.09 82.435 ;
      RECT  85.56 80.785 84.63 81.335 ;
      RECT  85.77 82.675 85.56 82.915 ;
      RECT  82.65 82.675 82.44 82.915 ;
      RECT  85.56 82.675 83.16 82.915 ;
      RECT  83.37 81.815 83.16 81.885 ;
      RECT  82.65 82.055 82.44 82.435 ;
      RECT  83.37 82.605 83.16 82.675 ;
      RECT  83.16 81.815 82.96 81.885 ;
      RECT  85.56 81.575 83.16 81.815 ;
      RECT  82.65 81.575 82.44 81.815 ;
      RECT  84.63 80.785 84.09 81.335 ;
      RECT  85.77 82.055 84.63 82.435 ;
      RECT  85.77 80.785 85.56 81.335 ;
      POLYGON  82.79 82.055 82.79 82.125 83.16 82.125 83.16 82.365 82.79 82.365 82.79 82.435 82.65 82.435 82.65 82.055 82.79 82.055 ;
      RECT  83.16 81.575 82.65 81.815 ;
      RECT  84.09 80.785 82.44 81.335 ;
      POLYGON  84.09 82.055 84.09 82.435 83.54 82.435 83.54 82.365 83.16 82.365 83.16 82.125 83.54 82.125 83.54 82.055 84.09 82.055 ;
      RECT  85.77 81.575 85.56 81.815 ;
      RECT  83.16 83.395 82.65 83.155 ;
      RECT  83.16 83.465 82.96 83.395 ;
      RECT  84.63 84.015 84.09 83.635 ;
      RECT  85.56 85.285 84.63 84.735 ;
      RECT  85.77 83.395 85.56 83.155 ;
      RECT  82.65 83.395 82.44 83.155 ;
      RECT  85.56 83.395 83.16 83.155 ;
      RECT  83.37 84.255 83.16 84.185 ;
      RECT  82.65 84.015 82.44 83.635 ;
      RECT  83.37 83.465 83.16 83.395 ;
      RECT  83.16 84.255 82.96 84.185 ;
      RECT  85.56 84.495 83.16 84.255 ;
      RECT  82.65 84.495 82.44 84.255 ;
      RECT  84.63 85.285 84.09 84.735 ;
      RECT  85.77 84.015 84.63 83.635 ;
      RECT  85.77 85.285 85.56 84.735 ;
      POLYGON  82.79 84.015 82.79 83.945 83.16 83.945 83.16 83.705 82.79 83.705 82.79 83.635 82.65 83.635 82.65 84.015 82.79 84.015 ;
      RECT  83.16 84.495 82.65 84.255 ;
      RECT  84.09 85.285 82.44 84.735 ;
      POLYGON  84.09 84.015 84.09 83.635 83.54 83.635 83.54 83.705 83.16 83.705 83.16 83.945 83.54 83.945 83.54 84.015 84.09 84.015 ;
      RECT  85.77 84.495 85.56 84.255 ;
      RECT  83.16 86.625 82.65 86.865 ;
      RECT  83.16 86.555 82.96 86.625 ;
      RECT  84.63 86.005 84.09 86.385 ;
      RECT  85.56 84.735 84.63 85.285 ;
      RECT  85.77 86.625 85.56 86.865 ;
      RECT  82.65 86.625 82.44 86.865 ;
      RECT  85.56 86.625 83.16 86.865 ;
      RECT  83.37 85.765 83.16 85.835 ;
      RECT  82.65 86.005 82.44 86.385 ;
      RECT  83.37 86.555 83.16 86.625 ;
      RECT  83.16 85.765 82.96 85.835 ;
      RECT  85.56 85.525 83.16 85.765 ;
      RECT  82.65 85.525 82.44 85.765 ;
      RECT  84.63 84.735 84.09 85.285 ;
      RECT  85.77 86.005 84.63 86.385 ;
      RECT  85.77 84.735 85.56 85.285 ;
      POLYGON  82.79 86.005 82.79 86.075 83.16 86.075 83.16 86.315 82.79 86.315 82.79 86.385 82.65 86.385 82.65 86.005 82.79 86.005 ;
      RECT  83.16 85.525 82.65 85.765 ;
      RECT  84.09 84.735 82.44 85.285 ;
      POLYGON  84.09 86.005 84.09 86.385 83.54 86.385 83.54 86.315 83.16 86.315 83.16 86.075 83.54 86.075 83.54 86.005 84.09 86.005 ;
      RECT  85.77 85.525 85.56 85.765 ;
      RECT  83.16 87.345 82.65 87.105 ;
      RECT  83.16 87.415 82.96 87.345 ;
      RECT  84.63 87.965 84.09 87.585 ;
      RECT  85.56 89.235 84.63 88.685 ;
      RECT  85.77 87.345 85.56 87.105 ;
      RECT  82.65 87.345 82.44 87.105 ;
      RECT  85.56 87.345 83.16 87.105 ;
      RECT  83.37 88.205 83.16 88.135 ;
      RECT  82.65 87.965 82.44 87.585 ;
      RECT  83.37 87.415 83.16 87.345 ;
      RECT  83.16 88.205 82.96 88.135 ;
      RECT  85.56 88.445 83.16 88.205 ;
      RECT  82.65 88.445 82.44 88.205 ;
      RECT  84.63 89.235 84.09 88.685 ;
      RECT  85.77 87.965 84.63 87.585 ;
      RECT  85.77 89.235 85.56 88.685 ;
      POLYGON  82.79 87.965 82.79 87.895 83.16 87.895 83.16 87.655 82.79 87.655 82.79 87.585 82.65 87.585 82.65 87.965 82.79 87.965 ;
      RECT  83.16 88.445 82.65 88.205 ;
      RECT  84.09 89.235 82.44 88.685 ;
      POLYGON  84.09 87.965 84.09 87.585 83.54 87.585 83.54 87.655 83.16 87.655 83.16 87.895 83.54 87.895 83.54 87.965 84.09 87.965 ;
      RECT  85.77 88.445 85.56 88.205 ;
      RECT  83.16 90.575 82.65 90.815 ;
      RECT  83.16 90.505 82.96 90.575 ;
      RECT  84.63 89.955 84.09 90.335 ;
      RECT  85.56 88.685 84.63 89.235 ;
      RECT  85.77 90.575 85.56 90.815 ;
      RECT  82.65 90.575 82.44 90.815 ;
      RECT  85.56 90.575 83.16 90.815 ;
      RECT  83.37 89.715 83.16 89.785 ;
      RECT  82.65 89.955 82.44 90.335 ;
      RECT  83.37 90.505 83.16 90.575 ;
      RECT  83.16 89.715 82.96 89.785 ;
      RECT  85.56 89.475 83.16 89.715 ;
      RECT  82.65 89.475 82.44 89.715 ;
      RECT  84.63 88.685 84.09 89.235 ;
      RECT  85.77 89.955 84.63 90.335 ;
      RECT  85.77 88.685 85.56 89.235 ;
      POLYGON  82.79 89.955 82.79 90.025 83.16 90.025 83.16 90.265 82.79 90.265 82.79 90.335 82.65 90.335 82.65 89.955 82.79 89.955 ;
      RECT  83.16 89.475 82.65 89.715 ;
      RECT  84.09 88.685 82.44 89.235 ;
      POLYGON  84.09 89.955 84.09 90.335 83.54 90.335 83.54 90.265 83.16 90.265 83.16 90.025 83.54 90.025 83.54 89.955 84.09 89.955 ;
      RECT  85.77 89.475 85.56 89.715 ;
      RECT  83.16 91.295 82.65 91.055 ;
      RECT  83.16 91.365 82.96 91.295 ;
      RECT  84.63 91.915 84.09 91.535 ;
      RECT  85.56 93.185 84.63 92.635 ;
      RECT  85.77 91.295 85.56 91.055 ;
      RECT  82.65 91.295 82.44 91.055 ;
      RECT  85.56 91.295 83.16 91.055 ;
      RECT  83.37 92.155 83.16 92.085 ;
      RECT  82.65 91.915 82.44 91.535 ;
      RECT  83.37 91.365 83.16 91.295 ;
      RECT  83.16 92.155 82.96 92.085 ;
      RECT  85.56 92.395 83.16 92.155 ;
      RECT  82.65 92.395 82.44 92.155 ;
      RECT  84.63 93.185 84.09 92.635 ;
      RECT  85.77 91.915 84.63 91.535 ;
      RECT  85.77 93.185 85.56 92.635 ;
      POLYGON  82.79 91.915 82.79 91.845 83.16 91.845 83.16 91.605 82.79 91.605 82.79 91.535 82.65 91.535 82.65 91.915 82.79 91.915 ;
      RECT  83.16 92.395 82.65 92.155 ;
      RECT  84.09 93.185 82.44 92.635 ;
      POLYGON  84.09 91.915 84.09 91.535 83.54 91.535 83.54 91.605 83.16 91.605 83.16 91.845 83.54 91.845 83.54 91.915 84.09 91.915 ;
      RECT  85.77 92.395 85.56 92.155 ;
      RECT  83.16 94.525 82.65 94.765 ;
      RECT  83.16 94.455 82.96 94.525 ;
      RECT  84.63 93.905 84.09 94.285 ;
      RECT  85.56 92.635 84.63 93.185 ;
      RECT  85.77 94.525 85.56 94.765 ;
      RECT  82.65 94.525 82.44 94.765 ;
      RECT  85.56 94.525 83.16 94.765 ;
      RECT  83.37 93.665 83.16 93.735 ;
      RECT  82.65 93.905 82.44 94.285 ;
      RECT  83.37 94.455 83.16 94.525 ;
      RECT  83.16 93.665 82.96 93.735 ;
      RECT  85.56 93.425 83.16 93.665 ;
      RECT  82.65 93.425 82.44 93.665 ;
      RECT  84.63 92.635 84.09 93.185 ;
      RECT  85.77 93.905 84.63 94.285 ;
      RECT  85.77 92.635 85.56 93.185 ;
      POLYGON  82.79 93.905 82.79 93.975 83.16 93.975 83.16 94.215 82.79 94.215 82.79 94.285 82.65 94.285 82.65 93.905 82.79 93.905 ;
      RECT  83.16 93.425 82.65 93.665 ;
      RECT  84.09 92.635 82.44 93.185 ;
      POLYGON  84.09 93.905 84.09 94.285 83.54 94.285 83.54 94.215 83.16 94.215 83.16 93.975 83.54 93.975 83.54 93.905 84.09 93.905 ;
      RECT  85.77 93.425 85.56 93.665 ;
      RECT  82.44 59.455 85.56 59.695 ;
      RECT  82.44 60.555 85.56 60.795 ;
      RECT  82.44 62.925 85.56 63.165 ;
      RECT  82.44 61.825 85.56 62.065 ;
      RECT  82.44 63.405 85.56 63.645 ;
      RECT  82.44 64.505 85.56 64.745 ;
      RECT  82.44 66.875 85.56 67.115 ;
      RECT  82.44 65.775 85.56 66.015 ;
      RECT  82.44 67.355 85.56 67.595 ;
      RECT  82.44 68.455 85.56 68.695 ;
      RECT  82.44 70.825 85.56 71.065 ;
      RECT  82.44 69.725 85.56 69.965 ;
      RECT  82.44 71.305 85.56 71.545 ;
      RECT  82.44 72.405 85.56 72.645 ;
      RECT  82.44 74.775 85.56 75.015 ;
      RECT  82.44 73.675 85.56 73.915 ;
      RECT  82.44 75.255 85.56 75.495 ;
      RECT  82.44 76.355 85.56 76.595 ;
      RECT  82.44 78.725 85.56 78.965 ;
      RECT  82.44 77.625 85.56 77.865 ;
      RECT  82.44 79.205 85.56 79.445 ;
      RECT  82.44 80.305 85.56 80.545 ;
      RECT  82.44 82.675 85.56 82.915 ;
      RECT  82.44 81.575 85.56 81.815 ;
      RECT  82.44 83.155 85.56 83.395 ;
      RECT  82.44 84.255 85.56 84.495 ;
      RECT  82.44 86.625 85.56 86.865 ;
      RECT  82.44 85.525 85.56 85.765 ;
      RECT  82.44 87.105 85.56 87.345 ;
      RECT  82.44 88.205 85.56 88.445 ;
      RECT  82.44 90.575 85.56 90.815 ;
      RECT  82.44 89.475 85.56 89.715 ;
      RECT  82.44 91.055 85.56 91.295 ;
      RECT  82.44 92.155 85.56 92.395 ;
      RECT  82.44 94.525 85.56 94.765 ;
      RECT  82.44 93.425 85.56 93.665 ;
      RECT  66.84 62.925 85.56 63.165 ;
      RECT  66.84 61.825 85.56 62.065 ;
      RECT  66.84 63.405 85.56 63.645 ;
      RECT  66.84 64.505 85.56 64.745 ;
      RECT  66.84 66.875 85.56 67.115 ;
      RECT  66.84 65.775 85.56 66.015 ;
      RECT  66.84 67.355 85.56 67.595 ;
      RECT  66.84 68.455 85.56 68.695 ;
      RECT  66.84 70.825 85.56 71.065 ;
      RECT  66.84 69.725 85.56 69.965 ;
      RECT  66.84 71.305 85.56 71.545 ;
      RECT  66.84 72.405 85.56 72.645 ;
      RECT  66.84 74.775 85.56 75.015 ;
      RECT  66.84 73.675 85.56 73.915 ;
      RECT  66.84 75.255 85.56 75.495 ;
      RECT  66.84 76.355 85.56 76.595 ;
      RECT  66.84 78.725 85.56 78.965 ;
      RECT  66.84 77.625 85.56 77.865 ;
      RECT  66.84 79.205 85.56 79.445 ;
      RECT  66.84 80.305 85.56 80.545 ;
      RECT  66.84 82.675 85.56 82.915 ;
      RECT  66.84 81.575 85.56 81.815 ;
      RECT  66.84 83.155 85.56 83.395 ;
      RECT  66.84 84.255 85.56 84.495 ;
      RECT  66.84 86.625 85.56 86.865 ;
      RECT  66.84 85.525 85.56 85.765 ;
      RECT  66.84 87.105 85.56 87.345 ;
      RECT  66.84 88.205 85.56 88.445 ;
      RECT  66.84 90.575 85.56 90.815 ;
      RECT  66.84 89.475 85.56 89.715 ;
      RECT  66.84 91.055 85.56 91.295 ;
      RECT  66.84 92.155 85.56 92.395 ;
      RECT  66.84 59.455 85.56 59.695 ;
      RECT  66.84 93.425 85.56 93.665 ;
      RECT  80.25 87.585 80.79 87.965 ;
      RECT  71.61 70.205 72.15 70.585 ;
      RECT  71.61 72.885 72.15 73.435 ;
      RECT  71.61 87.585 72.15 87.965 ;
      RECT  71.61 59.935 72.15 60.315 ;
      RECT  71.61 83.635 72.15 84.015 ;
      RECT  80.25 79.685 80.79 80.065 ;
      RECT  80.25 91.535 80.79 91.915 ;
      RECT  80.25 63.885 80.79 64.265 ;
      RECT  80.25 64.985 80.79 65.535 ;
      RECT  71.61 86.005 72.15 86.385 ;
      RECT  80.25 62.305 80.79 62.685 ;
      RECT  71.61 61.035 72.15 61.585 ;
      RECT  71.61 62.305 72.15 62.685 ;
      RECT  71.61 78.105 72.15 78.485 ;
      RECT  80.25 80.785 80.79 81.335 ;
      RECT  71.61 93.905 72.15 94.285 ;
      RECT  80.25 71.785 80.79 72.165 ;
      RECT  80.25 76.835 80.79 77.385 ;
      RECT  71.61 91.535 72.15 91.915 ;
      RECT  80.25 84.735 80.79 85.285 ;
      RECT  80.25 59.935 80.79 60.315 ;
      RECT  80.25 83.635 80.79 84.015 ;
      RECT  71.61 74.155 72.15 74.535 ;
      RECT  80.25 74.155 80.79 74.535 ;
      RECT  80.25 67.835 80.79 68.215 ;
      RECT  71.61 82.055 72.15 82.435 ;
      RECT  71.61 67.835 72.15 68.215 ;
      RECT  80.25 82.055 80.79 82.435 ;
      RECT  71.61 92.635 72.15 93.185 ;
      RECT  80.25 68.935 80.79 69.485 ;
      RECT  71.61 88.685 72.15 89.235 ;
      RECT  80.25 88.685 80.79 89.235 ;
      RECT  80.25 86.005 80.79 86.385 ;
      RECT  80.25 70.205 80.79 70.585 ;
      RECT  80.25 92.635 80.79 93.185 ;
      RECT  80.25 66.255 80.79 66.635 ;
      RECT  71.61 84.735 72.15 85.285 ;
      RECT  80.25 78.105 80.79 78.485 ;
      RECT  71.61 71.785 72.15 72.165 ;
      RECT  71.61 66.255 72.15 66.635 ;
      RECT  80.25 61.035 80.79 61.585 ;
      RECT  71.61 89.955 72.15 90.335 ;
      RECT  80.25 89.955 80.79 90.335 ;
      RECT  71.61 63.885 72.15 64.265 ;
      RECT  71.61 79.685 72.15 80.065 ;
      RECT  71.61 76.835 72.15 77.385 ;
      RECT  80.25 93.905 80.79 94.285 ;
      RECT  71.61 68.935 72.15 69.485 ;
      RECT  71.61 64.985 72.15 65.535 ;
      RECT  71.61 80.785 72.15 81.335 ;
      RECT  80.25 75.735 80.79 76.115 ;
      RECT  71.61 75.735 72.15 76.115 ;
      RECT  80.25 72.885 80.79 73.435 ;
      RECT  73.08 52.385 69.96 52.525 ;
      RECT  73.08 52.385 76.2 52.525 ;
      RECT  79.32 52.385 76.2 52.525 ;
      RECT  73.08 101.835 76.2 101.695 ;
      RECT  79.32 101.835 76.2 101.695 ;
      RECT  79.32 101.835 82.44 101.695 ;
      RECT  56.02 61.31 56.16 92.91 ;
      RECT  56.02 61.31 56.16 92.91 ;
      RECT  96.38 61.31 96.24 92.91 ;
      RECT  96.38 61.31 96.24 92.91 ;
      RECT  63.74 28.475 63.88 60.51 ;
      RECT  87.42 93.71 87.56 114.85 ;
      RECT  64.98 28.475 65.12 60.51 ;
      RECT  86.8 93.71 86.94 114.85 ;
      RECT  64.36 28.475 64.5 60.51 ;
      RECT  65.6 28.475 65.74 60.51 ;
      RECT  86.18 93.71 86.32 114.85 ;
      RECT  5.41 3.045 5.74 3.305 ;
      RECT  0.685 2.69 1.015 2.95 ;
      RECT  5.02 2.29 5.35 2.55 ;
      RECT  1.845 3.46 2.115 3.78 ;
      RECT  0.685 2.69 1.015 2.95 ;
      RECT  10.37 2.445 10.51 2.585 ;
      RECT  7.84 4.355 7.98 4.495 ;
      RECT  1.845 3.46 2.115 3.78 ;
      RECT  5.41 11.095 5.74 10.835 ;
      RECT  0.685 11.45 1.015 11.19 ;
      RECT  5.02 11.85 5.35 11.59 ;
      RECT  1.845 10.68 2.115 10.36 ;
      RECT  0.685 11.45 1.015 11.19 ;
      RECT  10.37 11.695 10.51 11.555 ;
      RECT  7.84 9.785 7.98 9.645 ;
      RECT  1.845 10.68 2.115 10.36 ;
      RECT  0.685 2.69 1.015 2.95 ;
      RECT  0.685 11.19 1.015 11.45 ;
      RECT  10.37 2.445 10.51 2.585 ;
      RECT  7.84 4.355 7.98 4.495 ;
      RECT  10.37 11.555 10.51 11.695 ;
      RECT  7.84 9.645 7.98 9.785 ;
      RECT  1.845 0.0 1.985 14.14 ;
      RECT  8.88 57.36 8.74 59.97 ;
      RECT  1.085 57.36 0.945 104.77 ;
      RECT  0.685 2.69 1.015 2.95 ;
      RECT  0.685 11.19 1.015 11.45 ;
      RECT  15.435 3.275 15.575 3.415 ;
      RECT  8.74 57.36 8.88 59.97 ;
      RECT  18.49 53.085 27.23 53.225 ;
      RECT  19.57 31.745 27.23 31.885 ;
      RECT  20.26 39.005 27.23 39.145 ;
      RECT  21.59 24.675 27.23 24.815 ;
      RECT  24.32 3.465 27.23 3.605 ;
      RECT  145.88 137.035 145.55 136.775 ;
      RECT  150.605 137.39 150.275 137.13 ;
      RECT  146.27 137.79 145.94 137.53 ;
      RECT  149.445 136.62 149.175 136.3 ;
      RECT  150.605 137.39 150.275 137.13 ;
      RECT  140.92 137.635 140.78 137.495 ;
      RECT  143.45 135.725 143.31 135.585 ;
      RECT  149.445 136.62 149.175 136.3 ;
      RECT  150.605 137.39 150.275 137.13 ;
      RECT  140.92 137.635 140.78 137.495 ;
      RECT  143.45 135.725 143.31 135.585 ;
      RECT  149.445 140.08 149.305 133.01 ;
      RECT  142.41 96.86 142.55 94.25 ;
      RECT  150.205 96.86 150.345 49.45 ;
      RECT  150.605 137.39 150.275 137.13 ;
      RECT  136.275 136.805 136.135 136.665 ;
      RECT  142.55 96.86 142.41 94.25 ;
      RECT  133.22 101.135 125.59 100.995 ;
      RECT  131.45 108.525 125.59 108.385 ;
      RECT  130.12 115.405 125.59 115.265 ;
      RECT  128.46 136.695 125.59 136.555 ;
      RECT  26.8 111.605 27.13 111.865 ;
      RECT  22.075 111.25 22.405 111.51 ;
      RECT  26.41 110.85 26.74 111.11 ;
      RECT  23.235 112.02 23.505 112.34 ;
      RECT  26.8 119.655 27.13 119.395 ;
      RECT  22.075 120.01 22.405 119.75 ;
      RECT  26.41 120.41 26.74 120.15 ;
      RECT  23.235 119.24 23.505 118.92 ;
      RECT  26.8 125.745 27.13 126.005 ;
      RECT  22.075 125.39 22.405 125.65 ;
      RECT  26.41 124.99 26.74 125.25 ;
      RECT  23.235 126.16 23.505 126.48 ;
      RECT  26.8 133.795 27.13 133.535 ;
      RECT  22.075 134.15 22.405 133.89 ;
      RECT  26.41 134.55 26.74 134.29 ;
      RECT  23.235 133.38 23.505 133.06 ;
      RECT  22.075 111.25 22.405 111.51 ;
      RECT  22.075 119.75 22.405 120.01 ;
      RECT  22.075 125.39 22.405 125.65 ;
      RECT  22.075 133.89 22.405 134.15 ;
      RECT  26.8 111.605 27.13 111.865 ;
      RECT  26.8 119.395 27.13 119.655 ;
      RECT  26.8 125.745 27.13 126.005 ;
      RECT  26.8 133.535 27.13 133.795 ;
      RECT  126.02 42.615 125.69 42.355 ;
      RECT  130.745 42.97 130.415 42.71 ;
      RECT  126.41 43.37 126.08 43.11 ;
      RECT  129.585 42.2 129.315 41.88 ;
      RECT  126.02 34.565 125.69 34.825 ;
      RECT  130.745 34.21 130.415 34.47 ;
      RECT  126.41 33.81 126.08 34.07 ;
      RECT  129.585 34.98 129.315 35.3 ;
      RECT  126.02 28.475 125.69 28.215 ;
      RECT  130.745 28.83 130.415 28.57 ;
      RECT  126.41 29.23 126.08 28.97 ;
      RECT  129.585 28.06 129.315 27.74 ;
      RECT  126.02 20.425 125.69 20.685 ;
      RECT  130.745 20.07 130.415 20.33 ;
      RECT  126.41 19.67 126.08 19.93 ;
      RECT  129.585 20.84 129.315 21.16 ;
      RECT  130.745 42.97 130.415 42.71 ;
      RECT  130.745 34.47 130.415 34.21 ;
      RECT  130.745 28.83 130.415 28.57 ;
      RECT  130.745 20.33 130.415 20.07 ;
      RECT  126.02 42.615 125.69 42.355 ;
      RECT  126.02 34.825 125.69 34.565 ;
      RECT  126.02 28.475 125.69 28.215 ;
      RECT  126.02 20.685 125.69 20.425 ;
      RECT  38.48 3.045 38.81 3.305 ;
      RECT  33.755 2.69 34.085 2.95 ;
      RECT  38.09 2.29 38.42 2.55 ;
      RECT  34.915 3.46 35.185 3.78 ;
      RECT  44.32 3.045 44.65 3.305 ;
      RECT  39.595 2.69 39.925 2.95 ;
      RECT  43.93 2.29 44.26 2.55 ;
      RECT  40.755 3.46 41.025 3.78 ;
      RECT  33.755 2.69 34.085 2.95 ;
      RECT  39.595 2.69 39.925 2.95 ;
      RECT  38.48 3.045 38.81 3.305 ;
      RECT  44.32 3.045 44.65 3.305 ;
   LAYER  m3 ;
      RECT  71.275 95.47 71.765 95.96 ;
      RECT  71.275 58.26 71.765 58.75 ;
      RECT  80.635 95.47 81.125 95.96 ;
      RECT  80.635 58.26 81.125 58.75 ;
      RECT  77.515 58.26 78.005 58.75 ;
      RECT  74.395 58.26 74.885 58.75 ;
      RECT  77.515 95.96 78.005 95.47 ;
      RECT  74.395 95.96 74.885 95.47 ;
      RECT  67.795 76.865 68.285 77.355 ;
      RECT  67.795 59.88 68.285 60.37 ;
      RECT  67.795 91.48 68.285 91.97 ;
      RECT  67.795 65.015 68.285 65.505 ;
      RECT  67.795 78.05 68.285 78.54 ;
      RECT  67.795 85.95 68.285 86.44 ;
      RECT  67.795 62.25 68.285 62.74 ;
      RECT  67.795 87.53 68.285 88.02 ;
      RECT  67.795 75.68 68.285 76.17 ;
      RECT  67.795 93.85 68.285 94.34 ;
      RECT  67.795 79.63 68.285 80.12 ;
      RECT  67.795 68.965 68.285 69.455 ;
      RECT  67.795 92.665 68.285 93.155 ;
      RECT  67.795 89.9 68.285 90.39 ;
      RECT  67.795 67.78 68.285 68.27 ;
      RECT  67.795 80.815 68.285 81.305 ;
      RECT  67.795 70.15 68.285 70.64 ;
      RECT  67.795 83.58 68.285 84.07 ;
      RECT  67.795 61.065 68.285 61.555 ;
      RECT  67.795 82.0 68.285 82.49 ;
      RECT  67.795 74.1 68.285 74.59 ;
      RECT  67.795 63.83 68.285 64.32 ;
      RECT  67.795 71.73 68.285 72.22 ;
      RECT  67.795 66.2 68.285 66.69 ;
      RECT  67.795 72.915 68.285 73.405 ;
      RECT  67.795 84.765 68.285 85.255 ;
      RECT  67.795 88.715 68.285 89.205 ;
      RECT  84.115 83.58 84.605 84.07 ;
      RECT  84.115 84.765 84.605 85.255 ;
      RECT  84.115 88.715 84.605 89.205 ;
      RECT  84.115 92.665 84.605 93.155 ;
      RECT  84.115 80.815 84.605 81.305 ;
      RECT  84.115 65.015 84.605 65.505 ;
      RECT  84.115 82.0 84.605 82.49 ;
      RECT  84.115 63.83 84.605 64.32 ;
      RECT  84.115 76.865 84.605 77.355 ;
      RECT  84.115 75.68 84.605 76.17 ;
      RECT  84.115 66.2 84.605 66.69 ;
      RECT  84.115 85.95 84.605 86.44 ;
      RECT  84.115 87.53 84.605 88.02 ;
      RECT  84.115 70.15 84.605 70.64 ;
      RECT  84.115 71.73 84.605 72.22 ;
      RECT  84.115 68.965 84.605 69.455 ;
      RECT  84.115 72.915 84.605 73.405 ;
      RECT  84.115 67.78 84.605 68.27 ;
      RECT  84.115 93.85 84.605 94.34 ;
      RECT  84.115 91.48 84.605 91.97 ;
      RECT  84.115 59.88 84.605 60.37 ;
      RECT  84.115 79.63 84.605 80.12 ;
      RECT  84.115 62.25 84.605 62.74 ;
      RECT  84.115 61.065 84.605 61.555 ;
      RECT  84.115 78.05 84.605 78.54 ;
      RECT  84.115 89.9 84.605 90.39 ;
      RECT  84.115 74.1 84.605 74.59 ;
      RECT  74.49 95.565 74.79 95.865 ;
      RECT  80.635 58.26 81.125 58.75 ;
      RECT  74.49 58.355 74.79 58.655 ;
      RECT  77.61 58.355 77.91 58.655 ;
      RECT  71.275 58.26 71.765 58.75 ;
      RECT  80.635 95.47 81.125 95.96 ;
      RECT  77.61 95.565 77.91 95.865 ;
      RECT  71.275 95.47 71.765 95.96 ;
      RECT  67.89 93.945 68.19 94.245 ;
      RECT  84.21 83.675 84.51 83.975 ;
      RECT  84.21 82.095 84.51 82.395 ;
      RECT  67.89 86.045 68.19 86.345 ;
      RECT  67.89 79.725 68.19 80.025 ;
      RECT  67.89 66.295 68.19 66.595 ;
      RECT  67.89 83.675 68.19 83.975 ;
      RECT  67.89 75.775 68.19 76.075 ;
      RECT  84.21 91.575 84.51 91.875 ;
      RECT  67.89 82.095 68.19 82.395 ;
      RECT  84.21 86.045 84.51 86.345 ;
      RECT  84.21 71.825 84.51 72.125 ;
      RECT  84.21 65.11 84.51 65.41 ;
      RECT  67.89 67.875 68.19 68.175 ;
      RECT  84.21 89.995 84.51 90.295 ;
      RECT  67.89 89.995 68.19 90.295 ;
      RECT  67.89 73.01 68.19 73.31 ;
      RECT  84.21 92.76 84.51 93.06 ;
      RECT  84.21 69.06 84.51 69.36 ;
      RECT  84.21 78.145 84.51 78.445 ;
      RECT  84.21 87.625 84.51 87.925 ;
      RECT  67.89 70.245 68.19 70.545 ;
      RECT  84.21 61.16 84.51 61.46 ;
      RECT  84.21 63.925 84.51 64.225 ;
      RECT  67.89 80.91 68.19 81.21 ;
      RECT  67.89 74.195 68.19 74.495 ;
      RECT  84.21 70.245 84.51 70.545 ;
      RECT  67.89 87.625 68.19 87.925 ;
      RECT  67.89 65.11 68.19 65.41 ;
      RECT  84.21 74.195 84.51 74.495 ;
      RECT  84.21 76.96 84.51 77.26 ;
      RECT  84.21 84.86 84.51 85.16 ;
      RECT  67.89 61.16 68.19 61.46 ;
      RECT  67.89 76.96 68.19 77.26 ;
      RECT  67.89 63.925 68.19 64.225 ;
      RECT  67.89 69.06 68.19 69.36 ;
      RECT  67.89 88.81 68.19 89.11 ;
      RECT  84.21 93.945 84.51 94.245 ;
      RECT  67.89 78.145 68.19 78.445 ;
      RECT  67.89 62.345 68.19 62.645 ;
      RECT  67.89 84.86 68.19 85.16 ;
      RECT  67.89 59.975 68.19 60.275 ;
      RECT  84.21 62.345 84.51 62.645 ;
      RECT  84.21 67.875 84.51 68.175 ;
      RECT  84.21 75.775 84.51 76.075 ;
      RECT  84.21 73.01 84.51 73.31 ;
      RECT  67.89 91.575 68.19 91.875 ;
      RECT  84.21 88.81 84.51 89.11 ;
      RECT  84.21 80.91 84.51 81.21 ;
      RECT  84.21 79.725 84.51 80.025 ;
      RECT  84.21 59.975 84.51 60.275 ;
      RECT  67.89 71.825 68.19 72.125 ;
      RECT  84.21 66.295 84.51 66.595 ;
      RECT  67.89 92.76 68.19 93.06 ;
      RECT  72.36 55.305 71.87 55.795 ;
      RECT  73.8 55.305 74.29 55.795 ;
      RECT  78.6 55.305 78.11 55.795 ;
      RECT  69.96 52.305 79.32 52.605 ;
      RECT  73.8 55.305 74.29 55.795 ;
      RECT  78.11 55.305 78.6 55.795 ;
      RECT  71.87 55.305 72.36 55.795 ;
      RECT  73.08 50.61 79.32 50.91 ;
      RECT  74.68 45.885 75.17 46.375 ;
      RECT  76.61 45.885 77.1 46.375 ;
      RECT  76.55 41.695 77.04 42.185 ;
      RECT  74.74 41.695 75.23 42.185 ;
      RECT  76.55 40.085 77.04 40.575 ;
      RECT  76.2 49.755 76.69 50.245 ;
      RECT  74.74 40.085 75.23 40.575 ;
      RECT  75.09 49.755 75.58 50.245 ;
      RECT  77.075 29.185 77.565 29.675 ;
      RECT  77.175 33.935 77.665 34.425 ;
      RECT  74.115 33.935 74.605 34.425 ;
      RECT  74.215 29.185 74.705 29.675 ;
      RECT  77.145 31.265 77.635 31.755 ;
      RECT  74.17 36.12 74.66 36.61 ;
      RECT  77.12 36.12 77.61 36.61 ;
      RECT  74.72 32.275 75.21 32.765 ;
      RECT  74.145 31.265 74.635 31.755 ;
      RECT  76.57 32.275 77.06 32.765 ;
      RECT  73.08 50.91 79.32 50.61 ;
      RECT  69.96 52.605 79.32 52.305 ;
      RECT  74.68 46.375 75.17 45.885 ;
      RECT  71.87 55.795 72.36 55.305 ;
      RECT  76.61 46.375 77.1 45.885 ;
      RECT  74.215 29.675 74.705 29.185 ;
      RECT  74.115 34.425 74.605 33.935 ;
      RECT  77.175 34.425 77.665 33.935 ;
      RECT  77.075 29.675 77.565 29.185 ;
      RECT  73.8 55.795 74.29 55.305 ;
      RECT  78.11 55.795 78.6 55.305 ;
      RECT  74.74 42.185 75.23 41.695 ;
      RECT  76.55 42.185 77.04 41.695 ;
      RECT  74.72 32.765 75.21 32.275 ;
      RECT  76.2 50.245 76.69 49.755 ;
      RECT  74.17 36.61 74.66 36.12 ;
      RECT  76.57 32.765 77.06 32.275 ;
      RECT  76.55 40.575 77.04 40.085 ;
      RECT  75.09 50.245 75.58 49.755 ;
      RECT  74.74 40.575 75.23 40.085 ;
      RECT  74.145 31.755 74.635 31.265 ;
      RECT  77.145 31.755 77.635 31.265 ;
      RECT  77.12 36.61 77.61 36.12 ;
      RECT  73.8 98.915 74.29 98.425 ;
      RECT  78.6 98.915 78.11 98.425 ;
      RECT  80.04 98.915 80.53 98.425 ;
      RECT  73.08 101.915 82.44 101.615 ;
      RECT  73.8 98.915 74.29 98.425 ;
      RECT  80.04 98.915 80.53 98.425 ;
      RECT  78.11 98.915 78.6 98.425 ;
      RECT  73.08 103.61 79.32 103.31 ;
      RECT  74.68 108.335 75.17 107.845 ;
      RECT  76.61 108.335 77.1 107.845 ;
      RECT  76.55 112.525 77.04 112.035 ;
      RECT  74.74 112.525 75.23 112.035 ;
      RECT  76.55 114.135 77.04 113.645 ;
      RECT  76.2 104.465 76.69 103.975 ;
      RECT  74.74 114.135 75.23 113.645 ;
      RECT  75.09 104.465 75.58 103.975 ;
      RECT  73.08 103.31 79.32 103.61 ;
      RECT  73.08 101.615 82.44 101.915 ;
      RECT  74.68 107.845 75.17 108.335 ;
      RECT  80.04 98.425 80.53 98.915 ;
      RECT  78.11 98.425 78.6 98.915 ;
      RECT  76.61 107.845 77.1 108.335 ;
      RECT  74.74 112.035 75.23 112.525 ;
      RECT  76.55 112.035 77.04 112.525 ;
      RECT  73.8 98.425 74.29 98.915 ;
      RECT  75.09 103.975 75.58 104.465 ;
      RECT  74.74 113.645 75.23 114.135 ;
      RECT  76.55 113.645 77.04 114.135 ;
      RECT  76.2 103.975 76.69 104.465 ;
      RECT  43.475 63.185 43.965 63.675 ;
      RECT  33.605 63.185 34.095 63.675 ;
      RECT  40.22 67.17 40.71 67.66 ;
      RECT  40.22 63.22 40.71 63.71 ;
      RECT  43.475 67.135 43.965 67.625 ;
      RECT  32.245 63.185 32.735 63.675 ;
      RECT  42.115 63.185 42.605 63.675 ;
      RECT  42.115 67.135 42.605 67.625 ;
      RECT  38.095 63.22 38.585 63.71 ;
      RECT  38.095 67.17 38.585 67.66 ;
      RECT  43.475 75.035 43.965 75.525 ;
      RECT  33.605 75.035 34.095 75.525 ;
      RECT  40.22 79.02 40.71 79.51 ;
      RECT  40.22 75.07 40.71 75.56 ;
      RECT  43.475 78.985 43.965 79.475 ;
      RECT  32.245 75.035 32.735 75.525 ;
      RECT  42.115 75.035 42.605 75.525 ;
      RECT  42.115 78.985 42.605 79.475 ;
      RECT  38.095 75.07 38.585 75.56 ;
      RECT  38.095 79.02 38.585 79.51 ;
      RECT  54.545 75.035 55.035 75.525 ;
      RECT  54.545 73.06 55.035 73.55 ;
      RECT  51.29 79.02 51.78 79.51 ;
      RECT  51.29 75.07 51.78 75.56 ;
      RECT  54.545 65.16 55.035 65.65 ;
      RECT  51.29 90.87 51.78 91.36 ;
      RECT  54.545 88.86 55.035 89.35 ;
      RECT  54.545 84.91 55.035 85.4 ;
      RECT  51.29 85.07 51.78 85.56 ;
      RECT  51.29 82.97 51.78 83.46 ;
      RECT  54.545 90.835 55.035 91.325 ;
      RECT  54.545 67.135 55.035 67.625 ;
      RECT  51.29 67.17 51.78 67.66 ;
      RECT  43.475 63.185 43.965 63.675 ;
      RECT  51.29 77.17 51.78 77.66 ;
      RECT  51.29 86.92 51.78 87.41 ;
      RECT  54.545 71.085 55.035 71.575 ;
      RECT  54.545 63.185 55.035 63.675 ;
      RECT  43.475 67.135 43.965 67.625 ;
      RECT  43.475 78.985 43.965 79.475 ;
      RECT  54.545 86.885 55.035 87.375 ;
      RECT  43.475 75.035 43.965 75.525 ;
      RECT  54.545 77.01 55.035 77.5 ;
      RECT  51.29 63.22 51.78 63.71 ;
      RECT  54.545 82.935 55.035 83.425 ;
      RECT  33.605 63.185 34.095 63.675 ;
      RECT  51.29 73.22 51.78 73.71 ;
      RECT  54.545 78.985 55.035 79.475 ;
      RECT  54.545 80.96 55.035 81.45 ;
      RECT  51.29 89.02 51.78 89.51 ;
      RECT  33.605 75.035 34.095 75.525 ;
      RECT  51.29 69.27 51.78 69.76 ;
      RECT  51.29 71.12 51.78 71.61 ;
      RECT  51.29 65.32 51.78 65.81 ;
      RECT  40.22 67.17 40.71 67.66 ;
      RECT  40.22 75.07 40.71 75.56 ;
      RECT  40.22 79.02 40.71 79.51 ;
      RECT  40.22 63.22 40.71 63.71 ;
      RECT  51.29 81.12 51.78 81.61 ;
      RECT  54.545 69.11 55.035 69.6 ;
      RECT  53.185 67.135 53.675 67.625 ;
      RECT  53.185 84.91 53.675 85.4 ;
      RECT  49.165 75.07 49.655 75.56 ;
      RECT  53.185 73.06 53.675 73.55 ;
      RECT  49.165 69.26 49.655 69.75 ;
      RECT  53.185 86.885 53.675 87.375 ;
      RECT  38.095 79.02 38.585 79.51 ;
      RECT  49.165 82.97 49.655 83.46 ;
      RECT  49.165 77.16 49.655 77.65 ;
      RECT  53.185 80.96 53.675 81.45 ;
      RECT  53.185 82.935 53.675 83.425 ;
      RECT  53.185 77.01 53.675 77.5 ;
      RECT  38.095 67.17 38.585 67.66 ;
      RECT  32.245 75.035 32.735 75.525 ;
      RECT  49.165 90.87 49.655 91.36 ;
      RECT  49.165 73.21 49.655 73.7 ;
      RECT  49.165 67.17 49.655 67.66 ;
      RECT  49.165 85.06 49.655 85.55 ;
      RECT  53.185 78.985 53.675 79.475 ;
      RECT  42.115 78.985 42.605 79.475 ;
      RECT  53.185 63.185 53.675 63.675 ;
      RECT  49.165 86.92 49.655 87.41 ;
      RECT  38.095 63.22 38.585 63.71 ;
      RECT  42.115 75.035 42.605 75.525 ;
      RECT  49.165 89.01 49.655 89.5 ;
      RECT  42.115 63.185 42.605 63.675 ;
      RECT  49.165 79.02 49.655 79.51 ;
      RECT  49.165 63.22 49.655 63.71 ;
      RECT  42.115 67.135 42.605 67.625 ;
      RECT  53.185 75.035 53.675 75.525 ;
      RECT  38.095 75.07 38.585 75.56 ;
      RECT  53.185 90.835 53.675 91.325 ;
      RECT  49.165 81.11 49.655 81.6 ;
      RECT  32.245 63.185 32.735 63.675 ;
      RECT  49.165 65.31 49.655 65.8 ;
      RECT  53.185 88.86 53.675 89.35 ;
      RECT  53.185 69.11 53.675 69.6 ;
      RECT  53.185 65.16 53.675 65.65 ;
      RECT  53.185 71.085 53.675 71.575 ;
      RECT  49.165 71.12 49.655 71.61 ;
      RECT  51.29 82.97 51.78 83.46 ;
      RECT  51.29 86.92 51.78 87.41 ;
      RECT  40.22 63.22 40.71 63.71 ;
      RECT  40.22 67.17 40.71 67.66 ;
      RECT  51.29 81.12 51.78 81.61 ;
      RECT  58.9 76.785 59.39 77.275 ;
      RECT  51.29 90.87 51.78 91.36 ;
      RECT  54.545 71.085 55.035 71.575 ;
      RECT  54.545 86.885 55.035 87.375 ;
      RECT  43.475 67.135 43.965 67.625 ;
      RECT  54.545 69.11 55.035 69.6 ;
      RECT  51.29 77.17 51.78 77.66 ;
      RECT  40.22 75.07 40.71 75.56 ;
      RECT  63.475 76.865 63.965 77.355 ;
      RECT  51.29 73.22 51.78 73.71 ;
      RECT  51.29 85.07 51.78 85.56 ;
      RECT  54.545 73.06 55.035 73.55 ;
      RECT  33.605 75.035 34.095 75.525 ;
      RECT  51.29 89.02 51.78 89.51 ;
      RECT  54.545 77.01 55.035 77.5 ;
      RECT  51.29 67.17 51.78 67.66 ;
      RECT  43.475 63.185 43.965 63.675 ;
      RECT  54.545 75.035 55.035 75.525 ;
      RECT  54.545 84.91 55.035 85.4 ;
      RECT  51.29 79.02 51.78 79.51 ;
      RECT  54.545 88.86 55.035 89.35 ;
      RECT  54.545 78.985 55.035 79.475 ;
      RECT  51.29 75.07 51.78 75.56 ;
      RECT  51.29 65.32 51.78 65.81 ;
      RECT  51.29 63.22 51.78 63.71 ;
      RECT  54.545 82.935 55.035 83.425 ;
      RECT  33.605 63.185 34.095 63.675 ;
      RECT  54.545 80.96 55.035 81.45 ;
      RECT  43.475 75.035 43.965 75.525 ;
      RECT  54.545 65.16 55.035 65.65 ;
      RECT  54.545 90.835 55.035 91.325 ;
      RECT  40.22 79.02 40.71 79.51 ;
      RECT  51.29 69.27 51.78 69.76 ;
      RECT  54.545 63.185 55.035 63.675 ;
      RECT  51.29 71.12 51.78 71.61 ;
      RECT  54.545 67.135 55.035 67.625 ;
      RECT  43.475 78.985 43.965 79.475 ;
      RECT  53.185 69.11 53.675 69.6 ;
      RECT  42.115 75.035 42.605 75.525 ;
      RECT  53.185 90.835 53.675 91.325 ;
      RECT  49.165 67.17 49.655 67.66 ;
      RECT  38.095 79.02 38.585 79.51 ;
      RECT  38.095 63.22 38.585 63.71 ;
      RECT  53.185 78.985 53.675 79.475 ;
      RECT  32.245 75.035 32.735 75.525 ;
      RECT  53.185 63.185 53.675 63.675 ;
      RECT  56.775 76.79 57.265 77.28 ;
      RECT  49.165 79.02 49.655 79.51 ;
      RECT  53.185 75.035 53.675 75.525 ;
      RECT  49.165 85.06 49.655 85.55 ;
      RECT  49.165 82.97 49.655 83.46 ;
      RECT  53.185 71.085 53.675 71.575 ;
      RECT  49.165 89.01 49.655 89.5 ;
      RECT  53.185 77.01 53.675 77.5 ;
      RECT  49.165 90.87 49.655 91.36 ;
      RECT  53.185 84.91 53.675 85.4 ;
      RECT  49.165 81.11 49.655 81.6 ;
      RECT  60.985 76.865 61.475 77.355 ;
      RECT  32.245 63.185 32.735 63.675 ;
      RECT  49.165 63.22 49.655 63.71 ;
      RECT  49.165 65.31 49.655 65.8 ;
      RECT  49.165 69.26 49.655 69.75 ;
      RECT  42.115 67.135 42.605 67.625 ;
      RECT  42.115 63.185 42.605 63.675 ;
      RECT  49.165 86.92 49.655 87.41 ;
      RECT  53.185 73.06 53.675 73.55 ;
      RECT  53.185 88.86 53.675 89.35 ;
      RECT  49.165 71.12 49.655 71.61 ;
      RECT  49.165 75.07 49.655 75.56 ;
      RECT  42.115 78.985 42.605 79.475 ;
      RECT  53.185 67.135 53.675 67.625 ;
      RECT  53.185 65.16 53.675 65.65 ;
      RECT  53.185 82.935 53.675 83.425 ;
      RECT  49.165 73.21 49.655 73.7 ;
      RECT  49.165 77.16 49.655 77.65 ;
      RECT  38.095 75.07 38.585 75.56 ;
      RECT  53.185 80.96 53.675 81.45 ;
      RECT  38.095 67.17 38.585 67.66 ;
      RECT  53.185 86.885 53.675 87.375 ;
      RECT  108.925 63.185 108.435 63.675 ;
      RECT  118.795 63.185 118.305 63.675 ;
      RECT  112.18 67.17 111.69 67.66 ;
      RECT  112.18 63.22 111.69 63.71 ;
      RECT  108.925 67.135 108.435 67.625 ;
      RECT  120.155 63.185 119.665 63.675 ;
      RECT  110.285 63.185 109.795 63.675 ;
      RECT  110.285 67.135 109.795 67.625 ;
      RECT  114.305 63.22 113.815 63.71 ;
      RECT  114.305 67.17 113.815 67.66 ;
      RECT  108.925 75.035 108.435 75.525 ;
      RECT  118.795 75.035 118.305 75.525 ;
      RECT  112.18 79.02 111.69 79.51 ;
      RECT  112.18 75.07 111.69 75.56 ;
      RECT  108.925 78.985 108.435 79.475 ;
      RECT  120.155 75.035 119.665 75.525 ;
      RECT  110.285 75.035 109.795 75.525 ;
      RECT  110.285 78.985 109.795 79.475 ;
      RECT  114.305 75.07 113.815 75.56 ;
      RECT  114.305 79.02 113.815 79.51 ;
      RECT  97.855 75.035 97.365 75.525 ;
      RECT  97.855 73.06 97.365 73.55 ;
      RECT  101.11 79.02 100.62 79.51 ;
      RECT  101.11 75.07 100.62 75.56 ;
      RECT  97.855 65.16 97.365 65.65 ;
      RECT  101.11 90.87 100.62 91.36 ;
      RECT  97.855 88.86 97.365 89.35 ;
      RECT  97.855 84.91 97.365 85.4 ;
      RECT  101.11 85.07 100.62 85.56 ;
      RECT  101.11 82.97 100.62 83.46 ;
      RECT  97.855 90.835 97.365 91.325 ;
      RECT  97.855 67.135 97.365 67.625 ;
      RECT  101.11 67.17 100.62 67.66 ;
      RECT  108.925 63.185 108.435 63.675 ;
      RECT  101.11 77.17 100.62 77.66 ;
      RECT  101.11 86.92 100.62 87.41 ;
      RECT  97.855 71.085 97.365 71.575 ;
      RECT  97.855 63.185 97.365 63.675 ;
      RECT  108.925 67.135 108.435 67.625 ;
      RECT  108.925 78.985 108.435 79.475 ;
      RECT  97.855 86.885 97.365 87.375 ;
      RECT  108.925 75.035 108.435 75.525 ;
      RECT  97.855 77.01 97.365 77.5 ;
      RECT  101.11 63.22 100.62 63.71 ;
      RECT  97.855 82.935 97.365 83.425 ;
      RECT  118.795 63.185 118.305 63.675 ;
      RECT  101.11 73.22 100.62 73.71 ;
      RECT  97.855 78.985 97.365 79.475 ;
      RECT  97.855 80.96 97.365 81.45 ;
      RECT  101.11 89.02 100.62 89.51 ;
      RECT  118.795 75.035 118.305 75.525 ;
      RECT  101.11 69.27 100.62 69.76 ;
      RECT  101.11 71.12 100.62 71.61 ;
      RECT  101.11 65.32 100.62 65.81 ;
      RECT  112.18 67.17 111.69 67.66 ;
      RECT  112.18 75.07 111.69 75.56 ;
      RECT  112.18 79.02 111.69 79.51 ;
      RECT  112.18 63.22 111.69 63.71 ;
      RECT  101.11 81.12 100.62 81.61 ;
      RECT  97.855 69.11 97.365 69.6 ;
      RECT  99.215 67.135 98.725 67.625 ;
      RECT  99.215 84.91 98.725 85.4 ;
      RECT  103.235 75.07 102.745 75.56 ;
      RECT  99.215 73.06 98.725 73.55 ;
      RECT  103.235 69.26 102.745 69.75 ;
      RECT  99.215 86.885 98.725 87.375 ;
      RECT  114.305 79.02 113.815 79.51 ;
      RECT  103.235 82.97 102.745 83.46 ;
      RECT  103.235 77.16 102.745 77.65 ;
      RECT  99.215 80.96 98.725 81.45 ;
      RECT  99.215 82.935 98.725 83.425 ;
      RECT  99.215 77.01 98.725 77.5 ;
      RECT  114.305 67.17 113.815 67.66 ;
      RECT  120.155 75.035 119.665 75.525 ;
      RECT  103.235 90.87 102.745 91.36 ;
      RECT  103.235 73.21 102.745 73.7 ;
      RECT  103.235 67.17 102.745 67.66 ;
      RECT  103.235 85.06 102.745 85.55 ;
      RECT  99.215 78.985 98.725 79.475 ;
      RECT  110.285 78.985 109.795 79.475 ;
      RECT  99.215 63.185 98.725 63.675 ;
      RECT  103.235 86.92 102.745 87.41 ;
      RECT  114.305 63.22 113.815 63.71 ;
      RECT  110.285 75.035 109.795 75.525 ;
      RECT  103.235 89.01 102.745 89.5 ;
      RECT  110.285 63.185 109.795 63.675 ;
      RECT  103.235 79.02 102.745 79.51 ;
      RECT  103.235 63.22 102.745 63.71 ;
      RECT  110.285 67.135 109.795 67.625 ;
      RECT  99.215 75.035 98.725 75.525 ;
      RECT  114.305 75.07 113.815 75.56 ;
      RECT  99.215 90.835 98.725 91.325 ;
      RECT  103.235 81.11 102.745 81.6 ;
      RECT  120.155 63.185 119.665 63.675 ;
      RECT  103.235 65.31 102.745 65.8 ;
      RECT  99.215 88.86 98.725 89.35 ;
      RECT  99.215 69.11 98.725 69.6 ;
      RECT  99.215 65.16 98.725 65.65 ;
      RECT  99.215 71.085 98.725 71.575 ;
      RECT  103.235 71.12 102.745 71.61 ;
      RECT  101.11 82.97 100.62 83.46 ;
      RECT  101.11 86.92 100.62 87.41 ;
      RECT  112.18 63.22 111.69 63.71 ;
      RECT  112.18 67.17 111.69 67.66 ;
      RECT  101.11 81.12 100.62 81.61 ;
      RECT  93.5 76.785 93.01 77.275 ;
      RECT  101.11 90.87 100.62 91.36 ;
      RECT  97.855 71.085 97.365 71.575 ;
      RECT  97.855 86.885 97.365 87.375 ;
      RECT  108.925 67.135 108.435 67.625 ;
      RECT  97.855 69.11 97.365 69.6 ;
      RECT  101.11 77.17 100.62 77.66 ;
      RECT  112.18 75.07 111.69 75.56 ;
      RECT  88.925 76.865 88.435 77.355 ;
      RECT  101.11 73.22 100.62 73.71 ;
      RECT  101.11 85.07 100.62 85.56 ;
      RECT  97.855 73.06 97.365 73.55 ;
      RECT  118.795 75.035 118.305 75.525 ;
      RECT  101.11 89.02 100.62 89.51 ;
      RECT  97.855 77.01 97.365 77.5 ;
      RECT  101.11 67.17 100.62 67.66 ;
      RECT  108.925 63.185 108.435 63.675 ;
      RECT  97.855 75.035 97.365 75.525 ;
      RECT  97.855 84.91 97.365 85.4 ;
      RECT  101.11 79.02 100.62 79.51 ;
      RECT  97.855 88.86 97.365 89.35 ;
      RECT  97.855 78.985 97.365 79.475 ;
      RECT  101.11 75.07 100.62 75.56 ;
      RECT  101.11 65.32 100.62 65.81 ;
      RECT  101.11 63.22 100.62 63.71 ;
      RECT  97.855 82.935 97.365 83.425 ;
      RECT  118.795 63.185 118.305 63.675 ;
      RECT  97.855 80.96 97.365 81.45 ;
      RECT  108.925 75.035 108.435 75.525 ;
      RECT  97.855 65.16 97.365 65.65 ;
      RECT  97.855 90.835 97.365 91.325 ;
      RECT  112.18 79.02 111.69 79.51 ;
      RECT  101.11 69.27 100.62 69.76 ;
      RECT  97.855 63.185 97.365 63.675 ;
      RECT  101.11 71.12 100.62 71.61 ;
      RECT  97.855 67.135 97.365 67.625 ;
      RECT  108.925 78.985 108.435 79.475 ;
      RECT  99.215 69.11 98.725 69.6 ;
      RECT  110.285 75.035 109.795 75.525 ;
      RECT  99.215 90.835 98.725 91.325 ;
      RECT  103.235 67.17 102.745 67.66 ;
      RECT  114.305 79.02 113.815 79.51 ;
      RECT  114.305 63.22 113.815 63.71 ;
      RECT  99.215 78.985 98.725 79.475 ;
      RECT  120.155 75.035 119.665 75.525 ;
      RECT  99.215 63.185 98.725 63.675 ;
      RECT  95.625 76.79 95.135 77.28 ;
      RECT  103.235 79.02 102.745 79.51 ;
      RECT  99.215 75.035 98.725 75.525 ;
      RECT  103.235 85.06 102.745 85.55 ;
      RECT  103.235 82.97 102.745 83.46 ;
      RECT  99.215 71.085 98.725 71.575 ;
      RECT  103.235 89.01 102.745 89.5 ;
      RECT  99.215 77.01 98.725 77.5 ;
      RECT  103.235 90.87 102.745 91.36 ;
      RECT  99.215 84.91 98.725 85.4 ;
      RECT  103.235 81.11 102.745 81.6 ;
      RECT  91.415 76.865 90.925 77.355 ;
      RECT  120.155 63.185 119.665 63.675 ;
      RECT  103.235 63.22 102.745 63.71 ;
      RECT  103.235 65.31 102.745 65.8 ;
      RECT  103.235 69.26 102.745 69.75 ;
      RECT  110.285 67.135 109.795 67.625 ;
      RECT  110.285 63.185 109.795 63.675 ;
      RECT  103.235 86.92 102.745 87.41 ;
      RECT  99.215 73.06 98.725 73.55 ;
      RECT  99.215 88.86 98.725 89.35 ;
      RECT  103.235 71.12 102.745 71.61 ;
      RECT  103.235 75.07 102.745 75.56 ;
      RECT  110.285 78.985 109.795 79.475 ;
      RECT  99.215 67.135 98.725 67.625 ;
      RECT  99.215 65.16 98.725 65.65 ;
      RECT  99.215 82.935 98.725 83.425 ;
      RECT  103.235 73.21 102.745 73.7 ;
      RECT  103.235 77.16 102.745 77.65 ;
      RECT  114.305 75.07 113.815 75.56 ;
      RECT  99.215 80.96 98.725 81.45 ;
      RECT  114.305 67.17 113.815 67.66 ;
      RECT  99.215 86.885 98.725 87.375 ;
      RECT  74.49 95.565 74.79 95.865 ;
      RECT  80.04 98.425 80.53 98.915 ;
      RECT  54.545 67.135 55.035 67.625 ;
      RECT  77.075 29.185 77.565 29.675 ;
      RECT  118.305 75.035 118.795 75.525 ;
      RECT  54.545 75.035 55.035 75.525 ;
      RECT  74.68 107.845 75.17 108.335 ;
      RECT  111.69 67.17 112.18 67.66 ;
      RECT  100.62 75.07 101.11 75.56 ;
      RECT  54.545 65.16 55.035 65.65 ;
      RECT  97.365 86.885 97.855 87.375 ;
      RECT  108.435 63.185 108.925 63.675 ;
      RECT  54.545 78.985 55.035 79.475 ;
      RECT  51.29 89.02 51.78 89.51 ;
      RECT  74.68 45.885 75.17 46.375 ;
      RECT  33.605 75.035 34.095 75.525 ;
      RECT  100.62 86.92 101.11 87.41 ;
      RECT  97.365 67.135 97.855 67.625 ;
      RECT  71.275 58.26 71.765 58.75 ;
      RECT  71.87 55.305 72.36 55.795 ;
      RECT  71.275 95.47 71.765 95.96 ;
      RECT  40.22 79.02 40.71 79.51 ;
      RECT  97.365 82.935 97.855 83.425 ;
      RECT  74.74 41.695 75.23 42.185 ;
      RECT  97.365 80.96 97.855 81.45 ;
      RECT  100.62 85.07 101.11 85.56 ;
      RECT  88.435 76.865 88.925 77.355 ;
      RECT  97.365 71.085 97.855 71.575 ;
      RECT  97.365 90.835 97.855 91.325 ;
      RECT  63.475 76.865 63.965 77.355 ;
      RECT  54.545 82.935 55.035 83.425 ;
      RECT  76.61 45.885 77.1 46.375 ;
      RECT  51.29 63.22 51.78 63.71 ;
      RECT  51.29 69.27 51.78 69.76 ;
      RECT  51.29 86.92 51.78 87.41 ;
      RECT  51.29 81.12 51.78 81.61 ;
      RECT  100.62 89.02 101.11 89.51 ;
      RECT  97.365 75.035 97.855 75.525 ;
      RECT  54.545 69.11 55.035 69.6 ;
      RECT  100.62 81.12 101.11 81.61 ;
      RECT  54.545 84.91 55.035 85.4 ;
      RECT  77.61 58.355 77.91 58.655 ;
      RECT  97.365 78.985 97.855 79.475 ;
      RECT  73.8 55.305 74.29 55.795 ;
      RECT  80.635 95.47 81.125 95.96 ;
      RECT  97.365 73.06 97.855 73.55 ;
      RECT  100.62 67.17 101.11 67.66 ;
      RECT  97.365 69.11 97.855 69.6 ;
      RECT  100.62 77.17 101.11 77.66 ;
      RECT  76.55 112.035 77.04 112.525 ;
      RECT  40.22 75.07 40.71 75.56 ;
      RECT  51.29 67.17 51.78 67.66 ;
      RECT  100.62 79.02 101.11 79.51 ;
      RECT  74.115 33.935 74.605 34.425 ;
      RECT  58.9 76.785 59.39 77.275 ;
      RECT  118.305 63.185 118.795 63.675 ;
      RECT  51.29 90.87 51.78 91.36 ;
      RECT  33.605 63.185 34.095 63.675 ;
      RECT  74.74 112.035 75.23 112.525 ;
      RECT  77.175 33.935 77.665 34.425 ;
      RECT  51.29 75.07 51.78 75.56 ;
      RECT  73.8 98.425 74.29 98.915 ;
      RECT  111.69 75.07 112.18 75.56 ;
      RECT  51.29 77.17 51.78 77.66 ;
      RECT  97.365 88.86 97.855 89.35 ;
      RECT  54.545 63.185 55.035 63.675 ;
      RECT  76.55 41.695 77.04 42.185 ;
      RECT  43.475 78.985 43.965 79.475 ;
      RECT  54.545 77.01 55.035 77.5 ;
      RECT  100.62 71.12 101.11 71.61 ;
      RECT  43.475 63.185 43.965 63.675 ;
      RECT  100.62 65.32 101.11 65.81 ;
      RECT  108.435 78.985 108.925 79.475 ;
      RECT  77.61 95.565 77.91 95.865 ;
      RECT  54.545 90.835 55.035 91.325 ;
      RECT  51.29 85.07 51.78 85.56 ;
      RECT  100.62 69.27 101.11 69.76 ;
      RECT  51.29 82.97 51.78 83.46 ;
      RECT  43.475 67.135 43.965 67.625 ;
      RECT  76.61 107.845 77.1 108.335 ;
      RECT  51.29 73.22 51.78 73.71 ;
      RECT  100.62 63.22 101.11 63.71 ;
      RECT  108.435 75.035 108.925 75.525 ;
      RECT  97.365 77.01 97.855 77.5 ;
      RECT  80.635 58.26 81.125 58.75 ;
      RECT  54.545 73.06 55.035 73.55 ;
      RECT  100.62 90.87 101.11 91.36 ;
      RECT  43.475 75.035 43.965 75.525 ;
      RECT  51.29 79.02 51.78 79.51 ;
      RECT  100.62 73.22 101.11 73.71 ;
      RECT  54.545 86.885 55.035 87.375 ;
      RECT  97.365 65.16 97.855 65.65 ;
      RECT  111.69 63.22 112.18 63.71 ;
      RECT  54.545 80.96 55.035 81.45 ;
      RECT  93.01 76.785 93.5 77.275 ;
      RECT  74.49 58.355 74.79 58.655 ;
      RECT  78.11 98.425 78.6 98.915 ;
      RECT  74.215 29.185 74.705 29.675 ;
      RECT  51.29 71.12 51.78 71.61 ;
      RECT  51.29 65.32 51.78 65.81 ;
      RECT  100.62 82.97 101.11 83.46 ;
      RECT  78.11 55.305 78.6 55.795 ;
      RECT  97.365 84.91 97.855 85.4 ;
      RECT  54.545 88.86 55.035 89.35 ;
      RECT  97.365 63.185 97.855 63.675 ;
      RECT  111.69 79.02 112.18 79.51 ;
      RECT  54.545 71.085 55.035 71.575 ;
      RECT  108.435 67.135 108.925 67.625 ;
      RECT  40.22 67.17 40.71 67.66 ;
      RECT  40.22 63.22 40.71 63.71 ;
      RECT  67.89 93.945 68.19 94.245 ;
      RECT  109.795 67.135 110.285 67.625 ;
      RECT  113.815 67.17 114.305 67.66 ;
      RECT  109.795 63.185 110.285 63.675 ;
      RECT  53.185 84.91 53.675 85.4 ;
      RECT  102.745 89.01 103.235 89.5 ;
      RECT  84.21 83.675 84.51 83.975 ;
      RECT  102.745 75.07 103.235 75.56 ;
      RECT  98.725 80.96 99.215 81.45 ;
      RECT  84.21 82.095 84.51 82.395 ;
      RECT  53.185 80.96 53.675 81.45 ;
      RECT  49.165 71.12 49.655 71.61 ;
      RECT  53.185 67.135 53.675 67.625 ;
      RECT  49.165 89.01 49.655 89.5 ;
      RECT  67.89 86.045 68.19 86.345 ;
      RECT  98.725 65.16 99.215 65.65 ;
      RECT  98.725 73.06 99.215 73.55 ;
      RECT  67.89 79.725 68.19 80.025 ;
      RECT  67.89 66.295 68.19 66.595 ;
      RECT  76.55 113.645 77.04 114.135 ;
      RECT  119.665 75.035 120.155 75.525 ;
      RECT  67.89 83.675 68.19 83.975 ;
      RECT  67.89 75.775 68.19 76.075 ;
      RECT  84.21 91.575 84.51 91.875 ;
      RECT  98.725 77.01 99.215 77.5 ;
      RECT  74.74 113.645 75.23 114.135 ;
      RECT  67.89 82.095 68.19 82.395 ;
      RECT  76.2 103.975 76.69 104.465 ;
      RECT  98.725 82.935 99.215 83.425 ;
      RECT  49.165 63.22 49.655 63.71 ;
      RECT  84.21 86.045 84.51 86.345 ;
      RECT  90.925 76.865 91.415 77.355 ;
      RECT  84.21 71.825 84.51 72.125 ;
      RECT  49.165 77.16 49.655 77.65 ;
      RECT  67.89 67.875 68.19 68.175 ;
      RECT  84.21 65.11 84.51 65.41 ;
      RECT  102.745 86.92 103.235 87.41 ;
      RECT  53.185 77.01 53.675 77.5 ;
      RECT  98.725 78.985 99.215 79.475 ;
      RECT  84.21 89.995 84.51 90.295 ;
      RECT  67.89 89.995 68.19 90.295 ;
      RECT  67.89 73.01 68.19 73.31 ;
      RECT  84.21 92.76 84.51 93.06 ;
      RECT  84.21 69.06 84.51 69.36 ;
      RECT  84.21 78.145 84.51 78.445 ;
      RECT  102.745 79.02 103.235 79.51 ;
      RECT  113.815 79.02 114.305 79.51 ;
      RECT  84.21 87.625 84.51 87.925 ;
      RECT  77.145 31.265 77.635 31.755 ;
      RECT  53.185 63.185 53.675 63.675 ;
      RECT  38.095 75.07 38.585 75.56 ;
      RECT  109.795 75.035 110.285 75.525 ;
      RECT  49.165 81.11 49.655 81.6 ;
      RECT  67.89 70.245 68.19 70.545 ;
      RECT  84.21 61.16 84.51 61.46 ;
      RECT  102.745 82.97 103.235 83.46 ;
      RECT  32.245 75.035 32.735 75.525 ;
      RECT  38.095 67.17 38.585 67.66 ;
      RECT  84.21 63.925 84.51 64.225 ;
      RECT  74.72 32.275 75.21 32.765 ;
      RECT  113.815 75.07 114.305 75.56 ;
      RECT  53.185 82.935 53.675 83.425 ;
      RECT  98.725 75.035 99.215 75.525 ;
      RECT  49.165 82.97 49.655 83.46 ;
      RECT  67.89 80.91 68.19 81.21 ;
      RECT  67.89 74.195 68.19 74.495 ;
      RECT  98.725 90.835 99.215 91.325 ;
      RECT  53.185 71.085 53.675 71.575 ;
      RECT  42.115 75.035 42.605 75.525 ;
      RECT  102.745 71.12 103.235 71.61 ;
      RECT  84.21 70.245 84.51 70.545 ;
      RECT  98.725 86.885 99.215 87.375 ;
      RECT  67.89 87.625 68.19 87.925 ;
      RECT  67.89 65.11 68.19 65.41 ;
      RECT  95.135 76.79 95.625 77.28 ;
      RECT  49.165 67.17 49.655 67.66 ;
      RECT  102.745 65.31 103.235 65.8 ;
      RECT  49.165 65.31 49.655 65.8 ;
      RECT  53.185 65.16 53.675 65.65 ;
      RECT  84.21 74.195 84.51 74.495 ;
      RECT  84.21 76.96 84.51 77.26 ;
      RECT  84.21 84.86 84.51 85.16 ;
      RECT  98.725 63.185 99.215 63.675 ;
      RECT  42.115 63.185 42.605 63.675 ;
      RECT  67.89 61.16 68.19 61.46 ;
      RECT  67.89 76.96 68.19 77.26 ;
      RECT  38.095 79.02 38.585 79.51 ;
      RECT  38.095 63.22 38.585 63.71 ;
      RECT  53.185 78.985 53.675 79.475 ;
      RECT  102.745 63.22 103.235 63.71 ;
      RECT  67.89 63.925 68.19 64.225 ;
      RECT  53.185 73.06 53.675 73.55 ;
      RECT  98.725 88.86 99.215 89.35 ;
      RECT  119.665 63.185 120.155 63.675 ;
      RECT  67.89 69.06 68.19 69.36 ;
      RECT  113.815 63.22 114.305 63.71 ;
      RECT  102.745 85.06 103.235 85.55 ;
      RECT  53.185 69.11 53.675 69.6 ;
      RECT  49.165 85.06 49.655 85.55 ;
      RECT  76.2 49.755 76.69 50.245 ;
      RECT  67.89 88.81 68.19 89.11 ;
      RECT  98.725 71.085 99.215 71.575 ;
      RECT  49.165 90.87 49.655 91.36 ;
      RECT  102.745 69.26 103.235 69.75 ;
      RECT  42.115 78.985 42.605 79.475 ;
      RECT  102.745 81.11 103.235 81.6 ;
      RECT  98.725 69.11 99.215 69.6 ;
      RECT  53.185 90.835 53.675 91.325 ;
      RECT  109.795 78.985 110.285 79.475 ;
      RECT  84.21 93.945 84.51 94.245 ;
      RECT  49.165 86.92 49.655 87.41 ;
      RECT  77.12 36.12 77.61 36.61 ;
      RECT  74.17 36.12 74.66 36.61 ;
      RECT  67.89 78.145 68.19 78.445 ;
      RECT  49.165 73.21 49.655 73.7 ;
      RECT  98.725 67.135 99.215 67.625 ;
      RECT  67.89 62.345 68.19 62.645 ;
      RECT  32.245 63.185 32.735 63.675 ;
      RECT  67.89 84.86 68.19 85.16 ;
      RECT  67.89 59.975 68.19 60.275 ;
      RECT  84.21 62.345 84.51 62.645 ;
      RECT  84.21 67.875 84.51 68.175 ;
      RECT  75.09 49.755 75.58 50.245 ;
      RECT  42.115 67.135 42.605 67.625 ;
      RECT  53.185 75.035 53.675 75.525 ;
      RECT  76.55 40.085 77.04 40.575 ;
      RECT  76.57 32.275 77.06 32.765 ;
      RECT  49.165 75.07 49.655 75.56 ;
      RECT  56.775 76.79 57.265 77.28 ;
      RECT  102.745 77.16 103.235 77.65 ;
      RECT  84.21 75.775 84.51 76.075 ;
      RECT  84.21 73.01 84.51 73.31 ;
      RECT  53.185 86.885 53.675 87.375 ;
      RECT  53.185 88.86 53.675 89.35 ;
      RECT  98.725 84.91 99.215 85.4 ;
      RECT  74.145 31.265 74.635 31.755 ;
      RECT  49.165 69.26 49.655 69.75 ;
      RECT  75.09 103.975 75.58 104.465 ;
      RECT  49.165 79.02 49.655 79.51 ;
      RECT  67.89 91.575 68.19 91.875 ;
      RECT  84.21 88.81 84.51 89.11 ;
      RECT  84.21 80.91 84.51 81.21 ;
      RECT  102.745 67.17 103.235 67.66 ;
      RECT  102.745 73.21 103.235 73.7 ;
      RECT  102.745 90.87 103.235 91.36 ;
      RECT  84.21 79.725 84.51 80.025 ;
      RECT  84.21 59.975 84.51 60.275 ;
      RECT  74.74 40.085 75.23 40.575 ;
      RECT  67.89 71.825 68.19 72.125 ;
      RECT  84.21 66.295 84.51 66.595 ;
      RECT  60.985 76.865 61.475 77.355 ;
      RECT  67.89 92.76 68.19 93.06 ;
      RECT  -0.245 6.825 0.245 7.315 ;
      RECT  -0.245 -0.255 0.245 0.235 ;
      RECT  -0.245 13.905 0.245 14.395 ;
      RECT  6.165 96.315 5.675 96.805 ;
      RECT  6.165 107.515 5.675 108.005 ;
      RECT  6.165 85.115 5.675 85.605 ;
      RECT  2.485 73.915 1.995 74.405 ;
      RECT  2.485 73.915 1.995 74.405 ;
      RECT  2.485 85.115 1.995 85.605 ;
      RECT  2.485 96.315 1.995 96.805 ;
      RECT  2.485 107.515 1.995 108.005 ;
      RECT  2.485 62.715 1.995 63.205 ;
      RECT  2.485 62.715 1.995 63.205 ;
      RECT  6.165 73.915 5.675 74.405 ;
      RECT  6.165 73.915 5.675 74.405 ;
      RECT  6.165 62.715 5.675 63.205 ;
      RECT  6.165 62.715 5.675 63.205 ;
      RECT  6.165 79.515 5.675 80.005 ;
      RECT  2.485 90.715 1.995 91.205 ;
      RECT  6.165 90.715 5.675 91.205 ;
      RECT  6.165 68.315 5.675 68.805 ;
      RECT  2.485 79.515 1.995 80.005 ;
      RECT  2.485 57.115 1.995 57.605 ;
      RECT  2.485 68.315 1.995 68.805 ;
      RECT  2.485 101.915 1.995 102.405 ;
      RECT  6.165 101.915 5.675 102.405 ;
      RECT  6.165 57.115 5.675 57.605 ;
      RECT  5.675 96.315 6.165 96.805 ;
      RECT  -0.245 6.825 0.245 7.315 ;
      RECT  1.995 96.315 2.485 96.805 ;
      RECT  26.565 20.965 27.055 21.455 ;
      RECT  26.565 35.105 27.055 35.595 ;
      RECT  1.995 85.115 2.485 85.605 ;
      RECT  1.995 62.715 2.485 63.205 ;
      RECT  26.565 6.825 27.055 7.315 ;
      RECT  5.675 73.915 6.165 74.405 ;
      RECT  5.675 62.715 6.165 63.205 ;
      RECT  5.675 107.515 6.165 108.005 ;
      RECT  5.675 85.115 6.165 85.605 ;
      RECT  1.995 73.915 2.485 74.405 ;
      RECT  26.565 49.245 27.055 49.735 ;
      RECT  1.995 107.515 2.485 108.005 ;
      RECT  26.565 28.035 27.055 28.525 ;
      RECT  26.565 -0.245 27.055 0.245 ;
      RECT  1.995 101.915 2.485 102.405 ;
      RECT  -0.245 -0.255 0.245 0.235 ;
      RECT  1.995 68.315 2.485 68.805 ;
      RECT  5.675 101.915 6.165 102.405 ;
      RECT  1.995 90.715 2.485 91.205 ;
      RECT  5.675 57.115 6.165 57.605 ;
      RECT  26.565 13.895 27.055 14.385 ;
      RECT  5.675 79.515 6.165 80.005 ;
      RECT  1.995 79.515 2.485 80.005 ;
      RECT  1.995 57.115 2.485 57.605 ;
      RECT  -0.245 13.905 0.245 14.395 ;
      RECT  26.565 42.175 27.055 42.665 ;
      RECT  5.675 68.315 6.165 68.805 ;
      RECT  5.675 90.715 6.165 91.205 ;
      RECT  26.565 56.315 27.055 56.805 ;
      RECT  151.535 133.255 151.045 132.765 ;
      RECT  151.535 140.335 151.045 139.845 ;
      RECT  145.125 57.905 145.615 57.415 ;
      RECT  145.125 46.705 145.615 46.215 ;
      RECT  145.125 69.105 145.615 68.615 ;
      RECT  148.805 80.305 149.295 79.815 ;
      RECT  148.805 80.305 149.295 79.815 ;
      RECT  148.805 69.105 149.295 68.615 ;
      RECT  148.805 57.905 149.295 57.415 ;
      RECT  148.805 46.705 149.295 46.215 ;
      RECT  148.805 91.505 149.295 91.015 ;
      RECT  148.805 91.505 149.295 91.015 ;
      RECT  145.125 80.305 145.615 79.815 ;
      RECT  145.125 80.305 145.615 79.815 ;
      RECT  145.125 91.505 145.615 91.015 ;
      RECT  145.125 91.505 145.615 91.015 ;
      RECT  145.125 74.705 145.615 74.215 ;
      RECT  148.805 63.505 149.295 63.015 ;
      RECT  145.125 63.505 145.615 63.015 ;
      RECT  145.125 85.905 145.615 85.415 ;
      RECT  148.805 74.705 149.295 74.215 ;
      RECT  148.805 97.105 149.295 96.615 ;
      RECT  148.805 85.905 149.295 85.415 ;
      RECT  148.805 52.305 149.295 51.815 ;
      RECT  145.125 52.305 145.615 51.815 ;
      RECT  145.125 97.105 145.615 96.615 ;
      RECT  126.255 104.975 125.765 104.485 ;
      RECT  151.535 133.255 151.045 132.765 ;
      RECT  145.615 69.105 145.125 68.615 ;
      RECT  149.295 46.705 148.805 46.215 ;
      RECT  145.615 80.305 145.125 79.815 ;
      RECT  145.615 57.905 145.125 57.415 ;
      RECT  126.255 119.115 125.765 118.625 ;
      RECT  149.295 57.905 148.805 57.415 ;
      RECT  149.295 91.505 148.805 91.015 ;
      RECT  145.615 91.505 145.125 91.015 ;
      RECT  149.295 80.305 148.805 79.815 ;
      RECT  149.295 69.105 148.805 68.615 ;
      RECT  126.255 133.255 125.765 132.765 ;
      RECT  145.615 46.705 145.125 46.215 ;
      RECT  145.615 63.505 145.125 63.015 ;
      RECT  149.295 52.305 148.805 51.815 ;
      RECT  145.615 74.705 145.125 74.215 ;
      RECT  149.295 63.505 148.805 63.015 ;
      RECT  145.615 52.305 145.125 51.815 ;
      RECT  149.295 97.105 148.805 96.615 ;
      RECT  151.535 140.335 151.045 139.845 ;
      RECT  149.295 85.905 148.805 85.415 ;
      RECT  149.295 74.705 148.805 74.215 ;
      RECT  126.255 126.185 125.765 125.695 ;
      RECT  126.255 97.905 125.765 97.415 ;
      RECT  126.255 140.325 125.765 139.835 ;
      RECT  126.255 112.045 125.765 111.555 ;
      RECT  145.615 97.105 145.125 96.615 ;
      RECT  145.615 85.905 145.125 85.415 ;
      RECT  21.39 109.95 27.23 110.25 ;
      RECT  24.065 129.525 24.555 130.015 ;
      RECT  24.065 115.385 24.555 115.875 ;
      RECT  24.065 136.595 24.555 137.085 ;
      RECT  24.065 122.455 24.555 122.945 ;
      RECT  24.065 108.315 24.555 108.805 ;
      RECT  131.43 44.27 125.59 43.97 ;
      RECT  128.755 24.695 128.265 24.205 ;
      RECT  128.755 38.835 128.265 38.345 ;
      RECT  128.755 17.625 128.265 17.135 ;
      RECT  128.755 31.765 128.265 31.275 ;
      RECT  128.755 45.905 128.265 45.415 ;
      RECT  33.07 1.39 44.75 1.69 ;
      RECT  41.585 6.825 42.075 7.315 ;
      RECT  35.745 6.825 36.235 7.315 ;
      RECT  41.585 -0.245 42.075 0.245 ;
      RECT  35.745 -0.245 36.235 0.245 ;
   LAYER  m4 ;
   END
   END    sram_2_16_sky130
END    LIBRARY
