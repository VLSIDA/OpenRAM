* SPICE3 file created from cell_6t.ext - technology: scmos

M1000 a_36_40# a_28_32# vdd vdd pfet w=0.6u l=0.8u
+  ad=0.76p pd=3.6u as=2p ps=8.8u
M1001 vdd a_36_40# a_28_32# vdd pfet w=0.6u l=0.8u
+  ad=0p pd=0u as=0.76p ps=3.6u
M1002 a_36_40# a_28_32# gnd gnd nfet w=1.6u l=0.4u
+  ad=2.4p pd=7.2u as=4.48p ps=12u
M1003 gnd a_36_40# a_28_32# gnd nfet w=1.6u l=0.4u
+  ad=0p pd=0u as=2.4p ps=7.2u
M1004 a_36_40# wl bl gnd nfet w=0.8u l=0.4u
+  ad=0p pd=0u as=0.8p ps=3.6u
M1005 a_28_32# wl br gnd nfet w=0.8u l=0.4u
+  ad=0p pd=0u as=0.8p ps=3.6u
C0 vdd 0 2.60fF
