magic
tech sky130A
magscale 1 2
timestamp 1595931502
<< checkpaint >>
rect -1216 -1260 2348 1750
<< nwell >>
rect 380 0 1088 490
<< poly >>
rect 77 182 136 212
rect 336 182 408 212
<< locali >>
rect 60 164 94 230
rect 203 130 1070 164
<< metal1 >>
rect 222 0 250 395
rect 720 0 748 395
use pmos_m1_w3_000_sli_dli_da_p  pmos_m1_w3_000_sli_dli_da_p_0
timestamp 1595931502
transform 0 1 434 -1 0 272
box -59 -54 209 654
use nmos_m1_w0_740_sli_dli_da_p  nmos_m1_w0_740_sli_dli_da_p_0
timestamp 1595931502
transform 0 1 162 -1 0 272
box 0 -26 150 174
use contact_13  contact_13_0
timestamp 1595931502
transform 1 0 709 0 1 354
box -59 -43 109 125
use contact_12  contact_12_0
timestamp 1595931502
transform 1 0 44 0 1 164
box 0 0 66 66
use contact_7  contact_7_3
timestamp 1595931502
transform 1 0 705 0 1 362
box 0 0 58 66
use contact_7  contact_7_2
timestamp 1595931502
transform 1 0 207 0 1 362
box 0 0 58 66
use contact_7  contact_7_1
timestamp 1595931502
transform 1 0 207 0 1 214
box 0 0 58 66
use contact_7  contact_7_0
timestamp 1595931502
transform 1 0 705 0 1 214
box 0 0 58 66
use contact_18  contact_18_0
timestamp 1595931502
transform 1 0 211 0 1 354
box 0 0 50 82
<< labels >>
rlabel metal1 s 236 197 236 197 4 gnd
rlabel corelocali s 636 147 636 147 4 Z
rlabel metal1 s 734 197 734 197 4 vdd
rlabel corelocali s 77 197 77 197 4 A
<< properties >>
string FIXED_BBOX 0 0 1070 395
<< end >>
